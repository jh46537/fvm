��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���c��ct������H���{�c��ݨި��^ΊZ�9�:��k�m�4�@^Q���$F�o`�s�_��}ٚ5��г6j9����gc/��g�Rմ׾�rO+�D#k- ����zyrV��� QG�":Kߔ-Ym�C��L��Z��:[_c$�����Di�����$~�G�~*����)[��-cͯC���m·eȰsD�X���)	�u�X�wA�<�K6�=�F�@�M?�ף���LOc*��A���Iӹ�
�,D.�Cs.)2�X��ph��_gʭ,v�X�=�}5)���;z� ��n�����GT���5�����9�C�h��[����H�m�]9L1-[>�~b�q?I6P7✪Nc��Q��4���9S�s���?�G(ndu��%]�E\�A!P��	�c�>B���3nY�C�f��xY��\�v�5��K�.����B��4ӛ]��9�%���J�kǨ�SZ3y��E��%H��x/�����<�S��C��lh��3l�����_
���<tY` z�YR�_FX~���A�"H�?�9I���oN���1���*���$�2"�û��z� "�^�
�Ѱ=�s9��OjR腶.$e �}�,�he���{�.9ڗ�D""�	�D/Ѵ֔����Q��� ~8���r��[�U{������'� g1�S\h���|��J���8�.�(�۽�����z�� G��t� P����a�Ǹ	��7��\ѷս�.8�U�'8Q4�&W}�U��,
S��"��=��{?R��O3�� �j�d���d�J4M��ޕJ����xF��*���xK�c�ʥҐKG,Cp�����1u�.�.G��Xfq��n��fk42/�~wՄ�ڪ�?\�|t�Z���ބ%�ֆ띮˧0�	T���#���m��&�9�(�C2�� �\H�c�[�����:�<�� x=��I�V��H�s��2}�׀�Y1E��^�|���WT�`��2^�q�=UW��d2��*�
g�<;%;xF�;C֬{�F&��smg��Y�w�����(�Yt3��?��-��������s���Sfr�.
bR"Į�G@(_Y�z�2nv\ҳSh0^�Nby��C"��k����j�d���c�qd���I9:�L�����_��r��~�ZFh@��"0��b���둈����xeť�x�qw�Id�,cwkT,M+�w�֩{B�1�zj3�g#�A�oz��!+�1	4��2�*R�n/��(c�5��7g�<�W�h^�
^Jt�ͥ��������~����`� kvm+t�ޝ�K���@�;.�4��0�U�T��@�֪�*-�;؄4���-+�����{��o������
�.+��m:���9ɾM�Ć�}N�4��K�19�,��K4r�6��z�C��y��D�u�9<kIE����M�}r����_Z���D���J��F�M���Zo��&�9KA@�E�E���j��e;�R
/�Z �8lj�N�e�+�\�̏�VPK�%l�n�i�ɯ[vF�̆�z���X�(�Jzc3Z�?k1(0�!t�-b���v�>�!f]��cՉz�Wv���2�����0b��������ƫ����
ۖ�)�Zz�j
����hL'�:�N[�4�ы9d�����4z8@t��L���9V�a���<K������H�ϋ%p�\ޛ4UC�`m�CT�@���4;���0�egԃ �%1�8�K��a$�.@��+b���焐 �x���P�V������~�;h�R�����l���V&�������s�n��s��Zl�@�Ζ'�%�=B�M�ʬ���M��P"�vk1x���`��K�ג=��c�}����a[� H��J�-�c2d���ي�P���3>x+�wբ�d�q)q�
�$l+�;\�t�i�!j������A��(�wM4�bm֪֋8#cP�Ǣ�\܃^��+:t`�h�)�3Ԭc���$ƣק���	YPG����
�i�B�}⟍�F	�\�E�k��}���s#$5�E�}��N&��y%��m��yhϕ�XE���ϓs��$ɖ	��4G(�Z��I#(�J�?jU,���YAur�Q��)'����RoX�y&z���Q��
�s�e5_��K���2`��U;�՟8:��+�`�Jt����P�Q
��o^[j���w~5�X��F�����
��ȴ���3��� E:��\>�7!�N���,�s2zĪ�l�kɞ7���eH<L�@�=k�iR:>0�WO��K��5���;n+�i�
��kG"�{�c��R�Fک��C0B?:�����uU(D&�y�y_��gu�0ΐտ��z$pzY&. p����Qc���	jw��ʎ��0�K�?)�Գ��Z�+�;�eڮϾǂ�	�[��k:x3,�+8Hwfq"�~��d=�aIE�O�`�6�����KV�d"�rף7���5��e���ٕ�!��~��Ty�8M�u�<X����&�g 9�<u����ÿO�s=���-&��a
l���w��fa�;����[���q��>,��(<PS�ٯ��+� ���=��+�D ��E&��u��5���j�Ⱦ��ƺ���x�X�í�U��뱷��o�YL���'�J���!��Ǒ�tGZ�E��=�&_.�u'J�@e**�xd��#_d��k�j���zj���&�_"�_��P��aD��]!z���5-g*�^Ϝ�e�����u4D���zs(~�s��+����sl�P�x��0!3UV���1Q�X5�V%�N��@	Z���1͠6�d�.:n�#Y�v��Ӧ�y�"w����lH�y12�{��>�a2���@X�1��rYd =�e�� �1Q� xE?�FY4��J��3V�H^7SU<Ǹ�N��-��ɺ��˖�8���*�B�Jca�mG��;�U�
Q'j���]z@�uW37u����_cQ��o��-J�-=��Ӵ4�ڈh��e��w�6ǟ�t�P�>g�/��AA\
c_i@�1(�����~�`|Ԅ���j��u�8����?�MfA��o�Y��	b�ڢ�8doH\�x��i��(]g��C���Us�������|oJ ��]���XVEkؒ�V':����C��P����k7:K��b~��V(.��cĢFc]� �O��;�-�����v<��Sdr^^�'��J��B\��=��c�I3X]�ޅ��3��{l%a����j�J�"���#(dHW�vD��o0�$5��k����*���p������=|�a��APc�{����i.���B�ZuK��]maj���bLi��Ml��<�Pͥ:�G8`����h����yj����b��.�\��VS1��0jt�|G�#C���Ɗ��������+;㬷^�*O~X�]�3��c=��j�F��^W�;�o �3���J����0rm_6���+���D�Ů�k��)Ae)"|���@+�(@_5~�1䨌��<L�é٥��N�������4��s�%�u�9���vOo![�FH�I�ǴCqI��<�#!j��g�l��
E'�����L͐�[,?
�6�eɮO(^" �H��٥�J	���W?���&0����v���Y�k����=<��Y����Cj��K����b	E�N����1�c��<��8�N��]�O�r~x��ݖb�^�?��?�����������������j��Vt㋲6��S��k��$Z�g��5�>�߰ ���j�����A�{���P_�R�߆�	�.&�.7���͡�NM�+�ze��(g��8L$�������T�Iͫ���b��u���dT�?��=��z$��l�c��΂_��k�0p2�晚�tq�V�����vWȬ�D���Vq�?�/RMv��(��w&���U���';twC�EZ���I����X0?S<�\�<�����P�8�S�ES��y�M��z�K1*X�
)��c��`p��l��U�Y*�yr��s�F\���ݎ�P^:{�)wJ�m�(�	�����V�tk&
V�R%C�r��n4ٛ�-@+�4DR2PU=�-�z��ns2e)cB=��3g�5l��Y��a*�uy��Oi�X8��2��\������E���%�[���
H�#_$_�;�AF�9m��lW���jO{�Mҟ�qn�Kۙb�>#s�,�����0徵_��p�k�.=���q�ɹu^�)4T1 7Ę���W=V�R���Eu4�g��,�MJ�og�^!����A]��%���d4�9��1,(���pW�b|��$}�~\C� n�G��k�����D�����6�ѻ�Ś;���8Z���t��g�
5�D��&�H-6(*I�&/�����*]�پ�
�n�Y}{����;S	������A�%��Ë�XH��V��f��_�,����
��۹� �.��Iǘ="�*���tJ��+"410�X[r%���x2.�L��=�=ݩ2�K[/ѿ �ָ�h��]��85��)����j��gr3��o̰�
�~K���k�Ϫ/�_���pzz�A'HqUZܬ�A�M:���,&c��-�f	�����[�U^���>�Z[��~�9R��տ|�g�J-���SRkS#�]�$����Z��{��o��s����B��!8 ,����,�J���V5��N����o�+����$s���ޝ5y���/Kf�p��}�&���I�P.�*l�s �}�������se�b�Bag{��,��t�Z��kyCQ"׽�O�P0��!���|��j�1�7���̦�!�=�MS�����4�P6l��Ik� ��'��y��NǶ��zI��j�_=�e�k �ܠV� �oo�}���9�np�+�"P=�R� ����������'�@���Ѭ���^��f^0Iu\�o��d�3"Mk˜	Z�4�i�\c����r�c���8��o��,�J�]5����3��r�nG�����e��nQ(�;�2�B
�5�'+��>��g���m����#&?�ъ�|�	��k.\Ы��|��k(�5��e	)����M��65�E��q���?]ж�//����c�� �0�� ��t����7�|�/�Y���B����j	��REL,/'~�ρQ��'[���u ܶ��I�L� 
>O����`F�@����bk�&D �:��IR3�?�a��`��6l��Ɨӏ�\���	�jB�W�)SuJ�ʅz��K����F����Ҏ ���M`đ���J����2"�����ǔ�*l�,�zx❲���s(����z���'��4=Z}&��U�ս�RxX�����BRq��M�6&�蘕DD3כdIY_�����>���>!�s%��6Q*	u��v�g�(���}c��	 ���.Йn�/�8�����N��<��:��
��.��Q�-W�he�����7Ղ��V7?�t�|
�K�l���}��C��n�?o@�%�g��2�S�oIq�vpE
��}��"�nn�ѐ���[ds�o'3�
{�R��*�+�7���Zq6Ǩ���"�-Ŭ{�������hzK9Ğ��
�:��{f�� �Cd�#�{'�4_��m�������'~?����{>���I�q�6�����]�I��Cm�ܰ�;/��m;��Y�th�G9!�l�OE�zZP��8q��:��׮w"����_Qpc���:�1DX�N�s��� a����,�[�mf	�O?8���B!�1r�_d���l�>n?F��z\LmjF�xJ�x�8.1�?�z W�3�Yc�:���ќ�'C��+[���bT������CD9�z���%���(��"�rD�g�5f�Qx*{]k�\��;���n2�؎����"\��J�`�������9����� �̀���BR��rd6�(�S�~?~��R�?.}��z��PQ����c�~h�+5��G���˜�C<Fۯėq֧��%[k��lTO�狎h���1k�"�c����l���K����)���%����ʩ�V�)�Ъ�H��� l h�z$��� ́B�E��O�R���0:���(C�6Iv��k�'w;;d-���Z��@J�4ņY?��7��+ǔ4�d�"���P�ԓ\��$)g6�c4#<h;�Y8Y�Hi�(�af�yP1��9B������Mb\(��>I?A�E�f�~�`{6�[�W<�a=2}k�T�Q+[���?)-��a����i��x�ϸ�&ϓV��W��d��_��}j���S6M�3�I,$�n��z���k7��)9)k;m ���
��Ϣ�E�V{'+Ĳ�
-<�������2�WGiBR_K�Q̰J=X��5��6��Z#��>Z�ʲ����ef���:��ޏ�:���J�UL��xT&[��1Kl0A�*ä
��~P]|m�Gʄ1MZ�hA���zPS`z��%�����hMn��d%m�����'õ�|X�Ɩe���Sy�ħ_s���Rr��љ�հ��n��Bi��'"bb� �Ü��G�g�t��U��h�p�O���v�@���X���|[g[�*יL�M޴�\�Z
x\��Z�CW�$��xv���3fJ�����T�ɻ�>Q���2�R�6<�NNc��e���f�N��1j���O�F�{D�Z�2y�zK���#ǰ\SY�X��i�u��cc#��PAr��v�"�^.A��<�/e(��"3)�F6&��O*9}r��[[$�寿����F]3���.���R^�����b0���|��P� _�,�lĬ��V��� h��(IV��ڴ&�ޚ�<�'Gގ��_�uK-}�o�u�����6�
1hE1�W �a��ܢ�rp���uv�#�U(rG��WWm{i��V��-��;���H�#��]���ғٓj����Nz��u7��\>2��e���p f�H��\�k:;�G~��S��o��;l�|�������Yl�Nm}5���%�t�Ax����1���f�#�i(�2V�Y���D�iB�Lbķ��1��ޤ�0C�e�^� usf>��gE���(��ݥ9Z�M���9��V�X�)3�F@H�W�����������t�z!!(Eϒ?zÔ]��cPC��}�Q��*a�'�u�s.��Z	B���2��Ls�9��`+����O���	�q��Y��D�A;ju{�,���5"*Y�ÜJ�*M�Ԫ.y,4�fOU�L9L����$,HʪO3c���ؠB����i�14��A�3ý�A��ٮ�ļ71/�R�5[��$ e�{�1΀���'�wL�$�V��Xw����ٰ5�$l�6�T�𶡹CY(b�~y5b�o �}�5�㙍c����a�� i�"i*^�˶�y�Gs9w#�Wv�43>��G�c+ P���:\
>1g8�[)�aV�Y�O�7TG���`~�'P��,�8��HW����6��;�����΅��e��[՝R'y�d���^֮τ�
�ľ��c�ox�޻B<z�$H�ݾ�Y�H���7�����������$Ȋ�R��N�1u���������ZJ��Q<d��i��� w9aVX$�f����_���)C���3��Y91��r��O=�|��IB+z���!\�̈�Qv��+���2A�]4�|U��;���������4��������ߓ�m�W�Fǥ;�i%�񅑣45��bN�z��������� !��W�Bɮ"$�����}��z|�3����'��������`JNB�`�N���ٽe��Q���XXztDA2M��7�s����^����p �)l�-���y����bt�-�<@����Ow�4E�B�W�����t�(n���ɪ?!�\���Or��U�*m��Ӻ���J=\$���w��3�W_"򣄰�r��� ��݉��ޗ�W��MOх�����׹3Mv�L�,pzu).#���U��H ��P��%9�X�f/k�R%��Ś���Kz#{D��T��Q���!S�=��9W;ުO�>��A��եߕ�IC���,�xC7a�<􋍏l�u\���[\�1��I,	�N?�LQ�O)�ض((k:v5h�|bmu�	����G��� � ��C�"N��I��_�D��i�������Z���-k¾v�E
O��,"�ƚ;������M(γ��/�\R�r��ˢ�S�B)�����I=���c��� ʃ����OD�G 6T�����6��L<�n���� �u��ڄE�旋�]Ȥ�+U��~�a�6�������Y1�ѣ6�Pr��'���u	a��,�y��w;�	�.�'��#~��@�����0�
����3^f-j]��4���Yh�9����{�A��rB~�m�˶o"l� �,��(��d��a���-�˲nc۠p�X�.N�� ����/����K���={���K4]��'�,b^��bjnV�E��+�+BD0yh��^�^mftz'��x�������l-�ڹ�GS�v����F!:ʲ{�ă>�x��R�/�T6�Ƹ��?�/3ֱ�_$	����;,(Y!'��f�.6�{~|�>�IL?���¨��Q>><�����k�"D�gڳ������Z7�u�WP2�Π���0�^��{g��$�"�B�
�?hMF��pm���8Q6?���*Rk����	�2 ��E���@���c��c���C�={Q�����Ki��'����ݑb�'VI�J%͐ˆ���{�Ci�*�h�ư��U����-�)5j�1�^�y��,Q�G�G��c�;<�<ӡJ|��Ώa[،2K2 F[2�i{G��%�֦����Wr��Iڤ��HE�>��΢/ݣ�$�.4���5���2EI���	�k��x)��:y�1��2�寍���m>3�~�mֱ�N�]i�i�kBi�ߑfaC�SSyD	_{P�+YbL%T���W�)DbY��4c*G{���Hc!&�<��?r1�H7� ��EC����շ���m�s�����S�"�� �!_6�7��j̨^�a���ʹH䊗�� ^-���kT��+m"�E�ކ�8��EJ��w�j���%�B ����1	���eZ8�ۘ��a�)�b)9V_#$��}����07���s�_�@���GF���R���3
Lk=��*WEV����k3𗲙H�|ڂ|瞰:��y�����=8�u������Y.��ԸIp L`wC#�M�� h$7E��+E��"C�+(V8⤳���5:E��A�v�%1�"���+����|�e*���$����T��m�m����:B�6�p	�]����=+
g�?��m���f�=b������iE[�@�
�^�#�)#e-`yv�ǈ�ѮΒ>��=�7K|���_���P�R��-��)�!��E/���{���b"S{����׎�V<�rݝ�K��JA�QQ;�af6.���|��Q��L�����X������!������
�u��yKv���Ѱ��m-�m`�q��H�3���.��5oz1��J��u�ۛ�H�����X[v�I��V<)���H���Ohe�%��C� A��3=��6���d'�����wFAG�;�K3�2���S���/w�-=�H�}�&���c���C]L��3����w��8hsy�kJՒ\�,we-Y�����F�l��^���(4��7��_�_�wHV��ڡ���|x�'ߋ � ��t�ނ#�R���i��Q�x�d���
���ω/VN'	 � F{��x_?��h	�钺>4�-H�1ԭ	�ۡ��k6������g�x�w��4ފ��r�F��Q�܌UJ�iB
�|�g��_��c��܍8�uUa��X�v�B%��f�j�����&�l&�e���*���Z��i�^4��j��t�O8�	���Oe�0`D��8�5�����K��������Qd5���&�u�����Dh%K�(�ɻ����5���v�-c=&�"ZD��'n�Ts��z{ui}�A"����6��DKHmbf�d���U P�����jZ$���U����'�wd�E�z��<pP(F�%ۮ7��3��'� Bl���{�B�_#���)�9o7����Ub��rL\Nm�P�~"���0W~͎�Ǆ�y�1U;\3c��/�Nd_�=��҂_����Roz��#��1���7�9�C$�k����s�/���U\��A	P�r�����+�z�ٴV��}4�ݤj,��CFx��HGA%�inkM	~ތ�)������=��v�F�.��[�hn��1tߐ�0���5�ߏ�2��������q�}����C#����'c%zh�Z���q�7[�qA��O�u�|�������� ���-m�ݐ{��X�.��5w��0����0�&0L]��G�qm��T��kΪ�6��uxR�̯7�YJs�HWo�F���:!m��n��(�mɚ1�=}
��T�6�*WuUGF2E� �k�VWy�D�Ѽ7K5�ɿ�-��\9�a�,�),ϫ\�:Z4,H�v�B<erwi;�����v'"W��ý�P��=��j��rox�j������]bϢkV60�ź�sԮ�+��{Z�d]�dT�S�pbwv����l\m�DZ�㷗���.|j�MZLx�w��^E(N��3��*sej��|ձC���x��iO���׭D����n�%�ʈ�L���i\}�p������	5��`����[�\�V�[lX�0D�9�� ����n,�E��t>�j{:�����w�����_(���$c�I�PA�%�o�����})��6�3����M�y���>}��p���0Lh`��I�ɲ�]G$X3j�%a��WK}pM�5N���W+���N�D����֙\k�~k𹓦����5���������ԯ�X���P��ʂ�2��H����8-d��eu�S]�۱)�r����_6L��)SJ��2a���xm� /�[���Z���mQ�<A�n< �kN�`�� �-t�%�s�&~C��h[!E�NUh�xnӬ��fe^�kδ�u����Ŋx辌]N���f�J��f>�MWly5���-��m�V�~a�*LLy}����!���xEͰ z�|?%7�7Qb8�X��q2Ï���җ�uM��<M~KWC/�<G�=�'�S��E��pN>��|�[������oV����|�Ĕ�A�bhl�+�
w�f5vղ�5.RBrd�)���)�ۛ�4���g�ˋ�2��gDO�)H�?���7�}]���l
Q5^�Lb�k g�����%L�m0�؍=��
-����E��:�8��D]�����ֺX8y���` �E���)wQk��םkh��=�ٽ�����*}nf���$8�Ls_���# �9��a��U]���\�ɯ6��~�\� $ɂ�ZEK��c#��jy��(6=��L�'�
B7�m��Ct`rk���������K�W� ��hF�eO^-��hA�|�ۼe��g�:׏)h�'��,���s{�����?�lQ>u_߾��SR,��#[�y��>�,�t���W�;�oR�	�`���j̟���a)����e�"���i��'���$c �b�T�bH�X{0+��1C��n1���`�����ȿ�s9�#<�&|��CN����=�b���D�qm�g��f,��u��]�q6�b'�t�y߮]���ݥ���4=�g�~xgh���Ԋ%��r�g#v��[6.����2.�ߑM���*�"X���A�}u~ˌ6��v�N(�h�)��AĎ�^��J��<L͑�����	5����Olܹui`;@P���������ү�������8��4�+e��3&9�������sc�0�?3z+'��a����~>EK��S��؋�?C�p�q�� X�64��֚Y�&�H������3��Z��Io�	O�!\"�/�X�}�I�j��V�x������4y�=�	F4iR(��:�=���Xd����;���]ZQ����)O��[3�
B�}�d�`2먕[��ϢZj_[��bxQ�ϖ:����V�Ȩyw+H\s{VҬi��lķ�ZD��Cw@*2�I��� �����trG������mLxBe�����m�~Sc�3�\7�l�rHo5+��.n���Q���hn�.�E��P{#hXj� ��|�P���t7�if��bF�~�M'��U�����?>{0��>%��As�n��2�R�m��A~��C����ρts�Z��c�r�����ST���<�]�_m�@X�����Ċ�7Dt[� Y���7M�����e�z!�/�@M�@�2l�=���YM1�g�S�c�E�C�H�����*|?�����JV>8��:N��q2c��f�����.���C�	W3�o�/-P���� �́@�+����6�Sx�o��X7\c"	mf:����tÙ$�aΌ	 ��J����r��Q����=������#H��Vĩ����DTIo�� &gUܫ5�=pU��{\�_B9�,l0��-^y�ؕ��D�1]O���H�>Z}Wة����w�]�c/�T�@2Q^ ���o1���Tkh8Ei	j�6s����a��k)Lɾ�
a����i\������7�K�����/$������@M<5���[��RE��G^��U���@�2Q٤Kr4h!�IWl�p)(�|�	���*�<�!F�r��.&U睽�6>I�e0�:�]����9��hQ�Թ�m����c,�"o����g_�QK8:q1!���ǥ��S�� �x��wS�4��?�����)���@o�����Ȑ'P���w�n��=_)�rq�9>�Ugk4o�<�G���VCV)��J�e�#ݴbI���5}��q"��;����l襥՚�u"Ј�/ۃp�<��	�T����e	�lg���?xR^�����:Ҋ�.ПbCn�C���b��8�u�W�(0�7���'	���>�bC�<�W�P
zQ�����G,^IUǬ���������U��H�6j�?�=Gh	��O��we�R��Fǆ����;~EN黖{�l{1=1w|���%���ۘ(y2~��X�8�
#��2Bs��J<~�bG��Z�j��E��X��{�0C��E{O�j�ܒ��t��4.y�!��;Ij٘����~ZX+����I~���#j��vi@�����[��z-���ߘ�JC#U�%9zY4x�Xy�d����F>��`��F�m�������Y����!�����}N���� [�iߗ:���[�*+r��ob2����y�����������o"1Up���T5級������o����b�\�v�^�T�[Ok-��;��X1ڕ[�܌��
��;c	
�������X�1��Ե� �%�����!��Kg�Qh��Z�F��9
>���#�Y�����И��s��fF�`�+��hd+�gꪫu���k+s�����Db�f:+@�]^�(�,� 2ڧ�Ϭ�dS��aJ IG�mKs�xP<�E�=s0�����_�8��S$rRZ�]�{ѤP���s�׆���Oo��;3� ol�jϙ���� �9�U��a�?�Xv�@{�V��'�9:�rxï�_��}�	�x+"�f����C�1UI��j�~�0�S��	x��S�G��%���D�b�F�����ެ��A޶�D��썆�>�-V�Ć�X_�=���W�e/���!͏��
}㳷�O��Z�%a���k�3�Z�t��P��.�k}{�p���M����o�1c	S��@��n#�z����<�=�x���q���>����H�4L��[D��K����힩w��$����o��/�5��.,��[؛JX����Oi��f�w�H�6�ܣ��p�^����ѫI��=��fu#�
+""t�0 4=ƅ�`���*�̊$�vc�v�^�I��D��Οy�!q�Dzq�=t��C�Z,���E�Ǣ��.q-�����*��n�ߣr��<�t�I���q/.���+�ӿ�����/�D8��Ċ�0�~]�'��<ύ[��k�N�����/��XG�vdk��ɓn6�xƄ=��W�qm
�ZxB�p����m�ie5=szcB]�W�M��[���ɏ�Þ!EL(�9ؗ�����w(�s1�zC[su�6>&+��˧n	S�L��EU�x֥d߬0�0W^�E*���,@��t7��x����jS[�^.	2�+U|Rl����sCvib����d�Gl��4��#�n��;J��zw�Z�\5���|5�����J�q<��:iJ9R$��_7ږr��*sn�47���fn=�W���h��:�K>��R�X�y���1t�?�W��퀟k�����.(�F 63�#�\��K�И٫��(�V�?��X���ǴSɁ�$�A�lי*Vpĳst���(�I|�������4����;!
Nԯ�	 F9�0yd�9l�V)X���S���:�k󞨋2���8���'T�)ѣ��{�rfî������ӕ�Fqt�o%��sFO�����hb����-��)e���~�A)r��3'�Ba������ͺ.��UOa7�����cJ�{O��_���d����5?ա �h�	I���a^+n��;B�f�3�2��� ���XYd�%�c���vXO�P.	g�|�(�q��ς��>JRݝ�8��R���U e���ׇ�](��>�$��<=㽀tG�	����
��- �(R�?gS^LQ��Z�(��VA���������V��Np$$�R:�=�.k�?�y$���|%�_ �8G˖�4<#��K�����Ng��D:ua�-����9�o(�i�%=��_��r��k3o���ߞ(I����C�H0�q+";�G�5
.�D�T�ڥ0�V4�'��5 <�8�ݙnsl�9���lf����dD��(9��r�����=�+��E��
�cl�G��&�m���� }��iR��[�9baO�������M���l[՟Բ�7ݢ 5W���� V
��/����XY�0#���I��i�p� ��ӹ�Ҡ�wa���%O�jh��_0��F�x�^�.�ϋ�=2��������p0�Y!�хd��J=����Đ0
�u+�� �V���;��+�o~b��~�˪G�u�_Ey8,��l	�"Q��f��xq�4��*�S�	�.�ғ6�� ��1B��V|;Y�=A�V���/�:2�HD׏<�b�K��E%v�M����]��vAcw���G+��bJ�l��,	1�UO�S~Z@.�b%�]Ov?�Ě��}���v���-�O��]1�Y���ô p� ����A�u��9_��hb���J��ТӀ�C{N�=��	 �h'}M�w8�EY0#֌�佐]+�����:.䈀��W4�x4�
�~���}=0��4b��=o"0���Z)¯�at��L	n"Q''�6S�cSJ-�ΆK|_�Es@�n'IQS�wLz�{�У.�S�N�l�p�"p���g����pm�u�B��m�C,�%y�jۈ@�b�l��hvY�:�]�KP^�ѿ��*�$�k?����
��`�g^�S'z¥	rB��;��p��"}�J3ț�cg7�nV�;�1i"�-�����s�>J^`mw��2ft��,���9!	4�:
lm���L2P����QA�bZ��o��f4A�W��B��0��7����!���z i��po{̢�����]�/8��@WH�x�r�,��}"ѣY5� ��8�5�e4J��sǸ@�](�3_4[b,�y&ׇ,<�*���4Ý����żt�I��M�
�����/9��^J�9�7������7�Ȗ OT��n�T�5�vK@�Šz�#�X��P��q��N<���;��l:�Q�6�g �QO6U�5�=|��g�̨ծ5.{��:f-��ƈмw〘z�乹!Gr-�r��.mv,ٯ9�!9n�[ȗ
��VM��'�3����EAR���ܔ�$ +U�^ĞقL�X�b#G���x��@��G A,�΂F�unݱ}�^�^Խ"̦����<T���oW�ȴ9����I�d�ŏIW[	�e�ȏ���w^+�5NV�IΤ��	��Q������oFU�Mt��N�a�X��2����q#bS:,�����|Ə���GD$x����7���}8�!�,�4�W�6��E$��(�:�{��V�����+�$���NG�����Gdz���� ��0W(Q4�.����ޒ�<*@��<J�>�����R�Ȁ�&}*��	�,'�b!�\��y��|�ً�=���1�(��_aw�p�Tbo���]�3�꿎��UTRq��B��R|J-�ͼ3��/*�8BeoR�*1�J�>�sg6�>����H�/̑��Í�;����v\�t_�t�r�E��|w����v@��^�|����VQ��"��/�ߊxpPl	V9xтf)PL��$�ؙpx=6���F"cJvw�_�ռ�uNOg��hyW������uc]�⢵2q��B���㑧��]yU�q�6�ї��lJG;y�+�(��Z�V-��Ky� �`�n����k���&a%$�Q�h�V��YC,����#���,��E��_)�E����E��*k5SK}�_l��]�{�����` ��rEcY�]�p�k�3���㬡lH�R'׮ L�O����i|�~��%��*�{7.2��}�Y�,s�_��5(ζR�9#�yF9M�`n)�":J����G���B�D����x��>��Q�2�~���ᯠ�>#�u��z�Em�a��S��]? ����-�v��<˹�g��ݽʟ��<��/f�t�sTn��[�Da���x�+�w��7���f��Ĳo�g��Z�.���D��<'n!���M�h��9�_� �� 9�_�[	�"���A�����w�7�W�r�Ǎ���zz��KW���eWz�]V�p���k�5��*,�+iWN���u�N��p�g}�;�ǚU�?,@��'!h��o��d^?|��VD��_����2%��RK'[�-S�ˏQdj��3���\��[�-DLj��p-xF���0�i�J@��e�KzW`-ז������i���r!�j]|P�b'�&qY�Xޜ}��#P"�`b���Y<K�'��	�AS�CI�L�J�!@���j"x��O�A��C��{4l�����}[C��I�1�m��Ȩش�UBk�r��b�y���-�`���}�/xE,�������aP�6}崨�����ϝD�9P��o�$١������֔OCA��<:M��>O��I<ĩ�#��>�?�S�*�Uْ���-~�X��!�&�ݎ[V@���
�7o���b��J�w�{�h�Rk1���@�K�w�7
�HoƤWĤ��Pr˻ ݶ?tZ�}��l�Y@�Z�ivra��T|�(Ox�uI�M�Ƚ�ǥt����iI������}yP��i�ZU��{6X�PH�^���J/)�P#p����l@�8,�O;��{�O`Y�ߗ�����n����D�����άk	�cYX�J��ډ!�c��Hkו	�-��� ��{��D�0��W�D/r��ƶz��iN (m�W���Ĩܮ1����9 �c�qX��7�.
h��<'a�z���+���`�r�vN�{?����7{�>��A�V�����[ f�S��b�m�E-�ٝ{k0�N>����K_"q�Q%:�烬���P?���v�E;.�P{BX�!L�Y�%H�������]�	8}cT4A�_�C(g���*YmOq1
�g�{ƫ�����?Qm|1	T�D'��z",(MA!!"4�y4��o֧�.�1��?#����B	*A#@�yV��KzC�!H���x�H��P%�(���X�=/)�4"�+�ڱF|�1'�A����KM�ף�IJ%�*�(��w��T��?�>�I���_�������Q�	�C�@Az�_�O��#:�^�T�V����ט����M�C�������;9�-�-�^�T�%U:�!�M��яw��KM*-����/\�((��`��Q]�ӕJM' h�ml�\`�� K,\�Wd�[ ��~E�E��Q���G�Z���N�D����@2��m"꘩�^�ԍ=0�d�u�5y�C�
u�j^�:lG;Y�VKJ�"��l�.����<�0�PXC�؄��Vv��%R�
η597ޫ��$0��i��n7yJ�2�׉�*�&��t��#R����X�^F' ��_p�%Ä���!L`_<P����C�B����p�`-�Ӂqک[�ǆ��v/6��?���Q�3e�SaӠ1O�P@�p��Lt,2iɜi$n�K�>�*�
���GO[��rWd'V��}�f�Q�As��
)
�����|�u����@����|k�W�/W�6g/MQ�]�p��R)²���xI�b��@<TK��\���13o	b�j\�q��Xv�b����lt���1Y|�	*�d�5{��x+))�T3�	K9���Yg�
�~4�;i7%�7 )M��@�`��~���E(k:;��
��o.����d�ħ�7:�4^-��c���n�;��츥0���O��D�tp4��M�B|���ED��W��o���e��T���)Ϗ��K�n���v���rl�q���j��d�A$�)gDZ�浪{�#~�x�+�R�.��E$����֩�d�{Uk&�u�����۲v.��h!�E���r���A��S����%�.Pl3P>�8���j��W�7aׯ��Iz�P�v��t� ��Y@>��9�!Zf/^6�ᩛ���|��w�Y��������X)g2?�k���Y,��s��h�k��SN+��ȍG2�%�\�e�	�P��.�14s+q7-��Jy�O��}_o|��-Ć�0˘}s1�����4��~��W�V�J�o��O坡�v�:G)Ʒ�%)��г(�!eO|���gj��P���f�s�e��>������i�!5�k)�	���DΧ����Ť�#�w�Xa2��*��6JG�9�~��T��s �t�	49K'^��`(��+�۔~4M��%��76�!DL�:Vԁ��N�u��F��� ^�Y���;�?g|���D���ݧ���႕TM& 3����	&w�b�!%�z){�JF��z���g�-�'`��a� FO�f%t1����g'ɳ�S�+\� ��U��'�)�hn!b�"�Z�����9�fB-�`a��]�V��E���1}�?�s�w�A���u3��sS�C��z�^vFM�aDu�3q��I�$F��|��X!.�Z��r��l��Ƨ���L5��;;t����IȎj]���A~b��}�qkTG�>����~R�"�~񅼥w"v J��J�v^[�͋C��dh`�{��>��h5T\46���0f���4��S�<s��w���PJ;��d*k܍k7�d�I������'��=���>���`q���:-Ce��sB�%b�'H���n:�6��IB{��_0_�R�[�I�a���� �z��N���wR�oC�"5���vLmE`����W�wwQ9+�(�/>��8a�������假Sk�I<<��W�F_�9CI.���{_ښ(�����+FKk[�_:,ޝ���yb&�ߪ�r��ܸq3_ˬS�T4\�4cu�7����m��V�s�9eM�B���?�m����w�\(�H�� #`ƂB2U�ͱk��	^�=��(����}�b�RB/�i^�RoU���<|m1x�թ [���X�p3��_|�&��!z��yP��^]�P? ����W~��!Og�c�LOu��<���A�#Q�	&"a��ޕZX'�<���n���"���[&0ԋ	�Ct� �`���TS3�^~w�kc!U���<?�.�lգ �`�b��YEe �7��d�I6D�S(U�7�,�4�ܛ����+	4'F�b����j�R�N&Uɟ��EY�:�<J P.�%�����j�Ϲ���	�l=�TK�GЧ���u'��U��̷����̏s<�;�Q�$�jey��y���i���b(Mi6�·f�ኝ#.�S�
��ۘ'�o,��+��rB�7��KV�~�=zKP�����g��&CPZ��$q�$�Z��qI
-� .�ydQ�0W=�.+�IEyY�մ�y�3"(U���\�
���U;�I��ߥ���뤡i��ֽ]e$�k/��4�,���9��p��#��+�RZ����z�|�|zհ|�]DY�uJ�*L=���&��\��#�}�Ϟ#t�+�ȬB����������2���m[��7lŋ�}CO�p�A������h����p� �ӟ",�3_�'�1�c�~���:��٬-b���;&�=�+�kG��Yn!���N��Nm�;:B^���Z6���� ���{$�� ��	�D��}He#�vu^7{���o�x����X9�2���LB��g�Y�����+΂�׳���R�i��%�HC(����<���4��l�8�j�� ��6g�d�Pb'PGB����W�
��ve�����;�Tq��V�g�*k��9��8��w�{þ��,O�e�ݯ�߂��o2Qe����H!cG�@��x�_M=��9{���!�����؄��PK�/����3�(��@6��?It���d05П
�K$����fO�N��O�ɔH�@�7�0�l��)���z�O]���G#.��l�7K ��)�� �#	���NUפn�X4l�3�xg5��l�sԐ9Ҫ��uFC'�vdupqYh��z��e��J�M$�=�	�7�*0�-*CIDn� �!@��M��_kƊ��V96KD�Sk���f�V �EDz>�X��G����̓p+�c��ON��5`�%d4�%������o4���]!���26[;���7s3�>����z��&�]줓4�����f���A���{�a�Qڳy`��:��MU�xa�=�_���d�AXD��������fǣ�XϬ��~�v_��Z4 p�	��c:}��߅��"ca�oU�2�����_j��f0ْ`v$ou3�ᴳ�}~���m�	��N��'����w��`�j7A.�q.��=1I�w������SE��yhKh6�Y�yl�؀�#F�����X��>�y"���<&U!�k�$�
P⌀&�%���k M��ST�A�^�b�r�nf�K`���yT���
�|L>%sB��*���HEhU�?/�z�M���T�E�p�3�+ͥc�/1�m�ྦྷ^C��K����_Z�=K5�ѱ����tO��e�w�
���X�v4%|<�(6�v�Xr�8�������}n�9��{��Z^�!�[��Q_\wD���P7nQz��7y�e���?�z|r�����_��3��7.`!p>w�h1��W��qb�q_�t4���T& "�����n�R�8DP�j҇!�Z��bM��� 4Q6�'S�b~�k"���x���I�,/���"�u��$�]ķR��l6>~L���I�5���������ӹ�P[�s�.��o*!@�S��JV��u���+��
G�����،lU����M�4���g��2��𑑽��_�%�42yq+����f ����7|^9�tm��>�~��:"���2=�g��3��-)X���t6�i����`j�g��b���lbԢ$�a�-_k�OY�_��v���,���[CU�~x&�xoi�"�.*m��-���`tj
�>�fP�S)�z���£/㐙L����Ǵ�U��GWk��I-�y�/�O5?����DkAy����y6Ӥ ǎ��0T���˼�
~����A0�}x�D�X��c�ʀ���"U.=��(�爅��6��
E������a�`36�7���_Bi��[��<�n���o����a8��O� 7��j���W�����u@$�|4�|�bfw�����_>����q@}��LWN��.1����n-���{y�\�F�5h���n�ŕ�hp��d+\�㤵t��_b	�W�Ҳ�|ÍmSh�`����+���?㾀��e�T��N�w��ܱW�WaWB`_rQHL������j���R���V-_��>�F�uڎ�$p�w�qh�K�-�T�l��.[u|����<z�7Md����eH8�3���.[�\d��s��T>@,B�Wy�۟7X��"�t�E��Km�@t�5�����V�/o ���z�*#���6���a�#���#�D������u��"�s�i��� "�$z9��>�C�v�q�o��'P#�
N��n��hͣ�z	���{gp�Au���=�4�j����Gwg�h��ϟ��\���q�՜��ǋ�}��-���X����Z\N7�x����5(j���n�8�0KF�s\@$�����jK��y�|^��G��Lp	����d`���M���R}�K�H�biC!����Û_r�P���ᖷH��0	��6��t�+���>Q��,������$����a�|q���� �(�a`��ᤠ}Q^�\�[�#�,V��+�5����V;	�v�gu�߷s��f8���Wȍ��,���)�2L�j�<���3[;\(��8УmӗbDy@Z�ަ�\%��ulR@S��Y� B
Ѻ����٪�J�_	�T�,�OJ�&�J/��0\�艀���+�^A��l��4��|��K���>���.�/_�A�3`���K� �E����n�����X�;��O-�4J#nk�+�d�BF��A��2����$c��b��p�9�_p�� ����h+�>��J(ʱ*���;�G��V�.4)d%ad�r�*m�HD�c+<(nR��U<(٧�Τ���ǒ�~ӟH�hD��VK��\��]�llp��f���`�x��EQV����U��Iep�S��u&���T�$j&�ׄ�vz*=|�qH̥�gM܅�9qz�D�u�t��K���6W����|J��_�������$�EB�d|I�#�;S2i��e6���JQѺH��
��:�:�ܯ+�uc�'9��W��$Sg�9!!dU�}I�������wv����n�b��!��! {)��,F]���BI�=��f@�ӊQ`��E���n=�� ����>�u�����r�s�ug ע���45��~�H/v+8CH?�,�a��gI>�0��I�H���	�PGνE<����-,U���l�#��{��Gɏ�ʇ���4�c��#��	��ʥ�e>y���i� ���Tn�f�B�2�̊���yj*^��x("#vՍR��L�=��z�߰�F ���^3�7U=��G�`}c@4\�$����@@fns����m#��S�4��7h8��?��C)���ϐ�x:��f�ޖ��횇33���jW_��:��l����H��Z��e۠�l���$��p!0,76�if��1�K�_~�G��)�:��z2#:�ڎp'��7F	V6�!C�� X g(�x�M,ߊ��>���Y)5����/A���ma ƠTԮ4�����*U���D�_+?�Ʒ� �\@%�3h�u��R<���7x�(��d&ڮ�YNTS��r�,S��-m���,V�Av��d=@���.Z���v��1 ���S͍��g9}��8+���|g��Q�f'����+-�6Xr�Q��C�\���V��d���e���
	,J����gM����2�<�i�G����Y�.�d~�c:	�L�o�xR A����d'L~�����x�Ƿ��^���h�W̍�Ex��-1����Pwyk�Ԋ��Bڂ�gQG�O�>,.�`e�Kp#��������} �6;�/�����\�S����]^�\M��a�1ڭ;+y�����,G�/�,t�zow�N�V4��Vw���D�IO�#��#�S�裪7����M/Pn*�i�/!v�A��Sd_{(]1����K�=I��;�7[&��J�L�en����x
��[����>�LWw�:��tUЧ�v�v?X%s�D�E��"�v�J?x(�gι(����r��r;^Ms(�J	�(���+mx`	r��,f i��:��u �O�\�q��iT|��*�0�B_����/B+����X!: �NW=�~$�ӱ=�T���%N�����g�z�^1��}�N³W���!�Z�s�8Y,n�f��ۡdJ�J�3���4vB�Pޏ�{�4!�ޣ2�?ժ��7xc���x¸�(�W�e}(-��m��'��#
"�D��]���Ʀ/��8ߪ\�\|��w` �J�1�%X?�q���<�P
�&�P�_��5�}�	�&Z�5���tq��s!:�x����P�f ��q�����;Z��ʽ��$e�%����%@�a����G� ���� dkQ��?g@Y8���a#�y�zLDV��#便�&���bլ\<�h�ˊg9B�����3x+�/	�+nQ*h�^-�q��yS�W2!���a����o,�Q��¥K��i�	�	�'X{�?��A6騿���8�f�g��t��t�T̳/�k	N�(1đ� Ƽ�UGΗ�,уn)�bb����8�#�����)vxK����4��}�vl�.�7�78�48rS��!%���C�r|��R��;6�a�1�ʡ��z4o�l����2�����&~?ϣ��P������\q��,%�'Z�\y$�a�}Y������ћ\��$2XC��K�@�\ ��a9H���z˔�9H!"����]��b��ɽP��"O(r7�D_gh"�{F�ƻ�Q���G:���U������X�3w�b�w_�FE���p��A�]6�|s��89��7�۷B	h�1Hz:A������N.J�i��4p%��p�PT�b������!��B��������UW����
��Q�^�F�n�˕�^�H�*c�ؾ�����UL��6ZCy�D��\k�^�[kZ����>��gB-F��2�Ǡ���K1���ES��Q�L)�����(�㑛�=���-W�-gD��7�{�� ���I	~��J�yd�O2D�i|]�'S��x�	/�$~��`�}8�4��\�?���H;�|�\�|R%��SQ��Ckq�ġ=ȱ�1�?5��!,���ԓ,.��-����V9�,T���&y�<�j��Qwg[E�P�cZPW{���8���D�*fsm����� �Z�v�hm+AqN�<������X3';>;WHO����;���H�7z���Mm#�4����<�Ϸ���Q�7��=�g�.��H�T9���6����5��<�,��鄡��-
pn�G�����\����(�ܰj�X�&n�r-�D�?̽�j>��M���R,�M��WY�
�Yd�>� p��<ms{�GDF����j�����(5����\>��P��ު<94�g98Ȯ�[��}ǳ|�S84Ŷ�|�r���r���ěQ��cW��< ,8��NG,G�E��']�+>�"��E�zלt<��JM��r�bfG����z?%+ǅ�W�W��l�pX#�F8J��//(݉�������}s��Aّ����q����Yj	�r�t������W�+��C�s�ش�Rݵ~27����C]�2_u��E�S�`Y��I�Ɂz����
E�w4��C�l�heM;+,H'�	��%��/��aʤ#������;*�A�����|��� �u5�J7�	�B�v����|�
6d�v�D嚞�Ofa	��u��Q�4��m����+�PT��O��q���R^C�SBC��!��3x�! }���:e�¥f^�seh�ҋ/����ѡϕ5n\�WpV�%��X�����_6'��
�37��g`F-����'`�.(���W���P����q��{z����n�X�����}�Z�;:�x`E�=������P�b�Y�^�?r��`վ���>(�������x�;c�:�@�Ve�4���U�gey{��$Gz̩�h��!y>�z8���{]�14s�t��B,�܉vX����+��<5`w�'!k�\�p��|�xW�V8F�:�s+6{��|�
���ub�G'����JDh7 �����YU�nF�����5��[�1����t�B��D�ڌ�כzǯ��7P�X��k�ma�3?�n�,�z�߾�v.)�:4RG����7/|aa)h��%��玭�^��g9x�?����N��O���dK~@��r�n	���%Qh��bC�H�3���[	5�W�����K��5nB�^t�L�%Qz� �[}�
բ���^�l�ޙ`�#�9־L�b�}2Z��nl���m�L��Hk��'c �-7�ކO�{x:��qm��s�tEa͛���b��IP���Ŧ�͗c�>Kh�=�֕�Ob�[c&.s*�@�isژW�I���bF=f&Ol���q
�>����2����o��DҮ�s��M~���k�5w��c4�FCE1#���V������Ї���_�+�M�a4�Չ�q��ɽK�NO)�'�	�D,�¶sc�=�F$++�'#���f�_=��\�j׽��X�5���Y&L�!�T�/�J���`vi���)����0��t�\v�XE��[�$24�AnC$�\�b#Sއ��ѪXV}�r�39���6	�3pvw�-F��(�*xV�(�QcĐ�O"��=�05���Ĩ�(\�mu�E7l��w��)�5X@4�v�,���鍌��%�x)�����0��)��"�o�T`*Bm��X�X�[�ڤQ�:+��H/ܯ�Z�	s�C"�������,P���*�dZ��F���2yĩ"�,���7oȔ��KmAl#B�D�?�g���~?p,I�����a���i̎B&�:�f�:H��׵��,q��E5ܒ��4%́&�v��2������2���-,2� ��# 8��4�}�$�{D,��.�A�r����=�5*cA}0�;�YN���<{X�_���Q|�J)r1D!�%�x{�"���S�u�~���a!�l�][�(AO��4��}>ܰ�YD��b �y!�oO8�6�<�*Jn��M�Q�O��Ĥ�:T��;��%	ϼ灮1��@Rd��.���5q�O=۾B����U8�_0�˳2��'����Zx�'7%o?���53������L��	��|�۹�
QU��f2������y��)�h����D�Pi�X�~�72���&m��A%��wT荁�|�ZqQ��ټS����7��z�_Co	�b��`��j>wܜeW�c�]�J,c�N�?R�^э���.�+���w�?3��ZGd8��xV�<\�!^'X�V��s���;����#���tZP&�����WRߊ<Y>x"pc8Ds۸n�����֒�2"Y,�b����H#uz놽ً	�����H�5�}�Rd�i��24S@b*��j/P(西	�fe=W#�7�I�c�T�M���{B� �2��_�<�� |s�Cx�q�vlR�ھm����W������������1u�"��@�	�T��:;���@Dj�0�"9z+�u��������Z��D��'�̦��D���a{"V�JvZ�3��2�i؁--�VX��Lr�p�$��=��'J�<�OՌ���el�\�S��E��W�8� 43os�3v1x����V[�����A*����-8E��9��Z�`Ъ��ԙ���|K�7��u9?�ꚑ�,� D��E�ǂkȠz���~@�w�Ff��ePKK�v�)f�`��9���� v���^MۙC|Z�R��usn�O��mVE�fs���+��KP�︴x���2�_�-	��(-m឵_��R#������G�ڢꄋ�����f���;M���R��Q�%\@�S�2՘�Q��7
R�>{���I�rN_ޢ�b~ƾۂ�/pqy��!~� ����F��Ob������:�ނ��"�!!p=�T�|�=
IA���.�,�n06M�]��1a�}�[�Q?Q 6&f]��������!�	D,F��~�,ͣ�`9��������D��[����27���2�j��O��)�[<n.ٴ3�iV~�ې+�q��t�wr�v�.��w�³�/�_mp8��-�J��Uf�Ԝ���e@ў�bE"��Ѝ�4bQ���lϹ����Ò>�y.�l�22▭��~����m���� �x���ȱ՛�j4�A�[P�U�OuG��$H���[�������J�����甊��E���M0�x9�Bأ�0����*䁤�[\�p��Ug����*�����Ka\2���E�<�.{r�y�'�NqY�J�ң��4Dcu��$��S
7U��� �����@�8���L=��?L�SV��L���~���~�%��/:w=��������i<�0�`�>��>Ҍ����케��_���NCڰ�K���/Y�}���S$���e�T ���,9yx������{RD���8 4W�3N�+ٌ|K)reVN��+�GF	5�Ȥs��O:cc]�!����O[1,���=��e$z�D*!�5��ߢg�A��7�$.w�zh�5߶��{d4١6�|���y�s7�u5�g������/Fp��F��"�LD�ʥ�)dniq�1/uU��IK뾓��D�\俓6�-�2�-wĐ]����?�%5o����7͝�����eT��)E��`of�E&�=)���ְtw���}g?P�� 5Ma��%҂⁰7�����3�u���)�0�l+Vv��B�tC4N�� ��I����g���ZG�v�'�O�1ڡs�+�l,�蘮lF����e��yB ��W�K�&+	��Щ��aŨ�#��q�\b�&c� vG����"�H�'�l�y5n+x���Q�nB yXI��d����"�֍����b&_�m�>u�U	0����c!N9񬒄��� P�$A�����l9��N�'0@,9t��9�b:��Jm�����L�G����c+-.=oI��1}��(�Ц��Gr/hO�R��?�cWa�5��>���`�R�sd؄M>�|;sWl[Uʢ3�!�k�Eʑߢ�����I�[��a!�9�re
�*9/VmV�u�x�NsJ���]���y|_w��d9����v�c'x�x��6�h��7+P`���W���(�N��d��f,�V�|��s��|t���Q6����7�E�պtwA>�<����gT��^�F�Z@�/2ٙN
5:/��a4�-�im&{@�9��&�u�#V���Q�̰�p����W�v����rK�5�*+���,���0,��C��.Y��,Ƒ�b�jJb�5u��哪������s��b�ޡ�NiBĹ���ۈ��c��(p���-F�3#������#왾�-�!�A��n�I���x#� �,��a0�DO���b���`W4u[���}w����[~��@�<_㽵ߓ�������c�o�q�� _�0i���/���6݁�]~�Y�r���ؘ�y�C�P���H3���`���3�m��{��.��,���X�)ߒ|IP�P[Oݔ�P���ga��&emy�TU8KM�1aJ�Мa�}?�脩��_[&�徴�]*x:���*͔����,Fbb��0��V)L���[/xS�C����so�0�A[yeƜM��/s�R?�C���1<��9VTkx�05�� ��r��|���n�(!��4▏�%�&�?U�3b�Q,��*t�`�~Y��IVF�7�]��Pr�T�B<�w~���a�QE��u�8�����s�����8ڲ�x�mWx:JA3���X,���8����PlA�`Z<�|p�Ph���D�,d��f�#�T�j	V�m]'��T����ai�����~O`}4i�O�\o��>�G�>�#�+�5�f}"�/�Z�ys��mg>��7��H2x��G�w�����W�c�Ǻd:��sG�U����gV6�=*N�ĕ��j�w�v��]�F�\��S���H�� ��뱵���[7�C�S�_� g�����H�څDZ�*ѹ5k�)��0o,*����.ۥ�Y�bE	{;W�t�V>^y���� ���	N�If��4��f��M=T���|%s��I��6����������!�ߜHh�u������տ�H�g����{b���A��َ(^y���btt�~�sZ��n%V_�*6OXs���-��Ӳ���o�Vb�ZY'u!;E���67�'����\k��1[���㥦�G���J�x��� ��O���AWd���<'_�l1�J'�|�@��(��M׿�	ϻ/�g������4p�_}���
��I������}2�cx�TՉ�XFa��\�/�tp>������rr�1���^�D�#��y��u
L���������@'t=�Q�4+kh���FTk��΁�q�^{	�l�7Lls���X̾Ѡ����=0�T��L8} 8�� h/a��K��Z����Q:��289�<�Y���K�э�h�4Rmcyc�6��hg���|�}�����x:4d��p��l��gE��v��r�|��k��0~A47f#3OO�q��0��F�d��7!�d��ū("���c<&�I8�M#���f��(yq��5n��ﭝ�mT+?W���+s��^
LS�rrs��+��� �5U'aj1��8��D��'��C�K�"�ZՒ���d�S�D�i���{t�I"O�^ҽ���0��"�7�R,9��p�^�r�b�%s�}�B k�|�V]��m�\���JZQQӃH E�D�~�af>��d�?h��:��m2�{Y���A�����v�YX gP�-z�@g�ϬV�HM���x�	��p�������O�P;����!д����)H�"��l!ҋKH��/a& [_Uz�g5��p]�7P�7���{k8�vo윦�~@���0�2\�y�`jn�6�ߐ�Bv���ք��6��H�FB3�lt�T�3)7Y�9U�03
�UJ�H$�N�����/^�{�'M\��!o����m�%X\Akх�]������6?���]Ff�Af��t������NO �s��9���&6��0��4��4��j���o)��@<�+ �U㧀�xQ*iU����YBM��~О�`���G��ڞa�dFI���>���9�b^Q���$|���oڤЙ����&�o���C��P�	��*={K��M�w�@1��B;�\�3=43z[� X��*�����2+=�~��QR�:*��P����{����)4`�IֶJ>��I��Z��[󯆉D�	=�,]�P�v~�v���?��g'/��
ޑ,��^������+p�Yi��i�B�ɨ���u�Q�O�כ}y�MB�q[�#k
o���+L�e$���XZB��7և�`���@�5�f}k���B��9Z��������� ̝I�"7Px0h��ho[�m)\Q{N�р�d&?h��B^��J�4���̩�q_s��IykCk��o|��b�x��m�x ��ik�c�A�WD:o�:j�o�䕥�	��[�=5�,`�K'����7#�bz[��I��xI!�"��m�2 ��'t�v���kpoqr�w�s��R��[�w�����
�R.)�c^� �pWA�Uc��D�I'z�o�d�}p�O�J[��d��\ȥ-�HDW� ~e�	-v+�P�?�,�G�	�L�Q���������JG�Q��jK����Q��>M��ױ��*>�V�@�d�/%F��
��C4�E������D#%��=�����r�:�.9��T�B�O�_�ENOX����Y���q�{�<+���1�e\j�������O�K_Q|���y5C��m�6Y>I�{�Mk��x*G��$qG�^DZՂ�}��d���)��7L�����b'�5̴MIѹ�jQb�ee1�1��e�2�i;�qG0�IL��b5�~�M)@�0�j
��.�1�g(믜��r�tq�9�w����E�ҨT\Z�	]󵱐���#vX���~H�p��kb\��TN��L%}�Ͻ�MF�~i���]�oi��TQr.�of���e�P>Ԧ+�W[Ms'������.������)j��fd�y>.�(8-��p�F�c5h�ű���R	Iz�q�������ƣ~b$gh,��0fS�/pXyQM����ȋ�H>PJP�X7i����#P���ieP	�eٱ�@��~*9�b�
�PR��5�t���E�3ڟ��/�uL�9�~W����+���㘮$���_��]W���?+��zi�g�!\޳9�ۃ�b��T~���=��m�zs�58ލQ�'a+,�<�g౿��
��	�T��Ï��-ȶ��R��h�ى�tN^��p3�+
���u��xH�:�B(��+�I4�iH�keLU_�"G��2��Jy�*ס�!xŭ�_�y��4
�~���ˆ>1&�n�E�j�ܙy���a��)!���4:��3�E���,CTN&L�����^�~�d�e'£�;q!�#�&�u�Ч�0ȿLsW�<���MwO���묮WW�G@O���M���M?J����.�V\��\�D��jO?J�6m��.l�8M׊��ɖ�3��,�с��
��Be��rdO~�Eb�S�*�F����R��MpSV�����>���m�k��L~v�'�V�V��}�hM]f-��XvϞdJ�]0��σ��͎X�Đ ��eb��)��4�˲��V>�,أ��4�\Q۾���r_���LK���&.ur��@[GD��&	��5Ĉ��nrhJ��9��
U�U%V��}+��nh�4�}@��������
:~�V�O�C�Wy�*�J液�C��(���~5�l�n�Kr�*�3�7����~F�T���ye��O��+�ŗ���ƛ���,���3ȟ�\�Jy�����q�G�$u�Nc@Y����ñP���g�'��oQ�xaa�?6���@tѡH"~��R!h�g��yiN�# ���q(���<q�GvIS8��Q��曛|�uo�kKC~Z����x�<�z�Uy�%�	w���/c�.��b�u�Bq�����~0R���ԯ�J����`*����p�z����� +��:��E-�Otjp>������Z�?�Si`Ϟ�d���cV���
5㲽P��������ȡv��ppC�Q"L8�]3~����O*d>���W]���u
�	�[8��h�`���Z6a��e۬K.�w�?d+�J�����U,�=�"�w�13�!�(DA�>ԟ�Y���r�R��������|���z	�F]'r�׊��r9�!�7��E�D'�
��%��[���*d��� ���4%[hR�ϣQ`ި�a[���$.��K�R�+E��
'�>y~��4�Eo��[�h�8�CMEAL��A�j��م�������y��B�_��	�j?jU�<�Jd٘��yaC��	������9��u�2�ĩޙ!;�o��9e4�E����EJ�9-��:V�;UZ!bխ��~"7O8�}~L�hx�����\�U��*a����5�@��[�\�bN�D��7uַqM"�q�IKfmx͒��W���1;4)\�'�4���ċ���c��,] ��h8�fO�L��֍�m�Vf_$s�����
�i�Nb�O#.���Hns�?fI�H�Ȗ#��tއD���;�o�$O��2ٗ�}R\�P��W������gg���_>��p�����S�[v�zdT��O�fP�Z�:�3t{����jиH��+��Dn�����"R��Y?Z��W/���F�-�{�2��B�p��(R��c���%���M1�޺�έu�[��k��ۀ��_����>`-q(���Ԧј����c����pZ��[n�ܯߺ��*�x���!�dMET��,:�MEP҃zp�!$q��h�[;�Fl4�϶,��H=�����/��M��Z���`��%y��s�_ڃ TC�R�1gA
vKg>��6!��\[^�p
��t���F��yv�D�_P���Q�$@�6G�.S�2%Pٖ������a�S�G��0��=�f�N�Km�E�]���B��M��e�˜2�n��v�B?�<nk������ʾD�
xq���X�oEm����S��d������I�i27�>{�`e�a����h3e)b���|�<��W���.��6��[��qL��Ql���B���a�	[f�h�C���	��T��T��{���?
���?a��y���֡�nIE�̡ݸvO��8�|���2K����"A�)��X�4w�b�=�d�T xɫ�4�;؈״��ʹ�5Ǎ��ҿr��.@��
�p*z��������䚡�h7T+h��#�l5WT���v�@40_�t��:�+ ڮ֩�V�!l	.�^��A C�l|����M��>��`�9r������l׳({lp��<e�,�g�g�?�[��|F�s��	@��T*�W��L���Z������RŠ1�ʇ�ְ�I����a˲����[�>�}�R�dE��������]�v�Ƅѷ��`/�D�1��ʪ�&�-O��C4��;��,Ysi�~&�L�R�%)����y�9}]z1F�O� `1�����P�q��S�p�OtA7�2�J;���O�|�1ף�=�=STBjG����s|�bЌ"ꤴv����q�{
���D��H��|�G�	�N}3��p6߯BXH)R �
�I',�m�(������}躿3.`G�.3�$��h-�f6*E/N�(Q0�">��{ZI&��v��o��3�H]����7 nO��q�03 � �u��eI��Ȗ)�7�2���d�-�a�� �Lz�M8�V���[CL��>v�Me}��'�Ľ��In��Χ\/:�f���>dq�VO1���=.ø�)��u���I��>x:h�.�W���)��/�N��%�q��]R�e�k����{(�ce�?_��(���$���l���&�
|S
�<@4�^��p�J��l�_�y��Ij���N��e!'����<�3Y����JAD�V�5M��-�~ �+��C�Ѣ\�����l�X��4ӗ=o/E󌫎���x��X����l���������o��l��V�U���5�?����| ������W�w/�$����+M#���y n��d�8w�~L3ikg+��i�U�b��������rO��#�y�����%��Y�j1�K�o���ճߠ�S-���Z8��:P*>Y�D�/r��j?JD����H$s��$(C��\|���P&�|��{(�O����	��@��rk�2�"x�҇�60�P�*LԕU�H��Os� $�9��#�)�q�j�'�3_43������cy��oA�Z���g�OgN糕z� ���v]d�)#�/)vm�A$�wkcء���Oh�3°�N,m`9A~�?�MK���?N�d����T��l�e^�x�ܧ�����5��S;|��QC��Y5v����8�Z�aVu�=��U;��H��7��:GsyHDu��]|ŀl���-���T�>FB���ڀ��RD빽7��6���i��~g��Z�Mm*���.�]�:`_�zy���M�
ܶ��U�4I�)	?�/�5� ?Z���.]�2	�+r���L�)'[��F�e*���kYXb:��'n�D`��Ԋ�^x�?kBHX�q��N\r+���)>�֏����ӑJM��N���C!`"��Q�L�O+L��;M{�s����@�̼\��`$�|����ۻ7^��-�[@3�d
�5�;�մ7�����9�Q�"%�)�������х��*�E4�g��~3�gx#<vm�GB#��j�k��p�F�\Q,����XA�o��n|�5_,h��r�e��W��)f�<v��=���	2����Ux@�ҿ�� |�T��ٌ)�T�g�>�|{�76C���~Ʉ���S�|�Ob	?P�3H[�a��bQt<8�В��cYC�V��5B��L������1W,(X`��gthH���w�)F P��O���Ch��,���d]���1�A�m�����$=a�	u��X��T�:͒�/)E=T��%��J�@���)�E�@U���J��'co�1���Ӡ�mxp��� 5�_��+�ŤO���0��`O͉*H=�Xv�VB �5vF�+F'�m4�X}�(��
I�L��{�x��Y�fX����K�#]�P��簊p:�qb^3�ř
]�O�jf��)����>u���o�<�pt3��ŗ��*my�V��rU�V�a2��Q�D��+}��} UE�$����M^�b�۟/͑5���Lۻ�	�is�\���5шa�Zs	F��p�Ӛ<���^�s����S5r����,��ޖ�/��!��UY��������Z�3�tw"f��l�Ӡ���$`������ʙ���
(h���0��9	!���{7�W�C���\]�Ҝ�������V��*!�3;��1s��y�%�Д%�mXEwq̴�or�PQ3D��Ȱ�^P�t��L&l՝�z�1r$퀛M����QP�J�~I�&,i�IN)*���B%o�{/�N9��I�[����7H�9�ưgК���1�_�h
���U
��6;�ݵ��Wl���b�����G��P��ز����:ض������4��1�r��:~�|-E�q V̻����̽O$���N�с԰˪�ڕ��=չ;[���v�}�젺��w�D]Z����1X_\�3� -%#�:������J��jF��ː'��}��m�Zc��	B@֡�|����x�����.���F�յ$8�[x�������`<�d�jD�{�l�+14�=�&n��q�>m=���:Wn�p�8k!�b{&�o��0�{t˰��f��*�׀ү��J_���'���Ά��u��4n��,�vJ֙����1|:���\�a5��O��g,�:���=��	��а˛�g��-��찝;����D:�*��e�~z�à�N�� 3��]a��H��JَS�nJ ��8�W3 f{��֭uւD�&N��`g�%�j������(�_�IE���8�SȾ�g�@
�V�復�C�d��i�TD>2�������/��9</	+�SV��CޗB�g�Ժ4Ì��ED7rlM���Zѿ��Ȯ*��1r�1!rhTOS#;�Tf`���Ȗ�KR�c���1�� �� ���_'D�m��RAc�����KM���իg�>������B���#e��=3j�_�"��S�k#�Ĺ1r�N�I4��؀��]�$����;�f�d�[qt��� �<��6��J�X�N+�$�]r�EFǅ�u7/+!�o~���-�����ʸ��'�nMhX����b���I����*lB`l�
�w]��	�k�ðGF��]��4DQtH�{��ʜ�Xb�k�̧T�(�aC&hl��l����4��o���~}�,ca�p���TIgV�/@��������ve4a<��ᥦ:9/����YH�?��J�t3 I.��et�6֚3t�F+"����"`��CJ\� <3����׎̲���.�)��^�6���1*O�	9��r���[Y&����!�g�勈h~���ueb��wQ4�o��� �c׼��;��2�F���+��!�&~�m�g�k�}��
�����lZFX+n!1�j��玼᝖%hGi��qA��@{]b��8l#��	�]_�Z}�����|7ȹN�ʏlJ	T�p8�w���,I�f7�.��Muo������V�7�^d����� .x�Z�8�\'�����W���}]]����y��\�\������Y�j"x @�u����~����\��4x�����*+I�P-�:og?�#�v��=:
2D���u������"���\z�w���?��\��NLn��m�|$0�j���n��.i���Ӫ����Y:5�2�?2�`��5�m�w��q[TA�t�"qY���S��͘�ǍF�^���?���RPJ;!�Iwʤ`V���8w kw6f��1j���s9��pŨ��f�ͤ��
"�aF�3�M�W���J��
S:Gr U��fy���^l��D��:��&�95�)������F˕۟�C�C���_^�͊��Z�����_���g^������B��Mb��O5L%��[ʞ��&Ĵ�$����`QJ��3� �۬���U�,/I�r�N(�mrm����3��k*�O��\��m��G�*x��ut��z�4r
C�⦽���`�=�����^��e�4����U����wف�I��\��'m�F��G���	E��ǏǸH���m@�4�٩�/+o+[�nkLAv��!?F�x~i a�!�z!'�OxYjӚ ��$�����G�)J
�~�@�T���"�|ж����5�u��^�:wE���8�;�_�/�Ρ&�2)H�k�)Κ�~=!��o �xm���J&�D�ZVi�y,{�v��	�S���Qj���,��H��̊>�0Ϝ������t��F�����u�y�x��h���6O{��aA�YKd�T/|���eHؽ�.�W��C���)�ͣ�e��I�ri�@X�^@F��? �:��k�(���eX�6�Є��$<���h~mvv�Y�	��_��{X���_4�eO��[y�䖀%���Z O����+��C�����̆�svU��D�U���@��W���?�@�N�|�p<���|���N����L~�g�������u�a��-�'T�N!���i���m�j\�'�N�+�7��!<p�[f�������Ѐ`m����W�*��/���G�3z�_����Dj.��a�Z�P���W����v�g��~�w+^X�I��'��Y����V2-$s?�`?b,��e�/���|���X��%/g7���
tu+�y���d"��~m��,\��$?-/o��,<aς��R��Tؔ�⴮��"�7[��T��4BP̧�В����dE�Q�Q�?o�-�B[]q�"n����I�b(baBD�z��_DCE��鞽Gンs�.�=�Ej�U�
=fY�Q|Ž�1�v�
�QZ����9B��-8�1����= &ͲC¬��Z=�B/��OUh0tD��Y���ε�c#���*���e��|3W�4�{��q���������#���6͗���e���J���(�C�OD=ǫ����<n��H�7*/d�FqFF*$�K� �N�\{/�74���S��b:5K����{�7����<���Ol2=u���}�g�S�_ȐN��{ĂB�y~-��-�$G,$�R�L=f
�?Ȫ�ً5�-R���"<) v�1�P�8͟�'`���)���NV^}Bl�_�@M�Ǣ�d�g\�G�����d=_9�.�a����	�h�������X���l/�X���x ��Q-�*0ó���_gY-®ln~��)���x�1����_���C��&mT#�r=I�
p:;���+�ŲK�o˝��d���KΕQ.:�k!��NU�}5��H�c��*J-m&�P��wD!|*Ț�c��c}ީ�}�Y6���<+q���������qň���R����B�U�i����nf�\pC�c�?�� .�䗿��"D��p�K��gEi�1��Z�0�ȍ�~4��(p:d>��W(��[k���g�	;9��W7Pξ�@\��Ԡ������5ZN(�����C;v�<;�2�@�RE�K9��'�3�!2�=�P�˼�6(��9ϵN�&盙,�u���w�"���{3�vac�{�.�+���
F�c0���p��S�hl̠=[�2W2+޻b�[a��?��,�w�Wt��Ro6:[�u�7�3����Q�,�:Re 2kŹ�ogZ����9CH��@Sm���M�(Y�K@���  z+iv�`�{e�Cgc���{���?�_��B���^�b�C�-_��"u���T��A1�S��H"CA�3ѧ�~^h4�b��(x}��6���!j�Uk��/��l|�Ԍ�i��q�5T��
7�HW�쐴\���Și�N~C���C�>�f�.���=�q=�=q���~�UPRl-�����'���^��8��?���@�ސ?��ű�D�����M��r�j��;ݪ�zE���������g�2���W[�LΨ`�Sń�Ěƫ�'���fIYB�d�7C3=;�$�X���}6��sx��}��<�/���{T�b���9������N��oa3���UwŴN��,7�,��~B�7l�5�1ǟ?K���Dt�r��8����Xg�T
�j����e)��x��e��RJ�>�Md+�ڷ��u�])�A}����a$�6����W4Vk�_�)݉�I���a�ut�F�&��{�X4��A<�\�42y�Xu�@��-�T?�nF���� _���Г��c�a���NA���*�ʃ��e��늼soS��*/��|��~/��U�w�dKs�;�ߵ�C$�~TS���[��@2��rxEH��ŷ5X��v?���FrRg@��y�m��25�2��fc��L�4g�bT9��Q����=�~�Lf"��>�N���qrGq��F��j�	���2��Ŝ�_-Р�Ż�(�5��T�,c�e�)(;�WQe^Ѐto��ז���B����(���L��W�3���)U�7W(�ܮZ�Iu$w�AGL\Q��;���r8蝵�����׵W|X�n�U��˅��� ��\��m+�h�ف��m���:w�o�ϵ?(/��刅�yG08�!�woXm8����b�i<t�E�:o"�A�{!�,�o��]�����;Q�m6)��{�՚F�<6�������I�$�� 3�"g�)��<�W��Ed.�cZM��2Y7��?5�`HJ�ٌW:�FةA)9���S��t��Iw���"9��5�i���~� w�n�'�Q��$���05��(��d�:�9p�)���fZ��T����~@H87�?�Q0�b�B��ր2cW�[�P�	)+�q��mntФem���s)0B
��"��^%���b�>2�?&/�>$l�40�i�%c�U�}�mٛ�S����R+xO��_J����RL����JA�<����p�ߖ���+��nd�e���4p�%�=�����Z��xpҧT ��<z���jm��!NF�s=g�����u
��K.]��o���O;���yqR��0G.Ef�0V�9sØ�VD�x�n�F�#9�lğ���'�1}���w�;�*̊Gm�5�eL�F�_'��I?�UQ
�[�'�����I���zJ�@�
�<>���$�����10
@)'�W~��
4�zd'�-d���N�����1���A�i��c��nk�.��� �\���|&��O�/䓎j��p��ڍƎ�Mw��|�Bw�7_.{<��)1ܣ�q/�܇�ؽ�L�|7���|K�>W��k$,�_ǯ������A���� UB^k�C"H�hh�g�ԞHʽs�ͰK}T�%�]�7��j��~����PeDL���:��j����+�̟0�} ��%��g���{��X Pq���N�fí'�o&�}�ݥ�u^$!*0�����Uіޜ���i@���l!��>(��^6P2��� �튌*���� ]$�hl�=��y���t8C9�%����(��<�\��֥�ZW�&[��<��ӎ /v�%_ ���M7e��$����y� ن����A�ݦ�v��IAO<n�?�/��|�I6����,��{i��Z��E�\���l�+��WNC�x�F�.
B\awִ�)����?q��dk�*����P���u`�>R���֜%xLb�Evñ韔;��������T-��\���.���AV���/�~F��ƥ(�xB����O�E���w�|-�O�����}��N�#�6��Qt=��p��Qm	���dJrݙW��^����}�Y*;����k�M�S,zN I���t�H�@V����?ĉ�@2���9��k���]s��_�k�ll쪫��{�ڟ>�<�ؠI�Hb㒔AV����z�}u��{1g����_��s�z4�^�W����f�S1�L�|�j,����H�s̤�e[�
8 en�ج8πl3��G
�/[9��Es��Y��԰;c��g"�b�R���AE�-��Q���u����J�SyJw���p��7Ղ������1�����ʰ�O�M>�����
�3�\���[�4����HN������\ih�j�c�r��#*����L��	?'(�#	ggg�����p��d	��y�.dL��Yjy2�q�2@�f	�'�s������\+Ĩ�R��	�#N9L�GC�yZ�C���n��W}�A���g���p���X\���7Z����N�!���G*JS�O��_�eĘ��#�,�^%:���,xna��c6�0�,����V�&EJ[Ȟ���%�r��K��g_�J��'�A]�]�1�-�a��G��̸�۵�&�|H4�a	�:����i7
t�z3I84���!P`�HP�P��G�> ��o�������0��C뼇��d�%겄�}t�P�����d�~�]�>��M���9˜\D�y9����m �-l�3 
�+_�&AB�2t�n2�tw��n`"i�y�K�������ɽ�V> X�5p���I��}��^��_y���JN܉��\x"-Lh�x�ZYOXح���PI�>c�ن~��{%���H��(v��|�3:�����iۄk�.��Q ��u1pP�y�G5�ϒ��?b����O���K�!��&T1��Cwqt٨,�(r�Z1�����\�Q��(�"��O��g>֞w�c	b�<��o��;��*-k*^���z�SQ'�J�ϫ~X©ke <94��5�[�F3��s#�ݟ���-1󖙈|h%�R��P�@�	M@�; ���Ս��i x�.˫�B_�t�nb_�%
}l�<>)P�u5s��ǀ�}3b��ω'#P�W=����}�)��o
��~Ȇ��_���m����o��xy�
�c4vE;x�'&ə���=͢�E��kޥ<�i2�!k��9���λB�����T&�O��oS�Α��mf����g(� ����a��	��ĩ�� ���x7n�R�����W���L�Ӻ˴W©��C�l����Eo�{~���YH�kj�rUݺ��fy*Bz9L<��^qgr�������o{��	�ru��T�#W��1�p9�_Z V�ۭ>��X�Q6�8��m:�8v����E�51kf�a����B� 9�w|������e�:4�����.�1{��ÿ}7{��1�S�P�ǃO�w�a(S�s�������d�D��Ĭ���z�ū�%�y��Xt
�(�	!*�?'��%Y�.�=���E��<iI��f���*�p��˾+^�6��fY��t �SE��V� ��zb�-z� �*ݜcB�;y�3���w�=D��Ne�0����ew�WE} .U6:�|��J� �����h�1B�m�B�aJ"�{��)zxo@��9,Gx���p��R�^�!�j)�1�^7�/ԃ�+I�ms���m�!�r��$�a�����b�1�,r�n�N�Ҕ�:��Ē݊�f�܅d�����AH�0Q��:�U�����g�v�,`�E�C]�;Z�:�&K��e~z7~<��s}~-�-�*
��m�.G��$�ܡY��W&x]�A���Ny,.�];�ۚȽY(x)m>�@M߇�'�z"O�"i���n/'��D>5>ȄP�#�I�B�{:�¼
A����R{:�")U%�/�[&-jY*�><<��'(/�;���w��L�<�o��#���l54.������<
c?���C����_��C=v��IU�5�Z Ͼ����T�׹�?7E^%^"%L��y����+�2mI���I��rOA���b��ȸw� �_���kM��H�{��-�&�-BK �!���9:��2�%�׀ͭWe1�}��0�A=>�q�z����OB��A�6`�~	��X=cM��j���;1��F�K�A�g�ԌX�^ً/hk�A�)���'>��3�e.@ǡ�H��T�	`����*��\�9k��R�ٷ𣃾'ñyh&�J&���;��k���	}�����:��Vο2�L)�:�0X��Q���/��kP����պ�Pw�c5 C�`"Dq�+ 4��>��X��j�O�-f����%���O'L`����G�����/�g����z:�%����=���}�s����`X���b�R=�SB��8�em�:�d'��ϰ>�d.���+��c)�B5jq��݌���}�PL!}��0ў����j<[Ɵ�����P1�Db,�q�ī��/�I�@+`��LJ@H�v�K!#����<}�����z4�8���2!�YQ�!I�,W�qiF]����ΏX�,3�ą��Pֵ8�d������/}�� �In�c�Ձ=g�_�O���f��xl�=����Ub7��Ì�hx�|�pz���y�V��ma��V��A���)�*��iP��x���l?J��߇��x�h\�J��7҉��3�	���B� ˈ{1UաmwGC	%�A�w���5 ��aS�,ۖgp�1M����أ�n�,Z L���ӐJ�;�D̶��@l8�i�m1.��� ������_�rT�ɩ��>��+� �
���
�x%<_�^1����8Ǡ�w�͞�49m>�@�}za��x�+!R�~�3�|�W%�pp�y�������AAY�9&?˙F*����s/��Ɓ�����H�r�{����h 9&LƑW0؉��Pߒ��:T"�қ�Ъ�G�֌NlC}��vnu��������`����+j�p�E[��N|��^\���㉄e���W��h��- �e�;�wkvh"��s�岋��YC�cWl! ���!��)(�#D���4rV�4J�lV]��炌��9HөeD����p6��?�TD�o���ִ�9/�����|@~&������d$z`R���؁������%�5��:Hz&BU:�EBv<��T[�m��2$T,#[y<�_��0f��z�_%�Cޡ�}��C��:�y�<�|��PXmU�w�@1B���Y	�9-�Šm"�j8����ɉ�V0�Bw�Ǐ �L���1�@z*��+�_1��X��)�/&T�m����`i�z��d1�W���1�P������Im	$%�]�A��m������,Z6;�¶�\ۘ��P뿣�]���$4[�D������l&�����&��RYUhUЬ�y�3Ăf���vǋ�@<� 1�_߱
I�ćU�1��׊%<�ǖ��P�4�F���}|y�3`�_��+��R�%D�F!������>/�U0�l&�r9��a�R<y�����ˡC��o�_vXO��אָd+��B��4gd�w��i������1�s_��~�f��q�[���r����Gk*1�>����t��L�A���Z�:6��q*A4JR�	�8f��^ė�����>I�l�R��HRvָ
�����4ԦH��9}�JO4-��X%���>EXD9?��]��@ x�n����<y�ܼ_}l[�&���[�
��ù85���w�٬�b�Y��;+��%�p�po�"�I�� �
�"����2>'�<Z\H"A���D�׶�����1;��2�����.N�B��:I�㉇(k)aJbw�1qK�V/�H儺��]�!�a�*Ա�(uA���݆��I=�M��X�;�zmϛ|�Itc�;5&�����r��DE,��&΂m6CSk��!3��~����N$dqk��'���R�]S����̝�X��"w����i���96�srn� �j&6I4�b�#Hp#���>�8��͸�2Ox��8%��o�ܖ�a���ԏ�d[ �[�t���絗�
��LҼ��&�ߏ��˕#��sǞFG��\�F�#�G=�-1`@�:�Y�k{6������~3��|?�4N�n�6
�� ȎQ,m�e�P��ga���v D�wd����m\ �Y ��V��[ҵrxNG��e}�\���s�G��Y&;^~9�hH۱��U�O��̝�_�(8m��e��T�
�yIi��F�c7:�p2R_
�s�ӭD�w�1ʤ�r���f�`�P�T�WD�kt�r@�q��h��T�T�~-"�fB�Z�-�5�{���\Q�.����KA	��$�$X�e3{��Z����z\g�ݞd|C ��?��L��Qݜ���|kn��ǻ����I#���I��g�+�� �e��O�V���L2:���ÅvMလ�=�L��s�~�0O!�r �P�z-z^�aȔ
�[�0���1s*Ia�;�3�?�"Gt?q'c�;�����-��ݰ�-ݵ�����/Jϋ��xk�?��0w��������DRb'��fOp��&�p �������6-h�ls�S����S���ᐣؽ;pb�k��"[\*/�]xAq��d����
k��Fh̋_a���.���+M�����=�觠��c�s��_�/��{�����`�I8�߭�e�C����nr)���C�{j6s9x["R�%^�����i��>P��,{@����B���j���ǎC������zS�O7�Tq4�u,{0��l����va���&��~F~د�C�2۱�'~ۻw�**h����-����ꊓ1`�.�ʡ0q�H��Cf�df�X�.�����;�I��Q�/�Iel0Dؓ���g���8 ��S���n4!��1�h@�0d%�/���Q��˳�JF�� ��t �#�ml�D�,F#bh����B�O2�=�c�������ɴ&����ʃ��5K�XA�c���$rLڦ�>�R���GH'�O@p��TH�iG5ཪv�Kv���%U㒳0t�2%�A��X�0 KxՇY�t"��,|�T�4�E�Ræ��q�k�\���a^�(~��8}�oxzv�՘mD�������|d�C�!h��k�Xu�X�� �B��욘<�QA��3` ��ġ���-�D���lS��.n�
�����l.jtǐ[��YU=q�	���1�XD�r�O��2{�6S��g[-�Z�O��:2$n��uJ�
+���kې�$Oe�Oh~�he���*Q{�-�߃��ڪ��h�Z�9����$�Z�΁RZE�7aoN/7�@���b� (��N�O�4���N���ңnJ|� ��Y�{HL�b�#�+��E��|&�Ν���&y�K�YB��T�:�X�" ��^
!��w��)F8�Hz(�DK��ZQ2y�ekv���-ŏ�r�H1k?v�@8{f�1T���r3�^�9Wغ���'�p;�1%?<�K��]�����a�U[�n�ol/�)��_��t�,Fm������v��!\2j�h�I����Vpɝ�d��Z������vk��W����F�#['��@	n]�vB{��@f��ݰ�F�	p�(dc�Ҏ���KD���aF�}��B1�e���o�����n��L'�:���N$sɿ�>���_G�Ψ%��E?�����f����F�6�6P6����D��ʨS���1b�i�����N�gr�N��s>��	v��sM�8f[�����٪יtV��������v#q�*���X�(�3��fs��*u�2c_�)�O�������b[���<��dD������N+S#��+�ŝ)b;ۑں���f�oJ>�ka��wh��9��|/? rc��Y�C�hQ�SB*��s��%`Qc 2�CO(@u� #��='yU���|��}�v4ԋ\�LS��n�M�:��}���ןŧ��1���̰h8����Z�^�=ۄ���nm�k	uǾ��4��ޗA'��*ۓ$�;�MQJ��*>���m'p���b��--��H}��	D����=��j7{Acm�O{���ܬ�����M���j\�B2V�Y����GR��+��[��.*�g��_��*�c�F�)k�%���"q&�4�#�t�iR�E�qxSD$��t�Ү�ݍ�+�WLqh ��upr��حШ'v��(�6Dڂ�ت'�ۓ��` �sU�����w#/"b�PE@�(1��@�����n�j)�x'�=����jP{���͊�*�-S+6o��al;kCظ�e�k�mF�#0�Ɔ~��ÃMx�<K2���n��ɭ�L^��o�r���g������"]���]}�I��Pu]t����H����u�6'�k�j_!�r�f�����|������6�+�i���C�ˑz�.�[�*�'�Y hA|� �Pߍ8�m��ڀa%˳�ԍ5U��r{.�2��Q�����,J!7��fr:�6���z�i]���zx�˚�c_̝Υ|I��1���{��nz|�"���zm�J��K��բ��f�I7��a���1
s�f�^�-q�;yc%$�99��"�<׽��҅Ω����n��� �ǂ�4��ȜR2�y �>���x�ڳ�i���w��QR�{(��z��5<�-J��m&_��%���c'��K���͖^0�4Sq�ʅL��c� W;U ��?g�x�����k������Pܿp��2+c������k�6]��i�Aͮ̏�=���Or��z�<i��y��a�(+\Y�b ��*ZfG\"c��I�Ǯ"Z*�4Fg|?�J0�i�_D/��̺��Ñ�|�οXZ�bG1�c�ύ<tu�����ߋ�d�Pt;�I5�s�7ߧ��Sy�G��&���v��TȢg�e�.o��{BT1;�(O����x��>��n����4 g��B�e%��0/vh�O��gH(�?/=���W��*.�bo�����D�fZ'�Kş�zO���lA���lJ֍�3Ս��r�F��C)���޲{���[/w��F�,'�k�yP��1&F6=�#Y�n_��$�f���Q_���g�ϵt�L��z2��;ǲ?��5�L!����H�J�]Pޖt�HO�J�[�K�2�ɗ�)�;ʳ�y�#gU"����P+(_���E� �A*��'�8�o�K������ټ��M��x¥qV��lw��E	"Jc���b��>��s�2�w�ׯHƹ�	��ptb|���p�U�gT� +�3����UPk�]��x1F+`�S�)�:j��	�a����Ԉ�9�� �е��*�=�	�]&$��:c���F���C��t�>���"G7�HS*u��9]�ݠ���[��uV����ik��GF#�^�b@��y�3���m���A
_��y̐N	��|�E^���q�b
OX��0:����N�*��Q���B;��w�wB��h)�F��PX�,��*0��u>}�R�r��˓-���!����1�x=庉���A�O��&,#<�}A��e��Qq.��	")�1
�M���4&?L�$�ox�ߵ��X*�x���ȕ/�U��1p�@�ch��A_�-N���jy�{��U�(�3q�fdW�bt��c��qw��C�&
�eU��I?C�K�(�
�ƋJ�v��;tv�ɖ(���W��a̹��p'8-�����b�O�鲑��_���8:6h�;]��!Q��0ru`�|쌗η�`�z��h�n�UE���-T:j��5�o�zv��T��qN��\���R����9�q��V^�j�ae�U�'=�@==y�G؏��D%@oo�U��QB�Pg[��h�����mc��oк��2�zB�7c��%�ڀ`��dd��GX�5��<��)_��g%	�jjZe˄*��<F���J^E
�O���QBYJ���U4����������6W8H�ux���ݎ�;����.�+/���<oZ�<��5/7�� D:ص��$�n�uJ����V�Ѵ�Xȑ�y>���S��>���	�b+W?�Vb�>��.�����W1�PT{s'�>ͷ����5Y���5��|Q:M@t��tŻ���Ҧ7���(��(�õ���Yk��B�eW�rf�*_��k�LS�pe�~zZ}�,Q�w{1��K�\)�L� �v�v��-�ӰR9�d�@��ݽ#�|�Dr�уE�2�WeR�3RC������H�Z;�g��T��`��S��ȕ��Ġ�7���;B��rɓHqA����UI�0wlo���V<���x������,,obB*�";į|<^u��f�p����1� χ�ĐQ�ɐ��b�w!�Ca��i���횉�O�s���F���,s�?<0���4˥ě���vx�� k��6��3����|�݋J����aHFr.:��di�}�@ O�wj��P\�x���/p$l(l�`��9�{&���<Vy��A�J���=S���sI���EVM�o���ҚmGz*>}����{x~	�%�l�E3a� Uv�?h�q���W@)����}���Q��<QM6�4����E���B��e�;6O_qPv&��k����d&��w��(�k%2�CJ��%�D���`�D�Kvᢦja4˄��*�a�D���𲳐;���t���d�t$��}�.��QZ���V��A�а��~��� r�xo5��E��S�BZyz/�7���������,=����º1�l9��|(�x0�T�H.%�j�u�ѩ��XBLLY�W%���V��H��c&,7e�f/���Q�*���}�aG�
�p�/E�R�n�eK�#�vL�����I�>Q��&�wb&��O���.С����-rTF���I���`{��~��ޠ�H�(�@���ŨK�^ttѲ��No��6`�^���G_����N���|r��|je�z|9�Y��$�����G�pj������v��
@��Y��L|jP�r��he�1����z�q�[`�)���6T�7���?�����4���v���!��+o�7���Ͳ�ԩ��{��О�����w��Y�9�m��EM� ���<��@������$�X�d�y�-��fY�$��@�<��1T�ˏ�ؾ�z>��W�XZ�Ȉ���P)&Jy�/���{+����X���cŃY,O�c�k�J	��˖��E8�����aM�&p�
v?8l<�^��NX�e�����˻����o,%1�S�`��Rnp�*W�dd�KӯqN��/���@Q��W��-ێ)�+���
"N�,��
v=�������� �G����.F�.���RL�i3 'E)��;�ev@�<&�2�Ϡ3����"��h# ����ji��(�H�lJ������B�,�x���+-=fy��}�]Pĕh�
���o�m
���`'(^�c��Q�/�ȩ�����x�L��!OͭN:v�h�q2d\w�n�V��w�g�<�����묝�(��hRh�-��L훲%�:��kQL�2~��V��*���y�&�RF�7����c[�&�D�`:1�s��F���4������5�s����.+��~'A~a4��3F�a��T1Mf�X{��2,%�_p-���D�x��	J7(	U���.Wkc�f��+|�B�J���zk�<,2�)�.Y��̿X��s\��x��j�P�����R9�K���/&�-��G� �F�m}f<qTJȊdm����J��i:�Y~aY��BY�lS�u� ��o�1�����q��<S2]�t����V�HӐ�T�t��btl�jUO����[w�����A���ѽN����\�;�:�>���6��t�rs/۸�t��s���c��	�Т"�Q����{*Qz5�3=���>f�
e�9�}������G���O���6v����Y#c��Y���@�[�+?��p"O#�ܝ� ��� `]�|��������S@Ms]kܜ����!�DuEcI�'ù��E�hS*���)�xa^�I�!��V�M����[��2�����_2�޷ϛl��8Ӷ�V	�Ò� 7~�=����2N��­7��i��b�@u�L�r#Ο�����,U٨�)�;b��$��-��H2}͙�1O
�� �vH��)�I^y$WcEA�p4���.���9���U���7�U��ڊFBC�d�_��ӈn������`NGI�\��������0���x1b���q�����Q��A�(G����L�5*:픟�<������,�V����F�Ùm�8��)���#��M �7�8���"���/�z?��6�7�%k�8��k�1(�/��e�/�.Z���~��r�ٲ�<@�s�M4Q N<�� L0o��Ex�U�.!�W�7��-�X��6�p� �h����?3|M���Ŧge��B��6Rj*���/j�U���b��w+Ef�9�5<���<��L���� �qH�f<���S\�s�?�������0�V<m(@���� �ɷ�x���~�BS�D�K/�\Z��Jj��}
��S�K���%�����υ��O�o�ll�f��nI����G>:
Yo�^�Y���dA����'ǟ���3���DHh���.p9��VMR�:"�<}ǂU g��!����H�{���ǗfDo]��
�b-~�� ��,M'��|��m��%�0�d�m��|����K+a�;�h�DE���H �
2�a�(Z7&t��
��Tf�*�\�����,��#��i����|�s-�٢�L���E��"�]5�Ih�l�L�NA(�v[�e��}�Y�Q^���&�W�u�G��@׆�N�?/?����������}~N.��0Yj1
rW���!B���<����9I#V�10������!��#�8j�F�x��Y����
��}�Z��6;�kD����r/K���?q*c��|6��؊n9:���g(�2��F�9��΄}v�r��睹E6�ɖ��0� �'�;H���[�x�T�d��{����
.�~�G�O�g	��HTzn�O���%�Z��ٞ���JD|�)&�B(ؼ�C���4d��FAG5c>U���x�tA��m�j�H��O�<a�'8��+d��۳z!�����K4@HXx�j�<z���8���S�"���&*��3��E�������l]��9��;�Jl��.��S�:�;���N��%����i����WSD��қ��䅹�})���J�A�ڿ�b�[��N�͔ё��{�����\by��_�C�z���6�t춷c�	��<z=�?��L��yMs�ܛ�,�����b�t@%��������X�y
��?DΘ���&�w�7����}f���M&fb
9����0u�A��o�gT��@��]�X,��Q���t`���c$>�n4��r���P _�����(�e@W�e� 0e�������`8���n�.6�,�UAY�n�ēRs�)��{�����j��''7lt��(��Z݃�h4!M�L@!kb	��>�IHOM�B*oXd���'�Pb�
w4F���O��O˚�ZN��L*c���{Q��1.��m��@�|F-麟�8k{2����@ޡΦ��P�~�vdwU$KS�=*C�X����<��ΓEqJ!��@���*��{s�#\&�2�^�q9h����z�����'��}��Z�Ҙ�5����9iϓ[��ȍ(��F�����H,0�������h�˵j�i冾=3g�� ��/7F�+�~��nE@?>� &܂>�a[�OeS��T�8�J�L�a�\8�X�"p��ii|ȮޟĮ����\l{���։EX�15���rr$��}�)����ռ�FX�e�0F��SU�N[��BAf?Cb�V��KҎ��A�W~�5"�BU\�{&��-���M�e�$"����/g��\/k8�Cf�<⌣�-����.��U��C�}�]RU���]�ˮ����w]fߒ�W�R ���K�է�~6�SJ����3A��t�6��@W 4���9�-3����`1��8.�D��fEz,w�Q(ӝv*��&sd�����Վ�w�1y��d�	�	)EY[
��T����Dy�5<'X�X� ���:�� �gO��G秹���gg��d��s-�\�\] 
:��T8���O;?�sT����#]�7q���=;�:�M��[7���;|W���n��0��.�x/����Ͻ�i��QZ���Ӹ���6ϡa��
p�`�+��y�%��B��0�PŗG�l��r����u����ѭ؜�O�g&�8Lt��njZVv��2�"���&��*.��u8��!փ��+N�}��{U�pZ���:���W�О<D(�j$Do��X�|j��6��� ��h6%��{���cHI�&5��A�(b�������yUg�k����l�S�m��	��1_��P~s����Ny|�s`)T1���R�@6+ʃ�"Z�Z�_
Nl�]�Ɲ*Պ�6+kZ%nGe����K.W5$�0�f�:V�+OE�-{��Dڂ������uZ���J$k5�a�F<q4=���n#��]��`�4񚅎Ÿ�+�	V�A�$e���~����Wx拌���x+_�C C�ޕ�Ҡ�Vg�p7�wZ5_�"�h
�.��$#f��oN�OF��T�5x_H��m�Hd�c]�~�H&��<���cC�������b��>ݐbW
o�O`9���hw��
A(>��s-3]W�m��]�����]J8�f
p;��$-����uy�p�e�B�@Ks��<Ҹ�ߕ{�@x~܏����w�I���~��b��O����k��&�ry�f+�2v!�:��pCJ��?��U��0]��;a�9:+�U៹U�p��ם����'���TM>�@-c������V鸶��)�H�Sx�p �X+� ���+j���a���s�4�h+.�Dӽ�Q D-�Dj�ԩ�1/��d�dv�4v���6�ѣ���9��E:	��S�E)#�C�^ȶ�u��W����z[u"m' �]�8��)�;�sN-����j)�,� �����5������ZKYvs���;U �,��m�9���5� �
X���:��)�H�[�|�j��v�>Ǿ����e����C��PC�aU-1���8��MT"?�8ʚ��*uy�9(6)[���!`n��%%/a��G+���3qEϼ~:��5�F�1�$D�����I�XNN�lCC�zj.��~�}�3h��d#�yQ6u����7Y��Ԯ�g�]�4õ�"'�8�2�A�s~0f�;���N�xӎ��ķ�\ �\��ʝ��Qmox*��@t�7v'�ۻ9��>����n��$��ݹ7"F8�%m�<3��H��&7���P7����IL ��D�� �_`_�d0<�v�5�}Yǲ�?������?須�9�v��x�����m��EiT�{�۷����Z�L�ޮ�@cl��<��A�Mþs��^���Z�e�nƯ��䜝=�!I�h�z���'���A��aE=4�??�bp�#4g�#����(�FL[�~>��2^U'��X4rp��^�<��x=Դ?-%����05'��|��
�y��r�snh��B�,�M��UB��r;hT���K 5k�662�Ջ��F��*���7�k^�ʼ׿���Y�OFw����A;���0����|���[��qv�pBW��o7�Сy�o ��;J/����/"����l?=g5�g'���X��9P_V �;cïK�j�(a������b \�b��V̭��T24�����6�n	a�?�E*�HË���#�[�9t���~��Օ�>���紞?S�a���Qw(@���P�R&y�����؛�,��
�V�f]�H�K�$�gG�!Ƃ��=�:s\*W�U?��>x��� �[��2�ץR��}j`���|M��`��;{�9ۺ9��Zf��	����>�b�A�M�&Aw�4ws5�M�^MJO��-�"��.����*AƈW�e�[=ڊ8?�?P����+���o�pe��Uգv<E]G��6���^`w�&���3ۣ]��0�[1�W�Oa~���I�z��|/a7��x�Z�\hX6K�_#�J���U�ؓ"AN��
�O�
�M���q�\���e+��g�M�iӃh��Nw����t*� bs.~ebRk��8C�����D
� �kT6؏}�����Bx9�ͭae���0m ���`�}D�A�9J8+ DOep���;d�_��Jy��S�R0���ٜ���͡�ܖ� �9�~��N`�6��lg�qrie��
R�{�B��WC�Wa-�)4�y/-�WC�qi�UN���˭C�&��� �������q��Z�j���xZ:P�;�Fuہ�-��{�K!�LB��/�{��W����T>]m��E��.�'m.ХJK��S�Kq:������~���H�'�y����V�L�MՓ��sU��ds�#�e�7�>�J�j�0.����-/e���O��ջ�,�t`1�P��& 5eU�``u������㥐���f_����4�`��8���K?���jg��6�}�|Lr/V��tZU��l��E��f�[�k^k,׉��VB^66��B��g����5��d�V;+v�1�a���	�enp*^���Lp�H��&��<1��~mLn���9M�
�w������W�	�=)MLv�Ȼ�u{�8�����r���NQ�V� Vd�Gm���NA؜�����qN?������e	~eng�f�Qʭ����cA_�=òÒ�˙E����1�/C�F��%�	f�a%)�a�g�Vp�յ�#��A��K��qxP��.���4# ��K�n�
;Ȉ]���@n��g� =�/E��� X�0xmy�S4�߻�>��B�Xz�e�I�x��z�B�V|d9��W�O��R�s�+ V�'��P�����n��j���^3prQ�����en���z{����2-�qvs�ӹ�$	��b��-��8��k��zMi/���=	̼���#���p����%�j�V�R�&Q��O�UB���)�J�C�O)��[��#�>�,�m�3 �\�z(��}��0�²P�By�CC��
����Nq���3���u�����{��|ImX$7P/�~�Ҫ��,�Bi�J�����"B{x�7���X��ѕG����ʆʭ<��%A�I@��B)�W���&E���~�U!��I��o�oGjX�4��������|�K�[�I�����і��e]�U�~�-�\�'�xWQ]_;t��c8�s�Lp&z��-����L��Y��)p���2��bŴ��﷢�{���IL��S~���s��R�Ud,ݜ��t�!�jEQ����i>z�$:j䗻�}� �a�^�9Z�f�����vp�λb�+� K��OS���$jM�����9�x��j�8-%Y7l��!�K5_��A��o����nI���c_`�A��؛�;�)ϸ'��m��1��Y���� Z*	��߇�@U�G�VC��U9v ���kz� ޱ$��=�xR�ߢ�Z%����R��M�Y�b� cRᘣ�3��V`�h��~ �����؝Dx�I���Ix�u�ɖu�P+'�3�F����4�>?j`�QC�vݎ�����[�}@�dbL�`@�P�e��a2���H����F���-�Qv������2I����[װ5�k�L2��u�$�72�S���6:N2
K�����ORw�������n:ܡ���p�N�����`b�(=��~�}@��u�e87|U{�zhhM1k�~���Ȝ���F�ғzN/gP����f�@�䤓e3kIw���Ô	/���8ECi:�'���xDֿ�'�^Q�� Ԋ�m��{�pܵc��;I���)�%YzX�bG���p ���$�6�N閽C�~�Z�o�$�JYI�yk/��>js�Ϗz_
�Qɦܟ�<Ư�d�cz��}ԕgmT�2{I����*�4�@��������0�% ������{ꅶ��\����.�Z��]s��R>� jB&���w�lzv���8VgU�ȋ�����MNYs0��ʘ��`�y���
���}��z��E�~�yB���7Ƣ��������
��{��*�Tw����r��
γ�Ju-r������\���3��/j��}��2ʷ���x� r�z����7�%���K��`]��G.����<P l4����KT`�
��_�4[��G[����	>��]��n�0(�Jy�/_>�\ի�T���E¼>�?q|O�b�o�^���a�o1�J�!������w�D��4N*`S�o�l��l�UA	kL&�y3:^���ã(��{��|j��1���za�
��y�Ӡ),X���/�P���)o��2����S���Ҙ7T{����X��Ր�J�f����ܞ4d��\�����5'��1<4^�Gh#�����1��`Zɾ5�Jt���鷾�1�Z��j6ԝÒ�$���s�6����aQ�����{c /4p�J ��z�U���&�w+;wSR�J�1nڧ _>Ქ��[P�Z�a�}U7"���U&n3����ɞ���r���RD�l��o���p�h��d��ilE��ʶ?� �ڳ�;��ʔ��k�*��Y�_��5��˿������m�U>BolD)�]�[z:,���1�Z��К��A��r�mc�� � �b�"_�RXo0��"�WV��iVT��P�!\	&Y�+��l��Z������U;�����<u
)��Ģ&@ٴ�v�I�mY�hw��W�Ʋ��$� %�;2��i���[4L���Ė�%��:ܘt�\D�3�.��y	O+���N4���� T�B�1^����[��o��f����n��{%�A�M	��%����R�L����4�ϻ��%��Em{er/[5�N��3�K�NP�-�}O����'G�ܳ��Y��b�L�����'A�6{mV,����vh�2<�4M�r]R�|0X5й����\&5�;��_��Qd9�z;"��ָ�+�u=eB��#�t㖗u�{�vI6��n���:�b�ݞ��D (��ۋ�(��^�0n���V��cL�xk{XR�tY�3�Ħ�������H%u�8��>�+1�W6c��)r8�Ɋ���@gC�*XX �.dj�hkя���Fm� @��+ދo֛$�K���F��O[�Ċsi�EN*�����%����s�b��qR�G��	{�����e}D0�V�'��-��:�U������Lƹ���� ������i�d�9����OB|1�bxL,J�	��+�r$׺��2����xM~ߖ�;����`�C�Ց���ۓ���9>0ޣP��y�N�y��6�,���J��ee��ʝj��7C�ջjH���pmW{�t�<m>���~EE-co"� R9�WvĢ�	�����)$���r�Z�l�P�@ ���2��Ѿ��KH�-���S���|����4���.' �B �\�;1:�5�R~uXּ���$k�3]��F,�<��� f��Q�.���?Q΃��Z9�^K���Z��S�\���jR�>�Vw�(���~m4}j&�6}� ���5韌��T]�ۨ��Z�?���_&]J����o�1�rZ��)�$�������>+_���v8�tJ���vQ���B��m�fK]݅��Z��x6��S�`�dO	������O���8�������͹�6�x��<�o��cۖ�{yLt�t���i�@x1�c�	�DJ�k�Y(s�LD��J ����bh���n1/Ł� H��aV�>C�3�ЯM �K	��30(���#N��;vX,eS��&7����0 �h�2P_��$$�s7�F��ٍ�h��yi��e=�1IEభ���9D���~^�f�����*p���CE*[�1\�3���iy�l�/�����QE6D�����9�ـX�$�'���K2�O�f��-W޿�c93� lfÅi�dOw�s�Q�ġ�^����寵X�sх���Y4�.�G@����\�s'��ބw�n�ٱ�s'�Z�-�o�E�U��P�v�C���؂u����u���<��D:��!J�X��,�Ԉ���W�)��t�fI�nU�z,��q}�Q_ƽ8�MI���1� +ʕ@���iVGJ���Ѥ�;b�u�o3K�S������eDP��� �T�W�x�S%0T�})�.�2倻aF<��7R[t�iA�)/ �G2"��/|��X��X"ZC�&J��jc���:B�u�"Ҹe H�#�!��.��ܮ�)n� ��>��$����
���)5|Y�%Xc%�P~��O.�^�"K?l��;v��I�R�N������U���BzG����!	��#,?N���w�%��r*��7��m/����K�ϽS�C��P�mOȴ�V�E޵C[������|,�����Ax���w�y�Մ5
�rL��Q����r �XU�<z�P#�:,6�P8�M���~�薊^<�4��k�g�l��ʍ���4>o�{{��Id�ݧ�������':�%�4���Z�� ��W��J4r��_:!>��3i��/�3V�,N�:�w��o�A\�3�ڜ���&.f�IG����.:D�דYA�ԧO��l)�v%܋�K��
b1��c��4_���̸DP^ф�Wf;�w�=�
�c]�*�5��L���3z��Qq�P��mu���#���wV=���Y�οy�T�#�7�[E��M��T�p=j��/��w:)\B��Nw$a/�#��۠ 4U�
���V�*� ��B�z��G���ϯ�y�����q�GD���B��.��o�Z�Z�g"i���V?���⧃)��	�2ktN��!o%�y��r�3��x����5�K���}�=@�5��z7���G����*�_:`cK��|�#{�s2Uω�_#���=TJe�vg����K�R��Ƌ���Nfi?fM�1UH_s?<�K�ؐ��Ql�y�4|��h����
k�CŒLZ	ovsc�-,���|ǚD�f1����#&h�1F����;�H��.��GV�*��p��|���V��������TDv����Gu�9���J`5oUKO��?C��?'� ����!�cK�I���tr�A�W����;0��i���,�{��:)��t��.:��A,�x���Dj]Nq
y��.�KՀ����˯8�xz�5kd*��OD�yP��c3�	�٫����L��*��G	�����7U�EᓖzV+�X�l��YE�i�r.�c�Vk�@�o�O���>��B���99T,A|1�[k����o�t@m�H؟%�q�XN>��e�i�x޼��d���	'��1���V�&�� 㮘���7��~���z6ᶤ���q�%B�'?d@��>��)��WO��$�fi&H�S�5a �rӆܖj�E���qy26��ד�%E�t��1~x��PU]+GX��ET�,.;�:a����o��|�i��&)G��5���i���E��g�R�n�A.���/���NejA���k�����\��cT7��r�M�T۟l_�MS=֦�L����М+d�P��R��S�e���WB~P�i���c����_p���-��vY}��4�_��SZ��-�F ��%B�XA.݋��^Ί��#Λj�����y�L=f�%�JIB���'��du��DJ�6|�V��Βr��qq�3txa �)�t4�Z�O��
�|�o�A,jb3M����
�V�Y��1���H��cA��f���5u!�/���/�]d�c֌����*ړ�ߝʢ)3���{a�zx^RZ�v������� ��.��ְ'zv�k>J㼜X]�N)�ކ�佪��"�#�RiAO� ��M�a�|��/fN��S��Ť��z� �lҘ�"�*�fwlN��������٠�aJ�h1�P R���񍽐��`WQW!�:�'�J��rI�\j�F3�J�3�`齬=B��ݺ��D�>�������é<�h�B�t�^<w��;br]W�UJ��E���tD�U���t4	u�䧢�O��[�HO5IM�y����TO39H���L�m-ܯ�rcүa���Rb�������t,���B4����m������`/r�[N�ݜ�[DL�`�������~�J��(�K�\6���F��fx�8��� ��UA�D��E4��x��7V�B~�a^ID���1�/�O�lN[����`}�5�Z1�w��z	�9�&n�>IL�'����={)��:��JM6�vJT�p<䱝W�o�dS��s��� 7ЖW����a�`�QW`��4Oi.�%�0F�I�f�ʐ%�%�$}5�ag�Wl4��^���� ��4f~]m����q�NlX�b�P*q*���9>v������帎�_�ez�C�g�a �e�MO�K^�c��O��]���drNE�"B䄬����cH\��;6�'8Ŏ�gᦾ�JJ{���Q�|H��%�^�{jB"�ϭB7�>;�>c���������V�P
�Ŏ�mz}�06�yȺKp��^>	ќ�SkD��,Q8��������gH{ ��^�\م�g�gb�����o�6$n�{�XS���xU(O�d<����-��j2�p���_��E�oTb���{~E�%����X���W��`�zVg�j���<*�<�:��D�S��<4n:T>*^q��"��%�\AQͧ��z~s�<�.߲�N�����&�[͜��,�����Dq�S�(��}|�rN5��t}b��V���t�D��/k�NE,�eBнpLx�d���VW(�GAB����V=ᅂ��	�
�{�M�����<{�H�D<�Gc�ve�f�^R�3"������4>d�A_%��I2��MK���MJ<�؛S}���S����=BP�$y5�����F8�]��_3�J�5|����� ��3	r�c���_����'�a�T롧Ш�~Ƒr��RF�G���i�U�2�w�Cq��s���>��Ç!/����Ť��u�`����r�k�{��\�oY��YdOx<��Ħ����m)5tezF��:�$����|c'n_������
6��z�?W�S��+���.�+�e(�o*"}��A�*����-^[���-f!��ޓ�������I����)h�Wc�ŃA(���%���쭯��N���-�h%��x
��3��G�.�����E?��wy�cpKu�3b�;�l��Մl/K�q�j�"�(j~���/K� �32�}�e�#��C:��7�B���ב�!��ꚠ�ˣfp%M��ߊ���gq��b«9~��f���&��S xw�cж�q����^^�[T��-� �P�LZ*�o�C��V������UZ�������k�$�#g⌀�����R���严����g��m֑��a���p�7�� v�%�3�_P)��� /�]:8b�����|N!b�c
�!��l�{�{�<�S�����b��ٍ��Ș��k��NH�al���r#��v�j��K�疓������� �j?���M�Ѡ�I'��$��,>. O&�h�,�$��]�{�� 1.V4��J�E��Q���\^�*�m���j1(LH�G��!�A�9��l�6���J�F������!Ԝn�f�O�J�t��e(L����j�p�m»7�f�N�4��O=f����7H�Gl���Hl��j�������xIZ��'���F��)�4W�m<
�m߫�C���Q{���I)�~�(:�s2�~9W�ɞ���H�&�nH���i�f���"u��(�<��F�Ĝ��itt�.(�O��_׃�K�RE�=����OI+���n�c�[|ޭ1����[�a���C8Z��ҟ�m�LD�ׯ$��()p���?���W������UÞֽsdY�����'G�8[~�/�Kq���s��C~�>�D��O�m�e��98�C�)q w�&����1=������(�7��zJ+;�
;I�'o�:�C�Sk��<l1�t#�_��
v*�����B��"f�S�^4���a4��B��b�[&,���¢��d�u޲ʥh��p`�?�����ЫX|�JE���N����Y)���WB��4�p¡[�9;+��%9s��H�t%��H;�]�8?��}�����K�ݰ�6ҕ'rD(�hc 	���7��p�hҐe�Z�k�/���G��IK)h0�e��n�$���������k����4���Q�8����14���>�hff�~�b� ��tUM`�C���K}��j�O�!�&�Af�E�!�j�Kn��N*��[������k۝��j;�6ǻ�o� ����*�'����2�AT9���̓�l?�I��ʆ��d�P���4�s��T�\�=���H��9��P��z�f�ҌxeH�~BW�}���3��H��3��/������xbd�^(�k�ͅ�-�$�eP#d���.{�Q�:ª��5���'��<��.���۞f�SSH��{��k��vC�7��&Ry��>4Awݾ�(����6�s8�HU	�TEGƦp3�4G~�6 �y��{�KOrC�U'�d�jW%�_.���EǢ��&�����������toO��-j33�#5�� t���+��9ļ�!���s*#o5��Ԕ}�u��.o,�4e:n
�U�Ů�O�1�߻6�[���Y�JU%�#�u�n?����鴎�ݜ��1�t�����4']��U���<n7�߁>U7���j�_c/�6(3w��H)G_���
���.�Xm�(Z��FS%}*���
�I*^k���>av�O�}�@�7���?�S�8_Y:���%���'[����`����V"%R�X˫L�u�%"����eL�AP�2B��� �T]��YJ�ε�Y��A������N���<�Q��]� <#B���֠�h�&(�h攙W����`*ò�j^���ҁJL��ۜ+ko��T��-���!��^q�^B�צ�J�����pJc�b�eUNͦZ �-�pu��4ej~抬"E�N��Wӱ26�c�u%�9+��o��i���!�M�x��CLcm�wϢ�!G��8�j?>�������9::<�����m{dcz���XDx�3�Y-9�*�2N�NW7e����ل���VKu��`�tޗ�yC��n���_�y#�GI8~3�ak���@��v��-m�����������P��k��z�"�Q�.4ea�a��(��:���`"}1�Mn�bW7����Xmn��4�W���_��1�u�\$�f��c�`��dc�lM�˹�]^fG�b��,����(�]{�<�s�v��7"y%��
�8�t����qز�����>q1t���1_���{~�k��M=:���x;�݊��g��P��9�"��!O>�H!Y���',3���ܼ�A#f�g��h8xL�DH�Sn�i�FϚ~?���]e����Bm������<q��J(����˰�z�n(�C�9�mak�h���]�*�JM��R���a�(u�+֟�~ǚ)MH��P0�$٫s�k>�:Z���4 /%�4��������{Ȼ]����B)	Mߺ�� ��j�z8�.׳N��_�M�ф|�:�t�qN~�U��q3�A| �e��m�� ���ڞ�x�,�u��?�Y@2�Հǟ+�$�4�,\�y�!�D�0�e���?�Y����y����f�i*�? 㓨,e��BA� 9��a2�����*VZ�O93��Ѥ��5VO'����n�.e���M�XW�����V�T��ܜz:yj8-94�ïcP�������ٝ��~�by���0���q�f���D�v�d_����P1���k�\�S�$��XGccA3a����~���Ww��z������]i�6�e�)�;�g��ՇK柬�}d��J+��M��Ⴑ���X�Omr�O�$��r� ����8���}�S,����d�ٜ�cG1�j:�����ݰ�r3h����y�HMn�da5����P%�Mn~���}����=�je�Սۀd��������k�/օ+7�p}M��<!.:f\�I]� ��Ł�ڄ��޴���u�"߿���E�*}T"�+�\�B�����j�#z�f[���t~L�.K�O��ڼTT���������*Lo����Y��(��	7V�ɧ���N�nl�������ð�� F�-/����������vR����K ]ɶ|�T���]�.���R���WtSj`űAtc�Y�;��y�����E�,�`n�lĥ
��s�B���x/n��m�q����9v�&�Q˹����Z�a1�(O����TN� Bu�����*CU7<�U=bf�jI������"Z@U=lI�RPk�.��NG��+e��U��_H/����y�1ޑ�O��l�k��ѵ)z֘c�e���H[&�(^���P���z���:	��p<#��*_W�p~�^6�O]�2,�G6���Kc<Q��hq����E��[�b)p�5����,�Vd�����R�*Ȫ��	5�����b�B~s����H�?�=�e��Ԗy(���;��g�I�e�0�p���BK�ȩ\�,�����ck#�����@�Ej��ۻ�nw������c�G����}17�-D�x,�F��C�i�=��IłOH�i��ۆ�˝�TN5�oֱ�M�8pR�l
��N�qw��F���Uq���FޥH�T�?˷���;K쀝��΅L�C��*E�ίkk�5Ǐ�-�ߞ����苓��{4�����,2������x�F8��81�c�vx�08Cw<�~�M幾��.�M�p^�Y!��t�Đx;�2���l�Y9޻wӅ���h�^=��x�f(D~d��~����3�hP�� [�i"��r%j���7>�_��$���V�[�x�&�a��^���y4����7��K?�����40���[ c8�8u8]1�;�`����x���ܗ�:;����y��,�U{�qH4�E�y���>.sb�P�L���
�,�w��z�]OH���q��\2�g��a�^��p�U�pSx����oȻ�+��#,	�}$���E�e�u����!���s(=Rӧ@U�Y��CkdM���*)Bv���3;:?c���}���tk�Y��b�c*�3WT����ӓ���bx�&ε�Y�5Y�����Kl�C�&�������8EweT�^B�hdo�<�� ����g�����N��$���O[�Ƞ^ߤ��}�0��&����i�k���Y�8�Ｃ�&�9�5�V�����������(�2N���{��kiL&�-b� Q��bWx䔑D�ʆ%Kͽ'(| �4��b��N�Q_��� x.H�Y�n�v몖��r-��\�,���ō+��Prb"�o|���p��n`�L\�E;���mϦ��yC�T�{f�]kC�zhg�	L����/ �R�����v��rܕ�^��e�2u�D*I5qVS�Usi�P<���_x�um���e���~�y<D�,&Ѿ�F����^��p\�l��ٔ*
��)k�l�y��R�4����e�aI3��LZ�q���[t��uF�%���J���ᷢF���\��h�-_H2)4�2��zd
r�1M�� Ŀ��^���W�_}qT\Q��e&w�9���7�ג.��13�J�89e��>L�"3(�Z?1Ҹ��bj�9#��r0��i��(�T����')N��{��7˼�C��Ίñ�v/4Ŷ�%gU�q��	/�֝�e��������K��N@~�� �-֣���p����eC�%Tf�"ю�=����;afC��FWr��������U�ĸ�!wf�w����2�*M�g�sw�BO�T���S0�WYR��,z3S]�=��@8����m7D�\�^�Wy(�j�wK���e���r��gƯ�cYIgPD+�9K~�O���{�:\�!�p��o��(����l	|X���'�&o6" 	R�C�{�/@d`<h>�
qh�ޭ��[���V2�K�r邈��S�le|�x)��A�`9O�;�ĂT<>O;���Ϳz���ڳG����_�;�QZΚ@��^�j����Hȍ��RX�������� ��_�r���yb���f��B�cK#|����ؽz�k��z0��s�!ky�I(^�*�����٥P�U��+O��8��9H@�-���t桭����,��W~�}@��i���o�7�C��n[�h�zRo���91����G�sy���?�=�lH2̵������R�}7�+'s��K�9�g���`�݌�Aͤ�8�l�.r����#0���*�8�y���k],Tn�1�����I�����S~*�Kt^)x
�i��x��ȵ�>~�.���&3�۩o������.���z���h�'3x�a���猼t��u
mI9*	���i�+>C���ێf����b>�r�x#26��Q�G�9������;��ϙ�a��Tc!��nqD\S^�F���2����yk4�� A)%��R�LO�#��Ǹ��1�)S�s��Y��_K����b��S�;ѐ6��3�w9���G�/\�	���f��(E݄�囤/�+xMh�EŻ���$s���t ȒL>U�Ϊ
n&o��i�F��Gc��{Z��?�g��L�څ�|ep&�ъٙ�Pş������>�s���6�F�^͔`n�y�q�ᘢ8d��N�,@40�4�QC��wηQ�zA>q�#���Õml����t�@�b��~T�K�^�1M��� ��v�`�}Uu)/����"��;^�#q�iPɝ瑹���Pd�c]�3,�4ݔ�EI%����� 5��۲�}����6��JD�-a��k�gv��CF��cJ�X6���Ȼ`j�V���?�od��"���u�H%�r�m��@��w7�	�C��O�b���9p��t?9WG9O��|�0Wk�Cns�K���ݰ�L?3�'pW!w��P�������`�Ψrti�B
�`l!�E?��8M�����߯����F���>������<���cf�E>Bᚃ�#�Ϸʞ+�Z;�3 �'�aG�%��{B�b���)��d+�{�`��D�p@;��%��I��D)Cݚ5��}?-���`wlx��<�������aC�R�)����:��IP˫�{v�u�.��9�j$�s��Zy�r�3��Ԟ},��F�&��5����k�H���JpR��Қ3]�P��e�VQ~����I��p�2�F9R����^��· 8r˃��:ɶb"��bZ`ƌP	�^��3$қ���
�r%Ǌ�k��߾Qh%����^��#i�y���*Pw��̶�y�$8�:|E|=�^�����1i�M�P�X�����Eugz��P�
�6f�:qa��Y��
>Ud3�N��`H�2��U�j\���Y��u_���)-l�+P���H3�~�5����`4�"p=�1����q_`��>N��xU6�03-�e�yK�n,ln�Hs9�Lқ��[sa��
��[���?�\���P~�U]넼a;������,����t�oʄ��)���q�W#5l�31��/i���3�m6��G{�����>�Kv�B�M
R�^rbg����n�h9��;/+�\��W�,IO�vsěRƢ�ؑ�c���/�=�M(�c�on)��U��x&�_V��'���Ea`�1���;���i��@��G�� �kF"��>z}7kc#QŹE��/V_uԀO�Y�?���Nf��Aɵ���"j�,��`��͢E�6i-О5v��n|���H�� �Ȗj�?k0�[1n)a0=�jER�̊L�OOW�=܍�8���:ѷ�JRz(jM��J ��$}7�[�� 86��5�u�/'$i��cO�uk#�x[�2�7��϶�ۏ����\S��F�:2��蒣���%K(�g2$ԣk���h���*�MU��d����	��V�ӎ���(�����<|ݝ�j�ַE���\���?�&x՘0�d}��\)���&x	����d�)�1��_
Uqp��/}��R�{JY�ɋ&���f����gK!ˡ��[vΠp�pw���}�����l��i�(��6$r�
��A�_d������K�p��1�����٪�Z����ZfC'��>�, ZN��
�Юh�cZ���!��m�0?��.I"�<�Gv��C��6ܪ�*v�8���Y��|p���@�)�l��CyAy��) �D�THv�����$���������A��1ۊ|��(ԯ�f�����Ch٭;܉w5�21}�iz�*�ȃ�P�PP��%��U�T,"w���ٹr�&�7�ڶeb5�B&r��g��l�_�����`���VV�[tl�.�� Y�vW7�z8?�o���|�<�<�X�.�ϫb�E�S�l���];3_��d\&U,X�ْ�]uYg<Q���.�q+JdAU��͠T@Y�qi���"R������lNl�nJ��F.����� /�!.g�Q�)tծ�&��#J����ȥ��L~Z\����c@UnBP�n/����2ꚜ������J�!�%-�(%�����H��%��5�P^�}�7	�p��R�NP�@�F֣�T_R�/��3��9�]# ���m���
���0"O��_�Χ�|qG<?�a^Ш�MX�-o�\�5�'����^��W�ITm%��|�i$2l�)+���G�c�pb��S��[eo�7�K�w��7:N<CDXM�2�M�'=��᧔{��߳��9Ӟ���6�tg�ݾ8�w���FO��(}��I�R�'@
f�b�g ��!T+Ϻ�n���=��Ll�Ȉ'}qbx#�Tŗ���!��T׭ž���"%�nUT�h�*�v⼆�JY��}�rn6�now#�)VA		4}Fqt��1�H1��Le�*l�/bCF��Ȝ4�A�ή��;)���1/�y�e(�#�O��V�ݞ��&c�k��V1v�GC�q��r��ny^�$��ܬ��E�y��#+�~t���s�]�Ʋ1S�0�����e�VK�_����'j��Xf��;S���c>�AQS���q�] f�*���̱��.�!���"�Xr1K��� ��5ڦ_��+S����,u;��)v�������`7�

��,a�/� Ҙ�z�i:��pO+{]X��;������;��&-��� )0{*'�B/8����?���Y��$��]�nH�s��PS�����M��p�K.��z�DB'�3��g����?�lu�6p���*�e���O�u9{=�()�����]-��ь�|rV�ҡ}��~oZ��%7����V�z`��ˌ�0-��Jt
>N�(����>d�GlJhO/~�$�D��L)P`�N�73b�_��E��x�z��E�~�ִz��T��+����Wr�y�	�:W����D�L8t��@1�'��[��5���)J�����z������rQ �����I�J3Ł�:? �3�aN\�AR6�n�	dT�ɬ\��ZT��J�ģC&�y�~B�G����/��P��������2�B�T酚�']!�	|~�%(2%ߣk����F(���{���R4f8�b50Ǚ��
LD:J��_�/u�F>
$�m��		����>���>�*��g�m �����n�~;*Et�܆r �;�'޼��3S�>0l�G�VB��փ����HD�Å]�W@=c7��h�#�^���Ʀ�.�s����L����L�i4�,u�:�[�FpE�\#�'���ɥ�/�=���^w����+3�d@Sr�;�c誨�y��� �u��R��c�/��]��S�#���ߙX1�l8�t��/#\����̢{0�e�ز0�7�.ZwVL|��@/~Җ���ˉ�p(��e��'�f.Ju�{�g��B�Q����O_19Լ�#�ٺA��YѸ�c��򊥕���>�����m)Ծ��(��z���u����R�6�XF�2�hؕfz	�F�9J�
�\<��j��\o�t{�?4�v�A/<-o��t��%�	M?+�'Y��7������Y+���f�f�p4�K������Џ8��Yw��̈���	ī�foJn�~���>��-$��oK!��͠���9�&��ɖ�� �!��s�Ɛ�o V��Q*)36�5�C�����8CEƕ�&�%̟�O���/�s�6Z���e*��v�!E1�V��hB4����17�)�"�gW	j@�u�St!9��w��[�UZ��@P.��oqN�=¿_w��L=����1_�jw�~u�2`��Y���T�f
����{Ŋ�ݛ)�X���-�C�>���;x����[j\9��#ݶ�Ȯfz�����^�0��� A���±���a`}"�����V���g��_Zaφ2%nMS�T�4�F
�Ѽ[��	�'��L�pX����|c5���YiT�!�f��gf��z�"��E�B�<~%��J6���������[t�~��.
�`�v���纜��Y�F[{X���$?�V�t�B��_��n}�,���Ԕ�Ij�l%���B�\�zL+w;a�|������K��Lm�U㹈�5��6ܻ�� zգ��c�2�I�������G"vP�:��͢�ה�3� J��Td�u�݇Ȥ��o����������*V$2�BN�Z��G��܋K�-��"��0�����K�=l{�z�ې�F
��d��}�xt�^K�Sm���|\��=�ԡ��؛��g��Ǜ�O5���dS��1�)��UU�)/��"��X��wC��r#��q�#0{��Q�q$C�A��2�`��9:���V�r~��u8�y\MJb-��}��a ��q{+��?;`z��k� ����Y,�� ���o�x���sI��/ �H��s"���6�1Ԣd��_`��J�f���:�{W�j�;�?������(@%��͓b��5��v4ו+�� /�l2��y���*$Q�f�lS�����(vJG�:�v𥛱�c�ZU��c5s�q^��~���q�1���3xk,'<j(gWLR)@�+m�S����s3D�ϲ�Af���ڞ�n9��l.hѢ�`
~^��쯭�h���X����D�q�,�����Ejz�@_mm??u`nd�Q�l*������K0�zi!r[
�4�����N*e�$.�r�E���=忞�md2U���85�V�>�$��U����q/n�{�9'>r�q�%��[k�Us]����#CZ����'M58��߲ct��J�F4������(H�M����D:>��-
Һ�~J� �~�{y����}���S,DLW5|S�����FBJ>�P0C�8P�"�+�b�*��f��p=�Ƭ�"Ǡ1(�Y�>5�{/,6�^1�s�
ӫ� K�)��:X
���xZ��<��6=�l�����i����j��70-���e�Ac���}�y���x!�����Ui�ab�)8�=���<f�Dq�'ߎ�� �v�w���b��Ҁ3��Ԅu��WPsB�����D�,���������Ǚ̀w4pߨ��E�%��j�mQ�?�#�vH!��S�bґ�����&��bԸ�ٍfi��[�t�s\-�A�cI@���\�͐ZNA>6F��׉�~ɞ���?�O�k0�� ���E�����PEO(�ױi�O��$m�Ϝ�
Ѩ���v����SE����.$�S:Rώ%��hSQ�l#�8��>=ok;d��:H��(��@J0�1���1i�=_�W��U���)_Đ+�ν�!|^v`s�;��!*`ݼ�M��Г'���!�A�����B[l�^~l@�^6��LndBF%��%b/�r���^���aĹ��0�z%m;�Rt�t�o;#�I� ��!��F��JBix	���e���.�u�Ŭu�!<�̆OC�Π�羒���^��0k���~Mj�w0���Y���<��S/ނ~8�]��24�{?�>�j�v1~�����f勐y�����/�����c¿/N�'_�)��M��A������L8��+}�X��m���G�;f��v���!BI�X6�P�kf ���`p�� Ϲ�y!n���%`x�2/{k�/,�un9W����H�W�������<z?���TM5M���|d��5��s�?Z��{���?^����
�)U�V��o'Y��tdZ/H�T��;T ���L\+�d	%f�n;�ӡ
�+l����B�%�{������P�1���� U;��~[Y��c�H+=����O{�C7V�$�[{II�
S���r���\#��	V;����ű����/*�?���q���k�6��qk$����F ��`0��k�4���U�f��T�,~�?=�ȱȸ�;J&��u�peH��D�H��eE�Fsh�"�D���i=Q��Q����3��ӝ�� ���9	���c���D�ȳg�����U��,��qk���:�ZF���	u�{�}�{�O`��Ë-%���ӝ��8F�ly|d���1*��f�?���&�X@���N>���@��������1����W�K��}M�.����a�������-c�
�1�/�ޚ5�t�(I�gk�����w�DJr���psmd:�rJ�o,���/�a�+y�?a2�/c���т(��8]>sh���ZU�E��O��#�*��|�aN4$�υ��؅e���O�l�+�^'��W���Q&���e�}<S6���1營�����݉
]����WK��^r�/��|��D,\*��V�{T�]���H���,:j�L5��K�j�L�ν>��u�W����1B�^�>�%�?k�Fd��І�r�ЫRtq)������ؼ;t�,��x�YuB��4{Iqj�i��z�J�����]��fq�7�\Ĉ�N#��Q�*ҙ���ɖ	�J�t�*TE�,�s�K�o{�"Ҫro�_x��W���l>Q�����4�$�T?F�j8
?��I�|�u����#�}�c̲g[q�Ni���F[�W�������W8w-�J��1�0$']������h�� ������K�r5�k��g� �q΁�zeB�������,�k�H���L��+-jU���m�U�<�2�o	.� ����"��7B��֞]��ku���ߛ� ����˭�	�ȅ��z���B���U�e���M���:���7���'�g6��Z=�C�������*.���z�e���_ɰ(��GFcE�7E΢��Ǝqv�E4α�=���5���"g(|d�&�a��q�Wޜ�!����1W�+�<����&x��8wj��^��m��M
"�F1c����F��2�F�p=�Ee5k��%HHY!�x��i`���V��`���}����x:����R?�h�%a*��jqA
0#�<w��,�'(v�L������gj�E�>�y8׈r�_
\�C+�
%��gF]�_6&lq���
K�ͭ�a�Z����B�dvL��-��:Vc�O������q�A�(��9�?O�>���s�!��E�_)�N�~:�Ao���d�ID�ب��Zܦ��ͪGwZ�?o@�wK���@5M��N�7�V���ت$Ԫ,�;��.��#�4A<���@kHi���i��~u]�~H)�qQ��˃.�y�M��K�}�j�QI��lpm������QZ��fRP� /���m��[�=/�X����=�J3��oļ�wZZ�Yw��V���؂pl;���h|�(��������Bl"���n�I�q|�233�½���h��%����p�"L��L��p�<=,��N�E���][�W_G-O\�\c�n���� ��zx��Q�D�����yZ�	#�j���r����K�؟�6W4e���s���^{�L���3&���&�`gL�OÝ��� �q1W�O�VH'v��AbHIj��g|�<{�}�MԜW�ON���N��%��)_,C�Q��Q�嗯�i��%:A��^�����*�ZkJ,h쐏�rca���H��7���_"P�Nū�t�Xj�ޙ�y�w<k�ɸ?����bJ�)�ɴPFD@�	�b�C����΍�\H�k�7ی
����*���;�17L��{}I�K��2t�8��������c�^Į�(�U[�KP=�J�Z����ւ�!U�s�
K�����#�5;��Ic�~�0�: �� ��;D	v!wţf�8à����L��*Vbz�#��I���s�P��q�c��z�H�0V��E�-�uzq�G!�� 	�zآ��`k��1Ƴ�|���k��,�4]��z�_�&�<7��y(r�cI#�b`��|�����|U�Z+xG$���ֹc#���Vr8���m�8����������ah�QV�
b���������d�|����#�}����+r�">l��v�� ����c0��C86�9:/*���V`(��Ŷ��S��ޕN|G�6k�_{��3*Y�`�����8�lA�">���
�Djō�~�)i(I��\�~��NW���Q��
�l����t�;4���oj^��f.�����A���&��F\ n�I=�)ش׀��c�6B�_���P��L����4�2ú&��:�{�{��R7���'A[WU�
�O%����z��E�
�����eF��~H �c�҄'� T3	\	�Vu��\0�g��;!`?��ߍ���ڦ�2l����mnmA�$�co;I�Q]dD�����F�I��>��I�y�v@�/n�!��*������l-H?�����S��+�K	S� �Ϥ[���j�A��һ��Ls�5放�j*��M�`���ݭ�4+k��[�fp��E����
��3�??��k��p2��5�ַZx�#D�W�3� �4=�} E����e�����wa�����$J<;�V�����o!º����'���Հ��T
9� �ְ|,[_�C�\�	�Y��#��F��K��g�E{����������r�Tn���o�u{�����d�1��'۲�������SS>]aD6WI5E�#��5�h_�a��G�Gg�/�$��]-d�oY��,��c}�7d�
����9:t�\�(��]Ar�0���!��p��G������E�[�,˶Vv=�W���I���R�׏f�f~�z�ߔUY޻��C������tT��16g9�n�I%�Wt���|�N��̗q�Ux�.(}{�	�R�l����dkV�9�`)��FnX��D$98����[^�����'�j�|�*i��O��)��?U=���ʪvڙ�J�ŵֱ!�_-�y 7!�ϓ#�����C���!�Q��ڻꮑh�L$!U��C���ǽ�o����"L"%jWjr Q��4��	��>n;�F]��ؗ~�� ��7J9�*���(_��Q&!��}�V���G����]'����8��=��~9A.ƞ/ڋ�8}�pѧ�)�gxaS~ߍ-;e���
��u/�5ø��)<��?��ͅ���;VK�>��=�5.sy7�ز �H�jAK;��ZR/Gjv������七�!�ޢ2(#�[ԇ/x���]!#���A1���VyԢ˷�Ha�Q%��hm�" ��9)��Ǩ{k���a��.*��Z��k�����uEN ����q��E9D|�1))D+�tDT�d��5���d`��'p�O�:���|��-ϟZ���X�V�!Y �Qq��Zd�#�^W7�Q�[���0��� ����)OV=�S�E��9���P �u�_�?�٠�N�}������hDk�1T��i�+�[�L�Y�̞@߬Rs^��Ϭ�_�n?� kZPø���JXfn�O���3��?̜ǁ�%�X����f����I�P�a��� �u5�`�KHL�O���#9���]}@bl`��#��-��Y��.��tw>aOx�~�"1@����X�+�T�����F:��0�O-n#5o닾_S���S����ZTAb�-�ɝ�n�*�T�G�$�����Ֆ�?KpV�/�$�2�"ifr��� JylB.�u��eFʣ��:�[�T�]��+�O3m�s�Ġ#��9n�C��
���j�i���V��|�����j�h��\�E!�j��.�,�f�ZDť)�n>�#��K���4��=,����	����~9�l �P�O�ɯ�ds[kP#��E������0�P|��	":\ ����Vܫ�J����@�P��׹z��^Ӛ]�8L������&�DR[s���Rj��$���D]°�l�ǡ�1��+Ը�9pQ���{�#����g��M���s97|B#��a�Di���C�*���v4T��u���q�"�Z_5lw� ��� v"%�H�N��u�!��hQ��\%�z@m���{�6�TlQ��p��"�y�n��ŜR�R��%�_ZL�����ֳ���=�����^$�Y�BJ�Z�3w��:b��f5މ&�/8�t	\�P  �D�z�0��S�_z"�J<"�b�5%AWzby�%P|�Q�.�5�"XcvC�5պlԔ
EUz��&�~ƈ�",����Dжœ*�]���4���^�vT�=���hy���ܰO�G��O_[{��&�L3˲���<��NZ���w�L�'O���@��Һ�$7}���tZM�1.h��Y����;@[l��ZTo%��+���P�������o�#W����	�$��p���N�;��oe��يr���:��Ǔ�c��3�]���?S��Pb:�5&}o0ɀ\�ΩSCO^���q�V)�ha��|S��.�L��	'�H�8��ݼ�M�-;u�p�j��o��!TX2��AM�Y���^���gr�e����s�e�OX���u��S���q�o�&�-��+��Ƴ�� �>%MA��0Vy�Mf��w8�ʍxn9����)Ñ0=��:�����0�0%S~
%"��W`D#(��?�Jm�a�Y�q���S���Lx�_�\��=���$в�߸��/Hk���[3��b�� �L��ᝤ���K��&�ҩY����e Y��mW�z�������/H�>s}X'�7+x��E嘋W�.Ҩ/�v�-/t���:� �5:[vY6��?FF0�0�F	��;���D����(�g�#�Ƣ{����^��3%��V�����g�2����WW?���|SJ��׏^��2�c\��T�2��`qGI��!|�T$iL:A*�@�_�V���U��Ph��>z��g4���A����<�_d�����&��m!�^#b���Z�����_�Q����Ӱ��-r�L��D��k����1�f�N�i+H0�v��	���k{v d#�~�loi��%��O*i䠯�ɞ��Q�"J�fw臱�S��lZ�F�՚�	܊q�֓�E/�Kk�m<q�j��:����i�q���1�Ft��Դ$�]�
h��1�T�Ӻ�C���V�aOB���2O���)Y����<?mϵ��C=�*NyJ,F� C����@�d(��d�uͳ#7ѧ�τ�	�*�_&��8T��J���"���#��Gv���z� �������c�]�$㫟��FF=��P)��%�n錻Pf�U�j;�M��-�-�?��������q�l��W� ����ggh�����-+8��d:��ۿP��R�ɲ�~�|���,�K��*z,�yܦ��:�%�����$��Qq.�|W�Z4�9�c��qU\��:�]J5��@您Xu�L�2$Af-u�!Go���}C?/�CQP�B�FX�����#su�u��5�t�7�� $t�֣�ڋ�Bh4�f����[[�7!_��n��Lg�����ZY��^+s�YQ�Q/���M	��AК��\R��(O#����j�ܺ���_2$������U۵�@�`��M�< ���-��t��nl���4r�a^�w.\{�Ȥ%t5 ˑ��Y4A�<T�b����X�������jx���Hh2�;� ���S����up̭�4WK ���c.��)�y�ٜ>�ϔ}��R~�{*r�E���;����.�bc �\���ִ����M3^�Y�/P麊�r蕂�	�t)�\f�H�,�n�����GȈl����0����6.K���m7V**�I�&�3$ak�)t���e��C@�|�
�rL�N��-���;�h��n���A�
���Ak��Z�Aah�DfT1�:�B;Ɏ�ߑ\�C����ɇ��ϝ>�!�P���U��Y%� ��ȑ��=�	<�5�p涖�Zd�{�9u��s)uQMy�t��5mD~��'��&D��x�Vb|�Af�Q������j��2"+D*[d�#Պ��J.��J�J
�i.ˬ��]/��N^xg����㚾�n���W�����ye♵kv�����ؿx}<�Iœ��vh{A��\�{��*���-�dv�P��o��7�e`}	{�2�=��x�P��ⴛ�ߓ����u\�r�xlL��!��:�bM4���������6��p���5Ϟ����sK�
*�4r��f��6|�������w+��k�S������ח�e[4��U�C�z��c����0��2�h�/''��m%5������hO�*e)���}zv��,�}�	�lQ�M��^<��\��H^���czqY�.'�ȥ3挾6q��W:=��N�0oj/�ğ�H?�\:��J�� ��j�_��=�ćB�	���c���"�מ�$#��xsO�'�4	��?���p،��&O��@ �"4n	i���sV0����
1o���Y�fK(ќcMJ��c���Ά "�$�}���}�&:ǩE���r<C���>ð3�i03��I��Y�Vԧ
�սZue�!�	|�"qc�/�twr�R���	��J��l�I���@���,��件bԓk�z}�A�	_p��}�����O���;�~nn]V�����G�&{��L%�X�q |*&;)7T��Y,�5����.����!>s޵�H��NI���ASHUf���s^u��*u��E��(��`I�4~�n�b��ͫ�d��/ ��; ��N�ɂ��)��5{O�q�ר���	����C����d�	[[ܑ���
�����A�����6��(���c@�!�lJH4��,*����}2/�x����>٣���0}o�S�M�I\]h^	��7;B��M���d<�x[x��Y���Zs#	l��|��������_�"S1%}2-�M�����2�@��V	�����1X�2,��k5�G��w�� �B�������W��O�������c*�O���E���ؖ���p����$�������b]�`h�0�z���9ëD�|�=�O����=������?���`�^l��m�)GV{��9x1:�q��x�崺w��������?!�YF�4g���!�^���v�M����yx��1Y����3���:��h=9qׁ������.YB�r}���F)�"��:g	ܶ&����A���g��i����[��2�i3 �y�x�� ����F�La0�c���n��~�ٺQ����mH'��zҹ��li��x;De)l�d��0G��*�V ����_��dN�ϸ�-KX�~��4c�&���v��r�`w�cD�M��������t��I5??4�J�D���Kjf �+��o�is�VLtS�,T���`�5�%����.���
�M��ʬ�
���&h$Q���i[����M⊊+�Dѥ����W$��5���E1/>�v�[5�=��A�;�|oC
y��o�Q=2���N����2p����;��TǃȚp�g�6��p��nf�{�mg��B�q�YT��NW��|�p���tgܳpƾ��EcAIjn��f9XSh[IE�y\��]L�%�072SZ4|_��Q�{O�>���h�V��FtTEP��T�z��|Iҭ�u&��v�a�g#�R��v漋�G@�%��H?BYÛ�ҫM.�yF�'�$����*cV�����@9��:�2����ÆOL�Zn�� `A��i���H#'��"��^�^7���Q�ka�-�%��2t"���_�~�}�߽�͡��Eb0���&�抐�4 Bf�¾_��=F�-���[�D_�7${�+{�P�+h��
�����t[ ���xk��g ��<��ݖ�z	�)Dl��n�f�E�AjC!�1&]TF�g�!�1+/ƈdďC)�?I��u���Bp55�\�M��c���FO�!�]Y����6�{��OhE"�?�[�ґ�'f�P�K����T�F�2���\-�`1)/�()%�F�AE���AG��\0��N����z� nJ[	�h�m���	�``�0ܕ������*o!p˜12�܈V��VZGĘ΁�WF2����XF?XMX}�G�W���@�.$pM9���(H4q*�s�ػh�S1�uQ_ɼ?aǯ%>G�w�u�!�8�����b�ł&�KV�X3YV}�L�Ϻ�����zalE��=:+��]Pď)�w!kZG�e2���[{0t��`�qB�UK���̲~���p�Pw�hTF;��e���RB�D�i�跾@�Ê$ԅ¼��=��A]EC!�ٴ�C���t�A�`��4�}V�b���x�I�WF6�����?���|��l�n����o�O�Q��O��8� �:L_t-����Km�N�B��MY�eI߰7f-��hD��ߎ���(�(�A���2{�L�V���+�T�p�D���cg��!s�l�
����F0�p%�������|G7����p�%�by0x%�ϣ�[�R|�A�,`���Ë���0ra���l
�Bb���j�v�.K� H�gub�}{ʊ�|�M߇�,O�k�ov*�P�4�S��qm�Z�FMCp��S��$���m~#m�Gu�v�r( Z2��]��-{:²�9�I��@�jE㪮5��@g�]M���Q�p_�.�q���<�L�H�ŁϨj-�5��֭
z��<���I:cF�E���kN��O���{�KZ_�Pm1����󓲉Y\>=|�֥���dJ��l��N L�[�I�ށ�&_"�S���f`(�f�dUw�� hg�Bќ~�������UL������.τ8N�K�t�9+<N� �2~��y�gQ���9Ϧ�G;ͯ֚nC*M�%��Ej�@��%qو.\��o�}�'�b��9W;����O�[ӟg}���`�.w��x&f�GX���ş���.O�iۆI�į�]!~��}��� �+>��,aKx\v+?��JpWS
=��7j�z-�� �Pp���D�B^�N��[��l�u���͙DHe�4U�_k��iL��I:��z���%�p%K M��ż��sȅYJܾǶ~�ރQ0KRPW�V�sC�S��A��r�bБ�$� >c��l�T����)c��Đ�in҂!��v[ȳ�����V�50�� �2�8�G��sֵ4�ĐM�tA�N铩��*��ٰ��ت�9w�
���3��nO��H �� +�
�����\C������uͪ�<w���]���@\$��A�~����4�5�%4U��r�A���m؇f��1��J3�����Ҿ�nB�Ժm$�Ȇ��䮒zn\���!��8{�x3��}?�p�w�3@\e�#Z�|���vcw LWGd���Rc���{,%��L�����GyB���?���Ͽ���r~`�K7��İ���:.d�1em�$�D6V�?�Ԡq.J�p���^������U7�aPmw�#�hc�
�]�$ �Pq����W�nW����_Z�i�;�B�OB�{L2ٿ��8	"+atz_	����Y�:Kb�6�v\��C�����Ѩ4�Z<j#��a�f����t�c��D���K���}�8a��SD�xF�x�9&���"�5���yF�+qG�1@=��H`(@׮�D�M;�H��<?ƿ �H�|9�>,f���C��a�s*	�V���ql�Q{_i��v{6�S��'�ԇ���0�Va�Q��$�x���՘*��l3+�Z�k����3�����쇺��7Ox��9��jڗ�⋝���E�k/�E~3Q��^@�"� XC���ZX��=9��SP�gV"#R�<� ��"9㼽��,�+NM��\����t�)E��.�����{o#�.���|���&��Xbw�hy�u�P!a!��p$���&�K�{q2-�L������S�a�i�lA {qv4�y9j(���Ҹ��g��^��NO!� 4���ʮ��1���Ç� �w�m����l���1��������c%�ˉ�5[V��Y��AP���f��o��=��5����-���v�'.cx��\� �{�`���c��M
+�5�!6�rc��6!�<�nȠd���vo��9��|*��X��9��:�-4H��e9J��-���P�\VzŜ��"A���H��qy*(-���Sr&/&/�|h�rٝ&;W����׻�#9i�˞�3*�Mt�hfq�g���*�q�$���+p��h��u,d�밷���� �:y��m�1��ZO)���66�ݞN���|o�j�hO���dQ��#�hr
5��*X�r������+w���gU0$�W��-�֎�~Бhr[�t<��B���g�PE�e�ę�!�z`�0W�/�/h c#3��.4���*�=��ёM�	c�{���ڳ;#�z��Բ�Rށ"������S�)�XC��Z����ni`I����PM�QX���3f��c�կ�T��q��ҧ���'��To/��� Xl-|L_�ެ�`��CM������ǎ�3-���X�E�������?���ja��Y�O�n�V�)�}o��W0t4AL�9�1��iҠ�rY�焮۫���^�k#'�ᓺ:\}�Þ�2,�>�p�j���Td�n��Ϟ�I�Am�D�y�I��o������mW��ٞ�yX˷�V�L�%L�ΑO�6w|r#
k�jz;����.`�}\��ф��Ga8�=�r(�C�w�U&`�Z�/vhy�|���\��0kuA�'E�z.]�/�S
(���d��+����x#�y���fF�Ź�tG�Z�r.v����&���nq�5ܪ�0�|R���5�K�j�I*֡\]����<4R�/��b)o��75Z�CSӪ�qM��� \�Cٷ�6�K-ѻ�ju~@:G� �{�^�����7V���k��vp�K�f��Y�1D��F��pC��3��a,�����cDEp��1W
����}���*��P���8`��?�T*�؅���| c�;�:/�4Ks~6z~q]��u���X�V��?��=(jJ��n#���)r��юHE@���Mǒ�!�ŋ	W��/J�Ľ�����dN��J�O����b����C���Sr�Գ�T�I�����L>-��R�S�˛�u�]�oc�	�.3�-½�K�- ��Qs�҈,'� WVK9�.�ms~�	��">(��Zg��~��O���%��^s��NsjM+- ���=>����x�"pdt䗃\,3 Z<���G}7#I~���2Pd���!;ڶ�QX*��SU��{a\���� ��^��*���+.� l_�B�7�#1%z��c��Xiz��F�!M\5�W�����)��[�:pF3��(�����93�� ���	B�]��(���]#�v[�dͦ��{:���F�K�C�����L�B��R�_s&�v%�!��ml\c	��l�:�O��fH�DT�E�$�#X��{͢�S��4���S_�|�Y�]ý#O�Q��v<�����h6BQ[WY��?)P_�)&�J�/g�#��n�xӰ<��Q�1��؝,�@���Ê�dT��}�P4���)�I$�*�X݇_Т^~�,*T�e>1������̦RJ�7CG���a���ru�2t^��;�N'�J�fK�y_�[3�C�!uaC��p�
#�z�Mk�`5����jX���^62Y��rXw��mD�nV�=�-SW9��=
�u3��2=D�(�~�l8�F�Cs����	y��j�Z+ܫ̰s�Vk?΁�:lݵ�a��`��D�2P���GǓ&� ��1���U�c?���@�h�6����T������<���%�ؙ_v���{�?�W�jK�R�%5l��-]%R��$�����z�QN%gcZ��M/ڣ5d&��c#d�g�����|��SU�Xn9r�v�<�¤���_����":��^��E2�Lil�(�����h���'9m��\J�%[Px�b��R����������0^��t]��͹;�.��1w�g,��VNP�6Փ}m6p�z�4��'u�Y�i7G�.�$�k�'O�[��쏊*���ey>E��{�b���Lԝ�#ю;��L_�Q�𠍙cm�KRU�V>*x�)9��u,f)ö�y�ꐘ�aP��.��*��o��[)�Z����r�%%�F��&������d�K�5��@ d,����(��ר�^"6�j �=!���ڨ�Ӕ��u<E�׬�I��4��t�/h�����}6e)
��v�u	��|�\ˠh��������n��j�������*��
��������ۭs��x.����H4��GO��z|�#�Pn�HHƌ�%�u����l�N���21>.Yӄ_쮊7[�H�dS�� ���a`ڑU8H��0�F3<��U	-t'X"G�����=6:��]Ԃ��4% ��xJ��Bi�r�.^�@v]G�"���� |%^2$h�Ãy3����D��E2�*��ֽ�2���M��o��l,%\t��_�̟���̬mRtH譎zM�[��?����8
W��W�9��A����~�����/R7�A�އ�o��c��t ���PzG�_������3���9T�GM�����p����ih}����f���K�Z����<N:���=�4�J[GкH�ud����l�8�������l��(�S�֕=��g`8��By���&����
T����5�" Y�vG:t�3�ނtf�iy�M!�C+QߜЋ-�p,
�+�V��[���$��,ET��e����*����K�|6��X�c�>��F� 4.���T�����1`OZ�E�Ij������l�=�=q�ThxVe^s竹��p^�E:�,Ѥ���ά��f����c�U����Λ��>���Ǣ���%9)����W����~��ߦܰY(�u<�s��I����N�Bx"隚�Xxp��<uz?�/��&�ry��d<L��  R��}�ZCg�[|�u-E��w�2f/*�1ը��p�ӎ��yJ�H��f0"���е���Y6#�M�Φ�I�n0��T�B������|���-��цF�S�X�Ô�Ӄjn������4���",�U1�.J?a�H��H�$��ʚj��E�\^:ќ�wO�sO:�.D�Sh̾����Ը�ro���No�.��x
���˫�J"?�K7su�ݩ�A��n\�9'�@��6K"�a�-��[M�0XiX��������A�L`�]ϋ�t�AS�csA�S���fkMCA��j�C�s'�4� ���x���{?N��1����;}ٝ� ��k9o� �4�K�f	���
r�q���$��V�`s�hk���ՠ#c�����ㄧB�EP2���o��t�i}$p
0p��]��������WR�:}wHr�l�]�"�sEPF;��)��?ݏ�F��$�F�r sH�*��,P�P�=!��I���I�ܖ<��;W��
��H���Ve�ӓ�I�;�Ya��a�f�ޛi����K�>Me��r�	��N\I��7�I��=�GT}n�/�	����MD�R�D�1�K��c����b34 ����եt��.�tDd�_x�&;y�X�o`0�=s�~8��ꌒ�6��dG�Zt��&�`[I�PGӷ1�l�'�'�f�_�v�(�G���b
:OZVq�@	>����S�	]�:lVv�^����a'��tO�~j%����el�]�ȁNS�F%)���X����H�~a#bE wdm����M_�ɇ d��@�k�]铚��T^̮/�V�}���Ki�(L���R8%�(?�aRWak9��à. �rYӳ���*N����!a'����	�%��w�dQG)�Uf¶b]6
���Sk�(���C�}pC������ĖMbF�R5M�H���6��5bO�XaBj8��8��Ѳe�1������{dm@�
�B��Ev����o��|#ތ���f�T�i)�9�+e>��X.����"b㛜�p^1},m� ���X���D��Xqrz�En�ÓM���dwTŁ�ˌ��L��3���,M'�G��x�r�g�5���E�m�ݣ�p�g\��q�j��s*��&k���7�&���x����T���L�b�0��'õ���B��R��߅���<m���3^�宙��x)S��ĜfX5������&�.�<�=(�]���)Ō�Q%{L�ð�*�QD-���0��_)�`���?t@x_@�&�^7vj���GƝ�&\��ƞ�����r��R��)��I�Q}=�B-;��R�ś�����T5��,������XQ�#nx�>.����CO�PgC��B��{�Ue멜Jߢ�Ai/�1�l��}{ؽn���}����N7�Q�/A�H�w�V��HH<¸���0�,4�Y�$�hs���5����p�g^�F��N9=�<��;���*<%䯵����o� ��&G�MJ��J�j�ED�P@6�c��;.�s�(j���T��P�#��nXf��*����sr�g8��e�������M�U�h�N��{dz}���9�)�]���5gjݥ~����f����:��e�갶�8�c(f�GR�zLO�".��N�	x+�48�	Z�^.��>����K*�|{�m	b��U*��t����� � �3��V�Rٴ#��bLra[{�j�E-w?Kf�`��=U���a�r��n+l�Z^���M���Ig�+�D7�s{b�ҤNf<�H�fEЦ8��R i�-oD�\G��<�&�g��Q4 [�G|��G5X�L�Q.�K����b�}̂��"�@�ˀ��u�!r/0�9�w�bY�O�5¡"y�|�3�6�P��� �0�X����z�"��ۻ%l���i�x���@-�(@���+����sD�Q�G{)�#db��o�:��ݬ�1}T�Jl�������0p�
t���Ā�D&��(���|�Q�3%��bEr��ns>Gpj��zA�a�۔��<~��n����=g�����%��Q���#[}��Ci_���0� ub�X��g��!��3�@�S�v�;<�P��/ ��KF};0n_�p���D�����}��v�4�g���I���c�8�j�i�J���#ȯ��4&��aX@=ķ.#�F�%��y�^�ȊF����t�s���Q��u#jΚ	]Hb�
,�Jc+�5q���e&���?XH�{6h�Rn���L�W�$�@�߿�0�}�Qi�����S����
�ӳ�����^�y�ḌÆ{a�I��߄������s���*t���~�^H���G�ˮ����ϼ��D�O@dL+�~�n��Sǟ�i����r� �?�۞�f89<%΍iU�O�������7���Au�\���1.� �j#�.D�#�KtZI�D��C�y;.ä,�k� *�Zi�\�fGXx�c�1�V�*黹ʅ#EN�t�p+ϯ;涮��$�;#�h������0��( �v3�"]g��nE`p�=���L��5B �L�����};�&�� k��[}Xo���VƯ*��y�Z��dY�`���9�'E=aj�hLKǻ�A1���)`S�kL��ws2):t%�H�o�IGf�_���@�4*BE�0!>8'��4�(�dkh'$����i$謕0��nu�PǴR4�r�!���w����D�{��e���Ui����,�1ܙJj���'�Q�>�'Y���7���[n��+h�ߺ��A�0�tv�ʢZ���tQ��
='�="L��V�ғfH��T�������;=G���k�smO�g��l�l[JF)�y����@�;f�s0t���Q:>I�0t��lB�i%_���HC���Ld����J6.�r,.�e.����$�Sf��\#!�R�gضW�0	XJN=���K_�̔��7E��Scx�T'���:m�"7 ��شG��\2������B���^D�YS��İ=Q��7dL?�e~S�b�:0�������>�^b���� oP:^h�X��<�l�+�n����5}�7��yg ���}h���%�]�r62�a���F8��1Kӽ/���Z��v�mS����YT	̫ʮ�؀�R�0ڑ䝢q�j�E�|�v�8<bm�7Wl�C�Na��B���\�_�=�Pxtbs�5�E�x���fB���M��������j�)oC�j��YC���\>m�x�)딆�����&T�=$;P`�`�''��T�xĞ��
��N�v�nKb��ݱ��Q��{�������;��i^�%)�l�����F�_	�;��l�+����t:ޒ��k����$��1���q�
�I�m���C.�u�}(��h����_p��@Ȃ����BJ�ɂ�d=����/BP��������7#Y�����*��<�Q�d/��	�\>V���$:O��"�5��B׊^U1��ӊB]{�\�4f��i��-f�݌6��{�A���Yֳ,��jjd����_�]7~P'-�]�L�x�"f�A�k�����""�����{C��CJ���*��'+��?~������H�+��w�����S�~n�9	@���>y,*�9;��X�B����I?�	|E�I��<R�(�P��:!��a#����ʕ���xϩ����S�XI�I$E�R8��餯:��e	��~�4�a����H����6�?�Ӝ?|���\�K]�{�<�Q	e�َs�f�]�;��a#�P�Vj������;1J��J�ܐ�?��8/��Dz^c��2�S�,ۻ[�A��u��{a�/8�'A�%�gF�X�;�{��xDv����dh����������X+�%�X�=�9��>;^VK؂���9��!��)e�p4��2�&�/v�3G�z��ߛd�k/��M��W�7���ʎ������-@Z���S |2ЍƲI,gX�Ǧ��g�t�>��P���!b����h[妞�ݢgl$pqݧ�͕��NsNT�P4�h���:��(��qs+Ω���˶v䅥�(@�����V��eMŞi��&�&���(�^u���[�����i�0�����U�t
��κ7F��]K�@�������rOg[��ҭl�o1�&��A��,����u�nB��*���, YRy����iQ�;���PL(G�::-h]p��v�G�?�,i�&�G� hW�_�IS�q�Q6 ����o<�Jü\����2�b�է��
X	b����q�'U�X^L}�"�0�c�Sn�������|JT-�+Mzw�rQ? �����R�B�C��b3v��Em�Y`���Z���P�Z�f�8�I�]^@��O	;��͞� �-@}�4+���q ��٫i�L�F ﾙ�TByP ]��	��X�P���$<��?�{zclK�T��0C����Vey��o�M�=:�Nՙ���u�߫%j�� ����0��ӷ:8�ަD	~6R3	�����&m���7{�p񞧼�:��uyo�*���8��`��������1; ]�C�4��\׼{\�lN�c�_&[JYY����O!!��}��C�r$
nwb�g�IK�5������~�$�5'x�}�'b�b�kgf8�ix�8X���`��m^�\�"qyKE����L�AK� ��V�Zg�s %�A�E��]+��5/]eB��jI��fc��J�(�����a}���0c�7��)%!����g��}\�Cͣ���`�}�F̠���@���s�H��>_��,�p�\�;�~���ܸ?r�^���)�2��.�ą=}�b�f��U��Wr����s�ҟ��1׭��0懾�==U��	��0ׂ{��J��t�HaHq`��:頻m�f'B��k#�-�ĥ���Gc�������Nl���r���V��Y`F��F<loAS�҉CЧ$�DL��d���*�Y􂣔.JN)�ǁ.���Aj�������d����A��������x7't�#f���αG�g�2�忤gp�]Qek�1$��d6.�8-ͷ���Y�(:�^ֽ>J���VX��t,��t�&�6�B[M�?�������sqx���/� ��Q�t/�HI�^�_D��'�jc�dmr��]�R�vTcⒼ�&��kdW�3�0>��1}.�Ļ�;;m����u-��~�S��QN��U�t\2b�8dK���vĎF3��D�؟u8���<L���ɖ�/љ�t3�$�҇o%C�|ï!K%OG��ک��y�Ē疬���qYv^�g��þ���ň�M2 �M����z� 7�,�|L�����KK�͎��l�+��F��`[�մ~�����Ǌ�h�*��|`�O�Qm�d���zDi:wUɤE��1���6��2�)S:Qc���Vs����.�|n���>���3k�Y�~ykM�[�՜�?�`��Hu�z�����ϋ%��A��UH���3�;>�� ��"���H�K�縟HnT���O�mc;��ի묪g���4;��9J�3,�6I=���"F�f�-�=��H�9+�ƾ���AV��d�C�`[�"�ͤf&��`|��N�p��l�ܤ�%A�	��-��NN�n�L�_y��8��c_2�8��9���r���p���g�'���)�tK�4����ہ�_u9����7�m�����<^���^&p�JJ��`#YxC)R������I�Z��ِ����S� ���rm;�!�-�m���ұݱ玽��/-�\��_`����5�ydt���Ϋ?r���^���WpM�$A!�fp�&[��i�����*�@ : ����L]��o>��?��"g��r�ts���/��Y�#X0׈�z|	�Mv����1-JY���ޮ����eµd��h
<)�#��Ns��IB�l�N��e��DF�XN~����&z��q����t}�!�뻎Lc,�ʄE��|NYf�����R�L�A6��h���y��{7KI���ǡ�>��WLW�y�e%k����A2�jC.;TC�e�T�I3����Aܭeޑ=�����W"7=�DN��N�h��� Z�F `��3�]#1�ihG���-b]W!P����D���gI�[�H���A,.1R��
7���!��7]d��K��2��C�l�j���W�=�{+!��7������Tw����K�����K��o�u����T5
�g�^B�wYE�P[��\G-�yuM��K��QGf�K�ô����o��������3+&���^���<}"K�����R'�2fg�/)��fG�	H,�u�`�p�G�,ȴ���g�f��n��Mµ��7D=;�Ү�Y��5�R�4�y�4�g�ji(���ѓ���꿓�X���`a�iU�#�IJ���~�"ڥ�A����Q�N����F�_u0w�F��� u;QZ���UT
9��Ό�(�P��{Q�FnY��I�rf����9��>9;����yޮLU�e�Bm-$��%�>��a�5U�T]O���i����I�%�� 8Rz*?�&�l��H/dp��]�W���ݦ3���w�<ӂ)3|DclԒ��[zVς	Hxg׆���Go��sjY� �'�2�>͎ ^&
����RU�=�C�����Q���¹���!��@���|V��Vrn�|�,��evN�g�d�Tҕb��
N���eV1�k�ɑ/�����կK�}�AaU��p�"W��	�Rr2���.���Ds�?��d�B,�MsI�
#	�Ɛ�2�I��U�E��l
?��>�4p��H��ժs�X�L9կ�\�m�S�4�N=a�!�>��GC����%�n�K��j�)<�4��E284��jܯa(�HR�=
]�
YᲐ�������*z>`��1������ �-z|�T.���:_/a��O@9���Y6ǯ_~gl/�{v$�f�2HsP�v>FuEKc�p����ot:]	�WE�^c�HV(�L���+$II�?�p�[�C�O���F���贛�>{��,)�x Hk�^^�,rP�j=��b2M}Q�6I�]	EE~@腽��p�����15�
J�S�ͧү�����rdB��}��0E/!���θN����K�>�������)���4�v���L們.2o�����sq!aȊ'c��[	�0W��X��4 ���VK�`Q��Z!Q�g�.v�T�N��ã&=����'�2��@�
�|�}���ߩ��Y�k�g/���A:��.��oq�R(;�?z�?j���5wJ��^+��1}X���đJ��i1Bnj��"/��}y���:��S����'�wǏ�`W���� ~�g�D��4o�����L�5F�ۗ��QuLeD*����b�'�Ψx���;�j�p��i̋��b�ߓ�YVjp5����%C1D]I������9���=:r�����L�Qm�$ern��L6�cj��c�����n�̆ݚ+��y$�J�uc�,

��,��U��|����G}%���M��d��=n�D���zbH�E6�2�%��X�h}��8����	sw{N��}(�\u�K��kAECҶ���3��~-��LV�S�X~@���V�ғ5�)K��!�ì���n�l*�[N)2R�/0t���s�_�W�0
(3 ����Qz+��Ϯ�Յ ۚ_}2z�py���Ob��`f�R�"/���>�
T�Q�0I��)��j�:�m޾C��W�P)�<��K=�z����>c��sg���F¢�'�9���X"K)�D;�a��"VTO���3R����?`�R;Av��RH�m�����O)Nk��ʴ�{qB�D;GQV��9��.��$hđ��D_���+����dL�m'�HN�>Il�"�j��'���O���+2��$����!�zW�6�@ge����)���c��ظ[�y�j���u�PD�"ĵ�&��&��7*w�~�b���c���Y� k�� P���Eq����Զ����%(g����jF	Ke��u:$�v ��0u��X"���Z(G=��=���3�F= �UC� 0�������vR�d��n��8r��[Y8p�`(.�[<K+���]����I���Hu��5��^�qA����/#[���h++�8}�.��ۘ1p����#�	P;���m�Z(���Ə��,� �s<g�4��\Ӧ�1
a���R�)��n�����x#���`"������7�O�e~���h%9}��8qV����&���)C1�pf���c9��s�\J���C@-Ϗ��ګ���=�
�~F��S��h�5`�ڿ��n�w[{h��F/�Q���+�N��I˙�I�M�jV؇l(�{��,z;�!�,��:���9:3�P�9�	�m	��oz�#�?�����J��析��ҁH����q����+���O3�Ғk��G�K�lD���4f
�������W?�{�̏�6(߸� B������N1o�^��[N�C���貝�,=��*�*�Ѿi�˚L��A�4G�1]��\@������5�y�!6��'�͘Z6ݠ_��(CN��J�r�Qg�>Ѿ?஻�=%����j��@K���8��7�]�=��'E��6�MV��EC3lC\v8ez�r�騻��+��b,%��^�f�ŰZ%�k�l����=�YɊz�D� �$�,���,��͗��@(^�����[�q�諎w�	����ܚ����c3-���v�Ӹ�h;}�Ö�kƛ�:�By#�D���ۊК�
f!��Z�/д��7��C��)��i^M�uB��:y��K�ו/�gJ��[�t��颸lb�VZ,����O���<�v�{Mű���e
�P��
󰓔u�'�bX-0�RY��\1�	"�_���k��[x8��V��tʟG��w��*8z���Qt��^�0���u�,��`L�}�H�r��<T�[�꘺I�=%;������	�Ԙ��Z�W�\�ئ�^y�0��ϻ^�G��-�S��6��?�h�:�'C�L �R7~�M�ñQ�[Z�e�~գ�����*�~f�T'Nœm\w�k�G�Ch�6��:/Ғ����R�r���|�s��[Y@��G��b̿��M�}Mz࢛&V�ZSd��Z�y��c���m���#��	.�vb������V�T
l��g͂6���_�gfY�Oz����y�[]������i<�Yϕd��s{R��ߴ.���(�IE}/�#�y�h���c'ʲF���U�~~[�g�~��߬�� *j��@���^��?�7]��G�U�`�ϩӨ�9EƤ�p�3ͥ���i`h�;O���g>�w�j��yb�gV�%�t]If�
D��@,�_���kq���6F*�m�צ����c����3�!�17i�1�=����O����/������Q��*���Y�Ɗ���0a���;Yƪ��A�|6�x��<�!�eSk�O����k��dB��N#j�
X�+"����夘~�v*���{˳W��7��e>0>�Y�1�qWr�Υ*��S�Cݳ�Q�ʏ�ɃE�@�Ǥτs"J��+��+���Hzꗙ���t���~*�$%��qG�jUӒ	w�A��vMX%`d假�5�I��&<���r��$Fo��]�_Q(�\)� 2�AA6�У>E~<�^fo���>��s��E�rP��{��g�3���)x����!3�o	',��Ny��:,v�i*_�B��	��~X��$\��?��N(;p����yN� ZEN�ٲ�zu�BA��z��p
��/c��3b�]�8^�G��&c�u |���0p�Zi{���">���c|e�U�0yA�k�u��� ��A��5�҂��P~���]�]��ш���A��Y`�ҕL�����LVF��k�[�������??U�k�
/��ڙ�"�(	/��_��{�K�Ip/H����%��4�P��͹��f���	�+�Z�cnY�9R1ǋD1$W�/`�יi��f �Yc��qQأ=�E����{f��bq���1&��c�pab��o �b��=�-������n�6 f��$E�'�p��ե�GU!�b��>���j���=��� ���~X_�]hĬ�1äd�������7V��v��K�Bج/Lsu�P�"Vp�p��.�;�<]G��m�D.�2I �P��KTAs^nY���A�ӥ��t,�~&?$������y*�vaX�Z5t&�&��̵��I)^�0`:��4�%��R������-)Ji�ٍ�:ϭ�E���s��	��q����Ը��r��ßB���k#"-w����Ⱦο�>�����@�h
�R]qV\��=:���W�t�X)�5��{�ѐ@�(��:�f�π�������B�%�]�E��b@�v)�yb���)�#��
�%_� ��I}���s^�aT�)� �Pd	ڔؗy�O��%�yw��7�ӛ�d��^F�����#��{.K�+]��t c��ibW*�!-��է
�,A=K�û�2�D�v���~�@	����*�]�ͬ�&�E!,��&�� �#��y9�h��DGǶ�A�e���F-�M��Z�v�4�Ԯ����J����RIB��^е��}7y�Y��R�ϰzK,!�-�Ѯ��£7<K?�n�
gq��!B�UBHVg�M�'T(�U��o>��1<��a�J��C�r���6K5YA!N����D(8ɪE����m���ưƩa��vK`'P<��_�YV�33���Je�Np�I%��Ig}t�����YK6��$��EH�Wb򲤢�Q���Lk=�I<M���� p�Tt�hl;���'�isAtL��Q�k�%!�9uh>�2i˂,o�>�/��I�_�h��%�ͮ��1��;#��c��v7 Ƈ�G5�O�YR�rͺ�1b����9�M�
&G���@�%��}ľ�9م�TDb�\ �n� ���T'�*�oz�8Du�L��^
E	�����4���ù�?�m[%� ���E�o��'
�C�k�e��|�pO��A����K���k9]5���XA�=v�Q�i{�7^/��Dп9���"�����zd�T��i���(x���H!�<o���5yv"XR�\�jf h`=�s�hd��Uc4�0����H̝�"n��+���ۚ���z��i����J�u9F_vO�L�����i�I5Q�}N�L���Hq��@)qW��=��+}�P��-P4��c�7����%>�gkt�,�{.A�0����Gp��BRn�������i˫�¼�\<�c6%|eh�^4������w"��׸4V�|���Y��4��Q�6�jO��^H���Fb��n�F��1}-vt ـ��;�cb�����۳Ԝ]	�'kP�f,o�h�*��"�+sPưl������	5��y�b���<Ƚ��lX�n�r*�T&U�M��'nA�A��S�Im���9�`3��p�	��D�+hY��'�ʼ���й�:�p�V����NF}�DuH�*��o ,6���ʀ��H�h>��F��{�� �A|P,kH�����ؽ�
D�)�L����b��L��.�m���)�~�f>�� �w\@�#q�5�g���(��o7{�eGO��I��̌��֭�'u�]}�3��ؘ#�a�U��L�v��#2ex+9��z(hr��M��\�����\��IQ�-�%=~2�"B\W)7C�������Z��vU�\�m���V�	6���[�>�V=yV�^�>O���T������3]���?]��4��@���)�DS����o��{d�p��x���%��B!�NZ��}5�[��x4Ձ
 ��/�+��_�ǧtNw��x��Ʈ��ͮ�Y"�xX��X�z�8l����alcǉ,q8�w�#@��V�y�y����i���Zw��S�먱3M��DV�B�����I"ԡE�`�Js!�v��V@�:\=�o�r��F��nR6�ɰ�r���Y�M��d�I�/��|wT�V2쑝2�Ѭ�?�ۍ:8L�u�b�����{yn��'[�l�˺�����ew��5E[(��,z8�/�Z0�~�q����Ǯ0�6��Y�
�k#<c�E ������c���K�-(5�;^"3�w&l�6�F�����'������x�\%L�n�X�1�$?5-�{C����`$���ٰc�叢�`��=�PV۬C+rw���z[��o�٤���ń�S�:N֍�E��?*]����?VT��W��V�To��y?�(�{�{XL��@��}A�;yz��F��Q,�-c�"#��W;��֝eW�*g�Iw��Jm4G>Jۛŗ�F:R~p	�&�O����u!3�YPL�$�>���nג&�~�/v�*��٦E���r��Sn�X�d^�eӇ����ѽ�y������2��?�W	[ݤ��Qb$���xI��\^�C���}�
J
����Y��l�Ν�'4?�{j����N;�.��S�|@3��ǹ�3��g���sڻ�lw!����# ̑���vnJ��FA�����Q:_��8h��"?K�7A�@�)�$�<F�7Nl$����oG0X���l�_e�����'���$Ï`6�_�{|�$�kAҭ��ӉA�S�P}���I\��Z�E�=��C4�ċ���4?Mq1ۄhW�q�f�G��t^�Y�C`����u�-���ڨ�{��և���'?&�����~eRBs��[�[��S�����"�*L����F����Z�ӕ>�yYTR��^�~���%s�����r���Y@�쓻�͛�7<*����n���������I9��-�k���'&� ����m�3t����ܷ���as�ؒZ?�~gP�z#if9�N�-"=������6le��
���Ӻ"�:4�"j�g�j}����z�k2��8+١���(�%��I�l��
:e1�p�|D|Q�;a���[��I�(�����BC�Q�L3���B�,S0��4._����S35x�!��
�K�q������o5-Cp�9�ʇ��oh����FE��Bd��s\L��sp����D���Ԣ���,����9������rӦ*����	�j^�	R�9�jNu�b6�؃��#����������|Ux�Q������۞0���YQ!�8�]�9w�T�~�"*�1�zI�n�4�^���/C��ҍv&�2'HX���~�R�*�H�mr�n,���X.�_���'\wq�s����OB�z�	�MX����SǻX�nB(^=Y�Z|�&�}�l3�u~;~����E�;ȃw�CD��7�3(K#R�3�6�L%�0�@�<mg����?.�$7�^��W�ú��|>,�続��'���\Gl  558o�m1�u*J*��p�O���A��xkFɗ���f�L��0V����K�q!��2T&����� k��P`����Й߲8oq
�͐�fX�#x͠��=:���Bd?r93h�-/�7�C>%��!��� =`{�-�����(��$������_��D�6�_u{Ӎ�='n���%��3�9�Y2��ͳ㨥:/�!����1jX�3�h� cry�����u���R"s�q�֌�l԰�(���{�	�6��|�
��T{4C.���ۺ�!�_��,>��*,8�#jH��^��p�ϥG�ƙ���;� �o��6�5�O��a��Q㛻S�6�z-�Q$lW�\t�!ʚ�RPG��PPЉ��v�)kA�}eߏ8x��NЗ�c*A��N�)�й
�NRq�C��QO |3�9[C0��LМ��zK��Z�-����[!c~�	��a�@���HT9����3䕢�&�F]-��X�����s-eX�"Ӧ��V{�����Dj��f�EW�v��?y��'�4^�:W���,���}�����ȷY�)�����6�o4���G��������xY�т�cs@�gp��C)MN�X�䒰�|�'Ԭu�}`�T��ߵr��J��7�i ��5�|�l��	��b���V����F�%���U^�ء��H�d��5�6i:�����/�1�>�S�qJ|����3��A��C�}�������i4�^FZeA}Զ�V��#xWFr��7�^��>�}~ÿg7�t�6}��8����Ti�A��Ne�G'��t������ R����M��<�nsH��:���Tл���s��� K���}8����b�f�gXe��C� �ۅ�*�D2���P��ٿ����E�sԊ���r�)��&^�eRGo}?H�&� :䕦���`�2���Qn{ ��w����mrG��\湋����D�x��v	#3A�����Vl���4ۣB�Z�i�-8�%�CN��S�\-m���yC�K,=�y���v�ޖ��J�rj��� �����ICX���ݯ��N]j��J��[��蕣�U_<6 �Ӹ> �vJM~�x�Ë6�4�9|�"��8����;S"p�UQ��N6^6x6lX5�S��q�L^�܈7��ryX��^ ���M�����pC�D�[ʘ�qa��DZ+�1�:w�iVJ+����k�4���z~N���Ǟ��,>�WG�v�C� 5�w�!�����f�����oc�X���8���o�?;�^n���;��'͢S����cp��Q�� ���7���K�U"lS���&����6�p8ɛp���O��S,�ru��^�Fi�/�T����3��'�	є u	ƕT�:ʔ>�f��~>5;}����^5GGg�j���z�jG�����G�i�<�<�&+C@˶�U)v�s�s�c)Q����*�@Q<Q���H/άry����"�l@ݙ�<�f�La�a�}B��9�چ�&az14�hG6`	���.s�:��_�P[m�H.H8����eV q��]*�a�9�sź���R�/`�]7nK�*厦�甼���q4ٞЍ�=�ɚ1A�rI�73,4 ����G?l�7(^���`�3S�4�s�g#�����������g�k�v�)WV�ӿk��z����q��hyj�\�X����VΪĄVޯD��A�����'X[�JCM7����psUFgۜas�,I�%���%T%;���u"I�������C�֟������&y�d�����{�|B��i����iɾ@,� �c�L: �N�u�S� �Rz����ʓ�\N��N��a(8��I��q!�{Iƴ��׍��wy�5Uw���
�9�%�#������2��o�퀦�����
��0����R_��l{(ՙ�]���E����Ov)ȉ���҃��AW��)eT���A��ڃ��7�%Uett-�hh��	����M!��� �:G����|�����cA�XblFL�΅����{NY�9M�����Wt���Ȳn����������J��EX����o%�Y�"�9���dУ	|@K�ѯ��G��y3�G��B��ꃩ�f@?ƻs�s��M#o��������0��o���G�
��X���l&�bs�(
������]&w@�9�ź��K��`���p�f5�uB��;ϊ��&v���@�7��U�y�UN*�R���%�=�@��7��;md�IS5��G|�������8�cY(�Z�ڒ�{:��׽}iMD��I���Ѣ�v.zT��iM�n�B�5��U3����-��<��Du�����vtn���2���;����q#�@�}��W!Q� 1��$ɱ��_Һ����P������:/kn����ڎ�\�QH�����3��<�Ԏ��N��*�u������9�Ѭv�i�� ])If��EqП�'Z��{��Q;�roר꫗SP=vxq�/�$\�)���5���ŪLsRe���'RB��k�dm������b=���C�gz���%�P����MM΀ȥR��hk�% �n�g��?���b�[H rS��~���qA斝�E� 1M�1�������nv��ǁp�Qg<ٚ��?��p�;m���.%(��er���K����V&R�L��������pxS�Xio������Cm�,4��fZ=���yzM ����@w��S!0F�,DU(R�����EE+[�*�Pp�2����Ԩ�?c���܂�!�;i0��N;���x@D�H=k��{����̤�Np?D}�<$5�qߊ��/������Fӧ��v�ŭ"�(��;�j�P��@Ťm{mĠ�`� 6�D�^+���2�9{��	���\�ѻZGD���m�M����\&0���u������~����<��j۶э:* ��Ѹ��-4���S�$��n���}�VxYiW]M8-K 
YZ�v���w���ls�m��h;W�2h�1�u��!?���tw;�&m#��y�d���Ak��+��qK�'r��pEy-5�3�NE�e�if��ϗ��L�?c��a�W�T�R���1.Ͳ���͝�ԧ��OU�̙���-�w~����Y_� }���.ވP=�����+U���o��t�CG��uAr�u��A��DG(���[4D��0���GP��>����9�w�0���y7[��+��ys-&�f����	��?��0f1�����R�����{JkTD}�����ǡG���,~��Q��.mNO44�Z��UH ��࡛ޏ�F�۷s�|��r�C �V�+��,�o64_Q�
��s��i��|�H%z��ܜb�����a�_�ɯQagl��$t9��6�������B+��nJ��zX�]]NQ8��8�ND�U^��~�[��S�%�����Q�� �o�{XC�(>(2�/F�jʓmc/��	\}m�2aRh:I�gk���2��-�0����[�'9;�-�	"��E�J4�����QT�~@���� ��*{��[�$�v�����7[.tX/.SmtTk�E5!Y���E�������4KEW��[)��:��ˌ}x�Ø��i�aLoh��r��z#S��N�$���D�1� t?spЧ�ه�� �ϑ0�"@!D~~�Hq��'�+:���On�����,>��R8��������^I�L��yNK��}��-�ƾ����,��A*a3s�i���@��w�C�]����U0����At��Dĸ�{ب7��s:"�w����o��Q��(fg�%'�МbxX�BSGk���{�0��c\�K-�����g|o6�W��q�ܓ�;�^ ��C���v����Dz5R]���G혓?@�7��[�$�"7@���/y0����fL�Z�hQ�)2�łD�+z���Vܪk؟l�I^Y�w�ؒ�&��	R8���y�P	�c=b�*?���*�_�s�>���o!�<P�~��u4\�n/ɈM��/��&N�����6�Єˏi"�u`@DG]K�:�V�P�g&�A�=��[|���k���v��"p�M�G���;gt��S��∅���j�4�[��{om����f|�ro0�ms�1d�V���󽙵�Kt4��l�������i�%�̼{ŊTP�� ��V���/* G��V�h�4�mp��lԇ�.8�f��v L8�2��㳨�4c�n��6O ��� �t���)��X��i��rK�'���$&�6=i�* "z�y�6,�`C�Դx�Nv56�]���#m)W�w)��[�ftU[J�`���'vFf����rW�&5n�^27;/���.�}E!���$�B����6
��6<���I���%FW�`���:� �"Ӻ6���xƩC���1b�
��#��4�3H�%�S��U�ڮ�<�PSV����رpD�9|�b��^kD�Q��8���#9.VEw��&���ݚe���.�#�ݾ���~�b��