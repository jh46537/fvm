// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:44 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LP9AbNEUdwJANwnd/QaGqG1mlKPZI8GdIne7pEbod6GZeG2lFn5qegWWYs7Y1FJz
Ucf9AHMHxZS2m6CqfB9uCcMb17pDeGzbNw+bvbL8pbHZ2vGD2/Mzywv6n8QRqKmB
53EU/X4oEZSfRfNyRBKk7Cl3JQzMiwLegz+PYAzQ244=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6544)
Sl8w0LYEAFG5AysozzkHCHJLgt1SezQUsRoHdELIiK+Jz2YqNVVgaL6vm+z7KCrm
/fMDoB5VO3qz3Obpk9+K9xRpvwHT22lACdWC6B7hR6ZCQSN/QXJi9sZTFrinOdIv
cm4nxWnXq6TMb73sBisfnSHKwe1xjJaNMgXD04zeJi2gqPy08SO9ZvjHp4beMpfP
7qeIZC84x/ck90lCCfjHiny5ax8JdcsUONvpYSeCMuwhvRsXzbSMoTuCK7EOSGtw
7TI+bfsFBVokYZmojIidJ1mcoGsNqfEDzGoJ6MULl+sQ7mwV/y+J2OEJgTl7k9mV
n9Wyb/CAEKhNOyuNsb0k+AY/syflO+MuUraQFu9S81KysMPEU67Rfl77FnnFiygx
kYtBxdE5W0G3QpQst0uIUsBqyju9NR4ZTj63XBYh7WuABbMn2OyD8NlZHvpBQe6s
D0SwCbmMAkGyjOg2UBIPUmG0yuyLmKzzIKV764kRKNO7gwNKVizD6qXPo559l6Qa
P4Z0jxM//nJcOlgjcvGJRx7JDOM1eRhfXl9KmumPsmSMs+sFfFcZxv+LXgRbpj2a
uMjD1mvb7OZZ/9cV42wVLLcQXFhnQ2LuMQBOmIamDTSlqL6SoW0VuoqrIU+YhKB5
Ld58r0XdRXlMOmtenDY3iU8/47cj57ruofrxeWTKx6lCxMwlPGioPz2gHbsn4NBt
iCoNSP+Fo1eyhblxvQQZRasfYdSbFiSstRfb/Y6EooPhw8MH80bG6yRQ/u2l44BX
r2abFOHxabq5rHGI136Sbb0S0Z/VU7chua75V10Q296bKNqjR4n35e26z/+MryRJ
InxydUWxzBr3G1JAsXSX0GjMWqY5cBZ7bFN5kcPnKCboNaltNmMUbQAAtqx7m/rv
X8uzJbdtf5TNBmd9Fn+kJy9I8gL8sjGvtk4BPMMk8/7GK/JGWpLdYfl+VlG9futP
VWMmgG4xaOYGZjXLzMCnPsEfCXkE6l0rS23XAp2wEdiHaPFwdB/r2W/sREB70RT1
RHVvIbGdy9wYmWGs3Lnq+3hK/tnUrqAgh2lwdCIh2sGTYCW5YvbiaFkvyAw319wW
zBDmjGUBUZWenusPv0F9Ha/YwjhC8E07mOcThA/cgdXPfKNQGt2S1Z4FIROxCrDV
Ro3vdDwtSJ1/H9BH1g6zrqDBzEj1YlKhO34f30BNlzDVxmsr0ZW3ebB7di1v52Od
91NHMvaoZNzv/d21zAeOUt6f7KUzTmqtkq9s//t8zIR6lR5/JQOEitp4aewQmH7Q
GmWqzScoC9vwLOSYPo+oVvNGezmACa3ROSMLxFHf3OMo4f4wrywPQgq0a4kpaibW
sW8xTIO969AyaQCeGts5kKhYyqm7g0ack86p+dKD7YXkY/DoJcG0hCY8z05DZpsw
VsLWZvMZwmOBqeMFT/Z/tOLJVCH4rzDWHx0sLws4b+ua6lZ3cEVeFMbK9N2P3nLf
U5HRBNuJdoNH1D1Fcm69fuKyDrrCuyS9Lkdssp9x0fK+r15hz86ZLQTRBc6MyI/v
T5kun7dNrV70O0fPQXOntGWT0OsmS8JgQ5aVPo0eYo/J+BHELhL4oIuRAP29TI7+
ApSvTNyhjy8FFZd6xb4pViErsMbVJL4LL4HDKrWLDlzLvDB3AVMvWJ1XwpnJzc3R
/D9cUwszCEUowR73jc0pAqTNOl1Qt6lgojDZh1iDU6E/6NClwrVUlB1cQK0yBkLx
aRmM9RSe9wXK/JaVIk5TNrsJw0hIoVhGJFxU6VU6QEHr+nquaa2XW2VGITgcEyZy
F85Ees8PynfSYxXqdKcA8BvdmYCy78aTPXBTo+/TcmNiREJaLkON0lOxIPntK+/j
W+lQcdGElYjgnLjQibmc55g0IExbU4gk3yBf6r6z4UKhrlrcHa2ghwi5CcH7/wnF
A3GdHGucwmKC8DDykih1VPnuxwmaE9L4JutYfDdafdNfhT12GQz0EdR1vUf2WdcO
U/YZXOIV9z/8FajNO35jEl9ZMi4ngr70jY9A274NdBlYyQkL7d9qzOsBGZ0sjHLo
QE2oGNPthWX4gBo20NXSvJO7wDl20Er1r9m/rIJwzLWuNJd+3o3A+T+8/ZXzGcQp
+0Or+r76tZ6jRceOoUmkJZqcYn8MPMbDzEFIRdSxqlS3cvmpCA/OzCTDHT3VC95f
mgW3SdhDPkx6DwSpm3lYGODmxqnVuyc+gVUZJBPzpoW6zTzWEXc+6+RbBQFRAwT1
ahP8GjvZDjTkB2XuajkWXDSHlXoiHKfD+9BSVJpoNohtHw0TvkqOvYfV9Rs36zux
yrcUCVjaBKhcYlWU+KwQKYtC2OF2Gb/T+9aCxGlcNMMArwyKyOjvztDhmA5clxhw
4zb5wODS5D6wYp/2eJAF6gNltFrGhGsP8cqnf/xcXCVlmUJLK/AEiLD4j9Uks/L7
egvdP8f8bBOzp/qnCV5jR5I65Rex3oMRl/ze7qFoXJQcY7xlfUrIUY/3x1aqHL05
zlod2n6lHMYhXgh5Wmla+I/6zmvZl/lE8IEWbzEWFhXXzX4tFZ5BY7DheJEgeaAI
vBDsNHPoAQVnfvAVAccgHJtjFfCOHDTfbB+N1HbSrShTy+ExDf29dyP0US03SvEk
A8kJayjp6EYfZ8HoQ95pD7rnY2Gep/JIzLWfFbk3OHNkNwQq4HrUD8qd8YLzorVK
ZmMdpW9A1pKUMjjDpnRfwwXURP6RgCX/GHWwVT60RSKbT9UXdXPdu79eIUeweVcc
luEhE+PpBi1r26KwLv0zNL/csmk4FkLvxI92Jts9Q1xtu+7/SzT04M6ZZ3F41msM
UtpdX6XwoKkOJaR8Tg3O2X9xc3GfIkwWj1Y/DsbBVkEopFQ7LUXmrHWK9PVOVnZF
FT4lPUsg6Hgqo3MhVMA9v42XHUe7uGU1OHUIi+via/2353aTD81negPu+JM8TVJv
xBDZc6JjdSADIhpO5dh4q+0Y5GJgoIAnRPnnsb5Zj9qN3RgMW2Vrz4FNAD3EnfeK
txW9QAo7lO/wILQQv3OCOYXX/CPmd6PnhjdpJMlqMx55IWKaYtTVq0rP89zX/de4
+B93+OCkDLLr8Dky1uidgnU83dvAS6WHZvE8l11dqPij3lzUtesSh9uQ0XuuezM9
E/MYDoJDXnEtaCoP1sosEIyUOFyyEguGYqCjGdRfPX7X2JdFn2mA0fmyp/XaEKXR
gyae+yS2kSdorJKlAY8fODcNkRgYl3boltL3xNZrwLDBraO57/lwp9qXPKSvx0iM
EVI1FNIrTIQOE5aW35SRFpnpwc/LupbN2bBvD8DBOe49+lusFzjr/E9d7/NZaUKh
6t4GgZSLaVFDenfOlE6ZKCMONLYjF7FWhVkffGkmlqlRu1m8mJ2okP2WJFvUn4YN
4ZEM9dv/Mp464nmCLNNSHitaI/34bEazmCBMcjlWYSF3rejVhEimUPT5aBofuUDU
0k+CPnhv7y+7ZOIAOcPoJzE22V6ph8jJIqOpyObpE9JmmMPm7b2wIcjkUR6Gs8VO
nZyl864YCTYXrtpKDckUjH6wZ9/ncXn208SMReWaah4xnVoPUSy0iYTVhUVP/9gO
S8282SdZ5bEhs2tMBWuEosG4uvFlZCI1Hm6AqmyfbR+4nsBwh1kYVuHXNT9s5tyR
D2vCeXijAa5iScOA8ulU0+Zo8dT0/Hzqy+YnrZhA9v83qWGF1lL5uaa3xf+g4LRb
uzFe6n5pm3FcWx4yXVU++u0ucRDZi2ZjxABmDyuQJTG3bJa+hTBArGAi7aeIp2t6
CMfI9rNv6PC6kmJwSx9Dp+PrToOW9iFpXAWiZa2FTHF/wLqPTKaiF8q+8Oxy/ZZt
GWt3E+GyerkBCoJ547A9FjH3HqgFN48ZcYoWmMX/iO24i0mtdcp3eEq/56qptPY+
0gu9nJ42qf5MR+XMqJREqxbhYxzL+hHBIbP72D1RiBQObjlTgtZEie7Epv3kyfof
8TTBVvh6BlUTYd1mL8GYOFHyr0AmsG2KYn6qZycRIPORgVs2FDIqPMdJmun3EpVx
LgJ9xrTi5fnr8KbmK7wKFGw6f6L9a+oAuT07qsxyaUdBFO3r5XtblKDpNsgzjO3H
SgxAP+LNasmJqnGl2eEa/oyXygpv9yA1ozP4QrOhIZDcIJbO5ZLa19r0tkCFaWNi
YEcTl2c7Nm8bNxGNadQIWdBPDvlybjiROrr6pxkrV38miwgSucIJLvVtTz/trX74
6vk4Dqd7d8o2nD+2e5hAOesRKc60GEz0iV19CCKPN6YXNs795QCxVjxojikIVHjR
VlnU+4YQqsdRr4eA+c0vq7de66tsiF/r0Tjrn2DVFntN16g22yAhpQq4/5esBGeJ
lM8/1WNObeVY9/WOAiU65n6LKL0ymLKvtQyaZD5ypy+npDJLxp93c1IJIu0L2YVf
qBXQnuQtZybJMdQOA4uTwioAzMr/rZn0tWqbdoalBUFbTxYLL/XQx2RJ3Z+iHKIU
upfGSBvHbPo1W/1DTizjOnmxKHf9mNm0doTrKv/1E6wMxODwbTUWeu5XXs+o9CtY
PrkpPw6mRqNG8wskJofM4A9uxIoA2myemd03IfHsFwZuxlCt6y9s3Ts3YTwaxx4y
3564R2ydxWEfQ2F0IA5LBtUBCBwfVojaRNI6PACFlZIfANAEbsDCUgSClBC159By
viq1ZURhHbfbO3CCa1EHuJF7nBuHW7FJjLB/4E/LVokLZgwrZuawSQOriH2DDyoV
0+A4wnImcwHyu+9Pdkrtyh0LRLFA6hK4JgXcleONehu3il8KEKXJzPvXDV4OIMTd
BZV4Krlaef/UjFOdsOtNWrhB12c3H/eeTnLbtdV/8PYSL1r0SX1OAhUfk6DJYjgK
hfkBuUYg1ynEMAyJIbZuz3LKKXWErMpaoYMLV9NtjFw7SbZFtq8Nv2iuFE+e8R9U
I8Y7o7q54Ak5ZlTdGq2My77hsk2rkxXgJXQ5QJZ9WP3getiXF5MaCvtgybs9ndFw
NMFFZOvQZYMsI2MfveBZWe+tAnyzZ/l5iBhRZZoQKEssbDiXB+oHJCughP2pf0Gn
qKz0gVwqUfQvxT4jBZ+d5HxPi57xvZC1lJmCJlRzjrYGunWCUrdwIqAfmQRswl0G
Cpc33wM5PMGte3mWTVPH4FrT7WmHdnO4J4Rr/LN1ojFvfiApsE8+XpaH2gofQUeK
STqVp4QpxvfvXO4rq4PFGl9li6weeNAY9zNoJ9jxkmEv99DHrYnQDq6jAZs2A8p3
Uz4P51Tkyuj4g5EtWDkzVmC414HzASGfMLd9OCUUGNe31ysRIu+ibmxLhOERsCks
LIdB/BLWB3kJaciR7SV4ECPb/pRDLvND0C/id2vPSPPo8qVA5MIQPJOxF8b7i5Mx
TDGMphthbllGSBCCwElksOXcw3ztKFmailvkIQDXa7ELffyvd55eEUQanjEpKqNX
J0ThoTk2vicgE1RBOwItJyZOWr2xD2poaXSXGW2adqDOjcZDXLIMyS7cALX5jDMU
2E+0QBt38AcAyZ65ggCsc5v0bGTtZSNpqvw/P5H9nvAHUIyZ762d2Hb95cQHuryW
T5+HFmUgI5M2P84tib1nKlQfDWny0zTQBSrOMxjY/LT0G5bOH3cFdlOJMByVq4FU
+vQxrMOMn2OI2+2BiJtA7cNc0TvAckxLYGS1CSnA+jqrNZ6xIcNtjRLLJcacUaZM
pDZMJSSI+o7frnKPoeCme55ioRP4JkZmMb4L4wMqDYRUu+yGit1FQxkCNIUviXQZ
d0M3I7Kyu/XxhE7CEJGZ8EjwWbAsXtC9seh1m9nYGQZVcOw9VPmrgMDoVZWwynJ1
+o18oMBs/mWF1cSYoxxqRlvdoRgFNfR7LaYx+gHOgExdBJYRG+kGqs/tPSZzlgOf
NXtYvP51YkLPiYx8NohHDciPoya+nG5aEVRLqQdrWHp1D726kDf9rXPJf5iUq0QL
5XR2PEkp5blsVhww66UAeMFVVHQWBMUVUJfqCLA2b5mQyVCCv02qRH0EAdjjNgZ7
VgzEaRokycqK5eF6uT3h1gFexjgLUrhqURiCcVnSBMBEkubrilRnO8KPWj+u7irq
7Ob2reHblRT9Z8UlEaVgx715U1R7v62Sf4q4Y3w3yfcP8nsHn0dsj0tDJOEX2vN8
dka+NSceMJ/BU1N/IaRtkVRPcCrinIeQiMhSbh48D1qutKvRrgXK59oJUt5SdqLf
Szt0pbY5c29t2pMD/cIMzV2DVLueSn2NRzt0A7aaFa5tGxsPcgr0XR9E6WKYGBlO
C12jgbjPigusk+TlQZfwgHuX/Guv9cXVW9T7BAQcM2dt6X4H1h+AtAA5AGBdxuO2
wS+O+6B7ABJ87sJnjSFEoD4AF8ZxxWWyWE2tKPdPy4UQ5p+wEhS+rJyYGcNUWehv
ZFEAszbyXxig7Uy1fLubEUhbR1XTaqqiNpZNgX1HlAYrBpE+v9vxOu1IPAFQk0ND
gdsa1TZeDYCPsWuDirCPQUMTYXMnmQk7t2LgAL/2hM+doL8yFxrEv/lxTG3l2uSh
yZcxa2LDpFLWck4OssMxMqlOOt8vH9U8t7+sJlKoPrKCrMVL73vZgo88tMCi65f8
zumqub9J24qV8ZGk81swBxo3s9pPChdzZkiqalA19+Y5tazOALewtvcUC/fQQOMd
g2GQxeJsxvvaQvYXTm1aqXnddAkLtd/qqvZi/TEwJwQ7xBslogxwNIgnDx7j1KZG
Mpp194YmT67blRT1otT6QBXUV8j5DxatbhIwNPdVA3blqARsXtldK/NBmnrhnhqq
qHad8KDuAQzqjZub1UE5SPQCd9c6j3zUes0Awd/qTByPf+Ri88tgQ0pJD2rhKUIB
9oE5cfFWxC4qJsRZAeGKI7oPwG3u5xwJ0DPFbvUZtsq0azLdDLDSUHTnYr3eYZsU
ouys4afAImJRZRG7GZUaED8RgRTQWk4R6otYmiJeUsUxKUUcVfHajkCvkz6RpBG6
MNukIJUYUZnzBXUzVMXpXruHh/IyigZu2s+Exo/au9sq3o0XBVsEzZ9BunYPv+/X
CuAtYbwNcAzlIdWhN5++2elBqrR6Xzthwfsoo9lGGOvZjxF+PJXibH3Sw6g4aIPm
tasMVz87z2g8a7diIdtqrgBCzuN1mShhV0vR4wLgcpxJTA+H55kMqmeifBxfws2G
6phFb+fo+yxQsCYLlHlj7ehLKfnM+6j9kJUZ/GvIRyPFThp8EZ2GyAuwYJCzpaFl
AH9Wzd6fsOpefw1dCqVrNINjlEKa9d01H7i7TKBpVGcATUeLBFW+LQKFf9p8Y9aX
hYGuouVmfXNHiFDghyl4uk5l/3upWzxFvae3/iXa7R+9q2oMgnaxM84ygf5ASi3C
/NEmrsLxvRh3dpcAWWPPR674xpK0bFW1/9c12gRZuCzikKZIiE+9YSvr6eyRjZfq
c3fXoZx+ZGcRwSXNoXLMrEpBLL5LikfWKk108TxcEMDp+5JfBXgZn3u1y5MjbcgU
6/wZJ8IQI2ISkgjNA/0biLUuvX/cwbrJIUxqRmusZVwfuQkpkoE1+0w9ByGf6kjo
I8PDRqgYskAfc7OuZqI9VGG+Ftb+YX7XWPXz4wN7yLNb+nBMytXELlkbMgyfrANw
UwJ/tJdFHu5Ehkqy9KDdco4e0m3egQvv8YdvYGNYatER4GORYzr8mNNpUt73ItWL
j6GiP0SavHFL8hQ3PPjcv/WvRq7LwDema/riljFnarHNQFzUha2XZ9MqwWzEeHOS
5o8an7fT/vO5i+Ho5dpoH1x1FTT2CyM8xb8ogeSmQ5fCOpggYufv97ysxk/opP+G
wGpY8jgzENjQuOx/tHn8x72OLupuemlHv8lHc0llA3mhWHfCOMy8iNNK6ibr3A4k
aGnIPEcfc254EB5UIurm+FQmfjHKRR/CNrjfO/8DW9RCNVbgq67RZWd0YDNmpfFi
yiTd3//71RxAfpEK9XDQKJ/zULvuS+4KstYWcoLknQ6COiEMkZYlXwgYGm33B757
VSpm1FnBc0fr62hIdAnNBajN+AS40RMVXlt9xgrV8rsaq/p+1NqB7nwsKNC2hCou
mRVMKRnmt3ChscllZQbaxkpu4ZYqJJQZr8tu3EchmcWB9yVUb0V4bVlLC/iFa6+w
QtupvvENq4t5g2keXjNb5tYJ3FhQQK5zXfpYSaC9NuoEaqmVho8a+ZP3211e5nlE
knJ7VAgH68qEZ0+7bhonoDFc5V3EBkDrP/qDCJUv2g1Auk9QVu3sxMXLp07924oi
RPjT93AL07575DBH21+gwpZXe5OVVBaUjt7OKyN93utFWxipTNcIvHywKm7bIrHT
KxZBfQw0nN96Lf/la9OCugOorjk1aLokkBUQZReTbiLkmedthaZD5iB14YZ4R+rr
YdjjqBxdRYangxa/3BZI0bfbBKUE6BEmpRljZo8bueCYnr0ayH0yOig+0KkTwfn4
1giJFWc9v9EoH0YkVx7Dc6+SzDK5uXwrjtX1GvvMFNsWzLh7G/jQ5lTB7x4QbjST
YGangIbyKsqOk/aezFTsRlcfwjXSKGBuEMsCycGWKO+ihLj6ZSz9bNukV44+j25l
ftfBFHeRLTHJi+TjfRZ8uTPFOm1nT+KTyP5nrI/g8jBidbInOt61GBtB/N3iCkcf
B8SYuqzqgq92N9+ZfJAxkroz+I+wTRql+tljlJwR2Py1Cc0qBdJdBmF9qNCQkFhe
nXdd0EbtX8Eqx3cc6jy1Rw==
`pragma protect end_protected
