��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�_PN�2��,H_|O}��$7m�c��`�W�mZ��H���wz'�K�s<{(�*���w�%�:%�o��<+2?�=�l���L�G�n�y	�f��c]��g��77�D|��W�םfʠ�� q4���z��ص�n<S0z)��� ��]|������&(J��� #�eۑ��Nox��c6�)�瑹)Y�����sTt��p��T�j��凞s���<F��s�4����:.��� f Z*��R��?m�%�����Uf�ek�6��g���-���Ny4
�Z���l#ꄞ���-�Df�d�%��|��i�C��ٹ��o#��b�� ar���c"�Fۃ�l�9���6ތ��[�҆g����A�O4Q����hT�W1f��:
�z\n�s�Fz�#E:�9,���D������q���0h���z�E	{D�L�3�����ʩ@ q���I7¯���0O8��u�%0(7��f��i<����g��yʲ.�H��~T�/���H�g�؟�������o��#���Td,��P�ןEYH�q��<d� ����%�F=a����X4"
)QA-d�JO������A�����ִ�`���H��|��1�|��j���a�+M��#o�`��d��g��1����q��&^<�쑭w����ƫ�"swa"�� �3�É��\�$.��H�l���94���s�a0�%���_0@هp)I׻p�!�ꝗ�p�c�I���3]�U!�T����J�O�	)��Γ�y:h]�'�x�8�{{��иC"6���unD���L*B~���Lf_j��9����Qn��!��_X�����1�4|�w��Z��Ï��i^%anQ�@Є��.�{�I�k Ѐ�2u�Zēr�����֚0�s8IPfrf�y	��)�҈��X�����o�_Y�������3�G�T��.j�l�ό�+������w�lk�̈́�%�|�_��Ty�洭;��e�V^G*����V;����-����x)�:?RE���׀�A��34���HA�de}���!1=�e�ߵxq�2�+�JyW*#��6ZD�R(�]���'`x!�aY�X��C!v�cw��Lܛ�֬��1a��fљG��1.�r�A!��*����y��5��;�f�/[TВ󆅢�W�_�,\ס+bC�i�p=W�����G��)��0�T��??��'��fV����LC�m�6{s�x^������^nԫW���.]JJP�+#4����u_T&�b��9P�\,�k���l��^�Z�>��F�T���sF�FҠg����boh�4�)f"K���D&#�	y7:�6�Z9����|�.����^�����NQ����S�9�����Tb�!A������D0���X�J�
r{�-ek��A�X)��v�����h����E�-���ȗ�U�Z�x�3�}�X됍mN�ű��a6cJ=_��d�>Nk��N��B~�Y�+ܬ�b1<
#� t�2$�����e�k|B�m��^%/EL��҃�'T���!�RU-	���h�� 7�����{\	YJ�w��i2�&;�i2�b�h�vJp���	�Cx��&{G`�]V���s�CQ�ޢ)Q%��Y��8�xx�bo�c�18Nu9�$���5g��e����A��^�tb�zc�sR\�c�6_�ױ|~wY�b=� �nTi�g�/�J�O*��b�Ъg~J9�%�7��yC?�;�$���߀����Z��"l���W�yC����E�<����_
��ѡ�)9�-�}E
H��bl�?�m�V>���{�y
ei��Ca �ӖfgЩ�����қ?�����(�P��NBΛ3��@O:N��n����!�W����4���4�z�r�zITL�K�����6�8�|M@xKD�Mݢ�[��6�I��F�G�ҹ�`6й%��<X;�A�1����6��r�~��@���⇘;c|v�3�m��$�R�C��m��zam�����B���󓚉�W+h��^]r�:�m4Y�o�7��n.�t�
�Lk$?#�P����Н�^F ��.qY�ƅ����Q"�r�]�?�oߙ������i;��+���� �Иcr�n��E�5���U�72Cuz;�7/!���nP�����0�w�a��Q4yRK��j�W�o+^[��Vp�#�Uf�>��z`W��*������ߋ�G��J���1
�{7`'=�[�y*�y4����(a��G5$t�*��g������A�����7����^6�;��P²Szϧ3r��(��� ��gw�]��?8R߾0w�S�'?�Q��kIBj�2-+WX�^�uZ��7���Q��P2}A�,��y^Z-���vec�UR��I�@��-���z�R�0��8�tH��ӛLR�J&শ§NUq�հ��tR�tu{"�(�[X�])9=k��O8�p�rѬ��Ҥƨv@?+:�6�"�����=��K�ͪc_�R��_�`�9U�Z�J�P��ۇ˭A~�(�, @F��T�@�/�ÑBC�<��e 1j95/�0F=�cө-MH����ޥ2s�;e��?��["���y%��U����jac�$���N˾����(4ce�zkl�����(-ٸ�� m*�$��|������s�"�f�9�L5�6���7�t���7`f�{�rL�#�O�,zq�������"�%+I��bo(�_⨲e_��Ō~fq#<��I�a4�9T<�6�[G~	BZlX+�	���"W
��"t�u|�7D���nr�ie�|�ݟ��5ko�@-�+n����?PG�{����q��K���qF�-W�����I�%,�{ 6E).#���8�c%��H��5�j���c��݋��%��2{Cp��t��N�p�=�����W:�f�x���ކ��#�5yKx���bĤA�"����ŀ�;�
�䱸˷�/�|��y����4��1��N�����?@��I�:�"�Ψ���.̊�ʓ	e>XJ��A���wҪ�,n�h����D�0�${�[e�
۞�z<73[*�7�<37�y*�(#�DT��DK%&��16�
�d�7`C��[���U��ڋ娤u��hV&)"]�������wh�U��K�JB��4S
'�8�a�l�)��4�7��4����`wuMδkq��1J�����8�z�i�TR��ve����d1U��3�S�G�OzO�ͫ�W/4�(�N�˧�9����Ȧ��@��A�q:kp�&�lW���}�@�����
F�Q��%~�]�S2E~�6��B�������̥�fݼA�t�}�^���X�d��۹�>�b 1.tM9G�����;$ۤ�ͺ�E�� B����׀m�#�^�%	�����~�e!�h��Z�4��ڄm_e!G@[������gr�Rd�|�s�|ٞB�=PS%�(k�{y�2���-<EE�/.	�-�<���n�UW=ש�*}�"�Nq�ؾ#�lU+�4%��"���2�Ēl�f*є�.���4� �<�[�/��Z��J���gr롩/��7lL�y����ۜ�;Kd]��e#�%`̥H�(�\ڽRI#=F]JI��E��`�KoN Ή>GV�l�ƻ�f����}NQ��l�H��A�z�x��b��?���7S؆��u�(�g�8�Dl�\��sdV*�İ�b�`�c�+M�) ��3 �8�H�7�gE{�n�z$>}�cf�|���y	k���N)R�bYy� Q��Ru��GǄiox@v71<"j#BP0Ʌ�1Ś�I������n���R�!��6�H���a��x]�]['�f;i�_�Ҋ@���}��$&���ۼD����Zh1�k��?��	-b��([�� ���pA�\	��8M$v�u�)9$���)�/Kќ�G@1%f�=e�cE dls+Ow��,��g��0m��v�y�d��"X(I.y�5'�4�]��~�b�
+��f��4�k�8� ����/��T���${R ���H��8�L�����t!)�"5���ߪ����k���f@�ʓ�1��8΅ l��s��x�g@)y��I)��79�0:���"Âl�r�{�9u"��~�2�G��:w��@/�PwW�E��^�`�xi2£r��N�q��,`�J��y���Y�9�xoϻ)��W��^��p��L^����wFV]����3�!7��݂a���d�
h
[0ZQ��$��sZc^"�v�wt��0�:O��C�R@���~X濺3������%���%��;&D5�����NZ'�X'�ZI� ��"s��'W��9�A�����7�RRN)$�{��)����[�_�d�*`��9~A��(�{az��<�fO>ڐ�qO y����	-���?�d̳4�B�H�.P*WB�ݢ�qZ�#�r���q.75� �П�gܽSx3�#�(�u%���$�3)���Ƈ5"�wqWU�/n�R��+�����J��)�gI����E��^"2*��
�e�CVy��4*2���٘�͂�/�ώ�	�9���W���*}R��]g�B�0���tC�������k����������Y
x�P� A��4{@�x�w��M��E��P-��@�U��vRrՔ�[T�D5s�o���5��9�N�L�K��ً�x��ܔ��4�LB�̮yI!�$@��j�;�uH�tDm���VzR���D�� ��c��S���y.����]�G�!�S2~^;dGV����Vk�_�k_HwO0��tv�Xy���yV�$C��N8��JƵ�k�u�ˍ�[与���h��ՒuSnhD�y�)bg�y��7(��? 'j�Y�b��o�J��d�[�N�o>��=Ɖ�0�N�۷�s�v�z��R{A��[8]V`]�%t�nC�^m�7������� �%�o����@�T�r��
~6�T&'4#tF�e_H3�Ν.�g?���pB�y0�ot�G��Čx|'���j~g�8�X!3XL�$?v;�'�9l&�6*�T&;i2��W2�y�ۅ9"�"bּn�%��P&&�Gr��K	�ek��KZ�|w�>��|� ����mDV-"zË���������J���8�2aF���nh��$E����e�\��p��![e�,n�K9	�,��1ylC},&gS�w�vQb���;#�(7]��Z1�.udX���P`/A@=��N�Hm����M�Y���	%��_8�?�0���?%��k� �uϫ$����ǘU��"�	�Ę��q�{��u9Q�l�-��޼v�s�H]��N�B@VMq?�.*9sJ�X����ۊ��0�t�Y/3�wfql�4��1QB>�P 
�Ph�SgP�i�ђ���b�Į�����q��wlE�E|�W��`�)��(b�K"��źsܩeH.�Ze{�l�
�	:Gr�mŏ������@�N�kU���
���2��\��*7@Э�#mw�<��r����&%�a��{5��H�i�B<h�5�Y.Ʈ�~b�@	�[�Ft���q�zR�;�4�/��3�(p��q}L�|`��x�*�7=��@��. ��Ʈ�T�/��Li�-
��V��];b࿦�6���[M�4C��ē��PG�	6$�r
Jvj<���
��!=�N�����)���#)�/+�*�G�f&3&ݿ�-���3u���n���;Z��&`�O�}�rN��j���*3����a$�/}��-�+�B	K6k�gMQ8f�b_X�<���u���,A&��h���s�������ѝZWD� �f��f1��j(�,-���Zϔ��  ��|���}�sKg���ZX��
�6�V���b��'��gѤ4�!@�I�x����~�Va�F�a%�azt4��%�a���ְ�)��=9uϠ�zSr^�_r�lӶ��2�.M��C9,[�kћ3�;���u�|�rN�;�Zˡ�}i��W�d������g�mG�ZGF�qm*�����_>ϥ��x�
j��8W4m����t�;n)��4���N�Q�T��E���G���SWhϑ��}dXpB?��Y�_�hBB��	���y��7�ޢG�g5(U���9��SN�������#H�a��}��ۛ�_�|�~&jw�M��c>�rv��a���I��o�Y��DbPFn��(v2�vCQ-v�<��TS�%%z�ԉ���w��Y5����8��ᩣ\�jw(_��P��E�c���9�U����	�%H��3�#��no�$����~��+V�\����uH��2�3/�˝�GȾ�����wm�Q���|���(��JA)��G�U�N;�{��W��e��,C���ƞ���'ڸOǽ<8�X�~*�1ä�����c�)�YWAV��1�lӢ]cPe`5��$�Wi_v��;��w�E��GY^��w��C�	El�T4��Ѹ��~�xh���1�LZ���?���o4������B^'<ND�����n��yC#����dѧ��Ȓ������̃��/t�9a�<tr}Ι��T��A�ӏ@G��$�]�P�5���2eXa��E���y6�B�mo�ܶ�x�,?���-�5&@@v��,��+�u�-[�	|u�g�"��S̱S�a�D��  �a������-\a]�T.������� ��Wj�	?�7���%�r�>����\$y�� )��"m2���n�;Ĉ��ZK�~<�:@8����*�T����x������xd���
���:�wUZ�	w� ]���؁T3��!����}�o:��ma�qT�BV�,[��eaf'����d��^C?x04��R@JBz8�����x�Bh}�QS_�t+��n5��?���^H�vZm��9�A���|�Ý9*S#�'ݛ��KG3�ٟ�6U��q�I/[R����Hxc�cG]}=��O���+Ǜ��-IE�)N
�ǩ��^v�fp0������l��`�v<9;gd�f�3f5��3: yqܘ7�H�^BD�8�A�W~봷���:z�lf��ԡ�J��U؋�,h���o/� ����=�T����%V�HD[M$����A��\�����?�
B��>Wy���V���;
��K��p��%C�n�A7D.	��k���y��V�1;�5\�]�&���i���˙�����U�Z7xܧ�4)j%FQ�%#W�YFkƁvdO��1��A�Z�|�۵R�D�h��T�iY�Z��<�D�$.��*S�/cߵ��P}"�/�4���qH2w���^d���T���6U�.w� ��	ej�^���O��/�i)>� �*r��8�n>V~8�G󇡺Ll��Q����?0��Y�ۅB"x{��H��is��� 3��Z��n(1�|W�����ZfjU��v5���r.qol%� �ި�X�7w��s�#���x�؉�\N]��e�.��\_�3�� ��a�~܇ٸ&��#�=����ҿ���XQD��,mE���$�ȿ�co����� ��g���e���`�`�D�[W�R6�&u�}���?,"�1|?<F��Vg�O���]�~���4�e���I�����fV'��݄�c��ubw���˕I�V����:AF�¡;�BE���e�*����+���@9�";������|�����6´�*N9�aX�h2�0�q�D�\�d��B�wg���PqMLRU�_��z�+����p��!���/A���σ�Dr9g]HW����X*mFєU�5FV;	��p�pt���G���
�������^�ࡥ�������H�k���5��/V$�P�-��R8u�Io	� �W����?����3����3�������+��}�����$�m��'<��j�#�THr��q9 �ȣ�_t׷�t6��5z�R�ھ�޾�DXt�1?�C�9c�t"�V�Al�GOa���u`��R;�DDP��핍�E�1#1�$��\<0ǀY��ோ<��ڝ$q'Fp�4g1���i�QӁo�2��˙�D�WL
�L����o�a������p���G�����M4���4K��yo.@նS{ �X�Rg�0vb���2��ά�w5��W~g��<���6��//r
?^3)O����Ы�w1��O���'	��
��Ш�����XЃ�LV(��P@��(��\�n�&t{#XX#�SG�Vˋ^Y�v�[�5��Յ�O���MQ�nB�[	n\�6"����B�>g�胂t���ۦo,�D%C��Ӓ��
���m�#t�"�J��8N��?�ѫ��Ñ�CN.Mjl�+
�2��2�8�
���-�R�ϡ�ATn��<m����DH��d�@�J�2�-� �cJ7����J޸�Ѯe̖r���|�o%��hR���Z#�h� �Q)����� �9�,8e�T���L� �Y�l2���m`��!��>"L�
�0b����54C>5l��֠����ɴ�ѽ`up�`Ȝ����Y�9��OLoK��_M���5���;*���qC�}=[�?��ۣ	:��@�+ʟ���_����Zg��J�!Z�����R�b��{���V��(W�<Z��E�\S�\"��I �"���#gEl����}S�e��ӫE&1�8��i_Yb��l�-�`��\8Y�(����z`�{��a��	$$Ы�:��F�A�^�\Z�K�Nbߟ�����/7'-b3ɏ4�iR�W+c_�}�*9������E��l
�A;�Q���	�)�<�x�x2N�9q��^R�4=H0�t�2ig�}���5zvľ�0Yɛ���T8���2��*��4Y�{�竤����ܧ0�A��&}��H��-=j�n��Zr���d�[�����7!�#T�Q����&�(���.���9��i�f�	
u0��E������W���Ǌ󇮙^S��uh�*��3��:rI��[�hģY��t%�=Y�����.�EU���oZ�Q�q��$���}m�,�p6���G@��_1&��g�f��d,���o�9W�J�б$�6�',��D�������qܣ6ܦ�g������BA��)�����W�s1t��(|�1� �\�_��������"\��)%�q�K�s/(X7Ĉ�f��۱��>�Qu*+*[��tL*�s��3EP\k�7�/�8���Q�i-��P�$A�	�R��/��[w\�UC�
ğ
pK����O�'>��x����φ��M�sɓ�Fu��u�@��7�/U�x��l�d�aL����t��=��<����m>�S��@S�5������MG��,��7�L���p��^;6���U�M՝�ڌYn�Z ��Զlg�զ������Bx =<c��>���Z���Fk,�.�x��=���W��"��n/wpr���n�U�S��Ǫ��T���� ��.�LB���Е���I?A�&;��D�{��0�fq}�PRU
a4n��Q?�]�����ZP��GTC{Y�Y91�)�]Ǒ�{d�
��s�Yk��<�p�}�Q�����4� ��r�E��eӿ�]�>X��7l�\�c��O����������TX�B�mGQ�Wk�h���?{������8�ËqmYd�'�p��qS\a����{)�s��4�񚷽���W�[4A�/U2��V����� *4��%�8�F�L$F��󕤾'X"����x�V8���>u<�]}zy+��9K$��'ƙ����N,�����;5~���j*�S�axiW�\i�r,B�
���0��*.���1sR�k��ޭ�Q����Rt��s�a7f����7f%+c��D`s���Pw��Z�����"8�W�	��Fx�(EQ_R5l��>͑�#2f8wn��1�"��^A�ڿ͢*+��-�a����1S��̢�B���ha��G��e�հ��E�˺��4�y��~�\��)��y[˱��$�62"G��ZQ7����l��c>*U��ހ%���}Y�4�e�m����GU��v�V�?�5�Okn$k?�O��A�x^��@���A�v�>|��SBΙ��R%i�^�̭�L��JSJ]��f$D�1��S.C�I���.�6H�cܕH-�zeC!L2��XLx��̓�
U�R�S�CJj�o��z���z���)�ø.�p����\M�琢b��/L�����g3	o�e��(zO�h��)�c��A�t!�o��Dp�4���Y����ʚn!L�_�aî�����AÖ��nC��O�q��lnO����R^J���g�L9j�i- q��Y $� 	�6��֕;V�p�?ѫ��*�ĚC8��.
�ץo}�a��	�$tQ��B;�Jֽ���٬ɖ����?5��Q]R��s�Pɘ�</I����/��~�=�0��Efx�3T��b~�d���g�e�iy��a
��#$4��l�9�u������z����n��b
��L��C�9^O������ ,c����n?|5�!B���g�g����&��"���� -�|5��!{��>�739�2��t��G�G�K�\:�3鰮h�����K��U�MmG�ѪZ�� ��t�(��sкYF�/�@a
u��ႇ�h���m��-?:�˰Á�U|!��.xJlڊ�A}�Im����v�Q�!'��*�gm�9��3Ƌ՛�����ΩTT�#k=���_�
SR������L,>gN�Z@|�Ŏ��FL�B��Yi]$�~(���"b�Z��Č�"���E�	L-;&�f��T�fyb�ʡ��L�u)`�G��;� ��*f��V������KD�kҐTq���a�%(�Ye�]��u�b���0��R��șjXm�
K ��]E���q=�M��q���پ���/&E���ևU����%~gBAڱ��ڹ��t�A���Z@@:/{���r����V�2��y�����c3���'5�lo�ҏ���݃JZ�
�A�T��;S�~r�}�vv�=��{^� ��˭SS�C\bSz�Ar� ���A���A���m�'���aM<r+��e���3U	�`v ?4v���h�� ;���$� D�0K�!%�oR���U���j��y�3��,����4O)�%�ҮJ�Gddyl"�A���a��.�ѱ�P��j�x�t픓�hՍ���	�kx�f�/������UW��l�RϽ����>�����#��{���ܽ�l�ϗRNd6�:p�njM�A�#��%�py���m�Pݪ�^�J}�����ǘ_�7Ed]m���a���LI��n����d$,b��d��m�21c���vc$�V��y�� ��(~Z����
4_�9m8��(Cˈr��9�L�B?(1�*��Qk��ٶ����|�DMQ*-�:���F�w@�k{���KC:�N=���͉��`eJ�V���~q.{b=��>_(!XV<% ��
�֍��S������'�џu��J��L�$�.aC�.�C+*�"�&|�c5)�S�_	d`���CKP�$�����Z���x;6�p��4��Y��p�v���僮~A=E�%�D��{a6PV���-�)��o��6�;w�������{�-�E��gU��������]n��Q��������(C�36F:�*�Q�*.�,0j"#{ܗ���?h���B���pnZ�ښ;�0�Eg�^��Y��f���6��|�&f���t�Ð�9-��+�r&�"���.%��>��`<9Jf��4��=Ru�ڷQM�\�YÐFŰp��z_ڊ������|�4x4�/�}q�d��=���..��ܹ�2�`!״8Q��X����'�f�#' �z���Ǽ���g� qv�D��o-��OY�7��@{�� P����r�D% ���6����Ȇ1�5���5��4@o��I�_Q$hJ�?����;3���k��h���8k��'�����Ǯ|h�-]=�>3^�w�I �J��N���Nį���*��3l��r��k`Z�A߄�7�L�������P h�5Έ8�����ހa������-�Vi,d��p�B�F>����(�H�2�إ��oQ���w�6��αʗ�m�Z�PBuThF��6G�T(d������Etr*;�@��1�2�/���d�E��x�c�3���-���w��蕛0�&`��m��:��h^�[�]�9�A屮�\��	%:�#S�h+0;c�Һ�^�`h�e��3+A�oR� �2$J�Y��y�Tm��0׸1�\���[#��,.�k>6@޽��"8� ��M��E����oxڞ���f��5���['���qP-�o\��# l�$�*���70��C-S`Q9 ���יi�Tv��`�'��/'C�΁m�r� ����٠�ciwF/��LH��W-G�e=QQ�-ٌn�A�NR�1�k��=��4�!����h�Z!�XCHwG���p��V�_�n:Lf^����<�C[1�t��P�ZS(ː���	�������W���x� '!�6�n���U4�'?�T�����&�u��E�_<�҆&��Ny�ZC�4Ղ����ޘ��s=����� ����o�&����-X���ch�����݊�W��>q.�ָxItݩϧĨ��{t��rǡN6��>ل�>�W\��d�Yw��pŞ�ȍ*�,ֺ�:>a ���f�M��,ݜ$�-��z���n��I���E��tE�''����z��!׻e�ų�Ay��j��V��Ѓ�9$p��e�ԭ�
?���3=����or7�x(�I�D>���It��ȝ^4i:�ĿHV��P~씭���Ñ�����ĸ�d��z�]�����!��\�lvw���bV�	��芠�}9�8��Y�.�� ܋�J�S3����c�R�?�۷�U����ۆ�D��-�z�[�]l��7=��[��b:�3�khIK�y���RT^�1���k�J�M����ȧ�I�$N�*�S��v�N��  �Q��*�;[<G��w$��6�0[���c�=)�;��:K��1%ҽ9�<��"����p��/R�E�1lk�y���L��A�L�ۘ�)e��q��&�P���e�p�t7��5K3 b�ww�M�v3n0���y�����R����ɱ��������l0-�ݪ,��Dq:JT����s��nH] �
���,��:��Č`��0�Xo!��1��-��)XZ��]�"(%�Tn�̿���( �ї��.^�H<��o��8�c.�&<�s����+7���|$}��FQ~}�%������/���^�В�S�cf�R �Vy;XZIR��4�ז�0����a?Qt6��q�I���ri�FC�sUel��q8J���+��~c5O�7�'W(�IB���Bj��7�U��,��AL�%vJk��!�)� ���,ح�{n�?�]�p�.�k�4�D��  �kR�k����3�Y��5˲�~x�Y.Z��'�]�v�-�v�ui IS��2�(fx�zgX��*1~��7��I�������Χ�+��+)n�G]��4/1)jhg���|V�f��6'�\�(�ޏ����|�c�ul��8�曁c�
�Y��vqq,mnQ��i�~*w	5�'�k��]�g���G�s����&�J��@(���Da���'C<�uQ,�H0G�E r����������
��{땲я�~�$<Ns�2���:R��g>�m�B�w��\�Q����q�D��M�ET�N�q�J�����(]/�������E�7�[��rq8<�բ��nz[��	U�Q%A�^�J���gC�0[����Xpgf�*w�Ν]�s��̳86M���>L�EM17-��w����뤋2����t<q8�,;����:����S������g(g�%6Z�8�A\~� ܽ��п��%���[�b:�v44)� �ŷ��B�{���r�KM\h܊v�L�0B�д"�a���1 R���X��{\��/d̡�)y�3��i�f`Q��Ɖ����%(�F��,�(��n���O#L*d
T��p@	FQX7ه��xpSU,�W��йs�Hⴃ"�*�b�ߞ���t�C'9��+�� �)�s��ŏ� ��j�n�#�)��
�n&��s�sd�Pթg�':���j�'�p���y_��J_��n�2��H�]���OԪ�˖T��<��#*(�K��ֽ�D&���8���,�T�����җa:#֤fX�GJ3����;�,�>���Hɵ��PNVO녛�2���f�/�2=����ݡ�^�����ÆH�nB�E��`���O� �(+9Q"��ʙ�:y.�A��.��B���p==�ˎH5�q�,nV��u�D��T A�i[�z���}B��zFu�%ă�xLK����\������bڵ�#7V���lN���d��^<id8�$�E�o��4�qq��9���C\y<j��-"��Z�P�H�8����:<P���_V}��'�ν�KQ�^2k���S�MDǞ!;P��M&c�+�%%xm�\��S ȣ�7}���f�|�=��F�O�%�����{�U�������PJ�9.��ZeS�Ca�H��� �Û�L��ns�'�6O6�a�w�c�_*,{�{�� ��,�KRԇ��6��qՎ�psgn��s��RxB�C(�����x�O�f�ʹ�X�����IZK��6%�%w$�:R7�;Ӫ6i��[���+���h�#Դ���E��=q���S�C��A���
��!tC��j������
�c��*�v��	���%����٭���Bt��D����+�T��G�Vb.�fzOqMBY��XO��F��ˇK����IQ4l�\k��!@Eҍ��!W}�T���q�Z��FU�T������h���O�B �w�l��S������<�#J���'!�n� 6ՓR�C�e�J���q��N�Z&�e(�I��2����T��k���_$څ�\���+GgYSΗ���?�\
��E�W���Ȋ%̅�v��X_�{V @n{��.o+N�	�]�ՇOT���w��t��(-�o!
M�w��{e�]��!���cu�F�p�I��JV�h4	��M�����
Kr� �c�/�g�h0ˋF�1	]#J�;�d��'��8��L��� �Sn9�P����$˾)�\HV��I�?�>���R�u7�?f�û��Z���&��.�����H���M��A#ƅ�Pܶ�ee������}�Ď� ;������[o*0�xE8CEa$�۳�����=�x0�����5��d@,���!dh<�����Q6�[�W���b:8�Xں1��������SE���riգde:�%��D�L��T=�~�{��t��I��B�/��f�SuH��zE��2|ģ%_��>��%�c��7�����0��b>^��ɋ���+p�cT���E�\�Y���	��as�$y�tU�o�ۢ�t.�#/�X�+�9�&˯l�K@�PyY���S(��e��#��2���̄ֳ���$�������t��"���9)�kt��v,�.:���*��&�}�4���%h�RaүwT�K��/�����x�"t�lŏ+B��Aژ��ML�S=b�L�et�_F).�� �>��~���%=N{�� �`3@�˂t�zb�7�B��A����`�X�����M0d������&7}�M.S"DTP\�9���N���mje6,�S��ədaۼW�e�?u���G��aW�Կ�U���%al��F�K>ٽT�5�`��n�Sr��<�Pen1�y�jA��ӇwD�n�'|���&��=,Ƿ��;J{qܘnmH�f�P���b����ҚJA�NN�Q1fe��Yl&���H��vf�#.�T��I)v�S�~�Nl��O���:M|WU�S��FQ��՘8>[����2Y6訦��M�$/���/�ML�Ὶ��9M��AW��9�7܂��qZk)x���PЎr �S���@�^�f��â�F�ýݿ��ev@�֛�9�nRy����u�w��7�5�#��ӣ�7쫜4*�b�� ��-�=o����w���8.d,@�S��T�Y)S;y]�=��K��D���2����]���KUµ�Xt���;�ĳ�8|+��&wJs]��L�ƔV��/�jă%�ɶ�vj��80վ˃���x��h��M���H8���C��y�گgqb��}*�6�c���@-�rLD+�z�޶�M�Hl�b0Hß	�u����/�6�_�Y�i���b�K_#m׽�d7���-�<m�@��%�z�����T�$��r�1"���؂�]6,°2+*��P�i�9P�Rww����]ф���о�(�!J�(,���r:����m�/!NsOWA����}y}�ʀB�<m��!VSSO���7�:g�y���Txު6I�:g�H���8��B��F���}r�^���$������3��!�h��ORXA���@�V^�N$)����#�9�MI���u
�KGQ��}�'���r��aL�g϶����ߨYp�v�~���[쫪���O�8O�y&������=����M�Bo��[{��cK��J�"j��RN,O �j��4����ٿf�6}`֔R�'k��A�OR��Uؖq��<�����\3�Lh9��Y�5,O���v���"���&�	|���z~F�LF�Y�<�R��]7?�洍�s��Z�A`���u�~�� e��Q����B���
�*8t2�`��=���9��o]+�^b�.y�*�Y�}�f�"�%�L�'��z����m}�̭&�%bףJ�'�C��]�n2��N���h�h��2;��UOE��f݀y�B�AE�-�V�9�O��;n�v�_��0 2��iḭ̂p�oP�+<�&طg�?{���J��kNB��D���@T��
hM<���1��A�@�q^��mV��v�4�Qbx���zny�$IߣZxvv�~E!�x~y��m}OP�JYU��p�{f�ogw{'�ꪱʃ�����H��DD�Y�h3�k�V�<��^��zK���<C%�����)�)�I�3����~r;xRqӅ|}2[�J�F��m'5�;Q���^xa*��,+z<�$�U�y+�R�A��Ikڮ8:�>�WA�jbWқ�|q /p���=H!���\���S1tF�&X�Y���TCX��;�X�&Ш�<���$)�&�u��_��+i�+^֬����/��6������Պ\�Iw�Su�ڗ�V�.���w?9����r��\��ZyB���w��U�$[�}f��3�} �:����3$��w|hU�A_G���dݾ����i��P�̫l�_��滽	A��[�Yt�$A{#�LvV�T�I���]�A&C���	b8�MϨ��q��Ժ^�P�e�RX��)T��e.n�������A��(Z�m�L���yt�H��_@�W��g(��K5@��|]�\��҅0o�kI�>�'8��♎�=�@d�Y��۷�7�1��`�8����qܒ~�s�;z^�K
���':2F���U��i1�*=���P�K�O䎔�ywV2�����Jc>����Hr@'�������V��"-ٱIX:���׋Z2Vi�]���P
�at�ʚ&�jX�nX�i4���lT���J/�ں�L��ޒϦ՗��G-����AY�1C���8�X-���#��_,��gڐ\��8���p�۝RTտ�=��!�D��k�Tt�,�_�S�Mc�z�RNbrN��x���Xś=z���Jy���������c|H}+g������-��
k7��̡����C}_�y��,,�;#z�~O>��P�����M���8��xQ��S$d��sl`�'4�s�U�W�w��=4��|K�_�ˬ��CTY���H��a�H]\���nBng����ad5�Ph�n���6�X�9 <����Y:���2�{�W��`R�J_�@�7��wE�,�*!��p��u��g�k��(�F_"'�#Y�z�̨��1��NeF���Z�t�G��^{/)�*�`�I����Er(�s�@֬:��9X��b�'�~]����-Y@N�9�l/D�+�ߎ�`�&k�	˓"sG�[��攆o��6�����xЮO?;���nf��,��g 3�1���	.P�ڢ�4�s�vq�$��IS�s%GDZ��Ydٻ��o6�>�*��="Z��I�"ى}��R��Fd�i���o6�r��M�=�ӂN��������2��A�(�xĲ�K\�Gc�b�Y���l����sh^�zQ\;L��!�+��\M�R��T��{۵��.�0�F�*D�W��+%����iӷ�)�l�o,E����B��鍓��H:|��]�M%��8�t�Q_��ՠTKs^��HQRo�3�^��؈�LL�c�%��_U2p��]��W~:����#��0��E"�i��E��̥��"��Tn1���_�Um �(�&SAx+���7m����C{��wvd��2��� ̱����9��Y(t^�)N�mb����#N7���khL���>��k[�71<��礇�_��� ����hZ���r�(�!�fZ��C�z֜Gs���!��Cv	�"���]d5:��9=������r��b.I,�^�b������>��`��@`�a�k@�s�mxѾQ��S���'H���Hw݊u���M"����`B���nI�%,��gy���ƪnu��0�Y
f�?�]�K����<-�����fV~�nMu�ڱʰ/t�|����f��g]f�S��<�s��3�:w�J�Q>���{fʑ�ц�9vj���`ZXc���|P}��9��rvh�_>�h�_X^��]���b%�����Y�̒��� _"��ާ9���!bq��g���1̅�I��'KN�<ǿ���uYs���q&�$1b�:�soc�mF��\[��D�BIeNT:?��K��pƟ��^U?������|�vl�wL>���,�	L�}1����`t�L�&0���
�/ߣ�N�!����N;OI��|�Q8����h���9��F�������	�;JI늹�]�j_�J�StC�����.�G	+dǽ��tP33�W��=�����`#������.�:��/0Jcwg��%�)@���i�kD�S������=$���D����5]�W(����&�e�)��I���2������^SC?aY��Y��$Q�{��{mW1kŵ��l��!n�ޚ��}q��2xo�5�l �D?q��,HD��	�F���m������Ȍ���
$($f��c"�b�j{zǙcg~*��[��u~�<��.ԍ�|JR�_�k�QNR?��X�ShC��艩<���3��[R��pw�8ۻ�f\8x$>k� �?x�Ph�
u���
��ϛ@��<�W.��3`�h]��z�ԥh��B5ޯ;(D����
���q�=�?(=q]=c��h�H��,p>=ݭȭmA�a��u��m�˔ ����b��?�J�\����H�џ�P�b��I��>U��̫�|#D�"��~����s���[:�����/���=cEM��j�=���(�	�r!��2b������xj̳�r�ETc���M�ГQpQ�,i5;�}�k�`nw����6�^,g��>����2Q�1Z�����^��\��<wb� ̼g�̰��hvXˑ<bP�?��e%s���6'�cҘ����joS���ro[(R�o��fjmK�>։_�"Afd~cW�c>@2t���VK��]UB��v�ߠ�)	�QW��5=<�e�Nn���h�>���A���
ޙD	�����A�<^5�CȂe�d���!�����OM��LwF���r�-��&y����[��I���yM/O����ms���f>�{;n�F��h�ɝ�з �0��YF��ub��oϡ�61��.{!x���.���P��ȋ�(�$�������QjZ��@wnO>g:wp,��y y��B](�|v�<���%��
����FN<s@�>��4����'KyW�\����">"-�ƶ���0�B�mC���FrgL������]$Px�UU��6ںW�=�Q�*�|/8g�[
�W_1��}B�����KZ�p��Y���w�,�9�����ӵ.�v�ܣ'���"`ނ�Z
l�3*�(����K�|�"�M��3�P�[�{��8"�
��2�3w���	f�L����ˈ�E�L���ҷŮ_��w�uU�f�4)���������W���8��:��1��At���������͕�O�,m3
)G���H8jp�~�堏�!�ů�&����t�M/i�+�>E��\�җl��1@�O�fl��[)-I�}�ׂ����nGp�E=h5�*4ْ%�c> @�^�����u'Ɏ�e��o9 �
���sq�@ �p�y�d(�jrt8�(]�5o61��{b�q$�k�q	-���;�'SBC�� ���]�m��.�o��Rw.������L_��d��ʋ����F��k9�r-<�S�|�c��]هA�c��j����߿H��P�h�|��,�>��o��t��Ʀa�&h,���s���}���!�n>����l%?��K"���i��TfQt�l�MaZ �2EX�]]���~�'�Y�gm��e�kk��	�Q���~�QD�7,��tq"`�?� {�������-}��	;�5�Yw)����ÍL]`��]�$#��O�<c��nf�G%���PE�bg���\n��NhpV�.X�&�HL��������,j�ϥ�c_{�NXN���xA^�;-c�޶���t�����i���+�!��9>
k��yٽ��=p|�4�]�>o�@!���Ej%u�#��ͽ�r� ю���[���@ʌ���Y5�C̘0Ț�wSK�g��^�8B2A��s�ZNgAkQ�e�d֞x`�c�]r�Үm�tAH8&��L)�������Q�a�pf���Ƅ�Y����������S�SR�Μ�r�����I�zp���;&o�xP�. ��7*-5��}7�<��?�ǡ���-�1����֠��y2o�\��?�P���Q�\�X���#�.��Fz�;Λ!�x=bS���fB-ړ-ꄽ;=��W�O��ƜY��
���c���+q!�[ #q���m?����Jght�0{�q��#��C#ki��K�ȳ~�)�hm~�d����Ҿ(k��X	�r50�D�q����kGT�;=Z2�a.@H ���XRD�:w��vc�N*�Adɡɞ��5k0�p�w��9's�&R�)PAYB"���R�#��D�_���
؂gj� ���Ks�|��&33x#]��ȡJ��ȲБ:P�j\T��՟	� R{�ͼq�@6~��<��/ 	��vH��ӥ}@36�?�o��3�Ǒ�_;��nwƝ�o�r���M�����fZagA��e��|8���t�@�K2@�����0	 ���zf��<�%�;b�kޫ)�MF~��c�:���ʉ�������^��`x��![�]�[�K)$H񦺣�o,�1#�@���x���i/]�X��kk�CPS/�$��=Km��>~�u�P�Fº�/�{�r��,^�k߰�%�Fi���٢b7�cƶ���3��^�B��̒��*�^c����4�8�'�fPAu���o�)Lβ+�����}���P�C��~e����O���$��.@NsN"j˦�����i�ʀ��{�$����BD[G����o�N���ٓ�"�^��<����躖�y�2��_7.�ǎ�8�$�)����]��[���|Vy���F���sx�G�~�c���}J��Q�^3�5�Gp�f�J��9���bB*u��L�h�˼�YYs�.M܁+6��S��"BJ�?ؐ'F�w�n��:+TN�b��!aW�d�F�ni��a��Sx~��Uw��#�����
�2u�P Rź	O�S�1���%��t;!CuL��k�5YB��ǙX��UC*�'\+I��n˶��cm��/�%�O��K"ܫG]61��}�����&��m��>�j��AP��r����H"�
棣��ڠ�4�
6��.�����ɩ�8����J�t�e⬣�Z�׺��M�;��b�c]�,T>�D�g�lg���p�H�`(7a�a&h��1�	�ܛw�z�9����eK�9�՞{3!̌��:�]E�����t%/x�;g8��C*���uTO+bK!�&ٽPԿ �vA�_F/XP	_aS��
���Sh`4$"�,��&�Д��T���[���c|m:-���9�E�oNA�=�}�S
Q��v"=Oq���1U7�v�W@@�y��l�����{�|����2�0�c�#0���_�-��|�s?��Y���-�S��x~l?k��j�B>�t1�yR�Q?���T?5�<�]ҩI�=1���X�f�v��ǟ�#Џ����-+*��p��N�-" 62�����,�V\�,�\�kd��ecM��q=��A��S$�^t��D�݁ۜ�|	���_,�.)�ec�2���>v�F�r��Y�W,�?���~$F����tf�@c��t4��$J�<��Ph�H���u����Jj9 �ؿ���[�> }�APٖ�Q1���)>`m�<\&��< ૕�,��^�-�+��>p�tKH���~Q�8����rCDG	� 4����ᯗ	��O�:%��gb�*/nmv�l��ԞƖ}{��~�J�t���+v6Q����R�r1�p�y���s@��Q����j8`-�q^�H��E�?�t���$,L��z�>�"�a���Zv\�m�]�Q�n�m<"m�o���4:��`Y񱿚�Ӝ��vi��?0��`���a����:]�0$^>�F�PG~dU4M�Kp(U�D��YW�	��iaV�XPs���3QZ���ԁ�<(�)!�,��?���\����'(��m�S�����T��\�> �֪�{�I8|�~��i����`~5��F�G���D]Y��w��C��/b'0X�Ϳ���錑�,�	��W�'��������Vᥡ'�zT.�(�bk�����I@�A1@^�e'�����L� |fT�Q��4lr�WY!���f� ����o�hz��L
�I���ڧ��Ʒ��E�Og"!
E�7��� ۦJ�&ƿ��o2���A��~�{����dX�L�?@���ЗS9c�u���dF4�R���q��r�/�AV�.'�Rlb9|"����شc�Jh�|�0G4=���k:gU�1	����D&�²��f�u:�c�55G�Hv�9
f��\�J���dI�sU���{x����� ��\����ɏm�6�H��\ ~��`� ���dc�j,G1���GiEz;)P����.��Z�����5�7�'����
��,|�Pwd:��>PN���1��I�S�-�k�᧳row7�=�������J�r#0�ܖϙ*T,wlY����x9c5���Ky#�����	ʊR�����[��X�xy-�����0�~����¦�K9��0��1+���&�dn�d��T&�\�z��M�DO��^!�`�c+�?�A�O�i[�j5){%=�}N��/.��R�v��Y����H#2
cu��	���`_@��j�tY����o�=�Ctz�|oA:�����:M�`*�]�{q|���,���$3505��ˁ5��Ww"#��f0�����=�U�<Y�1?�uXk/;BG��=�M���/�}V�S�X��o%��
3ux��z-^�����R���w�V[�X�z��]X������f�G&ʚ�Ggx��Y�t���?9}u�f߮��fd������_?�*�r�^�[��^g���x��~xI�4�@A4Pgб�Q!��	�KI�����b�b��]�j�n�3�����J-}��;���\h!���F�w��`�Ȳ�3��b������( ^��@KF[�X�]	5rha�o��璬���=��Ia`/�o,Y���	�*��,�Z�A����H�i�n�|���5
]�1����Q�?�_��L83�k
5(�ɝ�+h�ٛ?���/p<�:bZ��.O_�䜂���7���?ݬ��_Z[��G�c���{uK���|���������"���V<)��Wȃv����E\T�Z�Si/���a�����9�� �п��kP��Eg�ғ�jⓡ��~��'��Bذ<���KӪK�1��ܼ��(99�崄ڜ�(`-TOj]67կ�0�ʫ�:l7��yGt�sgj���^=�]11=gv���������=��;VKeϺ�Vk�0+��(L�wX�狣֨���a�h���U�^1PI����*��8=#��,���0h���D7M6�H�E6�3����jXuU�%l�e�sz�h8�hҤ�1�ݺd, v�V�������`X��U���=��k��b��W��8*Nw"=]p1,���B��0�ԨhMN�d��3?�Id�wj� �{�$�B�b�	E(��(}�闍�?�ں}��s5o���h"<���s�{��ԇ����"1�2�� ������4�+c��/����El��@�Y&|�6N��������.Z��6&h�e��*ϲk�/���]w��V���I��GyvI"Pʯ��\6^��=����z��B�|�݄��r`�&¹縂\���x���a�ᬉ�1µ�&ʫ��b��`�L;�e��M�J����Ԧ=���g��Vw[L����U�פ�5-���\�b�����*@��b��"\�$����c���nO��ʰ^�:@Ӄ!l7�H�e�i��ߤ�=��Y9�h0�ݵKq2���8phD����������)���/�������o*�8-HlR6�w�����\֖�͈���!˧�Jˢ�J�V��~;�0.��>��(0 lס��a�MbyN;�eJ]��T�B�M�wԋ��o�Z�ad�]_����H��0��� �v�=6��'8YeI�ºPTeǬA�~�&ޟ�.֩a5P.�4ﳼB- M7���c���&��?��/��J���1z.|����u�7��-6�K�d��5�s�sd�5�����I ����]'�h�z�6�CY�����ѣ�3��qs�P%Ow�M���l�`*?���Ԉ�>N{���yP�����l��dk��5X�on=$&��B,����qO����&�1q����)����f��g{���׊T�Ș�ϗ��a0����(��à�z��}KJ���UyI�#ţ���u�V�V�(��-�J* �s+H���e�1�?̬�}���r�����h�K!Z)�W�t�n������&��KO��V�.�i垓�KͭV��-�]A���9ѡvE��1v�K���P�vL���d����y��sݣ���u(]E�8���ep��sQ�Z�Uf�KU���ɤ6a<��?L�ا���׹��зxW$��w-qxI1	ŭ�$cA-�1���(�ÉF�t� 4�'@.3�Z��I�6�7
�'��^���j�P饯8	�
��o��u�2��F�TodΦ�ub*f��?{zَ{uz��sW=-����Ó���˾�|H��?� �������"��F���^ؿ1��X�X��̽���\	>��P��,���α��Sd/�� �$<3�B�_@� ��)d�G��驢���ի6��/�k⎰ل$/O9:������P$E~�^�r�x���F��"�R)@<|�O��4�K�n��U��,AhˢϳA[8�n��ǝ���bN�i"f��
Җ1yg�L��s������'1Y3�_�>����M���-ML̘�n�,��7��N!nq�A��^��&��D�������aߡ�7%�"o:7��1��XŬ�^��b��2�9�%3��$��DJ���CN��	����(��L\���u��UR���Rܻ��|1Ǖ\W��	BؽQ�o���3��	��>?BǓmZ�nV�ƴ�r���2� i��S��c����:�S6�6H�"f\|{y@z�Qdl%�]�L� ��E��k�*a_9�3��/��:7:�'(>�&�Sٿ�ˡ0r
�F"���*�2��B��g�W'z�A2V���b�sbV������{�ݎS��K��!G�tQT�bo�U��p��V�tRZ��
�#bv�)H�
qԋs��� ��`>��X}�L^����{!5F����:F� �w�����>��GD���LJ����	���,�Z��1Ր�������]��o����ɣː�	6W���9�'#���Ǆ�����N(�N7G?��ꎪ��A�w��+�^�k�#����Wz��KBW�'�f�.R,���ҧ�٫���ua�.�FVI=l�x�1�m+<5K޽:l��
�P^ՠ*���3ş�fe��w�D+�X�`�=��8#���\y�V��ypւ0.k�r��*��$��HK���n��y�&!�4�"B���$��0ǲ�W]Հ(�����}�0S����eB�9/:[��3�%�>6�Qw	��� BR����ɏ��ߔ��0L��zK�x������6�F�Ɯ^�!ږ[*7���O���֨�Y�Xm��(PN}jξA�K�����q�5]�Q3�_i�j=�`%��w�o�Ӂ5������?	5�+NJ�$�ű��wRa\
���rY	��9㕜{��R��iȯ��V$��Q��B���0�op�F;vT#X��T��"e�c,ى�Ch�@B�3�Ư�N�br����-/�.[X�h����,C/d4Cc(�k��/�L����SP�r[�
���?���P`���]k�^5Y�o���P�S`���߉���P�[�[��7��Y��]>K��gF��&�1O���3���I��&�+*����i�c��V���x>�;����=�~��g�����7�֓��+�J��>_ْe.QX��8R3���@c2`�������������`����l��_yr�F|*HS��y=�n7D���b[;��i��Z��P�Q�����։'��L����9ޭ5�������n̉yi<8���Jh�w�`�lQIt%kb(2Sh>���Qz6#�^�Eu�Leĸ�
��нa��P۩>��g�q�ٶ�W#W�UY*��ʦM�{��&�xH�~� ˦^+7"��(�Mѡ�W�L�Ӧ���֔���z��C�PK�؈��a�|{)�7��4M�q�/�Ƈ�p���9�%3ߌ���NG�t�>A{����Y�;-Z�����r W��'���)�����$�'_Ǎ�tI	���ҕT�A^|�m�>��!� �x�{�zG$+3	,����wW\��lb�������Y�$#����x���U�MK�"
�ȓIN�,nm(-]͝��B���D>d+�q&�Wkw���6
u���j�����X��b�t��
��n���u����#{��װ�3�o��YH�%��.�x�Q;��,�wqq�d��W$5Y��GM�"ѻ��H�2�ؼ(�F\O�	��MgJ�&wJC%�þy������X����E�u�.w.$ $���c���t"Ϙ88m+I��c����p.�Bd��FE7��0�3p�:$xfY��ɾ�A0R%H�ml��ƛ�d��\Z��,�����'�M&��VB���T`,�����n�w�׹�}<��u��Ώ���z!�`��v�̈8l�43���{y_�קt1�;�(�ِ�x��P7�}�`9RY��:�R-�/��
2�#�w�ݦ=W�#A�)3�-�h�~"ݠ��ϼ*͙5"@+'���l_�D=��z��fk--y�����W��
���2���Y˩.�j�PFb0ӳ�X����LC��ʩ��
�6^V�"��d�^4�[R������x_c�����֏|P�\
���;��0����^�����vp��솗�:���s�e���&�}�񈘐�Cm k�
���s���s��Vq����;P���ڍ9*�M2dL_�Y^9�@\�:�R9Z�A� ���"�έ)1�Z�+�R��jm��a��~!k�����U�]p� 8�&�S��
�D�b�角�ē��@��E�؁'�y��*�|ʖ^؆+}�jW��~B�0�:N�w�[8"�#,A�������s�Ni��d&ν;�-��t�-���UV5  \N����tnu�����R�]TTѳ^tް��&�`I�&�=�������=�}������͊mڹ�%�>�ܐ� *H�gUض��_��S51�}���u��³�xQf߰��\�1n��+�;[����w�ٺl�H�L@[5�K8��p��͜&����?W}A�3�-2C|M��+n��O�Ӊ)#!]��Ƿ�k[*���{���"���u�u���O�⣙]�����g6���jL�w���p0#�;�ɂޅK5K��ȿZ�;���%� ��g�������3��{�2� �:�L�ǂ��:�/�S��u��2)\�dȴ3G�?��h�2��[�7E�����HgV�x�"����j(l ���H�ik^Q���d���J���I=e����nd>={3������U���lb�A�?�>eM`q}d�.PE���-��8;�K.<wf�kp8�T�L�B�:W1��Ȇsc�1sA�D����U�&Iq�^\�0p2��E��\b�Ϯ��/����|o�{6�ˆ�������R"N�zT�ok`��il\O�v;�#B�%���P�O� �at�&5m)����4E����(��]�!�l ��fuNqp3s�XR��7����ŒaS��!Sh��b�}��p��	"�$���G�s���0��(�PL�Y��U��~Z��/|Z��f��_��C
�BU0�2�7.K�H�� ����s���s���'�ֲxH�7\F�8���}W�'��ˁ)<�[�e��)F�ԧ:D�r��};v������O_�ƍ��v���	D�Q2�t�����$����}b�,2I��睈� �`�X�{Ϗ�;5�E�]�H��	�AHR�.�&lm�[�ݴ��d��Y-��+	���F�~�������'S��g����!����e�1�~�����tYۆF���˶H�S4���b�4m�N&�
<��NxOrګ��B!�� �yj�tx�9��)*�4o�Ҽ|���-�	��W��y��N_�/�f��@h�[�N��I�q�.��$"���/�Ȣ��r@�`���#��iC�tF�.�e��xd�pKЁ.T����a!���$�lݽ\�=�W&g�c}B�
�Z�R����q�{����1��(EH#Ȃ/�qn֓�m�vIT*��&&yU���8O�����7���so�9=� 9�&R���!�Ra��A���MV|.��avl�������ۍbD\���m��@�qy��P�懐�Ƀ���>�?-O� V�b�&o��W}���In`�Fk]؀<��{���u�?���l�ؼ��n_��G�\M۽��m�Van���܇f��Z���Z����[���;t x�D݊��悸��Tz�y"���@9�?=��#�ui��X�6�ß8���!c`�7�p���G:��!�'�~�%H�r�=J?�Ns�֔�c�����oI4����s�m�W�E�p8�|��m��1'�,*������h��
��$�Ho��	Zr��˖P��t����z�|�{�w��NJM�>�ɼ�R
��wa��D�39h��Q��hW#�b؆�����/@ ⵁ�LmJ��q����&�+�E��v������A^x��Ihh3<mP��S��Z��q.0X��X�����7��}E�m�ϴ7�ܫ�\1�14]��ξv�Ɂw~�ϭ�8�ǳ�}����-���~A���.M������KS���K)0y��st<ѹ@��C�uxf§!�{��2 ���?S�έ3��v�
l�o\KtH* ��|u:�NCn)�j"��n����3T>��.��]L�:ų��Rz�[Y��E8O����C��d���0Rd��pnǨ���D�#�AY�/ͳ��x(�Ʉ3��L�;<o邺!��`B�cuH��%l�'��\E���
����4�'Ɵs��F����L�� @<W�Aƾ{���%�K߰�r�J��<4�����@�I�b\3��'��]a��2,����SY�1s}���Ί:^�Op�����fY�I��ft� ,����6rJQܬJ��c�'~�
�.���ꌥH��x2���u��]���e�~z�	�.Kp�$��q��(����m�=Vyt�.�u��w���g4:�p>��5d�*<�x��t4��>���L����6��>p*Vu��=y8��`��|��pZr7N�Ν�|+=�C]�Ƅ�7���Zk9N:&4�5iϱ�p��#A�@,�ҥ�jY}��J��?�5gٺ4�Y����p��@H������y����5�Q�F�B����hx�mD�lb��wۻ�4�K'8�?,����\��p����d	~Қ���i����.l��D�}�]_a��vU����Hџ0�43�rޡ�<v�Vm�Ⱦ�v��yah�ߞ%�`�Ie��b�$�k��I��5�V��X��;V�I葯��� h�8�U��B�m�F�!t��,�լ��hF�u��B�G2��R~F����ԯ�D߰H�rg���\�-�NV�!�VT(_f�N�;�	�O�ß��I�tz�~�{U!�k��}��C���������W�S4(2�*���yw�+�=���NM�S�qY�Ut���)�ƭ�D�P�a�3(-F,�?�Q�w9`'�^>����펹��	�U��A� <d�yPQ�����t������h}Ψ���@�G3ꤢ远�W��ߥ�5�i�l	8��y6 &�2���Wi���P��u�$:�2Z&s�o*�}>y�~�d�>��X�/�����z�� IEp	(�,'��7)�`&�2��I�B����9B�>ߢ�wݯ]e�P~��}���|���~L�l�1�9�N�e9�:s�DZ��Y@�f��^�ޯFW_��II�G1��e�]��ۆ�����Z̉����x���Ti|ӑ<�sx[�{�Ҽ�� �y��&���1E�~��/9jϢw��~23uex��w��5�{~?؋���)�ܼ@��V�<��]�,�Qʐ�wj�qx�2l�e0�H��C���JMZ0�*n�����M���XGR�#�Z��t�>7��S鬿�`T��<L�j�5"k���E%�����/�M��y���d�+���A���@�tu:�A��&���$�VfgX�3"�ф���2W�C7����|J�o�/�����	<�/�L_�uyx�њJ�7��S�\�5c�`k�K��냁��F��}i�8�Nϔ��� Mh��RƆ����>�����_Jѣ��aHk��Y�:�ʸy)g��z$n���e�����q!C�*�˒䗛�`��+��"8�D$N�A6l/L��5?�[�ul�0k�l�yɂ�(�XDp�R�(��m���C>#���|�ӻ����)Ps�@@؈(;�x���ĺ\��02w�����v�ڣ�s��V����8y�Y?�V��A�1���Ѓ^����U�I�'ʋ�c���@tU�Di�R�;.���|/4]Iސ;�V�N���/��D�Ȅ�P���~i7:�� �h����CSl�wF��
��;H��ժUI������"���CY�D�C��LK��?K�[2{����_,Lh���ƿ�Lx4bd7���;vN�U�9؟P�� '�
�d�>�*1����ߖi�b����Ζ�	5~]b��Tt�dN���v����ɧ�B��V�P8B�xr }n�2�7�Rrb�W"z��?���_A�BƇ�^���>.�!���+4@狰��YF�Vы���*Y<ȡI�5��6$i���r�bm����l<糞N'�����E�h!�@b��[z��")����z<����Y���V�t�ԕ�M�C���!����P���uI�/ǻ
�pڬ���+��_��Ζ�$# �<�@�I���;ol!2T�P��Qҽ��#D�1�槚R�o&�͟J�= �>�Ox/����k[�]<V8nVa"a���6���}ۚ"$I�׽6̶���>���_-<ӆ�j�A�Š=;�'�cH5��j�1�:O+4N3��^ �I�w:b�(���
�rd��Hn}3�A{��B!�dV��|�j���Vso��#+��w��$�+&�#�U��[��
����9o^\[��Ʋ�Q�4�ż��#��|��Q�����}K�2��D�3�-� �iW>hެ�秺��qQAz��}�è[�s*N�Z�c�5����h��� ?��7;�q_�>ժ�z�yM�����LS%��&sG��U���ճ�h��f<���V�[ӥ����L���	���>����e��%77��S� h-}��ԁ<Zbs��$�U]��EN�47�H@�I�gCi,^O�!��`&|�]GJ�;�Qpn���M�n$�:��;��� �W���P:�y��講yP�/�o���J+ժ*N��/g���%����$�C�{��4�h�fM�l+z���_�]�''�N�E,�B�J�/�h�b��k��j���'1�Ë��'��>W{�vu�Kg�]FF�(%
���2[��q�
�����L�;!s0-B���N�7܄?�Ah��ߝ���l�J��q[�rFc���<���gl%��@	�rS qhm61N	9@�����2��c���Ad���G�h��0Qw|��YlЭ�����B}��C���`ʝ9s~0d��줌�a l��Xo4�+Nt�%4x�M�h^�q��H�ژ�pi�������ݭ��Ya ��th�~�Q�Rv���h���~����]ݹ���e/��竏Ϣ��}H�~F��ȍ[�T��.e*��=��P�=F��K#	j�kd���*��7�l�p���]�yL[FG�ZT�,,��,��u[A�~�5�G�����dB�7������_�n���dt��A�bޙ䴽�v��5(�>�EQ�(�;�u�+�7�@���*i�iJw���?��7|�-����`j �)@f�McFc�0�c��|�$�D!t���E����F��W�Mh?tCo�ד)zd�2�g���q��⍸}�JD��T岖ȃr���`Wx5�%�1�ѱ.%)d�w�j��Mf0X<��\6I�^�q�gh=rT�Y���0�i������*�m���nO��I�$4}�ׯ�;Z�`Tد���	�8@V�לr�0�F���
��SA6*�<?U�D_	`����xhvro+����� Tx]�e��Ov	�<Z\i��·֭�F-D�T�t4�!	Z� 퇟���2֐�S�� �]@�,��	etW��2v�?Xީ�2v�Wњ���툨g,�A�	��nx�[�;5W�'wT���|������kBG��N��z����XN	�O����YYޗ�k&�w�',�M,��6@���

%�8��0;�B�6��/�`�מ͜��ǷK|�gl�`�%���+S��HC����W���3� ��M㦴O�ֶ�MѦ%f5�6�CL�2�s�p���l\�J)71/���g�����g�H��ז��Ҥw�[�p���tF���=(\�!��2�s7`��sO��mT.��ko\���c��
�;�,�4��g�/�5f�Th�|i✎�B<����~���s�a溷:RQ�$�A��\F�@�r��Q�5o!�T?��?8�V҆��	uV�8m�O@����a��b|��6���m)�|Ꞛf���R�ћ7K�%mM7��NLX�]O�ٸdY7o��w�TiXf
�@��P^���Sya�݅�RnɆ��lN�#��}u�w�j�@�S�*���H8���0��x��#շN�0rp���U�Xg������gI���������A/�_��cH�¦��L��_�qF�O�za_Տ޵?���N\�3*�JW Z��[�H�<�Y$g����5�q	c�P9�S�<�nC��������af��qE��^/�)~� ��u��s �����(���P�g�sI�o��_|�%\(��-�И�A��y��J��c���Wb�.����������p���:$�SQUÂ?����*R��2S���7{�
�4?�KϦ�L��8Z9��eؼ�	ଟ�b�%�Jrb��<Z�]�9��)�9���Fv
���IY�JhQ7ӿ@���n^�MD4�p��ӟb�8��
���F��&������t��-�|�γ�?�fQF���\y���3�Sv=����!�u�4��B���9"\��r��kCݹT��ט��
��7�9��t��G�L�t�1���`>�3�LHb_q���N!����_~i�,�C9]/66�����pZؗ^H: $�s�w�1���I�t$<�H�1�΢���x�~(�ȯ /O�uۭ��[�L���l]��t� ��E�ɍ&�4�K��/��h��#�
�u���8rB^Y�Z�c��Ό'��ar�J�07dPK����ۤ+"AHV6����C��z�#0��2��Xps;���WX�XI�*��ˈL�&�W v%$Y�ƲvS�s�PҶ�M������^lc��buV�H7�4�LPiX �(��Y��t��񞜖���N?#<�8|� ��7 ��]t��Gq3����q��.�����γ�YmEV<�����i<	>���c]@�E[|O��,�`�A��8H��2'~�\Û"��!��[ �T�jqڬ�\H�@ʇ�Rg�ys9�����.�o�Z0�	!���*�/^g��b�3��>�mA���a��U>�m1I��܋�v�s�`3yFew{�j�<&�)�N�h)���rI�uhS���&�X����)��_�Z��.:�eFI���}
�6�p0:�f�+�,\��F�3$�*	�1Vh�c�S��NZ�ǾǇ�I�d(0����Za|)������y�JP�� ������_��7�9��"5�Q�ų�Z�K���*@МO)P�L�Sp�-^���I������W;��7�"�}��w�Yl7e3>X�lXe����`��0�¬l���֔�tg(+���pgE�=m�G��R�s����uX�|��E���g~�|�ܱ�K⁎:K���'D������>L=�b;����"nZ���Z	��w/]��O_�
�wO��z|�ϖ%o�$�;���J��e]C�j"4�҉,��c�)+Zy���f԰DD`��s��P��g�V(�����?|�1���\�����*/ �\�q�Ͷ�ol�������1㱶.�?f~�m(��
wa@E���]���1�o
��.�V�_{��ep�UV�]�׾�H�ǽ�Tj.�9O��h�%�ݥS���; RZk7K�_ec��K��\���^�ٞ��&�GN��r�G�2S�q�b�
Q���x`��˰G���ε�1x�����Py��>Z
ްi��ygl⦵?;UN\���u�90q��"����jq<8�Z��!D�d��
E*�������O$��ՈF�]�[�V���s�L`^i��!reݞ�h�M���Ɂ�R��F�T������f�/���A�������rg^E˲�e�|�*��-X��)����
㳌x�O��H����P��F���}��|�����d]\��}'���iAd.�'-FcV����I5�s&���=�1�L�C�R�hi����Ȁ�Q��Cjr�v�4���������d뙦�{� �!��5��QCI���K55w�"��ve��4�CT6��ЦO��Բ#v;SrP*%m}nSf�l��$D�/�� g�7mGJ�!XB�"c<���#�V��^��0�D�l�f4�r��p���(�tx��Z���c-������V2�.����K�î?�<���v��Gۗ!]�/TD}.'d����� h�* �b��r�}��p �o�%��Ğ���'�r�}O��U8�÷�vX^���ڋ*[7#��ݗ�q�6�r��Bd���	���S"�,"��D���C�OƲ���������!�u~�*��t�]z.Q��j������Â0r�+��������:�b^Tȯ�s�������8
ah*J����ҧ��/��M���3}D���������6ת�. �r�=����h~W�����b�����.��cp�z�Pe�)�-�U��v�#|�Ý!k@\��a���d���������譌�d�b�T��;�����g�.ȍ4T��Ej�&A�t�G�ڛ���:OQe;ZTY�&����b���8� �ߴ�\��\�����2���D�V��)(O֥.d�Ա�Xk|sFi� ���w�w�2��6oYy�����f*��VS*�4�2>Fw~d�ř,��E��,�Ft��4�~d��+��Y�-����	����Hʻ�09�����^���������*��ʃ22��s&��aꖲg�B�'�������A(�����O�e�I� �^�׫���Aͭ�=g�jCሆg�vbs�����O�*�]{��0��/sH�5��瑍������B�
\��%%���u�I0��>}$}š��tyz�{t$i?�/��g0��N���e�!#1E��rdG���
�T�+��.Z�5Js�na4�2LjVz���)?o#����u s�V��fRM�ǝY`�Є�5����9�-F��.IN��zR�%�CF��tfc��B�J#ݳ��m-���x�汬�{���E��>;�-�Cp�8�_=��Owb�! c6���r_.��G­��X�������a�z�3K�K/���?���!E�#�'h�����R����ORu��"7L�N\y�@�t�ij�1X�9ge���@;�@U[^v�-#��O|�������ZL롞\�XV7 ��h�'��Ĝ�+ZXP��%2�y�����@2흣@�s,6yP�M%+)�0f�͎�v��vqZ&Ձ��NI�C,u�i�5:��H*�RV�U�~�O$l��&��S{݇�>@��+C�Ur$�	9�q,K�q��c�CȘ���d�,�:���?��}�.co����d=��{�I�KMZo.9D�
�|~4�R�5�������I���bLT�ݐ�0�8V_��n��t/�h�R�{���W)��|6E�r
Jk�l��]��ed��k��e&�FS�K�ï��bb�9��f3��|��C~�,_���|��e@�8�S���s�ҝ�"��ْ�y+}����Qp��[���9�U'����I�	ye��5_��,�N6x�2|y�d��L�#z<3�]��Bo�������|��Q��2�Op�>�XP������{�^�[W�Jِ��w��,�E��<�hIY��p�_fb.�$o1�6�.m���C��6i�E�,���i�ESBN���6�x��C,����N��ꑝÉlu�]�����/�]����uR�F��]�4���8O�!jG7!���3��צcai��Lu��\Hq
bN�$��_'	Z(ZC\vm��}�T�-��ǀ�� �V�9S�o?�����?A��{J��D�L��7ꄮ-���-�$q�����<J�$$�� c�@f:};�\��1�6��ÿ/�
1���2Z��a�2g����7�P�7�ѺKv����A�R�UI���b�6��e��������R�%Qdw囉���~\�2Fk����&c	�e��L;K�:���N���Z������14�*Py��!7�N��ȼ������F�3�
\ߙխ���n?��s5uP��7��-�a`��P�jZ���M1�8��@��@H�;���ﻮR�9��ӛ*�ģ�������C�/��ռLn�'U��(r�=*/w4�����L�� �1k��#���/�2�fs��͔x��i�[+�冼��XV�2M�Fɮ�$��:7�ǔǟ6�<+��vv%^ZN՝�m��N�	�����S�Ȋ'��wW��*�ٚ	[��I_��X�)����Cт3Qy�K���ovQ�ncN�����b�4�݉]A�j�M�#�ؓ+l�轢�)I�C�2L�$��5m��e���9������B�o�F�S�? �s~e� �"Q)�̞��:5f��%�I��a�&���:���\aS���v��] �|��~tю��sԾ��J�����I�����UN�ӥ�k\�/��0�S},��m���g.�S%7��®���ى�0R]SQ�c�������U�9t_�r�|zy[s)���𦖴ٻ!�<S�i�Z�q�%i����/!ʺ�C��_��oE�y���j��÷�
���5��}ӗ�5�?[�"f���.<�r~�E���n�_)���Qa�5�����`��X��oJ�L����<j[a��P����*�:�	�,V�(�GσkCH����*P�N@�b�F�C8��[a��T�c�?�گv���	�V}��; ��w`~@3���|ŧ���b>cT��|+�i,��̯��aċs�����t�}�j}	��gZcin�As������i���ߏc6��)� $>��;ބ$�w���a*l[ꄕ�
}��:Ҧ�y.���(�t'�{��:Zx�\fM�%>���D����ɥ�)��w^;K9̨Z�%�imK�Z�mS� ����_�\����N��9�*m��1����t���,G�(��i=i�9�4�4l_u�6^���6i�oa��Zs�&-����HR��w���q��k���f����i���O�Ɏ�-z�f�˖�.��#\�{���O�L$��'�w+��6�f��j�&�6W:�*�ʚф5�/�q��+���-Z��t�y+�cp9fU�<Ƽdw�4���U�oW������Ϟl>��%�=��� ��`�`?�B֠�����s7�XÒ��n��ova�!��2m����a�b%�؂��h�<�ׯ�L�V�J
�Ě��1f�Od�E�ʩ��l���G�;Du�Θ� �f�Վ��跺��C=;��C� �����w�ٶ+I���p5Lܨ��q�����,�[y���̌@�+��C�{)���ɕڴWUP���e�]�7z^@ثy/r�g6pd�K���ȇG�e�;�btVy!a
wP���>ש�S�S{�M��ŷ>��N1�7E����"�L������yZ�<�b�^)�:r�f^�w�ҦX��q���p���.>��=wƺĻxE�@-CD8�ӶgI1����Fb�!�Q�5�r�V��Fu���h����P���?m�V9�TK�J�,D���\ ���{������1p&��Zu{�)Mt!�OH8`��c^ 5\��z�IVo��T�� �(3�};���k�;<�37��c���8�F�m����W1mV4��h|Ϝ�;~�I1��k�VR$���C�5{"�cTjc�DiK����6��`)`,T��4��|�,<7���k����=��?{�>������)/|���#�3��p��r=u���Ҟ��tQ�qE������	{�������j��&���&�?֮r��]At\���H�t����\�����=��f|X*�b1��Λ��b���y�],�=Wӟ�eʚ��I\aݽ*��w��J,o�Мj��(� ��~����y>�2�q���	#jngr/EM��;����k�����ݼrC?�vbZ�F�[�E3�0�0�$�ً_*���� "_���d���h
ܝ��=�V�Xb��J>����gƐ���|�	i����4߄by��A)�T��l����Doȡ�f'2�'���#�Øri� n�5o���\*�)�bj�̳�$Z�0߬�!�6ka}���ui�r$]��'��<@筏U	3��'n)��L5�6��>���a��ġ/�rٚ�oae(F�hZ�ۅ�G��4���N"�|kO��
P�a�-"��t��La��*����/�mݰ/�z'�*En���i/�VʨE=��וU-:�uϚ��U6������ޚq�l-is�p��R����Y2]y�Iı�3Q��6����G�_5��FC��J�r��r+�=�RZDZ��&ϙ��8�u�E��g2�8Oҩ�o�i�@�p.h��9����GmY����f�[q����|ע4���a����i��t�Dhc殒#�,�b�|�j�
q��g��P���������T��+3�&Rf#w�i�O�'*�����:�ur�ɪe�j=�Y�7��`}C��Y~�/��JJn�j<��B�p�4N3FP �< ���\0u���n������Z���w��G_���"��{��W��q���5��$�
]CtXxS�tWZ׎*N�=M��~���$�Sui�<�)�[F��q�Q'P����/o`�R�vY�*�aE��?`���p% � �
�\b\����	s��o�����""w,N��r�^���t���{b����M��W���G���0?��ɘR���#�������S�c�r��Ws��
�wx,ފ`�ΙR%�M����FBC����_Pf�Au5��0
q'?���\0DƏuJ��FG�|�D����"Z�V�x�u����^c̡;�!��#��1���9����S=?���Up���Q@3#�,�� ��7�l�
��C,v; ��k��a�q婋��-�0V���6�˸%i��Ѭy.� YIkvP�⚒���n�g��)��K�A̾��k�04H=!6Qb5�H���i��
��y�e� �΢�m�$0sBr[g�7;�%983����91��s5�E�0����:��H�WX�uN�\g��������Bt�����/��"^֦VbPe�(o�+&��G7a7
ʨ�
�bG�j2��ǭ���T�lq3A�G�"'����\�=lgy��x"�8�.����N�v:u'^��L�c�.*�jo�{
0�O"ї��b6H�k2�%��Խ-K�b�~����u���[z�9���Ko���*!b���]��6�y���q8Y{���ͺw|jMo�	$[ZUabđu�{WE�P�E��|���j�j�P��X't�⃙vӆ�P̓��N0�eCo,�r'�hʾE��/s�T7#���@ �Z��d	�l�8��U���%?��QD ��{�]H���R!Tw�h�3s�,l��l쏮�]v.l,eO%��w�a�����KÈ�S�y�v�À���&p"?̵_�k�����c'/���{#B|��b�Ň|�nu/�-v��O�[�*Ё���H�2-1 ���OG�3ûѓ����j'�y��yt>�K�r^Sin,4���l�V��H^�Ry%s��7߽qN��a�1�O�u+x~�PHA=³�ϕ���e��A�\�vF����4wb�L��Mߍ�����X`�Z@��	�J�s�S�\����zp���p��Q��_��f*�h��w�tb�HG�.��V�Z��䜰�w�`H��+��۠�O���5L�d·[d�����Y�{��N!Oie�=q^s������E��*�qH�U��g.I<�nd��f��:�9EHN>h,�R%����U9˃��Ԍ���O��������&�2�L$7�:�� Ӊ��1��%+f*���wE�^<��*�Q��~��O��!�Q�!Q����+c��]����1b6��N�5L���/*$H���
4!u��f:����dهH�#RPQ�0SΕr�Ki`T��h|�� �?����Wv+�*��x�)u���$n�M�n�-)�o��!�P�G������Q ���_���f � C>SN�F�+/���Z�N����(�C�V �`-�j�������� ��8�|W��sZ����o���0.(�*��؝稍JI m�%W�B�łٳw�#���%8�i�*��=�%��όJ(ĠbQb�I�<�x�_x��F��1��|�8�Ph�0U��Z]w�*'�$�-Y�{�=�~Ғ�Z���2ύ��4���4��c|뉋䰿��E�O ƺ3o���O�(�m�P��Kş���? -^�Hv[��WX�2�����Μ=w��%��3�}!�?r�N]�½�%ޓ�)!t�o;��Y0�Ϊ�<m�߂��I�S��j�7��U��A�����^I�4!�)�m�uv�l��z��ɢ���DpT�P���^��p!DY��4o�(о,=��Kd�Y��Vȯv�V���J�,p�W$k�[G�5{��(�&S��h�����6q�w}��G� hh� E�s��f+�#�%��S��I�m�c�����g�{��C�j�-x������i��4��uW��{�#vB���<X�xp$�~n� F�5�tۤ��&g�zwC�q�Q�Y+̸i��j��=r��j������f�Є�}�s��C=^��{:��#�a<��g����R��V{gA�ƒT���5���p� .'�m�WY0DI�"��W���z�/���]�\��O���-BL�oP�`��(.�y�A/�Q8�Z!Ҝy*!�
�` y��a>i�v!\k���WC��	��!�?~tL �Tcr>6&˒q�#>�,{a���*�B�M�d��r�V����ɧ�{4D��e����5$X�r!EH}���g�o����O�u@^��Oᗣ�!�����e���. W�M\2J'X�}��P�GD�oU�� l�m��kngF	��ލvM���-4�%�I�T�\��OEo�i2%Q�pY20�C� h���*��ҋ�����%"��J���!�h.����7z1Ɉe��cM�(��KX8O+�M(��Z�%��T�-���k���v���A��$v�m���Hu�*�K�8	C:W�Y�Ϲ�.�<;9�L%��X�w>�,����C���کM��g�5�r(�\U�[:k��|��<dj�ֿ_�Ev���+�������˨u��dB��Y�K:�Ej��ſ�
?S�������9�_X	�?u���92�Vj��@���w�%O}m�:���al�\��|Qp��(���Զ��]%�PW�c�����.�G~.CW 5N���<nr��\��5�
�!��1P�96�v��[�z��cf��(�"�I�כ�c�ǉ^?I=(���I���'s�;�ak������
h2`PG�����{u����B�������Yj��]��.ã9XP��6R���p�������Ba�/;甜��Z­\5��������-.E�r�'�y����� �ǁp�^}��Q(�Q���h�=/��[o��M-欞�br(+��	�xXE�AB�\05��x���?��<Rj�x���=��