// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:22 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sI4VqHn2WIb6AZF6xOxNKJMNPGnDMJDFZlDVjtZBboACzIitnM9yKWZ3fWdJdUbv
V8QVbmoO1cH7zN9DRSsiU+X0sk5BLwQKUiHBMwC25cr7Sc6pG/qeykspzhGiDPZ0
Quyu9yA8sYMBfXURDbBllRYChZc6v/yq2xvS0Ik0xOk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9168)
tZjsEjVjTVCfFz2FxH0Vazu584sx5M/EcIPqEqIset5IP9l64csXDL9UvGZfHJvL
D3V3Q4t0ROf5S6S9sZIKohZtYQUgyM5pO3ADETaNnsHyFutRgjrQTCeOoe4PRO30
jjSwC04pl78REKiJX5lvCpD00ZdCydSMik9NjrZiCUD/04MhHYsgE26kSx8hr+z7
gL6mL4TptgFdO+Yvvi4DfwN2/RNETAjCt5es32+eaLoNautDYH3xX2Cx3muKIkvL
ue240RAl80uBHTvh7r0L9Yf1tSK3ncj488Xj5n50TrPRVSxJtdbtzlQUzaIHHmmD
K340zOT106tzORxakBcpocPOJSUNkLX0yrEf+22WIbtOiD3kd2+MdN4uAnOL+1TL
dUNRxJXks1/tp98PL/78OzhcVuRcSRLqrof+l/clPhx8o9dBNLbo1GD+UFF6f6TQ
CIbBQtD3kuADkz69OM2vxME8lA4x3mceKFz5ogXuX0X7IUk4JzYfQglTzIT4Hi8q
UbKkTWm2mR4DMPRSTc2T+eWm6Aujv7UKnsnL+c2FcwmmvFnWIv+O5PFZrtObjOqF
cavK1EkzcCTZIdijb7NiardKJsC9WTe51hPGHe6tekm7iaqwtA+Y791uja6GETuj
um/DedoBlLy674PRhYEMvV4aK+1WOD3OIGDwlOJr40R58HVG1je1UaPbexM9sc+g
AHytLUtwACgrVkZbxQ2iQTZyULrdb0qIT6fFwJgZV7mKkhvhOpNXiX97LPp18prO
3d+xJAu8X/CHqDhSu9Ygzc2kmcTGtEssCAOtNhwJoIqsUo2NAJOhJTY4SL0rzTQ/
itrCAxUqsnTd08A1affLws6HvxbHIylGKxmWZnom7WK2+sn9EWy3qM8sh/v7pXP4
ULefNYLcS9VN3aYgJxVISgFaIcNRK+R9juqAfjNrE5zrLrD3KW1LKH33DurQ7of9
2kG4uod1JOkEdjvKZ0yrXjaJ1xoOhYb9YYH7aO3z220+oHo/2cymCR65cqT+OAq3
t3O6sgSrMJsrkwZzutR7fD+r20SyDJIEmoQLwDY5F8xDFeyUPo7X4BwXPEggwvRf
8OZxCUD+m5uwtBgvYG8V24B3COogrgy2LJAq1nLJS7AZm8h9Za2GIAj4tdlqHE0e
fupUa/sjjBT1EzcquBHTdnurWAm7s1q+UT0PuI3zl5YzaVNy6EKB4HlzWG2EeusH
2TJbmwKrBnAFCuGlvwONut6dOcHq+49Eem0atPHCrx4LgwbCi0kBOGaNu4iy7UYi
21D2F2Ru7GaBFKaQzg/YivfgEBuX7NOl6tPL+pPRTkE6gfhiLyR+/FX3DLwcmtOU
UkVEg25H/MN6OTT8Etl7CJKAOv6n9paYA1/8yCkI74mD/1kZvD8fY4v3HpiwRmBW
esJACe/DLXlBZ+G8rjUUShYcMiOp1YE/Lh47RevwtDqAiZaEnNslf1KK9ZZRiP5B
CMUhZm2HDKhEgQ9GxBF+ksm2alni5L6bK0mZaFDJcEypYsOCncbTwrW9fQOLyGpj
c6RNKKXRn5iaJ1fK4AEY4uQt0eOkXT4ihxIjFYUO9aArS8AsVMkmnOQVof9nTcbg
5pavhx0dmVKl+MAueMezrp9R41p7s4WFi9Fi5jW0MmgBlHMZrMj6H+4Cs/Pgt2Rm
9/RxZ1c6n9MXVQgxZIJLfe7zqX6kTIqXR5RPuVNNV6oQU0Z3TL9nrczjrbF2og5Y
VFvXZ4RntGvc1qpXuMpOrnzfdyu/hsYLaeg84do7fDtR8qeylizFFVs+HOCH28o6
RLF6y4S78F4+xwoSfUWx45AJqNLdjXbub0VZx/w98VYq25NNKpiKwsGD91VLBWGS
8ZTu4/Vf9pAmeF+3yNgozedKgw2kS2e1ntfOxKd2luOe88Gbm/lNuknMtJu5QxVM
pSM0NJH9uFBgXz9+e3YCXC5sa0zQFtAlINXWOz3mbcEZYzG+AfYlKPZLQ0c9S6Ya
hUgsFw0IE6Dd4yCJezuRhMmdP+aZ+kZbvNefazgWxRTDIeVaDlzx8LpRcH6/9jUT
r5a3HmmYkeKjtWOr7/c5bavbbTsAlS6Bcpkzg6BNHwZ2MswhILTjqER1agVpzi+I
t8HW8GfaQYXkpgKZBcYgHxl4TMV5BheSGBG+S0e37HNKIb+Uqn4q2DhmyoLFp9tD
N86bXXtPbWbiEajXYqvXAkSUJc+lvWkE6a+7MSVPon/avfoNbBiX4b2LEd7HZdna
PfyRO0V2OqddTfg9XXtqJ0VuwGJyJlHpljcJtVf0vWA+H6hl8OY7nV9JPY3Vr2s/
wg50st/B+G0g3ntikoqZxXl1SbGVf3G1hvwSk4ZX4gJ0LSEmGkk6P4cuv6zNyQXT
+/UiLL2Aa4fgv754DUjfV7qtOUxKQPQUv20aqBXxPYZZe8kF/TYjiDGijTIMFGXz
j+gV0CKSpxJb2Qx9VqZL3/6hqWFmz+Tkz9xC19h/vPSkClDtPvXXUB1zcZ+D4ryg
buwL7AU9JvKryNP1IhdlP+vxiptkn0tRgyA3jW+a3gldek1ZrjTvEjRv7Br6XGI0
vwA5M3ORQ9X/XIW6+u9fr9L/0phNXVIyx/uwsXszahTZgve9Xyc4BnRZww/CwXAB
dBORDYL5j/lvCRR0U6r45ZiVyDOii0doDcAyXC0h+1ptUa8t5YqCqoHkNFD4IZVp
w/3tbwCuO7BD/BmA4KVVCjq4rEnXgu0bnndDf4CDmOxSRs3EKPVUV2RYwCgI4dno
cOFvH42RMliWHY0jbdTNL3tXYZkbQaJ/iwBX70YofN/G6VZaO3tixKSFQtzZtVMN
vfTuxqaiZ67f7uO3PBsswm6oAyRmPpbIPTBPKFnqoTuCvwqoLMYL6qpUZuGPFde9
YEoPR838Vj+YXKCAZ9jIWUS4nNygPKYViJXwwg0StgO/pvEX6qA6U4zvZsBam3SP
SRnn8qEKCfa2SNALtnZXyD/ZPRamF1b/0Hp/7x9fRrTzT6+f06/joYjzxbF4mdrd
Eg30N2i+TU9HmrPpOf6CbtiY7TJ6Qu8Qq6rk4SKYI24JI3aNSykvYwDka59itycU
xzqYoc1PPSN7GHF4Syyab/7n0vV3SjEc0UsJ3TQqVubHWoUtBPxnl3DfVxz1mFEv
6mjuseaMqBsgFc+65Q8/RuVu7y0DToQNINXKcfCIIkKkLx1bNz4JvZyUP/L23q/O
Aim2oZJRO0id6Yx1yc8Y2Z3Pp2E4wnTI2C3+w9cfJQtufhzp2JZ9RVggLOR14Y+t
3jZJoSf9vC+gVnHXxtNDb8CbLj3Kz2L18Shie1a9vMsaJqcL1DdC8y/tgx706MKn
mBKkI4HjHEgKn8lBZmIHa7NIq9tCK5s+gu0T/PEAs1OCuNsSedX9wwVctcoZHSHe
Ou13PF6b/0p0f1hg0igHBH4NjniVG5VWB1+DIAcaOEazQPaOUnlUwT6wYS+rgCa8
abnTO+k0nnTm2dMYHICFmbGE58PvSm3ZcOpu6Gzo0X2arcnuRrZE55m8QIp/OBG8
LuWa1gF2T7wLEoNiX6tCMDkTubD/pkpRkcV7ewXcGFhZaYeKj/RzTODdOsgzAxiB
UF+rHBYXjfRviO1ZFx/6wwqc3dX169bPuXnRriAfrmODRVpj4/lO94s9oDCaURbC
Ri9CyMliEV2DfuNKsK0S4OBf+0zFg1+vhb55SMNc77tSvcSwEyqKfrzf8EruWDmm
+eo3Qk1gQk68koj279boGmmYS6uXpkxjSW3PwnJKQaT3dFaw6z6onIXT7ey88TnP
KIHQTOZSldaulOWPkVtMAVY2bKoYRIheu1lUCSpXZxI6Xb4ajxLew/4xBSyB0eDx
msM00YjHmC/+hGxz8lMYwgoLl8HlyMJyzEVWqdtWX10Bnq2C3QEzg3bn7E4UCBjn
We/uiqZFwYIPunSgxAl9lIdfNWNb7aQO0smBVK4z/aRED1J8STqle6/zSL2X3T4a
Zm6TkyW40ag6CKxkP1X7mQ6ttevjdQXRO+3fhd32KldYrKWTEX1C5M7PAgZQA4yE
MbBw1iGw959KPBw8NdPvjBUPJtIZLcDybgh0nmSe2De7uGP6EJMJkKIrdfxdiBt5
Ztw0fPPCK9ZqozMpsLdi3959qj/gky9ilnlRPDzmpI2jska3T9u0HCFtc9JghTZ8
A+v0vOpIe4lQMDfbeUAqO+T2YtDqC3xrLVCr7zr+HYSAy7GlECLTMxua8t3oIN9W
qLhYR9RKRq7MuBy9dTivm4zMGEB/T0DBonttXE40vYe1XBmozZAv+S8ioTmuOzXO
rN0k+Vms1/9La/+PVc7RpBdNWo9AKcr2P1qXBIu66YIqE2FFSVGcZt0cm9iRrGIJ
m68upowyhf3xbLGseRF3PCVnoFEZuPGGESACOHoLblgKVLlwZFSz5c2kzoVvwEIt
DjCOgX1jixgvEfS9utdxa8A0FZsasTxUwJ4/HokLqukU6BozZ4NCWiIUxtT8RQ/x
QDWlQ3SaUZ7WrTqhdGk+ha6jevZOEhfuv+fWpq7UIejDfzrTztV3A8PXMFrkiopJ
MfBK4Fk7TWiDLmMOD1Tjjmrw+fKJlTSeyENO2q+/7KMnZ6nFY3PoBOhxlhlmuHAi
0otgO4Zd1H3X4dyPZSMV0LDyzy7KdrNH9GiwQ8YvYDhnr0az+Q6972rGLAYDQUjn
sReY3HqTyvY2P2v618q8rv0R6bMAg4qqomy876b1kclDRlpHJNniNpJch5VjOrly
fe1/nX2AhA3wwcjYCy7Jb+LONR1V3xK1I0CRrtWt0a3fCe0P4UB1TASlZUNF3H4m
GiMOyjcSolhpCXeH9IQHFQRWmR1Svy3ulgFms+9J8R9T1eRlWHJ/44C5Y9l0VWvb
1s6I4h+X3lRmSKuw1lHKNMs6nZIoO6cao37KY20UvRECiRqhEauL6/NJUIbhkVPh
V6p8JOHGzoRijgE9LTLOqGHNjlh7ujJ+WvChjNsg9XohgQ7FWq3uNKfUjgxqsEz5
rWfhAiWia5wZYEU2RuoJd5Al9Zm9GECTG2jS8rGjJSz5tSR8pjfpq+EysW2SHmw9
FPP2J1q7sS3AP3Ag6dHkF5+0P2qBCiSgmR0Y4n+zG6lkagT/J/L09Ow1nS51QLwP
2q6ahkP9Sai0S7dtSsv0XqWL5coaqz9hRhPfAOXaa02Nw9jw5tPAmK3ofowONPpN
KSWWjnEqRJ5ec3JpA0L/Ds4f4nprmzeVJvHGIOTBWwZiXzgcFtggn6fpjRhHuiua
DKCSFu6+4EAJSdQMEF9DI6tQTkgOe7A5RI91ygP9/gY2VXXGbmUpCzVymV67l+Re
GIhq04ari+OAXvo8i8OX1Gh7PPU6maKIvpQVJd5SOMJ+Z+U4Qa5by4zvEYi2wCEA
1/CxOVcPwXnrOQ83RdA/eJ7Wh8XIqThS617bDcqIkFZnQyWNNDQF3OTMJmT/ANqx
PZSxFU9mN3/ILSarsGPb2udmcYPt2jFXPglf7ucozNtGChizz/1pb/sLdAS9BSWc
GDevASzVz1BfQQe7cC/Io02AwDvA3YEWsQl/bzK+bAoy7qisT/mrj3CBLDqkVBuI
qfNPEYeWBYAJ++E/jQZL6qcAfsHRMukIWTm06+aMO20pyWFdE3x156jzys444/6U
yE8rT3T6NvZKN5ddb1Ouu1IpG/7hPSvfVOX76NAe/0SpbeXxZR9FPfD0zV0x5tCR
RyI3DJ4h2IEKrJJUKeyuz/w9uATofBUzHeF5BUi4XxhcA/V4o0ewbeL+z4cayC0q
SXGbZXoXcXiXwkrOjCWGwx7XJE2IAWFnkahbA1W854t4IlHdLAXxSinoJVHKQTN/
Ia8LR1NJb/SZ6pIV0AtKQNM9exgzP8mXaJUeXKcOd9oUs8yzOmw5bsHofKXKXz6R
zgjUe0svOfGoW1rf393c+RIOH1DFMZEDLb4MqvX6i5FYfTPSb3f2vn+EgsJc9DHz
vxwq4WUg66X4U04DY/3wHdiBqGnvCu9X5NNWJU6h/GkeFXFD/nXFdDzJejTBFKFr
qn33JvmDh4wpjCYHnH1irfoL3QiXUv/Lb1WKY+xuxsRzYk9RdYQSmfhfRpOnmVd8
Wa3UgIF7w8W5FVl+2BQhEAOzCmifP96OJ0YZkm0l+IVQ+mQeV62ZbHPw3DQNJQxJ
9f77VYcklLYhJbBK29IBv1BceqAG5c0iS7hyaHhTXQ9Vw7s2LYOZOoyIMzzrj4S6
56CJt9uokzclVBsewpv7TbpCLmnZdIwqniWpgibK3O9ZEU91FLchX/MqVWNscC6g
N/ArGpEz1u8wPCuze49UGVM88oU/42ZXXUn/qvtSGLDGPlNIxJqARBUUlm/IFdPT
9M8eDFnkfNoVRuuvu4U3tB0awifDvdAOqYEkD44FxEPVafMGBsqvaaaHA4pWXz17
5V+5EPZgvErjTKeg2TwF7M7WdOx32H8CAuSbZwxB772E66A0eTZpE00eabmFrE68
X6vYW3AJkDLqP7K67ZAngWAaFoxb3gs4qyNxQlXHPQnQFUyIqmBvOrgaf69NeWLA
7RwRY6ut+sWNKhwqwr6BPHiVN2bj7TpdBZ/gx48q0bE4sMCryXaMnDsYo46LRYNY
eTJzFIcwTzC4yD7uAI3Yi0UgctoWFFLF3HZ1vvt+p3Ay+g17iwB7jWqOAD5pfxnb
cV86RrpuDwBhYnHGEkFcZfAWDjOr/KIxt1qSgdcdh69q3sJwAFzzW+mGG4gj6P62
yuaVZLNYNmTOJlAN4Zr262el71QOLSltVMdq7wV6kHuuedo7UcnmtjQzH7/N2Uzz
uxgSLyWxfDN/bV/ue/TZfVm2QUtL9Xmf8dRPL3rTGszip6O54/wXtS76rsKYTX5z
GMi9/M9nOaxwD7cSl/ay1s8myuY+uepZHxGnVAU7JNMsgMloaf/Unq3uL9zjUqYf
gM1U96xrQ/AY3b1Zn43riM2YlpDeFCU/j31AQsPztWPUWmgCm7GYAwGSsxzASgLi
RbKFzmTR1vgBljWr2KRdzTP5JYi8ZnV1RKSvAL618Qz65NcO/K3WstuuL5ACadYM
QFU3jlx9qHwzlq51J1lPreXQnLjPZgQ9yWMw2q4oKsXh0tiD4afJYxqBgAP9nO4a
UyXlkLUG7jZPT8EXJiTZSRoLgsu2Z5BCXA1HnsnWD6smH0L9Mt+jfdZP0igBx8i6
HJO4L//SPGHf+dh8s+K02uDPR3fgg/j1ZqHuh7W9Uq1Q7u3UH36Mtw/Fsib758TY
EXBnislvfeNbbJScb2xtUwdo3jtRdoL6Qf/a4PF2AjM2+JqwGvEsmUlXzliV9FsI
yPGbMog5VT6O7plfZuU+M5onQ0ti3PM8vRy26tbmdCWGxrtJ7ytzC14Z5FHvw/I8
IDsbuiIx+mT2z7zjnza9N2P5AOMi3NvbBUQ56Ctp9fUx9kTtjDkd8cMDihVMtKxY
t74wr8MNCmVR75DkZPtsRZw1pSW0BqDfVkxwaBgy37IGvCtasaDHXFrBRlL36+zY
rgAN6th/Y0VWInK3EPF8k5kI2R+yZ/zz8aXukeeEAwircBKql9nMHOFngPkbRxJr
10qEWw2if4C/vESFR0wKPLjq4s5cHxFHh0HCKT/8IijBN6cfFbxcmJrNt+TdHuIA
ICFu8vbzr8q+3X+yrlALa1NaSLEas6nhuekn71yN7K+Xh1T8f4VDJYPszO+y2XGZ
/0kIWBFkAoYwQZZCn2DybYTFQNFeeneKiNoffp5f1vPhpE99EQ2ATDifRfjoeYvy
VOnE/Sgn3tfbKTV2UAVh2dyyHKrOnoKpjYh59VJ4vj23U8xnLJk707Ne2PJJ0Zvc
3lRMNnsYC2tLlnhYijHFV3vK007JPUrFBiDIGtNtkkiAAVA/PTFwUDWCipMj/WFp
iatl+rVwPTc6wUzuIAbRziYpE9Ha4yLoELlnSoVjTVnP5FAn/hJjt8I1copSI41R
uJyI0qOUoKLR4qUy21FbVa7r7nXkZQryphzeR33JxmNvialdXFwjTxHRu1NJZGuR
5GtRkzmQrQIq39PYohcmBDWWedHeBd1OPFizfmV3gDdM0JsciOHwxPHetcyKW9aH
R5SfxAtoDHzJrIDWRWm4JX80qoc+tOyRFONyU93ezRiIROmCZKNwQMgIhPoGRzJy
0Um41OFCh5S2YYI5XNusWl2dAwmMWMjsz9Coiq50UUTPTj3Rk6C1e5wOhdw2Efo+
1+rdHZCmNHH0Y99ka6Qgtf/vzczYZb5qx1ey3b6Pvza32KBne5pWKPp1oO02x7yZ
fT7tVSy0ugxDf6hp3o+R8peCgpPIrnzSPZtLtaYX7SKLTw50RregYDIbuZuATkMp
a+daFF5PTENdlqcugHTd1e9uTw3Ggrv6u5NF6xZZYQbNxAwmcFNsydu272lTOGBP
5gJgc7D94Z8I5QXi09l3xHbowwSPPQxk+YyM5of25plUlf8Us0FYyZtcKiNcoQcB
XaUIBK67gew8pwAfklSUfjZz8+ZyYoonpIW85WvaQMKYU4H2JTQNhsdbsRo9NRy3
oFmSqa2CYHINYj55PP7lVAuOhrTZi2izbEs3wfpr1CDZhgx3O7+YL8e5GCC7/lkJ
rtTZhtI90lRLBJNRhDtY0JDXv4dipeB+dENVTUw57ZyaznuzTVe1HaSNm6mzW+Ac
wVrx2Pxvu1pRO+rF/yG9GwsfvMDGtoiGHtC48zSyhpOte/7R+SpfH2ECE1orO2hL
W4zDD4YDTZeV/LnjW9Tfkgn28soaFbuLaf6V7vHIVBa6YDzWao3DmUsefWkzOawm
28oMf93kgLBMgLAHQOBuXfui/3p+GoBH1JAdptIVGIiap+XsEmjArN2R2LdHPSW8
0okiZQdzClfB3HWR9zM6kCG5y3p6H6BElVJDmNXZKzKL3NhxIvapcZg2CjrxN0Qe
s05QvFBeZaiGeVqXG5gwECD3lfnpA2nhVeHSikOJmDhI9xHSzpXHsNM4CvOIZEvJ
KfbD0AtwFVQQml5xGTZ8ZAF8fRswKYkL1xGpmbtVFSBVgEfFLcqU2ybOOoySpyW1
WAAR5C2Xx7KhEbZWpFYrzXb6egwiSyFprUsO1kpfXx+lzF3rKoOB1wENPQxmEn60
Dxxnluev8V526PlKmqqgxk8KZJ1r3MtoP95fZn4ghG1hztQx/1zx8RO6bF+rQ38M
O0Tnp4vwUW+rcgilVScUwVzFko5lz2fmoJ254aySAi6m1dtktivZ6MaccYQYd/cC
UZZ/lZEQgoZTvka9O4BURLwCKUBp4XS/cGEzJRoOAHeVjXfrhgr+SjxHfAYFOjwX
6sLgZICcAiMeuElTBc0C4hVtD0jtd64Ouq09sfjnE4zUXWBJ+OiSZbTJsKI5kt3a
T1sF9tg53EDh5OyNxuneYOsvF5Ws33PW5PV+KcxP0MzPUPsvovuIejFSra34M2H1
5JHyaf0n+5VY2Hc3WK8E2dy4eMID6mnFLFuL+yGXdbOZetpuEgGFrc/7LLBjQ9aQ
CBrywoI8mL3Nn8/CFz2MhxYJj8cR1iW/qsytZSS5XxcW2uOhYKt+H+v/9Ki4/XyI
oE3M8rNcGfUWbxSGoii765D6Wxax+yCReZC776k7gOFOY1eVm/Dnl+9ki8OXWzYE
AjfRKuLwsP+ztkVFhvuHglIDRCv3XGaFu66b9hlwXFRiQnmtDrjIqAVMpLhb47Y2
9i04xd7CfxvYWzCYFbnr18MCiHVXmIanXOYprmIGpF2vKAieSgPDTPH/5QATapZa
Nj87J/83QPWSf7hIZIvnUF8lSUqKdASiONlWhEfzwjhmlfgehpOa+jAto3YqvF2x
t1MNtPGz4F1ANvmsLgnJjTzTZjP5ohQz25kxOybrnM5zgEjFPl1YV8Hh1f4TTjFo
xOmXMAgBcmB87GoByeY3H6pG+2qmzf4Gyc2JJ2L3+TFypQgQLqjFo7u7gygSB5g9
vF/U2iul/4kvKTBjDCugQqo3zY0lbUJ3Yzcf+fjOu7GYfMzDVhfoT3itM/LbSJnJ
HRZ7xmNshCZ1mwjo/fzn983fYMDep2KPE+5aCZBft2PSWaa2+raR3rBDH9szEqX7
NTSocRVIdoqGYTeu7uGYj920XLkBMhdgs3X0VLEv8wWqFFSRAkcsOzXzOLJiFu5L
uSqUIu7zNTbfmRJWRzL81wPU3KXRVQSwsiBE0b+fXybaG29a2h5AOcGqff/4DTad
Dp9B4Jwn7LmVWowFVfuRumcP1Yi6ZE0BcAOnfSkw8Ji+5eOnwT0U+v3AIX3sRIzN
eQYjfAu1JPHIzVmZTBd8xKHoP2LIc6g7OuyeurFVXzRBh6BPxfVx7C6NhLXUG8z3
mLxzkoncBDhOwXlrS+Ns3UqrVzRCn0dMH37aiYd92DieMQ9n3fd4AtEGBiL7rUeH
ZwasEhWA/M2so4mlcfM07DZZDkhpug6v5VwZY6OzHtdj5AnpwuB+0Mi8EU8882gg
nwclaDIvDtUZpa5hjWfCjj+Z9UtToqkg88Z2YEZibKGrEULVH+kQM0BxVRphDcpm
nY8ONT3gTGFlWxfuTEGw3VczUUY+zsRXJkS6W3nFMm6ymxYZmWu6nIC1f2hyhPmA
uSVUgI4fUJcSmtxWL3fSoWG0BHxBDZL6YtoElFoURbA/GhseR881oqt+0YbH5hnA
yx9X4EtcZkxWJEypxw3NXWXZ8FdldA9Uo4v3sLTxpg/GyKToEL8qezmxsVxb/Ri3
R+j9lydlPA/lkYm3Y2oLx3zS5orKSlB/G+l0bG1sBoKt/5/hpHWFXfrxOCCdrOgh
jgBxeREQbIWFTESD0E+4Q6jG0vR1120gcWDImvRqvfo8G/c1lqe34XOpbFsI3/bb
LP80jRuj47Q4snA8g0CGjVRMbtw6NfzSpoQfQjuRF56E7n1xuK4E0mQUr6FX+tDO
yEy21bdHsLe+CEBcKHAxTGePHlmhnNctcDbdv3OtafIyh3GduzPTMJUMM7pOIRTX
/OHYSnKidxjOhm+KILItQ6OFrpw7D2E3dvxSJ1KEFgP40oQBDnhqc7d0vJ8bDFWA
djQiwpJzi24HKibKf50rs8Cy4abJNiB11A5+a76uOMQN+358F262heTcalE7qvUv
Xf7GmoEge2R4yQWgXVfK+M0kuEID4iR0uCozMrnWY5Gz2ts9cEco9P31zjsXZBJY
9VQHwRxtTp5Gvw07aEoUO4WC1xUogS8R4GxjSzySg+h6cskgE83R2AVpHwy2HO1Y
LcOXDUjQi5xRtIMcOYbU9j2V2Hn1bIHeDGTBXb/sXFH/INiPkhP423cT4AR3gZOp
hdR+ZSYk0ISN20ALAiRwGhdV3bRMsXJHZLHAbLXS9TM/bvvMUYscWb809BUWeKFM
ShmIvp55x6XXUmb4Nkf5O+clnBi6HN5oO2U17GwLp5Z5+dx4E1CdfBZCNeHWwXr7
O2a4gl5v5Q1t6DLSL1a/ids+rEHmwmqp3L7SagPgvMZSMaj2qS4/w799KLK/+faZ
Ufwkoo2Fzqa0qYv3CEFO+y9/lWD9t13eRL3oWPR1Vku7axS4orc2lcoXYRsvDv/n
hxs3hNftYjcgXP9y1t9G2WL6iLYrzHyXAshMnhee6y6i2DT8VvXTKBn2SekuNBUb
V1dwtnCLRqIA8krPSTT3fKCIx2NDWGRtx8Qj4aOJ7ghvM1WlHcxSUV5MCS0g/T+0
k0BOdCRwi/dKMNvnbyapjpUjt9ydKQuMqfmQcRKP+thN092hW22CMbsdQTyk4nOD
w1v/+dotiP4igBRsafqde8mFbOiXb8JdZuzAV9cIeX19sHMnT5BNhMFCCmZ9dn1j
ld/k3DjTL8Ha+cIDl67OObtU/DtXyCSUDhj3391Cz5l9dDfvfboQsdqPLfj3tl4O
v9w4kcWZkq9uVbG6gW+9YmmijqkekQZoCjP6OURLvpCfji0hICwTK0LYK25s7pJ1
Je3WipP20xF+QoA6e+afUmreIT4o0miUoyFnbDxyjupoIrwVgUOki+gTYeFynn/J
7dPl9jvo1gmUknJozyrxX2f/7H8F5yYzpFqwzV/Ch0GvBcQ0ccpXJHTv5niqFvM+
ncXs1KYKk6E7NZT9ojdYwrOERerJl7FfBTUoFrkYAhsFj7vXVMWZ2Ns+QtVlhcAQ
nJicHZ/Tt5evLcEtBB61C2+uvVW7LE16Y1IJiJAUidRlhji0UYpG16C66Zx3cRdh
huTxhyPDhwg2P+IOTFgHR/LkRqDXl/Nn6HarUEu4UU7DUnlxbth36zS4RV6B4eHF
`pragma protect end_protected
