��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z]F�~�b6ˎv���O������-�v��UB0��[{�&#39I� ��Fj+���S'���&%�L�
[� DV��xPҖ7�k���A�9�+�(�v�
�ع/L\@�k4�u�C�! _�t�@��\"�oJU�F��[����vH�f�;gF�)8�޺�	O�/]�kd4�R�T8-��^(�;iq���=`�{��h	�
��'L�ׯ��O5��)�{��ϩ��qjt@gJi�ڻ�l���������n��	Հ���%��� �WO��^c�[�fy�vA��0B�܊�� �
�A���z�.��x�b�p0��/:	yy�^��݇-��o6�3FM���ܳ���gj߯r3쿘ׯ���������>q�*�Ϝ�X��bm�4��f�h�7S]I05ם-@��l]�g ]-���y������Dҷ�q��b�xk��el��'���P�XU��z�&�n�`HzAi���ᵳ<v�;
@�g��k����3$��o�5��!}@��X�X�_��$A��� ntT�Q��u�-�߉�t}�*-�7:��^�)�*��G��簚F���@�s��*e�P�Uك�{C�u�����zt�Q���A���0�ȫU+�a�5T}�V��Ս��/�*�vL5�H�_��r�0��*��u@0[=4�^v8Wddqo����XμP0C	������U\��]dD��˅V�6y�yʺ
c�����#�*�#vH����e��*5a��W���qSe�!�=��엪�_��(�@E��2��ީM���3ք��{&��Q�A��}ȫ}��AfUԈ�x�6D��ݒ;,�Mg�5V`��.}9��0��T�hM� Ҵ����ݩȽ�y��� ���bc䵺~��`�Eܢ���6W�tM��Fb^6��c;|�R̢I��uVgX�eoݛ?*�}�� �]G%��	����"퍤B;���	��	��,d�\���%ġ���!���a�noI�x����Ah�Q{N27�ה��3�&
�TxOtCGW���N�0џ`"&��֠�#��~I	፶gV�Y�N�.�ZIe�}J�a�T�}̕�#��^��KaDzK�TY6�8��Z��r�5;����y	@{��*� O����g��(a����o?0��k���4�{�H;�T/)�Ȑ�:=���������>�k�.g��#�'j�LrnԸ�@�
=�©oo���STz7�9�,/,R�?���'sz��t�+�E����:�x���2�ck"��f�+X���u\kv�[�y:*h���#�=�����������/��ύ�z���?$��v��T����NK*87*�1�T���:�#\���1&�0sM]�v�pH�ަ�"i%wƂ<��)���tI<��A.�v#��u�ψ5��U�o*��.$��O.����p�N}V3�".5'M	�"��6�0۰�N9r[CjCD��Yrl�Q04�_�Н�Qn�VXBom>�����b��R�+0�p �g����:� �M/[J²�B��g��*aQ���I��I��J�<�,���4�+�ܐ�����n]'ʥ��OU�5,2h�k$�6k�Ta���y��p��I3F��C�woC����2�0�q�ȣ��2|fx��n��<1�~ؐ��&QX�{�1��<O��q�����&�A}�ISZ��Q3���YԹ���	 ������ިN)�۞�B)��!��C�����J4�u�X��+$޳%�����S͝69G<^Q�����}_�NX�o��I��sP��K+���*E�<�EgU�r���AQ����TK#O6] "+ם,k	��0�[c=8>_d4E=S��'n�������F�(Z2.t���z�ږ��Ӊ-���6ݦ��'6r��������v"&Wj�r�ť1tҎ��Tt":7B;Y��[�9��	�l|ϷkJ�j}�P��_�8=�޳�� =/O�GpF��ݸ�����*ߗ��g(���Ʃ�K�C"V�%�N�_��@����V��E(n�(��E���v��>�+�8v����S��IЧ�O��P$�A�s���c�t)��H0/v� BNr.�h�����0J��i��~Dk��G�a�#��_ {���SbZ����FR[WO�����Y�έ"*ȕ�jS�.m�t�n��}�
��`~q��\n�A�J�]��V=�,T/��nD�[��U4u�ƽ��p܃3��,�C����틶$�u��ふ��l-+˂E=�,�@�C��쭝��?8����h8��V飓rA �^(Ʌ���h�ٲeqXn˙/�`�#a�>��Q�|]PK����[�o+�&�(�qv���>��$�Ḧ́��q?V�U'�/�>� �-��cc@��LL�����x̺��7#$���fs�.(��:�ZZ`@5�8j���|��d�kf�[��5ώ����;��2�P^�.��ƭz,�}X}�hˈ�n�_��;��u���� �I��`5�������@�[=]��Bup�\x�Be|n�y+���+�y�	[5�x�K.��������(�M��r5ʖPJ6�X���C�d���?T���LJ1��xT�վ. �5M��2ap�[�R�d߆OI�K�ק��)q�C�}��;���Z�
��/B�s�Ū���.�0��w���\�Ie�(=R�Z�W2U��	ƚ�'� &�/sOa�s~� lׄ�����xO�T�C!�Mp�����Q�£�2���r�~�M_"��o+&��,d�jWEr�y���|2�nz���@h����K
��Ty<�&��Ֆ����z���i�5�?1V�WX��2���Y�˧��P�C@���r�3?�n��'EU.YT�*�:Ⱥ8��l�I��$J)ӻ�no�&�n���֕�/uI�t��v'��i� Ӡ54�S��^(.���0D���H�jl�<q�|�o8�u�V�H8άE�(�����*Y�@&!=�q������:v���m�an�\��~�݋Z�
*�(�n+�x7�O��J��cE.d�4>2ƷEV*�^ /�@����s%aV�&Gv��k:�o����ص��f�ltV�5a�=����w���bT�O*�h���a�&�qF*e��p�W�X�46l
U8���a͆�{
��[�_n��L%���ԓ�~.o�v�)��Ѐ9I<U��>[%�+bN��seK9�����?��;pq���-5s|�@�I��֊Z��3������>d���ff��w�v�8�R��&�_���]�)�y�gA�e����j�t�ɺ!=O��B�N��<�>����J�����)���c��ً�M>�>$�&f��":i>_�_ޘx��U6Mu]���,���=��� ��섓*��̺�?ǯ�8����i���#+r2��,�J�fl�?G�b�xW����L_K��6�ʂ�՛
ń�?��8<�O4.�g=��B��\���G���f���]��Ġ�g�e�8�F��fe��j]	�&)ᕓX��v�����% ՞ONEb�q42���vb��0��*X�/�^����A)��
�5�H|R�@fחH�	UKX�d�՛ñ��:� �-���p��� �L���T�o-'n�l�}��N�n�V����G���໎3�F:i�96Z���h�ӕ|�MJ�_�7���x4** L��\k��*s:�=�Z��.��l֑�ȁ��zӆ���|�+������m(ݥ�js��]J��43�+���8]��7:�����z����!�!���p9A�s��3oA�`պDJ<NU4ZN��(n�,}�F��v�v˱���1�G�j2�l�F�H��m\E������O���$��4�S
�հ�R3D:~��Wx68��]7�{��������h��
��C8��XP��mĩ�ɝ��"��˷��1*�)[1�
�{������'�^�����ݿ�����^�+4��p��gE��B҇82������������h�z��2.n��F�o��z�Y�{�EGu��$���MQ`'���67�Po|�0�K>(��ୟq�G&��> `(H� �uM��a�ӊ��H>����x�Ӝ��J���J� ǳ4䑝������	J�G�3��t�@����"��3�����I�&j��JF�j�4o��l�&K�˙���A����#<�;OX_��~�8�F(pk�N|���\�i��rхmLH�ߢ���&/uU���P���ң��E�L�C�x���=���b�75,ҽ��QR��[X�*�V�6�F����`J�E�r�(�*Q�{/���[.z�b�x.w�0 Ta�)�V�X����U�F2�Y�0$���7�JM�_ϖb=���
9�D���%�:~�h�g"t�"����j����M��eKl��:$<�-o>���H��� c8�(z�@WJ���4� 9.h���F�~��r��˫r������� ��Y�G� �l��/�	4���.D�#��i��y��3/�$H;2j4TU4N�z�2��)RU5���J�i:)�H��� ��1=�	��̴�
;�_�W����1]��NS}��4��7�!�U;I(wN��.�K4�GW�A���]�X�-O1_H_�0P �Ļ'��/����ٜx*J�n��8�l{z��8���lU��z@��D?�pO�OU��wc���@㍪���H�*�,�H���)4��\iOua����oI� �u�Xi�	� 2�`�Cva�}�\˽L���8]s׽d��,�x���j�`�U��aN;wy3�`m���{��ǆ%(��Ǎ��w� ���@�k����P@!ɷv(���3�W"V�>+#��tx�:���b`��,ʕ�ك$�R(�Ua����y�#����换�h������r��ȇ���j��mq��7��8N�E�Pt9�@+�E�4�(��>��6���������׷p�x�3��R"q0)5���q�?Q�«��6�
.fzu΋yy�'
Ĺ
�>H%�7Т5̶����+�eV_��.��� ",b����**���^���W�1�;���K�\��E�[�O���W��O"i��]���Mq	������fy^�H�u�e=ԥO�խU�E�۷��E�t2�T�锕Y趒!]�3zU��hX�r�0�Kvs��R��+=sK7́��ٟU該F�&ӃY M�@;ft��shǘ/g�J5U��U�w{�Jfm3�eN� aNw�M@����&8moF2�}Qk�X�n���E���G�we���L��+�T��xP��QO-lH�F��<�v5"�|*��P��-�R^2X��O�FH��ʧ�M��jJ��Y'^}T1S����u@Q��?�~�<*�W�5o����=/��Ҋi�*}ȳ{��<1�q�$A!ϡ���${CBP%Xku��F��s�b%�S�� ;6�QUѶ>T�����M�t1��D"��@n��=�y�b`U�<�͔�c�}'޺�#-�g�{P�/�N�s�JH��,�f�R	������_q��Y��Gc3��}�?�@.��߰��l���=�(��6��`cp*���v�_��KC_�?�l�>����\bl�{�����������#�l1Rշ�j3�H�"���Z@]B����8�%��jv������h"����j�s+`���&�>�ErA6��'�K��Y��y\�˹�!N�nZ�)��=���`�cޚd}ۥ���&J�m%n����E_A�U���C�s?��h�%���`��[�p�N�!0�]-Z����w�q/�QȠ�H���1���E�&�	���@��/x#�I�Td���ć�7d�q4<M$�j��:(��r���2��{*)$8��`��4��*z�{�&�^}��!E�s�M��+}�*���{r|��%��1+:��y+�׳Z^�'��Ԋ��kq�1�֎�)|��og\�(|v�6p�(�5~�u�+�K8{���#�j7���e�����:�7��N9P���*0�𾎎b�0ٓ�
��Fm�3�ˬ]e����S�.�M��Ϟ�9��#ժ4�:7n��ӆs�8��!��:���k�uu�`�D�*�N��x����Y&�D�D����4 B`�r�{�����0����Œ??Eҙ��
g<lN @�^�h��(��y�K\����k�����f^д�k�vj��c�8	D"����.�aO�Ǌ�{��Mq[�Q���`�����7d��7�_�{@���4-�ε�3JS�S��t�������.<:���04����)��͔���h�vI�|P���<�`޴���L�[0Ш���^?��]w�%�c7�U�/
@]��g�t��)8�u�PHg>g��r �K4�L�Yk?�����
e��	��P.Z+	���	 �й6f2�~�Df�uIⲝ����9�b1��V���( ��5��y0f����Q� .*�V5����2��pH�V��_����P0�"��c�j����;��ɞ�� �U��i];Dj6 /�.����=T��V�sa�
g�%�1x|��v�3^�U���M�R6
�����r���]���3���2�*P�و?SQ�{��Tt^���Ӄ�Л(��E�rE���m��FS�:���&H�|@X��
�y�Z*��<�m�(�dP�gu�u��������')E���ɲ|�1��'m$O��v�ﶬD���NuD9�s�`��<���#>%
ka��!rI��#,髷U]����,�$c��
�5>fm���ṃ��}a'�nj�����������>@��v#ڳV��q����)�����W�݈J��X2�Ya�F�Ժ�	G�:��-��n�H^,�����h����]�(q���)�l0q5���0FG�Ыm��|�7|�Vj����>a%"nobx���W�ԕ.Q�X��5��@��E���8OΫm-�\�4�6��@��c/��9}�/`���.��~hj�-��	�%o��VV�	�u%��:��6��/��{L�'�V��V�p��R��v,���������p#��'_X���@�9c�=��"h�-�d5xh8�`������D��� ���^8Gh�����.��`�uY���x�2hgW��&px����V%]X��,6	|ƿLg&m���6���Y�ZL����!��%�ְ6�3tx6۫j���<�`ğ&<o�
�z�H��k���Zki�%J���),�鼷R�U2}T��8bƇ�VJB�a��ƚ�`�I�;�K���Q� �h)�<~���-�����5���˩l�Gh��9��8gZ��G�HK�E��χ^���{�o�g��Eޝ8µR-�`��nk�ۖ��ҧ�b�I���ы�S7�ӷr�%��ֻ�뷲
�Xb]^yw_K�C
r�}����i��K���!F�2H��+(�0*�hbΕ���C�����G9��� 9�D�AR1��HD�[S=�ϗ+�'&����x�K�K��ѳ�'�^��Z����r��[�N��1��<�y_�7�l%OoM#��KY��������,�M�[Sta�C�s-�V�q�Z��H7#H ��&7�&���t��&�}��R���]2��1]�fD1=���˷�A��Z��nm��+<^�qO�:�ܞ�EB(du^���a��Q+)d����R�e��>�El/:��=� �Z��B�of�r'����y�&4TcC���+`���yQ"d�L1��t��TyEj#P/��].��mG]#agaM��ݲ�f��꒘�%�Q<�:�����v���7 �f/����W�O��$R,��9x!��m	z%����;`��dz^�eݦ%�W�U������a�������|�ŬP��I�B�&�u�Yxx0O'������Z~r�<z3�����5���`G�����
�.�ķM�M.��m��lz���#��������q�D]��6�9��N8	�;�}�r�+�3�Ӗ�4���7ˬܧzWV�a�o��
;�-�&�K��\�tAsxZ��Z	��5p��_rw$x�jxZ�����ˇ�;#��<v�eGpU� @P�G�
��P�8x�x38{��w~]�b��3!�3��l�:~f[�"�6eXg�2kl���go�V$�-�꧛������;��v��5_�6�7Ϛ��:�Z�&���Y��R?f�U��/�ҷ�[�ȆP�\\�!��x�~�.q܆S�40�(���* \���Κt��l);��)�J-��m�I��5Wf���k�-N����L}k����%�f���R*Gضo�h����ê�������g���`F�w>���m��]֘��L4�)&��GzI}�����{E5�҂�WL��Pk�QQ�Qv0�?W��yK�Or��݇@�n^�?q�s��R�Է)��>z8��.H���vD��(p!/�8��*a�*�T�}�[�i��@���=�̞��7B�Z7N�H�%�&eޘ�M1�>h]D��h/��je���%6��d(IX��i�g�0��U��_22��G4�X�� j.bU�	��q�;����d`Nү�8��|r�Y�i{�yO�B�i � \I�j���^<~2��T�
5�C�asNp@�,Lu2�����Y�'ڒ�S

a������冰��'�ʞ� X�m�-����ߕ�!���gɗ^8(�坁@}�m�\j;u�P�킭�tu.�}�c.$�lmn�&�����g���q��/�wmԢs���.v-���a⼐r#���Bs��EW����b���t��q �<���]m�&�֡�ڴ�W�S���aq))~����}���wy��v|�y1��Y�v�?bA6,QP�Z��Z(0OM}�F?����_Ie�˔�m�,|���(բ�>;�x�+�qd%q�9��3����Q�ͬ|�I_/B�	�R��g� !��t@����itZ6�pGі:z�XR�h�@%��Us 5X���bPj������0��j��{	�ɗRՁN/PC��@����\L��0�!Y��n�\�U]�=փU��0�.+~� c�^�� {:� �=@k�I����Ь=c,z.rxW5��8����KI|����FX V�E��#�}b�? �L������MP�}G��1���-Ӹ��-�m��5���a.^?v��c�eV��[vB��ݱ�A8�JC�4��Bk�c�R}`��-���<��ߖdԼz�� |��FcSC�W�DU��,�׭0oHu��<6 x�� �"B�+��R���L*~��.͝�
�������5A��;i�ٺ�ܥ��	%���z���h|�*MQT'��ҧ'0Z ����G6X�o�h���|9��!Rw�5A+���D��f�~��o�Ѡzs�>f%�}�رrD�'�r���a��J�ꋩѤ�[-�K%l2���p��%�2�}U�qr��-f��/��ۿ��,��d�0S�֦M��N�B�N�g�k�.q}�<-8=�rd6��ǟ�
0'|!������|�,�����	�rᰄ��X=��kt��.��i�8q�6��(c�gZ��d,r��q�UU�	�p/L�W]�X,$�.[�S]^�v����Ê�_�Zt�
�P�E��Ш���w�{tPW_��.�>\��`�{���(_�:�1��� ��V�#d^���$�"�t4�ܓ�:�P�n]�J��P�
(@�t��KG0eU}L���3c�� M���D,\\�ӫgi��:.ۼ����N��E7c`|������!"א��@����<RM_��5B���=0�Ū��{���l�-T(�"r��M�_ˉ8r��e{T�G/�����2#�������oMg�{-�A=C]��{y��J�~=���V*�\,C���%,��,Y�ۧ�3�-c� o3��5psZ�����y��� ^��;����������A�����D��GGƃ�dhR(s��2����2nÇ�X�1��c�$��[�G����t��T*�T���虡(��g�v7������i�^uހ�|�y�|]z�7Hb¶-��-�}�P��Ok����O�ɒ�/��tZ`��߳5�؅��}>r�*�nT.�ˣA�V�T�pK��x�a��+NX1T�mr��@�v��u�*l���Ԝ�������!t�.*�}�G�}3XS�ڭ��������k`��2�6U���4�',�C��!��m��ZoR%vJ�Ь�J�Be��=��C�5&!�PʂGy�2;M�3f]��6鼊��q�*�[���)Ւ�^�\+�@�Ooy� �9X&c~mD���s�+��W��1:�n��<ͪ/R0��>�4���e�z�`��8��p�L��L��Gñ8/c���rNlq5I�7�1
���̈́.	�*E&pF��K��O[O��eq��J����Z�C+�5���P��|�$�+D�S�/�M_�a�ϲ�b.�?&�=����A|0:nH�������;fn �=]
��|�c�ge� |H6�J(�d����Z��b��S0Q/���0�ɠ`��]HA�s�RGJ�G��߰�3��L�DW�0���]Yճ�P�`棩��^nA�Dq=[H(���"����1�
	5#�g�l��=��\��MN� �%�b����Q�BL[=�"����D�Ma2
�'U.�����@�w�0&�p�j\W/����	������X���dV�:tc6XMQ%U)J!�R�0���y5vF�h��I��z��v��\�G^��5����J )�:I��p�+ۧ�;��m:�;$~�ї��µbF����i�ċ$�ܛ����,��a�`�vf�C��RF��"�B2�Y������9��֏\��ui�	П�[�A[�Q[���QDj	|�@f�t�)@�u�˄� I0}Q
.@���&9���Mt�pE��&e����y,
mY�%4g�4���f1U�݂� ƌ�Ppb��A����ii"a��[�C>���HI�=�O`t�HI7J��N�����(��^�4�Q��o�a/S.xH@J�:�2��k�y����#�ڢ�{���X�ߝ� �+���/��,�Gzm� 81��j��G�Y��},�oD,���56���em��	�_����?3�̮ol#��q��q�ܿ�L�����*/��,7t.�7K2���1`�����.R uPizUT��cl��P
a.ƪ�6�^�$��3��t��F>����k"��WehWGj��//���GMm���&]b���v�I�dt���a�O&����K�T�q�?>|����fwˮ[��z7�e�dG����n8QeQ^�ϯM��`̝p��]G^a> f��s�78��7ֹe{�pT���}�O�}R'd|��k���!!� Ⱥc3X�"��v�� ��|����q\�5H�G5�	t l�6�:P�B�#�����Ƌ�H�fO^/-.�f`��=PN�&zy��:�WgDʩ�9��C���[�R�CI1	Y�v�����ψ�����iH���s=��b�?;z��˸��ĺ,�<᣹��)*1*󕎟��a��U|k�{����h�О��B�.v�s���#�֠������ޞ�d���'��׳��w�Vt�=�w��FMƍM�D�{0�Tj�Q}(�)YxՀ�13�Pܡ"K7#�;�|ȳ�R�Y����G�MpS��%���φ~��1��P��k܅!���J/U����w�x�~�\S�ZB:ڇA=����� ��8��g���#dw/��3�D���zJ��P0�^�5?ќ�!����M��,)��0�a�?4k4��?�����sӑ��c.��"9m/��o�)`*pl�|KR��q(5M��C�5��P�9��='����?��!�¤�y�^�W�#�p�u �H�av,�kz��7�\d)�����!<����C�S�r�kK�ѓB s��\z�K�f`����Ɔzݣ�W��KM��.��,�1�b_ TF�t �K��?Q[�RL�E��q����Z�z�B �B@��z�o���kz��U�w7��қ��f(���=��W�z.��[񖪜��w���R����t���s��/��̷�� QkT?'s2�;�����WE��;!��%�E,�P�e���]�v�o[��5y�����X�q�.�CJ�����.�а���;Ҹi��ќ��Ȁ-"׈"N�؛SEn��$N{��r���`ޗ���`��`ʋ����0�����o�t��ݕ$�p�q�䖍�B��)G�U�[�3�
�@�o�Vi"/�����	A��K6�9+�3����a�?κͧ� %hoN\h+���diV�x_A�+��V?��E��
�����PcZɶ���U2'��vE�Nt���tE�?"v�N���&������ܩzD�Ri��r|ܜ|��/>9Y�
���c�z�g��_����i�I_�n-���i�d��\�� ��~���dk�����?*���J��Y���1և�¿�����Y�I�����Ĵ~ҳ�G|<>�L��|0ϪP�S�yN=�Sa�d����$G�3�duZ���ñ]�1�yǫx�q�2���5TzQ�[�s�\4-��伔�K�1��'��Xͷ��LL����� x��x�+k3`��S� rE�$"�T��u��d���*����D*�*
��Ŵ�G�.��&qCe�n��m*X /36�O�������\�Wn��%k�}�Y?h_�H��t%���"�?p��,I宯k����.x���]�B�T�v@�p��sx}I���5�qDs�V��
��Y��2X=m"��L�blO��ͥE�:f��B�.������D�뷞󝂪I�0�]�nR.7��Oos���p�>�s���cqs��\��ϧ{�+ۤh[v����[Z��.f���AܹJ(y��?�qE��DIGj��B��Z����D3�U[��X��Q	���"us�������������E���%ؚ��6����P1�{�����m�bs��'#�Zmvbt1Aմ@V�k�[����v+�\��J��i�`�1
�}�ͣa�;�ߖ�a��"5ɹv��c��?�OG�|yJ�!wŀZ�ۘ�bE���/̥��
���?�� ���,M�E�������D]/|��.�3�r��p�Kr��v8}�����o�-Մ��A�|PL|L���j'�o-QqG���(�A'�����_r�[�і��7e��*�T.��F�Hu@o}D�̞��ʉ%n֛�ϹW<�q�iBʪN��	(�m�m�0,����tX�J���RX7�F��R'�'�r��_��!X�N9��Z>�5�Y����4��SQ�+m��4�Q
��"�c�D�|:�}��=��ְ�ܡ��>��'�,��a��ٽ�4�B��n 떠bI|�[E^��**I�7�)"2�R�Q���o�'L �*＊8�G��T1����.�8�%;q}.��LA)H��^��K)7�^�kq{0���.�4�χ@J}/{���;��\V�&��JИ�1_��ɜ^�g�;��1�A��5��7K�����w��I��Ωt�/��j� ���>ȭKꋋăl�P���Qr{	�"+�Z�P*$��ׯ�q��:H���[�Y��V�o���ܛ���꠷�䐥�ÿ�'X�#_Y�'�&Ӽ[�tBn���^+W3���^�r���z�WWźzuv�~L�
Љu�b.������4���xWi�9��mbo���.M�Z�}�%�ɘ�&�����#���ab��h��Ӟ �y������z��ɂd0��X��H�y�#Ie�ov&J��հ����0U��	����s�K���C������E��^�I�������2��\N�mGۭ�j���U>�>tk�4�{?���A9M<w7D�;�馩i��uk��&Uk��Qr;k�M00�g�i&�-��jK��3�͉EVf9oK��F�ԗO���a�-�6dgOh&���L��<��:���"4�"^i�O���զb�X.�p���I+�B�t�ǁ��������n* ��op�XN+�!���r����&HݣԠ5{��{r:4�A
ð�nx���xh�+l�PiC�E�����D�;���=�?HP�E�T1�P�x!�=�M��L�bJP�N�Ϟ�.��e�_���hCX�Or6 �yd�TB޾3�(7ǸI2~e�'��`�%�n.��Z`�F���J��\�#I�ׄ��0vh�	�@L�sZ|`�v��H@�8�ܠ!��p��Is��^��&���%k�(� >����,�����|��_�E<�� ����iWB5���c3�f�m}�t|��U�_�N!49��������1�����m8?�de��I�l^��\v��4f��'K�R�Vh��<3Iy�,u�E'�>�D}9׆Ϥ��T�EV������}K�~~�c�����N�ͷ�e���ŉ���2V���@J5��Y�#�8��Zo#s�e�Y��AР�=�����4X��d�<)`���?)dT���i~E�\	W[_���^�T�>zh�8r�+�������f#���}���;E�q�|�8GX�#�o OD�A�b��E8y�eH�Y� f ���e��C��7?&�{$��L��G��v��^��K�N�RN�Xx,���8��b5�\�]���<FW��K�Xś4��զ��Og1�����K(�*P]C}��?��?�Ď����J9�l����?H�i�SOt}�ˈ2��q~zC����0=z����W=�K��3�ʟ����o%U��jƽk�I8�h{��:jW�+�������Y�D^��?�d>_'L%5k)�@E��ۗcw20�Cо ����J5�!�2����^z¬��ː�~�D��8k�XNv~�~�G�_�������@��Wi�Pⷢ3q���T�˘a\䯞�lsT�j���ߚ�֯;��#Hl�{�h�M�ueדn���@W�K.|;�ʠ��ށ��e7x�o݈�b'�V닔���)< �%/�u�8<Y�Y� �K�Ӄ���n)��~*(���4LY��L�#f���YV�5�F�(����RZ:-o+�(�:E.9�<]%�������ٔ&P�Z���sI1E�A#���r�S�C^n���������_��lK:$%#@@X}\�axk�p�C��k�)E��ϭ]_�"���{'8���K�z���[��mzGӆ窜?N��鼆���avE�?m����׬Ԋ���k11W5Ӛp6��y�	�ۗd�`��P��:��J�I6�~,Px$��kp��m�7�ng�}��"�Pܘ(('�P�}YqW+��Lq�^s�N���г�&��z�y�b�d�����k���E�'�{�e����g���l�� ���t��Oq��zÞ��h4��.��k�W��8�ayTC�T�!��<�@�뫁[ꜫ/�{\���Ml�����m0��������DQU��ż��f��Sf3!Τ�[p��Z�]h�s&�Q�[T�lf��nGnב��,�4��r�@j�8X�F���J/���ڳ�]��;�{d5l��ŉ�w�N��&4ӣhKl���d�����g�z�0���M�X0\i�RN[A.����c��y`������S��u��6�_=D9 �'��5t+ �D�;+K���[o�%�(�?��(����b�iY3��~p����m.d��}� � �����YC�Ԥ��f&�����`�fMV$ )�ﻮf���|��zǢ���3ȝB��b�s@�S��2y��3�ޜw���"Ey�>u]#E�a���6�
"���X`�!�1�[Ⱦj���Ʈ�P��飋ZR��e�-,������ҼY�enZmfO�ܔ��vpz�X�rm�E#�$������8�/�zlu���b�qx�x~_��̲,�m[*v�蟬a��*�����V��Ob������o�:�tB�}l\.)��F�Th��V��$XQx����o��A3��M�5����Kn����S�<����_��q�.�����ץ�[v}i���t.`��0���w��I�|�L��:N*��؈��g [{c������e��ed���K����EI=gҌOV�v�9��3�(}=����~?�Z�L׻��"s�!xp ��,ٮ��t��u�9�.�J������5������M
o����>YD��ʭ�����dځ��^	�ƕ�����w��L$I����_1��Z@����UOr�Q��	�η�7��H1"X��%����[̄J@�fE���?��/�r��f�����+�� ���G�s��y�1ѻV�n�g�T�H����a΍�C 6��fY�´VW'�U���Ew���>��n?{�༳ors�>��F�c��nl���'P�kͨe-!�p>����D%�g[6͑VאO����	*���j�=��/;[��BA�����Ă���υ������E>[��8�V�jx<�P�5�����2v�������B@��&Tv�&�3?8w��md��rM���g[�ثa����G�3$K�:ט/��B7�83���Y��25=�ERf�V��L-SG���BS��n>삫M�$��i���p�DeёA���nBy��]���Ó~�S-�5Fl^ z���P�%hg,l���M޺���j� ��o���\�Q�'s�!��d�}��E�8�;SVh�o.E��s���*".�X���'�]#��wE#ڢ����XFz���TRo��͕|^�	W��o,��y��j��o�d�0$�quM����zպ�0�Y����6��W$ʑ[�"��{�����d4�[
2P��5��1�-ⅺt�g�hX�Ц��TF/�B�\K,��6��S�|c*ҬȻ����p�oa� �ӑt��6-{0�+m~�u0/Y�h���%�_�/�D���2/"�@k��1�&>ț|�ue>� 
��8�4�Q���˛3ƶ��7�ԀV���zތ�����H��pOp4|��%�`L��d�<SmqAu���d�]L��ܤܹ&(�R�"$�,K�]�g� ���S�t�*�/IRը�QN�S��A;3[��Rά��b
�5��T�]W��Bs�F���"v�Z$i�!?َ��I�H*b��_^� gX,�Y�@�e�VY�Bѳ��2%���=e�U{�>H�,�e�a{��ڹ�mfnb��N��/��t�^��rG3�z,���P�׊��1:t����!��v���9��Z�l�t8�Qڐ�+k��E���n�n)[ ��T"���w�t#����1)�1_V�Jm����(��W���"��^�+=���+��}.����[�֊(M�2��XF7�o��!�U�c~�����\����tWh1�xp��|�>WR
���/D5�f��.r��Q�����?�.O܎y�:�)�G|K���a�x��!�K��<� ��=��|��p���Y��e!^T-�z3n*�\�t�	ג��re�Լ�5y���wd�c·��?��|�����v�z�	�NP�����c�R�f����U������E��V��ovs

��3����Q���W!��U��!G����^/�Y[��<*J�ㄝQ���d�%cU[�mPLpm^6�>]��$�Wq�Ͷڶ2lc��n��;�����Q�a��r�
�$�B׷��SD⼁�x<��s~;͏=ђq�P�j����q��_O.��+�����jD�F�(گu3E�a�zqumS����J]tPI_��3����-��"�X!TSn��Y&�ú�V9�v7
��IW"��&<�~
�H\q��\3���xP�tX ϓM����-��?�i�Ѓ��;��)3[�Z��o�r�����.��YS�5@�}VEx��~N{��&LǢ�Bp2�/���]���t�>0�nn�3�1/�K�C��~��ѱ67�o�=~�m��u]uЭJ=��g���@n}oG���k�(.3��f�M�^K�����,��p���.��{{�B
ZGOZf�s���1�t�� K��8/�F�4�c�o�S�W?[�Υ�RО9v@�,��n�@�"��
AY���zj�3Y��_���	E���'?���-�1�:u�쎯k��I�!2�	*��IC�����
N��E_�:05�^Ƈ�,ճ1�k��7@� ��A�+�����Ozp����C��n���A�ע,Ap&�|�Jǁ��(����\���pYI��o�SJ5�N�L�~�~x>M�	x#=���m���ݲ�:�x�}�'7�.H(�|Wg9fuf�?�ʒ��)X{�n��5>p���w�Lx+�����w�lrPC�{,E���&1��/R|�9Y�T+ �B��'�Qp��Ȃ��Il3��\����~����/����3tk��BD<O�7kR��v��#*f�llqI�q���-�hn\���5L��:�VK[��Z��n�"p�@�'��j{���~E��s��%�z������Z�8���x�Ɵ�Sπh!�bУ��ӹ���A��o�8�5l�5��7�����NK?��fT7��e�c��A�w,���co�u��]Ġ���W���x|X��ze�$Xb$���8?K��1�P���k��D�6Ӻ4��{Xq[�G�������*Ϟ��M�v�Z��Q���_��[㿨���΃�®;�Y۳H�+?"#��rϡ;b5�뇕������r���j	�|ݬ�y�`E��px�����Q
-��T��^ ���đ�����BV�W�k����ߘ�`!��σh��unul����7���^���\])���2�9�1%Y�O��0���-p�5-�i�K�:���h�Lx���(	�e��^|^�t�.e����O1�.��!,���4)R^m�,r/*�&�[�Ϧ�J�Y!Ib�oN���D+x=�N��� ����`��K
���ي.�br#4�5���ȯ8�4eKnQI/��J�,.�N�;L����'b���t�OVr9h4�᫫�v�X��C��-2O�g������� �RM�ߜ�����ڼ�|G��<��#8v���fq؞cX[���8~i>Ae�"��+����d0�����4�"0iAxE,8�Ϡ�@(�(�O��wB�@)���G_�!�[b@N����R*{�Ǘ���Q�i�#�h��o`6��&��+'��p��Í
q�����T(����8���W��mF���}��q2i]u���q\}���
/Bx��<�����.�7�[����E~׆��|Y�r�^��\6|�pM���^�p\�;%���i$��|�K��%�}�Д���AR(��1 �X)T�j�q�Ӈ��?'m�di,���e:��D<0E���CX��3p�Ud���zM� �JT��Y�?w�C���bk��h����̤-1Tv[9])0P����H��ɛ@\+е�r~]4���Q�u[|M�w؝������J6����0�Y������G�E�Ԇ�$�����4=��7V[z�&#G�����U���l4�1|���d�*��/4V<�i5�{Ol+?�<W�/���/��{����@٘e+t�K��jF+~�S�Ǿ�K���}�%<���c�Jk�Ú�zy��v�b��ʔ1Ѻ���I#S&�$ʈ=K��L:��H40��G�z��|Vp�4�?nwx��kӝ�/,'+�]�R4�MS��`���&"��MrL�/���+[�R�z@!j9H����� �;�P��������/H�g��A)dr7���mF��Z�]F�e�cv�^��n�.�l9O���K���&X?�U����D\����f2	�dTU��X�;��͞*)��1O�k�ErZi3"�Q�h��1�a�'�r�f�M܈���C���Dց3�%���k�f�aI��H�Vm�>�{L3�K�$�|��k�9��S��9A�& |���Z'�V[�M��a��1**DC���$�P�\�!Q�>HˌR}�z����Uo��<��.#�]�Sh��qy94j�R��X���0AtҴ{�C�J�'�s�벁���Ĵ���Az{��@����*�:1'���1H  (�y�ʞf���`eF׃M���b",a�:P�r8k���r4t�yC��oyBX&3v;l-�P(�8��ޡ����2��2Fqq|[�z���.����Y�a��9��@��rx}]����*�Ӂ�0}8q߻�|�|V���Y�Q4�ZB���Y���ǒD���zKx0������Y=_�,�Sy�D�\c��\'�3ĩ��kՔ� ���V%[�^	-�8�9��P�~Y�=n�<��5*b c�%���'T|éa�SK���+c�D,lGv�1<��X'H��UC\� ��@�������mcka�&�/�
5�F�}	�CYt����}��`��Tw���Q��p�׋�&�H�+�d��Iz2�qߔ5��'�k��t�u
Q[�!=���������aP��%���B2 v�mHƙ��?R��G�0�LO�4+�Ǡ�����$&�}_/���__��}U(��<����`�Z���=�xa�*W��	E���Q�/yW둣p�N�I଑at���
��m�%��M4��8���Y��Р��V��k4�K; �	����G����}B(R`��[oh��Y��oZ�9f�K֣���o��<8v1��a�׹d�|3δ��tF��%3zi]V^A(��KVP�ۑ���!P�d�u��u��a��Ջ���h������Xg�6�����v}��(ϗæ�]褹�^�P�nHy%�H`D̾N�k�^�Z��k�������HU�Q��=^o�{�+l��G�*u�8F8 �c��Ta"�JR��"�V|x�N�����oB*-x-�7|Iq�g?�ŠR�"�����V+�.(c�⟪/���d�$���8�1Y�a}���BٴIڹ�v���Xt�\uO�s�����  K�./l�胈˪����ǁ���|��6�xp)b��z�ڬ�5
���~�\�@�� ������]C�E9K*����K>�ȦlyxN �a�/�\��|~�7Z�L$��5�wIG�L��+<�Sſٓ]/ � ��� aE��1Q�=t����w�Ѱ6T�u�o��|gq۩p�-�K��,��|L�%�솳�{�����&Z@n��g�O��|O2 (@�W[��q�g��I+��Pk۷��CaB�c<l7ǜ�\�F�τ�w(�G
=�i_ҫ.����Q��L�6|c�F����>��U���"�6�GX�K�_��-�ȭ�vj,\"Vx��
�
�pa(����4�:j��s6~�@攮%W*��=��ny�z���e�9M�w���������6���ݸY�괇��@۸jY�[�$��y�5N���:�13Y_4&�ԗ�F����T˚*�(R09�^Į3^�B$!�&��[J�]�\��6�Π#H���(�@�U���"�`�(�`AST��;�5K�ϧ�{p@�ܗt"���VN�H�|���/��o�ޜ1�{�$��ٗ�H��)Nt2������մ�.��O�w�.�������x�~���<%��y�)�5\e�y����ˡ� ����u�쯰���M5*��p�Y�H�47񴚮�`a��3W��r�z�d^=a�'[{Xf��p�cf>A�����iye�����V�_&��T:�OS�4�]ؿ��Ɛ�4���^"����{�˶�TVHh�LzTqH珡Ae��'��A�� NJ�����xW}(��d�3i�����ضl����7-4���^��x�9D���GKѱ�/�j�Ą �Lw&O?�`��-�����k��4>mc�ZF����N�(�g&�-PX�Q�0A��1�F��>�Z��uWk��]�p�0��戚�#e�8���	Gt���휕#�2�pa�ї/��_�T`j�r
>�v��M@������8�(J�����d�1;��<�fTj#Y'K����t��"7E�#&o��5F���Y��'��A�?�~6�b@~EN�C>��n��`!0n�a�z��1z�
w^��9���Pu.��'�,�&�۵a�c7����J�Ʀ��@��^5�'�3� @>E���x�@ �z�x�`u/�����5:��dW,��+nq�Ƌ��G��:ȪQ����M���i��:�����r	<Î�)��M9Hd��Du%��U�s�F|�R/&���1!��f�ȟ�6���M��{�9�.Eqö��/;�=Ѱ?���'xn&����T��2���+�A�ȣ��4�!��p��]/;p�r39�l�f����� i�ưSLqp�T����&��b�<1sY&���놽�.eV��}���Ȁl��3}��T�5���:�n:8�:�:*��V�@�X��Ү+K��8!��Z��T:�~�y���X�$Tہ��%�l�U����op�pG��;$Vv�0rO�`	N�u�{��jgM^FR�,�`)��t.��ެ�����J�%n�
�t�s	�<|��������~n��ڰL���"����.�1w��p�	�*���MX9H}ٍ��M���<1�׊{&��G�m7U�� ��G����|�8��U��8�v��8���dt4������1��~�^���􈆶�T@���;8ښOұ���0-������S�-Fىr6��ȰڴF�=]��hL��?���_�Zyb��s��wk1�;p藒��Q����Y�IrL�{����Wx�r�����6� ���^��o e�<N�+9�ͨ�C�o��c�4�E������x��b@{,�-A�VLE�Xd{z�����)�#��fk!�Q�3nr���%ޡ�AND��Y�[.(<E �ҚZ��!6t0���w�}eo190��uN��g�� �9����um._��\C˅�V-���K��,�ˀ�E;Zc=�i��M����͐���J��<��\���;G�n
��E���(E��?<�7���ʚ>���G���(i�1�O�l���
�$���~����)�Hx�1�n�m8�8��(�J8����9�`�����Q��JYD���2�����݃g1������_�!�@�Rw�{B���2|g益}��W|z�(3᪎b{�V�!�ԷSu@M��,���� �k��K19�P�1֬��i���������Tե�����Y��X���X�Aaھ/���IB}���D��,A�g)�,�+H�zA!Ha���_8f�5�"�䖴Z)}�wlYrmJ��Χ�D&t�Xmx�=ٌ�s��F�ݥ%�c�h>�ݏ�px7���q=B�S�:���c���|wd��KƥXG3@I���l7xr��:h�8���U�7���/⽰��pY;٥���Lub��uWn�q47+$M��ȩ�{Ju"۫�U|�nR�ܝ�M�u�� l���)�s���z��� y�w�WBR�ݖ�`�dj�AR�fg �e���xO��Ip�t�k�x�: s���d������$���>�������jTon @�f�S<k��'��W�nwvɬ>����VoX]�` ��E�b�P���U��YLt
�w0W���*��r�֙ ?���jG��I��xh|4J�惂�}��.�������C0�ߑ��J�����=�z�]I��-|ŭ�]����}�_��
=GY���Z�&�[����LKF���:�=җ:<?;�����Wbnd!���+'	C蓂f�0Df�C,m� J��\쬔�q�x��g]uל|,�i���j��Kr�rA���^���C����C� �c.�$0k9��c�t���&�h����~�/z��4zݣ���(W��Y�a�|��I ����n&�5&w�N�.g�uڑ���Khw��h���$N�q�%��֦,ȝ���^T����©�1$U��Hί��@ܱ�i��H���~�M�H����F(4`;�%���-�Cis�C���w_�=�tb��*��N�`�I�h3k{K��0��OP�GPs|�����{n>jp������ޱ�Z�1��%��93Y���*?!��S���+�S��~�J���J�("�)�\��Ʈ6D�pq���	i�o(4�F�bs*�.2�'����ބ�c�}5�H48~hYly�&�Ԅ�V45
oD�Q�9���B�����	�c{ف]$��U �!�e�(�Q����:��]�� ��[O��LD�PP b�,ڶH#"���ߺF,.xn��$&-K���Eit��]�E��:��W���:�.����a�Ɔ�Oc@��(0-�Qc&g�bf�V� Q�	�PV�%8�d,R"8��x�﵎��fm#+z6���g��jt�@���
	�����)o��+���x��%�P-��_L��M�H��t7i7F<���8�__ڒ)ڈY(q�n4�iC������N]���7�_|�b�&���Zs��˻���e�銳�5>���4�Og�HX��l�b�*�x�?�����1S������~dZ�;N�wE��mAv���>���*ey�Y�M�m�� �!}0!"��A>�A�Y��n'<�#
�����ơ�pp�tJ�����vB&U!���8�D&��p��*�K�N�rޏqn���^��8Y������b~�a,�|�m`��
�uS��� ����N?�ɖ��'�_�'�
6U
o��w0�����*i��^�[��M�����|�v�s.���y����S�p8�т�����м�RCt]��ں��&�R�E�ʉ;R�4��PW�1Rk���2΋*Dyqw�t��f,��?,Z�qZ�%P�w/	u���%�]��_����!h(}����������t0�]� ؕ�u��J,hvm1L��%d�֚R'��ײ{�\g3�7�{K�[}Q�N!vV�gM6��z�{ª�d��8�ᕆL��5	���Lj�m[|��@~l������cw�E#��U��e��_S6q&<��2??L�ׂƕX�=z�{њ][v?��e;jkZ��*���r/yR]1j[�-�s�O!��2��߿0������ԁ~)��'D����m�-p	�V_�~IHr �D��?vs�`[�p\ ��r&pڛF�����r�m%t�D��l�Aҟ0R~��KE�iY��f��&f������RyO�EcX45c1�x��hJ�NK
m�ש�d�+�~�`힃{�SGA}��דPπI��a4ڳ�۳��T䚉 �~����@<$�u�:q�?�NM�z�W�O���}�hpH��=2&�En�j+*���G�[�jQ�O�Vi��~��хΰ��O%��1JNtQިi[��yԙ[?n>�j�΅��St�x�F�Bi�"��l�XO�����I]?_M�u�_�9Q��Vk�+.P�0�F��=]��KՙT$�6fa<�~AaC�YY3w�z��P��9g/�+�Χ����k��d�,�N�k��~-'J]:����Vq�	��&k]�(��0~L�|8��D6�[]xI*�?c𠛡� Y[%ƥ'O�Ӈf�@y�m��A{��v��B�LVr�^x�b���4n\�����%َ��cWS�)�ѫ�"���S�b��u|�P�(@+���(�BF��*_(� c��z(�(㗶�3 �O%	;������_�
��`ޢ=��0��tX�^@��><k�UF�*L����
*�Q�K�5� ��%�������\/��ȳ���
�}���H�5�9 k#�u�3��Bf�p�\�6���
,�,�٩C	��B�����:p2Q,ə��@"�h�\:���?`��;:�(�A�'&k������8*����Dz��Q�+�o$�9Ҙ��H�I[|��l/S�}��S�s��;B�z����@��c�� ɘK��[]��N׳�u�_�� ���5n
�B�Ҙ���(�e��P⿟���?��}���H�N�,ͦ�޶����lRA��TVOb�7������X{���X`q���,X!���Њ��tX�\X�PW��K���ױ۹~�j��ab :�v ���K[5=���U�G����yޅ��D/����龗�V�K���a�� XW#��9��֯$��A`��qc�^=��z0n���.EAB�-A3�*��R���_��l�1�ZEQ���{�@���� ���fv�K<ʥ-hoP�Je�
��}���H��@#�P����r�,��yi�R	�c1��4�$FOf��ӎ��ī�(�tEm�6*~0ѧ%:�a��3cx��;�q��P�I`��_�9X���Fח�e�H}>BP
k'5����M���Xh !Ļ71&�%���{�ѻgb�}c��[Tu���xhZ3������l|ʂ���ѻ�`�����[�S��i�4�8;���~
�%���5���������}uP�/<��vEZZ�B_��+���=����<��b�-��Lh'�L���G,E�z����B�T�
��8����xp��7E��U�xnc���^$|<涛:�� ����1'�#�x��4�,Q���΍C�אԾ�aF�(	�-��5�����Ya��ŷ��O��e���HepW��l8��0�щ�1"���",�>I��Q�6S�<JZz������Cbmc˃hcłs׏U!�2�,S�
Q�j��~Z�"x-���]��`L.�V<�᷵��*@mV�L֤�W��7=moGa椢��H�r���2tsn5�2W��1_딉)C�
�z�I��4V�!,-�
�M��)��>��Vqp���`��!���]L/kW�f-e��8ZY'$�����4Y�hXı���_FQ����t��7��)��:lO�>���qؙ��O5���5Ӯ��7,n0c��	J?����m'%�H]�wᒜ�ӿ���(�xZ&���/K�?V��G�6�o�� �圦,��|>E���v�XIBB� ;UK��pF1�����M��)���d��(�h1�����xp�$�p�[�T%u -)j�ؘ�A��E�e�e�(��^,p��Y�_��9y�+f�\=f̯�� s�X��Ɂ��h�g�nR.a�Oǋc'�=�R�$h�۞~�7�)V3|%B\%�C Bf���
}՟i^B�x�Z/���l���+c��g��S�.��52���OJ�(�c%��������N-�w؈7=��Zd�L�hـ�p@mP����͎K�%U�|^c�����?Ub#}�����D[ް޹P9�=��� ���uʪ�ˑ�����!�8�T1v�X�8i�;E��>��3r�z�Y�X&X:I��8�9�w�����7Sh�&�u���;�_�:��dV��nJ�~)�,NE�~��$f��^���n�x؎�]�þ=ޣꉿ3f`���E �/�c�=�-�c?�X��z�H�Ïh��uB���u��,	4�G���l�^��W�n�H���w�s�����lT��2"|x\]A�v�s����ٰm�䳘Pē����`����M��&�Y�p���_�R�9����ni���\�D9��zrT�A6�Do�"GL��(o�*�+χ�qr��a#���d��Ao��2P�Xץ�<J���n��������Qi��#И!Y�q`:&�
ܥ3g���c�n�Ѩ�jEjsfA�-5.�C�X|��KG)�X
��Jc�#�f= ����[@r�9{@3�L��Cx �y�H(��wx��՗���zcc��堩�\~�T�#0.s���)�Z5��X�5=��nB�=�"�S!��!$�"�=����Y ��+㓮����&�^F�j��V�M"	d�O(R3��"{�MY	~��ͩ�፴S����ŭ��P~[�'WG�9�1²�b6���Eҏ)��̓-� ��6PT�`1�Ȯ�,���1��� �ڂ��¾e�`�oCT4�N��������x� �3��:�`�3w�S�^�TK���>�׍Y2Ҹ�C��y�5�wCp�z��%�{�Đ�[�H�$�D^���#�ݑ��g����b��C�Y@��'8��H{S����f�q�'��A��Jy�=S1⼬s�	?"(����wX�D$�*ɣ��/C0
o��`s
��H��'�g�@�e�;����A]_�t���/�?ɿL��a�Ϲw��I��/U嘜�{@�H��T 4��E2v�Ϛ��Շ ��n�R?Sn��e6%52��g��b������׫�Q���2��mq�����(������}��b�����)� ���lB �Ll�#y�+�e�y���n<�u�Y����sϩ~YɎ�Ყ\ؐ���$�q{J�p�sT5�t�
���$�Q"H6m��6ɑ�RKs�Θ+������R'i��$��of��BJ��uM����W@�V_SG����݈��^�M��b #ùJ�T��7 q��:��n|xT�_��mhe�HvweJ 䐜�*Ȥ`"��A$tg���j�V[����"�)�������w��N�?�1[�x�yɘ.N�-��<�p���	gvs I�R%V�"��Ceb4��<$3NS�����Z_��+��j���#?Q��uE�cP7"���FҴ�*trWZ�M�`�堈���J��D��W��)��W��j�S`��U��z���h�4����j#-��FJ�co ��>�;9LT�"XO�����+�Ih����=�c)l6�j'�xܗ��*)���KT�؋Sb%M'?rh�6i��i+�!��Ѧ��	BHJp�4����n�vwэ�g<�f<��>,��&H?~�7��MW��=��[-&]|��	1�G����z!�@C��}�@O5�߮dxe�c]��?1����ۼi�s��]��ԏ�+�M5�5��%_~:�]��A{
��,����%�7<lڽ�5��Ln���wfc�t�ش��i���_��X�ޱ����~<;�?�k.��LZ��#d1K����p��v��v[er�����Q��"��3�����*�q��%蠎�AW-�JK��v�����Vɠ-�9R�g�I�B�MY�����66�+����%��B�-U�I̅��?��F%g�}�`6�ȃs�%�L4	�{�%�C�Ա9S�Z6:�U��'�S��怌54�$+v�i��i<N���A��˝'�ȐK��� ���b�I?�9II�A��v����~��8��
��ܼ��(ؠѣcV������܍kH$�fZZ��=~޼#��Gq&AB��>� �,2�r|�P��.�L��ab��D5|99����F�W���Fo(HOVeF$��U�����nB
���u��ިX3&D�J��S±��'�u��Bx!�g�}X�&F�V���|nĪ��x6���d�x<���l��B�����ox�wS�̕rA��ʦ�2�$�ȇ��heK�9%p�`2�Xno-����!*���tx
�]99;P����p�^��M87*��&JyHYLB�.�K�N��6/L��o���o��P�PD�-�j68�LGG�wȓ�~@�2�#��4R��LZ�-�[�ǳ+�SO%-�����1�=N@�J�^~eJ�n7X�j)�j�>�F�ۍ �:IC�����\GO�~3s��p ��iZmM��0��L�y���=N.��ݺM�$zt�o����2��ݲ@UhXlT�M��trtv��l����
�sd�X�_��n�����L���wr=�-ߠg@�饿3�ʬ-�n�u���g|p��/��%NU���Lhf2��":k���3h����R�F��S�.���NM���%�|Ԋ�M{4�[���åϞJu��(�LO&Tt�lI��=�>��4f���ل��g��j�2�/����Roy���6��;�!o���x�j@��+��+[E�͘�"}�bX�ÊՒĊsC����i�����H��?X�x U��81��4Զ���7�M	�;pX�Wɒ��%7~K:����������?L0N{�G�pY�����ľw4�w�}��G��4�̸�����W���*�kA<�5���u�� �Ml��aBB�
�����c�c5)�kCB���RKT���V촻~����*�ľ44*����
s�G�*�00􂷱�
�3<���>����g�2��rR�	/E��t�
����)�[N���?�5kVf�o14���d��k��z.
ʃ��!6zQ#���XD�勛l���:=���C1!:g��W!���l���!�h����d�{x�tk=�(<�bJ�b�.�5=&_�u��w�`�TE��qul~
/q~OKe,g/J���h�ET��^t�u�v���ب��%[ ��<��,ٰ�sS}��j� �Í�A
�
~���Q`N��N5��|9�7��!d�߸~��#<�ƈ��PjuU� ؽcجj�a��d#%�u�Є�)9L�1�:�m���M�@��鮽��J� gl�yپw=�XM�pz�a�3�Ȫ����������j+�,�_����Z�:h���iݓr���=,��`�7́!q�W�R�_�,�Ʌ[���姫@`����_�r-��r��c���r�]��(l��l
7�۠P�&Q��d��51_�a�,�)8��������c� .&@�k�I��8��A�|:sx����db�E.��&/�N�GHEr]�&����� U���%5)bl~��v�k�j+�m
?��,�i$���=�B��r���u��t���7k*� �l4�?こ� Sݫg=�b����Ğbv��X��>�r�źp��������4�p�� ��ڰ��ho������������<�����#X!�v̻�j"(ݓ*�V���ƈ,A��E4V�0`'�����'*x��G�v�
3w��s]ls�ME&^���:�}�b��Wk�sT�(ʑn�������W��]���,�a�8�ݝ���溱uG+�vĸ��k�x^���8&l��G�ȭ����l�T�Ӎ��<I��CGP�;���Z�p,W��z`1����W�*H/s��%��/��']a^�6<�n����엖qĕU�o�@]������f�7P@��2�㿒�C%���#i��peZ�89C)�?�����1^��*��SS_j�er](iZ�(�'��)ؿ"<����U�i�b>�q�qRL�|J���R�8��+���l�����,$��[z��h��X>�>��oM��=j��?4�$�R冁l���1M5Wm3Bx,���ĨS��;� ݿ6G�:���,��*�!@�G��&T�t�7BG�5��EN*��s�T��)2�!}`�ͽ�`�_25��Ph�k�\��{�w��T�km;4;�7��eDD~T����?��ʌ[�t��vɸ�-ե�z�p�ͳ�G��_�dƦ`��֗��z48���pW����7�9��d��w���b�U{����u5#���J4��@w���:!���H�{U�*2F2�CY���l��5�H��������t��qfA�(�����L��"�#��&'�Q	�g����~��э`��O3�yY) �Sd��Х#;o,��zb\E����{^��D����(���a�Hb@"�$��9�ϋ��z3�oO��oX���[��|�C���<~�(`���	W1��qYȢ��I��վRc蛏8���P��K���SBd'����B����>x�zE� 
�P������?�T=HvT=-7@[+�6I|����x�Cj-!�@���+�i��c�Ƚ��E�!���|��^^͹��K�>_8s�	vF��+�ާF��|�L���r2�񛰕�۶�[B=cߧyD�����c��b6u;:O�0��Fu�Nɥ5���o�\ޖ!��L�3���#�����V����M���w!o���k{��i�~RZL]?pAx�I;h-մ�����8+�7'n��-��竎���x��/��9s?j����A��C��E� �o*��xAS��Ȭ<9�}#��}�O�ɏ���o3�sM�<�R�χ�Xg�!���t�7\�O�TΊ��z��ʷ�AizV��^g";|���X����e�T�0O���5|c����ʴ��-X8�а��Vw[Di ~iQ9�[�2Z��e���'	RC�V�	W&~u��^��M��������>@��� ]Xx$Cn]���8�76��8�2���S�E;�ͼ�X�Z�OW����= eI�g@��٦��V���,�f(�^LJY߅�j�ʐ�>]w��_�����7UJ�����k�����C$��7��Ľ�rup��R���X�PV��Q�BH(��g�<wjA���.G-�~c�FlyU v@Ӓ>�4d�lWC��8�-T�MZj:���5�{�5Ӟ���9f��ߕ�i��{%�~:.�?����0U[<;XV�'�T�s;�1r�v��q"l�Gp֜�}�}<�!A���'�;X�u�3�����̊(%��f5&��V��\�k��� zA��y�l�@}��U�9���ɬK��u��	cVA����n(��b�jG��ό�i쉃�&�[�7� ��:"�1}G�u͕�5o����T���m��4��-W����h�Ǵ���ԍh��cZ�����q�(�����0�@�"������4��,�ͧxR��&G;��L'���[��Yb~�B�G�.V2-���M/'K� �J�	,���/���b��'];t�`l[{!��ս�k���A�9�X<�)����ʝT��@p㕶�1�.(��H�\�uԑ��]��3�묻Xd��|&DS,�����X�@[u}��ћ��a�������lH�T�K ���W�ؿɆ���5>ƾ��"�k+�9B����!��T#�ΰ�q@J�St4�c��^-׽�#ӡ�ȃ��7�am�"��y���蒓'��M?��2�-'���Yp��Y�>��j������Sq����jZ/p��87H?Oi�d˟P��9���e�Q�c\� m��v�/�>GJ���[����ߴ48��ϣ��=��|I��Ar�;��+-y,���M�P�?��|�G��^����(�a+U
R|mm���l+vʩ�������'< Z���w^?{��;�*��6�v��T*�OW@=��=b��m����u[�1L�m���%�wi�传�o�w/d�ͦLH�7ӗFp�DՐ�����:����+:2����	Sw5ej�=�����ΊBI��O���$���|�=�7�^(�m�T�iv���O����i�΋�(D�aB�y�>�F�n�C�{z;BV=r.��w�h�(6�+��Rޟ�����.�5am�zsR�R>k��W����B����G���>d5��
�3���Eu��|�k�����$o��?�MQ�:ҿ]���'��2$�fk���ֻ� ̧���E���Iy����5z(h���H ��/x�%i��Ua���~��M��'����Z�t���ȩ�|�ma2y�6%����Y����)hT]�b1�\��j�-��'4�Z���U�(CE��ƽ�jw�fxQ���,���3��Y����P�s,�d�KÇg�g�5D�7ݘaV����m#���l�f�8�,�r�M҃R�gn�l{p��D�x�rM��]8|q���,��
�s��[�*�#^�R�{�&DfL�/�\��h�s��Q�[��r����9F:z�^:xkر��ٙ,�^��Ë�:��$����\��zP/�ۢ�H��j��TG�[�KG_��� S�k��9(�����1ĕen���1!��ޤ�h��e'�X?����T��FCݎm�,!+(���(\���_�F#���9O�@���Me$c
���s`;�Q��!Xc�6�޽b��a7H�Ju�qQ�>���ߧ$��t��em�1�~���e�+�7Y��^v��PȺ��e��O��(�����}w�����>�?�R6K?z�7���c���IW�3#�~E,�]����#�9��Ҋ�I�X������=�&�ﷻ�jϜ]q�?̞�c��-sԔ:����6�2o�(@Z=�ׂ����DF�W��1������w8�����j9`!�]�Pe�Q�TL�rIh�@Y|��X��4� ؿ�R���dG7'}E ��	9N0���:Bd¾�g{�A��.Y/ɢ1:��73�\9�F0�/�S/�'����ʰ�$sy�.��f�� �(Vk�����ho�%��G�>0%r�uJ�G�����	�`�e���[�J���)c8M6�`����"�y�$��%�?��%�_ެa���+X	:#�Ԏ�sqNG)^�U׊%n:w��&*i�~��ĺ�r3~]L�^+���"����I��B�g��9r;@JZ���ޘK��~D)���a�}�$"����.��h8��k#<�������éŬ��y,rϑn��a�b�������(�@�45p$��M�B�R#r�E��G1��O��1��y�ք��9���?��#� ���	��?�5B���-�i'�0����=�f�~uٿ~���*3\m>^qp/%򺿗�=��B�l�Q��ɸ$���>�Ň�|��"����V�|!uEiq��b�n���r*��f,��aL=���
�Lx�R�dX����>�m.&]�v�O�>H���ȣ��Nґ��tD��ˋ����I�ʓ�=d��myP)dv��#��Y��^�y��
C z������gk��ǟ<Ȯ���ix�~y���v��c���,r�����J��xՕ��槫q�)9��gT7�a��@*:L��5�zj��r��bzCQ)�x�m,���x��:_�o��;�2��rQPCKI%�;�a˓���-����Y hr�©-��kS����NHK�������}���9�TE�#�A���E�%�Q?�]�x��e
�H�����m�w�Y�u��;H�u Ӧ[k\3��a
��¸�G�|W��r�U��(��҇��o\�Bp��#@r�K��&Ik�Ěf�����?ط*�N�Cy?����چ���R�eO��&�>m<���A܃{�Q����q�D,�h.K����
��i+� 츞Gj��o@�,�}��Θǯ2yc�J�RĽ�����%HK���UC���Y=��呚��@�	!<g~a��:�D��ړ9���*j��UW ����B$���x�T��Ԏ��k�:�`ݝ.wZ��{�|LS�JS%ق��ʿq���63�6�2�s�����Xܾ�
���%4�VmW}҈��-���»�U�Ϟ?�Nh����O`�k2� ��W�f��kVFu6�ܻcCsez����E�j�1I���ST�b�~I���$
ȬH{Z[H�l7�_���ouY���#�;�X.Y�N�	����x�,�ʤ w�*UxA�l���t�J���ƈC:��H@u�h��0)xW��<��A�)�2E��"&�׏�#��1���{�~Vj�A�U�%�̮<M�D����EY�Rt���.aK�ɦ#�c��/��su�
����$I�d��Fa�*�^�uX�M_���V�P��3��d �q�^.\ ���hZUM��^����;�S.�M�&���I�n��֒���3,�p�^������ܧ���AC�����624�.�%���X��`Oq�Q�c��6=)2ΨY[�����<'���RLt�O��MeF�)%�E"�@}�&�����.U����!b�!�XSJ���(���>'sLK���%�߶GP���6�:7�x��5��W��]jWvT���}}8��8��;�ި_%�����z�U��;��"�iT6�Vڃ},��2�D�s��z��+F��|_�-5��f�@�3/�ԇ�P���15-�R��e*���x��]%�`��f_H+�W�Fu^֏�%�����KJ���)4^r��%�L�o���F��즥N�G1���D�ʏ.GŃ�a�0�7g½���O$g�xo>~c"؞=�Ғ=G�r&$Sʀ���!s3T͌�.cڙ�����/$�xP�Bߏ�S'Uw'�y�q�<���C;G�߬�����Ђi������#Y�
v�Ս��!G���[�����w7�|\u����R?���SK6%I��T"�f��?&�i��:7Ew�;�9���-��Ɠ>�씌F��:����������N��-6VI�P�(���h���V!�
���z��׏�nG��x�`Iz2Xu4��z�9�,�7�F '	*Vf/2�������`�f-�|-M��gw!�l�ԏh�y�p��f��̕�sfgfn��cS��ZI�y��#�*IQ�J���$���u����
���8F��m��Ѓb&�K��I��p�>rn�ȿ�]�wֵC�M���m�{=~�k�y�a�+s�����Q)$eh�`���S��+�v/��Su�,�����Gܲ��p���~�	r9���(��	$=ɢ�%�ǡ���h?��S��H�@��7�wUד�${84����r�&bP"�Y\'Miú���-p��3���(�1�s\@lPs_��3J�sK���K�UǣŻQ;�'�zz�	�3
8xE<:�#��5�\�:�[�+!뫱R����#=�~������>Q�<u��	n�aw֩���Ư� �wI�k&t(sl�P/J�Q��D]]���v-�K�ʣ �!o#q~:��[��h�ES�T�FgT�J�~Q Nͷ��2�WfW�p�D
�B%f{���X���W�bU�r�q)��*3��k�_����W�m⿐M��_������] �Ķ(/�3��4�֮� h�Z�o��*� ��n@���Nb����dtקt��>"X`��y �9�!�D2X%R���a1��@�p1�6k�"�8BNm�������D�䀃����B�����m�zOm����-�-�L��c�΄Ao9�=��N�W���l���>:�������&�Bs�^J���X�e��UyZ���_���UF9�!q�$+Ne�)�C�L�X�gF�S��5��1�'7�� bPn��y��A�e����Svv�>69�O������k��n?Ԩ[xd=>||-cX�ǡ��υc��E(�dI:�d*+�,
kl�1�z�%�Qx��mv�ߩ�_�m��}�1c���'�`MV0����bt��b?V�Ǵ4�/�@�MN]
�t��M�-�����;(�0�F�Yr�eEv��%>9P���8"`���d����R,��1�^�/��Z�:g�½7/�[�N�[��ZQ��w����L|ˮ�_�9zU��gg_��[ș Ym���������2.����%�q����ڗ)�].]�x��ܵЈCT�C�`����kz�B*����H�Me@XM�� _ |éم�)�n?i3E�P���U#� �E9�B��-�6r$N�LZ#<�BМ�=U�Nؓu�J��AI~�J�C�W���F����Cb�*���hNʁYU5Zy<0�C�ܚ��O/r�kw�P�EN�,�y=4��КY���f�;� :��b����w�x���E�c.�B��ݷ+EP�{��\P�~G��,e�8��Lc��.�̹���#	ߐ��'`��"�S�M��x�F���E3X	�}����F�-�<w	���óUGf�p�|�jµf����J�}dvD�vv�&����\Ը5�i���8r�2z��SAA�;�ɿ�Y�]���󶌼�D��ń�K�lk_3>Gd1��C���/�R���:�#5�M;�.��9@���7+�w=b����*�8��
�nUX�)����㉅>��g��I�TM#h.os���R*��R�2�6kqx�#%o4��0v#��M�E��G�FFJ���Իh�@�;}���P���E~k4f���k՛���Jv��G��iX>�6��za/>�}�{^K�t��	7��X�_�J]Zk	��,8㔕,ƺ������[&>��-����F��l'nQ^W6���(���!�z]|�e ��V����(�ㅸ�ɪhұ��h�Lu��2�����'�?p趒|D��-pfF �AM ��}��Lʉ�zA�aN�^P�iZb��eRMPå�ϾduA[��U�Rm:h��֥;
���Z�����|�S�3��P���T%��W���%Q� ��t���b��lZ�<�p,�r]�q�% C�V�dp\vi�b�d����{c+����(�5�4�C./�H
'W�`����Twa��:ҿ�?��D����B��/ߦ:�&Ή*g���V<��+���Go/&�mg+�7���S��GH���_|3�v��J�`�pW�a�~����R�5?M1�g-��}���%@3�F+v�\׼'D�M�`�b-�����[�i�,>����Sg��Q�AR�O>���O�ȝ� H��aT���sQ���<�ໃ.L��B+��\���7��*�.��Sv����.���̿B�CV/L��8Fb��:)����	2�
�0���J� 39�*Pa�m���T��� ZO��w�K�eh�UK�}� �Wu+})p�JC]��/`�u� ����K]�oVVT�����c�����R^�%�籪��:����7fD_�;[s���fB�1Usv�)�{����52�O �7s�<mS�]c����}�C� ��73�f�r����o�-^0[��>Pf"�=��&.��g5A��]���}����]��{M#9`�H�f� Oz�H3�A�{U�	
�k|��ֹ(R���RP����2�*p�=%�m�+`��f1U�1E��4�8XTƝ�D��s��%�%��s�&�nXpa������>]����'��Х�EU�������@��$�y�B%�YO(��1Bz#�im��N��h��XV.��x��NQ&��j��_�EMiෆ_��d��Q5�(r�߮�qs��~����<=�4Aah�%ʔ&��M'B5_*ol ������]D
��Lf2=��O�
i�AM�g�>��؋�w{�s%C~��8,�x����Ԕ�#�F��*���T����mz-F/�QCXB���x�V�J{�{�	:��W����fq�+A�<��׻����.Z�#i�~�uZe��rN�҃�Q
���s���K�s�]Ƶ#ށ�嚙g=桐�y�]�D���ǤW�SGA�0q��Ĝ3c��Hyn0��pj�T.��ʤ(&iZ��V���#�Qn-�wv��G�s# �r�5y����0�\�=�zLX����_g�Ύ���e@��e)^�H���{�΄�ݼ�c�qJ!�������uM�J���I�l��Ý��狀ߨk{��w(��A��塪`^O�7m��_d?��c�y�;�l���Z�;����Q��N@c��M�8c����B��M���d�H�Of��\17!ɛf�g�#�Oh�1&$�	��8��������^O�%�R�ɸ�P�Α������]࿜y1F}�nr��zbR#b��\
:�I�~-�]:,�]("x�;�=��x t_17|P=���	q�2`��e����2� rZx�V�颉�:|%m��p�����~��D" J�;ўJ�s㔋]��E�����X�O@���L�W�r�v̭N�<Rᜲ�93�e8~#�8$<��m�&�7�?@v��{���9ouX8{���2�2�mE*O������nQ6�.��I�ޣ�W���D��A��s��4��d�2��tuQwe8�qw��ZmW�/�IrI����.)k|A���kJ��Ԉ�;��ĥ=��eJ�� �\��4�&솞�P����Po�)��~�����T�d/i���~��?�Hql�i��=��ɶҹo�&Ƥ�rl������:`,��AHY��7*`J�����O�����kJn�[ m�2s�گ��4�@W�ŀ�5x��!"��*of[/r��օJ����v������@{�0{��p��~��� FƠO��-��Z��W~Y^ĂoڲQ��C��8J����C4���PT�Vy4�`�!E�X>m�Hn��AF��4\t������|�������[�~��k�rx	ˣ��:�Ѵ+b�?1<��/pu��4]T�H�7/ɚ�`���c�����b��t�Z�$��{���qe-�V����t=Ȑ ����xtm״�!t���Z�du��y��X��5p�y�`��R��:#�
�@��p�D%d��*
�����?E�2���+6���M�@hڃ��@?YN�A��t��*�S�ךU}�P;_����ʹ��D�'�����s����s��'��[�-g4]"�N5���t���H�8F�AY��\��p�I����� oyJ��Ҵ4�������x��߽�{T��w�[X�,���r*kaZ���� jMT
	��\�y�ړ5f�e kU흄��U���ɸ��hT;�6��}�s	��>!X���KlL �k���W�_'_z���(#J힯������-l�n[��Qp�'�W�j9������4�o�;wg��z� ��<�"��(	���X�)�<U�po��a>���U :ɂ��V�H�nck�t�W��u�_�3�u�
(��	s%�ڛτ�A��K���<[��AHp�Em�&X��ujO��{�L�������큙���b?�2��L�)cAl�_mG������o�a���Ջ����0g�]��C�T�7��]��7V�h_>��α*��ԴaZ��X3V���1�8I\��D�c�Tߧ�·�T�I)��C�I<-3r"�;
�oz���ٍ�\��u�}V�	�L��Ƶm�Fɇ��n{5�2�r�}L]l����-�y	nl1�uB"� �8`�U����єw��x�T2�̝�:iK��}�(}A�Ku~/�e���e�F�L1�v-�N��/��V�u>`�ƾ� >���"����}l�٣#�A�iL��K?4q�^�^���x�uMb���O4���lS���I�&�'�^�4�+��n�P�J4�.T�W��3�)�@�,]m��DQ@܎�'m*j�f1�{����T�P/��lhk�yػ�&�����4��t��}}lz��q֝�"P^��͟tE�Uo�]��Y�!�&ءQv��Gĵ������J�M���e DkfB�=��,^�Q��0{��y�n�LBC�z|W*�Q�L­���g���yb�pb��/
�������H��(�+1N
]B�y���#}^�=÷�7䞍��1��/�#�6�
�0O��ThP9l&�-s/�#.���{����S�7�\����ĳH��zMI@/Tzc�exo�΁�߆4�,��Ԕ��$=�}T1O�B	l���Z�.&�@㫖�_�B�4[8�ꚬ3�*dq��/㟢�QG���Q�KnZ�ѧ#esi^�rnc�XZ�o�	�����m��@�S����'1���b���v�wvp��o@D1��N$�PK��0�457V��/$�5�ں�\��L
����l0īnO%|8mf/�w�����U�1v����t��.�+ami�ikL{]l���E(<�0mU�=n���� thiF\U�0=�������QѝWP!-�(shʹ����y=R��Ą�ᄫ�6�HN:{�3;Apw�[?%�+�;8W�r#����ˠ����b��-�Jj�w�������?�T��+�su%�8���76{�J����r�Z��u��QÄ}�O��in��#�!u�$�0%S�֭U4X�P�u���m]�1k���W.��8��W�U&1�����J�	�T���)���$쳬gk{��������Ge�3�B�l#zq=	ӡ���D�x�p���� fz�7,"���8�;��sg��m�k�P�A�<E��L��6�J������2���4�B(A��wk��N�1��_�ϣ��)|9�#�m�Q�{$�rS�-O�S�����(��7�c�jX�$�'��wh %e�C4�|Q��K�9��ag��f�Y�>-Vf�%�H$��l�|�v����q����߮�J<�(���saL�FS,y���{���{����fX��>�窢�1�L�D�_d�Ʈ��W�G~�+��	�j�C�zﱬ}�i� ��Sq�z�A���ʆ&����9���bS��� >Xn�_���lM<L;��t,.����!Ihg]28+<4`Q���Ti��ͻ� ��K	��,ƮN���,o��U�Er�&�o��
��34@b��
t��p������6�HDW7�s��Y�>�
M��r�lq�j�J��y�HgmtE�U3p�X��)<U��R�����1�F���On�4���Mc�ۢ>z7B�d�z@?'�¤=�!��nja��娘r��A�v��c
��
���:-���6��w-uV�(a�� ;��M�8W5�LX���$(\��j��uP�`.A�w�*P�����C�3*C0=9����Bw�|�h�0�ii����d*��Pg��wjtI��Zc)��f}O�.�~�宽
�/D�豘�d��^��''����n;�":̘�12�90�&�i'��y�c�hؗr�)������O�E���F_�T���� �刅�Ѿ�>e��w��6� �B�%�O�u��(��
/�U�R9/W�����<���Ԉ��T���<��[�(��D�����Y�k<E�S�����l�!��h	i�]�1���=Q�v����J
�� �.秤��Tk��Q�����S.�w_ܮ��Sg?�M�,�Fw"6`��Z
�4�V�X�#�� ������e����0]%�
��I2��� ؁KGE���2c�]���ɻ|��>��/�k:�Ԁ�1t���1��],ߩ��u���޵��@�йȰ_����&,ӥ]�Y�h<�*���ud�#w���k���I
�\=˨ɔ���ǽ��]��q�G�R|�=k��߄9A�����V���Ԣ���ΝM[�^x��/�x��1}�&��6RIb}-�Y��ΔD��'����s����N�!�!dAre�@����P`I?K��~������˯_ci�M����L�Ҡ�E��x�okv|�	�!���E��/�8�%GqmjJ/�|$��@�JJqA�8,�%��00�>�J���m[e��Mg>/VT+oG�˟�fr�����#�I�a����P���%��n���Fx�9&�t�8�L���z4���_��`1?�(_�jC�Χ�-�X��dbk1ؒ�3�w=�W&"�W�\G���������,��6}!����ѕ��ǑW��>�ts���)�`�ʏE��B��Z�
�"Z�JB�C���������`F���m@7��7��}��w�\�����;O�R�>���X�d��򬕺�2x��X��]�R0w/ç���y�)@�������g-⏩�j:�MkU�rM��M���"J�	$�<���,#g���2UK®h�֔� ���d�ݎ��f,Y��˶��9�X�@!ڴ[x�����]��º`�2�G����f[rf��������,���唙��9�D5�z�J円		q!�69�MOd��ݜ X?d��`�W;H��=M-~b��2 �@'��׮�Fs�{Z09�z��R2��ÄbnO�����@��y�P����E�7��<��5�۽kZ�h�/�@
����ļ�I��OB}#�Zz��n+�Ǖ4��qj��
�$!�f%"�~��-���GA��~"r�����K���'��oW38zA��S}F�M�����!��@V��2(�B���X�;�a�	BO��'s�ֹ(D�ҟ�U._� �����?��M�Ee�<�?sG�MW(L3FX��1�7�|�S=�������L*��SfǁQ���
��N��pu\��'��R���+�0�'���v{O�sC�C0[1�e�e�1<x!�Ҭ���C�@�n����m��=�~��e��Ṵ��e��}���=V���k�g�"7�_�!�D��o�WcŞ���{_
���>��2��3�����h�yZ���g<�W!� �x��Q�h-�����L@l�7P�HUr1��Or$ˢG��*G���E���-'�a����ur4�M-;�~��mW�Y��,�B�S���N)�ѿ�[�%�Ʋ%y�g�l_����K-�T?��<p�12[N.�q��e�c��}�E��}���*Ǡ�#DC�d��˲�����%�撱>$h�+�v
t�a��〚����,h
p,���"s-!71�|���JO��T��J���Iq�Z�u�&x���>�}9��ܜ����F;�������43��p��
���6R����Ƥ�]��pi0�w��0cLk(����ʎ���͗Z�Z)��%},��U����Q@����[��3S�Ӕ�	�O��-{�0�wc���=Np�/P9"=4-�q(~�r��o�!��ڧ�OG�D��[����7���ۊ���y�$%�.K<&�}��)ہ������PR�@	D���KHJ�!�Q�n�+xZ�4~Yo]�E�O�;-4g#�)�d^�X�egB=�� (�I����t�ԥkBc�A��Jl��sr�0��>X*�In��/���*1�Kkџ�S�Ӈ"�[��)?�|c`H���;���m�����W��n-�VPol��Y�Bï�0x0�N<�y*"�d����T�Ő��t��N��Ư�]p��ג��f� )�В�!'�>�g�yT�:���`���� U�H���x����bΟ�}��6���?���E��?��]�
�n5] �ZyqT�OQ�0�J���#F�J3�a>E�~hx�m���帼�2���'Z;T*��\�Q��F� a�a������ȗ�DF����UBp���gaw��uVѴ�4���0�������uI�
^q���A�3��Ǧcw��{��O��7h#�ʹP#�=�P��u�ǘm��e}��!���Q�$VG����RG
Z��*����]�>$Z}n��m�j>��E�Y@/���mH��Ȓ:oh��ug���˗w��}+�ԕ��k������+.��f4 m!�e�N�> D|A$ .��_o��9��j>�x�e#(��:��f�M����Q���t{�����)QJpwY�T���	�7��>� �tYd+�)�rB7��jIXٱ���
�����n�-����vB0�&Y�d4O��x{�[�C`�H'?�*b�'�o����-�"(� �J�ˢH(�j�
q�&���>�(�I3E���1�Uq����֥�W�(.4������R� IG�n�t3�~ߛ�	V�7WD^ ��ľ�8��p���|�(Í9u�9ʃ�([��:�����_�Co����le�=t24��uN� &��fˇ�"�һpag���j)uK,�iv ť��
�(Z=��v).�k���tN�@�|	�-�������E��m�}�7#}�u�_ �����7kfc;`�m�%%u�Q���}��j���s�tAh�[��� :�)u��Ě2���@��/��ҾF�q3$�M�E��Pn�ѯ㴴�	L�_+&uFrK��Z��������^kX�O��H����NC�2�w��:���UFG�u4�����h�����8�w�ɈrB#ȝ����ݲ�Ƃ���A�,r��� ������ �>�<�?�.�����vCe�쿨�
��d7-ǁ�`,����r3�'_}�%��7�J��^ޢ���K��_T!Ɵ\��) q��k�{߯���1�����}�����5�D0���,��i���)����6KM���n�o@���*����,�dq�j����)B��F��[��Ca��"Xo�m1k*�����L��.�1��S��Y��X�: 4�mp�R��e`����?dNT�yT-�/����VK�L9&�N�	K3AaУ�c��:��5��Z(I�יx��(�o%sI�ś�ЌCt��`�8!#�>bH%x/ ?n��b�BW�^�B��%�kWJ�n]���t��7��#�1Rw7�nB8V�0H����y �����.b+��i��<DtbO�>��~Ӿ"Af�ۻu5����#�u���v*���q�o��e��'�\6��.�Ҁ+Ds	� 
��B���Er�d;�<X�e��|�������*��8�z/Z�տr���e|!�H�K[�w��^,���kI��dH��f����~]F;Z3%-]�����-�H��V޷��G0����xn?�W�o��y#_�j U��誅!9C��g2��/A�k_o�i�Lݵf�˄/�{c�������A}���{Z���V���W���o����A��ݰ���K>P��@q]m��fpw��(��k+j͜��f��k��4+T���|̃D�LQ�z&������:pM�-*�a��s�� �)Z;-�B�S����=�{٫�
��.�rR�(�Sò�J.&
F�"���D �]�p��[c�������(�y�Bs�����yy����N ^Q=�u��_�� �]�iǏ�.��|��6�w��O>Fi�ie�-��:.�@��2�7��imwc�[D"�C��|%��H��/�Gg�9���K�Q2�jz]&�ڊ����oV?@i�c�tȧӹ!!�n�}���:��V|a�LǗ-�j��?Cp_qmg����x��_��䐅�=��Br�h*�k��,Nk�ǥV���<�-��V��@��;z9�)˪��c�BQY��������A�����/|f{�Yh�{=�f�KH:;OL- ��!�	!��7M�=[��?�~d�ց�hP����ܽҚ��YI�~t>���A@�=�1.u�>{�y�3G"bK�z� ��
�BU0�6x�}�~�LG�%3�^(Ğ̦~_�um�y)b�d�}�%k��i�br@q����H-�X���@e�³��f�*J�b���q�_��H�c$~�H�9���(F�d�PJut�g�P6ע��r�Ȱ4��_�ڙn�K|����B'����ѥ����$���L��B-��<뺉�,7/jؖfOV��j�H���k�[���9):"�	��f;ʁ�s�����?)��u9�mf��?枽Sɳe)����P�2����Kvr��~.���8G����}�4c!Q:Mi�!�v�e��	��*�� � �~,�K����n�3&�j�;X�9��Ĺ�_��D1��K��]�7���C}x��x��1GB|T�Xh�4��OU��0i�y��IMj)Y�R'Aڕ�L1�k�N��_^�]���ټ�iJ�`[�CW���p��[�r"`38<I�w-[�ہMv�"�b��ZG ��y�M�=�Й�q�rMr�	"f�*�j���3��m�_��ʞ�m-����ԫ����t�lp����u���-�����y6ԛ�#���5K%�����1 ��T�/y ��M�.�Pg���v�@|c/��S k�T�m� ���5J��~�%�9v��bF���(�4� �2Tq�=� �D���
���V���f אn>���z�F�Yϻ∛�}�P���X�A�J��%�>2r������v������"l��t�n7���1�3gB�"�{U/�i&��mz�#�(��-?��H�,_��=�>�p2`�i(�wg�(�rP���'���ݎ��_g���;��v-�}Р�Pː�fa��9������5�	V}��4�����w����M������fz/@F�Õ�ٌ��#�����ӌ�Ȗ� V���G �,�̫4��("Z�kb.ZT���
���.�������c����\V�Ec�-�"W��b���
|YK����+SN��4<�Uݰ��g	*ݤ�31��袊�vԪ6�q�Ca���3�=����"�ܒ�L1PPAs�hr:oAU��a3���h|�B�n9x��wm�>:��>'�w�р��\�t	8�~��,�A�O���?X�4N�u��9��>8��?Z&wn�A��ѸY�9��uR�͝�ޙrkh03����W��1��l�x�$)WY�����I��q�q �L,��!=Up���F���ą�j)vīg�S��Bs���J
��k��y��Ŧ@�p�^�'���-�ʡ�sx_�=��s�n/�� t��1���˫[P�P�H��Z�._;��ԃ0�}T�/)�E�,pb�1�R&g�ɴ��
�'d'vr
�i9��t5=�^����x�;\�@uw��o:�������-Z��������P�҆�(��7@��7�&�K�������#�BYB�B��n!r����S.�r��zs��	���-�)d�z��wsvQ��WxY�y�s�+0��^I��S/�����D4�4T���T��Z+-周�G}�M��	Y#���z1E�;61[�8��(��CGmr�d4Po,�C3H��9'�̢z���Z����+v���\���n	BUf4�Y l�(A�Џ?�{��m�B�Aॿӣ6��{\�>u,xx���3f�U>���<ш�E���*'ڔtA�{�!.�� � W��T7�M��7m���y�7BF6+=B �����mP  �)�'���5.��S*&���QI�3� �[��i  6B� ��|��������cO������G	��C*����G��o���3��)��t �BmH��Tq޷�����7p.�� ����!�_�w_�_�ڨ����+:a�v��Jspe��A�G�Zfm��5�������?�P%i�0(%��u�);U9��:h�8�c1�X���ۻ]>�����V0��@�l�����s$T�uQ�hp��Du(vsa�A�Xԛ�O��٨���jk�ō)�V����͌�.��pCL�#�4��&�����w�6Ǚ��Z1׭�'}`�➛݉�����t����Ҝ0��=z�_���ŵRդ�l|�)�5��r	A�BF�+��[�����s"��P��R*�7�P|"��k��qM�+�s"�9���|��+K�^�b[C�����^��9H���'�����8�[�vL)Nǧ���)Be�sPOu�.�Q��`�%��0��ആc�����KK?8�Ve�r3k�W��ץ`����16LB�kE@��F4�_�v���Ιa7T}�6�>�`��TO6�X9���q{e�&�\NT���35/�Y�|�G|n������HU�J�C�)����8�KE���}3���~FqY�_�1��˹�����฽8���
�RA����ͺ��h6�S��OYtp�eaA��H}�Q��8�����,�򑃾���#�(D6��պU=��� po���%{��mD���UfS8��w_\���A�t�P��6&<��t2Cx�h���*��~W���s�3'��8>�R����\�0�C��[%��ji1�=>ܩ��i�o}���̐�ߘ�b�i�T��Z�V.^!����"i�D����GC� �}���6��ot^���fxsrk�k��s�U�sa!���-F9�˄�A_�rzU>82^�+��ݢ�q�Bo�B����.�V'��a�]�$�����b�0��:Q#D�zð"L=	o��#�J�ո�{���qH���!���-i�磵�����ۿc_E����Y^?�A��"�ρ4�E���l�)��d���y\Ż�m�������Bc<s��"��w�.N�&��V��t�0�i�Sȼ�it����m��G���׻�>���Rm�@1�]����Qj\����l���Wf�{F�����������H0��'47.>��o}�ծ�!#䴢@����o�H�\���.��&^���ʣ���?>W>��n��	���⟪�K1��PP�4��&������PɈ|0u=_�\�f�7.�~´��N��ʏ�s"	ǼT7V�0�L0�5 ӽЇ�B� �b�-�M(��!2+�3Y�` ��i{�����K���7���M����=��9�8{yx�_Ș���o�v����˟(e�S1�Uщ�;�Nk��@��^�t׭M< H9^܄������l�J�*徕ȱL˱a,0�-�>zR!GOY(�+W�dͤ>
��a(ZdW�4B�m��;2wC̒��ƻ]���p��%F�*ʀR!���h5�P3�ܨܔ�P��p��9k3�A;͸�[eE�������L��w�~K�DfF����E�p���)�]�2�+�%.P�R���Mz=d�Rg�����A@[� q��b̃@zQ���#ݸ61�qEde Y�xHl�1�H����M�~/�<_���B3�%�\�s7*�<�wX���5�����D���
�����f��X���r�L�!���D{�p�Y� ��ڣ}�!,`A^4j$>ֲ(�8�E �H�?�j`�M���@����I������ڊ�V�s�F��=�
y7�����[C���g�V/ȍk��
�E�p6/ҧ���K�U�#��s�gm}d� �g�/)%�L�rD����!X�%��Kf�q/~u����
�5�k�nnM�h��y��|����#8�-�Q&�:�/S����ڣ�<Yb��t���/��)`&U0�S�V���^v!w4 �V��.@0M)g�����
�$�D�A�jW���p��U���#�L�Ep�`+R׸o���Ll>���W�{N�P���֣����Kur�,��6��a!�U��{f%A���@�}��#�'W[.��P-ӿ^@,,Y�=�ʽ|lO�;�=�yDBI�I�JI��t��3M�Yv�K6
e0q
����qt��q���w�(Sa��&��J�0'F��뺥r~J;�ͳ���6IN��So�ٳ|��e\��3R^q�f��`�848?��$�&��A�?>��p&3�&+���?�{T���TFA�y���%��9��dt*2��T0���ϣ>�ՄҪ����W�F���@��<F�sz��Y��a��ϲ��(�i(S�GU�m��w$c(R���`/�� ��H��l�d�Dz(��6w:���S��iEEE�p?���F/�6a�u��8J���=�������� 1b�L�K����-�b(,�L3��fBY3Y9`N�%� ��4y��k�v���5C�r��0���䐄�u���>G��l���fYoN��E�x,���4fc��@(��,�#�/��a���v�s93�������p�I�`��N'�JG�� �]�;�?�����،���g�%�-�|(��j� v� �4i����N=UM�?��`,�w�����+j �6}JH~L��_�+,=\W����<PM�5��iߡZ��,
�6�(� �G:�h��d�z�l�Z)[�nr�ut�3����l>�S��$K��Wy1�pXfΩ,��"�p��OMj�v6X?T�D���ɉңPa��1YC��p"�Gz(�#C��qL��P�U0^��r�~j5�)0T�H� �鵨zSn�GBj���,�Y�,*���)�@������?�-�P��H���d�!�%�un������I~���8C\U��u*��N����V ��|�}���I
qp:�ʃ�wlifC���4�j��7�@d����Gr�W4ڹe�&,҃J)�B�ₛW<����|��tU>g(E���'~���'"~�I������=16g��uc.d+b�J8��@Nr�ː��6� �bz�u�P�;��ą�tǇ.���� ��zN�4��gr�K�&Yp�<o�e�UCeӏhFS�5�R�Ŭ����?q��WV]1rD�
!��#w�KAG� VE�o
�ȟ��!�)�?��܌t����1��PX�yg9%�Z	h������9��Ć�����˖Gj�<z	���?��қ���y���i!�|1�̴Z9��2~#2l�����L�B0��S&~g�:4!̖�Wi��PHI����;������&X��xЊ�Q��1����'��uˋ�i��B�n��oO�v\���uVI�۶9Џ��8���UL!%Ù��2�E��~{P������<`���Aˮ��?_2q��Q$��q3-��zhI9�}��Q�j�_dUӍiT�38sk��%K��	�RJ����7R�,��i�E��J� ��_�jߺL�u�/�?m�᭟;�~F�,qO%D���&�c����˟.G���4C�=qf�;�#����t��KVѪL82I]�O��J�Q�<;z�&Ӓ�Q&��
�BDk��u��1v��^$:��������|�������hb�`7`n�$�%)��)֭��e�P��e\�@���#o`/*Õ[.��35k�V���0��L�	 �c��y�����ea�m%L��F��^�����Aʲq�Iy	)d+*2xذh����b��T
��ePQ��T��oA� ����t�˼�����pP�6�|%
`��I|�\��)���^� �7����O��4~^w}yS�TI�аk.$�ɥ�D{T��g�<B���X�$zKA��1�P<�,���s{k��#�(� j���x�y�J�]�F
���y��0���<�Y+�j�b�h��\���MSFt�������u���-���O�����>�Z�!�"0�%���JBK��A�W[����_d̙]��@Z����M]*�4}^J%�}�!G�`D5�I����KP�����o�@y��gx�p<D�gw�b����3��LJ���eB����S9�$��u���� �����@�a?���ނ�#!��O�#�'���d3x�y?n]<m�ɡ��]iR�X�ޥK7��cY�h*3�+.^�S��{�7<�ؽq��_i��t���0�ԑ���JjH�Z�~��HΛ�o������]��G�f#|R�\[���}NvR���ˏ��^���0�s�.��0i��6��� ��0�>�;�(�E�Eb��~������]��ޛ�R��Q�*e�a���j7�g��(ߪ��D)	S^6%r霷��SJ�֬*��R��}���m���&��� e^;�ϸH1��>�;6������fI35+��94]�����fh��lH|S���J�{7j����C�u��#�"�;S�K�n��[YpD<p�AI?�S@���Ë�6C9܉�ڙ�2vl}MN}Ú�hA>���W���bOoR����7,����#',�s@��=�0���7��٨�(nB��p�X?d� wL�#�@��{B�17��	�;}�'��n�0���>岦��S�ʱ[�7����t8*q����
�y��M�A�4t�w�*���<XB8��p"��iL�!��C�������$h��M�җ�/����=ӱ����\ߖ2i7X�xi�Z)��3�:�-�T�,j��A/L��hO�6R,@goLٻ�G���=�gPRI"�5�@y���ܬ�(��%l�:�V����6MF.,��J�DKw�\@VˀR�l�s���qK^[�.�7;���h��}pF%?�pȨ�ͷi���NEg;H���D&12LG}�=%��M��D�gl�Tc1x�$����l�(6�+Gk1���wE�Q�����?r�U�j2�:��Fk��f����:ɴ������,זv�V��s����h�S��5Gtx|��	���ŦZ�Ԑ�D�XN����k��fNl'w_*![�x���?��7��������N��7� ���iu��y��	274�F��i�yl���(�����e�K���Z�u������0g��l|svQ&��w�6P^�ً�Ń)�1�A�˩#�%���Ϫ��+����N��Z��\�2 �}MaKG�u��R~K�:S��N�o��SExywp�>A�,l��v9̃s��o�	��19=�@�|1H�Cq}�{W�9h��(���wxiC��è���c�Cc���3�� �!����J�Dn�du����n/�tO (=�H(B̄���{��ғ��E��u����͸5�)�Y�2�2���4pw��ՠe���nx��w;��^����bB«|UF���-��eq��,Hg�D��.��"����T�~�d�7��B�m�����\�N��<���Ҳ�.�UF
�:r�ԣIr�Z�4צ]��9�h<޷yW�R6�):�D~�j6q!'�O2;�7�󭄜���iR����Y&���KU����(�M�p�G�VȂ���ؽ(�F����zk."�Q���37
�|�S��'G|r�� �[�Z,��D*rɐA� ���Z�Ŗ���&�)�n��=���÷X�"�HZ%x�x�φ�0:#ˉ_�ՠy��f���B�_qC�Ï6�M��?���<��Z���T��]��v�+�1ؕ���ҭ����ĝ��@�a��Ζ�����F��X�̪��N�cP��g�,it T-��/
ŋ���}�l�sk7ؙr������b�6p}�"1���azz��x��FE���Q8_L�����Z���?�Xb4�]����a>\?��n��Mxmf�6�����䯂C���-�m츪��/�6W��SV��_22œ�`lbt�'=�F�N� ܁�!��C���p���A�Ak����6�E���XX���k���[�J�(� Ʊ�P�����&�c��H(�u��F�&|��	ݒ�3:(e�+�٧>����޷�Ҷ���?x}aw+�\AMI�?��ẁ����?�5 >��t9�n- ( �L��dy7:an/����NR��I:A]�ɇc�1�f�������o��u!��t���O�Xr|�*a��<՛q:�)�$s>A�=C���BТe�e���v�e��>]))=�b��U8�����E��a������&/�p��7���rJ
G�K?_S��3ܨ��+��O����ɷ�we?[J���V�ާfVk��ObX��I��hU���	�E��'p �Ә����S�k�X*0c>a�N'�\4�D�����4V�X��� ��Ɨ�ֿ��2��~��TfP���?�(�"�rz<&%t�Ulmod���sK_���ld�=���ZgP9��	�� C��F��=R��{+��U�HL���,k�"�M�b�3yqF�,�|'��O�^
�;&-UFu08��a��v�8۵� � �j Ɇ=��,]	��)�d16��'�)+��h��f��u�KS�$���ȶL2�&��H�m��:�#�w"Ht��Q5�!��P�ѿ#/�d���F%(t�}��KS�8���&`S���h}�+�]8���H��<&�2((Ȋ��0���:m�Jx�[P��*l��:o�L�O��ѭ⿐ފ�Ѹ�%�V��/��g����H��(f��y,���� ~1!V�o45�;<�(�6Б^����O�X %�;�k��n���O�vd���Oz兹⌑ �9J`��XE{�B��*���W���!8�w�G�6_���rJ��i}n��Y#�(�TE��%��t
���t��z�ҎM"_�#f"��kp���w�"�}a.�I:�s�m+<��C��lAlWϯGڲ���J�*hH��2��c@���Ww��2������R����do��q�����M�\O'�b�ֽ�#q�H_ka���^��K�ti"��|�"S�V�1���0pZθw��-�3��	�! ��������)����u���
@�l���M�qٛ(�߸Ĺ�{���*e�H��m)�︟>_[e�7��xR=�up��o�yc��O�eF����G�@��."2���`b�Ph�t��) ��o�]��Q��PI��^]���ȥ�1el���2�����ad��v��ӈ)��++�Y�h@+[�L x��[�����`j@���;�%�3����~�8t[lJjS`sbn��ff������V^FOܶ`���%��BS'���qt ���s�%2��0E�>�����%�֗�5������ͥ�MI��s�u�pV�i�a|Ab���)�
�vC�*�&��|p\Qq��Y��䧟qF�@�ľϓ��6���|Gg-a\�"��	f _�\��R�����&]���y��ѺV�crY�>�� �سvjwnѪ4(��5+�/^'�ȣsȴ�a�*g4�A�9F:}�r��a�Y���6����(��E�_��mU�ۘ��"c���y�l��v�N��|X9���3c�/�"؉A�c*8J%rsh�g���)�~74��=�
��V{�&XV[�]d�ǖ<q˰�`Q�8E7I��í�҄
�uV4ܛw
"`جs
���8y���Ft��e�y�B��I