��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�姫�gLk'y�ЎEM�AɬA<!p�o���s�+Y>:��h�p1	�A��KM�1>���;�Rɏ=���0�;�[ �p����4��<�������b �~�v80+Aa����ARV�e�E�.��곒t�"n����g���+� /PQR���i��ͳ���S���l��V�ށ���s�e�B�<LB]�/�ܢ' �_oe��P��.+�*B�,��8�����o ���M�$�g�5��R�� 3���Su$��Z��2LF��G�
�g�L��P��>Al;�o��Z�s�F��T9��
��hݱ�.窧���?�ʛꏌ�+�,�l�j�!ZQV�p¢?,������,U�H�Oki��t���7�IzP����r������x� �vaܪ�x9�7u��~�"�L���{�}d�F��Z+�7��Q �1G��< �IF���]��n��3���=r�8zeZ{�=�L��f^2m���k`����U�dU���u`��P*�������;��g���U��&�"R*i[���$�4�?�x��T/6h)3�t˶$��pY�w|Zf�~������u��6�#��E#,�-9�lX�R�q%��D���q��N�D�d�`D�y�@����Z.Z�)�(r|��6�%�Ы("D,WN�ZI��$�����BR�ۿ\!��a�[�8�
��J�]�tvU-�׋;n���ٴe�p^�ܫ�� ��Ʒߠ����@%�?3Cs��ka$��&���Sp�mN�
c�zA�I�jQ��>�HI�	����:�K���9����R~���ؠ���)��:nD�c��K/��eD��S�+�)O�Ӧ8��;¬��\vԮ�<�I��N
��	Q�
�a�vʁvN�o�Ր���N��TA�$�?���,C������ ����^^N�`R�X���P�,ݘCA�y}BW�i�t�/�59o5�kg�dƮwY������|cX8"���Dm���pϯ�N���Z��_X�Y�n�t�l����r&���� Seg��_�������s�0%� ���C�yN�K�f�ڐr�(�o^��>Z(o�q�,S�G@��<-3b�Rc��ᔼ	��I��r'Fe�c|Z)Az�	��%�؜��}-����i�Q�"4Hs잣�s��P���Z\T(C4t �]�F��i9�|��� ���$�19K���R��d:��.��'�!�h�e]��~�hT�M&OF!y��l�(����>�VX�K��MנW%�U��픿��a���IB���^���!�R>�D���RU)�,
N�N����xN�,6VC�G���Sr4)늟��HQwd���ie����#��`��d1���Q^� �5�]�,$��r������2'�4�Lh��GG �q^�E��w��R�@�'�L��U�3q����a���D �Y4�J����M���8]c��M8t�N�p�g)ob]`s6�U�t~k�N�6g2�����#(��̖����`����tZ9��-��ɋM�HdD��DRd�Q4&��+�=&C:���g�εS�g,����%�w�v�D�r�3��_����u�B<1��,Emќ��TVE۬ø� �Y�R|����T�d5N��P�%�V�'B���)q�nfws�%��y��r��([�����:�l��U"`���6	��������������<�UQ��+�u߽��3��j��h�9�M���_��Fs���ɪ���)N�L���Pїj'H�k�]��.�C,	�a+[�yް�Pb����^���|BG��e�/��Y+��_�e)����V�$�CRMUف�j���5��8���
͜�b����)�Z������&R_���� �w�����;ڂ��zʻ��9ZK������4��ޚ�?�y g��n�o�dW��#�J�͊)��6#SA�����Z�m�!���㉔W�j��K"�L,�5�!��O߾D�� ��d�$�ߙ�-���}���ي�G���o>/u&�2�(��l����,"P�v7%+�7Y��U��,|���>�r��*���9(ݭ���
_��Q���9?Q�/&v|2��`�F�������Gh��3n�ߗN�4��P'��-��<�NZ�rrr7��i�F����7!�S�^")���f"�/�F�����B>d�ҽ]�f\Im�g����I�+���"-"'�5�#.,QV��6j��@.Q��h���DJ��΂�/}4�p&�3�IC�h0};�O�A�7�:pG���mT��M!����7+��KtT04�+ԹDq��l*YF���a�(��1o=�JI�Jª��E�y������y�{����j���$���:�Mܭ~�Q�T,�l�D�N�S H��	��>�@�#R]�aEz,+�ұwL��i�M��h����>����k�r8����Z1Q�d����ܳQ��}���z'����jNHC:�W�C���ϭeX�5��31�R~5�48|n0ľ���=� �G���A�I�T���l�oU��s�Gj�N��,ZM�2l��4��3�����^��t��>y{�G��є�01S�L�=| �~�p�8�#5m�����R��LK�� Iv�tjj����w����fa��^@�$U�^�����%��d+873�l�*��>��lXr9X�j�sg���̀2k�}�O6�0-�{����;�W�I;�����3�L�ͧ4��P'2۲p< �/-�<�T.�a<v:M��o�͌�V��0�fd4?|gE"鑅�S��ӳ��9�e6j�� ��.�P��VQ��㋯��o%7�c*��7���'Jg4�DM���m=�<��W>Fu���0�T1xԩ��4uC����R�?�B���;,�]Q���ic�1�Ѻ��5�6cWl�r#N�ě���_��PH�zrC�U#�UFړ�	԰��Sz�1>��ygRAD�I�*>Ks�ZzaZƯσ�L�W�"�ߌ��/�Q�Ӌ/~������p�u榙��H��`���K�A\x�Q��&���s���꬜��K�)��u�[+K%�.ݐ��g��d������j�I���6՚��G�-p�O=D=��	����7"#���넠
Yo��ϩ+�������qC�����c�������=�b���8�i} ����U�RP�K���͠�fc!w��t$���x��"��X��r�C?��%����?I��|G���9�M�8�o��=5�ؽLRP��	SĠY\v/l�)2��c3)4�T�@�M��'�ǋӅ%K+)��%��D��e�P�,�&ӑ���K#�}��")����UP�PP��k'��
�m�o��j{�$
H�J�QF,mw�qf��^��ܭ��l�.u�uI���%i�d�RIM��e7R���[gf^�BS�l��X����ía��h���kc�a`���+P��N`�H�������L��l��\#ƃ�������_�xty�-�A	:��ݶ�x�p����������.�\���3�������s�'	�g�l,����Mw(��X2�5_��	=1o�3����IMM��4��G��]t�����Q�L����_H{� ��ߟyb�E��lL?�����#���`i	y28����Q�����.��A�O�������҈��Ϧs���ۜo�^{�qb׀������@�.To'Â���k��f8���,05�o����n���U)�t��Z���dm(�`L:�Y�K�FL�� �)N�rzE���pS��a�va�|": T�o1�RA�i�~�zN;Y�bI�$Y����9aE$�݆�7�5ҨI�ԯej�탠�˻��#�׽|ن�h�N��� ��&�HW�ަ����RU�`�j�cK�:�! 1g��b
s���|��j�n���$3c|�C㭑�?�Q��5��H��6e�� A.����ߚz8^�~��c��a��}�f��KB�q��]��yE���}+f�n#�TP&�̠۵`��D�vX��J��*-o�J��n9���]��P��ٟf��γ�xqt΢����O}�1�	V��FQ0��B=4B��w��t�m�
r&�Em�h��$<@�mVA�!2R��ǵ��J֘b�0B�1]�6Go3X9����M�H���ӆrTԕ�0۸%���~�W�GIs�ߡ8ᢉ���:����S8�����Xl�h6nf�Wh(�3/T\.m5��&Cxж�(_�-4�q�V�O�X��@r cy�K`<�yk=��tp�ݗy�