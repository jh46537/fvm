��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�T���g�?��L�X:�O����V��.U�;Q����b���`!�Hz���(�$h�65�X0!�����r�� >A���L-{9���w� ?�" �a��h߱|��Ӎ�:���|��)br����*{�SPv�+��\�Q҇��?���{e_��@�p�?�߇�)r��zM��-E�U��eT#�P�_�lh��K�	"T��b��I� ��qJ��;����N��}�Bj峇�;֓���n�{���㝃���� ����1������ǥL`s.����f��:�����[ ��M+!�Y%���@�0
-З%pZ�q/��'������d� s�k��H�V�(F�K�2&�H�RfJ�Y?d��s_ �|g���{��+.~�����{�RJ ��ޓ�*&����<s3RKk�x*�8�&�yo2�W��f@a��B��FX��O�kL)h����8�P�4C/����=���$:�T���%��^`�w�z�T9X�"P�,�,M��sB6K�B�c��������1�@-w�d���V>L�״Y'�"d���2���c��T=K�f3�� �g��\a�F�PjEN�iNYv+�t���@x�y]NI~�^<���咢����3��߮�n��Am�,�W;^F[�d�L��o_����c���iSQ-X�QA���}��d���ٔ��(��-�E���&�/>���M�*��d�t���N��؄�0\��C�.��؜���ۯ�_�2�=�'��8�T�ؒ��ar���F+��Ç5�Z�Jr�3��] �� UI��Y�xn��u�{���:KB����;UA
�'���è�68�B=����{$�ʦ�.�*|6֝35��05,e����|B�� ��}I��t��\3���\Ȱf�aMހ��TMqO�@bgL���o}~���d���JC�w��M�@q�^TO�D�X����l�M��4�S�����Czpռ��oN��1�c�^1[����;���ML�=�$B��(\	�"a�A������Fռ������ϭ��&7_��15����(z[�s�����v�Ճ�?Ǹ�OڲC�Pa��T�_�9x�.�h�Ş9w܍'/Vw�e7ȴ`���#I� ���:(X��[��=_)g�x���[��%� ������y�Y���v�I�6iGT¹��Ք����6�@-�e��0��׌�6_�=DÙ��_!^�ӫE/~��-���}�c�],��w�۴~��Z��"萸B�.H*HC�5���-�@ˬ�m�&"!䉏�	�a5��֛���n�-z�h>�tݬ��>q����~(��S��
�#f|�DƁ<����dE��{�9��ԉ��K4��-
�����KN�p�TE���n��OR4S�����tO�Lx�n��m��wM�5�+���:�/�8Z�%#ML���4�:��u~��E�j�r���/����oB���,"���|�%D�1)6Xo�h���)��<� ������I�nO�����̏2���z��Y��{\p�v\��Lig�ڏ����R@
"��` G$���,�O?1"(�	�Vj�`
�!�9/�5ki"┴�C�ب���i�0�5'j8�g�+�Zq��&�wf/}��߯��h��Zeg�\��
�� K[�\?R�t�F�{�
�=@���F�6��|�!'� 	)o]s!֩��J�,2j��;� �&���>{/��5�]幔>*F/�"Z�[hyC��A�A��n�H��ׯy�U��Cw�d!�u�j�°6`�A�rBB�!5ӞO:7��lͨ���Ӥ�����,θr&H"d�̓{�[@��bT�lnKX��3�>�O�^��}��S��!��A8�)���K��L���9:�P�y��	U��p�,(88Q�����>o��N�����na�W��jl� �&�h�2"�P�J��<��8h�/�jH��·	��������T�.x%<����J4ț��4�z!��$�z�����gX�m��W3�^2�]b�讃�=�A���t�Ur�ܐ��J��p�E	?G����!_�]^�O��-�.�#wZ�P��v�C^#I�xә 3�4��0�e�VGyw����'H0<1m_���>�(>[D���,	4�\"��EA�,E��G��EA��'��{�ZwS[>	��O�@�q�>d^��ƻ� �Է�V=Qـ�qߡl)�"�z�G{w�������1S.\Jj/O?HAյI��g�D�u�rZހ�㌡眼����h�v5n`�/�W����]����	��`�#R���DK�XL��N�?�a�*J�O�=��G52�6&1��s���.��Zz;��ږ_���Z�S�ŷ਑/���Se'�AagބJ��y,���=BI��v^=��Y�;�ր����9�G�D�<]�����6�l$P� o���r�����I��~Y(jfQ���q��{H}�4bW�'s�	 j��m.�= a\̗��ir�LcSw٫���~��z�OѭD"���!4�B�g��z��"�(J�ٹI�������>S ��2��H�i��]�3�SL[� 9~�4�������Hp��~^[���L��a�d�;a�$;��[F5�;��'����"|3Gk�H�\$ �T��mq	 N�x�����˪|j� %�Me�����*�TF��R^���+����������%į1�E��VT��Tz�kbU���^[��<�4b8�|"�:d6��+�Ǜ�=X�Ad��pd:v{�'�����б��&��b������(>��$�|oٰ&�2|P��CM�I�(��u��7����W(gty������^j�3��m��Ml=�^-��cѓy���D���α�f���C��{,�n��D~m@A�x�dx��.qS1<}R5!�@9]���o�Oe�	э��HOn`eZ�j��'�����{|��w�#������$u(����2���ȳb��]��^\6�<��Hz'0�2��?�M;�w߉9�[�12��>u�T��3I������=��s��D4���xi (m�B��2b�l���N�&��!4�-oG?Hʍb�=��9�Hrn������E���v���}ٟn�O��Z��wh�������27�y|9]I��@�H)��[IQ�gz��v�)�-���\����V9�,�7��G�"�HeGXR�CfV�K7�ɥ�)o1�ѐ΁B�"��uEGW�D�.C�MhT7v�=��G�!¡����G��u�o���P#2Mz��a�/�r�܁��e�˖�u�Y<o،����/pَ�럗����<B	}�;�1���~e�����=�� �
~���Ś�;v�G����vv  ��7�sӀ�(�^z>�lu��	�ޣ��R1��e���{c]�EcSqf�㓞H��(E���f دv�C��GV���V���A�d�q�D�^\#�MJ��b�>��7�y�>��i�ŨԂ/P�2)l$}�~���>|E��g�|ń�Nu�B��t�>C�:}Ʌ4.M��̗飦?"g׋����������2<�fB���y�����O��@A]���m
�Pf�L�Mɥ�����CRh��=F�����ӛ�\5F��A�:�\���MYb���豼ʖv~���7��M�G���Q�ߴ*�A=����y��}��.C�!JR�	:�rR�wՎ�P��1��è�ʺ''D|*�@�u�{0T���Y�gܚz�Y\6�^���8�or&ߝ�K�!������,�+������4;0L�I%�?�?��80�%
-��lv|Z/�����st��l孀$���	Zx���)�q@r�Qb�a��M��P�]kz�˕eJ��cnn�����k˭�/�{jv�G�����Q�Ļ��/�l��g���u�(4���*nL�C��A��I�+oQ㍨�fPW{T�L�Xo�OZduǆ߻2�VU�^i��V�w���t�t��������ݗ����4Knq�d.)�Jzɕ-�yVΧlR�S�eʔ
�
���}�X$�M�=��d�(-'q�0v&��*I �ƃ=a�g���6��?�HB�Ox�<��9�+?QQ꼬��ܩzݭ`}r�*L'J�Y��-?w�n[V:"�����I�v!�M<�v�D���O�E�a�'����ؙ�4��6�����O��V4�kC�)~��ƕ8;G��]�M�E�z�4��m	�0~���r��'��&��ǔ� �<Z�^��T���'":���ɷk�
�Z:���W �4i�R�c!�<�,�yPE��&#�l�|M���� ��h�4p����R��[/��DC�¢�2/��>(�莕��o��0��Z数�_���oxK�ɩws^)���V3���I�4�Kn��r���S��Q��] !p�}�P��U/;����� �nH`�'��J5��;́��8bc�	(�J��t��Z�33SIg�P�CUh�#�>� 6��l7��i��G4m�p4�2�yP�l%�*��<&%#0[�|�<���e}������?�%��;��S��js�U:�?�f��R U��SV�'_���_˚�N�Q�
4	� QJon��IU��ֆ�$B3��М��0pO,���(K>5j���ɃP|2�������]�0Pm{E6���[�lw]9 ~�r�}TA��AZ�Qq��L0�z"�V"d����$���B���8�L	�mǻ�T��"U����� b��)I��}X;Znt�Ǌ��M&#�h�����6D���%H�nN�s��T�Y%D�����l0�kgLB�{|�4��hn��5�P'�=�k�f�V"�Q�r����GS�hˋTK��O��4���)�E �_S�߰�w:ߎ��/~���{"��X�	9�>�]��LK�0�2^��z@�.u�U3B�=G%n��r��!�{��-iY�x�tq:h�&��l��Ie�؈U����,(����l�S�v� ��07��Oљe�}z��URL;W$��%-J�7�ޭ�^}sry��%-��Rx�slf�F��ײ�$�������di��&e8,.1�8�cB�z���Mc}=�p*����O>T�3:{<f�}�ٿ��eV�%�
_۲6h��'1g�A�u�M9�t��v]?��������Ț@�f`'��jڕG�)VT<A)�*H%6瑦e~������wy]��1[y�!}�X!�+�Q�]�Q"r���t���k��ht"�����G�:��XȎ7^�����a?�M��a�0&�}��TKKTQ�����Oy�M�L�	���&.Ԋ�[$X�yR��钝�V%�|� 3���:ӘT6,�A#oG�y� ����@�4�c˞\��Gy����;�`[WxC��� Bi�	6��^ӎ�]���+r4�����O%쩐����tA���0X�ų�-����B�2�߂��7�C���m_n�.��B�UqD�_����	�׌�OP�@�oCR����5H�*��ln��� �)�Yt����qPF�f�����,����������3D������>o��E��!�11]y2��MT��t��\��|�E�̊&�F]]t�k�~���i֓��Ee����K��/�@T%�Z���!����k�S��H�a3�!�0]S�Rܹ�p���|��#Pw6|3���{��.�>�`҉�K��?�.�k#�\�٠��d��|���μ�|wF�����zVH0��f����#i��ݹz�aX�^dX�xg��fe.�DA[���춐�!�!Y�=Q��{>T�<�p��t�3+�w��y�	����9��;,,�X�`�$Rѭ��ܽT���*�i��o�9�C��h8<�Xr��+�{G�cɬɅ!Y���wD]/�uKC�Rt43r;6�}8�U��jhx��B6n2e�W���O�������j3�=��o�q�;�}���D�m��z㈶T�0�a��1AAh$>kX�߼w���H������Hp=,$��@�5�O|buL��3ִ>��p�d� F�!8Ŷ�A� 0�����f1D���M8*dDF�Һ��h���~��_H;A�����iظ��3���Zt$R9ȿM�g��Ӑ�P�"�}������s�O��Ik5�u���Ox�2!�Ww%<��f:��a�x;�<%��tֲ�Kz:�_@̟;E�݆k�65>ca�n�� �V@��?_H��[թQ�w�>�J�ѭ��	�)m��kw�6�G��@Â"0��p9g��S�Ճ|ȕi�W��'t6�Q��j�e���x��_�M�B������kϝ&ۧ���I��j^䧺�E5 �u�ś�/�\�~�a^��^�ݐS1��D����A�?Q�
��0K2x�*+�q�A���h!K{_�3�[�>`��(���j�.��^���Q�%�C��S���e�+������)�aR�dm�ץ�;�fE%,o�(6={�s�)�+8�$W7��o�|� e�Y�A�K��]�����҅ ��zĬ=����k��O���`��˹1���~ �� p&����ʅ�.���� =tT�΂8uE��;j���)����J\�wO�xH���b��E8��l�`T��K�@�	2�f؏�j�IE��[
kDӇ�}`�A�s��)��{��q�6Y�9!��5��ʟ�f6��*e��D�0�B.Z̋E&���������Im�4&���b�����
�O����
̓A�NZ���C!�/�vG��;�\>z}۔ކ!^,Ox���EG�x�S-r�J/J_�w
��qw|q	'�۽2����4mZK����uT�qi�'�׭�,JG���_�����ޛ��d_U^:V*�����w��\,P�g�hZ4��-�#1!��˰���3D�` |�!� �V ��)!��E�����/L4��X���n���ۑ76���K���U�2���x��c��3�Vd0�<綇������G��%��#�I�O�ox�5��_�K�Rq�&A:�z?��O�p/>ف	���(#N������F8rB��,H��Ƿ�A�z��i���l����^ �NS��Y�lV+���,*�#ʨk�Y�����T�|{���.t*���0�1�10�84���K�Z×ɀ(G�2���u��I_�tl�]bV����ٷ,�m��R���Ia����� �:X�����4��k����]��k�����l{�	g�%.Eҹ��)����}F�p�k��m�-5�rb<� ))�o�7�|m$�w7�κx�p[t�DK,f�a��$����<�ޔ����DU�*,��(��T[H'?D�u�(Y�I�W���C5r��{	� *�mZ�7�"K�W����r���˖��Cr�)�C6���Z���~�˰��>�Ϛ�+0R%:�G9�� �h}ۙ-��G�B�����J�V
f�-����Vt���޷]�Mn�J�Z3�ˤ%Ͷ��&\���`�8�d{��v����� �{��QR;NV�..�ac�6*� ��:7R���J��(w��Z|lw�v��vAlzGn��7���R8�E+tN��>�8�?��&L[�ѱ����iW;bǓgЂ�V2�?��E�X"a�1��S�Omq8|1��[�x7���t�T�7�K�����j�A�_Qi�9�$����gw>��l&�eO6�B��]�-�\���5�������$������~8h��.R%*I�FU�*��Q��
����+�H0�h��=��P�9�X��ki�x�¡A�����e۔�;@Ɩ��e\6���B�E%Fb(w�k��'S���W;���-ɀ��[5��Pf5�ל̸�j��Xx��{x�����ȿH��m>B_o��7��)�_T�i���W1I����;'��D�*�Ӫ�鏴�5fEW%;�w�W%�4��H�n�*�CluN�C0D��z⫕�\���my��H�,��^����Q�=+����+�K!���
��i!��f���<3�&(�e�ۣ�"��+�-ͤ���1#|�Q�!˸CWV�z��d���&�Ō���䗜s�������ۨ>�>V�Ӽ���(��w9XW��p��_2�G����9�ojU�m�0±�_{7��ʗL�F��ˈ�\ĞCO�6�ja
�Q����?�,���v�C�c�9L~�̽��G�)8B6�v&���6F�yحą|��}�������"����9��O�Yit�1�{��	���-qst$	��}�Q�o+U����;�6o<.�Ѵ�>���q6h>s�O�s�P��[p�q�I1=�Ϙ�Ktf���P�[���	���])�BY�4����]�sX�_ꙂOrmm�g�R�@�X���gJn���S�^"�t��h�'�9��%�$j<q- ���g 4i��\�9t2^cV̀�/O������s��n��fP��Bҭ*&�o�ڄ�a�H���`s�є_IeK
T�xb*wY��'���T�M�ً.��lF�Q�$��*�D�G