��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>��������ّ$�*X`F~�������><06�L���\�D>�WҎ�����r�.~O�I�V�X;w�G��ts��K�5���t�7��R��пr�.r���x{��}sbeq�XG|7 ��$�ڳ&�e
�=r�$��!錋"���ۆ[�8����lr���8Yi��9���eIE�(Z�)��VJ�j��?~�	��c��R�6���/�WC*��B�����-~��R���$=��&����O6�F�~gh��\P:�w�o"Z��{��ܪ-|$�EA���ٔ:�_JFJJ��S�B	*.�a�ꇔ�@�/~�WC(���&q����?��V~��A������(}�b	ѝu�%k!gŝ>�I8�s)�u{��>kp�Syʰ+�� 2����=��D~0.i4��SJ~��U�h��ERc;��@�p&)Aǳ)��� hU�`��ߨ��a���IG�\�A�0ߝ⢹Z�E���՟�9���p㍑~G �.�v��W5ڥEg�o�e�긆_�%�4�9�)o��4j�?qx*5��x��л��&ɩ%�:�6�����w�[kl��@����9h5=u�6<ڷ�@yX�#�X�M��wN{��|
��&?�l�BK"�z�~��#k(cTf[��i5h1P"C��&T�~�J1���Y<��3��ؐ��=�cʹؕ�7��$�`�v�%���S�#�����M��oiM��;�М��O̻��c5g�1�+J���l+�zz���^�7�G�ɦ@��n0�\��! ������q���P��v߿�|��D~&&���$��I��=s���S�$����]9�^ϖ�L�[m�虩�kI%r�>E�\,�;v���� ���ߗ����kQMP|�d��[RD�-X%��Co��.�Tr�����a`����-Á�uE9f��>�i7~̂�{�?:�s�=g5����ׂ��j���1-�zW`>�����K�if�Hn�'Gv���4�>���
r#ͅ�(�����i��Z����_|���$Br.I���N﭅�NDv�q�E���' ��F��*�V��=F��Vc���̆�N}@d��!�NI��Q5'��=��mW4?^ܗHz��t�ff��ઙ9{ĕ��Ĥ���L��T��rl��?�ݛO�*ޭ5ސb��O>G�dx�HE�	��8���%�|C�_���22/s���?��p)�U���tO� +PAd���\n!�jD�/՘[����t� �V��X�]������������0=C��OXR���Y�dCh�g"���:�k����	\�����U�OZ�x�Y�c(kI�X���A��c��N�em�}lsg��6�t�I���E�J4ʴ��1��M"w{��qb�[-d����x�V4�c���9O�z���J߿��UK��IB���H�峞Ϙŧ0����	�r!B=�(���b:�)���2Ca�`���L�e��dmn�j{*�۱t�pyGa��8	
�T����5����a/�U�L�]� ��ݡ�s�U��b	����l1�@��Z���&�������i�.�$+�Pd����e^����c����(n)o���,�ԅOj4%���C���Ean ko��Tn�lbs|����Od�1=%zb�N�%������T�H�sF9
����E˞���r@����NA��<�"�Tgd+NLr�b�Պ�\<9�K%�a���S�&M��5v7x0���$� �&�$c��`W�Y1k�qU#,{�N/ ؓ"�({�%À�֤����������%19�Н�X(�@���z��WL�b_V�Oͯ����{��8؜�7Z��|�#�I�^=�o�.����7[��u"�O� +��U�F����cK�V�M�޶������5��^Ό�7�ڲ{�:I�C�]�h5��̚1y9h&
�s��EWe���3#��l�+�e��D��M$w�d�
�{�&�^�GTn0F�����NƵG���D�Z�$nO�@�F�:�K�j�Eɮ���z���qHe�������y ����u�9�/{Z��_U�`���!	U��<��u��v]�P�^�?����㉿�c�])���Cy'I=�X����[�i�ʩF���b�N�{�f���i�\�!�O<Qy�hA���Ë_ɇ��r9?W��{�Zf�� �4u,m*��aCZ���-���xdj#����&gUh�WV��hsq���2sn��W|�(��t�O����؎����f��?�[�ʈP�p{�1�8D���ۋI�`팛��M��=�?���	
S�t!�h���� ��0+ֵ3�;�2V����`WןI��ח���.��5\QK���	c$�;����s���,.<�L��q;���L̂1�9ZZ`Ӂ$�h��#N��
i� zA��6Ї�v�\���.�!��E:"LfL����*O�k�s������S��e���Qg�j�p�]Bȿ����̮�pI-��p�?CW��S�r���~��y�)h5�&/�ƫ���T�g��
��G���Ɵ/��)f�`�ڐ`eL�͔;3�Ͽ�KM�m/��_���*[(شi.�\V5=�}R�4���j*���ǖP���׹���ب�t���]K��bp�����y�P�+���%�f����iD��9D.h)Xl7��.��-9�<���t�����9������z����S�N-��6�]��4U���.0_f���U��IA���z,�?S�H�C#$!L58"����+Kl�X������G��UN�0}���:���rJ)��f�1Y�)L��	
���HMﳱ��3i� 0nXE�r�0t�b�d7�q%�nqK������&݉TV�n�m՛m�U�f��ɝ�-Y"Yݴ������d��4�.'��۷f`���<�m�˗�Ob����8)\�]�d�!z��LS�Ρ���$I
Pa��L�/��i�qmx�]��?*l㌦�-�ke�`��+��I-��s�֮�Xg����^*܃�#�h##��;MVL�6�b`�/���b3~��9W�w���Bw-���	�-k(/�1�<~����34��S��av;���Yo7Āz	�,f|$;0��vz�`�g5>�Ϙ������H�!5�>�]Rϝ��nR���S�i���������u�J,���E9P��цm�F�l��_
N�~4�������G�^<Ȳ�1�Pne�a`��"�|h~�Idxnio�$�m�է�7C��X�ӑ���"cJY�?=(3ThZUܽe(��j�G�1��}\����=1�h��>8X0?�7�!�n�3hK�T����K	)�5d �ב���/?���<�P�;����L�mdΟ���p�G�#��?#�Lh���̙\�ɟ�Դ��/�v:�X�&���Eg����s���2�\);a}s�@�A ����d��k�d��!{�����l%�0kD���C��&E����.	��(?����i���M�n5��AE�ظG��ӹW��Dw��4��ma�0O����	���� P+��T�=L5�=r��Ν�U*Шa�v|�1����
����Թr��>�$�Z�_�ܤ�%���si2�WpK�"���Kg(K�����b�~p�V3^�?��|b����؜�����o&�}��e��$G�M���q�ꨩ?U_&�D=Q�V�+�2�(o��4x1S��>I�a���	q�M5;`M��EH��gΡ�\��OJ�������W�ͦ��B���%���>��8�������Q���'�����pc�7Y�K�|Y�Frso�#�T�ݛS�t8�^��|�$4�������lu:�����=ϣ�ĺ��J��8F�xJ{�t{����m���</5�����;rY�^�j*�D��F��ɠ�<j�a�PG蜣ܡ�W��G���u |z�	�A��D,N}2������׳�����r,@�J�^	h'��u���<{��	�>!�R�����־.�m�ا������
�٨� �5>֠{�?$�+�K�N�>)�-}��|��p�����XB��'��l���l�,�U��'H���&!�ˀH2�˴l�x*�Ohz|!�랊=l���?�R�Z^Ͻ#Y�Y��q1���6.I^c�0�˷)���/UCw}�/� #5:�5-�$T���~�2^hu��Q���8����ȩ=��4�|Ix=����4�sn���LN��Ph���m~*c5��g��g[�)��������K��o���w)��T
%-~h�gc�#�<I$�2я�����GE��@O��,�I5"�F�U�����\�(^����H��Pr0*��a�@;3+B�Y�G�+��mU(���ZC�ZRW�ث6�ꛛ=��9�h����m:�	�� O�N���Μ����j��m"9&���0�d�=b�Jt��ٌE,�Q��(jv[�%�D��^��#�T#����l'���VH���ŕ���<�8��s8�@g��<�_�@�~nc����x��H7�Dpٸ`��AR�c4�7�4�$b�;o<Ê)c�9����f[�fשE'��2�a�c�<m ��N6���A�;���ob��U��������T����H���*��%��i��}�H4��S9��t����&^"�����+�u���	 >{ߵ�H	��gM�MW�E�H�'MB�Ho��o�J|�U�E��/B�8�;\:���^y��	D��&n!0Ѵ[ǲ0���ݟ*]'��)=�F��Q\�R����f03 �&���ڛ8m��;��D�v��C�ď��;�g\i%���@$A����b���^�(��CJC�w�\�U$�uj�"�����B 5�7e_pL^��~in7�w�<�[����OX��ߋ�]�F՜l4~�h��.�j~@�p������`����-����l@W��>H�2�M������f��Mqt7\v��6~�`�1k(�@b�ٰ�����P��	�T
0�t�0v����jeE��e��.���1� �&�[Xw��>R_Ӕ�<��ˠ���
��K��J��-K�3��x �x����h�0w�׸FU�"!�7d���pt/�bCo�O�����ڽR~�����_�{�p�Ks���^�\ѥ}��}�pb����ܶK��U^,�H0��� �V���Ff쭜K�����wY��",�'0އ�`5i̯�Շ�FC�6 �L�Ʊ����]i3���rqK1�%ix(���-�Fܗ�K~����mJ�ѽ�E� 7:7-D�Q�q�@Q��=�a�e��7��d䈜���rs��kw���u�Wn�#� �2t�!� bٺ� �_F��ň��"u������ �Jq�"w�I��~�5������Yn^��*~sN�.9��a�1�X��v�P��-��ڰ���<�}.�X:%��0M0��ge��>Z �#sM�����Vi��a��Vk�B�_��3Y���&���̤�����Z��>@�miD��}��(�jͲ[���Q֦��4����S����!�,m'$�n�7��M����sAуR�t�8�QE� #4 �n����H�)╁���ΨVc#)�ld�P�>����ogV���j,)���0�+��A���n$�Rf��{��S-�����پf|V��������!|}�\��SL�~�r2l�*�]�Uzq��n�{2��.첳���-#:�ݹ�Xo������Vz���*�~	K2yep�;���ā ��ï��[�!FλB�b;����1'��������yق��(9ݴ[Ĵe]ʝ�P'���69�Lj�dy�����a��X�4��X�n��$�%�L)~�VV�?��b ���þ�TZ*�;"y����$�N�O�o��.z_|(s@���`ȜE�2.JW�u��`\%��^�`���Ma�I�d��q�I?H�u�=���� ���o�i���jХ�o��|�*&޿bq�_���`l���$^�JT.�r���ա���5��	5;��]���V/m*F������*Ъ�
���P���#�@2{�e{�'���}�U��!��È��Kj~/a���j�����b���Ot��ߝe��O���� �`>	�;�O���=3-{x���$��n���YP���M����M2���r���-����j����^*U���(��l#b�>4ZOK+# �E4��=���]ǡ��d�'m��n|L�.���l�/�Z��&܏���Ͼ4%mf��b��}Y�QDĒUoD�?({�������y����;����#�������k�Nkr�_���c��˿c6�qb�7�����21�AO��yޮI�K4�?�`�?'��x,�p��)�u��O4 X�����\�Ҵ�ϣ�y%l���=��,�1VjvDZ�&4�cυ^
e	hoi�a��Rԛ��d@Y�p�MڲB�?�g[9�/���"�]�hnxz�ge���(�z��:4��X��vJi2����#�&�_~sA��~��m��b|�C��a�Fc�9k����{��8���R��M	��鬕
�/o�����4O�� ��;8�4LN��rw�+,Dp��툿��QXǓ~��~��C�>�s�_��������ݙ������e���B��d�7�3��s�5Ikp���\����/R/@_ �JV��"�5ua���u�k3_�S�37` �Ј<[��qg���'�"�ܶ��;��h�y���&�Q�pIH�
�Z���wރ�l���^�xn�U箠حQ���
4������!{��vB�5����o���KE���$�������y<y��7��;]>�f�\�y��x�&�>��@YԶ�Wc�k<���(�����S!Ӕ^;��!�}*���@�����K����P����81Q���� �y��]S��>���܀>ӃG|�������b�:W���`��+9�Ge���!��:r!���s��̥����a��������u7�݁�O�V�N�>��U/.*N/"��ڋs�?�W$�#X*ݾ����
F_���d��'�����#[�'����WAkּ]����hb�8>���QI� �u�����v�h�Ν¯ɅLDvNhO��Z��A\�z��iK�jJ׬���:i�.F�Np�h�_�:��}��!B$?=W�R�gW�0��!�����ohf6[멌G�w��ח�ٻ%x#8K@q�5�DE^{�_j���vF����C`rvH���8F!�ؐ�ǹ�o���=.���x��s�����rD�����?=�x��h�ǅ�X�#B��Ӱp?�O���f�0#���V��J��n�T���h�~��~e��Ћ��R��,~���o��t]{ߋC���X_{����t�:́Ca1�/�ਏ:7�Qj,(dl��j1b\��>�^��<�������>Y���/�����4�1��6	`q�g,q���?�b3�g�v�LlP�ߗ��~f^�Y�w����>�����dɖ+����x����I�&|T �Kӫ���z���+?=��5�o	�Z�p�g4s\y&Ȯ�󸘧j�¨ �&ܘ�:����C��뉼�2I���$#8d;�j�My^��8tTʥ��R����m�-���{ٓQ�/��WKZ�����Z�,J�|/��	���g�"ι����MYy4(ʧy�h)��`�b�$�Ea�D����!�tgΦ)Y�p�]���G�o��d�)R'^n��s&,I���`" ʣ�fk/��E+�0�l�4'�x�ݝ��gCO���E�I�5�1_1���sl.�(]Ȃ��n�g/[I]9�t�u-�BDOc�7��M�������)�T@����Դ�+�I��,�4$��C���f�x�E{�Y"��l��Y��™]�ˬ��J�4h�E�Lg+����oo/B�\_NP*��LO�bQ%�Ƅ�k�B��ʧ��ДotM�xiw�_s%�iJ݅�Bz�K�QԊ�j������D��|�;)	Z'AF5��v�z|gq @� ���Ͱ#�����O������UNl+V��đ������YPޑݷ��n���Dץj�ѓ�	/f���D�k���8��?�Ha��o�5�C!--+�m��N�]n8&5�}�%��h����?76Q4��J��l�7�t�O���V9�w���jH��K�8�@H�M/������ːuD-80��bIT�@�n� hw8YZ�@��e,�����M��\C�A��?�����22'#Ո��!Tg��_O5v;o{���I�� ��}g�*�(���ؼ�2�~Ե��Z�'MF�X{�}�UO�9��]&��c�qډ����`��ƥ_��{xm��ms�-��B������x�+kj.Y ����/�<TMN	r� �!"�9d�_%�r�(?��#��>��ǁ�pg�S�㝯!5A����<ߙ�3�[��γ�f�΁�7�∌0�Bm��˥��gİ�`q8crE���Q�t��38�����U�)�A��~BY���lF���򹈆��c�= $�S;�7�" ��-Zߠ��5�t("?<g
�ap�N�!X���K�2h�[���|^����}QrO-@���.N�?��B�X�շ�-82K��2"���G��2�F�ki�.�V?�i��ع��[%s���ʥQ�� `����`���y�ڃ���>GLEYA-�4�s�r��DP��+-_[R�'�0*<�_j�L���KT /J�~xF��|��VRp��ٹ9F"����z�|GcN�Xd��W*Y�k�S+�K}~"�t��.a��ނ_����rd3�uF\騕Zk^i%��F��8U�`+�-�T�P����O�n���u�\v��0�;2c��m���T�fYm��Y[X�rN}����CMWj��2���R�o��b%+�z�x\r���7}X�d:��deFk�Bi�V� 
`u��L�3�VS7.FN�HI�3���$�p�����џ�O��1�{~ZO��±��8yMp���g{�NK����iXÖN������$z,Q�WH�;��S�����y�G#J���Sq��_�������*����;�p�XXwJ^�G�"���ܻ4�
d�p�I�
Jf� ���6�n�M(���.H����B�b�m}���7�=U��^�Q���c�i +^]����0�.J��E���X�^��{�v��im�0{s&���h�A;4Dڙ�Zg��];�b�l�+Zl�8n�r�UO':�(�������ǐ�Jk�D���ҩx�ӊ��Ut����~;�tJ̅��d^�G��e�শ7�C�>O��3añ��.�+��%<�\�=fر�C�J�	Wl\�AI���1��hO��=��;V��@��8��c�9�u�0 ��JMu��f��I>�g���\[?����8�}�����[�7,1AR�dߚ���i�t�~p����]X�g��uKA�a��Xo�۰
�D��J�ˎo-x������#��9�O(�������U��W��Z���ӌ�ޓ��cE�B�Uh;�>­O�6	4;���E��)8�A�/��q���=Ṥ���2d��3zN&��V0#�Xƈ�=����j6����� ޔ��R�˾P|�^��x �HH�o��"]�-X�Pդ˽.k^|è��Mu�	�Av=��a�Xᩴa]-w=�x`}�k��	���ȏ���Ǐ`�~1��r�����|y��V�&m��ɏ)j#�y��$�KwOA��Lq����+��°y�1?&�b�vWq����l�g4˸h��LH�o�@�"���_r��!� ��s��]|i=��;8`3L�e�kuӎ��١�x�����|���!=�g�T���$�~�v������\��e�'�H�:K�s�HY����B��zYl�A�#1����˟7��?<��,-q\�BB�!�&�[���:��8�چ.����%�$,Cy�D
!O��ߙ��Ы1�tt�[rS�yA3pZ�̐��z�Uk��f���4�<�Q���6T�iG�����z��V���U>{���r������l�f����f%���t��1�E3�G^\l_��^u�s���&c���:c7��iY��;��L��*#�t[���������������tJC�o�P�Sp��t9�@�y���s�kϪ`��k� 6f8�
@��`�}��;5��`��`x� ��x�V�ǹrK�N����B��y3�ȴ���K�s�x
4�	Z�V��$\�˭�t�(r��_��M/d�h��e�v``�l�)��a\JH��O��dh+�<��Hb�,`Y��;��N�~�*ʺ�0�.�b .�
�(�@�M�+٢�H�4�~�?����ʄZ�	�X	X����ˉp�N5�D�ߕ��J�b诲�=��!� �UV쥑�ےD�2^N�Z����kpodk��5�`gDpA��1nkF��נ�w��'MKw��{%1f�;n�_?QD�c�$�Ǔڧ�t�JDe:����N������kcV?0��_*�̢��}�2�M7�ፄ��/�й��6������j+�K�7��`0�~�Ŀ�U��<�M������?�M]%d��!g!)�Te'�T��T[�[)����~��`��غKm��4A�x��<��1�{6�^�`���1�g�>Ow?�ީ��)w��.�Q�ݓ�5&9����S��N@'����!��"?��y�l{��A�O֙���)�旅����->�D�sw\��W���X�م-`��u;�
�c����L��D�|`�M/��6g,��5��H��`w���|x������)�I]���_��RB@�V9��do$�r��ylÕe'��/4��б�Ԡ�-�UXH_#�љ]�d�
�r�9N�{o�gt��\?�gÉ���73��Z��K|�]ː�ݰ�Z�*)?�-{��)rX}S���H��Z���(�yJ '��6-[S�P�(S��vʘe��ӌ�(o_�i

3Vj%.tB1��m�o�t¡v�tG�)6��T{W�v�6���"�D��B�g^�>��Ō�-�fh1�� �����(I���L/�綁U�o�wʜJ�i@�S�V�+P�M��
��1����#����:]���y�&a~�����|Ԅ��F܌��ñ�	��1��ag ��'#H�����ti;°M�{ǧ@^�
�S�˛���ܬ��YC�e�RP�p�s�ŬГC��a�ߠ�����L\��6����f���5iRFx�8����O�_ D΍K&�"��G�y����U���]�2��a�7j^뇙E�ےK�=�;�3|�r	�u�f(MW��@=eӛqϋ:�H?Qpb�����a��S��Q�H�1p�n�$YA�17D��G45��qj.�@�'��󿬲������Q�Tm�F��Z/Fp$����'s�?�ҷ�/�4\����5芶��-���0N�[.����P�9Ëbm=u�����T�G�:j>��B�����~���`f<p�F.���� l}�&�L}"�NV��ЏAZ?�J�S;o&>��$v�a�Ocq��[`�S�{Vt���r������Tgl�%�j,y�1��~Q/��4�ry���\���s�o�!.~�bB2f���8��ّ�T����縃1T��������n�Js�i������귐a���R��#?����˔�����b�E ��8dДmĔ2Rhqj��9#ʭII��6U��jh3����k�W6mXb�"b��7��ݜ�`9��J�&��2W��]�(���R�{�iA�g�!��Xo���F�%���EQG;*Q�7���B�G����'M��� ]���+�é�J4�i���U�h�vVƜ��y��IvO:3��	����Nq՜�L�]�e_��A�~���n��#a����wΈ$��Z�Y��W��K2H��T�n_/�ZX����BȦ�Z �z��V�7J�K�!���:򍭃6��%$���&%ޫ ���D+�NZ�������2�����8�E|�� `��.f�,*���c\��2n���I�rrn��Q،:�3Z_N���6J��˖��W:*��c����p�����q��~l��,�!#�6�6C�H�.����C�` �\ë4ṹP.,���E�O�?o��W��|�`�����2�	�[�=�p�u��&ɀ��L��:W���Z��>���B~>s��'<�^�0�*p������/*dv���A��_��E�R�&3���*P����6�SDpV�dƶ��E˺v�iCm�෻��	��M�De8�������� ��*�9ц8n
tqDG��d�w7�e�7�{q����=c2����4�껵��Cw��D�ˋ��n���^Y����jjv-q��.��:i�͘�͓'kr�ٽ���p֢�%�GCE�{�<��p��JP�z��T^Ր����%e���c�3 #�Y ���j�O*��]�g�_a�l5����wY����%����B��	���Ì>mV2�0/g�MS �,K��eY͇rdFG��|!��Ĥ3:��j�VCφ�+q�h�@�Og8�}��>/n`!����2h��s5fʐ^>Ň��A�zf�K�$�v�S0��Gm������A��{/�Y��aQ(����ɞ�jH����[xD#��C>I����Dȍ=�z�� ;�p�L���y�"�mYrQ����.���O��8Y��h�`w �#�S��(Q���L��"��\Rޏ��� ����`���Q��R}�t�T.�����h.��}0Q��������������P���tHG]~,A��x��u�T�2�D���Xm��d�w"d���Q�Js���1c�J
�&��g�0^�X7ܿ}ή�>*I��sԕ&`t���n~ {K��@���X.0�qV{��Y��Z�n7��O�b;d�Du�q#E���^�j%�k��T��г+#��J�a��q�r�ćU�z��~/�r�	����ಮ����J_����#z��v߭u�reE����E��S��-L�1��.|��Tr���IR�-^���ZiOq��pV��aHA׀bizM���N���]��~E�����pQ^���p<{XFy)V03L!O���{tҵ93؝���Qr+���6`����X=o�
�k��w�^�J�8����=�h�e-W_�Ėf�A��B�8U%_��: ��
�K�6���[���5�`�c2��Rzv���՛��@�p|YS�L��E�s*N�aYC{'n��tm�5r9��y�W��"��,�_�G@Y�Ծ��A4��H�W+nz�XeK�'"�c�����.�,x0�< �������W#/�N.��ʦ�԰�Klo8t��m��T9N���m�|�;�+_�!��^�M�c�i�D��粞t�������a#���Q�ٵ�\G�B�C�Ϭ�/i}���^: ������@�j\�V3������\�SQ��W+	�!��I�*>�Szd:��^��M�k���zd�i�oV�@�᥊&��/�*A�J�5 r�rگ2(��p�����@�>1�~�wzCc�,�r�C�#m�þ���4a�H��p}I�9A�h[!��b��S���l9#Xد�<F��u��餹��_. Wbm�w�`���'��"����u"D^ػ��a�O�(�S*)�X���lh��wPN�ی���l���*� ���(�����-@{�`�� ]�ӳ�B�*�����*a�15�Nmۇ��t9曛G�0QPy��?�PU��⊺���E�z/��T��	��2&t}b~�%T�*5����45��S����i/݆)@�!o)$=�ʼCQ�THק4%��X'0�k�-��I2q4)����+���1��j�4{'�м��H*;��^�N��)]����J�52��%��M#&>���v�靁~য়��'ePW �߱�Vx
�)_���v1�|Xj�M�dxc#P��oo�Օ
@�߶�b�R�x>jΚ���T~W#8����_3)1���M��i�W��W��7�?�����$42f���<jHEQ�4�Fk������,���r?�\�� `������2��>k*�ilV�pEԃc�3�8���P�}���^:�O֚�/YS�<�9�F� xs���2$�S=Cw��
���3���ǘ�W�<Xfǩ����?ͫ�ݕj�ָx)�gE��zMK�`
����G�!Mf=�)�Ko��/*j`���f���B����j��?�Ug�p��)�����Xm�C�˥9���طzc�"�4^1�п�ۀ(a�%���W�r��ݬמ��(�o#�/�zG�@�PD��J�b>�W�lB��J9(\�CQ��ej�(w��g�&Gz��يpJl�Ly���z�2�z��%�<��j�"�7%���f�{n3D|>G���u#F��7#��d�o{�A�,�_p���^~�g튠;
Ղ�Qj��q�V��>��g��������n}�eL��S�fK�)���p��U��}e��#?2����,������Lt�Ξ4�T�!�F�O�Q��f�PX���v���0[`ĉ\�<:�0	�91>=�êє~qu��0�(�
��1"�8W:���B�p�#���\u�^Cv�	67* �O77�'o:�h~�8�g]B��qb�p"y��@���ښ( 7�=w��3��N�dX���֪J'�v$�N��g�&�A��$���#X"���W�aM�� ���L��rݍ"�LN}\�Nf�\`@��'l���q9#O�'�/���`��TU�ʑF;{Y��Ndam�� p�r�������I��NvnRh��/$u8�hRe��y����h"�����T{J5��'p����~잲�vB���ͬ�_+��I������Y&�����A��q{��#궰a������s�]�f�S_�yk���a�)�'hG=;8�-��ǵ��rp��'��+�N� U�/��f���e�TP����[��I����!ϐ>S{����x�
�Sd�Lp�k���1�Z����)~����< �|�<#H!�"
����V�b[L�7��h�Ԭ\��~W��Fj���)���j�p%�D@W����E�����:1���:��a>�#
%�ǃ�\Žuhh�~��6E`G�سGR�#�}N�||`���%'� ����`�K|�=⧿�=E�G����'��e?=]|�� k�N��m[��	���}���T�TD��ڮ���0anA/!x� ����/,�p �'�2�blP���NK��xW�?���u��4q�����X���s]���m	_���ՍfZ]*�5�J/�jä�qw$��\��.A��c)�\Iꡥ���R^z��G��Ö;a\�t�8a����V���C�c�z��x��"t[h�C�ޱ��+����Fy��>Vj���dƔ� >@���+��w!�=���mم�h�c	�3u�<z��8���']d��"C�L�0ѤxT�#n=W$��`�a=g�����*�n�1���w�}I��C��gnv��ׯWH��"��b��p-�n��m�qo�:��㓙�`fO��̷; ����r�.�ћ��X��Cm�*��:�%5�G��������.7o��&mE\
ۡ�W�BE��m�3��umֳP�+��Ut�ιZ��e�6A#�V�]����3KZ��O]A�Z�F.��N-��_ْ�`8�����5���A��M�j�P͹PGF��}[��F	W��-�ݦ�̈́��s眹!-�)rQG�RXQ7g��D��fQ���C~R����G%ŻQ��t����	Ķ������y���F��-�iЩ!X򑘊7j��Sl��A|Ua%+�D��nF�֬���'�ޝp�禳3&�4��"�U�.�F>t�@�ry+�`I!��$}~v�!ٰw��6��1k������ih#y�'���-Ӑ�Xp������hAE�+��aS5.q- .^,�l���H�F����X^��-K��W���_Y�&@�*���YUT�I�����6��lÙo�MBx��7s����#�sO��!�i���gU����#�h�BX�4�Ǯ}
�s�(�HM�e�(";�����ݢ�!*�K�m��LQ�S����Pn��e��M�+s���t���V]�H�����ւ�%�xd��\f Ff?�<�r����X'jɹ��)dǫP���3����q�
c�Te����#�hF���L��cưb�I��Qā�}K!��h�Œw�^w�w�D�03Xm?�F=^��fs̤5�9*H�q���X���4q�\�+2`
%�o�eW���< �]c~FR�Ŷ��C�vEX���T��C�N�XPl��O�Bm�o��*^��F���2뜆4���������r��3_�8h�(�O줈r��Wm�U���A~Ǟ\��A[
:z�P��\Kz\�Լ&{��@wg=>�t5�7V��13-;3���b%x#|�\������
!}�~#���ݜ�Y[ޖ�8~��H��yV[<�
��s%�i��.����{�VK��piؿ���:�R������ٟ��ք�QG��li�,rm�CY�<5yg8��d�usv$�ҍ�r��q���N"��o�pC^��5=WG$P����w��S����_��[qL���{�J�(n��nx�z7��ry����:��7\3�����2Y�P�:sҎ�[�-��2~	�C-�ܘJ�WGQxr��o�d�nrZ
�,�'�ǵ�h�[�ߢ}|���
�9�C@�%	��3P���ҩ�;}���g!~�z����F<Yk�Y��Y7X��
,��ha��h������!C�*��Gb��-g��� :����֏ H'6g<�vXşV����N���3���2xM��@�[����}�S`K�7�W@iKC>ai��;i�귧/�Ď��*��F�nGY�癭�@Ҝ��S��-=�	&}�`G��� ��G��JA9G&�P/�1��H�Y!������N& �X�~�=��K�J��/��
J�;�hD9�J(B+��a�R}*UU}C������ 
�ծyƶ�bp�p�N:ǭ��KE��ڃڭ�1�5!�o�����)�k���qܚ�#"|�<^̸�-e��I����|��I	���2��s������-$����:�h�x˧w1�s���.�WK�a�K��=;���������z��ց����l:׀v��p+���P�0A ��w�[�|�k��7A�n9��28���%�Iu	�IR))��P�Y�傝��0qk��x�jt�wZ�,����"�ċa�Sv�v��Z
�-�$�r�f �0p_��j�CS�eĐ�3��)q�a�k!��MJ�s�T#�7jK��|g��+��6�$UL��)�27o�0��EP&���r�ɸ�s�i�B�W ����}��6�+�L���9�C��,OQ�����Px�_WῺ�#�⡚���{�\g���AK�1��O��Qr��qS���X_�Yʿ��X�,ly*�H��o �f�J�/�G<4�����A���# `J�*��6j^���͙��5o�w�鲉Ry_��~�,S]&��A��Y� ��㍬6�{�0a�y��3ӎ���8Ű�u�*��i�u�����];��pJ�v�E�U�&@�,�2�|�Sk�sE.۹n�����։['=;��G�b3�x�R��^@�n����3� ��'{����(��S
��0Yz]~�˯��}�%�\k��SVЃP�/��~e��Vq��kQ�3����mМ>��p�L�����׺��Xu��a|xI�X��$aՉ=1Z�,�ӈ��؇���v��P
�=�]�M�4�7��Kݔ'3�:�@��4Wh��.L��4K8綹��?( �w�L;7+N�a�:��z��6�R�Q�� ����(D�䇳OWofH������J�q�b�i��o`�vՑpS�;eapF)�Q��h���6�X�=׏��O��x3��ѪȻ�|%�����lٳ�G�}���Ś����c�?�[J1r�K;��>�#<w���xhG�(P^sj/#1d\ķra���q�sMk-���upLK�{�����5�wc��|��U�D��%��x���l|R�ؤ�O�4�Z7%�/m�c���ڽ�,v\�Hi�x��G�)�-�*�'�������P.�C��(p	p�λi#�ֵ�^������r�K� Q)�0
~���B�p��!a�"_�l��4�k��A*�j?�7�?�Y�J5hU�9+z�87����B✦�_���WJ�U��kl3�{]Ib�"�v�qg�FVx�L��B�^i�AKm�v˵�#��0v®�/�1�AY�"�ʅe����]m&��czoݿ
��ܯ�Z�QE*%h˹�迊"��"r���Pu���D�t�a9���b�,9��a-m���h	����aљ̏���]!��TٿKp(����(XgwZ�'G�q���)6�2���*������^��_7i�X�GS�ڰ8�S����&����R��L�8!�����V���(I��^b����*�2��0�խ��^�� 13���d��iH��l9�Ϝә:�W+�MO��skH�'�6�Op����w�� �8 ��'a��4Y�p����{����7��2˲�il~6��@����=SV.�kA��h��`�<��]�˪!�^���p����޾BA��kC&|×�����Ѩ���,P���.e��MM�Di��lʀ�W�+�3��/���1S��Weh�I��FbmKi���l����5&�!�єI�[E���b�C�����T��@�K�&^ǲ�����I���e� &�_ܒт�����1x�(Ѧ�����{:cJ�G�)����qņ���C�Pdhv�q��FؼN�
����q���y��p��^?��r_k��@ui3g��!��S�Y\��;
J��~_�x�~���(�_ۺ�w�-�W��^��Lv��!ܾ�zn���'OJ���0E��F���n�M�[�t�$�D�	�����_sjud�s4F���'p�[���A�^*�^��w��Y*1�p`@��[8�����*�<{���)��T>�D�<a?�������zҢr:v<�*r&��S�T01��	)q3�_�)Ղ�{U�x�!A�o�d!��m����/�x�z
������ �o��Yr�jXavZCfP���^��7vr�e5�;�L��h`�O�A�'�q��j���������է����	2O+%��8]w�����@"��4����r��I�/D g�	J��5��ޣ�/�>�?�����vbP;^�B�~l�C!E>L� C�%��8�R4� �ܽԺkF�j�vC���C�Ѹ^Xc���ќԩ��B�G���k#X�́ ���Xg�,y;3��ё��i���b���6��������\l*̪!���>�����$�ӥ8��4��!\���W���d;�}���b��ؒ�� ��(qY'��������\�����鉥�c��9�Oh1r���]��z8������LV(�`�R'WO����[�ʋ��=�v��������v�����$�.�)�h��A�b����SpnHgI��
������_0AL��:�!s��s�{��� 2Ѓ�[ƹgD�
��ȣO	��[��'"C$�N����p�/�¡�>�C�R��?yU��v�뭧S���R�})�j����˳o��M�@P:�*s��������$�Fv�1I4g��iyT��zD�&��5d�n�����R��Hϲ��8�$ �8[�uN'��yg ̷U�L�� �HFr�(�����^[.{���	���~/�w�.�����vI3�v�F���	���_�T��Hk��ss��A(rOI�cAH'�b�@�Ϩ��>�6Q2�"���]�w�E6����V�?B�ã+��o�EL����F��h��nWa�7e���ᾦ(a4���b=y.��;�E��݅�/X�Jڸ�U����̊f[Y�TG7���2t�k%(��t$�BEAO������tz�-4�ȓ<�^?�Y7;�2���Y�~�7��fi��Bù��v���)R��x����5!�֢ &N�K�oc�Н�o1���ϣgC|�Z�-��ӣ�i��l,Œ*7L6�� i�T.bi���*n�5�W6yj?�q��:-5Os#�ݞ���'��ͨ�XUg&�<���}�/M=>r��ќ��靋]�J��6\o�tD�
R�q;��Ϯ�2k�8�j�΢��d|�EӤ�%퉰�NZ��1vː���u�)�f�Ǥ��6��8��(�)."e
TD:�Q����>W�_��/c[g4y̿��8�-�L�@>��B�����vV�r�A_���2�Me/���3r.6cU;A#����z)Bt�z��LcF�{T�.)�,���0���=O
	�[}�e���Ǹ���n`�Ar�UU�v䡩��{�6<�B�굧�D2��W�������(d˖CN�9�����>�p�������ƨ�f�A��G�����xǍR|�Q!����֦������{+h�����u�'<.`A�P�w)��f:{b,�,w��RUy�4�ކ�J�|t��c����N�p��Qxc8���N��GQO�&���:pʶ���
1�:��18(��.&��R����7������mP�w�o��n�/QD�#�+m�1�f[:�\qJ�Zs%�N����h^/LŖ�E�x�~F�y)s�1��]�'��G���Y� J]�k3���C�@����¡c,��z����ٟ��A��nz���~�H��EF�G�]'���S�Y� nJ
�ܯMb{��頨䝳�R���Q�z�}�D6���=��9�mM�c����m��w����H�pAEqxx�G�r^�G!q���N<ewZ�"�;����ԷJ,9 a��o�w�YO��f��t���e�
���*; �����������W�-6�$�[�&��1V�R>�k'ה�`�!k���k
Ǒ5� �����m	`G�&�{�F2<:9w�Q8 #V�x���"���}$
t���-?��4鬮�3a�à�� ğ<u���Ԇ���>~���>%��^wb5K�=ې;N��?���K�>�W�F��Î�@�A���Y��c]�X<C�+�+dꮒ.�tN��nG��h��A8M�=���h�ЎD|��B�
����>�k��H�Yp���O��SOG�\�/|$ �N%��?��#�Xm>��<�dژ�����i�}�	�3���!�P�����Hx�^Z��s�	���׆tTw��T�¶�E��f�Ʒ٩�5yV�~�63!���Z a��)#�/��g�2��H�f�s��d���A�f��ChO�<�`��^�n1N?�#f|j�?��Q%�.���)�۟0�8�8d���H��+=�ߨz� ��*��~�����J��50"�B�_�s��S��8@u� n5�Cl9JUz��cςQUk��Y��+�����4W�oĜ.��aS7g� ���s�z-N����J��;�]��C&���C]�*%�GL����/D$�M�c�$�jQ&�?�I����W�e�x�Z*��%q�ba\���+zǈ��P	,��ԋ S@W���g������q!I��טp�Ӱ�B��*~����k��'�������р��c��]��"�]X_ϒF&v	�׻(�Rq��=j;�V��B��{-V�^��36&�H�5x�2�` &"ҰJ1xaǙ�b�Fr��ݲx�e�:���4�^�(��)�e.��y@gD���m��%O}�EI�'$ڶ��h��<�v(Zժe{� .u��1Oz�莶��'"����7GmC{LR�?dav�א�8^p&�_>`�T��`�i	6B�f��P:"޺lS�>�}�2E[��hpcE'j�æ�vÙ�'iB�F|��`�iP�I1_��+4�˵o�$�XGH-�tdV���菲;���ءp�ހ!���%$�h�J4�����j�x��h%5<$��� d��W��4�	�b9u�+�c|��@�wo��ou�a[)��&�kx%oυ��ugIH~^^)��q�.㤉��^�zȞ$@������Ď^2%�!uX5F��nQ���z(�$Wq�0�A�O�K8,̀d�(G��"���"�mՁb7�D�D�e��I�Ib�I[�[g��Dj�z��-�n�cH���#���5g�]��9�Yk6�P(��'㜤�YN��&Mh����g�k�X�#f�b�LC
�9�;Qb�7\Lx���` �T]��ցh4j����_e���]�����"��7��V���^�q�-d�=�fܹX��PI�i����$��
���E�Ȅݴg�J2�Ad	��vR��7P-�}��`;�m�Jm�����p:��̶H��ƈj�sA��k����:=׌����|e��W\��i�P�w��F��/��|3��˯$w ���B	nɇ�k��,~&��Y�E��'��\�6s��`��I�K$!�4́�f�ұ.s�:����ԑgF�L�N��%PO����A8��U�g�6��n���C!T$*�TM���)�����d%����ޏ+Q��CN��� ��B����Ϭ]9ұ��S��GCVۃ�r�m��K������y�x���ozb���,�4~���s��|4�G-��bO�s���Ǩ7,d�uڏ���d�s
9��@�!�����Z�޾:yG2����!l�tu�a��V �S�_���YV+jkS� �`5�rA�L�AF��IEU�.ġ�˖�O��Z+�_ˌ`��=?Ř�`��<Le@*tz_�N/Jo4�]=^s�j��0��"�.
k����J�pw����j�.?�j#1�mc����ū|�T���|�Ҷ��(�c'��_GXϚ�kïآ�&���asq<�~{^���+����V����|��s��������Z��IW����=ㅉ��4aЅ��=^��<���1|}_��2̧�~�J��������!���@�2�^8)�QaQ7��&kC/�5@�0���m����Z1!Է�$�<5۟��xE|�e;m_Sb�m'X�A}���8�Gc���1~k�ADNSlQ.=$^��>]�:v �:�=1/CS�"�us	G�����q�H���O�ۥ"�t��7j�ՕT���p��NN3����$Q&���_����G����"������ H�s˒��B$V��3L,���5oM�3W4-�w�qE�w�Q���
������y���K��׾BNLϖr�oL̾���T9�)S��2�v��,;���2^+|�Ҙ��`��~&K ��󦬸��h`�{�Aij~VQ9��d�����v8`��H��e��g$d��<�$,w5�$c���[P���SR� (�4�^���D�V�=�g����r�Loﶘ�׺PrȾY!�9��f�"n7�8�H�Hf�I�Y���M�&��ZU4'�:�]^�������"���A�ȠK��4�d�O:}\�7��[�^BNeV ��I�
q�Q����VT)�Q`�Ũ�Q����?U����Ǹi߽��t.�7,�i���˂�ڈ@إ,�}��/2j�Ɉ��2CU�JJE�X)�x���RaY�n2����!�	�h4� �SF�a/V(L�e9^�A�wH3���f6y �1�G���*GO�$�)�"���l>7=Y�-?�Ҩ��:h��ڌ�;�x杳�̣�-*gC�r��CKW�p��z�%f1n�Χ��n�5����`��'��������T�Z�u>�7�I�܅I?�C�^�Zˋ�ѯ�����Y�,ٸV$���n�;�W��Dl���"ʁ95C���y��Ǻ�����c��/��,U^]����kA"�6>����<ҍ�&G�9�R+B���w�fW�E/�ev��=�>ȁ]zxh�ґ���ݖ�ι6��cj�(�=3��.��������_�a�u���>���m^L0�n�ހt&w�p\��Rm!a7�1ֽ�ErOU�)��I�%�z\� 5B\Ȭb��i�3V�	׻�+���V�	.��G����Ťb��h_pI\�.}�
�+{	�?mM������f�L��Ȧp�������dJ�(�O���e�?�=��絸��Z�l�H�U�K��U�Z�>*�p�X�xk��p��淃� ��Y�~mw�/�Ou��*G�GP�
܆�����io3�:�1�Q�:&�\ю�&�b�k��1�
���8?�D��ǔma�S�R�I�'j�1�\о�����b	s�*	i͒U��:|��pGG$�Z=�b�J2>���y��JȬ8�0�];���(X�+����比btpo��>C��S�_�Ľ@����~	-*��p2|6I��ޤ�5���+�fζ��K/'�no��Pҍ�E����0������ݣ�Y�W1��O8��󸋰`�g� n�s�&%�~Jd����op�D~�]!�_�1���zK��:%�6q�6�J�L��L9s�F\>���S
��i��������5��ON8>5����-��umA��{�d��
Q75l(�����}��Gc�y*�N�C������tM[.ߧ��8R`<:;V��
�W�)Y�X[kG^�)֧�r�myƯ��V�$�!l��J�ksSi��K��Oli� ��'���3�0�<��Ǒt������!�n!�J}D��9���3n�c��O�}$���L�@�N�58X�[�w�yL 4\�Y|ߑY<F���M�S�e�P�v-�X��h|F1��<���-�>�yJx�u�ĳ��n�8�Jid����pɆi
�!H���ҳ�e&���_�}b�h��`3�e p��6��e�w#���Z�yԝ�c�m�(�ko���jU������puZu��r��lq��2�)�$X��|�X�mpV�-+]K ��m�>"B�槩^�&Q�Y/��@�����۞!�%�@�����r��䴵�mޥ���-Y�X��k)//���a���e�o�{[r��#����07_�� ���4hkeKߚ�(٫��I���*6;H�UPH�->�u���½gs�4��F��ƭ�
���2�$Ǉ`��K��?�n�:hǞ�r���DFd|��=�Y�F ����hB�$	��.����5f9g�tǹ����
Q>�Y �:_h�/�0�wmߖ�c	�=On��p�TRD��eN�;]��]e�$zd�����@��.��q�*s~�k^v#�6�A'$py�t|��LR���K;�?�� �/��)'_w��W�=!�i;oĝ��Ԏ�z���^��T?�`��н���\+�]�Uj����p�r���g�1^�eԓ���|��k� y�L���p�Y+ܝ��1'��.d�i�&�UΠ0��%���r�I&�3C�D�3�"�d-Z�v��pM:~�
��DQ����C��d��������(S�x��b���?|i��\�m{\L�"G�#L����q�g�&L�VZa g�i{b��A�+���{�eaM��n����A�6AR���筡��g935!O۳�S�"ލ&���{ֻ8�l���
BO�&�`���eT��A�fg=����J�}C���l�%�D*�A{)��i����&*|��/w�"�S!��ƞfS��^j���F30[�wt ����W�!%�Od�M�}��v�_O"@ %�-�-Fׁ����Ëg��mv�3+z���Py�Ff��Q��ߒ�������Rc�F̈́i�ۙ|WyY� YA(z�������<��`C4�<�6��fܜW0мQž���Z@�@���3GX-��/�?k�X %u�^�5_��X���H[�X�Z�Ȭ�6螨�0u��<��n ��j摴�̶���˯�<�Mf�l.1�g��xy����bz��_ <�
�x\	DZ��w7=4�OnV�����y��״����^"K�.窞����Z`�Z����-��l�Ѥ�aR3۟P�������|���\�D/���B+ �������N�@�o6�L=��K4$ e@awYTWa�<+���ϵEU��sE�k���_��;����ywF,�@"3�l6����fJ�j��T+�p
���w0����z4���vq��͛{��)���Uc|��'���}n����5yV%n�,�.���m @2�}�y�~مmr��ʀM^e�0�@g)	A�>(�[�t(��MD�a��o�˙h��ͤS�{osX���^q^���W�� �I�HO���#�E��ߨ}����%'K'la�Lꖬ��������1/&�xn@O�P�<�C��� Rͨ�g������	��0�(N1
F�
� n�,��@�x�k��H��Y�����B�$n4Q��]#?����[\�M�M�6C�鶾�' �Yϝ�
$��f �A�]���	l����)��h���C:���U%[d�5K�x??���Q��]���z�A�B�i�-CG)m~^[A0���+�0��]���˞����PQ}�T]�.�\�	��� ��ym<�'3�S�n��ʇd?%�r��y�<ϻ$Qbs�T֨K(�Ƿ{�� �����%:������ �$�{%�4y�[`���<�5�S�c��ɤ
u��īj���`��A��e��T���f���&�[�0��Y)�qᅡ�6�)���w��a\�=�z��Fy�ݾ�F�V'n=x� !�#���^"��wja֙��GĲ�W1�G�u��ȝ^��[��4��1�˚��m��t��ͷ���c��j
�Q�e��v5~oһ�0N1��R&��yD�A?V��N�?�@��2b���b�9Ë�}��-�k.}t�a&q%3���ͣ_}d!�㟬B�z�O8Yq�t��}��b)���>8vO��.���2�P���u�vXf�ѕ)����S�C���ǒ��t1���b�i��ϝ�Y%��{A)Y�e�t��i�����)��L0������2���h�]�����>i�PC��+�<U����*@A�g�/�ڷ���x-"MS`������:d�e;�=P"K�&n�w�{"�a�3��v��M� ~�f�]����E�\t*�,���*[Ȉe�*W�7gO������jڶ3"�C����LO8.r�LeM�7��U.���Ğk'צI
AB?��=;Ӏr��d9+_� W��R����*Lu#����`dIto�����`���U�l819�p�n)�X�l$��ah�����6��Kf��W�6���\�B\���)G2@�����8�&�dt�����B�$�����j�L�vg�Bb^�1VS���UBk�Ԣ
�޺�n%�-����~q#	y�i`��kkV�e�m	۪� c5S�OP�~���otz+�t�յ�9��)]/^�����\��q}ߞ\����~�L
=ߤ�a}S~������QkXm4A&pD���y�@(��^'����>,ӫX���,�vI)��Tv T���BL����$^3�㪇 t"�B�}�#�bB�rYv��c�/�@�6�g-����CW�"mj�)}l鄠'�4�{��߆\r���?�N�G��X �,xmX���ɾ6�qe��n�%�X�@x!���gr�@Oa�J�7�:�{|��|���=�D�|�(e��3Y᪅��p�4�r?R!��?y	�����5���\DG����ۘ�� �C�8�3.�  �Z������˛w�t&��m=]�WL:�[�5c�H"_�!���:���;��F�������Z�j4ۛs�&����%����<��3�MHU�đ%���u����*N��7?&�DE$B��Ra��-�+iwo������&�/��8u�ςqU�D��M�e��-`��؊i�h���e�Ln��j&��� ��[���_I��&K�M�9��2��ā'BGO5i	b[�o�m@�ɽN۟ﻬ`D@�3(O˥!��7����0���t��(!Ư(Ho!"�X�gX P��������Y!�T�Ќ�5�wX9�L�ؿ����{�]�� ���_.�
�� �ҧ` `.������N����MrWZ���	��*"����d�1�V���с���k�q�
���[�%�	ȶ1�O���F0f�|��KV���ٝ�C�d]P?Z"H6k�M�����r�l�����7M�u ��A��,�fO������ݣf1'"Ԍ�Y�&bZhMCm��zCB�/�������Ք��Ji�a�;�ֱ�?�z+��!��̌�M8p��G3�5�
J}���7�H],�tZ��ˁ26�#@���;:���w���ؕ�#n�Tؿ��X���C�$\�������
C��� >�Mv���a�h,�uW��N��B�1�$TTv����!��
"F\�� G�.E�az�b����Tm����}]_�A//��K�20����&:fl�]��0d~���5�R��3w1B�U��W=�4
�����;S��=ɸ����FllQ�I8`��@�mߠuûx�+w�����2��1�=bC�S�6z�gB�]Bqf����s��Z��N��[�%�#��A�$#�t����PfI�a��n?hm�G�vU�6A���y�I(F�������FM��0"�͊�krJ����D������h����l�`ֆA�t��o#�nl�O0���}2}��z9Rx_e<��/��ң}}�V���+�=��,\�-�֧�m,�i���;+e�:�V]�?S�G�/6%����R�Y�}�gV&�3B-;n�K��/ׅ��G��-')�Nu��&d�2�SEi��W��>�b�j�z�}����#;i��Γ"���9y�ۭ켚���^���4%��Ki�;}(�d/��ź�QXtJ]�h(ʒ"�$�Qٿ瓿�fu�C�F�S,����'>�],!F9]!�~E��'9�[���%���*��sq.{�@űA����(S����O>����R/8m��/��>�ДU$��6��g�D��\ ��S������KMm}������]���m�j��s����e�D�62���(--��$oC�&ʽM�B��1��4''ڊ�P�|�$�ؔT��X��hw�%�=��H��5�>nƧ���W3ȧ���/+�E8l�)��%�����϶u䕺K�򹌩����4���.j�	�_b��ֲw��� zyw��7Gp�l,��v�V��8u��#�\V,g5Rj��s���޳�8wN6r9- ���{�`D�!h�t}q�լ����8}�)6���4�W�"����Ke��0D�%�C1pz�7h�s��b �Z�.�'	%�W�� ����W��O�d�ذZ�'{K����؁yP�r�z.��������n�����{6�s�	�P%խ��H�[u.�?�!L�G��I�%c���j�e (M��� �,l-���0�,�-f�,���t��r�$	@��voNU�j���T�7�#.�1�k�j���.�"����-*T�rx)�Wh7�A�p�:�b!V�Q�֯�	���7��MJ�V-���2B��� ̗c�t�)���Ŷ4\P��r��z!k�|DO��7!��.*���@Q�o��|}z��e]�䞤6"�R�A>3]sti݂+�o�1^�� ބ$�Y'����6� ��ޓ��]������U����b2��"+��D�4#	��)��6�D��r�J6�7���kք_�(��3�� �c��t��k����Z5I���5�J/�!N��e�������.��gz�Q_��G�n�	�[����ǅ er�K1���^�r��5̫��>7���;�`��ѻ�u����/h�sW�v�a&�Bl����}�<�4�o�Z$ᶘ��ɯQ�U���E/&x��$�%q��}d�vy�Kݾ0xu5zb7.���z�>I�_�2�.��*��\xHr�ɼ`�y�C��G�|lK<!�..J�=
*G_��*Ǔ��֝)Pq�G,��S��ر��0���%�1W,Q�59���]�fq.�VNδ��:�n\0���_w����e`j�嘱O�B��ζ�m��pa9���f(��(��C����	�8��>�M�<zm�sjW��}�Η!ھ�q�a��r��������=��o�<�R�h8]L�#빅dql���O�h�=@�U�H��̘�.��
#j���Q��������
�b)_��R��瑸*`M����ԉ��|d���~����}���C���~�WS�"Ȣ�P�,��ڑDR��`�o��
�o|�A7v�l��^����uA�g�� b�Y��x/�+�A�ؔS��R��d����7�@'��4Shة�t�	^�#j�U%�ֱr�nS��+S��D������B��W��H4��H�J���lZYSyD�ȡ��+���k�������ݖ�*�-?N�7 t�q�Z��տU�<�e�g͝���%��N�ߓȤ�I@�"�����w���e��M�(����5��ѣ��U̙x����W#���(A�s��:���Jj)�/`H����P7=��/�����e�YC�	8ϊ�S�q�p�D�4����M�J������.5{vǜ��Fq�ɹ٫����Uu�Y������������z/��P�����̄��NAZ�Zh���8�G��C���<�\���?fAGx-s��3�)NI3Tl��bϑ�nI��p������h��K
ˈQ�F+�ŝW����uyj�2��d�lsb��Z��(�"�.�UoXv_���	��ӤT��w�/�;����Ll����F��pĽQ���R���T���Ӎ�g�86 J����vA����b�M?�d�`#)���ުC\�s��(���]�o0�^��2/;t;��,^��F���_.��{R�	�nޤ |�h����}��Ŝ�f����S.��,��1���k�`�/��/��>2�.�=r>�}���>,<������GGL)z�bv�L]֊���n]��4�Wk��h<Y+��7F�"{��Ć��(��PGք�wp��'@���[hQO%-��C�[����:EѺ��� ^����ht3�O{i����q�>����L2
���KNX.��ǧ� !�$ %� ݹ���Na�G:����R��m�i�"��$��s�P��i�P����#RL��&{@�y��o��Sn��!�W���TW1����
��;֞�nTߩF�e��=�ǅ�`h�K���U�m�I<��0����Zfa�n)ň�I���ʖ�z��M^�d;�g��m��=uu�v�rj���]�Q��&B5�y���\~:Q\YD C6�@�"GE��8�<[��4{6�x��M5�5�!z|�j� ��gZ�oʍ�`������
E+��V��bi[����C쨞#���)���\[$�}==5�L��hRC���Λ�ȋ��"N{q���~-Y��&[��?O���@(�M]�f�e^���. �l'ڰ�X(g|J����ȝ�g�ɏ�]q<Uxq{?�xQ���N�˩v.e�c.�?]亖K�O���)h���LB\�]�GR֬r��cPc'��!ZxV�^���Uސ�x#2�Gߍx��9�J���f��)ǃ�NC �� a~�����u�Y?�Do����Ki��s��ߚ��핵"��됺��W�>z�	����D!Ga��Q�/`�z0`�gF*-*SY@+�;��u��P~���m=�f'�]�d=3R������p	K��[��HsZ�D\�k����Q.mw�,�x��&�|��O�=<���G�i5�2���������ā���;{��GQU3�)4⪞�NV���*bhV�&�~6�.��(D��z��c��S��q������>��MpM4��/������� ���p�B���hcA��`b�יP7a#a�q��u>������ޘB����b�/�J��%��Մ�+�y��*�������@�gS^¤舱b�iX��(�94Ou�.)5=���[�
��$N8����քT����ٻQ;k=�� 3a��鸲�66G%*F��&��부��O1�ТO�^+�x�}N�B���b"�3�~���H����w9$�z�N���-�\�x�<�5X��upN1����}��;�)�iJ�,յ����!���7�,� #S����,����pW�][�춆��m�E�@�=Ma�� Ut���O�Q�z���pI:t�(�av��u�X��J��o���2ۃ<.��a�\nƭ7ƉH�</�Y��躋� ,7Z�#=��YsC�����AX��Kjي��:|(��Hi�|q�%|���G�ޜ�m�r�=��af�3?�����W��'���[ �t˂��ُ�	Jx���y�r�-z{3ro[md��Lޮ�'RU�V��8�\!����:<cvW,�����暼UW�!��DV}Q�$1 ��H��`��n�@qn�o�`�f�V���$R�x
)�S�T�R�
Ձ��;�R҂�~���#h��z����LWO����_Mɋ��D�*6��ci�i�Ee���U�@!�A�"�GY|���y}m�fB�U�����W`�*�t@��/�! �������u�$�
q����ʞ�$8�)��Z�UXl���g��SRj�g���Z��(;I��걹�vX�	�3����p���v���$ꬲ��6��C�XEJӤ&=�;��$�f��Gb����n�9�B�;�a��`�LB��bAQ˟�q-�'=����u�6)���l*fQoe�f������Br�m�UC��0��'OM��a_�Tx#��8� g.3�`o�?�l3B��DPi��Nd�?T���2wЙlF	����Md����(��uG:�AhM~��s_{�J+�NÛ��:�tnW�5z�I�}n0ъ�h�_� C�R�O3F�ix�O؟'�6�m��� "��~� �e2��86 {pY(lp�Hz�!���$���i �IQ���zr'�ǒ��n7Gov�v�9ݴ>O�s3����@w@^�b ���,���f���Ͽ���BW��`�7���</���-�P.c���mwM��Ҝ�U�5�C�����KI��7kd�`-����h�_J��6�q�b'���Ƥȱ��\��poe�w�omW�������ȉ����y�`�o�J�Y��� �����1[�)sbԦzF�%3��0���Т\��`EAvw6���>.��D��̥� �T}W_IC)�m��<|w�˳�-�&m]	�K'C�^cԛ5���J��f����b����X��IZC�S�.`9A佡L����:!�9� �@��"L���*d���\L�#6��̀�2��sSWz46�mak"�U��05�t�Ǳ��;ջR?mJ��_�Z?�_r�̞���d�^ds<���o�P3�y��|F�A��a��}5>�ߜ��d�z���W����W��gݽ%g�_�_�ղ�	F������M)��u������J=��H���b�y�&�'\߼Ysj?�������_(c�l�ո�+�:6�G�.F��=;62.qv\�7O�B�RĂ�;�QV���(������F��M�q��փ�1G|�f����)#|�����tF ��|t���M<�,�ʊ��{�׷�p�Uj����g9����F%:9ZT@Ԇq��p:���դ�$��p%�!~�M��2�2
S���\��.��#��ˡ�����_]��Q�N�����2�J\��ư`�Ӟp1�������~�C*������ۈx)����;3�#���ͱ$S���!!��	�-�2�[�*+���*�M zj�&�6f�<�4*Z�ϛ�ep�-M���������혃'y�,���0ZBW��ެ�6����H��f5���#�~����	�PI�Ԟ�4"Mx�Y�ٲ�h�8L#�iS��DK��f�|d�!����T��|�Vž��s5�Ҡ��r�ɍl�Ig.)ۂ��'۩�?n�v�%�AΠT�=x�e�a~�\W\�0lf�_�� �N\��;3�ܑ"���Bۭ7 �Y�a��$'��:���y��Ʃ�z�,R��WW�]��L7��0��ҕAč�;��G��+-Л��tӄ"=��?�$~�+�p���D����}<���A��@:&��a�A������M�a5w���c��i�/4���:���vv;h�c�����{`Q�����)�n0���Y�Z��+�0�ýJX�G�/hW� ��j-�k3�/��W���3�M�m���	��=�!�
9ʨx�kD��w��x�>C��ر����OQ�2	k�F .А��{��8+��3��#�&$pUR� �%�'����Y���l�	]�L3��#����@���[5">������Ӓ�5�����Jx`���n�¯M�X��}��a�ф�`�SL�6z�Q%$K���$�����X�?M2�\�@4?�mYMr���|�VB�..�ڤS���(RP��Y���џ_�ąo��T�M�]����v^��N�_@=Ј����v�r���}�.��#�?�O2��xDCjLEW��E�;=��r`FH4�[I78��Z�R:5P�,͜:L}h���+��MGxBNĿ8��\��~��e�m�� 
)������?g)CW꫻j](����l$�Jz^rQ�L������	��M{��Ý�ط����ö�lw��M�'U㠔VO�z2]Կ�����I��s�J�k�nu*Fo�6�,�����\A�Z��6���(T�ԭ�T�1%<��V[>���AUL���_��`D��9_��bQ� �����À�*��hI;A��7�:������.6��}���9�xΗLT��K� !pRFj���Je�����2���y�WH��$f�J����-[r��Ӝ\���^k�`BW�/]�Y���
�lv��"�J��Sȍ��^1v��<Gz�@舴 ִ�0�w��z+!6'��5�BIU.�9ފ�^ċ鹅m�V��V׭�[Ъ2�D��Q��D�_*0:��E2��_(�L��<{�;��E<�rFc�G�]p��(6�c^���l�س���c��ҙ�Ko�Q5�.��k���3E��S׮G<��M�W�}��H|�1���4Z�	Jb�����!�b�4�W�l���s��k�m+��DċK#wn��~��U�r��i�Ђ�Da�]Ͻ
!�<}�}+����nx�௭�/����ՓQ�M9�"���}N�\�1��v�Vgʒ��[�S&p�EuU��_�\DU@C�\�$�{1���3���җbr��+`����m����Q �
d%�P��Cp�R";z�~]�s�Pj>��V�j1�l�q���e$2Kg���#u�M��6ZEϗ"����ܝTzQJ�?w��b:�<���/�9���0��^��V��wG��j��d>�C�Pl���8��	�� ��.bфwB�������Kb�̇pl�.���[�/�}����r����s݋��Jf�)��e�@kCK��R���Ӏ@EՂC� o�FKb��8��#z����T�BU��_;����;�Z��hr���kGP�*Xj߉3�[�3΋[��͎g+I6�#���l[#��6}��&��$��+1�҅�$�<HQ>Cj�J��I�53} w��