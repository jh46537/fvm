��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,V����i�E�;�3}��Al(
��9��+��W�Lfc0Cp����'�}a�$D҂y���sM
�FA���V������eX`��/�n_�IP�s
�g:��-\��ܧt8gA�eUԴW����W۝�U׺�L�+D}�CM��&�NEu��,�j$d�m�Ս���k��v����L&P�^v�آ?�I�(�
'�����XD�����d�ԇF[D?zS0�L�w�ϛb�I���U��٣��� �	X<X�q�~kD����iBѸp��u�Ȋ]�������	��C�<��]��>�5zAQJc����¶�.��v=��K��R���S�x�e�q?���)r(De�L��Y
�eZ�rx��@$�=a�9[[^����ǫ�+L�W@:�P������-�W3��ei��9\�@c���E4"����ypT_LS�æ
��ۼ]m?Ĳ$��.���8}z��_&�(�o%;SMo��VG޵ͦ+R(LG_�o���v~��
�X]\�C^������]��
q5U�x�_������}�F��/����F���EXXJ�0���;ә �g��g�/Y�	ؘr: ��������Z�<`����90@�~�8c��ڀ0�hx
_IR�|��K�r1����.�ĥE��'����2V(3&�J5�&%��h���*\��6.L"/�}��`���b����� ���/e�%g}Ȁ%-"�0���k;L�1L������EѺj9�\���嗴|�S7�#I����h>�
ws6�`���$KV�c�dk�N=���-H(���ǡ4�Ml���ȐkC�b?zV�q�bg��YBW�kF:j{аd5N G�D�9���s� ؏��:�px9
j�������:�O�jc���Y�6���~s֔���`����/T	R��>�w�\�ӏČZ�&�aVV�*U}������ـQ����R������f+��ʖ~,fG��Vu��R�^��?M�.�P-�m�f��V�x���@�#Q>�q��q~�Xҕ!��[#Y��Z�[cZʟaG`�n��}W�-�k���~=�ArvJ�x�õ���CQ��$�B����&lw�5*����Rv�*�["���f�'H�A����ohî�X�j*:{\�ckﮘgGS"���*D��#�$�#mH����5�\�l��e�z�K�;	�x���t���\ ���FEp�܃��E����՞> ��Ph��2�&H����}�,�g2/�hF��[X)X��>�4=���qN����4�}��(~G�=���{�'�r ���S[�陬�{�h��[v�V>QJ�~�mt}�i�����Z:X������2Bd�6SaB��o^F�����|�\�[�ɗ#�b`�� y8�f�#q��($�*7_"^ۣ W?S&,����J]!���CK�
R��ʳ� rpEp�t-���A���%��˽�t0�f�tz�:���_��+j��9e�<;'f�6;E��E4�?�W�\�}Q�7��kM:ѽ�����x 0awd43��a���R��q�tZ&g4B�I+�?�aY��<����cp��!A���g�U&(�M�z��G(Pj���t}FXт����#q��S�x_������X�������{���@���M
��l�B��l�_�q��|J�2�"�"W9�?�u��ia����@}���"�����T��X3���`��j=����-Z��ó�?f���/�C4.���%�W]��b�'X�(��Ϥ!g��COdX*�m��(����+��ֻ�!��Ӗ�/��Μ:pb�1�E��>c��EEg�$���j��ƞn�������nS��m.K�{?�|��2";�3l@��R��9V��0Mc����dW���\�c5H�R�o1S���2�C��R8a,a3<������P������A�8?|�w�%������6�	�T�2wÿ@�S7���ՀW&�|n[�v�)�UF������xC���,�v��̒�w��E`���F|LL�J߹m:HW�?/~@P���*8�Gw%�H�(�Y��!�����h����``�ʓ�Ԃ��ό���F¯!{髂������D�s�en137��9*:Df>
Nx�`f��4�Mt������)ȿ�e�o��u B��ru��Om!�E6�Zfl���b���*u��D�ʀaf2�4��.#*�S`���)��f�*x��j�3_��lv��73[��y��
.l��t�N�4Z���r(S{�HX�B��e��x��釈�����v��h�w��@�窘iG�����EG��sj����5$
s	csd.X�T��[	`!L����PҠ��ED�f;զ�*ZOt��)�Ohl��6l�厫��a����e�頚)6�3�V��/J`�(�����5��j�������~�(��R'����)��@����綮q�{k}�WBP7���W'\<\Ac��5.\���6�ٗ{s%�	DV<�Y2l2'ծ r̰��j9oz��n��b	��@�$� [>��pԄ.�==*戋��4���q��v.e"��'+�P4�~IN�c!�J�pl5�S���������Ƀ�e�D�bU��k�`�E~2�`U�jxUT9��h@��"R��W%3�@��
s<��^>��>�(
�'>����"c>c�H8���Rb+��`���(Np*������o�Q�z	��f�!qQ)��)B�����J1�@<��w2P�D�mK�n8����[[�8e�Ɍef��>����� �E�T�V�m�S�^r�	���ז�'��:�ק�l��1�}˸Zf����^��e#��ȼ6@3.T�s�:�b�+�5��7�dUܞ�$��plf�>��adc�+���K̷&��g��7�:��Ǳ(k�<L�c����
��CϜ��-��>�u@
`��rerc�EF���*46I4��s�)Bc��|��K<���1!��@A�02�7QEx}���]+m EW�a^=J��t� �*����+3;u�� ����1G�uڗ�"�EuB��	��C�8f+�g�����Q�(-��1�~��?r�A�I5��ّ�n��C����-���p�/n��kߚ�0K���ej�Kp�sR7�X�id�a9"1Za�J�>E'JBAc��7G���;�8W10�����΂��=�ޤo�%H$���4.�p<��[���`�>k�;�����y-G ����(��ܯ��@���5t)�u�:�GLS�t~y�*��XnD���B�q#�E*E�a�Up4�7뗿 q��k.��q��"���O��Q��u�J���ܰ��NQ2�Ӆ,	/ ���Y�w��r}����W��7"Z-
�-~ӿ>@��:R��Ύ4n����,s�~1{�����w��ȟ����w��vn+7��y��u��F��s�6���j�%��7*p��y�.�I�hs�C=�F�<O���J��3dކIG�ep��1�9���\Q'�	Fj��B).}gV���,j�Q�{�j�<��Ȱ�D\5m�����O�U�zT�@��ܯ'N�)>q�yoB�Y���pG)	���KC2͉7�h9J�#��`��##�֛�T����L��{Wvz@��!���[E
5b_s?Fs��n�&��D�1���t��g���0��h��^��a�$u^m����	��&:c�]����.A�P:+��>��ǚ�Y�t��ܻ�ns�-�|�R�ҩ\7�V|�(�D��)�s��d Km{A������1��ãR��tb�u�(�D�j�Sj�K�w���uv�����o�g��O*�@1B:��oY�l��}R�8�h-�ۧ��b���Lm�����M�����YUłj_+"v:O9��E���6l����O��R�Zf�6�躁w#>d׳<ȗm����o�_�?
�c�?Y���������k��
�m����B2���d��7%�2w��i�ɇ`�Fh����f��5d�R{�[��ZB��!D�\�A�I���|�\ޯ��~=��2�W�{��7D[A!���M�~F��*���F
�U�=��o!f�Y�G��y������������U��zP��D�S:_� '�E���X1������Ҡљe��(a G=�N}��� �k]�F��������B��uRI��82Ty5bb.N���l�!�4��zL/(�;�1����3�,xը|�$����X'4|�s�j7����tx��X�3����+K�$:5F��d��G/u=�e�Дym��Q#�`�zi��-���7�SB�$�%X�̀;���A����"u���ab���%�ʷ��T��"Ek��W�t��i�Q�DL)��� NJ��B�7���k'	�\�nM߀X|��oo�m��������A����#����޺�ai�
μ��1+/���\�2hx~T}}l
��8[�'�m@-S�������j��Y
k�����-�Jt��7@��I����VCZ����6�>~���4oI:Ju�w���K���/�$�uuC�|�4�"���=��0��݁NN�|�'���x���3pApM9Æ ����o�/"�1��ۊ�"�r����ڪ� /ý4#%W�b?��]�[�9=����֒e�(�=��L-�qUـQPc�_�~����?A�c�Ɩӄ���*�R�!VQ[k�QX�\�����m�`�a��ٻ�7��EO�������Iv�=Hz�?��-���B̂ 	`@Έc�;B�����o��BXdo�,�hҚ�_�����G�3�R��Q� ���Q[��J��ZbF���ߦ������!`���2�L2G��W��_,5�����gp5�L���$�4�c{���#u	��jj�c^��C�9:b�h@xB�
�P��Ō>�=�#XX��R�P~41��;�}���^n�>%�x�]ҹO�g���Wt5%RoN���"󐅪�{�dfB;�=�CM{.�"x���O��y�@��Q�x�J^����ّ���1�Ć9Y�#Rd0��>�;��9�+n�dS����Q�{���$g���V�>�ظ��4uX��@7�+�o��(Թ]�HH�X��4�FY����H�9�;�Ֆ�;(�m�"�&����ij7�g�I�B�}�J_W+H?��BIK���U���x�ݽht���xu������T�q���ܬ���*4Bn>-�(�$��ζ