��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���;0���[��q�N/[85��1d�nޭ�!oX!�ذ��p�ޥ�4��^H��*��i�f�m����l��&�<�]\�8e�44���k�t�CЇ�+Y����^���($�?�`�\!��?>���l3�d%�	�]�_�J��^���׿G����y4����bI���Ѣ �4�L�:�,nmE��HHDJٰ��B��A/Y��́\MD{�+��<�Fb˖,�r�I �����$^�tL v�z�ڥ(������k4zV�%Vd\�l�̽��b6��C<�������2�	��ډ#�X���sYag�v	M�¥�.���9��䴘
0����m�}d������W�R�S<�V�j4I0ҙ�fd���K�]�іn��$]��z����}�7�O`��r\]1E%! ��)�)ua�(x�= :��i�(�1 �K��gl�����D���@a$�;I��XE��ܰ2G��w]ИJ�uEr��
4�ey�e��I�U1��Ӭ8��{���v~k��?v�`-�C�Z��T�+�jY����m��Q_4C���i�`��S�M:)�piz��::�����r�n�,���_���U��weD��N�Kȹ�@��=�c�e3�c�$�^�~���ļ��S��̲P+j��6�uzq)��t4U��4�����;���?����t,˕0�8�� 	��IDf� ��رq ��!�T�: !lL�'t1ʆ����)xs�	��A�j�L�!�n���t-��݅� U0ҝAqq��ۧ�Ű/���n��=��£��B�=2�&��Ed};��<�\5+=֒l�3U�*\f��8�""�M��"6�c�Α���ࢗ�d�F�	p8A��cax�ߗ2�Q�^��XȡL�+�ZN�<���E��?�p ��̴��I�E�V�_�i�q(�!������#���x�k��]Q��^�*mS�ar&��j"�W�#PA8��?{��^L�L�s �,�-˸�#�g�����U�����L���.j� ��,���	��(q�����R�O�z-9;��������LH|���#	��6�z]`�nנ7��5�f�h�y׋gg`}�T[�2���z�,��5����	EI�Yp�o@<UA��f=�!�S��Ee=��~p�XK����U�.�}64~¬���������;[82��y"=���2m٤畁<�rQi2v>�T��ˆS�Y߲�
��tv��.�p�(c�[�$�x�k�z&�b��t�]���:�e��"�ള�8�.�>��üu��kL	mr��<��Z>ay���$Ħ���uV����z��z}��_qP���<p��Ê&L�*[?�?��p��.>��B�N����s��tzN���AL{h��Q��O�Ǧ�	F��([�l�b�������Á�C�7<�p��1p#~|�:�NV��l��T�Ma�$7\M�W��ߢ���L��'��"��XO�t��Qm��'9Y�Z�iÐXy��b��	��jS��I���!�m�㛰��F��h��Y�R.�f��cţ�JF$�&@�:���\���~�;Pv����܆`��������΍�u��ILGn�h����bv�dDp̼�Af��{5�KLCp���� B15�4�po�-���B���˰M���5��s�jOy�A)d&��D�U��7��i�/�m�a�ʭ��
8�$�)"�]~�mu����F�W�(}ٳ�.���,i�~ĉ+H?��ڂ�����H���<���}jcG�v��y:�9��afcL��R�#�:Z��J"g���lP0�E�*?�#��X`�x�zUʱ�i��
��ȯ-�W�,�faq��hQ�~��Vq/I�&�&F�Ե)�e����eY�\S)�0`��m/��E|��Ws���e�Al����pԌO�e�*����$�z�z���O:�RL��+�G5�1K��[M!.�:�n��/IV��W$�;:�P__A)ؠ�QTĝ�P<�4Ȏ�u��c����N�]Y�%�>�F� �Ag=�l�3�隼���|fk��9����F1��l��#-��Q^4��D�Gdz�Պ\�b�z�Ѱ�c�㤟Q�"	ۮ�Y읱�x�VU�������ྏ��/��'�����z#kw�t>@��qqξʉ�P���")�F�{�ji�jH��d(!K���.��,*�ya�̔3��@C;�T�Ȯ���M���ֶ>2)6x�פv�g��Ͱ�14 � |��q��"ϮF�J���-�*�$9}�q�Ƈ9T����w8�=�vh%|RXp��?�|ʣ�%��^$�=l���G�ŋ��f�����c���/��`j��Z��Pq�����Ӷ� 
�NP���J��1R�5��^�4c-��t0����]�W,���.���b��ȹH[�jOy�|�G\��c�&6:E�T*�"�p�Ռ�*���c�8Zv0�v�Bf_��-l�B���Z�^C:�����|��0�7oQ/W��~G鹍1��U�{	�=�]����+�-�R�'��hȕF��[�����n�q/���י�_��5�1�s��~,����pf[T��L��N([�Yp/�a)�MpN)��!����s`��r��\D'����b�$�3�⭮�@^�Av��
1���w"E*Tr����c<��mb ��/e����m�B�x��~��ɕ�ǻ�=�W�+�$�8��̩V�X.�Pc��Pl�|VN���WE�S�;.3��A���B�V6+c�e�Fԭ���O�NU��.u�z�%W��9��}�(�*Wv�?n^�DQC���-�'5�
�5�Yd+�i�Kj�v2y��Lsl�����P��KXda`��d�orA!*g%Ψ&����ԉ�I(V����L^����-Bs��H�5�'A��6��aKV�XTY�Jj�7�����[�FMY|n�(��[Y���7@:ƞ�]W��3~�&w�tu!__�A��+�O��p�o�|�푩c�c�).E�f2�v��X�M���"8��<�~ C�Ia�>_�8�i'���[��T��f0rg����͞)���E�$�)?�.Y5����=�>����GǺ4���(��S�pid����
aQq�D��I<�%H
AR�D��4bT��A�]Nf�����;��u�sJ��]��
�M��>@yC��ᩞ'��O�=+����&�t�S��S��w��.�)��{]3�;3�Ka`s��}���@��d"�Ae�k���$>
Vޞ���9�u�����~�0�rMZ��RCr�y��c݊׿��ux�����;�q<\$���"�ت�6�_b~([ \��]� D�&
�	��U;�h�V�O��V��Յ	�sTn����a"�K�BX�u�p����X�[GD������w�;SJ����+��k�����)#h�24f4��E�j�4+�4wZ�5X���,��s ��ꏮ��:M�X`��7�i� ������錥��?���Lϼ݈-ت��{�pֈ�]cZ��>�B������Ŵ4�K�&F,ڔ�U>c�J�p ԐN��\�b�=���͒|+���=�s�/.���1�s�C;t�w&*j��^Bvt~j�6GU]> $��`�D7*�f���e��㨯>�����|��7�L1JW�u�����^�:7�s�g�#mpں����k�O2��<�Q  /�2�$�W�q��)�)������D���G�]�+�n�#��n������0�E|㜴�}e񟒧ƒyD=�(b(����b�i�����>;[��h��E���o}��G�YBp��r6�^_���_sār�:�$� kr�P���^��.@Jlk�s��C�۬{0� �JZ_��F�m6Ҹ+�}�$���ʂ=&�|>�&5g���kG�np���8�ӯ�a2��8G�E:��命f��hϽ���Q�p�a?���d�\%����=�= ���ŀ�p�t�̈́��m�Z�&�QB��d9�e�� �؅�y:�)���GNִ 7���s&��n�g���`�PTٍ��c��om�Tվ��0��M�2�GY&)���Gb��Z�1�h��}��6/�b���'&f����Ԇ��$�È|�F1�Lp���K+����*��y̧�sd���	[�2��)�:��x���D��6��u/J��mxn�
�R��7��T)��s�ϝ����)�}�����uW���Xř.��st�rATh&8O~hn��ϒ��n��}d��7���=N�Q�� G)�'�.cL�*U��W?�$L�9�>dؖ�nʽh3�0�ֶ�O�$ ��F�������0HY�oN�%6�5���Vj�K7+YŽ�g�8,�+�7`��=W�3NHs�oGj�A!5M�������MtrTQt���%_J�$�Q�5�0d��I�n��Rp	V�+�]^� L1�!����U^�h�o4Y`�2	���-����K���o��R�T�%i(W �V2�!YM8���AX<�W�QN�KǢ}�z�t?����I��3-���!6�#_�ku��`<�/������U�r���z8W��h�V����7����1җ���>t�ў�X˛�����������������!��q��Q�	�r�rLI8����sZ��ۢܬQHK�ɒ��_�vVDV(����~��ZD7U^R�^�q0_r���^Ƭ)n�)�=Bh�\���eI��il��xw����m����raLƾy���Vp�԰�:�G��E���>��CL�&�!O���ؠßg�v�O`Lpk�6g��?����i҆�"OTz�W�k	Zf�uQ�o�$;4*��м���O)/�LHP��|JIV}e�x��K e�6������p��I^!BKD1�~w��*��'��*z���sv�R��˟?j2�uq�P �L�b��gъ�uC��;Rt��M�w����)v P�Wӏ{?�
!m���< <8jm�0���A��>N��<��G�d����<��&��$U`1�Rr%wx�_7��-O,�>����"���j؋F��U�P�&�\{� !%����o>lǝ��K���yN�͋���=�п0ہ�ۇ���֍t��E���G���&��mp5r�����Q�j�vxQ��(�j�o�.]�H T	k���U�D0�Hƻ� �W�902Vh��)�Jb�p|��;wo���Z\t�'U�1��ZU��z#g��d�=������'�-Y�&�^@I�� �ė�e���k�v*�Z&!�([�8���^��Yܞa������h�����NK\���Ȱ��I���� �ΖRh���y�1�=�2��ɩ���'�k_��99����dy�秬;�Q5���k�B��@Ժz���K�*����p^-�ů@%x�A4�f]%�R�l (f���;,����QAsU�_.��~I��G�@��HM:Y0.9��3I~1M��8Bt�ru5�r�ɴ�J�=qX��H
��9���a�Ea�]r�\��ͧ�:	��6z�5�
�0�ae��J��ߒ;�b�j��E�3㇪hG�	yY��ud���s�hՑ�T{ד'�oS呶�r�(���$R��8�lY���J�8�(�l3h����+)]�a�؟�T��Q��הC8��t,]�A����q ������8��'�/�mh����T�h��a��?�=��J��
�7%�ܶ[y��� �su��j�n
��qZvrR�d}�&K�.̈h��"��V ���uY`�(�<�T͂�c��2/i�M��r�<t�3P�&%�B-k�������&z��0�,'�pWT�f?Q��N��6�}��b��|]2;%s������Z�O�h��/St
)ڒ�d�7uB��,מ �i]�&1���H-w��AAc�?��`���g��r��	�Dif{����Щ��UƉ��1�o���I*Ӧ[a�H@@1��2⯆�B��J]7���l�GgQ�<��Cc}�f��[�!��zPV�E�Q���K�^xa�����8 ��i�yKצ!4�8���8G��V���3���������d~��9�J�������x
^���T_���d�^$�E��E�R:��(*�e(��>5���붾%Ykk��c�p�������A��Qsq�rQ�ܜp5�`�k's��U�#��sh	�6@��"�l�wU�������(����/������j������#�a_�RGQ��`������Kx��X�<��Y儙|����p+�v��.��p�Ɉ��]u<]�Z�'�����F@��m9l�Q3�w��#��f/��R�)�4PR���oJ-5�|A�,�����ʼ3<��N$� �&1 >� ũ�z��Ѐ���k��M�c�C��hٓ��3�"ɻX���g�:�+az���b�D����m�\��~���Նhdfeu-�/O�h�U���X�&�P�E��ľP���_C�xq^y��O=�Z�͑أgd�?��
/����>�5�JB>�(<���S/ǀ�䔼xȃ�ګ�dt"�H��t���<��h旾�(�y��VtL��`�f�krmBF[Є�Fb�%'������2n�*�XԷ�#j��ߎ� ���.2Jg��"�k�,`W�9Ӄ[�;V64��5߰o�*�`�#��.r�2�*�}��It��Hk`^�>%�_t��`H�����t@e������y0�� jOIy�=��<��f�fjb_�7��"i��e*hVs�v��>m�g�&�u�%� -Y8�{K&X ?��a̖�8SQf��Ę�)��۩���̫ �ы�E�q㿙eEW<Z��$Ŭ�!��
�f-�	��1�4t��^W�1Ȑ.&CP��:��B�8 ������O��e!�y�>P���Rhv~���n9��<�Ҏ��%���1$BVڧ=l�x�4��L&c�ĉ܃IM�G@�CZ*�=.\W� -Z�J_�Z���t��O��"�
��۷��{D�AIl�
<���Ս�y.�	䚦-oK&n���ȅ��V��<���ȭ���6��]^��ȱ`�GB��Q/��\Z1�vL����y�����'�q�D��#��=S��R��
�m�#���۾r��b�0LE	��5�И���A�b�O���~� �AI	�Q��+p��Tʺ�w����aQ�LǬm���5DmV�����k��xe��O*W�z�=�a��XZ���*|=�^�_&b�z����C�)��ׁf���Oe.5��eGL��H���C-��x�NU�����;��= �j�̲��O��+U+;A�uc7�ES>��kt��6���?��Nb⭽7:��0�Ul��Lv#�₍ut��p�q��\��u����ǅ���-�g�q%@:��$ �H塟��x�*���h� -�3��B]���:o���[-�)A���CZ�d���i�ˈ�Gc"����k(zx�-� ��i�;�ˈt��{�D��؃m��2�CҞ���\�MM&!��H�ׇS_c����wb%����8�	��C�c��0��7wd	j����\P">�] H!rM�{ݣ�Y����f~��+@�z� Q�\�5g~��}�ꂤ)Ŀ�n��$B1-�Q;�ʆ���\Pa�+�&�(��b�~����{���L�{V��� {��k�f���Ox[�����l�A�������KݘSIL��"N�X�	����(/�GV�Bܖ{�a�T�BR��,{�����n���ʹ�Ieޑ�	U���@�9/T"Y�����X��z�\�/�@J�[�E<4Q�z-��c� a*ܵf���>U�a�����эuNo���0��K0ZP�'�Y��\>b�b�$��zC�c�0���sWA�T�����R����ǎ_I�s�iqA����ГU�%�N5���8��_�}g��id=��!U]�h���變.����`m[�L�;P���;��
 !Ȋ�H�wB"(Z6�����
4��!{3+�ɜ]l�R���Q��N���jB�[6M���_��Hf������	l��@�]`h���!D�����ul?4k�u �b��U�Jfp�ӷV��R�����R��5����/��E�<��s���V�:OD�S��@��j!�ş|�ͅ�� �׌��T)�s�O�<ДHA^%�h�o5�K�"�Z�&���o��������M�j�W��Ѩ�a�T�s�۷��4�샽��R1|v��	i�/����4��H�ߵ��!`�Gc�Y�m�ex����Tvw��
�3D��Xd��-׻���jѹ�E�����w�&�^���6�/Rg���3ڪL�J������aS;&SҦ~ R"n����ޝ~+�{6^8%���!N�ob�$s�D�f����A�ݱ(� /��שX����l�G�%v����/���#l��5#�?���/��I���Y;-Ɋ{&�G=CZ�{��2�G���]���'�r�k��%����^��۾����b=���s6�W�G��|��
��L-w�Ί�Pm0|~!���Pl���:���،�'���Q���z�b���M�ع�h%��0��9We]��#��,̤A43��<�[�x��@��'��o�$o����$C�|������35��jp�MM������1O��Xa>YNC�!�0Z��7��jEmШ��_�����L��0��`�Ύ@�f6�	�fU�t��hˎ,�8P�E2Mf�\'!����9�DE�B�����%K��L�3��<���;���nݞ�k��i��`ߵ�P����Ut7�(��렵��܃��P����`ڿ3�c�_)��:��|����ђ�ԙ&8�qX�)OuX'.�3�A���	*�w+i��c���j0��m����7O�/��G���\�^�y�I�5Vn¡T���<Z���sLR�:�.Ջ�j֡=Όzl�?�J�)��_����(�prLѣ>v�Q��s�Oe��.l:�j���yҁ@�̒��{J�G_E�� 꿝;,�p�I�a��	E��
��
&�vfq���|����m(�T�ͮ%G��`�a��N6L39��9���n�����31X���֋�~Q=�:,jf_	����<������hd��GI����Y�'z�ٟ��?^�v�)	�D���@X��w,Gi�|�b��)�V�	��j��W3���k��K-tJ���S��V�LCi���9�������B����FV�Fw���%c��o&��'1 뉤e��MSV!�T�oU�x��Q』�	�P�u���?����E~���]��o�<i4�vʞF|����~�-E-��G�̳z�X�N��I^\�U�0���H��"�|��7�l�T	���$bNJ������������"_�w��yet�/n�yIé�!�������~Wd���f��wѮ��wy|_e��5�3;���:&�h����&2�M�|��i������ju#���}IJ��W�Q���*J���:O��հ9H���2��U^Z��
�R��깮)�٪�OTǅ.���&�e�(�@�Mf������a�_�7�;�C��'�5��
gP6��H����
�M�/�L2v x�%�A���Q��	V|Q�u)�k_1���0���H�RO:��E��k"�͓�gj��d���h%����mj�gp0���@|��@�-:Y�'$� ����9��9B��B��`gцO
�u��/��ZH��瑴���L��9e��Ў��q�g3�z�
��n�EB| �\����5㡕��L��ݚ5����	ՄTK���#QJ�,�h۬���x"�7�}�<r�06.�*�9�u�?����*891��̢�+�����\#��TDsΜQ�?��}�pgI�h,_�m;|L9^��v�q��/'V�{���CJ%�e�=�:衣�A��,?\�F��nImo�V&a��-\�'B��[��@],���EDL$�E잯�0$�$|]���35�>��A��9�o#
����ޙ�9����MQIִ�ʂ�����@}�8��K�dqԖ9i��a��/����zN�uG/B��_?����G�����I�[�DZ�$�e�%`&#�6v�]�����(4e�j�0k�����n�	X���䓦7W�ߒ��������X�s��=/MڛP#����^���tș �I�h_0S�:g)� Vg3y�*�X<*��R���)��3�3Ħ'Uw	ҥd��"�x�� ]�-\~R;_��r��S�:�`s
3dR�`���_�qo�$Ӗ�L��m衒˛&nꝚ��-�}��PҶt��lsw!��0�����b�֗7��-�/��+���SOи�F�}	@���Y��|�M,�"vt�J|�h��s/+���ޗ��D2�h�T\.����D~�I�v���3���m���[�Ovj��|4]0ȋQ*'w���O:���N��t\���\�� Z�[~��$���:�O���!&�ց�&ĝ[���f�����T��_���*~���%#�Y|3���z�p������cހW<X����E��m_�}�8���/�m y�gL҇�s��dY6y�ߞ���&#q�e�I��4��7ͅ�g.K���gx:���V�O���x}��`��ȟ �X��N�kziv���Ϗ�=	���Ƈ��D�;Co ~����Q���7�7�r�U �,#�.�2 �%DX���6B>���s�h���C�"x�>���)r����Tz�c�*Q�,��F	�ib��^	Ŗ�������h���<akKj���h9*-�k^)����/~��i4��˅���=U�.���Z���
Ǎ:ww7�vY���7�Ħ�� 3����?%;,`�{�U��c��jW��2a�Y$�VO�4�5�w��Dy򐄃>��5�p.�Km�9h
@(�|��*84�S:�l	�Ʈ�Niz)^�E�����߆���vj#[������c�U �=�i�2�tKe>�� �C�Ќ���F���:D�QğȖ�z��3a��d	���A�@j�?	��:�� �S��<��[�O/.gK^�����w�]m��i����>�̍L֪���v�)x'�d� -��N���|�!���� {,\r�W��5[�`�~����tME�2+R��X���Q���1��p��2�]�G`~ƚF�uݝ�����2� W	֭�cVā���e�S�?l��T鿢b�Zk�]��qIjQ�M�@F�Z%���z��ڴ�x�ʣ�ՏT�ĕ�"�*'�O����q|��hx|��a����yW�9N��_˵���Ђ�	]����#������ ��>uM�� w'�U�^�s,&^��ɪ�-����Bx �h{H��I:�s�]{=�NH_�2o)J`�A;u�r��8�U�b~��bf%��~��u�9�a��X��YK�(�	KDlu�,"ͼ������^ڑ�2���?�J��*��yׄ/��}Ӷ��*����}4��6��Ԋ��k�U��,�,�ܙh�q��C@�"kY��ʭ۩1���!ʗ�8�|6a.�w�ݭ��u�o�~�R�Yш|���|��%�Ƹ������|wX�{*S^���1ǹ��T@�\��w�4k��zꐊ

���6`:��:�n�aF����ǁ�zMTV�At�����'�ӕ�p%_Cۖ\�V�����Q�&�u����b�*w�:���B���GQ�����5�� K\Ԓ�E⤅o�b&Zҡ�xz
62�(����I���Z8�Ol°�!�B�f�S���N���U`��0�%%لGk�\�깣�?Z��& �a7Y�}�����yk�UƩO�!X�2I���j���`���Y��/sc�n�P���`
A
̄�.�ͷ2����Z�ڠeg�s��Q�C+�9�y�k��طc��yy��g�Ew�-��E�b�ʜ$>^�Qr<�Q '\�6��;�750ݥ��Ύ�!1��%5�5��H(jM��3I��6�� ���8k���1[U�Iag=���I��ݍ�2Ԙ�y�f.�R�k��n�� ��#��%:���p�eN�o3Z�:�)����[㇗S˘�#[�|V*Fw��44�7'߳b(~=����2k8�����PG����pq�#�������8���4����=�K²%��Ij-Ek���E��"�߫E�~��S(|���c	ɛs�2�ev`�6���B����Vc}�!U�YRqؠ*������$1Kh�K��hjQ���iIk��K������+3�ԚoOƭŽN�աmׁU$�'=� �*�d�"�8��4wŧ �_����������o\,a����[$\:����7#��6Z^d��u�(���P���N���ì�Eˣ�శe+b��	<���9�������7�E�k���f�O�7�S8�_�.q�Z�k�"�RU*7��df�y���_����������2���4(k�:Ud_6��hł������'�%�>a��������:��_JVdR6�۷?��_��ߩ��ߋ���=D�f&����p ����DpД't�>�'�Q�0��xI�V�\�ư�Ԇ��}b�M��jV��'��	�Y�m���n�%�x���B�k�׌Mf
=�ha�n���1(H
*�gE�l��U���7���My�k����{x�[��/��
v�Y�c�yeD/�ߤ�F8N>:�b]]��G��`B�^��y!��1U�r,b��ԪޥGL���6V�f�$V�l�g��w��qbō,2C�c��?�X8G}�V�6���$\����'^�`�-���DY&mGH%���Ƭ1x�l?�	��)2�B�\R�ĿI�_�ٛZ�o�j-�j"�C�w*���@�z�t�5o6b�aDd75,T���~�d
^�`�JhT[͎�hs6�/jC�%��Me��L��:
� L*;�CH���SL#�efL�5,��}���jg�8aF���Æro�>���(Q|����"�6��C���w�Yl�YDc�Q��󆥏H�e.Cy���g�����S�Us����u�'��R����٢ldR��������4�/�s��]�j�]	�0?LH�,��`����CP9JK�ڰ!.�(��f���l��)����}���+ <Nŋ!����
,Z��X�~��_qD	�gl���0���؄�{T��K^߫��\���&�r_�=�T-��^|(�d-/M�a5����ͷ�{�F�ɯ\���&H|V2��� �4"�����b1�`��ʝw�\tVI43�d����b�5g�T�k�=\�8���ݨ�18�r�����ȑ��Zfc�H`�j�H�&��nvC��ʠ)�zu6>�ݱr�d�LJ�T���,��B;�9�������5e�}V��֍���9��h����T�ʴ?��!�k-� 6����FJc����>g�K�����A"�T��J�9:U	�s �c&�P-[���&���+秊R�)a<��H 8�v�Ƙ��Fˎϟ_zx���j=�T����o���B��rf1S�3E������o�a��^���;pp�u~��;����)$�Hu@���h{�B�k���D�q�BK̫�gV��iŁ����rA\ʖ�h��9��s9s����pE�F��j��^�\�iť�@�t�œ����c�н�K��_go1��1 y]Ϩ��Pl,��i�pJ/���r���Rۨ�+�:�Z�Hc$����n�nF�5߂��~ѭH���x�R���H9k�i�-y7��ÊM�{k���c��lO����$M\�]��h�������ХTb���"{�m�F�eO2ýE�jEJFN����c��aXMe�cv;�ͮ�
6���?�?#x�HnU>���W���o�l���hq�T`���������o���)+b �9�Eą���Y&���fÞ�Ѽ�w4���ȩ��"�~������1K�D�-�y��A;\TkwV���{9r)��M:5q�p�b5C�y����=���\S���g���_,��-#��,4��j���	r@�� ��C��R%�r0�Kw���е�p{ Vvq�b�Q��#4	n��P^���`&�S�|�^��K_1����i��%���Vy%��u��k�����iK�Q� ��`�o����h��1��٤��?������D�bd�����	Hó��tZ�#��ވ�z|l3'��%��M�$V��O���vs-��)��)�6�p$�*b���b^ �'qpו��+p5�uw�!�&�{� ��QF�`{?�ț���$+�=APk��6O<�Z\x}�9�\�k�x�c��}��O�e׊����ݘ�0�Z��#����{���Y���@j����H� �-��2(����>v~j8��`����3�E�d1s����7:�P��h�۠s
�' ��r���q����y�5h'�=h��Rr�_6��%ȡ��@_��+�:��ţ�yC��V��l�Y&��ؾ܌�V�e�9��;���V_�*�_mŅ�6Rj��7��D���E�7�x3/��D�>a�e��Vl�B#��p���~WL�"�Ǣ��c���Zu�#�� �{rP�@V[�Ck�v�x����ƿn�a�"E� �y>�ݯ4�3#?�Zq.[�(l
�S�p��.v�qDw��O�z�¬�N��&U�H�}� �glJ�eT2w����-p�)όB�݃�� �90���/K��KYPr���e��8Q?E��*���J<�p�\sO��M7�|y���5�1m���aUb���߭:)�y���*MV8��-�y�bu�Sd<I3m7E���e�h3�.&�vj�(�>�,{���T�����D��#��4��;>�N�3X+�4��s���@܎9���ؔ\pM�n����di
�հZ�Q�t�l'@��)d����>$�S&0�Q-X�&Y �,#>�h�,/ؼI	�a�wOR_m��`��L��bl@�j>7oEtK 3Tʬ��Y�#�<ފ{�����cxf�/����j���'d�T�I�}v<�6�VI 2`�:4�3��o���r�&x�#�����fw�Vq���?-4��\�J���0��a�;M�U�l0OYz"p��/����Џ��#���:��|Ҫ����Lz�J&Q�K���Yh
0lgu�Ȟ��i�t�0�� �L��㻭����K�5�Y(E�|eG�QY��*u>ʕpE[D� ��,�b�	l1g>�a�π������erNj���}�&��প�:Q?��r8X�w���i�Ю>nMXʽ	���v47��_����� ��x�UÒ�FUL�S|�B�$E�����n����&�^UM�|m�I�3�o���'���"�/i��m�%7rx���yw�����P+�Q���	n���=�ȝ
Ć�T�\	3]Ѓ�p�� �f��]]�U.�~
�u4�#@ſo�~����BQ���h_������8hz9�>Źk�81���bG���s����~n��U\�h�q������O�x��q�1���am���x�Ď��H�rqܦ�C�mT��m�8�.3�b>M?�J d��0)�1j"��H����G�x����G�ȸ�(N�Jy�g�M.��O}���%r���L�d����M#ז�Y�*�g�I�pv�U�{tD+ ���A+N|�Z��B�J����e��p���+ӗ��	5l4ޤI�6��e�u�5
,̻��]c�!>��D$�a�ة*������О�ɯk��\���fZ���?��K�$� ��|�{�9�
��-��:��	@Q��g�`��dԈ��}��?���8\�ay7��g�q���!�D���9��vk�	�]���O��j�*`�L�� nv3_�����h�Ӽy����/Q2�ڿ�a����T�lk�ݲ���$(� ��Ƈq�[���Ty5��_��?uVw.�/2��ŇN�b( ������#/u��e���;�H�pK�}HCtB�z�Ǳ:��|����W��^��,w���@�e�U��W�'u7r��(��s:�8�u@��_?0�������?bR�(�U�uP�]��(��u���K4;o��t���7�e�X&��~m�y���[Z1D g��'+xMp�\[�TG���!.��׽wZ�-x���(�X�n�*N�w�T�7R--(��ўΖj4ٻ)�Vd:Q����=ҍ0�<���ױ������;�i"Nܨ�i�=|t��w�0�cd�a�D&sT�S�>x&& �5%c�S�[�@n!��1|��߫�t{(20�:MG��H�PH2�|�-6s��os�
���0�?�:R/��.n 7��O&�І�I�\�{]��s�>�]0r8��q�^;�Mr��Nh$�fS���=޿��q�1q�N9]f�^3#���c��)T�b�q�v$8��9M��W�F���6� ��Ϛ�mÊ.u/��!9������ԭD����k�5h�f�6]tz�Q��{�CGi5�(�j����]������L��~��Ȫ�pvh��r����ӵ;�t����,�mj�4�Ɛ7�	�)��P�����_^G�gr)��.goe�uqS��'�H'�(�����G���"��L�H�!�t�ԏ��܋'M���+�%�Հ[J�j�Q*o�21�wp{*d�E���6h�N�#w��Z.C�u#ޙ���X��g�����y�g>��Fӈ�`�H��F��`D1���Lw���]�؆B�Ci���J-��:���r
F���W>���,<V�������/Ko�ݏuFťkiq��T;4'o�o�V.$�'A��	M	�ۯ�^![�Gg�L`.�[^������������B���Q���[d�AL�?=*G�?��'I�f�&�|O�!�$�U�!���E�GaQ�bU�r�P���F9"-vŅQ�1�4���>'��i�� �ڐ�f�9qf��ǅd'��l���I 6���Z����¶���UM�b�t�&S��Kn����Vy�J�R>�S#�w:VJX����S�~!clW'�5䇾#c�C��cݻd�-X��h�k��&�$�T�����	'-A�ժsޡ�Xb��F��=b��a>M�#���I�{ٮ��o���5Q� �g��ؓ�S��2�4]�b<f�,�w�!�A0�*d��Z��)w����]^<о��f��n
c����_k(�'�)ޮ�81�88yR�81�׃���:��C�8-a�mB��l��	�8�1��yp��'z�pJ��s[6 ����9"[*���7�v�B���ю?�]�bi}�x%�zP���B�8.�߯B�] j�dg��$(r�3EU_���4���ټf������$7�x��0������}���Dc��U�����`U��O��dԧaRBU^1c��L�Qdzw����¡~;qۭ�}��6`󞷟�:X�w`�]�h
3�H�3�]�&�,K����MF������o6��Dbۃ�ms
�*�KFO&'[��R��R60��%�����Q|�B�P�q��8I�p�;��ˤhY͵�t�Et���}0R����ɟ�LA#'3fgB 4��ݯu�{�v�9)\�W�s9@�G���5��{V>�2��^9����������^?x��E�"o�&8��U����;��d��/������𠋌Z�O�b7b��ׂ��W�^�ȿ�=��`�"5" ��^�:V�KFDIk�p������2������Y6����0�T`i���Mw3) �P�~,OB�hS?����-�Aǅ_~���KJ����Ō��IT��;/�*H��A����M#�W�&$4���^
f�{H#�
k=f:��K��|�����>(���+��A���ZΖ����MÀ��;�0�N��Q�_�FWh�X�H�_191t�/QSMU�cI�h4&��LN�@���J��4 Zs��?�?D�A}�}�=��T^aX��hA��E٭j�$�/�N��xK��'�J��4O���g�f��P��I�ϒ
�]�O�͘�n�x��V��K}>�G���+x�3��ے���K���i~,��I�va�Ek	��Yr
����uv�_�+Dibr�.J�m$��)Rx��$� �& O��U�'�8d��� )���AKŅx)��s\���D�rH��q�����irɳ���BWM�,��teӪ���hyq�;�vdX��� j�+�+]��WHS�U���	��4�hM*!�}�{����d3_
Ό[�r��v�'~1^�e]޴�j �25�)�J�`�/�-h��7a��}�'�xB���b)P��r8E�hC���US̓�y��V(�:!��_R"�2����rq�G��z���1�ZR�
���ٗ��w�z�a�~Cz���\���WI��j����4Q;�LT2@�}(��yi&�gխu�Ox!{�ͭAC$�;iғX�Bo$7m�\�����T�X)�^�j��t_��������e&5rŦ��������iމ2�)e(=��J��?/+�з��Dvn�6��Z군�3�+��p3����R���LO`b����L )� m)'�$����x�ǡ���W���َKk�М�0�_<G��!�Ҙ������N����-�LX��;��}�wE,�n�q6��g��
��������mX�HcHWK���K.��X���*B�������:��a�Ѫ�Dۉ5��FFv b�B'�B��竤��L>Zz������g2~Y���	����Amkib*P�:��AHH�ߥJ���:��o�^�-9R��p�i�=ʈm�S��P����:�`���n,4N�Ȣ9�,%�M�wJ�� 4��o�n������p+D�实�. ��5Q�?6߾(E>�tx�.$�#"H�­ܙ:���&1���x_m ݪ:O���r��ПR�nSI�p��Jmإ�1�J���^w?��_p�=���ra�l��e�G�}	 �1WK��LO�Ëa����)ƞ
��(�/��J݋,1S���S有E*E��+���!�;=/�l�qѱt]�1����' d�����s�q��m2�w����Z1�e�a���(���$���a�)��0�Z�Hp�T@bo1���a��6�B�ת��#.7�����G5DZ�Ht!Ӹ�A��<{n��>�y����g��$I�W{&<C 5�I{��Փ�sI߃�s��T��!8������
{h���?s/}��]ZHG\J��9��_q��W�J�,��Y-�{�ԫ��'�"Q�+|eo"���*>m�'j{�?M���������:�����u�CX��������ǘc�C�%�/l��\hOy��^�srڮy��K���į1fǺ�ld�����#3�R6k$��RYs�a��Ȋ�`wG�WQ�XA^~��@���^�3rϾYcm�,��%#-���ѽE��V,1�s��џ���P5�	P���o�P\�uK%@R�F��'mU�B���U��IA0���p/���j/�0x���	�2Lg�=Ө�^��Xd�=�z���"��ƙ��0�-��"�S��%?r[.]���g�����i�Y	v���� =�v���˂�R�GK1��[���Ɇ���0]�R@'!L+ɛ�}�c�r���[2s���kX�0 �-�B�MwS�n@hgT�N������(�̅Ϧ��d��;Qz�M�U��
��Z�gw�E����%2�}�����,Lݑk�h>g-���/Fv^����P�>nU�@`40b������.WibV U\n.������̊�,lB����悘��%���TC�w�
̔�N�X���^*��5g0lP�j���;`ö=�������za{�3����A��^NK�.����j���'�3X�<���⡧�>2`&Pcao���i�V��@�M
O�]�ƌg�!�c\��P��c��8��#�1anK~�qns�z�u����t�kma�N8�k������az��R�O�G�����ߕ]-!�J���^�ס�p.���@�B�;F��2P�~�@nv��m�(���ڡ7�r��5]��H�����т�q"֖��W�jP�������~s�u�8MxK)��j*���.�~(�:�HL2��n��J(��E�:ITy�y�"��cl��0�D�ػ����E\��%��W(�����t<���ܬJ���c�Z�G�20���:��$*�b�0�"q����h)���}:Rg����[� ��?��#�~C�/�@��KV�9�*o��1+[��9w�e�%�Æ�t�>,'��14�#��O�����N�!������Vʰ+0�M����hKe�w �߆,���<7xʠ�*��y���;���r�p�ܠ�"����PE���^�rrP��ҏ��f	�$o5�S!�/�w����0;��˵�s�>������C��@�e���)2����&>���6���׫߳C�	�3Nh��s�����^��&��=�|vj6����߀ÝձK�|�2Ew�#a <-c;�1ޜrڅ �������}���6@��p��+xۉ��C�����~�� �Pݐ���)��Vv���q���V�d޻i��!4���13��@�!+�MT�UOک͓�T"�y�
���t^SL���A�M�`���3p�Ht6�0#�I�M�?$���i	�
�:�4���ֻm�1^=��/��˽�Jd1�Ӟ5P�4��U��#2{��(E�.�$�m����pHp��l��r�앨1����o�OP*@w�X�Zv��7	it�3��w��q�6O1x�[�|������myQ���O��#�:�?i5=���Q1��d�?��.g[(&�2�^%�\e&VO6
`3��=ΉW����,����e�N��F�p^_U!6�D���"Al�t�{��(�`F)O��չ*�8h&���dʐ�Ap{N�O~v��ܓ�������!�XI��
�-�ӫ��%��M�e�>�,u[k)���Ș�l��6P+�}Z�_�����HLy{��?W�{]��yy����9���:m��qȜ��������T��PU��L�{6��xM���:p F=��5(1r'h8OΝ+�� m�<��K��@�N���� U��m�ϪN��p�mh�a*�/��`g���ݟ�C��p�����S�� ϾB��4H�L���5^��3(�%E��߻���2±�K�tnۑ���^��|�����\�TӰ��iڷdi>�l�P8���l�Ԑ�����u���/���s'�Xd�Ɨ�n�ߔ��cX��NƠa�� $��*��D�� �-M�Qu,Ё�3�^D�ӊ���hy���[˹�23EK����)�����Z��~�gED��t�vY����^3���85Z�,���b�j*>� sTo���<'8�N�W��-j_A�Ut���}T��~W�2�IX��]�ߚ̉���Pɤ����F��aY�|*�&+)��>2��~�{D\��/���Az0��s�+|���Ӵ��� !'�QfU?�C��!�.m����͕�;�K'M�u�[d3��j���I�hс]s���a�� ��G{�Q�{�W����e�ECgE�8E��-O��/�7�3��DI�����S�"/Enٲh�[�Zؽ�B7�<�?o���т)�� :Z��tՠ.Fpykf��W����N�'53��<5�XM�ڟ��]�����d����+�w���u���̋�O��Q2$�򔰰( ��_��G��+Y��������~4@l���Hf�L	o�*σ�� "	5S�]����镤t�f���o��cl�]��vw	�x�F�!���w������N��<!�u���&T&��1�B��G~4�#�u���c�J0"������Ɣ(���|=���_?�4C���C!7�ɲ�$O9��>�rK����"F�L ���	��웶fo->���+6�~�[-v��f�V2�,�����<U�@�jӟ����C��.�����X򌸫I$���[P'IuH�B=�����'�OA(y�@T�1���23U�����؆���߱�2��7X�_s��HY�i��g��	�/݃��j�tЌ-b��_��5V�"*he���~%Ao ���<z�qŷ��Y�z�C��#�����S~ �ԍ�r͞4�JbXP�o��Z��>�A��R���u�� ��%qВ�os���$�(��ӇM���P`[q��Mϥ*T$�R`���W?�*U�T>�^�jvQk���O���eB�f��+�����ؤf�ϑ�}w�y��]�x��/�=(m��ԟ�{��#ӣ֪�o�n>	8E�4ܻIo��2o�������Wm�rθ��Д��~:�-!�	ŘM4�OnPn�ͽ�������2  ��Kgt0�K3d�j�U��(�X��#��,]i{G)���K9g�����_��#ŧ�D�tG g��!UJݐS�"��}.I���;�F�"����E�Gb��|��Gދ`�]@F8�'qF��!E���?׵{�r`���9�<$9�+����xg3�m(�t���E9˧�v�{����$��pݢ����x��RM΃.�g�+�u�66�%�s����a��!Ϝ����1�ʗ���aS��"�/u�Ly�`�2�������o!�Y��Q7���t���)j,�89�T�B���P��M4v�Oxe��^��s���6�5�q�h=���9zS�40)�`�����A��$�j�-8�~㯪���E�2?���B���K��xi�W~2��	c�#j���Q�e/G;35c�l>�W��LG�!3�fi��|ip�}�"Ŀ����"�+�a��I=�fe��r!����z�C2?�-e4�b��.�
6�ؚ����3nPlj��74�i�6�]��r!Q�U;�mv�Z�n�Ë��~�A],1E*6��EVu�A���1����~L3�h�9ٔN�]����㳩=��"����G^��,/7�'��	�TsW&�y���L��!��c�`|���V$I�X�C�P.�B���U�ؓ:
Zܽ�Լ�v���#�(0���&0֭��m�/�n�<}��DWB&�s��s]�q�$]�x�z}3�\G\�֝�o�<ob�e�k�n���!�����7��SL�n���[% 	�gw4�#0{Fc���l���I�����sM���eW�3޴�a�4]H
�/�5���?��EGp��B�Va���P�<�,-������9�v���VΪCq�kS�t�ʐ�1���ׇ���UN؀3z�Q���h��������f;>���R;0�EB.F���}�d����Γat��x{�HC�z �4�'&���%�4��)�c�F;c�h�k���DG@@ٷ��g�1k��<2��ڛ
���4N�z݋#���~z��@HXA�Q�=d{��[�r{�EP�m �P��RS���\�����XʹGX�ά�m������$��~�Q�O�����ؘ�� �:��M8�2�? �}B�}[�l
^C�
�
*B?����-�'(?S�Zc��������Y������q��ҘH8�>���hW�7�����w㙐s��6��tT���T