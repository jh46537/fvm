// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:33 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CGRWVjbRN2Fp8FYGc5A9DWb2ur+ffmXKck6VbQnQWvXYjYiddCzy8Lmm0p3PI2WY
1gEiq+I9FXy+cfGG6uPV32eA3iXDPEgN+y6JjPhaXNp3AEQdP4k+j+db0U9hEjJt
T2kYQe7BwqTHQ6dMRjVUZioXMkAAW7V90QSZ/H77Dqw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2864)
1U23r+wnzbRgLmmQ2R8AjdsIiPfuLMXmUhTSumZNiDZ7nW4dBs8cRTJk8PTAMB3i
xK80szJCJByzScLq0j8c4jvCVn84AxIgHWq7FnwLxPkND1pY2acCuAnpswL8cLRC
osFph/i5qKsyUT0kshYopw7FtxlrwnIYYKRqkWjNrCd4KJtn+xMUOfqcFyZWm9M0
RhJkvSTdDkQrmRLCL6g+G5vxgJJL7a4DlnmGwawf4QA/CJoODGho/0QrmXyoKQQk
m/Mo7O+6G9s/cSbFQYIemsshj28tDJ8xItVDzBbPD8aC3l2PjQwZwJoj3CUtRr2M
eWaFLgnlbjq4xvY/v2AiiPLLqCWhrBrZufnSS0UsuIMAyhs1aqiX0QIXZMeaaadJ
PBTtRkH0DQnv3BMzym5VjlpDfDcaK5lJkdmwr3giqrSzX2/TiVR15qA5rYNaq5vj
e83U6t56Tis1+ERMdg47EL+4KNSsbU7fKGkYySXh9J+S/3aNJcxp5UpSl3Sh5KfQ
E+DTdjz1kwPxrv9DVFTUQ17NU2PUEmcCtG4IySrjH5cATz5yhjNZoeyjgxZqyuzX
+8mOi+YOI5gkG++4FSoqi9BSizWfjtlnqYBqgQIwUSzgReYMeqbYRk8dPTfAK4Cm
TZDRpdCZAgQ0ZuIfUCUrCX8fLRNs5D+6Ft/3BITGiaFYR5R8/GUaBB8fku2yfVIQ
7jmLdwnRb8H4TWsQuOdY37ghHN6RXPWGY2EdfkgsrIdaQOk3tvvmD0SbfdIsCz9B
gvF3YNuJy/smdQcs2Mirb30ZMemzdeM4CNE4fHRmiWQRCk34hFTYU74U/MMp9+9W
RVTeAURY0kviXAXaZMtuflJApqOHa+SwZz0VuocYRYrc8lsQ9EIXbzgfl+upBoLe
6+5RLX62GY7Bw4A16nQW7jN9zNFtMYkJDcd/63upFW0wjh/j4LXuG62Bt6xWPpT1
9iNZ8ZtaHDENjD3DSI/vvX1QzIjYWL5Q5QhxpSgByqgNttDNb40cyW02neAQN9CO
AIR7DZ8xEcJqBsl+h6M8CxGtSncjF57zuxv+nBD5LSTgu8RNnT+eTJRrfgjtntSa
bLu6rP8aC3jr2FQbcGVZx6qrAkCyyFDIOe4lYTxsviGS66DZ3+T+6+jFdzZXfebZ
cEVhnXDG5a85Fd1HUvVHWGIO9nEAGPVEFEkZjNI2rcxAGJwCD3IKK5dI8wideSnX
OWpz9j43DSRSM+lUc69BSd0162WGeT2c1rQOe7wzCtWITck5K8gyISlgQ+1d1/r0
oyIsDG5iW/+TvOp7e/avvmkYeXueK3IJM9+q3UCZ7bPXSwj5xy5+VMjXzUHyFtsN
Cfd97W/WNRVarX2E7UsiBpYGoz4pqhuQMbbMUPWHfFbsYfsEiWKa8OrzvWjASSk2
Ce9Ur84i2VDWb93jWejHl/xwdaWvFDtNhixhklRzN/GK9/RR7zXbBQJR46sVb/F3
v+vu34b3PxqF5XAa3YPPuLw1uF2gEyJg41D7CLiafTH+JfuExp3aSWpXynf7fTbw
nfuOSv9COtEI/NZdI8MIXHREIk+ZaELNMYrMbINE/qF1SGlKAhVjaERm1LhkRNH3
2RK/P92WCL31KCawRdfegYUZZcLPmj+R41OEE+nK1cMs1eVDmhutO7Dfxfhzt87E
TW3owhpQK3GiOpvXKdNkPYdAe36AsK4xkKlwn/8evgvJ3nsIQChzSAd5YDDLqlKT
HwLnkHvFkfupCjeDQuaD38gx7Bn92mbfPLRGUesei5CRbe8uw9h3u49Q41sJZHhQ
DvWOPqIAlR2Jv0GLmqicNJLQGsse2YukgMRGN1x8wEUGx0UvmqqDZzmCShx3LGTQ
aZ0D01pl09ZbSz0Atf89qeNO/Mz5ZW6WqTXliKur87VsVPvY+rqpBIcfxxWQJEv5
/rsz4gPyWScRKSZlgQMYdUqSHMnxCFJRSJVEZvpn+CDfllFFb8EBcHcQn0uV572U
GYeQv8xp6J6z8sFYg4Gy+kWn4fiUtb6Y4UhLXqnD259t43Oyf714vRaFzTwJm9RO
EwFhDWIKqUrf6S4bLpmIKsv528wdzZhty8E8JYVJaXBiFJFTBdPZxaPlqU2/fc2i
9hTMBwvnp94ZZzyw1hYvBY7vYLzqLqBwnjd5KWXpZK8sTgdxbBO4NUz1VfUf6Fhy
Ua5XuVaxNNH+bfuC4QZ3MLB9SzZSEKJXo3HlBCo2c/NuON/gcil0sAb338eEK1I/
QYHuyOxOS/PimwSuULK3ectkN/1s80QyDBBs+uJ+W/CxeSihXXS+p5obEeouyFEB
B5X5qeQdJbhY0elbkVILk+g1qBHSg3eNAEfZ0T4qkZn73dHrlVAU1pvjkTy0OAe6
V57dYYjxeDKqpjQlgwkw0l5UZbH7ZJOfm9Ow/kl9VY6SPzPC+uCKp3Mk2jVfnj+Q
nh4VzHQzCecXKDM/Kh3ONv/3nhPaHu9qO4z40sFO4IYazrlk8WTvtZNP16M0q6hN
4TK+OOra1VKBvmc8bWak8PDTT2HiUzM8TlKIWz3Ntrph3SQJoGRIuo8mCtazCSuo
PSNm77PweWOcUvRHSbGugrq8UvC6WORhkrjA9WBJRmUn2n3GmL4HSWV7fe4aDxEB
QHneaMBSihjFcs0UkpoM1wgDt7Xx2eGyX8vL93mFKyO5xz3VPWXkn9Xq+X9OHMsM
AaIVTSeqstLjfv1U4gL7ceEhYxOdMFVHdCOtE3ukx5EtisJo/iCaWzY+YOTeuvw6
RFAAlInjCTEew05It5FsqHWhHz3Ra/hZXiNS5Q3mWk2MHYYhYYgvVnkwjF6wR5XD
oDVVn1iRniiwYJpG4lbanqRWt9sUv1C2wmCtJ8enQ8BR/LmZca5cZXTlsTrhxFwv
FW4jditGI4NYC9hHkgUd+gdm5Z5psqpKgFnTdgFzR6d0nFuEimW4niolb+RYaWxW
QqfjhiYR0U3dP+1gmF/CXSAgiZvOdDw+ci1H8jxyRVXFwla/zilM3/qecJhSwL/4
E5cf8U3DMfAxug5g3U+/2/6nJKDKay5R+VL6N6jCRbS331nT3jF6lP15Vo7mOwNq
HKQ+2dky8abEkPhV1cFUvNKFyTcRDn8VDHI4bC/o19A9ljgsuSPcbvxhkYpfUfG0
f3Iy/TgM80jJdfKpucyeMaMBbo2lMP34oZfQJERxfePShc4aIYWoi+JMAPYxJ/PL
jmopuPgRigljyvRKmPeyQVBO5aAt7Ktj3bg1TuKgd7NYjBjcLdxS/BGNwzQSz9m4
D0m1OCUmXq2ldzlJDs84kzKRkyd824L5OoOzAQQkyLMeBDJ0ezfII2Vj1mpEd0RZ
Gvc9db28FRvzPiZlhifRVXh9JRljtsDpRBRZu/jsK6inbuTRtrdZ4H1eJ6rrEizC
RHOL+NDZotfF+nfqiYouI1YeNIVka/gvMvHyftdzbuRvouiSrbxHMVWGFfBq5MA1
sqlnv4MSD5GyiHAC+Mp8Hq8eEsA2lDz98+tKs9h0eo69AmkzkrnAa3wvE1ZuwvdO
ayngK8N49hrJxM4Sj2QHkeWIaY4+RqEhs9z9vG30YP8zCAUVKiEgKOw6gQvEGxVj
UoHYx0gUwWol/dF8ZLvHm1Ey78ZwED3D5dTYlOKYtsxfFQk4dhfIrs3qjQDP0Oig
pGypKw71QfMwsvQMzUYFu4G9aUI8m7wrLbTYSZg4X9DJaAkP4mHxhlWIEOyFg3bs
vi55I0TR121R/sH8J87y2x6iWpzVcE7/P4z30FxLpkuAOitqnNth+Rbrj8LZKD4f
X/naK2G6ohMLf973L+Khh4iV7gNv5zjqdbmV2kRxtck=
`pragma protect end_protected
