��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�_PN�2��,H_|O}��$7m�c��`�W�mZ��H���wz'�K�s<{(�*���w�%�:%�o��<+2?�=�l���L�G�n�y	�f��c]��g��77�D|��W�םfʠ�� q4���z��ص�n<S0z)��� ��]|������&(J��� #�eۑ��Nox��c6�)�瑹)Y�����sTt��p��T�j��凞s���<F��s�4����:.��� f Z*��R��?m�%�����Uf�ek�6��g���-���Ny4
�Z���l#ꄞ���-�Df�d�%��|��i�C��ٹ��o#��b�� ar���c"�Fۃ�l�9���6ތ��[�҆g����A�O4Q����hT�W1f��:
�z\n�s�Fz�#E:�9,���D������q���0h���z�E	{D�L�3���r!r�t���NgӺH�%�������;��y��_�4���~�7N � ��b_�RfZM�����}��(c�lO@H��-#/���,{M�R��4����Q
7�H�3d��EI]Kc��Nx���s!�oG��)�E������d�ȍ�� h�n�N���A�po�K:b,,8���"��fE���G�(̜$�������ݿ����_���I���*�3%ȣ)��[;o���2â�vv�!�\��a�E�q�_mL>|S#���� S�MYP�h�P�;�PV�O�s& �-3�βF$/����K1.\t��?|2l���|Ρ��G�)﮴e�<��,��ʃ�%ϦA��F[�/=��+	|�m��0�g��@�xZzO='��|w��4�/��%�T���b^����H�*g��K7�<E��"�K"K�*�G�q!�
����ΆAgV9�l=�A௟an3��	Z�������&~8kwFQ�P7H��ܓ�-�~�ݢM��PJ�p@c!N�5���N@Ê6�ͷ��x�}X|{���%�O��d>&�Bw4�b�k�n�0�߀���� � �g�e��Αp��p�N� ;g�k��cN�ڄ$Y9���ò������Ug��O�N��  �k�:;�ѼV8�t5�hGʌ�TYI�a/<�ͣ'qYY��63J[=4�.���0���A-!O����=��W3b��$S���S|+3쐽H�KbГ&�,.!�?��3�oI��bÛ�뫸�(���T�	$���Q�鈋���E-�'=D�8�,w/޷����EO�˝�~�$I'�x.O5ڧ�_l+�cq�n�[$�.a8ܝʂYf��$�Sy�aCH�f͐���g���1˚�l�I���H�9Rr D�2G���_�=��R�v��ĩ��ηLX~ԩ>�1\]-�o'�^�.s3�|}K�.K�|鷚��uy�z�)p%b�s�F�N3��d��5��,�&>�n��gR|�uC4������;g}���^�թ��]�Ao䟽 �}MC��܈�WC��ka���좌�h��r�^���i�]�6��ƻ�4�����4���_�n����{��h�J��QL��<���>��c��k�)Fj�/t��ɰ&���ܙ0����A���4�g�>�=�����U�v3����]1eS�̭B&�?�b�p��������ul���?`~� �s�α�S�q����y�J��/���v0u7�Ґ��'��qE�<5��]�H:��Q����	F���M#��_�?e�|~$�E9:xv�zR�ȼ|cʩ�*�T�X�e��P�}�'�if���ZS~�Ə^���K�Q<uq3�px��N�g%D +�����x�0�(mG�4��Z�nPVn�к��jz*G_ǡ�<�]�/�����h7���2�+L��V��<��fym<�m�⥐�]��ERQ��s,�*��ĵ�8-3A�p�up�oC��՟L�SD������Bwȭx��� �S�4y0���YA���Ψ�ۍ�P��Q�u@��ꚴc���ܭz1M@Ea�F�(���#��a���V�N�<IĊ[�*�㱐�{����[�T�`2佢$��#�0	�"��+ee,��-��Z ˴:�?/�1,�<����R���'��`��n��T�����{��% ��_9�v�-�Ebl�Gp1s+��\'������t��u��/e�&�	-i�N����<���zE��U�V��PWS�{h�9���[��uE�|�ݙ�,JA�p7cw��%X���r2k��S���Qoꉶ�-6H���A�N*�˻AE��c��6��pk��q�?�zɾ���d�C��&_�;`J�$��hzk��-�`2������]h��݌oz����Ջä�t2+����s��U��vI�
��W��g��g_`͚�x���}kM� /�ᑑ��6��9=���\g�@F�����P��������z����T�]���!��&�rDW��s����e�+nWٚ.o5����5����rIA�=����sl���ˎ� ZP1����<tH2�=�,���v[ͣ�<�O;�eF:8S��%����c#��9����Q�|y�`k�5㶧}{"
�h���y��<�m�3	0W��s�',4��8liT_�4����]@�;�Cs�]�����Q0�{�M��VT�g�*өc�6]BM+W��1?��	��p�w;YO?�Lx@�%�p|��\�l��0�;��gY{uqPFi(�J-�������i�����	�>����e��Ŵ ���K|k�\.7�J^�$?)�C�.�%fR4m�4��;R�@���h�/�H[�d��.�4�nr�v�>F�ѵ��B�1U��LV��$����Q���n_*
����.R�/�Ҕ�������D�s$f24�^�T��
X�$F��V�2|��c�����*t�D�O�±r��d�K����o�y��]�OˢL�H�2�8�P��:jn�c5T6/�w�͒M�2ɽ�c�5�d�N�hķ�KXZ�F:��:�H��ӻ!�U���E���/S��ft�v�H�ȿ[(�=6!$y��?���F�z��:�G9]gK3[�c�Y�.t�����)q�!�r��@���rq-�Y�������.^⊋qmF�ߡ_չ�2I��;^�H�
H����C�+��'~}lqg�1��Kٽ�oZ�P<%Ą��nyr�^�p�e��>!�m�{.o���9,���$��ٟ����E�����CY�_�D�ľ�������:�u�Ⲥ�Q�jk����%:�I�rΞv��z���	F.�E�13�
�K�{�f A�o��:cRq����U ݮ.��U���o��Q6�u�	�/<���ރ�A �L�������f�`�krVӻLu�nR���֍ٞ-֕!�0�3�k��<FCI�Ӟ���gQ���O��,H�~�/�����w���Z:vC�w�Dx�% Y�pw��HϮroD�����Y����{8^�0Ԛ���[:Kq�]G�qTB����]�Џa�������������#=�,V�����٫�=t�VD狸�6�; �h6�XXW�=���v왶)��l�j���닜�Y�8o��<f�h4D[r��&$@�+�*����I�m,����c�E�.��*?W�ظA;��b��7YQ}'C�H5�O����ye!GD	0�H}��z�|�C�v�^���,4�]S&?��*�BH�"Q�Zʟ!�|�O/\׻ � �rtτ�w�4�	�9��0���4���˱������ak<G���~I��@�2=( "�7H&��O�C��d��G��dg���|�o�fG��[�!>(؊��o�*�²]�qO&����q雗�p�M�ybl�H�XX���X!�L�Ŷ.�,�����m��Q�V�'7�qV�ҳ��sb��� �d�iģ"߽9��x[Ԗ�	|�nNkI�KT&5��Dk-`�����޿�ڷt�����a�0���89�󕕨������V� Ҏ��)e��l �"�l�c�N=_y��
�P�F��(��p�sf��MU�n��Iyv�>��ԇ�Q���Q�C���Y�S��W
n<î�6ġR�]U�v!�(����`!�{�*�Q���?C(J�`��J���*�5�p��iy�t����������&�z�6F����s휖H�T�%ĥ���sV��9G~*���3Ѐ
���L���a;,�On��'���@��dTa��0�����Z/�\j�G漧��w�$� w�z~�'��A��a`�P��1J+�4���6���!c!�x��ǀ^4���/op@�I"C�D����'�:Y:�� �7F�3�V�zF�pl���R�����;���@��(L8���	�k����`Vt�I�� p�=JnC]{O)��R5��$b� ZUB���������Τ�%���z4-��ϟU���g��H��`=0O���L<�#�����l���ye��B<>Ks~uШ�I�b=*/�fb}z������G�.vC�w>����B���5%��t���<�(� �����tr�;�]�s7��"j3����v��v"���<E'�WPH
6�>e-�e���e��KO,� "ڱV�X�w�lH��`);rU>aSC�dW*h�H�̕����E l��=/����|>���&����� �<����	x�f��"D4ߡԼ=�{X���/+ʢ�D�U��գ�|z�qwh	P��훆����M�(ITr8{��ڳE�C��!��RLn`���=rL!�A�փ)=�["*���L6:��O�{d��ҙ�x��1x-�"���pȀk�@�O��U�����P�ZEE�(Dh�U��e��aiX!��>T�&� n���=����Iئ��)� _��+�pCL� b~�E%�=)��e|�m+�V���W���6�72��K����%�M��$#�h��Tu���@�DWk"
�R�ߏ�I�m�M���V�1��D!�Sr��>+��V�4H0�+��<.j�h�*I��yT(O/J2���廬pr=� ��Ҷ+�[=��N��J�b�Kq���r��J���.r?=�,��f���V���/!
v�!ԏ�%?�p�I�h��}x}x]��J�NV�dg���=d�2_�㡃�����6�2��lT��#*�4�ϖHa1ٟ�d�uzX�Z�gj��xd�eX��91գ�B"�)M��:=s9���*0_�x������dy��'�y��1��;l�������Җ,w��������eL��7�����m\R\���w֥�J6M��	% *�j�/Z_f �ά���� �R��m��]���tk_�A  ����Qyn��"�k�՝q���h&�CH��P3J-1�E@�F���D}e0��&�0��y�6 =N)2y�Kۅ�H�mVQ��)_O��̎���"nS{���V�[�>7��]��[��|�=�#�}��})����7����VQ񔭷�yj�QS�Rt�����4�0��;m�P��x�Dq<�SltJEA)Y ����� ?=�xq|�.�h�j10�,�)YP��7̤��e�,+��ϰ=^��Q�KY8�y���Y�����ʷ��M�����:�]����59���$ly�#�.��9bd{?�z�a߰��-L�u8!g�F7��'��%���6%��3���R�����X%�7�a԰ʴ�f�a�&,�j3Gveu5~Z��d\�1�u.� -�e�i�$��'^�����[b�1h�r��=�E7Q�6��߼S��f1�9�����������'3|k���26r0O�"n���;��YKG'+ Ix�/�%v��1�v6���H�\<&C������h�j\�1���FnG�QP���b�qOX@`y���Vd��=1�O���QŅ�B���Q�&b�m���ѷ�WU;9lڔb��oxm��	��jo�_��Qdd��&�:�"%+]��vE�:�rq"r�.�twpa;x�N���%v�Y�<��%�i�t�oX�Dc��g�ߥ���٨(�����UPc-�L�F���焧A �����
?a8J#�	�|���g��P(�7mX��~���������?�I�ʑ��C�t��aZ���̑i.�Fy���*I`+����O���Tay��Jv�Cˊ���(���Ӄ�� !h�(�6�L��ۙ"H�M]� (.��2s�F�G���@��G��	Ϫ:�>~y��8�Y�tm-����SZo$���A~'�s'I|�>z^t���8"{���b�H|��qáq�2������J?���9�w��&�h	M��*SqyB��l���V�Q:�!m�F?s@E�0`���%����a�z?9J0�hC�L64�*WII;�[`�sFwK�\�i��e�{�*W���?f9�`�a��9m�^�Z���L�b	L��Xr�r|+�AE�\4T�R?пJ��%�����Ŷ�*���;����p=��X���R�<u����u{����&Z�����uZ�\HW:�p���m��D5FY��ݰ�ڻ�]�}�2%t_FoA�.U=�KF�80���X�s�!쭸t�5��q$�|m�C���D�}4�J#d�VE�l;�<���_6̃���.K���G��/�:0"��~��!�y���:i��%����W���q"�7�J�jp��YL�c�w��z����#~�^�|��x���;���8$�7P_�~��i�PE�#��i �����N/W��EЬǆ�P3��F[�Xu`������g@�$��ms��2����Yњ71���'��l���hY��=@��K�Å�pL�����ZMH9��*��Y�=���.�Ƨ���d�������2�8W�Pp&-�~�#�����ӻ�-
ڻ��x�����ᮺ�}`]?֚��{��Q�&����hf|�>Ĵ9sg���p�5�J:6�+��GP���/H�s]��"������(M����B7<��B���X��*��\������H5U�Z�E�%f}�W�4F����cP]p���5,�o�����	|�i^b�ґ�[A�#nfs	f8H��W�M�湦�y���ә����t�|@-v���~��Nϭ�T.\�$Uk�Oٜ�	L��1���L:]-v��������� Q*�{	W4�L��,�Ǆ$�Ygy�&��b��u��N?DR��H��M���L�gm�uiÙ��]Цs�g7䇯��T��8ɾK+�����������4��Q}`�F�ɞ� �$3���u�f�"�Rn�U������r���c�|y�9���y�ʃ;b;g.ƈ��<�z��L8f���"؆�B�bKj� z�c3#n! R�-�S6:Y`�We;%<��G\���7������L/8uA��&�yf?y\�/? �v7g����_B��?Ck�Ga�o�U�~˹D���)���������a��=��x�Al�h��*Iʾp&�hSeV.�.0`
�d5�{�h-���|�͟t��2�D�|'r��T�K�O���q�ł��=�ѧF5��-f7��>�X_=�:#6��P|W��l)V؍x���%p�k�Q��O1 qF类��=/���^Zߗ����g�����:�����'"T�C�,��� ���:J%������4���B�=��u�r\á��,�\9��@���ݢݸYj�И�E���^	�5����jY��B�}���9�2�+����\%�ۗ���>���D]�ۈFc�7���a'��55#r�<�H<or�L�����D�i����$`~:A3`��BqqRn��'�����{p�9�8%�|�4��\��A}N�S��A:YxmХ��y�X��2����8D�Em�T�>���Z\�����3�)�pAl�Q��r�A�R�'��8�x�Ȱl[��^Sϻ���Z`w?�������T�/5����Q�Y	w3��;��w�|�K���y��5~���e��b�*4�bL����ჳ<APG��Dr[?ϭ̌M)v��;=��@&`�MU�cw|�$cfi���/{2��<6(��s���I���n��'����X��> e���L;��ˬ.Ƙ�>���7t3Ǉ.�	6�i�Y�y�Ddg�0j)�^��V�7!Y�*foVi�m3k̈́�tc�8��Ԋ!�����.x�q�Bo���-~eJ�eL���>!?*t¤��niDՠ�C��(d���hQ<���-pey�'oRe�Q	m爵��"�� �	�� �
�P�ȥ	= F#��^p���,��B]�@����g�a�[֕������1�d����K�j6�r��+7�u�[o�/˅��z=tF��A��=�Ӧ�*��Qi� ̄>:���#�-��^�+n:�hZ)���m��c��%��L�Tw�!&�.7L���� ��Z�_A`}W��7	�5��)Ыil-b�IĒ��IEӠU�o^���;Z�������x�m����ح�f��b���
���A�<�uӖI�"*��%��l�r�dL�!.�G�S�z�I�?��!K>[r/��,px%�.����xH͡®��qW�_/K�9)����3�R7$�[b��c�.�ZaY}ٛ8��J��� ���:MK�gZ���|��ф6=p2�p�k�4�G���5�ֱ5�j����ӕ�~A��6���s��^���H��ܓd�~n}��(ڠ���0���T,S�ͮ��0��b�f7�Y���Cb1*�H�?%���o׿��]��Ο1I���킫�X����6����$9=�qr����D�=/��z�V&�R%J��RQ|���{r�8�x����]�9��x�9�֙ �V3�ժ�<�fxo�M�4ڤD."b\����Z.җ�{w;������\93wuI���F2���5T+a�iRb:���D�o����3�X��)�쑊��;�t�PJ�!��N��i�0��ed��±��q�I��5���{s�{���\��O���g_	sr!�9��������@�mz�S��1>����M9�����P���i��N�x�ґK�n}et�F=�g�(-i�0P��޲�W3S�d���0����7���������s7����Sy����BJK��B��CU�-W�c釟`Y��^r��7�U�� e���kN����)�X��w��kHQ�d�R	�e��jpG(� ���lD
D��b�b��Oi{�E�N��wt+�$ۖ��zs��j���4B��N|�o߉��d*�T{�٬�:ќ�����wo:��K4��->hkE�����vӌo#�or��:��i؈��"Ȏ�gPX���(�Ƙ�F���8���|���j����VT��G�cCQD�m\��>0��F�%��;��C~���1����>�p�5�����t�m��%o��	,�j����1�� R���'�1���$-�{)����6�ӕC�ʥ�`Gv;g�Ϙ]�ƣQ�J�R�&�ߣ9�*tk���]�QF��'��Pee�D��B�J_߹�U�'1䷸3�I!�l��y�0OC�Ԫ_���@��_\�ol���
�O����AK����s>:�4�������Lg<�{�
���O�%0e�}U<Zק>��J���	��ʨ�v�"٬��f�k'R���y�/4���a¸Xi�"��jT������jS�Ge}\yB�I�^mbld�f�>̔�\�kټ1�7�L�!p>!�u��po�B�.A���nŮ��b	�'���j~��"��x{����NA�܁$�r��z���)���HM�&�o)+m�@�@�Hp(��kI��T#!�ˤ>�&�Uo�\~x���r�R�Y�7�,�\�d����Q��|<��w�Tw��%��w36�ط˫�˘��	�#�{)n��)��_c��=7'�I �#���K�О(&��m�|s/q��; V��o�d�� i��d�q�b��Tݮ*\�����r���"�G�U͹�B���� n�����*`����ڵt|��i�J�P̆�4@�`�$y��ם�od�Ħ�yOq52}����%�F\��.������^3D�N�B �rI��'-��@N���]�w��^b��o�.��{��ÿ	E�&�D[]_m�k�Z�K����9��E���+A��ٸܛ��[��ʪɂ��dz�b�$L� B1>��u�ܥDA{����9�a?z��L�V�g�D���K��[pz���txgR���"���L$<YX�3>Xr�����cYQמS{sI��w�R^,ǽ^f{3Ѻ� �Z�K1�R=�ț�12�,��z�Ĵ��ħ�p3��_.L�y�ۡ�w��+M���ř�����/��# 1�k��3�� ޷x��1�-��m�e:�%�q�{΀��s��"�����1��Gz8�ͧ�IoJ��?���@@Vj`�7�W-�nP��Z)��@����]$8��i�*|PJ�K4���p�rs��[�jƖ��
�:r�LW��~��x@B�h�O΍��P�.l�4��&��B%I.�Z�е_�d�L߽?Il�O�����K�2�h��U�+k�z�3�D�+xZ�'Ə`B�_t�d�Y�r2�C���hR��~A�~�Gvq�����~�	O�7�'�(D��;��C���pg?Y�����8�YS�D��!�i1/쇷)+'�MR�X)��������jͬ �2⪰��Vsµ��GG���01�)P���-�(I����,�ә�?�cFҫ�}4���h�?�]�WW�"���Q���R	��v��:w}�\˼��i���n���#?�n�Q-�>i�#F��j�U�* �����Y;�Ƿ�1���g����'lU��`h��/H�-1MA�a�cl��1q��R�S*e$&Q���7,�nknH�-58�xϱ�i�N9pc�]s�����正8���%��G�a����(EL�k��Ka�P���ժi���
�61#�ó�lĜ�+>��C�� ���jY���b1A�!��b���X_���#����)���`\��^u��5W34+��@\9�d�Q<U?|���lDj��L��4Lz)4 u�躲?��4��$�9�l(�S��Jo��}?�����D����nf�ذX1{�e�'�l���3��kʓ�����|��PP����O�?-k�R[D@gTطo<&y5�!(�M@`���|�Z���Zw�|����gT��Q��S���,��%n]`v�a�?L1�w������u\�6%�α)��frqr��a�RF>8y���YŦH�]�)��Nr�u�,��=p�dL���rbWAw�r�m��<��}G7��<���2�6�]�Gw�� 0T$�\8��};��gxN{�?�V�kA��=z~Z��Y�Ż_���M`�|�c��<q����J½�����
љP�9�3^���},�j��P�Z߬�������J����{m�O�����}��&��R#xX6��x���s� ��@6��'���k/?%���#K�.�� �r�&;�+�j�EaC��V�쵥�C�ʝ����H�g�f�J�)<4r�_ґ(M�~�?�JO�{�n��8��]}�i���O�(4r~s*c���>�i�C[d��~�x�,D�[m114ò*�v���{���ß