��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[������0\8�J_R8�C�{B�z��I{iE9�Ъ�+�x	/q�{̱7\j�2�/<^�~I -t����o��1
�Y92AY���u�)H(����͠,5P^�V�Z�u��rw�`P�tR!���	?vM�i@YY�h�S�i����ȬNJ�Q;��m�ݸgF��݃Z��^oC�g��g�`;�'�gA����v`��#��^��PD�{"�pnfN	C)�=/Sd����I�V���,m��k�CCQ�q�Y�����ٰ�]-�aʿ+���rrI�Ҥ5ՔY+�(���ae2�˳x@䒺QdF�4�D��f�@��4�P8�Jm��zÏ������bUO��Y����>�CO�e���݄0�BD-��`�K�P��v}�{L8�>-�c����3������$��X�~ ��=3�y�$�
�El1P4o���W�����VSt)^��o[���SmCƝyZ:&��񅣚�GYx�K��1����ĻS��֡)�*B�wǡN�b��h@sv���\��|�fw��'-qW�Gb$Ȫ�*b$H<�t�Ӌ��?Ɠd�?��B4�}U�uѨ4R��q�I|	@��Tm	Vs�G0Ֆ�쓖V>��w��Y��s1�]��ǖH�~@ȩV]W�e���&!���۲p���!�WT�`����L�KJOW�ry,l��Is�%��SLB8Z�!x���-��p���4�!<�2�~��&��ڬc/�V�|4�[~=�Jq��/4�!q��k�ɡ�דC��7����Q�[�0��A9]��F��M�x�}�w��i@cr&��V@^��_ߑ��gM���PZ�G\e)� Rh_��}a� pBV����F�ū�^��Rዡ���Y���c6�'0EAe-G�- �n��*pk&Q��&8�M��	%f�BX�e!i[Xn���ȅ:��R������H����89�p����F�q�
^��2�YT�m�*���	�����A1�*<��k��Hp_EЊh�󵈏TƷ����f7p7@5�бdcI.^|rw�����ݼW0�}�F1�w��w��G���$~?�Ѱ��H!%�ϲCW춂C���Ք����L�)*k�v���:D�D�b`-��\�]���6�����N����H{�쮒-�ǞIDj��/�O��JK@n��;���kK��sc_0�0m�m^�KJ�M@�D��� n��?��X�yC���Az;�����$A8}`=��LE��{��兔T��x�$	�TT��¶����\k`�!��},��Ť�²3�肛��|�ʏ��C>�G��:e����-P�q����С�>���]_�5��ηY�|�����8+���]A�l�L�\�#d�1$c"P�a�[��� @���q�)���'[���ُ��e�!]s]T�_Ш�K��U���xq+]H/,?b��E@� �6p��>�8ն��dH��F���a�`y���"�P}6����S얕j���u�]�yڜS�]��]��<���A������㬨ع
���9�Clo	r�Qw���<�l7��ݰ'�@������g��a9]�/�Ûf;.�I��vF�B�V]$��UU�Ə�ŗ*G�/��/������O�ӂ�X�ڣ� �ko3^q�ao��׺�fb��x�
?�6+��%�p���*�Ⱥ�(xW@6�ݘT��&�;�2�h:�ŢZ�����UVF��Q�D��IbU~��#�C6�!MXڂZp�8�A�o���K�<]n�\B�'�]S��C�����@�zJ����'yn����٦#�\u���^n�u�
���T/��QVϨ��kt�f�7'mݝ������U/��늣�[��]��)�U����YpN).�ay��1���S�ݜb��s�2ބ�\p$�����}����g��� ˝�����Yj���Szkp��*?~�c����I�����.�d�^wc��b7��-� �u�(�aDu���0E+�D���X��.{@��0���k��1,,�1�%���П����
�@�jj�g�bl��=�f'�i"�oGI7hL��)^���?�}o����~�kP$���,���w��h�j�0�	B�BU%|��`�����AJTEe[�	R�nn�5(�#A<����S��'�Ӄ�4�Z˄�[��B��&;Y�0l��n\�a��`� �^�ZQ�����n���٭�#�-i�Ꙋ�D�lj+��Y�^���Ld�yr��9�YRċ9�Ƙ���\��c܍Ga���j���3g:�~wG¿��Ä-�0�],�5��>��w��#�Sِ�(�y��`���N��P�H ����8��Ye��ߌ�l?��:w���N��ZN������Hg',��D�Yϫ��%�7�{�l"�W�_Vn�@d�����m�hj&^6�4�ޛč�+�G��rc�I�?2ǻ�Q��{��B'�����a^��ϧ�h�FյC׹�M��CR+��T|����ns�^�˥���@h	�P\�{UDRg�`�;�n*+s(�j�6gς���P� p������"5ޟʗ�N��Xէ��ǚ_��rB�B�F��S�`H=\r��"��;n��������-b������5�:��belA`+CM�>���mA�$�F�F<'/#�#���m�K:��jȆ�,���0B�FҌ}ձ}����pq3l6pә���'�+ժܱ��e�'2h�#�HT�8bx�AW�r/}j\t7�����^��0�,���k�g:R��Wk�:`
x��f�vB��jX0��=6d�+��5��,��
�!�@�v�4V��h�����(gO��J�YP�;���-� i��B��ك&)it+�|����u�Z'�_�x�P��ES!�����W#��3��Ĳ�u�U҉2��-�H�����)�,Y뿝��/5��~4�e�r�/�ꄆ��͢��~�Hx#�T��/Jc&��F�@�멪x-���az�]a\�{�Q9Q�c���Vˈ|\��0�D����W��h�<�TO��7ʸcd�KιDM-$�nW��(��.-����v}uA`R�:��%ܞ�y��dri�*�՗��ص'{�u�V>xQ���Y����*��weB�.1����?�r�D���Qa�@hiK�d�
E�%�kF��%� ��ɠ!�ba�$H�� @\4����;�aq�s�/I\c��ƀ�=��N��.҈	ԯ��ɴ��7���9����W��jG;U�v�����z"�����d�o���rf�=���:�t�ib��il*;�,��*ʼ�N�?Dx��B����e��� �t�^���jG��L/
Ԃ�"��<Fw�p N������H�S�n�b)��_�'�b/��jV�ޒ�k�v�"��ᩏ�'9t u�V�襆	�sE�CV��:`�13T8�A䇱������w��]�X��
әu4���Գ�)��-�І�ߧG�5;PL����R�xvO�Bh�h11��*m	��Q�څ�P'4ޟ����t�z��U�y)�VO]�����#mi�͙�W`�E�-��VY�jFA-���T�"��N�bLUC*FU$�G��aeP�3a�F�+�N
ա���d��5�� ByԽ�S숂Y�����/Vzc��೬}�倜�����hS��R���9�Uǋ��f)��_f���X���&h���
���P͒�[I/����Ĉ�Ķ%��IZ�ƽ]�#y)O��>��^O�]Ė��k��Ͷ+�S�̂�=9/�*���ԧ�+�-��d�u���hL�ϻŽ��'��L�ր�#�W���.�(ϱs�r����xS ��M�W���ۖ�E��<a�w�F�)�w!��К��!,�	y!B��{�R�Z5+�~*�O���c�;���yY�5+���&7�C��(�nO�y�!��R�|�$fE��˃�j�����;0�h
�q����%ڠ�N� ��M�a9���qEy��LT4�P\첔��g�[��ˉI�����x����G�d��	�j��D�����K��)��%D����GB;�9�@�3�穴�!fԿ����XP{XO(�����s _�YK���\�f�;|#�x�'�Ad&�ע9'�$���ΰ?1����+�����*��L��~_-���
��W�F*ۀ�z�;�ah15�y��B����~�(�ݡӫɗ7��L�����c�!�Ů8)�-���c378�1���+,%}l֢�u��fi,�q��+=w����$�2�P) ��W��]����rp�]�;��U�=�O F�a:��T�|N΃�8s)�8����*���I�e)�wCNq|��R>zдJ1T�lk��0xք�V��f�m�{7���Y�j3��I���Y��8�r)�a�EGxc�3"#1u/<X�[����χ���ؾMȗ�%�};��	z�V*q	�!�-(F�@`�b�e4����p!8��ߓ	�V<�0���FՔk[�W��U���z��EoA�s'fטd<�k�!Z�㭥-�Eλs�J�i#�i��=��ݨN/���y��(GNs�m9뼩
��vvp0��!��4nd��񌽠������W@��rt.�&���ڱǀ��ޯNq{�P?���b�~�?E1~e)ng<j�+�������j��hN�}�D\ 
����HQ_��!��<�ۓ�̓Ќ��}� k�Y�#�O <
����y�@��Nk���Ln�qvs@5ao:L�0x�Պ
ض������}����7��c~ �ݽ�Q~aip�H� �n�&���JÍj�<A�9@�0�k1~򱔽���裂�4�[��(G8�˪D��������S��o"@$���g͓�]'%�UN�c3gy�ޮ�����U��� ��>��弙�]��y�k�F:Kz�j�x�%	4����缮�-�eu��c�.@�ٮ���oq�2�'��#��;4{b��^M5��k��c�<�A��mHR\q+埔:ʹ��~[�pb��z�i�Mk���Æ�����
3�K��RǺN���wS����z	�^P��,i��U�W�����*��T-U�.Xr���X��*,�f	l=v��G�X\�W��P�L�7.�Exu�b���\�hHbV���ǉ�Ĳb�Z�:;P|e;�)T#��)蠱���Õы�  �u	>/��?D�������N:�*2-+<qR}<=�t�% `
o5�w�/�&�Rx�m��"��i�*����6��
��pG	�8sE��޽�5�@K��+
�{Ù�����_�kێ��.>|���k�ЎŴ	�bvG*f��de�ϋ�r�5�����	��{�?�7�*2�^6��G�
��XC)�;�U+�S�酰��}�.�8��'PpmKm��H��q�ŷ��p�cx��M!h���0k�ʥN"��g-����c�NT��;�{ �0�!�r~i��=��RĞ2.����2�l�J;�<n����4�������`7�Z�$A�)��&]W�	����p�f7l.̣ǌ}���ڏ|�Z�n� �k���?�6o?�Q��������� ^�wZ�t3K�ql��ӱ�lM�s����@g ?���,����Z��v�EX��-��\R���:�~^Ҕ����_-�6
:h����Āerc�x��q�lP�˒�Y|F��K��˦ mb�=i<`8��#��vaS���%;\���cT��EM���7�{��X?��#S��(;;"JE�I�?m.�Flc���S�L_��W��Zc�� �Q���D伻���_����|7������X�y�	����1����,��;���'��as���3$�D�~w�G�F��#���G7t��ä���x��x�ڏ��["��@��=�7�收����H�J�pP%��v`:S��;�
�
���G��i���X�z����͎��#mEc���b�}~��R���Q������Ww\�n9�u�z�����.5S��-�#�H�/�-����^�g<(�7)�K�)k��iI1ˉ�k��X�RoՠP�d�FZ�����E���ӹU���;�q�#��|�t���7&UF�V�Rh�����hU����V�P	���n+cU������lN}X�T�M��Lt60�8jk�"{���VE.�%�ƥ���`�����fTb|����֡��o��iN���a�
��L�w��鬼\L�c�}�S{5�/�s��Z�Ѡ0t�8Q�����'Ȥ!���x{�5CϔRq�o�͢��_�с���!���|�
ͨ=�5��0U�rW��v�$�{�E�bII6�9��������?1�W������na!�0�p���P�D �u&�\C��U''0���/x��vo��]`tQ�-�׬�pQIy�3l��Q���m(���w� ;��)�΋DNfRC9�>-��g�ꪼ$0����1�2W�BDQ�^��s��By��I�8�;��� �����Oi�l}ĻTG^�|PNF0B�����Ӆ(�T�ɫ|�`�2*�3Z6�|������4����.Ǫ=aLSj��Ù��y�u�9Q�~�ɿ� /n��r����x�^��%xW�Nja�.�zfd8�a`��yZ�W!�3�붯����Pwʜ�*�6��"�n䜓StB�7~��	}Thͷll��g�_h�7Z�l"�Ϣ���XP����D4�,��S7�%�H�׸�ei@>p�S��&��,F!I���c����X��9���h-���t�[$������E�TM�=��5Y��7#�̼�Nؒ�2����9�z�~�%�N.�p�m%n�����ح�|�oV[�≐%�y�S���n��؅r�?}!�~"Ra���_$.�Q��R=��gH�O�g���e~Y~��ƻ�C����jKg�V����_0+�q^}Z8��	�"M��]O�C�5��n���nU\�+#>�J�cjm�_UJ�׊�"E��s��gĺ?T�J����ɰcw��H����e#-�팼_0���1ǚ>fjq@��UWr\���6���f5�y�A��5'�\��{�8h�+8�����6?c�2��k�v7�i�2�5�h-�)�F�$��Ġ��&��)�.�BM� d^�ao�wjh��#�v\�.�>�?���v�2���Ef�<Kx�V�|[�J� ����h-S�=�
��g���BI��8��S�c��ݺ�o��U&㑲���/;
B���k�R.�z��F��Qz2���p��<�j@|�l)GI����H.d���l�5�,}<�M:�����L]���S��#�2Yp�5D?/�vmH]�vP����p.feT�u�E��Z�v��`\ʺ�yc���ex�o�g9�=�&�xj�[t��~p`Vǝ�Li��M:��ҷ���m{�܀���R�NE+GD�F�Ҩ�ڐ)��̾���mTr*´
��8~i�H��{��+M3P�V�8�D$���/�HB�W�*e�~�מܭ&?�U�,|��g1�Q�[�E�vU�t�����{��\��e �oH5BzRl<��L6J�ȗ�G�]���5P�GUg�)�X�R��i��*u���c'���7�+G:����i��]Y�ƛ������O�%y95V���7�E����l�����^�v)/��R\�~(�w�foh��(e�$bCs?�3��h��H��<w��_w3KEĳ,T.L	r�M���X�"Ot����!�����0�9Y5�KL�+D���o�0>:Ur�W�6o�%�D������aUxn(��"k&�~VP��s�oH����id-�m?����@�xw焹Q��\l���4޿�3~�ޜܯ��/�{&�Q�Y�.}!
�C�!���{�SA�-c�m�n�/��?x�e[a$R�7���a��{���*�e]��h_�/1J@�Į5Ѫ��!�9�a�c�'�9K��CN����r�j�	�ߨ�$�m�C��J�Ҹ!ґݿ��Q?^���/+��H��,�zԭ\?���x1�DmJ�Iv�Z�<Su��+</��>�j#!^X�g���������4��-?� yRIq�u.n�f9�- �{�2'�f�=���T��W��C��z 3����Qy���gi]�����:N�âƤ8(>rOU�u�ƨ7�NA���2�z�s|��,mb��'c#sRX�	/]b���^p��	ob�Ĺ���.Sࡳfә��HX�Q�]���D%�L3���@2�s����\�s�#;�ɐt#�_��M���Y�b_"����ܴI��}��	}� �����da��as�[���St|ou���~.^�P��pj�sD���-�r���q><��ĕ�l��$��ء�����{�rɢ.O'�T�v���X娸0�Di�g�nȓW(�g�VN�_�	�p�Y"1`��v�QJ��r�j�,��j�!!M���Mq������ (�4Wќ:2d���WGD2aH�}1�1R&:
����].�C�q�-�Bpr�hю S^�����T㰎E 2"�6���ˢ�ͫ#��z��;V7����&�x�o�e܌��)�
$tw���#�K�M{n����[Zn�l�u���W��o�+x�~�2�+/�D�^ր�� ɘ����2I�/~;�-�����
�W�#�IF�7*�'�/w6˛�m��U�e��i
�Oy�=<6�эvÏ����zWd�"\���<U��[��Qs���}S-L	fA�g�[ҹ��uŒ��n����eF��5�*��*���xzm�2݌krZ�\čk,&Q��i�pyct��т��'�q���%�ΈPdm#k�Y�b���iLb�~��ޒU�1m.��y]���]\y�B�-��%���}Rh	lfc�zd�M���H K<ʨ<�jӖ�)A��w�u<�X� $޹�{�D�Y<�����M�)��i$o�r�	lCLQV2�fs^�3J_;_	6j"���6���*:�J��L���vS�b��z= ��9���Qw��B�n)�,;W��)�XD6ґ���Z�(�0�d��G�^
M
R��/�d
շ]�|����s���*aC�%�J�?��
zxot4�A@y�̉L}V�漨�S�o:�-J��}=�#�G�j::�>S�#�d�ǨT�Qw����><>�����[ƛ�H���F8�F��^{������ڝ���b�2�R�������ĕ9�a�C�{��d��v��@6j�v��5�����������ɮx�"1����a�(7cz%G�j}[���^�#�|��$����DRΧ�H�Y	���W�齙JE��n�3����B�v"����E�o����}B� ��w�f�e��m�Z��P���'9�v�@�&S�i���+p�P��� h���B���]�Կ�O�|�K�-�n��Ά��(�ɇצ�uTs�,Q/���-Xz*�v�Ri�`��!.��-/�Ȕqƚ��){�$=u#��__�1�\��[��(��w#+����9�$,H��NJ>��cf�n`u�ƭLa�6:O7c!�Y�F �hя�G�$�}�RYn~��Q�C�aM%��� 5�d���yv��W�)��-|
�+c@���$�j��E���lW�������'�<��|��	�&��
R�F����OH�4���sۡݷf[̨t]_b��Wr@� ��O�^XLe���&��:=����Ĺ/J?��j#�pa�<ൔ$������$k'�s2�����'�Cqk��t�T�Dg؂dʺ�J�?�?��x��]у�_  "���h9���/��G3^k���p�5�S1��W%F��\���4��ҡl�_��E�>i_��z6����E� �_H�m�m��.}{�ȏ8u�3o�x"OS?�s ~�Rr� �#@� ��3k�z�����2�=�ä��&y�ք�+����W�� �`Å*��g2y�%�5��d�p�$��s!5�ck��}��c�D�2$�R>����,��%t�1��..R�ǿ�9c#� ?{kU���t��T�����;[�$�������[����A�������I*C�u�GI%�ь��\B��Æ�'EJk�h�S$�_�:�
�_���,bF���$�]4CDm1�m�夵a��4�ӆ�uZ�ӦWI��	A��s�OP��0�Ͳ���J(���!Pg$��+���J{,e�`t�͇��R``��	���o�DyO�L�����6eǲ�>Kc��L��$�A� "Z� w��B	���2��0��J`|�s+h��Fe�Q�z�A��y�5̔kre�[�2����{����%�G}��5TAǿÔ�y�����֍1�2ȗx"Upp�-������;V�xkD�x3�-�̠VLҎ:��.���DPDAׁ��ֿ�&-��n�$�Q�f'���`�����zP��(�U�� n�<T�%�{</>��� �ŷx�A���ｐK޼����<3�2P����z=��MLg�k�#<���Bm{�E��x�
�J�7���Z�!է1�竞��y�k�&x}��ӀY&��>��$�4%�����&/k�����E�?����a7��)��4<ї��f�qڀ�
���S��d^���j+��!�����p���s_������`��c^��mz#V籃/`_�i��ao�Y�D����*�,�~�����Sސ���I;1��������-�(K[�u�25)W^*��)�����RBl%�3���$%���|{F��o'4�x#��|&CAOHﺳa��'9��$��0��A��a�  *fN�K���>~,KkC�c�hE�?!ґ��F�xH4O����n��I�eF}[X
�U����b����;[�W�L��xFos�Q3=�DJf/�S�x�T����@7�
G:T �X��z�d��)��#*{�\i�R��	�������Bf������Sx*u�UM���L�ʨt!�KlL�?])m6��wA��Y{H=���܊*UB�i�MU�t�D���КP��<�ݩ�z6���{��vp���i4J��&�/O�H*��z�$��mpٱ�ӂ��W
����r�ڈ�N®X3XmDG%���7è�����D�$l���<�oW�K�ݮf>\NOa�fm���A�j^�H��'��J2��y=�5r�5�����*�=z��c�md�4Uw/�N��%3�ll�%,��~I����JoX��~�jL�q�B���Oy>�qe��0�	SL]�����r;�~;�Mk��Y������X�?�q_��
�CC=ۧ�ĸuݽ���cB>p��\k�3���]ϕ�W�F���@5�*��VMd�³.S�$ع��՗�ǰC��{���p#^�y��꽿|Wɍ���U.E
�#4D�#���8�l��^v3M%U�5t������J5�;�:JT͛SƒOB�a����4oS�#�|�;w�K;��C��l���]$�Ԥ�=RC�� �Ӫo�ф'�3�c���R`,��H���L8ž��.�muQ}1z D]�:�Ր���^����/���n׌F����~��K��e�?0�L��b���+/yt��7n�#�o�y�:	E �W�C%K�o!3i�NI�<3G�FUQM�Ƒ�gw�������=}F�����/�4����2^ho��>��b/ȶQ�Ɲf�<t���aP9�W�e��g�FR�v� !�y��cr�i8�s�����x�.�p��q�|�p��|Ie=I�ö���`.�3H��L����]� \|����Kޓ(���0
�2�+���K�o=���[�� �"z���-��|����N�tS��d=��y31�vk�����q����2T1a���� ���|��G��u�𢧓��L0�b�	H��d%���X}L}|�R�/6*#���/�i��	N!`������0��/��㑂�G���/;K2��H�I|J����j�Z���K�=VL�����=��J�@�|�߂��Pb�`ÓD��@`�JO�ËL�s=aVˆ�̎f7!�KTq���Lm�B��IP<{Q1�B�<3�{�l���C������!���%���<�M�}���by�y�J�7�%�|��U��6�	LZY�I��3?����	q@/����E�+���/AG��GC�u��hж<Pz��2��������w�Q��3�7h��&��G0fj����2Г๚��a�r���svƎ���8�bCU2`2�f�}��}S␚ԽP��D^ͥ؅Ȟ,��~�6�&<���<AO�6��#��Ķ�u2�
��=���b�<+�ʗ
Z��܎^kCد ��R>�u��ի!������/�P=q�cJ��H�S�0�l|��f�W��\�D�))���e�Ԥ���~��a9|�&U蕼�5m�ڪm���)|ٜ��b�.��0��:��%>El*Q��Ӈ�ͽɄީ�վ���r�h:9�̻���o�)�Y�+)O���0����y�������4��7�����v�k��տ�@���8u?��ŷ4�Ď(y0V`^�=u�j�5�I�i�u�GA��[p�
t���|���r���KixjqZ�^�qh.�7�?Up`Ͱ'6����M6��pI��2A���%��:�/ ⰻ�\x<�8
��@�Uģ
���M{r���w��8�GZ�Z6�Y�{:��&�zf�$�X+�=$�U�����֐1U���%_�=���k����Bh?-4�_I�[٣F��2�@�Z,ϟ����&B�J��l)��%򜤦pA<BԘ_E�m&52����� �e������lB.�m(���1riw%���mѵ�+Ea#�A�RE�'�,uu��U%���Nj�{�0���;B6I��#8^�Iu�45(o����V]�V�`��O{�@�"xm7*I��+���S�Q٢<a��Z[��"�V�E)�l8��&&��@.�ӫS3�88�Z���yn��τ�o�^�:��R�
Q��I��*�D��~�aL4uN-��z	���O��"7�N}#3�=ZUz<b��"�������b�ӯѪe]>�+��C���Vp(��vƒX*����GS0W�%�`�-&�QPEU��D�}��T^��Ea�`����d�����3'�1^��q�"�B�#��&�0-��XȰK�,�M�z�*�l��{:��(���c�^����c`D{ d#�A��rw*0��t&Fc$��r��^�{���=r��qEG>�*���U
A���+�X�#\�Ί���S�!s?�7�OZ�&���]�3c3��ҍB.>)��k� �j��l���O^|(�ǧ�r�C����oB��%��Fp����Z��{��U�L�>�~�se	W��'�1�M��=1����޺~sde�M��Mʢɳ���5?��X�W	�^������6~�u}�7��\H�ˏ7M�����e�5:�/X���d) �WL+�/�$p����e�I	5���'K�Z	��?���7K�I�����ȳ�{�?k�p�-����RU����>X->��r��.o�2�!�c��ٵC`�9���W}�3�C*7�3�xi�y�1��Ͽly�:��vq��]��_v)`�;���Ȟ)e\��3�9��ox�i�5���o��9��p�e��������ER���~`��g�L�9�0W��!���9��@����-�s�= ��t+�#����.��J���ӆ��n<`����oQĘ�~�v�1+�H�Uz�Z6`���'�O֧�`��l�x�#,�a �MP�a'���E���HE�,v��]ƺs���Cq��̜#�J�+1��Ģ,��N���O?��z��&ϓH�8 2rr��YQ�uq�YgD��B��C��_���V'R+��#1�48�
�˳_r���d^w9� bn�:��%Y�������xK���	Dܴ�w�@~>���;Z�kN�,m�,���f���j��'�M�z����X/R�`T"�@�e��~N(�h��p|]�Ԝ�)�W��� �=��l6����T��˛��ު+�le {P�A��p�&�t��ϚZ��mר*�e5����|&#�Bhj.k'�--��pn/�j�&���qiA^Z�h�GR����y(o�>�F1_>�i������+�d��z���h�����IM����B;�ƣEM]�f4=U�I���+�z�?==!�*��"��Za>lv��6�}�S�7�עMPS�����N���,~�N���G�P��w�'���ֶ�	�����c��ᴹ�d���a�F?��_%�B���h�I:aĀf>�7�&��ؕk�"<��P�P��r���)!���^��=m}XՏ���LįS��2���,�P����/�sm�b���?R۫��˟f����i�Q��t-5hKp���[�'����+Q�%�pD���&��n��_2��\]�"��a��13q��ArT�Ԓ�ῆ�E�:�d��bf�|�P���װ��m׹���� *�/>�A���щ0v�fj�ko�AQ�H!؄~o����$O,�N�k؆\�mTJ@�;u��?��/E�@�y�
�d�A�Ͱ�n�.m��`W�����z�noK�4	��th��� #������̖��E�u���»�c��&-!�p��U0����,x��N29!޻��7/����Zk#�C��n�'g�F��M���V�"o�����?>`��� `�~EQ���uMq��k�#eٵhC������V�������WY�h�C-�(��<��s9itq��>%�5���F$pո�9Y̗�NqM�3C�������Y7�&_1��~j ��(��{�h7��
�SOBr1w�L��@d����:�S4%���L
�d�w�b�߶8"���2�|�ǆr^B��K�NYc�F;j��\G�6}����Ir��(qL �z�����3�\��F���/A��2�`�Z����s�MrwD$�[��W�ax1�L�9p/�f,Ze�2DH�,��#ZZ�+g�0(¹�'/?����yt1TS��,R��sWs�	�4�瞬v���$�F�8dqT�������zf�(M/�g_�_4~��э�R�6�\���le��WB��_*w��~t�
����1��m����A1���|"���{����>8�`��+�7���%����&6�O���j��n&8�h���\��c�;=��Fg�0��{��%�m|F:�=����vWt�$��i�e�ۥ��I�^�K/Z��*�Zض������%��Y+�ߦWM����(>��U��� �]�B��w��E,h
~U�z7�S�7��mOQҋ87��s���>����T\��!P���f};��17ţ�������$ �}Wz(����c���I��!��b�U��g�S���<��E�V*��a��]9���*��������\hב�^g������|��;�:����V�����.��8gs�������˜ũN;��AF]r��,q���\xO������l^Ɠyo��+�X��?,���A����b�Mc��3?�Z����ؠ����
��.�\?��$�B�"�Û�����4A@���u��W2�h�j�a���֍@s�Ċ�63��l�����"��Q��<�:�.3�ʺ���XU��;��ӣ[tʌ����s�"l1?��Ca�?Cƙ��m
��W@i� ��XO{�B������j	J�ƄI.SCnş'�T��w ����
*,$���n�?VSm�����:���F���S��� ��峞9�b?���v�q��Oμ�����*�_��s�/� ��>	��=�&Ns��_�w��i@l��Ʌ|b[�)N�ͩ��:Z.v��"])�?�"fgo�Hv#�ho׃|&�n��"҇u \��6.���
��#��T���N�Y/9$�h��blY^t� w�2��@T����-C�_�%���|M'�F�����>T� .��K�n`��t�M�_��Q�K�{�:ȴ�0�v�ݥ�t�����	�f��M>7j����	��|�1��.��NO܅���	���X�;����Ņ�N�f?[��K�����e"Zo�(ڤ�q�un}��L�g�ɸ(T9�2J#S�]GN����'h�`���6�v5����'mu  9V��dm�~:Ř�Vt`�^+PH\J">��6g!�R���Yj���V���ơ!z��?����{��R��p�K{�!7�m(pO���យ&��`G�ZV�=����T挐Ou����䇢.���/,��5ol�㬮S�xĮѡ���ųxX�>�x������-oS\�#���,>�֛8[���������K4�.[k��1��k,0�cG:$��nz��!Kܘ;ӛ�4I�� q�én�0u��ِ��Db�	#>��DL��l�T�8�DJ��C/l��|�=C��d��x,/��i�}x�c���'/�o�wn����e��J:�{��b�жG��5��m#HN?�|��	�7-���@/{��sf��Z��l�Rw��c����R���� **<����KN�fs�H���gN�DH���Z�x:^��}I�Rݥ�olF2ޓ� ��G�9��0��W֣=���o,�� �#�y7�<�	#�6V_|C��O�Q�7Ŵ���F#{	��^�w�R��JZk�4q�k�����<[�>w�;n-G�`�͢�Z_����ji|��:���<`X�y�xH_*G݆���{̔���lQ[�i<ZH2 Q3�~�͹Ȭ
VP=�6ȽP�u7Ѫ~� .��6v�Ծ��Lu�޻�d��*����@��I[Xl\ C*r���Gה�E���s�]�/X>�l�
��?s澗9�=�m����;�T�Q�Y�b���f�#�e\xY�2�x�a@Ǡ�H-.�d�B z�h�@hX�����t�O���o�}[U�@���p�H}&�ڛ��p��F�NE� _�|������e�Xo�l��f��v" � Ja��5��Yu��]�������3���KA�F��R ��q������w!K����]�	,�(�$/� �����n���&�\\M�њ�n�ǧ�
'���~����H�V���t6!=�NDK�\B�0^���n�;L��ǩ�(N�܇=HI�3��9��ܱ�?��v&K�Uj� (T*OgM5�@0��HU����b�z�B-��w��;cî��4L���F��^̉�^�`h��`"��~r�{�m��+�m�%�L���USI���Q
����n����9��[�C�CJ�ܗ�Ԅq���eޏS:R����hH������q#�o�����;�xo����4�u����z&��r�u"��oM�g��]D�>��H��-=�L����kq
)��M���U�Y�u�&�.��$�=��?�
�
���l}Y�Nw�΢�M� ���ܲ��r��ݐ�����];?t�q�����D�Q��_��sp��Ӫ{������ �a�xw������\�*�f��V���>�c��U�p]�!�pH�
`�B1�>(�iq��.��R�#����9��z9�GmA/�AͬT������_�6���N.�n3y B~�-֫l�����΋s����^�H��7Z+��&�M�u��Y��!ƣ��v}���̑���󩰃[.2�N���y/R���7aTk����
�UDdg��,K3'˕[*�XklVU#9,6	9��M�[Hs�0C�+q��Nld9�A���J4m��e<�Lr #�RB���i�|Mƕ�_����i����`��'�I�PUɕ ��%���GMs�,��йL�KX�C�A�_��cY�I]�w�.���òp�m�i3����]WLS�*8βSӪ�öaȣ�|w�@*��M2�g)�Z�+'@�a�϶�Ji��)Fk���re+�l5#^��Tdo��
e�N��>��c�MyK|hk��}�ɮ�3�bĜվ�F;�A��*�X�3�ֈi~{%l��AhD϶�޻�����f���yX��1�&�[���)�����:̝Y���	� �ˑ)��N��g�76��,�K�2�h���5�(���b�NT՝Tڣ�����e�{�RT��گx�����F���f�U�����\,�mN8�h���(Q�IA9��ۊ�)�����li˛�͆�2,!�K�@�x�K�`s��K��S' +X;�_��oU����T��Č��3�)��@��x}�Z�d-�������͸61KFM���tp����;Û�}�X���+46A�<s�`-C�o9{g�j�/�˖K����X���p�@c[*������%a�lf���m+%��Z@��\d��f�c�7��9��,!胬� {wr�Y�a�F�]7靰B	Р%����e�_ŵ�`Sk[�A-!�%�Yp��<�%�bϝ�V�H~���Ay������Q�-XUٹ(�LaK�%�Ϙ�9P�N���D"����ha䙽�������9�1�Z��@��Ǒ8��C�|�����,��xr �l:�3\,kE��ߌ�7�рO��6!V��Uo/$���\�(	���I��B�y�ע�����>u�	D��K,F���c��^c�%;��x��r�16�2�-�=���ÞQ��CC�٨���ҋ>�k/+�k�$k{���[M��((�߀���8��S=Af��#�"�I�혍�G}u�θ!I��5�d��sy?n�� ��[$���Dƙn�s�׵)��:vF� ��6�~ߺq'bF���4�o�f-�iY�~Ut:@d˄lq��E�������ȗmfb�ւ`K��N�j��D���ZH/Հ�x<׮�f��p�]�xB���4Jځ�4q�\ֿ�͙�]��a����H�{��Ă��(K"aof�a��	���{�G�,�
�Kn��_�z�>j��^��\7�x6�LL��#����L w*bU�#{��A���3�{Ucx�����Ruj�"O�ٍ�ڳ[�
��b}.[:�E$!�ڢV�:#ۨv�����DA;�h�>7���e��8���^z����_� ��.41�0;�d�H{Mz*D��»����Sy�?;��!CDC�sC6@��G���n�9��}�w��ϻ�lxB��ڏ�?W���e�V���4���t�D����.��N���Sfֽ�V�2"N�x���5��mBo5Z"*]Sf�"��7M�cm�k�q{x�i�wx�OO[���V�O)�,�g�>���0
���Յ�����Z�
����V��*f�8�'Տ��P�����V����.�n��ζi�mZ�h[ĭ�#��������^j&yލ��0�� �C��n�k�v<J��rJ���C��:�X~IB�g|�����Iq�x�B*�>ed��#�x��ތ� ��!����^�����r�u�3Z��%[α�J�-&$t�ߗ���蛴*�E����FNZ7I���==�@ҷ60�ua����1��!� �n')�`�$c0ۓ�����w�b���n�/Zk��IV��^@��j��c3a��`�����zt~0�s)�BO��͹�#�ϰ(����"<����*�sI���X������ �T��Q�a�3�ǐ_�%ۢ���� W4Xg������,Ӹl��H'������2L�Ƃ*�"�@�G�qc�l��ް(��ф�ZقI�+�}/_�f����f���r���������*���_A
�?�j�@��R�:�~v�X�`=�x�+<�1�,p����l�ǥng��L'�c,u.�'�����W,'ľ��U��j�YI��^t�L��̜�>R��9 �����f��%0���lM�.���Ei���g�ml6^pF�	�H82���X��Qv�p'�)�'��eM�>� ��ï������vN�E�4�� 5Q�����]��c咬�	-��e�D:�����&j�U�N�֚]E�m��*�^��ʷ�{aߚ��p)�
I�p�y�a�1CQ\r���X�bٓP��(�g_T�Q��	��<�/�Δ���*�K�r'8������+C��]2��M����R������v�,c�t�m$��,�ɵ@���Xr5��~��N^�%��SƘ*m��	�;r`s�x��󒞴�i��:0��'⏚a|��.���3�81n[��3rJ5z>�G��)�S1_��Kَ����h��B��'�a�(��rh ���{�ܘባ��yϯ�i�;�uuh>�ti��M�w�����P)g�e{ ������E�k]H�]�H�D��K�!u;��W�]w���D��eyX_�ը�c�)Ā���1�X`���$B��wަ�~����FGV�&`x_�O�A���ύ�sȻ�oƏ j��fMߜ�Yu�W��2�B�E��	�>�?b�Zw��
3Ñ}Xa="����3�m}7ί���{�%B�'0���}�,�:�Ph?b�1i��c=���HY=$/����:���.<�͌zf�uS+��*�ܸŬ�7��aOpCo�S&��QT.H���)�ox8��O�0%�C�H�[7-�*���)�`xO��� ���}߿����@�:Vd�jR����VqH�l�ۜ�y3S�I�(W�"�b��@�ٕ��v�Ld;�]��V�e�<��):���8G�6�P��������9��!��o�O�A\A+^!����J
*�����vcߕ��vI�'2@����_K�YBy�Q$���\��H�mP�Y,��������&WS���F�Ï��		���K��;;͖�� ����J�^�������s�s
sA�vE*���'m�VEI��)5¡&I@������4E����)�N֓��(B��w4g0=fΈ�8."�g����Q����d���F�������"��~b=�R�Ҕ�仪&I~��M��~j����d�����=o��p�M%�]�E�ػ۴{���e�t]���Jl��1�b�+�x&��nӒ�^Mv�|q`�8�zRo'$��ڀ#�J���T�C���.�4��#c�"�_�y������u`.�EJ�����VLM;�Z��n��B�����S��kg�sy���M�??��£�1.�Mq9r��F�M�Ld�bd�C�H��&���N��q��qh�C�\{��qF�RF�����@�"�bڑ-ݗS{:*o�K��!�2	c�L�������C�v
����\��)���F?m���D�Q�[?��%zv���WK�H�(���@l^�n	@��:b�9�j�)�ki���i�<*�{�\B��+�q0��gM��EV��eH�|��ͪ�̯���S�e�:�+y%<F[�VH�;�ؤ�x5��J�i�M�ޜ�>6Uz֚~
K�U�f�`;@����zu]
�
��BŮ�r�}��xϐ)����τ���tecFĆή��~ط���$`v��=��/QA��z��Y��{'���'&xv��s|H�OT�m?M'i�L���p%!35��������<l��?����]��H1�#x�����i@��جD��FX=R"�}�p�\6��u��ed+4���0uls��b��H��3�ih|->��`6�W���b�T�F��cQ����B����y���Rm	D��uCB=2�a�# ��8�����~ʬ�mM����^�lI���J ����Ƹ���$U�R_�:h�%^�߽<�˅kڕ���a�%(:����N=��|>���0�����v"_$�P}��%`�Zg��pL������.jrdk&�_[����( �)P[�!`�2EȕZ��Ф��(���1G��8���Ș��*6�W�˫����uN�9-H����C͋Tt����� 3sY��ד�T�B��)6,~Tl��w'�s���d'S{����j ���#i9TQ�.��h�|2�z�'����q���I�;@yt@�a��B������9H00�$A�����9}d��)=�^�62�D���������MBH�Z�i�T�}4}�ΐ�e�`�*���&�GX�)k]^Ě�P*5�>��	 ����3�t^U��qFA�݇��aѣ�r�%�w/���8fx[٪��g�`q�i��13h�BFI(��s�i��ib�
f���2o��5��Gpa�5��G-	�x�
f{ܵ�)m� @~ �RT��:���\���|㎊ꊭd���"�۶®ڿ*�f��*z��+ŋ�N���H�q7ސ����q�뇑�?/s��*V@�.w���Հ�Z�?{���76��E�:@��4-��x�jZH�<<��K�%s�ZӃ��r��J/knR}����*!"6��8�) �����v&j������"��T����zF��#o O&9:��vX_�L=��iYe��H�n�.������I-\�|�5.��=�ۖ�|?�$p8�a�%\��i������*BZ ~�e���e�F=�U��x�n�^Ç�ȱf�$oB�N�@H3�O��h�;��9���U��,_GFq}#��&������Dp~����p��� 
/Zr�x�	���9��'x�T�WslS�;'P$����2���X[T뙱B��}_ ���t���c�}�Ú���ed*�H+�m��ޘ��r����]錤����,^?��x�y��I@��^�Zݡ�x-�Ǵ�Z @��TrN�O�gA♜��U�S�tW��rI� 
�D��>�M�w�no���R�,d�p̒�T���/���cQ�֋�Դ��[�-����E�BY��!�4+���O����z
?HXE�����A+���w�M��dD��=�ފ�a�7��(�� ���U�Y
����-槲4le�2�OR�J�`c~,ic�y��Xp��R����F$w�k���y��@�Sˉ�"���b4
tj}�"���QX����#h���`����KK����>y��r�?Gx�{����C��P뇳f���b�=k��07J�����UA�n�=��6�ݭ��	��'����6x"�P��2���� �]`-�7��
'��{{mK_d�p��;c���$<;���tp�l�$��z����H﹇\dђh����"�'�������
�MG}��nn�떦#J�OR�m�84IJU�xѭ�4�	Kd��)H�	*���䧇�/s��6.���k,~�6�=��Kz���S��Sڕ�xx��N.�Cu�(�8z�G����̙Y/c��`�14}��n�����ԣ|/'�� ��{��f����M��Vr!��	OgT��b���:��>�T� ��~�SF�U�Y)�uc<�A�����=�C���&�;�[ƹ��)E]��{QC����bn���o��
������*��C���:�ig#�m���:��e�����.�]Ґ��$YEܔd��~�"2��U�&2|�+�3��"��_���5j���r���Tښ8B�^�����bѠh����D5�%�%ߛ������"j�}��%2�.�u(B�֫TM
����Xy�kKh���ݟ+t�Z��6D�qY��/�?Վ-���z�:�G�k���T�%��!p{�Jx��L�H�����`G�V8#�
�,$��������T��|AԾ?�`���z��7p�����+[v��J�J@�;
,����,m޲C)?�g<�)4����w�-7��e��c�T\,�̍i�Js�w� A��Ec�_G�Hz2��3��q䮡��P Ì�(�X|����7g��h��X6�V�WM��Ϳ���PBC(�Y��Zs�EFz'8"1p����>̈́����[�}2%�=~Do�T�|u�X%1���2�>�mX�F҉umS'�����+6{z%X���F���
[�Y�DE`�a���Iv��`�t�4~�V.=W�9�P9tfE�*Xd���щS�SZז<�`�d����*z/S]b���}Th4����<;��'�pO�+܌|١�3���i'D#C�G�`r�RnI�CL���1�R���H�D��y���Fntw^����7��W�r�(��m�/�2Z.�p	:�4���Z�i8�Y�S8�d�E���<�0lAl�a��P5�9��^|�/��bdԵ��;�ci\�ZJS-	paygZcݍ�&a���/U��mc��3|^-N�`q��g��`�0�+�2Y͸�٥����c_����j�U�j�FA&�>"�a�q�[�t����@AH�Pa�� FH�U&G�{[K\�jc��9�O�X���j���@'�B'��Of�֫��Anb�/k�
�;,D�6��e��!vR����f�_���� EA
9�l��/(դ#�vQ���5N�{�lqK� �|`fA�Ϊmüv��2��ow.��g��h)���t
���ܐ���)��Z
��S��l��1K������0�f��&6���O��O�~�f#;z:(�!N��*��{N	�����fX7�b�@��>�E����GX�CC��g�>��k��JXgiֵz�c��SL΄1
�n�?�a.�g;��=�?X}�!$/D-?6����+��^0�v)Wkzs�8`ؒ9�֯�F�3)��*�`�oM_���S���i*���ͬ�Rh� ͢^�ff6� �.�����å��6��M�^Q��f��z%C0�[�������
��A���[�����l���;6�r��{ڶ�6��=�j�1��f`;StrJ�[H�����kK���(!0n\�ޗ�!}�It�Hs���8;�R����#E ��u�L�)2�ŘN��_ʙ:p�!�9wÜ*�z|R����D(2�p�PYB����S�4,�dllZ�-"sGg�ϳ���1[F-��%2����z�m����8�.���ʄ+�"E�k��:�M]�|�uʷ8~]���*5{��Ό��a^C�B4��H�{�;(YC�������2{]o�5��r���~l2Ŵ�Gy@��u�v�QUE���M�<�z5[\�t��}����W��5�_���bƏ3��?�݂��-(��'%`S^8
��F����LŒ�ܒ��������.���� �@�����v=����Oi�)��$")	��2Qޕַ�=z ����C%20r1��Z�ݰ�V�)�P����`3��4����Zhƈy�QS��ȩ
��)>�� P��ir����u�b$�J�g�3I�wx̃r>��/L�Db�CNM}��i��5�m�z���B��2��z���f,��������?�YZj++���p
����M�?�D&Z+���
5'�ۖ�H��i�g�°(�R�Q�@�R5��up��Vıs�I�o��;\�oH�k�=HueQt(Q"�Ȇ�Ʈ*U.9ָ��,�0P�ٳ�>�fCk'��6X��~�&���t*J��R��I�02��v�Qu�ǶY����|:��L��q�|���Y�ǁ�J��Z�,^V_�����Ҧ�B��j�JD�l�B����.���>�ȣ-l�@�Sxo@�w�<�v����N?���|��a���4���*���!}P���p�<q�p����&;ң�,�#.%�|c�p�>���8��Ev5��̵wH�|�SȳI9�W�z��A{)��h�F���Q����v�,���6���<����q'�>kF�>f�����yfod������c�������*j����	h�͌�;8��T	�u˖ �_��Ҥn�z�o�[����4�G� �J���<��6���D��+A���I���]��˩Pv��.�:�Xz���C�;��ph�|OP�]�
e���5G�U��&�_�*Z�\)��`6��x���0�"���+w��ێ����M��3�����ͬfN4�f�w(�:Nl�w0 ��(��̆s���8�B))��g�I{�a�n��u1f&2j@Ms�͘��2����ѻ3g���� ��~{b �<[܀(>J�6�;�c�`�Y�Kr�xj>K�(p��֝�t't2v	��*�嫮�U�
Ԇ*T{�U)� d5��qͧ?���a�d
|�Vkc{��|��T���_�P��u���/�%]��G�G,�ɰZ�u}i�2(9B�_�����gCf�R� ��������:S��!�t��6���7��P�"@�!��k�C���=G��k�9F�5@4�!T7/��X��`w�����c+F15�ÇG�)��]J��SG�i7�ĴH27b�?v���`1�Xɽ��B���q	�D5����|��q�}��)�y�4,�p�� �}�Fy5��T���@i�R>�Q��4L9"��Ū֨�K���O'���,���0����{9��*1��d*@�����|������_���<1�C���~u������)B]����������QLe�%�>�r*�n���-��|�(?�A���-u�O݂fW#� KP��g�";�utn*j<����X|@6��@�H��2���j�bi��,�D�.{[��F�<ܰ�<\�Yw<]�"[��{0����}mt␢N��DX����Ð��u�"�7L����E�Xz�u(/h�QJ�3	�?�������A��Ԉ�/���N~��"y]/�/��F�,Bx��}�ˢ��P6�O��],�X(����н$w�BY��C�x�������ͫ�R�ب�1��&�Q'�g>2��(y��{��Q�<癟LEpy�P�`(�k�T%R;$�C<+�ᗮ��Q�`�P�[`9�q4�;N}O.�K�_F�²|��<IT����� }t��,����}�F�ZifA�̘�X�T��$N�6`��[�S�b��Q��N+f�2�+����-������%md�_뤌�I����� ��G]j�P�},����.�ߑ��t�~
�K�gLPU���c�7�t���8��ٮ�C�n���:䴮�k��%O]��F��	�"�2���'�"�k�	����\�H���n�4�j8~��<'��w+�HkCt�_b�OE�B"���_t����QFi�;~̍�>\�}U���Y��&MAx皋� ��j���pu��lxvl`���,��2��,�?�ֹ�3�lN���g�/��U9|��������*'�m�t؆.2����v4ij�x��'�a�%]A�j�L^�=8G���ļ��P:T���%�e��A��&ċY��O8�s�$�����0�oҟrKD�:4\�\u���I���X{�G�d=l3x��M\�)�,�q{euz��y;�
d�H	M�"�%Q4��a^���r�N#ּ�(^!ݢ��2�}�מ�	�|���.�	�꽴��令�'8�WR�UyS�b�9��p�
�(��52|┌��^k��Q��L&1{�t�K+6�O�CL�:'��|N�5�h��B)����Q9��d��j?y�L�buE0���		5@��<�f@��7rW#D��셊�s����X�6?A�w_4jh�-��THGzZv��ᶄ������J� �GB�g��g�lbx������=���V�J�Ϊ9}�q�Uo�FEO�+�9��v2�kKݪ��L�\_�Ul숻��t��7�3W��̧�GBT�\z]Bn�>Ҷ@��3�;m\�����'s�N�%F��~�5���~�#�:�\��NW�q��Y4������=�!8vrxp?e�}��V�C�+�4(p�q�6����!��Y�WA��/7N��0�u�l�>�U-|v�ց�O��l�M#g�|lcA:��{�O�����z�N��N)`���@ů矹�wo���z:���>D�9q�w��,��>����=��o� �vD�g��� s�y�5�@L���0�=�m���F�|��"&����s,1�[D[�.���!۳��x�,N8$���M����5;Q�&�PP �^S#.�4�����^�Rr^�W?��4��xo�_l3�6�M�1���D.f�?��&[6�H���&L�M�����%���5� �g��x�v�����fh�H�ftb׎I�S���ͣ��E@��9�ۭ��d� 6�bZEq<g+d�D!z��������	gY��e���I�_����$��'yBT�`X�8 
��مm���Ҟ��Jyn��}|�y�]$�ux��%|L�pF��Ap�����Q�ḱ!a�K�8Ndu��⚥@�����vE� ��E�Dr��aL��,�����M.������+ȏ�N[DbGX��UD�,@꼹W������"��K]t#�K"H���fG��.3�r^��x�I���o"���@����>Ð��`��wLW�tmJ^_�Pe+�>�p�3�C��y6�\��L��[���o�ޓ�c�[�ެ�%q,O�:1����(t�d�訋s���o��}i�;��Q��2Q�d6@��ZUĴ�)
9Ы��%���&������g��y%5)��Pj".C��Q�j��J:��ylU��&�Py+�����U��=���3b1P�<��ᕂ��[ri�d�cVM���OT�uu��c$�bH���V���z�vNVۡ�/̚��e�"W6�Hx��/S�ן���
�e��ޣ|p�,'1�<�����R�v�R�-�Ӓ�d��jh$�FXw��M9�e9�h�0^�k	_��ߺ:ѬR��U�Y�\�Ν]�2F,v��8����8O�쑋os��B,���Xы�.%U�le#`�NC�'��3��p8h��M� ��Z�u��Ύ��t#|�_��S5�nj�י	qRl�(,`�n�Y���ϩ8��C<~(�ѮZ��R��ml�c����� �Q�*�O��}�]���m��x\�T�"���NqL?��Ʒ��LP��!»����~g8/~�r� Z�V,���F��2?�����p���\�_0ʁ�Sy�#��
ɊG�����e����tB��~���r=�n�����;����dF�d��=� p;�c͉P<N��t�l)0�y�r���\�*���R;"�J-���&1^�V�ޕ0��gi����R��Ǯn)!�1��e� i�qW�ن7�����"󟣂��2��~de�2Ч�|��&�Uu�C�YO]`|@�Sр�����?[u'���xI�ê��4�c�_�Na'�f�xR�}��6�1�71�%�$Q<|ެ�4tO�	0���/����C̞r�5 �s�N��>	�����%z����UH,��F��w������bF
��x���R�,��׊��p� ��tv�xE�rz^^[�d�xPS�GK�uY O� �}]޲{�w~ؾ����ra�ch����Y.�lev�1cg����v���IΫ(��\@
΍�t�Z�>�c�q��s�蝌<�;Q���Y��$x2��B�����.T8ML�y���-:��;6���΀�8�wq���p�3�b$P���"�ɢ�p��o��v���7r�i�f�d�F<��I ��rӅr3g��H8�?<��
ūJ#���Oֵ{l�u��ڇ�l~��$��o9�]��Q�HY���n��RyC^GcDǟ��]�ɂfNz��*�8�����UH ��Ρ��$�ݲZz�o.
�u`Zj�ϡ�k?�n�2�0dV�����ʊͭ핥��c���̩�/MSȶ��&Ã������ }�Q�`�x`K�@uﮮJ
$l��b�#��-���ٿE���ߥ:&�_A5FPW�o��[}T�x[ih�@�8�	t���0�	�,8$MhlP���ƭ��B�GK0�#� _�wW�}[z�g�38_��Bk��cC֍���Euׂ�M��1�8j
W�~|v��vƞf��Ӗԭ��r��ݕ�*����&��At���9�Q:t�c�&��a$�I�K�UO���|�w�պ!���RB�`��aݱv�IQQ�x�3�:�8Ei�*-�@ד�N_�ו4�x`��P�QB.9�����R���p���s-�Ӭ�t E�1��Q�&s�s[��Y�k��>��H�����	�U���O���)"�n��Ob+U�rӲ�d��2k0j�v�w�-�W>a�|���}����F�D圼��G
���3���FRiB�~����w+u8�F[2ڇ�,��z"D�/�g�}���`�Ř.��/+.W�-	g]��sI\�>�)�A!/OM��X��᧻�n�hPև"��;UL��� ���CV�):����`I+s�,�}�(�z�����>l"�UL!hC`��r���i���&&���@t"�J0k�aAߖ8�>�O֖x�c����?�?���(�C4��,1�|(;P�B&%�Œ:vS��":�v�wɺ��@�"�`z�$iĜ3�E��p�g�m:u>�C.�cjG�@p�{-ʥ�RUEZ�F>�����y.{���}ܶ�iy-���J	N�(��7]]���#�AV�Fv�a�����GE$BE���C�gg?��X�K-��?N�(c�.7����g�hf��m�[R� �H$�'�>;+ڸ�7��)���,�Ӳ�Kl���|��]};2\u�<���g<V�K1��E��������숃�,�V���� ����i����x�E�Kzw֊��U�2ē��˅��қ�RS����j��b��[X�CC�-C�kY��}9���@�10�Y��0�M-�Ix�#��w�����fE臸[5>~��Ϯp|�QN^�[2�<檧T0z�/�'�!�]���\|.-�?$0�������/n�`]-\�ND�[:{n�� Ȝi&���%�q'���\�5ӊ�*f�M;���УN�39ѽؘ�1�x4f��2,-�Bo�����v�λ���/������D���P�cn>}�)���Y���~	�/�P�sc�k��v`�\_�p�3�vp췊;=�qy�S�����ӥ�d~���� ��F[�۪DE���llO�����E3�������7sL�Xc^�y�Nn܉*?u:/�6Vx��O���̓4�k�P�5w��DēOp鹀٫���*A$�O��'��Ȇ8��o�,යE�����cӏ+��WpT l��Bڬ�<��n��W����A��������Ht�#�I֦Pj�X���)M2��� ��(hr�0�V�g��y��}9�����
3u����S����Q<x��ſ�D@c�y�$T�>Sǿd� hIN[�����>�S���<'�o4��Z�Ld	��Z
�`��b�H���c���/�Z���8It�%i��}���Vh��v�a.ގ����ּ]e�� ����2���ۑ��[���Ċ���S��$t��B@T��Xm_��nK����אߨ�{�
@n�����6�[4+���O�`�3��z�y��	�j�����c�&��2s
μ�0���'�w1=����mux�G���w�Y�g}6r!7ν?*@�DEfE�~m�@iV������ZH��,X���	�����S� �ڰ�a�Ǚ�R�a�EJ�f�M�>]=���Y��YT��ds�G�_txȥ�M�f=������]�g�e[{�Femh��u���߮y;D���SDxЛ����x��n�L������&��KDJW��W�@ͤ&�-F"�����j��1Gi��Ϻ�����N�M4�������1oؿ?F\o�i�@!��vn���� >�{H������ �j�7S�+T�`sM9^��JRj�3������B���M+^����^oQ�ǂ�F��se��Ih6�YP`�i�hݪ�Ol9�m�q�^����2��/\1�Ӏd�$3������߁�X��";�,�6[��7��u����Ԃ	y��($e3h����N��H`A����vW0W��7�鎒ڮ�U����χ�N�Η�Q���bzՋ�wq�F+(��L�H�g&��'��^�vf���Ȳ��������Z�R��;<���#if��pgG�4��4t[ޤ�k�IY�AO!�]4=�r�'�Z���0Fi���n��VR�}W�!V�Ҍ�׮|B>>�O�����-���^*��wa��K��|�{����S�t����z3CЇ3B����T~Xf������V]��H�^2h���,��z�0;�TB���h">����^�(U�LB04�yL����������A��C�. [�����r;WR���))�&���Gf��2Mz-h=�XH�+^�� 7�̝Q �#��G?��j�f�%X\��}(Sȸ�D�?,�>w��X
dp�)��Z�p��x6��0��k�9���Y�3:ri��35@$t��m���x�f�g�7��:uK�g
$�����u�H�GD�S1�ݢ���	��n=%�W8_�Rp�-~i�������O�O��]�D�rbs���E��C��(��,v�#&{��\�A���XS��)Wdh�ĉn��\f@��H���5�}��|��E��.�!���&�+�V�N��m��P����=XK��T ,�롚�&�q�V��z���H�[��<qGy�H�3V�� ̐���!����M��֕���]��gjY��lp��%�����"i��4�]�za��q������6˽���t�[j�v�J�ZR�ՙ��ݳ��vk���kż)���6!^�� ��Nc��T�E��R�n��ݓ7�U�
�����b�}D/�mR*���T�V��ƒCH�"H�_+��(o)�cC/���Τ������)�v'����F}��3�FH��� u>����rq���i�f2��!���l}�_l�^"jYKr����NC\{�8|�������b��ZC��_H[��<�L�7�^f�4�'�{��9��Ͻ��F 5��I�pV� &�'k6u��"��Y�c�ī��Y��.�����㲗�!?Fc� x�����m{C��}���O����
�UY
�a
L>�>)��fw������4�����l��;��"���%4qx���Ϲ��dL�	3�	s،�~q�i���QO�?xT7��}�T�:黍��Nҳft�W�D�-����(|���֎τ��_���3$bk�������������/���l�F#��Hk�i����@E�s8����\���]��_��h�<��i,�&y��g u;΋/@l=�k�m&z��8#������=.B��|��Zኑ�C�`})Q�-du8�U'A��1?z�*MZI��c��Ps�|u�4������N�����#�/���wq?�7�-X?DEy���\��T�Z/J�����n���N�%h?	��W�{l;��G��B�:�<��BB \�������?z� s�&�
���m��!��F�"����u����x�h���ҷFRJ}���0~#_�Wf�j�W#3�_٫OWUJ�5a����6�BR��C��0�_-�����/�����u������G�z������)�T�
ο��`kD�k;}��W6!Tx9�3��e\#띜��������I��0���?�x�B!��\;��{\߭W��Sg���\L=�Tqqի�z�2�����м��y&��d�2�o'!�"�����O�8����½ĝѻ���/�s�j�N�#��_@�;��9C���U�����^���Ċ�J��˩V�G�Q;���-�/�+��]���P��ԓ*�aZ�"	s�orx��e���)�nK���i[�ĀI�s�(��/ӱE ���(-7�6�_����wGm����r�0�� [ �mx}&�u�A��pJ���U��U%[��ܔ��v���ٖxڊ02�H>JK×fA,Q��X������y�����*�5�zK�4p96�Y~��=����"�	Y�D)�n�)`{��m�*p�eKU����[��z��^�fѵ�y�� �qkx{Gֵ�3z�y��p� :z���U1����yp�	�X�a���`2�9{�p�C-'H�Q��<ɶf�G��4͎�8@�t";9CE���-���/�͓���;�)dĽ�����X$y+=q����k�Ǚ\��۾4GA��O��%9����LKH˶,X�^�ӷp'�s)]���$=yHH��Ɋ������F#i�8LR���V�L>"Q�����h7���of��&��?�>$�!�Kۭ.=FCn��Ot
�C9���^?�%���49�5�ߊƀ��wӐ��/@�h�l��d[�4��7�ā��oǢw_%-?M�9W`���~�vշ>f���!>p�	c��E���p�ᠯ�=��owV@��4X���+��m���T�B��3�.B��@�4#�;��,k��T���������(�GȜ㻅��l���p�	��l�NE`#
���9�V�R���HI�Ih�hV��+kR&^�1ԅ��X��pg�b�%���)�����wK�H`�!��۸�ӫ�R����;��H�̨g<Og���Jҗ����Ⱦ�	����o���h!]�(�y����6/>G7����k!P=���X���_�X�mM&�1}��U�w.��~X�|H�6Y�1ޢ/qx�}z�a�~�����Y�H$��Pd#�q?L�ۖ���UcL��oӺ��ܒл4�X�Rw��A�]���J�ş\��j����j��>���Ų��hS|�zXnˣ�ƀ���w?/��#�q1��6w+�N�#�X�g](j\���]x	��G�r�Y*��J�YX���7$�а�9���!gf��.H��L
Vy���&<�@;~�f w%��n�/"�'4���ڂ�R�2$o����8����[��Vo��r��X�`�F!�G�^Vq �J@��Ξ�M� ���3wl�,M%b�])3��R�^���IG��κ�� �.潢��T�J��+�R�F&*f��A�(n��DUXR�[@�������PƄ�d윸[��s��Q�(QO��i�y����y�PLH���*���.~��}c��Z��fn2��}���eU�na�3}Pw\���J��;8
5-������,-Ŏ����=��'J�[9��xX�V�gn_�-b��x��$��,���j$�Z���ά����4\`�o>�4�N��1�����X9�����|V�B��ח����WE�{��W�uZQM����ls�Mr�˱4��mD��SE\�I<|��27����?����
P}�s"�Mhu������HL�����檬Mp'��01'�Ssg�v�c��Y]6 �����;A�t��j�z%�$N6
�
$��Te25�k�7ƞ��/p�d�=n*B4�7థ�����-�Dg��:H\�����L�@	�����J�޶(�a�������HT�Y�ԛ����S%���h�n?H�p^i1���aha]�����rI+ķ��T�@���x�W��ʖ�v5�^����KHn	w�6y8a��x�F�L9;�l}�f��z�̯$�(j�ou�M���_+݀��b�~Ц��N]�:�n�)��o�"����Fj��Cy�\A�y��ph}��2a�n��`B,���kQ�}X�+��"[9�7�!�=������7��$�G��{������aF!��.f����0��/<�vG���e
����dDI���G6�r^פ^1;F8��<�k�%{�|�D����C�q���Q��T?AhU��:���ā�ʹĽ.�RȎL����2 l��ի�������Q2���M���~�^|q�
���iRޑW6�>|�h5/�J:����lwd�R��Y�2�=���{�wL��c�MCzwe��h��WI���%?߇V]����x,�Ku�Bmv��$ov�V�%������8�*_�sZ�ׄ%-��X�{H�axmF1���}����$���ޝގ5ϩvk)���^���(>�0R���.B\,x�P�`,0��
-8�9��<�!�d�����F���y%�L�Rz���X&6L��O���9����ͷ��&3IV��\� !�O�Y4]���C{Yb��ojT�%�yx���Ɖ.V;D@�L,0&j�H�Vp�߼�%+&�q�����Z������3c�A��+@�%�-)UJ��T�G=8�������jn�*}�t �3P�wn�	T`���v�X�D�������2~��_��BiPU�X<�)�or.�w� �:a���u�{� 3���*T�ů�X��}�jr����T*y�|k���c$�hp�~s�#[�ؒȇ۳�-�><��M �D=�pɀm{\�u��.y�����#�P��ϣ��Ui�)���������K͝��]�[8o�]#��RH*L�N�%���D
(v��[g+���כ;�΅�e��1�%�n���]��,�]%f�pY�{�&�7:j"��~�U��{Ȧv1)����׭����NŰ�2��&&f�s�9+���u��\�#�ؐɗ`�Ys���F��I�4�%�����z2�`�M�K��ʢ�SCp���'A!�3���877o1,}���*�`�pP�.��臾���߂���o�
�A����Ǧ	���C0f��'Jѻ�ڐ{B�c�d����b���~�,�ݍ��U�Q�B��YB�rw��*����ÜD�
�^}���/�BK�õ3�#�X����p�S�l�1�2m��=ޝ:v��睼�N�^=��'���:�������|�t7��JJ��LG�`r֯�bӞ-�'����J��1=�$b�Ή��ņC�����7z(�����}����;��U���P��"�	m�#���`4����d��z�Y�Xt����;��6���W~­��1d��·�� ���\��4�� O%P#�x+�+{ů�ړb�
��|D�JVF*o�g�q�E��耋�=�|G,d���VB�Or�@���2�	���v{��;�>	[�dZ�?|[�vWqR��yl��)��,����엌Z�>C�2�g��6��m8Lk 0=^��C�|���n0uI a��9.�'a`�OԾ�֧Lb�s �2���,�[+��8��s��kа�x��n>�Ćv�苼5mNR�맾��b�}y.����3��c;�lZ��z�n�.��:f	�R�n�����PQe�
���n8�C��D~Z�h�cх�ח���]	�f�J�?�E���ը%�JB��J2�[�/a�k�Dn��x���L������G렒�V�&�ﬨ��F�@D�����g�O�G�!����
��;�)�7��p�MN$]�l�p����A��6��*'+G�K�A�:��U��ě�M��(MhF�ӛ>���h2k5PH#pQ�Ll!��dȬ ���^J͛�����S���Ik߭M��mRW��5�|'fb������86��T�l��:,��аCx2۸1$5�_ވk#1��4���F��c�̔Z�c����>e:�]MUy���L��H�:� ��qO��ᶜ	��4%���j\���ISjHS�F�KZ�����_D�=���,�G�0>� >Ȇ�t�U�U���O�Fv�K��,�PZ��_���M �n�� }0�~��< e�
88�I\�<D`�Y�	qu��s��f�ݾ$Q�g�}�=�g��_/��ľ�`U��'���}ȇ8D��A���`�`�2�G�� ��}�f�&���1ZRx�֢�d,���[�>������@'���Ne$���QG$�����7�4м=���N�n ���q'�sƴ��a'&u����q���c�T'�_��w{���sv�;��:u����R90fT�&!�8��P����?_��S�!� ���ڍ
��ul���OF�>�&/_���[]��2,�}������O�2ת�T�Y�������*��W��oϣ�ޘ�	�Ժ���[L��u�p�ƌX�t?<⣡ |/m�8�A���2@d�����������+(����ݾ�2,m���a�ׯ����7@��	�2��m������^I�$F��L���YYw���F��f;C�jA�!bu:>^j#	TF�+A�������I�Qfp!Ƒ�!#ڤ���Vv���}��r��מ� ������{��&j:��O�]~�J��E�M�X�P�(Um���*�:p�{ۺ�X���5� ��bGw���4`_<��b:���P�.@��*�lp���:CF��� (��ZΒ�9�K�V�X�]���"�?�W
hy�b�]�t�� ��Y�y��^��
�<G�s1ԩ0����ͤ��tWB��||Iq�$��\�_zY�7���`����A3G�P�S[k�<;7����&��۬�tҨ3�q8�!�s=���8
%��ߘG����\���3J�$�/*fSH8EG+?��  �KZ��)�xmE�V ��@k�>���]JV�#|���X�HO����ŵ�_^���>�{bg����!$r�:�J"�A�t�?�����Qq"�7��b��z���=����l�r���#��q�������=-+���-�	��*D���v�62=��g��>\�`g�LW�>*[#�Oq#A�騪�����;��{x����jM�jŎ��Ӕ����y`�ه�P�{��n�Eh��"���ɵa�&)�T9�[�e1:D�]&�]L�.� �\��KK9�-�H;/��ksL]`K#��m���D�?��X^�:��g����Xp��	�4y����@etu�8t���W��Fn�xb9��.F�F�>	�b���wKF~OD��"�#���N����������([L-�ߧ
?S�Zg`6wpFS����5%<�SU�5�0��HTk�6�3��������dQF�4��
���-�l�bT�0Ik�*���b-v��/�?+���S� =[�;wA*}����\�}n����}�dࠊ|Nu���p�w(9����Jm׭�pr��w8��X�v��t������lM�7����h1���+���zo�B�cB��Q��37�U�K"���+*�۽�q�DA�y��dD������B'��,���2c�S)�b3�}`��6X%=4���)w�`�Y^{���Z!^~�����t��UŴ��cLyb^����(�؂�Zk�ȅ�l�ITN���% {�a(J��ߤvx����Sq��ʞ��A���L�XiV�X�z
�s���Ĭ|Z��K!e�i.{ ����p��η7��a���ST��&k�Y��b�Xf�玔$qP�j���;R7I�~�#���/��g�d�����k`h������n�?�Fb%?�i �;F;�;g��y;냿�ͳ�q��ba#<:~��?W��]���{��7>|�z�LkG�����^ѧ�n�-���cu9��ۈ,ѩH-�����0Im�8�0H0Ks����L����:/����`�"k��muE��z�ԎH����Ϛ��{��g��[�ӆI�R�0�e`��)���"G��zz�_t��'3KTp?��^��F��	�E&�.�/������uh��pyOy�����J� j�b�(����ŧׯ뽑�^_'��r�T�)���H�w�Q����
f���Q�T����P�MEE�<�o�7ӄ������m���/̵���a�n�l�O�I���5�`��Ƴ$.\}��#5m����/MTDH���6H�"m4�A��
߹a/�[_�0���MV�$�Px2���!r��IkmK7�����$'Qb���xC`�f��ݶA��&6�`H�b�_���������5��
��`����z�����'�4�D���'�2�0 ���!���B5�q�4����45��9f��kZ�/�4�mb�.ھ� ��PQ�;v�,z;�Z�.�c�.��>�����%R��g�.�U�e1RlN��g�o���E�����#̬�F�e��#$[�t&{�J��|����r��5skq�C	t��k}����_B��X���_�F�uJپ5,?����
x�fs���;@��3yrt�I��
\�+ݢ�(7�����ވk�)t��2Ưo
��NE���8��h4t�Z���w�)Z�����&l	�*��6Ak/��f�����"��o�.�c2�hp�s�5-Rc���2���6ݪ�j�G#-Ґ�ㄧFh6������Ph�57��MXz7jx���c{d���9�!+�hfIw��6�%��B{q�Yre�� ~R*��Y�i�lz%�9tC�`��d�?F�~�/b0`g�Y l�"`��pH���1\��u����	5q&,�zg%�I�'yx��:�'t��j��0�:5����_�hsVCݻ0ѩt�QX��~F�`�]oH3�����D[l�{)\|���(�gF)�v M��]�t�N�J��ӯ+Y���eN��t+M��y�
s���$�ДP�>o�M��"��a ���D6@�'���Wre Jk�(
�Ƨ��R���98�C'Bs��e|�^{�Z~��n�IW�MR0p����;(�l�;7N��P���:FI]�h�y��T� ��'©���׳�0VEB[5�ra�fw��;2���E�2�w��,���<Dj���?�5������]���A�@�s����-
�'���jG�0�Y��_c@�R��P��R��w����j��v
-�+��g�Y_r]
�\�eA�o����M%G�<)�n`,�\h�6���?���g)�c�eU�?PZ(�=z^���x'���52s����Ծџ�J{����~L�?�B�Jy95�_?�G
}_��O]��6�D����p�uc̩�UϨ��ʌ�Eb4[�v�?�
���7.�?4� L�s3 ?�K��� �/l�/O2Ȝk�R^��A�릏X�0�q�:|-�Axf:4� �/��-���`��"��9'Q��HF��
P��[Z�$.��=L�m�&Ud3���48�m��-�V�!���YN����3_���t1h���e����z�����^*���G;-)MɈ�\d���򺻠�����@!2}؀��g?4y����8�Ί�K�o��E\{�6>F�-�CL��01�#�u��m�g��]�U���9z)��?P�cm��E�c?y������A٬�]�d�`3t$����^���<�X7[��z�J�v�TR�X������謁� ƌ��-�O��RU2ys�>I�e�@z{��_}�i�T�a��;���	
������u�o���k�\�з�nH˲���M!��#ff>���]Z�� �wl"�ЇZM zU�3���Ԝ�5�K� N����ޥ��+7پ�?�䒓�pkͅ��G镢V���fN'H��Z�b��>��D�0W�p�n!lmaM����z�DasUsF�5�#��	��*:eL�?eNQ��� {cc �ִ�2+'���:P�wD��F��l�oDZ�)�T���bt��O�aq�}&��&�ve��L �ӕ@*�/���"|�ͼ��F�NY�
�>6��A���w+�%�uA�V{�X�ݧ�̲�e+Y ���J
���edU�x����Y�z�����X:����
�n�4�ʅ�թɮ���n�����Kw�P��;� �n��� ���si��߼���A��m������C7��	�B8�@~5Q�la~�V����A��+ �m�A4�
�	�Io��Z�@�.]�1(�^yfؘ�FRp��q;nlc:9{Ѻt���*��#n: }3o��Cga٠���S瑡_�t����lk���8BP��9g\.�|��?��D�l�
C�YQ�J?��<R4�}��|���JY��|�h8<f`L���cog����T�Hwe�:H;9|���@7c91���	��~�ě۫��1�� ����S�"�*<o�	�0OWx�M)V�%л3���K8�$U���G�Zn����򚟲w�����B���;2�5���|��Y�Ŏ,g�_��]�Ŀ���;7�2�E���Vi`|~?S�<zTG+�[��MS��D
����p��=�j��s�"w�p����[>�%�J�ɳ+����?���EWõ� �){�>������v*�f�%�I�/�{�ʒ���#<�![P7<�M ?�í g���ȣ;A��}_�W
�^���k����S�U��׺2;%�t�����N�'��Kd'�E���
-U���X֧��H�~��2��<��&F�	1���!�t*�%$��st��II�U�e6� D�x�*�N��4L־l�|M��� ���ਡ�<�1�vT�J�vA�}�Ꮲ��II�g�Qh3�?+�� 䣓���]@xQ��?��ԑ��i/op��j�~��A�bh�F�[\7ڝ^(�"�"
�sy4A}\��^�����=u���$�r��)o��r�yf"�#f�Mr�O.$=5�����{ Z{z0�H�,
+�,��9�_2.�C^�t�2-"��q�ei.j���s���a٨Q�<R���*-��7�dޜ5V<+.u�y���*(FxpH @ ��^�;⚭C�E�g��H)�܋K�x.w�T��ww� �sN�$�[�F�u�(ygy� �ß�򒓌��͒W8�Z�&�� ��(�e���*Y͑�
J�/��#P|X���=ծ�q������=Ն�C�v����oD��{���oQ+0��4hBX��t�y\���t��e|�p�3�h=& �?K�Z�)�Iֶ u/~4�s�� ���H� ��g�Xĩ|j}�93�A3��0߮��O���1��>۬��s�d�O�A�Ի�v��ݨd��@�֋������ANc�C�O�;��7������p;��z.����D���[z�y0��&3_�RgYθt_�/��E�ۑH"�N�2ET����5�|n�g�Hv�WMzP�*~����H-�R��3Nkr��\�凃!���92��c�槝Ѕ�;�By����\���0�{lDY�~���6/�&t�0�>ftq/�3��f!꼵a�LPQ�~�?l��`���[��ZO�Bn���;a��t�
�NQZ�Ȩ��M#��Wp���`�<J0����'b+�oK��KH;�,�"��9�H�#���y%���X��m8�������ʕ��_��Pj]���P�ER�N�6�I��.�(�z&<�b���u��N�4ĠE2[R��2����A���oU�8�ks��q��T�_��IK�������uI���:��0�g2����0�h���d�-v�m�>|x:���:���*�u��NI�$���#��::��l���f�8���4-��I���M:i��]�%�ݜ��2��d6n$�T��}���,�~Z�������h	�K+�>��2��h��q$}�OP�)sX�}X�}	DO�r9�{Pm��;��TiFN���RY?�Y�5
/�T�xF ��'R�2�R�cΨ�#'0��RP�d��YT��fײF���ì�(G\�]�J6�2�ث�[U^���9W��JM�?�W��J�:q�����3�N����W:r��?e�3��<�/Z5p~�NЦ�?��.9��ٖp��������ab{�#�C��ѡPT2����(Vug��D��|@�Y	�_�L�i���p��d�`.�� 7�qӭfߖ��W:�Kn%z3�b!��gM�_�`Eq�ok]U_�Zyo0�݇TJ���ПC�|����;=��bPG���� �'���l̊����3��Mi"|<���`/:&��$�nK��$Q�69�3!|21���딝j�RR�Y%�f����p��ǟ��_��l���kͯjChh��t8rÊ"-rY�ur�V�p��t6�n���
E�x��7���@s7�5K��bo!1[��j���5Կ\_��)	]���`2�ҝ��|�����b�p�_[x�>1@:6��`�t<�E���T�i���s�C�kU!K�|� �w#2��ߠ�����,���v��r���9����}��Ӛ�fJ06��
���by6�&�3]�~Ĺ>JK9i���rz�#]֘����{���O��x�� �I
��}��*��'�B�>�_�K��3�]�����)H��6�m��dT�+`�,C�ݩ$��O�������.w�,��IP�d�|��݉u�I��X�&VwT���6&�$
|KƓ(ٕO5^Ir`t�{}p�I.(2�}��7w�phd�����."��4:j���
}�X����j'5B�0*9	]Ļ�����*��2e��,��& ��s�D�K���@��ѽ��i�4��a��Kb���"��@�6e��:ӌզN
�_^��Qo�]2�yjJ��*mFa��=�"V����w��p<Z�Y�-0p��?8�%ZR�p�տq�9z���cI�V,��㮉�3�2P��ݧ�k�(�a����o����^3�����.u�f�"�;� ���|�ӳ���p�x����	(��+���d�����Z���QE��8������u6O�F�_|���T�-�\L�S`A^��˺���Rh(9���0�� ��3���Z��9��z�:�EHv���*>�xo�^%�e�gA���ۄ��(ht���[��'���R`��ޔ�	�V����<�>���;GBV>�{��A���S�kSŭ�q*��JI�c��rma��}�v�+�I&P��%2b��L���\O7��0��!�R�񣘤qE�B����ɸ��ɷ��+�-��3�Vw.����w)W-<��@������X3�����m�os�+٘h��gk�%����P(�P�9�:_�!���L@�1�n��9�Iڶ��0�H5)l���j�D�����j�Sɰ�;�p��},z�^ף�|A��ɩ��p��.2�@$��hW����,�������X����k!�$_q������*Z��;X�-�1��*�9*�e֦�l�e߼�<�L��M���ց�]���W����
�!0���X^ ј>����#��ڌ�Ƨg�^�茕g�;�UJo{~���e^7h�`��;+���������_����&�4���*^~�Y�Q�ت/�^�[�[7\W��r�xL��ۛ�����t����Y���p�>s��e���R��R����LV����M*�"ӌ�\��:�H�|O&��+�5m�5?%��� �R�	��he=w�Ej������|�FK�TL�
���/��`�8=D������Mi��ؚy��i�fdN<�%�ls�\j$��>0���X�~���"�z�������$A��I��{��0K��M�nB����)ג��Χ�F2��f�=���g�E�
�\B���B�MՌ����������<k�ulx��cNG�n��gN�O~�@Ko�