��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[������0\8�J_R8�C�{B�z��I{iE9�Ъ�+�x	/q�{̱7\j�2�/<^�~I -t����o��1
�Y92AY���u�)H(����͠,5P^�V�Z�u��rw�`P�tR!���	?vM�i@YY�h�S�i����ȬNJ�Q;��m�ݸgF��݃Z��^oC�g��g�`;�'�gA����v`��#��^��PD�{"�pnfN	C)�=/Sd����I�V���,m��k�CCQ�q�Y�����ٰ�]-�aʿ+���rrI�Ҥ5ՔY+�(���ae2�˳x@䒺QdF�4�D��f�@��4�P8�Jm��zÏ������bUO��Y����>�CO�e���݄0�BD-��`�K�P��v}�{L8�>-�c����3������$��X�~ ��=3�y�$�
�El1P4o���W�����VSt)^��o[���SmCƝyZ:&��񅣚�GYx�K��1����ĻS��֡)�*B�wǡN�b��h@sv���\��|�fw��'-qW�Gb$Ȫ�*b$H<�t�Ӌ��?Ɠd�?��B4�}U�uѨ4R��q�I|	@��Tm	Vs�G0Ֆ�쓖V>��w��Y��s1�]��ǖH�~@ȩV]W�e���&!���۲p���!�WT�`����L�KJOW�ry,l��Is�%��SLB8Z�!x���-��p���4�!<�2�~��&��ڬc/�V�|4�[~=�Jq��/4�!q��k�ɡ�דC��7����Q�[�0��A9]��F��M�x�}4���R�䅅�B���er`��]D�,�	9;X� 'k}�2�!��"���,���r�7U�z�uJ?���rUfW/l��>�|��{����W��Kb%�՜�>/,����El{baɔY��O W��0G7Qݿy��!*X��J�eG�R��~�kq��A�0�]3�w,�y܉iH/?T���Q�h߾^�!겄���>�F�V� C8�[���n�4�,d��9���Ś�I�D8�^C������4�¬UH	Nm�|��2���D ��|��<GB�l�!��A"#ě�%�C]q_�	Y�68xM����y|�_h��򤍅�����?K�a��k&i��m�1Ӓ��L��H�C}_4�5m�MC�nX�[#���&���$g�S0x3�>�=�����u�� ����nuA��Ӫ�s{�xt|�x��G���gy���Հd9�I����I#�����g���`����ߢ���#Twy����I�)H��%;�z:��]2�A��eD�A`/��9�]&��������BD��D�!G��`ߌ�ب��C���%��Dn%���)���?$ˑ�4�_<;�,���of���'�ν�ɻ��d�P�f�p�|��mQ�Z+��Wd�,>O�0���+9�
q�|ձ��O�#{�}�A�#�j�Aq絘�g���icw�y�:l�H���qn�>@P�vȾmUȩ$p��c�=�}�n��қ�]���6ӝ/i��*��� ��uح��sm�����VI@lH���(�����v�Y_dz;��iJA�AG2BN�H	�6f�T�ܣ�����;�LɟR"*��x9��������KZ��vM�87��a����J�WP,�fޱZ����1&�0	���
�n���ū�oJ@��Uy��L��  '���)�F�Z�"�_�2���F��đ����\]�o����Z_��3E<��kʬU���wq��u���O���B�^����V��������*�ْb\�SN����"�5pq���CJ�j�%-δ��p������-ױA 
)�Ne�u,�DYgu9/I>E6\>��� ���!�Gǥ���&�W��ev�yP�D(-���z?�1^@CDw� �t:G��@��D�i#�X=�"�~�`:�SF�*��
�8���c�Mvѷ������Z~���`P��_>��u%1��6$IN��?0��՛ �9/��O<� ��YD����8�Y5�K�7��~+��G��z=���=D�y땮�v�_f�sJT"���č���o�8e�AtPxc�k7���}��Zbz��3�� �����V��}a�� A�F��<�r��3��(gJ͖��:[8���ܢ.٣\e�*�2E���fD���ao߷��b�c��p� &��ͩ[��8�n�=f�ƒӽX�6t�P	��TeR~�����,7c�e�O~s��w��mX��]N����> -P�X��*�Ƀ.p��lc0��]�3�8H��!؟S2�w��J�����*��a1vg�p�� k�j�yh��,n<V�
��0n* �$�Užz�P�{�h6 �j/��8���r�b��%�����U� ��^ё�f�g��yL\p���L�- �D9��y/k$GqR	�*�K����LH%ֱ˞����5�1��z�ֺ]�q=��h��;3:5Q�m�6�?�D�\�(z�1rk&b�t���D%�u�ydF�� :�L��i�/Ot���P����1�����X��7��;~�Dn��IqlȸMݛ\��M�C�Af��{�.��,_l��X��[��"��Ep_��S|}��S�*��4�Q�%⺝=0F��2���-V$#��4"�\����UW@��G��	 R�y4I�d��r��������0��m~b2����y��U��~������ß��X*mF]�O����/��jbv�ySu�2��+F�FA�.kY�C�3K�������ߠ2V�~nw$�<ײǛ��Z�/SE��%^��
%(\0����yd�퇳���`���?��G1��J,}d ��W�9�5��`��!dI}� ��YYP��;F������:s%8��)�p�iK �v����<G1���q,��s���-��?���l�T`��3 Y�z@�G�K�ȩK~қ4��]�c��1��
���\�<Q��x/[	��U�#��Ldf�a�XB?j�����4C����p�^�_�G9�T�O�Aq�CnSqK�N�e9W�9�2��M�}��[t)� (����i><Ŀ}i~@���|�H:!��7H�U/䒼���+M��!
�Ni�n�0MY���z��m�+K>��K�E<�*X�5ƋY�}�Y�\N6���1����`�v ����_����re �~��hH�K�P|��(������^��� a��C4�d��u��މF��^���00M��m+a���>H�6���A���(�,0G�;��k`qt+7���q8fɩ���#��j3�����!��T$s��0F+"���+H2��?�:���7DӘ��d�]�l)1�o;t��G]lg�F��⋦���9+�"��мX�Z�<yc���k�mL�M���	�6Q��`˭����2�Z������4�kW�f �f)��I�g	��^�Y� ��xXY�G���aa�pAoY��v���YE�C���L	�m1�ק}��3/4G&P����Y���<�=��?Y2����iz�U� 0�_���JY�a�O8v�Jיĳ'Y�-o��#(�<b����p����Kz/k��:}��r�u�7v"B�9�S��������N��DR�qE������0�{z�*ii}�����I��ޭ��zY��#���!髼*K���AU<�A���U�;��$��m"ɚe�?[��}�63#�wv��ۺ�}�'�n�{�Ȗ-�2��]&��N�g0=k��<DW�:A=�*��뚫O/�`Q�r���(n!;3.Ͷ�S��XJ �K	B���E�j)&e&#a��lR?z�A���[꒕w�w�������S���3�R7g���F���W]N�V*F<2��鸧BB	�,�@�����pX�xC�����`?�7��M�����41�}c�@n����/�a&^~�4>�BG�R$-�����S�TAƿ�{�<�Nq��d�c�����R8D2�ٟ�=�G0���\U4�/��������ùk�wq��U�p�`����:Y����^����-��@��g><h��2ǥF[7gN7<����>)���T�'p ����uu�i�Qu6~�X"��lC�d�1y����I~�m	�"z��p>_�o#�� S�>kG�C�H���8����舷�c���z���`�����P�^�v�.,!v���Fe?��г�ʋiq�L;搩BFp_��坴uZJ��v"��%4�E~��+�������0:`R�ɦ^{^k��g��Fӹ���3ֱ��B�gH�;�܍\2��\����7=d'��i/�Yb��R��U�xԶk-�m�T��U7�ιZ s-��_)#^��5�0N��1��7�\񈧪/�{U0�-�g���4�:�ݩIO�+�2���|��aH�L�h/R?v ����i�����1��p�P��uki�cy�����7��iA��" (�<d��ػ�����Ȏ=��dT%O^m�vɯ����{���gͥ���9�����R�p7��0<V�-��L/�KU��2�݋b*������d=�T��zL4�F ])�o{���?� c�y����\c��B�݅�S?�P˲�+W/��93���?����@�R�R�B�A��ߎQgCC�ORmS枼r�_U?��J��%6�]C�Cu���YS����K�Ԟ�j��̟h�Yn�-�o\��յ�G��"����Z��� ?3Y�H}Ӓ"wƂ�e9��K�u�>qm�.�o�����ǔ_a��:��DF����B��Oų���(
�Z聡�W:�z�0�K1������	�"�d���P��i��fH��i���@Hǧ�ܗ�P
ƛ���j��&(��R���^���8^ �AXʏ�S���h�X���h������mKf�+�Iòڪx�j��˺�3Y�air��<�T	��v�w/�qiveҰX#�|e�e�������� �@�ڻ���p�
�E\�M�[]A2��t%n�hVb�,!�f-vo�o�#EfM�)4P>���;�E�b���ߗzL��GTU��cIQ�1";���=!�s��0��\�$)� O_7�1񨁼Sz��4u��N�� �"�:�:�j��V	�߾C5�~�ay��^�sd
Q����H"���	Yn7w�G����W�%c�CB�2Y�y�;uD�M���UA7�����T�������dku�M1m;�?��٠q2W-�|.:
�Yo�>\���A�%�{��'� Vݑ�����n��Do�$ҕ�� �φ�ߝz%��v��f���a����|Sy��sc�U�##�����6��p��d���j˃�懿f5�1�CP��U���)o�J�>�D(������g�ż��?�:y��OR��7j�g ��hmJ�O�����'������(�#w�SR`�d�k�,%/�qS�k�)L�hHb��7�C�]��0��U��V���(
��S����#���#�����;\�H&Q�u+k����sr��	l��FcL��,��L'��?���1h[f�W���7�R�Mhp�$�Q��>�Kj�� e��Q���h;)��2|4�hQ;EP�G�y��u��8p(��]���*c�_M�샯�km�������ʚ�Q�`�r{�*T����l��r������eJ�s�<.m��+�73
:8-Xa���Ӓ�$9��f�K:�4�I+�ܩ?�����21n���M��'���"s`-������H��m<t�W�,���HNI0�,�� �������ޑ��R¼UM�7��9K��M��I�����u4�TrtO{!��D�3�G)p"�|j�Bx��hs�����:��A�J,���q���Xj�8�jL�9_���3��c!S�gn�z�k�|�%���sI�p�M�O�B���+���6R��61�P@�!F<�y��$*�(ec8)ޭ�gT���q[PF�9��
�<0+��Ѭ�s�d��M/ ���O�:a""�J���92��j쏊�aw�����\I]����N9?��<�9��C�o��Z"�nv����AfJ ��Gx�4�ݕ6�F=PFR�5���Oc�2ˣ���\ ��Ū|d��(U�=���Q��9$,)��V̒@c�!>�n1[�*v���vܝ"��VZ�U�LC��Þ�}�D�h��±�"���bm�f�|��G���������*naw�W��fzG$�!Ű�
S�oϓhk�`����v��:��lo����cRX��ZG6����*u�_����ǌ�&��	�t�2j�C�j�hA�Im�
3Ͽ ���<Ľ6M�d�hr�<Q�Ӵě^��yJn�� i|3����n�P��;���:�{&a(�=�7w)bC-��q�9%Q����ڡk��ʪ�թ�7���@�w������\��v롱�����r`.��fq�p~21$�h����m��zV-��z�O.���+�_ͷ�W�1�59ы��Da� ��*��D۫�J�!	�\��|�����C�<���R���ACJ�,�	� �j��O�c̡rb�2I�=-J�%7Ӄw��v����S%TU�'���"�۝̺x�����Q*�9WRHax���SNV� ��J<���H���o���*lmK_�mC��GY_�����>��lMĝPү���M�ã���IV��\Sr2��T��}�n��< ��� ^���[��)��ckG	�4H�b�KWq�gG o�W�Md��<[�0�����3�����+9���%��J�����7�UT�!�����Զ٢y�:,���䭡a�}�S��S�X���h&�@�Ӟ%8�}�6�Q�ɼa� �c�������Ǹ���F���,(kEH[>I��$P�Z�����ś�odd}��	~K:N���L�W��������G�ѣ�
0�¡ǽ�J^`C�_\w&��n��'0���g>Xf�N��~r"��M�o���<��,�u�u���ߋ^2j�u2e�؉��;�����ث�E֚M϶>�sUy��G�|����=/dc�hJ
((���á���i�Mi²��$	�ɗ	��F��C
	$���l����D���cz}�%Y��3�/�7��; p,c�$K�[C�g�)�xv�od�n8/�q�"km���$1+�Xe�V'��Z����B��rl�aN�>��������KL9�U�������T������(C��3�@�����S��K�+�@�b=93�4X,�~aK�#ӹXҊ1� c�x�Ґ�@���
�,,-�2&��L5]�n���zR��N���褛AJ��8��PCƊ[�&���P�A�*��q�=ŇuA�G����A䵖�MAu�W������]��Ti�q��`��x��(\d9��}��߳iNJ]���{��eg�yp5W�#�p�E%g���`����`�ma��ܡ=� �/z�K�����V�m>�&P������ca�-w�P��Y���D�킎h~������s���oi��~j�(�23�[T�qř�L;(��{wB���Q�d���:����bC!o�0���"�z�W�M��{�~��@��xҾ&��G��S1��Zy���7g��=�B$E�g!�����J�?%��.���Ueĵ�5��O��D�\1�$I���z��\�����q��)~�s�Q�X�L�'_�b�WjmiN'�lo*�7z����Ry_՜�p�@<��
�o���[�[�qLg��o�d���zJ.��C�&�2W������ἇ�\%	t��jf%E�!`~��.��l��Ϊ��Q,����|B��L��;�I}8e���`�e/zR��X��*�ݻ�*�f��-ӍX>��$� g�g�`�NN�
�Fp3�1��1� O�}��ű�@*P�Xv�ڗ���S<2I�j������BIz�h�6j�}�rٷ���c%(s���^�ŌBv���=�W%�\����'���"%aA͑�7�j���hs�8�V�b�E%��"�h0����͖l�����C��5�@� ��;ܶD&��v	���}O1L��a�� �9v�Lsg�2������}�HFҡK��#e��t�h5�����E@���B�a�1���x�����B�d���\���t~{��Ř�, 䬵Y����믫V�]@J�F5-P�iB{D��']Q.�.�e;��{�!ʕ-h3��BP�y.o� ���?F�*6�v�W�pSo�y�F�f�?�z�Y�ͧ�d���_�m�
���CP7P�K6�Y�ٴ��bX�t"m/�ͱM��p�	�MN�F���ru�:k���v���R�y��
��-a�U�Z~�ӸU��[��� ��p���Ϲz�S���ˤ/�k#�9v�X"^$��.0̲����g��E�����ܴ��gq�@`��v�]�)んE����O͝a,����C���׭��i��HEҋ�M��O|�JDlܷF�q��@��1K@NQ�jr��t��Q,�[�����g�2C�U��KL�J�f�B���ߨ����g'�3��9hQ�Rp�>���oͥ���$r�h���E�q( ���sS�٥�,��N
	�F�*R1���_��)��b�*)WXU+�	��Y�̃��w����{�-�"�B̷�r4ν��Q��Ǐ>LW�r&��0���B���)s��������3R#��ԘS�����r[�}������m��w�E�K��%BI�Y04H�/�����]�hd X�^�D�a׳{!�\�o����W{�y�M���@�>j��a�Z�N�_yǨ׾_O�C���g9�K��w"����4��/���Fj���>��`4.Z0TB����x�ȄEEq���L�ɤ��������A����2T��~�2�>"vl� �/�K�4V�M��5bx���=UTq؂fO��K�R����-mZ�s,LA�k���ҏk<�6��]+L�gbsmh|��xm%C\�YS.�����rcZ>{���٧(9���l�n;7��A�\l�֌�����E�`�c��@��$>ףT`��L�NKR��z0.��z,V#�$�Kc!�O��D�m�ye�YӮ�(K��������0���A�ᢋF�jz�����%J�{LΆÂz��F��o��/��Rd�܂%6�;5E�F޲����إ[�qn��sbm�̰ѻ7VE�o����Q@p� T�c�#�>߷U�8}c��1��O7Mʈ�ݡ���n�|�5���ذǲI�*��W��_3���Š~��tQ�-8;ZL��x���Z�ˌѷ�<�*�dZ_KY�=�Cq����#�m�:xTvJ#��F�B *(����"V<�g8� �X ?�ۃ��@]M|K^�)�絢+��½u���(`��1�L�<�%K�'M��
}����1<\h��V��4U��-@,��>�@��&�_9W�3Q)�e���k��p/^w�1lztK�݋�������`d��5���8��W��v�U�7��=8�^�Ȅ�J�sP���w�19�[�K]�l�{�H�*5�6o���{e�p1�/�lՕ�K��ށ�.�/<��Tis���#�9��j� ��9lp�0���T�I��@�HB�*����{\n��a�U�7���~i�S����]}�W���YeH�-[�X?�-k�r}���SaW�'t4����)�22�8�!z�CL�{���s�0���q�Լm!�P]�>wuH����"TQo���,���Qa>��>ۛt��?Z��(�O�X��~$��Ҫ1�S��?�aW�)Q&���\n-�m��ϩ���oYu�̯�l0�J�[��a�F{�n��L("4���ڃC���&b	�S� ���v�����+����tS^16��8�&D�%Ǡ��:��~��'Z�{Sxy��h���f����8�Cۃ�Ƒq+r&V󈃔�Am�f�&���[H�h!�h����h�<�ޯ�:x�"�p|�~|u|��"�@�.��6&Ӆ!�B�� v٨�����#av�I����aN��_��谵ڠq�h��p�@�RP=��vՈ�:0�V4�r��
0(��nHAz�Mq;4"	��'�-�e�޼`�6x&���{�]\r~�T��y�Z�n��
� v�ӷ�s��ɴǅ	��B� �&��[���v&�A��:�H�:҇����7*ȭ)�*�Xڈ�R�7`	�@��}��4�?�����u��͘.���!�`N ��Z/i�k8uT�"�3��̣���3 px�#�@7']�0n��,ڲQۣ�jc�Ev�SL��}Z�(�۩UI�i���H�!&j<�D6o����� �����D'��d�Ïd����՘eYE�~h���h��>��������5�V��p��<z�o���I�{'/�~6��bJ�,#i�ҹ<)⻠ m8��j�L��RJV�r|����0�e^{t��6�u���-d ��A�o@n�o���2z�x�X`�]@t*��3^37��5��KJ�u=�~�Wc;�PP;�r!�K:�P�[�L�H)�,�3A��̛2&��ܼ]<��g���Q�v��ҙWN�uh��b	�H�2e��9�.o�c����%�k���y�OG��Y
V��"�D!��1��c恸ro"33��p�ޫC=��NiZ��O�/�굏�B�υ^���+����`����(����Ȱ�ᮍ���LP��D����)�V��|�c�c7���"΁�fv��g�i�ڝO�{Xob�P�G���ydÃ賠{^�	$���P������@y��jW.1�����tM]T�����v@c~ū^�OK��t���2ȶ�=7��.�%������B��,Vv2nH@���,o���Y�����ƻA�2,�����HgWY^�'	{� qo�'�Ȅ�Ag/PR�_
9��b�۲�n*L�yM���jF"m��r�	b?�X����g!yM'��1����j����e]By�(&g�����h��(G����.w@�#$�	����;�#��up�^a�=����
V]	��b]8;ۡ�Xi����̾{��L���9��\$m8�`��i��� ��ED���!���
j2�̛m���+�o?��5�=��V6/6�B[y��HQEC,RQG��	�#k���}�1E�B�Ð�o�p�K^-A$�!w��Q#�뱪�2CI������n��˟�x�:���tj,IY���/�#jBg���ܫ#d5�B>���0�^s�9�.֭t�[��p/�i0���y�����3?�?�����n�%ׁC/6c 3�fh�D�I�ֿ,<[�Of\#�r���Ud��$�����`�m&"���:B�v�|�`�r%��i��&YR	.+����TI�jA[n.�	��i�R�li
�-��)ƾ>�󀝣o�N8R�Vj�!��s���ȼA��(3�g4�Wz���@tJ��J�1��B� �?y�)�W���ُ�A�kV�tm�ż��>4>#����ɹVW}op^d�M��|^�WҖp�,ɤ��*N0���۱�3���PU������j�<9I^fއ5�
A���e�B����{�ǯp2ƒ��� ��T�Jf&�/:�>��?����_R@�ܠ��
�����2u�D��{X��m�
�D��S�LI� �]��ge��.6o�PE�4�u�#��=?qJj��= �8'��A�������ا�邍;�8�����оĜDp���Ü�y�E� =wa6�4 H�UL���V��9���Y^�[g*�����qL��j��(���O�ٵ�����	�]�*���,�%�`XjJI��TqrѨ�5i�r砍ɣ�Ɓ�ۣ_��Ґ�tI�=��r~�����S��Qm��шʫ�gz���_o�}LU�r�2Qd�8�@�ʈ��>G�1J��ڨ��"� ��4��p6�к}�$��N��{����J�H	��4��������nr�A�H�=&�uX�H�.�i���<0R��g0�,h��%�<;˔+dEQf�r����r*+��!���qƛ��RT���k�c��U3�x�����f(�9�����x%���n��`4ܗ�+�n��A�2ϩf�G��o�`8E��,��w�mx6���NLQ���.�˦l�qρ��h�7������ޑ桙�ț��0�"��$o�I���l�ި�4N����0�4�7��ܛ�h~�%镩 G-����C�.����I��-�0�!�G=��+t�.��ؽ�6џ �EI�>.J��Hs�a��i�f��G��
�;BƼB��xη������L1{���Ϗ�`t"}𜊺|Px2V���I�j�J�E�x�6֦xw.��>��ö_�	�[�gFnj-']�b����ވ0�$�wN�t�R��(A�;g����ׁ��g���Id�+�U����F� ��09(A����G�މ ���T�K/4�ן�`�F��j`�ub�".���/����������:����6�_0��E���Κ��Jiӎ?+���T.�:f&���%K\֙��>2�>Px����n��{$@b�3�e���s ~̔�t�9=��Kg�߂B��!10�x���&�B*�FMy�&H	/�-X�[̝V��3�S;�o�U��z� I��8tT+7l�5,w��L��͡��9�M�@0�*$�2�դ�8}�f���Em>�	DY������L[T�Ն`ԃ٩d�gzN�`(����*~�'����!y|�l���T�%�kd�Zہb�O!�Cuj}��,?�])*��<L�G�ov�����˕z>����3���N�%Ө���7E��ˍ�s�v`w���f��8VQi�w�+����D��`v�d��R���/��b�W�~^t,�-$���h�#�d����u���s��<����s�-a��e, ߾�*Or�Z-9�/]"���m	�oJ�������i�d�D�_�0����=�wv�`���ܫh�Z��ڥ0�M�C�N~���L�ۻ���L�*�{ ���[^�@����8�B' �Af�=z+\\h.������1i8н@Ԛ6s��G�Bޏ�u��)Cb_�4`^�Л �(�������0
̴��N��&j8�<���N�pA2("�џ�'-�.����2un��(�
��EP�$]��#��Y�nI�)ZgX`��ƺ:�[���r���dI�r�`��|�.^�r�؍L�����a���q$=9/^NИ���*]̾�Ǿ.�u�'�}�����f�w�m*sg# �y�E����)�i�� �<w��l��hđ�I��j�)U��FrK[ù7$n���*4�FVjW	�2�ȸ
*E������Kq*�P5+m����%�˴��
��4!a5�G�/R�����pt�+��6a{z��b9yr�m��5P߇sҖ��O$`�s���[C9O~m���e!x�e��?�~F/
ysj���q%�G�{��������&�6k>�W}��"3�$��R%l/��� ��~�>ʎ�r�d�����2�u�O@�r�����^��.ݼ��T��[X5%�Q.<	�-ݸ�Uizq��5p�'���t0C֘d%�㷠y��-�}��N��sb8�����Wa�-��Ms;��jD[\Ez�M��#��{�b���3K< *p��F�$�灭�jW��
2�vu��d��n�׸�6����"�E�����B�7>9�����A���m���Q6�<�3��9�fR+UH�4�v�~ P9s�:��| ��;-�����UN���ۦ،�/�0�����|��Ot+x=A�,���Q1+Aֺ�5���vF��``N��j� �-�m�:����W��,��|ʒ p�k��J�#ے��u Nf�\|��y&�$dR>J�@��:��J��$����C��Fr%A��ad���J��F��w����~����ݞ7X��i��qx[����pm�Vڱ�ӡmB̷�=����Z}Z��v!���ep��Z��.8R��Y�$�7�����>p�"ԛ-��oڸ7D �����},���l�r[���ρm�L�98�XM��Dc���6ȏ�	��?b�}��1^����\u!�<�o�e��i^tO�_T&.�1�F�6�T�8�����\�P���*	?2�lwINUF�m���yMɸO�)f\�Mcߞ��q��s9X�<7f�����*[ٛ�!��1��q2�t
{�m0]�ש� ;%���k��X�0����M�%.��v�5���2cy�/Fs"E�����Vd `X���1I�4�Qt���xDv���	j��m�۞����u��L�;��%!J�qpwc(�b=r���V�Ö{��1����7���'O��l�4�'X��ԡ�<���ŵ���W�[��"+�QL짎�>zǫ� ��l��hfM}o}&[���z�I�'���%��4ԥ\K ���I�L&s��"����N�e<p��Z��u:��R��#�גC�_{��U���V+��`�B��YEe@���18�K�"e9��Y9}Y�"Ė2�/Qz?� �Ă$v)�	��c�e���@�8���<��]1�eÒ]z��%��N�קjHo9Ri3�^c�DV�F]|����sԲ�ue0�L7
�&�/�����-9^�"�y�oq)�q,���c5&jڿ���h�&:���l/�P��*dڎ�o۴�:���_�^9�z��h�)d������ޛJE��_����0\&xY9���xF�k�%G{Z�Jy�s��K�s��.nҕ��(��]U�`�q��a�}S�d�|�l���ʦ��U��U�S\8o�F�����2)��$kc���E�K��Z�uڏHЙ�$����@�ײ���6��v��]ћ`H���@Q��š�q�!RC^�����f�s��| �B`�������u�`�d�ڿ�-�#ؚ�L�^�c<�	c���X�J��"hQ�O\�����j��i�ʻ�7mB��j=oq�*�B7�u��J,i���׋-��y��]�'��<f���	v��"Vv�e��#Ms�_L�}��(�Y��ȼa��\T��8w�ks�2��L�AO�l�Y*R��(&�����y|Ye
%�+�r�<��~GJ��҇�^���2Ljd�ut�x��xl⩲��R�JrЯ����̍����f�2{Í��pz#)L�r��-}b�eE�����s�@+�oB���4sh�\|��HO�߼������ʐ�6V�Z�K���f�+ɤm�%BT�D;����U��2�#�=Y�B�s$��'��FR���Ů+�|G٫�i�z��u������6�	+ǩOU
w��L��'�Jf�+��Ys��GC�h�g�	Mm��j8# ��V<L��u�򠵝���8.~%a�q���$�=�ވ�/��NƾʕA�[ߺ���\�d$>�g�!�V�R��꽘��9zM��Š��Z���_.X�ܾh�EP]MFc��<@��dE�׈˥u1�W�Ȕ�I�y�]��*�W�S�B�Z��u�T�eR$H+Z.�� �+�&��LC��ϕ\�|���}#��{�QS��0�������n�R���?��f��M4��m.E�Z�5��v9 JP�Á�F� ��E(7�cs��Κ]e+�_^��6�9��e��ធ�o�K/�v�X����H�>D�k�\�H6I	|�7��D3\ �F�#i�3�/yM϶B������Q����%�>�2$�=�A}ꧢ[Y�}`��Q����|�9\������^�fd�Y�����>f��>�ƌ���o��K'���R��]~	�!e�#��h�Ucq�^]}�� ��ź3��'��fR�j+"���	��P�	ab�mQ��秹�:s^ҏ�7=?�P��i�
��f�l����� �t��2�O��/g7�~�	�H���/̄]M\"�f���f2��e�� pD+?|m���m�ò��CEw�8���8Q�^�ǐޤ|T.�g9.ډ@�m5�S����mM�3�Υ���i�8R�XI۞/��fV��z�9������`�d4�����~��V��nVE���A?��u�a��jh�m`Qm1wa���0/d���g��s4�������&����?a0����"�Tkx��ӈ�WO+��ّ��?ũ�l���Ixw�8����Yͻu��320�����R�I-C;|N��2��{��X�@.7����S�]��*� o@C=����/_}�<��`!�ۊ�
�A��e�{:��r��k���Hq��w-�S�W��E\�Qm ������u~�Ok��%��͉���~x��Di��R���Ў�I9��KE��>Yw�y2Ѿ�x�BQ��kU�ѝ�3�i4A��.F�'�dᇏRzl�Sdo4�[��7U�cJi�$֐�"�NWx��C���wUd�(> ��h�Þ`�ι�_R�����j1�Y�dP��'��-f�χ��#]9��ն�v��A��_?���6�z�'|�抡f���ބTi,G�<=y�%�=�물*�p5�x���d���_�
F�D^+SE	@�a�h,�Ǌ���-�]$�B�����vr=��aF����)6���ʑd����^��߸�t&&��	:U��mf@>!L�^2y��@}���Zv��˴�2ڶ.L]e��>�s��9,�ep���W�C����������wss;"�_-�W��	�̅"��ʖ��z�WN ��J����]܊\�U�Il��4��P	 D7����& �@�'�����#YV!�թ�'�&��,e�7.�Da���Im�C�x��׾͚�ʶ��Pj�A1�_�F��а����z����J�sͤ�szB%^}���� ��	# D�\z�UH���K��=�ZR~%]��g�)e���etu����*������\�oppS�������g\"V�����{����6�ӳ4lz�۔�d5\��p#V�g����95��w7�F,E�!I����X�R�p��^^J�D��|��I�ۀ��S!���.�^�ʷ�SG*�د"�ٓA��(�꛼�V}�]S�`��4�8�D�`�xǓ��/�
A�D�h��f�N���~�i�П���6��EZ(�F�/�o��V� �AN���#~Ū;W��˩��!�����ig����|��;FQ;�z0 W4�<�6�4��ZKx	$�K̫�~�)�lR�z�T�x��Y�ӟ�N�B���Ҳ���Tl,W?��d5XtE�ɷ4���P�|����U�9��y��<�˘������K+c�wv�3�������!�b�Co��0�����
�N���ݿ�^v��	g��f�&B�1��#Z\�6�gq�wwL��H#�7����E� *Y���."����������	��u��*�dK��3GI�!#+�/��ζњ�����ے#u?ߐ��xt��,�)1i��/��8�<� ����u�c�Y4yukn�9��m%8s�gnd6��粟��ڟ�9EW>��(�6t1q�|�&Â�Q�T��,n���0ʀzN�F���d�b�_�ꬹ��<��3�a"PУ�wt"<�>eÑ�o��O*��F(b�=����nGx�]{>��b�+=E� �<h�8��ّ�gK��Ecτ�)��p��f����\7Bz�_Su���~��e�O�S�D+/���p����&�S3 ��t�#�>z3�F���2\]�K�|[���c��θK)��-I�t~�5@4]���`��u�lU�M������Ӂa��b�9ӆc{��l��?�	�������Y��C>��K�/h���mː�&�a�?Zcw��̘ǘv,&����،�Z@W;�*Y�w*s���K�o�ZH��QW�`:�К��&��/�5_@;�A��ǳk����W&��<��M�R�U�B�8��1��
�H�1���tu�[�w����O���W�2�7o��-n�;;ź�U���(�����4:=Xc�f~E�z�>+�o��1eD�=��Ѵ�F-���W�� �����S��Ǥ�d~�M�2t�dY7����K�nK�GR��*u��Nd�"8	��x�9�X�tU<�c�"J7뵎Â�������N�pJǹ��v]$��C/S��ֹY�
m�ep��~y�2^ �F;y��ن�h�9_N��|Ǔg���a��Y����d!�P"G9����N��w����3!x��қG�FE0�5yZ#:�.:����.�N�n�A}� ��l�ˌZ٦���,���g�/a�\�,��=nA
�����sR��x=����ww�9w�.B�^�ۂ��'��-���(�T,d8�I���\R�+���v��&��
����������K+��r}'b�&^�L��ˉ�g�k��v Χ<$9Y�`U�tw�;2�_�5�UU��S�K%Y�����ʂG׬�܄�^+�=��/bH�**����pt�;e�K�.A�=W�d�����$�F��޴c���j��g�P����s�� g>���/L�� 3r��w�6������qhmq�h�?��ԝH*cn��:5��SI[i܃a�ѭent����	T\P/�N+�g���
�[�annA���a8k�$�u��m��4��("�F�X/T�t�8^�L��n����oSBգ&��	�B�r��!�K�[��D rǎb���_�v� h�|y��t�����4^�@��.�H���1ψe�*����2f8ʁ�Ʀ�3%p���P�BDU�H
�t����g�t�чP�¥�0>@�bu��*��� u&wm^]1,8M��c�$���~�E5�E�W��::)�=����(}�FJ���A�Qۋ,Q5ysC�|�ؖ���{eH 3�?�����lԷ,�[����<0<��N�\��1|��>{�$j	1�%G�GFr���iC:U
'�/�ڣ�)��ȀVъϘ��T�囑���2�1��\��	G
LȊ�dU�A@i</�Fb��u(
��֚/�P.�.1���������"Y<xZs�����5�ܡJ��MC�lc�,Wk���Y�Z�L���d����@��[��d�@�A�s���x�d���~Fvh��k�+n��Ő��ke4���t�&�/�H��)*�u�L
�9�d6�@9��ٗ��UhzrrSȍPÁ�EvZ�.wu�JVB��$}m͡�b:� 2��z��u��嶣�E���3EE6ԩPU��� ��.�^+Z�'FL��-��&R
`D�u�Vڋ���w7��6eM\2N���Lr���\�̛��� �
W���uYP�+�F��Y��I2w��h���)��8f��!�X�E��冏��}U���:�εPS�y3@�0OPK]x���W#�+�|��a�������-1P�!�G�@��P(�Ȇ�u2@�w�6OD�{t6����!Ou�أ�7��|޼C��S��d��N�~"n,Z�Z'v�Kp';R���(����(��J0��&E�kRT�O��ݡq�{�Ys�{���M�ξ�'�����7�F\HI.��T����g���9�~D��mb�|<�3�X�E}�F��x�I(���G���7Ԍ��9U�����P���/��ߕ��K��s'!��ވ��W���اA^]b����=��@�t@��×��Z�{�i�w���NQ"��͓^Uk��DJ za�������dp��{��`�?�⁽�����J��c[+0��U�+�%N�Lx�R~p߻`�h9�ƶQ�gT��h/������`��呃��E�Б���[ zH�i�VW:O�eَ�=V�����<�H��<���-�\g�1Lmܟ�N#`�	�|J�����+�����Z�W6�3��X !� �3���4�!2��I`ѝ�"�Dk^K1y���i�v�,����&�?jq�%�BΑ�I�b���K�,#� [u���=��hIg�~�<��Ӎ��ʲ�_�(G4;*}s��@�@�GQ}+����E�)�`֝;��a��V]�s	�g�>�,���ԺK*��c	��{�w5�9���5��p��(��yl<ϑږ,H���ތ���S�w����g��U\ ����;��'�[���`����o�\�����q�R8��Y�LRQ� V��AV�����SS�A�Zc���r���{�{�Y;+�|&B��Q�j���9�Qpk2�J��Ҕ���J^��~\��tz����P6��#k�$ N��=���0�0�O�����*Q�v�?$֎�9rc֎�+�<lמ@<]�f� T��I�z���M(��+'���<hL��Á5����$$j��T����36:�4�?�C���P�s�����4�i��F0Rm+k9���l,bT����ɐfmN]�U�-��A�f�a�B���/�Hʉ�~u���֘f�qvy��顊�k��!���Ԃ��i!ϕx.|q�&	f�I�u`
�8��O��Ŗ�ֳ6p���0U�#g����BsS�#���~rZ�_�ZQ}z� �� Bw7�x��q�_[����H��/c��5*�X̗OT{�Y���pGH��3E�ڐ�#���/ԧ���V�� ��'DԺ�q�|l8H{����P�ӵ�E��|&Yw�\� p(1�z�>����H��b7�M����y�ˠ��n��
 �H��n0hD<nؓ!�O���Pl��(8q{*80�����O���pi;D�	����l�֛�ߘ>Q�t-"L�c��X(:���w���G�yFn�u&�vbǻ\��~�t|jn�(u����$�i��d��tB��E�@�
��k��`l��2���1����*��hD��E�{(�ڎKE�)d�i����㿣�v.�V䢖ƾ�S"����I��[��~B1~�=D5x�h ͦ���w���.��`p��"'v�bE&����RVÌ۹k��׫x<�2B듶�9��u���uT�ָ�/]R�#�j��K�cnҚ=�@���*Z���T��!��ȱH��=y�%�\cs�9��x[��\PD�� ��P�{n	C��V�*ݔ��j���C�A�o�m����8��˿������;�+�<Sʛm`�.a�f��6�:Y{X� ^a8��ߑ���S��m]9���x&��<VW�y�-f����"0��0=���e%̠�A����gI�!�=���>)�H��F,+=i�f��ޝ��m��z��O=��x�C�	����c�%�.�1+�o�KH_I���(.N�";Y�:*E��:�>��|�\|���4�Xy����$�G%S���W���i3��!]Ӊ�S_�Gy1��y��Ђ5�6bV��l�K#R:�0�p��Z8"Y���36��B��:�NZ�1x��=L۞���Iy42�N�m�R&�օ��U>�ѝ<k#�wӍܒ?x!�^��Nݯ����3����D��P|��kJ�oƼ� ��c K"*A�O���:�g��!O��J�[���+cDwp�[�oW��v5�Iu�qb�W+�w�/�u=�]��O��2�9�u*L>WK�i�0��p���m�(+J�$B��!*��v���z��AuKA͐k��Ļ���agi�:�D@����">7��gX���RC��6l��	$��Z��>��qV��o<�N�>b	P<�$'�5�{sk�p[>| ��G�Ź���� �@(���?�%�yS����m����F���c�UrJ��D$��b
�b$zzuo 0��4���(/E;�][�	��a� ,|�*���6RFz�o��	MAb���xJ�
�zf��������6Y�ҥ<�Ӥ>4��ս��0}J����o1p:����}},�[.��C
 ��E	]
/���;��M�R�m$� ��8�����|X�'�ބ�^M_�����-,���t&ӧ ��`GN�/�T�U+;�ǂ6�v������G(�����6�U=���z?'ټ�Ə�n��Ȟ��jj�X���ly:���w��,������P.�f��r<@$����sW��Cx-���_�߽�B���a�7��p*�nQB�{��c��Ol71�hK�8�䘟)˯�'z\��{�]/�kXXF�n�E�}���"���IPO����qN�ol�X�v�S($��\��Eq�L��Rh�Ov{�W��?�S���|��츦{���5�3�"{4}�[�
@��Aj���T�%*�U�9A�Z�l�(KZm���b���k���d��E�2�VXn 0{KK�;��uh�nb�2�24�v
��ݴ����K5�%8idvMӳm��R�}�ɭ�sxl��[8�x8��M�╴�\�^uUd
��<M�P���(
��a���N�P�RI��e�Zm�KDY16ɦ�X�e6�I�X_f�t}&CF��*x%�dZχ��gj���7g�
��3��&�W�-�
w
�&s$_�jF�n 쇁�ӣ��R�b�b�hZ���惾>Q;�I$���4��n��o`���!�Z9��v]:�tA9$Z��2����_�Bt�΄a%�E%�Z�pX0 �z2�=y���M/u�f�f,�'.~���zim1�K��FgnN����fY��Lz����69��0�s�2�r���>c)�����&O���j���Ed���ʄ��&mm�v�����+��e���Uew�Q�9��I7|>��&�����PP*�pF1@��[�{��$+�k�!�<�-�E��
Il�|�޽n~�ל(r<��9���*I��$6+d1/v����јi����nғ�݇��C�ۭ���V���3�.��Ԗ C��ji���Zr��@=7#^�{��iŁh"nE�R�#**l��\�|�� Sy�T���l�c��Q�љ���`n��^>��q,p���#���kM��!<�Ի�����NA�(��^+���8� ��'�R��DD!Q�U6�/%�_S�a.	�1L������Z��n乣�S�;IEWc'�J	Șߜ.ڠ�8�#W0���%�(�x�|S꼿`����)�$b����΃ڈ�"�Z(b�c�҃�K�$9����"'Z;����ɣ�:�����h��B���/�hfNpu��惢ӁHIV�q��Ӭ�/@�Ѿ���,i�K�<1�>?�[W�`�.����1��;8$Yʊ���K�2�o���h�����K��	�N7i?�s��uV���<!��˧��'�w���V=v?�72}�~c`��Ħ����畊�$��6��1�?^��#)���ْ�=�,�	7�e|-�7� @=p%l�����'ub���V�d�Th�HO#R�l1uS��q��k
�pĝ��"��$�k�ۉ��l.eb��?�f��1}"BV��ML���	s�+��� @��)���ړ��Z�1����]�z��믟7+�'�t�{N���b���3B��(���\����ShWcb�%��
)�� @�S�_c�v�|���m_������L�M�w������{�!�].� ��(���ʋ1C���� ���8�"�]�AH�C��3gC��'h��h��ݡ�!o���B��7S!sI�~�"#�fX\҅sF�g���8G�B��qY 
jmq���ʍO"�r)���m�cV����ކռ#?iH�ք(�ይ����^�ѻ�Is�oOU�Q~�3�z�h�|>5�v�,2�ƵsA��ƪ]LN~���ӝ����j�m)�x����`=m(U�( y՗�$z|P�is�V�A�e�ܾ/���-LąR'��"��򆋖\H>���9����ؒxHr����f��2,n��ʒk3����n�R�j$��u>&EN-5����0�qJaF�]�N
�QaaD@miBB1��Q�&1�|h��~m^u�˻�K_x�H֭�)H1o'��SHi��͝B�|�>p=0OE����2�5c5=U%��F]�h_��������d,���-1��B����Y��������x�o���@�-�K���,�/���O�,&O��=㩜&�:y��SÀE.��Zt�_a��(���� ����![N�x�8|���:������i~ ��\h�-a�烺P�]�����&�>����8	 Џ(f�Ϥ�"BNjl�+��Ӧ������;�|a�����,�$�"`�D6w�J���jxK��l����-N`�"JZ��z-�>�2 �����"Vt�k��tE
P9ɶ���5#�?�����&�Ǫ��	���xy*�x���%vw�qW����-ڋ4"G��;��	;�k����jis)z�%+cQ��q�����/��x�P.U$1�����g.�½*6��T�ϫ�J!�"�m�l�QB�"T��  ��b���ÉHA�^�w�=QR�ܬ��fŽ�f�;
��b�c��B�*�-�T������w�ezN	iL�?k��գ�����J��D�B�c�������C�s�������s%�;[ƀ+DF<�l(Y	�\>��Lsg��i���<�hX�.í� p�tߌ������]��>��7���Q�t��,aL[�b�����Ƈ<�	�'�@yi]Z��-ղ��j�P��Z��`��uཌྷ�z�����ۃC�B��S;��j-i�w �`�������̔킴S��qKݶ�_q��_r+�V�_�
�7��2('M�ny������=�����<��O࣯14��h�o�A��ٞ��~ =������/yCꂡ$��r�k}j ����t#X2�c�"�\��`���\D�!5��1}�'H�Ƨ�#�;)C�D�L6��0�Z��nU���	����"�{�{�NTZ#42�ᄗ4U4�F�e��ۖ���=���I�$R�PˈR�^q����mFj}tddDP �'�|4��-ҡs]Q��^����� ��q�>��4$��E���A��Wΐw����ei�5|�e���PօX���"HC��&Fe[���@��w��m��Kk�C�$��@�z�`��6�%�j���c?��x�[I#�vI8$ư��W�*n��bc��5x[������ �I+�i��}%��`����b:2Q�� kb���B?�:�1r[s�N���#���J �\��Z%;v��؂�/X`��ӆvP��h7�Zlna8��O��[#���crČz/<�F�t��.bp��ؒ:4�¯G��<Z}͍�d:'s!|6Ѱ�0�5�.*[n[
��h��#��ݪ���"���	�+�m�\�>�'#$;��W��D΅CC��n����<c�Jg,�����
P8C��$xmL��,ng�ך(���̲o= ��_5J�a���K>^�w���#Vop&���K~KA?~���š�S����Ð�ktb�6vF�r0݈	j��>h�׺W̄���r!�d#>��-k�Y�B;s���a�����vYCUf�E�1�Im��$����>e(���s{D!�`2��z)��֪R�٣EY��E�z�������밚��Cc�,��⫹��#����4M`3��(ߧsּOm�,q|�5:{$��|��	�}C��(
�!�s�7� H��(02i�������:߷�'�?`Y�J�������|
tn���^�%�Nzb�I[�:V[��Q�$���|�2+��g��xxG����7�� �	���e똞qu�`�2+��|���.�e`OyqlͲ�����9����%V��C��%�e�n�9�NE��8 �n��+g�^z�#�hj�/�Qbj����C\-0Ჟ��\�l-��Qg	�� h\�JW~.���0����!���m��đϝ�Ի��MW*x�	�a�o��b�vˬ56�΄K0R�l�+����v������؆j����{������ֵ��K<e�@�p���X�#kaQ�Ά4:�Q�=_�$z){�6~7a,�����x9lٻ��P�	�W��(^W+l&Ļ�[�.����w$;N�%��^�&���ơ_vֳn_@'�:��w�� �r�T�f.��<:Q_Z�R8p�?1���e���8o���u�L�C�^��ٮbZ�
�tU;KEgi��������Ff賩K��D���C��d$���݇�S�;�A����U���:>�3ʮ���՘�X�뱀{v��,6tŉ�wV`�u�;�A|��]���	Yh<���
�?���-qn~|�خ��b?���n���Ӽ�
�wb��3����8�ӱɬ����,��
ۘ������"���z�Ów��a���p��P{�f/T1�rf*�	L��19��b"т�vH��UJIR��v�ѥ���sE׳�/�K��#ܱ�KV��cK�2�����8�l@U,�Å��(���sL#�MH�<���Gխp`^�%��YxD� ���[:�h��y}��d����T��zWP�*����C�Hf��7�ᐘdF)2T������j3.��[��Ӌ�g�#���ɗ�M[d�^M9�m���r�:����d_.Rp*.�9}��hqrY"Vm� B7��ǵ2#8�]5����J��ac͉��|	�O�:��^w�u&�J�	^ʝ �<�+�.��e[k�J�yq}��W*B�F���Y�D��er`����m=K�}v�8��c:��m��RQ�mv�U�3J�7���s����bFE0�u�ּ���槾*zsT�Xw���TT�;ۊC��3m}��J�N�0c="��_��<��������?h��N���fCa��_�#Hir�r<y?����g�|`�5�%�[���/u!6�/AZ�G���:y��l���pp�8X8�҄�ؚ�*���!���C� ��jN��2'q���b'�b��*Bk@�����&��)�d�LZ�Ը��Y8�*��Q*�{�%N��X����xp�8k6s7�C#@�p�8(�4���P����H��Q�ʐ�Q���̱��/q�����P=SI��?�W�ۑ1S䝪w�6f0lD�W��>��v��^8��V�"Lo ���|dּ�[���6��Y��\�))���)7��n��Y���9@:���\[���y���۪1���[���ɗP���,�Ϭ!ip�qi���y}3g��t�����0�ˊ5d^��zL�{	ceZ��6nAXFn���чlR�y- c'�|�dDm�O��2�gՋ2Z?�s��'������3�0V��{�cf����Ù�1�O�E>�ċ�����
��*64"D�,�D�Ҟi�tA�rT�r7`|Z���w�!��@�SLr��]H�$FD���z#��3��(�Φ	)�6�M�+ڔ�1Z���ѷ�LC<���ѷRxl�MEĉ��