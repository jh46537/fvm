��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0�����
����'a���en�,�=y��~{��i�#�sS�Z�àx�WW�Bg������𓇴r�b�ex�Wv�c���V[�4+9o]��\�S�������_���]U��J��]2c���L��<e�@�&���jX�3r|~�SrOa�{NR^����y�R�ΏD�|����m�'�m@�q��S��Ƣ,(�jݎ�4��>X���w�j2�)M��&�wU�=�a�;�k����K���b���ʎ�\������E�\��,D�`�������A\]��J�o�A�����^�.�c�mC5�h�9����N�
�.�C�!�V ˘�٬.#�]�	ޔ.�⏩� j4pTMt��U�uW#�����3��ɐAw����/5���C�اDt�����e���#�h�e�W��QyG	��,ct��{6k-���w�Y&=pK]kS�g7�̝WJ� �
�Y�X�K���L �n��ӡoQU�Iy���r���o2k�aYDx���v~WX������+��xe|F\u�R��0?ked�1G���U��'i��Q8{���=X��c�H����Մ�t>�"��ĵPD,H"ʞ�q�m��X	6f�u�����
0�Bl=U{B�1{��!<��·U>�4-6�8J���0A��L8G/���\f��W������
1��f �X>�"�<�M�x�1J6
�B�?�1
�H�=�.q��|������3DB�[G�'0�=w�p|J[	*�F�zz�aV�B���d��PWpm��O�l܍��6�_B3�/�|I:��(n𣴋R� 6��H,�s�"��d\���S��������(���hR0�ip���b׋Mf���r�e¼c�b�ˆ��`*��,aQJdk=���I��j_4�E�!���na��Ҽr`�p�&g�,7\AwqJS�V���E��&E�� ̄��l{Ҫ���2���Q�u��u�8��¶�U2m�}�5� �wR�T��q�ڟT�Q��ݎ������Os�n��j��������څ�ޮEq�� h�3��X�е�n������H�^v6�6)	g!l�~�i�!�b%&*���3B�����?`{�i����n��3 à��^�L�섂��*���@W}a�WVx������'���j�PZ"I:c�Rwr8YDX*"y7P�T>ok��(�j���[D�G�~��	�hL ���#������k(�:u8Qz�[�xN\���3�0�����O,E�����b��Jx������BWSXP�a��={�$�44��)Wu��E�X���!�������Y|�=s=�WL�	K3���|�ZXjs��:�3�MS��{��lʍկ_��6�I��H�].����l�t��+�� g�zG|DT��^m$xB/�~���	�2��r>��������2��'ta�v����v�uu'�Si+��n(�jԭȒ�-)����6�_�2���mB8(��o qX�`��M ;�]�'9"��eF ��C����̓�!3����xU2��z�["qu.a)C=�gH��Ѫ��2AvD��0挾1��5#m��6`E>���+�	��,Ք��� g����\@6����	��è֞2��ONԣ�c3���y�5�^@��f;��8�D�>̎!�#�b�(�Jlp�%�.��e���Qw[U�0�4a(��D�,�3��HW����ٓ�y�n�Z0���w����C��'�<(.����M<�.��^�xثr��B��T������g���/z���'� ����1��=�b#}��q|�@������ ?��	���%���A�<�#3��)NcT�h6���Y ��b)��,GD}�Z��i��*^>J��P�8�TH�ʫ�'>�&%'�����BT��쓭i���V:�P��O�;���F�fJ]Wi0U��È&�j�4�^��g��:i������;��s)������?Ut�!:ܭ��%L�sI�kls�14�N�L�g����N��|E���H�en]�K�:��_��Hݔ��R�������:i��.���$.�.⚸>L��%��L�O�"ѿ�����wʹ��eBq�� �݈]1L~���?Sq6V��o-4SRW{��ߧR�Xwq=p^���lܨ|�K"����M��wHq��KdS�=��r	Y�t���.MZo�9C�a)��}/������;�g8���m�R\�)�!�3<O{g΀��`җ�~�õ &����O��������Z���6s}�fCS5`���|l��^�G~B���u��[���gJ?Mc^�@�5/�11#����R����ec�4�>��]7����iKN`[�q�Y0W2�0%Xஉtz�{���|�/1��;�7���(�R���U�r[�����tB���)$z�S��llRi�1�����}���'�\R�f~^n��'2��JM�(UP�Ec�E.o��I�����%ٜԦu��e
�s`��ɉ�F�k4r����Y�y{ش�=��y�����+v�4���J��T)�5��r�����S)���p"U���ߐ�#�E=\|�+)��=��Y���#� G6r��ކ`���*��ѫ�궡p��V�>�N����}����Ψw��:�x���1dJ�H��`�қ/�i��z�	�lI	Hc�P�B��v+�t���@G�p�8�C�HJ�s�7�+~���*@���^�Z�*%�"a{P2��R9��}n|���v�$%ü�)�� ��?�E�.l������"�������uB��6e��N��\m�9��2⸘o7AT�,�6��2��J�-N�Ōv*[��B��5�C閼:~�i�	ΨϞ��y��2�x�Hz��a�r*��j>L��+�]@
]�\L�D��?:ظ{�ߢ����bS�j�,i��:�.i��Y¡ۖo�|�r�9>M:-���_���j�/j(E��a��q���]�^���h0���$�z�'��%j"�SI��ȳɥ�(b�cA`���.�wH9T1���	]0��{ȆZOU�k�Q;|Gh�E��>�ɨ:e���4!�Q��@D�<D���l�+���b����t F��]�������6�eÁ@J>c��<|���������)X�̄t�f.eI�]9�t`��W�}�-]i��R����p��j^N���B�jÏ����N���Ln�h:��/�1%��V���1���݂V���8�_%!�y�͙�g�F P��0����0v|[&��*������a��	��� #g��]6-��[��^GE�>���4o~�n)�řf�Kk |e
Mw�s�B8
��,�gY#����K�|�@�k�!����9��f��Gj:b3o��i���v�0ۼ<�� �B�7�p=�B�ġ��w;H`F��ؑ�*ok�OJ�Y{e[��'�yƠ�ҝL�&N��rc�	����.�G�LAF��ί�9йL���|�o�����rJݣ�|7�"u�*��G�����A���5��u���q�����)�Iѕ�(�?��.��sҀs��'g�s:c�tJ��|B[҄����'�]Nfyj�ڽ�^Y��mm%Y�_u�9C~�W{E�g�P�5Y'^�E�r	��]�eD[x%Ā6F]x>b���.,�B�X�L��S0=���x��M��Dgd?� ��5xv�08O�����+>K���C���*H�r$+h����yk��*���=�Ij���&�
?!D�B��؁�L������k4r�,��8���Rt�B-cA�+��pf���n��ŗݑs,�e'��ԝ���^X��´��:��}�W�K��ˊC���)���ƾ~�ɰ{9d �1��!��D�%��S(ȗ�)|�h`��1F��h�-�̕�lLX�_v�����#��T�YO�A����h�"�Uy����Ir�"���)�Y�O��zC� �і�IA	S��jIoPa6]� >u�أ�^��R�Q��:7����� (�W0Z@���b��C'F�/tW2��o1<��N� ��95j@�Z!��������@/�9�8)��#�g�b�W�B@��]���zJ���%0&�*x\�R:��8��	O^s!�}�|4p3��6`�K�y��ox ��ѻ]�g��3��Ἄ��}Q��:a�aD��P���d\����\����}�p���W'%���A��15�rp�g�E�P重�w���Y?ݲl��������[��h����7�*:a_Ǻ�>��X�2�� u(n�-���i����=��{z]@�-�N�����A�J$Y����:������䡓�����Q��*aLj���R8����"6(E�۳���/Q�z�˅�L��U�X�jÁϒ"��C�H�n�[;{�_������b	ݓ��:�̔@B�G�	�pt�ٳ)�