��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""���᤬����[���%rl�ϓ�6\e��b��o�)�֬��+/!�ܒ�P�m��)����<��k41�Z/�T-^F���j�κ�D1�3����9�a��B��ӧSo�aj�Bq��G�BpG���I*_����)���3����
����cAOj?v�S�`�$�ۣ߀d~�Tz&T��O׎�C��K?Ͷ_x������%M}@ٵ�	���[��Н+�5�:��~�+��DZ#ޘ��=���E��}t[$���o�`�%�d&�|�5�,�=��N��7��}wu((���js�`P�WV�>{;���.��ܴ[����u/eDɵ�"Vex�K�x�3���-͚�fN?���?����������QR,8�y@�����]=÷z�Y;!I�13���\~�h�YWAq�/J��,�^0����Ů�΂���n�UW���}D���	�K�<0q�{��ksw��E>�����0���Nz�K���Ϩqk��&8uj����aDR�|,����j����g�>��4Q�I�T�^mC��q�x���]�Ϸs�RK[8g�,�xi��ʶ��i[�Q��WU���<�.�z�<�g �:$�]V:,�KM��mq��5;��V��p�,�K�#�{��O�N�_�S㍞��F�q��'���IҨ���?�:o����xg���ѻߛ����{�u\��N��C*!�Ux�Wi*)r���E�>��UA�d>f��]��&�Q�
eG;R5hj=w��xZx?�<���0��าufR�&���Ytd�Zʤ��YI�[�c�>��t!!��)�%��ǅ��rWK����A��Q���H,�1B_��Am�*�h�m�2,�I�E��:�.�:e��7�u��5]Z�G6m�-�S��I��`�������8yi��J��a���������V�%��Ec<ܱ[���Ee兣��V$y�d��Iq�����вi}��D?�9&��{/OAWU���xt6ި�bXs������&��m$�bpX�16SZ,��M�?ԧʽǝ��*�kށ���������釆�?�7��g?A-3���BA�Е�mQ<��n%|=(�$b{S6h�ī�Q-�i����v��6�OOej�$K�_��N��w�@<^�Q{\�#�����	4�1����\&$�� 7Q�|$11�@ltxV1�N�:d�m�y=,�Yq��VY�J����9�O�������;n���O��� ���,W��������w��/�3K��&��9�8Yܙ�>�=bCJ1a����p��[Ƚ�
��Ŷ�:^�I���E���;�8>�Ng��7͋�RK�Hp\0P�Y��?-����ϗvW����Ώ��I�G���YF� �2Xd#���4�Znt.mO���:mzq���R����k�<K	�,�@1U_r>Hiv�v4��E^(o'��t��g��zc�+�^{b�a<ޝ�&�6��I_%;e��0�ʲJY��͙�)��MF��Dڱ&yI���;�#. x4S*+��S�cбu0��&v�����f�Fq��������`ƽ����<��de����q]=�v}-��H�'�۞K=A*�v4�J{X��Dd=!���$܁��`Ep��vK�Q�l������uQ�^H�F�c�a��T���X����!}@m�����:&[<MU)3p���ց����3�����JL�Y'	#�M�~qY�'UZO#3��*��IB�^$�Lu��uq�p���K>���ٵ�rd�F�d��\2E7(���T�c�!������j��(E6� ���ʌ�4h�,ԑeL��o>6����>��D^��񶻼��#�K�꤇�˨B�_�5�f����ż��ޣ%9�ݘ�6�u0��Y-x���u�`�*G��pS��@��}�uR�$��V8�w��SC���U�͂P,D�=]�&�_q����TQTzD�t/{�؅d]�����g ����y�)��ŰeO jxu�� Y@�s�7�T���s�M�ؘ�uȱ��w\�S�L������p8�ځ�����%D �(�����>E��G���&I�� ��y�t�7�Kqe����liJ��>��i/0���ѱ ��%�b��=W��ׯ�r�M�dyB��PF�l>�_F%�&u>AK�%�@�v�i�sK��r�V�1D���n�9�B�)�y����(a.��3�U�|��>?��Tyc|��,�s��sk�$̀��EZc��3Y{�In=ܬ�c3%�橉xt&(��b���2uί������r����/?���% V�{gN�#� ՜�:x�m�?���]�Cޘ����9lJ[x��՝��������3~��h��i�5��z�f�J<��w�*xpeBO��f?Z������-pӉn�]Č��Y�R�x>�a�hAM�y�*�+6�
���d��P��8dh'�Q}nB�����^&�΃������@X?���i�h�ѝq	�)A�;��_�8�6�gA��M��J�Z��t�G�+�_��ʵ[�ں��?C����$ء�@����$N��2�P�.g��`R�<G ���EΠY��4hs���î���ҤK
#�c��C�
�EJ]��$L(�Af3	Ӯ(���큣��;+M�ݪ:G.(��gU���6�y����K���e���bU���#"�h�z�j����o��~U�Rϋ�7��K�<�%���0�9J���\3UTL��8�	���U�6؛���&�!�Z!O�=������k�=8�͗���x����^^����^gr���]���D����}Zn^S���QB9q��!=�N�hR˙�VJߌF�z�s/��l�Z�.#V��w@5?@��d�s��Z ���:�8�!]�|����N��L�q+��y�9>�~g�ӎsz5V�?�jm�Or z���+� �/�gC�MXH�M�i�Q�0'�#z��Z❳�#���L��I�')4�Q��t�,<LGT�wm�0��=�u��l^2�f�������I��_��ft��JN�g�Eɽj��m����߇��cF9��c�h���"����B�*1Шc�$�����6��Cy$f��-O���ߜ*im��Y 
�>OֹQ
�bZp�� 4��ۜn�L���v�?l�{��ykq|%f���l�H_~�]�1�T���N5YKݕ�^-bcq��{����ٺ�7v}_�#	��x"���Tv!1�o�גz\W\d�%\���C�*M���������(�&ȥ��-WB7�QF�١xg�VO�$����hl�0�K�F�ol_$ш`μL���XX���|��*jQ�ÕWVtc��'�K��W�q]?�F���A懨�MZ���:;�W-�J&,ud`�� �G�Z���ȷ~��h�:� 0�N�}¼갎Q�L�S� 
E@x[w̏3�5/��q6}P챷+'�ئ㟫�,]i��Tx�s4�d���<?r���b�R��݁ێ��z�~sσ��)�F�w3X˳����^�t���ʔ�"�D?(_�R�M*��ΒNr�	�^W2�c��6'a�楷����GV��'�Yt�YoFutIG�r۳q�^2���[�Z�tϝ��J���� I���/���E�6�ك�/v#Y��܆k00*���g�5-q�4�K`�K0�I�v�v�/���
�F�bb���*�(0Z~���оo�!�g���;��Q�?�AfA5,�5�tZ`�5x3�r��L�T6;x��������۱nt>�H��6�;�X�U��i;�n'��J�8ɳ3 ����	����,(<�Rg�!���KԬ��kZ�!ؤ:7�C`���T!|�xʞ,O�ĉ��4��5�eRǚuq����I7r�a	w��J�=~�8��>IKֲO���UE�v0�>��|�ÖƭO[1B^-�\-]�Ӛ�I9��,�'�V.�ep��;;��H��/GI��-��k���8'�@[�N^�]t&�2��A���������`-��I�d��O�/k�ҟ�����Ǝ1��O[��oV�:����N)X��E�T���@����G�9�&���0��b������>�ԏ�avf���#��ƅ�������qaɍ|>�?�A|��W(r��ʠ��^��:*m+�Rf�9�z��@Э�i$�p��"qr:d4RAU�)Vr'z��*4�Nj��EE��\��p��%����۠|oI���2[���@��G�VB1(m:#�X�"��*f*\�2i�����Z@����AIj�IQ�4����H����S�=�$}��e���g0���ݗ�!o�d�g2�@Q9#��p$ �	��z�5y�~ߌ_Ӽ)�~��܌�$��E`gW�B��_8���EDgv�9�IN�5�8�N�4�x�X�3��;��HA��m q�(�40�S��.�ٶA��(�^}Y"A���j܋�	�bm�b���S��k���sQr��8]ԡ�l�@��_G��z��R��
�����O���F�L��'1'"��V�V���)I�]�� 
H��φ
ze�DA��3�(�mW����x;�p�!�����>e��G�!8�o�FS_�q��0�{���(�	%�ak{W���P������K�h����qɇTQ{Uv�_�^pve�N����JL����Z�AF��ܥ�4�jr�ޞ~��u���vi�r~�Z.��M��s\��Qe�v-���E�-���Ib��J�<�3�*���K�{��r8i�%C����;�Jw�p鎕�&��/!n��ٜ��'����!�*�{[g:�p)O�$0i�r���@�m"kw�M{��z-��\���"'��#��p�0��p��?g�䜍Iz�u�C(B��dWv칾=,���h!:����k��L�����Ĥe��l�%�]Ҏ���KM�1��o���K�/޵����P/���������J����o�Řtlu���6|��$���M5��0A���ɲ�ʦ|͟�����������*��}��AQ(&�SG���^�(�����xT8f{��6���4��g�=��i��*�)�Ű)v�ׅU��$�?#衎�Z��1�0�2�S�,���tʐ�N�<�1�\0�[R��uμ���l����\>d����w�Cᦶ�T�s�>�[�?�}�S��� k�pK:
?�}i���$��7O{���G~�/�#4��F�@�"F�@JG���/
�$XOid�F_�H�\G�Ē}����D��9�n>��ۻr�dyȌ.�7�GS:Z�����;�֡���3\ƨ���U8M�s�W����o�@�k�������ؙ?|^3�`0��Aº�����Rom.�Ħ��k�A������~���G�l���=Q>��HF�����_�3�L|@�7�=�6�3�޿����Ɨ��Q`�CP-#s�b��CQ-�)�XaV~TcJ��׮�[t��Mg("���Ӫw�<XH�Tyl��`�/Q;�l�y2�X}��>:b�I��pf&ϴ���B��VDX��u;�����cՙ�j�Hq'zc��-����2h+�n�#��<Ű�'��T��T��kW]r��)n�*|;'�Ұ����?u8g��^+�EF�FC���w�צ�9s���l�8D��$�#�Q�1�7�`�!�|������R��鐨���T�b2��9�!��@�i_!��\�&Eq��4�^�m��B�L����:���-a��4�N��ǾS�����g�	�E�y�Б��C�2���^h�a�%ڼ|��[k�6��Sò&�$b-EΖ:�AQ,:j�g�@�AK�3���������.P��%�ZK=S{�*.�n��G=����i��L<6��q�L[4�����Ґ)�A�Rț�ax*?����f��"�E�oS� �4&��A|$��q,�-���� �bÃ8�Q}8�E���#�T HY��3N�`1v�}�ͣ�/�I�)�޼}+�)��v<hLW�G4�0�ˢ�=n3�)��m���{�2�׫�F�|��d��p�w����d��<c�b��>S[P�E!��,�Ӳ�>� +pq!��
�(������J�Q�"�uW�捓7U2u��^���L��p%SN���A^�8�
�V6Be_�O�Tl�ᗶ/o݌��ev�_�׋�b��y1@L��#�h?$�����I���{���p����t�[����J%B��V� �=�5v��gmt݋�ȵ%6���΋�'��^�TS�9�Ee�ŎF�Z�<E>�e(�,z�QIH��O�/�b�E��ƈ����b?�wN��A~Fs�p"aXh� 6�ݞia��%*���$�����N.pҨ��X�y}�������jwE�m^yl��������,	1)S�/,��/#jagR|���m�`'��_��C��[ٓ��gj��t���G:��*/��]���t�*�)��h:�����̈́WeSd1���?{�ӯ���Т��J�� �!�>/M'5��J|P�!�W�t�h�B���3�TJn@&_r�AHda�K6��G��LBz��5P�& 4좘i~�6�1D}&�}�?MD	`�aY����6��ҧ�����9.���[u���`���җ5����xe	h�H�f^�)F�{z����s���I9����3�q��c���rx��_�j)Q��$'W%�s�8�t�<�3'�	�:
�� ���7���\��	�eKκ�~�(�����.����p��[ AM��� )��V/6�;�~�Q��n��TlT���$o�,��'�J�UP?a�<⒎�I�k���J@Pi���~�t���'�;y��ϋl���'w�a+=Z�t�Xf�|��\��Ov�f��a�����Z��4��v_�~��N��%�؇X��_���� H�����hCxr��T�Dt56d�R??���y�Z�	׿ >w�����kQ���6����v�ȏW$�ňrΤb�56�P�_�)_{}rQ�a$Sx���JFj������s톴h�\o�bOW�׷�*��1ƙ��3`�Hx�t(���SSᓻ�|���
*��������H�7��b�	�JL|��d��v��(�_������XQd~������1叜}�X�,�J�(Q���~3����5`�m�Ev]@D�#6?i��I|6q+.��Wn����6�~=��4�3�e���]{iG��Q;�=M��I���Ar��.�A�O�pNr��Jż��J}ٞ�s	u��d�. ��*�mA��ޯQ�9׻mv�K���n@f���n���6E�99��	�Q�n� �f}��;1ψc�s�f�k���r�.�
_M
�0=�o�;Iq9.��ȕ�Jlr�h�M(P���@���E�����9��mLͯ#��
��8k%�t�V����vb׸C)���B
�7��Y�ϩkA�@�����O ���e߈�JjG�Q�]���_�v�A�YS69�X�vM�#lJ����;�vv�P6".ߺ�ſ��������~��}HSXd��|�$�-AK͓<y��ܒQ�E��}���}�r������2�[���$��p.
BH����*�#��F9\�y���̩��O�5���/eĉ����
l�Z�+S0E�dH��z-}C��H !��Q�Rf�x�F�rQ	O����Q[v��� �^�
G�s�w�]�"�+���t,䙩F�@�a� ���E�c]V��C��3ŁˌC\��dP-��#���J��[�p������֫��*HF���jī�T��?��^F���(���7��жp�x��u��ĩ4�d��\-.�\�����������}��A%#172�r�Z�.:�T�66T�>���b�R��k�e�L��Q8N�O��t̪GJ�)���35/s����C@C��ѳ�Ԁ��Y�����J�c���l�Ӭ]��$�_<MAé� ��߄=?��;Z��(~�(��
iuY�Զ�\ IߚĬ���!��%Ƥ�����o��,�%�[��׊�W�a�1��T�������@ÀQ]���Z�u%V���1x*�H�!um�~7�a"QQ�ե���SQ'�C�5��_:�2
��^�:�ziȳL!.Jn �*��[�I���*���p|�j�P����ea��ְ]��ᶤ�wLK�uؽgup��jڂ����Sz�8�?�p�ӭ�)�~U5�}���Tɟ��B��sB��� w��z(��_���wΠ;}Y�x[�m�::X&�&�J66�!�u������>��9BI	Az���J����Qwʔ����o���'t�]���A���]Y�#�z���^��M(F�vvG`��t˞m���҃����ղM�f,!�� TgشR���o������'/ҿ3%��#���
��I��i��yE V�lHo�N4��:��y�ƃ��Tl�k�Hv]Of�1�m�����W��F-J�mPi�߷��9�hi�q���a6�Z���'�=_ӊB��[����A5$ﵰ��8��s1,�wm,_r�c�G����(�sw=���,lgI��sP�.a��j���J����_�9vP�O�=��%n��� /|�4ʜ
����Bt�P1%��n$K�D�)�s�G����9���{Z� "b/+��~�1c�(�^����QF�	0�9ҝQ$�t�8���T��d���^rU|��"T�8��8:�b;@ꕑ�$�Z�/m�.���/+}�$�����ut��2�.D1�/��]�N8O��Z�x�����O'��؃ǝ;a��3�M���G$�ڐ7$�6m!E�����!�W��;�y�b���c������r��R��>��AQ���@����Hn����L8�g�?B��b-Ŕ1N��R5&��e�W�`��c{��h{���	�'/�$d�lB�+[ �A��ꥺЃ[�<��j���À�EU���4iIsu}��yH�5�̎.��[����(ըڌ8�S�&V�;��`2ҫ�A�a�:��(^{)�o��iG�k6e���$��)�%8I�3��؊�:1�K,_/�K���]3��g��r�pO�7��[D'uI�A�
�Ü#��?��z���Y�	�O���ǹ;2��?�ɀ�\����,3���{rhA�X!�v��u�S��)����q�������ߞ3�/�B�j��Vm�(���y��=}�Si ����'�l�E����\h0ow1��&p;�׶i��N�}�`rǜy���00\=�2FP�&��\<�t9�"Ie��}n|�s�r詀-�"��խ�s��	��=٠�%ҧ��#��`;Da��eS�[�`L_|��%__�*�n��rl	���KF��p�?����8�8LjD���`�.=��@`+��p-8�Kь��h��$�8N,?��M�ܯ�a��9�
���� �,R�� ���Lz�N*p��\q��$1V�F���nI��@�F�����	�r��$�ǔ�*�ټoY��; �Ĺ�j���P�cg�qi�#��)���3�ܖ�۝a�%�?&�/\�tb)��%$��f�3�D-%�@UQfɔ��Ce.w��l���a�*,�[�`i1���7�����iT�*�	y��lG�`��M�x��!BF���8�#�m��v�k�~$�w�9�i�ϓ��4��^�|'�o���E ��Et�&q�G!��G�[�:�͒��q�ǰ�������k�NEm%��l0�h�t#��'��������v2��q���j���H��tu���{8��0g4x�Ef��G�����b���b} ŒQ[y1]rd,tF<�:˽��ԭ�4�%�����+�;;���
X��"�����NE �>���op�8~�K�Gbϙl������t.A���<�)]П��K��c{yL���q
F� A8�NSv%tK��G����$I�p �����-@�] V&��Z����"
��k���{���N-�܋�R�0#`��w��<y�'�9N��M0�.��5�2�6㥇��D��{8�=�����<�|��ܿA���07u����^��L�7�U�C��p�2��N��k�����|��"�a{\�Kami�_��6�_���*�yg�Y��>����f���%�@�c#뿖��<�<�w|oR↜{;ct�0n��33Y@C��b;5��.O6�z�Q�)5���C�.�HDBV�A���S�)�;�u�Ů+���Vv�ڧ$�Q@>�/���X���Z=;��%p��/;�|�\K���AyF���k�ȱfez��x�D8nW���c��sy,r�1!�S����g�Ŧ[U�9h����s��,�u��U-�,7:2O�V֑M�:
t�Y�� B�g-?j ^9a��`���ڭ���q������m�5���\�0|%���E�HD�ds4�\��3�H#	�i�pw���Zb����Ū��<� (�p���I�i'َ����m��у�I���Sr�Q���fƃ�@}��b64�O�-��|I��*b<5�k��,m9Շ�%����#��{��:�j�(;F�Cβ�`Șp�ď.v]t�3Ġٍ�a���	���[�?�p�V�2�T�6�!MQ��1sӮ{f�X1&	����lg\zy��+��3��sd;��]rU΄{޽�w�,��{=�`|���'�P��b�ĩ���&�������p��1(��=z}E\"%.]X���c�c/�LP�&�2�Fp����VI�^lAt�=��,-����L_�%��}J�]�0�F���n�Hj%�R�o*(7�oFX�e�K��nP�_���������{���Y/�)EdX]��Ca�g�v�HA�lh���i`$�of���3L�k;��0����DvEB�oP�6h#Π��[��׮Mo��V����y�a��e�~[�D@b���8�&U��K���Abnd��_�L�˽l4!?�yYe�ߎ��*yo/�kzc����Q�+���)�w�2�JS��izl�xv&��!B~*J��TS)����EmYx�a��z�c�B�m��9MP���n����9I\�g;s.<�������Oe��k�5t���_�`�ʑ�v }~1�J�T�M_;uR����y͒(5��YޱlR��i��Q!�2�1��2�}�*XǛ�5aܴ�G�:��\��2o4׳6���TC:}��1��m�[5�y3N�}M��v���/d��/ȑ��|�]��a`����9��Ò��`�!m��H &ڶ���i�{u�ڮ�j�_��8�P!;�9�u);P�IU�	� �