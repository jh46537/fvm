// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:36 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PF5+FVNJeSk6D0nNJiKrWp9cv/04r8LuHDoOLsKQoo0vbyrU7Ls0uuOeiqh5qM8x
JAF/kSbcLRjwVX4uJ4cT9RtFP3NQZfvKkiL4jCVeYlr6UXAzx9+2cdO264LiBVMe
BMVzsZpA51VtKnUIgJltbdeh4YeR2QxGfQ0NV12OG+4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9600)
MoylX+NacVxVm7tUJICNNNRs1UXmgE0LAs0HkpjFUHhdBppyJGkMPvvsk+1e7q2U
T6PEJcS73FegHGGM6TPp8HoM4sa+s2lqA76RxU3N5scg1+fNEJ4oTxuk3DmPIwno
4IE0fMPjIdQ/+qSNMMLIK1uUpiY7LWJYpnqqP4iuhY60Wm9mhpc6ueKAOUl+/DIG
Gjt6178MW/ynmKlpm1wxpy6x+u8NYliXdk1dBUMIXVKfGOoRn3wrz4HHmJos5WIi
cU5hyW7yOUQ9H9FJESCM9pUfqTA73ytaMlEr6EOLYVpNFpx9tbtrxkeiRlPybWy2
5ZGYVz9bOoQg/yVfbCuOAdqfIj1u1oAs+ry2Fp3xo+1V90wbojDBJNk5S2Oq1AYh
8i1QHKaZu5RlSyqCSyg3fcB9gzvx787idi6egBBhKytb51m7tWaVrqtVgzkNZYqZ
fyaZ9clCW9nL7wfRVZCsrROoMRnXziIOkG0mEXrIO/7eSIs4K/sjc2lm9eALIpkz
42FA2NVYIQwsEyZM+uqHSxngVb5HYsMjazzrpsG+oh0703hwai5IDR7S0YVnVZl3
5GU31Y2qMjLEuI6Yq73ZdewnNA857mW/929krv+EizAVaf89bKiyoqY7veJGWtys
dqhPM1NadH3b892NDDNwmdfow8bRGhi3TUsvhvpT01BgGQUrWpROwWbFCP/UaVuo
zT0f0ZoS658r+BHGP71m866bNWjuKjaJnj0+CYWKgiphWglFaAqoQ/9tIpjJFlMl
AKlFJ9JmRIwCg0i6+r5ATg1tgDNH0aeDWnERkur7ls93y/u8ecxR5otWDyxIkrWL
5qAdH6vKpomOhGGM37M8B6sW8cNd73yAadVAGCVSlz7Gncs+Eoo7WdkYzif4G4Fb
6pFZoTSSDoPWUi1PhH76R/gwtr4rJ1jmCbOsUQRBnob51cbYFRE7sNQeo4icefs0
JX7+6t3DyxaflJP1KKj9E9Ztj3rxa5qSm6b+6ZsL4TqDfnrT0wUMspfF9zjcAim8
ZXCWu7zpgVeFcEtaO1H4/W7BmvHpOuiMbwU1niIx0gkD61KXkMEgEfkYYsSUgkd6
wfqSdmLJiChMtCfrQ0tAKXn2TQeMZcr86pheRtFr2Ti3ogHt3OjQVfephgp4sUP1
8inseQ1H2Cb+MZ2iD/Y9JoO0CSlvn5xWZuRlv1uBBijydV2292cNtQYlpbZHcT7G
aFWvJmG2pbMkjnqig5Fpb+UfSPTVevBDEkuo/f8unII5lHKmZTdmw18hM6GQhfBH
c3QEoFOllJLKkuwFILd7HwsUM8b5EJ+ocKGEWogdwWqeb2niu6L0ZCsyKZLTIPyv
exKB437FXnFUhocdm4ucOm+r9yvLDmt2nMxMwqJk7mNMVkgPOJguFFxk/gGPBGdE
hSGhRA9bTYJ7cfjJC/8tjxe+Q92fj3IQKZFM16pHKyBJuLhybzYVIAOnlXIBDZqk
8LWy8A8locn6jAAitDnX8B425VANpwt1g3/DC6SbjQO2/2d9YsUAb5LRnImut6JC
DBUOl2TrCglyS3+jQn+GjGxL6OiQjsMiXbnohkAxSz1Cn1ir/F/+cxk1s6NPo0pc
NfuKWNjsfb8Rz2DatJfVnQaS+Te5BGiiuxwpnFPI8Jgonkf/R7GdI4OV0I2ejR5d
WaH4fBHLzHt44OQGziyUNO8M1xW2iyGlQSg+QoHEag1/isyvrHB/XrYSXIrgKYQK
VIv07MIa/x9T6voaQsvffQoG7aSGEtVJInNExuaQAqQd+xFNz0CqsM2n5hdUFhO3
ww5Na17F6vd3xqQ/jT/AXPVVq+ItsI3D2jlyw32H8lr9Bh2rcO2/LkBhdMhDuN5f
SKKVsE9pTHW7WoCS0wSqlRtxGB5D87vrSHhVrtv1iUh3yN/sC9ZznBt/GZLUU/+I
3DnIWxS1NeXPezgX1cRRaLptFMJRiGenGgIT2kUW/DViCf1kotmAVPZg61IZF9Vx
C8u+mf5fpO9DPZcSanumTVaG6NKas3xeUVTxCf7tLjFfST55qRxwCvmWLG03Ir77
hqT3si7tXAZqQhkBd4SbC+tIS+QrveEzT2knV4RKJGeCNFcK4XiEYenw4FBVjiQp
tYVmB+fNU5WU2qsxGyg0K1x7o6SBcExncFYWfn0/TArOOTmrYyIeVqByL+oQrAX5
18Cynw7T7PoRdKxCwpagx8GAoEBHVtZgY7tkGGJZYc+3AKwBSNWiKC0YQGqpu/EF
F2hcCbM5V6GahlgeNrDvro5O/U+1nbd2lUZg5jvA75qWXcPiKLedOUDW/zMCHoJq
NNeDPCA2x7SNkoSh3Oe8Uw4U1cuyQg/s4KJWlCSxujVxguFU00DKTabpi4LUPQ0q
/CN2U0ZZGQey8O2KJLapGA+KhGmw1qqB4lzcgoaAacC80GR8rpFitcPv6QZWg+Ox
Rx1xG8cyZvAkee3GP1rAwL33kCtUEwzj2loKaG5wHVgz3WUv/RI0n7AvcA4nT7cq
rq+8VZQOnEZ2LuJaI+QYxdDw1lhVXlBboIEMvgPcCOltP4JcXh9M9U8QgtW8zKnF
wMETnFy7D/hlom2E08ca+714Gt4PEVVW1q5Z3wyTx5EgcT713beozPc4//H+pyhz
gquQZRP+Yr4dzBmec7i2sNKpxiZbHmyujfw9UD1F7MPQ2QXq9ZINayECP5MXpUW4
ELW+PzDQKCDfUsr9iEkgyMVtBPOANdNXx2daO8EovdyUGPOOIgclytHFCe9nsiY+
5nhpXLIvbaysb9ldoI7jCM+7NIkVcLqvbtbZZRTSUvbGLZlwZesjy+ILQIZRhY8a
zTeTJ/jxPGRYTXLkGnb/V1qa5RCpuWBN/1fbuVab5tXdOIWN7vQV6IDZJYBMdSsc
1PgLzg8Od4XmVoRVaXXIOHcKPN1y3T4mzG1VJNi6ZiOqxjI7g+lO475WCptrRciU
+cwNtz8W2LE0lJJO5gWIpHszC70eHmor9lo7e0Q+9L4zMBTRL4iQnfo7t+MgIePe
8nksUN9e4/+ATiVn/p0SHxB+NhRu55QqPhzm7OfXorfkJlWAib/45S59JtqyV5xT
OAg/cwxHn/7z7LelUu8RTkqGtJ+6jRzYzZSZuKxTkKst7XtQCzAIOIWcb8JSQFAr
7jqhqlxUJYpedwA9/cZ7TkwcIloL0NWFnZJ4bS3rXEeXqv/sRj+lVzPuWxTXqIiv
EhOkIV868KZMamgcAaysjFV7c+WQ6I3cRHdTZJyyG2Bs7pB6peXlzTsnrgtpmToq
SwKyvLs+PadFt2WD/P4g1RS20g2tJpdWiPC+IgYvP1eX7Ut9hr4GXp8tRCt5AZxR
57AAoJE8UTqflSU1AUNhQomLwAh/yNIepW6Us5/nWWCN6NKyiPdh/lby8s6Kvqbn
GUU2R1qPtBFPDQq+u7lNpEC62vNf5AWQsPdGOBqOL0r/ZSy3UYViRuewNM1823Gp
WHQaIpWowVmeU3cqAWFpGMeLWze9TZe14++UM/RmPCOmmt9/cxV6V0knaXncS70n
Cwbp+1LktZRL2MPGGS9X1sQIUt47ynA2Ob0PLvtAtQuK69fL0wCqMQM1LgK5Bp+E
6CucUb/+T1UwR3kjbGqJJUpZWTHlkFzrSDyu2KyVq5bj3K8b2OJ/TLcfEUSJjnqD
VX4gbyUtrt+oQNOIW6nbgQXrqaEIOxlUgyT1h1RpGS8GHDIIsfZetG6FkKlSifv3
3WDh14r91EIOmDrtV8kQqcfmrr0PcfK+FunGME7dglOI1GaWzFGDXsG8khRdxWxA
iuVypT+7kmTJj4ASK/CQbgdgsQ3W6Jat6Qw5H2MEY2w64Xp48zwOrrF7Y0HcDvVo
QJP2LlusH8LhPjW+j8qUsCKFHf0j4jY/U0eDnTkV3u0cm1I0krYwGu0RhcWq02aq
EoacaswjZ+ZLPmy7+qf4QotPCT/cIcz9uRyK1r+NR61LzXi5x4KpGW+28rimbmUb
e2ZpUhQOY1M9VwgK68v8ZECeOpS/Y/zEIhghhg7Qjz7rrD4gHymAhonfLhyRV/gv
CzO7gx+iPHa87C6SKNcZ4g1WBImEBE1yaVZcwzH6RKqAZyXPfpCl+ZurpbfavPVa
8gmUwR9ChqYq8Bh3q4XJPBl/n8bhjtwjsN9Fr3DfXxysIwslQHDFn27g7DvwCMGW
hyUFzkEGdHnayXDs7nyjVpnJ1QalTWF3HnIseTTTEWfns559BovOTTKg+5B1Uip+
wF9IGImPVv7d5jf0jAov+nfT0ty9jUu9RG8zc28GfIfbZLr7rD8qrO+RX8sXfAxu
Wsq0ctJXlCwTC4T8k44STjqh2ofkX4J1+YTWPULo7o5OyGwA9zZEYIacqK+tmdO/
SLS6cMBhClP1CxcuAXmOBoS4TWtraHFXpp8i5an2cTKd9/v2Bb9HXB6/7/ialuHS
mj0TZJsjG6x6uq8ijx7e7KDOjwAqJ8DdMmeVBTu8TGy4B2PAnDPL3hXW0sMT6uHE
KF00xVTNJnKfwZMDIPvqbVwd6MWgSOeKwx0DHlyDHkfLQfr7lfv8AERRXUqoUKDc
lV4/acIdSQUHSWcidWck6cMT0Ihotu9FtZiDHovHbWMiyMkfsrkUjd/zMTsKFnYv
jHZ+NXYDONPNEssHRUffQTTnCx6aU2MzGVt41CapHKrz/dMVudtiJdPIMXsgRPsD
npVc8CR/H6MiUlKWpCOHn7jKbrY4Cxn/IewLBQKBvc39aUdl77Wn72Ktfmx9zJl0
/x+Rqe5PcmvJwxSKpjnYY70RGs5eUdViqfmwMStqxdeZrxT68tisPH4OIgZxV9BB
ija9zmCZ47V47IvgFeJDWNPskDhHzMCWQ4BrV69ffUI9qCziKs9huQeHvQ/qgYPL
TPlQdL2UqpsNHEN5jpB6PlhFzjNVcOSVla5nNEFtLI/b8ontIcvqlNhcxxhSeAk0
7BsUk4ip10FlcU5pPiergybansvnqUDQsb2SKfnr6cL0nk3hQXbJKFJbW9m5jswE
1BE2f1ppzEoe8n9G0fQShkHYqE05QDT7jHaCXA5ptGU7BIvDzfX6x/5lmahe+Qbn
0lzIbNA5IENLXRiZXFD22n2UgZYNsZOZWGu86FcCPylaNCOZ08gwSWOqfytb5bxU
Cv9aveZN+WrSf25Ogsa1vGdH9q95Gsc7dwz1ZiT9HXuRJwrGtbwrrW+iznFG68Xv
zE+9Pks0zCDgZ8A+9nf6Nfy7cym6THUQe2Yh6iqcdF5CWC8mz5BczM5LeqiHSuSR
XBb/9/KZjPMHtlp7IKicsLd4lKmYUp5s62U4ze0kePkNAAK3v3VxnFZp7gAKYHDm
LTEDqp16JiwMkkywKYDomOQdRsQ5RFevhxK8Y+J3wgGp7gnAfxVEsGWU86cDu7y8
ptW38l4kmFzAAGaxfgUTbv4uqcBxtgAq06ontVjNI6F3LNj12f8FhE5cSlVTqlZX
jyVLh97Oz9fhNoRPOit1y4k7vGM9PDJjWPh1e+7dJyxvjJCtWOd6uJyBUV1M/R1V
OcHus4de5FlDU5U2bWP3tYL9Jyx507+OcgoLalUerm0Z1La60b9lDVQDrKaOX3fF
IkqWEqAKdg4eGWOzdok7dUUGNhXefuODiTJ7juLbPGplNvqjmciKu1bHFZYrgp2G
hmrbxtnX7AJc/M2l+bJC2HXoxOssZiWx2lxrNZSG0kPmvDg3O866isPfJAkHWYtW
84I2xWx6RIwjFS7sYkfT485rn/jBBhz6Fg1Xlfmo7CokHE4Q5ksXFTsNyHyeCp+9
GPHmH1TYUxEbvx5ewEuKPsoVzeWbqUS/xKPc1PYQ5jXPxkmVCMRVodEBb7ssxYAd
tNm3veC/5D2MUPVHB4yLafJ4WwMay+84tpHB+PVHvKV8iU/q91+6PKOW5uOdSLX9
v8P8cD5PjcfVi6lz0Ir2520ff5LGO+RjvAU3M5N8SuPZrwPT9pOg7022LEXkhVNU
PEy5qGGzDzCEp6+21mCqdNuXBdzghHsAWu0c/gLoCNgc7IA47xYTLwtR6/JynxQ+
+IKbqqbW1rHEhFGXOjJCFlSOnHDjQ0rhiuXbgYElR0H+fZrKRS2rOF/Ce/0DSwp/
za6E6iYq0qy/fXLj6U4sCJpBu8yNUkacjHERY6koiytfUXsk9s9Y/qLJV5Fl8T0A
+6c4d739wshw7j3wQCavBeg3umpLbHQtgXMP/31WXnV8F8kq+XWbEPS9RKCV9g1t
bk4Dwvswp/F+08yIQdfUfLjl052kRsMepfINKqoCBaRYXP92qYc8XkH3W5b8mX7k
LvBMt2Pc1HSiTzHHEG1xrSmdezdjCq2PkWNkXjEDubfY+Mec0hJTJMvXJRFhC5+g
kMkQ/Jmp5EYMBlWCw2Axpqmd2YPlYx6ROlJY4UelVMDvomewXOV/hJ5+5lJjdD1N
hy3439kfaIsm20aViN843xfwsrNyX8Op45zyc4KIaNepja+cDHMUu1xml9ZDJWH4
IgJLfszULqkBZrvxP2obI3/1TZkIcF2CBYawblXEJUoppWtKS4z2S6tsB0V88Ie2
oFKguEk3hrSwR/HadaFpb/HZ3cBgQDfQhIMDvTt6mQ3ZQUJiYwwRj7LIhFfR7/bz
3ybxQACT0RhS+SDTS4NVmjsa2CGszTI5OTkJhhpUsdOkzivjUjOm/+1/94OGAPao
Kss82LFkW6R8Hh7mBfXWDa2rL2alkGZRL81Ib88+UXT+IAthvTN02VCxhxahUY1u
wc9NuiQ/ZxFZAKvDELaFw4CRvOp4PR+biYwH7rnaWbxUtpaBURwfHEIAUffVT3QU
/LIsYxu04l2h8c0hQPg+ryficmS/lYv6qwDB6NFd6X5LIXkA7700NkS0/k5aS0ey
U2t3qEKT9RThhC0R3Dlpk5nRPRu3uqIWz0nUhLwrLDRtwnrC44Amy6XfdNdIqdQl
XKEYDUzZ8Z2PbeVuXbXz+rZiCAu3eNGGY/XDF+4MnL1Q4R0+X+pHI15SZjSXaZNu
lE0BX73prwFyAO4sh/lYDvrpomc6iR4c95g9UUsAuMu/Nq+0SI234/mqNBCfHEDP
oveXreRGkY410iSkG4Tkdd43ah/2G4p6PSOxRjGh8zZuVMrINu+pFW+SUgUkEcT2
OvSDEnBPkqBBUvVAxv1oldHwAQgXyxZOuqusGvj7hBR1FTYhpgaLQ3SOG4H1UTIo
Yd6Xgkn+Rx7ADYh9uiwhqULX0QutlybA03MAfnhf6CIY8wp+aRg0V7IojjjYcs7X
mrUp0CoM73Zuw2qRio5GoHSA7iAFfFdvnLcNr/pT7/M01/gGWAIQtMmYrDRdTUgF
u15XSQ0dj5VmwmTkKkxL5uMDWlU16MeuqAgjVEdHEBODgWDEjVWPD5CgniTFXfuK
kWBY7kLUHI4RaHo8I0piCWVwOjgYxcza/xyU2wxpH+Rj56yMI+tDYySu81jo0hJo
Zc2TYJlbp8cB0rsd9uT9ZcxQ6ESN4qWtzuYjfRbWqJC5hDFW0JfL6DhakcX/0Lw9
pLVel0H119clwfHKh7VXnLG7Q/gcgJ/xL+kG7RtPp3Jmp3EKjKfvQC+8+GNh2H0z
kMNQuVUKlGdamID29se97FgwJs2pEfPGYdhl/9KkAp32h+BG3m/u7vyq/agKE9zj
CpBnpFPsQ0iz8ep5R9PNA2H47H0UoiBS6ecrDa3cKw22hDEVtPyKTVBN4KqqmmgN
DoIoL8pOwjqJKqjNP2GHNOsQxyJAMkQHfXoCxuCaJ2x2+eAiiSnXSGvCU0/B2+ui
CuRFfyx+6+uDc/WxwPBbbhy90rRJeSrAPK505DegU8Cr7QHmsMeaMooF7SobD2Re
QBnfVQrjcDLin0j2F3Iep3wRg6A9N+zTikpdBIY0aTRmGd7ZeQA/YRlFlFJ8KH+A
T1JQMMGUtvc6Plb3RB0fq9aqf1tPpTE64cJveM82sVfURZsXCFQp6YD8O5vrHwHx
+R7KAn5KnnAZkzTEzTxHAf9CHs65hGX2EilVATGa1dVYQ23nrzomzM6WjkXGsskU
e25hYc83gptieRaV53HJKoXrpMhUF90heODvnfdCemKCveXCLpm8Bk2k3i5/KDow
Ul/TGO9psckKiBqvNBXsiRMMmfbhoDrbH3An5ZNFjRBMde3ODMAboIxWL9E1tm08
8/Rx4g4IXrOcOD925ng3+4dahkHO5S2NtBYFkdEUbxrHoXvIX+Crje41+jI7X2cD
VcSHGpUggAMrDXBWECpeJvMGFW4b69G4dNOqIjcKo4bEBHgxJwI7Ita80IRFU/bX
cNJhlLOH5aNFFALBI++H1/8/OglIC9+TiaEfvCJf7COcn/7C6NA1Tz5kqH1h4Dbn
Kf0rEkmohstaRKsRtiD6ZNkUAlF7WsMj53rlv9Evn3XPQRpFj8e7vPoJk+xBqaan
wq79cmPcjwUAl0roN/RpZtqYCUxqfYAZ0+v/dlHXHJYEBPylxkWMUlKGjsczKcN3
OkDFfO1vgEa/iZmKUbOtsmJgyZXptTLjHSvDQ1RZ3b+dyqvUoRx7+/J1i6XlnWfU
R1Bx0YD6s4XxKn5I950SiJxMzbaUh7it3+2wV3fI3WsmzcvYthQGjvuzcO/HTZAi
qHVDwkiDAjY5/FmnJVmgcQUIFjfBcy7bQa5ks6l0aJfgOmO0uEZ5/Q7eV7rxPBbF
fdBR+ygTP91JTlNyZPVs0UIcLb1R1JqwsUmosAnPa4++bHklulGgSZby3nWknJAH
UPyHf/p4FzjGvrVdCxkaM40QLzFOjmmhFNgnQjwFzpGXLSjmcl2k9+ZgGFb26mfT
5MRO7ALUSxNkNRucQ+UgOvtYU/TjQaQ7yCBy1wlsdtOyL6b9LwoE4SFJMcJzKkjy
ykYaF6p6OtfosiHBvy+ru6IVncuaQQjeDsEv6e9FR7yG432wvObHzrugwWOdCu7C
Nm8mqo9/NzY4UNK5iRBX+qK3cPuR1o44bJEtacRabBTPtpiiuoaBFo6MPJGsyKHK
m3xuG2Q54L+Z+fIuMCkP7L7+EsafdVJGRsl9bHm1oUCiaPA33fwLb0WKSyoGLX3p
Lq6+OYHj8wVPaTtoeVa5bwbO8ImNY2YFZdm4wfn0bBWkEdLcFP/3zKaGbmI74bQo
GWB18M2/4Z5/twejEuS9dt6cL7Gvh5abf6D7WfuV7OY5YlqQpbN27rrfoslF7YK7
ha/PAWdaP4+vFFU9pocTwQsH9BBhxIVpgYDSIaAC1T47Mq7pV9XRHxN8WEVdOolB
i2PKItOwswg0EyE6J8GzeJq/G0ms+s7OAAH1RKOtxw8quUvdqFy9i2SPCFk46lii
vHbtRtTiolSCvYDONFuiSe7tzjZxf1vz9wT9ZX0EdKzEDFffThajXfG8fX6zVrFY
wPBzr5IAc1+2eptJGhGt04QdRlEUf40jJi9mNCrwWGrRq+sIRvFi2BznsRkcUL9Y
3dE9sjxjJooXL/zkfm7wnrPx5g0sNf8uVNfus+S1k/e/AilT+LT03dMRhZ/DsOPE
Rj3rxKouOfGCGOLLAxiJvnKHx4oyMKodzqTj9OgV5gRBH1IEa0UXQpIrIlyaaQkJ
apK/l54rDrkAp0AjsMofVdgQYVjNwozatbrwsemgGzvJR29WFKYbSej44xXew+yZ
VNB1S8RO0/2JEBYP8mOyGUEce/icesFK4lZvpzn++fqdZoqHpwOtOPF6ytXc0EyL
klUoCOFwS7lP0VPZcxNCLdsYWxQsbVbdFgqjU+6e0kdHNynvDes8RkS9R8/TUX7n
5b5SnW9Ld9PUmcv6YUjTcvcoxXsavzKxvsuElCBG9CgAIjaNL2KF82f3chX5dLIS
JUvBCDIB6nJBc0J/J0Lwo/iKeweI7bPSBh/8QYyCTD9zD7DyGgjQyIHHbNQ9K1oi
BRCbtNpHjxdD/ssv4yKF4LxoztCkmJxxEHKe/VbRxqdUaxhs89iFwXxMej+I+bCV
KnbySPTJLPpQ6H5oJEdlmPGvADUBPIzGi8CIQSUD5s7erpMKsaaxAgE3YStiN+Iy
06Qhi+PNScwHC28uvurzrImploxW8ET2WkNVeBlKW2HxjPozadZshx9Rw0795PuL
v666oUo2Mm4fC2WlA5lc8bDpAKhzEkJDX3nct6lHW+rRlgeWWNDCBYliZ0eVnxi0
JUoALrgBmInOlpSFq+IcfidT3WSn6VVViSBkFCg4Auws5FLwFkxPlazDX5DfpX5m
7o/Cb6tfrrj+eAx/cLD+Ns2E8eWuLJAApeDxNI8IjEuvYB0cPnFdfZrXfNc7R4XK
TaJqSBl3rJXG0m96ZMcnUcHaW15Sibmq9nbweakcKnn30kd4omCbgCBYNV5nUpkp
+6sD6P1dyZMS4Rao0SpvTE2zeajiB/j6KN1jOtwjDRMtIIlOzoTh6QfS0Zwlxn8t
MaCsFMkWj88VXNderMXrJkOvOMlGbf9OZuqLelrTTGFjU2wjFWbuDFuTADf6AtPC
Lf/S5FvRFvz9kJwmFlBOJY1QLio5zqK7tmS83fb18aZY627O5zdP9RSPfMp1snK9
xPaTB5/Pdogw3OWfDrj3ZY9PBc+QPMcc1BnW+LvDuP8uLP0csQlzMiecv2yEq+M7
lUrBVO3iGytXTV6z+FaIco1og63LWDvt9l96n6XJdJaLQvnpuu0S6v9jvUuc23NI
Kxxp0kmCe33T31raX5Fq7EiiZIatye8INIy4Ey9Y/67n89ZgQplCx875iJQM5xPm
+yJOFo4Fm0paJoszdAsBUcHvpPy5u+E9wIVnkiUikemcR7Ag0dTO5xgqZWCycGpz
UraSH6i9sRSoVHYY04E3Y83fmlZMPO8N5y0wm1IDru6GsKV3s4wt1atWNGNBSzQY
TY9mEbBNgJjQ6bBb8Atipl1GKhzXvduvud+5Eiv/deMMMTn4tgBjBLwENJiiAnbu
YGTKYcb1UaF5r0fsAOnTnqAbGDPl/How8XLgwOKbJyx6bePUd2jjGmBcaTVNPak9
aYIyGFxwBJD3zK5Sum50Usy/SwX3TOXadWNl6Jyiuxo6fNCYJlvtUeRWiFrsGZtw
YfBsRMtHQeNLoUOl5Lou02E8Bakec4JmxEj2PqyyLwL3UiqT7IwCY2htFoz94gyD
TPLXKq7FCNp0CWRlwydWsyMI+UZqQ5JRbqnJMuZh6YGcn4KPrVS8GjOUZctkLNyV
UuFGIuxlM4ihkTpaHQ/45uT5SEM38Kr+b+294PGJoJAfDL0FF1Eq+hc8nwlkcaT1
GgvU6KViDjrr2da0ePO4FT3Ib7gxzuoV0e9tnxwr2cJqPsOjw8PMYPmnUUkQ5BvZ
TAMSN4l/rNWArcwZlhmz+IUEr8CbkYX6tBFWYGATHMZ+1mCmkxwFECCZ5ret7Ar1
jlP0rt0UAQ/lWBmJDfOhX80IA9Ib4/hKVK8TXE0weCrZYRI19rS4Zm5qQlH2US7x
0jMGJOZ+IGrhQGoY8EcLvhjkajHaQZUjRvSeBR+mW9SFjq+NCsiiRAF0CerdvlPW
sMPo85vJeLmt9I19sWJKO8W38I988oZ26o/iyuJ7TMwiNSA5slEpkr9M9EtVLyBb
OBfzpPlH6Kc3Yzujz339OtTnchVHSJPqWadgL3eASJ+YD+pnZEjqKHntnUwP0KvE
XJmyOAmWoVZe/2v2Vz9VukHqHx1+V5OtamMT1bS0gonVsySauRzZOIJuCnCGOaCv
AMH+gQpCDwjkk63+uhn1AB82L26MaHAm3IJ4Cp9v1qVWqoqoVmyPsOUI5V3vDRwu
3QOGi7b00eypNulvkCCEVJG3CKD142lh3paTzY+XqrV4YFwB5+mKVUghtSqnkL7p
nTPXjJAlSmWm1Iy4PgYvzmUkt968JCF1SxKiXTAnmThbaaadpPjfL4SrXXlCOIyz
SGZBIHqASnaQFITtnribQFF65bSLDZfwBWNOZepKBUATPb0sWrgQPUl6UsRosw9A
k7yiQ1TbO9AJ5L2JBDbO3AbQkQ2UsRmC7g0DkAaRLRr/xOst1REu0XYvXb1HFjgW
/NjfTVLRudkYQWY2YwKmmYBTtwSPZxDSCDUu3A69OgmlGpZK4+/FDXdB4RMuUOdI
i0ZMlHWqNw+JZQdF8JxB9MS/ggRdBcrXncOu6j0leFtLNhGlnbUbtHDsHLA6R1re
wwqGU++qXIKR5bI6mut4DFw8QtloRqPwh2lgdQskgvjqkCf4jzUgoxpFyLJ1Lzo3
KZAWTK6PTCZL9ejIVVba7x9Vl7vzy3u1iADXjhOhbN4/2VWkvgRGTUn/Muyi6bF5
8sCDRAYa6bZmrJ1m6AiWTplXuNxx8vARsDGj7Zt/pjKGBAAf1WZHISdBVSAwbmGw
StFYCTDHIuoDOjk7l5kHcLZZfedQBPb81Ntld0t08mg1ly86YFISQ7QG9xTdFvz4
XtvdO0W675e0ZFLbFUMeVp/fUNLBWxBYfNTW4A02LcgDWCvi0SaQziJw0U/DI02G
XRrsI/FB9TIvBkeBC2Z1Kd6w20wJX4FdA6TT4/lYCVdk5SYfoiyQZH/Rzwv/lQNj
oJ4wOsH8hy2ExrK1Nn7vfw5ZzCh++wrF+pB+cX0jSn45aKE8CZuK+pGPhnKD9Btw
EuG51L1SxU1KUfLJplqrcbeOI41gIHr1OLuktq6sswTlN6nM4lujPTYg0b9fJtyt
RR5mxz9SfBcJ7/oGaI0q0CB9cjaru04JjrutGi/79egCjDifbGdGbftttH+quVOQ
Zr+jUrDWZdyx1WKBTsat9m73pvow+Ipw3DnXZHOpfFkJfWXbQ+3f+ULC8YvTCDg8
QcVGqRp3KGVnP5ydHqKBd/jLYjonRJDAgjByKUqVbi7Mr/UCg47XLdKRcNIHMvCo
`pragma protect end_protected
