// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h4qsCpErvLYYNKyDKjoYNXGr6bYWmDAptrg/Jex1zqNXx5A1Mm14qg7cc2a4zGU7
BIajpdt5vv1Fm0MZR0T4N5QlEYCAnIcCb4kML5ljZUGjLsOWE/8A71wvFwOJrNSb
x0hKlM+wFTPQSQFMQPP1q6McsWj2Iqfz3W2ZVofMd4M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7488)
GQ8E81IdlMTsrFNV8b8Ycnu4SsWQwSx9wwV6pwQUU1F0myo/e7x8NJueTU9kYr0a
TK5rZZXWjSjRmt/qK3zp8pI0QaPKwHKY6hHXvI/7rpQZeQ0sCKZzYNdgM6/dffbU
FiuuBCJwGOfyP1mvv2QSeBf2tfL1xnem80tUhcIkySBttE/Tw1tslFS2qZ4FKioq
HmV0zxc1RRhFFoXFpfVaX335iXFfLxIKrFF+gTFs6bUJjUvV2+VbefWD9DR3/nRl
hQKXPesa2xCMAJ2GVmYMqfXDHwZeSAHB8oA7T/IuJVQc5HIJWomDkFI7vtUY0Ncf
cw16+7lBgQPJtdM5Dl3j+WXNWOz5doobHRaKccdxvJOOZZEtKs4h4v1Cq5BqTcce
Ux8tmx1itsqJy+xUlXQg9/RN8QJ8uHEUSh1qL0oVTynMMWCLRsiualwlB9k1w/cF
NVl157OzqO0TSXNQ7wHWJ3/KZpacTwVIcfb8UfB1OJSB+BWHJ6TtcQ9rzJoucLl7
XD1QnxaisOPrwM2/3acEEQ8kTiXins9rLgoxSacoV1d5vdOOr9laGGI8YMI1pu73
l11fwTUGEf/Tkim9Wk8mlNHkJ9SpUmLOOHA/bnPy87EBcEfXJCpTWHTxcLOJsdsD
OMXjCxSnPO4/nJJ2o9W+qUF0ZkRe9cLgB0rsMPDwj3EJ2g0fL3yTGZJaBJTVQIe2
+heZTcNUD2n3RThRtYqcTk0fFF75MNooUXCgw0nYtCGskLOtE5iGFmYC9d7msbzn
D3b1kvIL0wWEh/n0grC+o9Q5EhAvr0hH6+D/QGicLoY5z5sShdxh/B78UlA47hbh
bShcCT6U/uPRHy2wX9Ei02zZTbdwgGlfUTugMUJQeHX375TA7zTNlLxpZOW9JvBi
0+YyAn+FEaQH3BPrv7wd25Vo+gOZGYUfTNlIr7IyoGKgcrB99cfdsV93Z35szU/v
4JqTqFD3+YyC4ME/gOeU+W7wq4vyz8b5sez7/fx+6r6+/G55Jn5zXLkJDGCiHDEU
1UTJhOKghMSo+kMVH7rKJVFIChl9NaZdUcFZrGeS1qGw3lGJkizJ9PqePFfimINs
g3fxIeYAJM6uZVuq9RoDNAovRS7c8T6uVXsQSL3MYEm4WeBu1Jkq8DIndfCPkXZz
MeufCbLFgwdp/x+QmWFK9RbjRrwdc6Qp/xFm26P7DiTKiOOWCVKtG6vkQLqKN3HE
dLC8J9QvJBXtbu7vERitkSSZtnLDG/SJZsvCn4X5VnmTsu4Hii49N5yOktyAaui7
zWrxothXD6c5TGjDnlYya3Flt4JC2xQkt/ltjbZt/tnM61nPSP8JG0On/o4768tp
Ne2SNJiihWFH52Qh0fOyh1r7++wvFK0siFSL32syXv4k4Y9g36IMUMxnq7kYZ7Il
TiGho/q3LI4iRL60nCkM23DXGy0ESFlgsVGB5yi4Z/R8ZXVnGO/EAyxvbPCke/Yx
fRZmun1yBBsY4xBb32dxguwagxBJOEywQ3pxDRtO8pu/YOdiwPnBUIGxn21E/buF
DsdDXcvL6ERpr4EdllPH+JARSB9rcJlcGqV+lhYoweeQVu1puP9cyXM069PglrEE
laivYX3PT4KDYlARNiU7uk+XfKF/Tv+42mv3dwIofHsxgUWWVG66zuL0PPmJUTEb
TahR9Q4qReR6YQ4UKBo0ZE8Z/0COZDuUnll0osy2W9SL5Fp97gJ2Ke2Llt4Ju8qL
PMKzhG3Bvhmk0+pdllZz1Wv/EC641n/dMe7BMoj6sBqw4Jgn2vrEW33FqYF6Hf1z
ijLoqaae9LMMZSrwMvzkn6CaNPmj8DRPoqNhrRlTJiU6JxWoR9EsKwl6aVO8TEqn
mm5HNJf1u8o4mS3RgVXIpm2KSOJgBecHdfpj8t59n23pJuvwCiiscxGg5fMz8AWS
taUaQ67oegQPh2D46IOiH7vOnaHl9mffRiI3n7aiLv34Q5TQODl6Q3EFurznE01y
nh8aX6EQyqeKjcRP+ucKj3tfU7LNwHB9Bv7Rc7OyVWJ13ATb+k3VdBtuP7ak52wM
MvGPvMH0gOF8QDSNPcQ0axC/r6DQUyqV9nLZZQ+3Q4c2qhZVmyFac/ZOc9Kwm1/4
gU66SXmgS3otc6I+AyQ+e+DkTq/NfDUF8P90fmP15caWtkIe1sLNF71o4EAbb0mW
TBxraCaZMOFU/UazscsAafR2XzXyKBtaNsevUVMRxpJEH0i+lWJQoNFI8HHsw/rK
ytwwK3DohOULokmS0PjeyG4V2mKJL/T51+G6WbcjScY0GoPNR1B2HN1sIVMbiC2h
lNt+HrVctUJCJqEUc5mqUjnbnMAOVjmVsVtmB4uGB6K693IEhKczxxnEJ7o2uGGW
gO+T10eR06PsElcgmv7kwNDQcZ7ZvZ+0FuQmYXFCa6grnuUle/nLVp1sLvMBni6j
jANXCb1iwsRG2b1qCNL4k5q2LglYdFE9nNfPYslDonO/GDAIwJMS7pcU88zoax78
R3FCUZK4qjukvadlVd98tEf3pTdLn/9ydqudxz3RNeHHw/Ev5Yr/VvjNoivAw9nI
rAwUjIsL9/Obpb8quEMv3dKS2U5VRV1dmNz47XMTEz8a/1pU+xC6r/9+ZVn98Qwl
SWu6gzgL6s8MuySlhu7iVLOFVAfpkg9zDYSwgs1/+1Fop7clJYiojNCHFC1BO3zj
KfB55ebA/2kVY6pJhTOXN/DapAApkZ15SrkIbFx53T1/nPmZwIO8QPqrpsZJBrMV
OH6C/EV7CJeX9qJloA5Ur37KWE2rscBkwRjQzbiFSlRy8xQ6SdQf7YL1FTP4J7zM
n1sVZ7zesjMF62YstVT/v5Q6dg8hCl/35ToU959EiDaViUb5+7qrH3pXHGehsSIB
r0KlglaZQWjLYYjQBYFGBtJ+VJN5zklhoP9XNCN7IDAF7lRLu1RgvvEDRx1V/Fii
5yxVEIZhPf9I4wz5DJSsQ+p4x3lW5OF4/+cFw4lItbI53nhNmPaZ+JCok3CEjneV
p0HN/4GrvEOQ5y5k1fyuZQfllec6bPKU3GQ3pgwsfPN2fqfi/ezzJ2rIse9clnF5
9uOlsKw6J5192PUNMevt0Xg8B7JaQNkfFia63GEo41KJiNHgyn/3WE1yAc866/Y8
Ph5O3FTzOuTZhuY+JvjUND5CptOM0wLIJLm4pwvNWR43VSbiDdG5Tu3YJC38AfyN
y1O5HKbVR2xEJHEuFkR5CCcBlumnGmzw9Rc+xKfw1ChhlGJYPf4noBlEa//V3hKv
FXixUXUKbckgJJ3FTtM1REb2B4IVX9YOqFCIOWCsJECYNdGpYTaJ+c6VjFBL2n7C
G24vhmEOm0fmYZxs8nu0RrYlxfkWsfOTs5k5Um72C4DUcFHu/nA+4Z1zKMczRzCQ
DJqP69C86DDNbR/SZDuUtTsZd4R3N6p5Qva6/JYAmz4FKqr9Rhvz7z+zBM4alOzb
egcMlP5abe4vGvugTKyva4eScq85pyzD6Os0zO4X/lYYh84z97Y4CDrzzCXrabu+
mg2rhMkf8ZmYucc94PGSYpbIOy5MRI30dTg/MsZ+GF4X3/vaeuF2P0ylTV9WndMO
D3RVo9CC+Ut00uruOeHmg52Yu6sKgea1RCZxWXva5yGTeSjh2USxOlYN+txAFMDn
gjZBD+vhRujC5gCwbQj3PceFZmV1oSW53gCN7XMB8BipwaNIuVV0kon5qb8qqt2u
KUwo2ZVuSHBhTOWtnOYjRV+7J78gA1ZwuUCDlj9iEyKMCvFQHEGT3Igqm647tb68
NoSZwHzksza1TPsmvCOiT9KmLl/Y2vf2/CxqAVmCI2FVyi4Bjk7hXVSLFnLUpe6H
9l856IBvpTVe9MRSkce9Q/vn07Yyz32Wp6KS94EIA51jxxMrbKK2+mSZ1N++Ps9K
SL1FXMCEfsWOfGSPVwEWS24toZhJFGypH2aFWBdk6mVaVCBjPUPcdG5cFQyGz3YO
VEq9yYNoO0WMVHQp5Lnw+xE4Ys/hNQiCGpszA6HzacPvYKKSYhxbolCmfFP4kFV3
H2O0uREZOKoKXUz8Be79NyhVXlSxfrJg2AdQ1tMfNQAmj3jX6y42OSi8gBfRIs1M
HqB0idcm7S7q20QVXWgZLmQ6oo5760v3Adj2K76+eeo12C+YjZ+7fku3MeP8P5ec
IdUktf0en6A9phopczv5S0I1Mj8lqv5WF/GUhjNlI6BiYpFRgxJo6A5sKWjShOje
nc5alxeY2glb86qqJ5NNSiTvfgCRT/iabZm5XELMMPwKDPpSw0QZfSomXKy1KHft
9MfkMJYfz1GtvEJc4n5Erjekaq9djTY9Nt7JPyl2kNDl+4X0TqVOLXEw6/cRpc+d
Q5mnITNgxVBjJSaRKRZbVf6V4HqMnpcOZB2vEVzCzYUHD1QQPtI+R++b6CxMEpf0
ac7xybxELEIT2A7FVpgzzLgZOrAtArbSIbanIonQpTS1H5Kg4nX8qDGT3H22aHv0
bxGBmlMzvBIUY+45JvLGer7T6mFdIVHW14VC0t8tENaM3JJrSAQFSUNwMPKzMqRT
XNS+/VKm3pQ50vz+VcXlF7VsmvMNPwiYmIOEpGlU8xOTzNrYJ28PhL40xjhyx1QA
Svwx5IGupofg+2umkY0WqgmKbjmlo+6X7267DZE3WkCbZLH/4NYUa0kjmvjiGzED
l890M3/k1I9OVmOYszS1S1JU/VvCDj9yquHpekt66phQc78FjRzxHGwflZoh6/rT
e85YiOw2dCdOjEZ3UXwc1cSoXOvrX6A5EZKYgwkViMdVQDK6QH6A0B+wmKcw5qoC
POPRp+YFdB1IQk6LAOEDkLMvhrYzD2vD+4elCxiY7ZAhY6vNFm4h1RTpxVAuXpTb
cS/qezJHoRxAUOmJTRyMA0Zz0ekmywS8MIgkcOd31jMcbPFuuPUElNhhS69oRQ/Y
fSotVeSp3ZgOTj1I94HcYlRag96ilX84TLvkxuutjQzt3kihnKMx7EWdlzz03vHn
zxB3rR2eOUxF1rygQHf+YyddhMRx6bJBo85T5DMe6C97p5KRm55Gtuhc+A4mxG8B
FgjQqRvKTO+3AjEfxlxy82T1VQJdJvKVvgeAIWBRYG+1Y9c9NSwBsUt/WQkPl8Pj
B/gl9kBzHEgTLPWiPzALK5uuI7FxlXEv3+8EYPFu6Cm6mOMbW13UiMBuP7+JRfqM
qKavmH0Ld3QTtXT/BIiMLbme4jgo4j3zlZ823RYbaXXyecMwMtUsONmmJe1UfoQ8
8bYqEpzCIkVxgqG28m38TozsXfUJ+raqMcFMrnOsCRpG84izZVmOWai6D/kRPsmX
VwUE+fiE8p+FVX/xg3+WbRKlmFNWwtbnU93z70qHoyJQZ1DxbRB7bbOQK/dAd+Os
uLKMuSyoQ7bN4p1T8ZFoh0s3rRETpLjiYQyaB5RkHK++CqoCKybwMwiFABwZbksL
iDqmFim2RAx+rBqKG5HbOxPDEIi3ZFt3aMsiWrW4JiWlDLeloqE4OlQDru7pAdKw
O15XsGl7i+y0EfSTcNg9Z94kxdcgY3jMBuPBhI3o4ZCb/NwDLAHLaNgjQzfZfjw4
GCzccM0hFGETaO3Y+VoH+FGtqmxk/Hn5WKeWfhBAEmMDWwLt5ZVq+45gUps/Yik0
dswamSoTawDFJWiFBmDeVE8wxKPLf/6KRVmY+yCDFFLS6AuOOQ3k7z1HckVf0m6/
DZAHxyw23KucHDFM+2dvRtUpGhOkB/9nRRa6nJ0OyiEjIzgbqs2F/4vP4/WbrFwa
cFBL284LOlqMoY2aC14IFjD0dA6i0/ApfTGfrmh7NsjxVmbQJNmNXfaX3KTUWF8Z
E/IWj3B0nfWhafISuq17FPFrxb7/mAl9jsV7gwXdcpzIaClbIEKkC0VedNVOUU6N
bAE1hPWfmg7DmBpEvvW1OvTdasJWJ8qTsER1Fsmk8z/ijVV9PKbb1qckMAVmSUZj
BGMaXgzNrIGqUBB+h+29e/r8X9EBYRoKzU7TI4cOPMrfhdamJ47HAR7CMhQaLy2W
NztUQ6uTMflw9cKvNqllWTGyDO1L2Hdn+DUeIu95W0j7/GJsHaAYDHWeynjDnbmR
+BE7KW5x31JMuPEaUpgr5Ip/xZYxxKMaUUlV2Qg3pjsvFwQngPjqC81KUW4xNtDd
H/h5+kKSL6Vtc1ZRMwBJ6l92pEHdDJtmJa0CQPZoTZ/kW8T11xRwMsEmbI3/qmTg
xZESpwSOxwA2BjYfwccTvwWBHA3NXja/nX76NiMv2GRrxoGoxdNYQIuMVptqMG1J
ZhXRRr/hA3GM5tw7uZLI1wNqoY+OBqhTSq0bTjy5m5XGLG9kGOcs0Jc3cPIWEQks
L9tdGPPFRmea3TyvZM+/TkoeLBR97v6Md4sAEmhQKQJb3euqcoXNRvxOxTUIm4Mk
2URaytkZbGdcegJBpZkyUmcrkyjYBWnB61ls7M8s4+zorR9PeWXN1reHrjIFtY8L
SCWCgdJ7MB2sT2Vp4Hgz8+EEuux04sbN5Qb9OfhHD9JVONv46VymGtWOZEtuJyVi
VaDjhpW3QWZNv7WVu4WVDrydjlWSIBw6p1S26lXK8bLadNSr5rUJxt5vmBsUOw83
aivYqWjSa9KIAT6FSUW7OhXgAPPb0/zIdgocIwwFIqa2cVCKUuw1eVxN1+WUY7VS
GStf0iaGcPYnuYrQzodwBU/whVBeqC5wAKxgj3cd3PU5+edgQGrMvqgvD6px4FWI
1dnNWmmXJk5dN/+fRFGXk0Eqp929LfT/LvsPVIaHtQxovMgFQNwSlrYZgp1x/2eD
6WySjKhLNfmN/6MGWhWzbHs/zzYfgUhy81gdSKFC0PGJAGZYjLF5C7sKz8io6BaH
zktsxds3e83CrT2gQborVf8B2SR+zGIpgNW4/pxpKC4FmwWRPCkFVwUYJc9ZFc4h
gSUYcXAalOIXYBZOhfCoDd0z2Q++r3sHf1dhKE3lck+zoREUcGeW5YZ9nhS/U2vW
OyY/4axPfYLrU3rpqLpp0MeGIemdeHjbIpcBG7PUYWUbhU1QzM8JLOfaACcsnDJ3
R5L0dYzXIr31g4ZH3luYdTtGN4ZM8C2DJocY6AZjV4/rgDTWPi7A9H6r79irqHJh
d+F3l0ywNDEehW0YBLUVMCXLCGTROB89jcngVx2WIYlSOiuu4iFruoXDi+9lQI2a
VJpj6lXTp6dfzQDWhE5CvSGhMfJQh3p4M+vmSjF2h0DJdS0QW9Plfzd6fjxdDknv
oyelY07c7afyTp9l7BM2+ucliBIC2WYt9EiEG9nmAs6vpJ7m0MwjmcP45+SRg/cr
cEqgCfUQSzytHKnmj6P7+q0V89nyo9ilcN/F5PBk+eoFYDlY6X/qXsTNDtDJrsXs
UV/vm6756/zcGICxOOujASI2rDTV+oYniUxqghfNCcu8+nJbVBIH49Vkg7MbJncg
0rmCpZooyLJcphUTcccCQTj7usV5/vCVCw/wFq98hh/ZLmkQxzQh5KibZWr86GrL
2C8YAa3PJ/SC9vFU+F+8gdAJSeLcN26RRzx6bDc9A8HrsooFnjllSj8DuV6QXnJ5
zfp8JQNIQCNpNi6LzWH/EjLMfM87JjST1ICZASwWY8G9bz9pIZYFIgJkMJLrovKZ
Cf7acrBtW+MscxdxT1kVNhEA/dVDCsT2FLrSRkiAuf7uepsR5ZMHaisfvJTw4SEy
dL2p5SD+irrRkLwZAPRbfhqCCpbxVK0o/6XBdGJ2ZaFU2ptaURvqbwAWsRqqY8P6
E93qp7+R4uF1Eu3DAnz9A2oHKPpR+P9enoi8gAjIEoJE/Rjaz/xTYxH+KumqfMR5
ADeBCm3KGmHwjaHuSKw37fdv08OJEl3ajpSNmoU66JPM1jG+9qQVmZUcWc/Mx5+R
OlyeCicWLb6ZMVe8EEv2sI5J7P36hXknQHQCch6pW/trQOISrRPUn9wc7Tp+1njk
mCtr7z9+8dFtz46cbR45wwOIA5F7QehM5PcJff3+NMeeK4NFJIYLKSeTyOaaZ8+D
Lo5L6IBFrAKI6rDSv/Kk33cK9YHgQNmEaWu9WuwHI3aw7bL/CZfFm83zUFiVj20k
2FtX0bUsH5Ca6OgYZjm/MmLRCJxrDGvojojsiLjtMpHDyBqGlHm+5v56X43n2JP5
FRTFdugfuDfOwEefBDRWfcWhw5KkyrxasH3+tCik4Ty3DPWSiI2+xl4+pJEULmd7
bqkrmmAGeCNS9KsotFk24Cajri6CBvZjVnid20tf78fH4CcqqkQSM7ldmgOhrKyb
+nH6Nnf7xm7vR+766rmQ7cOL8IYqh0F/n46fxU4Yt2i0S1n+fFIXd1tDdX0pu+05
eLCp2MAIHth1jKQsXIs9XQHUSAricTWcdGPohuSoxqetNbgo5RpsJry1h14NYg9s
IKyToTFfY6fJuuRTjGPU8kU+XvthlYqkUb3nQBkp9WucisRix4G5+ry7QKzHObsQ
xqjBGa6pFISqVyApuN7JdGIkZJFwB9abU6zs9e9OYbL2j+tObX4wtps12SngThRt
9CmdvfQ8qYrjmxI71TELnBb43l3jQ08XrKi+Of13mbOF/fcacj2tmsIdWrJSt99i
kXVrz1gQ8r1CVPHQaEjDiOam4bZHYOj+eOUowY0sZ7VbESfZeSD6i1vggLv9HF+3
guPXNV+xhG/UbqXl5kkOggSLFoCudGfbR4Jzcg5QZusq6aXlM3b/TVhQhbratz+D
PwbRcHOz7H7WBSNsgFLqH7FTR36uWIcXV119GGTIT/Ml6mCXM2/g/CXAdKbXQjNU
52KTWkwJ+giACdmrKmHhgLUDj/AzkX6RcwFo6CYhdjDeKCWIjHELAwliU553zGCW
FZzO64tZIVlPql3xXwoCGXtgHmSWfpBMLwBdltEFoS5gsLWV87VHj0rfhvduoz8U
qgGOLlAzvzM+3rxvgNk70lDwrNfsumcVlOVd/Z37WFTCzO2ref5aJ4KmkDZVUjXs
OhiDrhwhnlfL1UdfeYlpTCjRUZ/dWlv0q1rjwNzvSzmGzIzGSweXDJgZhwRG5t+r
eZ9grn8H0TDz/TRY8V7uvdTucDSDPnJtxGIAfhzsNdDMKURdlZdmgpgWj4GMm/xI
SuvRU+TBZpZFB6Rv0SqtMaphda7iWRXGMY0s428UPFjSbSavpp9DIDxbhfy78dfh
odOIEJzJbf2t+dH451pfZ5AgZDT9SriAXATMuAb0pOBtfRaj/XhVdmPQjb0MJpl+
TmJ0A+qDKHRPhKbHcfchXF2HhYY9Hd/1eQ0LCyx4RkWa3wpc4RXnpWfSFZsCKgQn
z59Pbkhdw3P+0i4LJxJQrJB5KQMASJf0QR8dWRb4dLRazH6AIq8VJH8Q7ESQ3oDE
sLaEH7WryZoLQiVTMpoCgM53w7PPyziozZeOPXaIIVFY9hP/aaKNgO7W7AxAHn9i
fChonEkVUXhL/udYAzSzpOGQMv/qJO6q9psLqT59V0Jw/d9zNXTyloFyLCg4Gjmd
PblHkmtDE2Dsji7Slkkqy63VDJmWiOjzdStUy13C+A8bKYJa3RLpYcnV2VYM4ipn
irhB85N5OPZVUOPUGJJfDVN5vvjE/aOaZZte9Re2cYCgPvB1gt/jKtksu0WRRyQb
XSD4S6pebd7Tdmi89uK5144E6PgmqRUIeSmk2tBbYappdPQHXu9+dIm0oLXFd7MD
BKMYn50YW9HqdBeFySvhrRP0+HLqf8Q/ThMIQ6b0pBfnFEq98fwOfXf/OG5yAueN
agcrIi2nwK+QAtS5MW67iB7TNoYs77/yf9uAV1Qf/xX/RRwXZbX4hxNMVyuM5uUG
EkYiUgNVJTeUpF/AUQtB4tSVJEYkVVfVDPtMr8s8F/kq1g/AiTMtfvwcSy1t14Uk
ukQJZooX+gp/AR3HAjAru8ewncvy+VLInJbtka5L8hxQWZ88EfwqiF3xZxD+L9JG
xWWyVtG4iyMEWRv1eMuvTIZJj+XLtoi3gQGW54/J/7FbrBF+qK+eWV8lRbbkUmyT
`pragma protect end_protected
