��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""���᤬����[���%r��E��Ka�eB&n%�������M[��.�%��T[�#�Y�g%Vh@�;�x9��3,)���yi�M�+�;�̾$a{�Mg�"㈥Z����_S!X�ú�N#��´�1�yX
EnO6�Hb�-�0��簐u����$�S�~��� �:R>4pY����W)_۸�KSQ��R�ƶ�}g>*w�r��e�ؙ3m�ؿ�%��}2��'T0����}=4cֻ�hb��l ���i�x�M�k�A���wɺ��79
� �˻|`��b�`0��%˸�:��.��#�L\
��so#rz�_�ձ_��H�ˎk6�� 	��p�E[�
��(*�9@7�nF�����)����-�����j��T��E<���Қ'��X(�ac��g��߫5NS������gɄ��nW]��A�.~�!�r�%#2k����3�����6��nT�kr��E3�l����(�,*�+!j��wx�F��-�I�3�����0B�l١I5w���gl�u)�"��bc�7���g�4���*c	,ԮV&�]���6�X�}��)[��	�&���`��q�8�ck�ϫ?U:�e��v�p;[8�|���<~ۆ���$ECE߹��C�坾@�&UrRh�Gi�����bQ��S���:�S@�p\�.xd��w�)� ��;��b�[�"�%�>���!�0�D��_(;Uq3J����9��nT��O�Ye�%�7L�b�,�?gl"��9M»��-�uME�m��R�B�6���|H���ztb:��|^S��=7 1�c�ĳ$�F>~�1��FI�V��􇣲ޢ/qp���c�A�4���λpE��^ڐ�k��~����ֲ�FA�3��iH��-e����s}�T�<c�ռV'1oo�)���E���ӪX�4�˂���a|$հE(\��k���u�a��l��Em$ �����:F�����ä���F�D�/��s�����Z�j�����Z�u%F�j)o�u�=u͎\埍QA����Z?�}���yqּ.�T�y�����J�x*�~�#P�V�Uy"_�\ѬW^G��_'���Q>�nh���|bg1�5�Eg��ۅx��cvuͤƞ��V���X��ˉ)h(���&�q���R��3��a��w�Ь�;%\#/�M-L}���U�Idl?��<jlgkkA�W��D�yмΘ�c�E�����(?�ң�;��ݧ>�-:\{�At��h�#�hhA�J�Vї�)8�qV/߃=�+AׅB�˥���l�7���*/s��M��jd�V�|�<q��|������_$�c�- �J�`��ƾ���h�
`W������&�GJӬaUG+V1�,=�ɞI�j {>��M��BL+.�W�s皳���O���KS!EY�ש����W�D��T��4o��4����Q�9��xj��w"k_ 5e݆��,.�[>�v�?o��aǃ�'-bπ������GQ�r�%0K��Q��6��^��w��|�s���Wi�%�U�{ҥ�ʓ��J�d���BCFRV�]6��b�Y�<���+��?l����f~q�'��k�h�7Yr�h�M��(T��~+z�+�`Xs|�	&�ŭ��75���=PQ�aaLޘ�'3�H�5L_
{����̇��-�P���aľۙ�9ȗ���
�t��`}z(���;k�tp��[VM�3���{�U����M����;,�.A��<|YoF�<��o���n0d7�lW��b���5٦��3А-��C��'��#�YF��w�n���`��Dc������YE}�`���L�O(n��C���PR��%�8�j�6�� ���C*�7����JB�K������,-���n�c>LY֔�9O`�;55 9Ws����G���G�J^[��+G�IO��� >���ev�H�1@���zhY�DX+�rJ���193[�a�X����UF[Ƭ�A2���"X�bG=�u�Y�-nȖ��li��k�E���0�<_Ka�s��J7��|h"n��6�#P�ܭQ0��<F4~R۠��"�2��XCC� @­�9j��GG�"C��:��~�D�W���3�| z��ix��6��\J�������:�,:��CÜ-�W�#s8ޠK�&'�6Y��L�0f��CG��K/���ܘ��e��ɩS����R��u�c��{p���Hu�Z��}�u�v����F �Oh�a�K2�"wrˈ�j��@�Mң�P��)&t7�Zc�h��LB/&��w؂���稊L���g�_�X�2��ޞ�mT�����6�7��=.S���\}����q��v�:`v�}��~��2r�|.:��ϕ�n��gW�߇��<Z�}obq���B�pu%i	�)\a"r>����8�������~�������;�E	x�P�ȧ��e -�}F]��c� V�4&�W��;����yOQu>^$ˌZ�S�&=Le^�����Ũvk\���^^N��>��;ŗ��Wq���e��6����_�,Y�D�N�rM�>k�t�*�qaT���]��P馣��ۥ�yË�3���zc9�(��D\ZQ�s!u�FM��q3��PO(| �2_F-��{$�Q~������^l�s0��.[6!��ʀ؅r�P�e�����2�٘��c0��a��j��YΩ�|�[�↾M�p��$yq��L��n�	t����Ne�=<-�	>#duu�7=$4����dx#w��U���V4������94�<C��K�޼_HUR�=�-���.�V�z��/�/�N�rx�F�Ul��/�ُ%���'/GJ�{�� u��%��f}�s��o΍�f�;[�N(����.{��Z��38���W#���(*,e��/� F]�P��4����Ǔq�2�l1TzyJ�|lݟ��%�A:SO����G#�*v$Gw
����h�,�rk�lw�b)F.��dyiYx�?�2��(����Ͽ2x�l�$)�o�xh���(�"�:>���]��qD��?����h�mw����'BO�݆���S���VV�ucs�ΆVvy��g��k-���K:|��e���������)���*O�A��1Q�����9��i0�K;�^���b���uXT_��2@�&�
��S�.�#�'���v��+�v�"in8tPt���ڱ�� L[�*`x�7����<|� � �x�k���Lhn�y)���ٞ�rH̲��@�3S���?]5�rbO�GTGջM+'��'�ƻ�R�\Y����ql����%#�-��������ԁ�R��?���NJ:�N�8���2���^���1�W��v�\�Z�צjT̩w��zsTʱ>C��^-��x��ϰ>�U�{��w������L�Z�6j��:D������|(7BFp��&�0��{���� �]P�	��>q��:�P/�Z�(8=��|�j��H� -l��e�th�2��$2*�a��h��z
�t�U��2���`��p�#�������
<�� �a�9+	��J���"UA�0�}���;>-x.."_e��XM�5�B�]�A>�V/̜d	�~f�TV�r�x�d������H�V���3�n�r[��Hx�D}�^T5�E�[�L6_�(��
�j{	<\�����'����PC�*T��,lt_���Ԅ���qUr'�֊lbV�"Y/D�����x�2�~\�#g��$�j>I�{�/8��1��"�t@�|>@t�"�^S����	���ɚ��;O���v���5$��MN���ʀ�& ��V�D�T~�Jk�灼��I�I�4P9�U[�X;{���-��ؚe������I����P��!�p�K�_�^�a��]���&߆эCH�>��?���J豐m7���8��(��́8E/��?}_�=/�F�DŜa�u�G�AP�Y��{y�M�R3�����9��ۥtA-��[����X�TXs((F���cⷌ�����ɽ��xș�L���`S�k��"���6�]���V'����	� �e"��e_�u��Byf�T�v� �Ȳ�6�5��~
��nK[J�x����8E&�'b-gZ�s�*%���*����sV��c��@Y^�d� Z8��V^���V�5���oD�O���ƀ/�򷠟}�6ke����U���I�Ø�2�1�SLiPW�}�O���d4��Ks�c��Oh[��kJ�][��hnuQ����A�|>Qz�#�?1�w~��ޥc�]��ؚ�A¸]�!��ƪ�i3��.��fۀ�rt\���OӐi_qD���	Z���P";����N�;9�K͋.��`lx����kh��:�'�6%���T�q-d��F��[�T@�0���`�a-�KS���^@��:2g��9��<3�^;�Q��2�j�A�Pj۵�|$q4�n��2��z&��)�������Z�(uZ�F��^����:)�Ћ�Q6��!5�O>�lv ?4/��xF��,K	s!O�,��\k����݉.��]��Z:��U��g�(��Ù����)�/Nt�L+��Ҕ
'%w��r��@eʐz���	��A���%�hCa���?!H��P�I��̄/+.]qp+��V ����"�RyH�B���c�*�� 
`�{�8��I��<ɶ�.@A}w�"���I����{ِx��@�H��-B �JV+C6Z������b�dd$�DLa��
��!aњ�x�u6~7�i�6�?`Ύ�Eߢ�Z�[{A�`#���Ud�0f]������>*�^X���p8FC{w1l�n� �^y�Kg28�����?d7_���b�: ��� I,v�b��G�}ܘ-d{�%�y��k�:�m@~�m#��A��� ����\�(����&��b�K�@=�Thū��9�9Z�FQ9|_�7�.5xAê�b����ww<��;�G�8
�e�J~R��s��'���Մ�-=S0����֬�'o�{��i{�d���nx p���)J�����`EVS�Q~(kR?�B�[��#a�~l~/��/&�:^e��W�����|d:�.Y_̠xS����{mC�ޯͿF��;��uGC�*wU�و Uދ�PFpo��k7�Eq�jB��IA�2����HV9��z�!�?�1�¯��S�:��[�˄*b���N�c+�M�	=֑�ܼ��6oێ8?g�W\ގKN��ȷ���E�OY��Az�j|k�#B����e~Z�~����>]/}����0!ɪ�~؊:g:�Clh;���� ��m��[7�6�Dw��x!��"��r��6��4@;
G���4���w�"ipC,���9: '��[W���<�,�4�`ٳVUޠ�˹6+W�����ަٺ%�j1#�GA��reK�rp()����)�h����G�b��%^����L�{������;�`���ׅ\�&᮳������{��"��b"�5����`��{�P�­� :'>Z����/$Ӽ ��N`��(�Q4���fq�/�t�|7�5��	s[����<�^�J�b6wj�&���ŝ�Y}��*�W�~wnfl�5��_.^d%����\��=���
��i�d� '-2�JI�P ������Q�+�b��0�/w�	v6�T֋{����$�X�_�g��}�'�P�5�pn�"Ĥ��W�\�rx�`�}v��s��UU�3,�z�g�k�rQ��'�3����.e/h��W��C�:��rX�}7���Y�Č�u}��)��~s��g�W;]4iu��lM��m%=�2�3��|a�#�	�h�co�ER�LGN���q�W��%��;
cu����UUK��G�I	Ʊ�*��n��(*�.6"���P�2�gd�"�||��6�g�����B�@�r$�z��)���Ǵ���C�e��)�i��8|C�Ugz���8�~�V��c���
�v�B����gʭ5����W�7(���mj�����������֫�V	/l?��B	��̱���m`!��ٻQw�B��&�$�A,N��X�d�J���b�>�k��Eo3��q	�2��&}ҞM�ޣ�<�6����<n�`�L�ƨ� �D�o�L�㺮����R��g@��9�N�J�}�Mq]�s$�!ְ��~˽A���=R���찢<W+�֐7dݛ s�1	���Ԋ��}�w�~����X |���!;'��0.RqB�~cP��1�&V��nߍ٣������v �a�{��4[4@�����%p�2z�&�����go�~�$�`J��B�{$I�����-�)���z��)J@Fso�7o�����En����JZ-_A�g���&�ېP�:Н.�F:��>���~��?�IN4u����i8�K��Z8�Y��$Z�F|e�D�͛�}D�z�2梍$&���� �c�4�ޓN������<���8I���O.�MԔ��H�tG���>�ʃ���ЇMp�����Ӓ�j�qU��G;	�������{���"�[��Ə�,��)����*e�������r1
ä3W�I4���m�QX!��W�]P,m�[aY���9���,u��\zJ>�7a���Ę�3�`ܺag��g�V���8���f��'�Q͛F���h��^��:|)B�3���q�,�t �rXo�ژ����1���oP
���F冉�w�7�)dͪ��<����NPB���cy�)�@�i���jf�g��x>5Z�]rh�w	����3����x����R��7t'���'Cx�ITL*"�^mp}���2�Xs�'KV�J����y���@���_-�!���*�)e�xRQ�7�&<8sJO���k��c��\�i��{!���l�$�ڳ��n�nq�9�+�������]�����
M����+����U%��?��h�����M�S*��yUW|z����`Q�&�\V�K.|7�0'F��
6� u���6Zu�[�7���&
�i�)0�����$�f7�]��B�[�:7�@�������]\=�Z/�?�2b�⻿~.U4�{�C�yNф=�����~��#&�~'c�( N�J:�t�$���t��Qv掀���!�k�`�E���T�4�a&��-�tU$����dR��2�]҃�#��iea$���ǀ�}���~S�w��:���d�I"؁�$�	J�M�@*h�8$4$.)C:(18��l���
֯)c� �B���M���`�3����F1'�����Bܽ{�$��Ԕ	g�R�5��M��|�sZa�b�$8b(6,��P�������ݛ�אe(��)qDe1ͭ����3,�zK�$c�"A���*Ԥg�����2u�-x𞵲���Q3��I')W!�����ȅHM6���0/�U�Z�}{=#<ϺU�V���N,����͆�z�њw0㴻(�����{F�p��КDZ��1%(�&Bޙ�R� ��p���s�O�U*������v^�9�ѯ� �%O��϶�,J�����L�bK
�d�v���[	'�1��)��7�/���3�ٿ,�q�u\�a�Y@�g�/�Pu<�>������u��Ҭ��ŧ�t�\uA�흞�+�����T����,G������Z_\�E6���.U�)�/����Nh�k3['�e�nw��cx������u��q+;{��a�ۂ�0��,��mэ_ˀs�A�"���Jy�&�Y)�wV��:T jR�EC���|:��H���g��!X�8�s*��\@��r��ף��5���G�BQ�a�mPZ�=����z��fQ�Ѵ���!u�bŰ�9R��(�E�b2 �P��	?Zh��w�̔j�u�e�$l��;���H(�d���]���k@�t���h1�t��!R.$��w�"�#K�/���w[`.O��g��ւ�[疕�\�b��f��(E�����>,Ì�d�vub�����=`����$���Ǔ��Q�5�
$���TOއ���ђsVD�#����e�JMWgL��с�.�4̧z'5! ޕ)7t��W��+'^��>��F`��qxzx�(?�\Ͻ¦F7 �Y�b=F�|�ĂK�9j�{����.�<������fڒȋ�a�A}1�\3#�	�]�酟'.�a��9D��b��ﰯ&[�2�uk���6%� m��/��v�?~*�|��``l�wEP�����V�y�@�T��
,�>wg��\��"x�:�����"Y{���F@��֗4}9��P���bN������( ��,iY�NT7u�oH}
H�3f)A������I�e�W߁������>� ޚiXT[���,~��b*Z~��Q�1���il������qǼ�0h��0��μ��q�:��7=ql��8z֥�Z��X?��I�L����J`���=it�R3w�#(MTD���־�{(iHA���%5F�ul�U����v�w�w4\�_�5!�ws	y���,Tה��1�+�ִ����~�J���O������B��?���	���Z'�����z.��{F�o/6z�,�c3��Uk��ħ���aB�í*N�X��y>V����*.����Z��� ��iuO�-o���xt�RU���Q���z����{z���'Q��N-�Z�ޏ��#�[������m�Ғ3����0:T!�i�f��XD��s�~�r�><�E���t���Z��n�i b��A�A�M�6����N�ƪ��|)��aR�E^k}�����V��D��Ԑ����.���j���O�f0r�:�N����P(:ZZA���R��8x��q9@Ai��Zִ�3߉��X~߬���ҹ?U����Cȕ3�(��Y����H�CR���Ʈ�����e�j��� ;D�o����qx�����22�����߹��|Fa�jq�o����0wq��T,J+�.�����'%Nxs��#)��/m�"j1i��*}(^:u����l�ɫ�:��?;���+.�m5W�n��N��p ;H[��q�[W'~7h_܂y2�����F�!����}t��ǎ��o����FI���|~�x<���|u
,���+h�-�،m��#}�-�y��`��PIXRq�';'��w�F���;P��e+�>z`�#����f��f�2��h#���_9�WC6�=���e�CG|�a>g�జ�x��e�̈\{g�'��j�ܜ��Gc8�������x���8�k.(��V���q�-�^���gts^,��y�:�im��89�"G�]gB����C�>�0ӿ'���zdr���]��<I��H���%��� ҒpԦ<��2�SW s\��1��{긯7���9C� ���e��Xѵ��8�U�<1���s^��gx�D`�f�� F*�[A�~�����N +��]u�I��a&��fqe��=�1k �0�����UV��#W~U���'�4RS�n2�R��������L6�X5�Mx����'�0���{ΐ�P/U��K�?�av���gt��y� �=�x��!@7�i����K
b���5k6��D@
�2���4��w�ը�v�2g�Zd�����׎�7~�1���RN���V�y
m��^���6�>;t�3�V�SZ���k�Z�����p/8 ��XF������<�p/(��44���8�`��=�;oP���ڸ��ό����y)����9�b��%{RJcԡL��������8𙞲ﴶ��gW�ʱ/!D�*�WV�ٿ���3`arǣ$>���A;����	w;O>Zf5�!}��dKį�S���0���[5