��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""½�c��ノ�!]&P{��v��."VH����Ħ0������<m�c�ǥDE��3ֳM��ڞ"R��d��<
��g����M�d]<0@�����i�Q *v�Q�aK-��U�q��`�nh>-E����8���G_#��̗D�--D��qg�7>��sYVN�om���4�G;�S��B�]�s����3��+ֳ����:���[�R0X����t�/8�����>�3��$�z3�!)}h����ey-�/ ���z� ¦�g\M4y�i���#�{y��KVY:PE�2����y�՘_���$��Oyſ�Av��9;�z �@����w�Gg���3�h��)�vW��xB�FW�ج�~2��$p>j�Vm>:r�ͩ|�+�p?�=՜b,����hG6 ��Tg��Ws�(�ߙI�P�(~�]N)��<������?���O����&��B�n�FWT�B�������'���j�����C�&@>�҈�8q̝1�3��y��mÉ����͸�h����U�+�#t� �˭�ϑ�qU+�.axkJ9�КeC6�Pv�6m����d��U;��S�ұ�����RI�Ut����~�N��AN���ӛ�m����I]y��@ŎQ�U#d�=r�V�N`;ܰ��,�MRS�K�8J��ՈK>��[^--�C���ز?�Xdڸ�Չ���r��sˢ^ͷ����Jw�G+�B0f.J�4���U69\�9� !Λ6_���s;^L�`���ݳ���c�O�J��!R%d`�k-��8�xe�Z�f
@T�Eڟ�v��Y� 1-�5B����j#��_��F��?�z*o8��O&=S-�Ή��I�7��w(rp��9C��C@F��p�&o�T=
_*����~�8��3g��B�`����i	�\r��B���iL�������"��x2���j��ͱ��^*��]�s�(,�N� ��R�@�إ��G���r�+��:bj��<�3B�����MgQ����F���a�8me(?|J3�@.I@�2J�20y�������0t
u���1��M�6_�Q�k��V+�U�h.l옆�j����������uv7a2�4��13����x[�Ӊ���{�!�"
�R+h�q\�v�oq.�H%�Dp5���_L8�bbSHƽ*X�:5�\�X��-�@	(l���ox3�SLA�qWf+F`4&�#���{��kDqϰKL�a\��w�<o�K��	�:7*Q�Ϩv�~v8��g'Jl���>2sB�3a����r-�͸�P���Qn�z\�_q.��ģ
8o���D�B>��Ao� �o��uލ�W{r>(���:[T-��U�0T㭿	$��O�$�$�����������@���u筨�����qB���kYK�&��_�{��f5�P88z���*w>�a	TN.G���Jγd��"#r�t��r�Dh���O��4>�5#n6��w�P(���w�6��ҋӊ��I��N��e«��f)-��m?�B��<�o�))c��_�Δ�J�����y]�\�q����d;
׳x�Q�f��O��e�bm�m���	t~���k&�Vq�)���QQZ�+kXR�X��X�w��K���u����jL��[�������� �0����V��ߌz94�D5��|z��]��� "�8zm�6�R��nՏ�M�uE�x�E;�s�$���"��p�!bϷ��ߢ���,Y��a�%MڪT��s�]���:�W?U�?�X���Bw��:��$�D	M�X�&T[DA
�7�b���Vh}�1�x6��K�*�e+k~��[����p��턽��_�r��w�$!��y^69`�n��ɖ%�U�P��|]OL����=+�Ƭ$ �{�)��p`��۝�1��~oд��T�p�:/:_)6�S'�;�^|�,c/f��x�`q���!p���|��(�P��EɻykP�K�޵�᪩e"�R5 �Pp'2ܛ҆qrF�������3�.���)X����9�撗|'b�N�l�@�uF>�����m�E�1xD�%�-��><�e�%�M8���Ĩ��X/6��p�+��������.����[7�hċ<J�������d�F>��%`�������b����6��,��·O}�0�݋���~k'k^��nZ=�i�D��U�*�y�[,�svW1�T\$��=j��&��%��tF7Y��d"zxg����
�uU���(�l�i����CW-�v��]�A�ةk-׷l�� ]��_��<���TV^���ׅ"56���=AHİ�	�i�?��y���C2�_ڒ=�"�HE*��N�S�ڌ:6+~�Ƣ�A�-�6`,�V!�`:M�ȷ��!���<�rօ�1����`J+GŰ���*c3��%�ެ�4�+�~&�p]|q�ݿ�W`��f��2��]Ki��}x~[i���Cj�Y�4�RK<���Y\�z*�ق�:g���@�7w���<l�@�yl+�\�pR;a�A�e�f�q�4��6��r�|�+�D�r�.���<B������BJ���)4R��>��������Z�x��i8pѰD7�8u�>��;�0BΪ�?$��RC��k^$5�S���VƯiD!4���X������Yh͗	7Tv`�	�fB��x�bQ�6칱l=6�"����xp��a1��]�����w0����<JN��3����LWJ�zeO�).��h ��: ������A������T�3�k�|�U-�	�|�1�ҭ_F_Dj�mр�;Zd.wğ�%ۤ fD�uG�X~Ȉ���)V��
@����q��{��[���;��P�sr��댐յ@w��V�'c�V5���RY����j���A�ϒ�Y�[��fa:���~�+N�3��HڊD&�@����4[j�q<����Y&�e��7x����A�5�B_<=�d�b��<`#�������2u���Xi4���l�<�̓��ܽ��g��#NWVl�yLۨ�=����nbX��)�'y4�tÁ"�|��ӋZnd�`�v�D_P9;Ŀ>fnY��	������V������9'[��ʫ����!������_+z:0�6[ʻ�Z�����5hӄ����@�a��t�ev�_-k$�ܮ��7~���v�n[-�#��u|0��>r)m��|2GK�ci0��#h��=�`7�_Bo�*�F|X���h��ܣ�[���01�vV@�t�M ���7gXk|��d���d�I�	n����%p���D�.Uh��5���CЇK�sK�>�3F��I��1�'tda�H{�ыy՚�TT6T�c�n�H'���	j[h�6����f@�A&EGu"Q])D��]�q�^(��A�A�	�%�XK/p؋��ȏE�/�b�.�O�l�J.%b���e�'�2c�Xa':9S�y�F�܃�2n�����*̸�@��pNVw?��0������-'�t %)�������[O��tg;���')@�i�w�H��}q�<.����Ms�ݿ'�����^�FLEad��V���m�Jr�6����L`@����_�'��G�����J/�j� �4�¶`Oc?�*n;V��=1ǼE���X�/�,��-LX��-�چ�U�;�[�#��X���uɻ���=�0��PnA�ov����fԁrK���\�=��=��!�Ѽ5[&F&��ۣ��H�i/K�3kA���g��j|\��1���;ՙC���������j^�������<��q���B�Q\�.�m>x!��.9qq�K��
�>NV�o��ȱ�gE��i�R�z��\#�BR�2�$͹�{a�صO�m2�)�Z9�(�vL"��xs>z�o���3}	�3�k���`��P�a�d�a7_��]]�p�`���w������Y+�S��J`6LNa�+v�O��V�xj#�g_�Fu�T����X�Qz�Hw@|��sV�q�)������N�"D�W��e����I���,.�ױ�Ę�B��ګ\���Lآ-�0t�0fz�y�(,�+�2^#��B˧��WhAqR�i��j��XB#e3�� i�4a��گ��I6LlF�S��*�9�:ц�m�ܫ�}g� ��=����~�Ŋ^C;c'�8��LȎBbewN�^m�0tw�]���n-�J�Ȥ*��j�Z꒪�c=g��� �ɣx��(2[��7��B�3ى� ��Q�ս��C�{�	@��g�&��2B{By�}��hv�m���o�xc���JU�B��ݨ�Yj�o2)Ub�a�g�\#��W��)qTvN=�mT�)�ɗ8�
��?�fϚ��7�����;���ԍ���}w�G;�W��{z�G6nm|�� g����H�o��6N0@�yuFC�Η�z4�|� ƍʈ�'u:��i�-'�|Fv���������ԜN(��F����l� BO>@|ŗ�4��T����TFr���:�B0�����2�.Ţ_Z��Y?�	Wϒ��,r������$�,�V.�g�1����B}��� �H<]{���̿f%H�J�p��K��W]~s�b�Q���I}Y�%�F�Rc}��eE��� 0�Ζwf��s2�h"�vB����oT�=J�/�x��l��D��0�-�f$�H,�LX��6�r��#�>煡Ț����k|�
�@&؝���5N衂J�r�oY8/����rg0�Y%��T�Zt�Z[�(�p\
&�a���7g���0�v���'Z�ǰ�R��2����a�/����ߌ�hd�̞3�uj�IbA 2i�t���ր�gh&�Z���f[uۥ��T��c�P�I�&<��ν��y��K�ic2Q��n9�e,C�D�볹�4��^�����#37�hp��v���>�v8���ʒ-U"�l��̥�����U	�� 'l�HJy������azьkT��(��-�1�I�������u�����!�`��ci����~�C0����(��0���%�Fm!bx9>�hI��h��$���~b��W_��u��%f/�(H�SwAиk��|M)���i?̊�BS��j*2(P=̒���o�-<Og��h� � �!l- �D�4Z���o��[����)� qz��7��I[S����$�ń���K����B|t���!��2��EGW�@Քx��q�0s����n��w�w(���_�����mhh�ag��q���]��xԝ�0��꧸m������$�e�[���2�C�G�����	��ا>�k.�|Z�u�p�Dy�K\��� i�t�2"'��:Gv�f��`�Z>d.1��Ip]֙�P���]y���:�L�pJ8�>��@�s��(�Jj�@�DI���x��>�����=z��'���/撏�
M���t��U�
��U��V���`��(��KދO�,�<���<Υ� ���Q�I?�u����s�c�X�!~<Kك2H�T�\9Vv�$sݼpwS���N�0�ռ�y7+d�ٚ��������|����=w���^cS�'�*.b^��&�x����D���s��/h�*�Y�QHmH_�)��]KOY[��OQw�j7O�@�C�9��?Ӳa��8W	�~E���I\qG���5.�G{L�^]�H����*�ؑ�0e�B�ǚ����?���|�P�̾���P�{��c�v�D<��QP-H��;Ң�ߧ�b�Xұ�T���i\B�sg�Ƀ]c��Y�*:���qn�ϔ����N�7�%`}r �>�h���h�������'�⛍~�z���G�����ͣy`��Ǘ
!&�k	�$t����h��t��7Ђ~B��ٖb^f��A�"�VX�YDYY��n�.W��� +�Էn���\"轜�`�9��ŏg�&���[�j��@�gWk�e�ګ�2UtwB�B���4��t�+R���Ǝ�f�z>Wc9��˵���ֶv�B-(�ߎ���`W�K��������BWv��=����'�2Y� Rr�:zA�������t�Py2Uj�&�VFI5Vh��4,�,�����~�|��ray�$�O~��0�w�ٮ���T�҅v�v��ӝ�8��μke#��6������)ڹ����O�e�M�s�,:}�ef¸��R�9��Ž���v�0�Ā�Ahc��K�$���+���8!w)�=�(�u�������J��T�t����'Ǩ�B�������]K�(3;F]�%q�ku����O�#���#���(���̗X��6\=PQ:�1$�ơaF���e'ܭ��r�����@p?I�bq�%�ӂ_�<N\��e�="檳 ��S�W$���̰O�f��3��w�v�e��ȘRNAᚠH�� G�P��s�8�zB��O@�3�2�35�� '�F��S�gT1؆��K�l��������nG5�.8 ��h���\g�H0����]�7}���n���Y�`y��M{\�j31��=�c�=�y{�i�������(�5�>�B����K�p'r8�z	��\o�Zԧ��{i4]8f�k����ow�{C��
�+��q����WzY���~\�����>������
�--8`|��R���V)�J�:v��V�a��Ȗ��ͯ ٞ*+5 �mVU�t�G+fn
:���ϱ]EULGIg4,GkQ=w6��
T�lh�D��7~�U�4�Dګ����C��P���D�����/���X>T�cI�U�g�b��l{��JZ,@t#:T�2"w��S��$��<w���!���G�
b�9S����i���6�C]�qFV�W��ͪ��Q>�Ң�Fы�@���4��46��������D60������AKAU�s�w��.�}��)�D�D�itr�.�Fu{�pR5��[��=����f�0�1���3QZ���S��j�q~��}8����yj�[������:�VU�gݜ�5�H��&'�4g��[nY�+,���J
����67k$�y��_�p�H�Sh7��;Qd�,P-���9�D�_�'dl�!tw� �D�ь��/)-����;j��qL�'��GgG��%�ؔ%7��gQ��M=��>�Tb\2�kR�ۻ��ԡKR�VN���)�5�	n��I� �$6�����c�^ �f�r�e�~��|�z�J]_�~���	}�cc{�ƊH�h/\�1UI�fN�(5��qµ[������Y�AN��fú��w��+��yk݌2k�LM
@e��9*aJA���<�r�p�#���N޹'��lP4� ���߮ �t:�#��c��<V�rv5%���u����x���xfM�d���x~}�I��.]�iήv�"�N�+\Č��qp�:FD 2�3"�U|5��{ΰ�$3����3;\/GዪR��vx@�d$g[|�
'�:�	��\�S����?��
ո�����J�><^��z�
f/!t;	����{abĀ�y�pj�[��^��F���QA��{�J@z���!td���NOs�|�c��
8�w��Do?>73��I��t9$�Y�h�tD������t�
��AR�1���OW`��3���^��L0�����ɨ��b}U�`���0����^�>��JS�|�.�h?� ûM���qї�p���!P�I��bB׶�nwq~��]�Z���B�;��Կ�s�^�m���?�P�x��o-�36��K£c:��2≥�.��\F��o B����=�P3���Z��]l�Vv��?�J�a�L4KQ?�wS	����.j����q���x���[׈�z�O�UT4�l�������AE5-I��qN���:4�|&�M>��l�S�1���E�~.#J�f'F,D��N�q�ӨN�PSyM��~-U>@�PYYAՙ�|�ΰU�����N-���Z��+���D��Ai�]+��v^�հe���B�~E�^nq�_3�go�O�>#�����i]��.ҼD
i��"�NH�3�Ma8t��Hz�
��VSl���"`ޛ�ɢ�Qh�,����RbT��cl?����+%N��;��AU���e�v�K}C�� ���I�����o�s��, �Y�� FL��4��AbU���ϋ��L�YNku.�IC������2�i��
����9��%8�^#O�8��*+�F�����N8D޿��"�Z��B�x!�Ċ��񀎍Jsn>�f���(̚�}��{G~��>ѻ�K1+
z�>�n��b�պ�n�*��_��@�5�rRd&M�RsH"b���9'��#�$��L:���?Yw�H����3��,�B������N�H�������]$J��&ʼѳo�SW2����,wk���t̫�?�~O�
��]E���6�S��f�<�*J���ٌȤ����7�^��)'���ڃ`�Z%J�zU^�ȸ5�2n~2��xr�-�� �J�Dx�9l�O�g~I��O늪��n5;|����Y[�.�
���#$c�`Ǐ�Ի#(RU{_�~�;� ��Ԙ$�g* ���I��A}��u���X��"+�&���JI�v���H��=+��Iz�o�M�̆Ŗ�g��r�|�L9�K��S���8z$6�Q���P����kmZ��eP�VZ0#�'�$�%��;j�=]M��(fj���"��V���Eس�,�؂�U����
*
�#�dN�P�.
������!�����b{�_���<����8���}��77�
�Vq�u,��G�b�rN�k�"x�:�3�z��s�~1cC��MPm,�ʐz$aK k!]������~����}e��A�eæ`�Tr�_Ʈoi)�2&������̒S�י�2A���]�+'I\��XTO,?c�8Q�t^l;��,�_�ePә$Y۝�kȞ�fRd#	׊T�P��ыĈr����j�i�6$���E�Y�w�l�vB�X��)�N6A:_Čwڹ1M��З7^v${5�j���PY�`�	.(d^����G�;��E�L�>���*��DQ{��.�|[b_�{�ѵ�8�"Ҷ���*WE��4�nH�ek�2zrZ)^��r>ׅR(�XZ�8�1g1��QY1�YÙ�����PKEVjQFG�\s����	q�KkR��B�/���2�H�:�h�Z?���Ee���ކ&��zB�dE�V�#[tu�nt\��p�t3��R۱��r�������ؾٜ<��r�����q�m� �����rk�KN��i���u(U%+�W��^u2	���a����M����ɲ%i��KϘ՘�Xݮf=�~z1l?�F�\Z�R���G�=����'Ѐ�m�J�L�MzX��J�"�+�:8>[�Ԝ����sI����#����&j�D�@5z�˛W>�T��˚�����f���[N`<�9�5��`%��f������)X��_7�m)?����\�"��*e(��#��3Ȗg�<L�"��slM��20�<��ӛƄs-�q��Zz7|8���<�s��K��m��Cw�=ϼnG����xF	��M4��z;��6鉍�$u����G�m�N��bB����*7�2}+�������z0TokB����.$/���E���.���
>���u
��~w�Ջ��t�ǐ1��	�9v��u���W̏��+.�|�)k�%�	;F�F�d5�[[K�qu	�]��M������#V�U��Ki޾����Z+\%	
�$�AJ�"%@l���M��8��Z��ɥ�
)m]�2!�\d(��D�s!�ƩVo~�1 IF`�bK�`rC=�yV��?S��1�e��7�t&]\���z�^�r�gFz�$�]&��[n��L��Qlh�cG�u���&���H�W�=�([qP܂�Y:)������:`�����;�"G�Xf"&�
�?�1�s4�fO�����SIò*�B�[����Y���?��zA�_��f��yˮ^��V�vF��Ⱥ��=��v�/
�n+Z06;sl�r� А��	�S�^O�DSγ�n�ia#��z�?��N�>I^���?C�ռ����<�}�G&$X^������`蒑��V����5��۩v�%A����������&�(;�aEl¾����UY��e�5iG�������X!�&A[V�{�kޯ�;n����hF}�u�jo���Vda_��C��Y�tVE�5�3�6!���]�
������5��𗗊"���C>D�[�r����r�u/o#^2�!Z%#;���,�Ncvl�\'�]�Tܶ[���LE58��M��K7���"Q��I0�d�����V�������w���_���&\Z\�i6��,�W��.�|��<�]F��0�m������=v�$��ݻ��*@'e�K �����7��o�x��'�=������Z�;������4�<CB���+.�j���h����k,K࿼��u(˘̹��K�8���CDG��9�Nv�D�[�G�c+�#[�ǭ׮���	�&���O:�m���u�L����N4Xv�U��n��Ё��do��.C�?��Ô(F�A����]�����B��Å��s�����q��7�G>V���1h�{�}������x�}�`���Zz�UdD߲ڟ6=���H�*�������'����1,oZ�/�'���W!�J���K��j[:YYax�cP�1�sNC�ʇ���0q)�� T	c@�D�(G�i���{�L�Hi~Q|	�m�gD.Q��ݒa�ӥm+9�|ב�1�+W'�/ �8���,qhn�v��Z���'��@"p��!x֦/�y�0�����m�{5�p��'/�P��Ĕ��LM"�K�n���Hs�WZ��YOW}TCv�K��;i��/�t���7�wT��%C֗`/�
�!�?BYL���њ���-C�֙)�V�������L?�42;�o�AƤg��Om��{�l,޾�itm|���
��d��m�|  ���G�[�ܒ�_��	1;X'����?�3>1�*����ZXQ�����h�
��^�:�7$֕��^��<^����H����e��'+Q8}G�c(�`����������S�^��1,�� �<��i~�����Uܣͤ��762�W��MDݾ8��E��6�"��#�88@�@���:��9]�#��W\�
���M�g�-'��M�k�{ �tk1�b�/�y���@����Gbx@ g���_f�i��������뗟S�<"���Z�