��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�Gf�`x��S�.Ao�vZ5��]f�(� !N��@�ZP!¶+����	�6�L��s��o~��x��hr��ӄ,Rf�H�����Jb�g9�Us~����`���d�Z��H����)��'�=t�Q���l�kגe�#��\�ܯ�����oI����T�EY��}w�&/Ф����y�͖�z4���f�f����G3��u�i<���*��$A����0o������ ,�~vB;9��뭰PL�6=�{$���	~I�Lѭ�97���O�{���v��9��sDt�%��׎���nfif���P�W�s�5.�o�4�Sʘj�(,(xn�h��𮩸�M�}@$Գ����)+2�v�8�X�o5�#�ɻ�,���gB��y��m�SdƄ��`���X�+���8�CRZ��q��8�/�8�����C%}��؛Qf�ji���V�B�R�n�֡=��{���[�ىS�i!�\l�R�X�N�O���~�G���K�dv���	�,E�呡�_�+yr�5�JԪ���#C�+�S_[i�9c�?�p�x�	��l��z�zd:���pj�ă��[l���RW��P~4O�Y�ܳ��\�� �a~��b����g_����������;��ðF��
>��A��P��p�
��Ü�Dd�����oR��m\=�v^p=�.~q����Ud7�@J����%A���1�8%��;F�bZ��Q�p��gK����]��U�߲����OAf�p���Ei1��M�����=�!�H��4�H�P��W���f�3���̐�RqJ�N:�3.YH%��"P~��O1�H����]�Ȱ��Z�_s�X��`9�\[�{$��	A���Q@S߁<O@�vvT���~_���0��m�Cv�=��때zt���q��_2�>Aϯ��s>y�<i��:�B���s;���Su��4����.����zj���ő�#�(���~G`��)ۂ]U;�Ț�����+Ab:#����?g�%�?���N�h��?{��V���E[3G�֋�;CH͹qP���<?�0P�v����ʩ�:�us����wР�ùGڒR��DX�����@����<�TLt!)��B�De����8$?K�a-�D����%z0�t��W��C�����.5��c]�M�C~��}�\�ص �+�x��T*�+����<?�(*��OR���Z�U޷F�����K'��X4��I��T�y���+µ�L"0�:�[q=R����M��Be*�m���sJ�ߪ5 ʳ��R��Ț*���X����8�q��B���?jF���{>7��	\���+�8*��jH`�wv��0�
�#�SJ����qA>~N���݂�"È���[9hqfl���xdU���x~�%ƭb�s|_�E*���J��sϤ�m�<����0"m��Q�֖"uT#����U��v����Y�JJz�{ɳ���]�۠y�#`��H(��x�;�8�r p[����̍M���j��c:@�@Oe���)3pT��Mk(�2�B���`q����m�g���T0#גT����>.<`EM�Q�ʗB9>�h��odh�dd�H�]$��3W[x�o����K�����ΰ�lL$Gm������+V	��&a�Q��a��&��Kom57��f����k���q5�K�D���^1� �K��2ɜ��jY�����͑�q'���/�B�%� ���UZd\R��觌��}�!=7�>~�b0*_&-����V��+x�%g��I*C�
�:�v� 1K����i=A*��/u��F�j}.(�~׆8���W�5�Y�5Hx֌�g/غ60��������Z��7z��gQ�8�'�Ǟ;�.�v��5���Ұ�e�QP�"H��	�p?C�`��b++���Ҧ ��>I�qL�
� LHJ��d��&{O�As(.|òA��}а�:Ә�4M����C#�0w�Iw�RQX���B��n��I��	]a�n�����\��@Ԇ�q�}��1�|���C�"�}���Q�U%ѽ
�P��v:��*K�]�͗��C��qw���S�M�>*���DGY���ϧ\q� ���͙��P�=���kE*Cϛ8>Kdf�E��,Yf�3s�B�j��y$�2�G����_������{l���-�$@j��R������D�ߨ�0\nr��y#�s��kǧ$f��g�ߑ�|�U�nR��=s	�w�C}����N�$6����P'rԥQ�����Ԩ�*�(�=
$7o�YځESK��+z�q��S'���x���3l.:��X.��6�`�zZ�n��u�[�z�.�t�V:i�N_w0����M0�Ջ��h�cf?@g��s��Ƅ�ޫzq��&V��Ls�8z�̘k�Uӝ�b�SW�G�K'wfL�u�P�Ņ���@'\��?M)�4u�f�ObZ#����>�#<��C���Ct���N:7�ÇM�$b�(��0���������X��az�)G۷��o��'/�m�H�e]���Q�|!_�� �>*�3��qY�.�ņfM�w2U%��"ʝ�1a����hS�1C���$����0Q]��h܎̐؉�&>R��Z�z@����ޅ[�jۡ���1����ƚ��f_����ev�o�^S񏶥Y_Ͳ2ɝ)�����^5K=%o�<| z��gӬ�9����(�3`N�E�+ts2�t˛��A�	1c�TS��y��q��x�	^�D�7q�{��U	_
	���q]�C��Oo	�Z�f6��H9l�!=F[4�������_��آ�n;ιJ:)�=F�E�p�_}B|��Wt`+8E��\zEP�%g��<;~�N��g��vr@+ޑf?�+<u~�[�B�����RGryc����-�Xx˓Q(�Xo�Zp�~���w�J��i����h?���|z'
����F��j�� � ��3Z��l�0��we��I��M'L 9��9drh[�\�Wo7����`O�Z\a�-?�	4�5m[Y'�ʫ;E�ƲT���'���W�'���'-�L8=��E�ժ�=g욒9
p��2["�����A�cUy�[�"������}����i~�����C9Gv/6�o�yj�k��kj#?H������vD(�x����_`����ɏ��_@�vrRo��V�Z8t۟C��jA�+�`
Դ��\$�W��;�;����+D:fa�Hy{Lm��~V�Za�;���z�U"�SQ@E����*:N��0ct0��-��s��';V��`�PR�w8�hz������*)�&����� Ϳ��c��n��)�lKL��>hś㊍���=�L�&xf�;���s�i���iMyi��/�<7�������uB~�v�p������_�{�C��-�H`q�fۀ�Y��0�DAJa�1�ClQ�	(����%�`��"���Zi�Il�/ӻ��"ŏ���-�;�R���$���+�l�(,���D��=�g�Fv�_���^�6�р�wb}H+�38�{��p���/�#_�ƒ��=q��c̫�S�Q�z�����Hb"�oL�Ec�{�_��KT����ц�����I�� ��o�4�N ��k��O6�ꑠ� �'�e40�BY��h����
kxgU�����A�yx�1�sBKq�j�X��Z�/9'�_x	 � m�jPRE׀���	t¥��,7wj�i��$KW���o;?����@�QL�\��s�O<G8IU?�ʟ��SԌł'��X5��To3��m����<�SY��	,6��t�	a.X�ϙ��=i���/�30��Ա#/���Ա;X^�Ez�9�QL>�|)�k�y���>�M�)�qrv����wnt�5O���F�_�r�I~���M?��AۜP����V� Vs��t�_X
��ٰ���Fd��X�|ą{!�'{o�.Q@�~e���֌�������!F�o��ߏ$m=�!�n�u���Ψ]��'��j�����v#��)y�G^�	�FӤ���c`BQ��D]�E�/W"c8��0����[l��w�ݷ��3<��i�&(ר�2C����Ğ#��)�4���4c[GA�]jX�����K��m`.`O�&����D�z�j��GU�d����r]�KE�kL:R��W�]lh� S|���V��)x����+Е0>�ߜ��85 ����-�d��y�mI�R�~��P*� N���"�v�Q[3�Ȕ5Q.O�3��4��_�(���5�}7P��x7���hDF���E���0�3��W#8z�m��8�?/y�J@!#%�c���9�\��]~�_;\V����� �D��Gm�,1G�J���ɦV��,�Ͳ(-�P���ʒh`n$ш��&��b���]�i������o�2#�+8���Ez��zSS)�6�]�ɨ��)!���b[G��Y��	NS�]�w�̜˨��+�$�}�����SH��Œ��o,s�I~�I�Md@�P
�0��D�|7���$�#��5�i�'{#y����^��d
�8@)V3Y��#9"�hy*T0r_�[�]���%��<��EQ�)��c��e3���Ȓ��;�W�E��b���3&B�����)U�$�������?;B_(y^l]99Lt����A�7�!�O��媬0�}�W��ʗ`%��;��`�Qn����d�Ġ �m~	��0l�<x=�kE5�̃ /���o��s�&��9�u��g��;�n^�4��WN�&�IҊO��غ>C 4���m���oێ�tx�3���~*R_��/x.�R�~���q羣�Uo4,�h��X<�Tf,�h�Gk7$$� �U�NƇ-���\pm_f�&D3��`��i?�)t&ʕjI��܃��P#��߬P�>KQ��L�xQP���-6;�Y&��;�7�R�z5��bMFL߭�J��F�5��E�#�����A�`�HM�Xc��w�s�y��_�$�a�W�3����@;��oݯ��Z���;ؽi�>c���u�܆�;���}�9Ԉ�����x��ن�C�$�_�K`�
��'�ҷ���=�	J�j�p2����;E ϓ+Al�oYZ/}ƚ�
>����(�LG��n�d8�+��P'�v��AȂB[�^�W����$3��H�:(�a��0��������m� ��h٤�s�Z�f�q�%��e��=��?���,�ix��PM�;��۵�O�~�Wb��i���Db��ek�#{��R��?ꡋ� �mC�����dᡔ7(�(*���T����L��J��ӋG��H��@�l>��Л������JaI<�]����u�3���L�b`�U����%���[����<���+�%{qK��Sd�ȣSO+ �N�`o�kd�q��J������*/�*�r�H C�Z^,(�m�L5v�s� J�x߮*��p����\��{@LÙ��ɚ�2����V[��cV�U�u2E7:�F��Q˂��j��`-o|���H�U�5H��@�x��J�2"Η�#��g��	Ο���h���k�9��ڗe��j.�i�<���䵁d*ڪL�㶅e��F�nl�=��Z�o��gfvt���,��_w4D��.�g�����Lh䷎��粈 י�k�z�Q�g?^Fҏ�l�f�);�%5N B�X[��7�'�A��������4�C�&p�3E�f�&� !�!�2՗�r|��Hܫ�����������P��ਘ?�c��$�Q�g�;4r�5���v�S��XIe�!��9�d\�N���]��IA0���%Y��A��
�,�=�4Z]���Q)
( �S�L�D��w���5��I|��Xؕ1V!�~2�\+_<�ٓ�B�;_*LZ�wV*nJ�=6����ȯ���������������+�L&�D5��z�o�����a1��W���{�"|
CgH��O�'�+�E7s�yv��1O�\�����w�VG��"�ۑ���3odS붝̥��҂��υ�l��,�E`�Z���C�
`]R�&6rvz�Ʀ�(�(]�;E@R$��_��ν��En�6����Y�՛m�-D<1�<Hp+��+�!���=�A�����w8ߟ�����%�Y�;z�n @���k�'gt�݃�b����xC�P?�Ra+�3�3���T/b&C��޶+q�,�O_XI�TI�L�8K�'ą�kh���v��P5W繶9�I�JGi�[]"��&�VB��'RbTE��Rz���fzc�o�b	�nF��V�i��ڹ0|�lc�g#�L��/+��*`��:n�X��9��'����df���y��Ӥ��z��˔��¨#�b�E�S�q0-l�#�E��"=�����%� 8� ^�>�Q:����������N�7T eYzs���w�e���8���+��Q��jy��LtV�Q,h�~iõ���~6c�A��<]�/�<g�����Ո�4s#�P�j����� �y̫�Y���cK�w�J#2��~��>9L7d3�|��(3dn�R��Ģ���Y��{=ۓ\�"Ӱ]ŋ�G���w�	s/��O�2L�!扛��^r����dQgK���WA�ȤВ\B=�FC�[j�/��|zl�z�,�W�ϩJ�Z�T��<�8I���<�_Z��$�c����6|ɶ��n#vD6ߟV�$_}�@+<e�%�'Ú���Tږ���1N�=�F���[�p�%�r�<`4lna������C����F���"84����
COB��w^j�CE�&v��9ԁ�t˰�4P����F��)�_��hI��?d��d�o��iQ�\�?TW&0C;�PM��>���cAf��>�V��	ôߓ3*4 |�O��a7�]j�y���~��#¤?���ӛ�:��F. ��8Oٞ	a����o�b�H^��oF�n�8��R&�_7��qp���M'�YR���mRd���fw#*R����n-\��Pg%�����z�]0V3���:�.}�B��82��ԽS����C�1��&�����_7K���%�Z;v�3�e�/�u�[�lyK�)��O�m�\`%H:;�{-�}A�OipN��]�p?��a�ۋ��_T�J��9<��W�:�~���O��²�79���]�����������?��}c��b���~ ����&��]]��k�����rR�0+��:� �SK|9�r@�{�F��6�Co�:K�#X�ͧ��f �Hŀ��)�a)������(؂ʰ�f4��N�/�T	u����O���ݟ�����hT�!�/�#,.Xf�e�U�,\��>O����2��7��Av�*"�]���X����9��L�L)?V�\��T��j+Ә*��6&��4�*�N�ۿN�J�ȝ�I��YHPPٯ���<���P!ZǻXp�cBn>IF �ꔃ5����>2߽W���/E��pi�љ(��hn���Ff��!��r;�#�wۅz���������j[M�/����ȷ{([���ɸi��QRKFJ��
�N��]Dy�w��l�Ll>��M�	�w7x�y�%S)A�Q^���u�u�����ќ���O��@r�iI�*��
aKjb?�Q�Ln���WH]m�~Z��i���l�6e%"�
��Z�ڡߖ��m�N�n��b-�xP��,�bT_�i�s��$<MΚ��â���T�tFWd���}�����)ۄ&����Z�<�y�/Hv�H��"BGyh��\�����4��<���)���9\�L�5��_c�$ȼ�嘘;*aވ/�c�j�����"��z��h��ο�x�4f���J�{��]}27����n8�d[|-�VL�~���%��'rn16�Z	�Q���@<�I��z�c���@�/�s���O1Y� mD�0lx���C�RS���C����1�H~ t��Uf�E���ZCs���{v{j�0&Ǳ�$�VU��ߝK���4��{�g�-��E%x�F� �̐W,�y�U�In.3��Y5��oO��-@����-��6p!�Ux;�Ē�y��^e<�P.�TvP�f��gi4�ekeҘC�|��\��^�*LH3�E62ڨ�������rk3Q��6��.���3`5�L�F��R-����H��M�u��˱�˱�L�č�SKA�%�ϊ=y�b�`^�+�1�S{�����]Xˣ��WrK�:H��ڻ���8�B��e&��K����0�a���ANu7?B���ʑpN4!;�%�����]WƦ{B]���,z_���Ϟ����\1}*��/�f�Et���P�qGޖFX�����Uv��2̪�г����g-��j���V$��em��l�)L�W��&�z�C�kĢ��a-��=��������y������z2��LK�^3;�uq	��L�Ļw��d�������2�u�y:��+��}��|��+-()���o�<�R��I�����+� q�+���"������ՑVҌ�U�F�o���V�f����zK����S��-�_o�V�c��<��I�Zu~?��"�3"��z^*9}E�����W4&a*��m��[�'����$`n�k�
qu��*��J{�ȝ!%�a!��򴰣R̠��׫�����,t�����+�7W�G3�%X9KyZ�/98	��o]t:o^0,Q׃=>��P0�1OF�uĞrZ����Ѫˮ�Ljس��ͥV�_/�s�j���7L�лg.8=��e%^,������)��*H�G��QW��8��}���Q'e
����>�l���,רE#j��eĢR�H��zBL���r�m��b����EGX�v��9=�����z�wv��&K,��Kq# |IV<_7���R�jD�b�!>%��ұ���G�ג�V�_�X5�(��$���BN�4�;��H*S'�ѳ_X������o<fa]����h���^:�6Fi;'x4
����;̬I^�O����%u���6�Gj~��z��7��3����l���s�����<���1��o�%����K��ƪf��"��g��ejN+P�ƔM�UI.M,?*J)�8-Z��Ket����Bdڎ$�?n���d�"�Ļ7R6��:贀�pwJR@sU�>v̚C���g�o�����ǉl���f���7����o�j:�ղ�FGF�K�g�O�
nE���ꟘF��Oʴw������������ь�ePi ���SB�[�K��,�	K�n, z�w���C�����Vy�j��$��;ԏIc��m^����f�M�Ս̈a,�1���t&�Dd��گ ��Y�ŷ��b��w��#sa}%��ES�Ez��e]�7W��nM�TI��˻`�?F��/V\�1�
�2�0�n�8�v��	%~7�~�C��߻sq�Y^z�R��,�2%�^=�Dt�
Cj�8�����MhF�{�~���*N�e��A��8���l�&x�5#�ܘ�.ȴ FS��t^Y"W�f|�9�`f�ߍ�pԼC�
�9!��s�x��Y|�@.QC����0�-.������$׻�p�Z��@�d3i���!�%�e�`�Rs`q@%r痎P]��Cl=��6��e6�Ľ�3�j�3	8+�S:v٧��=�*`c�S�#���3����I�H��(���Ǩ;���m˟�jV,r��z�F�~�� ƾ8%V01�bu�����k旵;��)��QhDucy�6c�����D��r�{���O��4�?�/�З
���g���9.��`����}cU:%�w��Qi�ݬR9G&|>`-.w �(U�CtMV_f��R9꧑\T+:m��g��4g�V)]@\�#�I:-*w�}�db�N��8@О^�]AB�"l�[rq��P��<��������e�y�)-Jܰ-�|�М�ڶX׮4;����5@�x����?�A'e�fH�<'�-�����du�!%8���������Ժ��ٮ�����Y�v>ů`��5ϥ
l�%��w�d����)��gM���������KN�B�`��d�s��+ط ���G�I�>�U�!�M-Č�\Z'AK;A	n��w��v�VY��d�QR�Ԫ��&���r��fuL��O�U˴�H���^��m� ~Ŕ)�M�IR�#���P�����v�9�P�7���q[�j��Vm_x�����H�,y/�6���m�g��M�޿�h!q��1 ZQ�{�,;���j&�V�\���5�	��ME(x]�;RU��	�=��wn��CD��n��<j�[�e�T[��As����-����F�O�L���9/n�AnH����TE,`���Z$W�#�����6���:|oQ޵}�+�'���xu�������fÃ�s�zi�!���gAGB�']�u&�)�Sn��!��4k_�`_ڔ.)��E���a����V,