��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>����rhhm���%�ñ��\X}"y�GM8�,�eP��:h�Z�{|��L�~�t ,������DN�F�	�:j-��u*�zn���{�h^���C��zlC�Wg1MH����{[�rx&R�+0,@Q:/��ц�?yU��g_b��1���C��M����훅�[�>F�?X�	��ϟ�]w&A���E t��/y[�x�b���튟Y}
�]�w3cGTe�����F;;�A���|-�¤��^�{�w\e�+����"-�v�E�`iӆH��n1��Z���Z"9߸���֦�}Q^�t%��$w��=6�e�C�?'G;n�F� O�9�Y�,Q���X^��"�p�񔺖�3ЄQ���W*�'0J��kq���>|6d$j���V�+�{��Yf[�( ���_��qd�pY�o�4�8h� 
��ɴ884�|�?����g5�9w=G�۹~B>m?gU?��f=������W,M82����q���@<��폶U�ټKq��s�sFz40,�t�>&΁��Ã���Ǟ�u>�J����<�<��A���s
_�m���8�IJ=�;�Y��H&�Z��CȼG�o���?����\QY��H
j�&��y#� 14țJ@�:���!�ȄS���`�nҦL*ɈFC�2g��T1��d����?z�ӵ*%7�P�82HO����Uϋ�։���u��'#1 ����=Ki�`� U'$��0+�Yq��(8ّ�=/�mN��fmM9�r	�	52$aƠ��m�q��6�/garL'����8ZE�1u��e�zh�]�g��C�JT�h5��
�#A:Iz?���Z]��dN}r)￻Q$��?�)��gh�I�����M7�Ve�p�I�����o��!�s�2��A	�Y��Ս^��/����/¾�R����B�3�J[$�tu�^�[{\h{26;�_��(pz�2����ʄ��k��f+���Aͳ'?{���F�I��Vʁ]��r��]}�s����Hm��b�B��j_w�\�X�Q��_�E�J� �@t�|ͷ㬷�R�!���C��о^�؃�U�^�|p >w	!�������Mq��Y�5�^�P�K�pT]\ɉ��S���诱��e�V�+�>ݛ�Z�O��҂���T��QX�$��jW~ƩbC�Gh긪�-^1�<�d<σc�k9α�^>�� D�v���Sm/�	���yTSGW7<^���˸��qt��b��}�|{ΖSf�Q~��164�G�\�$S��
O��?iҌ�mw�:�@�yE	�>+��������e߱n���S���Q���}�G��մ� ��I��}���L�S�mw���Mp��ܮ���ƪ��:�Ktp��[en2�܃���7���[Ƅ�/@� �q栂���[�����x�x���Z�[	/ĤJ�5��7�4��4��M�د�fMыX��ۆIC�՗��S �B^��;
Խ���$ېyr�Pwa|l�T$nhha�qN��U��k��	�\k����X1�A.��"F{�xh׋�
rޥ��U�����1����}ƕ�4�G�[���%�Ȕ�&����θ�C	II�)���U�OT�����SէĦ��f ��ji�()�a�	̲S���u�h��gZ~_&��q�$c�	�4��7tF]����\i)�_|�0U$;�~�x���֘������EE�]��컹�L)��9�תo��b�Fxȸ��r]�|���[�	�[Β+�_��ԑ����i���DV8N���&Ŕ��F�T�t$U�o���\�Jn���Q�ȑ�Lfi#���տC�%p_ɍ��&m�@;O~�(.���h�h+��Wdn����QEΣr���|G�؜���O/ՄE��ǡ���k����"Y�����Q��kg��J�D���������Z�r�{\��Ag��� �,�u�41?a�4[A�L��:a0����(@���hS��l /}�WZkF�$}��9�*��T����O�M��6����\�t)���(�0�i�g����m�2|@�Art�	܂&@��G�x�60�f��>"M,��t���KĲ����r�'�8����t�N���Q�$��'��o�<v�ȕ�a���B���tY�Q;��٫�H���r��������*����ҹJ��]�z�h�j�)j�)Nd L�ue��Q��^�a��Sc[\?�eص�S�)�r�F�� ��)��T�l��F�*���Q0v44��<~ڎ����I���_�8J��_�!R��)<�L��ڟp�[��TYo%T�ϱfs�J���U�I_�*0���C����A;�w���K�;��I��*�CWK;�'${	cV��!�6�N!�;�'������g'��etw���ۨ�}��K��mF1[�ؿ)���QNa��6Z�;�0뻚��C������T���~*B�fc>^̔�,��#{�s��\�Ȫr!�}1l���n��)��/���n�,7����8���kdXB��R���_���>��@�t�V�2�
����A�`7q�����L��͍
=�?]����X���%q%����,���+�C���G9��|�`��h��������"S�R����K<rV�����Is��2v�T ��~�x�AM�ݽ� u�>Ucq�s\����t��=���|�t�I��,-46�G���A��u�QÍT�	�	���	p.�s</��-�a�s�A)�yx9!��֫+�����1�`�&"���[�+� ,�.�7*��[����PK"�.H�I��wb(�+����� L'JU������0E�7�>9QI�����ܲ/���0<��lQ�>TͿN�W�д�Y=��Es@�d��ʌu#��m_V���ߜ�p��=פ�H��_>4������B�ݏ&2�^>�����T�jG�PA�&lRz8�ko�oI:�?X?��j��d��[��I��ַ�!K�.k��N��b�6E8�\.;�WM���:��d���.&r,E��h4t�z�6�N�H�n%j��	�onIX�;CoE��\Mt�O@�K��&.IP��h��@ANA$��n���W&Q}/k�o&��%�]��[�2*ʡ�|�B#�"FWY�a�\���,8P�W	jj�rQ��9�&(�d��6�<��0��r�Ԇ`h�O���^��{�fSJ[�9�k��@U&�ݎ.���f+�:qLR O(����3Z7ƈ���µ���q�0\ ��zJ��1t����I�I�<3Y��d��o�S��<�)���߿�l���������2nhV/��ݔ�4��v�C�[�Kd�,���-������w���q}!�j𠰒7.���<<t�!��+y�����Hu�7�4
aZ
�@*Þ��/��Б�A��L�q�J��_�4
 �M����_�{~�u��`��8<�P��:n^X��Ǵk��xd6E7NY���^��K����gW���
'��xA�H�;L����NòV7�Y;��}ǁ����H�-�hm����,v-exM&�Hh��Ϣ��C�tQQ��>�	= ���d�Z��0H����❕�X?���V���8U�&q��Z�PP�g���)�!P�T��(o޻�-�=�G�|"e���]rUum(���[���L[���W~��X����M$�c_���+�?HQ<�Ur���Wj1�&��b��&�iu={+^��e���vm2Mi���@֛�oXg�]���J�[]FF�`�A�q�0J�q4$e���b!Wa���|��M(u27�1yߡ'wmX���p�u���w{�3ɻ(�ha+9s�~:u\�>�%���M5���2�z�Q�բ�I������`?C���=�3�ݘJ㠃Ԇ��@9_��kI������d��)��I�VkE���%�-jG`8�1@�>f[�����_��A�3�hۑ�ShR�3���j����^�a��G�[�����:���}�������&�����q���� �Qk�^�Ѵ�ϟ��O���J����ӝ��e��lST�=}'	H�\����Bx��yG�씄~t�/�J�����P�[���{
1��S��l&b�VoQ�<�poZ�V����V�h�-K߫P������
����f2���� �ku���OY�����W��[*�~��5��j3��s���ڊ��)*
�;Y�+� ��i��~V�����]��4 +8o�'��$��gx��E�mM�e4�f(���n�h�b2����Y�F��xL����B��$�`���N��A�����|�����0��|!`.�\(a�X�|��Y�H_};�]w�+�����*dM���a�~L�6���aֵ��D��ua�"a��nh2�K��':���χ%����������K���q���B�A���mȍVMߩA
�2�mc�/͉c�r�����,�s��>k?���ά+Y��������_�_��zs����� qB��/�x�T;�}��H&�������:�"6=��gA�q"E׮R�߭�5F��:��I�M���;VǶ"���5q�א��aXc/ae#�)qv��U!y��,rOq�1����V#d;p?��
fHTQ5v�:�CN΃x��L�����!�YV�@��L�����1�O����I�'
=v�'��P�<p��z]���X���D;���[�~h���x@z&]���H�齊s`
4(�p����?�3eݣx��Y^��(z�ɑ;-�j�o�+c2=����� �R����@����7�ocҊ�;-�z��O3ݍ�&\���['�uk���ff݃�Y�T��k!	�Y��m|X�؜��z�XZy8�'���\�.�h⣕/#����u��<�B��wk\�o�Y�UU+!�G�xO���TIM��8�����.9���~�:�~=pz15C����A���R�i��C!�Ѹ�sM��#�SN^)�N9�Ҡt,R�f~q�G�+�"i�u.�|�w,,n��P�(?E�+�_�ܾ�C0��l=z�n?oy�8{{����k��z��+�*h��6]Pd3�yT-���������8�D\��C4����D�D;�ؽ؜'�a�>ii��m[�2��`����u�,����(� �Zѷ߳=��%"��1a�>\�\ʶ��Td�?�梑�5��؅�NQe<o��������ʟ�do���H���Ug�J<�Y�P���q4�c�Y��&+6��NOl�ܶ��&�_��2�G8�Z�R-]�l=����@,�Ld�DZB����@�>`�G��QU���PAoV0��9Ya��h�՝*���攌�ˬ�-z��x�aw���-�-��(
�/�y��4�{y� ���[ҊTǇ	�O�p�,�Ȕ�+��cR�5t���A��Ͼѹ'b"Cg&r3Fj������$�%�vJ�{<�ւ7�������Wä��UI�|�1�kԙ��@���&�܎p���
%ߦ�9�e�d�
R*���i �&2礬j�c�@�I�d����75�h��l�iΨ��"o�_*)2��ƹ��QO��ߊ�1���p�c�����ɆаP�D�қ��ܒzZ(u�jy`��	�'���sMA�z#�hlbnj;q��PM��B�
�E<�$�DP~/3���"�B���l�$�0;W����u�*�<q�P�����pd훲����CN�%�H���z�Z�
9Fm�h�Y�oڌd��\�6B�97t��]����7�Ob��~4�w#�;�g�6&ñ�#�"�%����OK����@j-��<��f��	�ja���n�<�2>�ϗa�[���3���?+7�d�'������l�)�Zޘ�m�6�ՠ��Z�o�T�r��[L�����q۱2���U�b����eWU����3���İ��7���}�1L���3�u���J��9O��GFVw��;�M���_���@�ś��bމ�p0zS�~Ww��6�PC{�'�[*���o���r�k�9��I�v"�+Ǚ�<�}G&� �vP\bx_�)�p�Z9.Dy����\"+�MFW��z]%�=-�Ѱ����v�rU~!�]3�.��h�؏Ծ�(F����o>����=7��XN�xe�UK���,�CeM�˲͋hAg���aq�t^|^���!sK�ct�L�����
��~ESP�j�j�a����+Chf�&�2P�W>��X��yP��X�x���]���m�̍37.@�ӭ�RC+ʗ�����N�^E=k�� B���eLK�m�	����t�;�������y�_�����D��r�<,ű�EX�k~�ė��װ�H@�����>SdW���?����e �J%eJJf�T"Ul�}�}���w�[���*�'�Z��ao\��V���7;`W��б����J>Oq	)x���8F����cW��"���c(�1�j�@{M��ڴ�B$��*��o�PK����|�Z���j\��5J�g��z�mq��ժ��z�@q���(Dxv�c����D�e,\��,�p|m"rZ�o~�����Y�=�2!�W\�l.�'K:DB�.��@�Qݷ���OG��w�xw_� �	+��v6�����R��sMM /6��{�=lɁB��B�K��	��e�&�n�G�
*��1��\v�`��Vb��n f��>T8�[9vdH� U�σrt덿�ce�;Ӎ�pf����rD�BOO��-IfK�D�7z�_w3ЏΊ� �%���%	����NS��N������B��6Q��l{#RE󓩭�}��n��<��3:R���[�2E ��f�\�H�Ń�K��7x��fo�(��M�Mi���R�U�&���g�a!+H#�|�&1F�M8삍��6�lp�_�m�bE��kĈd��]��V�.�g���\&o�i:$d��o�����WMC67�j���:��,?I3|{��yR�q"���AFoT 9Q��;����L�������tP��f�m�
Ģ4��#�r�q�^��2_G�I�������~�b�fM�=�R�;(�*���`���B��[�)1O�tK�R4�+��Jm�L���K�cPH�?���Dsz�@�/�FͫD�����}����e�q�^'y��xǻ�O�jߺE�K\��t����7ܯ`�����/�����]�@0�Bk%]5�<�Ȣa��#3�%�V���'����	��[	��d���ƘF�7WE��^��,	*.-�/(��0���+��}4�ޒ�򱻔$����p�w^�G���o�դzՁ9�g�����7\ T�_���?�Ia����k;�J^S�@5�Y�}WЯV���A���e��O��0�@�ѺFs�^���	*��B�Z�A,J�@I����z��#�A�!3�9�N�$��|�#89�_):f�6¼�K�Y�����u�mj u~�k\ -.��$'w�4���G�Q.��B���]v<�(	�B�Ϝ$g�R���ڇ��Y�$�s���n�}��8x�J��Z�oַ�)a�����=P�}��V��v��`T���X0�I�M@J��T��S@��OO�L���×�u��җ�����sS��Ϯ4���ӭH'_�i5�SP��.��P�׬nϽک*��w��t��� �A���F��Z�i�jˇ��t�Z�]ǘ�*�?�~� p�����Y�8Ne��#�f�5��췧|bq�K�	d������$�jꄋe���퓁�ɂ-/ ��{��3'[��<d�"ai�4^�a��"^�|@U�B�N::G'c@M* ���ۋrź����{��rS5���L���&���I���hi8�K�kpH+