��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]G���B�X�x��x?ь�¿Y�ij2��}�$,�M�?�_[����O�D^P�ώ'��PJ�!�}XO�+��7�xЕy|fzc���wN�h�M&�]*t�p]_�-r»�nEK��,�����n��x���k��p4�[
�-�V_���)}Buhr������m;?���9����շ1[$`�AL�'>q�d)��Cb'/�.s���٫�#�]ǎ��D�?x�L�+�ʤ���i��6�[Ϧ7]`�-U�b���r��qt�F�Pk)�6g?��x�ۑ�;�iB��zE!�ӡ���TrԆjv,�`�2��;��f�&$)�4v#�!�W�
��a��ū5��ϐӪd��Ǘܰ.2zN�;�D�͋bX'>v� �Шw"����ͅ(�pq����,sӀ���oM���a������{W�o焳��\�霩�{!��΍X��R$QԬ�/�t[�R+��<�����J?�e	f���]�����C%ED"�R{���B�Cڛ��Y�J|����N��	^*s��H?����]#��<V,��#���E��'��Q<���~��9��7�nt/'�KcOjV�=��t�����_wn����v��\<����"fQ�ە���C��(4�W׏Ԧ;QfE�3=����y�"���eϣ���W����n/�#��Ks�$�r�?�|x��g-"��N͡�ה�l�TR�髋����6o��a�5��Тy5�������u�s͚RĢP<�W�8E��#b/L�����iٚ0��㭵�}��k�'�6�t"Cn_�D�Q��]��Dp!������^u	�K&��=��М�Jy�2���(�+g�������R�C�>'�<}d&��X?hF��\ߥ�O3NIw �n2�οz���v��P஀b[���RsGf&�JM�Z���̛}:'"�BX4!��}4Y�T_p=7іI��نm!W�>XC $~���<���@)����D��euT�[m+3��5%�W7�z�~ ��f����6 ���œ6.���1���t��B0�b����,KNWe�gF��@� ˯�f]��dV�%��Aˉ�^*�|xzP|�,�&uo�]��W�=&��H$�Wg~���hTHI��m̡�uojo�:�����ԋ�"������ �d��ɗ|����LTL�Ͳ1����o��ejQ6+�Џ�pq�y`���4[���l��)R���~:�a�BRk�g)ɰ���]ٕ���5v�t�d}�ӷ_Y��N�ķ��.�%A���t��Gܫaʏ�R�n������ց��"���VDB���:Ă^LeᜌZ]��H屛���& �}�~�ܤ\�m��wɁ�ϫk���+K<*'@ ����-�:�h��د�̯J^�7 �ڪuA�(;$@�\Z�o���V�x�T�:��ͦ�
��Td%�VL�](��7�@ξ��]@-I2�E��A� ҆I��3X5��x���9(R����P?����p�qfD�݅tuCy��PD�h7Y�h��/���Wĩ���0��G�v�����G��C��SO����u��j�L����8	*�o�zB����!i�Rc�S��{�Ք�=��oU���~��X��N�;z����4�>�9��8�U覧(�B{���X�x���<r�xu|f��>"ze��ں~غڲq�(��z0����b\�2<��	F�h;�?M��4�F��2��.թ;̊�ˆyw�>k�6��ԒZ�g����Wv��G��C�Q��ݡ��+'D�$��,����k��vu���f_b,�K�1�n�-���R+�ksb�"������vޒAs�٦'����}�LQ���\��.«{�9>�]}P�^Բ�^}�sD�}��i��j��F������VDh�ot3Z�X�U��^;8��ub���=��Fk֠�nrp/��34s0)��p��e��ŢF�

�C���Tġ�6
�n�y��<�`σ&Y���53v<e��}�X��
��Єށ�6��b�!W�Os*�.y��S1T�Ϝ�)G*�]����� �A��@��qzJ7���>��W�J!�-��{���\3L�$nEygP�1(gKWD���B����z���և̶JO��/�O|n���������Bݪ؂�h1!����A��'�P�Rlܛ�g+(I�9�j���h�^,F�ޥ%�P�6 �����f	�?\	;h�!��Ϳd
���~�x�'И�~c�_˼�k�?p����$t����$@��a��.H�-v�
�{:1W�%֨��@ѡ����[�*��o�Z������"عc3��N[��T����>XF����/�i���t'��O�R���XJ���ӳ&��T3�	�J�%��j�жQt��/<,İD�dK�;;P������m����'B4��3����Vk�����ѐ��n�Y���uT>���%x��
�x��[גR�?�e�V5����k���@Z�~c�ֻ6=m��c����~-/�^��	�I��J\'?0/A�~ϰJ��>F2�|�I%o��}ʓ˿>��ٕ ���#ݔ ������>�y�.T$��\��ѭ�:S��$#�m�{"��L >���F����<�5��-'p�z��u�;|G��R�
�sQd�^б*����
c�8
qc�8�����6���	w}N����)$�dn*��a��qL�!{��
(�ؑ^L��\�	<�Q���_p���$��q��|�ߑ,���p��S^Y�c-����2�XM�Imc�xז0�U��ۡ�{|��(�KÇ�žl�WF�ێ
^�Ȕ,���w��zB��2�
������s��d���3nK����Nў`B����g�9�z@�g�'ޒ;i�~(?#�3����jK$F�9�GO�?H��˚%�M��mW��U���g�I�H`1�v�$��"2�ኑO5��e`�U��F�&�`�����v�٢��|�	�9M߶B���]��ٯ]��d����SP�y�l���'|����x�6q5Y(���09�&s�%.W�z�4O�1Xnt�KG�2w5!­���h�dv��
)��}͕�>E(�-�E��=�U`9��I��E	T�-��F��C�x4�Y���]n��+h_Mð�)����Z�R��TmA<�
$�_b��D��?V�|�
i�y-��Y	]\��a!��N�>�C�&�������q������̶И	��.�WT�B��g,0�րZfߍ���Ɏ3�L{�⡴��'͆/���(���4�(�����<ᴶ}d�[����0/6�>����\j�zci-#�5��{�����ʶkI8m��~!���/&<�=�	�����%�o��bNV,�6ϔ�ѿZ�H?�c� q���EƮ�C$c�����<��#M�ƹ!��_c4-�}P���bߪ�Р��U���(.��;\St�g++��~D4������{�eL5єy��8������ԣ����5A�/Y᩻c�1�s���[]x7z���,cƫ��,�E��'�'�Ɲs.�r݉÷���ĄX��