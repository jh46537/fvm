��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}����M kC�}0��E��t�r^����9�=�����r��q[����QHz\~6H��˛�y}ԙ|C5/�Az��X�\:X���)np������{X.���I�G\KV}���G~��v�h3Y�?�/���ٗ_�x����찍<�z}|$|��a������0 8�D�����u窤>z
\�٢Bi�I��/&� �2��q�Rz&���?昴�҄�zG�E��d]���وwSz��fXu��a�c�U�;�>\�k�t4+�z/Y�dl\�O��
��\�b��d�\k�2�������IP��{��E�|^�Wuֶ*��VNZ���h�U�r�wՙ"������iB���,铟m�!�:���s?a���gdl�ՠ�B?v�s���w1���(�@���-����ۋX=B�N�hp�iC����č��D�����۽wߓ�N�Le"��j @	\���(,Nڄ�R�N���6Ҋt���޶�Έ�UG�<O���K�4�����u��nB.,�<��9R����f-�K!�kn���QL�9y�Y����~�&�����`���w����И:Q��Q�hoG):�ix��׌�Om���Z��0�����}�*�G��gs�K[r��0���k�-�4�to�g��\��X+�˂�/H�����,���6�dS���\>�!6$�b8eRo�Yɹ�5Q1ߍǩNswF���P��Z~Hu](r*
F�
iOȂQ�����\�-��_v��,�e�E�r���C�a�Inf	�U�x7��Z�a�|�����15+�e�Xd���'4����m{(��RU�F�p%l�RXY��+`n�@M�O�������`��h������S�9�I7����^>��KM����������,�':S<�=�	��p���~���aN�`(cbW0V�K��'5�)�|�~�?z����:uC ���Z'l@�2��[���+�Ǉ�i��}��g0�M��n>XU�z7>�+��z7)���f�� ICf�K�r��I���z��C�	%1Qi(��ۧe��$x*�t��ªzZҘ��:�ذ�(�B���ˠՂRNc8�sZU�^w/'�\��)=�z�����0Y���k����D9�h�hi���X�����s����Fi���s�<꽤�+Q{�wB�	�����N���!���7�8�^c8�Y0T��,t�f����+��& �/���L
I�.��FS+hu͠���ף�$nV��D)d+���C#e<���`"h�~�ex i	�7��kMĴ��؃)��R�#����㸣�ZRwed� �z!���acV�	�����w`�s�^���� i����苼�����Wa�S�8��Y���'����u_(��ls.�@=���?�xUZ����vp��~1�?��J\�u��0+N.e��b��>�u:���Pj()_"���0��.��l=N1|92]n��Q9�&�o��J�e�,r�Ǳx�M]��CT�j!ڀRG$"v�7���4�{'�#G�H��̓�ʄ����F?��0�'/�v��X4�R�K)���o�B��`�Ga�O:�q��Y�Jp�M�����
k�JK�Py��~��04���v�F�N+dl�2���X�T���ך�2t�݂�g�� �硔]��3���]Yٹ�h����>��|��$��"��Ǟ��P��pl#�� ]bFY��
�;��(A���A�j8�����U�h�<������^2�D[/��0ɩ��bꁊ)�uj �&�ű�0
Y�3a�-&`��nH8D���*��t�1�a��������n��?rs	��c��VZe�r�.p�
�o�	5��7�P�_�J�Q6��w�32i�~���>qqZ��d���+�D�<(<�MS�K�T�)��|�M7U���L��Y���lʗd�Cs��kwڌ�K��Ct󉙙Z^�4�֞��a���j���.�iOҤ��QLKw�����kZh���i�p�M�q��R���YԷƋ���O�1�{{����A�(����p��5E��U0�^h�C�g���1R�����N�'㌾d��bfhX�F�WY���<� a����.��W��f�s~F����V+.��-�>�C���K�v�O��k��Y��L�ڦr��Nh����.(l�6k�K)�f�nY���[�z�����!\l�;�˦B$���>�7i*ĸ���=��>e���^M��LPD�[���&\ݼ����S跛�%��UK��,�aQ0�PV���P��<��,ѷpL�Eh�`�̳hl��B,��Z,��(-� ���nfo�MX!�D.��U�A��tX�X�~5�3�������^I7{�L �א�1�k��K,Z�S#G�O9F������21��Ŏ?Xz>
RQ�����tRĭAw����K���Z�;ЍZ���|�7"� �ˏ	u���j�U���>8m?��|��{��W�<�
* �ș
*y더v�fN�:ޖQ���0�i�m�*������by@�p\e��T6F!U��Dn���?+��>�Vp-+�7���K;������S^����{�'�� $r�6T*y�8���$К���tY�B�Tv�(j٫�![�P�z �:�b��6��:�Fr&ԭ�����5�UkA�����fK�LQ]��������,�<���!k�f��(Qӥ��7��������B/,��6BY��O���'V��F�b=���$kd���9 9�3#}�L��漚V�6"���+;��T�o�q⚙cDMU�M���M�r
�AC."6Q:\�����f�ν�������ܘ��w����!���&��Z�/Ż]�tAqc�?����*�;eSN[+@�)q�%��,i����fꘔ���C��#�_	�S�����JUml_��ʱ�䥃��3�K8��rʩ�(3ݙ��Ma�3�j��f|�H��e�J��j�I�bѫ-������-^BS���6A�H�_�?�r7�?\��%f?<&!@A�k]�H�W��ʹS��J�W�,�HdN��$�&A%�ƽ�>ܼ0EO~Ȝ�7�e��>U�rL��k~�����㿣���DjcP�i�/z������$4�mL��J_��{�s|]��T2�lDS��W'�f��0(ߏ����T�M�m�En@���gу�ao�4$3ӿ�A�SoMw
�h{��?��Ɋ�->�2���x�d̽/_���T�}P�1����R!�{Ey���9�C�^�0���:�U��2�\"�&����H{͉	��	p�`�jO��h��؟�r��!��<n�@dT���ƀ�I�O�a4�$6>0���x~@.M���n�R^���%��:�؟��Xї�)��o}o�dtZ�x�ᄫ��X
�,i-V��rζ��Әx�Q6�@t�6nr47�؈ʙy�� �9�8{6���|�}S�?�ݏN���޵�ְ0C��h�wjǣ5N���o�����k {v�y���P�Z���v���sO�D���\��4@�qPO}e�"J��Z{Ɵ{�,��z��4��JT�7�h�c�ڞ,��P�E�89]B9���tծx_�\���M�o�]�2����XFk�͖�>Z,��FO�*�"��B[��<�G�R�a{ʙ����OѺT.�<�F#���(8hh�����r,��X�"o�zб��Ҵ�d6`�CT�zj��Մb�<�1s��?��QX�u:���9��]�n�j�nz��'M��k�����Ӥ����6p�#����=��v^S�=�R��9�o�����;%��-0$�ߖT+L�����GN�Dʡ�-�,�/@OA���jj�_�hQ�!�-e��l�܁hBŉ�5���W)���໡�u��$d�-�<�-:�:M����b�aDO��.-(0 b�h>�]��lU���*�GN���(�~a��-��ǔ����=��F5�Q�O�!6e�y�������L�l?1HP=�1�p�{�V_�߯D�1��ϵ�7e�s�?���+�@����)R���5�kB�*����<�>,��S����s�p%/���׽�g6�7a�گA�E���͍�Ju�Ӗm�Jd�dP�9c"���Z�l�n)��.,<�{\<=Qp�����E�c�/F�.L旄�;(���~DQ bA���gDJİ_'�)��x�jdt�b�*�Pf���""�nW���	��@:;2��!ĨvV�4>!|�A	fߺ-a�9��2jr��I��g��o?�����Kۅ�>9�*-y � <��u�@���|k�Y�᪹LJޟ%�u�
\t,а�q��fb���$ԗZP��&��9��FŘ��]�0_�^�������Շ���R���[�+^�%�* ��<n;��:��X��T�qb'+�a�����+_@@d� �a*w{T�sN �HH7�O ���9�~`Ln-
��K]�"��oEK��t@F�%���q�@�B��������
eI<օ�[�Q!&vIU�N��->�� �uUOŽ�����4+Me���R��]-�܉k��w��mk���A�t�o�|x䬀P#�,K��Yߵ�?��5g���2L�0kN���@ZJǡ�Jz
2�]��������[s!f)�����q�X�ܮ+��խu��ES�`R��/��zB�������u6�5PK�JȤ3�wɪ�Ԧ3�;Ma-�7i��%ҩ�Dbd�K�:�H��UK�g�~�Uˉ�rN�"{�" �j�<Wr?]�WH�Q;|��	ו��T@S��g��tB%�Uʶz��ĸ1�<�Q��do���:�p��'�W�? 	���[���3�P�M�p�{H��
E(͌TTɐ7�?^�_��s��U��.
8R�V^1϶)=� "�.���iS���V˽:�'�m����ݏu���MfuOO!��o��<�	�]��.����`%ߞ������:��m{v}-I�YA�'LfM=��".'�/l�tɼ�t����~T՟��N`p뚸�a��A�a�Q�*j7n}�k���X��V�Vm�37:����x^�6�#3�E�r��1����x���u�J�vy"���ڄ�5���}#s^�����Ps\ �Y����E���]��"ކM�r�ME�`q��ux�D�� �w�������$7u]�� �a���D7l�l�w4��v�ߙ�*Rc��Q�wz`��Q�ѲM����,f*��f�QԊ�) ���Z�3q*3&<���Ȃ�V#��WP'TQ����t�+�X�!\��SWY�S�VRA��_ȏ��.�\���Rri6�]Gk�����l�`�%sHR�(�$)�~ OdU�m��!O��>k���l���٦���?]>E�h":Z5}�|<����zh�a�1�9�(<$G�&ܜw�жTJ_�*k��m��S	��d��9>��:��,m��t���@�ҁ��[�B?�{�l;+Xg���F9��¾����3F}@S�0�^�N��+���m��Жj�+���e���S@�S�|����9*0J߱9F�LЇ�wpcT`����辪^�~_B��GFp�t����eYl.��6:KmW~�_��i����(+&є-�*qW
� �tI��{ ϖM���{�WO���m��S�����!m�~��Ұ�^eh��<ʋ�fI� m���e��79�;���9}�3��ʊ��;g�].K����������}\��;�P�������%����і��z�ή-�|ң����[~���!-Ln�97��Ԏ֫lP�Z��&��Vo%��{����S`S:e��oE6�g�=����;R��D������oϼ��G���?�/�#��+�K�
�u�aDÙm<i�q/?��/`��vWߩ�#d��=�e��j�/,c����^>��?ϣ(�`�đʴ����zᮛ��׌��TX�fgj-4BI��?��t2���`���E�2�^���i�W��*U:;�J�����<���䲐:T�b��7��1�F����fM?6�s}�Vn؝�L�F�X6c�E��'ţ�[i� ��/������3� $��*Py���%���u�WU�
6��:�:J��b�����4S^:UU\�ٯ����`<����i�� �w�L{��/ZƏ�[0:���㠚I0I�#Y���|����*�����O���T"M�$����OI5�����+e.�0��!���j�>b����8p'l[T&C��aw%���26�w�m"`�h� �_��Pt�Ҁ�t���#7�����Efj��UsS�l���F6�6�X�#&+T6�� G:l����r��B���`���������H�>�1b�ƖS��g��Ɣ��r�䢜��u$K�0�V��Lȥ5Ep���*��XgA��}T/�;��̒2Z��"���,��p�NoPe ��J0�a(+��>���KC��xwgj�1j	V����o���]�BbO�
�y�.�߂NΩ�e�+��s����TC�{�����76�pZ>m�<���@1e=�r�M�VO	#m���fC�:����&������5�t/��0�@�M{��,j`F �����~։)-�����G$��		?���'b�Zme����_�ž��.5/Ϫ��$̊+P)��Υ�|{Q>����PI���Ar��v�tA.�	��;^�s��p�)h�-A�]6��qq\�v?>C�l�G[����޳ �g]oE�o�@*����c�^�4 �pF\�ͅ�|�y3��=-(�OX�&�}B<
)�"s�-I�GT�������#W�)_#���.3C�Ɓ@m{ᕂ�\���P�������Ց���`t���i!h$�'S�}��n���p7��^���?���R�l����x~�g:����;Y����7�f����y��*��pҐ���L3]�/�O5h��P��Bψy5�?Dh�;F��SLr�+����*uPh��OG!�V\�x����ۼ�o��a��	j��\����r��f�E��8���b����z��&a:0(�\�9U�>���g�6/����L��5f5Vv�G�M2�����A��
��4� �ĵ�t�X���F���U�XJ��B�-�l'���U���06*i��9�G�R���zߢ��c4�;g�?�@�P%��ڞxф$�y"����
T=��WcM\eo���J�{�I�l��F��? �:93�)œ��n.�Wj�dP )�/�d�fs��G	� 籯	�Ddz7i�#�:qt]�od�,9s��={G�MI��S�ۑ���'�b6�A�gY���OqlI�O��3�<�#�ң�p9���Y��I���a�L�=��h���#cxz�t���n��c��#ҖA�H���߰q�[!T��ߐ8T�m������oL��u�șW�Ce�r&̉#�pd[��E��q�23_לH�k!�#[��,I��m8��:0��L���� w��u=��'�ѯ����o�4�^T��z��ʲ����B1�L������JZ���/5��'���[�i�Hy�d-pc;р���6��:� ��m}��S޵�l�t�^IV��o�.���G����1�i�>�"�����c�%�G(�T�������-���o�Q$i"�:��*h��|�ܫF�@�����*q��HV���Xٖ�^0TS�a��7��$��FAN��o�s)/��a���_�w�ɲ�+\��/�n�&�⯂�2��t|m.�fE��L9�1��Af�~�"��;/�Q'8�4?�ZW��^W=�c`Id��n[��/p�� �<�^�������8ڑY��J�sr;I��te[�O5�+�OS�'��Vuv_![N�A����L���I����=��b������Y;��ҫ ��x��[m�8�V�|�E���:k#�Y��J���n�>	��X��ϳ]�Z��*��ȸ�D����1�q������n��3	��DJZ�0��r����^�"{���QhU���e�?��_���#<`��(I�S̲��"��)c�ۜ�q�́Am���߉W��YFxԔ9h=��,{�y�-�i.�#�ݭX��u�M��=$����w}i�\M4�PXD����_F�e�r�����{H��h�~�q���wIf3��)�.FU����������X�yj�y|i��:��r���U"��;j;kU���0�I�´w~�.>���iM#z�..g��q�Jsjmlh���6h #�3[�V�ʥsY!k`�;X !�)�e+�Z��[��F��.׫�)C@
�5,�?�y���?�pE
��/���X��%��Z�L)��|���'T�#��d�h�Y�<Bw:9��(6��2b�i�8�Њ{[B��ɸ'�Li(�P��������2u��1�v0JDo��)�s��y�i�Y���ܽ"���������y@j�?N����_[�� 'SMkB�~d���V�e����$��W&����ғ̟��t6@� u��]M��1W�3��RF�TR�:0
����Bχ\A�U6W��9ƌb+/;wr
��mWE��A�8OqL�H�~Ѡ8X�J_��7�3s^��!zN�z��,3�dx��2���y4���V��&С��:��6Bc"�SA��W�U�%�����1����]k9�Τ��I��#'�o�&cQ�@'��C&c��}��2W�xhL$��e���&�F��Pȍ�� �2�:����;ln�����u��;}-4@�C��A���O~nf�v[`�_��)�iT����]o��/�ͦn��6�q��&;��*ݦ��w��(Sظ �D=�]B�R�n%?c惯���)����d�>��4���e��v������B�uO��0lq&=P�FbRMA�$̩�BR�������~9jw���#�dU�����m?�����ImKGL	`�]	�� ���eHA`�d�Rpy=ՍT��[�e7q���/�������U�p��i�%�>���*����[��G�n!�8��Tu�aP��t�Y�g�W�K;��͇5��ݵ��/褫�EIR��7��`�x�R��X	��A/����Q������f��!?AMfǝpx����MD)�����@EDQ���F5p���A��l�\
Җ�\A�OwܺÝx������ s�]��Ka�U~g|��,�v8�6��E ��]o���'�.����:�B�n�����ƻ;�(�l����p���˕�#�z �I�3c�A��u<%_��z�t�@��{Oى���x������K�W�j��z�o�=��C��Ֆ%H�����I+W�:���ٝ�����0hԛ�.���;��_#m�h~��oZ�a�]��.�%�l���q٥ �'����:�>#�����O�A*GhN7�h/S&#�r\\�	)������n����%xef��̛&�HLDH�� ��C��z��v@�B���;J��(e���Ld�'<���krb�>|{0����}r2���ƭ�A�Z~��k����@����-�L� �E:��r�������ܴ�~�"C�5����KC[@��J�ݮp�T����V
M��8������ȉ;�[�ތ���<>?������e��Y&�C��[��ս�L���s��K�{��&]�㉎X�Vy���(���`�����ߩ�fB���A���x尯������������~�%�����?`����=�W{@���7�f�G�2P����½�G�ᏅA�Fz=��^}�-.ߌ�����L��'����N-�ї(�FL𨢴Q��GA�-Y��9���!���P�Օ�1r{/P�k��eKS��G�����*�8�����Y�!��dK�a�;nq#,��~���iY���jD:2N����ya&�����¹��"��Bq�­��%��e�������SkK�R���M�>فo�[|��V~+G��L��=[?fbn�\��Rsތ#���
ؑ<ȣ���64t����3��{CX�+ɩ�=^A�p�j�zdj���k��ɝ� ��ȹUd��{p"*I����ռdޣЖ��O��ޟ;g��"���mz\M���"ʼ]Qj�6, ��u���cP?}�Q�]4�����D�\dwH��ݓ`YR��'��>Ω��,��J�k��4��m]<�1X4foݧ�d�l�Z���鬆^�*��!��
�U�,)�	<??gt�bb�I<�,q��3�b�&^0+�2�nS\~^�qJ��X'�ihg�$����%�i�p|�h9���� ��2�i_ԗ�)u�z׆�f�P4,}l��0�吗���yuBy�`����ls���(��U�	jļ�-����g��j�P�9A������l����&$�_�5�G�i��!����G��I�����$�F��b�q"�Ԕ�DъѪt��8��|E>��W�?�W���m�y��q~���ڛn>�&��՚|I�Haw����^���4KaC�v�������Ҙ6;3�� ��MA���^T���p�3ߧ�sP����Pme�QQg�t�PH](��y��+,����O��=z��h�91>�:�u��쀈Ց�f}i�����Ѵ��&m*oqXZzxW��`B۽W���睱*�����O���w{K��3���}�3XL�"�`P�p���gC��)L��8�ͦS�"���]�u�OX�)���e
~ 58��Q���l#b;�I%d�*$ o�1'�[�����}����Z���W���`ރpĜ�_[T�h�`�IV]+w��fl��� =��ӛ��-�}6��ҙ�-͹u׀�m���*�2��R���ٟ�C�"M�ݴɦs,l��b}a����1c�W���7��hX3�GA������!�e7�����ې���HȿD@$
��U�r���-���G��X�/Q��0O�%��Ѱ�Ge��n�&2��C�d���H�#���q��N��1uZFc�5�����ِ��
_c0\e���� ���aH�$p��wk�i���}�L{w
�{�)֮`�2�T���J~\t/PWɑ4�IN�gQ�jnp���!.��A|!W뢿�l*�^*-PQ׿y@$�e���G6,����흶U\�LP�'���6�8]�q��9��7�D������*&�اe!n��x����p9ۼ�+&�_>�`���Y��1$�����
���ֶ#��,3ܸ���*��S3�h�|�����  �'^�݉���k���~E^D>�13�M���]��3����uZ�\׸fka�8W��X�`�rZd�SXP��>�ǜ6�e�U
ZZ��ٺʬ��*���A�}I�]�L�Qz��\���-�<l�P'�1Bq+KO/��xd�s�ӈ�|z= =�Q�`�?ufk���1�Q�G���\i!��H����Qۂ�!,�h����o�z|��B׫^�3�ة���ǣ�u��;�G���Z}��?����n�#}�����]�q}�ed����ɔF��0���&�`D-j��}��"wb�$N�_�2�𯝢q���:��e� �G0HF�ӎ�98규Zf�,����[�9��1FmŸⅱ�Ml���-2e�}G���1Ah��*������j�}k�iV�g��$�����4y�>�]1<��̐�}r���p�g��Q?���h��>��i�S��CNT���V��bYi���`�����?��ƽ����0`ާlϦ��.@��&3�UG�\�jnp���H��L�`h��MUI�8�M���\�N-U��j��;��D�K�D��r�65ʎ4*���_2��\�f��Uck�)3=��#���n�8�u�1��/�7�������J�KB���^� ��*���.̑�t������T�a�$ES;������*�bj���?d�GB��o́*9�?X������r07�����Ɖ����Fm�l�S�̤">@⣛y$\�>Ȁ�&�?M�/�c�_i�	��:GP��s1)r6vO��-r��R];k~�e��z c�
S��R�\~O�2(�Y���[��Y�4����7^�(�[��M&9q�!��<��G�F�����{���
�T�N���xn��'by�7��,�T�µ���m��&2�D�æ�t���GPz���K+ʶ���f�Hv�M��.�t�ה������j��7���@��R5�#r�u�K*��T&��/*A������I�C��@cb!�"�Fq����%�@I�gƗ8��Vr��^�^��D�̏��ߥb���OL#W ��B�;]��뱳������6������(��*�K`��"W�.��F� ���'�����^d#�A*>sߡ/����yܽ_HVq����,s�5�W���4��:���\D�L
��؉3(�w�+ ���YLR0k�����)�d��,�z�+�۠Ղ���)Ϫ�6t��Ë&���1��V�Ï�d�K��J:3�8+��|^ݜX]�N.ݡ��a7��I�'��ddr�?�'���ɝ���ˑ�K{��Уt��!7Ⲍ�T�k���u����X�A�'+�	��<��J g�2�R!���jȶl�|SUp�+���Vz^��1oo(�5�fRd=Ә����4c�(0�f��<W�h�l��_� ��0N��Q��%�L��J�i�2+)%��l���.�SW��H��R���G���$+��!��)� ��ν���y����IΛƲ)��a��t������5�2���{�W/wv��r��_��0�.��bYh&��|�v���@y���l�?��p���^>�ĳ�u�}�a�b)+�P���EGE��\���o�ึy�|�W.$��)p�aA����%T�Y�M^N0]�b�6F��[=�Ꮘb�+.)���yN>.���j��a����ebF�op�nV��J�2�����P��Dk��Q�%T�l�k>����"Ї�'M����%'Q�Z�bp }��i aFN
���O��8Kf~���p��t3oD�Y�C;�$�0�}Nĭ�����#�"��54"��*j�=8�������*7nɧ���#�&��'�Q�^s`=��N�L-N�����
e����y_�)��J�.F�㻭�2�e��b�y�nO2�F��^���d�'��%�.�1����R��T)�$?����e(U��$7��M������50����?�B�\h
�F}���ꏓB�G�2.=��贅���݋�Y&s�YE)�N�!>d��T;��(\�d��~�2��́Q�}����à�����\yu+]40ګ;c�7<�����J�������9��4�MKϮ<�X�9}]?���{�v���L�]���R�����F��]�,6S�&��0��;���ʉ�&=�%�&g&���<�bY���΍�,�ܗϴA�gN��	�ܪ��r��У�'�rl2Ĵ6��@ӬyES��i��W2��No}�n @�.�>�I{��5��ȿ��t���(�K��|�lH�cF����R�WM�>XVx�����"�'�t�����괓ѐ�P���q'�mÐ�~203�W>���<~��`�G[�d���nH��YF.�{v?R�/���� �y����C����-^�,�\C5�q��޶�N
��tޑI�G\�ʢ�6h������0r�{����|O0��'I5�Pb��e��'R?BV�Cci_�up���l`����#���^��i�n{{�Ϯ������F����l�ÚbL軮>�u��C"fG�1$�x��}jV<�\o�|��x3ƫ��ڠ�D���$��/	ѻ ��:�B	�bI>�щFKt���`�[mߖ�թY���n�Dh)
��ă���#���WC'���tL���z+~"�9�t�h�m�Z�(��!�cg�s}�:�8a���i�@�m�o��������3��?�XB�@���ϙ�@���U]*t�}e�/����U���D6�}�E�q���8�I.��nL��!Y.���4�Oԃ0�� v������t�W(a����k��~u�cFw�� ���LT�sqC�K��.�N0��xej�Kb�l(���~�#���Z�#��y�Q �V��qw������W�sp*1������x��4�v%��%�MCW�S��@"�:޲_ɥ�C�D{����8t�/��I�] {.���{���pd�v���(�GX�H[
]6�@6�zx���%�m��Þ�&KZ�u�@/,����ݺ���j|E��i��q�ҜB���5���Ҋ� *f޷T�5��ƻ鿬���\���:LO�x��߂9U�5�}_{�r���
�{3��X�˘�о�£���
p@%~�4KhY�r��y�j�U䧏çN�ɻH/��l�Rؔ��p�ۼ�
���]b�k��m#���O�LoG��
�Et�s�.��y��*��yU�\�{��^&�_�e��|Z��rJdQ Q��9�Z�G��Ò+5T ��!W�^��?� �f��E6+3p�b�GN+Q^М�i��������y i�H�.�v��iThCZ��K�S&-9�B ta_� tN�b<>-�˓t����l M��>���FT�"~js�$�{݋��f��/���%<1�vvˏ�T�}�'�;�SZ%S�=M�|�[���0�l���c�Er�RpA,�����X�	܄�-=md=�������q��5ȳ��-��4�~�eΨ���B]���1���֒+�=��T��2	y�+RXWN7�WS+l����w����IL�|_�[�I�j��l�Y(Eڂ�RF�^�A���|��i�؂;YS1B���r�Ț�%^��^O�����lxv��L)���w4�Ͽ*����ħji��U����]dO�9�VB���(����O'���+�j2�|���=z�Mɬ������Vt�����m8�*�P��J %>N�O�i�M�IN;���8��V�ZIR׸�h����C&���u��H�߾&V�¿�|[�<�I;����_��y���uG)R���I(��#}�����H�4�-3���#���vFP��(�������X�
L�Ǉ���qm��T��D�3��Q.���m
9vep�=���K��Ap҈��UE�\��Ć(�hQ=��2����s��{ǎ�A���ݥ�b���GD@o�.���O�1���h#�[N�!0���_�B�7F��~�-�N��w���8�%�t/d#���Luk�����?Du1���b�S�hG��w�.z�LX3w���V������&�Ӣʳ@=!��&�u�ZE���h&��[S�@�`H$A��K���+�9SZ�_JJ���x��3�"NpmzD�aN��{����G�ON9O��F{�("�
���w�\��d�M�밐��Ơ��HEe߯bE��ҳ�Aɟ�c�����P�Y�S��\�y!�������H�9dr���o��$Z�K2b;��o�����"��v��p���ioRx	��������P�����i�qB�����k���R �q���z����e�cR��L��T�>bD�^�<����ڽ��u$�j�9%���i���$��7���<�:1H��~�a:�K��`�+_�L�Q�P�m6�݈�����}&��ܫ>��^ybF����R1�Z�ܗmY�j��~����<iP�J`�D�~���A�m�m�O�+��?�������%���3��7�S�!���̲آ��QԷ#V�������p_E��7azl��;mI�)��	4O��g�����!9V�sؕr��d7݂��>� ��<33���٣�OV`N���)Z0�WaQ��g�k��Y��~�G�|�[��xV�ıwp�`�Ϭ���uRU��R2Â�{�eI�c�2nxJix!`��]�W`���9,�Ĺ	����`E�	5C�^J��E��2W���~l%e�M�#�^�R���iR�B�R�D�I�zO��8��SF
@؈YvP�0@S�`���c\܂M��3?,������2g	0ʢ1��7����� �D��:I��gA�՚�I���u�84��=�//7�Q��ޫ5I7��%���	�fo:�{W��ܟ�D��)���	 ���8�������
�i�����\�X3��C!yyh�5L�ʬAP�Q
�#��`�sQ�2Ҹ���F�~/ĤB�HH��6M��|����t6>�F���
�	PH�I��p��])彛�)�8(��py�`͌A��&���)R�73�67{(��t�'��S�ٸ��<o����J����Bɤ����d%�N�{lm�̓���7j|�i��P3H�a��
��1B�cc��1�E�c��E]H�g.F��Y�Y������n^��z�d�a�N�Iy�I4<vy����3�<[��وB�߃qf�>(�d(�h�X�ww�
�>VZ��pÐK�|�>BwU��_L�\���6
�d�c�O"���6a4����
޿c	u��z�֡6�,�B��.�3�~Cɗ����[�,�t�⡅]��x[�l1oR�����K�8)vl�{��+���N�fT62�=#{B_kW��&�HV>T0��UO�Ԅ �������L2s���lK���+�D#=�|��Y�`Zz�˩�/�ܕ���UoeW�f������8�Jq3#��E��3>>BF^�����y`oj�	
����E�I��I����lƖ�GP,w�j�@��|�Ԕ5}蝊���wq=U^ĳXŚ�"`�b�l#�M����x�kes���T<�Pzh������.{��R4�x���n7�1��K4�l��{�t����U���M���Y��x+��@g��Y�6��}o����I���G �^ؙ�K�
�&�|Bq$���ݺBz_3J�ܚ)WN�<Do�%����<�U�����J�q�癰�T�.�Q���Y��]�Ɵ)[�%��g����� `{�2<��5i
�zI���(�İ$�USď���$���Sa2������hKW@���M���k�^�'��DxCE��wp������	˩�h�)��ȷ��kL����κ!�۰�ݽ^�������X�gx�6h�A���u�-c�����,ԠBm:'�,RMO���B����OPSZ���`b�����\lOg~�Pw)Ȼ�C��#E��Z���@��v��T>�P컙��̾��b��=�m�4��F��-���J�c͟'X�8Ÿ_'-Q�w}P�V]g	�]�G��Ћd�^�n����J}�����X��Q��7�ӰT��G��_$�h��Ұ"����4e�Zp ��p��X8��;s6v��/r(��z���^M߳��u?���8w���}�%����r�L���K%00��%��@cb>�@�DTI@��T���ci��b0�S^�=��ꖍ�s��ӛ���)���xd���g4f`�/?������e:]�#�$)�<��ߔn�>�B���e&��%���UW�B@�����)��hʬɒ�znB���8�*�ZH�J�?*��*�m�/��{J#����1���Vm"uw��wcr�7Lh|<0"[�^m�~fT�B#gp�C��-h�����:�������Vߵq:�M��0�6F����7#���p�EOH��i�!�i�*�׍T��.�d�Wq�O왚��G�;
��H���i������߇�(f���7?ҵ���eV����/�C���J���9��
�tw$�GU�3R���`�@�8��oY���nXT1���l���~�	q�J:�X��������?�p倓�i�d%R"JN&šǖ�)���Q�`(���H�Aν�K��I��B������E6��$F����1c��{5ɑ�.l:?-<ލ�"'��i���ǻ��F�� ,��œΝ6W�/�q8�������+�얣���*s��c ���������p�-�ԁ��t�L┰����ֻ�#/��u�l��:#1A����0v���@��rP����Q���yO��V�imA����U��u�8EiM �!|�L���B�P����L+;���Yl�\C��R�p�F�7O�2	����2^�d"��͜����n�
e5� fG% +�F񖸕�J���7�Y��<\�몊t1��u���^��̬�������"�A_Z�Z��ٹDPz�
,���R�Y�������.�*瞫��P�����4�Tc$5�1?��ʸ|����X��ͱ�;<�:�z?<��p��܍g���+�"�ո�Ux�wn� ��5�+��#_ s�l�ޘj����ې�pͣ�s<����P��P�wh�6k�{&d'��N��(�^D��-��j�{~�+mVq�Kf�[)W�E����S����зr��z��>����5�k�n�h�5"3K�.�M��R�
�f�މ���'�.��Q>T��~�*Nk��x�~ (-�r�c��.ml��_���b�篪����8I�_�w1����Z���8Z%Z�NK�O��*��&������O���ʑ�Ā��ln��Ă�y��锓L�˾�Y<9�7�g��N�BJ��g��N�|B.�cn&��L��fہz��#�r��搽n��b�)��ur����=�)��X\� ����ф}׾n۰株�V�b@�x�1�t��}尛���T(|��F�x�Y�F8m�{�
FÈj��	�����z���#�@�0N���0��L��P�(eo��͋��~���g�n+��U���rTl�ccF��� �A����)+i��#�'�qԛ؃��|����ipq�)l%�8FֺE &.eF�(6/n�%pD�/B�ݺiW���R��s<X7]WW��F���5c��PPT\*͕+��� wţ�W�z?3�Y��5���t��8@�JUȷ�(ݕ�-&�	�Wv�+�~E8���A?]��t�
�����e�߾�)�
z4��]W�@�RD�k$�$���4�=��
��I��t^�b�w�y�j�C���	n5�}zkg2e��Ϻzǹ����ۓ`Z�Vg��?}`��	ume��J��t����T`�<0���yѮ�(�7��^b�������}*b?7�!٢+���p�^`F�i��5!v"����.��7v�����`�pA,��o��b�	�OT ���	Eϓ�a��G�r��_�VW��"��Gs9@�G@V����6��*����p��v1��	���mdz�tO�~�poC�?�Ã�1|vJ��M�.sS�1C���ă���Q��}'�:���\HSV
�g��G#f�G��p��@����>��6r�����0�u�+�����a�Z~�}��:�H
�Nsѫ�N��DYL�;����#;GJ^p�S���v&@�%�u�:z�����6A�������Av���e�ϔ�������ݨ 
gt9\J����������������jHv���{^�`���Z ��&h*��iwd��Q�a�Ď�I� "�7�t>���4Q�x�­<ʣyr�`T�`�I8���<�*|SAԺ��(��q�^ß.�����Zd�����L����JݦcnQ�{T^��Z}�u�Æ��Y��/�xW: H�u/�j��1���4�*R��i�Ж�i��m!͓��!+h�V��
�^H�9��<�`2s��B%�*7�P�{���q�zQT��B[6�=]yb�)�^�o7��B0iۊ2]:&�(ty�&��	��!����*s����@��"�����4Yޫ!��8��k~��M(l�qwe�2�R>j'�cP�=A/�GlS�/֤
jQ	�юJ��FЍ���.4ɯ�:Sa�di�AVԼxs�DWVa��5]D	!�V�$��%ZN��9~"� I&�Eh�9�%����o�n'/�iGIc��M���{V��M�ഊ�-|vjc�P���~��q�*�E��^���/7�յ�r��A�؛y���W�z�	��I��.P�`W��7>��\m�s�A+飶[���1K��Q�VVr��J����ܣ)m:��pD7>�cgdl�|�ĨeZ����Ű\|e�<>�`p����E;*��VQ�*o�]w��2̼� kͯ��Ƭ
�������|�(NP�F�AT>�Tpf!��#�imL�Pu$}�{W�o�rd�U��x,m֡d��,E�5�<�J�P\�=�/��t�=����E�HavJ �A)�!wGQ3�LAE(XO_�X՟�j�[d��	��}�~�Sęl�qՔ����'vbE��#5��QRA�"Q*\��?ԙδӹp�4�Dr�ۻs�T��j�1j:]G�8��E�M ��/��'��6��*�Um�
�����R"V�������Ze���?�1�6�<�A����W������Q5�>xr�(�1����l�4Bu:�&�w_{u&^�^���*�`k<���yu�`�*y�����8���� i�~�q��2�4����|�ya��O�~d�,��~��p�a�p����e$��1���P�� J��4�p���f۪��2��eK�u7ix3�	��]��[)faT\[��C��B�2|sq�(1��7:yj���Iu}�y��i�g��XW1��8�KD�>X���D�-s�tr��y��C�A��d�;��ÄB��-�C�A�~M�Aw	g��|QIeHKH��J���{�+�=Yҥ���9y�+;�=��Q�WT\�4~Q��\�*Xu���rh�`R�o��$�O�8Q��i�SZ������V*��=O:��6�H��)��2V�q�Q X*�93)������f��PQ�o��K���C�><�N����V[*� \h;�&;�r(�5��3t^��`����
��{]"|�
�r��Q�$qf��B��3nʶ�� ~6 ����E�J���D�7�Y���c�Cv��y%y�.u��3�yC�C^�A�D.��j�j�s�|�����]>�p��]�o/뱉�:��i��xމÿxS�cه�~�N��"֚v���꯺&���6+PDbk߆��ӛ:�>,�w)������OȦ��O��T������T�+(s_'e��� E��A�8
�7U��}�&����Z�����n:zDx4$)�u�ت�BVm�p$̮��5���gUc��m�,����O�T���B�劘.
x�:��o�x� U����O{
7v�Y;�(�����N@;[L�k���8(�lo�	�n��5��x�]0,�^����90����3s~�W�ˏ�aCO��o�qO��|��JY<�b�R泦�`�֍׃�nyO��lJe�ȸP�3f�_�!�s0	�L�-0c&��[��CO��/U��^I&Nz���a����T�e�[��s*�煀�4cv�nƶ]r]��Ź�ϝ����!t��$-�e�zy���h@�6^ ]n���KRb�A_��Chr��#rW��$��&mѕa����P��q�B�Ks�(�(�L#�T˷^�i�f]�(��.w �4&�a	jq��լ5�1��y�{!?(�Q����@�b���S+���>�Y�ʷV̺p#���dt�@�MT@��0j�<����DR���O������3+�9KI,�B����rgB�mJH� 6��H�W$b���źa�x����-G�x�����)(��@�Fj{-7��(;�E����ת/�n"X�g "��,�,��N{}E��{�*=��?��})㿳X��:+�I��mo�X���N�"L�?ϴY#o�W�,'�@��Ql�R���7'���b�t�r*��e)�JK�K]&���Һ��<�񒣾����'�1�*7Y��1���H]�Q��Ju�JI��I��y�&��y ��P���ܡ'�t#���Xr�8u�\�rc�;Ё��ʚ������ i�;N�ǀ��W�ܬ�� �{?0�Q��x�g[硝j�­��j5�vGn!��AE�2)ZT��=)T8P�v�����	O��xn�������@�����_jm��[����ܿ�~���c���E�a�XE���p���v�4uKԣ�x>�찑�aۭC�;�O�ߵ$$�.9�+��K�%�wj��M'�B��>Z*ۙ$���٧�G�ݖ�щ���|r�@,�ຯf�pg:�y���Z붐x�28�Q�Pj��*iԝ�k�O�i�U���I��B:m��A�묓�}��[T��E�����{3P��q�0� - E�;' b.��zn3=T.�ŔXh:��XA�Iy�e�C��b�\xn��;l��@1�D4�+�8.�>�(�����P�����޴NvPE���c�
�en��C(������DsZ���Í�^Ϯ���6Nz���S�ў\a��.�HO��=�֬˗%�d$53�j冀� �Ι�P��xX,�cW2�JU'4�?��?�b@<c��._�N����%�[%��u��C.`��r�����|z�'w������_������G��`��U��ʥs%����<�dil�п���戀�P�ڗMz����Ф��xX���i����H���D�Z�rƯ:<�+�iI����!P�P�������2�Y9�cBD����I����)�͏»����>�e%�ֱLR|΅ %�q)
�]A9��8?u1+f���/]�Z|
&C��)�<w �#r�����Y��{�0+�r�%V����4ng8�o�lb�K���l����kd�+j���yi��<$Z�i'fL���#�$Blg�VAm6S2}��
X�dn����̸}'3�5�I�֢�W��E�����F>S� ����6�6ON���5:�e�%��B/��~����<�:RE��Q�K�V[F��׹Dp��@�u��Q��08���裐Ķs����N�t�J��^V�Mf�ch_�y��=6u��!F}!'�`{�'(8�<����PG{���>�=ߦ3��&bS�.�Rj�)��@<Ai�Z�O��x�ֱFQ�0_�ő~G���]�E.N\.Ց{L?V�P���^�w��@�q^f��kIzt΢�2&F����C��M�y%��H��*���=0�.��:����lKĄS��5���-����{9��`�^��;�R6�ё�+�M��}�X�QT��&� ������۞���'�b@���ֱ\��M\�SMf��'�:!T�LVһ9����4u�'����o��}��y�o4ɜbk�����l���ß��'��έ�q��MD�(���v�,ha��+y����ְ�i���+�Q���PEl�;�@g��{����쮚����=#޻����{�:��^�K(��s2�Cń�<f"M�8���}�p��R��V��: 6i%p7N�>�#�zֈS��_��l3��NL<Q��rA����6]g�{8^~��g��#���y�؅ʘ���H�v�u�]�ڟ|�a��ʅ��b���0J�'�h�Q��/�?1t���]������)�0�!�y�$�r^qU�;{/���g�
�CA÷U�v�h[PZc�"ibf*��ֆOЉ�����m�[݆��X�}x)o�����h9��n��4�ed��SM���w�ig�ا����;�6���[֜0�u��
r7p��R���8ئ>ԋ3�m΀�����b�K�����yէZ!��A�"+��L�q�}^3�e�����'/�'L��cJ��NU�����K5�X��/vw4�R���O�9Yk�	_����Q�VL�H>am���`#'��� Yn��
>~�a*fb TBK]�����_��=c�������<U���%]���4�ԋ^����O$���8�,~~�;�0���6��毥��S�6a���@R��ZUS�KT���c�4p�4�K�:AƗ�_`���0?L3��040�xos7<�@���s6׎��?Ёz�*�;���󂪩?�R�^������������E��s"`L�ArR��>�����x�ے|;(R�KHڮ9.���V>�F��oU	x�8?�zGVk�]׊�ŷj)4
ZM����Tnk��X�ޮ��=�e<n.���r�v���Kn��� 9����}Lt�(�H	�wu����H��ˣ����Ai���á�~���}�����@3���؈lU@�]zi��@[#�h��'�k9W�`<���s����k�Ȓ��=My
��΃g��1�ԧ��}��5u�S������cG`�dc�z�6lXas�Kz�Ȯ��z��<�G���n���B3jf��,v-�'�\.w�G��"d��s�"�.x����E��_��	��x;8ěs�R9:�]�e6':�!���~~�޺|�m
lTs���މ�T��]�/�ywI��N�W�������S7U*��%4(�DC#K���P	���5�]�E#s���C\�f(��6�ۄ=��:�D�L�\��"�:Z^e��Opۚ�bdY��������/ �=~]i�j|HZ�?k��|���b(�KVhaYxjo
�n��]T�$�T���f��oH.b[�-�p*(G����4F~B"(Dó����}TZAy�bvn&� ������i̹	���@	N��=oKF�NkA�(֖L}|8e��� ���e�=�\u���+7a;� ���������!uA���.Q����L&��q6U��A+8*w%�胭�p�J����Z���p�U2>��,ߔ���R�剐E�5���5���=��:�5��e��G��8�p�Ⲡ��W#2����p�@�9ۙ
*�����42-٠�)�w��Yt�<�
Mo��mI�n��l���(4��4;����f�V!-�;��-3�k�+���(aBe�3G���*$k'�E��;b9�灣H6D��O�/��<���m W�3-���lP�CO�X�e��WF*��쭥�����tɚ���G�L����q����	��qҔq��>�v�D�U2���̀E���
f����RUd����c���U��.7��k�ʚ�sSr���%s�.���̟��F@�%o$<5g%�8���LAU_%1x�ni�7NGN��#s��I!|ؖ�B5i�+a�}�$��{�n�#4�Ž)p<��y
&���q)ݐ~͵٣
{3���4kI!�upSpR`�Ĩz��`{,�_?�����k�ڒ�T��n��}�,���o:*�AXtb�"�K�X��3Úv��V9ƫIO{G�u.߭�F��?��Z O�������+6��u�b?$\p\�n�8���:І�������9x���
9��D�i"�:����^�O.
s�_{Q��o%/�U�\oiZȭr�N�മA�␽@�ZQKj��!�'a���>��7�#��n�_;����S׍(-���^ï����	zi����^������	�W�]wA~�k�P�" ޅuF�w��1̹d� Z���==[c�� �׀�l3��Ē���x���t�jf��VE��Ȉ���Y��\�Tzǫ�������%)��������Pd6�V�Fu-�oX'�j��ӝ��Y}S'�e�k$(�C����`^K@v:�o��������y%�c������Y�nO���xhiK�a�4���UFO�H���on !��y&�F��3�ӌ���8��i�/'���A�'���XǻA�A}�������~<(P!n�~ �UpT��i�����Da�����I�e����\e��1'_���/1���3�z��
�Atl�	��U��~��F�H�K&a�hLX�Ų��,Y�jR/�ۖ�=�V,��q�v,,���SmR�����L�4��������4�%6��e<i9���q��I��1�x���)�P�)LWMJL�R���_��in������<E���#,Pk]1�OA��e��1��6�i�M+�}��r�r����h�N-��^��3�"�������_A2�"_�4���������M��&����9�<"w�`Ǵ�_8M$Bxa�޹Y�~~ ��zR%y�l�	��H�gX�y� �D��QF���o�K#�3���p�qڝj�Z)֪-��D'�����kO���E��+Eq�����V,V��an��DXs�F9ۤ�C����xq��gs�vY̤���Ӛ�{�n��F��u���V���X���KM��f�x�w��K��E=��Ͻo��WE�T�Ի"�h���6K�@��;���\@��t�vR|�A�63�ߠ�X�?�ј/ax:�ν5��b�W��h���v'2[�]���������6�&��zM%�L͢7��_G�U��������,v:� �;�昷�l�Ky�<a�Lҭ���	l� Ψx� �"���%��!��d�3�ZEN"c3�3�yA���l���n�5����}�A�g���YX������L��O�
-|/47z|_Fa�:ծ����7ahوʟ��J�fN�&������gr	�W�XtS��#>���c��uw)��=�86����k��x��^ö�%��E���6�c�< |��;��ӑ��B�Y,l���ǲ�#4�����2p?TNR6��xZ��i=���Z���u�y�~nZ��ܺΐ�f��h�M2��A�H�1��1�v����A�.��XC��m-��g}�JY_�Ls{��&b�ysfFJ�̌|˿��i�8��-/���ٸ�8u��ʤ��ft�J�M�ʐ	�W��׉'7I��{�|s�� }�ӿ�!�S�&�5 ͅ���T�MZu�F�ƚ��Ŕ���7KG�<��j����}����yq��UHW�ь�2�;�ʅ>t�Pe�:א��j\Sy����\�yt!��(���6 Z4WA������wv\r-Z�"{̔`3�F��ru���31	����)����@q:�U`�Pd�Q��ݤ�&� �Sv Q�#e�T-ϝ蔋�-eA��"uo-\6yWA���PwQR!�fm���ˌ,���Ν�T���i��f�j�ry����Z\�;�׫�VϺ�5֯6����ie(�Pn��.(&�%/I@%M�$��4�|�BP�j�����D��顫���w�QND��w~�OM��{- �l��Nܰ�ڔ��E(����;�r/��_)�_����Q	���ʠ��(���t&jf���L��RRoP����}��n9�(� >)Ȉ���oV�_������G��/��X�$���7Q^8��Q,k�b��E�h��0-P�Gu�HM/֊HK=�����3���'a^'x�n�2�3йM�;�Eϊ��E�%�1�Ou�����5*r��v'�m���j ��/~O�S5*���Ci��Z�:l1ĬWhySw'�)��:m�,�e�hq�������RXm��V@O���8�L	;���b��tzp��V�p
����%��|��Y[x&g<��ԠG?�����d4�M��g*�f�V�	�M`�)w(P'����� ��� ��Y�Z��!�Y��X�`�C�^�g~te��?�˳UW��v��R��cX����-_�R����g_&�/T�"��ʝ����/����)K��Hq'��� G!]��,���zQ��m��A3!����
��#ɱ� ���vD�/�G���j�'�v	q]+��Sh��y�2U���N��d��������`H�V��k��n0�%t<Y
#�k|����5�D�����\����!+�r#����s��#�\҆���[�p��o�G˭q�㙳��Å�@������<X��Û懲��
�px;�F򍲉ck2�7�C�2V�G����)��;��������!߼�lzA�m�^�?"U;w�3e�R��A l��=�^s�7>ڮ��rWjUuL�:`�)]<kً��x�<sx�0�vh���5Lt�Ŵ������p���(�@�us��u�Gi�4'�E-*��3��%T���NsR��b}7K`�k����a'?�N'1��HՑ��UI�I*������|�������Q�s��T�ߴ[�[Q��k6�9�'M�ǯr�n�q�m�2�q"���eJ�NIcX1L������7e���oMTu���p�q��"��m̋(��I~��x�� �k���ҙ��J��<eW�����՘X��ld�.̺��jhK��P:�UC�\��?��C!I��0h}9NZr��hm��:�����,y7�QY
n����2�
����f���d�u���yS��ʀB`��k�.�t4�=(g�K#**�	&~\�sѴ0W� 9�'T�����~���1v�@ؾTg�k����$>J�k��p��]�R�g���G�f2w��BH�H1�5v��I�_ě������Pm���|���JL�	���/�ӂ��k�x?T�����s��ԛt<�,^�zm�+K�G���i�)9PD�vʱ6�(�c��2	�L1ow��x�(���j�	�����}J��*���]R����9Do��;[؉g)��=���,��wr��C��v>�b^�2�÷44�~�,�1"�����Q�'�4����7V�+�<�-pJ���z��Ԛh�Z�! 6�*~�2R�aDZ�њ{�ƫ<� �t�Ie��r��$��
`��]�����%ޫ'���&5�]ZS5sқAk�	��M�y��{v��0U}SXWd	bL�G�����
n�t����k�8�ˣ�״�ل��֌�v�h{��x��S�Gt�M6MP*Xc�]�i��A��3��vq|�v"��IU!Yx�8��n�aTK0�˃���� 1RV�Z"�V�7W�h�h�b-ł�*˂eF~Mru�Q�vݰ��ϟ��>g�%��uA��@)�7��D*�����g, /᪓J=w��W�G���6��d�]�O(u>q���0r��p ���7�w�rJɛ�5xM"��S$[SY�����!9bn��7X�q�$;:��dd�$V-5��G�K�k�c�L��E�]0��U�mQ�8�aD--��v��_˧p=�zN�z���#��a|8b��Ҧ���ϩ��^�:���IǣmH�8�E�5�	*���	({�"�0��;���p��+����&V�S��:(h=r�/���6�L@Z��).�+"'?5���S��3����~��ʟ4T���<Dm��zP�=��aq!��)9� �z�����������s�a�a(����g@-��'���L��MT���]ow.�Y:��w��W(�Ch�P����]�Y����F�l��K˖R��~g�O�0�MR���u��6�0�ڶ�/�"�j�4�q�H9��j3��^8W��C�<Y̟�M@y����1u���-��Q��7�����.ר�t%�)�',�Y�o��3dmQ�+�4�+�vA٣�0ZK-��K0�.A_,[��#_ｽ�+�a�'侞�a�
'��fi��Ş��<dN&U,��sJ��c�-���>ĉ(���%��x����
H�zvE2`׉�%v��E0�sĀs]�e��&44�Sӗc�ȩ��S;ݴ���c�cKv��%!���:"h*�� �%�e�sS]ۂ�*���c�9��ٌ���3��CH�u�	z�Bއ�)��>[��q����x�I�XFk�ej߄�N�U93<9J?��`x���g�M}���6z;"��:l?�A���=~v|���N�1��X岼'l�o�X>�v�kB�e���y�������@�[��'X�'���N-ƥD\��E��8��Y:t=�����Rxw��V�+�k�a��5|���^���!
 RE��ے:�N�dm72 qqK��]�cIZZRx�"��Ѡ�X����f<f���a>��o؋���(vѬ�`�B���a�DX�-"�u�[�l�(#(TV-u�U`J��@�`;s���_R����q/���"i-	I���#K�I�b]��Ԛ��/�kj��I��n�+���tj�(�9qS�LwV��ؘ�4�ɳ�F�h���9f%�{�Q)P�=�!��0)-�W4X�*^����u���!ݔ\�kR�R�?��0����`�Йꩄ7����n��������O§q�- �U��jg)�:�� `�ʼ�2+���Sx��q|�i)!�����ŧt�u�q�<c�n�>D��|�0��@�o
�3�̀��S�Qy2�����N���3��)t����r�����抧�=u�I�z#�����㥭���yP}zV�BX�l/��p���t�\��lL�x};��r�ӬmRO�M���DȜG��q�d�Sv�Yw��`}X��kH��B��X���V�d@�1�7IC�ϫ���wP���y���U����R�/2���98�ѭD�d{t�ɱ��b!� \���^T���}l��T*��d}qve!A�ƻ��\�Q���M��?���NF��*g��z��|r� !�����&�i�W>~լ�4a��YK/.����7P��"�p����� �3�'�����Pc媉�F𳆑�'���aZiK������+s���fL����`��*c��,sկ�fb愧Q0|pI�A������/��X�M�����C���X�yv/��%x�UX�i&�2���/�[��g����m��beB��3�r#Py p�j��4s��0�K>�Rk�+՛a�cQ�+uf��0�����vc�KҠ�O��}J��p�L;�U%��>+	�e�+��"��L`����>Z@�$ݐEW(}�U��(�y�Ԝ��6d��eC����%�v��;������ �}����	M	��~;zb�#A��t�B����cw_Q��:�}9~0����"����hP�� ���K�EHȳ
���/_��98O��V��΄��T�.��'rm� C���~��$~Q�!��q[
�m�F4��=��]�O(k�儝j*�5�\�	_�y񰡨E)��-�ŉk��&A@��Dz)/L�q������h��
8-��K\.��:S2Tϗ�����-Vz
��T�Z�u� H�.�;A�;Aj"��	���-�'��4֏x%��	|]W7Y�e�O\�-+2�>;j���д�a�UA0��*�-u2�$�H�	d��}��Hq\�z���]�1�n��L���y�T�#i�C)��aO� ,��c��*����]>d^��NG�f�I�
�����[�����x�����N h�_������M@����Ӥ�2>`��&��eq��.{�7I��o����4��â m�fz�l6_�'�#��,����P��O�$�;��W�%�h��S�-M�>�xA��8sJr�C��E�w���a��W��ҋ=��h
���2��VoW�:d�!�0@���0��W�ߜNO�z)"�7��9��:�c�<X�����Y��/�D\��츆�n�h��i��1�Kqy�8y��;5k�h����%Ri�c��D�M����d��Ir����f�^�/�)��^��,�(*�'�St$���.C�-1���[@D!���Ň�;�� <!�l� ��H�x{��tVt��N���ݽ����� cʙ"�:*iK^΍9�2��+bG�osn���♏ր��V��:"�Ѯ��bk��ٌoſ`b��Po?��m����5�e��*B��4we`p�MX��.�0���6���T?���v��_�a8�Rn���{�b�H"7��p��L�"��H�N�Q�6����'�k��9��dy��I�@?����_�>��lmH���g:��	B�+pMb��>v*��B����:�I�PUfҞ�[�:��U�%x��b��-j����B���+-|7�s�P��b�@l&��/3�7ut��Al�dAnM�_}�9<P�8��#Tf�JQ/��d<Y�v+#�Ux<�U-�\��C{���w���ú�U�c�-�Qs��a[�G������X>T�̭��M���S�p��>^,	mBժ����^8P �	��=�i;��3�9��Ͼ�CI�e�.�jX��M�>�?�8}\^���!���=��f(�����m�m��L���DL�� s��M�@�N
��f�i�6�0h���s�L�+�+B-����̜�%J`]m������C����"�{&B�h=�75�&׹���K�@
���*a몬j�@��d�E@s��~*i� B���(.�1dՔ���uѲ��)8���r���$=/�`﯍��Ľ�6��|;-jݕ�K�d���	w���`�L�X2���To�aya�(o��,��JY��]'�w���-�un!��9ѧ�m�Or�
�ށ
�1�*zf��2�V�̷S�Ѝ?!W�dZ�OJ}���$�4�� �{���
���6� []>#�J���N��1�
�*n�S��̶���G��P�/^i�T��/,F�"`0y�VPv�$�}� ��DG:Bz8^@M�xl���7�$�絛�~�Y�7����#��5�@ �������#RB���Rә2��-#�~���Ja�4y�D��~��2��C�SC�-���s�Ku�}��p��M�Zk�J����3g���u�|^j=�����Ņ� rT�o�@uG���ދq�Ȃ�Ɍ2��������T9�d2|ED������C!�5H>x?o �zs�D��ψ̽��_SJ���u`���ж7|O��b�P�#��9�v�5�9�3���>��z�0����|�8���G@�2�:�1�C�g�|> $ʊ���cڒ=b�bP|7k;;W��ȓh��Q�g�owB���� �jJ�V]�C�C�c��N���9K�T$�h�	b�����/5�3��?|Ŭ��j�'yZa���� �+��ͻ*n��fj���sz��F�H1G���k��9`��kΔ���t��w&h7`\�ق@J�:���P�.��$��+J��D$�V}D\���h
�f�'��di�W1+�����͟�>��n��4����>��`1@n���?˯xx1�%��D�m��������l$���S�ՙu�/�3�v�Z<�*md��E4����Q;��㦢W���&߬�|Nk�Y�C��KX)]ٙ�M+T܍�
.�V�^��/֬n<�x� ۬q�*��l�G���tR@��a�̾C}4�#Ķ�]wǒ����naݚ�`�IU��&���ˣ��LWY�զ5_��+c����W��Ԩ�UsUr������dP��{�{w�4R�H�)FX��ˮ�⒋e��:��)���5o���A7,�g�o[�y�`��Pm6}0��\�c����X2�ĩ~;�g��Ξ�0�%�E����U�$鸘�+jR�Xk5i
L$=a��_(8��$%ǁ �W��H��������x��"�`������c��Y��4�����`g��f����������:�*7��F�)��҇n(��:���P{
;A`\��<��8>y��(���)Z���pC%���񿕡j:ϹxB!E�ݛ��#k����d�HW�
!�tظdNm,�!���1�t0c��/{^�υ{�"�Bc��]-���Q�g,���]�)��
-Q�����H	���]M���M�Dp�ݬ\�gh������~����^h��jP��!�x>Xb�E\-ߑ��� �?R�1�9�c�^/��V�R���7����c;����]4��U]Qd���9Č�B��L<"�TV[���3bj:ւw/�͓S�&a�Oy�Bb���]cTݾ(�ى-d�E�d�5�
�_��$d��&��p�u�w
��I��Nw�k�oN�����M	bx{c3˪�cٚir�F�!�ޘ�t����o"�C'wTh���<�B�`\��5o7�	�j����f:�w��cp$�qc�{���xav	���R�<�%�_�X<��	��B)��y�K�xTX-���E}	�c����x�`W��K+Q-E�>_�W$���OC~��З��ç�l	@�B���h=*���B�@A,/K�4i�f�[��Q������Y��?V�aDp�i�y�0t���'1�F-2���a�E3�؍ԏ]xS���m�F&Ybo�&9}��q��Ӏ3��%��XKL���ݍ�%m!Ba�D��n*��/�|���Y;�Y����^��0��I���=��wr����6�Y��� �X�� ��?X�%���ܛ8#F�zğL�&8���2Ck[m射��^ҤΘ�,4��ł�����*W��I��i,#a��}�~��?��L�3��j�Z��.����yGv��N o�q�ըm)G���D�Z�zn�#�"�o`���h��4���5���AX�����>���f#2_�˸_㪂'� ������"�#x83�W���������D�!��r��`CR91���FQ�V�� ����Nc}��]	�^P�f����f��l��v�9�fЙ[����ݥ�����p�R��ɖ�S�}@hO)��>�4S|��ߞ�nv$7����Dr��U�W�9&t�9��wXN�@R�}�> ����9=?�����
sCU#I�F��=w�g�Շ���ˌɠ����ʣ�ǣ�6e����:�H�e0D��6���"�.�U��A���1��g�6�����L�P�M`-ʞ�L7OB��c��&%l:�~2�a��頴}��q+��k@�1��J����u=]�߀N�i��Q�	,{���V�
L���D~�(MN�a|�)?��5����.q��ÕsT?cr�q��tq��Q�<A��8��E�C���F'	��*��a�[��eo?�����~F/���#c=Vf��=R�V[��6�{~"#���,$F4=a�5ճQE�2G,(�>T���<l���{`���֜+r~��=e��@h��cdڂ�"��4L�^��Sm���P���vct|�D�S��+G�#8͜"A�.8�<�@92O�j�\ȧ���r.i�h:
�VY�n�cg�,�wh�L��Ϗ65�P���].*��a��b#���E\Z�eAמ]~gM~t�=�)'Z�"����UeƋs�R���G{Fe����J��F6�-,��PΕ2�P�U�M6����[p�6_�O/U�K$�#��^9�� �^��]$@e���6��Й�+ɬ�0�H[�)��#M\�-D�|nZNd��)�|�4/u�=����gY%ϋ"IB�M��i��oҚ��R���+���׀�[7ӯ೰Az�N�b���'������ٍAv�k [؏wi�N.�ht��`Wf0{o���y	�Z�	yz�33Hϰ��͕���a�vyc��<J1f�-����;����ֶ� �bpwxU��]��w�ߩ �b��r-�3��3t"��z�����-�'�LW��9��q,�?�+�FPE��=���瘀�2���QV%T�����/�O��Uu�TG����E����.�=����ǧ�//K����F����IA��}�a��%�idޥ��+�i}���/��]?B�/�n���%���e���d[nS�!c;�/)��{���=����d�L���#�G��!� �|X#u��?>�z��˼���mm�E꼔B�0�nӡ�7~R��JE�^=P�(�QO���a���.S�p�"J�.�
c`�������3�V
>�1��=�6upGj��!�*�{� �?h�~��)}s|��@:Hf�;<��m���	��tX��T��x8i�ؾh=0"���b�J.�EA�~&��v�>��a ���މ�Ӿ������&��8�oާQX~l��h���_�ĳpI�p��/.lH�"��|� q�)N�t����N�i��t�0�'�Q&���Gat���-�ڇ,������z���؃�"݋w�F��?ߏotF|�G�����#qT����Nav2�5n�@�j��'��0��UL*������9��o[(��ڇ�³����|���叀�G��f��(��Ɵj%�G����> }ao;K��K���>��;�eŻu% �	˩a��`�T��ė��?e%��0�5������~S�0�=�}�8H�ٜt�֭�����L%����0I�:&�O�*�?EV���ߡx�S��dv�
�PC�}e���j�����[�VuvG,ar��>iJ�Ycz6���7���K�_4������q�䵃�a�dT])ńysJ�(=��hG������疚��n_�`HG*S5(����զ�yĥ��P:��d�����,&K���J$�2<a�`-cdNU7r�۝�=���M���Lh�`�ju􁁆��3h�Z\�з�Z��@K��da���3�2�|(�XO:u�]1пYqV��չ~��϶�~�!��2d��˂� �6��>�=�\�|����)��m�H*zB���R�-P�1s��?(Ψ�xJ��o�;�\۽3�z"��b)S�Q�Am�-���N	g�H�oH.�y��æ�;˫^v`/�Bf�S��Dp����[��ޚ�#T���)99�c�K� vB3���ͭ�2Gm�Ʊ��R����)�\D�X9C���\~l.º�Ч8\�X��4�ϣ߄�tn/�Z��Fc��e�U��-�F��L�PO��J�^�P�kK���1� ��� D���X�}�[�|�R��z9�)���c�~)��g2͍��^�nbR4���W!��~���+^��s�n�}Q�è<96�Q��^=p#�/Ώ+[m��g�T��ɳ���.08����;w+m��qA�St�3s���j�h�$v��'�b�
��^���!ƏK�B�~����Y���hn녱ɉb�}o ��P���d��.�M�{���
o�a��,�s�!N���#N2}�� ᣙ�	%�� rb�ɂ�VA��[q[�
�K&����6���d&�I�@\�غ�pBw��X�����} �-i���4���,j̺ �K�oC��	����&��.�a�?�*�~�$�a�q��n�q:��Mgm�np� E�Ld�#����N�2�o�MK�}�bcI�Kͬ�צ*a�=�Ci�N׀�(:w(�d]:q�w�4�.��Tn�l���a~��+���/���e��H���r���Ĉ�o�5BK& 2�5!�v����z����^����i!�z��	��'z�I�֐3fs;���پ.��\?L�Ϊ��2�t@T���[���	*5 Y�"Eo,+���H �L*�eҙg�
T�4kh�myFw��Ļe��D^7
el��j3�f�6g��D��c��2\oR@�^A<�ؘra����f'�'�J$C�rmp-R	VmL�
-�%�hA�5o����68D��X�>�+�a0�m‶�_���;ם��4$���(�T�Vk�E��w�R����}�奼nH�j�V�6�~�Q���x+E�Uw�sG��59-����f��ČH�?/�4��P�����-a3�Q�3��a�b���BC�|S�u�wN�>I
�O^4�سe�K��R�~��0� �J���1yڽI�zeNK?�y�G@؈�;O���垌٣a�f�K�c8�!��^s�����m�|��Im��e����/?�d���	��Pn(��E�80=+^�����L��R��Zt���;���pt�c[�{ F�"Z����?���������2���p�غ�$.��fJZe��-6u$�:̃�v��n�փ�>�eH$#�Ƀ�>+h��;�h�9$զj>�&��)�R'5�t��t��'��z���k�-��z�b����Q��|��T ���#+�c�W=gm�7L�aG�p��2C{�)��f��835����2��	3���?��pL����"ԙ_�p���?[�wZ"4|?Pת">��q���K�4ZE	ʠ�#��Y�s^(ܰ�&H	;��Ж1�K��AV�HL�;ĭ.�:�Ԇ�#"�I���;�9��w�[���)�ɊEc3�%��5�����'�������GҤ�8蝹d�_*�5�4�阠p7�"���
]�/�8&�H41ӌ�Хe�(����+�,�J��Q޵�6O����$Spu���z ��B���W��<�X���k�����h4��W��J�������f���;���l�^��U	61�� U��E��}�cJ����3m��G��,~[�j��hn��sӈ�,�lU s�8���(��`8z���+�q*�����_��B��l�Y=ٕ�W�R}���괦s�W��/�s3��Q|((�

%75I)~%�f��L%�tq�dZ6�����&�j�R��w���1�B�j.O-�
� Auh���ßG�?���?DJ�{y��
�~b���2>XN�m�i6���9p(�/kƤB��ͦ�A Fe�\�g�>s����C¾��8����0*���ϳ���3p ?X�>�FD��G𒙢��tYI�R1�Ԅ��a���W���w=k����鍥���㵪~�0mmݱ	r�l�P�n�m�����r���C� ���$��_�����2�-�
��z�P����\űyNG(;0w����T�h^g$?�z�͏TQ�rj�z�x�����zV��ϣp�/8@��Fjpf�������9��G�H+�}�,�K�z��*��R����ӈ(�*�cㅲ���ym�a=ǅ)���z����LQ'�\�G��� 訝���a��Ѱ���.0܂*���U�@������[�������k\�ؑ��A"*���=��S0��6m�ݛ�#��q�c�/�'�����C����۱ă�R8 �)� ���ۭ��LwFNᕜ��d�L<��:-O1Я�Pցm���;/4k�D%/�����i��q��s��� �fm��~&5ٟ*��U8s 6>V��ش�$њ���!ௐ����I�Uw)ǔ#g\a��A�I��w"< ɟO�� 4��E|^���8_!�|��U�R�Z|��[���A�:v=G :=b�1����Q�RS9�v��@5�r�$�c��I�~�,�û�յՊ���P��EC��W�]��V_O�S�^y�d���d�H�lSţ}�*W�չ&�b�ig�x�4�٭��_Q8ʏK��fᕕ�Q]�����dG�YԹ�Pz�����1���>��d�ކo(�7��H�ݗl�m_8�}�)����_&zF3�zm����횚���5 Tt�"�d�Xjn]��bz�czԊxD�2�>f�x���C.����2ڒ��c�I,��4GJO�}�f��j�	RJ)��H�HC�IRβ�|Q�=�j(���ZO.�Y�u)�~�t�$�~�J��Qch��YC�F6�뻆���NSoDy��
�U�z��X-N�lu�H�D�9zhjIS��"�-��96�
R�|u�.Oa<2�-1�IrU=ngb)0�xH�
õ.�e&�f�Y���{�JnF��벚v�R��V����A~�7����7�ɍk1���}+���S��$c�-�Y���?u*Ad��d��'Ɯ�xU��������l;��9�[��
�|���-��Y�[m��+��p��e��l�,@��,��I�f�$R���9u9f�:L�f	��a�Y9eᶰ�މ'�֧�ߏ=I�V ���zd����sա�X~`�%�y�:�6ss&>����&�X��#�#�!�>��-�D���'������6.��R�8�T�$�\�_H3�d���-uh	@A�~ �R?*=
���ȣK-]|��(��(�զ�J��1��b�ϟ3��P�/�'����'�u7>6��{$J
���'�����3f�y��m�Ĺ�%}.�K�S@����&�$�I���*'2���|M�EQz�+�>Dﴰu�1��M2I�r�}�a��_`���ƾ�_��ʂ�";�xv��gAB5 ?T�������N�����x�Z���{} �����iVG�(�&��41Γ���.����'�v���L�#�����I���c�aS8��%Pc�ܟ��D;�Ij��I��X��[�$�ק�?��p���?�A�|W�y3�����\�#0�C�?ϛ��EX�]�>)ᢧGٛ��{�����e�����O�UU�w�l�4%����f�~l?C�/r��ͭ�Z�,�<�k:~��Dt��^��G��S�Z�
�G���
�:\���%w+�Z��ƍ�� �pbY;0���0����;��fy�Y3f,��h���PF:��	����[q�=7�z��Eq�ܶB�:���ג1���5b���܇�n 
";�-/F���y���X��V�6kZ�������Ԛ1i�?��`�7�
�ɺ�nG�X4�n�h���z^�#��v&�	�J�+��D8�l�� ~��{n%1��;��x�^���EŲ�8$��s!������t0�4i�+�#�Èu ������FX�`����?�8i��Psj�k�`=X��-/" N��Z���M��/8�7� �tݟ�1�R����k{��'S�#�Z��I\*�Z�^�!vn���Wk�RC�|J����хx$� ^<�n�<���9N���c���i�֞r��'|�i��3���<��y�deQ��@�\��Ax�hV$��e6��. ��_
&�7�@�ۑ0a��Ň�q�N� ��Cf������%�^�dfM�6g�@ ����Y�wWo���L���=��Rӌ��f�I�_v."X9Y��U����c���K���m��B	�y\S���-m�c̓M 9�\���
ywF�g�!*mG�����8n�zx����w���eJ�g�m�e����2PS���/���]���16]����Fs�أ|6�(��j~���*���WX	<�q(�1|�U��M���w���I�Ă^$I��$� �	�?W1���K=տ���7"u���RV�ۜ��~*��e6?�j<X����`xd�����/&�O���}ea���eά����5�����(��en������ ���/���kg���t#���"�bW��A�Bɿ�t5� b��8?P^�t�)kgR�{NLA:�}^�4�&��	��O�Z��4e���/V�8�hu�"�8fI��3#�GiT��<�|�O�=�ԲMa���@9�䡣Vt���?�N���*Ո5�����b��Q&|�lH7�r?�7r��n���S��Tfz=�):��n{/F(�H����BX��%��st��+��c,�z\\�M}YfB#�y�ܚ�|�]a��&�R��ˍA�y��Rg�[G����]���^��	���4g�HQM�"ߙ���%��^νtz���8;�h���tqq�l/$Τ�s�(�Tl��*� ��B恜0���i�����O9[,KR;*����g���}�͙O�f�T8]�f���p��3jL��_�Z}^���:��*�'��S�M���jR]Ǧ����S��Y��R���Ɋ` ��(I�"���m8�< ��Y�hY¢"Ȥv�kz�8���W�:Tf��K0R�w2"�hNƟ��瀙K����|9c<B1F݇Y�HdW���p4TP&�>d[3;K��F�L}&�#��睅7�
�|���D4r�� ~��T��a
oJ%��u��p� �
m-9R��L�����f9�c����O)q.�k�2��ęm��Y:+=�X�6l��Mpgbysy g�KP$z��>�?�>zvt�j�l�W��Hѵ`t(�-�!���_���+�����Y�jD�����c�χЄ���gGY��B��.�:�VYHu���kࠅ`u���V?؇�:z;�}�Ma��?�>S��"��VܒP���.�ly���X��Pj/�$��4��dX+�-�8�x�2�ȟ�|3�1����iQ�����l�[�]���o��C�ʹ��\ͧC���>�k�JT��R��U�$L����_�E���&{[��4N���Z��&�XQr���~�ѡ����?<a�p�ԗ�gUj�P�W��A�$gN�����f$B-юT����6�J/4�S��ġrm.��2�	Ԋ�ӻ9�1�V�����3t!2����e`� 2�����Qvʹ��lL��f{�	��kP�-B���o�:��*���׌S�a���F��Ѵ��/㑾�O��>F��\�JQ��Vy+p$��6���`�˕s_��lR]ϋ����k��YrJ6�����x�t�y���a��~m�1�?����8A�@�*��'���ԬZ֍D-�J�����Ί�>e>.q�|�8�o�ͽ_�N�����9t|]�)��*���5^�SD0�¶�%�- wTjp/qz�J�M�7�
�!��(5z%�ACx����A饨Ʊ��j_e?q/��0�#9�c��g>�LZ�u|=�6���֦��2.��p��=��<P"c_K����
e�CO�A��o�?�p{�^�3�;�+~[k��{��HR[J�?[hv*u�|}�j�\
��_/M�-�c�N9��Gg�������<@	Z�<6�Nk ru����9W	�=1zBan��/��H<hE��-)����.*
N��y��zd6�$�T$��b;��Kha 8�&����-���Xa ࿠�݃�|�K͂h��U4���iʲ8_-�p֊�GS��#�w��NO��x��Z�R��3!�]'<0�����o8b�k�e��!��Ԉ@�ˋ�)��.m�)-�������-2��]����x#���?Uh�ϖ	۩/���;��W�����<+��m���)�`kk�I��E�mpA<�~e(��S����FO�nꔺwT��ȝ�ϲ�$�c�V�n�g�ܭ��(��`1�E$`n�ıezp���U����]�G�|�tc`�'{��a(o�H�9�dȮ�{�� YW2j�㝰9`����7�mn"�Wn���X��ݒi��'��R����8��2y�{���wf@����8wh�v�Zu>v��Ԑ��+��.�%ү���
���.�͌�+�$b[��b�5v ���	����广�#̬V_)l�L�@������L��%���E�.�Wߗ�2�,d���1��G�0���*uڝ1��i5�*_{'z�V��n��&H��eOn�������TZ�D��)�rL��hSe�Tc��ciqu�>J�wX��S���x��(G+=m�3�������6��u<��E�~Nx�Q���&�Z�8_��d���d���le���p+{�
s"�r�~&~�)=D��%��~��V$͙:���>ƍx�*���ws-e�:Ep�$�������K2�g���_��)�F�K\A6Tp�O��͵��(W}�
��Př�.��WH�2�yʛ;���ې\q~3rږ��]_#K�>����ժ�.(x��ϣ8�=-�7��:��6��.��3��J^�g�{��������\��M�!Ķ2E:��T)d�y6�7��m�@p̺f
�z^L�V@��WQ_|%���YZ@)YW�2�b�:V=���tJ�O�0��;72=��f����3�ņ�yH�B�V�Qv�a�n���z�6�T���cc
��bf q=+��d���9��?�U��P�c�^+K�3�F���%Y�	�r�[n�MrQ̇=.�8��~�Fb���)~�/E����Xn�paT@��QG9�_�OA��xڃ�F��?�u�(ɢ�g�&����V�w�;����{Zt3����,z9G��[�3�LL��)��'��j< s@��s��U%� f" �t�[zT;��EI�����[�F��M���I�Ŭ�y�������I.(��:&�J���c�� �C=��읃x�g'A��.��,$�\��^@�W����Y��� �h�CL$^����WҰ��1��.P�zOD�@o���Q�^���Y�;�0�Ϻ&7=�Ǔ�֨��/�[�HP�T�r|\Y�h�x�m4���$SO���\:
 ��#�ko=��B`���j�m3�ʾ2�`V�~�aH><�	���kjo]ڨ�l\x\c�ٮ($M� ���{Qjq�pK�����(P��CtHfe�2�q�+;��� ���<���\$�����? ���5�,VI����.����5]$5�$e����ͭ��^��M�V��[E�&��(�qi����O��'vҮ0* 4_J=f�`��j� I�&U�s]�^�_�%m,��%ϻ�<M{駛�D���)�m�����9oE���x�B�<O�����N�����@��K�gp��X�RV~�H�u�9U�6\�f���-\�� ���[�����$F���A��ok�2{p�fI��6[�����1)Όg�Ed٠:�>�gQ�<��(/Rr��l�k�I����d���m��+_��D\�9*bBID�Q��T��Y\d�Uv�x����+\(/k73��@-��|�1c��pxo,Y�(8Ub�^����E:�_��������B�'�FGbK����ף�d��0�q���l���Ѩ��_��s�s>i+����S'~f�C�l�p�^XY��SCC5��X��@��i���j->o3��`�}����=�.J,B�g�z�r�ܧ�7���x����ة�\�8@�kau�����K�,�\V�|ܗx�9n��E="`��a��7o�Z7>G^�qV�f:6�k���
����R�L�!�rǉ�i��V�R]� /2c,�����^c�L�؀5�c��t�"��gA����X�E<�PVx�epQ��w���.��n��>�RB����Z�����`w�&��g1Ѳ�: S+j���A��|�Z[ڽ�8�h	�N�ǵ�k+�7 ޞ�U�A�3�j���������J�*�����.r~� ��X�/j����W �Z=���9�hL0�C�i=�d�i(91��+a��r�F�~JLp
�ߎ��������/�'���OnOQ��)��[�]p������&���Z�/��2�2�Wk&;���W?�y�b�}��W���K�sg�P||�pާu��d�����9�G�m�Ƹ�r9�/m:<	E���<:�O�uSe��`'�A����wF��1]�4�k�v���U,"8�)��H���j��>��	f�:E�����e	k%E>�.�7pU
�s���>�+��> ZHiya�,>~�j���Q����8տm��J�\ 2����\(����C �	�Ƀ$]DI�*�1��ծ��w\��.膆���u�kP�م13�2w1�:���u��e�=�0-|���KCݖ��]3�ډ��[�Rn���g�a��+����e~�dgKK�.�/�zod.Z/n��I�^�"��[��j�̑G�+�+M_X��v��g��������th��^x�Li���(ohev�Üs}-�"GW���8��)ؠ���e�S�N;��e2%B�b@�0�ԋ%��FAfSMr�m_-30�ڦ~�֮|��ڏ��Ɵ{�=�w����$VB�ֺ|����û�s�q�V��M����!�+��.�b ��7�nc�@E�!I��?�q�>2�K��\rf��',�HZ��)�姻�Q0��l�����i��'�������~% ;_R�Qn�J�/(ٹ�w��/6��S@��̔E� �U��ۦ��r�b���]�j^��Ez�YO�"� {�m��k�.�JA�DP�}TN$Z`QR<��{>��*���f�ʲ~���_�(G��q����S�n�_%�~f�d]"����J�0B<���HS+� I�ߕk}*Od��7�V�-�0��| �	i��:�fPR*�*M���r���Dc�^�ޯ�aL�_�;C`Ӻb��]H:׷���En�h���d#����0�e.Rl�G7]����Έ�$q[�Q��s*���E���sd̜:>�XuLl3�	�^��
�GJv�~��z:�w��L��a͔���F���B+�4;0[���Q!ǈ�<�*�d纖����*�����n�1Xzn](f��y��(a(���]� ݥ�̽d�|�uR_d�t�B�&��>�
���������5�t5M��V����o��M�Ԥ(,���\ѯ����F��p�(��n�}k��+�`9�hSII���"��������K�'��4�)��{v.=�U�r�앜0���Bc��1?\���F=�q����r���G	�_�" �_�����b*�Tc4iR���@t�c����)|A��S�8_�%r���}Hx�o^�D��uD�l�9}(�����G@}*��%G8z_�aD��BE��x�Άz�<�\R+�(���{����������'��#mp'������9H�{i�D�	Y�,P�T�k�q��Auhȉ1�.��]�PnYk#3]�wZΓ�G>-:��JҴ��&X���(I��8��qm��a$F����-��bY0��'>(3�B���&��l��;���b�ǻ�Qѳ{Z�)k�o�����^|�L�"�O�����FL��h�yy@m������d��5ި��n�*�/"+ZT%�����I�G�ӛ���f5>#$:�+TO��H�������^7����	.~q5�	�(���Qx����n��[ ���iD.F�v�GJ�K��!�Q��������,0�m�e
���G������%������h��4�L)
�@����ʩݭ��Xy�ݔ/T�>.mW���Y�sa�+��ޮWZ��V�x�f#��R�Q3����)pq�j�����l�U#>�$�>��P��������Vn���Z����vN��ڝ	�U#>_:G`��ɢ�V9f�D��Y3��/�v��1+M\�/���/�?� h��^8%#�ˮ�h��S���ܐ��2�5^�����?�7����3�#󃻈�Fn_�<�83����'@�4aO��q0%�����w0V,@���{����q��f9i���2�g��Sy}Q�$�ڗ�,�$��60<N�'T
��� � �zA�H����<��ǢK:�BR]m�;V?�����?ӥH����i�,	��sT��9R P���|���-9A���{�GTk���+l�{��O��pe�.���*κ�BQ���C�C�ѓ�8����a$o>?��5*)��X�Kb�m�;z�x�4lCWFA�,e;V�[W��%���������op�=��m�mþ�A6'Q�y�+�=2?	��Ee}�n\�z��1��v$�V��IO�wj�7����B�C�T踿y��� ~�����
���E~u�tAY	t]�^{�䊐�������.�����["R�s�b'1J�[�(>����z�E&�HW��͎"t�u�	����"���ȋ�tY
�MU�I��1���+_.�k��[�{P��:*�)��3wN��	���R/��z9��v�	w|5�2v:�G	�AM��������|�I/jI���T�T7$(O���.��EbI�;��+��:�9rO������8Uut�L�`��� ����G��#{��qH�SŽZ��0�KT���u��GTQ���اwQ��5��&��И�s%�[M�X�@PRmx7@�V�\F�׈qŎj���p�����m��S�Q�v�2����=�'���P�4��+��i>>���-Y���?c1b$*P�Lp�t�-��j�'x�u,Wכ������alM;��y����Ңݵ!S���C�'fsk;&�Qp�9��2�q�F��$1��n}\ʐܝ*� V�,��cF��$�VB��ͧ��"�;��׾H4*��-Y�2���y�N����f� ��y�?�͐��KY������O�iN�>|Ѳ�t]�ׂaq*c���c�-d;	Z	�#�Q[�^�K*2�E��p#��-�QER e��i��>b[�Y�YͲ���<}߫�k%GϞ'���Elq��y���$�u�r)���.��Zj$rx��I!ki?򃱒�K�l-.􄊂�@���1�������v���cI2�5T)�.�vM���Ȃ�|.��z�����/�&����r���J�g�oc�(z7eT��dJ6s��*ii 1ih�����;�֩UNB��
��$q�"�6t�$.^�.O��+j�w4�G�e�r
qd�xS�@��/�^�s��*UQ	7�y��I�Q�Rz��ʯ�:�|8>S�'t
��܂d�Yvр���
������4]bϊȰ��r+�V�����=&����mTĚv�ZzQU��b�t(O�M�����)G��NmJ��8��-oƳ�X����oN�a��S���=p
�X�ɔ���4Í��Җ�Z��ǓB�����%���w8�U��D��&�&V3].l�伟��α��ÃIZ��6�����[O�倛�D�|�Q~|ICQ�ٔ(N;��Y���[��DgQ��9n��m+Os0}�*�i9��E-��P� \$�x0&�/�-D�f"��杣J(�T2�@4�x_h��WP4!�d��C�8�$�Ӓt�bWX]e>|�qv��V���bQ���g>632�Z�G�ʄ�Ѕ�Ŀ�b�Ė�3U������ �uI!)��'P$b�f��ߺ���@P���;��kK��@�xfۏ@�b��[x6�����ZZ���铆���;�oNT�JF~VQn�ob����0�c���7"f�6��S�w���3	���l�VAZr��Q�p*k��^�K�."���A2%��<����O�>�#_�'E�7��-�qP��~�D��7]�cI��jD6�\�+Ϯ�8����$M��#e��7|�]���j4k�`I���䀨�]�`..1���S�T�
�G��% �U X�!N��/�c͹��Ypi~�eЋ���3E�R�0��\���Zd�����ʧy�h*��@~�<����@ypS�.�?�_H� X}K��ډO�	ؒ���	����¿3�"f�;4�3e6�z�}�A�f� �'�/���moL�����/!0,�y]�L��&��
�"U^����A�a�Q9g���3�N�$6��\�L8��_C��s�&xI�~���D_bB߂kmt?p�z�b�]��K"�^8h��`��������z�	��Y��(��+8{���'E�UM3��7�So�����x?��$�i?Y�e��z\R�h6�%�Q g� �9��y��o���rL3*T?$�l	X�U0J�!�9XG�?A��&����1��k��:�lm���椸�`���7��e��J����w|i�8%�h���F8�'Qb!r%��� �~��y�]�|ry�k���gߥ��k�7'C&~��{�V+�|4�ȅ�<���v��U��L�`2��Zp�c�����j�V�[��_b�G\������	^�D��)�(B����5�m~����F�t9Ӌ�ಛ[Qe�d�>��I��g$o"5A Z��=�{��0*[��򽞢C��c���r��	c����_�z#pY�9��V�+R(�]����c[�~Y�S~io�����q��)�0y� �S"��j��3���E���u��}!�@��!sl�KM���Ji](�_NE��C���|��_���	$��Q�f���Я�5���,�~ �;ȁ�[���yz��G�:�y3[��@;�9��";Z6u_a��� ֳ��Fn�=ga�������k�HǠ������z6�B(��]�٬Xׂ"�7�i�'�M�����z��b1�W8^�pz�O���+D��ol+�DP߷s$��>����7�����Y���"(��R�o� +/#��v �%�{w� ��d��������fYJ8k���&5a����{�@�N��Y$�7������]*_��K��x�wb�l���Y��5���3�nd�����z��$ �t�fQ�x��P*-��O��J��n���(-�?��P%f�h�v#M�<J��8Ӛ��V]^����)�d��c!�<�����c���s�ԯT�n'�]B82�펄zp���W��Q�����������7��˶N�`T�W�F�:�7�W&EX��e��� ����:�%�HZ%Kp=%v��iU�}϶ׂy/flN�D������[�|�w��0�	�����g�^꓇L}��S ����k�^���9�b�4��ڙ�@fE����^tsI�A�x���À`a�
��=3��
ā�(����^�)~F�4���s�z��	F��x�;���9V��{w5��5xN���{�ivڨ��~�{.�/+ݏ�a�5�o#���y�h'H�%Һ.]x���`�����±�v?�Q��bm�����q��˯Z�!��'�������By���8QT��Co��{�Q�Q�Y�+..Z^u�Bb]<����G��_�D\(NE�@;="O��Bы�Hm~�ܭ)����M���������~�T����(������{�Hk�� �����J�0��Z���Q�郱�~~K3� '/E\���:��P寢`��=��`�����Q��d�׏�;��|�.��E������o��;0���0�ϳ��fT|
�dE��^r�9O����XEW����~���ʫdd�b��6���O���֔c�-`�g�m�q{g�@Z'P�Ύ��Ȅ+_i�X��z�]�ꡉ ��Կq�����Fp���Dl�<������Q�^�ɹo���ST+���4��N�EQݼ��I���q�CQS�|-,� �dl��5˻�~�XXu��-Vq���^���0k_\o�-���S��~�!�<CcO1Pˉ"Ju�D�%R��s1������=���1�ʁ��cTh`�!���{��
�$d�#�W�T ��T��m�<R톻���Kc;�g�e������,��IMO,$��3%l���Щ��A���F^6ε������t����:CT�=;�)�t�k�
$nZ�v1݄������l2=�#@6������7�b6�	��qv����y��U��'�#��T��H=ZxE�Br�C �hޅh=cy��eJQ.��ڔ���Ei�"���C4��>|=���3rӎ_lзd�TUq�q�<�%�w��ϬmC�,8��ى(��ʹ���+��JKux��.��%Z��jX����$m���p�����I�����r�Ll��i�pB��G�Y�ƃ>֝a9t���I �/��0�#�K��E)س�|n�pz�? eZ X/�n�� �qٓ_�#^Z��e�";����j�:Mi스�W�(>��w�W�9��2i �N�
n��)������/o���d���w!��y��.,/(�+� ��"W@�p�
�a��),����S��BW��S�����CeR��	;���O�0�
�q�ihI9M�S)�M�I�Y��xT��3�S�p�0
����5��Af�Qe�z��u����3U����䓬6�-nyT��S�#�4���^���qu!3���������A���@�@�¹Y�B�8�8L������6Q����#Ȃ�0b{�F�$���~o�s��X:\�S��V|��#�hNR2.��`�i�[ �I�れ�rw|M)�B/�:.^�F�Is��W���ǆAٳ���$��J��j��b�c1� $�֖�ps|.�Tx�)c��k�P�����uB'�k8�`88\��A�d�^Y�Oy���m����.��Y1X��>�VhBb8��;�]%��f�����!u�IQ�'�ڢ�����QȰ���
�	�j�Ni�ǖ�}{pY���X�6F�U�m����Rr��{!�,�,�AZ��|��r�;�SτA�)I������Ob�~��9b+/��.�f"TҴ��K=�λ�!R�5��r�U��%�-�
�5܂���Q>A����C���e�"}�è��YӺE��m(y?��W�i��bHP�S������ފ�9 �;��� B��N��ɯ�)�h��zY6|O�x��.��fhk�]�8�DF?l��A�w��sz1�����fw��^g�056�Y4ݣ�c�P6p���e�kyB���{S�5���4dR��Ohe�X|8{�sn�X��/[Q Cr[x���O�ό^.l1��~�o��D�f�E�h���0������@;^l���{<�m�����?��?�3U��N8�Xl`��p�M�Rb�$��O>��S_�9�g��ۆa�\��m������Os���>	�����7�cbĖ���]����]Ф4��k^�h�۲�]V�tD92�ǋW��23f:|��n�z
�̃���6�d�nvM����$�y&B���d��d1��Hj�&��5������x�M�|GJA�Y���Wr[�08�s��DX�e��b�����y��4�Å��;��a��Q�BN�6����D��u��P�ҽ��O�%��t�F�e]�̂Q�b��كO�6�7¹�,|-;��������	Rx�E�� =�9Ë_�9��<���H\J�B���(vqH�$	�O��Y��I!K���Q�!N��m��iBk��鿹e�!�@�etJ�^��_}�i1e՟��F;�X�0�=�GL��d��ᩨq)C�N��g k�ھX��$�0�j�U�po�9���F�gN2 �'�YY7��N��z�!rd����蔧��N�o�O_"9���T�(���\����
���.�	�|��)Mv+BFz�ނ�������	l(��'�����@�ͦ%�S�,{%�^ò�K[����i�k=Ep�uQ�8�̈́;��Z�ݙؒ�������1k�a��C��M�%*��bJd�|h��w�E�o�O���%�ј��~�<��
�Y���Y@�;���ӹ+4�4�amtu�׏v|k�Al	�k9{lE�	������&��^�U��k=4Uc��aj�4D�S/���Ŝ�&-�uDm�����*��V�:%��!Dv�r�;�&/�uv�+�_.>>�6Pa`�8�wֹU���'���-%����/L\nf�Q��=[���f*b���P��q���M<#��Dш!�t��'@�+��w Ga���%׬�%���?qC��xC1O}=�!3[A
V��tD#����tF��
|;������^	���d�/���aA^�d҆z��HS���hە0����%�q���*Z�<�fт=�l�{ 9N-�Y����gb�+��Bz�|�������c���!�0Vb�bq�`�����r%��ry�ؕZ��*�����܄'��&3���q�C%w��W
<y�j� _�{��,Y�]����~�s������ʙ.+�l��h���m��1��0���l�����sWxݿ��b��G��3�K�%ձ j%���bH�a�˳�zl�G�:8G��a�,s�9�������/{��mJq����@s=1�{Oz��s�f���8kc�-���j/5=:�=�kjwN��_��)?��QLG�M�läyS$�=�Kc׮Fg��}���_�$BĐ�"@�i��#�ophR3�����q��T��[��a�A�ԉ����@�[�f�[��Od\;6�1��d\��N&�	4-7��%�4\
��q�3�Yo�H�-
���I굸�c�$=j荿�d�N�ێS[�Y+nPx�#4P�f�>8 ~/���𔗦x��� ����nO�M�տ\��4�3�i=�U���$+c]D�b��.6wP�d�<B\$�� =ue�=y'$�U+�E��`s����^f��63���F#k���R�[Z;=QQp���l����'y��j6��v"&�n!�����7�J貐�xҎ �X���Bh���kܻ{T`��{��p���1�5m����[�b>Syh��.8"P;hK>p�nh��vq=FPi�6P�/�����bS��M��>q��8���Hc��Rߎ�y9�4���"I�����J喡Ea�>��ݯ�&fIc������^���G�>J�;Q�/g�R����be�D��uo�8�N� *��Ϊ�<��D���#�3�lC{~٣3�V�L�\�I/�'1�����?vR��|��2m�����ur�2U߹����2�a��Q ���jbA���M��嶳�unape9��5�d��ȶfN*�B�&%c<�1l`��C�\���Ό5q��c{�Nw#�X�A�,0���!���hQ�b��\o�˧�0�) �Ξ�G�#��:���Rt��G{RF:�=��U^������@׾,�O��5כ�{.��NCy�M�m��v�0^(Q`KM�ǒ�J�%e❊�7��*�t�~�ҜD矴��V�#R8H>(�>�w��%1�-{�H��R��+��%�c[�5��*�5�c����OklX������}97ʼ6,�&���B�Q{I�]����-�d}�c׍̈�6���;��R�/.�ժ#չӵWHx��g��������Tƅlմ�����sd(��Bi��6�L͹���FdE`K���2v2�?L��{��[���uG�� ��YD�e��<�� ��nG2^��T@p�]�3�g���@��uvf�LXM��+�X�D�����෶�wz������W�(��
"��o	EQ�d��������"��"&���g]��d�����"����w������!gm�]����խ�aPzHMS��J�h\>�Q�ё*b�3g�	q�ԴN"8+������T(��
�*�h��`�<a��\�����!�͵���&i5]sW� ��ܾv����~��8]گْ�G���<t�ejG�@�+�♷ѝ4�xFw�Chja�D�T�)c�q�ۻ7���ڞ��6�]M�K�3����f
�8sj�������2�RMf�r���h7�j�"��M42HwB84X��rp�^�ǿ���'��2�:�
u#U�x0� ����7���MϺ�d�Z�t:|���pi�IB�� �I�|�`3m�Y��Θ���ػI�rZ��I;���ԫ�&��Hr>�x�������,�_�n�_!n ��� �-�ݖBt�HB�
���m����GЬzE|<���c_+�D�<���\��ê���]x����i�n�����_��_p1�&i�^���	�Eyx����(F ���i)%�tw͠<B
�}����v��Z������TO֠���q�@��q%��m�!X���Ì97sf
$M��(->�KGc��(��2#@wuQ.��R�w�C>`)�<�1�Bi�W9�eEx�
h���Ѧ��̠L��#	_�	� GYg�"�k�-�cR�{P�^۱ʤI�h+T��oF)������+QՂ��Ec?�����
�c`<�����<@�l���GuX�ĩ)pP2`4V��a��9�*z7��fܯ� �0���V���&Dl�}\[�S0�$���/-9aMS�Z�6������m�-�ٔ��mv�p�`�y���&�+i=[��-�@��G)��&���U��m��cH�p�	��Јd.9 �}�@�D�@��>����ظ�z�ca���VL�`���?^��	�q����Dx�H\��E�<Nd@�[2�uR��{t�2/J8Z�E���*Ot�Ct��CDʓ<I��y
k��`]7�L$Ϙ��-@ h
Ƥv�v�\�w4E"�����ݸ#;����d	+�Y�eGy����-1� PR�_?O����A�-}D
%�gf��V�'����-j���V >�s�,O36�$���&k�Ō��Չ�S.l��Da%����{�Y��+/��\e\<Δc(4��LmV(
��㐪ڨ����Z��R;7U�O�[���)�#��hs�]�ӖܗsT0���,�zY������(�i��e����Ꝁ+�DG�W�e�[���� ;srV�J����lجQS���
f��:�A�G�X����]+�**����>�$�&ya[��ꀧ��'Y-~^_��U$C���W��-�*���\#T(�̘_'���"3C\�r�o?`��ò=?N�\;��\�N,�w��m��F�7��J0�!����j��:����d�>�˯8'7���H;�<DC��%ܟ�����މ�í�Rp��k��](ű#������8��&��,�u�l��M� ���ExG�e[�����XR�s8�!>��/H���'3𪃇�h�j�X�DZUiɠ'��p��T�9�u��(f����"ƽu;��//�k�r�@�Sm��"���r��ЫMy5fb�
"Tu(���T[t�]̣/�Po�S%.lzC1||��mߥ��/�_�+*@=y�gI��N@]ٲ@gn��!��'ВG�t���_��c.k��Fz"cp)�� f�f���#����V�U�4��B��T��Ɠ�铊`�W�{o��=V�*�dfyO��~^la�-��\uU��<� ��n\������S��-�u?�
�����i��3��?�����8��}�z(2�{9O�>w܋�G6-`�
rG' ���<����b03����򤓨}�,��&s��ķ�yY�Ax���P�`hߨ��Z%���kW������+� ��W�B���ν@�o�}�� <�c3#��7����f��O��qwj�
�h��x�G6�F�+X��$��qx~C=�˜o�\Ygv/(��!?����k~=��ڷ�ZW�LIRܐO!�OS�0���]q�����"N�Xgp�9|@��dQ����سv�r�CD�`v�q-�����,�}=ҍ|%���\�C$��<,��2�����Tl�
�>3���ZK�wĔ	Md�D?5o7�H���!2�P̦!$�����A��а́O;��B�p]'� �*S��X5w���Ul���8B���zy`� s�H���Pz��Yf3�9����]P0 <	Q�P]q�d��~�B���/yd��k2�M���"Ө�}5�G�D���^Ƙ�~��	ZѠW����ß�Y�y?�/���R��X
C,�U��_���On,�F�ypx�u��K?�������|�^�ڰ��&мh��v�v$�=��$��2X�>T�����Hܣ�����[%� v^\ E��D��ңL�JЀ �/�w�Ta�ɜ��\��Q����4@���j��:�O\�9`�!�o�w`�I�{(!�Y��������ߑJ�5"��W��h���C-����&��j�
 ��s��@bE-�vw-� k�-O+S{(0����v�������zh�}��,��<ڡ6��Ry_`�PQ�pJ�%#��������<��]�U��������������'�pm��?x"��0�S��Z�P&X�E[V��}E�"�H�rc[=NM�⛊�BPO�,�23X�×�[�m��Q}�Y�8�8&}ۋh��_�	ǁ�!x��ɋ`*�@��A�ӄ3�����H��V��r�������x@���5/�n��&EΙbg�'T���N���-�ͦc�f�QV��͹���qV[���p����5&�(s�C��P�(���!�%���ݪ��,�
�^����A3X�U`kt��f��Q��k뗛�e]:�bRYcB��z֕u�
w\~�~��'�;bb��C��c����- ���F"6���5�&~�3�y~��K������Ԛ� �.���FkN�KQqp=��� �V�fqҍۘ^�lh��J�G���/������%�
�m��=0(�E :��35�c�g&��OP�Mj0�!Ԛ��_��mG(�
%y�Ƅ��d��@���7x�	�ـ����/�%),��M/p'�v�l��+ON7S�g���`��H�81� ib����hoO|&v*�pӠK�IX�Q�Oe�v�3����dp_	���5;�챸w���V$X���`�_��Gk�S�5WTSF��y#o�����<�M6	�fM�����$fz��g�� ����T@;3>!�t���,�2@
���KiX�1���,�`�]�s��� ��Nµ]������PN3z|2	�d�����Ԯ/!������i�(�f���r����7��H����F�됑{E-��ʷ���r���{`�m~�Y�=R�k[�`wۜgn��=�?�_yt�'G8�w�_�^F!-���E���u$�S�w�#��<T�w5Ǜ� '7-��q�wX�*`yX�$d�p���sh;SV��4/TՐ#����8NMS�)�f������3�~�N&2P޽�lqȥ���I�%K��\�e������R���f&r�`��?4[�/x��5i�7�a���rX�B�	̮��n�efR��{����5�y�'���1�U�bj,�8o��
�L�d���O0��a��쭇�jwv�K:۠��旂X�ٛS!��;༱���I6,�&l�+��ܰ���5�A5|�΍��w�� ���Б���f��Wv�[�b�=e� D���c��	���IK���f&~Z�v%�9G��WeIJltY��S�K���z]�;z��;�����6��x�Z��[������Ĳԇ	�:O��$t���C�� \.-NA��܈��,�&CT�Ä�TP��ϖͥc ~Ja��/z��P��ߤy�Y	�q�x���g��!^�p=>����g���A�b�C�
��9	��T塏�4ڹZ���7^��`��K;ә���vG�0⠩���K�xnUL�*�$������~��D'7e0Ʋ�*0|@�+w�n//]9�oh�!;S�lQ��)m�ÝWǉ��M-e��=/P��&	C�@$ ��/�[�S$g��+=	�n�$�P.�szi�l��K1/7��m*z�g�+;h���N뾩�m+���~��V?^S�L�r��I0���ӆ�l�NI��1%ɨ�<cd�k_�e9�! �	�v55MM8���p2 �!"o)���=<G��*k�26b$@)���`���>�OHLKgR�;��KrM{�������/��5�l����f6qt�o\��(d_%euq���
b�e�s�D7\�y�no�;*�M������Ť��}xQ.\��#>2��s�l�A�dv��rr���JX�}��k!�p� ���=ID��x؍"�֛�������!��*"�b�����"r�Z�.�mX�_���QQ\6�g��Nچ�Wd��Ǒ���O�a��G-�7 �LsYk�]�ƿ��k�|:\|��(�Zip��
���c�ڰ%�O�bm�oM`��)��E��DśЊ���wY}�:oB�.>Xt�����wx�Pv�~����0�M�t��7��������^�/jڣ�L�t�rs�.�I�1$�A��f1": ��+�gB 1�;׷Qdz�(u~�%��ǖ�/���ȹD�3�w�%��f��=D�Az�I�E�N�K	M ή��x��Ǎ�J�M�IR/��l�p�'�8�%�w=>��������|�o�L�[��FZ�y����7�G�{����YS$DeS��G��OT�֫<����RӀ�,��ͥ�V܇7
كm�o�.�m�mQ�*{��nF�<ǩ������R�l]�]����6�S]���n	��*ˤXa�U�m�:,�Z��;����~Qp?a
<�r��t�^�R��L�C:I6�&? �%���o�Tq�!|�s�f� B1
��J�|�����㑜8�~-]��-C�}����D2����m=Z��^����0K7��Ԩ��":��ňS�gL�F���R5��]Qd�Nk{1Uj=����?1���]9;��$mY�O�7k�m�f�0��i���.��,���[�7�|V��A��+ij�S�F�u���E�+�.�Q@��9k8�:in{JZ�x���O�6��U�]�.�aaB�|�s�~���5W�$Vq�ո��@��@%n�ڢ�@Vq|��*���>S�7��,��+����D�b�a���CI׷�Uu�W�s'��9-�x�h���cP�"�t)P���1������1�qI���G%���s4�<�ˑ'��RN��	hzײ���G��F9�XL��κ�H�P�[Pd:&�B%��I�1���\��� ۧG�!9�u�6<�&��ͽ��Y��ͥ�ei?��P����؞��I��)�/BB�6�r�fّ"8�zї��i��S�d>d�y�V=��a0�[K�<���/|�xr|̢4?E�z�]�\Y��z��h�.�xZ�*�tВnΊ���q�K0+�s8���&e6�IW1���k�E�kkhh�̊Ѹ�7��!��R@R����VΖ�=�P�����y����EQ~��'5�! �Z���%P��O1�i�l`߃o�y���q�����s]A)�HO��l6g<��0j!0�����@��U���%y��$��JV^%2�هH�+9������:�N>�:��)���s�l�.y�s��y@�O:f>�s\	�iԖ���s�kAA���_Y�b��s�p{��Ѫ�?>P1���cq�%��{M�;�Z/�>?Wo�J���F~A\@Ȉ�� �����B@�é�v��@�^���ԋ���1�NǸ��ꌾ�?7��Sf�*T��
ѡ�F��&*�!��� zʖӀA{D	�V����b�H�#��%�%�������0�b$�,�mݿ�sM1�4G|��c�1h���x�Sb��,,��Е��,0��z�����@g�z0����%�L-�
�r���ZK7��H������ /����Z�L��R�T��J��rV��W4����,>�f��XA��M�׻�;谬4w��
տN�IL|�^��3�̅���F�1�*��vS����Ф�ҋ�!���l��u��$r�0A����|<�/�������&{�E��ً����w4Jq����1O&�m�v�0�m���_��z��pD"B(`M��*.PAc�� *�6/�lp1���$����{�Á��&q�F�ׇqSS\H�x��A�`u&��3ceWHz��4���a�<*������Uc�c|ͺs�1a���6˹��ܹ�h��͇�+p�z����9�T��mZr����UE��i�w�SY� ��'�FnJ'^WƎ2����;_�׊��}2�:��BG�v��{��S3�U=(� �! I��O�����b�]�[��j��aʀ�(���Pc�LJ��R!YhX�cl��u��1���M��<7�d�~���v$���3�N��WZK�]\��<��.vf�e���I��a<���&&�2Eϋ�M:ؤ�M[oWI��@�Ϣ�|��]'t��E�����ȑy�&{!���F�3���*	�DզI%
%a׎��%�����Ҏ��UoVX|�w�,&Z)�7���>�Θ5��ը\T���2̟DB�w�M 	�<���<7��AT�fMX�[���)�Ԉ@�KKP�w�����:�8�4]�̿�����D�|.c��S�'��6����y�Dy���c��K`7n�s+al���*���n�-о�5>�V���';��QD_��%\M�8� �$��Vk��81��	�S�&N�N~(�����ۜ���͖v�x�fVm-骮�h�krt�/՟���Ԫ~��׮6�h���8I��X�N0L
Dyg�8����a��Q��[��֜�C�߫��]
r���xg �I�u�0c�zea��~�D�fb���JĮ���ߕ�?�u�rd�Wr�W��1<Ng�vo`�%�t[Z��CY�� Y�E�6�~P�v����/5aL�mP"aȹ�	��MU�������uYz�5y�R�R���ڊS���4! �х����,�0Fz@j��0zZ
��x-�^n���s`j���q�mۓ�e��ԭ��c�T��]�+̛߳Cb�J�~����88��|11�Q����tm��Ģu�
{� :y���G�>�b]��:�n3�h�����n��FFO����0�B[x�ֶ�U����k��X6��[i�6��k��e�QvJ:�N����.#^d�7�ԃ�݄��I���d�5����d�!�	(�'A���,f�Y�/�*�:�����K���N�wQ��x-S+{��"}�	s�.6��������|��4��܆bK������y�Tu��6�u,Z��+,{}W$:��� ���߁6R���'�O �fO�i��:��-� 3ڲta0'��|EJc��f�B������@�9f=3�OT{L��"/Gl�+�vﭙQ ��ń�v*TBo�'�@���|�X�\�E[u��jg1��Y�o}�j6I�~�a���K� Hctp��@e��U�|u��P��ڼ�n�X����Z�.���&̟4˾w�T��~n�^�D��������>�%�d'H���������)�&*+�&)|�ы_�&G�Q[N*z�,C�ޜ�2��T�x4]�S��?_�M*��V:��<
���w3�_J<�҆�s��6���-bO��A�e�&d���kn�⇽x��d�	���vEÅ%#���on�Q�u#�E��5E�KZ��L�����!5�C< ��I�Հe\e&�[FB�<�Ҥ>^�	l�g#�6�y�oP*X]j���vSLү�n�քL�j3Z��c�����Ш>�;��Tz>â�T~�k�u��:�pU���MQ��{R*��/~}��!X�ps�;��o7(�p���u��L�lu�{��A�L�՛��@o{�/R0��@LKiPp��ì�wCDЩ�Y���j�p�����Pu��i�\��/e����;�|�v��qx��;�O>f���^��Nd> ��@mcs*��d��"!�r���c�AZY6)�����t�HóIsZa�iӪ0J��r�kCH���>���k���ib���d����㇗�
�y��~�{��2�N��#�횜-���vdk�*M�ۻy=!�t����%�\:�E�^
Tɏz�g�X�J <����oH��ۏ\i*)��k�`�ɡl/���M��[�c[AP����.P�ߊL�@i�<ٍ��l��K�*��%9�|�;�����.��f/�S�2[����t�T�/�#2��l�����H�;k�v�Y�$��@���	P��Q?+�F����EZ�GA�
�%I;����D$4]�r��,���\ְ�g;��?]�AK����o�W'��s���3��?L��-��H�k�!���b/7��H�g���**2����W[>M'��K�C�]�O���3q8� �Y��h�X⯐4`om�`�Pq@�k��KH0���@*�^�|W-�q#���M�������Iwrf]�gNab,%�Y�v�:�:�����[x�4;HY(�P
�$�ZZU�����4��t
����k����/��y���	��{N�.)���h�\0e�e?���[md
}�#��L�'�I??��� I��"S焎�kof4j'�I��:�i�:�v+�q�؋��~֥���Pt<ۭ�ΰm�c�O��X����\w��yԬd��y�E#�&���caZ�I��p��G�(��[�*bO�Y�!�;`�X1���E�c��q��m��ox�l���o���N}�	8��ܔ���Y�����	��g�8W8���Jt1�85���i��1�淂9j��NSM��j���YV){htȝ��6/O�\p�7�\��S�L<�����Iv�\�=X���bQˀY�-��_��<�&Q]h�K�q��� v� X�´�Cq�(������Y���t
�-��fW}�0x����%�P1)`~��O�"��d`��}��# �����{F�S�3�B�y̕Y����w��N�mr���M��^�;�rXG�����5P���<�/N�����G��d�Q��*�.fp�H��8W���Ө㢄.��ꩽ;�9T�'��������
�SF*��1��3��Dw^�F���l���f_2�¢�ǿ�2�NOލ.(�ne6�m]``^���؈��Sc^�*�[�K6�zʆ��_���O0ދ���دjTM��^�8��+ 14��
��< �(��'�UMC�nOՕ�_��K���-���0�]�,�@E�f�k��l�:��I�96��Hku���h�M�ms�<��� %تm�A!��l	�E����E��0�'�E=�τ�.V���y��ƿR��*<�������=�QՏsb	�eK��c	�7/>oG!wjՂ�uGVq�B���+�7�,����Y	5�U��'֟�"���7��`�4��>p��kT��|<��\�c���G��flF��AD���6_���R� Y��1yV;=B��Б��qP^!�^Ջ��08Yl[��?,Z9.���J�7���tye4&� wO�Z���"��d�\�y���F��1r�'��p=����Ӂ)����8d"V�#��ϩ��H��`�:��Wt��x1j��,�k1�r�J���>�y.�)�E�����:���	A)/�I��|_�lT����0�8��血'JX�+b�f(�^Ǣ���Iȋ�
ܵ���
Z(�P5/N�����S��Ie�C�O���}Hi����5I�.Pue#��bfl}�G)�[DB�ڧ?_��W���_�ŎU�9��2�쌇֜.�Ԍ���&����BANw7Z���\|�+z��3�0I�G�<���r\x�Ae��;���[����4Hf�su��}�bhǾ׼/��_ڋH�5G_�#�~<���x������/�[ɟ���D��0Z�A��#�BV��%��F�t�P8vU�;ۇ��[a^����"������g���V�x��MƗ��G�{�dU7�k�O�78kr�-�bjW�&�6~
�4�ڐλ\�E���M/Z�wY���-��X>ş)F	����!S� 1#�j3�����լ�P���=����ш����vZU���J0�-,��1t��2����~S�e�ҲG�(\�6�8�������$�;c�=�����g$`y�% `hĺ�:9�[��Tc��2UT 8�fYN��� 7*;@?�}�K�8u�����1���X��ǭg����� _�`��Y�1��cG�-���I'��_sEK�+��4�s��di2#kυq���_���KB�%{c�s�������5)��y%��W6������W?��Ϻ����6s$���ϪM�s��]�8%#S�H�J��"<M*]ߦ�>WM�����/�v�G�֒�C��z����u�0IL�sn`��.�r�0�a阛��I>�@χ+O�+�Car�T���%]+ŧJ������ZaFvƭ��U����BP�����p�',���U���Fk���t�x���4\��b���g������/5
�e�zX�KܒA[���O�-�ީm�cv�֐i�5�	Z�x6�w-v��K"�a�<�#��a�,zwW%��R!.���p�P7kL�p <���7����*?�s�\`���� )�ݘ��pV2�V��k y2��C�ԙ��@D�a�1y!"x\C�s~G���y6��56�b�)I'O�ʊm�XR�����K�+ &�%�g��]�u4o'��<a�}��
Y����T��K�*��aJ����l�o�_ws0��.?ﾜ��&FɘC��������"���>&����o�%���]Q��7Y�`�c��u�Vտ�y�	'!Qs��"���>�؇�o��a�z}9��z���� 2��9�5 0�	�c�b���|��A��=�/���)����j�5�u�@A`����!���&'S�Dv��8�|�ߤ�N`�_f�NX������A�zR�c> �L��nlEo����:�k���;MGiKR��G&)�Rf�՚��8E��϶	Xo�����W��8C`�f2�R�dha�YU�3*�F�7�∢��0�zQ�˳�������-�i��`��f�ѹx�Y��V��Of���L��Ҏ8 �b��u�"��	�3)u��O8���-���	?s�#$�Y&�兵��Z0a/���2-ϲ���B(�?�aK�� ����NC�L'�y���܋��C�����x��b\��8����Č�_s=��vؠ˩�Ls�ga����X9;4�IL������NX*�#�2�!��-�r~�>Z���.�*}0kH%km�	�X��I�_��>��Tr�}����QJ�wR�k���~^��d>���sZ}�)�qm���K��G�b�C'�T������e2]Q�L��!sX��DL5�$�-��[�k�C³��$�?�����քshy����5���hv���>���i�B���Bx���{�c)���W{��󶂙_�O���m�p�u�+��zͩ: +���-�_%�]�,Z�¦s�oe6W����y��Nv/#Y�	.�, �!�ձ�y�߬sy�+��YȂ�]U�4b��5�e�vf��ߔ?�}Y<���à��7�Gf�tirO���,)Y�?K�"bO�F]K�P��/wZ��#��x��o
l�C���Y*��"H炈�	l��@J������F�B���K��v�(G��o���3Vz�Y�M�Z�G*~�<��4��]����8�~�J.�tG6p�K�xʛC^��i��<������\����`{�����ڣ�?̓��
��}�����P��
bء�(�gL|'.�3����]����e��s���u��mJ�+=o����-��a��VQm�����,�<5��<ppa��6�<�f�頨��J<��}	��4�����*6߽�X��,�v)f��������é�C;Ho���������; �9�����%?D@��T6���䥷�{�F�,̗�JN6�Df��Gв�Q�o0K���q��%�Yr����|���`�A��!�*�u
Na'�$1]���.�{����O>��=�ÏC������N}��O&Y-�(���nnGu��(N2�2��$�ڏk󠷭&�H���*��T�z��{#B搿�+N�@���V[��%/��r�z�*�Y�95AS�H�?	h�IV�,�"K��5��L���0�L�ա0g�
5�'���N\X9���tu�����:o^�mm��ϯ��߻.��xkB�~=�,S������.>��N2��q(M����$6�rS��Fq�}�aDR~@E���)у=N�X�\��W��(��Mz��lh)��>&�$=.^�%	�Dw|nH[WLͧ<F,��&^��|�R�iu��RG��ck�)�˄���A5�	�0�Q8����{�<jg������uS�AYGπ�?�������3z�٘LG��jtZ��H)¡&��������B�v�z�5�K���g���"��6,ㅞ$o_00��F��%Y(�[4"c��<^RNi�էm�l�� ^(�wc]�J;y�s}�t@q奯�z�ǆ�@֤fbesn-πy�%�Y��������+�/?z�ɪ?��~�H@een��Z�$ˀ^dYt��͈BT���%��{�e��_��x*g��Ը����'��@GkSM_�A[T�]<�V:I��d��v�A=�[/إ�n@���2=$�C��*,�RZ�d�;�k�4N-�N��u�-�}'�`��d �,
!R$z�h�;��X5����V{��/��0��R�;���_O
SC�<v]��,�(�A�I(H��c1R��(�WC^��F�t�O{m�9�=m����3f�e>��X,Z��ϘMղ��@�R�������T�~P�7�L��Q�{Y�)T��2H��k ���.��������(�u���G}�r�έ[�C��M}�J�Tb���Y�x��k���[ �;�.W�5I����<�M�7(U��G±^=���1=΄�d���/s�J}�s��k�X� ցk�{������~o��DƏ?�cD2�1i����U�)�U�|������[�'-,�/�l�g��#��20{Wu���y��L`+��:}ZW%$#�S��w�11�K�_e*�_����qJsnݹ��:)�|�Y��U�\�d$+��@(��r��L��x
IZBT�\��W"A072�\��jJDiƞ�"�A�%.D:8.�q�D���fu����j�{Z�&��q˻p�Ms&��+
�rW�&�3�Pi�Uv��P2Jq?��a����V=�I�f�R�R	O�.���js7oܽAEGW�m��}��M�S�e�w�h��zۊ'�G�/�!8�����z�������D�J�I/����]�3�[�@/��dX:޾��4�i����mr�B�D�^�8G�z^�0|�4eV���k^;�MpA���f�@�y��3���LfJ|�rw��o	yc�=��ů<vݿ�[�z���(�� +�6� �P�JiIu�d�#Ǖ^Gjg��ٻG�v6.�ܑ �O/cn�}	w 
��Y������H�p��/.j�fB�=J�c�!���U�Go�]鐶�5K���2v�t��*��N�� 1��Ǖ�C�;C�8�M`�ŭ��}qF���T%=ņ����ǐ�&�]�]�\�>�T{vҀ��A�\�� z*y����dD�o@֞����J۩m��\�B$K��⁌��$�dq)Ɉ)��c,��R�|qR�S���ޜ�@A������"�j�<����X����%��6�%��%��/��(�Wѻ�u�M��c�͸�
dp8w��W��f9�C�;�q)-��6��D�/wY�:�����/I�}8��&:B��kf��u�8pGV ��<�-�������h�o�0F5c�k��]�ܛe���vO-����8��\	�Qd�X*s�As�����=��V�L�UB7؅$����J�W'���s���I	�0p��5���kN�Ȕ!��X��}��=��j]�/<�QB� {��ô���LB$�	�G���)*U^'�U3�d��1�<R�>T˃����3�.U[���OH2��2f��Gd�_����}?���Oȁ=�b3��=hr ��rfh�0Q�v�-�,�L��b���X�"m��sl�_�~�!h�{K�~sSDvt�������mf�l������D�7$�6"�wt`�i����!ۿ��Yb\U�r�$T֣�V^��(cŁ�˓ϝ�M�:��_M��_�̻�]A�(���x'�b`ҿF�E�i�A�w�.��4%�+p�!����ޣ�/��g';M���/$��c|Sp̽D/�A:�^[��y�6��^���%av�����k�/q���}��uA(v����i��� �����!��II#bm�n�I��OE=0�DRF�(e���w��/��-�:/A��?f��*j�c�TЋ\�c����1���G�B��j�AR�,��B����Cx��2�!��X�d�)]u�&����d�8f����(�N�1��Pe�����_���U�S��h��W�]��5p�m<��d�e�0��e��Q����U���0�{�M>T0�W�ؙY��Kݑ��c�P�A�L�a��߄��r��}(�ح| A����>f{�˖��K5����HVG7v`ȵ�n�̯%��hj���J5Z�}�0iK��� &�64�'������oC��b���ؚ�cy�5wc>�I{�؇�Dݴ'J /�}�)�����1��L�J����8��x�l;�)�z������9!-�z�* ��gQU�� k<�fl�*��鹊�?�~p�_ֆJ2���wY�7�$p�r��d��y��+���Oݯ�ޕ��3��y�[�+��֔q�a���jtRK���[���^E�Y��ɼ��m�T�-i��2�@ޞW�)�AƯݧ�B]	I��o2����\���LЏ3�i���q�CԬ���T$���;w����qy��bx>,`5d�\���c@Xś�l�>{el�޺V�#tN�T����U��&D��ʄ5A�9�e��� >?b0}�1)/֔�9��fSL��Vpg#��l��� �ª�&��}�5RO�R��@t6`m�i�1
�MNx]]q�,K�$o��;e�P�y��Q>�/Ab������x}3���p�A�LO��p�/2z+�nk�̮JZ�1T�5�ü;�������O1'�S`���iki{�'�zN�VJ*I�q�	���;�mb��$G>���]d�� T�f5���=V����,��O˅`o����1h�'��aM��������ᡕ���07�8��i1�Z�J7��"���&q��x�w��DA����ӵ֍3?�Чm��ء}��[�-�Ρ�y�B�Y���-����)uP4I6�e��˼9K�{ ��:�&���w�D�K�kz��M>*��v�i�q��D%� [��$|$7��m,�L<�#����(nf��)��5�? �0ސ̌�_Dm�h�bDl��WYLi�G���U�Qe�3B��,.F>��1QdF�[r�e�����|���r�Nʹ�g��
%���ǡ�Ǚ��ϟ.����Щ�n��V����>siUTG�h}V����ج��{��&�@J���-�IPvWOu��u� q.��m~c�����2���������jݨ�u��uu�sட���T@?��<�v쭊��Vn�e����e��`Nм.৆
ʲǥ���s���U���(����z(�F��f�e)otl�#N,q��#)7v�h�`����^�B�-{�v��	�R���k)������|Wp�G' a�?`�ĆgW���aM{p�[�e���俼�a�	��tMaU/v��8pXr��(_�<��Fz�Ư��	���#��;�br��9�����g��qN�v���M��[[�������.zL`T��*/՟��K��N�9j���2x*��5t�f��i>�;���Q*����&v�h�_R7�N�/�U�{T��?\��|����d'Ux����	�ɣ�_筶lf,���,���{��$� sƳ�$ۊ��G~_�������EA�?@��r��W�[}�M|�����h}����z/["�����������~�c��i{���V��Cg^��8��vr�^�T��$XLc��MP+=�`�g���s������?�UNʙ��� �D���z��XTN�p�,�?��2M��)Q�W����@��,;�-Z�l��Ȕ���d\���c?��L�<��_i�z�U@��F�1��F��>�۾�m����h�����Qw��ܠ�Zq��&1(¿�#`z��~k�CBm�9&q�?Ya&k0P���^�{w�1��˩mվ����1j�N�����Ko�H0�6V!��CBM)�yS
�ڋ�q���D%#HY�Dh( ������ɵ����O
e�l�B���]�oQ�n#1�7�s�ClH	v˸_l����\{�*Eu��T��������C2�`�������0?�_�v�eG_�M�5���d�|�9��F$�2�����=��/�q���@���ĤD�݇���&0Zd��^4 �pk���f��O�#� C`�/m�ת��ٖ#��
Es�F���~�=t�J�i���i��!���L���Br3�L�PΖh/�+�# =�ڪ����Xyn�MElr	�}&�����v�a@�*	(���1�x��'����U=�/�FB�C����Ũ�7�fJ^bYs��S�}����� ^�F5����_A�\�1�h��j+�u�Og���r�m�)L�3�A؎�$��"��F=�XR+8�����>�/��i�K}�Pj��8�х� 5��>�ݜ�8D��������J�ɸ��P-�0wN�L��	W��eP,ȁ0�`�D�?6sn�rL65��x�o��nFXX��3i*BjJtd�t����oP�ae�r`�+�`�U�R��09#��6������)o���-� ��t����1%�Ƭ�|i�XK�P�o90�� �b�?ߗV:{G��ץ�t�C�&]c:�͍XM�n,�sΟ6P',JA]8u��%z`>v<�M�;uIs�*ßԮ�������%2�T��D�i�P���cJԇj�(f�(���RHy��HOy���S6�(��������4��؆\DP	�N<e�( EF�˻���:,� ��پ����r�ȧ������V�����i�����Rx)f��9�J0�e����.0�@Z4�W���~a��FZ,z����(�QȢ��:��uNp��ʛKV�^��qD5�0���{ߏ6T�5g0�z�^�|��������؁[il.�P��++�9�Sf��c����u�o=�����X;%ϫ�����������s��}����R 12���<��7��psQZ�̝��w���N�i�&p�<SfD��ȶ��q���%Ǟ��(��>`�K��n�B�����XffQ[_�y1�n�Nr�]Г�iq��:������Kdb�vD�)ǆvN��ͮ�]Z�<�yv{C�VG
1}�A��ה��2s񷃃[=�	��#� ɮ�#
`���v,{��E�����k��.��y($��ށȰ��]����c��!�^�i%�\%���y��.P��(W���+	U�<���d�����򝳧&�_�f��e �5! ��]y�b�	�J��_q3$�d��:��~:�:zES���5g�Fs)|	��;������E�Lg���c����y^��*�@�&
hA�"&��e� P0�M�6/�g�&�d�wb����J6��P^c7jZ�*������iw!����@q˥y"1�]��>�a��c
���
���t[a�mB�y�\!.q�j��5�o1h��:�B�O��S�͵r���3"��B��{}��m�$�;�3L��a*�a��}�Pwk"�U�i�q�g�����j��;������6.�U����t[�Fcq�*����F�j"φ��f�"X5�S�R6�mKg��u"�.���W�Nh�\���=i�U�F�\ޏy�� �\*�Ec��B�H��ݷy5(����ڝd�гI�8`��D�h%ܥs���k��륯ǅ�zO_el��J-�5eY����m�^���/��}��v�붶V�6���Q�ﰟ��&8��F#�O03a���.�3��bߛ�����ק��[���.����e�t8�s�bcO�)�(���0�[���ќ���vR�p��z3c��[集�w'���y��V�[c����K���ʐ.��&<�L, �v~��P��(�ίע��"+<s�-���K��HC��޳g��ߋ̜�g�<C@�h��#���-�NC�X���5U�R{b�s�]<xYS�n�� 7��鴮4_���4�p�e,h��Z)�\�#�/p��p�6�Ώ�mplC�7J�pI�O4����Mq�N�I��-Bm�?�2�B�U�f�"(Ѿ()��Z",#����7���-P~S����@d�����5���zAd\h.տ�>K��˿�?��F�j_4�.X�$�6�b��4�P��ͅ�)Ͳ�><�3=iP��g��/�ߩ1%�փ-X�"A�1S?̻87X�[�+t�p;��Ra�0�@b��N��n��J�A�cI��0��+'@y��8�ў�^�)�ɉW�'"3"�r����ߍ�Bl0�ȴ|.��ȝ��(����z&a(S�{o��)����0cs�l�v�����%X������|�ʴ@t�!��p��9h��$��,gB�<���!���O! ��`��)�@����^<�{}jmO�0Z ˹�շ���.Z��ދ���vL�[N�}�Pb��
]�ޔ�ղ1�E[63��J6��չ��݇��w����kv�r�)z����{�k�|dʀKM�_c�#$/�*��ֆ�}�Ѐk����G�Lأ�2�z��id6\c:!�{B�Kw��_��,sy�`O
�x�
-%"�r����V�~^a�m*P���|��E��U���E��-����#(��*�JdC�:>�����:��+�.�*X�a����2�͈��KnԎ�4�3{���̛�H�*�s����鳁�I^�ǫ���E���'2�v�愓6��r�#A
�_��|?C
�F�E��\��Bgx�:E��H�g�*0���8B�sL���r��7B���L�����"�m,�%��1T mE�t��A�u񩷴bR@��R�4��7�Gzu���y�(��BhNN ?F��dʮq���X�eQ��݈�W���/�X7�����L��F��w�"vS����fi����Y�:�}�T="^
�_��o��3��������W_G{sO���j�N��X��G�lh2]/�)�A F��%y�2��}O�d����Kf�Y|��ps`� w�O:Ȁ� �Ѫ�Ȳ*u�e� ���-��"fV0F,�����y�6�־�
��r٤�r��#��x��L�E�?n�ۚ���0n!��7��y���{��pG�Jfr�F-��=3�דV[��#>.A���Ul��ѝ���^�����l�*0<��F�h����֚i%~�aQ1�,�e!��J�#�I�AO�L�t���#p	^��<G�h��#9�}�2��I��=�����W���%�^f�Ov�ϙ���z @�.�̥g�>i6��T������՜/B�PP�A��)��㩯·��10\,P��v$=��0����w0��	�Y��D��Qy컑pA+���Lu�o��=��F+�oI���2�,�YX�D0~ۂ+���쟼��h���
���Y�F��F"8_�<y3�>Pf�M'�}"���dz_�4���l�g�������7����?��HB¢�	r.<bd�9��a�E�ѯc���ST2t�?��(��T6@�v�j�9g�gp�m:ĝ`�{	}UԪ|©� �W�ۣ6�A0T.�V3k�W�Fk'���3��aH5gy�j�]v>Χ:OW��xR�9���El���h��{q�1`��I��&h�E~�j����~�N%q�H*z1�dS��tP2����ҍ�D���Z���ڼvD�ʬ�^�Y�P�� ��|���ů	�6�|��,ps���m�xrR7���ڴq:dN���x�>����5���	�q��U�qۄ�&��+�"�ƾ[�!�k���ܦ���g�Xz(��2fFi<גϑG^>�u�\�f|gG�w��Ću��T����Qh�<�nFG"&��}�m�[6���_}o�An?����	�윍l�0]Ed�{�#bYXr�������?R��ǰ��_�&&��q�*�($:�i��*d�ՑOK���on����x(%A(�b��$d�d���FĞ�XF�1q"��K?h�ϝ\$51t7�\�^D��m{sw��Y�M!���)��L�׋�rō��$��A�'��\Wj��6����+Ɔt����� \�m2�O�����ߟ�M�|�����^J��@*j����r�'�i(�nWt��Jܰk�{ܴ�Ɲ|�U���u"�Ivd��N�ᡑ �d����p4��D:?{�0�M;o �3�L�!��u*�3��ӡ��GN��'�B��{�ܜ�A� k2Bf�����.��2lH�z��+�
k䨎ߌX�t�]���Ԃ�"ި~��6��+�}Ϟ�;��9��=�"1�j���x
ڲ��:�=���[�9��z3���,��o�v���H�@5m�*갈b����#rj�igA���$ܔq��_�è)�-���O�������2�B��Y6p�0;Jl�k}t��T��S@����{|���3�a�wQ����*Q��Ɣ�s)�[&	-�N4���:���I�y�q-�0�*�h�W�GY
�+�OO��%7��j&�o�?ÞDRʟ�FY�{��oªD�Fn��B���ߎ��W��~�03Ȝ��[�9f���Y�bܦ�v�Lk�t�AA���#�8�5��-A�ws5G��l
R�����t0aJ.)[�1f�\�E�����\�w�rY�^�@��T�ȎBk�~{^K�AS?����BA6ֻa��=�fǋ>X;��u�#a�a�B*B��{��2-��m���󿽙-�u.�M�+��H"G;�����H�EWA�o<�_/�j6�D8��=�U5�1����/^u��x�ף�B��0�������Mi�w�E}�30�� ��4>_ej��Z	6�X0�����*y�S����5��E4���3���Mf� i<j�f��ٵN����F	���Y���6N�<[D��j`o��-��z���6�0���X�z6�Υ�n�0?��ܛm�,�|(�l0tqf!P^��Px2����̅�M�//a�|��B�eK���ͻ��y�i���qZ�Vc�f����0qH�CT����tH{�lJ�K��]�#��/��+���*�,�߬��:��<���i�GaZ{!h����u�!f,��\���Z�����jȓ���w=1���'1��>[J��
����%p#��|�,`̆FH�&A`n4�授�y�;7bND� ��Լ:���8�+�?9�:T1��Q��iQ�,dar]>>w/���"��+����*����(r��*��k��z�W[k//����7���˛���ei�1m�2Ɩ��*~�K湸���R8�d�*"F��[` E�>���i��I!u����iC���w36����Ә<%���}]�i�T�(%��%�Dp�N�P櫕/�ٱ���R-Z�%�%���Ǵn��묽��j7��򠧦R�q��!��J����Gñ�/�0�7\jl��%�	>���Y�C�8�S �}��9٨��gHW���5�0�pa��l�R'ֲ9�Sr���������P҉L�4ქrUi
� 0�DÌ���7{C��Á��K�2�a����h>a-�Z;qԈ�45V�L^l���t>�t85�*)ɒ��xShc״�rz��e�<�禃���vݾ�Cf �a�������������@��$�V��O�fk�k�3���j�]b�؁0����wL��/�0�/A��jfl
�e��.@+p�\����&�o�^���Øyk�� @]�B��@.D->$zQ=�r+c��t8�o��>�S����KO�����q��� �� 6<}"�.�C3Zⲓz��E�:�a�w�^c�} �O��DVm�qD{�8��N�{�E���8w\e��"��mR�1���^��Y�݀��"A���FkRX��"\u�j� �T2���'jB	���հ��%e(b~G%��1���>��M�G�PpS]�A�ụ�Օ~�CX��W���ǘ �D�pW�/(r~�W�Sagt��%�6]�n.��g�X�n�B�p��I�1X�S|�1&�hC8~`{��#د���k�S�a52QP�w~ m�~�=Z��Z�3����٦���\"$�+	j��hV���Anc��lZ%��Ly�ܔ�{Y�w��|�H�H
^x�>({ď/۩: ���K��к}y�Gb�.���l����qgՙ��g���'��&װ#�d�Lm�M��V�D�
��bѸlL�d)�`S��s�֗Q;KZ���(�Þ�~�P$�r���Q�m#E�z�6�.pF����C}�P�V�s/��].��ΗҾl8���"2�8�����7cv�p��0I�vv����`(�K[���TG�H���fC�1�w�d���.����\{�T蘃<H���?[�����z4�-��L�7�L���&ڡy�J��y̮j�J/&���D!\�.�<L{h%�c�C�p���j[�9a���bw����27��������=��Q]�-6	��e�YO1�]��u����z�4�V@��0 �d1"�2]>[^��5-�c~W#?�bD������v�'g$�+�v^غ�����;wͮp���Cз~�X���P]��mԃq��&>��H{�]_oY]���[�k\�QکULd��S�jI�|(WRS$��ʢg�v�?�<�����{c6^����>��X�4�>�}�2��n�/�81s�Wm�3�ؙ��@�����,���5���d�`Q�-�"i�]p~^<��++�I��!	�t��Sg�a�2�o~��8ަ����W�m��m��������>��f]_Q�a&^�&��}����h����i��;���*%��10�,]*��)�?��!�-;c7��5s�����5z<p�������j��?&F�L�IԈ��f�Z�.�����i;� I���N�N,s����TB���:�+�e�oI��A2O�&dE�(�"d)pD#G�'����cԁb��R6ԩ���(D(�o��&E�Pd0L��
�%t��k��ʋ���L�Yc+�	�YL�eYi�.Nj���A�F@n�&[I���Fk�ljWzg���j�s"����\����]����9��czPy����=��]sHh?����l��E_2������z�#�q�Cƙ��pܣ8MfNm���T�#�e8;��?g�}f�Hs�|+�Mn�IU���{���#���{y`�؏-8�T �nK��`&oi��!�<���%�(�<��u~�C��ӹZ�5�K#�5K=Į�~}���A�I��	"��������������y=��b$�+�Z�(m�}g�MB�	�e5bU�,�)ͭ��'�:e��2e�|1>�Ϛ�e�"� !߿�O����X�<��Ѿڒ�7ptN�AGH�v��8=���"�d��g�����,�e�ᔚ�ĞYL�y���?k��w��{?�`�n�M���P}0��Z@�ݠ���ٻ����k����m����5K��:ݘ$��A�1���m���ps�b.���tͯ����=�(m˥HT�y��]�����X��}����}����������+P�˽�9�a�.J}��F��&-��K&{�o1�P'2Hl2<��G�����'��`w�ʚ�=��7�'& ��@���^�+�8a���\-{��_�F陱��-V���{$�o�}�b�3�
t�e`ez�g�Aˈc��|�����!;�ri��#�X��4Wiݕ:k7x����~u�����"K7�{2�����f[��f��j�ξ;�٬�=e�Ɖ.��w:&��,���-�;��#�Ҷ��?qA�Xq�,<a���x����� f`��R&oj�`9�	��u��|�/lf`�z|T y6

d� ��Z�Ml��J���肍����io��/����E�cKm!�QN�@����t{tƭ��f�!!�HI��Gh�(F�����b:0Wb�'�[���uF�@�e^G���ɠ<�����¡���Q���֛��ѡwfpG.f��7���B��â��/t���%��!���Ww��e<�F�ׄ�x�I9�~��4m��.����j��|ct���McR����e�L�`���Z{f�"K�kH��v6��ݺU{�I��С �Y�z����7@l���?8\�/�I�h1&����8�.�,�==�4*����D��H�9\�.���.:'�����
l{d�r@{�������p�<�O�Ed}��)J7�FE�`V�bHXwF�Ж�c>�B��-@�W����u�/!����Νő�B��� IV�)~l���E�����:�a<mJ��Z��)>'}�����g�D �w5��Ny���-
㐍��}��h���LN	X߂5y~g+ՠd��J&ȑ��[��0��-�O����]V����p�u������u�ӧ^���N�2�0.@������Q��KND�=���8��$* ��~%N��ە�Vb� Z�SƱ�lxh���y�=�1���,��rV�j�CѾѯ�رdu��$����FC�#bn4�Qr(92�8�����&A�>�F_���~%�^�W��Vm����v��Gvg��,�bY���\��l��-��� s�U��2�x�i_i��p_��H����N�K������X����E��`s��"ה�g����!�g�e[iD�}��Ǳ,	c�x��8+	�aW~i��'����"�>Q�������y	pS�[q�� �(�Z0��~i��~��?��)7ˎp#7`�:��G�5��	4�}���S�0�2�aa�n1Z��g O̵}#DA�Gt��1���5�%�UN��ͣ8^��Y�0�V�-��L'%z{���J��
�?�6lfiȊKߟ�C'����}�Vg��R�]��w��}�-�a<o�4?ω��?\��R�NH7����+��u.��_\ۿ�	��mIzF� ��ǿ-���;�K*P���c�U7�`���E�[^Q눻d >Ra�^:Vuqu"�69i(���~e�W�x�Z`�L��@�T(��CgoL�0v�n�߅��;oj��K����}�� �U�����,�mڪ�7�ur������K��B�=�g0�[Z�lĄ�.�/O���GV�e����0��9�9m$"(	�= �Z�d���@<�l��1�B�\V:�mM�"��H�j�O�@�a�/��c�vQ'�M�d$H�+ie�"7{�eo���_�B�i���Q�]�-��Y�r1�u2S�;L�>WЊ�'�l?9'�5W��8n3��P>[z� ��0��Op�"��R�#��2whɲ*�(�˒`�2jY��w���tW;*2�I���j�Ꮧ�7B(9��!<��I��E`�1R>�/�@9:�{�.N�z|��������* @�G�zd�+g���V��z�X��+P���"v�����<Q��_<>R��m������h�L�SE/���ϙ��Q�S���_y�th���2 ���w�y;�泃@msqs\&����.���\z&�M����Wʙ%È�*�t5#��_����U�ݽ�RRX��#wWT�>��NK�YN���Ͷu���kko!cZ���� ��S��QR�q%_F�L���zu
XsqCh���̍��6@p���3��^���U����:��*3�݌D�����T�yވ�3��0/3k���k`�u�����TFoh�=�0؍���f�9D�͉4��sf�_i$���f؜���JB�ɷzC\F;�F+a��*���K4�i�?�BJ�
��:�JuA��������i�$�x"�%r������4*�Q�h����������{�S�Ů��:�<_N|T���k�%4G�ʠ[��癷-�6���pw
6��#/B`[r�����Z����y�a��;�� p�U��uWq%�X��cT407���V�M\�˒9�+�Ȓk
���l7����{���|��b�}�FSPT��?W۠���%T���dr��U��]�*��+��)Y���fٺ�%C6j����/7,�:�1!y'r2`I��cĝ:��- T\&�=�(�� �/�,$�)v�zo���Ϫ ����甑ި����a��9S��pv	�[� �w���7��H(���\�^��J�`n}��D1b��TWn�N�, �j2Tƞ�p.e�5��i�nrX���p>��i='W�b��zhw� P�|&t�YF����k�@���(�\�d���>���,ʓ��R�Z+���d#ff��oc���bI"��'r��j)�ə�Ws��5�,0�dZ႙���a�� ���~�>��8���R���V�
�Z6&�q��DWG��N?����)ٱ��������[k!x�(���;2QY��n4�Z�5�� �G^���&;���e?�>>Arך9 �x�:7�ut@��ng�c�������zVu��v���m[�~�ִ��G���7W�n���`s�4(S|;�������q������`��c��{���N�*���}��w�;j��zH��-n��_�J��e�.F���r����R:7�� %,4j.A�A�����F�P�n�H�d�'  .��`���~�_QH���3~�v��힦w�0�x�����}|��@e�x�3��j,1�s����<�C�?��X>��=�>�m�/�%���(�޽!���Ö��KFi�0�+)�V��O��I��M�����_vIeq���wd��b��*뾨K�[��0U�FS%��\�B�6&S"y^ڨ1��CV{�F���qd�$Ȱ�&�E�!�@Y�ё�,�ԙ ۗ81��2Wb�cx,�>d
'�>�uܙl�hv�H�B���p�AK�*2�4�#�;����������i���" ��0��S�4+kH����L��,���_�PF�fښB��Y�Iw֪}��A���[�vF �
����+��+4�r,�-�segɉ��	'�$f7-V0��ph$����(dK>L�g�iM��fkp:^�[<y`t^��"���}?u`�k�pRYh�7��"�b�S�x70;t$2i!Z�?�@\�2'�1�ĴB^DR���Q��n+<�[#�����9Z@���B�����;�_�T��d���ގ�՚Q�j���V|+B��ppͤ��K�O����^��n�ʂ'Nې���5S��$��"��9���A�C�0�2��j!��j%^ӯ�Z�,�fB��9�u��0{p����,�9��K,Ŏu���������T�n4���5Ej�O���v��^)1�$� ��k���~�꘤-+!�q��;O8m�#�-�(�.b�]b�v{N��d�`�"�v�8(C�L$����pO�-{����f������@�G��Zz��ו������Z���a����	#��
=�_�p�"��U�����w�۳0��q@Kȏ�
�&�y�R�cR�������|RKؿ�~�3�[T�纭1�ς��K7�x2�uA���gvķ��o�7Im�%�޳��£���*�(j�Tx��6��Oa�{���@��}��oA�~�>����y=�������,Ts��g1��C0U��Q�A����������a�A��p�{��g�=�t�A߃8�[֪�&���0{�U���|��ؗ�������V��w7u�n5&O��0��L��~���I���[���d]��e
����2�K#��2]$aT1���D��T�<�� �-fw��aLP��������G<��#�'�A��ߋ���'�X��Z��s�W�y����|��"���Q�q٘�P&�8�E⡾��%���j	�ㅑ�g��6��z�|D�C�o貪�+�a#\h��v$�)��×��Y��,-d�.c0���sq�貑c�H(�����_��F��^��#i���RZr8�b*�sA
�]�ؽF��X�2�z��K�Cd����n�Ѱd��C�۪��"#/��cxh�@�/ ���S�fкM�J�}�,�"p'�I�
t�.�dI���P^���Ȁ��vG����w���&����69�蚓�g;BvIW� �M��6���.�i���3��jl���W��%KM_1r�o�O�����I��}�N�E#�t(�+W�X���BI��ɲu�K��A�\c��Upʪ&����}���F ��ga>��kor���hqm��|~9 ˍU���O��r�u��U�twǆwuj�(����a��Ѹ���cE6w�<KF�܋O���s�:Ӓ�ǲ�&��YН�g�Դ��Q�z�IWJ�KS8M\f)J��}EB)IZ�����;
�ۡ#_RTz�^SJj*{f�ŢZ[���ER?.��]K¸�ŇK�U�^%�r���g/���*��X��C����ǧk勊Ƣ^mhQ�	�G�uhE"���jLV����w�� �צ�a��z��!Z�� �h�n{�xpȬ�en5)K��Y�,pUE%����1���i��tL=���5^BboN;���5%%�1������׉�(g�t|���[2�V����4�8����kB&�LwJfC�hE�!|�m�,����|��eUDXD��깝-�����v-���8���ܻ]!*@h�4�Z��6���"/�ʶހ�C�ѷ����<-���~S���JC�t�����다����3�A%�Er"��+��1r�g9�&C�(��`ygvG6N�{�9�8���@�;ư]K�ʥiz����.
�?���a�y�	�m��B� ��&�w�/,|5��lX�t�h濽@`�$7�L��,w8��s	��N�D��y0ο|�j[�i��F0)���q@�.������ɋ^��Ť���.WS|2��?��e-�D߻ �cE�,�L�_��ք�x~�No�T�_5D$Ѕ��'�����+�T],3��~����QZˡ�V���C$mQ�q��7k8#�
�$�-�㦫>6�b���nܘ�[��2H@��U�z[�R��m�ӂ�9���2<�����o��l �����A������޹7��=aw�T=�[�3)�^��5�{�j�BJ���F��j��ƻ�n����L����\�ӫ��D"7��U�§<�ֿK��Pn��b��h!��R�S"��L���c�;Bq�ލN;\�H[?j�O��t�[P�N���1�҃�q2
9�}���[1[ �8�?_9�^v%!�*���`���]�_d�	/{�3�`���(� 0��/�_q ���2}{l�1��d�pX?�5����ɝ})�G?N�t{$��5�� �,l��ы���'����O����@�����ѓݪ��~u���b�mz��c[g��9����ߧFr�(ǧ� t�f�P���%F�Y�8kz���ߏF�R���7/p�g _�Y�����ϰ���j��P�0�M��^�5�D�Ȕ��=�\c�f�%�ނ[w���f|�aIo�Pӽ�w�4��Ω��2��#���w;�/~)]q:Ā��M��������i$�M�QEQU�Ϝx�Hn�;7~8�{JH�s5���E�4\p�v�F.O�����o���O�aʦz���L�'�R��6�~�O�1__�<�0�oVA`��41�3��4�࢘ܜ�7|��?E�V'j2�e��i�A
�n@O����C�)��57��|��`��/n����;���U�z�d��o�*(�}���[�Z����($��J���TI*
p�Z0g�~Hu�fl8K��d���ͪN]*|ǦS������(�K���g��j,��߀J呟��h��=b��m����i尿�X���WR~�ע(J�(�i �A '��� "��`49�|�(W����^�֮�Тgj�����"Vm},]�+d�5?�a6N�8j8=�o��DFx�!������t�޻8�����D�L&��wsV�L��b��^�J�~Cl?v{��"�]�ɑ�_��93�#v!5h06Ţ!�6���%I��L����z�y�SX�xE�v
i髱H���G�8�fFF��l<&4���{ʇ�L����L�S���c�E>j��Ɋ$�
Q�I��Ncl.��P��=X�!�p�����Ŏ_�S>��M,����B�F���v�0E�*�"�Θ�O�`Ը2��.	��i�Nc��.w��by+����4��g�#*����*(h�_q��z�2sF�� +�� �.Ķ`�4�6!ک� �7�z�'U$!��n[-L����?P
#H7Ezw�xs�Rps{��
4Yi��.J�o�se�|l�:���Z����Z#�X��`c�Uv��7�5�Lp�nnA�.г�M3uw���#낃��
��l
f"��R� �N�#�bQ�OG_�-�Gޒ��k�a��H��6�I☫,�u�I��t�m�3�9
�{Eh,�D։7�S���L���;��<C%�`nmQw�p�Whɻ.ةw��%~�U��yҎ9��&i�R
)o�5���1���}��9���\G�3�k�sHP-d?՟���ߣnwÌ��u�������-���[��^#��ث=z�Wֲ�l a��� �!��N��F)56��-ʆ9�Z���a.#o8e[Y��������d������@�Vo@���Ʒ�� }BR�3��ʏ.̿ve�R��[H��jD�ZK�&�xF�m<%o^.�1�AǗ�@���}�	k@$�m��h�X�Tg��\�����3Z�#ï_UfJ���Z�+��01wq�����V�V"�,/�P�$�*	b�ݖ2o��J҇�G �R`��/o��A�j幹��r�0��OW����.�󨅌N?��0�cƵD|�1n�'TS����7(3�����B�	�?SLqͬ"|݌�D�v�S���v����2�u�Z��KGK�CV3n����L_����Z�qq�WQ. ��o"&�f]��%�4�xG%.�%|��E�����)?���J;̱����O�������v!�;���/�$�����(9�H󛉱PX �СHB�����X�O���*���GaI�[)W�zp��(؉�΢< 5��.��'�H}�H� $
03�;,��NV�!�ٞ7TE��>kj�hܬ�%��@��{免c*nI�H�8��xk�৾[O������,�wz_/���&ҿ�Eq.��?�Qc�	f�м� e6��bĮ�l�w�J������?�H����B\��􋚇Hl�P��U�r�.���f�7ȿ�)H��}�A�ƲI1��$�#�@߉�ˈ;ĩ�WJ�MW��`��8�c($y+�+ҳrJըKݔ�e�1�e�qD��U��<�ǱZZyI��%��k0$�O�����+Yn���N�@Y����JS�OAk�Q��+8��\b���D/����p��S+�c�c7f%�	�f�c�r��c���"v���i2o&I?�����Q"π����
�������ژ�2�:	�k4'J�ȃs>��oa����&6%_��:HR`�K�v ������\U����|mL5�w4�y �$�vLn�:99kk����O�23�C������h�|E�t]"߀A�� 7,�w_I�Y�u5��pѴ�1��jd���gI�e9X��׼\ЧV{��ɘ�B��8���Fތ�7K}[��Y��LUC���� ����.,.�5�x[��d��V�ﱨ3v��UM����4���U������m-t�TO��w�J�$Zh_�E���X�Ґ�U��/v�}�N��}n��d��p�E�@2�^<H���� ����AsK��l*���|&���ox��w�g�[;��*��<���QNL�tN�З�eL��mV�����c���_���Ԭ^F���i����AeE�i�6�2f7s#�WF=��c)td�V�`���üv�0�˗N\�"�f��ZQ�T�8���߆hXE�~Jr�sGuI��?��{,8���^�Ώ��YV3HO�^���׭c?�%1�m���1�drD���ow�X���/��Iclfc�3@�'�G�����v*���PV��<T�����KC"��_��id(,�kG�c����5 S3D+�1���1~�21�Ʊ�H32x�Y��
�h4����NN5����ὄl^�u@��s$�^�+���cG�w��av���E��j�T�x�����@�t��W{򐉺���f�gd!�NT�89�H4����z��K�X-�~s'T�N?=���d�l� s[�UB��������m��?���Kؽ]��!�c接&P�Ƚ/��5�L��4��M6n�_�W��2!f���]���{�����D��S�oA��nV�Ï�=�x�?�0V����|p�Ri�(DS�#�M��LW��C&qM���=����Yʠ2� e7��'�!����ln�΢g�vD�Y����$�e]�ҋ\m`�M�x�Y>x.��9C:9Ǚ��g$�(r-h����^;�rk���h�s�A�8|rƭo�
.{_�n �dŀ<�C�]���J��S[�d��<�rũ�hd����q���1��i���P�B�n�D��Noa]���P��P�XU����|��P��	�4rc[��٘A���L��k�rLM���w��W�k��_��
�^�z/��/�aY�"6�D9$f�:a�J�F^��U��m�f4Ei�"���w�U:1|��c.�p�h�l)��lmi���[tY���6�FU��6�� �������{H0TZ��w)��S�$Ew��R�cn��m='a�-2�G�ԍ�o��Y�����UՓ��\���1��y��2���P��">��ń#d����֡P���y�lڨY&ձ���Q��+T(t�J��l`5�f�Hi��!/����F9|אM�P|����U�b!ȧCɢ٧4����9UO���
�� W�~���`�7�����n�6�_=����%	,����r�wC����NG������ u�gݝ�����0���qn�����}�y��Aw�Z��ÖB)8��T��ge�7������� �'���"~���+�^=�-��$������Σ���2)�_���KE�6���)g�5��#=c>e�[�yi.�}�೹c��q�V�B7�!�%��#h�D��.2O�"�����S#\��y+an��Jk���J���y}\J��L�r�^�^0S�t��P*�!�!du,�.~ؤ���p7~�or���L�ۉL�M���d��2����
m*y��A[��Z�q�|�b٬�v�I]ŝ�^�@�zI'yY�a첀6�aŒ�}������t�6���UIB�����bΈ5�k�R�K I#�Vb��#.�]?�!�\����m���z9����*���kZ���)����b�#�WL�x��� jX�t�]2��Gd�^5o��۩HB�=%u����0��5�)"pz��JmL�!����*�UeON�F�7傿�F�O1�b�\e��UJR\�5ǆ@n���tTgZ ��p1K:ِu��Wo�ɻ�?r�/�sD�%_�� 	�寿:���L=3���,V�2rmP�����e ߚ�1�:���c=N��g�/	���~�pnð�/����a���Z�(A��CSd��Rğ�~n'zT��o���s�ִ�ui_@ēU���M�ߡx>S鶌��KW��J!g�l�[X��F�k�����N�ܽ��;��ZIej�@���_a
�ҫ�>�Ou�.���b#{�����o�W$2��뼹���NRUox����f��O���7�W��62��2�¾/��mQ�KǍ�!&|���"�����[+�R�f�$߈Ԇ�	�1�/u��8T���1J��n�)�SpLj���7����pO�	�>��T�p��ŕ%���wG�Ȟ���$�t��zd�)���9���_p.,��Қ:i�t����z\*ҏnP��O������A��cf�L2Y�:��m����%�?��g%�ɥ]>�}�{7�Y>����ۀk=1Շ�\��UC��s�F��W*.J�@ $D�{lM�%w��,�!e��u�!��~[G�h)m�vE�(��ӏW�����l����p��4�Y��7:�&o0v�%+�|� �CI�����G�0�go��E�c$9�!�s�6Yf'J᏷Q�ֈ�cn/L�/Jq��6�hp���Q��G��2��,M��m׾�iA����Cm:Z��B���C)����K9�-#k��"��-M&��ܖ�������K�$?� c�t!w���ށcM 7�!��k���_�1B"@mGK�lVs������Zw���~�����S٠�fMuXǺ��̗���l�ŃِۥG܌�}٪A�=^(��D-��K���=?g3�'1��3G�j��%�r2X\����O�����f�������	|
���Oc@`[��3��9=�B]u����E�0��YL�e�3��cTN��r'^�H	hE�˙�T}͢��V4ǋ��A:'ђ���h�#qSU 	������ڛSHjS�+�5��<`�o�GQrU�.fˢz���+ka��F��Hp�2J5�)��q��S�E�ҧ|�\���I������+n@�邷�za_V÷���w������+���ߑ�Bh�<�7��������.9j��_�z}}���I���#���כ���{�
8��u��=�r��K���ftX����'����:���ET�B�	^ʲ�0D%5�{��趢CθRdz��K��T���e{�[�1�\\�_�6Ҥ��b瀶S����2>������Xq��n��\�~��I@m�Lh�^�V؏�w���GկG��O�� ���t�����i�Ť}~�q�O��P;#�Հ�#���J�+��+l��CVڅ�U���^
`a���u�U^��4�j���|F�{)�n�?5+�Zs��d��QNc�g�NȪ���v���O�),Rxs��7�0��음����0��q�#	|s�砶\>�ˌ�п���u� H�-49�t�#/Od�ŉ:��A�9k!�y��nqv9���˳��-c��2G!�Ǩ+wk��Rh��ڨ�A�=+���a#����-�%��{e˸�A1�XH�Jo %��!�Hť'�on�E��,AU�D�u[`bS�ȸ����}E����˲G*5De����F�H��e���O4���&�OflG���o��j�j�;= ����JQ˥td�`�ʇK�#x�2bM�?w:)��v'2�*�>\A��NF�G����#����j��7)��`�o�@t
�̯ O�-����5��1P��L�W��x���ۃ����0m�b����H|��on{II�(�-���0�8�k�h�>-�� �i��r��eī��hX��З�ǤF�!ż�cH�Isy�f�gQxd_��SNō��L��6r2�嶁�N��:�C9�U�M�=aa�z٧Hfc��F�y�<Cg�$�<U��"W�MS��s������.;e�O>V�J�ZR�C-�Lt�sP\��T;�׷_��4� ?�\sy|�3���Ts"�J?��kN��$C�����?8���X'��#�uԖY|ۿ�/�CW��:J |�J�(g���$6��̯)��g�Zv�;d:r{��ɡ=�[b�s����xo2K���'��iz�.�j�y�E�(��]\u��\��H���B|�DHA�ڼ���G�����d�<0hMݭ Q����"���R|���l�+9�\*�#R��Ő �2�N'gr���(>�L|>����ת�i�p�s�Hh.IeF��^�x>��*��$�߂��S#.��:|3Y���.�!��9���:���nY�yWw��\+I�nEO_��I���vj7�G�YCUt���9�uZ}���P��f����J#����	��N&HЦ5K���y�!x�OE�XY�E�������r���Z�}Փ`S��,�1�o��g:�q�ڪC�HCH~8-:���O�Ӟ�8?qW;X���_�*>J�������2`��aY_��x�)3V��e���DbQ] �O�	��`���9\,����(���z��*5�RF�&��6!3�c�Y�b�u�F�u�����oǗ��z]'���+�\c��H�d��<[��N�9V_<�a�� Y�����Jb����J9@��C��WRCBs�7�d��@�Y�����w���gX��#E���\w��r>��y\�t݀s*=���,����~BC�dx���}E�Bz]\�'�c��n3IeQY�lw�c]6��wT�y���F6b��������V8O�ak׼���	��0�$B
^%`\�8��y�@s)�#�Յ�N)QOr�n\�N��U��Z@zQU��n?����<���z �TI�I�҂���r;��z�0�����l�>���q��L����wH�e���/��%}��^���L�+IM��ίΤ���}���HA���Ӫ��������V��f~ԃ�<'��#/�6C��� e���[�oG��|ä�+�4Z"�yz�K�����L��e�f��)��eV�7O�v��fY�V���fܘ��ܺ�~b�8�S��g�L�������3(��8ݴ����<Ƙ!��&����,�9�y���M�Z>�h�}�
J�$�-���Z$2�U4�k������ �Oa������a-�㱦��J��Rq���̞,ߣ�u����]�Q���J��%ɪ����]<�hV�� �䂦]r�5p�n%d���!�e��	���ٟu�a>a"�ײ��y���mj+gX���Z(RP��1�<+����~��2���iX�tGCrS �4�?�����Cl��zH�q�qt������`�>e!ֆ)VS��g����pm�{��pۄ��B�I.��k7KB��Z���N�|�-�����U�/I!>4~���7`�$v����qx� #��h�U����z� �z]Q��yrk]�8�[�F��H4q )2V��K��&�!�<=i�m��Эet2���û�?��Dl�W�^�"��=���.a#\�4W�b�=A�l����cr(�+�F����d�ݨE�%�]Q�-
R�~4[x�O_�r<��5?Ǭ�r��kq��Q�$O�fZN�M@M�`�A���7��P�#q
z7j	AF����	M(?�[��£�y����T=7悼��&<�M�tp�h<`{ j�j�P�Hd	��vl�к7J�N�����pp���t�P�x�b ��]9��>i��Wd�y��3/�?Ic����ZV�h���NP�&(�f^{}�9�i�iv�Gt3hL;��O罂tG��Z�*��H����v)�v��!$c0�k�ԁ��2 �Rؾ�R�
㉞��c_�=�'�5�|�s/�0` v$!�8���ao�H����|�-DB}Iv�ĩ�k�j����8����8/�E!�pƨrWy/y��N�F�x7����q�$��oWe�c.P�ζ�Y�9u�>G�!��:����z�!��ʂ�DEd��E��D��G1q�[G��B}q�}�ɕ��BQ4�TrD�"҂�Q"3t�a�煓�U���o'�x9W��[��� 5�M>D+J�NL�-g���\�p/����f��u&����xD`څ+�"��;��'�y�>��#���℻������*{	����l۱����5������jLq»r?���?O��-�����j�\m�X6
?��A�X�,rM�P���M�k�������_�o��{bh�6�,���[��|�L~�7��L�����[u��'����Y�>�hr�>�n��zձL׸�f��/ۍ���=�F��0����R)���:_׺�vbGK��`d5YJ-E9�4�
3�8��0>�S#��p�#ˮ�>1kE!�ѥy�ئ�>L�z�QO�i9X����y7����3�/C��|n�+7�>��k�.K��UArՐ걏'�)����Ym���j���_UH *�O[�(c~ikc������4�{��v;e�� >�&����ȵ�7#���,��{#����5�W�
׍�S��z"
 D�t������ǡU\�3�V��M��8�����|
K8��b�ޓ �n+�_�W�-��O2s�U�5�nPZ˦�j���G������\z�[�y�5�����i�+��:�uF�v�-5�su�O�����C�<4���`���M�q�[�H����%�#8�<Y��tt�S�eC�����у{�թgɡ\V�4O#)��e�q]Y��mZ��q�����h	6��g �ԯ)vw(�����:0�-��J�n�e�t/B�y%���5�|�Vf���JA����{��5�і]=t�!#�`�$�G�j�CN���Aru�e���R�����R�#=�X�|q����Ҟ*��]$�*�k���$ƙ��GR�L0B�r���C���y-t!�%*��h�[�����ȗ@NQ
J�k����K+%��Ƃ�?\���K�r��b�=���'��g��w���aP�u�8��y6l��".'8LB�}�V��֙���ɣG9#��r(J4g����"��!(z���[��q��[���Ⱥ���2��M�;Bt�(C$o��i��9_��hO�H�MK��Fy&�&���fU���&�^e}YʤS�>=�0CO��#��X����F��m�H���9B	D �L�F@.��!#���^�R�߂�#����E��P�Rŭ�2E�kB��:��iMFU�� Db��W�V1�p~v��x=��Bi�Ν��[8'7�"�r5D|H#��A��Ǯ<�D\A�X��7[*��]���w����]`��I�o���S $����5��>[�F���6i�C����w��Y�"p����^� ���B8��0��K9���}����LtP��cў�Ө;N������o5Kt��O^��?�4а��v�F��(��PX:��'E㌳��D�m9�Ǟ�i�r!-��~1z^p�T�p��[�+J	=�dT!�q�j�cD���%��[�7u��p*�h�tM��
�h�yRLլ*U!����{�՘SPV$��0�G|�2�kB4O�F��0%�߲|a������E��*�V��2��:�o�M�(8���,r�V�c4>�v~��J��+�|���>d��� C�DYX�v��-GAU*�Y�ܶ�!s�5����Ӽ%�g���m�"�	J���ƪl��2Q�� ���-S��{��bv�D�4t���ʟjp��>���<��}������H�Jù�<|æ�Zʆ[n2T����:Ţe{V �}J~�����B(��D�=	��1��ŝ�df��u�ь^t�G���H<F��a�Ga��w2�P��\����z2��H�lpb�T��U�ٟ5o+}��;�Q���B,d(�e9�	����g�e\9��:@?�dW��|zW�ŵ���>��VW��4~�;��`F6���G6)���@D��%|���*��m�O����Ғ�a��+��cs��Y��ه��ޏ[[[]��se�O����'��:ϼs���w����?0p2�)2��pX����>�?·+e��s�H]�{\fX�B��h�זS_�h�:�Y;�0e��V�8T������M�7�g�ԃ�:�S�
F�4yzU�3oU;�\����V�K�-+��b���P��c�����(}�h"�c�挗�����U�	A�4�uW)����0����v��'0��7V�� �e:g�X�oz�%������0�:��Mj���r�O�]��zA���'W���`�Ϭ-��%
�r��,�s�	MI���3��M�n:�q�[�b��1�Eq;�6y�P�_.{��R4�g�o�uI��.��*�}T����zP&���7��P�fq�CV�n�����xͩZ)eڌnf(�wyx,�y�O?�T'�1 `X��+����D��0�,��E�pqe����kA�1�Z<�L�qx����#�iڍ�NKtu[�5��,���V|FR%s�������I�ښ�m�`�b���de%e`�%u�9%��,��N 0oI���r��s|p t������@߬��]�:�����gH�H���ҙ��:X��D�����Q�<~Px�B�9;�oK�r�-�)nWM�^D�襤���ʎ+�˥������l:���R�/խb�C�+ŧ���h�|�y{@v���˖����k���f)�xz��ǕdW�Q�w
C
7����^�/q+�Q�7�����YĳV��""�����mL�rW&m�ٴ}�e�Xo/���q5��6}� /A7����y�/��Z�ύ��+�~���jn+'�ங\�u�V��6�U������T{���Ċ�o���ƒ|��n���mĽ;!�LRdY]�& Г�q�\'��V�a��btR�XGGU~%��B�J]JFw�ks$༑�$��j��G[k�����%1җ�yϷ�^f�1���f�7"�Bq��5y�o�y�C/�!3�����:������
��;�р�W��`�E�e�\��8q����@k�\��<c�aј�z�^��Kҩ�p:�?�Nd��%{~�0�fĎ��vA���hd�t��� �`n��=�(R��'re�Yg�I��Ef} �f��Dd�w���	�݊�te�R4nk�[���R]��G�3S�ۙ.�U^O��x�&�D��\Q,�s�$9�a��M�_P!�
&�Y��Ǆ���Nۣ�gZ������ =(�.�z?�Zua%��B��Y��mvs�D��{�5��v���LK~�㛠���4+:1�u+��z�RPG:?y����o�.HQ��=i��X�]i�{�h���P�H�u��A1��֊E�����]7fJi*�L��< ܩ�����R��'�cs���vW�N�v�`)h�P���#��/�*G�xR���-�Ш�?k��T�pc���=�&m�9�1�']�l�4/�L�d;'�z�H��G�o�$T5k%3_�����l$Bs��#�,Dkv�g`���l�e�?"�:�����q�d*E�	�Vqj���Dl/e!�#%)�:����I>⦋��)��@�F�A��� զ={�u��� �X���r/yu;��b.��w��*��j���f|ps�~3}C�|\���Q�b2�������E,��0-|�2����{&B�H�E$����H;'��*M��Y�!;ӟt���=����Z��+x�lz����ʿ�|X3��@�e.&]`���)R��8>��^��]#���ե-�.ߦ��y�>-48��'?�y�>^�m/WCd��H��&t�W�W�8�_X��.�Z��v�gC��G���{0�_3bSɄg�Ď��߈��Q+�Z ˊ�d1~���V��%c7�n.uW1L��N1C�և<NtaTj�y��� ɸ/�(����7vx�\�� ����c�w�����;ZnZxY�]�ʶ����%��%��Ϣ�=C�5w�)3��;��R�ϑ���٩j�=��~�~�'��6ʩ�iܾ��UOx�R�@��;�����]l�¬��;����ɳ��(�?띨t#���Ij��u+�y!i_k��â��`R�pT�s����k�tc���xmCGz諥��kW�3��ʊ�U��CJ��-����mUʏQ6�ף�et�Ń۸�h�ß�
����s�pm�g�X@��	�v�+��g9)�/톳m �6�A�q�̌�r�� ��Ъ�=��×��-�c,!�Y�8�n(u#)"ț/0��*�#�[�@�
y�f�\��kU�C1�(y-��.Q?�z�o�(/���W��͏�XU 8&bit2=[�Tʺ�Wo�P� �`�����'&���w��t�2��B	�� ��S뵵\��N�ڛ�,��k%*�]f=ڙ�m��%�P���اm��U[���rb��v�x�39|�F��xV�ק���
��f�����x���� yx�Rܗ�f��{���BM�8�O�b,��z鞲]�Ԛ�]�r��zLM�`;R��i�M�wJB)�#�*Y�w��$�R���L�y/�x�߳Μܞ�ap3�7k@go���얀���>%��η�J�`�!�{̾��]�~�=U����~�M��-��o���ø:�`h��1)��t&�g�r@����y��fn�J}�T+�&�<�\ȏX~�M��@]��
���>;��[h�TJ4@}�"��]�i8&s�.��8D�ҬY�橮�X�������C��%����k�,�Oh0J[�Ћ �8[z�$GQv����P�qn/t��"-�H��]^��c����j����(��X�C���J�<�O��X�!7�vj:�G0�U�|�_z��k����r�a=P��D0*X���3(V��*��z[>Ag8m
�,��Ƿ��#�k���Ĥ`Fh�`�>#h�D)U�ӄ��U�y�K�݀oAl�k1��9s��c^ ;#�p�{tU1{{�).�K���g��/��,y3���b�Z�P\��b�qD��Z��ÙMN��8\�JJ�l����jﱟe^��p�Հ�͂�κ�f���R�?�>�d|�k���nb�DFP�;����m激Wp��1g��/¹D���玭J��/ƤPv$$��@��<��)쀨�Hs�h1�x^f:i"����
�x)�xa�������0ll�j�nq�<�m���mgX��%M7�.�J�4ZvDǾ�=���QO�i�}�D�9�{��z� s%O�ͅ�T$:��m��Q�:NxPi���j�V�8�6�"��Ժ3����ȉiH ��,7�F��zdv�Ѭ�E�	E���f���db��V�#�G�w&C�l��Vݰ���ť�(͕�A͍!.��B�
�L#6������'y�6wb6���M|q��TX�����g�BGO���#���
MLC���k��!T�т�C4�h���-�_��ׅ3�=�/:&hX��I�S�a�/���5��U]�0�%?�ե�U�v��:QA���R���˞�w�N �o��]V0��D�W>������uRj.�!/a}��8�0j����;��Ļ�mw�1���O��_�j �s�/��L�f��4�.-�wn,����!�@[�y�p�mkU	xmg���i��OÉ,0�Z�j7H��I���}������~D+
?f�k���K�T�g4~�o������W-$j>�/��(�3��,��P�*k.#BP��=2�ӎ�3ų���EX{.�N�$G!!�� � W�u<��l�_͖4 G��tה�?���l�!��}�&�"҆^8���k�YCk�V ��Z�_���Ƥ��F:��g��I�ٴ���Q���o�ѕ7�3$�I�/���wyĲ���P#S�r馺t\�p�~��k}�a�A�T�i��ۭ��zS7p�Z�sB�铞�WzW�ġ�y�D�jfЮ3'n��`В��3�cĂ����10VɇT7�3�ԉ��FDz�
�i�0%;�ì]����F�x�[Q7n���K���ˌ��HĊXߕ�2�oF�p#���
���(L��/H��8yطe��}��M�{<_/��1��\}4��A��>��� @VI-q6�9u����h������h�?��V'Wّ���
 �y��d���t7Cl�+�F ��\3^Ʈ;A�Y���E���-�k� tλ$�������ʽ�.���zi
�bS������WM ��~�����cws2#S�Y����[FY��cihqT�q�j�o��r֧�fHd��ŽE�Ú�=��ɨ�*�$�ַ�$�GC��B�m���t���s����=7C%�޽�Az�,�F�F�A�!!v�V��߳�:���
�O�_~�y�d���D��)Q���t����NC>�̙GTD�`��݀�@��#~q��L�Vy���j[+�����S��I��oR�a���Q��,
X�T��=	�W#��-a߯�;0��Ph�>��55�j}E"�w��0�D�T٠���$4����j��x�\�%g��?��=�S'x��U��;�'�Eh����~�*��?�Kl{�Ɵ���=+�򥠽=:;{\�g��3/c=*i'���Nx5�������T@OH�oJD����[<�?�i�Q�����jy~F��az�����y:x����ܯ=�zN��;��u��
X�߅ZD\���+ %������"	�C���fjf��˫J����/²>�O�����`ˇ7L��w�RY>޷i�I�$������l��fM�y��L�x�	�\G�� g��3�1�i���;&�����@��P���Ry
I	N��u�z���.��pՒ,qMC9�L���+�ĵR��VO��b�#�ņ|�"�4�����Rk�Z�_�t���2���c�ƸJPY&�y�^�ǜא� )��]�F b�
X��@�
~�OS����&{�a���_�����V�kc }���t�
�Nz+���oy���x-Flv����>v(��uF��x�6�d��*~��8OVm-�U�������������py�~�����lS��vC��O8���$�����A�$��S=�q�U�@��r�f2���h�GFAu�;R*�v
́+|d��V�L�T����ē���K`����Js��/�:!܏nu��$��
�5�2U�δfH�.�P�iZ�p� �\�z�E>Fݾ����ڵ��p��jY6�,�������+�`� (���)VձD~\���vX&���5(R�'�k ��������S+)�q����lb�`9nq����g�bKq:���z��n�njSi%��w܇L�7����m���i���2^�QHw���"�C��A�i��&m�_�.�c�>z<Ǧ=��ZN<!M��L�_��_��YbL7p��sD'~"U~�q�_~gt�����|���������Q߳�Ta��lX���v��p�1y���$jO� <�s� ]ч?����;2������
��g$\���d����������ю���_w������+;��S<���&��B�T�{���DZ0��m��X����G��C�a�^�>5�&����Q2 @�`�~oT��Q�g��E��\��ef�W3�"�#��/`0�e7�Xm��N���+�Ͷ�X���.\p��**��c�u+�l;?0ﴹ�|g�_~wƈE��&��C����a��#^ʾP��<��U������m�`f��Z��ۀH>ϋ�؁��Wn��J�:�J̈́o��_�(����)��N4�-z"$��jGӧS�0>P$�|��֎�K��P������b�c�z��w%5z1AsX��c~�VґS\9D�|��5Ḧ����m��O���y������%�a�s{�K��@*�����d���+���g�iؑt|�9A�̾bm_ꪆ��6��)��w����_GZ�*_d�)dg�{��)���g�g�b�W"{%k&x�_�ev�a{T=I��?��Bc�.���N��6�b��s'^�з��7�A�c/�'ުg�,�����G����DR-:>�@KWΕ�u�m���!WXr�sMwUɲ*��HXQ3�����Ҙy�l��*���&�����V�ʖϬ�~._�L+b�NZ6=\x�8����,`�į�b�k�?=U�� =k-]��	 ��a�rNo��7|<�h�µ���,�v���g�#�܂2UP�?J#�u]i�-���j�����ړ,�D<�>=)4�rsk��C'R}N��k0��l���ΦK���I7�e�Cd���f��h�L.��:��}�俰����6wA,�+ahn5���p��@ci���?�<�H]�O��q1��ڙ9��dy�9)�� D����2��
|��((�� �Y���aDga�����ذF+��V�!2�I2���������J�c��fE����!�Fq'�\K��']�#�S#��]�%������3ѿ��������?0���� ޕi������𢛵��:�q�{�ۖ{�ףtK/�q; y�	-���&���S�R���F>ܬ+양VS�@@(p���{�`L��C��E8������)�,d�У�$�����K)�7Kx�JBƱ:�b�ӱ:En��t��;A	���v�3���1 ���幆\�F$�����Ig�KA��tX�ԑ��Б�@	�Y&����{^�"ϱ��*U�d���>m��'''��X�T#��cfo����u�l���g���in�0��uA����7�*�hAН_(`�9�k� K�3��9�۶�ų��\fnZ���������5����ؼ��15��K��Oqؽb�������,P������9,3�3PX|؅YH�I�1{�ލ��Zhł�o]̷G Q]�>qؚ�%R�!��'�s:e�̃����w'�R)>��	���5�R�f����x���A�_ܑ��Qo�R���e����R�:��o:�qh	�W��h��R�#tp1���
~��N���m�5]v���눙�LݝJ����Y�"r�<�U.e ��ǅ�8��S���-�����qlG �E􊒪B�E�o�M���#���k{�	Ɇ6V�j�:�������)��'G��V�����r`�,*��Q��ݭ?�"�Ѵ�g��D���'VC�ǵ����jF[�P27T׿pUGNJ7	G뺵�������%�#@�+�P^֩c6�	֯;l޳���/W���tA�Z�g_�k%U�x������C���R��?���-����]�|���ԈoV���8��wI�Fkpi6q�.]��IC�xײ�N�H���/���J}�X]D�c}Q��Sw��$�g��}3���a�3K�j�Z���:i��V���7��ړ`�΍���yѪ�+���G�Q��Ü��i�R,0�۰)^�ۨ���\9��o�uL}�W�Ӗ�8��u��l%�p���9�O\A���bx�A�������R�.w��H���\�][1p�X�*�ԋ�O��ʴQ�#T��Ρ��E��@�K����#�'��F�`$zk�һ��i9�L7��.p�S,3�C$���5��v�N|����:1?�Z�ܟ�޿-,0�\-���y��y���s��Z���s$,�������?r�
��Kg
��c�S��`>_2�Ia�u�S#L�f���{Y=����n�`�>�v�5l����y� ���Ƹ%����C[�BI��T p��RWdh�z�C�������﹅I�ӚV���+[��z`���~�B��>��ȥSa�h�9�`�r�{���Z�Mw��؋#ۃ�hG6�0�sE�����Dm�K��F��1lF��Y� �#�1ſ���\�Aj������H0�x�j�@�3���x�1p��G�dԴ�~t�C/�yV�6�����,�ȳ©�6ć)��C��u������AJ&զ�_!�[�&:��j���r�I4����%�9�A�Ц݃�{S������y��N��h����-��,���9��3` �'M�7�
A4݋�9k���:Ub흁\7�� $���Wc%�+�$�ed3"���`����9�$�o��xM���&Er�VR_6���k��:nʱQ��O�����J*� `���!1�cb�nqJ�Ap��m�/(��F��A����a�g�<�C��DL
@s�$�w�ݮ)��/�|��0&��b�ؔ�<(ЏF5eSǾ���$���������lC����@O���q�Xmn�J�t U��L�>~�py�$%P��Q�TY@+lPf�1��-S[·�,�4�,P�يE�N!���oEQe���7�hSv&Ńj4�A����4��������Ie<<�.���7�Ulh�}�kQ��ޫ�lP�cb��O߰��<��G�����@���oWN�Y�ub�`ǃ�9����Lw����u�z��� |E�_��w��<�T��L`�4e���p/Q��w�D�N�凋iE: �S%�[U�OP�X1��������`���>8��]%1��h?m�*�SJ��Ow�����*Ia�S�N�<�2�0��0v6Y���+����\θ�nBF��G���5�f�'���Z)������nj�՜�{��kV\*͏?v�9I����I������e9�V���ga��ᜤm�����{��yD����іh��[�Dy�F.���u'��QBd�������.���z��k��#���+�,&_��c�{���r�y���:�H6���`��O��|�7�������N���j����I��R��_�@6���a����aE|�D�/�$�(�}Z�?q7^d免�T]��r��wh4\GZ��7	� ��zY�$8̓yW�� ��UP�%�ep�_C�^��ګ�aye[.M�oF&v����́����:߹�����*xHw������!vIm����������5���|�#|��>/%_�Λ��x>�d�i<�����t�c�m����X5�c皐�~7���� �S�X^3��$ҏ�L	�~_3��ڙoJ�,�H놕�SX�قP�;C�!E�#O|��v�o���tm}z,�AV��T������t]Y�P�*U��\�]�;OL4����)��ei'C5��A��̨_���kʰ�w��P+����\/W�J\�D�Y���JV��*_�U.O�җ��/`5�՚�8�l���[19�j�
v�@FW�*��>�Е���Wv;ť-e�=�S��X� 1�u9Qg+Ĥ�=a�*�%�IT���]�����,��y ��l�쀔<IX�$Q��1� tmm{�=��5&\�*r}zC�1ك��s'����A�Z����=����&�>��7�Lt�j\:#E�n��ϋGK��k
Bq�Uq�b�����ω��r�I��]�����N�K���Z�	���W>�)��P{N�zw��{{)/���fWf)d�p��m%�a~�7�o3a�M!_�)���1��JPy>*\�+V���|�ȗ:�t�#�mZ��ç��0u�[/�q�O�z��K�ו��������i?��y��9�E�P��g�������A{�.���s��N"�;]gK$sG��΀Ȉ�yz��3��k'����|�B�z�r�We�Ch'-~�q��6~�Yt_�ރPI�~ƦJ�I�EI.+��]"@�`p9�q��Q�˺��I8?��:�؊)r��羹�zC�ś��6�h���/��e�X�l����"���ĉ��q�x��W�g'ȍ-�F�
�����W���c���g�pTϞ3�ɱDF"����,���6�׋%�Իie�i:*C���HWx�ٍ��4�.���+�m��)gȅ=���Bd���� ���nCp�����}��%7_�oi)Ӕ�-� ,d��V��M�ݿP���)��a�ҝ^��gu v($�X�#���\"�������n��Wc ��A�<܄v
�����T�D�(�rA��҃$쯟�'=�6�5���˽��e�%�Cd����K�7�v'*�E|@WM���s�&����ǚ6z���$|����͓b�����ThB_�z�M����`��SI��b�Ob<��X@����i@�#��(9�z�KH�g��$�u\6LY�	��O��|7KGі���ɗdv�&>:���و2�����F��!߯yRgx#i��H$�Ώ(���Z���J>�6�]��n��g3��bD�',��������J���t
��!)���,F���Q���nZ%nm�.�~�ǧ��@��r������.�z
1?�a��w;>��3�YD��%ߊ<������_gl���ok+�@�c� n� ^�S��,.vZ3��Q,p����a�� �P��&'�.��3���mUg���]z[_�D0�C�΁�P������*�r*~Hgb�~tp�������_���APA���34�����R=ZR�'���$?�P���W(k��aG�!w8d�ll����-�Ā@�,���k8�kg��!I�`N��Ȝ<s�Ǚ��(}��Z�X�;g����/8�y�Ȳ�u��ɽ�wX�C�gG����r�%1��
��T50w��A��Ч�Y�����g��h���Q}~V��]顔�E���B02�e�w��dd�M������C�oa��<��@MٺemV����p�05�����&2�@�~M:��bT[�3������J��M$n����k�	@>u�w��9Kv����#"ˠ�7���Zn�C�z��� �ui��Jz��z����mUl�;}��܇K�*/�O�B�D~K�␊��AbJ?��5~����lh�s�ӟϞ[iB����i��>��t�I͑h ;���V7��030�۝����J�/�$L��C�g��J�,utE��s�6vE|a�٨{�E~�M��c�ehhu�ȝZ
��w��PR�k�� ��U�^�9Cٖ֜���Q��޸5�U8��HG��2��Q�v�B�\;�J��9�fA$n�Ԗ������z�^�\�mub�^8ah$�~c�*K�3X�/���}�CMo��E��Te���MLy `_��9< B�]���c'q�H��rp�H��Î�k���}鿹#��e�a����	�k�aW󡽦?��[ˌɸ�6;ãQ�y+E�^I~쁓���o�˭j<i�t�/�o��>c���_GFG!5щ���.L3��>�^eKi+������!��`��g��k�^J���J����#�(�
T����5� B��=�nrS�M����,�[���ݕ��Z��˞3��\n�n�0���1Rl��%���}�+u�-�jǺ:1N�͕­�|���K~���#�������]�VSXW,ɸ��X��XC��\�%��w:����(�hGN��ä5�~�?��"	�M��t�����r�Mn4�f�t]l0@9nO{�b�ګԹl���ʞgI��ڵ�З@r���(�əөD��9̧�ɡU)�k�ߊS��X�(���=z��տ�%�� ;�
�1�J�0g6F�60Q�>Kz��N=�Oj�,�ix�F[5!�Lr6�?��� ����5T�Ow�&��X�ʋ��Φ�k�������|��? g�8���t�T�(�/���Wq�H41+�
��K���8~u����%p+0�jG�����aj�E?�Ƈ߆����T�!���.���bex��(%x4E��a[uD�=�19��Tt1�B��ϳ�q<3>,����(�3|~Wqqt�'��/VƯ-ޞ�?����vBg��'���jl9�C����m�Χ����j��H�T}&��n�����1EM�}�'��
�ĭe[2�u��)� ׅ��d�&g�s�C��@��3��5��h�Ok���SU>*5�O�K>xK�#
?����Z��Q(���S��D�-d�^�6iJy>��fN�њ�
�,�s��M��צN��uSj蒡�(G�0��nT��<CdS�~рςa&�#HgW��͎���P3���B����"lb��9��"��p*Pw���;����,��:��_��C���/5��h��(V"[k��3�Bb���G��$jzU���z���(t,�Gӫ`-g�`nE��>�^�)��C��O\P�- Q��U �4�Ԙ�h��	ol ��G'r	�qM���7�u���:�ޓ�� �h�۸_�� ����N��N���]Dw�0;������AC+�|7b�X"�h�1Q�D��\�����
$�2_G��l��j�Է���ws��9%o�:�#�w�~'����c�J�����Nq4���d��턁a����u �e�sd/�<��sG��L���#}�\�LS���n��i[B�����$E�ÿF��Mg�[i[�|��}n-�Iz��.�?��f�]Zp+�?��/�H�O=�����4�2p�[��x��S��	:�>=�!n։�ii�����C5G�-�c_`6sp�ԜKP���âX�R�[�������1G���ԵzV�]�u�O�\#L��G�Vҭvh��_ȉJ ��"l�3���߼e㖎�����N$/;`�D
��]�	�9�/�����F��p(UaKhP����Z��n��k7���,���F57C7Ņ��?������P��.� ��4QTw?G��<ir�	2A�M�t���Յ ~�i���w���Ԑ�G�	S���>���	�_,N%'�Ipo��=dnvh�U��E��u<����W���z���s�v!�c�!�f�VD��yD�Y��Br��<~%�Ĭ\��F$A�<� 5�m�.��Y?8T6p�nj�\ˉ����fʅ���z�jĹ�gO-�ܰ�
��vY������G�o�b���!F�Yه�0�ijY�2I���%:��y�'�E븩��>���݈�ʊ������}գ9�T{��#��9S�x�������oݐ(]����(D�U��nN��&��m����ڗG��tw����󁸕[�)�FIJ���ܑ��sN�gMY�|�B���H�7tT�F#*?�����z�l��2�̪�ip��&�[oy��x6x��* @(������^��"Ԕ�K$��I����3A?��uNe>*7�;�~2�K��#�����`>��IL�GB�������f B�1��1y�&S�i��@Lم�w|���2����o�:���)�K`ۭ����E��cR�7x�s�!�����#?�����"�,�{�۝^S�i@��(�������B8�k�F�)\Y����%$��bJ��I!��s](a���FF&h]d���	8�ޮAZk�p&;y{:�c�wj��v�����\�4�[���,ڵk�<i`�(�ԕ�	l�LZP=�Hg�i�/��z�S�����x��gӆ�{?����нE��C�J0�eZ�ǡl�L��4�T��������Ww�3Hl-x!|�9J�����c��+ �A=�[4��C��e)ħ��:���� Y�;3R�N����J��A��#����ͩ�x��4ͻ��,[�^��[����y~��)��[��CM�k�7��)��ޖ�-UI�\���.T?39̀d�"	G�0mO���׆g&,�'���=:E�ӑT.��-pQS�ٜ�@X��sś�\aHo����ƙ��u?�>����������i�zq.t�S�W>:��ր�Y�!�^�$���T�"��ɭ�!)�os3:�CǦ?kާ�`<�(	g����n��$��Ϭ^��}�mK=�K|~u6�t����#�*�x*w��6�"�7�c	�ymf�`��X<I�L��榳"P~*�6�b��Y�>m.���UL��#T\Y%e���������GY�ǅ�)�3)�5cRI�qk�.��g��Q�U@"����~`�u�Ǿ�Efy�����*�",b��T����G�S�Qb5��A�ˠ\���Ry�M���5K�K�zMki�{+�;q�B�%ը7�Iy�V��<��4>g�M���x��#�a����~�>U���?�:5}V
�J�:���!o@�@k#����E�B�����=U��h;^�&ىH�xrWK��.�v��YgFz0�A�w�[�u�@o��|a�_��!ֻW'��'~�w��#���Ĩ �N�_ܸ���	s� HҒ�z$oÿ �w����|���D �F-�1jՅ|��c�]�����#pЖ���X�k��`B��.�6rQwg�zL��e=�0(ÔI��bR� H?4��8ũ��O,�y q�}ٸ"W�v=�Ǎ�
o2�HX�8�R˪�����ùgR��-^j'웣C���`j�#cC�vq�_�X��d���[�E�m�Jxc���X������Y齯9z%굁�c�w��`R��̫�H�&��c.�����w,�s�V����d_dK����x2rY��۴; �&g�kD;\۱��ϼ+��X싿�h�ݦ��Z�
fs#�1��u��6���E���)\M�?9�$�]&�!�f"F��adP?O6�B ׋,��HN��y�aF���g�+x������)s��4�Z�&����7��; K!y�ztbL��&M�i�.�J�;"f5�i�|��Ö���a��O�\9��ˢΛ7�(��KH�#a�v܅w�PV���X@�:c�T:�n�cNL,`�Usu:,!��G��}�s���[�ME�"�bX�&�sx�ױ�s�V���H�V���&P��5F(ޚ�o��E�HC�U<�q
��Ϣ R���j�i�b���U𴢸���ǥ�Wzb8e����z����2��Ƞ�S?]�p�MP��t��d�Y�M����8zH�cɞB���O��?�ڸ/.O����9�<L�@_u����-��䭧�d�⭴����q���XP� 1�``k\ ��8�e����Jpx�<����~]{�T�>����!��O9���T�1�ОB&=�nf��f��
/ō�$B!��M��oد���GƻaG����G.2Dٹ�\��(G��e?�)į۩��'��$AR��P0uH-�h(�����e�4
2˲ٟh�ǳ���c��v-R�B��1э�����(˂���^�
������}�K�����#�P�N�\�J��d>�uKO�-¾B�Mt�τo �Ak2@ֳ:�����F*�ڟ�n�M��ϑ������pO)ԥ�̞uuF��-ld�������yp�nƬ,�'���*0�Ĳ;�,^�v�0���Bޟt�<�Ŋր���B�ίP������1 "�w���_+V�jѐ�l/u9Y�ݞ d$>~��.�0�8A�d-s�di�mOQV,�a=��&N�$���rYD4�A_G�Y��A�DVϨY���;%ؤGDS"�Dx� ��v@6?<�Ş���d�m�\Y3~mLWc��Tw?D�LkW��ڳ[�,���{z�f�����͐d\�+����"@�]-�oT4�����z�n���`���M�ź���G����6��$�(9m
�`��tO� A�Ok��L$&��'�*pȣ!%���o���n���P�x1�9ز�j4bIF�����Ǘ�+�Bћ��Q���9"Zh�c5%���Ue&5��i(�d�߲~�:Y�t������ؑ�~#]�3`�;�U��;�w4��2������AGq���=��^��$�x��^C^j3X1Jw���x@�l�ɡ6����=+��C���XOҎ�qkE��]_�m8�T ���"��xA��dNL�L�t�0%'���Ny��D�k�C�S!�����"���ԟZ�\	[����I5M�Ytq����{#�����.\���`R�I�?�O�!�S��?f���-0V@����u���4��u8��W�Drd/����d[�+��\A�Zsgp�Ʃ�>�WS��d/IyC��4����QҬHZ�e,1�%׊�����HmT���o	�!����_�����>>-���v��
���=ω�O�*�>�GG.m�ÿ� �Yb�}�b�,�4��0����)뜝�[Zz�R]�����]�U�@X-�v��n^�1d�|u��R�p�6�y�-c�S�{'*�:=�jX;��F�C6i���Ix����}�p� K&�P5�Na|���:�^P�s+F�O����}����\&
�21K�e��%[W�� ����m�ڹ&�/vq��k�֎�.��eW�	�b��U���E������)���.�S@�`4��qO@ry^\- �����T�WԄ�E�Flm;�ጎI	_ɳ�	�X|PY�5^l@J㳴0E1�:0Oi2�ơ>��" ��0L ����|�}�ݘ��[#������R�����͡S��ѧ3��5�B�`]Ց~/���>�l�Q'(Z�6�w�Xz,b�n�W��_N��C�
�w	���b��1zػ��Ɨc�z���Fs~�?�eX�	T�|�d9����VO�ǝ�b ��/ց��'��b;��O-��ڤ�wO�"�����T8KA
iOJC�������a󛠹q&hx���3lg�w�h�7�$�����d2ϗ�N�~^�O�
�`�b�_�I]
�����`�nH-e����DZH~�ﴅ���������o���u��Ql'�P���ZN���������\ �X�O����,uy�/��F��g�S8n��1�EuF}���w�u�����4�j
 �q-j@���u�DӰd0uМ�Ɏ��K�u�Z�T�LN����2r��sC�5k���HIL��	8����?~�g@u܋��M�ҭ�.�8O��o?S������_��ǐԾ��|UIhW۟� .qx��j��鴇WP�B{����P��g}�F&BL������I!$Z�˵M�ּa�/��n�9B�A
��Yf`�{E�ߣsw�.��V!M�T�K�*Ӧ-�fެ�À�Uj�M�u�(oG�r=S�D���Ap�`�Hn��lFX�+�R���]�vVvT��������>�q5�`���� �a\7k��� UmM��C<�o�[��lP���I�����U�FN����-K�dw����,!9����y������Ԉ�q�ˮ�����Q����U��
�
j[X5���menr�<h���������d�Y���~���Ԝ�@��3a��G���i��%7zP4g	���Ug;�߱X�Ldm'�0+L/F��-g�(�!��jȊ,��i�s��\^6��E:4���L$8�3	���;�����Ix8M���ub�c*���*����#�@�� ϋl��9��%���i4}@�iz"��`��4?z��P��q�r����-�-���
Z��,��f1Ҩ4�Ĩo�,b����/5��J�������xX�� ����o�A� Hb+�; (�� ���SY��7*73376\�rߎY *_��\�K'6��-�S��j�^��\JkN��T"��oY�pN�ڂ�n�G ZL�T��Ҋ��;M�� ����y>3nD�L���m4�Wb��7���wZW��uԪK����E ֎�߮�k�y�CAg�~`����ǿ~ڃ;"#ڙ�î��0�K��)L�FR�902�	������N��u|lЗy�c����!���nvS�ѴR�W�ӡtԺ�(��~�ח��r�/��ѳɖ��o���*������,��	,�0�m�Ǥ�#`T>˷sM�ɻ�)m�b��n��w}4+�v�#���+w�f׭҉�DFe��@X����W��u�N�~�Z�l�U�6dg�]� �ئ':�Y%>\3�.�E\�;�Q��~R�X���=X�(g��@�=��,���	�W��%{ӹ/?�d�I%Oh�Fr���� r�p��p�~���Ӆ�'�MX�.)8�;l�����z-��J�(>��L\�݁���W�n��?��J�� �B���}pm�4qg�������h8#�H@unR�[i>�f��/������C#�'�ϲ�-ǹ�]�t��������S�[z�����!�$��U������\����P��������R�OhH����Fn��!GRDI%m�Am/0�]y�Gv$���H�k���Rh����v��`�Pw�gh�!9��Hf��7�R����o`��EH[���q픏9&X�\��3����&	�K{��\�eC������q��<������&�?෨��$�{[���V74�À��!:��9����j��Շ�y�!^�[����d]��ᵿ��̚P�n���^���oO�PtK���́8���-�v��Ü�P�|�U�'P:1�BY����D�yt�&���"2֫c"����S�;�!�è{0�9���z*�ZK?*�Dx�͹�B�0����}�}+�zҺB�;�hVL�Kv2�b���oA���\���5z����x����f�k8kPoU��=r��%��W��.D�`v�Yc�|L-�4'D`洶 R��y���k����NO�M���%d�'�G�8�&��4����b��X�����61��i]�u�y��+������l#�,��͂~�RB�S�&k��Gz_� �ٓA9-��%���ȕ��I;�� ��|?�\�
9��v@�N���(�RKa�P�/�.U)�n�s��j�r�E/�u��!:C�s�;��s/�t��?<�ZZ�&8��=�"|]�!�:ՙ#ӄ���&1d�%����1H]'&�A�[<�뜓�H���bh�q>�	�ֵ���\Z�E�蹧>�'X;Q+�Ha�!�iY��w�O4.�`6��O�lJm�׀�l��O�+ޔU���=(I�j����P�x)/�o7�8�_��R��hG��n K��fw��X��N��gJ���}C|� `���b9-J����}��{��z䌠Q��uP<�I�-���i���<T���e������)��9?�����17��Ȣ�5U6�/�f_;�{Y�>���40�e(�i�{T�Y��T�+�=ː�<��,�Vp�.�*����]�
�Ȫ|���+�u��7T[WR(��h�\X�=��_�W�:��b������H�iٛީ{4������;W�Hl@
K�o�ՁG̚ �&|@��_B�m �n��D����d��	=o�#"���ļ���.C$�F��0�4t^�莭����-b":3�\)h�"'��:_4��PZj�� ��ȏڷ��~:d9�GS��%��I����"*�3*��WVzB2\��rU,D��l�V��w������NŸ�����z��Dg�uJ.�����/Y�h��Fr>o�*��#��C�{��6���S�O7������O�ڱ�� ,�$�wgX�Kq��J@Q_�L���%]�0��2%y'Ь�o�8b�s|V?�
��M������'�{|r�>d�Λ���LS�� �γ>�H~)+w�	�l�+���B�T&�A_#&�jG#���%Q �!m��R��ۭ�	#l��|� zwhRc�����|_OI!#q<�=�i|���E|9/!��F��(�X�b�hM�N7��ĲMWy#|����v�d�����R3K7�9�8���w��@�0�J����D�;/�^V�`���.��0y�"W/Zi,��ۡ�p��S����r�}�'��߂n���Ԩ�֡5,��fe��q�_��r��白?��)���+d۪6����|�:l�*�@O�a��:�)���B�G1�!}�ȶd�7�2(7E(*����*���k�{�MӚ��o����S��c�UJ=�s(H)��t�m�[�?̇ܣ�NHIL����'��N$����V��`qDfn׬!�	ݷ%1c��b��(ll�	5!.��d{�`G[/��E�ORj
O�V�$Xb ��Q��ഩ��C�H��1WfB�y�Qq������b�*W]V�{Y�7L�ڐ���P��:����k��OZ�K����;Iƭ`~�J���e��,\�V�\�~ı�Uhbڼ5)��֍z�^� ��|R	���U���0V���%OL��Wkem�~M�6�|�1q`��M��Vuή,8u��X��j�ih�;sQ�L-t#ɉ)�����W�O�Wt���@�ԉ�XS�����ML�>��U�"�K��μtv��3aI�Ѱ��E��`[^����R���gAR˽a9ڳN��
Ohq�����]IR�����q��Z|!�B����>�W��y$����Q!i�a�D��;M���^����``�٩� w%2��
�?)��^��C��9V�^G��t�'|$����8�E06/����_���Z; 2�W�NG���j'�^��L2?VU}�h�,�o�9'qQ�tJu�0�Rpb\�쟴�kXO��� #?����d�,?�8�<v׀��[�`����tf7��"[/��y3�_��!?�^��[��md�S�v$܁�������~DE��8\�z��3�
�I:���$�MN��/Xv� �n�7d����7�����,�t��g�M�� � �N[��p�ڭ����R�3exx�D��;Kx�����^��X�y�P��2��7��?(�\�GT���+8�A���������h�O:d�{^/����o�\�۟C�;��'������:��O�/EĢ榗�ե���Dh �5�3�N�	p]	L�=�W�FԊZ_x��1�MXoCMN�ZT� ��A��;jM�ߩH��stj1s1gMV?w�̄���Ŷ��xf���	i}��ή��	�1n�7,8�����!��l���Ȣ�Sj�獣�5ʸ��l\��,�����t7 �W2u�6�9n��c?(���+��o�����6�c$&�Vg����X̭2���=�����O�?QH��Ńu�T�����p�K�΄�ؿ9uJ�n�� �v_���k?���_���Eq�-�M�/�� �����zlɚ�G��=�;�+�]I�9 ���B�aL�W��G�A^�,�� �S�p��v|�@��e������R�7E��KTDn�j�;m�&��XA����D�k��nJy7�]Z��8��P3�*�7�m�~���~��Z�H�t9�ԑG.�蔸���1���ȋL�G{�I����KJ); ť��/�rX���x��k�0�Q�dL�昡����C1����$��%/��u���������w��U����ϋ��qp㉅��MUΈK(C @?k�q����T�B�r��%����fHz�Z�*ƺ�m]P��!�K\p)�VWm����u�`k b�K��ȵ��d�r���t�[#�ꢯWE͆0mP�`{ �i?�U��,\kᔧ̚����\��`���?�y0w�`�]�j�����Ԩ`���p��������k�� k�Q2V�T�x9X�I���b�əxR	 � +��)2�h��c�nP����է��{Ӹ^�mC���2'z�2�iP�&��'W2���G���@�U�V��w��},��$0��mŵ	�9��X.���K�&9S\���עS/��_�EC�	s������<�'2��=�쓐�q)��"�kd�q�	O� UTq�Lq�V���}Tr���u: N���0�i5��?�X� �-�-�n����*7�ep��3IX��gW�vJ����VX�_9�%^+so@Ҳ��[�n��u�'Ա!�%Dv}��v�"���F4�Z�"-���O���@���Ȱ��Q��O��t3Y9��5�E��\�
��r �|���^��ƿ8����w^��k�>6mÏyZN�(�����~&X�e��@3�ޜ݅u�Woظ|�/H
Z��,��3��K��K�aa${���U��Դ*rf���мpe�,�n7Dḟ�cٺ�ǃ�)ܔx�������%u$<z��?��ws���.q�����=��I.��F
#�2gX�� �������/Y�#F������x[�3߼I�Ӻ>�o_��Di`�g�3GX|�Li�F�nU���õ�~�Me<��}�]����xD&{ha��?.H[�oM��9)�Nj����x�d�CR���ܳ*,kgq�[���)�T����V¹�^�����*�����{A�����g��03ȟ#Rd�^o�>hՁ�,\|7�O��e�V�=s5D����՟���k$��`� �}�#��� ���V�SZN��ZʎҴ�8�NA�L�8c���Wڊ0�
|�P8\�	�F!��2�=�4l��e]!=��W��-Q�\s�zOL�I��TV�Ɋ%�U�G҄��f0A�-2dk��h�u��A�hQ.�1��y�oe�r�[{�8��x&���(XK�GR`���T��@w�pAޥ=������ �1�mS��a����\�젌b�ƭ��+���^��F�3ߣ{@��c�t�����?���~�^��z"஥y�ZomW������u�G��MNwW  s��2Vpb�=S1I�E�<��cR`;jĲUM�f��_�v���i>�mv�D=j!��Ԝ�gdRڜ�����1��s^��:թX�g����\�����c"��%:H�g��!m���S>�V=[�|��S�)��gM��2je��#j�=��e=�4�Z�R��}*��A~UR�g���Y.�.�U7�WM6!��"�[Sر�*Va~�T�_O���>h!�S}!(-Gb^t����O�k�Q�{i��jp3q�{t�ٟ��` �1�FŠ���D��H���R,�Ɂ��Pj$���Q��k$���<}��r2h�g�w���G�F��M0�+`*��e�����g�/ǜ�h�T7Q��&+�Ի��>n�vǯ��(4�vgW�L�� 3.�^���[������V:䜩0g�]�D�@�_q�����$M��s^$v�O���uy�U/U���8��T��Dtd��c�,�).u�=P��H���{G�	%D�;����in�7q��%h�q�9EM��)�����]ò�c�/�N�0�PV���I�
��`4����<D����	_�Dh0���z6�9�U�M�O���d�Lن!�ݢ0�=ҹ���"���}���OM�`hE�i�v�5�ZF��[s����f� ��~pɛqZ��hJ��h����?�i_� ��Z��uu1`��g�����W��	7��	Y�R�CZ��@S��QƏh�K����s�e���Y22�?���|���X2��Zz6��,@����v�@�IA��ZRb`����@!uNR�?��k]�]"�1����|X7���pm��h��a�4a���Yǩ�xU�>��8+Z�o�7���%� �#t\̋5;��O��ױ�����Љ�_�h#��1Ɓ�����iΜ����w��v���:B��L�ލ���")�0�*��B8iQNK�i��H��T���}���UJ����T�A����5��p�����4��\3��/˟�vY��c�rR���eM<���7.�(�8����`ƠS����3���=jt
��eZ��KJ��`k�\QIF��˲l����Qߺt�p�X����_�G?�Ϯ�2Ձ_)d=��w܆<�����T�O&�� �n��#�E�˻��D�3S�c;�+�
i[�Z���ɫ�_{a� HKRY��_˴�^{�ߣ���	�#�F��ͱ��Z�����ʪZ��
�����:_��wqo$޽�4Π�=3zl��O��v�����������H1R&�.�M3 �:��2�[�oV|�!��Rz=ã����JD���s��5�J]_+�E7F���a��w�����Kr�f���Ę���^�Xu��h�^J7AT�ݾ�L��S� mIN�}@F&�rw/|�?.���M�W�Ӿn37��=[-��sF�{(
���I���/;�Տ��~�^J�����F�1�"����c���M�?�rJ�������_��53��象UWm�ɻ)�L��=�6�Y�_S!;�:4�7�"i���.�OG��,��������I� EK� ��P�_�2iw�{���vH�3�g��=P�	Q.#a�[��v���!��A�7��i/�MZ���(�$X�7ne���g�[���y�|�Er�q����p���x�a��K�$�e��Y����_=�R�ώ�#֓��q"D1��@����OcV�qcv��`qoD���
�O��ї��WʶD��%vTe�r1����E:P�O�)L�D�`-m;{G�A^�X.�s���	k�	��B���8���B�Ք�!��-e�j��$�Ofl�W�u��֛˿A�1�J�k_���(�h�1�W\�����z�=Ql>u
�# ��>j���`0cҎ��(H�q��
������FʶKN��VI(+�s�z"	}���c$^.�����}���6�\ddsB3�Q��)	�O�J�����Z/��-�z���'+�&��8ڌ�aL�<��	�Nԣ�r�6˖�~dN5vQ�{�k�4y��<e���������5��R G9j�4�T������cd��YY=a�8_��z�A�#<v��>�h���F-��12���).�a1�
m$�T��,����3��t�_^�}l�*l���O;$~�B�s�f�)nWU�����S�C@��i(��e 9�L`&���ګ�}x�5�D�/)r��kC
��R�e�>��\HZ��.���һZ/00�z�,v#���j���*z�}2Rt+�9K���TF����!��sT_��"3��%2�1&��o�����s\���m������iB��+�{J���w��%(2�DJ�0���&��#Ԇu&���_LW��bJ(zD�F)����3�j��g���d��AI���]Ƕ��+b��N��@:�|'�3���y�O*8��\���^���D�)�{��\8���)4п��#3S�U9;����� �KI����U�C�>���tf��}� ���2���\(8h�����ܙ�f4�	W��0(x��;�r���0$�x@1��ֹ�y�x�)#h�V��R����Y"j�n)��g��'M�!��@����>����1ohh{�1���MN��D\�^e��5�n�D|"�X�_���B܄R �E���mR�g���`v�	y����W�G]s�����
�����nS��XЫ7:>N��V/7:��݃����| �U㳴�r^8��D/�;e�����e�Q�<8�hFY�!�QD�
�O8{]��z�L�4�ǻW1�R��Dm9��@�Oh�U�C�Q{�#�3��hy��r:�YV���)��ʵ@���B=�
�&�32;@��V�u#��\�[������� �z��}\��8XB7�Ci_���2��A/����o��y`�P�nN�!��rԖ'LC�AK��&����&cר��� �p5,edۯ/y�J4�X�r�{��I��1�=��D����d\�mS�Q�`%4�~�&������+ #�SbA����;���/��{��,��_| �Ǆ�~�,e���3P����Rf���]m����NTnV��nJ2l������q:��(������
�u8TӖ������kX������ف}�����T�f��P�h�/d5�(�>׵���j�p3���g��=LdRrT!���XJ7��p�P������S�H��<�]�F��J����l�4�ޛ$�5��ݞ�DC��!Pjm��p6�S�=��ct�Ӟz��l�H��~�?a-^��M�M���-�g贏(�y���.����5���DB8�ְ3�{Y�J�3?$WI�E�֞�e,m'1���/���Uuɢ�B;��D�H5���$%�9�'t�>��r��cGw�y��2֘�;���H�d~6��
V�|�/�e�l�@�iz)dBu+�[<��@4ɚ!A��'*8��Dv�>�R�aN�)�v��f憁��k�5G��*n���%5��W�Ӫo%�=u�W����u�Z�R �12a�>�eJ)t�+�6Vbyt���& �?�ͮ4�G�+�n���x�bN�pԘ�#5`��Z���^���^�׳4�o��UMIڕ�e\nr�Pat[�����_�xc����p�qÇ����oa}(䴃a��;�4�Ŭ}��iI���F��,��趜��
�&�������f�P�f�N.w����������NAv�a�%v$9K���q�фP�	�gFu��'��l�h��O�KVkE��Ix.I�Sp�L� ����R-��zl��Y��hr2|��P�h���Q���W�'��cƲ��[��.{]�P��o�R�$�5!GU������a�V���C���,s.�aP~�f��0�;Ѣ!��-�����x��x �0A���*mHU�߿���>%��n���N:-�K��NC���
.�yy�|� H�{19!�?����fV��)��]�hqbN���<,gY�&�~��@���Bd�\)��%L���w�C`�1W~8���[�*�D�D:����N�C2
k�qG��ɫ��d̟1�7_P,XW�u���@p8�q�vkwC?��sj]��t8��2�̡�'Ga���u�7i��ϯ���fq*$���7w�����A��v�Öڬ�[��a��;V@t�����M�-L�!� �O�N)�Ng��6!��_QE���nz9�p8	s�Ç��<5U󛩜��y@�ͬZ���y�,M�x��.�����p�(���ˎ�s9]�j���=
����v��I�� �ڂ�6|�� �tEP��w�Ā⮱L���ρ7�vi\&��*{_��4��5����6T��|�
��<��4�~N��/�w>B*$]9"�"��Qzc2�A!��\.�	O�ϝ�8�x��C᭮7p=�F4lB�q��9w!�#��*#N��kP���)E~���g�6RY@ur3=�f��)�rV�#eZ����Ų�	@��r;\�V
�(�%z���
����.�XAU;6��\���!Fi	�ؾcW'��ɞ3��L�%3��<�4�UN��h1�ݺjgnm�*���ֶ��:�O�v��3�a��*A[��@ʹ����s�t�A���1g]� ��kK#`pqFۨ9'��WʬDF�B�Uu3/�k����=>w� ��$��]ߟ�?���H�E�xi���-*�y�sWY�WW���7�W���&�Y0@b�	�>=v�P��'bR�<�*6�'z���Rx,Q�<#��+%BZ��2�K|>}�ۃ��KQ���������["�G���`k�Xb��"��|���$3�������a�]�$3?���Y�z�T�	��N�/wȁd�>o�[�&~���/��X����1$0��5(t�-ڝM�~3e����m}���P��,o",�t30��*��_]8dz�@G���q��V��%N�]�0ꅱ�*Pa�mm�İ78;���Ȳ�=�é~�}��E��v	��z�.�+J�Ĕ��#��K����p&!o�,�x���x�%������&�����+i�)�Erc��|G>gx��D�,Y�O��<Ԗ�k���Ö�鑶|��'�Se�m��=�'�Q}F+^`�!���Vp^v�l;���aЕ��r���C��I���d�-3�I�
�Lӫc�yۨ
U\H��6�^�'-���ڤ�
��y�"�B2*tm��e�@�g�����V��պZ����G�^�^�q
./~I������A�_n��!�ׄ-�^�|�U�S� u���d��1�[��ܔ�[9�җ�pU������p�ɒK��y/G��|f/Q�}7�d��4��z\o
� ��S_=�c��$-!���fG�1_�G3.1{[���'���/��D@��W�G�B�I�`҅njEv��e<�%�JF�_�Fî<� }N,j��7�}�N���y��<GH.�?|C��KB�� �D�H����B5�~\���d0����d�?��R=������ٿ�l����U-��B=�Xہ ^Ǡ�Z{s֊��Tk��a��a��W�eHsX��e��#�-�9��J�Vi�D��������s�-��Ihxpfl,)_��t��|i�^rg^vr���������_������񃁤���:A:�����V#�*���F�L�Ꙅ-�k�N;%w�[���+��xD4�;�2�$�<.�D�4q0���	|![@md2ߡ��k������[O�J�Ѕ ���lq��N��L�� Uz��;T��Xc�,Y�PG?����V�����|q�u��'۠,��&<Y:p�d?K�#bcOk��m$8�d�'.�Ҡ��y�	R��4���DG��� -�f�.�Z ���q��;��j�bn�>��N�Q ��8+3::��t���/�z���q�;V�����sP����5���Gϒ�?�z�H�)�)�'�L\�$Kq:Dn��!N~D~3Tն����s�4��3	䏰�Ώ�D6���4�!ĵ��*�uQ�ƣ��=���5"�gA-m;(�k�)�O}�"� ����Jm��7� �f1gf ��Fa��ŧ�UL�.�⵻X�&��\�=� �c���Q�(Pt��&,��)�����~�{AIh�[0�O����(�2v�2��T��tT��&Q�[����Zi�kA(޽����&�{�&tů���1@�\C�mE�Ü5�
3ە��d��M�o���/�w���569�¡K�4 �Վ��	t8lŮ�A�֌�+�ܾ~?�>ozn���1�䆛�]�'�d��)@�P�Z�+���ʨ�0�T��o����o�<��m/i���:����Tv�c�Y���Ҙ��� rt%C��c��G�(�ꬄ#���v�Z��Hjqy8���О�Z��QF<��p��)��V�cCb�G��q͊1�{1F9U���x���W�.���-����|�?�����J�x��VOĀy��t�$�^��L�zN�WO$�6�mP� ����B�k�?~�Dx�47HMd��#��eDн�G����tųG&�/Ld��f*��_�Ĭ����ݖ��倅Y2Uc̢��#��(���< �E%(h\}��jߓ<�S���Ca4�៪���𲸏��zt��"n���y���+��5���#0%,�>�vm�=8��'5��y�A�<<��[(^����%�c]�K!$�}L����=�+�µ>�.�n�	n��ƶ�  �C�����*me'W�ſ���0����N�	*�{2�Páw�Nx�et�4ntk�x{��`�� ����ߓޥ9\�)����a�0:�i�J�R����O�����k�}��D����k��#��O�W{�#U��ZGϩt�0����|�)�5�wSb<m`uz>�� u�c�<vJ��M��]�
�>�C�����ȉ�n����=#๩�bX��R��>��2w(�~��	pnW���Tڜs����⯃O���oC�%�`�C�Z���z>�Q�zէ�W�[������ɘ$��Fv�9���cBɒ� I;�a|�;��%q�Eo
*���j�_�:��m`���}�C��u	�@㛓����_��9:�d#Yd҂�{P-�xU���8�B���G��[���(&�Jiʗ��ق|�Ϛ�[<Vu�0����p���)1�d8��>1�3�� �,�h��;���B�K�EhŵKA�㗼�+�5�1�F=�}��dǣ�.-��-�`��n��"x���z��E�?4n���nGL���}X7%6H��4�ev�Hm��ص}C���	�x����Oi�4��T>n����[Du�"�&^���$Tv��	��[��yj%�YYc��B��+�et������S�ř�v��w1,T0ݻ!&�ק���^kK�F���K��4Y���8�u�����eӱ����:�&�R�rQ|
%Q������6��6���0*�eM58��i�J��0�(�o1e���?9��L�r����% �?�F��Ln��it�z���!��4�n�~��jl�j�6���6�;�̼�Nm�n����C�m}p�FJ,h���5Z�VF\��×�T��D0���W������V��5.#*B�0fA��o��%�-�I5�R�EUv���;BF�-H��<)�zLX� �oI�l(���xN�6;X�S���UN\�Z���k���g#R���+nS ۗ�蠋c�Pf����V�.U;� T�JC�/��Q~�`
NҸ���K>A���\+��;����1�C�|弒�� @3� o�썠�ģ��� ���H�[�=+�4x��%0k���O�W7�}�2N<u�T&�H+Z�t.�	���	���+ꤿYs.{�v���bD,�t�h!��j�~���0�֥��G�H��v,��J�F��!�����M2�]ؠؖp�q�E���`g'�oz�V�1+a���A��X�<��t�LtC�!��J0�~��#i�Ţw:Uգ�h���Xb�zl�K����j~�-�K���M����[��*0�,��{��s�LV*�0��M�c��F����*��W?�� �(U�c�[�9ւLR������x�!��%�,M�
F{�꘷�_�w��3�B�4�u�xT�cg�������a���l��)R�V��\!���s3���X4���/1+x�ߦ�S��8{w��A�O*@�p��ǌA��g����]��,���U‛�)q���6�������:E!�]��3U���[�8��à��x�nd����j�1lb���X�(A�KI�Lh�����v�WO�;4����N�j)�~�Wr�풃���$Bf��$$>5���jv:(�c��}uM�K���&�Y��nP�=z����tQ�e#|�Ok?�,i�P�B�9�~�Q$�o�ߗ3]�H>q�������<�R�2���a#W�[�"���,
��%�OQm�0���:���=�"��������w�2Ȓ#r��<��cc�O"��~ޗ�Z�Q�4�Rma�m)�k�6�U�۩Ƽ@������l3��*2ڛv�,h'�2��13�n��4Pv��,r�[�;���2F��&��m_&%dM���իF�c��]��B%����Q~*��}��e��dp�%�c./��Z���Ks�IAy�x7��	ڔ�wcF9�`:��x��6���l�ȶ`�K�K[���䢁;Ȓ$���*�R�$P��U2�~ң�kY[?�T�V٫�l�����V��b	mF����u���xA��17�N!k��8�A�&4�������̅��ݰ������7cq��׊5եp4��EVp��ܰA
šZٖ�/�tD?���ڲ@��wa��E!��,�[���ekU�Q�#]l6�Wt�k�em��	�2G���^�3�?1�ZG����:�H����*�d'�&��u5� ��Q�I��=��xS>�B�_ьQJ���h�ś�Iq5h�o�݀J��_�aGL�s0ba���/hø%TU@��Z�`Ih8���FJ�Tۊ!�:Hප?�%��T�ѕQ��� 1�Y-�2p`%yó�*�]�L$�t��f!2��y.�/9��Rt��ZI��\���B����*B��G~0���-�U�H��g��P�ЫE�'�$P�*��5�)�ЁХ��Bs�Q�K�K��j��޸b�"�x�lUZ��'7'��$���.������>Ž���k����sP��#L4����d�U�F<�k���L�u����5�$����z�8��c�~J�D��E�
�iѡ]�yb��)6�~W���!�R++\�'����[r���s�h;O�4Ȥ��2�8���6�>~E>�D���(	�MW���3Y
����0���+7��`��\�}4>3[�Vab2�a�Y���5|��.:��-�*�ڟWV�B~����.F��V?6+�c��b����P�W��� 5��5������ކ�;��Go�A2wIO��.M�qˑT�S��;����Ja�`E�X�cȥ �P����4
N��M@�_!���d�o$���=����m�P$�R�"��+�����׻e�����h�9_'�sNt����a�K?�)��*]���Q�B��R��{�rz*#w �2����\�Q߯�{ed�U�c죞U�5�v�y5aNb�;��}7�����r�T.�q+�����N��q��qC�
u�G��R5��B�y�<:�Ea|��5~I�,:S���94c�ׄ���Vhȇn�,��s�qѧ�,�zx��{Q`�-i�mΈ��S�rGm�\k׫m���}3�L�i�N�-�)�ykVB8{�z�d�?����W ���RQc}��Z�f�,=����2&<>�@f����s��r�nu@Gt�l(;�M�yL��!�W�͠�u1��Ԁi�^�|;�6�к�3nY�`��tr�d]ޑuZ���H�٩����/�T<�'�.�!{�j`ֶ������ f)]��7�̪I��*%���d�Y�1�r�:_�O;�7ԡH!0�V�*k���B�����D���%����_d �it8f��y~d��JcD_IMxt�g����A�8�#�%ƹ,�,������?�%4�Cã����<�u�Ť&��z��b�?p6��O��[z��e�A��<��W���Uu�e�U��F�!���� C��Sa�C�(��o����dI1�T�ij�Zo�AΪ$�5�VQ�v���wó�y���,�(PS��tTu�⺺$w�x�s�z8��5?�a�*��~~�Ӗ/.�W���a8k���.��od�6��7`;Tڎ��������[	Ď��� ~}O�F7�u�(�Lؚn��>�J~<���LZ��?c����(��/G�'��@a�Z�,rF�/J���G���x9"�.�Iӆ,��<Z�/�c	-X^ou�kF��ȸK`��Hކ� J>Ѿ|�	R 
?ע�k���"&2���"�A �G��8���1��"�"�J 7�
8Jm���f&��H�Hb{��Ġ$#��˵�P�/��4�Էߠ�fM�ܕ��_�����ee��h�#1�(�{��j^�e�=�c�jz����f&+�� ��cŒ��uk����ޓ��� �A(NGj�J/C��~�L���t�i{r��6��6-O������X�M��s2Y܀����̣�����4/�P��P�З�@ؾhhiV��S+m\d��������5�-��ˢ�q�=�w�&71�pF�� 8u�I7C�`�g�]�Yr����U�5_d;����"�J��hxX3X?�Zб����p��⋪늲�3�|��aG˫6�+"F���L�	xI�Ox5���n�3�a�qvi��l�dT��
pc0�a5?$*��R~N����@�Ĉ�ENFP�rV||p����CͶrG��ÿDk0Z��l����2��O~W[ez��
A+`0�K��>��)�R5�Ry����]!dY�����ᜪ���o}*M�3��U��Lщ�	�dMD�1޽n��w-�-�&�� �`�])T�,b�'��H6j�7��!{CT��M�J���Ȕ q�촺h���ܨwy����kGx�B��x{^2�%,�� l�$�Ea�x���Mހ�����j��J����fޱ;����m_L�[����4j ��{�xa 8^�������uPI0l^�'�М�D`���4���ec��,k!!˗����s��SX�h��粼�`�]�I=t�ok�9s.��-�-;ֆ�ts/D���'��B���0h��Q� ����EQD=���p������qc�choVX�^�T3f042��cv|i`>\S��O��V��R���K��#��֩a���7��_�\���	�/��G]l&�9V���l$t�ܡ�ya�
ϻ"�)ҏ�nт�+3�+�R��k?:�G��f�M'C��}��l&y��_î���)��=��3jl3\v�#�#�oSjp�eU߈7O����!�q.|�^��1m�\H���v�L��B��U:mm6��bɌ�#]�\�
�=�(�#<����"�+��&����P�ta. ߖ��wVe(U��2㞋��gԡ8F&�T�#���ex	W4���$�!�贱���!}��B en�
q~F�<	m�V�� � �(�C��$UCr��Y�������KH���;�y�S��8���̯�Id�;�w�����\��I��@���cm�hK��V�w�Dn~�����VӀp�<�`�;�b�1�h�uPn���Y���;�#��&*�������Z�i����%A��*~��YEk	>��:$���F
x�O��97�,/��1�T�/+�HP�*<�
t�����C@ppނ���#�phJk g@��EJ�SF�����o�Z��c4z��f����s8��:�Ґ՝m�3^=r8f�&�b��)=q�"mQ*y˸o���}��C�G���ɺ��ޣ�>zM�ׅ��uk��S��b�_C*�b�	�H��3�������)��w��Y�ߊ��t�����N��Ͱ�����zr{8P*7���Rv��<��"[S<TS�� ��͈�M�[�(�VX�_&���+�,u6J�����J�j�kw<a�AYЪzl��u�ŉ��m?Uf?;F^�?�d^O�>���R���:���wz��n�,��bJ�=D�����T���\
���+�9�|t�$y�h�KZ�|ٗ-�C��2F}�X� q�I<��h3Z����4�!���r��*]�Y5)�N��J���@����%���-�글����b�Tl]��>!&����_���\li1u�
�ۚY��s�X�X;�:q��ʤ3��|HΒ�r���f�=i���C9>��t9���m>�H^�+'�[SF{3,�JOE�j���.���I�P�Z�y�\#XF�d�R���W���S�b}���� ����>�ª�y�OS�r�[�@ ��z'S����F*A�6����@�qhwḲK#\�I7����KLk���MJ:�Uy�,�@��~v{H���Ue���0_�n���s)��D8V������)��M�,u$zN�q���A�?�|Z�!
�����/MD9vI�2�����M�����~}�RcTs�0u�Q���}Ԝ3
���<��A1$A�߭c�*���j�� ��	���S��t�F9T��"Ӣ�C�	jY���"���?Y�o�f�P+@ьw�ag�cЏ_ ���W�6�,�}CIa�ו��_���yR�XGFN���'c����.�n��/0�)�s��W���+����ӽ���Q�����J'L��BQU�"jX?�}��Lw��Q"��a�o�Ԉ��ץj���璋�WAځ)��%��0w���}�@����vY�q�7=o�4�A�;����/��]Q�1�d
p�t?��Q��6��,D��7R�0Bʞ��������k@��ߨ�)\���ҖG�҉^)m�����(��-��¦Ŗ>���-쇁�5��)%>��}��T�C",�M�4	I��%t�u�"�ݲD�bt�.@L���l�F;:[�6Q�mN��q��W����u2�(��l6�n.F�4q�'��]�.f�����z�;��n&7*�Q�����-]�j�L���ն��M5"�Eb�N�\��>!�N|~ө(�x�3Խ�Ȼ?�a�byLT؇��=�	�B�|_$�^� UމAB��6���r�¦; ���Qa@Ue��a��3W>�	�~H-`v~�{!�W�4��8�ud@���[�Q��6�+̖��P���Ô(�C���Bc7�!�J,�����*���*a���QC���[B}�,,N�G�]�x���W����6�U"�Hr�"�@�y+�7@G��О�Vl��εƎ��v��--B|e@���#��9X)Ϩ��!H�J��}W�W0s}��MFI��Vb���~W	E%�Ϧx�ʕ�?w�C�˾��I�:z���w�HҨ��Tg�)f9�+�Ѝ36�M)J�'1��e����4�=&��Rӑ�,����	X�FL_��V*���M�����(����S�S" J������&,3�P�s����2~���A�y�� ?���W�C��B��>\]�	����)\� ���4����(�����'m÷?�7��(��t�}5�Tsdo��	SC��!�A&An<Ά�t��-�0S��&$"B��:]�Zؠ�V)X�YzV5����"�]'Q�\L/��u�Zs�.	B�����`�C+Ü��?l�/��s���ؽN���SM~)�@�gh[�-.���� �!�`��:��Eb �����Z��������t���	3%
��H+��{Q>�i��4�_<��k�+c����>V�c�r:I�ԚGb̞H��8�ve�Q�+����G8���6�a&�bV\�[���+�4��a���t$�)�������'ĂQ���J��"�
ȃ�ه�NA�fB(�?th�v����-�Y7o75gt���S Ӣ���v��;���8B�VA=)�ݦ���=��x�kЫ���i)
�%�K��BHƗ��L����\�s���e�[JGC1+���U��\qI��t���6z�	�3]S�1o�i�:Q��K�W�1!+ȕ�������<Lߙ߿M�8�$v�qO;��Cx�`>9��YRQ0�T��� �z6S.M��~����g�ͅ�0�Z�p4wЅQ�1�Քw�!{��Rli�|7Sz��hp8����EOa��'u��L9��f�.��ec�˹(3]���Z����W�<�rm�^$l��)������%8�Fh3.���P��|8�GL��x�P�[%OD**�'%�S7���
�TF��)�����?����Y�$uރ�w1H�Y���؆���+�:�:[������:=���M�Τx� ���GD3��6ê��&CK	�v� d -El�.�Z"��vZ����B��n/���T+�=R� �r~��#���	��3N���z�E�lc.����ì�ٜʽ�0{{00�e�������p�?ƥ�I���� ����1;z^|pls<i8Py��3�Q��>��8v}��Im�jeqDv��R�=�����"��PWbG_D�': �y"]-�C�o��`67��`_X~�ǃ�F��Ȳ'�/eݘo�	[;�Tv��ܬ~+�
����(���j�)_�_১㺳�8)�wnߩ[�7��UF+��8���)�0� ���73�����@R�ca���������SK�=��R����e��bퟥ�
����O�g��"�A5���}D�'SgE��c�({�+G��~i%R�W(�YN�������7E!�x��;[!����V�Oi�A�,@�H�U5'�0bߝ:�4r6�џ�˛��^�$Y�8� �̢����墫����|@�S�w�;l��ۻW+��&v��+�gy�g�����+�֍Y� �޳��G��(;'.�� �.]��-~d�\`�B�-�����b��1���Yu�����N�=���K�UM_�5֋��g��%��~v���0�����d���cɂ]N��H$�i�+3�m��0���҈�v��=�� .��)�D�Ii0�
�T���#U���U��c�*�,�N�bM��sj���������춥�r�Q�Ffe��G�}�Q!�qޟq��>rX=88W���)�k�YB$"Y˩�GXej���c������õ@����$>�x���F�� 7Q5���6�*�Ձj��^��a�>���Y2�o����T�����)�1�ß�@��'�޲{AZF^LP�w���9�o)��Y
��0�d�@�;���O�c��W7yT����E5��V�d�̅]�O�7���-��h��Ru��J� i�A,̲��ܗ�^_���]�W���51���<B��=�t�K8�������Ase�b�;a'��
2��	73�'�,~���_�����L#fCQ��̛ePK��>	iP�+����B�?L�^q�_R��-6g�w�wt�k3ÈA�i�ppL%��c[N6�ږ�DY�������FQ���{KH�6���6E�3�P����ϷYe����H��"��2�$��[�4n٣��s�1̣�wK���+}�!��0c��B�"f���&ſl����w��&=�x��|�y�C�rQ��Ix���=��� 8q� �<���~��ݿ��˕��E�{��~�اS�ڑ����_�v��d�5FK��_��v[Q�|�fi�U'�i�8�͆���Br���|�ouVy���w{7D<#��.Y�%���6c��(�hN�Ɲ}cI�{��;j�R��� �!���p�`��k���I��_���1w��DI�%�SQ��2�B):�T���!���Rݲu�0�����x��H�IU�^���R��N�G7�_��Lu�vf��B��N�������k�H����g��oۉ
��!�E�]-o	�h�.����9�v��u�"r�6�-�c�(.ک���:�{f��b���MC��^
�������"t�ᕮ\�d�|�t^@�Q�{��g4^�j�������m���Ӱ�i�9xK�HV: .9�ȣODC��F,4
%L��3�u�����ˣy�O���P�2�h�U�y��5ӻ�2�j;ڊ���x�0%N��6��+Ο>�n.塧�Q���b�>�g��� .�`�7,&].]���B`�'���հp؜@��T��q��ͬ9N��z�:)vK��*/�۹eG�g[�����l�p���}�c�a���6��8_�^m7��mn(���ΣҢ< ���p+�%%���$�y��!G6�����
�n�F�s��iO�b��r��d�>z��Fq�D�C	�����!'rܱ�F� {��jӥ@~=X{�ۿ.|fz�I�q2���N.�	35�A#
Q�_�5�U'��<����E��\_�k��C
s�m�Waa؛`�K�����HJ�b�@ژ.F���87F2�\��R�Y����7�,�S= ���Տ�����.:&��\SO�4Cц
͊d�ٔ���Yj�#-uߤI�H�ԃ����zG�!{y�v
 ƣ|_Y���Ie�-��ظ�7k�}�"�ih����)�%k���^@3F!6�Nm�UN����i-ɢ�2W�}�i���:˸4<�@ګ:&j�p�.���<��K��p# h����,��B��ݘ�C�� Ut~�����	dD�i��I�[�3���Տ��o�� ���p��5��by*�K�Ojc[� �S�tf�(�Ko:]����m.	"��V�vt@�e�jg�6ѥx��v����AU:	���@���F��h�-���#��thz�.������I>OUzֲQ�-3��j�uǛ3jr�U��s���H�{1�����!U�*I�"�q�w���B�8 ��")���nƆ�%������C�e��.��K�4���G.�V��C�(~�)#�-�_b<$�x���JGP5 SiOם����!�g�$���BB���f�7���V��b������|W�R1R�����r9V�7����㥓����$a!An��"ߤ���"�!�9�|KR@�jPSd1�m&-VbNYMP1���>��8
�/-|&�(B���l"��gŏ�E�fL�w]���@��,bB2غ�.�p��f���%!��@�{IW������o��$$e�j�8Oϧ%i��&b��,�i���r�,�.�#3�Bb#�v��5j>�}����6�2�8�}��9��I@G�uj��۲���f�p�%f�)���P��V�p'�lŌC���1��?��`��Yd�F;̌�З��V�y@�)�#�'�bt��Z�x������ou��;���E�F��ϖ[X��]��6(�^��QX{]����EE��p9m�΅1Q������4)?����7�Ä���}T�s潘���n^��jc9�Q�������0�������g���y�ٱ�Ҍq�&!���q�t������?5����<a&�%P~�.^ux�f�\�&c�=$xn������_�Jt. ux�9c[h�~v��(�N=�:���)FP�%�*�{�i��p)f���hP��o���ղ�Y\�m�nS���+u������YHlHD`fJ�?kBr�5��z���۵0�K��L�bSE)�P/���>r�hI��̈́�m�Z����l�����tAew���<"ew��cMZ
���Mk��@�M�Y��]���p3�un�V�6\����#�Uc��e�Ww��:����d�:���Q��2���۰����ܺ�_�ΐ�	�°7�ۢ����xP9��B�&����G�F,�����yyG'5Z�F�������2�{�%��ݞ����͕S��f�
��t*U=�{��.؄���d�U����WO1o��d��Y�Z+������O����sF��l̤q�E���܏;ucU�VW��z�L��N9���.ʨm-���QR�ہ��(lj'r2j$�׀�r�Ї��cc�#R0�pZ�a|��c5�܏��畤�m�J���Mg���M�:��K���M%����D�����@E�������nS�ʸ@0�9�-�f ���jĬ$�|�絔�8�e��/UÓ�)V��dm�q��Vs$:k:�)��Oa���b��4	���!(J�ƻ�	���I�v�u�`��HJ8j�>�+۔��≚��Oo/����o�zܓ�T�g�E����&�a����Ʉy��>W�.r@�kqS6AB#f�ɇ�Ns;�T�z�~�kn7�n�y�;6�.�wi�%�� ���eQ7�]��\��l˱!�6�I���;�6�B�k�����S�����>�_AT[g@�����FH���Y���t>�5�R�bIM4rUY�I�lww ��Ԭ(%�[��P�h.���Nb��W�!fd��4�]p8�ԑ�f�0=����1(�`bpM��O2�Q�ȧ���W���o��.�{g����0LQ��Eu��8�nSŦz�9�⫗M9A�y����� �:�+u��h3�ML`�&4�����p�Zg��Ħ�b�UU�,b���8�����z�D3�9��F$Ds����y1��`͠�G�
:C[}�B����#rQ���*֛��d����#/���`[���噵��w#�Ѱ�����h �]�^ɗ���I���{��K[�z�y�x���b-���RX(8ʑ2�mӇ;��G|��Q:4S�0�� �m�bUD�؀���7�%��
�v���f?��4�+��,�����ᨧrZ�%U�x_��J�E�6ѰBiN0��Qv�
��5��n��"��Msj�O�x��-[U8�}y$�����!�2>�*H�%N^!]o��O���ݙۢ�]14�t��w���#�4H�/��]5���~��^@S������!}��b�:�L	���R�l}EKhŻD2� �`�n�?��"���j=�nT�ee���r��b�Aگ!�T�~6��^u%r��O�0��T�7��_�i�z���⌦��.�p��d�@�
�[i��e�z�Y���B�TI�Z��]T�Ì��8�|O�?t϶�f�^����y�N[d~(+߈o'�Q��]�"��;����[��>R��N�,��\=4,H�ǖ�u�W01<Le`�{m�lʏD4�}�l�uL�#pa}�OU���ذ��w���jDG�7�S�IxQ8{������jZ��jܾYEd{�v����Xl��F3�@f0��ATURi���X9���}1/v�C�s��G㷶�Ψ�̕px����%��� (��ID�ْ8B��kX5!�&�-�?���Pĕƃ��eG>�����Ne��=~�b�#��-lOS��v~fL��-����{�~<٧f|�S��C�M�V������u�z�61�C{p*l�uy؉/ߒ&�ɋ���N7
����1��|]Mkad &&QyE��h�֋Ȑ=G�8��{7�����3f���<���m�1M�'�m���� �w߃� iXG�:���#�Z����u�����o�q;َֈ4��6\3X�s\��wd��/"�Ua.����5
F��2bbZ��懗 ���� ~�CٲAl*�R沂��Tq�kB���OS�1���2��Ħ���vT��i�[ltDG��k�a7�T��$�:0��l�jX"ͷ�eu���b�:����i+4���HM1`#��aMHI�6ܻ�e%�����U^`�j/T�k /�[����8T��\�1$ΐmia��6������0���O�m��ac��l4>�w�)��8��§�
'��XA�+R��(�'��iW��������U��iFde�
�H����1ֵ����f�����F�3'��Uц5�3#��^��*;��	Dp�=.C��Ķ���J�Դ��w�ǣ��۟�<#�7�)��FenR�Q��E?*�EcZU�0���v�R�.�מI5��ޒ\�,�B�A�$Է�6�][��Ձ�х�kUG�va��'��^�5PzLR�����`8[�d>�1�]4'�wbs2��ɝ~"�Ɛ�Zt!/�H�M)��u4Qی�jQ�+R-�u^W���m���N4^�;�.˪!P3<i����K9dUJYJN�.{H�� ��G2��i�_�l��:�z�8_W�����<�s�?��g�]�[&U�Z�N͊K���L-T�A������-sMޣ�@ �L�`�C)g�N�+`3PL��MJ�Sى�2!�ᗫ�766h��bF.�J��w.�C9 ����YC�1ثUp!J�>^�_��M��˫h0 ���?���rGFso!�=-'#��GVC�"BЂ��탽�DSĝ\tn�ֆ���л8
�#�eR` @�F!0x��EKأ���D���x����×�sl�-���x���u�Փ�ǵZ��`�����e���m�	fqet��.�I��l�_�W��h���Ae�`���Ɇ<�=p�`��y�n���C �"�~��c�x��e[.��$A'�]��3@�l�1u����ue7�r���	����&�CX�O�����ql�~���g�t�4uM��eC5Pf���}�����r�gl�5tmP�ٹ)�ۼ�{�)�[��i���Җū��:�)
y����۝8úW߿Yo�V��=���;��BN�(6RP��cH������ͯg�Xp�#`LU¨��ąsu���-f1~��G<�4��|gET96bE���".�A�(��R�86]�g�r|�E�HAY1���SB��IY�T^B�s)P��|�i�6�jh|�:M�	˱�H,�O�#ȭ��@���j���f����b�xcXȻ?U
��|�O�nP��̓�I�!�n�]_���N<>9FXY����� C�����'aH�XfYժ/��������Q�U9�ZC��k�@}
�vS�ӄ�x��G����/b����kfbt��|O��7�[osT�609m��^��V.�&'�/���
"�\( �Z��[%��lr���v�]�}�I���1�(��黃��r�JI9Q�����?�Sq�oS�(p��H:�:�Ĝ1ɪW�8<q�t�ج@w'J�⃆�������iPLLXp�[�a�[W�r-��X�Dظ����u,�ט{
�p˚�[2�k44�kRhg3�]2���c)=k��0ݥ��-��ѷ��w��%�EA/; ��� M��<��D6��i24t�/-"���<Q/<z�+Z7��+F-�H1v�M�߹YNŧAߙ��V�I
�l�Nr��`���x��tFls~��[�B�7�����v���5N��3�+����P�rS^��`j"˕�uN��j|-p���[<?ǣ9z?םrJޘײ@Q�S`-����Rxf�r�c|�ܫ�a�Z9O�\���6�yhN!�TQR[C�0��Z �ƶ����Z�xoE�� ��n���G��f�3,�nY�2dr�	։���]�k/�b��>C�����Df�]�{�����V�V�pD��d��P' ?����5��KӚIA=�Z-�Uo�7�m�vOQ}�=G�L�~$��Z���7'Ϟ0I��4ݬ�"E��Q��g@�Z=4��`F2�a�7�G�X/
!	X� ��7��p�?~���9��F9���<���<�V*�/�RV_���eǯ��ڱ唯�A%YIhNQ�BD�k��5� ?&:�����Q���A���\���"����hO�
�d�Y�O	\R�Ȅ��0.���#o�wH��\��<� n4?�J���~%�4<QVk
;%3�95L�����z&�����!�W?��LN��G!�֙�٩0���O�.Ôr��wV�{�Eq^E�!bL��(}:j ��*��ܰ���qƿ�_�ȡ*��h����w��v�Q�����,��W�s�2��>yKt?�?T0{���3��p��6�g���_�jД�0�~Ɠ������B֘+��7�"�U������2G	-�c"��~�g�_���S�5���y��)L���r�]�cO����5ORU�E�E�^ɠד��a�p P2&�:x?t��������P9�>�$�9�y��0�(�>��"��:����E�	��܌��j[��d��F'k� ����-�}�oT��hhIqS}h٥�|����@gd��=��NTd�['��x��hb�3fU�FҸF�N���ճ����qu���ʤٽxZ� ��@PC�B?��{�r�Uq��j!����.z��A�չ� �Xb�|���ky�㍰fK�'��G`S�:B�"�Y/t74����k񵯥���]�-��0�jJ>����?&K�|9W���������N��t��R�S��d���n9�l�7�dq�hi�Xӆ����>ͷ~ۃG񺬡���*�i���PD�Fw�/x,	`�j��&槐|ڧ��,n�
e�*��Vޣ�����%5(+�� FC��#H����$�,> ����ڀ�v�Y� h���B\f�L�	���������(��  �P5_��h:q�^�ۿ"l��n��E���Yko�@����o�oR�`؋�H����	��}Q$ǓЈe4ى����vc޼��K|�ę���v���w=L��v\]��S?cue�Cy[�Ȍ(`(���3���N!�w�%-pe9��I����:W���A�~�2�;ďAش����-����V������]}�q��J��|�Z}�Ku���t���q;������WZ��&�	MgOIV<��JK?�ʞ�I5>\Ʊ|��9�͠�L��uk��G�x�����A�9/{v�(��2C��h���8Lmo%+�$\K8?/���B_�[%x9�.��L���dx؈��!��E2�OeX�Ƹ�y(6�ζȣ*�!KY+��%�2��4���]cD���9��C�-�rOH�Z��
^~���!0���uڎ��Y��A���z��,~���R�㜲���^����4F*r��;N���Z�i]��
} ,8'PsS*T~���_��G���Z2�Q-�c��&h����q)�Pe8�����ydy���Er��P��RN��D�D5���q�@
��y"H_
x�YN�@
M_�JС�Z����I!6ǒ=���Ϳ�0���gGx`�=x� R��D���B �]�mS�,�0���]L����j/��޾LN��J���R�[�=�p�ՙk�Aw�qS^��F��)�T%Pk�d��q�����VQ�	���u��j�~����Ƣ�9��@�k6�O��Q�d#�z|J(z]����f��G���
�9��T J~K�?``_��:z1�,��O�:�e���<��=4���V��;VZ�[*e�4�2	���=�A^M�, [bm'�3�W�t2����f�+}�����<�KV�
[{���m�hI�F�s����d+��M��+�|L�m�R�~�	���Y�7�A6�d��l;N��i^�'<�Y�95���-Oz���ȝi߬�C���&D^����"G�M�<J���v.G���v��M�f�nm���*�)B����t4~� �ǆ�&^5�o������L��	��2�涓G��H�$������uk��+h.
و����R�d�v����o�7��W��)��&U4�@��[AP�GN���x���4qhY�1�4д@1t��z�\ʄ�踄@$�3�{�D*~$�W�!tJ} �V��X�D_���g5/x�+=W��t���������D�z��1A�Q���SYo��=������vV���B+7,;T���}�\ϣe	O���w�ݳ�ʽPoI�}ה�%��W�爷U0��7��q�]{�D�6��Q�Qo��w��y�kah�*)!�z27�:��h#�z11Ճ�5DLۿ[�3�{��(���`{��rIB�n���C��-h�!~#�%�������20Sk������5���.Fވ�U���2{�l��9o��Z[��j�A&��+S����>����5E,(�u��w����c�ٛ���On�a��%��0*
�t$Yg�&I�r{���c~�����:��ߺe�����#���B��-�=6���tM�)�A��a#v�n���EL�g��7]7X����{w0�*�e�>)�p��b�����Z��	j�?��j6���w���F�Eb �`�w0M���U|�qm�h���_��5� ��*Te��f����2&�ڎw8E��`R��r�GX����-�˿Go�ӋKФ�x��Qe>�J��W�p���?0}�3�櫹���owg<��T*���%*��Њ����u�@
�@��9@�m���@��U_�ಂ�����hs�HV�wC~���,���n��mبn��+3Gdtp��L�gD{?T�<>�t�����:E�����/����`�X}�ʬ�{B����!�<e�{T���6�x��Fj����3���T�����̔	�\7�{×Mu�p�#�FiU˰�Y�:���X��j���z���`(��g�f�;�#��U�������d,���U'�E���2�૚����j������̹B�
'��7����x��zu�׍���볆�f1�
����8R#�0����A���N��N���+�8�6}
\��a�v�5���{7�e2�|�e̋�>���u�mr��d;��ִ��C~>Sx@V��#7�P�QGH��c��!i_F�LnD:>ŉ��`������E�'�i����h����φ]���j��<�х�]B>/!���k?�W)�oIƄ�C2U����H��b
�'�	3
u�������i���:<����[���ׂD{����uiUPU��y��(O01Vr���e����a��� �����I��`K�B+ ��$�S�:CJQ=��yh�f��?�7��~$����xY�R��8E{u��u��ne0��� I�>��a����gg�)�ƛ�MAp��Bù�Y`XĂ��h+*D5�S�t��	4��p��TES4ҵ��yg\���*�I	�Z=�
=wsl�\��"�2�F��������&+���@n^����z��)	�K��u$�g��_ُ19���4���81�IK��q��yg�� �cgٽ[�8Tpˏ�������	�4�wڤU���6�r*����BF	!������<�}N[�f��I�"{t]z�4�J�IEA�{bml�cG�5�߭x�Lʢ�-6������x& �ȇ��4��i2���BUKӼ#�l����X�^�q_���R�UzyuY7U���~��p�¾�t�� nXD��c�yBO��t��b�����2�[E�f��q䂼h)RE�w!R��>�1���N��V���%�U��aDF2��$Sח=�RF����.g9-	j:�e۰��cF]�m�w[�=����ˀ����XUH{��	�*~�믡osBэ�-�	����[I(�$�ḱ��z���|/8rNF��a�=��#6�C��}�L�䬅��eJ�?���m�a@��>�`W��ę��!T@��@$qr�bT��K�O�,J�w����<5��iS�۲n�L�,+�f���[�̖���+ev�D��R���ɫ8���S����rj}�ؿ�m�����<j��&~����Ap�8��M4ns@t�?�H�����ww�ջ�6	\β%)f��"����J���g���V�6�-���	Ί7�F}�C�"��ʘB%R}�Y��<ᚮSȯ��(oƵ��Kpn�]�Z�!��R�X��h�Q����q2<3V��V2	^�K��(|��f�v���c�Z����!��o"��:����ԒT;af�HT��c�����~���
?6RB���? �|8M�	��a�X`�ГOv�v@��}��m�cL�ښ���_HD�"�o���VR�l��4�m�9h���r��.A�%}����%�����8����������>!H�A*{#ؽ�y�?7��-p��Mn̉�%�o�y�=/!l���z�(!��$|�ڟ�2K�
�ףv�D�:��x��d���)�~��25Ȁ�!���W@*�^��%Ϧ1F p-�>�E#@�#���*�`��K��,q�X�k��'L᳴��"nE�rJ�6SM�7�*Q>6e�0m	�`ī�:�.y�n؍��o�s��ØP���Zߢ�vb�	%�ymHJ�����l�1s��{ �q��F��k��L�����^�͈��r����k9P��w�{�HO�wْ��ݏ�����4�#�d�u���8��g�3(~�OQ�yw|�X�/m1a`&��4������6�<�5�9mt�S�@.[_%�Yg�ex�&�ݧ���t\ők 1L�rA�ݐ���B	�'0�z��vX�Jx��F4�2F��~�Ñ�:�`�/2&zm�.M\��^� ���	�&w�6��2����g����ݳi��-:r-g� ֟���r����U"Hiu���y�t��;�PQ�4f>|��m$����mG�Dae��Y2zO)�6���H�Uw(�.��� ������i��Z����z.ѳ��7ҝSIl�6���"#��[�Z]����ݶ:��v:�oP$�P�rN1.���~��<CT�/����E���{lz�?��7_�N,�x�|+c�YЬ�W�lzQK��
���-}�]yxP��_o��6)|z��d��������
�+����b#}��/�y���B�/;2T���V�{�O+�0`X��Zґ�����>���/0�wy`�xJ��`��-i6F���>W=�Ӂ�e���K%��p0�ݏ�-����e�SX���e��K��e�e�)ЪK�P��q=Q���8��󾄽1��+���m��
��(�s� ��UU�+�o����yKQΈ)A�T���%-��`[��r糊���0�W=1G����{uS�[��KM5���!��� 8����Y�؊X�'(Sm*�T%̡���Vdyy�����㦱I�
ay���t-Q&n�M�����#!ꖍ��j�O@Rx���P���[�� �!�1E��.���yO�I�<�"uu����M��<X,��&�?Я6�|���}�$1Ǟ&���?*�P��ޭQEbnW�R�D
z����"�.���3S�2W�n�c�u��ͷ�vu{e�Kk�xy%����26�E�}OZ�%��rl�5���¹��b�4�`�V�H��@�JD]O�'gZ(��+/�����D�1g >3@8u�|�;ű7J�yP�p���%�СR��${��6*�����1����>����#0�${��;Z�Ғ����]���d��Z�K�5���a�Ǌ�L�3Dz��I�1��<�X�s�rUL'��s<��~�R��=Կ�Z�Uѷr�YY�����F�i� �v�'5ZΠ�����'�����0���5	���}�����i��x�[P�B���ڷ�/���'��s�x\��L�����q�v]UT��f�j8v&-���� r���YWBb���$6�׌"e�1R1�D�P%��i]�:Хrۇ�_U�#�j�Ď���TO�CFZ��*'f'<�������ERY���s��;H(�o�S�PYq�ը��56�fq�䦫�U��$o�ˎW��Xls{Xe���A�ܭ���#����Al�C�� �Q*�x�qЌ�]�Vv-fb,��&�kc���l����;�H?��]��'c�B�x�F�v����Z�餟eZh��������o{K�~n|�a0Z�K̰)�wH����.�rN�o���{�)�M��u��[G�㈋�<o�el� ����\�R�=��
u���-�W�̗|���ߐ�A�ru%�1߫���_Rr�/�F�7�-��\+���p*J_ע5�k�(�1�`Q�����E�=(���ȍ[��+r)e)�����2�B8�������w�#��{�! �P��ʑS�	��t#�/�Tb���R���:�1T��å�/чO]Ɉc/�Y6YA��D����JM�C��pФ�)Hy�����M7Y��e�������ZY#{3Z��ΰ�Qo�����+Wԭ����{�a��p���h�_C�4	�	H̯z���=D�r������?J2���ح�'�����M�"^s����K	1��6N�̦�r0��W\�SI�a=��ְŔs�7k��\�H��G���C �Y�U���̥!*�T�Pc�"��ށ%����=��ssRJ߬��Y���J	kI���i-9�% �m=r�.��诿��q�<(�j�<�\�U��j��l<��5څD��W��b�85�+�����Qx!���u��S_�|'�e�������i��nZ��y\p��J�N�/��e\���G>dT�=�b`��:"�r�c�<�s6�uB���M���zCZ����t��o�F��Q�i�jP��!���rq�ס\_��f�W}Z�����s�SJ�mvC�@������� W�a#_�*���+�,��-���]K�@�w_���NCx{|Qj�Q(l�1P�6�օ�=�Wr�=�͚�&���>(�G���<1��?'?^s�����l���,��y��,[���}��=/b�fy.�1� �NMt�<�����T糳��9U�<b/����D��D)��Ik;%���� C#ш���v�=�h�f
�x�%���M!�WiNa�AEyp�E����nQ�Cgl��K�b�_H;�+X�HDǷQ-�`4ʲ���2�rH(�Ai�4o�<�~�H�a�g�*`Ƈ8|��o"�(�g�ʜ��V�	�.��R����<T����{KN���P����ף��W/
|�q�)�O�c���A���	O��-�_��`L~����Y�bY�, �DGrJ!G7i�`{V��g�xW�{�����8[B^�= Q��a�S�A��L<A�SP����u�D\]Ƥl̈́Fg��b������()��!A��7sCH#�'`���)f�I��>���Ng��F!�8HE�[\��w���O6nxB'��=�9)[�2� 	v�.@lP(ί������E]�p��XC�m�������29Rs��.0��_a5n�5�� ���~���I	"B��e�-�C8�S�b_�t�Sx��`�?b�"B&)D�t֋���	���a�o �3�ȁ��X��akL����ZZ�k5*�D���dpv<]Jbpf�Ͻl�y���9F{J*����D��� �%���1T�o/=��U�h��N��l� �Y����.,�CCJrl��:\E��L�7�e��b���4Xs
`m�m-2Ϟ���~WM�,e��D���[�k��^������Gt�����2G�g�{D�\	��=�4����cO.�S�B!>
Y��`�Z��	�I�I9W{�	���J	=J��5/�
	���yZ%��������m+�mx�C�� ՠ���~�(z�ho,R�?�|=l��c!zz��s"@o��ǋ�'3N�Z�ڙ���G�y`9gr�<'ܜ�Ff ���Ĕ��i�EJ�q5a(d)H�o��dv�7�=���25���*�9��]�`$������	B�B��o� 6T�g��'$\����.�M>J,j�Y���Sd�U�b� ܪT9��)�_�
5f�����}Al6�íJi_R�xY,�_)�vB��p�05������W��!������tazS�E?�i��_)>x8��c�����ft��9��ޟ���2����)�C����% @K��L{0��zڧ��EI"���d.>n���|WK��]�8_	�Ꙛ�C�>R�2��VymҚ�-ˁ��,��ӓViZ�8a[�S�����Rɀ��m����G�6H����HO����,��MMO ��{��q�=o��e�5Ѓۈ�}���H){�nq�$U�jw�5���t �k:����xszIň~���Y�X��9p둽�F��H哙 b� ��Gwp1��e~�ߑY��"YWLl���]�·�^wn�ސX��FF~���myVq����S�wE�5(��>M�,�����A�
*���!��ݘ��/td����֗1=�Ӿ
���W�%^�S)a�!�缛�n�[�|֟���u3�Aگu�g��r���~jq�5	����E�KC^C{��AuaCu��f����9� zl�Ǘ��d3-v�o�I�#���?a#ApEy44r}�x�m���M-N Q4��@��
ḝ�!빆*��x��Тre�y#�����2-s��k�r�2N !'B|m���v���C�
���� X_gͥ�`����5�pX�h�i��5�ddMY�Q�~��#�`N|�q!Dj"ey2��Jr���<�h�X�J�Ǜ�f���	��������5	Ms�DhL�2Wa.�vhnϚҤ�=)6t���2���E�`0r0��zU�/y�I�3'q/����q�
:�Dy���S�H����F��7���o����0�D�u�G�H�p��# ��?Cl.��t�A&Ց���x��u���B��k��n��gj�.4I��0��Y/4����<��v��B"�ÞEh0ar��.�R ����>������Nβ��ckZ�'W�m:�y\��^��+��� �z��&�ӔB(�:l�����W4o��Z�fڑ�	�q��'Z�5I#N��g=;�Yr�]w�{Ȳl�ܷG�T��o:� ��W�)$�9�
;��쓤QFJ��J5���wL�vU�qD���$ �6��r⡕�V)d}a�>Бt1��in ��p� �f��,;yř��;I�"B������f#%�s�b��cܙ@"��m(L$c�I��g�ZsUȽ:&-!O箂p6�wٮ��J���p
ă!�5��M����'=-r�x�"1,�{NݻC�Ndg��Uo��G�tm�adO�N���!�-���������bc1��Am��B3ay��q���Y��0Vǉ4���v�T�xc	:G�����t�;��ø��e�e<�i^�}���*��� ��Z͛��`�@��+�]�~��ºx&�3�en�'E�5�&��=h��%�
s�����g�Rp����ʊR����ܓ����ޢ��&r�C�N�yrנYh�¡��0?����RFj̇�Բ���(�y{��XV��>(V��^Wo���X�S�@�}y�[�J�u�T�Ȁ�9ma�s�#>v~�*�Lk� ?�i���(c e����r@�!��v�X�l}!����D��+:�GO9+������mK�'e���>��ͨ�|f9m�xJn{N�t��o/�G/V�6hZ���TuA�pb�0�_��?*���.+���g��!��>j�������?o�.��	�i�G:X���Q3�X���!s�e�\q%Tc�� ��G���%��+����Ł���Z�N���dG�����YUź���2&���_3~�6��z�n�?�ת������of�5�(5�_k�Ս�|X5Hd��p��[w=�
@<��馓t��WX6�e3%�gN3�h�uK勌|}�ѽ$�`��P!����*OI�\E��aP� N}5���0muaz�jA�L^{Pѡl�������/<�v2|/�C�Ǟe����`���أ:�]���ITH8u�ei����o׳?�wOP�zsˊo *o��^N��ģ/������Hl6o��Y��ٔ�b�V�U��0�j��c��ܽ�$'q�[���R��^����<tM�Y�;WY]�G>�?��Jh��_�j��n�I���^������O.��^pr�����ƭ��������E���S�KYY[Ƥ>F�R�W��#s��$6y��@��L����"?�tJhW!�掚��ͫy�Nl���r�p	���w���!s��D��ن��ڤ*,��&TqWԍ|n!<�c��)]1�CE��� <6�$<��#-�i��}Y��*L��rad|��6?��L%٫���AhI�i��D-�x�~�f�aq=	U� �� �B/����+j.}�y{�z�
~�N�#Rj?q�ѥ<2tB>� >��٢
4�������p^��Lfԝ����ό��;&Zr��#�+b�����H��n�/s�JC�*�P*�+��wʙ��5�Im]j`CIձ�>�O~%ƑR���c�c�Ľ����mn�m������b�����ބ�6��L��n�%u֙��+��.�D-�	�����p�>aXW�8PX]kL�6'�3@Br(�@`?���ʢ�h�Lڲ5n�L2�4P,
3��'0֢���`��I|_F~�tA��*�z�������*�d8+~[W�?9\����V&�G�<�֔s�ΰ��b9ŰJ^'H��L��#�F%[w��%�TW�s�E�{���5���`�jr���rG���m��&��̨�՞�d��r����0�, >��+oc	�3�9���"�jj[h�G�Z�tH/y�w��į�csg�+}Z[��	���Ѻ8�㔚|Ǌ�QB2ȪB�N��'W�n�j��i��
�B�>�-$�7`n3��b�S�3.2��ϒ�Q�@��lW�>�K\`��:e�okj:r�v���6v�j���Z���Z��T�����l��.�FP���dK4@��<�
`O�׬�=���c���b��Bp'���%��EL���}1pP�8ŭm��U�������QރԤ9ʴ�m�D�U#:�G~�o�b��bFj,�mE\8_���= ֫�?JBg}��a���x�U�U?ʎ=3Ø5�L�(�4%�Њ���s�U��`01��W<�}���;'�����zW�R{�o�{[m+�f2bKdG��vƹh�uUg;v�]AU|8��_��~���W��I#�i*����뭫|v�'u�]i,>��#��#�k[��8�V�Q\*O��u8�BЄ�0?�Qw�C��������{(��T'�%�	02���Քp& �c��O4�F�6���,�.�޻	�m8����zs��*�Ԟ[�A�2u�c���L�	Rru��j�@�c+e�1#e�f���d�����GN��K���뗠NP/�(.,��l,��u�q��i���Z�ꞧ��f�j'
hS�o@���t�<��Y_��<�X`����Aj2�w���r1Y��T�l]�����&Ey������'z�
h�����rB���9I�{�tRK,�`��D���syų�&���^�nՊ���.8t�K"* �μ�{���2��&
����z��Ȏ6M�zQ�����Q.��i&�W�]8�|Fw�Fә�!cd�?�K�Ub������_po�9��$���Wι���q�N�����ple��zOY�� |eι�*��8��5K��q�e�1�ŕ]^�0��J�a6�~闵]�S����+'��i�.�̑�Ve�	:N�ݷ� �P�N�k�f��-�|u�6��h����ёGb��3*R���^A^��l��_�~�QT���Bo�U�!��g����ch�,����pm��	W�1ݧ1�ע��x�Ⱥmo����X��;c�ȹ���5�L�~"�Xɋ��Ұ�A��9���Ճ�2��0�tW^�z��f��Y��5�L']ca�7B���3̠���c���;��q���B#JJ�34`��7�d��zܵR@��Of��t���/��&o\��~4�������h)̱���։���s���A3^�u���;K1�^Lu�l�����T��W�+�(����CK0E�㸦Hqe4)�j4di����=�s9�<g�`/�����]�
�o�4'9" ���n��aу߹v������|U~��U��7o3C�D�>��\�~m���Y �{C��)�7� s��+����iP)=}��+��Ty=�Iu���k��*v��z���{�촙t���Ϧ6��r�v�<��w������j��!E\�ؾg�(�,�S��|cCԘ����.I���qj�C�)�y9�?���պIP�m��e´Z�^ݝ����q�Mi��'y�'�:?,�,kG�Aמ���hf�c��9���]���yW�^(�0|�;�m����,�9U��j��R�Z�O84=������<�����o�N�����ưo.)��Hʪ����6�����I�1��f��w�F�3��[���D4m�7��S
y�Q�{24ts;>���#���V�q���Z�V����>�q�� g�5�B�N1]XOmt����Q�݃���^%y�
�����ޑ�#N���h(>�[e*�SlG�ݷl��8X�/��a��Y�ղ�E$��{	a��]�j��S���	�J&��l���R���bq%+@5�{���U�j�R���r�w��{��ޛ	y�㊇��+O��, I�nϒoCOe��<�H/��������K�q_���\��'�5L�"��O4X��aT^,�CڌNqR�i���Q�ՇGY��z��Go�=E�/�2F��F�>s���M�l��0��~w�rws��5������IdD�<g�,^Yj����ڵ�b1�����,M�`(*�Φ����u���ŗo<!Oh�v0�K�t��.Π�Ӛ?Kb���ND�qԤXw�x�����P��j�Ɛ�¬x�+MI/=������2|V��pn��8���'!��A�~��'����N��z�+��XQ	q��=���a4��nO�^�y��V�P�i,���byM�[S���'��(M�����:��\����߱�2&��ܦ�:| �~��.��~���EUh��V�i�o�����1�z�X�Rk��Xb�P�%���Lz��c��m� �-b��C�R�?��i���A9�豐�����סP�~�I�	�#��_���X{�F_�"9D��ۨ\+$�x_�*wS�I/�\���~��΢.��W��B,0:�5�̯n��[v�nD���t���28�d:��͸s�zb��ގ�^�y}�%��N�y7`T�)0�b�gl� /*���(e�nmH�%Y�����Ɨ�7׌ޙ��KP��8%�	�g��.F6GD�n�87& >�P�R�<���Lև��PeZLj	w�~Oޡ��f��q����S�z�1�q�eu759�A�jk���X9;[�_.��5���}��_�˵w�2����%H90l*C&���x�ּ��`yiO�5-^��7=�d¾o�̭���?��y�j|dӅ�3��o��(�k�m��
�Q"!�:�VX�j�R|�<g4�,��m�����vxZ��b��Z��<R=�b��}W\4�H�|���?=��|4�'_6{�a)��ރ*�ruT
F���J���F�F9�� 	^�UҊ;���co.�v"$�2�4�@dq�琄�Z�tn�`9g�a�X�dt%P�-8�QN,�|�B?O�3X�����c�z�&�G�]��8�̏�2��H�O'I�M���#�Hh���#���P���,�s�P|mݕa�œ��{(�����H{o��!�KzFd��E߉*c�)Ҡ#'������9ѱD��]�2'�'���3�����@�ȉ��E5%Z��˯��X׆�%�,H(F�>�4����
ր�N*��jU�نQ���_&�CҌ��
8?�Y�e��Hn'��!RB�=��,��cg���"t��`��"��5c�2�E�n�Z�Lţ��o�K�A*��paƴ�-$E��~�^ʣ��EtCH�2o5� ��_��V�$�:ʒ.�Ӗ�$:���5����;��揶`�S{Ɓ����l��]`�����nZ��$?c���&>�[�%�χ�O��$*��D}�qJ6�y(�*�q!q��cr�Z�_4r�$ۣ�|HK����E��y({/�t*9��cX�Q��7����
`�"�wU��{��h'��;��ɗJ����%�8��T-^�Z���!\k#j��A��")����*{y��8���M*=�W���	lZ�������o�m��C�����
�<���SA��p�Jvʕ!��UnXȩq������٥�PZm�B�[���J[�~��Q��"Wn��y8��2y����69�N��7>'�Z�����v�9{�*��#4��Kٸ[�byi(�mg�<���CJq�e��&�#㉤��J�B��%����_�>�tFǪ���oJ

j��i��;���e)4-��\�:�>���!k��n/#C�.����\e�`C����F�t`�,�S�����ނ�#�o������ߔ��[^��tdcJ<ː��r���*��������=�n��;G�a�����Op���%����s�NI��t��L����K'��mC%i��RO*kI%�(./�3���蜸ݩ�N��-6cG��׏�ro��]u�i�L?*	��t|�oe���w�KDN��L���.tO�q���oǝYU1,q��H�ՙ/@|�K�J���f���<pHJ�\���[d?���r䥁�����춨Q(�v��;UIU����T�C3"UjE�.�Z�*x�3����C.P��y����!�%����7�Fku��/�3���Y4΍��g/�����1��#�<�	��lH�7�>v�1?j���6��n��;H���;p���Zx�J܂�Uw1P�϶��U
����%z��!��/�P���]lu�M6�Mv#���!=Y�t�/����X�'����˗�w%ǎ-U���� ��3%�k�ݤ���B����Z�]��U�� �V��r&��F�sđc�c)��˟%���05K6N�ܥ����=Iu���u�S����Kb�����ѳ�3����o��mC�;�T\�w�#�6���ф7�X6���~�y^�
}�D���<� �1��0
�D ؽ�73>蔇�#ǌ��B)P�,I/Z�?b>�e��|�X����4@ �nvUZ6�����63WPÔ �&��
��r�+���8�э�7 �
1N[0�x�z��p(;���ñ�m��Ϭ�U�X�3���Z*52�Ș	�z���2 ���[&�*L�崏 �q��8P.|�_��-��8�u��
>ק�Tck�O�f*���h+�2L+4��چ�!��I�������h{���޺6�<۱��H�,�A�g�2�?Dg��E��X��~^y��F��t@7U���2H��}��(�en�>E��[Dh�F
6ۄ�6� v2�p�T�%2�qܞ�I*�>����˹!��$�R�x��/ԁ�R&��6�ApÖ1�툗Ü&�,�'W7�FQi"��*�A�����=э�냗��d\t� ��F��$��S�[�e΃�����\�Z�$�ٳ���
�"�a�N_�6H(�vim��wq}��),���?�$]mv[��=KAsj��&�~U��h_��H��7v�p2����V$�W?�=��7�Z���A�AٺO�D�X>�A��R� Z"�Fv�3�����[nk<1�ا��1��2'{5��ww������Q�����;���6w�V*���qtO~ v���8��e\-�O;�59��-�n:5��u�8�4�C�@|?�Y����w��r/g�6&���h�G%�ö* �| Mxaf?�s�J�f���b$��n8�|���[P�[��,6�4��< �n��~�؊����lA����^�� �p{��[+5�h�mke����I������fc�<#0��)�H!c8�n1�>�����E�Y����#�i�l]�!�o��"[g�y
~������ձ����R�P�ꓥ�HShZ�L؞;ƨ��v� 0R��'��Y����v�X7�1��U���o�j��<�tz��v�ң�� ��)oH���������e���ep������;����R�څu��W2Ƣ�Ԇ_ƅ1lG����~����q�=/��� �\R{����чG�6�S��f�>�҆M�cd�P9�F�{��������i>W�黹 ��D6��8�5��s�F^��R&|�r��m�Q����$���I+�c�5�����)O�G��p. ��7����EJ�����b �6�l�nO[hb^p���G�Ξ�	�3���O7Hf�޲�5O1-��H������[R��ǎ��Q���<�A�_���V
�o�L�S��.i�[��X?�x����j���&}r��-8������� ���J�V�#��� ��G�vz]A�A�Nu8�����Z%�W�DxE
�[C犇c q7�1�Q�܅��h�_�%^s��O��V�4�_�9Sn-�X�9�������ז��JN�d�#<���t����$W: ]I5@bلV!{Al� uiϼ	E\^��T%��>�~/�G~������P,����&��ۺ�
��G��?�&���7^������*u���Nl�T�X䆉��_L��Ī�}_��~�X`p�Qb�/��٣��ޑD����P�t��y	��-+��H���F���-�.��H���*,flo(&�Vf�
'S�Z��Ti=�B��:����
���p��򾇏���eD��/ ��^zDv��N^:W��v.7�f��Mk�X,���&#<�E��{�Lݯ��@k'��-؟�f�mp�S��E����)�C3��Sq���׏��PD{]�Y� snşg mh�����79X����ZF�m�ʜA�ze�����6��uQ������� Y��q��n��9���Ŗ�j*��5����Q�7�����q
<ª�RV����0%�/y��iI��|w��(��9�)#�
e\��u�|m��e�X,�^���ʘH�{��Q�����)�*��� �9�[��]S;6��P~�'�oy. 1p����@%�3;��Ң(}%�Oj�M�h�������l��7����g1Ȃ1]��n(�u.�Bx���?W(�:A��({L��l$��q�_�{`Ϙ�m�Oɓc�/��l�~���	$��'��/�ӿ�je���)��wj�b�q�&:2��,8����Y!y� z���mG/P�u�Dv�r~;��p?~��*���cV�x���*��z,��t��)�oy�o��?Y}��$��^'�F�e��DVᐱD�tM�D���al�M�.��(᭣}v��>����!e*��a�����$�*��+����R丁(>v�G��2�05��}'�i�|���f�E#�����/�����Oϛ!��F.�{V�}|د����3c���O�K���p��c]n�)����W�Pg6��8����>JJ�C�B�l+�9p:8;�(��J��6~�T�(��Տ�v�'|��pbmP�	C�}�ϱ,_TΡ�R&b`_���U	M�y�M�eY�s��Rݨ�i��kH�wFf�ݍ���=�ӑj�Q���:�)��Ȓ97T�g��w>�UH�\�A�L��Y0�,�H�Zۍ]�J�Y�	���/�KU��mb��1ܞ�e��YI��Vs�<�bH��|Y�D��@���}��N�édLp�m �	]#��G�Й��m���f�V�5�k�y��/o�8亼�2xѭF|�9���ɡVe~��ށ�*܌c��q���ӰV�bE���+K�/��	�W��-"m��M��L���2;B�4V��e��{<%�[l�F�!��8�������T�W��VLR;"sus�˼kz-ƃ���; ^ء����5x�=���NN��o6C�0��w\�����Kו����Ķ�Y
��
��"7 s���Ξh"�)�#��)��c{mn#%�g��Z�ge�=�������Z������o��h��ۈh���<06a`�{�-H�^�\�S�hǮ�CϹ�;o2�8n���[��������ԟ-�j�w�v'zGaٙH�D��nY)$hu��T�9)���P�X�~���L�Ͷc�2}���Ė��z>vmI�/o(����Uڒ#�M
P}w�l�b?/�4j�����l���V`궽Μ�?�o���<�ũih��c�_�ӫ�R����Y��!�B(�{����ۓAZF@9�8�mHt�دU�d�A�]n�x�LH���*��lXN Ԋﴤ������:����s@q�4Fa�j��K�w m���&B¯/�F��<6JI8��N9�>KJ�5
5�|�uR�g�٠��&�|ib����l|��F"D�Ds�DO�V�+��J���W;���|��Җ�q�gz�Z�L+��b���x�؎�Hn��2"��A�G��/��.�k5�7dy�R�1����� �9����F���������+�z<#gYK9!�Il���jNrX4��,"�Nbmߩ��Cc��E���;�s����F�Ǿ�?������N��
U��O��Gܢ�����X�5:�i 5�
�������b�ЩfK)&8� ��i܆�Q� Ф��jET��з>�"#���=#Q�>��oP�z3�,��{�L~]o���<ˍ�zٺsfO���A����L��Uhʠ�3ӯ�mѨ��en�Izh��=�{",��j<@6����yf�q�ԗ��>3���ufg�����C����%�V�4�<����)����y#g}�}�Q��Y�yۼj�!� lC|�ɭ����
�97(����5[��Z/T��㆔.�>�ѣ/h���@�]:=�����O!�l�M�}e�LZ��>-�R�p5�>����%u�~g1KqU�ƹ��1��s�b>L��7�<�F#4�J����A����)��TI����@ϮS�(�[$�N��	%忣{�ό?q*��=E����w]�=D@��+H�O�f�ZZzx����_@"^�
9���$����0�z�(�7����g'.��<L�q�J��L֦B����"�^T�cm�,�U^�L��䝿:�.�F!�^
�3t����S^����mZ���&�a��͛�e�#Ꮳ-�������C�&��fe1�|�������pH%����]M$� �;p��[�[���Z�lgW����M�so��s��X� Y����<�߶���
�2��V*'5��4�#�"M�ȹg��3e���X��,Td�8��a��]�G㯜8#�p�V�P�Y%}����	����m�+YiL�8��4"���Y-�ø��v��T6k�8�I��i�c@S��HՈ}d�	�Z�D��X���}��H�!ȧ蕤If�E{�b� �R��z��m�M���8��*���'C8���+7�	����*\Ic0�'�i���k���Hٯ�P��k�r69��1�>nb{��I����XW�G6HǾO�Ђa�z�Oܾ�u4k��<����+DG���䔗b"vv*}Nz{Ǣ�@��i�`Mg�#|����T|w3'��ش��nܦ�o?�}J6�<qy&|�����l���u����t�0��y%�T��O��g��bO�'��N��Y�M)�>����O~�;$5[2��F?Qakpw�����\�>!&�'�gt�������^[������gC'n_���q��v�!�d�ۿ����/4@��ͷ�b.������`B�l��9�t��\\�5��ƚ`����[e�����¡MI�4	���F����7��ً���S���������>�
�rb��*&
��m�H��I��[d:+n]����Dn�����0���e�T���u���2��P�=�������N�h�p��l��1zõS͡IǢ[��O���r���Z�7Fd$z�C)�FN��I3I��-�#q��6�@���Z�_5�����5��Z�����?�˙��Gj}�Z9ˆ�+�A���~"�N����9�H\.�Lh��(�j��<)�?ڛYe�2���M9r8Id+�p@�cv7_/]E<��A'	n��5, S�b%�����Z�,���S�GD� �i�v��	�oҳ�k)n�!"ֵ�w��nc����I�p�L���iT�ZW�#g�'�eܓ����S������Q���ީ���|F�1����;_z�y���`2��������ơ���2�[}���(}`�Vǧ5�	�FDG�c�b�c5�W K
'�U��ae�E�7�����/���9���|.�N E��P^Z�K��=Ou�K��im����rKVX.p(?�B�Qq� � #�_G�,��i�쑴~�����,&;h^jʹ~�+�R��y#�b��/����U��]x殐qi��z�c*r���4��W(}w�8:$�Wz0�y�k�4��1Y�"@��z�HX�WDR(�w{�W�=�b�2W[|DkռI� ��D�u�{���z4X����L,T��n�|D�L/�~�a����i;el=rZ�;�5(F�穀S�(
��oڐ@%�¤���V�Ar�F�^Ď,��{1��7,�������#5�0�#7��h!���5+{��+�~��Vi��z�!�kCX��(��KmVv�%_ݏ�㔧W�;�y�F\n��'7������:��*�v ���i�'� L�7���+�,^��sG�W�� �)O��w�:Z�ɲ��>0P
�����[|pkrUq-���x��w�l��<@T$��Z�z�ۺ�<�?�p�C��[���}�p}Q�Yz�)��q8^M����}�9!�H��S���[��4�h����/֛f� �?g��G_m��H d�[���Y���(�-�� �3���El��D�!;s	^��z�
��p�&�lՊ�����Xc6$/��ìx�\� k֍�|��P�(w7������G`�7ߊ�J1
O/ r�ڳi}�[V��sQ7�8�܍�j����:�S7S�bǾ��~F�+���}k�ǁEZr1��6���Y��E;��FÀg��/[$p$�m훟��F�VM|�	$����>%��/g�����p%�r�Ad�7��!��o�q�N�6i��O�nt�u^1�S/t����\�-�\�ݥ��b�G�g\ti��4-�N����]�ItJ�rݦէ�kI�C�X�(���5���6~8z��hH���6���9v7��s�b�R�{U/U�L�%<�B�G}�`$�1��q-�m��\�+E=&�d8�g!��ߡ�=Y��p��h��C��r(��h��� �Xv�<,6ggg�0E�O���5l¸Zh�(�R�^�2d	�0�s�ap�"ݫj$���.��e?�~,�~"�'�bّޣ�ľ�n�nC���u�k���~r��
U�ܧ��������X��xDf�ϓ��|�踚`��W~�g/7,��J#J���\Ӽz.��0F�Y|�SgÓ4e��ٓ��Dp/8�+�2>��1JM�)l��d�/X.�<B�m��ub���5&f�w"V�J���|u��.�a��yN��ۣ��阅��7� 3��t���ۆ������)+2�D�S���ή�q��'�e�#2�	��?=%��լ�7Y�f� �@��hY�e�At8��z��U`((�\=��#?j�8��|�6���IO6+M��S�����
��ů`<-���p�k5д]I�`&��'��V!t+ �{$�|�_(?��l	� +�Pg��\�u�(jY͆V7�@�����1b��S)�>Eo?�j��0Ip�.�����xZܿo��^��#�@+�5�=���q9f�M�OO���am�")���O�F�<�=�7���r��qu�T˪��k����`~����+�q�	�{��+�pgF7���i�XõR<�䗘����i�����H�j��&�|�R�s����:�?\�&̂O0w��H��o�^���i8`�mi�A��:��V�D���'�/%D״�e�փr�!�����04�W�|$z����;4�]GJ����`���W�+o�55�ҢQ^5���#t��:+x��5P�Tc[(f� ytw&n��p���͟P�"$�^Nw֒z��N����X�O~_��Bmko�f��tNr[ßoK�#�)�"	gxk���x�krU��Y�9�ܐo6xQ�ڻ �cz�#v��"�z]y�'Ȝ�8��V}O�Q��X�g�e��͔���@"�n��evPt���l�?_@: �|X^<���
�����Q�Ì��7iP���PD�H::�rk�7��T�{���x{�9#�5�E���V�� �:$�E����
��>Wd�s\�;!#������Z��� 1��l��6���|�o~�/���&Ij�'�E,.�x��6E�2�h��]�Ê��(��J{��� �ꀈ�4;3��ۻ�R4���� ����Y���%����Y����!�w��m��'��Gd�O�$}�CX3.�b�sEsZ`�����,1B=�Ϥ� �s�Y�G���{o�P_�eL����������*3*��Œ BC�Uɣ�KnT\r�ͥ�Tf8dI1�^.Db$�c���x�����9 �p����Zxކ�Po��=qX3j�֣R�V�q-�.���(6�ˇz�^ �	@��p���E�)�J�Ҽ��v�<�B�&�R�b�5����D� F��w忔(w%uA�%�AɋY��0���DFw�A҉7�s���h�S*B{(��?"�^&��X,k�4�=�oC�)�0e�����@H��O��?�B�6�X7�C�.AR<MZ���VI�7�C3ྩv�p��t����,
z�?�f�;`M�o��q[�~t�O��+�n�9����7�t�|���n�m�����r�a�P�:�X��:�L��|4j�+f��k�ѫs@��^$<8�.5ꟓ0@7J߀�FR�W,��Ϝw����Qp+��?�,�ܢip������"B�{F⹦1�����|9�y��k]40z�npv����#j��X�8���9#��_��;���-dp�J�6M�hhd�����[(vM󒘋�o.���ܲ�<֘[s���1��GA��Uƙ��}QhZ��di���
�D
 �F�͚�'(|��v�����h��S�re�\��\�j
RX���5nry)�3z�
u����'�=%r~|�\��f�B��H(����N�'��|m(��j��S�����+xR➛�?��2K�������Z��K0t��1ǘtw4�ิ{��|吷�0�ls�dN�`"��������I�H�@�:M桲go��D�9'?����.�D�>Y���/��b��v/>{̰�.�K{�� �=��^�Y��UV�4!r`�}"�R����'Y�3
o��|@�c*�{���hӭ���W�U"��[k�iH-��&���Մ��9Y��iE;È�j̳b�`��fS���q����
�O��c	L��ɘC3�a_,�����I�#[�,'��<%��E�n���#ꂟ�v7m��߭��9M����(�o.r�}W���l��E��oϕ��[gi��xw���bJ���(�َw�{jF
EG�%.X��{��&dPC~�\x���6�Y�QŚZp՞< �m<e�We�͘�k�&3n������cw	3FbFz���ʹO	L���_� g��t��M|�zöb����y�+M�6�k#�$�<�s�o��Y�l6���� 날�� $�/���_����I���z���p.������q�[��fh���W�t���%N�l�N�g�4v QkT8�ԱK����M���w伒g��C��/Bϯ�(n��S�)U�2��7K���:��� �͸�m�i�g��Ȼ��O�Z�`��O��
�8��7�����!��H�3�+��+2����6���P��[t"�e�R{��t�%�E�I���^$��U5f���SF�p���@��r�=��.���ZE��5 �s5�s;dL��h���*Ug0t�D���A_3�b���e�vD�h�t�TG}��"��n-�KH��|S'�-�?o��XqJ���-�>]e[�%�<��/��D|(Zl���9�G�+�O���q��"�(/���2��MG���[|�v\�b�����UB��ne��9������d�A(��P�Mq%��^�E��$�Y��b�6$����KL�P��n����qH�fH�zG�^���tIؑƩ�8�ͯ�1b5��al�wxi�mU�2W��������y��0`�������W
�я9$3r��R� %�oQ/j����w�A%��B
BFB4�6�w�l�kA�q�2��l'�@z�rF���M��z�LT�4�b��W�H25�|ƶ�zB�m�s�e˅�a�T�Wyֱ�~B�`�e!.���&.2G��{��DG�%SR��<^oJ�a�
�{���a���˾͈�0�O�����C©�I���f&�r�M9j'p�2[�2��W�ۦs��<[c�F)���V�F�@S�Zʋ���F܌x�,.�єr��{&�I�f�qvGя��|��2����b"�lr�}0[r^;B�3e4�������d�����X�O4U�dH�� ��OH���c_G|h��[mR#Ja(1ۦ���B��Ěy��k��*���j6�n��v /c|"ç	����tjD^�k�H��D���]��d�L���aP|���ͧ�C]�_3Gv��h���FH4���7N��`�-�; ���'��n4@�t|��V��!�
�kO"��u����,d��ԍF!�itp!:����af����P�#��p��¦�1��,�l����)/�j+��j�^A�nU G�,�8��7
V��"��N�+#/-���H���r�)��Z����UT���~A��Z�z��j��4�Q8�݄�����G�xʬ'#�<��-�����ʂ3鳍AeC\�-�N�7���g��3QV���5�'���J�Q�]m��%�'�7��e��(���~���>j!`mm�����.�[�Ut���ס	���Q�	�JXu^VL�n�������R��m�n"r@S�L�6�c��2��L�ߚ�IE��}t��%�l 39"��Hd� 7`DČfr�<qW_�6X96XU�K1�#|���ː��N���pɔ�^&5C�	:�q�9�������	O�U�Q]���N�s���+Ye�|�ֹ$�7ZZx��ڬ��$�/���l��θ���(��ˀouS�6FqK�������b�_A�˖\������I2�le�x5��E�XL�+-��*a:^4�>w��_�*�Q��7 ��6s@,�~���b����L���~va�\Ǜ�Ih��;��f�x~��X�;(r���۪�˦r�h�u ���j�$�	�j�8֢c#<D�%���6`���)�Ό���#�R�a힩D~2Ԋ�����ʣ@z�A�?�o\�ygS�N��^�W���W����{��� 8���΍�<�j~�� Z���Z�A	�v�(��%_��k����!��[룰"\���$�a�j����5-����Kc@���_r� ij�?��]ny'N+���y��I�n9'(�Q�\�7�%M�@�2�2�23G,n���P�G+�͸���)��z+5��vk]�`ؙ�ѹ��.i2�sv�/��Q}�W�ĭ�ufc����RF�l���X	��i�ˎ�8����bL$�ʟ3�o�"c[}�1��_*K���eF:���8�	&�r|�ą7�hS	[#���J�L@3�4Ӈ�n+�\�R�<��6����|	�eG38�Bg��o,�_h�~~I-&IE��Y�@�*E����Ldˀ ��`c��z��2��1���]{�8�
'+��{�[
�� ��� �&w�Qe���<7�&����?ź0�J��C˘��rpsQth�H�*�ߟ�,$�X_�3�ٺ� �HmTؒ�K.�8Ԅ���ƈ3�ƨ����&��+��Q��K<���o�B��P�"�T��7H���k�iN�rDv���V�5Ċ��]g�N�+*��@�h@Mn��!��E�=���#�#�v��M�ܤ<N���C��	u�m�7G��R��؀.�������,O��q�aã��t�Hn=Ώif�t���<������lU��;z^Rs!Y��8�W��@Ċ(������X]T=��0u��b��1p(���T+-s	�ݥ������K�Bb���p�������>�����o�k@`�,�\���}�E����`����Q�ӥGW�{���}A�1��k}�(d�J�d�߭��U�'W��l*ݔ��{4V�T�U���td�B��61` ��sY���XG�p"�v!z�+{[V�~�ϳ^A���#qt���MGe^B�i�u��h���m�����H��*!������eX!Nѥ��e}�u�8�a[�h�9w�
wc'"���(��>��i�e�u��=��4�3��U��_�.�p����^��P�6w��@����D�$�4�ׁ�`�&wXDN��H\,�i/Gg�h�f���ٱsv�������5�5�j	,�ђX�&+���;B�R"��}�>�ia�D���)x849U�.�L��E���.s�v�~��P�c�g6j0w����Gp��[oD�����r��\�w�7�	��]�@�%eѶU��p��`I*�9�Bn�ai��(�N��g9��/mv~s�I�w$Z�mׇ(���%s dcV��+t�������QW'D��ZH��:Cj�g��;&���X�v�v�,�5/��!�O�
���N0Nm�����\��q��KKd��f.H��8`���X�3���舴�{�=d��Sr'('��g�fu��,*�S�(��"7������pՄ������ؿ���w��⢊W�����Y�P��U�:R�\�5ݺ���lֵ��h"��6W,�ɨ�X��\�謮T���Iys��V����{saڰ���:&2emMl�`u_n�V�w�v/Ӻ}k�1f�(�qYƒ�4J|
�c�wi|��ZT�J͘&�O�t48�n��E�q��"�Ǎ��&�����j��#�P�����8�z�Q���q0Zt	8އ���f�|���B-Y,%o+l{_�)i�D@�_�w��G��C/6���M\�W�q�j��X�gnh�̠,��)ޡ�}Y�
���7I:$�|2��">J�d�f��&k#+C�h��FGz�rѥ�lyK>�{q"���;�.��XgV�!�S����ǎ?S�<�Z�~�����ſ�̠@�+��7��X�K�^CC:�����da��B÷�q�Ӧ���;���2�}O�aQr���MO� ����C�8��Z��Y?.&�#�nZ��k+wv��(4�QX�`8��ݞp�0©͆�\�S���P$P#��*F�5:��v��J,�C9�WF�d5���}��d�{���'+ž����f�K�#ZJ�^2:�(_�Q��@ihpG���H���~���<�����t7����GvO�;@�n�e��!�e/.��+�zm?v��;�I��5��xOFc���\P����85�۩�N�o&�W��E�Yu��J���D8b�m�RS�2�K�-�,15�{$�k�.JE�_cӼ\�̠z��Q<3$b��H��}>$v]x�O��N���֙�)yM���	�ζ������9m�M�W���vJ7��X��51�Qr�IϢ��ʱ�z7e��>�|laq���Yo���?�T�B׵��i���'��h�/ ]j|��e�өMft�I���?'J\M-��1��y"Tl�)1%O0%l�e<tb�x�����h��/NQs�aM�t�ݴw�A}��(a1Qb���
^�ڟ�a"<
���]������yP]�7'H۵�[я9���4Tg���ʲD'馔���OBpm$i�|G��;�'��l�S i�N��Z+D;��jE�Q��i�B��x��U��;<?u[%�Z�51CPO�����h���|`�V� 	r-ʀ�Ƒ;h�D¿Ʌx��&�{w|�X�-	��1��̳أ�\��x��]I�h�oz.9M�:���ʹ��_������)'�Q���OV�!�`h�en�g��5����J8�v#)�d�|�m�Lt�#:GW �k��L4��r�fw�M��NY8VO�-�nʖ�� �X����p�K/�D�ԺhK��|��b���*�\��b-����p�����Ý�]x{��������x������J�*;�
�cڪ�|��ݹ�t�7�� �/���wZ��55a,�h�g��p�l��Uv���{yeuD����p�E$�--���z�W�A=� MV����{�:���IhF����/0�"�
��_����Y��#G�udO��ob|	1�-���n;>z�3mڋQ��-�^��ux�B�B"�4[AX*�����Z��̚�h�ᥢԖ��]#{��x��g?�_/0�V�M��%�Rq��;.��������[~���B����6ƈbK�������[�שr���!ZW>]�I�?�ɜ�*&
�j��N��BO�e4�k�Nk����t*f�4��co
|�6,V?�@rL��U9_+�����I���1OI:��-��3��Z�W[TU���D}nA�� ���Y(��I�Z�,5�AZ2��6'~P�)h����F��w����ځ��c,�ՋK�F������-�jt	$>�D>�T���q[��_��l�$�p�H��A{0b�F���J��W��I�>Ŝ�RͪU��H����	)�ÿS�mm֍h��Џ���$��‏0�aH�A��ϗ�\�1��GE1��@���<>f�2y��<���̊�b:͂�~���w�Ƃ�6�4�i�@��h�	L�橇ꖃj}Yi�EÔ�;7�#�W9G��y���Y+��>R<~XM���T�V���6D���#]�sRr����(о����& �䗷�n�(�>hԕ�+�1�2����@�Ryjp��U����I7�P'j��Śn<�&h��W�U��!i?����!g�6��|^���\GO��r:;W�C����ӟ�qZ��>Vq7t���O7|�S���OZ�9���R2��HD9>�ig�VY]|�r����Nc�������*ȳ�0�%�F�՚��Iݦ -�����o5p����MQ��k���Ai�����}�r�a��L~?r����]��<un�Ɠ��3D|�Po4�	��L��j��'�y ŃY�Z*�j�m#�r��B���s�����B*��������S�Ҧ!�:5	��G��ޯ�cNl>� -V%m��эˆ=4��s�g EV|�J�'r{�G�/�G�1��4*YH���.E�|7oY��e���)��L
Ii��4���";~�;�}�)iSb��F�"V!n�w%����R�F�b��	��1�y�4�������KJT�ڠ9z�W`LĖ^�K��)�'��2�у����h/�A�;m$p��ۂ¤�yXU���(�v�5�H����c&@2u/�mP��[ $^�+���X�r�du?#��0?Y�\v�����ᶄW4���F�.���
>����[+�H��8C��i�DDXx\��iO~ߠ�w��g����x��-���Gz7�ZsW:��.,�O1��'�g����P�B����׶%��-�-��2+j�uU����$�KU_<���j�?r�4�����3�g��%�����c��.Y�,�Jj�F���!��pXgY�_W��h�[�pP��K�u�a�q��&��
i�a�4����"f䥬m
���É+'m&��6�&�?�*�����6w3�_J{ׅ��iHD���gjd �9W:��u"Y/r�#-q��O�GS�=�R�г<Ӷ��<|�'Pr�p1Aj�[�΀�LF�v�v]~��YW��Y
�M��\/?E�F��6+���32r�Sѕ0��}!�R@��$q3c�L���T�U���Xą+�fվo�p�]cVB���`�� ��p��~�cO��{�#�
��1�Y��&�' ���#"U��9�.��j����EzI��c�s%W�$o�[��$u�j�H��qG_�C�S�E`�"��E��(������ID�Y���?��D� `*!]��oO�
h�Ѩ�#W�xvs���~���k_�l��Z�;�t|IYpl�P�f�|���B��h�i�Ug���>n���i�A���.��j�2�J�-C�x��<.���x`lv�"��z�0٫���d�����d�wOe�4��Z)#�����ٟǛ�j��!������qN�%����v�2:H<h�t�C����wj�VQ�l��H�k:gI�yQ0�R�P��K�ׅAek�qxk��:�k��{�ѳ� �nDp֙�ԑ�����W*�a��7���l�D����� �`���V4ϽkuP���!<��C� W�����Y���`P��(���F�r���]�^ո,�G)�i5�w��X�~���ĝ�����'�{6N� )R���-�$��$�q�
f�~��O����b���m�t��=��ｸ��jDn��=bkx�]JMw�p�MFD��{���ߜzE~�1�������������&��+yP*���\�hS8@��Zb�.�CJ�T�·W�ָu��)����S������UR���U��Kl̓����4W�s��N��Ʈ����Y?���.�C�K���͛��`�6wė~	� ���Z�#�=K��5\L^�:Ụ�#�7V3�{�7,��%}J�1n;e
.�n�A¢���&�����N
aU)�"�s��f������;A���tWz~��O`��8Ȅk�W}�j�C�K���ﴹ�&��LAp�şcԮ��	��L���[�A�1�`o+��AP~�P�Qq�7B�%�/X�I4���g�`y��k��j/�\��Ty��Oۉi30��w(���l?��?vrū��h<�F����n����r��*����Sh�t8:X�T��`�>�lc_x�x��2�@ǯ�e�.�jқ��H|1�s(z#.��8a�$�[�� QU�7}�3B����@�w˓�$���׃.ͦ?"c�rc>f�=�����ŦnA}�T����U;=a�Qm�cŝ���2�Fo�/�K�WB����\�?l�=�ID�QE�NWT�m)!�h[�h��| �F���:�I$in�}h��(�l"�B�$����NI�D́]0��A��-B�x<��*ޟ���&�(�"�{��r.:j8��Fc���>8���f1�V�y:6���mF8���k�G��D)fU��Z����!"�q��RD_����%i�o���6m~�w�$:Z������zLZ.|���>D�h���2����(��ˢ��OT�l��:�biZ�J�Q��.Ӛ��Q��^!�_�h��^"^2���
�������X�;�[ [����r.���j{���!29�*a���^��#H
as�.^+V�&�,��\3��y\�|G�f-5�*���R&��l$��"	��#=�	�ӯ����"T�+-�cQ�ӌ
 ��]~�>�t+�iqɳ����6���2����O���#���Dy��j����u�*U���1�{%U�w�C2�"�����Q�,A}���g��ID"s��Xi�u���8�n�U�Z�J�jk�R�u0ߴ���h�@���@}�"��&Q_y6�J1b��|}J��H�I��3zO]�)8woXl1w6	��g�#����J��o�w&�6[mR}-� l��`s���IƳ:2i~G���6��;��~U��]��S�
�0�>�1�_��s-�L1��~�U���w>oq��	����N9Y%+9E'W�1��;�<`�*䖼3�Pxm�߶���t�>I_Þ��I���+Q�/�Hc�82G�G�y���4���f)��שr�8Wy��F���y�G���:4�r�(&:�;���G;|;���_��	���g��^Py�j���w�<P�fHo��+��-�<�e���m�q�tSM��u	��h�;�n�7��a[$� Y[���1au���<o?,C�6������<��7$5S��	�M#�	�
�Gs\����A�X��q�ߖ����a�@}��_��SU49�I9
@k`=an ���L"���-���'����9�~_� ��u�P�^:)�{".zo��Ҿ�n)gf�ޏ����"Tg�=��N�OSFL|e��)��zM��-:�c~Th�oa���:��r�
C�WA��P1f�Ek����}��s�&{��5@� �d��$.�H´TK^0�xUy_o����cK+t�� -w),��Jf�j���$�K����=����&8iEP��T�C^ה�����X���zۛ$gKg�FYc+�t�J-��&ǈ��>����sUJK�'����`8x��F~��������G�m�Toz�OhO-mVx��5�v�)jP<-�(~���L͊����6���Z��҈=���"�'!���,�@�sY��/� �͒絏{�M���oV{(pn�ҭ��$cI�U���%�}���R3o�ܧ9L��j��x�sU5-���D�	䎌��~�a�@�pp���S���z��Ϛ�T��T"΃W�~f��c;�i��LD����:F}�`�a�4�0��Y�I���14h�o��ڡ�S�!��&x�Uy��L�e+�h��ă`�;^Mae������s;ݎ7��rc�x�0��q�@0�X�	�C���Þ���Y�vS�X��2_�5g)����BEۦ�����wIΰ�w��I
cz�1i�ec��|WLUr�fP5[�c��t<���颾
>��l�#��l�_�7S3�V�8O���X�+��"@�=ZX�@6������l ̣�.��q?�$��P���р�Q@������A��9���P�L�p?F-v�fa T1�3h!��=�q��	��J�?������gk�T���	��e_�+�g2=�׷$�Lu�*[��r�O��^ҜBO�Y��Ʒs*,孹��m�I�G�����!��04��-�%�N��8�mO�p׈���cap�u 6�����4C��[��	-�����	|�����V$�R�6�8���h��b�ͤ-
-o�{4ȸ��uo��?�2���]��z��~��#ſe�p)|v���;1�����wL+�2�R�&B�`%&)\QڔZ���cy��\8��Ն�^���1�@p����x��#<�ל�3�dRu(�.fP5��8g�l��6Zw�w��>KRP��3baB����hQ/bs݌`��M�p#�~|�4�9�0�P������h0u�gU��0��'��(��^+@u�/_��6�r��`�|���2���÷���\��_���%jW��Dp���A
�Y�ؕ&s6T���*����%���#��P�|[�07O����4�nޟi9��ۮ�M�
��& D�˒��٢�U��(-� yM����!T��Q��h8E����us��%�z��8N������B��VG��@�I7)�B�	�ӥ��+ BH���@�ڶ]a�sγ:&�[g���mf�7U��f�6,�Rr[v5U��ɦW'���4�|����+��X(��Dx�������|2I���8M�	$�)d��DF�]O7L���R'�����c�O�J.�h�Mu���D$]AǈY.�1��s��sھ�,��Ǥlq~���9��"����CK/���۽ ,�m׿�Ci��o�*����Rbߣ""� �ݢL�7���d(�t`~D�K_i�/���;55�0(?DD/W!p.��-��N��+���ʷ�A�ѓ� ��&�rOT���o{��[.��f
���յ�,���?$�*Ry�Hz����ITČ����Z���W�ʺs^�5֜i��k�%}�1)�r�Lr�n��^q�c�8�C�U�ŐNE!d�ֺ�P-�J�� ����iZ{�k+3\��T�f,��g�� !ij�H�:����ԏv�X
<��ʷ��_�VYo��ޏ4K���lMh����h���(���u��[�<���?\�6�����s����,�bC�����A�k@�+�꣟�,U��<���=�&�"�D���H͸iu�:� ݟJأ�*�	�8T�-9x[�57k��6 ��t��27Γf��*�d	-d`BW�`_�=�W"6�s�'�%+Y����6�@�ŭ�cb��h���G�cV�2��2���������O��jk<�W	8���}�?�V0�W)�ء�s��>��q��J�G��8��n���y;/�S+Jy����k�a��k�l^�r\l��D,=A���gY�O�fA�?/+U������K�S?���pir�f����/�W��]kw�Ԟ�����8���;���+�uV9�������e���4IKv_��U\Ǵ2
��-8�K ��dw�Q�[pu����\}�A/#)n���_��	�r��� ���5���jo�j�ߵZ> �Lo`,$�5UX�:�n,j5�egU�К�� ���c���f��m�UWG�Z�K.������ƨmӬ�������VQ�ٵA�"EDF�ꌕ���9��[��巽�F�%���4C�����w̠�G�i-��N�C�ӀjBN\_����)<��B�V�	(WqUN'�
F�UŹo�pk��ZK6j�ذ���I�{�0�(��KK1�ܞ�7z@"��@+FK�v5)*��:uS��AOj�7#�
�Ԛ(ǻ�W���p�{gg�6�te�߼�P�Ţ�Xw�i�t^u~��!� k�[B�8}|�����k��<�3p�$a�E��y3ޤ�߹��D�N�s
C[��'���m�0�Ham� �+� P��0��� �����aq"�����'�CI������_�3�@��I�M��e�o�/q��r�b�(�n=[� g�oI��j+R8��)�~�\2���q��[�
7+u��wz�Nl{�^�~����Q�P���03\ˍ�����E���B�H��ݔ�#�T�0v9�}s.���k[��o� !��gV�F/���hy"���ߙDф��H���3�>W�#�5"�����f����z
c>ėy����x��m{E�뮌��`��E�Nuҭ����7`��o] u��ni���V|!�R�d��.�9�'����P�y&��FH�^�b�W5���D��}�x+ ��'�;�d=�-��~?�
?k>Y�ޝ@a-��7�Xt&"�c��Q��c��kg%�E���'�%=%v���� �~�"�ZrE���:Xe�A�הΝ�FX����gxD��3[{b�5H,��̃G�md���4���ʅ�joQ��[�pܠ5JT0�/�Ib�x����"���_]w�)d�yq/�? �M*��Ji���n�ϑ�A�&���<>m�5n t�(vo������߿Q�ц�r���C�%ڐ���v?����n��_'r���!:Uno�W
(���5UH.���<u�ă~���V�����[�e*r���]�߯�<��`����4wI��#T�t!<~i0�;�p�	��]C���%iq\�<e�wK+����/�>5T�������3P�Om1K_G�{lvv�u�������c��v�S����&$?i�w����1׳���ln�^h�6BL�2���]�U�6;�#] �ᾡ�p_YQ��o�;R:�iq=�C�sJ��rZ��t�O{ ����+���q�H�5��}�*,�{H�/Ѽ�}���9lۓZ���^2�0����z$6砉I���ɣ�=�j34��ȮCA����5��1H�S�BبK�P�H@{�k�dlT~0���y�ؾ�'GM�o���?9x��" �c=-��,����q�3E��ڭM��"������g�ͅ~� D�t�m�s�&�߱h��!ǚ�ω�}יVi���0�z0%xB��{��>:9��c<	�\<Yl�X1s�Ѫ��@��X�:����j���	����*{��u\⅙`R��'3�����/ ������h=2BD���0/TH�Gl=q-�I�H{ >�S�	g�n ��t�X��.Y<�@��q��m���Zr`Xv�2���d�|��:=O�H`�h i?ϯu���ذ��.�;�㺭bϿ =�)�h�Ͽ�	h��l���>�Ab���K��x�ጏ#�3���	Le5Nf��&�m�/���Áz���uN��8��`7��J�ǮF8`�lB�q����[UNPn�_kS���E����67��.\̊��_��Wp_�|��R��߅s���|%��Ǒ�n�P�۳15�$bԂ��o�H��p� ����>*P�y�U��|�m�Ǔp��p��g�Wi������gI�6��ɔ:p��Õ�7<�½��,��@�k!����C48�	E��G�)�����>�F�Í�b��C�dl�Q�|����kA����Ra���4敡W=�V���K�߅��t�H���R��9(K>ü=t�ᨔ��ع&����#�����rFƠ�9�����iU�h��R��IR��9��-���^�sD�l�j"����s�{+N�&�^TB*�C-�6cz'�z��>Q�F:�!�_��6ԑr&�vX\B�0\��O��ng���_.�5�E���ٙ�K�����Ξ~!+WQ�
Wv�Z��/�=CF:Ý�A=���Y?9�b���:4��Vm<w��!��_L�{(@P|��P�,'��-'c�UB��'}��g)N����u,ts���n�^�:�^_WȌ�hP��_�t���^�������+E2l�#Y�h&m;��21.ˁ�1{�����#���7��w9�D��ݗ ��	J��
��NX�\�e��/�%A^������${˨jσ��5���H��=87��<z.�c��uݳ��.�V#:dS:Q����Rž��'���W�ta�Jw�H�D��<�hτG̽G�N����P�n/���&C� y�y�tn��[���\&Q�4C-����z�:W���4���w�
��@�Ô�o54i�5��i2@�	�Nq%$fK��>�戈����zm�1�u�W_q!vǈ�����nF�*com@c��\�/Զ���*���:(��)�;�q7f#�DhAB���3��C=����BW]g�κ;��Ǆ�r_��L�G�W�*2�2�<����GDoN���R���-~%�b^5,H5�x�sc�To5�y����D�"&��?Lco���^��s#����m�?t��=�Sv�dk�L�C���A0����
��}�W��'�uO�7i�l���y�G;<�|U�1C�ǜ�rM�0�{�_	���#ɴ*o�&�����-r>��F�ӹr����c]�>Ә
u݁�cs�ˮ��3\'<�(��P骑�,O��!��Հ��cGe�$�Fs�˟Xh��zmT+��GRF�
m�����=L_�r�j���?>ꅇn-�c�[�ݑ�(�ۯ�FyK�q�/T#n�9�O"��Kn����u-D��M��������#&O9��h8�7�	3�ZQ��_f��b4D�7�c@- 9E`ĭH>;� ���-?��x/U'�E���FV�z����#��
��'�-������q��e�wA��4��,��{�W�%E�T�ԥ2,��=��+�F6������u�!4dh�-Od�h���x�%�,Af��V7Sx��#%�v�����z���Pյ�t�֖�SM�wCe3e�%�[dQ�g�jH5�4ݠ�9E%�P��_6�6мt��
�����T/l��_�D�- x\�ى���	����D�f�J� �9�r��(g��t��Yԗ�_�i��	��a�;�VX|�0Fq�n4`�w����}�Ϗ�$�}��{�6t����&�_Kp�����z�]�&���F?Lӕ��u_��[H �|�Y1�mb��Thg,��%(nK%���%�ip��ZsA6�z����5�#�}��RK���	u�����~�Ǫ1�d�6H9Y��4x*�?�}�G9�g�>��R�H��#}�@�ĶC��j��C��w�#����@0X�R2������X#z���w"����JESb�M��w����z�E���(�!�fB���(e���Sb�*��B+O?q�/�'\�p�a;L�"�T�����_�TK6���4�!�W?����; �2��O�&��\sXh�oӞ~��%=�P�jSB2VV5�*���"��p�c�Rh �]�Ґ@�uP}Y\T�����aۦ �.!�ڢAO�)��!�����룾�E&��ģ�囂��V帿�7b�����3J&�Ӑ����&�ɼ~# �j۪Il.���$�m�q��;C� �(��������U.���Bg �*r۰�FN���1��(Ҽ��4���j(�+�gr�qx�w�T�#��d�sN�|��D�µ�wjk�qNL