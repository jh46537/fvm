��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbж��ъ�]���ts�c�I�B[��>U����ܝ�N��Rɬb΂�b�`��VfR��w��clf�e�����7(���g$� IF�.�J
[�Gؔh�\��3��*��/���nu���Ũr��b�R�]R�Ė����{g�ϩ�(�`���N�Xb���މ����$fFʴ��@���#��0�)¹X7#R�5%1X&T&���ܟ!�gb7������_$���xD	DUDT����B?(DJ��k	ܶ)1	�}����f�*x!c�4��R�k�l�-#Ώ&���B���J�����7
��8 -���OIH��l���ogd������սH��hʱ��c����\�0���AfX`z�?�C�=�۰Q��}���1�鰒\j���.������Ż�Nƭ1i�	��	Vn[b������c,1��V >�TF��I��r����R�!8w�	�g�+y�`��̯s\�dW<�aL2��˦f�������Vkw�%5�q](v���G�N��Nf�	qb���"�!]��`,��$N�QQH�k$Q�8w�+=٤5l��ɽ0�d�f�`���ӫ�v��L�U)��C�s�'�c,'6���R��P�w�OE���m�Г��|�iQ���bX�-@a(��E*uv��������R�@��aZ
Be��ddN���l��D��E��$
[vv�j�U8G�6��i<2��.G��o�g���Q���+ ��n��㽙;��9������`��r���RJ6��θ�s�*�j�|��ӞV��ԣ�i/rl�'�����4�8Fm�ߪ�R�)2l��aȥ|���1�X�=!u{�{����:���8���o�u����1��O����۳S��{���OB%��|��Ԯ� 9�j�0A\
q��� p*L!��"�h5a�Ӳ�b�����P���{���BI�lY���p�<��*��t�����zD�+�W����_SGC ����|�iҒ�%e��A{�8�����@�7I]��P�*���Q���NVkQ\R7*I�'DY����PS�Smho	�'�}�$J-�01#/����ߕ8op�G*�ۅ1�����m9m�\�h/�ʲ+�F|�k)xX��.�w�=K����V�f54N�u�Sн�!0`w�1E2X16Yc����!fb�d���F#T9A'2U�: ��iw��F��R��6t�+G�A���H�v&��/d�8*CW�h�U���=-��FAk�`�IW/L�v5�%^���A5�j0*�Q�8٤,���/߱���Z�ҫ���؂�5gsk�O�4(O��hL�q��߹)�g�Sr%p���B�Vd�	�N�L˔���6M�aс�t�{N�߉�e~XJ��5��j�|�|� �Dh5���c��K�a��ܻ�))
mj 2��a�� ��"��J��Q����,������1���7O���:�<WB�;q�6��:��Wk�j��s��w�ǃU�i�p��oU�WHe?�:�0��/�vH�����{��h�G!�n�/	�,�t埍���ta�`[�w�/֛̔\f�=�6Lqj���´Y���Ԩ	׶Ś�f�Bh�
��l��OV��i?5I�1����/�A��k���j�$Փ���L{�x}���2l"��������lq�g�U��AUT���>���#Q��@�,�j���;|��{���	���O;�1�6����:�N:�۩�n��X�t��?�[�TL�������