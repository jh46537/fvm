// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fmSNhAvlzHvob5CKFYrmu6TnaaQ3WZvuJI/HlJTxOGw+21/t8K0y8ErpZ/Ts0r8k
0lbMdu/rPcnGeGavaxff9EhXIEprasEIfN41iMiD/L9JA6Zo9vBhWjh/LvRlP1V9
Zlghm9RY5LZmg06F+5P2QJ/LhgXCRQAqFMvbOsdZoiw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33792)
iUZp56VlGjOZpKNMuuYU5LO8WfPvZHZ/aAfcU71/yG+8qdXRW4dlW9de5oumlJJw
wg60pvvCv5L/5NCQMZKXx0h6cFs78c81gm1R5ySHZuH6glvOO+trstWLE7jGE3Qt
yjGVw3ifPmSZjUNSC58b7f3bphUxEnIMra+bRdKvacxZl+pUmxVVk2mRXAxMCh2b
tyXuYN84ln6ISt+m5AQGmbCozG6Sm1WMew44mkq5jFiSWWxnpga8dl0Vsqd24Eyu
QyfVzUeKQ9V2ZMdacWzCM0HP57ns1vJ74V5CaGPov9r0yM23by6V20tNUaZeEtGD
vj2svdC2ogwGR0BUnulVu9zKRh7q/C6KByvd3EyLwXUCz7o8jNApuC/HfSwwyZ8T
3f84MrhgUVazcx5EhXpUcB8EfDgVXAx+1+kGL0m023Os6fJ7XXx/fNCNK42nxp0L
3Qq+cr1nzfF8pyTcqXRhUTOTk5Ey9NWEWbGsv8PGPIvhBhQSnT3u7XmAPZDQ3EcG
br7MNbTZYNLbeas6PZe8jf93N8u5p2CBxANeuNk2NERKV+AOIbWezdrFvd33dy9+
5kecCCPY6zBlZh2eMW9oRNStju7oWCGi/ol56xGNP6nkUzt4Z1Qz4w9CLpwfhtU8
EATnIiqgIlvDzf8A1R+xwJYAD24wfLX66RN18jT80gHvdwl6Mm6xIKX4E+16Njup
yeCz/F823c3d7CthTrvkNxAO1Wn5ECVq5RFzp8FRxkak29/R7lkH10c9ZP/+CzdV
QGl8o2vG5qIh3G2KT2niDrsH+iOslen43gsZ2ZOziLvKtQhERJdJGOR+5SvJbden
e/hQp3Q0M9vKupgJpkZGF3hgPoyGRMgsd36pwC7h1xAIoNTlaJHeAGrV9Ql/r6Pz
erSJm0Uw0Nj8N/+ZqxpPB4vBiaoj3g2izuWwX7WYX1Z8o0xXw8HqnEr7LAC38Xdn
qQTZUvc+GHzB/6Ur3aFC96XuHEzX1Jf2AX+HLOLjo4mM+ipO4L81xDIt2FviKsXB
VqltN/SeOoWkz5YvKwT0EkC9kpQbqwGAtoNUaHX67KO1XnEbJDl57YnTRrUsgNjj
3ZclASyoJWA3uKWGKtKjkawPn/argWL5rmUzW32S+aK8PzailMSpxHdTcAO/wIS8
mFr74HnYi7c1u9keP5JenKlLYmHNQavOkYqQ32G7uDJfUkEWi5nrgana/d6q4oMR
qky59c+UY3lfAMO4lU3gPkuam07i2fDftIaV7pDq2Fj3Dd7ySM/EVBPPv0u1jCIb
nSsa0YzSsQc6TtXoNnROhTIP0MNt2t97aN4av8hemnOS9HBJjjaqyUvPt+izHGHV
IjWFRCOfDz2x5/DIOy+k9Y6/xyFwzLU2YwXGfIqxUdlBBQDLBNlTreybel6NW/yi
KWhkc7rjG0EZRFnLzf9usX2vTtgfo3qdNvgBoOmeWbEK2xCvZWpOYgCRCj3eyDu6
/fKwpK3goYQXPbynI1jzqBmvE4enD5JqLql1WQZzAyocCXReVEZEXuxp5TiZABcg
9Ls3wlp9p6y/HmHk35SJw5H8EzWCjpDtOV970NfFiQyoDEiFxh41njmLYFFbROfl
5/Mx4Yh6I10oGV80ct3q2LUn1c/p88SC48FrKk2jUTlzz313bqpYGX8HHJAksYqf
Pk9kBgGAMJsQvzzNJ89PnV3NERJIQEG5zcN2j34NXH4PLPVs9ad0xaYfFLtcXtM2
ykhBE2mOQeM59D0nX6xy+rKXuDxBWq6g8AyiIkFjLRtuWX3s1vBuz6C2fE9a/RHA
CNcel7BWcctpmJWg0JnKEYBH4vpLNbar171L9A4UbGz+eUbpZ+Cvcf+7KT0rKaWZ
p4AzuOTgyZWV0eaKZv8Qh9gtqooZ53ZQBqxV6JMPphs1j4u5saR78CEJC3cBUWFX
8Fb1rcu1OmvwQcEzqspvUi3XA0TAGA/Wx4/iBJC7SjIwpRbbJUDT16hamxRLZIYd
JEYmnfms4VSeB/bLA5vorvfXcmssHVkE/c4ro8K65dBCB8tlaPdxrWO4VGKqPd61
D4aE/9fr7RvE9JxnWJ7hXY8meAAAJvokfPBAoLNHjXYGxEuL6KqLJfuIiGEhmoZe
J5FyKpDTiVK36ciw6L0bvXAnGQ3Nt06jjbtIeL+7RBOLHSW82muOqLPf34FK5E86
rL/bFQsTK6TIWZ3Xy1IxkQ45SqRiLKMKMYMXUVXkpKbq9+6RlYiZcLMrR4UZltjQ
Jk+B0L8A3wkyAApJaq2iJIZe36/JCj6XqcEwPY/F77W+nRPZFIRF84uf4cZX2HXE
va/lP9LhTewKadOl2HU94L+tqG8dpZYhRd3VmaTg2OntUM0jhgf+e44NPH5YOBTl
H7Znk0ctR+K6Ya4lm0iGk8NoIrZ1DqtO7RLVigtY/4T7jkz3hO7QEw0Z+ABbEtd2
OP6B/RSGKneez3tQhtDnE8L8ePNPVptZYTZDpmsfVTJSJfzC9MR7CyM0YJWcNge+
plIeoXVVNtklh1he24g6F/G8nl8ZVLBMkWX+WdVP+z4TVtW82Q1gwfq1TPW/s7Di
cPnaB0wn1PRMrFj/6CdsmaqSmtA8OZJjpRQUFXDSJzcrCUWdP/IDQSReqdO2fMKl
WLZRiW7/MaMvccmtqNWp5bZn4unOGicXBDCjPv/0D1ERKnYH8we/C5MF8H48Ko1j
KVoG1UihYoc67XKZmCZYHwy0ppchaCZY7O1VNaE5ATTh7yj3RN5tfcNZsm2cy3gU
ns5Gv8jW6wfqh8QJY+zCgAKQodrHTRbC+146nRQwTSd6AO2Uycdc7wguQPlz+ToM
ZwjY0FTRd2SjyiBfiIAx0SJOo9kzxv++fSOwAgjzmswdBB9HKURnyjA26qjrg4/J
BPW9yoW/RxfS7pWM4Kg5XGc8pLv4H1B0BTQQCADAOsCDtpEhGgGNVacodpJRVO4R
byEeIRWIzBrAdz4KXCaE82Z5VJp8jn+P7Wxfs/K3seCv1o3XrHd5YAU8AtWwLggB
TnPzlAnHMGi/22a2SmWFxq5riIKc7ziaU8Bi2aXxHk+cZ3VVmp2bur0g6YmfxCdI
jzI39i9dAh1poDQ7sAL+qu5mk4mC9HaNW8CsAKC1wHWqXQ9R7/Y3pizNtHk7tetT
j12GCF8jLpz9lkCZ3M4tC+nTYQS2mWZa3mVdFL/1cYemyK1PtbUReC4rxBfrdnjm
9CAtB4IsWwoiMeNzI4lXw40N4F5MLjmCi4nTPaqla26E6rClpEmUbDl8eIWzfJrq
yYvACp1wqY71pqDXmZZzjSWX3+Nc7ee43UWRZIdMt/Sm3tTWDzD5hckJGLpntyDL
G4rKulpkRHVKF/nhUMcqRAid5kVcyMd610BSGcanVI9d35+XOBPad/hpBAfVbc4I
RY1zMagxyhlFRPkNLFe9sTsQPauIH6s5egNHMWcog/hRFaxxn3MK+XEDmmyd67Ms
u9LMzMVyFbwkwRGXIyN32GbBnQbSSODWjuVALPI/s4rsiK7ko2xF3O0wXboD+b39
IOxBB2udp9conLmRdPrX6bw7PnKqLgVGKMtoGOo4Hp1Upp7u4n18lzzkDgnzH8KT
x6tNh+IvRuYMDSlnGBJhocuNXN9ZhR4xELQHLvbcGmKJ3OcxITjBZfnl3tyj/Ya+
jHrZMMpBSkDCBkbuu6Kyj5RQxvGMaQTouk8uUNONLgoCFfcfLbu1YoOzhv9Qop3A
AWj8+4xaXivcj/EiemmWZ8vWyV6CZwwZvIR2VKFZW58J+mvKfScb5QGLPOU6eLkw
K+LvXLLSkzIVEu/RLtbV7YLN0RzRTYUlfojwpF5aQk8l4C5RwOccMjnMmtZLBsRt
dHcSrqiTLD2ZFXmQzLKZOUnxC5hnOUWboLYVq6Te65cutGBbfDvrmaL2MQfCTkHH
k3kqd9P1R1flTkycv+E+K3Yt3tyZ3kurRz0i9GlO0eI8hqClH+UED6TW0NsYfqT1
mSIhfSufS2LDpLhyFzcTDYfuQLaZ8rEwX2UIFH8aGcYr/5QQvklVv2ty/7N1wcRE
zg1MVSsU0BOXR6nuVvwhIrj3JKMvbNOShJ4Vey5XHXCYQSWU3I5Xlb4f2gb6kSvB
wMpuNw0T25DxBvbbqxIaUB2TPgwZAwk9imfbyPrcAaZZ20IC8xPhLtEfM2+Aw8dm
Lg3E13LPbjeKj16eekKa208YU3wM16VBKWOr59MCY5H4bnDqPdNEdZn0tx6sRej3
cO6BL8RfpmKvUEQQHjra6SZJw3RCv0esJ1XElZ4Ac7PZpjFzTZydYKPTf5uyWyS7
uuP1SQFFunZHWiBaK1e3qE0CDiZzfdXghaN6pLDy74edVRxboedFsx5eUni8yZxd
krmki44DgGGhu4xzzBvU4e8xVhrdUcp+2EU8qeRuSel/0EIEGRvXYghUWmT2GZ8X
SAAo12sF/09igWxG+S/GJLadwnV+DbrYYLgHJoqpDW6ykx84fmar2AMJRe/OjQHb
w5CzxbH8PQbgIoC7r6NnHH1X+LpZ0tjdn7+nmgBEPcKnP3y+6FNkehCIgRewkbUb
FaEwW01ZushNNvXJazCMAYOxmrJLkeYiFEmgSwS9XjSIqtRCzZUT7NeoBCgPQAJp
UV35oOhnHJPEuuRyipieW+ej/qAxNVuPnJlhjxXRyZwJE6BWQ59idgPgxqER9pDQ
AbAW2IAGXTfslUpyIQMbqQ1Q3cJbHNqSLLExayN8F5cOZe8KRCe/OFA8Y6KlSUYs
vvrVXwW0y98Sdi+WdPH8z8Pi5A+yetiY8f3+uD/6q8zvgYY4oGEOU/HC3oUiGhJ9
xnk6eyFEmE7aRtbjuQoV2JqZxPJjAKdCjCP2iVu6oYogXrh4Rzc6yK0bpdlrnRzJ
FjIAQi1+RxjI4+ndbJTJUhhzm9xJNTG26JAa6LBVi+KvzkD32tde+T3cloXG0l2B
uv7KOyd8Y6uctH5yDiHck7oqJ6e6OMfJyoEY7M2VKMJYyJh48tzuQtPIRWzuG/pq
QBpvcvJXQu6U7nZAPKHFIh6+QZL2qo63NtFlzcurN7M2degZU0+CHm0BeRIJqix6
OViN5TJRq/Bt+dCFxm4cFWu6cPeUgO8mA46WTLnTx1im0NGfMptT5J1Zu0vfscGZ
h5GMksBQQixzPF6UhJ3KR80ncI1FPVlR2kfIiKHXet2TU6QMwXArLqS1AdIMwV7Q
r6Fexd4nK72VPM00j+lceo0kfSSyrKWf3PCkDAXzRc4eJULCog/YfRas35c//jFx
XFCXbHEscKlbgzAl5gXX9Uq/JFMRKQDwjd+0bN63B3d8H9+jjYGEyLvzeiu1h+hC
h2N+HvXdacw2GHLnhmmRANLUyK8Eq1tbcedxYL1ZYUXjP9uO0xEuNT3Lv0UcgPS2
Yc9QYaIAeTr1lPtstRu4vYYEa0U5hb5h13kXAbJR9favbmaEgN7b/Jw3RSAe5unn
xgE+Raq6pyro5aDOFmSsf3ASmbDLHiWmqREIeOpxyaW7CxYt+cnQUhril3c0OYwF
QO2Hg7+ON4GHnLakXDOB5Tf7zf4g0dt8IQKMF4oBy3tz7pvJ2IPsBcX5GqvBVmyD
xfe5oyePyYXa16lFIfWxAPEZ0+/wH1nl9nMqTQHwsSYyq4BT6ponl7D3TjXKzlji
GUVdAni6FoRbfdBDqmFCf22KxJRCSO2o04CUC1P4jpOYOz4zyWJIDqp6/2Mbreop
ELMxDZundQObtBnzgS1ga8h3bETFYOAkd5lQYheh8QVfQKgklwY48txujThj97Zg
42UK/riJpOSscc6yh7+riBZRZoD6drPB6UU4y44c/uhIIkIdC84NWX/3wlfWzwAd
5ZNh40YdAOKXgsaqcpcKp+YblabDjMQh4FynG8Q7PI6aspeEaKDtIgX9jp4tjrBK
+1MCcM9ZMDjYhscpa3AHX11D1S89JccVkSs6yv3qB9jlJK0aSnvKdbSGL7m6cKcR
2TtDnsb9okZJk+KJaSpo6g24NY4kxhUXubTq1MVgMx7J6oDPX9zbLsrwKKHZR333
NOMUMAjNuzVe2jgDx12bd67Xps7HVoznHilRdmdWxSoMDmphBWzoeTT0TObZ3tsP
OVnD89ja+/XAfAEl41v4qEiXOb9Yw7wavLoR6qeShdN2UoeHglo47mTp0SFVMV+6
a+HWd181VBKkf8xZqVC19nVreZmfe1JcAK+nFKhmHmpS6y7fnPP0jc+Ij+++uvPC
0IFY4Q63HedAqrK6cbzr7acpdi3qeovyi8jDqmM5aq8ms29t0KRBiuYpdPt7QiVu
/IxlhZWVZA/lPTdqXCVMtY2z6PDlonjXLSUgJiaivVudGaGkQYUoig5GLNoWnRua
L5M+bjGg1CDsSirstBeRtXjMhFIXRU+KSVSX8RTGPX+idCRKfl8alQ1MjmxsnLuy
OWkNR8Ah+lgyOmUHIFNlPft4BIiA8Qms9y04XU6UymvhbifD1l/5VcY0Q1iXS7B7
wvgd0oNFsoj08yv4VDkan9bj0j5HSiGnqCM8YbASICVYNED+1I+CT8qVYbz1lMiT
5BGlWFh/A5erXE7/w1L+h23R7tHGa9e3GYSXLxI/57w82mM4FbDca1EqEa11yEF8
HUoozls+a/5WsIJxaMCHa16yMNhGCk7EFABM5k3tA3zA6ejome0ssOHd4BPg76YU
HfFVVaM40GfpqsHbVy4Y95ESRj+EXrYolT+PcvweB5rEtX24blWrLdzD7hRUbO+R
cFhjl3AE9qVFGB61Py5TQUnTJ0GFQiyfHte/OJ+UPkezUbKw/FVDWVT++RxkSQpl
yu4aLqqPFjydnWgAeSwfy2KTDXPX7z3XXA9nYXPYs+GfrqAwJzFguLAq7OtQSFVE
fOSq4PxSLFkXrbsX/Rjs5A05zPIMH1NLDi5/Q4ZN1sqEQZDZfbRhfoiafjqmtCds
ORp6zbekDjrEBrfiNFsvPI9TFA/sFKVGOV31vKPiroR1HKwdYU2bmfjFUh09WC6c
EeVLNYIqRz2eflRZAA5Hw/Js5HL0mRyZbIWzu+rpPhY227CDe9eDtaAITok2T78z
Kz+t/lhUI66prm4AFP2pFzKwm9XMhJ/6ztSUyeg2FrohP8fe5va88IwHMHrvXlKw
6h0z+6a2+9oQVScvGd3JDHjMIMglOVAEyNwhuYCQMAPpjStuIHBAoCrJBxUWz9Z/
9lhDrvvX2aVAlUPLquOJilwQ9jyf/dYo/3UbTvvDxzIbPaORI0ZPYzWnB/7r4pld
BohY5RxSDMIdayn8A3/9qM+t/9ao5YK43HkvTAohz5Eg1sE7Rp8I/57Eq6FeNohN
Q5K62N4WS7H2NmJKQhXp8DjQU43OF5RUxLFvHer8vwojFAfVAFR5JhHx8zuemZpV
6PKnSe84reIP8/CM0SI27j/cYzvdYCvzYcokhJl+taT2ZCvWzPK849xpAIXZwQ3K
v6msUVTm0NX0DlcVmnHaY/8aZRdOIi8rrij9ThGmGpcQamNqLbOUkSjhrtcRUJA8
o3VOKqLycF2M0lRvi8vT2tJFTYD0hJLDc15ecTQAcCSc38F/wEr9GMNOc8CjREXg
JsTPCIuOG3N/S6n0sRIQSEz6ZhMm7vLU7ivheMoqosKgUwAx4+ua24P6Hj3KhkJa
3IGgul3xs79DO9M+BE6L3M/j4IVvXz/ovkDV7j6j4mDouz5bQX40teC7ycuGJAZV
1vdCzSdB10m4szN/SbJRn1IuinrhVJMW3Xh97g5aIJnQmwwLIzmjhJiIxkeyGxDv
2ReXBt04rP+U9GTt8s605ED6miuKK0VtJVXuUQw6HIR6/lmOE0fhhJwHPQ2yXEA1
OSyfh+v+4xjR3sRCyILdk6zQv2cvxxdqj4xU+JgOWJoFIRj6LrJAFZ7rq9kShbxQ
xcFkbHG0h88eY7X/yFmiU9P1kojIXQSpsQHYAnn5dAtT/9chn5GTIMxblIAMsbNc
n1/SUnHhrh4QAAmLmlx9lIPjtSfAUOePUgOBrKIqv1nUzf9/G4nMcKQDhQSitJ/M
lmNbEd4gTkQJ1rT1XfeG423mJLmu/1HWuv5R4Uizkmk/Rlp1ATASq9LwzA37OJKy
URaP9Fopm/xTUxiJIxymi2GkZJx0biO9ozBAhOJ62OCd9e3geOGl8D83rtfXjhOC
ylcLhMFQOGZKEVRRpWVc8AQMCkVo9oQ9Ta//swmBZB7TxHcgvldnKtkWF1vs12Wt
TZQBy6I/IfAwnW+3a5N1l4o40HpvCnmnJ2QzbKI3Y5yu/92FHuEvTGIrQvqa4b91
Z8tfi7qXsV3j0BwDG6KVxlUktz6X9vsc0Ny0ihBpn6EV7LjkRVc3mXJOXbWtxVi9
IPzo+bwwkzxKgm8sRTwU/W4AXGASzzDqtAHks7C76ATxXdIkFnKFTwpl2Mace0Hr
XOlwvzrPgcC/ebw+RVaEcYGYFdWHACFNLmew7DPuDLXBk1LGtc86QCvaRvT7R/9S
p3QNv5nOAfpAiTCLClD1Kss73xkFRFUuh7xl+BucpmLibdNHAFz2vYvB63QOtMLm
yYjTxt9BAuNUzn4tSEb/5IrM+5Z0dH/lBAY1eL1WSv048rOBHrbw95xHQ93nLFoD
gh+iZdFix1kPkBUI27y5LUjAEgJ7A3kdocAn7oBWsCYZW48XvlmDYsCc8cfLS3zJ
X+X5ExIt8ozV/qWXA9+lGPKJ0KG1xupv9oqIqC8iXM9jARP2b3b2nwhuGXLptF+y
dy7+7C/M2UMw+5NZqIszZ5AN+8D5JW9eqmLuDb8yaFmj2ey570I1x13U884pGwHl
GaaDiY634jUtX1GA6zheg8fHq5uCUtKbCmc+psknUzJCWWyKKg+yv+9yPvrMFDYA
qYL2fnoM/Q4OFK2n0R1kue6YmiO9LmHPVXjz2djzk7jzm9KP/11bTNe14AZHAf6N
nXYwjle3w0u36Md8f6TWX0trSd/OU6kqetM+x97yWmwaAVoPtEFTPUVCjYuqzQeA
hPtQFBuvvrtDDL/8MJJ2Qj/JIAnZDj8pDpYZit6k7x3qC48k3ULpMJGWoLrOtxep
+NGlLw8ZVUUVlSR16exMgoRXqHuD0Mu7th4LryQU0NBzsWrpHikGMaAMguXpvNE3
TDpVgunPPSkUNaVhVYJW34bVaCMpeTDEaNTDQ49U/WK5hW9tpkQ7WmMuAkLjBh1U
79gvj3x/W2UQ6c041p2kDxzRgIqkksKkbE3s9NYBgZ2omDaWdvB5MPq639NBNMru
FIwsENSV8+Z3gIm5zj0dmkJn+UKUhwTwnSkNcp0h34j7FmSaKM+qjbt0XWIEnWfZ
IRVx48/BKOnOgGW39SyFo66kg7iM6jZAPNM6EUtyVaAkvJ4TDsy7G41g/nO6J4GK
Kb99pvpkL0kSbmnOvjyJt/CKFQbNkQtuk2p/YzIlyAUvBzpS+ew8gnYykauqd5To
lsH13i8+Tz7GWka5hx6Vy2nPjJCSfiGeoXisGqkQyjS7fhgIENGmdI7vgPrXHvrt
eDYZ0Ty8ubwqfivzLFbNJlFd8DeWo+OBgl8AfOhDGpangnqZEGdOwhEqqKUp0V1s
8EazVOUFXLrZzxBjScDFL5foK5cP7BA9/A2DIxVdCv15Kzizsn5M7Nrf++cLpgj2
H9X/4tbae34dDKUTCbrvQI7t3M3uzYwrzatfrUFctvrPPEwCkjglZmV2Lrz8+za1
tSeZYX9t/sXOR5P4m/RjjS24qW9O8BbKgwGupGtQwp4/6tVzDuf7VF1oNVo3RroJ
HPy8kcyw/BHcGqNCgF4hEZEc9MLxq3s6tTJ9b9HDnGXQls9CAEfybCW1FfJikZCO
STHv+zAKM6gd5kXjS7qT+jj28ZPF0az5coxQrTxM4a8sYGYoFKmEKgMYmLLKFA7L
fC2hY2fKCxrgKb25WmmkEhq+lawS4QUEu/kFb7V/CRiToEO4SM3e4mFFOnqLFbj7
hINkh28lxS/Y+acApZcPpbwLty4jnxP30Pcb6f/SFwweBvyJKPiccuTL+pE5WrCT
2b8rMfyupvrFSrJWO1CYgEbqT546JxoHN17pq/CBeFBSN8ra6AahK+2lGvigiQgC
ePnlgTMdsA39Mvjaw4ZmfBQU3RoRt3exXQyVDvlK5XTno+ceUkMinFHQkk7pvEc2
UsNWJCf/XlumZa+JtKyHq+U5kQo2oDixNV3WfH264F2FS6V3ZBxLr+3cgKSjvmeT
wOV8l67Rqf4ISuNoSHDJAtwZlT/i43uOT5uEZ1TFUSVI90XECHqVXImGKSrMABFC
ncBBZRih6t5qWCigorPVSwJeJ1K8GOvVnIaTVLfnsV1kPP+1mUNauBr4odlvkcrK
um9l6Fpe13hY7OCSJwmcMMujIGKtJPFdHnjyZ83QcE54sqKFJIUDgPlCqf13Mli1
TIA7kPI38axEm9Gxsh5SE7IHdh4HMaaXpdVy4D41mbKcWzT8yKqOTa+J961DZjJO
/FMt6+tf9ygRcmXWIzvn5a1Ry0nn8qfboNkN1uytQeNwirmvB2U1ws/sN8/MXJx+
vVl3PiPsz7SQuQ2nup6x/dLizdfK46OcCn5GfRq5Si291oDzjIXuPTIYl1edEKbR
Uz4YrWj1yXGyh9MwTJJ01kAL9rG3rZPeuyHbt8dwY5f660I5iSBFJOMqhZsSN79l
lTI+6XC9QZ1qhvnet+D4o9m24P8IysWlhS8THByVB0N71LfEWeD9KoBbjUI6PoDR
1uvAiie43eBFo/EYjGvfE1P4c7sY5nY7ldOiLexkoyTkv30kL3pbXHWhdcv/HPrJ
u3Ww7YwHrguQhvR2nks92bsmLW+ie2y2VTeFEcRFgq4CIJBuj42v75GluDdld48p
0v6QyaItOemQ0UAdz5J7A0/N8THRqmbTaBcow7BaYVdDqmu/qWoTvABQxWWYjWND
d/r96jGWqfIO8hO5O7ubiI+qBUbU0xdZC78HDcG2grsaIyeTe+Q/JmHQP9tgzIFJ
PchbKv0SoQ4Z0i4FPQweidZzJqKEOtk0bSC41sEAfMTtt3TUuD+6yWVBSzkxKzMZ
Uy+S9oRATfsosdaVmwpjEKxcwdgBVskXqXMrqQcrPTEhkFrE6KwYz/aGA35w/2II
A7nRjVy34Q1IeTkBod9AYfSD+kBhZnWbn/jNkzq6W0btCetbWjvP2vPyGvPdsDsy
Za6EWwrV2b7xosKQEzAbdmU3qfnKxLQzHsOv3fKS/NXlvdMr44pPp06RNUIWltbn
nqip3kcVInYNc163LhXZozdB6BEq5xFcz/u9Af+y7WJ8Szq1kw2P8AJF1b7FU7DM
jHqL3HYzFAQxuJyLNLcTgE9Ya9ZgzD63zprBHk0QWFrS/6mxn4sPJoTm1o5YjTU0
u8Gj6KSY6wowMIEnthgPKIKvJSDQV2prHZDxLLARm+gNogW48doaFvB6GY6FYuKk
kF1Yg41F4WSU8HFCqUAxcTQ20VPqTQrudmHCBIV3oXGshlSb6E05nuRNQLvMHqzI
yGBwHzeI71Fst3qIOh0FxHQR6ikVWaoGoCX9DOLc9xFRZjgb5ZKz/OMG4ooC66hI
+p/MFY/X3ZiCIgg7YqckrWkxoVVEWsbufGta3DnUiaIdmleiMSImej1WWt+0/NL2
eutRB2iUd2nQ49RatNoQuYWbZQiNrNXtxuPIImfNYviLZvWZFFs8902KiLoivMH1
/s1Y43lsaqSPDy+m3W8rdz4mpEQo8iyC1JPPJkfuscHB+U1v2nlzpSgCjmwlK6sk
aEGuwc2GB5G1d/0yIJhd5e9ONJT7cSDhtm97A964M9WCUDtlTR6PGIkoq00iBIwE
++osHuBp1eNSidbMcpPLqFDb/NaoQ8fcB2JRGv6hz99NQl9NEr1p31PxYVbqR443
3pf38CvBdxeGVoKWHAg50tWsSKIFfl1ismnHUaaiuDjQ+TziEfh+1tdSJnOUvM8k
fdvDqqkMeADjSUqAKzaFUv+oC/4WRFP6dBKyhNMEaHlWRPcVVRbWoGrwIaCR8AgT
QTNLFoUAAB8UK+L3Pd/RQ9335hDPVnpKuFo0NvoLg8e6tNsXJwimEjTP+Odhese5
gAqCGjEh+NkxFMgJwrArdXrhlnwKfpJ5KtxXFZop0xlU8Jo6a2qTulXBstoMYz0E
xZZwaQHnWgZJGdSLBMrKtDGRCW59hd3w190ixlgUzv4h2ZUbWQDagGS6ToB7+WPw
bHr7gdPqhc7wNjhYJoIcEGrO4jqjQ3GlofY4RDg4Xt6eZVwOMO/bXfX3TpIbegWZ
LzIqPqWM7bhWSAp2iO7mHTNG4LpLF/Lhke4JSAM8M8FmFSjxHqZWQWy1Wh2Fq4gM
pZTrYDYR3Y3u3O/n1IwQd5Nv+htPdfY1nRvP5ayU8m9O+fCdA/FJDEYBlHcVGrca
tLjNd1DCRQBvijmsF6dAceVUV3yPRb+BO2h/iUNAJkEpRfTTo/BQ6C6nSYTVX6lb
+Hw2QyTbFLl39P1nYG45XIe5WRaB2E/HkpCAICaDFRxQPIiyTbZjHw3vKVAhuyIF
U6K0BrNPTcvLBW9yMI1Rc80kvJUcV03iaCoHynV7g9DPjNpSP/RcWQtHuLquUWMB
n+waFqQCQEFbaOf/uHS7+1K9oN/HJHZvzRUQsqpVr9lblvX3CwfA18MJ2eqe+XqI
nEVcm0iPh+bTf0uhaF/b13BdH8yiRrfRn+ZWh4timDztJaB92zLal0z0Jdv/2bfF
9kczhmISV5pGj409jS6MCBj+Onu36ESYYOTZ0A82A6zIdP06wyTiNCtDOI9jclvH
mKl2keM8Myr23RjhNd4fCBgfC0RmCINDOJoOK2IsmytGzkOhPSjgNhrYejNCsZ76
av61R+PI37G2AiouXO1tT2UrT/PKrTVA9B8X4r5go4XT14b1PpD4ZJw9hIdBepkT
cmjbD7A4CJJw4wJrYTAZeysZlW6XTtaLNVDlVC2G4zVb4shG2y3bG3tSgfyQicnH
oh11hwJtq5gW6zfy78KUmNpFK3VX6CjzJAJwGNZ7P6M1Azf6aE+xAVRJOnw1k9kT
q0PcKUV8+GpKTCKIgPPP3xzPoxGQkX0LdPD2ZbmZTncF+OcOjL5Y6KZZyC8GKe9A
n/HjjJWNKPxXUAJ1KoIWTAnBcPNCheODATGqmoGIpWrHGYT1rMCnJ+3Z7wDOpJlg
2pQEzJ+JXUl9KIMHusX2wscW6G8pg8WsxhgaDicwCAGTERSgOniZvGgVf7oUCaKj
2Zu8ITcLrUcyKwyFMoNdcDNAoZgOeM9Vz+QQGBgjEMgIxKMeSxo7H1fDaeijB5uj
6RWs08e56M9rsNUBBRzrBXWPoIWra+B5wK1hDbCpE1mPxcEMI7PCyyL1aB5O9FqZ
eNFA/bJu0frUXO3SFNbQaPy2VkJW8BwNt3Q3RwzpVIhK1HqyzHYdI5wyldbn4rF5
Qk2kv43BjcMZlxRda2bLbS0J9smN2uFCFbsshAnfIaKDJkJ7Ggkriqda9eRs84wE
BFNKS1vgeUsKUuZzwcZw9usawK6HR0sshOEVspzhe4ESHPyi3wguz3FzihEWRHX0
FtVuRzAGt6fxS4WduRcKjudihf0PaGCzL5wVkXDuEdGokS8GjeU3l+vXMFZAUBTZ
9cuDEMa/cpJmyl5o2wrBWJBMGMH9sNYn0E8cty8tfTQPOijTUsuTLMS7spGBIyxo
6sWvXhrs1zqFf5kgJ5l1co4HFbI8Db3MoI0/9+E4CjGDJPS23kbrD5SbnFLoVweV
GQ2mEXjc38eU+Fqckz8G4JeYVd1+3BSl5SW+vrzn4u7l+qp8MjdPme3x93RD05AU
TcvXrHq/Hz29hKMbnkEcy6SxHAsKwO9+Cz/b5eTwKbke8zpkGC8zOqtGQENDbc6z
bUY5pSwTap7XnCu7Tk2kaoPYSZcZHw0SsWZ3glymDjOTUXEq6PMG6RuDTI/X22nt
4Dc4nBQJr5l4b8hQqnBGTG6pyu+aYrUwFhocOOWZrocylCCpJN3S4bNY1UG6VJHQ
sLJUCF6arZ9MD0QP0qtKj1q7KbQC9NVNPUVe6Kiv0/ltdS5qCWF4P2T2Mo1LUJDS
l9sZ+a2X0PWaK03okeAMTZNx6Nu5bNvgZAlqZXZLGeZyA+QvaG639+3CVWTOsdVh
7mnugK6LKXmuNXuRtBi8VjTF2tprfHv/2+8+pDI3WlkiSRSlIcuIRLK6z23MoO3T
jpESiEcF13OHLQFK9OJ1AUzBdf3WU/+Lq9CEutoSA/NALJrLgucz4/Xt+YVz4lOW
VQHtKghf9YeKWVKnMTKdfguqRaEf6e0bHwZ14tLOtPkrlc3tmG4CuA1W56zIgfOZ
4QOOfTHs2V7uSdMQCMHowlr0n0GrOiwNcAh9VtMO/Hl0FgsQMCAhl7fqvZdfo/G4
WG93Wyz5THBQgiYmRusUs14sI4jgZHU4AmPGcu0b5ervj/wkkeUtpW9dB2nUgkKi
9UO0UXPnE/P4ZDuvWFI8pY6kIx+ESFU++4flS2XIxlSELeFm/de+DgcoHbUJ9FMh
BVmAmGXrbV8PhXb7cVhC6rWI5YYTRQ1/YcgkBz5EJMZWRPgABq6kINhM4CLE2/+1
W+cQI/rTzanz7zV8nE3orS+M6kb28plJziB1Slvb0Sl3fN59r/KWtCiY4P5D/hLO
HsuQa+PXNLsZiWwAcjEpGkJy3830FYSkazDEbZXVliJvOjOeWasLKLmRHfW3NQM2
xNOF/ewpqVWlE0nTOs48yyl28HjEQeeDQMXpF/+3MWEDL/RoE/r1oRYi9saMh7kN
x/J0+ORsqcwQeXON299lOEi6WEecqUJJi4AAgevimTYbSracaDfI30PNGoyaH0oc
PEjlMhb3KHwslzLd9vuV+IEGoB4p/sfSjJk+yHVz2dW7Md4zBXmRihSo7IXY116u
pB3haAi+WMeex0MljhnLKzg5QTWFX3MvW8oXYp4EyFFPY5Wb9qX+/uqiRj02JJ61
lczQy8bThWTkRh506FWcXWfamzm2vgnzzGz760PHV/nN9dkhj/pYuTXO/qQ5+sxy
5zfJnpfCwx8sr0WsmyThQFp50BZYfsW8DkFsVKdXolX0KHVvgol2ekZ6YPE8aOxY
zMtbxRYtk0a7JxWE76At2gHyDHXjQYxS5wJnqc5jbuzV8EE80g2aq4Llcmr1OKu/
9vd/0IsYJuOjDqIdE8e5FBEaf06wj2N2wWLpLe0zPPKPRuFHqowXK9k/ayptQjoS
GjrHGApc3tZRYm6XaiHYi9I+b3CClCGzdh7Bb7umxQMW1afarzJKMiA69jUaH+D/
Nd9/PCxqjH+JDqtL/wNM4FdyyBf44DEuMbab50JV2w27dSoHQLkpoXyWNCDXPF1E
Jczol+HSP0vSC40poX0njk5cUMlIjjP9XaVNh5rOxuQJ6RbR9Bjt14EDo7c77cBq
+CbtJQEAzmLs4frAvxKd1Zh1NNGOPPRYwuFEj0vKJXrC4+B+WFzNPjUk+XnXaZZ8
kDJoopoqw4PVoDdA3rKwbKyRqMgkrmYhYV/47K4fwOhVYfurrSgitoP5O4Ec85he
qB2zquCzQbrmNuTc1B8sLuQGFxvecJnBxaFes2p3OIJCn9X/Kumb9u7CzdB2Ato6
bC3ZSNOZpSVQ/llrJhq9V+x7iDFfmmYmaqNzpirZcyTE/2jH5DASV8fsEYLTL8W9
VKsbYCnyhHaNtp4NBYA/FUhqGJ4TjRSB6CvTDmHLtayfcen1VgOsAeMPSd3m9URo
Hbx3G0IITGrFfbIYgGZ17h6mu8qufOzlOirQ+S07Mn+ARBjKl3fWjKRaVY5qcdbe
2Dj/fXcrJkf8OwQWuARH3XUZxY+UA8m+f82fk07Xp+4BLzXn939PCVe8iXK17jC3
hmgsYeMbiq+FndBLS74mcZ+nYCh+xmiD8FgiNHnztLpUp1rzR6Brc9oWpZjENRWI
2zB01X+O2M47HXPe2GUD1O/UWE8cCpL+cXn2s62Cp7BEmX5HatBgMqcBst31+BXJ
0pocqrmAgwiekLAyng74KXV5C4MnKo4LtZjYHLJI0T/VnHba+G0hJ4W2u85lLHEx
fA8cW9bw4ZRZUG/frUUqWwHUCGYSKwhF2dvVY+wEkjyZ7py42Imc63F+C6Y/uq7R
G6QzvXjD4PN6zbyed+yqQaHb4OKdi3ttCDp9eBufO/5UKrzos7kmQu2GjXWYNfwf
fdAtk0EutqlIVipyEIBMiJ9BiXrlF/du9pX7QeAKZwee/P9wP2CDSFCfYiRfAoCS
OZrcMPkhGZGHYfQ4xUanUTfcuJh6TcC3ryZcjp5LIYHupu/9rvjmf3d0dFfF37mW
2g3nfG9XiffYN/LQviZUDN6r7Om0cUG0DX/DWqkqgwlpBYc96Fm/0ht8UY5YxQ4u
BKzYbnRh1tsrb7if6tUWDJ3ltnE4QowexLdbxIA6zh8etopFQy0EpUkQJBYcqdgW
R0CHbigoQKtl6s+M6O57rglaajoUNyVUiyvwqU3TwrnBSX4cHP4Tzo3IqcjLtKB7
S685tZG2CQMMjKScB4IItu1TgwIK22gGOGdvg9i1c8sniyOenK3W5jzQFRM19cKU
Jay8RYmcit+JnhMV399ZIklAaHZSFKy75UQ4lC6OLZP5faR+RYfllCv765TubqIi
ZxrwIBDHanaDnGhVwm/Psdg3s0ojG4uAG4mxc6B16EaCcGrP4np04z9thyLcp5Yo
AIrbatu02m8nkttr/ZFDbBuPbs5TVjy+m7yJgB8pyE1sTBwmMUSWjC1TD5xSxWff
LX0OsWt+BhRuLecowkThs/EGFRWyzSoZlpdGf0ZOtRSxt1ck5jwYG/GTsqxZ/1Kn
T44pDxqXUD9RaNiNRGUr9dhpvJ8m0RvJEKAczGo+c7B+ptevkPiWz0zRAyEsHXfj
/XasdiY1iETGd56WR9G7dRcvD1V2Lm921W/B4dBcAwoFwZx2h/SszV3udLxEEQHw
db//PkLjjL28OXw9RME4KEZZ3VrT2+LXfO/+5ci94TDYHlFy8iarUOQcIYln3UJo
/TxIuhSOPb4ha7E0qJ9QOTsUhQYIb6HNvfjkTaPyztVDr3AUhqiQSeaRkGZeYg3B
1QleI/ipOF7n1wHcPwo1GS032i9iovdI9lCB5MClVEIEZEW+CIqqFlFGG9lJaqWI
68IXm6oKRcJLncxFHbgF5bsxSAwzjA5bRvHZoMujvGwsC6VpvUOwcyEz6geUSGu/
vruM1NzptOq/+qnV0X+e64EKDpxn/TGDNjm5ft5vpX5+0Jpl39zcZ4pMpsc/CJdZ
DL7vGq37p6N3YT2sb7RN4pSOqprikebwgJuV0S5rDugcrFK3zUhOjf6ZFSZlWHW6
iLYoppAZB825kP2XMuqqZ8opE0ZlKF7Zzc3ZnSRx9aBGWRjwedF7rS7rEPJuszH+
uB/zo94neSAkMPSlxb46ekXRfnc03WYNsojLdiJhB16lFk7PodwnU2GTvtc196om
qf6jPsPQWJ7OMTM3u41Bg5//yBsb/1h1Y2Yi1gDOuvDrmiC/RBicfMyC+yURT5P4
lUQxYNQSRqiwvoVGdkwHOiA7UJ4uVf6mZDoI4KABISx9iwW87ra0E1Sk8yjCX6BP
8eD0pmvwgEcS9eRSieNqgFJdqhrHaS38ztmsjzKqH/pm6GA/rbXISHz7r0MwurPm
RGgVoNvtDJG+FQyJE3lzd7LXSEcPxNr+iSWU48vvDrkWGSGS4MYsBWcOVfjaVsAx
uyrJ1KU45pxlhX71G8E6Xa3kvOXnubmiVqeqeMmr8DxnJ/ZY2iUT995tVe9tPksN
A7QmcDFn5cOOX1CfYwAbgWeMHtwGuQ0RcaPWgqYBzTPeCbRqYPJti2LK//mc0aRv
zI5h94cpOyulw1kTpLowj3OXs6FVLPmiVpcBo3eSVOkWhrBelW8L5r3MEuhVTX2E
RGX8LL14bOjKggASpXVCEJipJR5vVXxQZmDbkU8TgC8DPMVzZHeqg1ddjCCHsAcp
xZROFA3gI2P7EMySWQqdEzIzOE8/a+ov1eguBSP2fWDbQ/MX00VWR5XdS4VebaI4
EyHSdZKC6hd7YqplWnwY4j8E94dYl0+awY3iJxC9OueBAHqbXNQvq0iOVoJDkqJJ
w37CcHJYxzcMaSJt5qDNIy7zvnTFSClPwrSPaoHV+TbSgGSN+NwXqdXJ26PNvQqR
W6hvcgbaJvTKPykk+1edLQ0xe7mMfonirot2nWkowFvH3YWTSY8haLDqThNBu8Nv
9SwExe0Gz8hzQDu4T22o8Dfo9Vyp/sTKUKDOXgirpvlSkNOL+e01/rgU5R3qoqqI
UflWx42mDcJH89ime0Byci5Ykepi2NKuRSyAnE6rEEkICvhwFv6vFOOwPEVcCDOB
64Y+7eFNEd3NOgHwittdzv5PyueBSJEbj3wtaRwggqqkcXxrTxqsIvMVYAbmDwtU
Pxqkq0NcvG/6z1BLA3bC5hQ4uJEmDFoKc9K4gM+D4oGah4hAb23Xpd+lFdBiWcPD
QxG1tJbGrMPDJoT7axZJKvnxcBnkyLFviaeqJ1b33nK5bxx9dkzd343vpQjtPRef
pOqjTJnzw48D4FUAHxdZ3yOQ1cNNzRnATo8+ei8F/AoIlXy+kt4UFJBQgMH5vEP4
OM8c3DtmsKWkNbsOr/UkJRfDG76nZKmhQKitzAb9+/B7USUA5dPo2RAIm3dGUZcF
Pbn4toInp9K/bpUkFbfxipyipG0YnohxaMa/4Ocomy6UGS2nhS4ba5D9lCJE0tX9
k4M6/ltoXiBpDRcfId35jZc8kW/mrxstccHtSYZtOMv0M4GuDBwraj4iYmPXBVl2
5iELIIHPLLG7nJt2BJeN2G30peMPEKSsfkvtmI14n2APqYbElezbYJDLIYeCqiYm
FSNwN+iVCxd847dMXx1ECkHKSIluT9XqS1FInMETrg4NWzA48OU8YqTXzPtyPr92
2JqCtXylrZcHtagUhRrRM4P94ybr5idHUgdfJONuEBRhE82IFCi5GvAqU8kiaeqv
ywJt+Fuyldv7E0OPkRcpKUhVYX1TgIIaTptw40Ebm9fgb0gXZNURsPVDfZ2HHXg2
xVve9NWSopaC7C4kX//30Z4lgj+HPvwoH9R5JyqUlS0ChDeMkWsU6hD8y099MACz
hm3XLSL91q8ebd8bk7nTsiZO84qCGIL0mE5xJdr+mHv80k8MmoTUzyIieCx/GhIN
nrB8Eo/TK6qLgSqHmW8d3v84cxtfZGC0DCqG+d5IJRxkgECcykM2SGFKobflbbCl
j8cwLsDjfNkQK7lIpHt7C4AgFMcRMrLyyljX81phSmd9I959K5nhOwybjf7tgFO7
Ode8puTRfnkDAd3kmzESEadtwEaor9ejDh1FiEL6Qmfa8f4dSyzZDE6Gzz/upbei
hg1HZeZY9xwsQuC5wbTo2fdWeYOrAiVD6FgBPJSqY9U6DJlwMbmrNxKXhpk2bNw/
xavxwY3YMrrGcoTa7VeA633agKVdTJVZTP82PTDKwk/N/LiB8zldSFmTvVo3oRHo
g/nYSkSw0ziifmNSqSXcLLMHi0knMg2dVVy0/tnPe3zTfn0gaV2Q7E61sZdZVxU7
E1T+hmFr5SjKRJk4yNos9pFBZg6juC9jz+LGYthoQMNhuiPFdj0OZ6weLOK5CaE7
I6rpUXWbMVQImyIhZf0QUUNUSGVpk9QvI37txlhvrn5SSsksgVDjxHUsyNVe/sBF
qdZ+0b61WRh3XQ1vbg/HHQzbLrrNS8nRSPFCmj43nvqWTpdJV6H5tpkNQcI+4/31
adXy9iNR+VuyAcBJuDVUbHbE3b8xgzSnxP4Oz7bT2u+Om0oyP6e924BrfDLayYBq
0azH+QLKnaTJknZxn+UPn3N5SJj+Kvol6iypo+mhdywbIuViBHnAYJ8guyl8LdN2
Q0aYoqEZwPu7ab+1qSVv5uA4jjkX3vpR9O3sA1tsMumeXoeJdfelBOPGhK05f0Yb
Hzj0kod7+SV2yTFChBEcCVqtNNN5zgV275P20NhEgJbW1Cl5vWId6xtL0pSsHoN5
0uvZeNLuLZrhW5r/x0qOaw6zn//cURcJBuq6efEeaOH7sUBC6vER54uSOMSBSaHn
tjo/tO0zuezYgRZ5/u/zArPQAE8v9BrYW5jpSZnA+m55qWYMnLL+0LA6U+wbX5rh
5pZu57Lo3apMAB6sWlcnrpyNm+1xldn3okrQE9o5zQE6ixNCIRvIpP3Ix0+26D++
aKFbtTU+lenWj625VPoC81NTVqtnncM+4TsEq/xHvXoODSc6yMlwIflgajiASPYr
m7Y1QBjk5Mxyc5VXDSSB1XAq334hVb8Z7dv+ZO987VpkXLlzP00lWGT5T1+H7U9H
AhxtKX7f4R0j7EEMLOJcROBHDWvEqp4hkykEJamu9vNy7aUJ0HEOKdaBJa/gMwZX
9jGUMKjLq2jgYKjtUydwaq9OdCdngDkTA5MRqEW4/lwSArofFQgUp/d8s0/o0xO+
rkWiOMQypM/RaAZ6hW09/fw3UmL9TpRPrrgaOapYxvQ9HcrrsC1kPMltXNJnKWl3
hAe57HvBEODCKgK4hOTt+u9evK4YmOCxphdThf0z9Dm58TkQ894bLA5VAPmbC5DE
tAi1Oe4nALVLq7Im00/4CgbztG0AoaZRvnej7P8MRblhC6jAWiW2Y1r/g3LV8Jzc
/6So/kuXzet0Ch70LeNLsvMFTZ/+U7yBCpj/0uUits5CwSUhHzWk/R+Uf8GSwWbQ
42YiEhx0mnazxEtx+MYfY6kl+/2kIfVU2VbHKmmeg8ALo7YmyEe+k0/rSCrUhzHp
11wO6xran95TNetclWBJh3/J3fARDvQBBk8AvcK8UMWWjteRR6MRF82rIQr0JPEc
wtjOmwJRwHS1vgxfC/yDBOmhcI46KXMic9EaEBPU4aAiyYioY5ztafMv7+rApglU
7Rk0uJOnbdGXO0n7ILZoY7tnfxAi5YrIUjVbfYF55QzpMCbw1JtIxUvSuu0CqIcR
cidOCWsZl3f5AMePMu7iFhZ9huQMeKO2/PO3T1jdFeSHmG8Rx+37J08bHZdvsk3K
mtVtqI2qy39eARdflD1Gw2fHcU5PQ8tWtXMdCuYzovdh5dwVerJSVW2NCl1Juee2
3wPJN4sjpnMyhZiY5UpMAUYuG15Qy0zCoyzsDpPdFj+Ab8QdSCHC3RBsSs604ULR
0/02JY5xoNyUahIsqf6MmY4ez7hA1a75BejqqUu3G0nu50jvQMDRb5pDASBY0oSV
4X1gpmPcDDubUnwo0B11sJQV6GScp88aqVAWyRS7gR7XxUlUZEDobkkGgyCumY4H
bbonYYgta0LvnSOJ1arfTuAc2uz7EuFbnEKZeQCoZ24IVYR4rsrCWXUqtd1JH4yw
rcQbWCMfI+h2r9ejzDfz2ACiyaN8xJd8wnliRv80+6weilEfdbMVhM55LHSAN2pt
MQIPZBGhQlGm4feSWOhv8gntVy5BlPd3j9DlTPbiAr7eCxD7JBUjV3AjO1tilUqj
DN4K8A+FwKVsUZRG9f5BpLtkaITOp3J58zDGt3acK3UTlDvim3LheOB7e+739ooP
7qP6DWX5hU3AOsYybDI/izwIDNQYRZDDoFPb2YJOLDGG0YOFuTmS8jNeWs3bWrNq
vFjxsnz8VwwFR+ko4ehqQH4f6atgNjPmL1OVftfyI+comwhKhQXLaQnxiIpyneze
FNBdoYtR5JtAkkHi7P/b7t4tdTqzW0prwvCXXZMoDaBtDgLEGmt0QmxAvIAM/z1l
JYGr064830UtsuHHNa6E0bXKzqVAzjfQRBC8syG7WqChJ7w9Hi6LWzqxUAzLh+C9
Y8qNAqyZSVs+JLH5rmuHuOdroNbCSrR0VUaF3pVY8IKKaeWJd7BuKliY7meVZbc3
MGYDTJgf7n4Sy54Y159TU6JPNkBslKLqD4+XDYco4IZNFY+5NPnF4N7/d63Z0Vd9
9MR3VrCad0HlACxHs6kFQxwz79lPcmv6WLbuoEs7meCWpPS+Ecp6Ph/mPSfB7cNz
EbwBm3PzqRmP+mrKgKMj2mpPHQ2XwY6ucADCaIMoik61AqKffIQq5y8DoxkAD4zt
Dh9LqF3N0fSTZWRCBzIhQaxslOmcXDtDW/CMEOtcSePkwAXHlZ/rFWi1sPuS81vI
SEaxdErpkUJqd5bPjlkAHzcGlvWPUeV8zdwhIOmaDdls7VfM0jW4L6XKwwz5Voyj
ZVdgQamqv/OUxQh4s6QH63QjF8v1gNC+c+WpWApdSx+pd+ITPc/NoRFif5iEeGtt
5D9SdZMM/yKsJ/0F61FUACmqWmvoOd5aI5bHJ37rmB+ntb5nWVPr4/Nzy2NYUaPK
LmRxcItAfslGL1zDEAtjRbMnaz3iI8i9Vf9OwbqCnBMX6VrDaNP+ZKPKZRVnwZYM
K3Y+Obn4p828L2WIwnodZuLE9u9oz4j6yYIH+AGE1tGpZOYmrhbHeLcevS5c2imE
1eioufszNce1ObIndGbbYAXP57kBvzsL6BPV8wFqBThOj/A3U9BH48eZ4L+WUoHo
6VybJpUpyMuSeQNO2s1vdFqz+ZUyW/EKIQ8uGXGbuvNkNzkmhga8lp7AJXOxAOdb
0vjCZUU1hCML6RzrUfQY8jgTEyT+Y2IocF9+plyBP4piUDEdjFUkrK40MF0ZmiLI
jdjwf3mWe2h5qoLsn6aFF+bppUR7XDd+qZCr865hKFaZVZUuf+OrdXMmqDwwyWyk
knqrxsk6EwosYm/gHRDxXFt/84i1U7kFSgiSW3NrjQpIhHibXkWGNZJS3xELU6mF
1TcitNLEri4k+/E91WjY+BVGfv5+Vf9nKv6xDY833aqlzIzW3FupGgYLv9mvCcOa
5q2YAWIfup7q1lr7V737JhUZe1QzdMnfo9SS+7utnIb/9MJJvBmZSwQWKW+EpMxK
ULE+xhY0SZS8f/SfVF2akpSRoqNFwe+Go36QyzAFaZIO1jfW7T+VmRe9SoTifq4u
Dbxz5UWE6Ob+CvKsu98iVbfcFGg5a+jl/gRnusoSSyDuB8hRdwue/BaE4+vlCiT3
AhTVwfhz+r8DCDPYCfN50ji3LCBygXCxSz5JOLuc34hoamGgKqatIZreAio+gpPF
QUWTipoDGRV+GgL06G46M7bCt27ibbS6D+m+LifjFMweI4OFgXt6VmRSEK4psdUG
gZxlU7dpEh5oJuBYNjqZ7iv6ypA/r3g1elZoqTsi7YZNes+bBcwRG0p5PJAr8JAX
kCp2/MjRQ70ilFVd/eWV5gF2ZPsnZgxqRqx3WfBw6zxaytfTY2oStgk94e6tA+29
PBAz2uSbZ4kCosBmMOIz2S0pyg/B7QaDz2oytQuFwW81qRNpr3mJLm+YwUO7bxUF
dXGVh6z2pcGYvoheXpQObyxJb3um78VrJY5sGQyWXwSWohk/KeaA0IfEQc+HahgP
HFtR64gBYweEBy7TIIXr1lfTw9voHUmOG9yfwm5y6aP1fE+k8ZfL6NKdVnDZbo6z
w50iVS193iTdN9Unb5qEFuB+W+7yqwr3S+98QH0pDdTw9sNn6STLxlQb6Kc8t0L/
ZhLmVZvtuoKIwVDJ39haQjgSTrU+s3Qf7aiSdBluiD/HZvlaYR6S+Cukv1CZCuQz
duEqszT7sLs59Yc+wVfpyTqlP//UVebDncQIqlhDG2MIanlr1haZAMeV+nQKRyjO
mKk8y6C51KTPABxCuSdK8l7OeJm9FdXHb8ZDa5VbRrhOICAgu+gljuffk1eX2+Hu
Rv2ncOY5JKBrh2ja/DZc2tYaqLES2CrV31cJM4iov9BRMQbNsJla0ZeM/9e1GJsE
1xy2WWOOg792ccl87x6RD5CVWQj1r2bBOSX4mz1cChoQO/cYo+ARA/WRe1OjG4SV
5TYOyfUbXg8lyuvwX3F4Anu6fzaR2tsNnhtfcOIEJmBIIu3ZqMfs8GcTmGLlnRcz
QPByRQda71jv3SeqIG8kCS7qjES8ajN1eoyiJ4iaCb8RM3CqDkjFw/fEyfq0Bn8G
oQ9Q7zC6b4pOxXsD2YyeBoT1eW+5MqsheWAdRGc6M6WK7Hjj+4Jrz7RwLwzT7jwk
oF3WzYCV+PtzJXhi4h305YmXMqBMAvOdJ0yB+2IM19A+AB9dfO8mOezQkmsc+kor
571kM12A9SvUNcqM5m+Bjh6cLGdQ+0UFnvdQS16pabc7/j+loVtjK9tCo6dBzezO
tNvgXv9E04pEh9Ahq5rdzK8Xr01vQ7YCm98gHAJC2/nnsCof4a17MXmoWgxiezMM
Z05nnzCvHf8Te6GbcOpT7JufmwG1CX9cFY04TcCcDdUIH4xcClRkvSG1P2yu+NlU
TbwJ9x5pMY6uquwukakWhZkD2Zy0IJ+3bc6WxpzBXcvw6SeGX4zUus1l/zuKpFTJ
e8Cam4Nq75OSZx9oc5FxUCZdzDbzjJH09d2Fl7mG9cDlphbrpkPJ8xZZl4llMmNh
zZAaxEshSmd+y/7zlf9ZTYpAAsj5ZBEVeeob8DVL8uJqzGGDe06FA39GOyr35FED
9LW38YbPv2BjMeOXwxaVlmvhELkgh36wr1eLICDA3iREQiZCfFZmH0kyHt7BFKu1
uF8gWhYlgtlLR//wigKJ8kr4vmS3h6rhqO8uLV0EZ8wzXTNJcgZg+45cbwDDcyG+
VIB4IBNidQ63pZel7aDXoC+JJqxO3vnCkBD4HlfBpztTRBtCMo2fhfwR9BSF/Lt6
jA02mP69ZdAFTjr6UGG2w76ErLjF/tK6raEV8wsH8M6Ztw/DwtuH3pm+pc1S6Y51
8AFNgFPtauti4a1g3YJ8FgfM1Z0GtBQ97to8Es4qngXXpxf4avvwdj45yUfNRBaH
UUdpjvKfhqSCtuNmj7R4nRyygHkJTg0jaCnhW1UI01qMZsw6yx4HWLXTmRGNe591
TD79aeTAYrgjmqcVIZXrdX+PHDqNQ6pryq0LTTtYH21xktGngKobCEq6U9O2DP0C
PoUxkEi75YBtGTobt7FUIAsrWI7AX4TzY17MXhR+dRGCCnfKBlqir58V+GdLx8FZ
fU2lBwXjr5eApg6zsQgQZPZy4wOiN/079SOYPnJr0hw0dd8sbBczRTkto6eBy16o
JAs1sktb5rLvExFn9v2PZUuh8dO6qjJMgXY8ZJ78s6pXADNJJoKZaGaj63YnEHVH
HJ96iYTYKHP2U+ummXem4YveBoZ0ymBPgojPOtpKlKyIt+ybEVFbFQeJa2ihi6uF
0Xxc4PjYacNicdOn1eNmEo0MwGfR+bWrXWyGGC441WoZAqVlO6tGye0yUtm0Ldgr
2EKdVW6fVRxKkuK0b/kaCfZoEkwhUMG5HMvsm+Kt02FQRQIyS0OI1V1OPmWNVEcH
OSk67A7OHviezLdJAL4S9JxaIEZvXH6Xshd1PDAl3y6Ge4Lmv32Q/wx5w2WX5lJM
BR5TUuXqBMCxVM6vzPggC9bXtQr1BoGAGtqocbT0J27qV28RPUcPJmY0vhXaanD6
7BkpmRzEJ8byLcY6qMn/KLa8x04KMRWtTAg/qPq11+wtLhJ7udFK6sUe79iwT3/0
th+xMJppaqnWmKo8i53d3EJpuICtN/+w+t6gQRLqMKEhAjTAEQdR6i88JGaCIOSU
fal6xv3WW1Iv27dolpWGtb2Z148MwnzRrt8xvrzoeaJMdPPl3bog4fMgsu0d97ls
Dtu9DGsGoJIJI/Ipx79/RKuMvK1qBI1dFuv9ddJRV8q29lO/BbChTKdNWPohpX9h
zMqeGIa0mZSFKd7bYH9UQBCMVTjAqOKBzQoPyJsn5Vcn7jfHTI+AExiZbkFfxARp
rBunp1SEpHxizu2kgr3icaKcSKnIj0F/11fncoitLz5Rl7G7SCs0rRnWOp2ZgD5M
IArcyP2A43DY3rTWTq5dIOHMtjEHkPRamGyY8/ax373b+f12GlK+OvQFulpocOaw
x+fNONvEyYF/7Dy9Gw8EhUD+5Fc6pVAplbccXkE7W8HWml1E6B3n3johoY72QXwH
LHLYsh7da5PrJdpqMevYrAY3h01Jnr62dDG+Y/vUjaaqyKSn5Z/84sG2tKdjggPO
4j7/r17MQnpzc86/Oj+qQcA2W8VvJRJy8/rbjPmxtaa8a9ZyHNX5nBnKns1NrSZ5
nRBIpfZXScnJ3bQFffPAq+//PnokhFUh7jJPdudyNNvAInB/EOKzyZBUTrU0X+4n
423/k1/BTdEIv+w3w+pScypHSAfMgKFFdomMS9fgRup9zIdv8tijTRld3QGJ2mi6
3MeoJclcJVuW0ntKxWYuIVwGpt3IoCzfhuBY5K6Q5IkEvNaek5k3Y2o+EWEmUPqj
UHkeO6AjhSmDxkhQz1puc8t+qLC+GpKOM0sHx4GrlWGzgvenZQmBhu90n3MBGPfc
IbRj4HYDBmAx/+rlKDObWLNZCEU0rOwLAFDIosEeot3chij/BigH7ffxiiC4iOUB
8z1NhyeMk4MlAI6rZj39sNRKrrTY1lIjWg4/6PKQ4RQ88jNU2s5XAStiVmLIiJc+
0W0LgXZSBT4bh8w9g+on25Ws2mIrVWA6+BVxDzZj9mMR9cCd0uBY2atjNbvQePBk
ms1+EdOuojJTZwz8pgV/320jHSFEX8pHVuxeh12tRq9XSfN2KfCDy9YeTmbTzBbv
PGV8YYZqy9FTQHDwiiiceeU+maCDQUNPcw2uMUA0KLau3gTk//HvgfYPjhfo1OMj
MO72zG54VQFIGr6NgL4P5zETjJ18zLomKLJDcZ7dHMqiAnAaA0YckxrERroq9xLj
Yef87XzQTnYWH0WtDPdSR56VDGqFbq/cBqq3pF76jYUnx/R/bh+w3a085je2XJoy
57hor5hBwiazAWwfQmVYjCYcc9FltXFu+rwZNFE7e4WakQgBYL4MyRVAAbEmBV4l
31WQYwU8Gm2soJiDyAVlWDyhbP3pMD8OuxWJlLuBXVso/q8n3ZLbXqsalea1gf+Z
eb6OR61RurWRalDnhwjhWf0nm4apof67WTvOfHg22to1mWJJ1y3wBZCEX4QnMSf2
cnrRZlIvKgvSSbNYUBexRe5Ab28Hd7XMtH0HNwmcNrETveEYO6NLiwlysFyEiPFX
7xwlHCJUgu6pK7sy+8L7WefhDL9pEa73uF66FlY0ylrIe3ZztW79TyBZ/tDiBXFZ
RwN9NLzui73JP/i/sYajzjwuPmGLsuNtttc/eyhmMGDPH0XaSsgFryKAfjCHpscY
2Y2XHrjR2N+Lto3BCtAkVnfhz6ySijvMXJDU5RMiIs5J4AwgSo8YvP6Ssetqj8s0
PqWlWHhmINxmUhv2DlQkAuBSz+QuIRXuGRMzqoYLbZulKN0tFxmHy1ES1LGkA2en
nXInOnG53OGpEy5bHa1hDk4MagngApfIr0/tpSpOn+GCvxlSrPLT2q++tQ1VVcHl
ow34/pWEgGV/mlo5djbYqqZcddz5Q/btN4peqP6iWkBh+zChdCy1NXyk9Ui/ZrQB
9LZJaN7qZj+HmDw18MpJkj/abDUfaxifTv6NwhDo/lQyl6YPwylGd4VZXybpE6iU
OU73kmiEt0LQDvvPfYkhY2Vm9XFHDbOVgG/mg+NVjGOfkX41NPo0UHAqnxPzQYLY
OaDKhLUqesaSf66xq2dV2F6dKKVvXpPJtvwliBebcvBDrqefFTFGUMX8TxzJCmdp
XhLunJszqwTq8u+b9MrJ/4XSV6bE4tDP81RvpZ9dulpcy/W/bZ69h8qVwQwkg+c+
utwdGjPZxkPJ+vo2NwuO4JuJzf2Fq09uRzu6BwB5RzrfS2NBHbdz0pRcv0pS14p6
8CMSv6YwHV1oOOf+JLuFyUiscKFCMuqIKMjIB/+dCX3DnkoC/1CvxcyEfxRCiX21
rjEe6xj9tdYB50c2pbb9+NyQn7/xsDrNmW+MsS0uzMD9U03pm8YTgXCFDX618OXM
+mUZR4RdAfA+mUwahaKDi71mXwgV+dNLCJtp+IvqxCZO8xklEfKNfld7mBig88zD
BWTXtyWWk9JeR3KMXwKeR+KfyIG4I0SONWfQ0Liw4rA0KVH/L9e8F6P+l2eAXYZi
WxFMMePwkWEiQlGvLQG9EevdxOnsqcQBImOPV1cDGusrBWlVZMmJ/yassgPpayXK
cAYGzrTg9q4kLRiHMGsaWWlCC9V+3Y5hFo5mhRFuzrbuWrh398CYkDlBz4VcMctu
/vRBY8tlhWdHHma05TDrWtmZGKk0/fRWOOEE+MwGw2hsl+QhK/SOwgowH0hK09PM
rla4hQw7IoP/6iMdLEmtOQLjmzJLqtozto5SGYr2iQ2kiL6YG9u/+mnGn0EYF6fo
+DvctDdF3k/kdshKCT7Ih6SPkZZFayGxTn2UDYKs2QbzJvfnlCXfjMjkroKlmXgY
uImputWdt8TVyp7x8Bsphe9LX3EbHidid/yS8TH9sE1SxYkdkg7+ED1TTGbLWuON
2Xyfg/HMUp7K6nnlj9T+MpUpy3qbUDk5ww30zw53c715ltc4LGw6dRU7DFNo+qzp
1tETrTXhrbxI4q/pt/Gz4uWKi7KGN3aSs9Q+0IVSj7+Sz57VHPBPHAtay/nWIhZy
kTCvWmGtMbOp1E6ragzPQ017nVi4ue5k3OurQE+nMA+3w7TqTV2sIol42719zpiY
oXAF+FYy+jvokvDH+jNjKcIHcI2AjClUEWsMKjpBUlw/M8sVf0ylB8LZHTdZI9JO
D5WBUXyG28bF0hDY+zK5xeder6x+MLnlJigpNip6kjoa3oIhU59XssLZpo1mxMmV
swjMpB0GSQSSlSaRYTc2X6vACsADOp2U01LlkUpJVRznVfYhm80f2k99J2E5BXlR
MIenSaTPaHbWs2C8LS2E4iyG//x8vZ764Rh0S2cZ1bFIYPlmFvHYdfkd51AiAM72
K8DHnDYth01GoDSOfpMo1RQrDBESbbhAq1T17tVZtwFVUR//cWghIFpSKDHwr/11
fCmI68ZnbwijtFsOPM61WDNR+td482m7P9xTeEe3i1BjRrZMvxdzSldFT0JYJxmq
jA/sE7T0QDptqkNJj1D1659A5JPVr/oRg98QEs47KMgBRNJtLSLTLNpgqmRhtH2j
FGxsBqzRNrjpi+9bGGMjtPLj4znaGJbqbF5Yq/VtFly0WTWX2k1jAjDS0VxkVcqD
DENAi3NFeLPjnehjvugEE2s4c4OzKLfvM5ZHNYH/PezNVdK1tsvOGaiUPkZePUoP
B1JBNkVHYM0IHIrpFgY4eO1N0QqqXrWbVuna3nUIPi/uBrNmSGIJjNYTb2e1qsNE
6mLwiYv2XAYGMtBMzSupApSJ8rfOYNMFdjXfHJs5C7OMcto7+DdsAR+0uVdS2jkH
zWASRpVXB4yYfof6JT5rslhpD2ioCBCkbGSQnbOSQrnMKZ6r0rDGIJ9bE+vVxaq4
29idgPU4CEMBKP639NKNzytIcu8je4G2r/lNN9tIN4kN6vWPG9x6UwCqsrqzw2+f
6bX0d9VgPV7dKPQJ0hrWFojmVdJLQqWIoxUtXg7Gc9bNP0weUbqEUUecJtCV2Ago
Kp1ai76fGpCL8657YQSTj1a/iPhaekMd39rcbJNPUc1JWBTguFiItkIwV0v/BY2P
9cDo/ZpN7d1lKCgUffJ/6Z0JrGyN+PJoxfohFvE5Jq5/qLbPrt+icwoPBj+LvBwn
gaht2dKqROriKtxXxfybFoVmGIWdqs4ZF00XjoJtJisA6r8Df2hDRPSwLkawfjFn
++/qeOrP0qn6fxMzTjrXT/O6ZLPTPLfIvXsoe5flU9OCfGL05p8Yjzs+J4u33gUD
JNm+HgeMUwcJ7oGEG3AQCaletVK2ltNxL/2uhyFXtHGWomQGctsdFjXzKrzyjS4H
V4jksi8lh6wYd/Y4G1W8eTtiQ4Zf7+l+/rvGh7An2BLl1LZwySLQJbkkT8rWg63+
KwZfEoKDZ5LZB/RaNF0POJYw2f9JzzAq5stJL1kN4NhA+YHJi49J2IJV5vNL3c52
/VrnCP0u00cYFFdqhUgclxziIczQd52k9dvYnzCxCiQTWLHrHFnW8/BMhNDWMTWo
2lF+fHYwl4lq0xpNmvD2/87ErzsWvtDP4d+waHQMRqHL3FpPXA7W7vmMwAGk30/b
loLYULFbQR7F9cBq/HEbg0Ov3the0WYGHyirFYW+EsF1XTE8YWL0DTFMuEjv3dae
UWTCe4IMwFGJlrYl1aLPwOq0vdZQO/ozp0OKjt3s6kMisMZTtQFmTmSsBENPiI5p
YVaBBGKgUNSJ9L6hgpZ5Sddh/YWj7LobmoT3VvXoYSw4/zgvaDKrT9H8CDmu4D1Y
UyqL75NppeHHUcRq0hSi6iNqW5b3C7CLjjJr2IfJ4WxA9UDlQqePHqQ59bAmEwMj
fOBC7nPlTfqYqvhMtMRF8w47/VhadcnEmfkvZALluZNptZIU8S6VN1gbcPNLgSyr
0qXBQ7j5xCOr4S7vCl4Db/k6DMGmdP95QreFLpZsypXF2mHpZ1EHNgcMkTmtXhHk
dRrCuJ83CJcumGcdyX+it0FstHtOs+WJjl6jWLeCQGo7YJC+oNyJdjES0wsETvuF
bfWEnhtk3cEAISm690B5wg3oaoTIQaF0azPteqjuGJ1wapueJVVCNmC04/rEFc4c
uFg76ZFxTTH2Sb09MhI0EQGlCuew9NRL3fN4gQu9u2R4KpbnBl/YuAq8XwIYi6Y3
UuNbiVADvVASFsMNLb3les7F2nL8TYAcjH3Z8nsTr7jzYd5ZVAWaLKznKsAGoJb5
HwlANdR0P0HaehTWFJHv3UEVjxBdiV/G16otR6A5DGdXKCzPEfKzQx++ePB1uaUD
ziqgacVl79gkBMy4uoTioHB1eGR5XYnyiUbHWfQcmIHVw0PMrhdLLhFP7OWFXefl
kUWPk4PFAjGe8Yvr0akmuCQia/mKKvEOnfZnIGPL65y9o8ukNssmNI/hFnUwodaM
Umbm9OR2S2U7qC3YzPi2z4nzygtcrH6MiZHj2j6ru2CIWmWZOy544qJXNW8kG2Lt
435Wlo4UuLEVJYbkbj8bKOsYFWRXVbUAgXdIdc22Q2JHtQbv3365X3PBMRHCl/6e
cIM8oDsm+vilY/zxMZaA+fOXcoWOjQNAEVREkCXD7+v9aTuUl3sFrlE5ihMA3JV/
td5uTxvC7vwNf1crevx2N+ESjEUffyv4MuFn3JwFCFPLVySEyTLy+Kjt1AcS29Wg
8/7xWGf6nsY1mR9OM8P0/uoBCouzd4DvlwH3aICyNSOchdrRpC6lg7uiviHnOF0w
CXrU77MEMJOWOo8+l+VaUh5udQpknGTY/hKj8AE3gXHfeHoavi2sxFI8Xkrd/xQi
1GYKWxYPzhEo6HwImFdHb57gfB4xH5oWdmxzfT/gNipFjShF7Lcqcdma5ZA5W67G
qHdxyZni4sB6OD0rh+RENltuhz4LHcwnuQGUD00IAoArg8SKqrzj1HjOY9vkpFJV
Oe8GggnBtF2DmYZT2S7PZGmfSxYlFPdfDy9GG23aCKg5UCq8Gc4K1jR7p0TpqRiz
n++4z9Sr2KbPqdCWY7guDnBvzwRxL0xk9LVNHyyBUhH8R6/AQcXd4PMSJIdrhCzm
fHo1taPxIvavxOExfct88aRPb6rR/HXTgPwCirii4BEaN3btKf/LhTyaj5FmkHl9
GRcLZxSnzAJr0INNIe42MVceriUfsmHMg67TenArSpkQBdMJ0ezl3RkGzJH0VreJ
JJdpAwXhVlR3tlWeTN/r7F6j9f0TfPARDucBl4qjQM9Xda8XPMnZ2y5hXS6qLdTS
Ppahjd8G2OPAwCB/rQl0kkj4/XpeRLuZPzO2sbIv1BD4gEsiPLb5fpax4av1F4co
N5rExBVoeHeIS+iISELOWtZxHq9Ef+23TTfQPaGt56x4HLjF5oPoI+RRR/2bejQr
sfCIBNz6yc6b4WpcyIOq3AvcHdukpX3+J/vwvkT58QIsNlYh6+u/JxdN/RueYdzv
ax1RQk08DcnVLeEunq5HACr70NT/NIq/B6iiyY+1E/b250gqwM79+4NjoCW6L7Sn
ZfC1MkiqsdRr7yhPYTogOBTiCxf+zjc46hzxG8CO+SVW+wKMMs3zCzhz1J+715JU
jO4w0tJ2V9MyM1nm0bqphoSX3XFGXVMJuNQt2hdhKEhAJbYAk759Uncl789H4eLy
POn6vGvD6Ha5/KLuaHjEPWoTNY4bs6D7UFMTLXcQxo3XjSQ/AvLmuBcAopJBhbP1
yYB6yaRxx5jsSqynzAkwN6qHC5k/wQIiu3PqyOm1j6fn5hMk+0P4yzTAol0uqdf5
KESAAh54OcKb5WyjoeaWNUWNxSyutsvmdT4w/IPfGlcqb++44Jc28bziilYMq6KN
a3ALaBD0KpC84UmKgvSSk7CrIaq8Z4ODCEiIkBxuWgcmaXdFKyto+tzBq8NihJyJ
ydXRwNdUC4zxL0hyn8wiWmSwOP/A2GOkmcbIlBvT3NDBVIiqUpzYjJL4OMOfXlHu
tCrXjbMWFSd7fr6ilveuZ8uwe1NzCR/G4WiJGVJp2E2d5e3jlZVd6Lqh+LOo6ivu
pbV50L2Zoi9toYnrXURAAroEal9FCv3/BRRICFytl8yjeSI6YCCtgm6A+n9u7Ef/
PG8Z+0Ft2C8LSLQxdqLI10EsOeD30Mzm610MAoN19HbPPOZBjbDzx8ED8TVJC1n2
90F+5nRhViUyVppYoTBsJ+Wxd2g5WilYKoxk5HXAN1F8wwPdWc4NIRCQpzV8/prf
8Wk6YRlXyqwpYSwedvI+ZhNOKzS0mh/L43Np9O71ojsl2IAK3L43hPrGX2px4vXs
TjwzXhnRkx/FS5SC5tsgxDSllI+jlTfD5GjTGM2tnOpfhH9TzNih01VLqWxBlQHP
M8qrBMkBLSvvB+zFv1WxD1IY0q70h09vMuLhlmzzBPysiA4IZENLinlMn+SiyDGe
+9jyCWxeIzfgH8fyszpGo9OuK74qpQHxd4lc4RYI2vDyDEaWTCaiLkfBqDRqCixr
NE2F46mAJZH+Jd/OMbTN3GaXmcHnLadtuG7l5yDe7yF40P3nmIZkSjX9FaPrPIk0
t/VD2W6Ee1qdvggG3j8NClZfcrXC4s8dFwh4DiTJZVcWR/NbMSGYtf0ULyEaHLuY
mfirmXoK8SS7WKK4fMLQwJ4vlklACD15eGl6gVYjxq4xkzctvwzxDCizL7gydTmT
mrwJiXUMAYvy6uESbQmH16fJedED4u73L3uwy8kovMmRl3B2fj9lHkp5DNaoPQxl
FcWY9jbr5XPh847iHvR/zC4Rk4c2rX+AlAkHMZt6aD9XSrFVE+4P2xaxw0tpAn2u
WCuSAVeQq2ALS+aQDxFCcY91PU2F6KT1NJaWY2x36W5jsTbp0Pa1jXLLMdt9sRo5
7LIaxwQEFgnG6LhwGv5fZXJxMiQmbK9WpjklNuENdYi2mjl05xi3tyRE6h1qLH60
JdQbMqwzWCBN7lDZ4o5nRtqltQHx25ns9h6PlLHVuk753IrD+1vxFvS2ZVmNW3E4
9YkS23/RGiSnBJRNZatPCXz343WyP4OIuxynNJKUkt3PCk7GtWHl1COTXOIYLJ+0
KM1bsPdWjUMsMXVFiJmFgxSlV3WoT4pCxc4RFytJSLIvO/fnz4/dMME84FU8XbDg
sXAX8bVZQfZ4PveO6zV0je+ZC/Yj9E/0vfXzPNLexfFOcR9V6ZaRLrguywPFI2ub
5d9sEJp95UmoDDr14cFhHb1JcFY85LxYouzSF+zQAG7GixeFqiqE9RVr8WmUgcup
kYOlrJ9QOzRSyzqTTJD+JfC3/QCh9x5VB8zOHeAKzVx7nGS0tusoDJc4yFR3ds1g
8Jy9eJQDDSueWLSZlGGpIGCM/A4DHQMezpZSWwDcO06Dih7VdefVtJLFGMhXxtX6
p8y0x1m4TI2VR/ZWFQT/+5cbLQFCjOGCYNpJU3x9hRkq61c3IrEk00p/mZQRzXYP
k+fQtUp2Y+htgZB4q27dQA2indp3wjR0yd061MmvxiO1o8pvU7KHL+1f8rtkPQ9o
h7e5qudBktHVYQMF7omxpI1dYwVvsmlSZ35Ot+wdKPC10PtTgbka1xFgAuvXZ6u7
mNwc0Hwo2eR7UtG+NBTS8IqdYsXhaKujOeTD+2GLFQeAEa9arJqKYnaD3lcDqbJs
ypCoS4fc62eRfwCfVQFRYyWBOEQ0MqZarTh03UyZVo/W7sz6h4TGXTtTyloho3DP
YUMDB06H2azZeRIEGB8sYVMr+Vx4JgpjSZg3zyYi8aIdkb846XbqkhnmaaxoAVV9
eKUnm6qctMB7H/v+Ex74ECQIM7Vkxrq76QRMpRpPJgOzLkA5C6YBU7KfD8UfY20f
jz81PobTuxZt0PukBerZFH0cdDq+UuSnPDhyGDKID9/cjjXe9h0TsjWAhrrp4ccx
akhG31qaIvn3F+HFANks1G9TQTXvyFaDCoWZYcDmTNeFMUQLSi+9UtXNDXlx2Fn/
Pb3TBfEuzr/yGTYSOvzBmiyD23bqL3R/Ve6JV0GSkdNsWqiSSmh9+kqWUQx6a8jo
CA7t4EYi1h9L3+x82OyS/hfzcLBldL2pT0umfYK5M6knBFM+bCl9tA3WN3EAI07y
n8WJPZs9A8U8Jg5fHGgn7zfToUom0bc3pLz+PTa7cnJPEYL9/jsam5sv2ChQYqZm
5z6Ki8H00CdqUsJYiYLbgMn1QC9zBzG5CEHNgRaK2xijsQuhGyhzKm+RNrLc1Hod
y9bj5EQ4WLx8pnMpQRUi+12inVz3VjAsMlPU+RhNcOz+9gxZzTbAz9wwaVXbrMl2
7tIo5awH+6ZHKC0DbU4ALxwareBaYfyFUoJLHSzpwjGkGySXIucy8FXn+TKz5tw1
ZjvgThEBY1VeJYkF2K4c8iUGdJgv+3sVzZAVwvORZHP4tyNBP6e27NUSrUg5mq7a
tEvSRmooN1iIbydBeGpsdjswfb/pjL0/Y8La1yXt8uNMunhIcQUeNzHMELCYCiUQ
X+6o3A8oaojeKt7zBiYS3OsLagdneLMfxc9pLObhCQJ1wEHQ4nweRupLKsLw1ccF
/gxOFDJRabHfsh9uUfvCN4y19Wn5+PA6rpWby0OU8vTeJ/2I9vRBG2JsK0w3HSXH
NSG6mWBM7fEIeLAh9XYjnndhSvrFdJ9r0w+jHuEHrUauePVhMAJ6X8VVG5vgURyt
9bban3Pd7DiWAtvt38Sg8y82F2o4SfWWxet5QJ8rpauODkE3oQCwkR1G9bUneig6
o/DtAGvWOuMHp3ctkYLfAWCZtdve3GrCJbk4I6Oq1NPJz+7QSMoQKIesmOhUtEyG
DfOoSWR5qLK7CxYE56XM3tI3i81uTLV6yQodrj9rx2UmMV6I6c432yZGAdaX/a9t
VBZMFdjNVsD4lCFY/ChKwtrAa+qCFcqMjX6TcnDe+oWRKgSzJGwjIxR/6yBs6CHk
JMCpy/ZBWqIto0TS8chBXyk9QqjJnNl0hXOPw5yb9D8H9tRugCP28tTUEUbjp2Ql
I9VrI7VNzejCqiMmJe9MYJvHnzxW4qzAwYdkmHTra0yE/ZB0zcN8ErE/KtiUQXzH
/Ek797YCvSAZ7cndq+ET997c5mQEnJ8TXPh4FLWPrdPnuEtfdSDszJ6hCC6NRD3W
EVppG/st/qkVKAPpYuOgP4hoWs0IeOBsiJxigwbflo1mT7mtB0h2Xs+B0PxGKPnI
JYr2KufCNJ7wZGIyVLUH1cfnTfK3TQAwuPMGIapMBgvcX4gupwy/ziea8uHxZtKS
yI9mCNHLQRD36zAc2K9Ac3OuNLBW9Neijo4HrCuQhEjj5rEFaWmc/oqjWmrPNzWt
jzTawhmLIb8z6wL5opvz/Cb4w38fOTL8dnWe/gFrLk04jn7hTKfipMVSmULCXoC3
eQ3hC6nNcuq3LJtG/BcqFpXeJ6ok2mSo2oMpwGCIlUTQVj4cUgDmUhRNGJZ/AtMI
VqM3sERXnhotTBRVhO5CEvYbfVbVzQ1UgY7eaYffe0Qa0CzgbISyw0L1dlclwAW7
Htn1S1eVCvxN/U1Xfy4eZQ2B7HifoFINArUAq4eX2f77Z6y6IuLSkWrWnJoVaDJE
VrnCoW8zyOUMUFINPlTx+hRBzx72wv0hh0jeWxHeTGIExHR1aLJdZHCqjRwB+0f5
iHw8ZmUVaqZkN9R6qCaUWpBVuRhZEbjAufv7TK24KsNgk+GFQCCuL+wEI94dz0mi
qVJRweMMcEkTfZBHqoJWw+0w3UVGzU8yYwsYywRuH8CPDR5nZ1JDZ2v1CtRG6CZw
ui6JQULgKHwClb6oBlfeXdK8gayaugFkMDzGeYlqdoAHix1LpQkLdTqY6JTHyYse
QwQtY4wFy84zyexh6fP1CR8abfvl+H9ESBLFG1i9gJnBzn8NekdzAgoP2qiSPQDS
sXxgX+hF/WKFzOmjYYFT09Fx6b4zP6L5ArRsE20asi7r8tktvdOP8NXtipejcJkB
Jj20S8P7nXnoVI75hkUWnK+/JVyCEq8ecWVmBc8Gg4N7KKpf/AuWe52FD/V5Ua3C
QPV7XoVpH0EK3VfqVcrN6lpelsp3vVdmK1AyUc/FrCPPD5Rz+hNN23fm+UA3SqZA
LoAf5Vjsw35Yi03A0EGzratqp69Wpw2J4Bga+68YBFYxEj8yTNtLOBEgydWQlJuN
qOk5sCvCcvBYA+KyTsixlcHo6056BY6O2uevb3BAXLV40OskjBH3qOKBVBzUjD6G
CCKlfcSGLTkKshuYOo5kfCUIkRM73++lteb28RsRn8saQ7P8AXgRsKfePERAIUr3
N95uGtHnj19BYfbsCbZqstHzRPRiJYG8W9N90qrT4/isEqSaRZrrk9iFSknEGadx
dHvK//ooBa6qSNx2sn/YgNIP98CxDQ+nr8BucpKAZ1ddlCWORmUTzWLv6ApSY2Ms
9iBDvZvhljV+aOOBHs8h3UCez/GiF4YDGiYc+EmwT7fCAYJhhAtOqrZF6Zo1/99a
LZQAwnU2PwUgAtebitHZrtJyiK7vcd5/oJoQCYldTKXJKEaNQwgDnGP4UngfMpil
sPhbnhEGxssMHYz1EgiHy4PEmhRZjoGIVN2xmVjZmXg8/GF8jyYfWuBYLZ8+cUPh
Ii2ZZqkRu0iA4OPqfGhWz+rHLZ92Uhbnw56uCoaSpmaID24KveBasm1lQS7JJTNz
hwc24YP8ssq6BNvIEAMpv5l3LqSSan9OrvaU7v38H9QMjT53UW0Q2DCaqn9fsqbn
AVyxSxVbZ+vEjmRIaYMlq/uc8QWDbOvZ5nyH4vxUOxw3lERvLx8eYTwKfWG6el62
9pzYahzMRU77ax1Lzx9a39KxAekNb5yWCO3mWtGWo3pxkUfgBJt68x4P77oRvUna
rmzkzKC7XcCoOazpQson+WPhBDWnzE1naSrlyxFU8wi+ofdP2j829Aqaz8jkCEeh
+HJJ00EQLVBm7mHDRfeoQ9RLTK9ZLZounZQNtF4ozA3pSSTsh2v1PxY0O1AfjTNU
Lx46sORLbjeurmlcRup+ACWk0D/PMUFk2p8bK4tPk6QBrllunudFrRB2jiBSlEhg
wz80IH5OTu8z2vgu/uy8frn4Gu2Y3BYHq/QvZbC1KTJstUpcAAS6fn284mz+3nwk
WLxU+6MIaI4AxJWaHIh2eXGQbCKYNQBCQEyp8vW6c+/1oLzI37T4clbPVko/LPxk
u41L6bJFwLKctcsWZyLL0KvCCnYz/6HJ+IRUeEsYN12GPSPCjykt3CM2liYs2yPI
eHP8jAxZYTM/Q7v23Sq0Wokh09FtQahuW6tv2rJU0WDdGJVB1rMOwb95Q7UggirC
yOXGaxHcOoI1wLXSY5ZRZ5U8OtEtifPtxNAUorJd0MfLacRrg8lIrS/JAaYvG5nH
H06tOf4utMBrNdc/Y8B0Qc7j62PjaqC/FxBYT8nvu4xcfscz1KivqbLfYx9VTmmn
dBYBm9lFhopU9M0uCi6r7SRwCH6PuTYtutCokpptJFQ/2xqEUMaPQwMD6/0pAImY
Kl3V1z9O1zKkGT3BaFW1k+9V9IZrZqBY/vs0VlqF6G9SaAWXitbxLhKcXfH+cpZ1
mzWO3614oBhTShRulhCirC83E2nepChP25priW3zZfPG1dO+lT6sqq9gqdgNW662
5qWw6tOFNwQSKv0/Bq/KjB+47CP6cEIEmO9l5fMcWt+PkcRM9vGlY2uOhFIwM5zb
jqIUd5UHd07KObP5o/Qh+PnX6mJ9ZzBb4E66StmhyWHJIcEcJ0ArWRp/7jXC6gZy
P2zJyB6sYaHT9RaHcrku7kDTXirGFkR5Iq8j2TgED22+9Uy7gZcpmDlz6/VyW7BS
xdXX2GujzP4h8y259q++gZOgmmweneZZaxZYA+zKuv2mYAZi9pEd9D53WyawH8fV
a6cEfQr93JGHgo086b1suLGOkmWxcMiy5/HQR6AWMn15obadXVSLOQBFYmuWNv5u
hFP9b5dGADtCIo9S2itdylyMfy8j60nehtKJXiB1VPEsncIWKKJWAF8iVO3Yjx6x
5ekTAjvREhJLmKISq8w/ceHqqCIMRVThb1Qf62or6GleX9N+L2Jkr5/MlsGd8FRg
Mq5bfOJpXCrWoQCOywaeYUK77QIn4bQ5WkOaRe081OuKGv5a6pNuFgbL9foTHZBw
jZOevZU+CJUEfbbcOJLM0R+3A1jCQ2zippaU9q8iUkkzvVTNg3KP8GTZLmNtRsHB
VQL9UUu6kinNbqzkv/isG+4fFAy71kFx6fC5Ju4X7UVcYc1ncMyY+EBh2cGJbreV
9XIvvwVR7BNWkhGbvxtmUMJRnAfVz4GbyvFlZ4UsjtiuTaWFdeT6iSanp0TyUAGl
q8nfuK4tP/ZQm3O9vc3N852HMZ1iqktgTrdgG9dhhNjPt+ZBXT+4ZO4xLmaXIjrO
v9Ecp1GDmhTCMqYTmkh5ldQSVijojIp241YMBxGfa3jiYoEihJnqN+coLRv4TakK
crOj0Z2QE+u+N1745BSdo9vJfYU1jebvInJ1jqmbPnfi0c6gHwQG+KTX5ITDNSy8
BEcTk/QPejlUTYF99Wj1XabVzusnENl21Rla5BZeCBWrdX+fK1pwW7ceyRhr3W2W
4xra2KOb7ARXwGaGX+kYbD7iV8ndn3wrZHIWNILRcP97/6shykXfYZ1sx7yARzRO
OzXtbTxrFzUvljRvGbnZUlWctKKiZXGd/bUynOYOxJKlK6lRRkRxrp70xKQ+I6IN
IsT1IYoS0QuSj8w8j2awrEQ+MTDEad6Jv7YEkSSQlNPKN53zo1XbB26agVTmx41y
AbKlhsYpwGkL/LRzh88LP+qlXbxG/JcihVFSfMmqpC5oxolGhpEwsCWrhUs1eYUd
9MvwUbtJilsR2LyxZufrjkn0xnZak9jmdhzGG8muFu3vv2LHecBOJNOE4Aom+YNj
oLV2S+N2mxCvG8UC6u2eJultCCohxYqkQryTZkuaKOsmaB4SC8Zj9eD/qrjYOlKg
2f2uChH9667zA+lOSkEwsHvqWT0Y/0stqA7YOoszIOhR/DMGd1I//h0TpyEISRHB
PWDh6edpiq/ZapObkIMSjiZ2HW/e77lfe96Cjn6xAoxjESQ4GpC8WFSIx498jIsP
xqqKhsenU13fwgYSY+DbpWFR3hQHScyLlL7urZcJL2mK1IBPj0OZ9KiIrYXq0u3X
5y4SRhYGnXWIdudc0NTJhMP/YZdJWddbQyBM2FXyz7OoUJGbCwqX6TlYvvecO+rw
fQwf4NfzkxWJqyM5fUgwKa4D+R97brszH580N1eD32XW6+Or4l77E3pzCbgiG6R8
QVjAWyuTjSTaNjFXIxjUE++203U8YbmcS8ZIpGkiM+gY9VXkcLHPt3pXro4o2Csn
XpC2byof7Fup7U70cZl9xbbLdaQTmK9wbsY/+bXPr96my58gs7ToEMNXDrOoJDe0
0ffvH2g7EywNAW7NJ1LOccR/xZLE6vxwPc3yylJDF820Bf0Y1UFQbT9QYqZnbHfR
S3Xswls7eQWbLNuKLZLOMZbiT9z0LK3DG1g8+6257tFuSB/j3qCo4/p1W6S/jBwM
c4kIx0WiY6mI3YyZAgZO+aD89U0zd22kMHe51UcWe97zSOJdrxPodz6zUBCKYlTN
d+55uc1JGhwvBFpeusCgLf3UUv8QawTZuzTPMT9xDaDlhMMO0GnkXZgtZvYMns71
NzUjZrOJsI7+61YY/zN3Ys3y+II1T7DOoebabo+k9DMF5wbOfaeX7+SjM2xbFI6i
bezg9o+jKWGj7o/JaQ82ioZjFDQwBfagU1qh46lyPXCqBFynRwCWqnp4eJbPk7tB
I+Jy+i34uAXwijo1oy9IG+a78Y62AHoc1JIxX67eqqwveWmkYOxvf9/FAO2Q906q
H1/ibVgAH/lb8eemC1jba7KxN1ufNb0tNNs+ORAakhqfk/b9sYJCvP+4An5IhuiX
D6kXJhQLMiYLHZzq7eF/mZVDDJcFE4xZMrvOXJCbDvWKJ4MfIaOSx24xl5+JbQaI
CDyPFKNXiYXtoNWILv9er5N4Qak7HHGbY5ef2keCG4/OLcB7TroytrqLQp5fzT1m
XzJRRMJOiEclhMLti1H5yiKg95m01/ig9VTGjhWTrakZz11t+geK6xOz6ewNE0I5
naOXq5TEr0vCT3KfRJXM83SNSg55z+fek2UybI/twaP4kvlSMFT9tmeWHZStTc7N
PKP1lYMXdo6tR0AX4l18RIH4NKWPKZKvblAck+YER7fMYyFfOsIfuRnSw91xuzmP
hdOauyfwcK65XpPPr/L64ZVASUWs8vtS+Ae7WdCdYROpR6xgjeqciIRD51IGUdZI
CaSeQp1Sxh8vbuukrVszRKGZo4tXMBpeO4vcfAY5xY+2ZWDtSm1NXbVDM47aXXc7
ZgZWb+RDtMRtz6t01R+NPTVi6t9s/tYAb2OUmPoV8sysyTGbovqKA8UkS0vjKv9R
n8d5UFkL6fBob/DiBGs2orHFTScCl8AvRySgjEy/KgImbvMhmPnHTsZXwi4ry7Cf
LwP/JRrU1blSdmkf3AAKsKuZw3Cbek2l7XriKD7NtBYE0JngZETRbjDwnjM4ytTs
amqJzo0pCzvii9KoYbanDao87GivhlTHrccM5o/Gm6TZfTFaIMGXVOpYZ9AxhTu4
RdYHvDScdlxRV5xe4l+1gU1vhXxqZEsFhrN8aXZoDHy4BwqhG4zKoXSgWd0gQ5HD
Q1u5mtEWwKe8zPzMWJdpLGtC2nPPKDz/ccBRs4aNyMq8blfckiYrgehJH+dxk4Q1
HTz36q5XBVhFPSUsocJJoGrEvYKU0EHYQcq1s1Sl5D2grjlsUV4PJ+KzV9paaize
PX3fHStaarMm9rZvU7ZpfCx82XvLUlSv65ChFH06uP5MM/8NnhQc4Xe0RAQXEYn7
7ieAAteL1uwtTFV9MuLCwtobCgQT+CHHZG5tF6QOxTgpYKwZGKwHs32aZpcWdrRg
CwAhbHoWU6DBWr5gE/zFKQ/X+1wvHzhUB3WUUmhpG06W/cmu0qbLHa2hLeG3q/ka
QxT/tgeyD+SAQknvYaJPS6IsFtMZtj22aDSx4zNtpbm3+JUIXPp1Pl//r459SnI+
ZAQoC31R6X/KL2Evu+lsdRYj1vHpdxe0SqkGfM79JKyFNwVVAly83rs7ywKfbeGX
VqMnkbdMsAKmzaoYJkcMiVd2Gk+QWUT8iHjyg38aYL0WDLtSQkGPrMsctGi4EAjw
+hCQsHe4lxqaDCc8mu82ogPqGgOnC/+BORKNkvRhgLEnKT2VHW2JKgQZU6yxzdYv
8n17f01XrZtKueMlnjljuVjPuZPho2EYFM4xlK90tHnpyHUM0xe7A7/vV668IsC6
XdPDraPpyATY4ctxOVdeWjEDJRDF1AOjWdHdCM5Hhhk590A9Xfr7BswZ3ZMightO
NIBvOnukDK19wSckagGH57JrlN9YZP1bf6C7fAv14HvGUxBvh8C7M+gIZYqbV0IY
9R089MH9rGsBo4eMhCPP1xwpLltWA3Eu+mTJnGtEbn9G5I36PsbO1tuBZIoZP1tL
5w3SoaaHQWL3yE21DPQYa2iUtZ9+LXkT8lk95CZH6K+S/w367FnoprJvAdkM/zTV
GOrtCFsUeBUJMDOCdU3iawSgv02zq+xsU85jVP+cA25HkADsznjYtT8CZfZQXLa7
Bhnw6hCQqmxAsTRnXwmM0aPWoVso1LCu/ZnPIPhK0mMJKhWt0SWsVjDnlmDEWzw0
bOTYfxpd6YQC4/wfnP71etj/VxyO4CS+Q2p17IbTlwucAEI7I/nkmvnpyv1yVoFY
qO8FbHJtJH14E6+8oJFJ2dTJxHWz4IAp8kPnMnh2KmJY1nZBh97qSgxoBUC0ukIV
qwQiYiWc5XMHtKmPtOkqAVgIZYyWNQvzfTtr4516LFQKdutfBTqp2UjJY7S1ETbk
gLl84SuJGF78iWQK/Tp2BbgGz8r90FTXwj9vQBUFeduDeFgG+uIbxQSHyy001oiE
zY1HTiOuBSN0oCjFAvmjwvEInlnpqxWGiaKzW6wtmOHyXokRnaW3dQomy1hAlEXA
nrEJXfynQk4MkpK6vGci+VL9R7rUz8oYWfIqXaMWKmXwDyPqXlXY2NpjbrQdwDxL
29ScifQd5mfc+23tkHJ1NGw8ZLBwvaJTTnbVWeVLDYVdIrRsuz8XDos8vwrGPUw3
AYRFVMs8IedpsPpR+moxWvWoBlSlbqkBFpGusYIonUHQENeRsEkfccsPDFGU38kQ
SLlKg84+g5x30qhYffc4U3NObrcOM1K6msuCiNj/OniGmEMEN2v8ZaH6et+GGKOz
uUEO5l3b5gUbtEJ3rsiw6BbnpMlSHN2qUR7MccqZORs4Phhh7ByIGhVEEbT7I6GW
3UY2EyfUWfIpZC+vUhSAEazuhLqzXeiAaK/ThjgIj40j2l5isxLQncnLK4PAJf9M
k1JD+N/LMpF6Gv0zwEMaPsrr9bOcstULLemh633HjVuCE/JeS6mzpO6FRaH4xJks
kwGgvTJxP0jqTcZFwWrdnjQv8i9fiLW8wSU0wZG8E0I4Rnqtn563a7bE+sbVfw9Y
Hjp8ZxwGzgw0YnHZjFiwnEpV6BpQJr0ARKXGQ5+rT4+8gfz0/8SC/Uvaedy6mY6I
SR9iGo9kun5fqyyc7Chh/yDNkaIbGZ32Cts144WCr2zgwv33E7YeHs8jMT+EOhqi
zRGdQbDWv5nOVJj/9M5z4vbXZAqwITDKo2mMRgMYFg3+wt3jUd4fv3eqaCjurfDH
MNvR0l4gu4hHbDV9anyyfo2aqFSeUO5MzPQB2L7O7s8IYTneD52hcHlL1j1V3VvG
ItxeKyHT/F58e3P/yy/Y+N+8SsH3cE4Uwa9tfSGuW6YQWsDl07wCyfi6hwRqB+VI
86LPinLzfPgp6FK+WwblOecsAofWYC1ScQVSsOD+lZEaXCMYyUo90IBT8FzrPYLB
J2Z9IaWnQCCzqQUb2/r2pkMPZHxwMj7EQ02CagAMhSppSU2hl5Gl92/1T2ia5y5E
SIskiBSMJhYbsgN40Ly/UzgXfTfTLTRcZLnEKCRjimpsmJu+CTcDgkdQnKX5VTiy
MHknc31rb9RtpNizyN3KF1ZeP2kw13XWNZ7MOlUS8TJ/INmx5nuYyYujPy6W+8oS
slD1vWNbXkv3iZo6Qb8zkvHCbRrfTzcJmPyYgIYliRSGmXT9ZW0zBPppj/HqLpfe
+E/HLcsBTBMHcO19/nTlDQUYI1K2CLNXWMUH5ljMshjXlQURgdmqHAxgqHTCciTM
Awumm+JeyU/r5U60GqXd449SaewPr9+q/G3tQ8ZkjYl6fArg2OfD1WNLZoJ/14oq
TsQXyg0eaRWo0bX8YHQA/lOiR6Zfq0gsqoqWjIbipJbf5/l7+1uibxNLg9qBJ7q1
DUptm3ZJXFvdocYwcSz4JmuuxS8trDSEJ6E7CPkJev7HDhtiwsiyevD7tuAABesd
9pmzS5+9rIRT1URqq7caWZ6Zv18jCgkv9Qk04d6jSRExUb9K2szf+so2/Fybswua
wRYpLIRUKUu+Zh/IhzNWyh/zkcELEMTtPy9z+1c/1FQTMtNg9oCtQN0rzgAJJpAq
eBmhoXd1BOapr27m0+OyV8JLrHJn8TtKrn5MNfOg32G4/lVjCHNzzfkxhiNxKl6z
lbxxnnpVDlw8wfcA9rQsPWspWBAJU5UWtciNuRpHty9/Qdknybp5pDjFA1UV9MvM
w4M1izZOVsoiHAp56dNGQc3u6nRedAKPHgyip887lVnqC4b7zThQCpwaZ8n6+MNV
SrYqgzbsmcm77U6M92nfOL2C9LDPoRLoU7d881Vj+SIG7UpBamFbKi6ujveBdnbO
o3O4HH7XHIBfYibFiapllkeluDPbtRKdnstklQSxbvumoaIi/YdJfrkQlEI+1hz9
fQCsIZmeSnvOx3LescLZ/9lETb2jDN3nFLRBp4d36dHyYhTgujLimOZ1hZO/3Ubt
wDng0PW7Kjvx81Dvyrsnn8/GwWedygoIa2+KXZkadIeMglgm+naoX9cF5YAv7y/t
YB/hL1IGHDHdNhoZC90zzI5EYpmNz0ejWSpJE9HmxOLnk9RdBTG6o0FvFdJgMFpD
lrtbsPV67mGCyHFuew/m5tnvfSygTjWR7tmZjNhhIywdu4mayp4fyc0YusvWprZi
CLVfaRgPsP21npJoFjwhneSP2st0PHirEhKHpLW/k4chi2IU6nwFwlnDLov4eS/6
47NQk9yGh1v9nYOluf+e1pRmqyCNS93GSWMXYjEw0XeJVe6AyVazP98fjJnXSG9I
3bGIuCd0QGCT5GYx33dks3zZQA6SfgnBjHzPI/9jPkuc1UCeHLWdmNxUSnTNm5ae
A18/w2ENhjHrTfKIV/B48pZHOO40Ekl+LZK6PLj9vvr6Yk5/pD1uL2w4sKVLcmil
IZhTQS2nRb56bhSlNN3u6lZKreVoJ8Qm0zbZjkKpHz2dVPsC/c+lKHEUJUM+hoHE
1ADZ38Do1Zy2obVGzGQv4rQXhsn0+hsTF3gknFQxTFl59Dpg5ZYiemL9aVhn3FAp
+TjxnI3rNrSn3m4DEHbbcu08ABVHGJ6j2+MYnVRINAHGtG/pn5LXEo+wXfQi4V/h
AnAnJacAzj1G/asSqEVsWgoi06k6FDI2uzTcJgu4nZUgTuJcCvVEbyV+4YitmyFA
`pragma protect end_protected
