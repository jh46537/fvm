��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbYIҚtؙR4U�y���u	�����pQ��8(�p��5*�4Y ����r�S>0��Õ�!��(�au��#'�7�A@=̓S/��N��$umޖ��	-��ąy��V
t��=�I��ӊl��`�0�iZ�񦫿��Ȫ5�1�BϐMH�Զ���U���~�	h���͆���;�rM�(͸��L�>F������<�G�< ��aJ'�4�H�J 6��߀�/b�N�ZCeLWܽC�{Ǵ��x���L�!v��a5�$���ϔ)���dY��$AW7��N�I�=qE	cT�?�0f�Q(�0kHE�$f0V?��^�NV���X��� �Z[L�O�播NCA�u[��/�.�g�<��s�+��J���K��]'i�p	��� ��KR�Y�D��xI���Z"a̿NPO�'�9�j``wN�Q>x��XWbV*�t$��i����]o;k8���ǋ���~�f��$�@.\�r�@ �h0򝝸���if��}�w�p�eQS�4t�k�Ru�!�*[�3�9�j|N|�Z���Q������JG5s�`��RiJ�(bJ,�Dk�W[�Fd��g�+j ~"x�a5�>����3Ƴ�_���&q�S7�@E�l��aߔ�o�w�^K$����{ys͕�s��N�\W��Qc$H�{Z�2���+�����x,�[@1��J(�*�Y�>74[N��^h!�&_�j�X�3";�n3���ӱ3��^7���+���s�kK�f�X�Z1!���p�K�#�	�pD�fe�^��s�vOh����߀KL�{&wn;a�P�'f]�kf��)����P�(e�/a�C`.��#�C��-�Jdw{��!L�>;0�og�q��FOç01�	`2���F6���sh��A<�~I�ef����LP͊�e?��Dă��d$�:]?IRHfM��-?iǭ:����	�pMS7WHwa�EbB3�ϵ�#�-���R3��֬���ʥ! ��p�1Π��`�㷖SR��]�E��E*��kٹRQ 1�E�X�Z�[�ެL�k�3��� �?��
O�y���i�d��n٭V(T��:p���s(8�'U��A��YX��O��)�_Y�XUB�b�5�R��������	S���=F��S���$ᬇ&�47�'�l�i*Ϭ�����F�FfgUT�0x��-��v5�U]溸��a$xQ��x'���I���Ҭ���[wz�̋�C-n����A͔j�NȀ�n�qY������*])7Ìu�"�o%<[? �\cx��{28�5�$��LD�y�F�iR����j����Q�<�'�5��}F�w7��E��aw���H|����y�(�g���Y��离�`H����Ϟ*�����`Xv��x��8���x��ZѦJ�~��*dP�o7.M#o�������+� ��D����Hp�Dc��̗̎����֞��1�gha��R�w�\,�G�з9���R���<���_�l�_]o��h4 6*t��6��YPa�),T>݁��<�������!�Y�MT=@�!�<4�T9pDM�$7���v�6y�ʑ||=V����dKb��S�3��ְ���WZ�K	,��O�m�G�ⲻ{�_C#��J"ߚ�_L�vò&�`��=��z���ԩfݱ��VO^S�,�WN�� �69�Bߊ��o�U��fn�:[K��Ww�f*���Z�(X?R�٭� �������!z�;���0����S	���Y�d�R~���ZL�{E��a���-��"� 58/n:8��g3�	Z�h�<(�_/��i�|u-�� ���7�VShnϝ�c�ef���a��v�m
���;�7���}�lCP�7~���c`�aO*w��P�����d��M�W�O�_wؽbo�;���[�?���գ��E�	۬�Vt�H��|��-�Ո���}_�1G[���� ���A8;�T�a4��ˈ�؆�J�R5�իm:�e��Ҭ�B ĝG)[ �o�f��v���CJ�Ў[{/=��������� r�~��R�gw���=���q>�KP��^�>�V�n��PĂS��1���9�k5j�~5�pa����(7�1��Ֆ��f��jf�l)Cc�QE���AH�(�a�������������TTg�?�B�#kU9z�!�P\���e�f��	)Srn?���]��X�>r�.�XǦq�zo7��N����@q6@�v�ysh�4�E��N���G���F�� �@m�2ɶ��vF(�eX̚D*�<�����?4�FE,V�!�֞em�/
3�g+�����PUi��Ud��b����!�>;�ojE�v���[ż�����u��U���d�X��JEq?�����Ll-�6�ج�Y#��� �A4�n�+�N8v L>f6�Fd�,�&�<a]�?����09莴j�+�,�rϡ#�Ъ��wϖX���PlY�g !�r�Y�[9U�<9������}��@<*a^��Z*���2�@=��;{����s�;�oH�4�[�o�2�TǡH�`?#�?��د�|K�����M,X7y��_����p3H{��l����]�����&6.��_%r���i�*ڄ��(�F;J�y��2��SI�It�uF�!Ȥ�X���"͞Q�i~���M����u�Rqk����6��g�0E"]q0��@������� #���_�9��E�c��CD��ͽq�M��f���^�_�����튨
[��(/�f���m�aX�I��a���=��ӵ���pj.��f�<������[F��Ω�$��60�}/V]2mEЃ�UU��n���t�	���J�{a�5�}C7y&����}��G�z���6~E���ه���fE���uc,�s�?�w����w^W0�K�sQz�!�����N&T	����U&%�}�0�Lݹ�\�J�J���s���6��0y�T��C��@�|�� �Mh{JG��zl�}�Ҽ���6�p/�v���89�
��B.��q�LS
 �^{�Y,Q��bu��a���Z@�ԡ{���1/\�r�e�W3�ip��sD7ĚM��W?&�����Kr��3x�r9{�9P�V5iu]��שMd<tyQ_�&lE�h�NP�O�]EN�4%��"�AY��ka���-=G� y[J��Z�;D�&��ڭm��bR��g,`�?,�6ny6ѻ�"F�xZ�gu\X�osh�*偫h"���#>�1�"^&Dȋj�t@7$Yt�fCtCDM�lA��|��c���특ݙ����E��d��]-�`_�(���ss{_M��g��cT�'8����#�J�$�(��K����g�����B�D�ޚ/?�ѤˌZg��"�!�8�<'n��H]gpu���@-ͤ�(��+���2}������d��՘�Ը���4z�z�>�M��΍�+�p��:�V�t�~�s��)A�Y�s�ē��y?	��=� ���0��vFj#o�,a8= h&������j�d�v	�ֶ��S~΃������: @l�6]zf1b�~��;�wh��v��b���<!��6����S�0Q2x��M�s��d��p����Ep��'uP�,��ne���:�u6^��*�d�h��K���T_#n����V�ƴ�9�f������)�U<���@���R=YYz�7?ӌ5��ڃ�ҵ`�]�����i��+��=���\Dq����ep:� ��o 7"�I"\yE$˙�kGo �Xݨ _�$DP�E�웤����%"wD���,qd$怜������Ã�;�A��޾��LY�ر���5�k��A~f@����_��!����<$�/zV�iX2R��v�%,i�i1���n��Р`
�71�q�r#�7+<�?/��X��Jנ���nR��e�u��EC��h `&5�;(�[�����CwsaRG$��Փ�5���?��x?�I����>��eM-�v(�u^�n'{��jtz3K0���wo�����wx����2v���V��s�QxL�қ�:��멤.w��)Ti_1Gek�P@"����Yx�z�	�܇��? �ٌ̺j�:�0�]�pK��TEt)�g�\��Vr�؈��/�B'�����t��Uy�ƀ��+��{�P1+����H?.ޔb=�m��}J�ٿq=��s����M'��oQ���;��]�1�a�l�B�w��򺃏��G�*c�V�'��W�U_����6�-�Zt[T�{�7�Lh$'�0��� ��j.���
�.�2R�N'�W>�a�G��Yn�}曶�y(�#��md�F�P7��.z���:(��YRl;YU6
�����Gs�O��}d���-*Y��a��#6�+�Ctݭ%r�U�3O�C6=��A��*�:0��;��[;>8n}��+!ݲ��/�o��s8�]:����Ãӌ�۪\}�.B|`AUl��h�9@0;"E�������@�Kle0�����T(��AV���AuU[H+Ov�TQ���NT��=\Ť�_��Q�i�j���\�X�d�b#.���7py&���g�Iž�"yK�'�oEBQ=���d�[.�\:�Ԭ
_�/d��+���3�9��_j)��Yh\zE7{,"�UW>�$j[q'^&p��a$��w��@�h���:�Ln�A��$w���Y��%��:�}g����-�0@����i����QdȒ��p�m��^��:�XKh��ym�U��gD�r�उJ�b0G��;�v`�~&3�{��i�	3��X�׶Eu��n����_�9����y�;(���۲�?8+6�+�ǈ�~]�R�r���fNl�Y�[pc�@8��,oiM���T�2M^�T~)���6��7jЀ�zGQQ��O�%w�΢XӲ���

^�7������z{��:�*`\윖��E�U�]�:Q_:͍w��􏻮���M�c�[��ks3�� '!~:��>n���g:!R�y��ҭ~T�y+N�y�r��_B�irf���P��NV8��P�Q��A���h�o�@~x�]��p���PG���� �
���1;l�c��MK�t��*W7lLF]C��P^Y|��2�Ъ��)S!͗^��¬���r�:��R�t��!]� zZ,��A�m�mi��%&�"���e&�z�N�R�m����z4qAOef�	|�c�
2�$>��y�B�p��nѱQt~'ܯ謰 (X�M�#Ҷ��)±��I���i� ���ک+������I�F���CB�F0;�Y����q��_�S&���D��R�4Ii򯁀7x����-AAsz��/��`��D�N���'NwX�B0τ�x_n��X��S|3p[;M����^�#���,�P��_�s�V��Mo�&�Έ��&kmgÊ.c��j�r��J�����m�D�6aRu��\XU��x˱�����i%����B����-;ǟqq���,c]nw\�����%Q+�3���1�A�4�;�����#�J)�Gu���)��8͚v2G?+Kd[�ݴq�&��5I�<.`��exP��I{�R�7E^�� �ɳB�W�vl�U�㖀B��Z�(�G�'�/��q�kt8��XmЙf��J�+�0����E�F�U�gQS�`����=�Ȭ���̏J-���B���T���ū�ч���M�YJ?�����kW��Z0��5�Le��OB�A 4ؗm_cQOy���/2uA��[j-@����\�����@ǹ���Lh�k]N>�sƈ��%B�v������g	j4�H�G���x��3��,"F��0��"����c��d�����Z�$��4��|���N��&h�/�^�Y�jA���cp󍬀�T��^�42�c0��(�@�n��wh�����}�xCOY�ԄK��VU{�UQ�R��
hN^(k֬��L�/�i&RIg1Ř�Rx����2������ �R�^�ݍU�0sΟM#�,}�V4|X ]L�J���0��Q��A��:��Kl0,�i��eA�qu�ݐ��_��'HW<('|^�����d�4���hw�v��ۖ1�`N��E���]��q��xu���-���v+�op�����u�W�l���V�^��X\��$�|��>)�V�~�w�����Z�Iq}ٸ(����:�ߛ��G5&��/������[=�C�]U}�"�
�w�K$"L�v�㎧��������p�@�K��~ҿ�vH�F
�A���\O�s`H"j[�L��qd�n�t箾!6��ئ&��@���mTd�x>�y��S5�h�E36ٞP��h���^ԫ�Ԯ������1Ʋs�ԋab�;*�48��O1̦s�n���=��D�%���{�lYZ)yx���wʏ�r��P�7��P3z�Ò�hλeE�vPK:�'hMK�A�߬�qR��sZ@�)-(W��Q�K�/2z�m�.B��0�H�!l�'�}�K%S'( �e}?���#�u�
�M�O�˅ޯ?P�Z��3��Z_�=�H&�n�� ���9+: �	��#�r��J�(�|��������m-G�a"gn6��E�?��5���۪���!ݲO���œ��{~0E���Ȋ��Ç�ɉA�� .P�������C�����*��g��G�>�%���ka 4D�Ln�,а��$4�Xf�C��iȂ���7�܀lz��[�����E�-c�!�Y��{咹���c�{T�&}O�če_1�DZ��!I0x�E	��ǏOIml6؉=��; `[�@��8��ܩQ��rT�� ����M��Q��S���o�O�n��y���D	�|���@sJ ��2�A�Z�ZD=mV�JBA��������F���metO #���e�j��Ǥ��{��]V���Z��Z]_V�)�5w0�'1����`��1��?i�B�t�t仮OQF9Rʺ�|ܺ�~�SvO>,�lH5���A�~
J�e�jޒ*�B�I���6Ǒ���3��a}�^�ze�9 �k�Ru�'�I|�ܮ�9S?}���I$�����bq��߶�F�ƙ��������H��k@:��!g~�s�:�+��.��E��=���.T���)R^��q�v��;���u���c���p��2��m*�gj���D�����;]Xd��r���̠�9J��$��� ������QuS�C��K������Y�=F�g�
'�ޠ���ԓ�!��h�r?&ay><x�%���xk��Iઑ��\��k[�m��	׿t���lp��^��ې���ذQxPS#c�&Qn٨�Y+��!�C4�,���z����Q[�v����� *!�� CD)�,M�^�'b>���O�+��K��Ŋh�-=����z5�ͨ�{��f��Ր9c���w���R*j9��~e�#l���\v�]��ژ�,����JԤ}�����4eB��{ڃ �^k����XA���� �Z�Q�֜1`q��.�� �7b0�M(z�`�����L�u�i݈�Q}����Z�����ʷ�T<Ι�.����5�c��@ٗ���!�A�p��<PbtԂ��Wa�M��[�8�nrB��Xin	�6��� 2����ڋ�U!L������ޖ�W���+�!���y�:h����uf<���9x��"��d��j���Z!�1�=�����k#�r�ƴ؏Z�Y1V���𯅇�`���Ş5�F��� '�b�ނ��> ��(�U脯U�  ��f!�g�����]��_����

���C�.^m�G?!\�0	�x٫1�/B�����p�����O�%\mw��2d$����US�8���ަhڅz�o�d�
Iᶤ��H�[x4^���}�p��'nc�X���Qy{�ӗeһ5K$1O(��3��ͥBxw5&JI��?���Y������S�fq�&�l!g��O������]ے�@9�Ԁi� ��8�t�3�#Y��������oL4Ma΁�e}G&#�xqJ�x?0�ůfO�s�ҳ���#���y�s���:�7�q��^ɂ�V����O,�Lx�K�H�	^ÊnX���8e~==l۽�'����Ox<.���FLvǍ��R򜿽C��Zy����� ��+���Ɉ��7Ko|�_�r�6^�'ϼ-H�¹���%�>Skm��q��~Yڠ��ʐ�o[�!���#�0^�|�L�PSl=ܰ.r(fC�ׇqQ�GW��֍�����8�
�Bhkߞ6�?%����["��z�;<3`e?���k �%��'��í2��(���:`q��5�>��b�!ŋZ�N�
�'qoR`�!��;|ו��W�:(*�\�h��j gHG2d��R݀�����b�+�J����Ö5��������G�j2|�G;f�X9�tDF�^�L���^�#K�ij�J�ܬ!M��>����3���֡�0���$�G����9�R�.y�
�R>�$�Y�i��UI�nz%
��H�u���6�$�v�x~���s���u�S�Ŵ:�N'�+�m� �
cC�<�%�|M��X&^uZ�,&3�2�� k���])�U�jn4��2zw��t��8`28���?�4������o8]�q���vT>����n+�Nzډ��ߍ)Gg.>+�C�������E��qr_�<Y���Y�e��q�.�U�����A}������
�2BWt�f���q���e�7_ԻP:^�hS��PjV�ne��$��{�Vy@j�F< m4Rl�����{Z�kS��A�m�����]�ڜJ�1�t\�7	�o��Y���?%�o�P���}_�I�X���Ӂo�w����+߁wJ]Y��2bs[�uJ��~А�{��p&���xZ##�u��)� ��`"P�y���.:َw��b�,&#���@޺Ĉ��p�_Ȓy%��2H
w�/���Np):	�ٺؠ掾���2tb�DV��T|��f:�S�AXO#�D�`UDS�w`cuP	D%�K!W���Q�"E=x:�E�A��^�ry$��4:���H�0��B`�.� ��n`k�!e��\��a�O�+k��%m��ɚ��nU��?�;���i�8��M3�����#y��d�>f��3��	��S�q�������PP��Ml�(z��/ �}�I����L�*���Դ�!CˠOo����ec��T���P���R�1�`��{��`Fo��x�b$�'G�-�}�c\[|�~��¯+7%��lc�̀�	�Cؐ�>u;X�Hd��J�ᔙ�>�W�M�e�6�5�:	R�z�8�2)�8��z֑��$c��7�@��h��
ٷ~�b/+�͍���w�$p�G�pee��6�"0	�CAE/B�H��ͼMs*A9�2;��,e&-����ݺ��N�����5����e�9�\ܨ�'O������_#p���i�")Qw�"�U��_�6:�gtŌ���3�k�xw��&�/�� �e��ڞ�����̐�d� +��&�����FfW��JoGA�'�%�������rk/�廨Ȥg��1&7��G�SCTB3l0\a{�-E�T�XyX0���~{���V�_n��z�%3��G$+xˬTc�x��z����
�doZ�9���Rh	}��HQ��B��B�P�h�R�!�ά,�wo?ǂDdYX�Eq������ϋ����<!Ʋ�𒫞j���ᢒ��1��H�^��8�`�^ꖶ;�:̊��W��	�Ϝ�M�lL�M��ߩ?_2�[���q��6j�b<��`p��AX�v��%!O��qa�y�|�{YGCn���ݤ-#�)�����z�+WvJ� `7�qܨp�(Sɺ��B71UĤK�.n�F&��5dd-�8�3�y�!���Ђ%.(�.l�)��3�/r�����	���Y�Z�WYf��젊�������G�'>�DEl�>�w}ߪV5c�Ѷn�> ����L�T{Cn 7+ x%ϝ?&<��Ѕ丁�܀��	b���(�n��ϧ|j]50~J����z(ب~�K�q�/� �#�d�4���}ߖA��
d!�2��0�Qy\���^����tM6M���k��L�ȋ>Va��]	3��-e��Ĝ`�2�]��I2�EE�!P�yl�K�ӹ]�S���.d����\��1�6�WEҚ�,6�I�aR&zY;7X�G��j]��%N	bx&�9Ɠ-��ql5��f_������SM��]�Z�c��	u�l�Dk��MBf��g�n��։��g�̄1�����4گ���b�x	����q�K�K�Ǎv�Q=�puCq!�+y�B�����]lx��F��������Ǒ�)�>�[�"����KX���A��[R�`��C(��,Ghސ5[�.�	�o��D���Z+ű�����	 ���l�Yef������pn���HY��vI*���p�U���~�$��\�
���GS' {�T7�3h_` �L5+�ˠ��������a[��������V�`Ur�3;L���"�gQ�%��y7w3|z�^�*M����(��X򟗚��D�#�;ϕ�b<�;�[0b+�p�*x��ҁE�ޡ�DF+T�"2U�����`x�e���P�w�dӪ��4��R��# 72[w�R�U�j\5b��a�,�+����N�T����N_��ݑŮT�E��M+�W؍v"�|-�chsX���j�)IbLB�Sj�x��qb�
�~�R�����~�ϓ_�h�A�S�n��7�a &�s��t�0�:�vK1�-��D��F\ؕ^HG���,����-~I6�uX�V-;��R](���>���_<Kf�re%���:/�@��.^���oɅ�6%���U�����������h:us�D��0��襜�n�E*N��0��Ux�2Dբ 5��}��@�����MJ;�/��u��[�R��Wiw�B�}�E��O ��SNx��������Pv��;�ȋA3e�ob/�!�R���
�&-/��;�5�+�)-�\u��kOW�$N �K�?��#L&t��@�St�-k���ݤ����am�{al�w�&��~�+7�?�֗�s'��Y��@3Pq��i*�����e����e�K���va�����M �W�$#�F��*Μ0��J�	�D���3Np:af]��{�0jg��~#�M�(�l&q�[��-� ���82����*m0���Y�4���G�U3��А*\S�0풮��\Tݶ\?�����zߥŶ���5���>����5}�Y�������6���t�+G�v�3��^Y�G�Ӧ��%����K�=�cpK�_�ӟ�h���yb_��Lb!c9��𙎝��Aї����V�ձ:�<t����y&�[Mh����K�L?�UW��L�I��=�0�=��DIR�_V���~���:�y�N��.�Y�c4���=�����'8�R8��\n�M�����q�����,�f*~�oq{H�(���@��e����Y���z&3\���|�N*�قIU-$5�@c�Ţ�^�n��m�m�y6E�T__ߡ�5Q��e���7�q���h�y���E+��)Γjcpg%�^^���/]=E�x�6]��Zf��#v%9!$o�R�&��W�Ip�1�����,9o
%�d��G�4.^�vq�>�e0�a�S7_��l�b�/a��0�Ɋ�\N3��,B��oy��dx�Hzxn��=j��Ъ ����)�hg4�)n�����s��K}c�d��7C��bS����Lŀ�%�9��3�1=�nS����(L��7�u����� 'jiO�#��`��0Z.�2= ?���p'�Y��s1�)��ɇ���ꆼ���'���Pۋ�ꇞ��C��A�5���=���'0Xf��}��Л4M�<�T#������I�!;g���iv@�z�  ��(�4�ZG��%�7+���n`���n3q��h[�PD5_�s����mlXA�ӓ_�c���b�`���ퟪ�4�Á��e�ū5��.����C��Ex�q�(7� 3��I1�Q	: �;�����F�2��`��!?�����wۿ��Dod�C-[�Q��R% ��R�A��Y����0iD�F���B��vjO(I���t�J�� -A��x��
�D�?"�]��%��S{<
����UN>�;Q$q�ELr�.愰E��2�#���^��$\�`�pÂaLPm(O�F}HGh~���[����@R�H���%��Ҝ*}���o�@'98��p}�ٱ���:"x{�w�NK�E%�2��H�����`�t�jM�ZwE�^������m�F8?�3\�{c���sPu�hV�iV5o̻�E	n<� [��y���\r����L�D��h�e��.�.L��4ȥC��#��Q~Bh�`��;W�䕑������ [������ʩ�Y�k��$�t�yK�0kc]ӵ
��.�tV����4#_�k���*6~���,�����0*Y�Z�8�'6Ǣ���G�T�8ڿF?�E��,����9a���p����i#��Espfx���i�-�4�	{/g޹K�L��l:�����Gn}Ւf�JQ�mV�c�~���m�E3a�?6�6���B��Q�O�A�)58[$��bG�a�=�˯L����~��1�Sѩg=�3�ƨ�sg��y&�0���˟Yn�җӏ��T0���T��/�����/�d�V�`���bMfV"}s�ҿ(ԛ�z8�jai��~Sh=��:[s��Q�'˷
.U=�]c{��Gp8�Y6:��X��1�v@=�P�u[UgA�����L�g4z���m�nӤ���!;48�*;j�,�m�؞'nF����QE�Ge�[�*�TJ�;�T�w�h��+��?�NQ�Ǒ���O	\n*��>��+�^.K���A��s*�|��ȱ�O�;�]���r�A)�&^��	�3>�5n�hhsD�l�4�{���a:�8��ڪ��ܜb'`y\W5U�&��q/�B�JҮl�7���2@��1m��酛O����%�˫�k�$��9~RH7��Ρ�Z��Y�'f��y��*I˕�֙�9BÒp��.�������	8D\-��<������ u�����*Y���T�cs�!8������	ݜj+ξ�q?�u[��K?�џ��aH��y`\��ez^�|e61y�"�R���d��҅\����]O4���pf0OPc�Ms.pz���@�ɟYl��{R������sL���U���$��M�h�Y�V�Ynpb�ym�c���J�Ю���'���r7��8R�.�t�&�bs%�ynh߈m�)�D+v�#��e�p<�P��Ȗ�E]�G���v,��U��x���)4�]}��46�,��(��f&���f�zN���":��,�2<�b��u�⽅����u���HƦ�`�r����n�FZZ���y�ĭ�;��Bz�njNUJRT�����i�cGo�-��NWt�l�C{X�j�1��	�噣�t��_������ ����,*ea���[P�����\��͝ݓ1d��j>��3|%c��ˊ �
8�_����Z�j\����	����`)1��%�d���j��������IL�rgB���u�R�����a�
"b3�[�s��z�V-|�}�z�~DΨ!i�|���r�Xm�:L�!��ļ������)�k�)®�Ni�DZ9/c�/�W�Gy�{�:k��w)���WWKP�i�%��Yg=��.,�5��X�|���ty�q`��W��2�c7f+�9�:�Ӝrd�ܾ8EZ=��Pl���L4]��&̈���vC-6*�K��e�� zvX���V�����a��M��{�H�W�l�5!�6�r��_��
^��m.3��|	��գ�uv��L��Y��	S���/�@U�>Tb큅8STG��(G�S�1'k�{����b�a�[�C���Ɓ�Ԍ?�-xt@�`��p�/~�B�L�&[v�q��=�������&b�rS�,�م��"U�I	5t1/d�n���"VG��������8RՑC�؀8��e��
�n[y-U#����9/�I���2���L������&�+�C��Q��"�Սv�F���4bg�!��*|)�!��ܔ��%�R++�aRRT��̷�d��Hø.�/��n��hqA	#��HS����;�����W�09g�����N� L�B�x�4M���:`9x�JR�q����ˤ]�V����i�� ���w�é*ép�iI
�=�	���N.3	Tqnn��U�G~2NМR���C ��!-�l�ɇ��ԙ���
I��:oJם*~�s�1���������Iõ�ʁ���=�O�"���^����*�k��F��6p&I�m�˭�;��S�%�;�I�0�3-��2�>��s�E��F��A㐪*�l���Gq#4��@�B�RI��3C�Lӎ�*ɺ m���OB�㓍��<Q�27�)��=� {�����P���.oH#�T��/�!����1{�/$hG2³$*�Y��f�`���(LU#�16@H7_�xgP�).�������ybǲ�?���ԁYewP�n;,�qZxS�1�5�a��uuH]�yV_kǼ���-�|�XZn����p�S�:J}p���U������jz�Á;}3)�`�q0?��}k+���WRx�͙�	�,��O�����DS�	J�Oۅv�Fe���E��t���s	)�R����jƟ]��ͺp���qv&"���5ݗ3�h��~f��ʤxq�d$�e	OO��j�X�R\5����n�GW���]�����iJ����7���a���d3�7��/d��]�F+��c^0dK���Ð]p�i��PM��j2=���k���~��X��(�a������6��o�;XS���	5���ja�;�H�	ss^�O@β*��.�8	�C:����8�3�fH]1@�%:���� F�ĩf���%��P�5:o��S�T�`��5�|�-qѝ��&�M��I��w�)�����[�+4�<�2���&�u�����c�Q��ػ�~<f����Ri�K�Ɣ�Ὥu�!���*p�*�v�G5�T����)Ð��R�D'�cY��ێP�+��G}�|���H�c�mo�DZ�zc�+d9���$�?�� �!씟��Gtu�t*J}�3%�7%��"�C�_�mQ�tm�9L���O�;�6Um����>	�����ݾ�	��:�Q����W���0�c�b�H���f�s@h�L�T)
y�<SB��D�0ް��߇��+�J�l���R�w��9���bZ��̻w���Y<H^�$�����oD����'�sߠMg1;Y��;�M[f�}�,�8�JI,�+����`	��}�M���m�!���a1,�q��2��BƬJ����C)H���'������S�ݱ������[���-򗣆��^����w�O��>�' �E�����i�!IG�MA� �a���5��� ��Qn.H��
��e��f|bu,=~��7��| ���0b� ��ro�����7�>�b�~k���*�f���w�~��L���Z�d��}ښ���*q�h�=����	E8OJ(�g����QHs�:!p�H`ݏ�<ʍuF���E�m�*�a�-��<k���C@Q�b;��vn��>JU9�>�f���ڥ��T�"\�DD�y�f�čO~���Q�<�{���-q���*�B������Ѽ��e�oz��ltY��2��d��6S"�o4/]�[�&y�$4U�%-�~qM~<'-�:;:2&�V8��et>�'U���_c�9ё��7kӡ��#�Њv#굷��jK��p���,�w?�D�g�T�OQI�c���ѿT-�_�P����'Y�� ���'og1���ϥp�Ni�KS����`R˯��L����J,�  S��@{�h���9�ة*]�{W	z2,sjq^''o�*s���q��-�k&h��~�Z��&>�X��Q�O���&.T��v45m<ah���֒u����S�|�*ps{�b�o�\Cd�L{7?�oB��(*���[��'�@ �&��=�\=�J�>���A�����2v�z*�|�m��eO':�.�~%��A�>+���;&�g�LgO�.q遹fi�-g{D��{�g4i���ߤ��%��)@t�1:(�'�{�Ԟ2���Bm�P�$�,�E0�o�@+�_U�
�s��+�mJm�� N�n��/]h��u�5!+�l�pVe�L���:�rm�Q��n�fD��E$bV���!);��hr-����K��gC6"��� ��Q/UV|f$�ߖ����t1H+��C�>k�����\d$��?Pý
N��������#�l,}c�gx6Y���
�8 {�o�̏u�k(q��nƚ{��oYgߦ�`�NY]���y����@AG���zBp�L��(R�#'8��07��/�ov�.��ޚ#������9�d��{2-�ONe+ͥD�O钖S%� ��B�VHY!?,���O�����>�"��ԫS�Hx��_}Q�e�E��%2���*��+͵�+��53t11̆N�Wj����/&x��A���/*⿾��갦�_�pY�wF��5�S�{��"ʲ<�V��_0"4�?��_2���(K�a��w|��3�4�SU�6Vr�MN�Qn�Q�v�c,�&�)��Ə������4��j1daHs|���S)�3-���K��װ�T�a����������T4�h�}�%��ORJ�s���Ӄ�R[�1I���Pʙr��)!O�Y�5�{�����Xٱ�7{���x�~'�/���xB3QRK\���B�@����"��ۉ�Be�k'�I]�La�;�!F������?[�cY�;:�bjR��0�ձ����1�E���JML�H 8����Qd'Ҕ��_��-ys"�P^�2p^��Wc�ǆ�T�uS��u�/�U�G$Ԛ�
ʟ_�~/A�!�?1k�D�|�'�t�֪��� ��(m�u�cgC�bG_6�	iN�R�:�v�5��T��*��C�uӨ(A�;�:Z� @h�0]Y�6 �����W��M���PcUƣ�pg�6���)��m�4l�ċ�q�S�}���fA�wޠԛ��1�`�ʬ�M�*��$;!3;�>1�Wǳt�-���.�U�._�F�j�!q���$��"؀oVA�}R����+�f�^�]�TR�t����a�6��v��v5r
�ܩ/o5TJ	rIF|�6��D9�#��/�>3�eʣ�3�K|^�s	��\�V�ɏ�wt�X����L""�E[�j�FV{mΛ?.T����z�1��tX�Zr��\�U}r���?�b;ȂM����d�d$'ģ���p��b�f�J_��\����W�k��ګdӆ*�f��Z� �u�)�PR��p�a�C�7�t ��������H�L���x���M�f�=��0��ߝY�!�X��3
/��1����Q�a��C Rt��m4/I\ aŊ�6(�(~³��O�+i&�pN	t�Y�3��C�<(�0�Nn�?e�����4�ȤQ�"�IHXN���U�w!nZ��H�"7&��KR�>Mi��V�y�a�4��e̢���O,s���[�d�igJ�@�qP,���+�n���('�ڸ��)'�.TK�}g6t}R񥖟6�M�����LX�n�n,��\i-���R+O�f����7M����A�)��7�<�kn9�[���F�l�bĥ�E	�LKJRjH�U�y,��Bod�]�Q֤���� �=��b��v��%>Ǩ���Z�n�Ԡ�|�@K�p�SbmPK�RC#���y_����ϓ�Z ��@A��gs�E�mڗ\��1)K���
D�bò�Q�8{&]�n�oi��`� Jy�F��Ϊ8��u3����l�P��j���K;>p��̫���c�t�.#];�����묠�P���!�<Ǧ���;	�(�"�(��t�n'�k�V�B_B�q���CnNY5'���Cʾ$چ|	��$����ժl���OO׾1�A�� `�^[)®��37s�j ����{a�����I��s��X�o��~M�Ɖ�� ��ݎ�z��s�,
OP��]�,,g���iM�:��M`��!<-;WSn桏�CL^c�L���� ��b�7�F�NE�N���\Nsh�y���,#�6��J�?�j%$��v�{\�+�yR��G�pN�h�xt�Cw����v��}�������	C<D���B�

8�CK���I�1��X^�<��G󺰅��-����X��F��_~�௭K�k01�9�8}���c�Iq�.w�ά��nу�<�
*�;a��Q���k����K2��$r��\����w�o�YB9j�_L���E��4�	)�9@��U���o¤#4�V�7����R7~��	[�mӳ��ԡ��F�%Pq~7)����o���'��Cy�N���[-j����Ŝo�����d��s��M����U��8����۫B9u��.*|6��5"Ń� J4d�u��ս�T���<�$16�����Ru��e}����^v�p��%��˩<χE�㊁��g+��0���H��|��j\/�gXg炽�<ٝr��c��T���͜'y	��7f�x�q;�+LX*�6-a����=r����O&����IZq�2p�B��#��fѻD1�X+3���z�Ґ'dx�C ��1xہ�rw��Йu6j[O���ܝ�T���ۙ�3���C�yM���ܘ��ڡ��~��YD��������rCޮ�pv�����
�v���{9��NO�b"3���TC����%�!��p����B�O4�P�P~Hٳ��bg��I��λ��b@��b��(.V�,#;Il^z�?�6��3o��J��h�7phw�_r�uiDk�u\��Q��<�sC�v�{��p<��vl�@��7�(�)�޹ו�N�u�������Ɋd�Ψ���AHުo��K���;��Lxv�B� hPS|�J��3{���">�O^M�3<,�5����y6��-8\��\�*8�xP�2J��/?_�@�J�� �O���H��f��t2{���,:�|ţg�*ilO%�:Y�b��r���O�&pG���?!��J��st����>�pz%��H��r�b����u���e��qZ/Ȓm�h�	�΍Z:Ɩ-��ɞ�)���V`J-uF��_l�}��#Imf���CB�g�d�0q�-�Kr��Jڿ:� %j;aҖF;�4���R�Cr��ԑ��9V�Eu�J�HlFR7(Ij�AFUr z
�a�mO|�����Ny�����F���4��e
�匕^�`։�?�N�C��w2��<�Z��cs%rJ(�C�Ө��/ym�F�&5�o�Q��+n�|�[[$9=��+`n�U����d����\�`��"�̸j ��>Ƚ�	�A 3��UkY]5ˎ�k 8��8R���ˍL ��&y�d�P6�J2�¥�}m.~�^��K�5�R���� �����q1 X�Cݧ�I�*��힋�vȏ�-��������UmN�H��E�l��,46���տv����~�l1<o����i��֫�Pe�n^ٍ|��D � ��-\q�|�Ɯ�=]���kV�7�b(d �r�
�ӵy� �v �7tȊ�l=����6�pߤx���� ,�Cؗ�-�_�3��ؠ���z^Tl ���Y��.ʋ�����o�?j�ݾ��GY�*C��dd��z"~"	ӟ���(��?��FW����y9�g�SA���nc�@������kͲ�lF���;��	��Ns>�X��VC�j�}��8�Iʙ�k���%�DOj[�U^��c���]�6�: �c��e �3����Y=az�49sl,L|�����8�^���8^�%	�?�]D����)�y����Ӌ��$(�[2��q �;0�!qVb,�Ȩ�77#���,�f�]�?�Y�4SYx�|��)�2Q�[Wp��}.xX�Zҕ�=��n53��	�/_�3��ȭ��"Qp޾�?/�3a5�%|l�吮 �I�%�mg�l-2W�" �6[�g�gl�����a�;xQ���2Z^@nbV��}؍����B�[u�v��__�[WIM�X`��"Y�q7~Aa�~Q�I��h��%��Mf.i�b<�2��/��Ҩ��.���ds�^{架�e_[x;�
SF����L��V45�p�*QKrIċWx�ê8?���m��5,P0�$�n�j�$Z��F	m�
,�����oDϙnU�U�Wo9��;�-4�}�B%d��I����>[ ����t�)��Q�M���g@���j���� �̽So�y!Ӊ�Yr$~�&�lDP�A��s ��'��Th�#�J�7�GĂ`�ߝ@7�L�u������66�1�9���R�*񇂒]2�:��At�O����Ã�w�{�;��L��J淄��Je7�W3T���P�C9�@�4�	 ��ݺ���
%�����I�[���5-�Xfe4B��-���J� 㙩&�Z*K�TF9F(��)4��ɟ��|@�lM���3�c�Q\zP���2���AC�$z���ӯ�h����JE ��k�� ��"�,��/D�7��`��+~c�{6��]��i�Q�������ͽ��P�v�čHW�w�ވ����h%��:�ˌ����B�;�."��*{����%�Sj4�C>��E������
a��q9JLӽ+�'��%4���ͻ�G_��-A.ר@���w�a���d.��ǳ�n��t�Pͺ����H���� 7�جs�%����G��IӁ�.��$��k@F]���a�^�z�xw��~4�;쪆'��B�ޙď�;���s9w�k(L��a�?� �o���.n�mAy�$�Z�U����3���U+j��G���p�Ǟʗ�ʕ�J@�M��f�3�F��}d���ݺ)9X/A33�ل	�B�Vx�A/�1�c�/g�#�.��m̻~�^	w��5K4=)�\7��
�9*pWt�(��pa��d��_2�� v����Hî���K.L�/WدT�v�Q��k�ϴ��ݸb�?ӂ�Y � j�h���H � N�oF�6O�%�s����{�ی��b�9ƭ-彃ru@ՖW5r�sl�\�����i�4�ē���nWu6��%�}nr��x'H	~��+T0��>��Qm;����;da�ʪ�����]=+`E>������5��|j(�Ħ��*>�74'��
�_kY�'F�B���B8\�3�i�����T�|�nr|2�ٜ��M-�3w$��)i#�^P��8�#�6�rA&X�~�G��{��f��.7A�i��	�7�~�0�^i�?�`���x�j����`Yi_�ݲ�`�z[��� dڛ%�%��È��;����u�a9�"��sPC�s�]x�HK�h:*����R&y� 
v�«�JM.�a!?�j
 ���{'����߼*HZ�c�S�*'���@c�ܐ���_���]m�}�]��bY`W���_�p%wi��%��}Ѓ"t�y>�G(WQ$M��5�V:�fd�!f&����{��s?�Sï_KN\���l�F�\}�k�����HNo���y��� B�5H��gy|ҳ��2k�mL�o�:H��fɯ�C���fy'+��E�ka1=m���1į�D�!?���X�0��6&��W0�>����0��Q���l\H�8b�k��è�ݳA�67t>��c�ܖ�V��:�z<���qP'��s�R�a5�/�q(�Ac^^�gכ�T�]{�oԥ���\FA�+W+;0�#��%g��xd�����{�ꁂF�|��*
!��Mj�R
�e�+]g)S1".{\�0aq�17�}%��}r*
��/�(�G@�|�~��e!��Ӫ&n^��~1��gT�)e�G��~
о��<���,�+��ec�6<H�W{�.M	���r*��88�4D����9WS7��o�R�òP\��S�r}�q�}���ճ��'�ݒ��B�W=l��X�Q@is�\'�,���0m�%A[)���*Ӷ�|��şs�rf\��qX��G�����i.6%�q�=b�.����dˎM�G�
������<U�0o���l��<�?c��:Rq��tfq�D��ց��ȩ@ x��/�j����XIt�26�L�pjw���;H�5�ûV�|?6�į�#���3X�%y�����+�B�ȴ*�߄@��XS3�(#A\c�� � >�ER��8}8��i��.�qWܓ�}�攀���Ӆ^ğ:yB��)3%CB����(�'qG�:��^��I�\5#�ے�	W����RG�S`���_=���=�__N�E��M���v���y.þ�%mʃBJ7������TC���O�0ĕo�C��(��^�J�me��qJ��j�v��x�� �G<T���UU�A�|G�JJ��B�tF���J�YP+`yU��r�k��XzT,	��\��.7h��w�93��ӎ�5'�X ��v֋GD�nSo卩�Jo�ĀgU.kWc�7t��%A��Uۼ̂�n]V������e�v9�Eb��ڥq��Jz����-��#c3�<���N�φ�b3��-O+c�k�s}F�z4�:��w��
�/Մ�@�z\5:�!QgA�k@*7:����s�)����m�Cz���U�FbҨ/��z)J\�?"�E���^o��ø�*�����E@~��)wx�r@̒�������ŴZX!j*��-��g���{v88�4���#�l��v\[�����{z�L1SO8�v �
Ԏ��gQi�1��1��U"�mpv�>��E�V3�W���C`���S!�eY�[��1�1�nfh\�#o�r��2޸�ac324 = cX��"I*s4�KD���~?{l(2ѫVdZwS�E�#����s�C�x?��?u=�'~d����~b���Ϩ�ڂ���� ��ɜ�+�S�i��F�g��h����~톔��_�R��Ѣnڦ��@��л�����ggw��1<,pS�=��	�T�������+`x�iۯjG��h���i����SI���M��05���Q�H�U�_�M3�Yڷ�{h	���)��2d̮u���*h.ː��.qM�~H��6]�*�<b�����%���~o�c����tx�&���co���So��%���C���N�R��تrD{�����B~!$���bUy�ϋ�4L("?������_��}Rf�������yQ�HVX�G&_뿃eÛ��=�Z����rl��w̻l��NK���
���䏓ׇ#��|�vR�ۤ�O��7��rD�Uŗ+y]�_B|tO NB��dǕ�����|_�2A���?���Nt�ӊ��#� �v�-�|��^hY�͂
�=�@VN"��c�N���{���I�>��6M]޳��zQ�{��,�Ű�bQ@����!邌���p?�`KGj��ܝ�9��7nR�!�`+�Z�����9�^�m�����ȺR��;�#�o�C��>@ ���3�OJ^�O�ˠ~u�� �gK˴,h�W�l~� �w�`[���Γ�I
0>�^�8�J��k<"�Aa�j9�oBCJ���qD&�d��?~Um�D	�/QL)�)��<G0�x�7��c�6��=	��]�:'v�̥�@^@�3 ��ѣ��d?��_�I�+~d�N$k�P�$�r@-,JW��A;b.��n��,r�0�	]40~T7X�/E��&��y�v|�ɰ��o=��	���>Y����ԯ�Pya�2in@v��7G8��sO�S
�9��m+]9�_�av�0:2)�ʈ������@���s�����k%_c+���k�M����6�3$��)���"��fB�Oش(����Kw����:(����җ����!�CE�!���L�0�}3��4l�
�k*�k�g�1ǭ��9*a\k������ F5�\5���F	�E�����F�f�ȺIAz]����1�� �o�v^!g�]��lU��&��%�6�� �gxj�W����9��v�l�whUpx`�H�ě�Y�ݨy�� �1{�l4}��uf,~����r�P+e�u��dh�~���ȱ�n�^P8�`Ƌ�a��� �,5A���[`�I#��>]@R]F�����Y�4��IBm�S��
h$��s:��O?oؼūa� zq��R,����:��<eף��]�S�`��kqa���:����dt>����c���eGל���'���A����)xO2��Q+3���v0��3S�3Ϣ@d/���c�u 2�`3�y+�38�e�,���ә�'vJ��q�dS�/�[�\]�\�m���4��������lB�|fb�l.E��AcE$UM؂�O�����)�Uӎ��`�[!�j��l�m1��p���B�T�;�({�:z�X@�0%o�{���	�҄�G����Ɔ���m�C9�G4��ߝ��liAc���.��%#Ժ���B�Þ�
�}����6Y[�76�Odir�* P0��C��|r�&xH�;����>��M�<��^�jw�c�0W������=���'�k-��G'�}	��0[ӕ�|&��ۃ�(K�#���`�g*�q�q
�v	���Cʔ����8������+�٪����wz�x��O-W�Ȩ�e��
v�������/>��+T�2����:*�fJ+�Z�*
.���ݮ������$
�aV��!{�|��Wj䩓�$ܶA� �⸙|j�2�;�!�.ȝI����y���\�iWT��[M�U�W���n]abSg,؏��iV��%'��>���Vi�H� =��]�mC��͕�_g����TG-�#퀒d�o�'���)+j��9�3����\��"!�o�,%=v�.�~^�w]��{s�;�M��Z3hi��x�y'���d1ܔ���-
a��i�nP V��4��S8��ir#t,6�,�팎x� �S\A�;2��R��O(cME�O �\��3���Q���c��� ��=��&�n�%�ˏ�E���M�l��ڋ�O`��B�{VJ0S<�Z�&�U��h����ң����vq��`���ׇET¶p%�p�{�;�P5��OIhb�"�9e��Yu�<!����7G��d�k���[�����5��4�r�YRɽ������0K�-����3�.C�����!���bm�61^��9Łx�O\@�`�����ʒ͒����c���R��U�(i�t	��Ow�\��B$�YR���)������D��̿:B����-����%zORļF�Wy��_ID-�/ȓY$��㸉�,)(f��(*�J���;�R?*�Ԓ]Q���'��㝌�[d��<Q盇?^,�&p��^T7��O�O�x��O5�/Z\Й���.���Cj��2j������	)c�݌�W?R��L��K��2U9����7�2�r���bC�1���y��=O	b�f�Y��	��2f�������[�_.p���2\���d�/(�;�z�؎��D�W���ֵ�PIJ�U� �vV1��Z1����F"�'TѢ�j�KV�	5����x �@��OID�����"*s|]�#�E��R�:zh�lb��:̒z��z�fU1�a���G�`ӟG� �V!��6��K*ű��DQN��;v�,5�	�	�4F����	��g���E3y�i��UE�y�T����sԢ�G��+�<3�A�Z���ka{ۉBH�|1lmP6n�����l��x*�L��'��dN���6.��iIrA^�e��s��A;������KB�Bk��t������kT��Xr3Tm��x�WOS@��	/uz<׼��拜�{,�
�]C4쿮w�9�m�[w��MI\��#�.A�	"Ԗ.�^?-�eq�OR�ơ�|�����BX���8�qh�~�vEa�^�2`woJɬ����-%CbVɭ#�e�-�*�mvq �Kϱ�o�st��%���ח@���AԼ+��YGr�=Q��F��ۤ�Z$�E>������Yx��Zʈ�!@���S2�G t{����ⶽ���c	_Һ�d����;���.M�(�7��Gd����x���w�h��A�x����J��fOr��x+@�(;|��&p�� .YP�S�-��|�^:��ܷ%����1�|l�| 2�h�<���آh��Nō)C�D�>��b��{p`�n]0�@)�>��:.״q�4��V�*��f!��|b�8m1
ăF��ٹ7�v�&v3����5Y҂ ]�%���Ң�	�O�~R�Ϟ���}���lڙM ߄A$�h�&��*f���7[mM�Y�����eN��X���^0��'OK�@E���l�i����޸=W?�����0�"�1��vv-N�!b��`�N9FGoho^�?�2�1�rBP&c6�5�ܠԱv�pA�%՞S��AU���~z��c-���u��y�d_'[0�	Ed��*^�[�������4��2����V�5�^A�$�x+_L�= ���E�~�� %���L$`$��d�g�:}�a� �i˘
su���:�Y��޵�W����%.�@����硌5�:.l��N��,R�{,R��k^Q��%�\�7mk�/;#50-F���͠��j�V�W&�'��g�w��f�G�ܨ�|���$��[>Ú<���R�ṵ��X���9\0sx�l�)r~6x����;�@������l7�^��w���v%E��I�Ġ�Ƨ��Io]mgCj/����#YL�<�G���v�ۇa�N��4�����wU�}���� ��3��S�ݢU@!�)��R
�ˠJ+�������ף�K�!0�2��0�^����b
Oج��2�J�K�_�B���s
�>�;�-ג5��FhX{
��^�u�b�wt
�2�	�>������ QM('W1L�|��Б�/d3�B&��}�n��iT��d�v��V�8����\֮�(6���TB|�RW�Z¡�����G�g�%܏��Ůkp��|�l<<��߿��=�ǰ�t��ը�J����ny��!k~O�\(��$`3.�iT���D6��V�F)�w��{4�G���rOUX�*�֔4�|&�����"�4B
��q95�qBg;wjt8�n$
�]�ʀq��Q�n9�M��:XRrc���V�#A$��T�i7�zBҴk�]�Q�n7H�tt��2��$�tW ?�6�d�%�ctwNj|,@J!Bߧ�j��	;{�>H�Ĳ���P����`jh���C\j<t<p;hǸ�ԗhlNw�y��������ˎ�%X$��`S����<)#-)����Ys�>�%P�����b������XO	X
�0C�Tose����F�j*�;!�qc5���@a�]u��Npsr�[˴+�ׯCɘ�;���W���mF�	,��[HМC(O��H�Z�$�f��Ե����Y'Ou�������׌���7���L���& j����~"���}y7m��̀�#b؅%�,EnԱd&y�SD"��.;���N��u�j�`���&�^�fa�9rƞ�Tu�匾�a�#f��^_]����M�`�t������$݌Ai��p{�����~'�ɃS��b�������P�B����5�3�{��t��m0����?�ߧW�N dV�Y�� ��0��EBJ)����Ez208QW%@�ɧ$�y���M�,�m��fn�x�5܀�¤�?[֣%� H."��[�U�`~� 1�E�����.0b� G�4��p�ow���n�"��׊�Ȃ �JU)	�Q�F�7.�|�YТ���4z:����jH�d�Ts(f3���=��f��sK�mȓm��Ӻ�J~�6Mje�K��{p��Ѐ�lkث�-h�l����?g�
g��H���Uf	_Sɪtg�v��yP|�N~J��q��	_�[K��Z��s���U_�v�C�>oAT	lX��S�Ė����LEs�\W��;HxR����Ic:zwl,�Z����G���^L}]�jq����JK�)���9DY�j�g�Ц�ß#���KTСK��ӌД��2	W�g��Ic�ۈ7�����|V�8�r�#<~ɞ��u�ߛ�5K�n�����H�Y���T3�j�P�S�������>�W�L�b��l��^� ����YV��-�\B��VK����ſuY��\�)-܎T�P�
Nb�w�=��O��~�j���Z4U�,JMl��6g�^]^sX�y�N�F�a@�G�c���e��A�f�q�Œ� V> k��T����;�r�����;��Y�w8 �m����觴���&����%?d!0F��ð�٩��c��8?��� � 	Cţ�^&4�4�MlY��� �('v���#r�N]o��B�rč'=]�VO̟��]f���JbG@KIM��0��Y�{js%�TS*��r��l�;;Шj�2}���67�.+۟����$"Vm%����V�{��~�(��x��7�p�z�������q��&%J|#�"��q�ݤ����ɥ����QuU�y�O�1�-*Y�d�^`��L�K�`�	�H��78�Km0Ur>��
�{CV溗$�,�/k%�|������XP����W˸x�,:���k���7ݝ�%�C�"�����h�xD��AFz6����%�f)�o�iyZ2�̗|�tX�/N��K1�n���r�.x59�-L�噙�o���%�\�r��z_��P�l�񐝠��[)��MC�BB����
��mq�",���z[#� �0�bv��b'��x$�ioO%l.�Y����L�0�O^���C#��E�Ⱦ��/�(;�h��@���ޮ��Z[����t!��Bhӷ-
(?d�>��������a�"�$B5��,U݃6²T3�5B���.K/��sf���̮��t}~&�Bq�����be@_uV2�jX�%X�/h��n+��.���(����!$Da3n;:��/s[�wrm]F�/I�NA&,����r�we��h���9[����}�`�S��mZ*�_;wj�1���7n�]h����G�]�-�l�)�Bf��]hUy��79�l�#���6i9�BX )�Ub�cc�k��a�Bgc+���TD*�i�Bv��K�������}@5���{!(���Z��g0�I�J��q�Z�/p�{��_K���k��{����k�����n?�0��!/��[D+w~5�I�>(Yq��j��	�	;(�
��g���E�Y��*�$����	8M�q����v��$�a�,PsQ��]�{���l'�.�1�����w�C�e}L~%Ù�L�f���k u?���$���������4��H�s���ү����ݎ�X=���|��Gkv�i�fH2��*T������{_"f��VH
��w�D��d�Ew/a�/�O��&'I�i����}#��q
L��O�u�Mŀe�5��j=��6j��Z�tӏ�W`�`���_�2�]���	���ӜF�������ffB*��/�uK����HQ�:�MV{h�z�3�tx�=�u����ep�A�Z�р3h]fH��1�'��ݢ>1�h�5�}Q��	e�3ؼ��$�l@3�ܽt���(0���w|�a�|D̀ق�̐,!E��/R��\�//-��s�3|�2�&4�Df�g#�+J<]�X�?�6M���.�"-P�Ђ>�:��jm����j�Y����$:�6@�]�p�Y�ϑ��)�Y@��KH�"����l��FQ4��/�q�I��,���`La���}�"����u��K �?��@?T�_�T��8*iq�+D���֔u�T��C2�'���]^|� �K�wy��&΄���x �������IW)���x0���~�}���u��%�F��KE\�E	 ��qO�~��/3#A�1"ؠ���45�O��Z��q�,Q�+x� lW���]�b�0[}���wcLI�JH6d�r��+v ������Zl
�����I���Ԙ:��#sG���a�w���,@����-Le�
�QJ���j�u�0���x����;VX
{f�Շ0�@��F��u4������{�Q_���8�t���v��0�ӥ�e�����b�rgA�O	��;A�-:�\;���@v�`��s�F��ڱ�%}x��nW<�Ԋ}<��S����z�l�6�ێ3c��Z#Y\�I�g����#!x=u��b�64$�6y��OH.O��Jq� ~(`$���*h�w]�U��m��@��"w���;�XG�a6�>��.¯�H�I+x�ﺋ}�y�YO�f,��nX)iֱ9?^�A���C��Ə
_o�G���M�WÙK��o�\beǘ�#�	����F����2Fy#�Ϯn�l����~>�<#�C��؈,m0��14�R�w_��+�W�hWr�.VU�'���A����#��?�����[�HSR)��*
��31�p1dx]\�DY���~�<��x��3 *M���z�1%��0��48@���ZY�a(�G4'��apRt\S���X�	�� pް���}g�ܜ���I���=�,�%�
#���pR
��[$]Wem�Z�Bi�q �'�}]��&0|.���r�
�4���u��n���Ӕ����AwRC?f�y��v@?�L>�6#���i�`Έ�$Q�x�Mv��U,MK31�B��i�U�S���{� �:��&�:X�HB����~��f.*<���b���.��q�D��,�p�&N�K;�7B��Q6�J����-�Υ7o�d���	?*��. �Zh�z�x����GsεJn���H$��K@Ϯ��X����~O�o�P�n�=T♯��]{ÐρCΰ���Kf,�q�@|��K#���X�uG��'��M�|�Q.R��:Ds�=%?�N }?�Ə�c9IUk;�9_�shi�
�j�,�;�B5���l�*���l�-"��jW}Lg�t�4�v�I73Lfz�`�x�A�B��ұ`�^,�B���
e��0���o��e��	'�Y������ܺa������3vn��J�$� Ƈ�z����oZM����Q���
߅��:Q�W�7�*9N���G�SkxU���7!C/��g_,-V�B��%�8���g�"������������bkG�X,�fq+�9[VKn��<���Ǩ �$�rS�2nݼ�*'n
���(�bk��6���z�0Vc:x�O���t�$u��C�~
,yO�O�՜$���+(6d��|�6!"�*�"����50�@�z�j���X��`V�䡼�#9e0j r�@ N�0Q���=ӭ���~Y�>.�u�&{JoԮ	�8�C���W`���8&|�ڕs�]��R`�kV:��n�7)�^Z]�)M�����/���'M���3,L�{Sp��H���)C����"B��eEz`������S�a�/�ށ�����܅#_�*��ٷ���v����_��_& �Ѹ�-o���7|8�O3��zq��o%NT��R��@K�����{M����V����A���PނI�4�\b/�e\;|̊�{��L�4��.�t���щ�"$�.Kҍ{#�BY��Տv9�)l���s���s�80ӲC��1"�H��=�~;��χkT��?�#�X��o�&�4Q�sz���#��\��މiQ���
z;�\�Y�;�����Շ�cz.R$���|y�rDG�+!ߌ��+�'7Lf !BѬ���zu}Q�b0����e� �<�Bk\� ��<��]f�9:X�I>�iGۻ�3i�fړ o��e��������FJ�P�w)b.���ا�B�Dgl8v�G��f�8�Q�F$�.��y��>5x���nz!͞������d;6 JS�m�HX�t�+H��<��ײ�$�l0���K��苸!/xS�&�&�V��R���k��JL!Bs�8��y��Pp>���͖�Vm���?��x(w�~�yK�����Á�P�m�z�����1_~?U�Ha�!Q��O0w�^3���J|(��9�MW/�9��$���o1����x���W0�J�E��{Ji�`ző�*��5�U�x$:�-"0����47��C ���OGzEQ�v�bl�d� ��;9�!$>ZR��Z����Ó�Iε<�Gc�����i�L�ܟ��\�(z�^B�&�$P����i&vr��_�V�����z^At}q�L�)�F�*fh�����U���j����E�a
���!����"ӷ�"���B?L��7ye���@K�ּ���H6��@W�Q߲�F6X��Zy�	����r��>1xI	
�	�N�E�)��c�.?껁P5�a���
/bi���c%�6a���Դ���C� $�D�R]�C��j�����b���t+�n�6n͙�s�%�U����������UţIҩ���83�yH�?o�fw����	��J�TyB�w^�r+��6�i�+$�>%��ۣ�msMEx�a��ڡT�L�UT��kWCb� 8LoĎ�s�~��'d�UB�r�-��x-%`CĈ@Xi�L���s�=��������������3CB�3�!��6��$�o[F���4	��`(�|������3�	3d�O.	)s-�w���S���;F	�q�ҁ�\��\Ş7�[A�ȧ�t[����н!�/P�-)\���5�Z��|�ŉɑ�*>'tw�B�* �-�B� q)��jv.&�>�k���8��8Jf����>j�u
��u���_0�U�t20�l�┄�e���a���W���t�c����Ң���<���i��ʌ�]P"Tm�bFǴ�U�^N|epWh��rӱ6H���C�H��I��Xc�QmT�alj�Se�}��e��Ԟ�PD�TB�b�i2_H���__�Fc�y�'�;Q�a��od�eA���|��^>��"Gʸ��B*�t�^:�|H#������e�	����nrv�Й�S��j-��f����s�zNѣ���i�K�60���3~�k��$yȓ������S�i{�Y �%֓�m�:�J�[ |�C%���Εbl�Ŵx��c���^�\���t^η5�qN�W��8��}%�-]�8��]E�`�z�0���.�.���x�7De���<��L����� 7z����]�r�57������\Պ���-�gM5{Wnla��u
�254ٖ��ߠ��2D~1�����d���1�J[E_�u�ث�LhG�.���Q�r\�9��vW��4�����m�$A]'�X���㦔���Yw�N}μ�U�bH��G_���ԪT��-D9�!J�V=A!QD_����.��-�����U�~�(4��>��� ����$�88K��ԁ�@�>~�Ι��PS���k8O�a,̳$�������(
�
ˠ����5<�x�\OR?X|�*u� ��^�6�u��Dn[�|V\���c��t��C���ҩ��F��Vc�ۚ���\�=tl=ު24�NĹԅ;tد��7�xI�`H�"�Uͦ�o
Mp�D� ]X��G���x��rvw:lQ��"$���ϒ��G?p�}���)�K8rY��lq���#�g�/f]����XT��7���׆�9��6n������QE�m1�����c�!~�*�T�Pe������S��fM��Ÿ��64 ���bǄ�E�M�`d�=/�*�m3l68����&��p$}��)25X ����zO&��e�^|��,>���Cz�.TSl�ԭ"�y6;"��+���ɰ]��I����7�To���r�? �<�r�2f���a�R�C9V�$w�p��Ȭ��	�J�ghv�i�C����x.���z�L��gC�~�����	%�0�,;�������)�|��x	�|�zS�~O��3��پ�@�q�[���~It��dו� R
��_��f��TA]:B:�!�@%Ȩ��[{�Ǫ�_*���]t��ȩ腈<y��i<%��y9i���Q�دV�3��إj{vGHB��z��_�/�X��L����ؠdώ�Ũ�?��jU�1��V���;�� p:s�.k�$:��;w�#&-s�g�9ݚ"�V�F�B�j����c9�n���ߦ��S���[*��)K "��J.��0��ߞg��i�94H�>J�/�ٕʞ4��}tf�1�C���5W/E�1��6�PV��:y9��抅���n$s��ē��P;:�V���9�̚
�7X\���/]����^"�L���]��-��5����}�������K;>&��Doy�������ݖ�1�� (���0��34�4'�:��?'gp���	o��kUv;����2)A�,4@��ԖK殾�t)�G�I �]=�|51��ωukBoX��.,M �}���~:�B�PZZ��C�nd[ls�����߯�DF! �LRq�ֹq}��O�d`� &�>���@���&8vb�5>�s,
I7P�ax�;��@&����?��}���y�~#7�hƴ[G�TfӀuΩ�V^�`�t�D���:�hG��u�޽NFfl� L�������İ��>U�]�����]���P�*�ߒ���\����
��f+��Y��%������C�W&���K�G�0]�O��(S����(o�.\4���3a/�E@��PI�oo���@|��i�X}"SO$�ZR��kdU����١ڏA)�Qz�A`��8�"����5FҠ$7�.a5���c�O���pl�AXb����.�ӵ��Vv���rٟ�Kt�מ����]�1WU��
q�qK5�w	��4�O�J�m}�h���zپ��]�k��֤��[���V��c»���Y.&�V�wJ�Ƿ�}ѫ�b�A�7���!g�/����I�O�k����Xhs�7�k��\TVm��~"z[=�ƨ�B��M�G��[m􍵎�j1_��J����c�����x���e�ag³�:�lC���A�l���[bhw8ތ��Ù�������Rw�7�$\f��#g����ǜ���r]��5�g_��RFm�l�h�.ﷻ�����A������QF(a��%y�׼�V�M�^a��V}��pl�X
t���E�m��7�ޣO&�~o�M�$��u�3O�����[�0��!P'~C�4aFc�mA���kQ�0�}��9T��7j٧u�9T��4�Ϋ
����!]�6����K��y�J@��y{<��uJc��-B�Z"Y2�D��*&H;
�t�S�{����M���UkY,e��Ҏ�g�<dR�w�p��.ՙI���n��:�ボO����]]P�#EZ
:�Jl��ٙ�e�� j� ķ{�������Ypw����#��?}�W(�wOA�;ؕ���v��*�ˡ�Z����V�'�L��!r��ʜ��E���.�T���
S��Ȯ#ER�5[È�+��}��X��|��+WE/3���Z��9�S3M
��J-`!�}�IU�	X;p��
c(���!��	 #<�'r_Yoa���� ��ɷMd2��!M�:��<�M;�ƨΙ�ڦY�\�� ����jkXx�5a�ӥ�(e�>��=�~�c&�U#��Y�µv�9-UC*�/2g�
��n�
9lqR�+�4�]