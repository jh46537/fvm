��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���tǐ-a�Z��e�l+�H�uW�Љ��Lk�p�@}5�[o�Hݤ|����j�{38��/qlW04\h"��=7P��2.��[��,~�����d���4�o��3%��!�:���&��G�Q5FJ���H�(�m���G	.��I�I�_���]�r(1��k��0��h�&��b��j�����Ǘ�g6Ԥ�f��*��9dS�>}᝟�i�C�C�����Ó�����RǬ�]�BU�����po7(gP�ݴrsе�7�V���~'�u�=��Y��<�(�;?}��Q2_�����-N6�R;SK8�n#1�d��0R*h%]6@�Kp� #�|�S�nj�C���� ,`�T��m7��O볻�ʗ���lUw�{�\�����pL����@��pEkR։��h�����,�Bf}'}'zM����B��,t�T6��:��� /���9&�����.>������s������*?��:�4�\�Č���)py
\�cm�b�T���ː�DӤ�:�Qn��S�c��*Xl���F�fec%����,����2�p���'���-�Q�̣@�Zv6��/��1Ǵ�����!a�]^S����.��,�_�o��(ߑ�FqFʰ��l<����9Ӝ�����t���$����8����  ��o��R]I�^"����o�`�*�D
�Ҧ�Ћ�.'c�Lv5(���#�����01+���A�������H.��oU���JT|����Ҭö��A��tr��	����c�*�r��e����W���.�o6'Cn:��Rj1zCXx%
�iA��.��3����v���vA_9gd&�{��\2�5�Q���D��}�衃P��ι��{J���R+N�L@i���	$.ظ�e�Vzr���S�^��Ö�����l��
�$����`I��B*�;҉F҆HJK�����\� +��Oc8@�&$�q��8���ʓ�$ �E�.؞F�Q�Ϸ\��[�0�!���jz-1����:ʱ��P�~9԰����-�oo���
���������`��3gh�}�q������`(W�P�Ԅ�����ڄIb�s��1}�Vr��ǚ���f+�b3X�
�w0<�Ɏ[=h��S��\0ɛ��$鑩z	_��GLE6X@�Rd	E�cpݪ�N[�����B&U�a]@-�H��L���p��C\�
>�w�ӛ5��Ne�3Jw�Q~���V�t�ϼ�U�v%��F��is1|bLH�A�	ڌO����׹^�_f�h皫���S�e��x!q��o�����憦�}0�q�=䵴~j����Pʣ�?v�$J[_�0̗_�D�������%�;�?Rt_��S��Z>pA)z��@�������~X��s�(t2��oDq�m+X+7�lq��ܿ�����~�����tKJ�����9�U���Xԯ�,F����DB�1�D�M�2�{�v�cX*�%5���c�դN�����hZ�Yx�m��B&�qIB<�cG��H���77u�YI�,��{��}�Ѿ@���B�U9x�|�m���~�!K��ng���ME��en	�@���ٹyV�9lH��|�?���6ܩE���C�%��i��i��&�Da��;��~��1��sɏ��\�����ދ�]� R�qP���&~��*r�Jh��i�H��r��6�!���,�*�R��tz��b��$�U��ap?��>��<u"��!�M���6� !��Q��Ǭ��Q=�� �R��i����(���IUGxS�p�_�rw|�������k���*�P~�����$�(Y4�PaYM?)�C#���6��N��5<�����ZTL7+�^��f�wƚ��W;ӘQm��\���D���g������\��������m&Aa��,��U�[�2��r*	8m2v �}��V��W�>i�Pk��]�=����,�7@@��l�����"w�ۃ��+W�= �t����O���/E��fn�� ��@soY�H�4�%f�\��CmF�֞bJ�8)W�K�L�H�m��ׅ�&|;^Wk�a�X^My���>{D��Ty>:�.3��/��}���Nq��+����
�0>U����5��i,�r��z@\�Q%���w��� �(ls<cx��U�S�� ;�Q���J���`���#�Z�����y0s���wF�V����5H�4��qJF,�#~R��&J_��m���p����Q���=L	w^�L�ُs
�A�/C-���~�������'��̡f�.NQ�!���^x�*�|�<b���u���8r�k������{��H+g�K�A4��6���E���H����Y�w��ۘ�Eo~��$�"���G¦)�swٓ�U�A� ��/Sd�4�+@f���B-�G������5�,}��*E������c����F��JC���o��2�C)m��@�E U��v'��vR�ZX�$��6@9��?Klbo��N�U�u~¤-}z��z��1�C-��U�eTs���ӊ���".P��չ���W|�g�Zwp�~1X�q�gY��f�9R�C�}��������\s��5j����-za3�H��9�og��'�I�-5�3�j�FVɭ��2���㹍���6:[�O�pD�O�`p�_�IK?Ƒ;���]hś�b�jm.�"Ε]!Bݏ&�@�lQ��q�q�۞k\]l~u	�l8�`3�=~��*��!G�Pڍa����k���
�p���3��"pT��+�ƭ��f��a�ڄ=YZ��>�tHg`$��ƻ
�j�B��: �Q��zZ=_�[[�k��=ŝ��'�_nR������T���*�a�e��8A�?_M�($/��Ct0)\Ԟ+���~Z[���\�����E�tn����fL��1	S�<WtQ&�{5��N^x��~~���%C9�h����:�4o�E��h��*jfwTO� �Ԡ�_�WBZ<�u�fᆌ>p�o�Q��[9,��b)�����3'}�&���S>�s'�3~'up�B���;x�h.��ěæ7f�k2���3f-��,��x���sP�=g�m{���~Ȥ�]��]
u>RzC@�3�۝�;8��" ��@�D~m���#J�_��qh�����,�"��_˰��j͉�lՊV�Gf�de�;ad!��]ł���(sE�5�鎾��iA�1�UaXb��g�P_����2��h)��.��ٹ[��<`��'l8����ZY�ۓ���f;����+�����E/ͥ���kf���`�K᯽m�<�6e�z��~C�3��T���*R����3DTUYyl��y+�O������< ��9��D$Frׄ�.�*�+�A*�s����p-��$�u�L�1�솀��Q�����Z��7��ai��WLbL��S�$��዗�w���Yl�'lyJί0������'#j�q���	�I�{�8&/+���ݩ���5�!5���:��m홪�B۵��X3{����$Y�@���.���G�4qg��\�:�k*��D꜎�+�Ɵ
AD���q�0��G��ʆd��-�����RV��|�|��I�f��0��	��Wc�L�UyJ�E���ZWす���� 8�`Y����>	�� 8�9CX,�A��â#'���p�%n�3���)v񠗒Y٪�Q�&<�Ε|�80����A�6r�=g���Tkٴ�RM�Zz����Ӱ1�x�9�=J��8b<{ǿ�-ޒq�b˺j��Rqrﴟ<�� F�I��	�W�D�8E\Î��"7@h-�{�*��7Pr]�ʳX:�J[��������sM'�Rܩ����N�Klҏ��&/��}��7��p�{�+҄��~��u�%�`�|�:�5)�Z(j���X�$,)�auC����W��^��fq�!���A*�����U��XUWg�5e[��ٝ�;�:V� d�˶fs��*�g^���i^�F���cJ�Z� ����\���~�3B��ޤ����k��9RiH�� ��}���,/���CT����٭��,|cs�K�&iȦd���PR�9��+�v�t�O�qC��N\·��j܁B?��=5�6%���0E��1�[�@�z������q����#ޤ�9�x](�+��j�-����v6#L$���)���g�6�=��`K�"�'ި���^�|j�d :�?�	#�҅#
��)���l-b�%�2b�g|\�'QI纱⃖���=V���Vb�cx����PFF�k��Z�k����"DG/�XҾN��"��x���s�o�NXo��@k�O�z�Z�j�lۄe�N=�B���ׇ���[��)LŞ��s4<v��:�W�z�	@�����2�:.���7ڿ K`���7�6LQ\Ժ4}Z[�3% f���KKb������:W�/��_���b�����窪�z��d�f���}o�WR�Z΋�Ob�>ř~=������d�u=?g5<�v�d��O�&�����ɽJܻ�_X�3�a:�_��e�[�^���u� ����RC���hd2��>A�2���M��!66
k7�SG	-�aִ�!���i`�>���m�]�p�NuL��-R|ɠ�6����,u�i��\~9�fP)i�3fQ���*ir?��[�m2����>~�Q&�5o���r+ʬ��l�+��ޥ�i�x�t`��5���`@=��\�Շ&J�F��>��A��&9��oT�1+����i����t8ux�K��
=�����������rt"�ޢ��^��1Lb�{.q��4���z`�D2=^ksP�e���T�6f`H��y�����{@&.��n)�/x�����bv��r�2*h�(1�%�G�ȥ٢�0$A����t\r��3���pR@"%=dQ��>�lzl�3�^3fI��bv��gT��4�B��ۛ���Q����_�J��Hm*���bW/9�6+��T-sŠ��{��/(�h�i˯pD�t�:���Ӣ9zli,���$:.�����.[�:}3f�*S�Ȃԝ��+#� ��?�|r�l�"��=Q�T��
�QV��0�e>����ס?D�7X�7�d�a*�L{��V���<��+���˪2�U��
q!`@"�+�vHi�lE��@�����_����z�Z��יi/�?��i���l
u�����T/���B�]����.d�~�� wN!aU�a�;~��;����t'FC�Q/��$x6m���q>�*�X��x�&�V�f��������B'?0�
�J~��y��=i�5�陻"z�&� �T�$[̪���T�|���<K�@�n���,��M�?�װI����a��گ�f{D�i'Ӌ'���P���ͥ��J�g�-���C6��:����o�:��@�w�x{E��[���k�� :		���A������99��S�م����C�',#�h4����E.�]�L�/�_j����5`�F�}RpK��8]�[��3\��jBfT�D���Qz�x�w��_IM�8fT@I�F�`�v*���,�%��^��o vyG�Y��W���Mz��@M�}�Jh��9���BV�끙�-�ϨZD�5v@�%PAdPc��7m[�
�U�}w�T<��t� �/��b�(e\�n����r��v�����D�KT�$�����WW�sO��Q#����ʍz����|����G��a#����p"��,��3Q�����3���HY���g�b�D�#W��
����j�> 1}}t6إ�«�eU��y�ۗ�F�֙i��=��h��W��ɾ0�����6-Mܖ�:tr./���l����!G�U��L�Ф� �{�	�u? ^_G�d�7ێUD�*`�r���:����`��bfn�Jq�V��ao����r��'���H���g�a�q�}�]��υ#�������X8�z���u������7X��y�J�fq*�]��X�7�dZ�)���x�3�_�>6G��ӄ��6���"�A԰������|��,��&|&�O��� �P�������uE��	)�E���� ��O�;�;��ɉP|z��q�_0�Q>��?���N񵸾��	傇���\w��M��h�ʹ�;�F���;BŠd}�=V!0��J��������:�l�#=  �%\M�W���˘�k����p���l��,��/�ݹ ���/�#}+�]%��`x:��{5�4�|��2">�.0�s��<��t���.f���C�>r_�x����{1^;$1�/d�� (�9�J<<7ie5t��踽>AvFGZ�I�;p~�6�i9�B���C�P�$�����%J�B�0]�40";�0��yF'��7�&5B�U��[u��v�1R��Ji)�ړ�-���{�4)��6^tǕn���PI�?UG��� bOĆ���g�����������.�),wlw�~`�Gj����xyI��3#�Ŀ���q���%~�.����i�P�$��TXrn8��q�mT%R!݌��o-�এ|��28��t�{��N]C'D�n�#eg����p6�5
c�h��"]Ƞ*j��w��:V��������yZ����N���B���	��h~����}D$���ɤyq��fZ���Z�~�3$O�,򞠛�1�#��R�
�0���R��$�F>Ni��<~��s@]�&�L�9�����\�S�z0&�C�����c��	��Q��*Gm!�%�i���(�\��5��)�;BI�"j�-��'F�)]󥞱�˙��Mk������/No$�b��߮ϫ}���1:�������0�.i�E=uap�+��}�)�҈�:4�$��ʿ&O�>�j��^䈝,�����{��X6F`�����-��]o�{c�-����F�� @P���rM�<U��`��o,{��-X֥�[ܠ�9�B��2�:�m���ű.j����$S5����b�������|Z~�\������ņ[H �?_X�դ�G�|�	�]��`�
�
oL�l�F'�P��_XV�&F��.�f���},�Tw<����F<�	*�QYN,�	*�*�ovdw*Wt���]4+��U�$� �sc�����V�k�^�py�[�,{�z�@�O�L��/;�f
;V,��gfW�᷇h�Bd�d�?CӶ��FV�[��"FnR��|@ٗ�����A�9�*������PW�xv��7�ˣ[���c9�VȩG�ӓ�`�M���8���x@�4��Q��_�
ʣ���6��DׂL�7qR���՗�AhɃ_���{�����
�ʉ�c�S�~����v��d��$��۵�(�)�m�|�,n�S��{�Մ~�^�m��7���(S@lj�#g��
A�����j"�ò�/���q�73�_[�������B9g�Ā�D�����;���;��=�t�̃�|V�e瑎B(5Fy8b�� ��H���$ȶ_�����4��>aT�J�[Wl��
�u���;G)�/^��넟c��D���w
"�=9=�'�+�pH�t(yKMxIށX�\	�dF��G�� ��l�������	�еZ(vxZo���@s0�?��,л/��x+�V��&���r����ʞ4M��@F(>`jN\!N'�hk����A����f����u�hնv�~Ь�뷲�P�f .;_b 3����R�|Q���ڲ�Y�K�I$(�_��j��+7���,n߻�5������D��S�,���fy9�uX�o=�+�'���H���d������P����ۡa��ۗq��S��;O�& u���8�"ߩN�C��v�a,ԥs�%�+ǿ��Q^!;\��YYbB�:p���5�hb�T��(���_蘦|���6�2�9S �P*h�Wֽ���<A�>�_�Þ]�k3ڏT�� �
�v��QF�H�I�g���F�=�{���\���&M-'����\�z'n��Ѐ��_��N���b�^�g�Dm)�57'p`�!�q��>S��3p�]x���S����;��C�>��&�A�~ ,y���*9C�.ǥ�cej~�H� /Z�j�z$����3V-�ď�w�o �'�A\����d�G�Y�yC�C,�VA��}F��hlL_��2i�����|���\�9nŃ*B��*����?��i��K���%���y#��@��1��ڴ�⒍V!��V����FΤ���}>R�k�0|H���T�݅�j��p��^7:���7���x�H����9½Rov�G(*�&L��>1��qCS���䘌Ur®�W�]�(}T��P�?#�RhSV���eU�I�N����k�"�戎S�6�{��6�Њ>�ي��<`��`!tԺ�,���s��VY�1�]�9�2�F���m�&a~�L��Y	1�\��U~��}As3@9뚍��«='��%>b��v��;XF6��ߧ)��`P�/�!>�Q�?���rQk�g�!��hH2O����q1h.?	;=��
Vp�y��	8m�;	C��3�c\)�cmd2�$�v�}Q�s�ۤ�J�)�ΑP/[s�<(�N�Cs' �a��_bk���dθ�Wl&I^�[�"=0Ø�q�9������b����	�4�]𝰾L�fg���g�A��J�Z�k�� �o�<��`X��]�/ ���:���ۨ4�����6��Q6�n�t�Q�^�}������C�x%�I�-d� [��,z=U�)����\��ĵ@=# /�}��(X�iA���p3��>�ˁ�r��}�7�į�Ȇ|V�1Vӥ-�=ĳ/Նv��hdwܚ�T��E2��M�D�s^#���Wt���
��7���ә6s謴���zhq�7�fڂ�
0��1� R@eV���̠����?T!�㹤[�<�}w)��H�:f�)ع��gH׽��e�t�`i��v9oeE��I�,T�,�g�kv�<��@�1�;�DiCKGa���G��xR��y^q��\�Sge��m����q��(�ϝ��l�!g@��?n#��*��1���r��x��d7�R7m9��c���u��M�������m�R^Ӌl�z��rf�3�����@�L�+B;Հt-��>"��0�K+��=���`.��Gގ����W�Ҩ̏,}�];A"Z$�u�:����(ڀ�ZW0ᛠp2uA�;�ѱ����]�-�����5X��"��p�(�zZ���-���x|%1��,t،��ʫ�~�N�I�Wnb�!�E����*m|ii���i�"l�i[�L�vCX�ၦ��.)�P��":�_�-M��Z>�����!��#�r{���_U��5�r9/��Z.�H�D���zG����fgQ�{�r	��?�ػ�1;�_�,[�bO��O�l����Z&�f_-�{*O��z�+A��V�����d�r�j	�, �Ej(4��=$�J��$ڍ�p�u�T��d��~��g��S��\ Z�m�?�K�*9$u��;^��[2�1��<aE
�ï]�S/��g�%����w�i1~�g5r$i�5RF�