��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,VI�0=�E��Ӫ�-N���=��_�@Q�:�7�����n�KyJPq��QIVC|w#�18������c
�X�e�n��8��Vgdz`*}��LW���$�s6�j�E�r�bǙ�����.A:�U<����Y���:�*��^#t�2�U��0��d�	�Y���W`�A�<���������(>s\�#W��Z���XgG�����p?[5H#PuD��SW��������C�|��:B��`$���`[Æ#�^�͖�b�l�3���V��C�VK���t��_���K�֐�!�?Ux%&�$���F��y�-I@�k���R9a�eo�Y�T�Axx(�>Zr��&�e��P�C��-%��]�bW9�k�*/l��N#���<�,��مaQ��-�_K��"z@�#����'wiJ<�0[�f�"�����s��|�Z�p�3׉�A}�A��pi�.�/D��H'	��&��L󲙜tes@ѹg&5�
��Jf'���׺,T6�2)�\
�����U���N��Al#�"����Y�D�tRZw[d�C)PQ�\�_u�{xI�7��\Jt!$����1������C�[qLVW�"�9��=�+$�Ҧ������<�����T�̈�WEh�z)�
�=.��ѡ�B�l�]~	RC�:�:��a�O��3_�%V5���Q�4����Ǧ��ȍ�3{�٘ �q} �Z�7!�XN�J¨�gR���������ڥ��P"��t�L����I�E��N�3#A���{k�vCxE��Kv�F��2��b:�Y�m%v�sĖL�nQԿ�Vwx��!u�隰����6T%%��!��C	�F�7�ᣰݣ~��a@�c�D@�to��i�P�y�I���&��$�z*�'�F>��R�x*�"���Kzc��G��-P;:�M^z���o�Bp�("D>5�78�;�9�[Ю#�˖x�Co�ɛ������t9�&�=)����] �&ΝQ�cy�^�@|�ں�W�d�oPrt��T]i[e0���H{�o,|ڹ�e�3�2�>$���|��Ra������!%���1����[��[�0���d�~	 �����JF��H�*]�WI^���G8,�i�5�y!�KMlR���e�K�Eb{���x�c�ߪ��
	�[���'#I}�F O�T���w�W0�h��]V��Pd��WdJF!�l�cR�.(�5��/�����e�G �H�F��xs/︩;�y4Zm���*���M6�n�c1����_�I�HJ	������2 �yA�q5	�/R ���cK�f�>H#Tm-V�U��{*1��_>q0� 0�GR��V�eD�Jn�=��rҏ����}���g�3+(}�QN���!Ϻ��a��<�'��1�
P9�i�+G��<=�r�G�1nSji_��*Z�I����: �D�sp��yX�)�c�)'|(b�Yh�MI�iQ�?-���9��tBn -�c�e�]:�D���݇ЍQ����|�A��/�f�9