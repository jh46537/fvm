��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��b*]���I��̞m����
��6��Tt��{���#�=��'o�c��Y*b����2�������4Tx'wiI2�^���8�ف_���岗b��,@MhNW���1�q���m�em�D5�5 ��KI��l��}��:�Y+=i���},�Os���)�������냁��fg�]�i�A��8����kO��q�ϔ��tP�tN���,�_XH�'RU���B!q���"��imn��~��5��b�n���ι����w�EWr�>�OG�;�e8#%
���LO�6���P�j�����A��#�4%�W9�����.^"X�"��r�f��?����h7~��ou��vԈH*��ڀ^�v�:��5�d��<iCGVa>P��OH1!��T�E"� k,O*O���� �ɭΫYl_�E���H7��x��y�N3�0IQ����Eur�"�Ӛj�{�tg�V���0�xj���z���[BJ�w�Zn�ڡoB���a~�T;M3��9�.9�U��������K���%��W(Jf��u�O�؄틷"]���#�����^��kA���l �bpq
���/�A��G��]_#��QD�)3H�$T|m�@�S ��9:~���M�S���� ][N��Bn�����ͬ'd,ȘjdY�,�@��x�A���ܙ~��싫����\,���\�A%�I��Z�ED�4�b�T�6���:�/�K`"�:�ǧ��4
����]���,�D�����F]�X�]���B3����F�~�k�BY�����^��m���f?��Ҫ旼*��ٔ��P�Ʈ�ɑ��Y�� �@؁�l�b��3O�-�s=D���_��#�I�A� w~A{��~�>��.˘+��J�Lidn.�Mk�t��^<��8���pXYel{��a�#_�}4�*͟�2��4t���7؄��I1�� z.�&8����1g�E�W�c����������}�B�[Z��'&*'����~���o'�1���g�]s��#B���sޢ��9F%Z���:�:�����.��
8E0��g~>�ʉ[�����Y?�W�S�ݝ�E5z���kv�r[>_��o}V�y�E	S�����/��S�8��r�Ь40S�y���%�s�R�Q���,E���=g[Nls�%�N�)�h�pX5����5�pi���@|R�1M���}�P��k �PY3��ٍ�ܐ�kp�Z8n:a�Na��bS�e�����ͰұQͭ/���O�Î�r͟$�PT���YT�����6�*���'G�$^���_h� ��N�vh��;�e����@�����e�K���U��	�<��,"G�A	+.�'��E=��HÙl1!'�t��=�e��/���Cn��� �K��c�t0��d���x3�":�`3+!�@Ibǈ�f2m�%N2Z�1��:A�2��]۹�	��Tט�;�G5���Um�����-��KRށI8�iM�{�w�iAw�,��ڤ,�0�L;�7�U��1��٦e@��_��e��N,0��-��>y`RO&%�zᏍ�T�,C��Dvf����G^�d�<�ׯ=rW���t̍�v��g舐���=��+���1�SC\��)��{!v���x�x�����\%����-4�'�`P웵�i��X��#.�7�f�j���Ȅ,�C�򸷝��������|<X̘D�$#������Ѻ6UPK�V�f��T��H
��o9��ȧ���KWl39����A��4�e�n"�[|���ק{a�������6����!/�:@��~L���+@⽋�1�����*�mk�aĤE7�_G��!����L�]�mbC��fjb��n?z��k�V�?���6�%��H쥐>��6�V$ �4D�G����6�_�4H��c�|j��lvh�A���}PW�Wr54<�ɷU�C��Ryk�_AN��gO��3K����D��e����<Q����a�*�%��ޏ)�Ql_3��gD�͉�l��3#�ALHLD�eQ`k��V_�[KWO���[�<��rǞJoh�jG��Ը���=��R_�p�#۹n1	Ai��ڤ��X��[@0���H�kU���L!���?��Z����y�~1BEg<k�"Q�JW���3Ώ����Yk�c���M�2�a:`������6Y�>�=Xi�R�ؽ��⾧��R�R�a=-����l�[.�ob%k�����Rew�і~�i8�M�}��ֱ��D:�C�{��1|g�z��Bg�H�����ig��w���;���-GK����+I1�� ;:��.�Z�k�]&q#��dI�$��}R�j�^ðiW�2Eޢ��>�(�����F�$g��?'pEDT��2t� ���a%�-z�������T�p���Ryd��l��ëA9���S���.3�U�^,_+��r�Ov�C2ʀ���7�-HC]j������X��	��\�A��r�q�CQ���A~�(���̛r�-�9�������WL��~��B�#�hx7
��(�'<�cJ��zE��ό<����Gh&�P#6h��
o~(�9��&ؙ��$ț,'���t��!tB�P��G����v��Ur��Z����o�3�~���	���6]�(y^p:�ç�m�S��4�|2h��¨ �HS_������m�NO�V0N"}��V;�+��K��1E�-1A����X�Fy3f��	�W��`�W�qJ�׆h�������[�+�~��ꏤ� P�ok�@�[�w �������3�$����D�䘄�F�5O��
\1�plj]D�2w�N����SL��\hMFވ�E����@a���+���[H�($�ڟ�U�������"A�����e�UP;��z]�(!o����qmP��a��p���M!y9k�4lH�J�,1"O��l�VUG]�Po��D���jx3z+IU������˲�=I�B��B{���Ɨ���V��s]�M�˅�Αf��ş@Aw�p#�dB�cPjjøaF<��Dd�;�|oY�(@᫨�
�{e�Z@�	���E0��Z�ů.r�}g7��\��"���U�N� }��.�YC�Vk���E���$�o�p����[��=rdҬ��El��fg���Ib6g�ūY��%�����"o(�
���P#1O)0[��I${>��J�C+�
c���A���	��2[c����&b�'z*����Y>$٨���M�F��#�2P��>q X�MYrǃ���1p���{�!~a0�F�#�i�6�#;��� �A�B��{*���~��)��̻��+�	�?3t���	p�����S������3�}��R�X�Jq����/�_Ӱo���R#x�j���-L�A��c ����BΦ7���k�f�yqNYb>9�"����z�)�)���,L��	��0k� �Gڹ�?o�i�'�e�C�`�{QB7i�:w�����5c��*���3v�]�8Y͍�(��i�@�*n�z[%JVk��{�ݭr�c �ܤW�<�n�i�Lg�^\2$�#�(/�#����n)���I ����l�-�vs�'�ip��R�13�#��b���H��9O#E��_��|�V����ɻ��U���l_�:d���x��E���k�Xg���"�ԗWIY�(����Y#I��D#����pj��������K�Z����=(����q����y+��=(�.ћTp��b"�g�u���~|�� a�t^,��m��M����r�}���%#��;�Y��W Z�l�`�q��6���>�Ss��J��]��B:g�<�y�G�^7�F5��� ��
H���{�[I@=4��1�	)���@#fS���hi3��b�ڦ
s�aG`OIЎa��C��}:)����4ƶ�pG9��W͒<-Hf��_�3�,�I���2ϑ�����nz(F��S0�mT����!�5���������H4)�a4D2�l1Tu�L�`zFS�C��u��`!"�6� 04���g,��2��i��W�D؄`h�OmS�dP�|���ry	��g��XC�M�ibi�۶�eJ����R�����^=6���ƃ��]L���)����q�;�59������9�{�P�d]��cbR�vD��=�S�Q)��gK�sƈ�A�4T�+�N�X���]Ԅ�녭y�f�g�Y���~�1_��soZ�GF�o��f���ܯb�#�$ ��t�������n�St���:��I�G�&m~�O�^��;p75M)m����`.��h�"������Z�s�>/�H���r���;A�
_HLJ7 ��g��.�8�D.���
�73�.�=xd-W�t�ɑ6��VsnoѠ��R�Ȩ�ZF���r�(��>�������E]>�d�%;����#�9G��n�pd/������J�r�8����(��w�R��!�e`���}OB������A�g[��֢N���EH?ѠkX$��TU�zP�;.��p������=�J2�l!�WK&�#����n}���|!�ܡ����>�����h���~
uC�D{��&?�[߲�w�a����-S@���vec(��?l\)&9:��Ț��|Z��Ҥ@#(*�v��p� �Hz����dD�b��INV�k;C\�Ɓ����������ᵧ���P��%Wzho�|�>}}˃M���8�|����Ή�3L�-���d�I���I�4i˙��	��~b+A��D��|��p���]>Z]�y��Vp���&��b�4���T_�1 U�d��5C!��� �k+��K2?U��nZ�
�j�����SX!������K|�>D��(�㘮�!?�������c��=m�l`S���le���9�i�J4��D&I��'o���Ś zĆ�5���_4�=8�/���ʼu��m��<���+ߣ&NN�BO`��M]��Hp~|k����4t� _/c�cB���&X��Rߜ&y��+��
��,�_�t���k������F��Ԛ`�; ��