��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���q����f'����U�S-Կ���Q@	�Z��*��E*��
C�~�� ��!H�^���q�[����A����(���a�)��؊IIb^�웻n�$~�����ɓ8h����FL+[�*���|BC��.�&a�xC,�ɳ��R�u��*eb���K��,��[�"���a(襓���x���pn���_���j�c~}*�\�����ٸ��.ۚԢ��U&���c�{�<�q�n �
���x�B��XAM !W�&��Vt>��W��)��M5Į���a��U�6��,ˮ��/(L�C{#�IOvE��[!�ƾ}�pK��N��Ƥ��T�h`h���ߓ�Fc��!B�K�[(�PA�t��յ+曂f�>�3�_��-tWD?y~u�K��&|����������3/+h��m�:e�r����K�M	h�݀�9�O�ڴI�*�m���GI�����TP�� ]
 g��I�>_�F�	��ڙ��J<w$Lޕ�)%[Tb�	�l��|Ā�kt�o�!���z�е����F'�+���=�<;	���D��kL�Ktrwm��zM�˭�8K;!9;��Ò�m���M�%�V����95F��Q�r�`S��L}�3�\k�������H�@�t��Kr��@ib�\��~4��U�^��S����5�Ttz��:�,�ʗY�HŊ���no�v�k��UԈ�|��@u��5�,�uV/m��0��?�t�� ��G%��2_o����۵��iA�dm��dI�{�B�g������t���t��_�¨PwfA{݃C -�QWg�@S:�F\��,����z��G�����Jo�'�P�TA:�X�W��MA�OR�����߱�X�klg(���d��k��+�:�2@��Kb��\�J�������w#�&�/����i
 V�CyxS�'���R�_N��B:-ē� +k,#[s�ꥻ���f���-E�����ߋU��8%���x�x@Ň��2X�#<�"�� ɇ<a�) =Oc���,��Uh�� �/�f]����,RP-���rAo�J �)�Bo����V{�tV
��f&�y�'�''xI�&�)����l��Jg0k���3m��ID�5�P�`/�z�aF�T)_�~�|�cZݖ��!���xN�[Vv����u��(�6!Hx}�'�kM_ &ʩ�P���)v� �W/)|�2ͫCp�����O�W���!�4š.3�A|�j`9��|o�	�SU��*��}�d��Ց��/�f�eRVALl3��st�d�+L���)&��������B��:��e"o��1�����J*>���;9��R�p|n�����_�@��k'��I ~;c�����~��mq��s� =氾� BY�k���=]e�D�N����!Y�n4�(0{t��ݖ�(���I��4a풨��E�2�]�=|���˦Y���l$�IhO����nݺ\9�����^(�)�e��@쐹�G��~i���۞N���&�n�!��knR�"9�PX�|���*LI�</l���?)Z��듦�J�(m�_��vӳ��s�]��i:hڪW�H�m�H���ۖ.tZ��6���KO��UH�͡FS��/;�Y!M��I�1V-�Z[ͤt(*k��n�.��������4̛W9���Sc<e���^x�:8�:����*ГN2#��aF��S-V'�6{���j���\��j�(s�ۅ"r:�������F�jex��rÏ�����4�<���C�e��E���o�g&5��׎�H�L2���Ƃ)S$�)����X?��r�Ե�Qƺv�5�q`�k
Ӧ/����t�#2�U�JE�P�?2܌��m��Ƌn1\%�?�b�>{�sx��3���g�8����'A9竬�%����.{�G������8%m��%h$3k�2�SL?>��/�v�P��6z�K�n]��1�"7%�l�:�zZ��s�������Ab�A-ٓ�"\$>�0+���[����:�!$��#W�j'���6�zp*C���x+��/pZ!6ZS�I&�b�\B������5]��7��#��a�'����;zX�U��H6�OO�%��K4�޿b�P����[���;��|�cul�Vj