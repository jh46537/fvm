��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�������s�h�qQ Ҵ�pp%�bs�!F1���|W��ٍi�\��չˇ���7Ge�+��9�*m@Mm��A��/f��XT��݌��GP�s��Ɔ4)c��f6�}jwS�����r��j����Īf�t�8J�gmdD����I��h9EWC0^����T�
�we�g 7H�����2�^/����t��PY��Ivs�b�q@>y�%K�~���*0p�w������
��w��{R�8u-C���_f(ZG��|���/zg��P�sIY+�e���<8%���⌚��8gn*rp,����_{���W���J��fM����D�~ۂx�Q|�hCުŶ�_����[�����������=�՞����6�����o��B�#A�����4��5s�32.�^�`�!c菂Q�h�;�wטvm���Jy�#�d�d��_ǫ&؁�	_��To@�7o7Rt��;�]�xg�8'�z�*�m$to�1��z�����ž=f�d8F�J���PJ���5d�Ӎ8�޿E�m]2�+,���X�)E�`��sa@A+3_����ǿ��n�A�^; �yO���'��فs�ݚ�W�/Η�?��C�:{���v+`��+""�>|G>y���X�bd�F�{�����P,����u�9�Ǽ���ot�|^��g��A���ب�YW�vƻ����_ۖ�1d+�fxR�]���)1hɹ�A�z���F��Wj��p��O3;d���Aiy�ܷ���)K���$�En�[ҁ(+�����[͸4���!��S�v�goZ`*�r}�[��L��#�3��\LrT��a�[��(�:-��=�0G��:CɾK\�a����sG�	p��
���企Q��`C�F�L�|�T^b^]��Z!.��/�.�Y7���7��v�L��>#,ާ�6uq���O���"�	v����`�L�2���9CS�1����m�M���N̺�\�ُ��DGTv�q����������6Pg����.�O����up?�A�xְ ���v�&(&ޅA�a{Q�;
�� �Xk���/Z8{����&	P���p	������񛶭�y����kw����o����� �YH΄�����O���
`)���9i}�y�#[+w���#E)e)R.ؗ8�
�/�����n���խx�X��d7��VU���b�7�?���}����<���~���*��y#�!�^�"E0��f�R�A& ~���.Ku���+n�������nXl[�X�.1��Y3���DW/����@~�g��I��t=�3](6˩�+�Q~$k��I��a�ݎ��5e��E*�&2�5諦�,��H��X���X�ۅQ�`)���{���5��2`Ե�J��O�-8ArL@�Cڛ\5�\�
C��_p�E�1� ��]L]�\;��k�Vy���N9m�|��OH��Ƃ�.�wRq9�`�F��"*R�i���O�nB�O|��OD�(���R[0f�HOyq�7<9A�`�}�rR��[^��щ�:E!��"tJ���(�ƒa�¬%�D������8�6+j ,D����ٳ��9;����N1Gu9J�9B���h���S�h�b%},�� ��(�q�Q�%\�%f�����3N]�.�$`6��kG3��4���E�.���-�MM#�¾s�x_5�5��_��
�&D��G���o<3{jB�(1��X�u��}��fIn�7aֲT'��l+�ߜ
B��
���4��o��Z0�W�q�r��3��x��� �x�i���$xz�[y��=��B?�Qv���� �;k���1	�~4R:P�/p�y��P��|P_1��q#�p7�Kh�EOM�k�N���c�_P��Y��� z7z�'ߺ�}���a�H�� �+�u1Y��Go:�	.vBQ�BR_�3{xL]©�Z�IN7H��ʟ���@��,), �*1��F_YV�wҴI�@�D�M���zpD��4x2��ab�,Zo�@��Z̊t�|��T=������>H얙��v�^S���:�UoK5�y3 ��W���J I�1#;h�&���9	�h�[l"E�����ӭ5��V`��]T=3kx��u�������|G��Vϡ���WT��N�K�p�T�Trn����u=�qhu��uJs�h҅�nk߯�3]!��#y�F�#�>��`ꅠ�TcN��M8��*�J(Y�D��
�ĆzY��1[���[��"�d"������a�L�[ڂ���XB���6�]�qy&�6QT(�tB�H)��W]�����!�����\��iLT�8o�߸@��!d��>���-�|+�BbRܮ����s���V�/�hM��E{��1�_�n�:�Q@�k�
ɀ{��;�ʁ��Yz���&��T��8��N�X��#|R��ǨY�X��-q�͠�U�.{l(Q�빏�C �\B�r�����$�ϼ�eZ�:�����֘v픙�����_��O�U�8x�|���]��M��*U,����] +���&����K�-�2jQ�'��0�0F�|
d���
]��� ��2}��ds1��I�̲JZ�D) �ǚ+�����*��L�p^�z�K�!����Жa�¼W�*	G����پ4�-��Nő2;��(Z
N���B�K7��qӌ�ix;$f�/���J�DpU��9������Y��%��@�l�EN��L��8G9�I��k�:ᶬ�F�4��~Y���*����^u}�~���)ؕN� �����@��i�����p62\�d�F�ش��6�ٵ[���U7��V3K� �AR�m�a;A�z�C�y�K�fc��;_M�D�$2��8�%�W4�M% ��Ξ���Vno�d�7���q�z;���P�����j�Q�~2��Y�	�г�s+�y
0͸2y}W���������v��1�����X큖~.y�����,�� J��&v�QG�I�Cd���S��-Y���0��ңD�$�	.*>B��My9�<������o;��!�
<$+��0{Q��g2.?�vb��$�� �A�$���i�r؂<2�x�_�`H�'7�O�_��/�@�|��B��&`~��a�g����gBߧ�8`���W���샩  �Mә�7��ʟ��'�1����,?މh�e�h����iR�m���F�eB];i`K!5Y<�͈�Ɨ��t��c�b�QT��k�HA���}IiT�7bsnHōk�"�b}tN�}��������^kf�������8�.�t�)�}r����%ZH�Y,�4�Q�Z�hȤ�=��,A_Ӗ�z���$k��5����tb���3�Ա�u�@�c�r�E��ޗ�o���?��l�_Lbf�.1T�#��lQVBc'l��z�R v�VAU(E��Τ�{Qs��~��G�	��(��=�Q|3Ҋ���F\�z>䜏LK[�gI^T�A� =���*��>�L�G/{�%]RB3���W�Tz^��.�D���X0/��j
�F=���[V����T���U�������_����!��Gc�j�w�>��k������K�=����`
c���Bg�����M7`���@�*H�s��c� �(��X>�e]P���P|��s�X��-�N 7���`�3�S��dȪ=rp(�����xﱻ����%��]��>�7L ��h��)2i pJl�4�C]x�{�^�P7��5|��[�*Φ爐 �t��.K��^M���l�8����٭̮R� ��!H��Ny%	����Pg�e�?l�n��Y���Ri��tn}�p���un��p������(MJ<�W���U�W�;ފ�)�t���^�5��me���6U�j	2�����u͓%���ë3U���&�"f�3�V�'G:�\�d�DK���Bs�T�Q���)H��K�E�R4�Vɗ�nH����c��n�0�e��5�-z���D�4�4(]��k��Y���7R�)%��k��=W�>�k�QAݱgJEq����B/v�B�zi��8�v�w_}�q,Q(dGM�����ja%�k�u'���q9�3��aV.�Kr�M)�*D�naҗ�I�z��!a�fږ0�������?�X��ZE��=��Vԓ	26h�,9f��e1�x >V�#�=�=�%���TD�,#�3-Z���,������u3�k��^P	'H�ܨ�1�w{	-��>��,o�&x3s�k��8^2| M�ʭ�5¨p�G�ݬ��3�1\Ӌ�>�{?����-�e��m�N�{cA@]{Z<Ȉ�!� SCH=�{� ��3���@�M	�fo�4���͐$nW�x�g��L�Q�{�t��{k�1�:z�Nl�(Ax�kp��wFD?����9���d���'���*P�ף�R�Nz�i�@:�|�V�������pZ&�j�*�7�?�>:0���=�#�є�>�:�3zw�����lP�<�@�Y}/@)�|�N}0��G�&����he�=�!��w|����г�@4��/%&�:#�x5w:*�栻�����q��Ca	e�٤�y�B(dԐ�7�<ȹ �DSj��u@=T��]���P�q\��b<of�-�/����WZ̔�u��p>W����9�\'u����m8\��;�_�1PT\��o"w��4�/�����Uu1&v�,���+A�i��EO�ԹE>s2�F�j��<�	_s��d�/�&\�w!MYp��0�71��Ws��`�X��M����z1-⒇6;��G{����i�~@(|O�@e��>��ك�'�6:��t����B��$S&^l������_�v[ЍcUhJ4���Tr֗ը��T#����[q�?�D�I��:q���ܽ��N��?��|F�8WS�2`���)��յ��w"�CO�+��&�V�#��&����I��ො��Ǵ�C	�V�8��4�%�I�T+f)��[}@�a5���'�^E��Y2�����\�m��p(��Z}���o�]��cȑ����fN�A�%�i���߇�U�T˪;��g:���>l���M�!w&2ך%�9n�Sz�U/ND���0��E�3r���~����W�X���'���p�y��l�����X��:u�d#@�N1�d�*�΢�?픏z�u<�q[���Mb�%X�{��u�צȇ�c�D��1�(��G�l��&��'?g�H�+Ǜ������<�P��߅�#*1��+b�z��BE�����<O����8T��!;#�]ɲ�����fI�Q�P�2��'��E�����S��"yD|J��F�6��L��C�O����Egwa����	���Z���*��z����g����~w��]��π]wI%�td�װ�+�=!9"l�dyɸ�������Y�"�3W�:�HV�3��/y�w��ـe7|3d`Q���/3�Ww�)�Î����9 i򃟾��{�-G0z��a,����f��o;���i`�ֆ�-����,V$뱰'�{��袟� >��������uiR+�aN�r�tOln^x�ͷ�hC�����{ѮP�{�/"����tx�5��ZI[��Zi��DV�)'Q~H2�D%ٕ5�%
-5:�NJO�u@��FݔBS!�����W�֭��.N�0,�s��\�h�
�y���lO�mTgi�wL��Md")?CR ��7��&�����1 ����5�`����]ǥ����5mG_;�x}��V�4TT્�M2�<���ᨁ#�MX��|bqL+Og�Z�`�p��T������Ψ_*m���S�F'�\
��E4�E}k��O�y�Ԯ��br�%�f�Xi���.2 �I@�kU�Q�Y{:ߺud�7z��az�g4cPV�v�������M*f,��E�I���y ���x�n���h���|��w�m�m �O�������a��4�iw}V�4��
ٷ�T��@������?2G�$���g����L��DOU��	e�^�1Oi���� ��@%s
����S���`�9��>t�0�Q�!c�oSF(��F����k����l�X��ym�$Yи�A���I\��
�����;G�X"�� �������:����