��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	���uYC�т��j_�M\��<8!��a�n2����b�����`L�W社.3S)��n�5�^���L���$fVVɘ�돭��g���~�|���$���Xj��Ժ���H��N�E�92��4T�S7k{:�^'DΖ`�-CV��&�^NV�<���Y���tga�z���>�:q� c��0��{w4I�6(]8�������i��'D�Gޙ$��=��vp���!X*\ס@)\c �]�AD���&53��e]���eG,Bww�Ez�������ÏK�1��;_1^9&�1'�9�0i,-�y�6e��r�ZN��QF��i�Y[l����^�A�N<�w�q#�_��U�g	l	����T�K��zP�;͠W'棯q0��.���F7�/Z�}�xR�lv��48d�i�b.�3.��	b7��I�d��v6��b%����Q[���b&MV��,��RM,��a&X�];�zy��h�f��rJ�,-)�^��|�WXH��{�Oc��0г��@f�,�C��B�Z�KsjK�S��ӱ��3V�Y�r���� ��0\ ��Y��ӯR̾�j����]��j����o�G	-ih��\�G��eMF��3$�Zm��A ��(���ǌY�ظ|6��1����F}I���&-�^����ڃ\F�f���%�Ћϐm%���n!4�)1���渼��/��*��V�)��ڢ`ԥ���� \vO�[PXt�:��� �OW���{�S�D�S^�ɺ��11Dօ�?DR�A&CN�Ww�vT.��@�^��N~��Z����װ�U6lL����\������8C�g[�olwi%���2e�����Pid�|@�"J.��S�6g���x66�C�RwH���4���=�o[�|���Gd5I����r1Ϻp��QzD�3B���P�I�#::��S>�L�Q:�N�/�u�Ƣ_{�)��L����(�M�*nAy���g�v��ȳ_�F�7��@���bIB�L,7C
����8|���5�An��q�/�	:L��΍,�V�a�ўY�����\K�I�3fބC%Ir�{QVE�G 2���~[�E�����E�¾ٷy2�8T�J
b0���9jC���_��U1s��N�N�R��b������m��sn7��35�>��Z�H���.�C�+�p�\,s��Nj�����q��\�V��o3�
�Rl������SV5�s�P����C�n}T�߄���2i��:~G;\Z"0�����5����v�����p�Ko�u|2�i:�0�n�����ܳ[��YQ8}A�	tK;�����+}��D�o�qҪ��i����5��ڬIhv�lp���嚳,�&�b'��?Q�F��,��=�؋��:��궛�q�QS�����u�;���I@�F�h�R�3eU��R���|�nN2�}t�9��.Ø���^����G܎��"�(	�
�ͮ�
�����M�Iq�3�$����4mzG�|#�����r��d�i��:2^^lRd��ܜ�ô� n$��DP�X���%�g���(�~��qcv��$x�}�?�eA�5��qU�˒�jʨ��)�p��[��P6��H?,�)(6�[������T\���8�n���C$���,��lh��� �Af[��0�>�|�A��	qֶ�ѐ�N��k�zx�K�-��@�q�@��U�fdC�5��k�� J
��?���k�0�^e�색ƪH�N�1[u>��M>���VǬ��D�nR�]f:�1ʉ��
��i������p��x=��*P&�\Ԟ�D<Vv��+Q������=���!�)x�FI�{�纤8����w��r;Q ���IX��:�7#z5m�F u��f9$x�
�.��KeG�-���m��x��	�$��6@>��un������_�}g��|�F2�PΞ��F(�>E��/E����x~
;+��'��M�-���ފ��v���8M@��,�����)�#	{,(�s��Y���?��c>l憫:^M�4x�k����a��YӀ��B����7<9dLԑ�Rdv��~s�͢�d�����র\�� =~۶�/Q5'b���_���B��Y�3�CE;Z�]�z�tCcg�����#�4�����m,���	��0$[B�W��z�uz �e������S���G
*	X��»��Qs��t�b.��<�Y�2{W����'f!Ҵ�V�=i��M�$��?�W�w^RR�+�HX29�;h�m�6�呬H����]��K}:�S��,��f��f`��4�X��c՝WR�)e%����@�5TG�p�վ���͡�R�:�2F�i%8�9f�2+ �DhQ��ޖS�픭�dm<�J�ҿ����\:VX�5 MrǓ�@���g�1D6���`̚�R�G�rv~�A]�tHi��,2��%.������sb����#0C	�,Vp+����6P)���^�߀䎯����)���u���>M��>�g9�X���lGF3`ߥ��N<o��m��r_`����{uZ�:�����21�cz���=�`,�Xv�� �b�o�sޡ�6�d2Ib���f�����R�`� ڞ�&@�D�#S��J�E���C��t}A�y8���5�K�D�<��cH��_�79eFpyG0���vF��!d�˱*�ػ��)�{Q�L4�^�ŒG��g�j�bHzȡI���8�<�2����Ė�]h����Z�.�{���>��6&�#�Rxm�nI֏tA�����b��jd�B�/oF�A9Bc1��B]���d{�������Jf�9��q-�f�M���󵘘��\l�[�"�dGN<���L���W#¹C���K9WQ@��?�kы�Iq��f���@�+�.�3������E�҄��C&�1�|Kϔ��-�Re��wy���%�9$a4G|1�wB�:����qo�&�h8���h|k�&�nA�Ǽpx�{r���r�K�����]FQi^��Y�;w`�>&��o��6�1y`-7��,�+$�����v~�Ũ2d��Ћ�l.������˿�с�p��X6�7��I2��Fra����;�f6b��8lA�M I[�eG+�#3NãK�wr��H�-x`!wu;�y�R��n�t��Rt���skD!s<�7gr�9.�M<m�P�^�"e��?jt�`4��-�b��C��X��0��8+�m ��#W����˒�`����o��(�<��7��:�Y�Ad&c�b��xv��;�S��@�3��|KZ@�n]��Ν�Jf�F�����"4����d����x�e�b~@��B�̂a^PNZ�f��j\4eWV��g�E�����go9p���́4@om}ʄ�q�`�w{�&�B�,U��8BȽ��J!R��M.4�Kv��ʇ���r0�W������������Ɨ�G*�z4#�u�0�����XL�Q|�1�M��߽��.K}!<nL.� 18O�^,RCq'����	T��n�f2jM
H:o��/��4�Ye�w�+u�PX�N�I��
���	��E�����;÷����3�-�K|R������]Z�n[�ю�TS��ˋ`Ǿu�R.1�o>����O��f �qmyc.�+=�&P+�
Ꙛ7�cd)
p�X&x�t�ra�^��^.;����k>��1A�1O�p�F�FO�_w\q��\��Fm��sP�_��}\��&+��ߐ�c$���si�``���v�x趯!Y��B�bo�\��gS��e��f�8NM�R<��Cmj>�@�JGX�����Q�bc��av�xeX�����T�.@pִ�������j
mh���{�����.���8�������f̸y|�֢��MaE���?�A��T�	��K�x�^b84k/f���c�#C�O�C	����=MQ�m44Kռg	;��kz4��Ğ���On��N΍�kH^@�eå�͈J[G�sU�p�&���n�����(�<'�0F��B�&J�^4��
\��'9�F��5dF��w��	9���!��$�;$���|��n.`1[_	�3&���ⷬgAp̨zJPk��#�u�OsVN���w*""gsm>�T��.���`�	x�Z��k�Y/ ���G#W &�%�
̖�ÚS�9����V�U?���i��$o1�95��jy���<���� t�=d7SǸ���9�H�K�P�m�F~2]��Ɩr�\-S�4 �E�x{h(Q�]����@�o�`r���xz�/���є#�%)34�-�y���n'~9�s)-T7��*Ɨ��|��˴<��KT�ZNcѿ�Aki���YHLm����n��T��6�k~�0#:��ٱia$���3Mpl0�a�`�˸R�:=�\1F-bɫ�Il���NK���2ڻ�"�v��(���&�{�0ק᯶�Y����
fG��u����h�F徆���;0K�?� aDx:
l���U�2r��f-�d��a�X�����K]igă�;$s
b�g>�ӥ��V�L�&�+������A�c��o�0�I�+̩�n��N;Pȳ D,�������М ~�z��N��>��~R#�Y�Ȳ��˓@�R���<+"���1�b�L��(U�~X���I��]ͦ���������7z06���Zh�l��L���S�>?�]�ȥG�0�Eq�x�����-6��\�D�A������2�I͗$�Os]��^�z�eY�k%�!]\���Y}�&?��%���v�¡��+Q��EU$(�$��)����h��?{p
�ͬۿX}��_��0�ᓸW��Fٔ�cq��~�����汵lP��	W�Z�˝�W>%�>=9ȝG��lY��_�3{�d��D:�o��e�V�T�c������ͥ��1V����d`���d�k\Y 7�M�"h�h[�l�P
�Q��'����U�NWrO�	�۩k�X���T���*���%�+�a�[�IR?�Md�b�������3� \�E��ׂJ��E���!�-y睰^���'S�TXJ�Q(�#o�<qe[��*@v��U�9�vr>Jd�h|����^��d���O�Ş�-j`o>6�*� ��D���S���d.��B���_ٛ?�c�ɞ��m�X;.��̋��@�φ<�'���O)��lv�z�t��|���emԂ�e����
��"�Q5��i��y�У7��;�����rn��Z+y�R�j�4�����x��S����U�b�cbU�3� �/�p����a��vg�Nթ(�"�f����ZK�>}ܮ3a�Ʃ+;�ȉ�pR��H�րc�O��W�	4�E6���k1A'�&\��;�>�����u���k%;�������R�a�1�#���$c�։�����?{�������j����2�}-WB��YLd�D튉�*�|v��1���7^���Xעb�M����&�
�;8�?2՞oR�I�΄7*�BoS�>+i�l�?75�v�����O�K��}(:qHt"(R$����5�F�V�υ��wjnB��a��gӪ�1.�FJQ~Q�
�Z$kr�������Yߺ��3������x�SCU�͑�Φ(V�Z�ȋ��5�0��]��O�R+�nߩswƍ�pw�B ��lN�Ow��2�Wn'�a����6��_��%�<�؞{��^��*�g�L) ��#$v�	�]�u��b"�o!~EkS�2�:�"\�6Z��*�h��p7�!���)�B �>�W�z�丅�S��0'E��2��������ՙ���W�]R%�>����P���g��1�9�ل2�g�P�m{|�>g�<�O�r��S��'�8Nǉ�0�0��jnC�-�J�U�Z�q��sL�d�~�WM�����+4]�ǉ$�)+��֗�m��+�V3%�ա�H$�8�����i ����k��$=-�Rm�`o�I�U��.
�-���?���m0z��,#�	(�W0_+V��|n�4�����x�`��M���1�R�����=1�N��V�a�-l���^����9�K��ˈ6ˀJ,|r��9d����S��Ǆ��y�3]�:����2����b��9��}��Ꙏ�ʮ�� �P�>+�5�ur��{��)�F�/��x��U��aP�u���^ �a�S�g���JM��|�ٚguĀl�c�ki�8�vht���}���S�e,-IA�3�N��-��,�,jqFnF��M�Pk�H>�b�
�_�NtvU�оe��%+�8�M-�ّyL��z�ׯih�Ҟ�*_�R)�Ꚋ#�B�<�Z�3i=�@�,fSB{8{���YC���`���>�I:���B�G��P�̔Ĉ�
;l�h�@�����1�͒~z�O���A��O寨'F�N=d�/Cd�HH��p� ��x�Lj�ЃM�Hk�,q��o�pX��e��ۦ9�孉Ϭ7���P6�R��gJ�� �nm��7p�j3䨲����Q]8�u�O�]+������[�Z�XE���Cհة��5���b]�Y��5CΕtj�����%6UM!O�	�Σ2�p�f��z#I�C�d�|�>(�� ?��1Z3�[����w_3Y~MN���c���j�C�\�}�xb���k��Xw�C����:���C]��]8/��
}&'�I߯���Dx����#���.k�ex6an_^J��n�5K߀��O�&�;i�ͩi&Sx�TL9D�����b) [�6��vC ��c��՝)=�=1�@��Ey������&v�`��}b�I�l�Y�5��F$�h�.��� �\��1���1�~�gF�|�n?t���?J���]<t<�5�zq�E��`��;�&�T��D_�z�_3W��B�ڳ��g�;G���P��=��I�q&|m�K�0;-���
#������c<ѹ�{d5�`�2j��Z�,p��t7�.H�e�K� y�]šp֨F�b�'_���]a�����H��z$R��Y9���pt<��9�CK�-������d�R竿�j���J�_�h�����s��q��c�B��fV�\�I��	�?�J�����Zw0�=NG�*�����]P�����Z�2������9�1��	�ݵ�f���Aז~�8U�Q�>
�.�8vt!6d�x�.���V �?v�5���'��Õ��|W8���=G��&��Bq]Lq�(�S�|��ћ�4� �팒�ﺓ�՛%�n�g��g�嶎��Ğ�<� 5,RM2%��/{|�m�q������S,?��o��s˨�;��W�:�� F�d�qE�;/H���>�E�P/�ד�y��4��FMs	�;V�Ś:ح�8F�o*Q��unL�^��K��������#���z�̷�y(���v�CI��rܽ$d�^�TO�
�u6N�NY��>:<� |]���d�it�.�Y\�<j3��v��q�X�HtYI�R���Õs�C�:=$���ȏ�Ju<礻��z���v���b��uM�#��AN(�E��c�>;��R���A�� �1��N��^@�U���P�T�#l�z:|2�Տ~�,���ԛ��t���mi�U�5\�X!������c(f/r�����WDLt��~���9'0�А#e�:MG k]�J9���iӤ�I��[�C�z��������z��g&NH��	������p̯iYR�z3Dg�t���h�APw:כ��b�
���*��4����* i}��W�b^�pJ�.��>6�j��狀���2�B����^Q���K�1����k���(¯�[��ρp%��,	�{�z�\������N�ǮM	��D�O®ޡ�/���(m�bS�<wJ~Ƹ�Z�]��R)v��e�9�8� �����N�^d/��2�\���*Ѧ-�bNmiB%��n����%��b�f#�GI�J�%��BS�����V��։
�%^�֦�t(B-C��R��#�]�Yˋ�LG�uC�j� ������[�i��_����!] ��Y}}��g6CrU׀��E]+��M;��_� �y Y�4ʌf�FH���,��ρ�8���H�a/}�z��w���U���HnN>�|�d+*�k�jd��}/dHTҫ?G�k���@U�8���7tj��&0�_��`�4C��J���¼�'��=��>?��݉8&��Ҏ����N����G��#�_��
j��t1a��;�����Ѩ*�D��*O^3�r�������g�C�Z
���M>?�x_`JS�P~��M��o�����}Շ�
��bi<�?_�|���gïOk �,2'��T��C��a�Z]������z
���ϴ9��x��t�ʱ����-��l����%�l4��M��93�N�"��  3<�cLSL@�Ln��+'M�rt�:E�̤�"����~t+p�)W�U�v����g���0�l�fgY����-��t�U�[�*���۝wY��g����%v%�I0�r�Ω���4Ł�9-������	���R�R���s0c�,��e���C�z�҉�U��0ڻ��L� �#_����;)����˨�*F޻`]#��v�Q�j�ǜ��`�
V=��!Z�����
�V��*c�Nz�!�<&��z���-MB^�urm& ̵���(Ӣ���d���*U�<�X�̚ѕ�ѵ�F�t�vF3�yɡ4n�ۋ@��yi�g�"��ؖ����Y��٥g���	o�cet�/�+��t���s���lw�o��>�� �ş��Y��S��8Ms9���RL��KwԠTQ��P��V����A��m0�`�fe�B�4�T������_!�|��j�8��TJ�c��2�nR���e��Ҹ&ef��	x�����<Gz�Ur2�3D�{�M(WX���KMw�=?��o�X�wk<.ÍS)C���>�8gc����S%�����;k�̐��� u�`�f�TA1L����qۊ
���CK���(��j	�`�]�fAQ՗Y���[������s�,�S���qf�����ϣ匡aF���뽙98l�udT4/9ؕ��V\BR�@y`Ã yr�7����ʧ�MK��@��ﻓ���s�ԭ_���O�0 /D���3���+�����/ͷ�lo-�\�T�Ø�Hvƛ`B�eZ����H!`O|����u㶞`�.?�#N�a��BT��&ۊ��̱��
V�qu���z2($�P����+��vMPJ]Z�o�Q���[��v�������$�nT�\�����R�mkwƦj�RnnI�`j?������m`��b���vhzab� �T�wEu��ׅU�CD*�zs)��|��_�hcz�g`���l��b�o4��{�8������j1!B#4��!s�Uٲe��.�Xo�0���Kw�"���[P9�g"v��h쓔�7���Ʌ�"��{DAm(�n�ģ��D%��ԍOs�ao�bj/:I/���S�hni�Se0t��� �PR�,����$�./]ol�� ս�]TW���߳�Q�烉�P	\���&8R�<k�u������*��8�I�Tmٙ�I�	��d깛��� �DY��q���ȝY�d-}^q@�'/]�_jQ��!��VɿI]��c��A}]+�Ǟ��M��~4ʽH�|���'K�C@��|D�֙��Js��.}��R�_���z�/O]��:�	[�
���ri���,S�~� @Ԥ��썗�����w� 4d�/���=`�	ￏx�-n����g([Ų��"���7�'�"3�i.�TB����eӄdԒ+&�����GXvY(��/a7�|,���=�� ���5�$G5�SB�^#U�c��+d�i�_I9��`�x.#���`�b���A�똷���,�F�ɕJ��R�O��W�ml�OyS�E�&�g�0���WYM/s]�B��aV2�\��a�ޘX�q$1L۪��U|a�~��lQg��#� %0�R�&���@2��8]��%���ܬL�`�G�+Ur��K���9g�j9�7cףҠ�A#'|�L�Ë@T늵������灎�����5X�\��#�y�]�EL�"ȓ*�`��	B��C� �Q��w+�x\�{{u������'�l��?l����0b�v,��Y��2}��ɝ��O
=OD��"H�M#9Oy�z4=Z���L�(�z��*�-Y:ڮMEyOt!(�t;G<��&gs2I�h�p�rT�1�\b�@ھ�, ���VP�}�d�n9�v���=�q�`�5Q���,���`��_/�0�D�"�R<�Q�.��>�g��_��=�����h�\��'���X����)L59B4�Qg�hHd?�N�g,��0>O�fgϓJl�6����A:en+���}�y3�Ý��iB|A)"+��ԋҽ�i �8������O;O)�t+�*w$�����ܨ��p��vN�)��eIǑ�^b��o�^	w\WC��$�~�*23���A�V!��6=�-�����E�~�+��ڞC:�7������^a}M�IM�6��`W�aE�l^��0�$�o�h�{`	�W��6�`T[����@�����0˵��=����'��l6Smˉ�ِUv�g��e�~^�7�ꏳu�%�����3g^Һ�8boV{��A�Lx��E���g#�T�zw�- ��������\�C���Kk8��ʚ���UK]�`Г+cl$v�M�@Ї8���TEY Hݼ�" %@3�H�μ,���?��Ę��D���vFY�L�0��u	�~� WLJ 1С�	9�@�+x��E��OP�Q�Q;v}��������w�wr�N$��DY:~X�M߈�Z�岃0p|W|0<vc�9�&��k4�w�����T��8%B���!��&��W�%N�`C�k�2�{�4TY����|������= _<]P�G���kMZ�)��V@S�D���2� 4�v���KR��D�����Z�Յ�����PV
׌�����X�GT*l�C+~&.���?Z۸Q�sÀPKĀqI��!
�&���u.IK ����Ѭ�_�rE���	�-mO��a�%��Z���}�1j-�9p(��k�m�f�z���YzK�.��ɛ~��5,u�'����yls��|&�l������� ��>#;W.FEGm�m�����t+a���^F�n�lJV��sW_?��F�uʟ!�8��֖~�١W����.��FB�����yz(\K+�^uIl�V�����]���^����o��J)��L��	(yF�D9k�H�7x�*˽ɫ5۰���¨�*��k���I��2�^<����DGn�F����$�2�#%d�m�Bǐ{{���4��{h0�a�J�ø{���{�A��D��n���ƽk���UFQ.�`�<R�NF�֩���8�ny,p��y��MG���8���!���D�Ŀ'wo�ˡl�̹�T�������T�������`8�ZA��`6@s[����A�dM
�7���D[I�m2�����T��q�>s�|���4�����k��r*6c!�p�ft�0��pGz��~�U�ݭ�h�rA�z�Z��
X��z}��V��=��! �=�:L���1���bsq��ߑ�5貵�
������W� !U��p�h�N�~����B;O�}$�e��<�Ap��gih$,��$�J��/М��X�����
*�1���2��n'N�I􋎙��t���;�9�+��H�!n������ps���:�K؁J(E�~h���WL�9��b��zޠ��Ze1�y۪��� W��&mkN�4xM�{|����L}7KvӞ���$����`ө�rB4Ce[QP�&��	����"@)��ʈ$��́��� f7�ָQH����ݴ�6yD#�p��/5ʉ�=�ˈ�D�"����P�Z� ��?s
H���p���o#���rᐢqn[����Lq"])"��(uZ_)��+ҡ+��E�}HR�Eפ�)fF�©cyW��ș�y�mV	��x�/~1����7`��/~Mv6�i8"D�ߧ�>���,�ĠVՈ���Q�`j�����VQ�U�%�_R;xh/%m�?Yf��._��|����ln��f�ZFե�zoj{P֒�?a:]W�c�������-��Q�Jg���9�چ��Lw�7���� �l�򽹡��P]�������w�p@/��= ̻I���!k!�j�>�	��a�YZ��Ƌ���Htw�b��)�D��G��Wj��U��!��	�;��,���[Ӡ��2@�1ц�V�B}��E8?�j���&~H���Ł]
�{�� ���������SS��uAR�y��b����9pQ~Z���� 1�Ǻ�Iw@�?Y�=��T#���xYL|.
ST9~��������̘j���SB�K5..��w���&J��.���5��dd��͒
�
o%V����3�1bP	� ֙{/�z`��`/l�,�!��Ҍ�l��"��Z�8۱��\��%3����;�r���gF�l2b+�H������#�89�� L��@�]�>q`�.`��"g��*��?kq�0F@�3�q	��{�Jx�$�T�Z��։A��Du$��cu��G�$��2��AlG<bG"Jv�[%e��)Z�	*�\a�Ǵhc��V]���g6�
X9�*�*~Lu�ˤI3l���h�>a��#@�y��M]J��Gr<�냋�U#D�Y	zX��֒��7u�7�A]E:!'�ﭣuVڢ���$�<G��JjS.��Β�E��X���Ʈ����'�QЮ8��є1�v�ds��s����YὄS�w�$�
���bBr�9P{3o+�������	%����U��z�!"/�%�'h{�qI�)c�
��H{_������hd*�����Y�Ѵ�w+Wzl��hjU�!�a'X�yv�RK�)��&w*�;;�}���:b	-Mz��_.��,w�.NG/cn��.�<�Z��ϔ�V��n�3%�>��|�94U?G&t�q]�]��8,���|(���,�*�2�RnI.79����f��ف�蟟7Ț���K�����(C  �$�*���fk(犵�>Iʹ-��!�ĦR�0HE��7}�
&Qf�����Ow��̻��Ϩ��o�f�3�w�|��:e�і&�"���Na"�M����wvi7���h���'��M�=�l:�k���~a�[�K����8ׯE]�'���k�^�n�9���qy�6�����|G��P^������I⨱7���F��e>��,�\�~�s�*�֎x�z�5�����/wS���q��B@5"�~�ӅOL����l #Lb��dB��:�68�๓���B��t�&��i��w<3_��:Sv�!�G)�����˒b.iq�<�j��>��oʳg�S����vЮD0h�qG@wB�4�>e9dK��ʡGe��#��n!��2F�a�t�-�'*�?MƻEIV �A���c��{��=l)�%)�o�$����� Z���lQ��9��":��3�ol��]�쑺���K�"�Y�����;�k�<����7�~�	�sQw�Srf忖�u50{⏬j9l��R�!�}EA�{Pg?�� 9����~Ӌs0kK�n�^�8�H"�(}O��3�^�xj�_T�H��X&5mx��롕vQ��F�A��V�w�pD׍$�)�w�W�5��=߲/�u=o@�l�D:�a������!~a���xeM�Gx�s�e�B\�E;����͎�T�(�&
�2풶����ܗ�#��������p�Mm���G�K�q.8!���4��V���;��`,q�1f���V�(�
𬩙�'$�0ܣ����{�s=��u���6��Yt:������܍&	��k��Ls?���ן���!���bcX�����<�|�e>Ϊ�
Y!c�?,�q�UF��eҀ�YW/��⤕C���6A�����1v:��n���,9K08,��
N�@�����IJ�����^����~�p��!Ѻ�O�:�Kz]BH��K�2����q��P�+�X���TJ@4@	Rĥ�Uk��XGi�PaZo�u/�M��1���`T�z(u�+�+�M5�]����w�\u��C�NRC��kq|����4��͕͗
h�\��Fhu�}n��Ւb7�c�8�3Kڑ@	Ġ��Q2�b;���p\3�f�7֕�n=81#CTI���N6K,U��F?����ń>�K�]Di��wBu�b#�t���}3�<�Zw3J;*�e��� �|Bl�U�\,Ͷ%����`"̛!�/���p`�Z��i��t�����b
ъ�78��j�W�
��Z$Z�=m\����(�f���o^|(��Ǐ]���������!=`�rt�$��rȏǀ���S�n�/)�|���]e��Jo�SK2fj�SyNt��ko����*r�W$��#΍ ������A~x�b����?#�j�ח��rv[Wf*|R�hJ�Z����-��7Cz�����y�=P8�-VK�Q���ǎb~k]�ְȞ�K�H�R"S�eƲٱCnzeY�(���]zL������ڮȚ˴@�u��<�k#@g�I�&����;�'��,�1j���6�4.�Z�����7)/�כ4g�I���֦�;>�	ba\;u�Ev�Mk��L�-Gkr��Ř	�6?#�v�6���'��o�`�¦��%��Q[z��1C�;�9C��pqH��w����\R�˸��P��8v1;�=����X*2���K���^�m�a;"w�։�d� Iu�Ϡ�C�����	ԁV�)���9����
�Q�:�5|_O����]/%"����u�~�_�����Ǚ�kO���	Y��9f��-��@�eۢi9Q)4յ�!��sN��ɾ� @sn4Hc�e�q�=�A����U�K�+z	�sZˤ}�rL�4Y%�K�Wv�BLk��j�q�
P3�ߌ�'h˩*����Oz�ݥ\B�Xa�V~A8|We{S��V��YM�ҽ�ޅ#�+�0��o�y���oޤ�`��*n8��If�A4���4 y^�
m]���@�"��-~ǤWG��I�fe���mL�_��fR�y�Ǒ�h�&ƒ �!F�P�y���]e�f�ܞ���b����Q W4���ʣ���sm˗lۑ6V�� ��K�^����2}?T�D���Kc�>b��2R.c�J�;u���Y���H�4�1�k۵?.�y�8�q�����P �o���'��5��^�K~b���fH߽������`�䐙����U��D�9k��w�S�m��a�1�����5P��0?�5X�a�?F��Q�j/2]Y&uoCi�,��*��V���)�xd���4�̂�y#׀8��˅�7<�zv˛u(�
0��m1N�U����3Y͘����tw7�d�y(bz��5�7�(�u�ED��'�����iC�..X&�q����[����N������\���
#s�����3>oz��o�a�)̛r���!�~*;e(��gn_�#'��M���$�Dh�O�X$.���(��mp̀X# �V~b�0����|<�4,5�I�e�S�ɛFr#���"�����	-��*��}�w�	�.gg"�Ǎ"���Ū�����G�]_o�������{�χ�������~:�$�j,��e��[�T<�l�fFT�m�d3$��w�7��	 �|Cs}K�o���LK9��q���sn�����	��B6�N�Y�?�C�q�r�t���zA"B�r[W�p�JƦ#��9B�lHH0�������v�)"�7�"�>���K�%gD�Cԫ-�Cl�=~;�2¾1�LF�W�t��g֨��q�m��ZY�5u�x��fo��$z��Pɰ��4ϭ������w�o Ke�Y�۶T6�?�]�=G�O)��x7���� �8/3��n��W��4o��x!�
��>ă>�	�ce�R5gŢa���DR��$b'�mj8�~U���N��q�#5��Iٝ��0g��Ư:#��5چ�oo�
;-�	 k���K�"�,�F��� b��@b���q66&e���nv$������7��N 
7���@�l�M@�$�a���,L!�ZMa��+#�G��na}ў�=�(�[��17>lm�Va��(��s-�űR�`�~��~
ߵ�{��\��2ׂ��h���#���64+أ뢸W�~jJ�H� 痽�}�s3��B�H��s����b;��ҒG��߁x��i��]q̈́�c�N^�A�^�U��ȵ���Ĺ�D��_m�ו-e��Tg>����~y1C�0JőA� ��zyƲF1;��3hI S��i?��|�[.*�&��:.����v���#������ P�U�[ڑ���N�Ԝ�i�e����)-u�Q�P6h���ZAJ�D�Q�f���_SI`��6mͿ�!(�`x�ҦkFY\Oe\������u� jL��g�@~���ldc?Y�Q�9ΡFֽ���$欗ke��<.;ȧ����CeД�zP���x��t����zկ���S��lWz����
�sv>��5��u005�N�n<AU��k,M1��|�=��/Y��P�m4�!a�{�P��l��� ��Z�s��$���e��/F-;�{�)�g���*'�%�ǳDy�w/j�� ������+���F5�]m��>_`TbY�ֵ�Z�$����G�K)���/d�L*4Ugᖶ�b���Q'\|P3̱`��o�XG�M<��.f���86,{-��GA��&��D�I=o����i��<I���E�gOs���[�:���
�����s項fL܈Kz�q>��A�Gt�E\�=���N^�̻O��)�t�^x`�T�y?W��8Łvv�(��wJ�N#���6ˣP���9.��8a��1�/bX^sB���n��Q�U:��(�{��ʷ�HzF}����Qq�������& pk��I���Νa_�����]&Y�g(�ǾA��8�3��c�Wx��˕�*k�ݺ�e�}0�lBlG1��Q;��w��$?��9��.�>�a�h�b�Zr$�\���{o1�ݏe]��U���S�(�t�"ܤW	�M$�Zj�F���#�^
���W�{�`��~�z�����{0�3CJ�ݬ����=l-y;J���po:9�����hvp7'��evKZ{�(s����)xBz)ƶ�@g4��yX8]17�s!é�QϞ`�����C�?��ծ�M�"Lt��H�~j�J��_�Uu���}���1}v�ȏ��#%ڎ�� 
��z�-�}lc��,�TR��Co�^�fr�����K�4 jY��I���m�=�Vأ$�X���{$�Ȳ�a���{dz|3�E��]�� �Pt�thC��JR�a��yT����Z�\�Fl�k�@��&�%��\�+����%dA��,1�.7��haV\����<��'�^��
�xe�5������4�#ūi��[A���>$�nGx9�+��0�	Djf�CJ�ݲ�x�,���A�.v3�m��Y���H��iN��^G�8���O^�?'�d���c�8���8A�.��٧�V����;n[񊅎����/���-!)J��&]"]ID��#F^:��z��&���QZ�ɀU�ץ�Xy��OTVrL�;��ث�	�W��l� �m�Rd*+�h�����IR�����!�,�Rh���4Q��/f���'I���x�&�Y
5�+0v��r��х�P�U�<� �1��q����A%�r�}4�������2��F=w�E��H�d���tNB��B��SA�;���Sr}����VP#/���@X�
�?+�ȉ�Cl�.�"�LOYy�����YJ������i�t���T��I��#֝��d>Z�Еcj+������6zB��&�iFn|�b� E��(C�z�P���x�3��]�GJ�rמ��TI1�i(�Aʺ˳4B�@�$YP�
�����WC �����60h�ɂ��(
������H�KW6x]U�9^�C�;�)f�Ҽze��4s��]��j��"}�$���J�\c�P��Q�R��ڿbs�)�{�����t�����Q]؜���8���4(�2�sߋ�K�nLW۬�Q����vѶ������+f��.��ñ�|�b�7r����^�A�`��߸��wh��śY���%6Q���qW��ܡ��I0	u�gU���cyb?�O(���Pq�����M��\����G�	-��&��[>��Ӓ����}�,bNz��FE�|���\�a�N�����@ȑ��?h(L�@r(%�;���y ӑyX��g� �tm���Г:���)-�:ƛH!�������@��ح��[\�Ӈ���菸j¹W��ΕP˖�ɱ���"M_�d��5}�o�XW��L���!�+��L�0���Q��b�~䟗s�����ĤX�[C�1��㌺�?9���]�k��;����5��j�u��t�z�S@��DR��F3H��C_�o4�j��%S9Bb��8h�Č\)o�j'G/��ا������-[O�YT{ .R�´Jo>89-�DكrSv�2/n�u�n&3���gР�����"N�a#��u�u�����ǰ�+lM�ڒ�iQ���a���L(���ͦB�M-W����5<Q~��30�FNV����47^DbM����Prm���?݆�F��s�D?{��.�b
���A��P+�x-��C��]0�CrZ"�wZ�,u�f�.L�]s�V�i�~lrtئ����������JQ��g����I��kJ�F4�����q�L������H��ӷDhh.U�G�\�>�A�ǅ�%�SF�(N3:��]��/:[:�k���mi���I�r0M ��s�.뾆$�����j�����l6zā����fw�1��������ݶ�����u�W,~E�ݭd7�����#����Ȭ�8Qkp��k��!q�KX/�i�=�'m��$��0ܯ!�*G��򪗳`���L��{�dϻ`&����c��ް�+b�bj�=թ23��%6�����?���^�e芸j���3�d�v�Kz"�	�׊7�\N��Th��?��A|�+![���%��,]�jGP�R�W6�8��
'�h��uya,J}����̃������YbZŖ<a��O JoO��8X�y�����H�x}#���^�6��k �cɧ����v�P�	�����^���m^|��/!*`�M����*'Q��K!K6�@���]Pw����և�8���mby��\UfҮ�@���o�?�`������9�WsԬ���������
�����.��ni �ٳG������I�1���}��^0ı���E1�i/U�΃�c�-l���ĸ~!��i7G���!Z���*p-�bT��=h�w��yL�Xp����A�S瞖��?c��]�;��~W[��j@FΆ�i�"�@����Q�`{����.%�Xh���f�Sv�M�p�}�R^�d��L~�cg��e��~k�E����_���1�[x�vN�bt4��|2nk\җW�������s��_%�3�;�R� �#T�M�mK-�Aȉ�71�,
GM�[�����[+Zc���z���qw��u( @�:���pl�P�:�qg={F8�l_,~#���7��ü��Y|�R�&���#r��2��^\-O0'h�7²Ckqyܱ��%?��PT��,p������}W�:F~�&��-n��s��LK���zd�Lq��[��;~̙���ϴ�2���B���7��U%š�?�D|��5'lf��|����a�S8�IT�/��.�6ц����qtP�CHPm���;ň����h�6�P!��Λ$ܗ��j��:<�˵�ע�S�2���\]�����)��P����LC���m��wR�ֶ�iɟ{��f������pہ3��m{�'Ȧ�KO�0�d}���I�U��M�!Y+�]-LJ.+�o��m^4>����hX8�rY��D{M�8ΛQ�^�M��Q:t�
��ŝ���`5�p�ދ)�[;Af�� ,m�ۘ���¾��K `����Y��-l���E=_Dq/`G��ȭ�
�@=�_��� �X��z%�ѽ[@�=�\�	�Q]Ǉ�j�&^��Ș`િU��w���1��E��MŘB]M~�A~|$�"Ǖ�"��`4\l��gX�4���=��֮�7]��:���!�;M7|?l�x�SK88�������U��|��8y��AT���D��'+�V 
BR*�C���t����j ^$��<�C�|���C�sR�38�#�&c@;��|�X�nߑ+���~y΍����E�a&��,!ߘ`F'�b.A�.�H�#�rFi�D�bl��-�\n&0l;�6�i��[�XH�.��,i��6�\S�Y��+UxTzs<.-WBi�����`H�Y@����@eY �8*U���e�{�缫H��@�I��A:\��P]���گѫ�"�QU\ׂ�}�ҵ�?j΁ͅF�����:�~�CA�U�Ʒb�q�/��C��+%g����g�n� ?��q�u@2k��v��BzMc7����S����@u�L�Y��� C'��bT	X��:@��jF��U���Zl8U���o���+����&_�^��>~��l'�Vö��K�D����]��LI�n�S�,���:6��D���Ak���T��5Պ�%��J�r0p�'�'�z(c�����S���S ��(�o�쪳��:yIt�q��=$����gxJ�v�?%�����B/޻a*Ugr�;ӄ�<�i"²^�S@Y������_hp`�9�y=�}����<1�m�3�#y��g��Q�)2n�j���񢟭P��S �v�"+��-�����.|���!�:z���?E��������\����!��Y�$ff�ʲ��`Y�fa�h�l~�k�ӫ�r��,B�V��7�O| 8O:s���fzt| ^��EK*��2�U�=H\	�����u����}�b��G�0����=�m����;.Q�i�{�T�i�Q�lԿe7vG;��=�C�)�5�t�6n��0$V��#����=�H��ч��	���0�<�ՎPe ׹�N�sIC?�1�geڄ�S=��j@&��07���Pd��č��L��� ~s_��n=x"�9ɛ��s���lZ��l�٘��1,����J�^���k�|ƚ4�r����;1��B1���;�HC���j�H��[�	WfhRFh��q��m��&�Kc�I����J5;M���[;i�G��	I�A�)ω#(N��lS�zt��&����n�b��#[Ѥbʲ�GE�9��uy#o��zo0U%Wš�`k���m={�S�(�G�P�r��E��ŒCt��D�̚�E^"F[Z3�h!��d��3���.N�%jp�H0ͯ��Hv�����[~^Qt�(e'če�-�-���.ũ�kPrp)�sw0��Ѩ/���5�Y�b*F�ה0],�]�≮�n_~��GM�����!4�+<C�;�z�g�i�ǻ�eߋ�`��2��/�(>��E�|�ַќ�m��ޕ3�L;O��p X<�p��fcσ��I:wZ�����,Hf"wK�0s?��`��ê�z1A�����D�_��.��p<U ��nѣ�Z}��y��ʞ)�L��[E���'�Q{Ri��_�FǄ_r]����'�h7�5B^���T-���14�s��/ɔ��s�T�'�@Z
�}�������ё��LټP{���
�pR�/�hs�^�|"�v��g��!����>#����d����k�Rz�j��Uی�𣪜�����Jb�<���Q9�