��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\Z�;�j�A�D���£�d����2��"y�����!���FU�������?���M�3�Z�Iʜ�d��YАVr~��4;>���9/Dن���B(��)U�YZ����v+P�LKwu��=]�,D���|e�j�����\$��xv�J�l!����{��MM��y!F��FC씼፜�ו��]�.�H��g=|�}�w������gB��f;�m�*�;�� �A��������j��������	9j�;��~�� �5��{� �|�2g	r�J��ǑU/�G J�Q����4�$�����de9%L��B�n�f'�g���r�vT5��AR	V���$4;�U<��7�]�bں��c��CZx�ȘZ��\�ҩ-��S��0Eo6W�V�M25-%@xN}�$k�i�2�k��9Մ��kծM��������a��r���|T%$بu�~.@;F�dڃ*�������� N�E��Z�Oʘ�J����>�d��;*)�F<��j; U�J��߈7�8qW8��>�(���e��ʚ�`��:4[�=��T�k7/���`�9 ,zC�֬/�H)BUɪ���}�a]�GjNfk�n��q��;���⧍%�w��m�ˆ��[>� УU
@�.8m�#��Z�6�/8����#�X>|o��}YrG�� a��HG���$� �q����)AѪ�Q8�.�� ���5���k��!���dW�Z9��Ŏ�o�ȩc�.x 30�n��� ������{0���1�֣̠1��X��tO8�uÊ�ޝ��3_�\�;�҅x��I�ָ�/l����%�\L%jK��!���R{���Ι�dL@}�?��C]3z�<�n�9���O��|*��?��z��SY�b�g��f *��1_R�l��ˊ�8sG<K�T���e���rKm/�%��+C���߽�?��D̥��)�=���i��G{8V�6��p�9f��V�]+)�W�uOI����Z���XضX+�:�7�`�����fƁ�"la�N�А=��l�����7|%7����'x�k��/�1�W�Jܦ���#�;#8ᡎ�bX��ĝ�8�@Y�p�R	�İq��1Su7�����U�:H�(��7�ˢi~�������#
�"�Y�������sB��ղ^0�!�HZ5�=���L�e
h);}�����d�{O����e��0TI�<ם2��n��y-�}œ�L�]�S4y22k��QEc�ōI����%�,�M7�V�GOG�˦)�X.�2�F���vp������"��خy�~�)��I�Jܑ��/����0��p� D���V|My�Ic2���k�^��uV����)cJ����<�D�4�1�0#r��z/�G�s��3��In`A�>�I��MH�z�F�*�������|�d�0�ѧѤ��$?�'L�#�
V���,�S��Aj+��ߡ�.B����sm��1w�p ��u?P���?8u��2��<8V�`�����\��o���f����<��s?Q&/D�|˗h�/DD^�]�>��v&P�'�!&_�E��U�P��rNX =%�;~a\BLU�5�-ɴIY+��(am\$� qKᝐ\�����[�)��Wb�$����6���ѥ<��,K̅E&p��ʐc���;�t�`K]	n�-��#��J��y�hQ1'�p��q��q#e�!�7�
+�;Z�>���h�����ъ��6����h�Go֥&GF��*��i;2w<&-��q�b�$U){�D��K9�Z���<џ(� ��
�M**�F�/��GR��c?1/a\�^�,��ӣ�
�z��/0�*�5X��hpaܥ�1���<���l�	�ł�4�H'8BRI�m�b�1���qʐ+���.�ǷZ��PF
)᪾=�$]������� !>�-��āVm��]m�>�4��t�=���S=r�|�@2]�`o%ݶ�����ar1���f�p��M�0��D�fEDDm�8��}��lUrY�q���m��e���nq�A����N�<8�"�c_.�N�g	0���Fe6Q���z�2�(V���^�����bP��k!��o�O#������:/��\{��7r
Ћs��է^��uxd�,)��t�*:�G����#%�a|�G�޼�B�&�x�髲?Ps�n��\%�� [�˧P�Tl��4͂p��Ʒ�F�*8�|���rZ� �����/��B]��$J�x���><�7��.�b���c�?Cu��.��ջ�2��N�b��v�&n�y��~$���a_����i!)�唦3Ƃ����wFm�L�(*t�5��������dY�H��n�E���K4���$���&��8��1��R��C[�.r��E{�8	
��Q��8��j�8�p�Kp��#F��>�wF��}C��Ro� �y��w�U����I���7�\����G���6�D*Ij��{�2�N:#(�1��;�����sa�]ikL����4�pL�-&����a�2	Pпɫf��"�M���L$����|�'b}A'����G�ϗA��Tu�v-��7�EP�}�[�G�������a�b+Bݵ�ųX�O�R����3�.;U��cDf��Z��k���&t8���0�C�)�*���$b�uDT��@q��/!��5�a?@ Սj_�
4\7I-�'��Ĉ1i�o,Qa���#���܁`�z3�k۬�1�^4ͽZ�sɃ;���) ;�{�;� ��>Ļ'���	���?��;:Y}Pn�2�[#*��{�G�m����[v7��<eq�*�����@*7B��� ·ca5ʷ&�����S��9�PgIC�:�8%�HM��5�=C�f��/���3LI.P�t�3�gm�� �]0	�T֨X�2�7���XC�W-��d@~R�8��߹\���n�v������a�3��v6bB����n{����0;���J�����-�	QЖ��T"�8�M���`��9p�_��6�^�¥5�`0gY��_|���|��i�7o��r�9�Y{�����*�w��Uy����E��9a�?~gt���/;E��S��srN|�u�++��S�9�7�3�	4^4I� �G&P���'T�g�k`ԃ���Fz�{���dNeI�Ϸi'������1��K�x�4[�7��ሄ|��ʊ�I/=���@���Nx���𮡠�hY���&EOBQ�sy��M�uuJ}�q6�j��E6���<aMR���[LL�m�/�j�dh�`��m���}3̅��q{�N�Fۛ[�^�S� ��n� �"$wFKSse�B£�"����L�*UF�yv��	�MIg�2x�t>f�؄r>�*-cV�帍���0�D��[ 0�6jQ��%����h��﷎4X����6���i.l�[8l,�!�
�t�ߪ�8�hH���� &W��#��`.�F��o��).F��}�����B��X��lg��=���P�>�N�>y�ӏ���Z��?�Ҵ6~�I��m�*��b�G^�f�B�߻ӓ��"�4EJ�؍���`]_|}g����|/�9HOkeZø�-�;�e�$>��2l��������"{E��dw��)�P0�V���k������=����߈#�u}�_�!���Ӡ�D����@P��&�Z���:��ؼ� a��g`&�V/w�������lܑ� ���k]�qD�� �o��i���<ⓔLl(����4ɏS�.��DDi
h���� A���x0��>9�����t��$�Ҟ�ZM��Ї5����o ��m�k�6�z�Q������!s7�$3�gc܌��ڙ�*���;r�H���樽Ԋ0W����3K�@�9��{��A�M뵵k����ֽ�(&����a���� Ԁ����%�5*�@K�G��ɟz@Z��y�_�DB�ǲ���A.�|t#ľ�3r�p�������Z��U�}��i��С�6ytE�z��v������ W<�VRB�l2��~$,�d(��xBL��a/سE�̏��{��M���zۡK+�Ԝj��o���S���F;Q��� �^	����G��d"�
�W�@�-��Z8��ÇK+��.�#�Z3�-����+B���z�w�ڔI;!f/�����6�HO����T��2�?� �D˹A(�a���h�ި+��?�Cׁ�������ꇍ^b����@��T��7�5_"ݗFř&���x��ǂ�4����kAlɼ��-I	�����+~s-$��`f���7%S
*��wRP(|��s��B(>"��h�a��YMק�Z~���9�-%dBq3@kW��~F؇�ޢDў1���?�����Db	�?���^�n㠠&�C:듒3N#��pC�&�t�j8[�ɑ�Ol����zл������(�/�~��7�~�a����#>�"�4!y񚙫P�n�G*���]$)c&S�ؐ՛\R2�e��2��tY��o�|-CAX>a,/�Q�[d�|돰5!r�� Q��l6m��&��ab���r�'�D p6�<±RH�(�O[����&�o�JL�����FD��(���p�3|�M��M(s�Ʋ|����N}w�g���q���Y\��zEy&4��(����DŇ������8V�\�XY�`�)���+�/�B���ў�W����бs�@g��	L>ō�~�O��I�������(4�t��D�R���d�F�A���Ϝ���'�a��j/`�)�zj� �mB	��?�U��]6����E�%�Wwh�~��Mw�j:{X#��Ts��_{�B����zʁ~��5�r���zYMWo�KkMZ���ȺM��-��;l�a4/ɯ^���.PW��<em,Q`��$�cʳd\��-OR֟	U�ebM�RY[>�/��쩽���/���(��F�%����@�%/@}��	t���l:9�ڌ4�
��%CT%`Qk����6��g��=x�:�RY��է���>���w	I޿����J��WЌ#��t%��mУ�`�G�$߯U��e�V��L7PV������k��*B���l����90�C ��v��cQ����@i���ȿ�'j/�g��U��k�rn\5��]Z���/+���yl� �U̴���4|86g�_@Jv���%ž�	!ڨlE�)�1T��{�����w].߈+J���׿��z���+�G~��|� hE�	'�驥6�/���eX�K����߁����2�ſ7�'��m�5����{6x�"o���O��U:c)��|�,���ʆH�D�~0u��5C������k���4�&#���J�F��n����D��.�5���&��H$n6I��v�pg-�]�9����o�Qn0��ET�eً3������LB�`�p���_v�;k:�|��mʟx���B��t��e���$.�n���