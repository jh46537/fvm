��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""���᤬����[���%r���dY;�uU^	/���D�)�&��
ux���26�K���al�N��hU��^S�]/����7$w���#�i]�|�?#�KRM�V����$85����G�������!�}/���2j}'W�mD�?���B������ξ�4���\�����M$��kW��U���v�:9���ut�*��C�ǈ��L�I5����aP��t�Z��D�#RVe��&\	4�'�!\��>-S��<8�>ߤ~ms�jCK�A��hG��σ��P���(�X'�X�_�>�2X�y�d�KK%��ق|
tk��p�q� ���g�����2�G�K�脠Xv�P^cL����c�\+P���FI����Ji�S�h �Ϩ��8�o�%�ӸNUf�Η.T.��d }b����w^�f�^]z<$C(z��9�|��M�D;D�R���-��5-���c���P+�!#_X�ɸ*�)Q5�9c��4�uS����d$k�8���T`�ʢf@��HQ�],]�h9��(a���}ڲvr�S=��O_irq�*�2{: �(:����M���@MO�I��,:�׵a��.l��C,s�T��XGa�c.�n��P��Q;o��.�rڹ���'K���9��'2.���"�X�h���v�}B�/j��=c�ʲͩ5V����](f݋-����]��X��w�@�PW�& �f��ټ��,�X���[���H�BA���(�v�<�qg�/%�"P��N"{��Y#[�ۧ���њ ���o�W������є�A5i��⩽ϕy�҉�b996KYcD��5�7�[����D��$�+/�^�[�Ut��e��2��O�Wmi�����������Y	H����`U��hD��纬�����/��2"F���MY�Y	�m����19�cA+�k�ĂQY�C�Q�
���}�/
�o)0C���޿69��f(������A6Cy�	����r/��+6�s[xf2��"ҷ�4tہ�D�(K��؛=_�Y�d؋���Ά�y�cWM����FC�#��	���*��3���|��=9jc��?r�f]d�^u�����}�>!��Z��(�Ah���NMOU[p�����m$\?P�>Us��s�}r|�	�^4{����$�z�'s�Le�do����w���d>�"v?��B�2}B/|�+g�����S0We�N2��b��L{m+�lv,�w��贙��䜾Yu��7nB�]��v�( 5k�y�>Π�p���4K7���_X��h́���S�J�&��~������;Mϐ�R���ki&m�����-;����RۈRֱ�7ovT��dp'`�y�vs���Z�l\7�L��G�����g&A�H����������Vr�2�٫7'.�w�L�6�xKX�re��F�z&"H�X�Xvʟ�ݪj)h%D6��c5H�77�'��Yѹ�e��G��"��p�~f]N섺e@�X�� >(R3�Vr^Ml
�XT~�;����u��qEF�w��yҼ4;�o�dAɞ��]q<)��(��:�3sٰA��O�UG�ku.fDHz�[�<�-�h\�`�9���	��W@�/�0orCmfmz?�9ufJR��m� f���K��� �c�3��M�����.���4f�c��ۀOkZ����"�!�:��:��E)�$�F=����pO
vx�c�u�X�;�}u����=T� �?^,(Cȗ���]]ڧ�D���W�՞6�L|�b<��aʧͲ�`��:���Z�bSz� �8�R��ɀv}A��\�J�ݡgI�Q̎�LO8OS�(�O�
HRT��~؊:I͈�o�O�D�7{�D`!S)�����o7��xs��6�=����F�"X��x���>��X�*��U��5>��_XE�L���y5%m��A*B���uY���x�|��J4!0��l��>��$����Xa����fvF���Ɣ��+��l�y4D���j6ܡ���8�a"�#�)���:_���oү!��q���]�a<2�t�U8�22�\K-��ǎ1 ���P�iL{���\�I�1uX��y�v-J�yK�06+�Cp7b�t�He(�6��+(MM�$��@)+Rtm�|F&�t���D�$�y�*O���%�/���n�4X�9Jp��Xeƞ,^(ى)�׆g�?�\��8^�����9�� �9��b�d�?]u,�~��/ahWE)�/�����Oպ�����kl�#5���C��H�@Ru�Z.U+y���%f��`��p�"F��9)����uƺ`����ʹHnN��<K"�~����q׋�����8�� z���N�"[��:B��W���2'�.�@?ɖ��% �56G�V��^�WGv���35�q�4{Z� �%����H����������>�������
�i.���.BL�W��"f�
`&2]���݅��^�����+L�U���FV���ƟAu;��	����޴��[%�5��9oN��GAeڮ��'/���
'�p�tS�9��Nv�k���?�� fۆ��%w'�����WT�ؽbY3�,Y���72��{��g�eB?B�l�#>aO�K
@��"8��d`�{��< x3�v;�@%��3�b�x�r;-��Gϡ'YC�r�җ��Hi8�[l>���ngݩK�I�kn'��fk@�ۇ7�wMG\�)��y�5����:�Tb�ehGz,Iv�LUw����{��gL=�g�n��+�rZ*	Un�"έ���B�#���Z��*#)��2�*���z�j�A����x�ϋ\�硨E����P���	FݱF�$q�-�<�Tl7� Ήlj�D�����n�����;���۲oi��p��F6~���1$��:G��mN��ho� {�ݪu�A�#�!q��RFY�,I{� 8�x8���c�s�x �	Gi7�2�G_Wu��ſ���R+}N���s(dF�*�ҥ������c�@�ln�Ɨ ,�Ń"DFnJ����g^g	(��#`9����"�W-L}_�] ��P>�x�lb��:e�7�?�AG�9����ׂ�0��8u vj|�}�gn�Й<������F�JFq�q��m����
��V�y2�M�v�F칬�[�~:���w��M������?x�b]R1��yMW��' 46��j��E��+x�R���ͳEP�-~´��h:,�;���MΥ�`�y�2SH�cG��sNx��懪�(Q��8q6�u>�߿��:�n�gu�J��%�]3�1V�-hW�y�S��Z��"��M�l�N�bo���i/�D�(���� �$`m5�,�����q\:��6D��k���H����/�s.�DF��g�[w��������W���Yeq؈�%y�l�60n�XS�Oo���֒�6ۧ-]3֖c[�C{�>�����M�N*�~���	���E��1��YԮj�E��e�qI�f�V́�?��y�.+0� ����d�tw>)���A=���A:�p��١�sWzZ���8�#\���.���|M
2��8kC9�:�	��a�栫4(*y��b�P���a�V������C8o�5/�r���ė��h��s=����Sb�p�fn1����,�l�.�2��H�t�B��(:l=��޼�}v	[��O��C��X��M�|���1G��W��������	Y�u	3��D!�H(]�S�bn�㘷��~M�O��@������ެf��aaT�	�]�kxZX��s>)H��V5�q�|��+�`��D�1X�l��`�c8,�t�G���W0�̣E��ق� �U����Ln��b��zPC;��@p�a��=���b�����v��'#)
:q�L��!�_�Z����)۳��&f$[K���A��R�T��p"[hG��^e!G(������ayE��*�{].�V��N��m�L���*��g����1]r|��"��T �
Ў��;vb����'���^�e˘���#�c}/�����f���1\eP�\D�Xx)h��{
-]!�X�O>ӊb�Y/h�1��eP�p����of���;�9�P��=Y�-(���7?a��3�#�C6b.�P�!\y�(�H����g�+ټ�DRqs�q<��}�MV��;�bU�t��{�,Gů� p�ȿ�ox�
���'.�n��lΠ�LL'�R�q�L��6���0�a�/z[ ��(�Ù�ϾTq����i்V@��������ڸ�ϯD+b)?�}x��m�̭���>��n���sB�z+K�k�2]�W�����#"�佧��D�I��C�z�շy�BI�Qŋ�7��S���'���<٧��'��*t���1]�D�F���U!p�9Ɉ\Ź��K=�O�
�"���
8�\cVZ�a��
����I�p����#;��v2���͠v�o�NZ�>��L�f��0x�	�R�-��0���/g8r�^�1���d-p:Ju4����Z�*,���ĭ����N�?FF54��!#�&�ߡ�i�ZG����i������������@�Cr��8�	�3/� ���W=eZ�y��B�E�J�k�D傒����k+.v*/����:�s��w�4ù�^�"��*�J�b�e���l/8��}#���r8�#��@�E밨+�[�[:?R�pw9DR�Z��@:_r�[bowZ�����4��{��s��J�ͱNi����*A���N��X��NlTԗi�♪�x��"�Q��`鵓g�Q��Z��ҭ]M]c�}#�!�0I���	Ƹc�k�sђD��ݭٟoM�`�+��w��R3Od�=D�ݘ�hj�Gլ(emFBv@��(v���u��M�$6h~w`�F����=�V�87��fŚ����Fb�X܋�[/�a!���z��P�V/�Q\d0�4c�$�g��dy�aA&'c�qQ����&x�(fx�(I�����xxj�5��=-�hzZ��Ȑ���?whv#�9��\.9��d`U0���@ܐ�����y���ٕ5��#PX��<�Ԙ��:5���2���V�4�4?Jqb[�$5��2K+EC���/\��;q�~w���{��j�?O=��\����&M��;/�=$�Wr���X|Jqjj� ��9-򝢙��)*������E�����f�$)
�k��Z�8DU/��P��#V�x|��kA�����6�|[->#h�ު�L׊�i�OA���E�/v�T�g�<}�S^ 8v!�ydtɲͷ�r#O�ˊ����R7��������P���L���iV����،�nY'���.��)!��c��+�6�/G�ɣ5��{���b.��*_u�A�X��U����(O9��(
rt�b�	9Gm2O,���J^�� ��+К��?�N�z*o�,J�@�?�Ʊ���;h~i��^�K�B�/����K�+�ՄL,�^i:�F�-16�-�\#�����mnz���T�0
e��_��E�CQ�
�&��&�j���	Nb{|�9o\C��lK"˝r��|�3 u�u:��쁾�'kHƁt����Z�!3몟�ρÏ�V%�����Ɓ���V�g	�b�̍���>b�"`g�S�j,#��2�-��1]�ׄ��v{�׬}���❱��K
y��[	�heS(�3��ò��Yŉ�?T�����b푛l��/��x�r���zifbM�j���C3S�>����>�?��۩ԢD��:Z�\*��ٷ�	Yv<���<ч_VR��_�X�08��=؜fM�%4��=W�*I�M�hT�?T�u[���<�c�o�����VR��:������Bb�<�@��{]�+�F�i-熘�6�_!AH�V�VY���t��W'���R�1d<| �{��v�8&�zۯ�6�qC�~����"�/�烃Z�	�{����l-OP��A_1�мg�"`�S�Zs]�Q����9��v��e�[$5�4X�0C�	�ZhVa���jm`�	
Y�C�Z�L��7��.G�a*�R�d��`t����0��@���I=.6K�����2X�	�$��!�#�MU����,��Q�mA�`�[@��r&*A�˱ �K����o�����+�1�$Di4,�[�(�M���3��Q-��5l̀��r�մ�DW*�'n���_5Ã=ydaJ ڶ������
�R���2�Q��;hn|+7G�����{�qv�I+��e�i֜O�p=�:΍�"$�|go�U��Z*P[���8UƇ2Y�נd%��gŝ�D�/�t�S=�^մ��8�	�_�C(6������dk$������Y.����o?�M�1���o{5���_2H�5Η:����޵b|t�觉����������3���D��Ij?�kz���-�B�Q�`���,��.i��Sh�)�4��	�FfZ�P� �L��?����ל����!x��'T7�7��?#�gC���T]�~w�8>������Qt�!�87-%!�y�A�[]�pۺ�A�q��h�r$j�t��j$��B���%���,v�gk��h���% 0̓��>"�_Wx�N��fl�����S��5�$!���1
0)R*�����Y�N[�'��5j˯�|��;ңp���e����;�3���E�1L��ɨ[���5tb�,Q��?�f�V�WU���y%��``&}0���0���}�a��Z�˟��o8����Wɴy�g�c��tPM����W�L���!�.'p�h%�+J�q�G�v�
���>w��U�2��c+�~�����2a���G�R��I�L��i������/����8���%�(��ӼsCK�b��Fȓi������7$��ǘ���9Uxp\2�#o�?ߖ�D;%[��ԚD�����;:c �`���Zy*�i9��%��I0A+I���J��Mh��ֆ��<J`���Ӑ����6�<��m�<E�Т���ӕ��;�]��yu	������_��RE��Aj|tƑɅJi^���p����n�	:��a�`�Z���`U�aƂoj�%�u�T�*3�1�,C�����\.(��S#C�����n�E��zuQzcDVX�l��C�@��i~Ų���*���&�(&�Y719��(�ktfP��i��̈́��[����7Ӡ ד���A��@W�l����y�9�*��k����}u�o����d�����N �F^�_.�a�p�> %-��s}�z�U儯�� ������pU���MT1m�a��W�	��D�N�3�N�{�h�Ev�����9N���1ס�r�{^��B��a�֛'���7eT��iq`:��#�Ld�E
��_Y��W�Q�����@=U�p~N�V��㞖��z�-��0��,0�z�2~m���Ut��"�;p��.^2�qo��͢YP_!������ 㢗sy��T��c��0*�T �:FRo���=�P�T��A�t��k�F�2����~>�o�_����s�E�=T.�L���J�z��W�[r��e��.�e�!W����g) �rK�F�~$�$��
^{G>�Z�-�Fu�ŭ�a�6��l+ڳ]��o&�
L���M�;��������d�>��P�����f{�Y�ƩQU���-<������Q:Pu��u]�+N~�Z	vKX��f#kR=�>������QƤdT_<��S��|����4�⌎�Da��\��8>I����Jv��-W�351MUw��-
��m�OgO0�I�"��J����{ΜJ�g�1��Z3޹�!�)�s��V0L�/�$�B/���렎@o����aאB�׃Gk��߷������~�9�3}=m��H��┨�B���)0��HY6�°I� ��g��~�C���
1IR��i���(��LFK�~�Q-�E��X�f�F��w�t����G���{��$e��$�Z�N$��'��M�q�pmh�&��'�×��'�q�ۼ��pi���:��Je�?�F+������@p���U�,���^�k�]h�tϵ�L��]�~����JO�Y������O�φ	�e�'��
N�$r�ڠ��6�= �(p�_�L~��W(�&�օh�q�p�|���U�ARprC��W��b�'��~��̪�3D��qX�����5u��TÞ���}�5����YɝKg�%��n�%��/�Fk-G6�!��S���7���w�1�6�c�z���^�k�46w@�����ɴ���Y�aS6in|�"��T�̴���*�I���8�6�� T��^�����b3x>G)v�-Db�A��<��D��B/��J�h�N�=�h���&��,�+�L��sc
��V��~[$��c�H����9i�7΋u����٠�`�~T���r���?����ϴF�@՚dV�U�S��1v���V!DA���M�l���^��'���\�A-��9�̞�:}�.��w�h�bױ���3*��.�-#ڧ9<To8���G ��^+x�^�?���z�����[��:����VpHڎ�F��%;8�!�ا�Se�a9�t5K������gX��e��:���,��������8Eo�����ri�����߻�]M��]���C�~�MߢS�B,�Z?�9�Z�����:1�$�v�_p�,^���3Y��7�5�ByVi㱣P+q�\)��S;Yw碲��8���q���=$��|ֽ/�$�e��:��˳���/!D��s����1����5����RpB&Y\ �����Ñ�3�s*��4�,,� ��4,�h��4<E�2?�T{B\Ż��7���Q���.b!�[˰@���!61�3/Ȧ��pgĹ�R�bD�m�ȹ]��~�:����ǽ蟝�0ז&O~QJ��a>m�d��R�`b���30Yő�8��4��m>�帤c�j�T5I����-���n!� ��%��ιe�V� �v����i26����e̋ܗX��d���3����qC^CT��I�� ��^�Fֈp�ѫ��)"����~������s<t[(�C'�����<!����~/���uGք���һX�i�S_R��C�{�.U�n�Ow�sISIƛ�dm�讂�pI�_YO��d3v ����Y/>�uRX�Ve�	mVF��.+�Gi�}T�m[lՄ��*��H�}�P���q9R*::>�W�I��%V�v��Lt8�����pLj��v9�<o��n�@��{�G��j�bF/_�}`lr�����1E���?�gX�S��6�oL�J�#��`E�W�O�Y��l�価GL�������S35�B��S9��d
�Rc�݉�wO�ek��@��BE��c/�E)���y�Z�gB���f�ǌ�ԥ5��w!?3�}\�N���c�h���]a-� +��
 b>��2A�
�7&�=TS!�}?ߤ.��I��5MI��M�j0��b�V���ȠH���0ͧ��a� ?�d�TM. �����G��aR�*h��Y�?Rt��{�#�_��W�O!�.J��F���I	������\q=P���'��E\�5��Zߙ�Yi0۬@��Ri;$�F#`.%��d.p����E��}��X���<��͙��%Rc��0�s�u�t ���1�,��?1}�	�G��E@� ��Zz��>~�І͋�G˗�?�9�e��&�A�t�
�݊i��O/���q+¹���쿡௵/V�W�ZW"��6� �3���A�;X�����Qlx�8��aSY����'�հ��ۭX#�g�D���$0��0/o,F�kc�N<Y�{�JB���&���'���A�Q�#�܆� 2�
�P��)�kY���w�VԪ���qocC�5����C&��!@
S��ʪ��҂�t~Z�X.y
��-j2��;�q
�H��:�5�B��R�Wu�za�G��0(^̂K�EY-U��3���P�̔F��n#tI�GܣVUZ��8H����C�_��l��s�z{r�M��£��b�3%nr#Q%4SL\���G6^�:{�	�:��꧞���Kx!��M� � G�hl��tP'Iq�`�c
�u��������K�WIxX���X�B�S�� �l��W�S��O"~�[ㄜ�C�
�g�������sN�b^>�����C5�4-tx�3���9�u���u�Za�뗐� >؄�
I�H���# 2z��}Yc�{�D]}����W�e�lIi�	��x�P�w'"��1���9�@:Y�*�q$�:Ɲy��w
�S��e�ԑ���R-_e_Q?ӞSބ����Z>Q����E�b����.��a0AQ�%����l�56����bpS�,�u��au0�uW��������ǖő2-�>Ȅb��� ��/������i��槥3Cr"�v�(��~k c�8+��
���8���X=���&�$�U-�1�h�ƽǶ:*\%)hc�i�*kA
e��
�X`in?SpZ+����=�V3����d^o����}�5�U:K�0�}�ܿ�Vy�,X_y��b1�s�K1�v�`�x��vA~_v�B���s���3ߏ�R�e!V�l��Ƌ��/�sNF�j�6���HLnC}$���( ��ά��0��>]�L����<%���w��1J �r���e��dld�*��w�]X^p�+#�+<�Y3Hz�Qoc�}���Ӛ�]x���,{|0��?3U�P�[<��'�
S,2JO�ǃ�1~���a�r���;��7k3�����a=��a7��D�=�q����O�b�(R�ڨ�F��*��b��=�5g6�Ć�iEē�L���]YT��˓ׇ:J-,� Z/���w�Ibo���׫'�����^�(�@�i"�&��y5t�+��;��_1����zf-�ޮ��̢W{$xʈ ��B�)�ޟ�L雾�I�_d�1�\�%^�c��T������kj�m����b�W�X�TgLrrb���<
�,C�M_}�43=�2Α,����+�x��Fd��p���e%�|1�  �O�b����`v:$އ�K�*���la��:�o�g;�q�.����$�Iyu�Z��_Kq*Czl_���3�%��t�7b0-A�AY��&'Q�N뙔n	��IzjW3��9��K�[ܯ���0c5beҞ��]5�@��9콊��A�7���J�􍒎u�_Bk�� ��y�H�R<��=P;::Cx �����=����W��8�����X�����ﮟg�(����цH� ��\�������΅ǪR�