��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�w�\պ}���'d��qx�Ba=��1�@t�loa���u*3������~��
R�:\�K,�ǉ."�"˞\Gr����[p*��%Z0*�)1�S��Idt�r�'q�)t�#U/N��{ZA��/�-�tTc�z���lf�XdT�cS8�1��<��[Y�b_�`��A��8Z�_K�g��6�F&A]z,6�>�_�P�_����1���IA�dJ���Ē	�����O	5���f�%�͊o�lR:�$�`���G� � ��6cC��T�2n�S�OJD�r��J�L�OA�<Qdc�{�'u �}<�q���' *|��C0�Del�l�a��Kxh�*�&D�Թ�x@��������s�^��X�kp��|���K�6�4�d�`�+8��3�!}f���7iR��X�l�^k #�Yd|Q�8��`�̻y�Op�\$���4H�|E��qJk_�a8�S�PQ!n»54'��)Kj�sej���𨐣E�%�.�s����~�ܗAƺ�B�P[K�d�{Un]5�԰�>R������qA���I�ǧ��um��.���ߠ�y㉽�W?��$�O �����C4�y��l�OIY��(��2�c��QrH,��ߵ9b'%J�����/��&�@[�N�`5�5	9��)+�~��;�.^���CC�#Oe~gz�?[.[O��/\ٓK�>"���e=��Q lT;ƭ��i������r�;]wG� rdjN(MZbq�3�'HH*��Q�� 7P� .�w�T
�&;���
�'�OpH�n�g6�b�	�{���,�'�|ꡞ2�y���vԕH�_~�6�,jªU����c�D�o6��8曋�7~u�٣���c��Lh3�����r����6�z4�|㌰>�Od�������,>P���x����С�f4=s&+��L�� ���}h�.��,9�s�(�3�lY��{W�H��G�cn|��&p�)?��Z��U�]*�7y+}Z�o��~�P���-`��"+�Gt,c%1��n��i��{���0;j�a���U(��k�8ll�������@?#��� ��hI��]~������bf_��}��w��w�-oRH'��r����32 \�J���$ ����Ʉ�{�^4����>��a�{=��g�0r	^��c>[ɛc~r�{������m:����y�M�'mW���A׭Xk4�Op�1�Wb�X�@�%��+VA�n���Ҧ�M�>V.T���{�h�7�����,�-�Ga���B�0�������]���}Od�m����Wl�S8����	�����*�ֵ2,����7���>=R����h��8�7��'A1��pސZ�K	b`���<i<�n�L��0� ZܓQ�/ߜ�;�DCl!��$t�9��i�`g%�پx�ڐ~��J�m1��8�F�����V$�����͡gT��ǚ��P��6��Mk��٢�Ĩ|�ɷDu� �H��y'N�:$���ie�LI>$	vB�*~����>WûD�n
�:�n�5}0��w�S �6Hy)u[��p^��i���U�H����]Q�ORWO<�_'YJ�#z�@=�v�rH��R�v�k�"Q�&Ѡ�PM�^�=hG�й3�y�02�ƭ��c���d�ȓ����L55�ÕF��lG�x��$_�JV��L�����ﳽyn4FJɐɌ�6/�lW'2������b]'OT����Z�?"�m�k�	��Y�}��Qw�!�pH��5�~j@"�!v�&=���ȿ��'�q��riM"s-n�����B�������<"&�D�V���9�t��mUI�3d2���K\�o���mi��� ���-%��uE����A���BU*�"2���m �co��ĪT���1V�EX��o��>�E�W�k^a�d�5���1q?(y�Hlubl��oo������U)����%\85�ٳJ�M0:.ax	"?�LJ=/n�ΝH��'���c}A�T�!IJn���;<V�<