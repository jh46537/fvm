��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�z吴�)b���ΡrϷ���	�J�`,��1B��k7׳�k_�f>��d�O�Tx���q��t�Xb���[����>�ͣd�Q��-�W�pvK}$�#/�У��(��z��r�e��iD4m�x�1�:vLS���
��f���.�=2��ܨ���l�w�mŠ�.�u-��"��� ��9Gk�C��u��Ɉ����z��#���R��0�?ԫ�=�u���6)~AǝfӼ����w��`�DU��C�Ǽ^G� 5rX�R�k����fC���X$�̳������\fޏ���`�;��1�2F�D�/
&Q3����p��@#�O�ARf����&u[�%GT�b7����m�ٛg|��![�,Ȼ
L:�埖|g�30�~u'�@+�N��l��;����.��v#��μh���Q!���F]�e��+���ր��	�n�"��i����֤���n[�|��F�̶,=%�	��Ee݁8�G�!��Ԑ�C~:�59�������<��gf>oĩu��"L�@�8y����d���w&�+ݛ�}&:�8�����첫Ǘ�nz�5	.9M�[�F�5�4[V����������[�ԎGv�bj	��If���3�_PZ�(�S25�`��І)Q��l2�,Fs����<� 9O��s&~�=�f�`(��dFB������a�Y���,�,�!4��Md�2�!GI��}W"���p6&�AD�R��ៀ^��[	@��<<����+��Tc�m�u�YQU�%�t�<g�2�& �~���Y���a&	�]h����D�6���TJ/��mB=U�3�u��ٱ�q��v⯡n#L���E��~��I���ɐ/���HBL�	i��l�ګ���WOL)}`����+ƛin�(�#'&��v4��T�Y�:@��Y�;a�vC��nM�U�Z$�$D΄�����R���V�=�J�I�	�槲:0k���p��HPG���i!�u�mXt�'�/�t;�*C���@1P�X��?d����1@.��Z.*f|2X�Q��ֆ�%�I������8+�U}�5��݂8��r٧����M�^����o�V��K��'N��RCx��ׁs�zW��9jj�k��]��_M��a]����;�W0�kNp�/����2�R?)C_0&2/�B ��ղ��HU���,2�8�<d7�g��H��41ф&��Qb�0e�>ۗF�=�8;�����Oz[]�&5�U� ^
�
����s^�j��c�a��K*U���0���`����Lr�L*�+	���P͍��#�BUGo�*�Cu�Şj����2`����.x�V�{o�5��q!g,:�y�?ZQ �QGX���k-�z���x�do��)�=<.ڎ��&�t���{��^UTZYdh�>0$�T��]�s���M��[��w���>�*��o~/Llw��N�fU�⛯���_ۆa��]p)���;�e?.>�'�!<'�V#�٨��Zzr�kC�2���K���g�
�����<��p���SA,htr����$��r��d];�$����f��~�q���P'��np��� �����!�ղL�#H�ub�#x�-��ڶiw��O.]�wֽr6�V;�D�Ί���6c(ʣ� �*�S�T�����)� �*�ZJ
<���e������c��]�A�c�ߋ,
2%:c��U�T]ڼ?/T	������l�5�½�>�L�R����8����T�"��Q�p�a������N�	$D�={$q���OR�����eM�~�Э!�]�8#û=y���fA��98�(�$��'���X ���@f�3;џZ�hjAMYw^�w�|N���_	m���KN�����"�.�?}�SdP0xDUճ�4�Qiq��ð��0��|�-��:|<:졣=c�e/�j9D9[	�9���F�)��R�c�n�,���iՕ�
t��8�������l�o+�'M�b<<u�S5|�Hq؟��M�G�LV_g\᜜��h�s�4�B��1�r_ǘ�p�r{K\���嫪��|�3w�`xu��u�sP^"��<Z����lN��=����S�ŀ;.myB�EK4*��z	{�V`��f�8�M�8r�ݴ�2]��'}D�Q��Cc�y��7%���P��X�t���?'B����3O�e��$\�'���i�Qmh�VPRUl��=��b~7A��4G��x� T ��#�dʿ����zoJ���~P*��l�iB~��,�h�Ѱ����>u�Z�@�hx��6�cS��[�	���hn�M������*��L�	7��l����Z�bF�p|'��o�����ʓ��q#���۵�"���^]�9�=�2=͇4�����gF�ݨd'(��1`���[�!��I�@�l���%�,�A�}.�/I�=��y^�*,T_\hۣŎ[�N(���N�B�� :PVc�-�/S����E��r���.�7��%�V�o��v[�*��>h� ]NW.>��U�����(����q������ª�n�w�o�~��T�v0(��&j'��_��x(rG��B�
�&c�m|����nʗ�Y�|<U��r�<���k���[�\Ӫ�>˸��	�_�%w�w{������(��-�@�X%���)�A�p����Wg@�#�s�k�4�lM�"�7�i�a~㠉RE���du^=�	E��`O�#�����z@��5�`�A��ޚ�&���.��R2�C�`�~4d�)��z"��֍$�ѫ��z*F� �p8�'R2��}g�����q�O����3Oy��s)DY�d�󲤾�U%���hB�� ��^�������l�r�n۸5�������`Y�I�CbQpW�D	��T��+�/D:<�ج&
�	����RY�Za����u�I=egg$��P�"�f�"�B��Î!#��P�
)�!c#�&.������$v�� (*�<Ϲβ�[>$����e����fI�
� ��p�RW�}J�B�Q��C�{bE~[I�;/f�M�Ŧl��/��A�{�B�����h7�6t	2V�9�=�.��7�AdC���	�Q=
�a�\���{6��۔]�k��%3�65���ig'�_K���(���t�毬p6Ix�gG�b ���a�+�5�#8��e�@F�*�q�;B>�(R����{�'?��q���IDG��]��ab�h��ͥ��]ب4�p�����ryw���������)׬m623&��GI���<sCA��+j�Y��y����H���~�h@���.����t�T%���m���{X��1�	lҫHl3�#�&�bpk���#Y�#��a�v(�FE \6�	p<Az4�<�h}u�2��~����L� {�����+r������"i�Ʊ��L�"ԍZ�
A���[؍1g3������Zi�{�#����ɣo�%�m���hR��z��v쬏]�l��_T��~����?���X�-R޿	IE/��;�;�2�ܞ����7ı|�0)b���k��/��W�DL�i)փΨ>�����,���M1��,QlE"�v�)��Ouu�dy5+�l�9o9Ⓜ�J۞u��~w��H��	AcP����ކ9dHį>UNH�ʐ$���� P ҭ�p*A�/g��� ��0�J��J	��A�x|&�Pd;<�r�=��۳^�]ʢ�����sS���!!��e�!�E��X�����3xj��绁��1����YlV����Y��=�e�.��U���jOMJ��gO"���}0�(2�X���IZa��tb�%�/~�hM�f�,M���А��$�#rs.@����_ Χ��p�s+�XG-@��~���{z���:��:텝ɤ�7��|���f���+�9��(n�vb�(ml[�����P�G��{�{���IW7�(0��@2�9ty
���L�`��P����pu\u��hp&X �K�1�����<CӬ'/>���x� ;���{��G���`���BC��W��֟�O�Q��Gc��.�H�^ą���?H�xSt̝M_�y%Ȓ�H�&��ԟqQ$��Ir5����M��檴�X�v��B٪����A8�ZTU�"�D�޴�cV�ƻ��0�XSiҕ�H�Q���Yn���g�ڭ��o���� ,t<{�N'@�^�
����-錘׭�ͻ���Ǵx�}Gْ��8�#*Zp�ǝ��� `��'�/��",�9~J>���c4��g�d��kK]�Í��/Y3�m&��"��
k�{����Go�܂�|����C)6��@�&漸�+�{�
��v���Oq^���?b�t�V�b��8���9h�/�������<��Axo�\�rt�QRg��f��v4�!��9:9��l;�"*�#���$ �@��4���6��';<2�>:*ɩ&$�aaoJWo�։9�?U�Y�I�F��f�eC�J��g���[��)һU���0۳�����;�������͑���dm��\>�*�f�\8�/�:� ��k����*�T6j��Yq�̳���k�R�����g��U�!�M�b^��)O1%����[t*<�eՉdbhG�]�OP���@KQ����.��+���c�)#m"�׊��,6+�4�"+�?��0+�{�MgL/# �'zK��������?��	��f��t�t�[.&0w���K_��D��)f��B�������2�b��\��F{*g�+w�Y��s�:�M*��.��a�+�=��[�		����@�P��0e\?��� -�����.���,/|p%�<��t �IVq|X'�u��N�-Ӝ$y�gqv����Mľ��9D�+ƴp����r���QZ�Ȏ��P��S��gI���=Nbvc�����sU�O�7댬1����d�F8��gV9#�Ґ��9�=��_��L�7K����MW�e��r��w˶XC��[F�ۚ���z?¦y��+ܢ���kά��E�BD���@"��􌳃>����>r����l��uH����~M�ōΖ8�&5�7`�E������x�3��ɟ��`ȺH�>�1�S�������-g$l�[3FG��W��htM.������p�Y��R�x�鵝����;�"<��|6�BCN�^�7n��S���^�f'd1w���dR���΀�|6�#�A��=�� D<�����\��/�����B�oS�r[]Ca������t�Ѱ�H��9e�O����q�����~���4�= @��0�y���0*�?\�S����>�**��/Z\����eY��)B���d�_q[q�C�G���ji����r��w�B��lf*�J	g�b>ѿ�="�*��뛎=i(5�v4|`��է:����'�:{@��E�j-`<��^�������3���{�T�c�ˁ����R#���f�Y��Y�p}Aqg�lr���9�$Q��Y?˳�~�'���\m��ۥ;��lS����V��5f`N_lyÌ��!����Ls2���\���\��N�^�����D[��e94	hV���i�[�7b�7T�~]�6��]�:�/����%�0���#�����̈́�����n�a���}��r
!#��P�K~Gg�&�j��Slc�n;:U�5�f����I�9C�����ngy�\�l2��	��	�Z��V��L?����}�����녊��E�H�#��Hx�� ��p���g�ɋ��A]g�1���;m`De�bԒ՘��g�������(�9a;�E���Mܜ��j���, �+u�'|h �%Z�>�:�Y��1�S627(��q�����4�%�+���)�N]� F~�+�W�v83U�g��<�KYx�S�JN}^���c�3$��������[�JEN���l5GI���F���n2?I��c��2'j2I�^3��6m)1��^��8��{�e���,8D8�]wdL��� W��(宐��R�v�!&R�O�r�5[�E9�qD7��W]�"3�JV�F�'6[� �����Ζ5E�95�	0�|u���c`3��J�_��nH�x�+�4���9��U���"x�i<n� �u>���D��i�<�eK��&�J�,&��,a�U����U;܃7Z�SH��� �L�I�"O<���n���"w�����<Z{�&#��N��r�~I��I\�1#-�+Aϴ�f��<8��3�5��Ϫ��"�.�>�MB�x�U`HA�A��?��t-r���@�_�`K7zDD$�G�7A�DD���O�ᵠbRT��̇�'N2�
�H�~e�&�-�.���Aw��v�lC�P)�ڌ�}��z!��l���u���T
�X�w]cI��D��t�T-K`�?�,���M*�>p���V�!�) &�g�@ɣS@KQ�|akO_V[���v�L��-��,��4O�7wcfks`��B��g]� }��3�m>`����
���K����������S�RP���ˣ4ӽ��"_�tB�WRK�]���d��I��=�� w���<M�K����<ri�`3�
y��H�E`'˹3�/M+��9�}���1@Ű��R�=��|Q2UEw�)�X�?��uQ�'�)�ijYHNӂ�D��Y	��yww̍J��5>�{���v��@�(��m�dƁrHH*�����k���[��9y����:�����/]��WO����58~'3��M�7���f�b�D����� )ɪ�Td�B��|�c�eX[�f�C4 �<�y�Ձi dߧ�4�e��0��
&�_�&�K<�9�$�	�!aal/��W+#=J��蠞��K!Ɋ�wť�Qq��"=Uf�'[�bȡ*�ͅ�h��'������BMMS�8��[F��A.d�dAƍw��3��i��lEr�M��{�9|3j�k�3|L���m��� ]�q�t=9������C/:����%���$����$/�>�X�%���3��N���;��T�l|�d�����Tyv�u���'��|5 }�!���G[>Br_���n#Y�9ZL�������Ճ���2�C����P~,�u�������?7L����P\�pK���ƃ���`�Ը0K���]�ǻ�"�e$�z�Iy���Kح*����"�y7\�@�����3���DA2�{@� rq3H�t���M��^���\����{2����\%�����$"E���e*�A��,�����]|�_���a��^������Z��m���XW�WhR-�C�������Zᔤ�$~������\�ϙ\s"b��8�5n���ߕ|(��4ɾ��:��Q��Z���1�u�$dن\C)Z��.��
鮺h����J�k� Id�d@b�H�*������l�C3F��\��{=&!|��*�zDL�����UI�\�˸�O�@�0��	@��c�+��
ڷ���F�ٵ���}&O�7�WJ�l��Q2�J���T$�e�u����2���\>r���U?i�+�ٓ+�*4[���1��}ߟ@�
T'�#�>�\�賱�8���Fo2�dn�EQ���Vt	}l)���no�"�K�~��� �h��=���~�f��2*,�L��0���a��`Z���=�ie����d&s�w���l�>����+��f�-u�0=2
^Ib�ޖJ�H�n�nW	2���߁r����:����!j	(��R]9�cl�/|���ѩru:���ֆ��!�o(��dX햧FZj���c��7�5A���J����R�1ɇ�Vj�@������٨��yᘌ̋dXPp��_��*B��@V9�rX��n�m��Rr�~��m��N��7�?�ϴ��p>0~���NC���Lg!��˄� d��JT��^=���x��R�A]�Sz�0|�C��́8oz܈Wf�e�lw��� �hyo/��Xq��>�zixMͰoP�\b/��IVC��%'K��6'����Gvmb7D�3�۾�uXL�gےJF�DQ�M����xy�칔0A��y�/�)�,��3�Y\Ƴ8	u�-����H�#L�ޛ�c��J��J.��>����Q؊X�������+�õ�u�+g1c�i}q��H���Hj#N�(�Q��\X�{��$.��b��UY�Y�6p	Ш�UX!�I�s:��jry˒�Yd��/ў]���рT���s�GP�Fj��A=���hL�1ƬƋErZL�
��$��G�b���\~�dt1��;��c����z968��x�7�|%6/�����ij� 9V}3V��Tu����A��`��:(��` �QK;X�C�Ǳe�6#BV���u�E1�*-���bӚיT��汫L���T����@��:�r�,Rm�//��F{���`�v�讼X�����l�{?F���HhO�������p�����z�U����k���@9�\)�G��4Cw	M����V=F�kXeT�
��g2�?�1����/�Y��>wUZӂ�ԇ�8��IշI$��Ɵ`�iB#�����L��̬���6+� �h;�=w �>�l�����{�ᾀ1��*����'$�]�� Py���Gf��a�Tv�x��K� G#|�:V;��M.rc��z�\ߍ!b�)g�
g�����I%��� �F�#S|�HGvk��x�&��ҸO	��>.�� ����f������'�B3O��3UY���ט�M[��7��|�^)�PO!��7���l�`3&~�W`hg�n�G������O�3e��ml�6t���0�\z�%�\��h��ѻ�~.=��mI�iȪ]���c�A����)�.�*�ȦGo�1���UD�j�2����1�����!P�{ �TYu�3;S��F��X�O1)l<ݕ��eY����t1��Z��$[�-ч�O�\SA���=�^E���	����;���	�(�Lh̗�l�!���� \(T��^��(���2$�>�����^��� �*|ܿ	G�jF��i���:��zr�"=mT4iۍ������eh"$ (/]S�Nۦ�j�[�Tr'Ό��:O4���<5�y^#�G���l���PT����� ����D��MA��,��3\�z���Cp$¦�2��7��uS��)0VG]���څ�����˿�}D:�A}��K�inV��$#w��hM1��]�O3-�S/)���~�f�n��H���'3�钽���V������n�^�؍dP��Ֆ�l�3�]:Ґv��3B~��Rs%�����<���!��e�j�_�J
�V��6t6���<l��R*��H�� TA"N06�ܮX�䞛���^�$����C!���A�5��c;OU�8�I�!�$<��Te�bDfZ}�@7��
�	w�8�B��J��A�:�� R�Wa*3��
#�|���"o�ﹹ�s�#���|�﷎�_D���z /����C S#��CE���[�b�~��8Cߞ9�=�#�?GB��LË�d�yE��Fs���|[�n^J�	9�7���7]�w�PL�rp��b�*�(N��=�c��?<4�hJ�!Y�������/|�U�ݣ_f2�(�Z'|�;:_5���Y��e��sr�⫛j�Ѭ ���hV%�/�`Mzە�~��	���J�Ă�L..�îc�i�'�;��˪��}�;��1�ˇť0wJƟ��#���� =A��������h���_��s��bb�m��ŉ�ϰ���VqhS��o�'��O��"��ic��jɮ�R��1�7$L��ۼ��H��uÚ/F�}q��y��:�S��H��B�����Jp��Ijh�u�;{ơ �P����X���,'�dg�^�H�N��,�7�^5.�n�P}1��a׌�+ʐ�1�.f*M~������^�j9&C�ԾS�(��M�9�y�ǄQ2� TKJa�� �IH�Yв9	�e�7�/OI�3��#��W3�BB2fD��nu�)Y{��:����+a��	����X���&{d��ݽ�@ⳇp3�4�]�E��Bi���|
;`��5U�g=f̩�y��RHM7��D,�n�2����}�jF������x�� ��C&"ن�E�㾗m�=I�%���.��(�-����i�,��g�WeoR�43m��`�j���-]�?gpd�~�V��0��H�,*�E�Q��þ?V-���LZV�g��y�l�U^xg:��,Ox���9,SД�+�d���Z��
9CV�E��]��͇�P�`f�f�M�� �(2"����|ֿX�����]}�w��hx�D�#A(�w�� ��j�9Mpحx���5v����3�i��D��0褦͕��	;��'��&��܌0,0�)h��/�6Jy��>�һ��d�����+A�q V�6��b��1]�dШ� ��$X��e��m���H8WY�����Ɔ�#�2�t춘���[����_E'm��������|�)PH�A7���6��|>|)H����%��8n;`���b�R�!���� /勂ul�9f˷�@{c3����C?*���~ʟ���X�W4?L#���:�X�:��S�4�\2�<� �Z4P���Y]���� ��2]y�]拿���6���<�l��L`�:-�l�v���gÖ"a��81���^�?�=kc��[�,�=�>�
�_�d���(b6���8NZ-8��J�\\�����HiG Vn��L۵�T�����dA@��*Y�{G��m��
�o9!�،��D�9�<N�@m�L��*���V�pl���TI�����L�z|�Z�2��p�nm���[E�/���:;���h3�(��T�|E"@�Sw��IBv|��c���\������A�=lUޝ��-�0�#�Cp�O�:#�hoݳ4�ƾݻ8j*� ���:���{����|&��O��F��r�o@ل�S_�sI�	]�2������0{��|��U�,�8�
ot�S�d���+�=D��Kq1]����9��KͶ�A����V�G�
�Ks�@�l7:T���bҕ�Y���Q�#'��"��[��Z+̅!�( |����
��m�[ޢ>�S�&	970b�1N�p��V+eFAu��؞Y��_�>I<�<��;���=ڸ�hEXI`M����/0~�h�<]<s�YRL_�\�|{�P5�ؒw��%�R$���| /�I#-�9����h'��l�_�)W�g