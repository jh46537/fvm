��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�P���|��S?�6�B��k�K��F%5�@��o��5�������� ���@���E^������ ��65�k�T���S>MG�=��g���I�G��]�[��=Y��.�\��`��?Ր��Cפv�Q;��]�%�;/�v:��Q�'@���_�78�?�UJ�?��1ŧJ����[�g9o�0����
��|tz�<%���W$L��l6��cf.l,��Y�`�Z�Y�>�h�׀���w���L�"e���}%��J)T����{]Z� �X� ��z���Od�>2E4���Q��J���8l$���	�F�sk��e�H�c���CܤD����I��W*G��[~Z�ŧʋF
�8�P�����X���b�c��
}J�*�S��7�M�n��o�UyRJ�f��QE���_<�8Tq��2���W"�F0e�<�E��<ZZ@�-��B�??��$*�gپ��e�:�¸�A������Q�;[�x�'�VTQ��Z5��ǀ�)]28��S\fŵ!	8�E��+r�qv(\2?Z~�^�i#i_yk����k��8�P��fُ��aJ%o�L����C��lĎ(|���e�[��X�ulͮQ�/-�"Jo�҃&�U��U�v��ҪϿQ��s����̌�V�f�~�l,�8�i
��mՒ�R��R�Zvd��@� �����q�'εN�L?�nkz��de��������G8�O4�)�R�B�4�Q�@��PIa��pl�6ޕY��o�y㿏�ѥY	h%�_�����@*ixDMx#� � '�4�%:��TF-��'��z$�� YUɘ�Lo��#�-�gL�L��$:��'���^�|A�}e[�P�H*cO�5r3x������ ��ʜ����7�~�&R�gU�\A��s?�"���>\B@��Ć<�Z-�c�BiPN}��M���8�xk���@�Jh+i;��j�iG��+�j����Cr�og��qDqץ*��k˘�������vu}���ݭ��f8�iv���%�L7���������'���$ދF+��(,�FQ��y� ��0Q;���6��3+~j�><
�r8+%��<��gg�v���p�"R��*j�����3yJm��9স�IX>G�qo�eI-��n�-���L��>6>ή�u�J��f����hr�9DE����Uz�
�)ҧ��%>���wq���u/L ���gE�yh�ib�{�Ռ����L�-w���S�i�fq���­�@���0>�=
��۹b�n�5�l��ـ��'�H�kF��!���v�t6������/���Ne�(JH��H���1K���M��=�fFK�'�tp`�t�q�ѥ�䠷bZ��
`hvC�����P��z��g$��$�d�Zݵe �;����C�=�##VL����mx�-�?�r�-�,0�c�n1?�n�(��2�����|�"�S��򚨌V�!d���� ^C6ME�� }�����N;Y6� �<�j��ȧ��(�,��d\|�Y�VQ�ś;����g�$a�Տ%¤]�"j�RW�Zx�d.5wse�F�;����.��~����T���6${!#�J�(De�)]|��'n{�3�z�Fw>����&���r���)�>��U6Φ���D�G�R$	W�j����fkY��Fwp�|��ʝ�J��_Ftw�4��A�&���}��q>�a�P�W\��A��(�E�SS�,��#>a�@Q� �Y ����5N)�����]����v"�Ύݲ�+���tk^k���1Lj�0ΰÖ�E}�J~0��6�ǀDG�z���b�,�p�X8Q�u�����6Z r�����/T+��9]�+�w0�t�M|�+\
O���^����z�&�
��j*����35��U߼x�;��zJ}�{��h���U����"�9�y��=� #<`��n/��=^Q�|��&�ĝL�U
/?��\e�\v���L�Pw��F�G�7`_ҡx����?)�?�M}s� �ڟ\�i����L .^�@���(�:~Zb��T�f���+k�!��,a�s�G��[o���z�Qn�e�8�������B�	��N�iiN*���3c�����(��w�;���������7�՜��m�u�6�ژ�k���¢~��:�_������֪���=w^��h�(��|����~�(�b��
�6������L<�qL����t+M��5s �j&g�eP�1���J��y�i�q���_�N��l�ѨeM���~��Fpm<9���,��Q0�#w��O�wc_B���1J��q
���W�ЃK��R�xb�G��ل�V6��"��{�����/kudV͏���^�����ړ���gD�eo&�{�:K>���+� �rv˲ea�>����a� �񹴈`�G�a�":������ ��h�����V8�R� U�%����"zb�nl^�*7|8�7^�q2���!17�q�F�|ݠ�FLww������Xb�v|>�sc�W�X�����W��R�`��	�z�=	W�z�d1U������%���u��`�=�D�! `���v#h�:ǆ�s.�,�9FbE��:Q�Y���b"�s�N���øw��!+���"z*.���Jvo˗�F;�(��o��F"oB�8�G^�a�hyҶ�ۊ���#gf��*�
؅��