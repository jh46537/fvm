��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���Ox���0��?T�}�D�yBl98�锛�l	`�ġ	d}�:��PƸ����~��R��o�K�jV�,R����vy���3����O���Z�����g�̼A��v�{�7
��5�¾����B�C����������r}�:ش)qqa���·����BW�4����"V�CL�zhXo�e��6kT]xl(���%lT'�W���'�N�V#�L�`�`�Xy�6$���:��9I��ì=P��uS�I�w��������F��<��s��y�i�u�����ml�G")�O�4����}�,r��𯴢}�鑪 _@�y�Tkt}��8!�JŜ�>9��C �gl���-����{���Z�*� 9�[�B���c�M�͠�+�G�Yy"TGz_'l��2/;��	^F�/	b2�ܕ�Z���./k7iǶ�>��R nS�}O�i|�y�����V�����2(D_��x�c��h�`e����;��%P|�N�k˻	2�{B��-��|��̧ے+�o�.��Ɩ�O|�ٻc�-�b�{�a�-'����]1.�+!�jJz�l��^fJ��.��r�~V�`���%��̡+b%J_g1ۢj</R$���ϚU���f09��^��|:%ZZ���sT�+¬��8#�[���)P�ت{��R�P�en�܀�	p3;����ǐ[��Cs�~�y��c���*Ѱơ��[#�Ӣ6�vQ�)�q�#��ҹr�3��;p��N�}����4�hpOx 	h^̱�ŭ����E�ǩn���!�؀:��*�f$dg��?�ZOҔ�%( ί}$��ػ�m��S��5'.SY0x4/b��y��#?�t����rd}�&۱Ͽc�q��a&�C6~l��Q�ab$��"Z�m�?�y�A!Ou��l>���r,R-��f�(��!>v�=*��~�E��)lQ��O�AQ����վ㪭��Xsc��H
����ۺ>&0+,k��sY��ޙ�?%���a./lv����NOR��� ���g~��O�ʤ&i,�FZ\�3�j�:?���ft2&0o���H��w�N�A^"��Bp�?�MW����Y=/U�/g�E��aO`�B��Ԛ���8�q�.��p������9|;�>�d��z"a���q(wY�x:)��B�a�2I �b����a�,a�4{��J�N,@CJ�@�NJG��8�?��ƫq�p���\��i��h�W��L�~�l����(x�]����r8�լ��A�p���-XY�ty��&Dv�m׺���l둝߅�o����ɂ(­��F5�p�a;P���@�I��y��'>M�HU�W��m�X��d#�d�r�}�fZ!�Ǿ�stŧ_^k�@w�]o���S�p��w�z!}�Ⰶx�\��q45�������O����5f���2������O��1��q�SX���E+3�f��v��+��	�������m�����٥K��H���Ht�Z�0o��2��՟�#]W����~��\�vT8�b*N�Zy���>��~�j�q&�ͫ�]Uk�i~�����y�Ed��s�Q����,u{�^���[FO�ߠ��D�#>��Ͽ�P;5�UMt/�����z6h��vi����Ҷ��Y5MZA�x�d���\=n�p	��	�6F�/��lo	�-S3�u�pE���*�BAK��+ۦ��%���0cj�����h��<H@��UK/ً )�k`����Z,ɸ�3�hw�O��K�����lg%,ce�+c�p��cz2�y4c����{�����]���3g�
ʇ ��i�8[��H����������_�9N���>M]�f����8���|6LC���9�d&p�r�!B���1�u�e��S�S	|�ik�l��Ɉ�m��<�$R�v\lN�P����FY2��׭�k�O�%k�)p��`���b��-��	����1\�I�U��a�ڈ�Ȅ3�۫��%Qd��τ���b�s�����8N��e}��+Hs�(3����Ā��FT|FzL��H�r��Hu\�,jN��tq����:@���dI��5���������ؒ���=��Y1Eŭ4���e��ЋW��T؞��Cd��4��p�	����W�~4����ԗQ(받��+�k�j/eg��Z���5y�b���G��F�r|�o M=[1^��U�����rd�ۆ4�b��ͫ��Zb�ki������hM"�y֔OD��y��ZΜN�� ��O�Fb�%L^�4��mW��p9x�||�m9Ĕ�#jd���*���y�;�n�M�ZΦm`wԔ��C`���j��Ո۪'����
Z�<C��tU��)�N�w���Era
Q�֬|(�	�����{��"����CT���S~Z�* �!2Ŝ1�E9Na�!��  ��֋��-��a���x!�8�z��/{W��Y�V)qh�20�G���s}��y0�͒d+�k���scI��N)�4��ہ�&�^��j����\�.q�Rͬ*lb�0 ��*�����v �-\�D����$���cZA?�ڲ�*�՝N�PJ�޻���٫���N�)���R؄�[C S۷����V�mnu bæ|T�ƪ�����`�����pd��q3k�+�����~������j�vmp'j��9��҇x�ԯ��{֜z����q��C�]�|t����������.~��~H�����$��_Zj�4�ׁ�d�,�ٹ:����E��K���ЄAQS��� j,T_q��)Z]�H�5��9QZd�pP��ʤ6��ɴRX���l�@�!�U�BJ�Mx���ݻ�I�����
�p���͂'""4���4koYW�6�"΀�Du[��dܰ��W�w�>�
?
��>X/:4hX���`l�;�Iv��@��se�pҵ����(�4��5S�G�O~H|��k@`��x��PV��ڂ�L3t�5�Tq9�W�mJ�$�����~�_���O,�����,��Of_�w~��8̎_lꛧ�K���L��M�3h���5�Fa2���O="@e�_O춺0�q��M��iVm�J��JT�z�/��An�u�'疐f�e��P-��1���K�
�̒������G�a�E�T*9�2�ar@��J���K�Fz��;�O�� �Q��EZz���d��C$,D�6��7/ve��ƙUW�w\m�����X��Ozrn���B�ھ�"�݈!�^: ��}��&X��0�`qx7����GUceWl���-N�^��WG���5��FW��"��վ�]��Dv��t3�7�R���K���\
.��2��P���m�Zrl͋�T��+�w�������v}4� ���8 �Zqc��P*ɀ/�[aa�׹�u��E����	���Ss��_�qB�b�&F��S��v���Af������$W\�vy���곺�Mn#�u�,�Qt�m��Kw�$t�yg�N�g�63�#CB��7Td78�p��y
�/N���O�=�)2�`��z+Ap,��*�>���g>��'�Љ���N���9�w%z�y�CӱHԫ�_�ͼ��H�"%.���=�Ϭ�����C�Sp�-F�i�i�b)B�Z�*1L���H��!ˇFK8�1����M��	�Q�2�h�s�v^l��#�����V�E�:�|�=d%D��f�����qv���pV�y����F���P��aC
tMHYF`j4�'OK��� A�mD}k��r��9ru?T�eK	���aS�:0�F����	@�������Nx�|�D�T�^�Gv7��`�)��`��0t��+��^�T�lf9�����G�YR��	�oO��5�5*�-�oÇ�v9��*�\�9�j�=�N8�x���:�p`s�M��q+����d�����%d���k�h	�c�v+���f[��"�1.�~o(�g��W-"F�
jP�G�dEo3�w����1���}:���J��\kg�Sg|��A�����=�Vyқ����9o�h\��f%�^6��ҍ>�:f�,�K:�U�}��5�7'��h�#v�T�VyQh~Z�8Ïy��]����[�a�F��)i9�5���IYU �r����)U;FnB�o�p��o�l�˟�Di[��Y&��,����7�=S���
U���.zDԖ^�l��=`��~�I\hm���f��-O��S��J�G�|+���)�ɱ-B�b��5ڵi�0JX��7�	W��̆d�x�a�!����UPU�\��*��"0s<��}�@���xHN������b����m]�9�R֒�4�):~}���P)�I��H8��a�^�3xH�)��S��� �u)S+mȠ�.*���iA��d�ܱ��f�]|l����w���[���g�V��cXX-vj��YK�ol5��᫊�=�	ç�CD�M�4 S�s$A�
H.$��'�J���'�%Wj0j�RL?��c�<��Lw�ڂ�u7[�������n��9)����X�Ed󝷒�z:���5�2��N�ԫ�B����9IZ��
k�<t���,D^w/�8�g6�xg�L���6t�9�@��=�X	�RJv~��&'I�-Lo��cm3��ۮ���ߊQ�n���<>