��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI���!qp�6ht����B;dv
�[�܈
�/���t�!HO;���;��.$?�'�-#ܨ��q�X `*Ƈ'�e,��Sg�Bno~����1���V�0HA�=/�c�����)7!/2�����&��������N��Қ	Z�G�i؈�7ХP��^��S�T���4a��I����Zp^�B���,��1�W�؂���K�U��=k{�LcF���)��Idᦿ�_�Jy�����d��iN"����#�,^F"��.P�P�����9���})��ւ}�?�T��;_O�@0�|&���7cgKD��PD��댜2�.��%`:N���n�@�8�ݘ55{�K�l��߆,��`QJ���ɘV��kF�B��+]�4E�`�8�`�-��a$�$$�.~T������n`-*k���_�il�
�J��j�E�@���tΰ�krݺa����K3S��l`�.����lP��>aa}����#p�T�����L����t�c+��1�^x �i<6�����j��08k���g]V�e��������eٵ�|����O�^�w��"[㍰dɜg������H��v�q<�vӎ��"n�����T+H�|T�VPR-H�69^��������]�t7`�a	�^�a�;Cs����6"v�]��Y1����W�BOO�5� ��_3��g=J+1)�U-���BVP~�ƥ��^�2�}nt���*w�G8��I� ]^�|��N`Űxn]��1s��=%~ W�r���DS�=E��5B%e�ʠ�YX�|�7��	ѕ�a��ͺ�O ˅{��" �/���:���Ž�6�Ga����$�=R4q"!S�p���C��|`!���� ���
B�����wS����$Ȝ�����l�q�z������l�n�A;r+tJ��Qz9\�u����d�OR^1fx�Qv$Ѻ���hQҔ/����$��� �Ӽc�}R�lԺI��ۭd4�)��k�I��?�V�G��J��X�9���R���1jZ�!�C`G;��¸���m_���LLꀵ]Qw�B���[H~q�˦�|��a�D��+R��?)�q1���7���TG=�a���cT31�Ai����A\��!)�Vy�~lD���^����
���Iy�b��)]��O�ף���y&
�'3�"�F3�^��������F�X�b�kz�/EG�ʪ�Q��λ �k���z=�@��Z���. Ѱ��+==�\N��Х�r$��/"TГ��V  �\X(� 1��s���y!�-=Z����φw�r�ٙ�����W���5���>�ׄ�عbG�B���}�g���9��n?I�Y��u��o�.��J�L���ہ �C���2�'�>��Fa�<0�����6$m��UT�aM-��'B�@Ď,�z���~��')xA��@�,�X�M����q=f�����T<=��L4���R����C�]T�i����l_O�tO_̷'A��pr���N��o�*��hs����xҡ�Z��W�$t�8]����Wx��@Z;�H�c��2��Gf�O�� 
,*9S��K���1�e��9�<?����>�vÜ��qW�mA`��G�������5�&i5�	��.g~��䎐A��$�3!Z��X�>v��_T�~��L���"�-T�o{�R^�}l��-1�2�7D����*��ڽ���n�$ץ���ٞ�ov0r�ԂO����W���.�l%ۣ�W�1>��1��+���z6���Pn^_Jx�	ڨ��"�ظ$�j\LC�Fw �D�=�N�K�<N�֗�1��$?E�{�~�~*�OX�௟��#�T𯫗 � ���׀Y�К����2^��C��A�7ն����_%�kI�V{�H�!#�f(��>JNa��Q�#&�~1��l����~����X�T�$��q+�{g6���o��2 ����� ���70�����N��߁m;���3�0ȝJ��� -������.{�{�V�q���ÿ�(�7 �!�\���1%?���
a���(�W)5�L�o�Q��%~�Q�?��R����-���b�i���JkN��mk;X�DB���h�z��(	H]��~M?��-Eh��^��ʕ�q�i�������O�B��9������Թ3����-���(<��� �/1�ɲP'���;���K���˸�	�F������j��dԨ]����p;�K'�qW�E��aa�x����Ė)�kŝKV�g�M0}����^��󻡸������f�$W�o�,��L\�ZE�����^�#~3G�vl��G��T&��n�^M�����Y�ک	hN�]X���֙��!�/���^�XD���e�<��`�1�\�Kn1�* ���3�}vT1�Ύ#��J>�N��>��