��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0����>�P@�:��N���F�����"X��7Þ,���S`3��Z6M'�n�������8O�����>���3�75��Q�%���ZtT���Ow/����'�vJ�S�dt�2�,�`���q����l�!�S@a+!q�q��U����0 ���6�c���9p�Ë�5��A6�����m)J�eY4A"��cW���ŉf9�X�g����E�|g��֦l]�΢�Y��."��7L��#��#f��]e$���� f����P����
#��q��7�f$�7:aZMFV���Nm�b+��B���1�?�-&Кx����8�\[�Lu��hʸ��f�����+��S�+FG����wۛ�t�OfGw��׶�X/��6�B��>�o�+�Q�N+.C<[9���fv�㏜Z���h�;G�BQ��)�Б�O�{�xx�1�E4�� ���u�l.�EI���l`�՜�o�r�¬�M�U���%k#��,`�� u��e�l����3��2o��k�\[G?��w'�@�xF�n����%��[���� ��)4"/��sx=~f�2�M/?�����kݷ�ԃ��s[#�����91�PēR���0�� ���uB��p�Pmd��r7p�n���i��c�>�/Ͼb������v,�w� r��㋅V�Br�K)ipU�F�z�h����W>�����`��B�|��&���Sʽ��Ϳ9o2BP�5�!Ѣ	t��b����x}�  ��d����%J��\?&}�Ŷ}%��#� �	J���.��|�3fO �w�٬�X.#W���\O��z)�E&ܝƢ���q�c��|�s��}zT�zu���6(�=�to}������3F� z9��1\Zu��DQ\�Cz�c���Y˘&�$Y�U{q� ���/�����|[K`�;��'��;�2)s�|�$�����=�7�*.�~��TЌ�luEGɅ�=����w�Z��լ��W�ҫ(U�v̩
���<��=G|�H�A�K� �E��1�<� *r��<��E������
6�����mTOv��g]`��q����+��8�;@>�l�/Z�|��-
���A�zf1�yP��V�5��P�)�0�5T����u�@��VC��פ	�Q�=j���|�����o-X�@m}(޸���"!�]�jD�CX�
Ev�n��Y�{�@����ez�$.
%U�Vo�Cc��㺱������^��7�lm����K��ک���<{3:�C�Z���Pb7v������:	d�in]�3�t9���9z�%^a����ӌs�Ӡ�:cn[|�@O�5!wh) m
�@�YQ��i����;ynp���>5Ll�2rCu����G؟l��b�`��/�b�'n@��hHw������Ҵ]fg(�
>��*"/������`���^-�����	1v9�'��\7�l� �V=��c�����u����+ku�yr�%��tވ8���U�F�U�?��"����wg>�bAH��cv��Z�<���W�d ��tf� ���iP�Y\���Y��C���& x��Vǖއ�����(��w���	����Y���{ܚf���{���wU"���0��[�h6+*����&�n�DR�8K��#v��l!Wo�F@�:(8'Z;,ۿ�~����w�옹NS&�-l���+��#������x���6�-a'+�گ���q���hG�m�J�F4��Gd����1�oM	���L�uG�G�m��~�*�T�e,@�٘i#�"c�ӝD$�礭��h����"����_���i����h�!)#1�?]��{R`��_=P蔧q`�^*n�t.Z�
��_�se�o/h��z9"_�x��,#�n ���܋Є��C{�>�Zv�f�5Wc�pt_03�7F�_�V��#�[݂��L&kFk7�*��g�)'W7�?Y��Ѝ��-
��}�z $�S�[#4EB>�))�6������Tc�a�KE�@���L�i���~�?��E�aD �5�.0�G�+����|-�.�`��f����꘩��i���w����m����`���9�0��}��5��r�v=@wB҈	�2=�j�,<M�B(��Z���W���Q�. ̅�[h����Z��Em�F���j5/���4*���