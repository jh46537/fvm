��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��!N;�?'ǝ�{9�1�\��,�L�B�8��V�R?��[6F+�+�4"p���n�d�#�$؍p�����.�{¯q��ěW�F^��A�S*��|��Ea)��sz�$��O�+�d(�W�n{�|��C�:� O��U荈PjZ�h�'#��}�Z7��-?D����͈#�26���1�o%3}V�9M5@�����s���F��	+�5�������S�/	��;;�~��g��JRyyҩ�M�'������Q����4�1_A�<�����E�s������?�I8��6U�3[����[we'C	�De��m�!L�����;ܜ0��V�~Ջ�r|��˛a�1X�=��
�M<3��(&�<�<���U�p�b��)��+1��+�����=�	�"Eβ�,�������pR�Ry�+f߮2j�۞o

�,>��������wX��2�:D�J ��� ��<���h�S[��h��-(��(�s0�9��5�[t��s�Lm�����S����f�fQ
���3��?�$7I��Vٚq*�T���8�!yxɕ"��f���&���4Y�v����^�re��F��������]���g��D���?��EH���2SM�>ZT�Ӷ����k��ֻ,��9p��3��XoS���,������vtD�S�Z0#���:0��8��Bk��{����7��e�ecQ�6~�|��/��8������y�dgO��4Y���S�`�_�� �8|C����6 �N�.���]�S=W�h��5_ @�WC8��#����d���.'4����'5C�'�Qw�V�m!DP۸2O��Gv��fr˖~l�2���^+��,H9j���@��W�r���,����+���,|��֘����ǢH;�H�xV��q5�nR�<��îɊ���
��r��P��5V�%�R��4{N5�1w�A�*�lO>��㉲��
� �|�w����k�w�'u��G�|�p�e��x��~�'=2Ҫ�y��<��2�!J?�q�؟ +��_K�2A�}���UM��w�-�w���R����R��g����p�aV?.�V�Y���Z�"�h�������3R{?��D}Jik� ��$��ĳ<!���>5�\�?b�䐴��,���pB�L��W/�q� �\d{��#�s��c(�����+7���.��9��d�w���d�6�;�H��{A��hɟ0���||x0��L���O��8?q�B�����9��1�!���`q�tQ�w��"��h�;v��"hb���ȫЋ�{��c+�z��Tt�zzͰ(��Վ������S'N�Z�آ&r���$���kP[���Nlr�[��]
���f��:6��a�.y`ܳ��!n�����3�d?� 5)̀��ŕ9�&o�$�r+�+� �SE�N
�'-��hG]R���#�2��Ŋ����Qh�����fl���s4���nd, �FM,%��*�)žHە`'�/9H�0�H��1��+��N3)�I�KT�e�s�	�䙼�S_���T8GGf����L��lqz4�J��G�r9��/iU��%)C���W����l���7�x�n1K���²�5�k
�a��V�]DT�e�0*KV2e�Wn���3OV�"p$���f1F_��g�Aיr�#ɝ��oOd�;,�l�G��=�kD䟝X���7�������(��Q�Z� A�q�sݶ�9 �4>��\mҽol�����׍r�Q*�Y9�o�KUa� @$�r�}��"\R?b׭ݿ����.��E���%��ܦD�)=sڜ��~�?Y&���tN�r��
��9�0���@��
X,���"��+�x�g|���M�\�͕��Ww�gzҿDA	g�Y����]a�S�,�B��B�sJ
g�� ��W>�b�n����jb�K�*����6[�]��DL
L��zFq[�^՞2m$��W�P�����'iWe��ߑ0��h��gIt�4q�l�����ٲ�;'2�Q��y�C��)N�0)�>�&���U;������p/�l٦˚��.ѹ����w&��ƌ������e���ۣ��<Z&ό��5/�W�H�ɣ|	��qK�����������p�T�	��C#��P�m���F�(�(�a��2�n�z��NJ0�Q��֨�d���ym�
�^Ŏ���-#n�5j�Y"���p֪ag��Q+rv	�d����P��R�A�Cap�N�9:V�?����bV����]�&�q4|
	K��w|�6zXl!ͦ��Y�kr�����H��9Ÿ�_Q{hB2-�;��u���>>��BJY�M�_��V�G�4����p1.�t(=���%��v��[:1��QF�'H!�_-~�������X�-v��|���*IO���RY�G�QM����Sқ�·`���ڧ����t�A���[�z�6ƿn�+J,,�3��ջoJ�Z=�v����n���/I1�#�w������.ܕ��:�	=H�o/���4�CYQ�z�M*_ ��>�ݹ�ר�21��W���u�}��p�E�d3����2��őL̷��~�!��	p�`9/ؓ�M������Q�J����