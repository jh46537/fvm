��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(|����	t!�εE�0,�
��k0���K^	�Ӵ�:֯d���e!֥Pl���څ����x~��ٷ��D���:ݻ �7݃Y+m�*/�r��U-E͋���6r��	RC��P^�۞�,��Oo�`u��]Ƭ���ӵYɦbEW�,���d ��C|<��!"Y �Ϋ���n-K��O0��7N��21x|`B'v+����>m1R�벽A�7a���'\|���RIz4�	bS�F�j����*9���oWj�������2H�Z�o>|*�U�7�A*�:�ӑ� ��q%�թ-g}Ǫ�E'g��TL���M��P�ߩ��ΒW���4^��??>$x��1�td܋*��������(R�!V��hAy�Mܙ�k
*55C��	��k�Jm�Εj��2W/.8�t�a�r��1n.�!�i��7RB�Rg��^{&�MA���j�8���+�Nv��
\���Z�]
�Ԝ��6���\5�ڽ�P�+�γV��=��i=��wB:�-�pw=��m<��Q;�M�fp�4>I�׮�$��/�p��:� )�^�T� �'e4��B��ZO>�%:���S�����1�bg�lb}5QD���htȰ,	��8�:t��n���p<X���)����B�î.���o�b�H�yΞؙs	l��n�:�g��.�b�����҄R�MN�~'f#!��V}����O�X!5����oF�
�Y����Q%���bꑍ�,&I��4u��!�䷳)��e�ys�T�v�X<��=NV2�~+�>��:H"}��1Z�h�E���2�i��b���WDc#2����䇾5������ݫ2Y���Beɇ�\]�Z�r
si����׻��r�E_-R�z��5y3�esa��� !A��5����� qk�Y�e-�V�u�lu˦�y���?Cc�J4�$6��1�̍�:���c	�g��чT%���2����Za��I8%E
,=R�X�X5�/��W���}+�4�[�6S�0A���aӴ�9�J�SQ��ql7u�=ͤ��)�t�j ����q^-LQ��h�c��VX���[�P�Z��F�N{��;�"�D߶��U�x�e�l��jm����/��@NGmG�u�x�w�Mb�AjkA��kN,�E]k
�j;������Ȓ����s7�����zq�D�����1��(Ė褅�WK�,�Ș7cͣġ�CNdۀ�����z�_�o��r�-����Ҡ�]����3������2ǟn���O��+y��"�u�\��^ݥCYV��;�À&��#�	4�U\��`�i���|���?↢k4�_��U�cB/�x�Q���0L��e7.C���k9�oM���!�{dNҡaq�`t�>����4����O {��&�]�vG�ɟ�'�1�-ѤP���m�G�-Tht��OH�Q>x���&2ŷ��Ƞ�
w�M�'�.P��XN�nG�{]�m��SC�1���K�V��t�i5�ӕR���K�j҅�yʥ�`����sS-M
i�u7����$�N}�Ch{Q���\ɷ��e{�i>�+�hϨ�C?2�Ѐ���ݩ�z�A$綎��r�	ʏiT�Yz��{b��6w���E���'݀��jTA�J��7U�@�Q\]Iψ���8f��r-��_���-VF������J��/�� �QS����7IK�x�s`�`g]VM5Y� ����UK�D�.�������D�SYl�K�Zɋ�^�Fl`;��.���Y�C��b�@�ij;����*T����4�K�K�L�z�W���H���9TVk����Ey
?,|��h��G�t._�{@I�oP�7��wp�������������)	?lg��/nl������f�*0Kd?x�~��p-f�@�b�����ᢔ	dG,�����g��m���!���u��O���R���\��p��0�>�a�e��htL��o,�@�':Nt�+{M�:�`[?E[��h"�'�����%�+�d��΃O�3o��	���ew�g����?X�)��SW>�Jb�����e�T��fUѢ?g���T����ר���!X�e\�u�Q[���4��nUL��Q�=ᫌ�v8%��~
b� ���������o�x��5��f�h�w��?� �ou�ݘ�Θ�@5J��M���O�Q<�z=�F� ��Y�~x��
�U����#�>�(K�����(�` L�j���\1�q	6��mj���˅�~�~�:�6b��n�_�����`�h.�j�i_Մ��u��Y0u:�;1Yi��8����D��lj��C�[��}�y[��窳��)Gr)h�ӟ�s0\���a�5�EJB�-_q��'��w;�U(�6�� �ƕ5�/����a�\ݒ�k`�E�	�	t��<�9�>e��]�+O������')ˤP�l.L���gP���1��+��JD�t��ᜇ���(}�5����K���Mw���Ɔ���}�"�����>�2|�0q�AY����4��gS6� �l��_�i+M�1�i�� X���qc���|_h�;����R:�'|��Ј"��h��&o�M�?�噶����0�1�ț
u��I�j���9�%�?�^Q�8����R��!�
���aEC�C�kN}�e���K�4(�&�I����� �}7�<��]7ԗ����A����Q��ۉlB<������c�S�HW��{1��ͯL�I6<�J��|~�S��v���UkM��nB��>�=q�|;���N �� 2�/�I�5h�)��g��˙��B���uIrҖ�>�+FZ;'&��L�v!�.����H��>��`oBCy�3��xH�e�s���I9*����<�!;��Y�M�#:�ef�V�/	����L��:�����
�@�����lW��
-N|�8�$�k�P��F�a�{���u�����/k]�Q��Ԇ�|q��i���y)a˥S]knH�wӁ_�=H�:F�٦�\r���qm �v
2%��s\��?S)��ƪ^|�(��z��5A�n����١w��!@��݌�c�P�4t�J��q������p,���*w7�E����:�us)�7�=R[Їj=� ��|rb� �������XΚ�Ar�c���߰!u���ޟ����x8�x~�sW"Q�����uXY�C�]��W�<HG"NOP� (���?@~���M�/��;��֚��OaMQ���Ga̭ѯ����$s��:Fy$��7*��-c}�o,�O�X_s�����f�&���*Qh�3��Q�\����N�]$���-��f��WϮ¾h�ǐ�+˲���s�rմ{V��~�vբ�CM���0n��K�����r�D�*��g�l�0O�L�iB��q�
��!�� ��T4���rB��
|��6A0GR�Ƕ�\ɜo��S���o�(�+ޫ�_�U̝���d��%хȣ���˛�0|���b�_V�SMs掵9�`�1�GQv��J��)'�a���l�8�+�"@R��-��u��\�W�m�A��<MZ�
��D˕,wa\��t���"�vd��b��E|Km���e�r-�Lvf"zW<e�F�K��ٹ�/�o���p����5&�ًR7��BZ�#��f�FOУ�<D��[�ߖ�N�Z����QLRU���e�W���"?b�-�	L��)"4� ��٦��xH�yV̾Ɋ��'�I2o�>�C���zC�%�KA�qz�������riH���m�0�T�Vh��^�v�2�ެ)v�k�I���9�D@Y�ߕ�S�b:;$�fz��3:�� �8ԖװS��m
��߰��l�n
�#�G��)0�)� <�ULSu00Ӥ�Hb:��.�yuڡb�cQ��'���jT�"IC��Ɩ^sR.�l��0�j9?�\��O��ou�����'��EQ��m	��0����K}�5�l{�Qɿ��G�mB��f��g���p' ��&���_sz��p�A��l� P�rR/L����݆��+��˺�zo���-</DT_&��G��l�d��ٸX�R/|�u�ZRd�1>�b���T-`?ܪ���M�T�z�\�ڒ�ih��-`����_Au�����B)aL�єS�Vgښ�w?��� �.�ER��C}���ߡ%i��g�� W��k_�S#6���y��v���v+��4^qF"*�s�WFޮ�@�F�t�-��}W4G0�fw�:��I��޹GLٕ�;�!
~�����8̙���낱X�1���$4��s�H%*.�@^u��mW���6�(@7 ���聀��tzE}�W��tg�������T1��D���P����=�3s�x��>��M��J�uj�|�ڪY@^���b�W׭Wƺ�d��{~�?^�"s�D�5�AITɘ�ޔ���J	����[fU"� ��̵�0���j=l�$'�� ��R��z����S�Qy���J&	����(k������a_�޴���&�Wk+r�gڧ��ZU^5 `�Cy����#ϒTZһ��
�� �u/�3�D��������F��Jł���l�[Jh��,b�#��(�a���Ct�j~	<��T�.
����0��^uX�JB��wJ���(䖸��8�I���F)F�.�y&Ma��:d�`Y�ð�]I�Q)����S�=Rk���G�X㇅�\�"�R �T|&�TO��PS��u���Ҵ7Ma�uՂő���#I�>#L:E�~i�ߡ��!&M\
���8�����"�6�\	$0�@�۔Owl5��M�x�O*�\��x��B7x�5���v��>�B��1�"dG�_p�j��K4Z�t���[� ��7�\O�dԺ�R���u����3E=����Q��r|�}��DDO9dM֏�l�W|U�nv�\�V���.t��]yꔜUs�]���Ͳ�%���#�J�Y??R�䋦�I������}G���i5 ���D�GM�C3�Tۨ�+Q�릀�-�V��;�P�/�/������2v��ƽ����r�H��
�����|��Q���!^ b��m0?֬���r-_��I[�Wo�O�>b��������^�ŗ�A�w�aܒ�q��A=�����k��U�PjvC_C��9o��g�+�NY%6�k"�'�<��������ν@�
{U�����ˀ��(��!�p"��?��"(ۛx���t�b�����~c���q��4��Y�?�ĉ1��R�%�휑<C��°d�k�/�Ό�q���t�YT"d�o�*�4�#��� x�\A�l�L�/�z�G� 7�}�jZ/>��]jV>Sk��g.6�-�V�2J�x�Cj��o��s�3;g��~̬Ħ���6T@G8��k�Y���Dyu��(s�0�F�#��@]OI^BX��{B�77Kp%�Lq���� ~L��t�j[�#�e�{�@����#�iW{�- ��z�χ-����zA 2av�+`˂k�j���l���ԆEUW�P�VS!��t�&�$�>��\���S_>c���lh�9��!��a�� ��nZN��Wq���5�P�*#j�h���ף���i:�G@e�fj��[9h�c1ۋ�)��[�� ��:a���!�>�� qEy���x}��Hm�sEeM�y�~ڮ� �n����U���z��|!*y�x��^c&��m�$���7��qd��O�H(�:�,�)�|Ү�k� ����%ݼN.��މj[��Bew&�݂6��ǏT�n��t���l��+�K���z0���旉 &��r�8�\�f�@݌@N% n!�W�k���(D�U����ͮB��Y�4��֨����y��,� ּW������S�"��f�7���YUE���yV��l9�KZ}7o�.��*4N����� ��]��4�.�L�8�+��7%�L�ff���E�m�<�-�5)�q�f�xl��4/�$ҊҠ�ө�CZ���Y�e_6��6��V�� �?_��[I���L�μ��5+�6��:,	��E�scs���t���Ã�a}���|��r���v�8�������sa��_� ��}8��tܸ�`� 0�>k�tX����Y{�^p8#w.������.��g;E����� n44����� �e�_�po��!�W�,:� q�ѱS:� �n�M-�l���ˉs��b��_n����iH�ޅ#l�)ʎi�ܬ�f̓�!aT�׋��aA^�xX�~ �X�z��k���-3��}L���(p��!��k�Jn����$Zߺ��������*�oi�� {eO;�p�y7�V�:�U+8�,��N�k�Z��+Y�V1�����4��T<ؘ��B�!��7#��<n�,�%��g��}�׿!���m��Z���4|g)q�@ޔR #�<B�=�k)<�7�?�F���d�\�"x�&�P�N΢:��5�	D@-����Z����m����MF��>�*�c�Xh�ك�̖���cZ��bc\dD��85�Y�Ϳ?����/ג�� �;Q셾�
бg�EG�or�/�,��/m�O���G%<x*�ǳ�BZ�����9�W�ä�����A����H�:D �8Jd ��+������s ������ר	��k1�t���2�	��
Bq \,�m���	�F���J[�i�z@Ƕ�) r�3��C��Ӗ�&�{��Y�2s5�;F�Mҥ�
�,*��B��!L�:���m��%҂,"u&�f�Ư���ՏAIt� Sh��C����A�x�l-O�І><�;.��g'�u��fυ��a�)����,k
)�$t7P}��#�nuF��%ȿI'{l�x����V����eB�?;1�ZF��k�PO��`�JE�_]�)� ����0�dϗ1>sLj�!><P�_V+X�TJ�����g�D�9������^�	��Zʀ5�i�D�#�*�d(=yB(�P!>.��	�K#���|K��ʛT����a��}�ݠ�A�?����Q�>�3k�(u>`��L�e���(Qrt ���%/���3#qʁ-�c��<g'�����X僥�|9�8#�6'�U�@u5��q9�j��~.a933�$ �gE4���v1ᦶ�����i)L;��a�_��1M���dQx��e�>^MR7�i���|�����!N.0$�	���8I{W��fl*r��)"��Q7,R���$����yt.]����(���
W�`�������_`��b�	ǽ0�|��QtK�]-��#�;�k��Gp�X�xPā�s�Ӟ/� �1I]�E�t"�8����Q�q�Aԛ����J���cK��5����.��rU̸9��a��^��ȑE�t�x�콠�:�͜JB�����m�:�y��τ�5Ws�"�5SY��~:�4ך���<�R(Z"��
�fA]�9uZ�M݃���?N�T���i��I�3j4Q>��#�X�����r�0�b����=>MkmwT��/C&���.j�Z>	�j�-w7��VmU�.�kn�� 7W���8P�<g�'F��U��4�������l!5�����~.��F�d��r'�7��X~⤠�G�=����WY-Ǣ�z9m��LT]���ᵤ���an�8}�|��ek�*���F8��#<;%�;iU^YG�}.V���`���@Uڐ��ʦ�1��Ms̭���pZ}D
$�~t#�-tf%�&�޲PD���Mf���G�vFlJ�����>Ө��1��+����Ksɡ���<�*Ѣo�mWRc�^���.-5f�����*H*v=R�Q�:�5�W��;��lU���I\�`����6	0\�`���,g�I� �*�f�i��Wo��󝿖��t)������6���	�CF�