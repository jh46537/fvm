��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O!) ���Y�Q΄�O��*Ȣy�dsuQ���`�Q}SA[�.���(��<
vɼ��;4���͋s1D[
�f�T�[��h�K�"HO�¤�TwƜ|�J�tR:����p�#��;������A&�K��HȮ�!!@<Ȍ��VV ��k��ko窿ae����ZS(�F�FO��2�;Z=��t�)W�{yo��r��(�K�StcN.�����s{P�8��AN�C�/��~Y����[#�z�bEB97�'���?�$'�����ِ��ǰ[�'�d�X�������%��`r��`���8D�]�At���w	V�򴴌���R����F8[4Nj7�-���ιFUEp�]c��$W��9P�|�Ԝ��L�?�9�8	^rA�Ƿ���.�He���n0�u�+}@I�2��P%p���-���6��f�8Џb̝h����喥e n/&ρ�1��ue��Fw�����s���Sܿq󀷀�	�~��ݒ�-i�Ȳ�G���S1	�g��<�ד��f�t0-I���:oۼQ gD1M隬it�;y����4_���TB�چ���thh�bL0���]q~�����4�Pw��Du,��8n�,�045��u�3`G��볮��"�W����`�hR�u��yI&n��xc���&����7���W>=���Ű��T��+�ς7
�73�ȥP#�lm��"8:�K4�j��c��<��d�eA����
���&c.�nP�	�hy�Q� ��l54ꓭ��ٶ���j'bz~�������,��������&l$� �+��D}�4j̢�0��)z���#ef �2)AuO�3�ۉ��p���s�l,��p�J\W?��sk\���k��}�a�.�.i]�q��W���o��9�����^+@���T�ӷ1m�$�X��<�j更�UGk�y��b��}���8uw�h�R�b"㕑I`}�0B���B��v��u0ۇ���A@��D����N�Zۊ5&] ����I��-�K���_å��HҚlL#��^�p�wo�O!�`'����^6y1^��m��7���s�5���"����BM�&+��#��_����'k.�A�$ʎ����ąI�4Nj�^��Ⱦ��4�e�zg�J �Ty�hL�%� 桐e�L��ɏ3�jyBh��ߕtͼA+�)Y-��Ż��/<� �q��e�k2���mPf8�^�!M�Z��a�q�t�V��݁�o��C�-�c��ո74�3y�Vč���0�?Nl�S��>�c4����Ӕ��a�D�<N�A��Q��gM〦�@�`���ͩPsl9�SJ�MHM�� R����Y�ɀ�B��2\N��P�F�?zh��\��㓪7��̝"���IR0`!iw6�
�w݊�X�ǜ���Z������@$MT�b�R�1~��֫�sT����Xҝ���H��6 ;�|�Xϗen)���F�f�`4�-�!C����K<��גq����tjc���$��}�����3<95U�tY�κq`�odL��q�<"Fw�"'�&��ˬ��<$^x����μA��@�#��k�Z����\�H)��3jFĐ��@�������'�a#������/�.i�%y�������67� �,��{ �u��?*AXy�}�)@}9 ��S�����07I���+h�,3|�%�,Zc�6a����	�
h´�x���j� w����E��0�Ƹ�ePͲ+�� �f�R(�֑�p/$��*p�Q7bw�8�-��s*����P��&��&�a�/{|¤nC�i�\*��Q�,�1/	/_�� L�i�S�)HE�F�E�q��	y�0��L��T���Ld���F�~�l��i�-ሺX�zNB^Xs��蝹�}�9�/`��S$-�1Z6pY�T�t*7�fO�5M<��u:W7�Ǌ7*r��M�5І3m���š7n�7�;_��y�����}Y���d����J�ľ��w&m�ҟ|^��-��F�"���\��K7�E����+{j_�k7��t����~C��`n򜔹*��z���[֘w���z����LD�ΩE�ȟws.�n�����ep���\�v<�� V�Ƶ�L$`!o�7�\z'Y#��76��3���Q����hG �0���O���X���s�F�gۚUP� 9y�L��4ұ�؍3�1��*��xb)9r�Ł����U 7zvB'Y�}ׄ�v��g#�@@8:rp��e�|AȵP4�x�R����b����D.k_�?�k��_��9�.��>/�HԼ�#���oj��m@qC����YΆ�T�aH���(�A��17Qg8@���������`KH�X-�@�= �`@8�������Sx�����Y�Lm��=gZ�:%R|��XGT���p�V��$#uQR�{~1(�@1��j��RbeDY�n�	A�Np4��<�P�K�[����r�\������1����7�ɔ�G�ݗ�L]�e��
[\� �}���N&�Xl�̗C�Ð��sgS��z��ͨ�t�4�v�9ᒾ��Ll�L�cЛ�[F,�ɜ��.T�z���ڿ�������UΙj�l%2w��T_�^B�����1�����)��E��������P�%�sN]�IϷ�����Rk���
�UH���4����h)U�ܷ9S��P�dC^��1�:?`aش#5z�	�����`~�Z�v���J<~��1�Xŉ��m�s��D���}�WuX�//(͎�d�t�X�J�7��a|FJq)SB��R��;�%�G+���/�R�:���{�y���Q-�g�\�}��c�ו�y<�{��l�F�`+���щV8��<�9Z-��(�Pp[r=�y�h�%콧�����