��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z�խbvwR�Q�0�]*e�z��Q�t�&��.�9��������e8��]v��ZɃf�˹�:�bG���%$�ud_T���_mm�"�D��C���z���1�O�w������q�g:�۸�����C&��9"�NQ�� ��T8�l����- S4��V��׷�B���O��uQ�XZ��q+���`͏�H�s3��+Y�eW��3�otz�3Q&��`��Zh_�E!J*��Cì��ծ��&A��ȯX����2K^p� u�9���ѱczp�-�愍vLL�RJ��C.t��X)ޯ LK4B����
�2��%
�S�v�B�v�x��*A*&|���mo}כpzu���?ٕ��B����Ü����1�l�:���l����5\��M�e�^ǜ��͔�ӳ�.���0�6<�m��^��.��H�	ڥ׷���<<�</��&�ɰ�6`���`�z^�I�������Tw�b\�R0=r�hGf䋊�T^��K>;��{�lRN�?��q����u	�r��`�8�$��Zz��KR(ॠ0ˣC���u�|�8-0t����}%}���q���=�����m��ua�o�CӞ�w`fۛ�n�ʟ^m`���j)Ni��ؚ��
՗	�z-Y9��^�?�س�0؁��5(^ ��߉φa%�=��/�Yx-�t��Knp��>�=���Q�n��9�
X�2os�v�6ǒ	'�����|��M�rH�٣��\�q\[i�q�"H�|�d^�Z�~d����l��g���L�7���3{��/Q��C�Z�ij�#��_��ً)MV0�eׁñ\�G|�8���j>���:r�$�1���m�c�'-���>j0�8����5�fH,�r��i��`�JM�)���E�W��[��,�jU�E`-��C,����qb�wc7?-�G����3Ӂ��8�<~'�,�8=���DFp	_Fj���x��E�
ڌ�4���٪�/F��>�|r0D�4I
�`-��s`6�B#��V�J�2��v�R���_iN�+�L���@�y�L����,�,Q�	���0v�zh��P�)�zܽY�%�g�V�v.�y/5�j xk�
k�W|�/kv��t:�jH�P���<�<[!o�P������T�abhO ����@D�S$�A�.��+d�����ҿ�\��b�t�`��)`���/����ⶬ�a<g� ���`���+�<���5�>Y�Gq��:���#����G��yʔ��>�|���[���;�X�hV���{�s:r�5Qf)d����t�17^kNJm<l�5l9�7�ʟL�-$7�md�'�7ٮ�R�n�/,�쏔��MZ�[�~2Y%3��퓖+��l��Y�+*��jQ����S~>g�56��y?�Ѽ;�i�ʢed7���[)������G��T��I��px�3# MF�_ց�&� �~^�)Q��¯2�,z�3gt@�{&S�ZdSs<�$��ǗX�X'j��h�':������bo��T*�rƂ�;pJ&�-2��g�k���[J�I�oXw7iD�s�z�G�5����Duf?�!s��;�&�:uS����o��:d���tc��k�_�f1i�k���[�׌0��B<w%�W�����g};�&R7�½R��o6�Tyj�M���A�. ��3B7n<������	Am��6����A�{4�+C�(�$t%vJ�E b�-�E��䩓�������	�V?��T/�ZC9�Kp2<��޷޸i�yיS��g�*��[P�7DrKr�<�z���\���:e��:&WK����UqC�)��a�ﰢUMCf6Lgy��"G�	«f��2k5�c�����%<�d4槣�%���y�d~�dK+Ҫ��Bs}�4�y}UT����7��{��>�o����;��	`�;�<�b(�:�i�(��7�E�"���#�v�(�X_T��5��1���6����hhj�&����k��f�7�Cs_��6��#�0����? ��M]w����=��O^�~���b5cH2�zƖ+�i���Z����>��74�Z�V⼽s�20��ڤ���|�m@�GF�#9��p�F���L�R�Ȣ�Jn�>Ӹ!8�V��f���h1G����:�g�>37+�0���u���ϐ��M�õ���D�lK���+;!w[%l�!��:��]4���޼ǀ�,�ۺ��qu��K�Q�5ˑ�^}`J�
M9�}�T���eh�v�> ��*Q�k�]���>��x�Il�XS3��z �#U\��W�H2�ņ����R�<5��/.(ܯ��Db�I	l �xUr����]������������膎v&�o��@Q��R��>����K��
�������<���h;�~ec�t�E]����)a|WeUD i ӥ�o0M=���n*�j���۷��)����tU�q!�	�-V�E֍eҿr���;-�`��S�G��a��Q�vf:�a��,wU9G	�@y�N�$��z?�EOC�C�齃=���D|�s��h�|=��r�`�zcH�=����:�y�q���nNW�,2�%.�Z��%f��sط�0��V���?���X~��e:||m�Wg�|v�6z��̠^ժ���Kl �(����-d���Μ�Ǝz��y�MZd�_�'G�!���1�v�cS�Pe�ЍH��'.���	�N�C+��-c�$���S��m8r�|^~�	��g�H��VS:8W�{���d,���:N3������_�5wV��š�c�Vr0[u�v��)�`���}���OzSy���@�ג���ܽ��W�W������=�[�g�%^!��x5���� Ɍ��4+'xG�[QGx�z;B<^^��cw|��ˍ�6�*� I���{ܺo��CߴhnA��������&n���D+-&l��zq��0i��E�d��(�3�?�)���]9-�0�B�`�}�(�m�.!�Y}uT�%�Ka�)����Y��J�w��QGl%��K��.�&)��
��rdJ�%��b�=��"�� �޹�j�e�+�|������-p��F���6�{�^Lz�kWv�l�Χd�i�5��7'~+��d~X�Cr"U���v8�l�A���q@,��PO���q(Wq�EI�>��#��%��o�Vĸ�+}4$|����b��Z���b�<���
�.���O{b�|���[.��T���k��C�{T����������'�(r;QI��ַu����w�>c; �KMG"v{B��C�`<H�J���A�d���P.�����K�`B̽��3C{د'0��4	�Yй��Jp4K��%KP@���������x�R��~�����ָy�
`Hn�Q�����g�ʢ�\_n�씹�2q�@���=�b���J�Z�����ԮHO����\�5���R����-֚��jZ����2��(�1;|�Q������1bz#A�H�X��.e���!�2��Ԉ�L4��
�Ǚ�V��|�0�Қ������0$���Iڔ4RϪ_��$.�b�v #·Yp�!w;^�0�I��<z�C|2���hL���ZE%ɑ(������-�P��3�V�,� g#�,\s2̀�7��L�[�C��F�F ,(&��)�,�`ǽ0J��|E �㈪:��	��	�)9p�^��d�Q0`R�߅`Q����K�v.;q&��2��v��x̟g�F��+��?e)Qe\@G�(]7�N���"�E7\�u.�X	E>�� |v���@�؋ *4���Z6��;"@�Qؑ3B�����P�k��.i�i�,c��_1�tq��~��1t頺'����)
�!*�e7k��iE}����|?2���ՐFV��xﳵD��A�̧���Lm����D�K�Gg;*��v6?C�/�	sp�mJ��ֲDW;�|O�JA��ժn��P���X�1hFydM]r��N�^�g�@\��ۼ�¯TF!�\��׌c���BK�e�$c��)L�व"4��t-?�s�.�4ے*��]�C�~�'��"���"��:�D��K��>��?W��A���Y�R}E�S"�Y�����ԁo����ׅ����bd8��m�Ck��Ͼ�,cF��^��D"_NΗ�"�-�A{!�s�����'!�;C�����<B�O��%�uZm47WB�O�~�%=
j'��k���5mFF����t[����n��d��T�q�x	��;�� Ӻ͔�*z8X��No�qq�C�d�]N9GG0��4rw���ҙ�ن8�s`���Յ��{�jU�wY��������NL�ovk������|`�
��V+���g�J�3��3Jz�?��%ޒ[-Tb�U�D���ҧ{*s������k�Uі�<� ��FȦ�q���;��$��x���Y����ϡ��dhڃ�I�0�G�����䔳6'��Q���YaM����a����y�&K�������nݷ�>�+M��� j	�a
��r���X�<t�VƂe�2e���^	��xOT4����`46�p��M���]�Z��[�4�;�s�C�"(*��O��Qd�Z����ue'h!�_�P���kg�e�fH�&��/��Eh*������2�F"���q�V2�$� ����2�,UZ����x��@Kဟ����ٍu 57�ghV"2y�}m�Wg� 1[���P��\}���2�I��@e���iWB�Ӑ��bv�����B=�㗯���q�Q�����|�)S'm�̻�c�D*oc�tb��ڠ���Rx�
v0��s@д�`�:^�o?��+�ݛlH<A^wNo�6��_��Ŋ��f����;I�;ګ)�,-(���UzK��V�܉��jb���g����RP���;�T3j�͈�B�t~Y<#�*��c�z����Y��� �K$����#V#E*�E�g��j�rj4Q���~�1v���L���UP� ���*��!O��X��u)iM����N������"�^a�D|M,zf�]���1ScU��;��������fI�%.��(نy�0A�J-����@  ���%�b#P��IF_u��Is�\o("^�*�f��i�BJ�\�T9]8Z�� C���(ז<ӹ���FMݫa�"d���S���@��+�w.
\��}\���A:{��
�%�ǁk4����"%��#���бҺ �0Q<C��t1u��qdg�k�����4fY������G���f�²I��!���oKG�u8�-ёi�ĭ�e�:�>�BU��]�_�-��b�Xq�(or]�_p���t�y�����⴩��ts�,��s4�G|p�ö/��)����3�O�[� �]/�mf���85r��@,�5��Pڍde4O�<�ϳ��.Y�+ϾzI�q4�!_�,�CM�����fY��Of�����oX�*����,���>�[:�:�-�����N�__�x�|]��fq�Q�H�ώR('!(�m�0񅗪Ց��h�U�C�"����sZ�l��k�F?���'*�
d�|�L�)��־�Iv�����T[T�����Mb�	b�rMjfD ϾvS����PyT�o��X�!�q�ZğQ�����BJ��#���%v�:�,�j��t�k��Z��&� 2g��8��t�iW��'�T�����n�~�������\F���sTG���h��g�6���V?��<D��3�Q�=���]�<�mɺ��ڳ+���m�F������M��`Ma�]D��/��
�8�> u愚�A��$�:�C���
��|��u��k���iT1���!�(H`���8�:��`�]A0b���Kx��d��Zw	d�ْ,�^?~`*���{���;	pg}
�o�w��@�ay�s
yyHC%�K�|��f~�ӟm/o16C������+޽ҵZC�E4���'Zv)����=GW�S7@3��E���3��L!�۹�����q\�s�{�,�e*�g
������̝[�V�h�Mj~����f8.�g�y7���w��$����4�n؝a�0��Gc�zV{6|�����n,p�
ɉTA%Ӣy=YЙ2g�2�()�-�g�*>��o��-�-�:Sc��{t�級݂5bXDA�Է�&F��Xs�#����q65���_;������ ��T1$x9-�-�i#dXMgi�Z�Ո��$��y�n�j�H�.I5#�-Վ�������z٭c	!μ)��M �7��Ŧ&:H�p�Hj�3��Bfޚ������u���	�q�Y�,�MU��PZ�g+H~�6
7�y��n�p����y)A�fuZ�Z���|%�4.s�8z5k,d����@��L�-N ��(����WK���R�i2/�;��)��+�6�x�A*��HxO��!�ܞzR���v�����#J*_sZ����t�(�|Hg�?L%���P]�����w��:\�՚=�1㬋��H'�$��D�kZ����(���M��A8�3�J� ������#�tH*'M�x��Uk���/]�җG&w�]K�w�V;єz��蝜�����3��ު8^�U�tf���_/Fzf,��� kI�XW_���=B[��v����20�B<�0���%�4��:���<9f�8Tƻow�� ����͝}3�&�C;"v+�g�qoN7��(@m�����H�����~pQ�ǀ>��)�-���{HR�qI`�:}&��=h$x��~�RS�n�VLk�ܿ��<g�4 uڙ��T������u}y����;�\Fqf~(s�%��Q)��n��X�L�D'��.С�x����s�x�p�WR1������Nk��^��(�>d:=F���fϭ�-�"%�P=>4Y�{�wGN�P�߅�_7�ռ�\n�*��dIv�uC[�6�&��X����՘:mqo�rwD�I.*=��v�̰�w�_gq���Zˏ|���Ѵ�h���<��;��~�*���L�NB2.���o�G���Z2~��S ��G�e$��z�I�?�,%Y�5���E�ϟ�̙싓FQ9�U[��c�*�xdi.����V�=) �X�x	^��顠,���[�_�j�V�����'�qxR~<�?K�|��e��NMK~�dUrKZ炛
��	4dS1%a��m$_R/y]d��$�Cȩ-�'�f��5pײ:z���vd�����D��5I�5�s���A��O�.e���D��ȋ^�_F���(L�	�e��"n��<�C-	���s�	@L�<�����WhG�C��
��Qr�#���ux<�N{�ϓ����Hl��e�z��j�(f�V�[`��C ��m�$�;�Z������v]��N��}�:�pyY���wb�T��oצ�i�����Ι"}��(�Ԓ	�ߝ���4C���q/GQ���L0�?�)���������K�%Q8`��E��3�Lz�rj��Y�	��G��^^tH�1{��[y��!"�Bl"��yL�IL`���i"�y����ܗ��$�?�L)���xGvG|���_l�(�=�&P��C��ʏ�/'3β)) ��,A�?l�0ߢޥK����@
w��s4�3��.`�"�p'̴yJD)�`z�;鍬��@FRv+^��wx����+_5d�S��[xH��F7����E��sIr���z��E��BO5U�bA�ݿR4u�sA�􅪁Uf���2�N	�tQS����jY	O�{>6��@H����|��4�/g 嚘8��r@!�����NfF���v���*����+�Ho���cl������.������̲e�ș����4�9��Wh x�y{ğ�|m�q\ƹ��a&�"�s�7m�����������l���j��_���2��m#	�5�����_ma|A`���6��M'���%P���X��r2�BL��Ѐ�ឮZw��*�e�[���W�ܺ;SQ��$��P��?�X)if�Н�BQ���>ɰfe������Dm�ư�<	r�@��-NMF#-��^�3���H��Q�k�$0<�.�)����c�N;���/�4�;>�؜�����Θ�l�&���"�JV9=MT1{�׬�K"���,����j���Sˮ5���du�X��&KM!�#�_�<߉�g�����i�X���Oujz�]��I���0i֪���}�R����xk�?G�j�<!>&�̡l����H�m�>���|���s�j�f������BM�9�aR�a
�:��Y��t����	]���r_����܎�U�{>ޣ���ہ���S��X�/���,uc�=xa�8��4�j�3^i=p�� �ASG"h�b�Lq�P*��<L��W�����9,*�G��j��t�N��Dmkw\������=n�H�����q;̯��m��G�|�t�H�;7��Z]V+��g	b6DP�+�'�&�9#YS=P��ю;���R��{%�y5QB��2��z�J!�ҙU�8fҦ�W�>[w&�+ƍ/��΢:��wP�^��'~�+ͭ��s���C��W���(��8!R�~~�N��$L�]��&��tz�G��!�XY.n<��]��p��mTR����J� �]��b�Y\�����È0�@NG�ϒ�I:����Pd>���:����6�I�h�K�z٪�+���pW�ٜP-g^��{G�P�;U��_OiY,�7��t�>��@0�^�{%;�G���"#�mv���a�
f1"�;3t���{Hzʇ�b+Gh��o�^X1:���T���w����Ͷ���@��P��K�v�H�K�U>c�	s� HQ�]��O�\6��g�I�91�C?�N�^����)���qݏ�_�d.<�I�[�k����CK�M	˪�جj4Y5�*c�o��7RyÂ�<�}�2���=��4��s�iN�U=�u�z1ْ͝���͂��p5�R&�%s�`5���.���X*)�����^�1�-6��pF�}ϭW*���4��m՚�]��4 �w�k?��xm�kƵ���z��L,:��nR|t&ҔO͠(�l�d�bv_+a:r�́~�$�S���1sB+A����W����R���,���Q����2�u��T4��Cas<7�NԤ����J=t��,hS�j��gN��Z��'�Įjj��*>~p�ޓ֩s^/��-{�n��V7k��}����%�&���m;�p%�i�/|0�{��'��M����2(��\��e��,�j�
���]2�'dA�[�B
���&�=W��<�>��A��I�e�2f�@L��sU ?D�VD����-O�'���*�c��=�VE�V�[��,��L�#S����
�OI
'�;�@<ϐ�7��j<3�/Sn;'�a8o
�Ծg�7�CF�*~��+%�,f`5�%�N��Xѕ֭���K4e^�Mc��T�q�8�1�x�>5� n�,�����7=�^_���-�sO9���'V�M��u�k(5�c����J�j�ڴ�wt {T���_=������
p�����'HO��L?�=�~�1xI�b,��Sd����:�L��LX�m7�H@"�R��<� ǃ�Y��[ 8���-������(#j��M	{V�i�J��N+!���o��%2�&x�.��h�\�IHY������Z�/*<�P'�����L�p�y�RP�ië`�' ���yS/��T�a�����ja�~溺s"�[޼�̴�l�O���43w1���,��5�����gTpԠ�ߴQ|`���K{��nH�NS��?w���O��H6wC���l���f�����S�>6͘�_0y:^w8��H�7:��!��f�M�x+�0*��~�)0�E�� _���Qm1z0�IT��K����f>g�W�$��), r*T���p�kۏ՘b��c��oO�Jz��G��Eȕ��!5�]��������֩������Ba�8\xǞ��)��<F�^e��I�]��`|g�,!��L!��/H�ʾR��B�o�'��-�g@AF���<Ҳħc�s�8F�9g��T�A��Ø����!r�[�3`���d��}9㟽��ɫ������vMQ�lmߟa��^��G7�Р ���6�m�!N}��$�p�U�8�Z�[�d���M�j�p>�䔨���1#�Q���*Q&�&/������Q�2<���!��#K�;%&K��F��~o�sY���!V����I�����􀠯�,a�{�z�iL�믿���Dhz����<K�x׭�3�~�o�(��V��4@�V�92�\��zUC�������A{��NZ���������oЄw)eJ�uI�>;�`��xK���@�4���i�Ah'��zOb�D�$f���{���x���J�8�]��n':�o&�$WK�� ����i\'슣~��T��ס\�8�4&�ka�$�Z��\�����҄��UQL�46ߊm�Ê
�>j�d祼'���Q@��ͩ��BC��64�D�Pֲ�ȗ������= P=Z���T?�f��o��"�Կ�s�
��n�(b���5tTA ��{i�[Z 	-@�`����Zߞ�=O�Ti��mMCj��po�-�A���]��Ɋ���p�kl/jP:3�d����;��隕 ��Z��!�}{p�G�uTTc��E�{�N���p1 �v�Jzڌ�(���\�]6`<�-�<��� y��u0�����Բ&�n�K;G��i6	G��e���U������L6t�v(�ޟq�!�w �emI�wG	�#W�|e
��N���Vj����KE�����(�l*4�ϵ���_i�t��
#�	қ�>�P JGx{ ;���7�L��?h�!�C����v�>F�'L�%i�S�0ru��3����p{y�	o��f��i�k�^u,�]ɛ��_=O��c��ASzqK�����[23�. f�B�!��/s��"��T�fy��-t߷�s�D��l�1�ir��E4�,|9�M�?@����Ċ�ۖ�( �-Y�ZqJ`Z_�zo۞i����\��F�"p}��ǩ�5[,�t)hӕ��+x�޵3U ����dޖ+�N]��1]�z6��on��p�~�g79��G�b��b?Ǳ�T&Aff};�0�����s1
%;?��a����<��{@W}=j��$q�Hpz���	�M,B^vy"L�����R��Уs2qX��J+�9��~D�O	S%zc�M�+�\����L�dv?�����A�eHI�ꂐh��%Q:N�5l��bn�l<�.oͬ��#lն�a�x��w�V��[��9�Ņ�K�m�on��{zEξz�be��$+=	�Ik�Pj$���%o�H[�W���v�0�L�tK`,tN������lǤ^��������Gà���L�F�~2��A�#��[��Z9���1���~E�0?L���vW>cB4w��ݚd�-��NS�	��g�mh�}#��SĹykvc��LY�1�PZ�!�s�
���"Ƒ�=�>*�;�u�g�6r5\��M�L|� ��sx��,iI����}N[����j�������צ�{����pq���J�V�:ޖ_��nwൽ�+�I�Q��D]�@vLv"<^�K�b�~��2���.��Ѐ��#�w�h�x��7D<�L����fs���p������z"E���L �ZmM��W#?�+	�=D���I$<��&A�厧G$�8��pv�F�?7Ǣ��,)��޽�����8��������+���m�Q]|��:{`��*̒sP�>��e�h�Rd���^ʤ�MY��1dxZ�]�	�����,{;�����K@E���1]���:Z���(��e��/G�$���U\�U߅,.�|@�5�k�{+n���o>Y�&m���.$�5�zf/Yi���ʠ��\����n ��.ҡ_�(�ۨ��t���c,�R�����oc~Ż�	v]���GaƖI����[uT�L��x^v@���0�5�ƿ���X]�=� ������C�/(7��C�v&.!�����Ռg��B�e�w���_Ƴ��m���M ����j��t� :�UnM4Q4x�n�x�s47���k��TN��9k�	�j�CP�s��Jv]���uh��d�'�;
�!N=�3���:.�^_�0�
F�D|gƫ��`�@$ml��3$�����)w-_F7�qb�l���wrh%NJt�W�y w6��,g�UJ� F{3x�%�Fq�(�I�_̧G�#�P�d�u}�t�t��� �k��M9�*���Ҧ�J����ڞ�����}�	#�����o6���?����Ж�̓o���_|l̟�-�VI��:U�uaR5@�љ|��;�Ɩ��#$sb�73#��v9ꌦ�Pw|#+�K�b��۬W���j��������������d�=�N��=ܚ�
;�m�Q�e[���H�vV����~y����"��&�36^�Cօ�L��������I�����O�X�}jFS3��c�=�Y�U�v�/�DD����މ�s�#�¬���W]&υD߸|���P���[��Fb��A����8��p�=��o�8!�O���,F�:�
��|HP�y�B9Y6���8q��?��n��n���X�k���/�my+FCFEZ��Y%�s�%��s��OFKzP��CVLk�l�^?���æk��S���㖇5yiZ�A5����3�(�~U��7�9�GE�5�(�"�tB��*��z�Y�%��q�5 ���㮺���uk��}u��9�{֞CsQdh6��;C�l���0ՙ��9p�a�L�o��[�_I%m&����ԟ�X��7]��+���Y>�j��v�M70��ĉf-s$�[^�I0��(�ܑ��i�{D9�-3�V��>g�=�iS��!c�+�������Q��t����B�a��l���3�t<�,'X����V�A�/�:�0\}��(k4;y��(��r�����9=�x>u��!�Od�G�o����n@Sd\l��=c �H�ܴm>V!��Y#��&��!�9��*.���{���_c���o#��vY+i����ӻ��G"Uvۅ��^Uh��~I�_��+c%��62��)��5ήK��П���,�7�|]��s�V}6�]�z[BO�����q⇉��M_0tڼM�������I�@P���K���N/��U���OH+(�މ����y�,>z�[��>6��Bv�1�UF��	W����NJ�}e`� f)�1*��ڪ��\���b-�W*�W̎m8�o>��a7~���q/�'��K�&���y��P�4q���_POk4�-�Yr!�lsi��� ��B%���汇��5�?-�luݼ���0��/�Ю��������J������4��An���~� ��1�*�n�*���ɢ	|���wݎ��_���������F筁�C�>^Y��q����zߥ��c�mO�}'4�E�U_44!���!�,�@9w��ƶ	��N�ţ��
ُ���y�:���*��,��&S�t�w�$���"/*5�V�\�y�K-����ɬOl�X�0���J�yJ�|cc:�н�r6"lF��&�q�������wY�,�@�v.o�M��7DW�Ź/H��G��9  $����3��Y��X=������B�3o��n��Y�Qt���YH��x�^�ʣ2O�T��Wy�0F���t�p�M�Q����&}xv�D&c�ȳT�0�6��{)g�k�l���c�N'��{�^U����::�?����jE���<{�U����JP�4��Qn�~ݓi��?��AB��/2/��r$�ݍ�1��>��O���7����x�x�߽�O��5'���b�
����h,����v�:�.Dg��䜰��$J:�v45�8,�,R�9��	�������S�1B�4Br)�i�ܶC��w�~��^���-_*%�������̳�0����p�4?x`x���>
�_#_�!�Ǔ�:��A>/;;�E�AF�s��q�{����Q�	 �#�OK��'��x��@�4��&��O�R#�v��ړ'j�,����U��d}�b�8�]�Lx�p�s��z_�@��ĹnBn~g=� (�A���s���4Oo�V$D7����'Une �	wů�6~FP\
�����褍�(����"�z?	E�X\>0I�s񭢢"
�`q�7s�3w��Ao�s���ueh����1?����a8�����[��?��C9��4����sĩ�X�ڑ��J�`E6��F2�:�Q��w�hZ�Dd�L�dӥ��>���G���	+��É&���~҆����w�aR�΂Pr{�����Ё�2��_9F�!Fg�	�M�Tp�N�i^2v�yf]tf9���cDh�  y��a�dN�t~%��c�d'c�f�"��y�.-8$��[k;D��������f�İ��u
&]�B�P1fN
>�Օ�ނP�)+}NS��?���{��i;��C�w�������`� �'���B�ؘ��vǐ��nW�����D4DEz{mj�0yOe}�
�eL5r3eށ������W�4 �6m
��i���O=mFc��k�n��/��y��'��0jBQ�@��	���4���������
*f���	+KEo<�.�^ov�w'�R�J���L��0�p�����c>�����TN�}��/C6��J&� �HV��}n�ˇ;�0k���L���*'�)6���	�p���&���+�	,fu���)tb�_X��+�Ǩ���HVf=I����چ��
M$�>SO�z����/u���5as'�i��*�|X��s�M򄛑;׼<�h�#e��m��l�؟CX,�q�L$	7\�F&���i�.s4�qK.�I3ԏ�+��_�ǁ�!�yI�_�Ж{]��k;P[����M�~�Ẋ֓�B�%�̧��rm��y��e!E-�E�� A�t��ת;��.iy7V�EB%*<;!j�(�M3�~Y!x���
��?�F��������e�	+l�N�?(�O�=�ιg%�[}|}�m�'D�l"l)��t�2�ʶƅgL�s�"�I-;U9,��w�q!:W:���>잋�͏�c��$�By4߮�qrK�_eI�]�Bs�ci3��v�B���=\��,���Q*/�2��e��3��2��,�� �T����Q�r�O�bEn�K��݀���r�7Ͽ��2L^��VK'_�r���`�)��b�M9���N�U ���^�����<���u�)N+��_��`0����n���ć�&r2�G�E�w�E��K{p������;�L��Nچw�+�\�S�W��,�{�@"z������d��F�����2bxUFT�L92��;��m"�ۻ��`�(�;0������?��4+��@��a�s�
+��}4?�)�)\��:��G�W�}�Ɨ��|c|�u6n3���@����΀䅴�'�B��O��UFV��mX�I)�]`~|�
xW�;鋅�����}�6XfV�l�u�~���7��v��9�8��� �x��X�ה���+a��_z6�#��RkN� �)���~W�N���by�5z�yS��;�f�S�h��+��0��`�`p�Z�i��:�;%Dz?Y ����xn�s}�4�ʁ%2��Yz@5�� �X�V1����Vy $q��<6�u�������{�RU�a� wJߺ�prtP&�����Oy���e'^bN��HX\��>��A�����sjǀ8�.9��{y�����k�3��#C�\�Z��X4���zэ�z���R�*�5t�L	җV'嚝(�ȃ"����b�J�ɹyS��ie�
4~RMk��9x�@��}h���>�^	7��}�k�����{Ǥj�l��dA�����"pI��ka49�JLGS�z2�N�Z���rJQ�f��l�պ��L~�zgd��D�h��;1O���#B����?ϭ���/k��F��_����]TĂ{Ztm�1����k#���� )����q��G�ϪM9S�>lxq}uC�~H@∌�H�L���q����(g��|(g������i��^�A��u�
�k�?�����.2:u�{�hV�E��R�Dϐ絎�s�\p����	��r� �K8�d ��t��-���\e�.����5�I�@o�&ci-�K4% H�b���n��<]Dո�-f`H`�A�11���	xI{��u(�SQu���"�Q�E����Q c`(����-�)[�B��2w6�n-r����&t�6R���+m��>���.`�����1��,�0�Q3�Ig�)Dc���@O֯j��~��Jd����	m�7�jϴ�7p-���d�֋���'0���!��]-�*�ju%zK�?�u#kq)ȁDK�V5k�ʟB���R��RhV䇤��h�y��U}Ab�0|�/���5<t��`a�����wB��|���Ea��Iʅ��#�t�������=S����:���;�?a�t����~�%к۵�|}ߚ�*;�m�� 0�ZkƝ���5�7�fX�[��(y�����63[��X5;�-�ّ�&��p�{-��ȑ/�.�l�,�!��
P�C抡!��R�%�C�c>z�aM����ne��/��+<�}-0q���;Z�n�s>	��Q�ᅃ�w��v�e���D;�<!;���*;�I�Z��Y���������4�>{���R[ܩsOu�w*v�����G0�hl�o��AR͛,7�DE�t�?�n�ԴD�܅�|V��(R�\Z;d�b��Ʌ��l�p�|RSa�������u}%Be'2j0�غ�DJ��F;;L��8(��+������ c�ʿ�p���Gu����n�D��ר�L��"�QN��PB���Ӈ���z���
Q\ʥn#��Rc�'W>��
�����s�|��J���YUn)�Y��[�W����{h/m�Bl%!)�δDȹ\r帄A�:���:8�+��q�u� O'�xe�� ��K�M�����}���5/
�;�ȋH é��.��'����\�0"s�jBF2��0An�7����p�^zW��!�*LÃ(�;b��K��+>��~ #��wD�_,�2ŦQ2�\�)B�V���-���[���b9���_y��#��L�3d��q�L͈2�Y��C 7<|\���,RJ��JDqn�> ��V/�p'��y�������	�`X�,��\v�:�U�D���)s��18��WE�5_9n�[:ސ���/�"s�d�&��:�~�HW���`�Ҟ�&q%���h��Xq�VQVy;j�)?�)멜���*T<v^ 0riv�P���6Ә,�S]ʉ��9��O>l-�ft��#�(aň^�M��t<�	 �Ù',Fl���`>3������Ie{�KѦ�n�������]��5?��m���j]m�_��BȽ+�}�G�"�������V<�Z~��h�hB_���T��R�d�k��M4�2�9ā��������i�1c�9�=	 O�d_��<}�Q��{�8l�l���֣X��D\�P�Q�������1�v���!�O�a�y}����<M�k�q(��X��L7��qW6R��?S��1�����l�1J��������k���P�z��m/�;������8?D %�J�����s��e`7N��?�x$����7��oRG���Uo�r�b,� ʸ5��N,������WM5h�уX8vfw���u��h�y�1���O�:+���4wd[�b�|��AM�Fr8w	��|A@�L�G3�Gmq7�Ia@C�Z֝�ڍs��bY�^>R�Z, kW�q&ړ.> �<��*c�+���S��>�������S��cF��-��՚5,�Y�#d�4s��(���#Ǣ �2�\�*=�|	�r��Tz��BO�o ���ӧ0����%Vu���v�D7+�L�	�3@,=\�.�9�0�kQ���`EA�\SP��1D/�����V�/U�=�r� >1x�w�����jJ�I¥HP���*����~�w�b�u����/��>Lm!-����v<$I!)�4�x�ˢ�_)]fь�mh3r�'��� ���
� In_�Ê�i����ED�����H�NƓ�B�����#No��5פ��e~���G0�nf=�fȼ�2�������+��5�-���o��k�x�~Ø%�GɔEߕ�w��t[��*�O����|�3,���Q�ZY��Կ?G0��	lX`�l���$v$h�J���b�hm����˼�m`욵�1H$[�~)����Z�Y� �qL�͇]of�ז�ج�����8Bk|]�G:K����~CԁI�0,ʙ��N��z���f-�w�[>�uL����Z���E9j�F��Ŵ�1�Ld�Q�P.�������WD
���P�QlDq�Ls�C�P.Qg^4����S'P��a�p��5�
�����T�ѻc�hhŵ���Ji���hr�7WR�®�>�]�IL�
O@Ug}󆰨c^8LȜ7=�S���5L�a��sB��{��Fz�:��:�@M���6��I��3��p:�5�����S˸��ٷҹw
x
���]���!D�m�$�l��D;D:xD���Z��x^������N�����lP���46g(�5���#JM���&̯�3��D�t����S�2�� C���� �U&��R-�2���^Zq$�ԔL$��0����r�Ι\Y~��a5���(àI�ZՁ��Ҍ�}j��1h� ��\�3a�DElz�n,XV���,0���vG��ZO^�*��r�]��U}W�.{��%���{H�!U�M����)~߸�GR@م���n�p�A��t��jqN}�l�I�}K�P�+5������u2/^������`S�o{�{�J�l�s���Oн���-�2�T?��J�#��0u�����p}]�{hq��U�v�qa�Pv�)یm�3�x������6���cQh��4f����iz�=��z/F�1���:�c���":Ι�v�
��)N;���ߚ=8��}�N�z~@�DΫ&Nߡ���6��@#���V��ͬX��?s��[̥�/� �&�ɶ��.x��m�&ԜmQ���Ј�E����b�;�!ȍ����-���}�	EH�bj�:�XD�c��I�a5Z����_����D�E�s,�!g�� N�RK���a���`8jjJ��8�{�[���k]�M��;u�o��&A���Zc���:T��������b ��~��?/���j�������`�EEf����3FW\�����N�'R���	�V�U�^�*�n͒`[�쌕Fs��+��G�|�zi�������s3��~@��@�������a,2Z��p�3�����E��z�e�ux����d;���]��!���d�܇��C�c��X�\>V2!�ܒRy��*�+�v�4���{��R}��^�����	QK��P�t�na/j�7��@ά��x���w�0��HT���� ��c\�L�w/�����ֽ����;�����:Mᾴ��cb�+4u�N��(綸�[Ik�Y��0�n�t@��%�k�M��|H��#�8&|E�k��J�����(�on5��:��)P1�b�}��٢1�km�EA&�E�O�Y��7���l�'i�#�hW5�Z1;�ˑh��ٽLqO��M!˶j�Vtu9��'�0t�gxwިt;�Ԡ����)|DF��6���抧z��)aϓ����/GkG��X]fnc�P>���W�t��t"S�&E*�i-�Zrin�����g�
�c4��~�3|K[1����#�0P����(ĉ~,�������Oi�ŋ�GAe�:~_l�>Tb#�G*�(�����&x��f��Z{����&0C�ǲnnū͖|�γ�?�2>���J�����x5��v�7W8 �i��^�����Jυ��?��gX�Ԛ����OR#�u׫�s��-��0d"�/���d�?�_΂t�&{�~�/���ɋV25*,���`i��u�����\���VCv0�̚�֯q���)�d��>�8m{.���o�u�Ϙ82�kwx��^�^�r���MkM�ov��D�5���rvi�������C�:�}#M��V�[�[G׵�����4K�0��9����Cj��|�9�K��KNC;Ŷ���,>��09\���� i�B&��&�����b�ۯZ����SV�*��_R����@~�2y�������$�ka�T ��n����Bha{M��5l��	��9�K�3S������R��C�����u>��Y���6@c�t��VƉ���oɔ�(�@8�QFR�?����g˿Y�-�#R��:m*���\�:*��n�+���&Pӂ)����Ȃ;�A0�a��f�:&�tGg��2����Z�d���cZ�v|×�U0!�+R�%�ŏw���m��5�9>-2�h����5 �3�+Y"�� {	L<F���Hj��Hf������c
y��s	 ����a�.]r��m�&cH��;��~������|#�#���8e�&�
5=��i���<9܎X��,���[�f��~A��vK��|8~�� ]0.�厨���5m՘��m������6�?�6�lɊ#���i�oP�TzL���ݼ��BA�#�ʵ_���ŚT(�
w�n��Y���C{}|�ċ>C�F�,�����KjAR��_n�#��L��>��t��q���]��t��pn �|k;ˡ_�+�EpVe�u��Qd]�-�$��Ǯ(N�V����;3��f��`s\Ù���y�������8��,ǩo�k���ꬤEe`F#w���tQ:R�><~!��^x����;��B���\X�K�A�.I�n &h��D��c�:н|�'�7�&mr{�P؜o��;���c����'���G�=y�F�����6����7��k��h)����7�V6��	�z�.n��+ŧp��MZΤd�{7+c¿�Mk��tEx�}3+�X?K��G�_�VD�k���`�%\�Ħ�}���rm!;"��cG�h�8���j���M����_�c��#��徰[Q�mP���kw���j	92��U~��b� �E��L�}[�y��$f�M9-b����f��x��ۨ��}�J�Vȱ(�n>]�#���|�?���KG)Ä�PXۉ�g��/6 8g?��Gۗ�f����6�:/Y��"!K7�v���ڹ؞�)�-��	f����`u��y����޽��N�ű,��R��..-�gP�LZ��c�õ�l
���e���2�3�n=�������3{Y�{h��(�v�y%]�W��[�G^.������$��A�S�m��v��?.w.8҅�
����y@�^����	m��&����f#͜���H �l�U�0�����?tn����'yl����K��@��wРN�fN��oZ��� ����5^�� A�>Fi����;i�H<.VZ��g�����0���\'��z3X�J$(BƁFŇ���J��p-X�_f?`�ӑ�##dA�ꔥ��ݦ&{�
]HZ==�T0��M��i�}"��Dq�'N�����"=�����U�:,
�89K�
�;��T��,/�N��g�l&(�@�1�A��T�v�&�7=E��oʙ�={�����K���*啅l�������4�����K�=���Ξɚ�ڝ� ��]=�lAZ�'��n[S7���:�~��E{H��j�1&Xs|��X���H�3��7�Z>��@�Uj������v��/Ou��#_�`rA�Y��W
M>���l$/[�A+��FR[X��7i�啉9�I��x��UL6'"�	�Ӳ��{Nʆ�,�DV;��<�A?(�Bo����Z�]�D1E�м�У��!�3�oc�V<�����������M_,;�R�p޲�s	�>	�������4�@	4u�j	{,�l�����O��Bu��߶�\ҵ���8�8�}@HUf��:���/������X���{S�9{pj�8n�;B�:��Ķ��wߒ�l�Bi=l��E��u±� �秪�ӟُh�zD����c>3�#,��u���ʍ�� ��Y����8�:���p��zS	(&q]���4��=<rvP>�M��<Q蓡w5�"M��h㱷,��K��qp���؜d�*���u�?�0!`�_&ׄ1D�.p�d��.����a��+�]>4�̖������2��t �O��ɒ�WP�;_�yB^�\�CK�t�o�b��1�.���:�<�0+g�&F�CL;`����h�1R��h�(D+��e!�˷�=�h��?) $�0�"�4�#Jm�=�z*2�n-��G'���Ǆ�4�Y	�U<*eI�'������k8B�bŎ�$t)�O�]$&q4M�݂�}�� n�R�"��!��qTO8�q^��)�;��1��gC0���̌�A�	ВUa0y�d����l��c[��ƙ�`�A��3�����-n�Ƌ�c��@�xJ�T$��,��evė�ūs=`���.ˡ�E(�|EߘA���
c	Ҟ�q�����A^f܄�T�=� �Y��=藏`���W@��v�]�b�.�x��Ҏ"�Z��R��Zd��s���7���� �qzB
��$ꀋArIo�� �����!~��c�BB��Җ!��Es�=��[���Ǣ�<���8���������9�� `�#�9;n�v�N���Խ|����
����lMb�-}V�R��9���� ,������P����($������z-\��1i����ȗ���5	b�Cg�hQ5�@Oj�{m�cd���	�B�9<s�&���v[��w�R (ם�;�r�п�_�,f��L���H	����'%A�낎��j2㸲�4MUF7�e��Dah��Zm/�G=|z�tmcռ���պ���~�=�
r"X&��K��EoZ�0��vo�賀���o����n�C��C<ݘO�J�|��������<p�X,#�M@ŬrkZ0�a)�GC�r��nG�eҭ-�c<;�Z԰K�L��C_�ߔ!�q	RxBC���s;/o�"���Pw#�~���F& �� �K�\�R|lp��t�r�����Z��H�\����A��=��*��b�FŐ�Q5��,]�J�jG�4ڡ&�H\u��;��h�G�����;�H�_ �����Z|5u��'bh8���,���`��ݭ(j6�,�D	W�F{��=5 *�s����2�����3�
D�h��u�o��4���&�FC-�/&��:���M�%���'�b�)NŻ�Ss�h�ȀOz*њ�6�Cь.`n���-����@`�H��/�����ә����of���%��O��NG����[��$�v!+=6�rՖ�>��K�v�(�5Ȱ��-M���C��~J%oV״���͚���m�c�DT�f��z=��n5�h��!)f �s��y�͟� �rw5o�L'��]tS;�]�L*E�/��J��j/T'X݂�
�#���V(��L�2Sg;ԈIE�3�Ĉ�>?>�V������L,��>ubE�:뮍�O;���	������d��߫���S�e{��o@T��d�d'N����#C�oB�է$��� ��q b���"9[�}��Ƣe|Y���0�@Hu��Kw;���=�|��y>t�UkDfUa�*��b�H:��\��4'�6G�#b� �P~f�L�� m?�L��[u�됨E�ќt0~��BT���q���3Xt����������5��rtZ�8q&�s��Ϸ�eZ	�n���rZ����D����Ü���^��
�V�l��؅��{��0�o�c
�d���@j��7����/��)�F���ȭ���<��)�t#xR~�b�~��'}Q̂��)�R�Qu�P�JB���K�����X����P��X�J�נ�ѿ�t�#��SN/O�T�v��%�d�-���u;Ca,�����l~&���������_�q,W����אi�<��)�D�eğ=f�����>VGV揙�? ]s3�S�q��]!:֗"�C�4��z�0
}?[��p��sZ��4��gfC��S<.��՝kc��������f��'��
��Wb2$�yi4>?�w�3_-��.Ǵ���<P,׾�"9Q���P\S#,��r���\�� �T/����%g[u�"���/=���2�ܲ��:NA?"�%�Z��-��������!Wqj4��V�o]חySxM��t���_(�
z��l���cP]C�)1�e�o�,�L�X�Y˲��(FP�}J�݄�W�/UR�"�>l���y�`��w��4d�9g�Vo�P�B�������رcG�t>�_�-�YF�!��;�",�5���ͬ����(j��m\Δ��Q���p2JO������]g�v��*�O}�5.�����<#,�����p��DK�b$C��>�Z����[h�tq�1��_�!���m��qѥ|g��K���W�h���1�'r�#�_����;�ԭ�8>�{��q���Q�z�{��Ր�pl��g�)Q'Sg�be&�a����A2"�j�yKP>.l����$�Jz���G���6�o�n��z�� �'�Ux��l5���~�Vb{X��X����V�<T�.mmV�U����T@_�a������\���%\��[����<��P	r���L\�1m�DSb��l�]���T�=}z�S$N䋙|�ɵ��N�9�K�b�����h����w�Bj5 >�>�yl[����o�[�_��B����j96�rެm� 5������,�/�'����iQ!Z�����C~F*|��.���i��<ŉga�ό8�o�Y���W��)G�ɂ%�U�h�'d�f�1-Q���}�aOLZ�� � �
q͕9\:��7����V_�ҕ�澁07�@{�7w�ɦq���4��u����ׂ�nR��'ۜnee׊4��Xꨴd�_�u�Τ�:�訹����D��;�|MUy��+�N�VF^4
[��&R%.+�f���b�b&1>i��KD	�P�O�������=ĩ�?kBu����V`X`}�%���{:�[�d���`�,+��jq{�r
U�q�#��òU��L 	+���%p=��C}j_����uX0�|	.ŴOM��2ڗz��#e�-�b%����s��܇��0��/��X�$�8]=n�E�H*L��n� �-l6�S�Q�ݥ��#�Jm�?:��cX�V �:���B�|I���履���Z,�G�������/�Y��s�v��g�`2�	u徕SsԳ��Ӽ��ʕp�1^��J�?�t�e���>�ıͥ��7H7�܇ҎCJ���C�c,�18��e�n3�5��pE	�;�[`�@�_,,��ik�@�?�}J�F"�����c1>y0<��m���ڽ�,$XAs�Eu��&v�l��_���9PL�PNZn�������u��*��N��)W�����,�d=��@dtP��x;����@Q��~!�½E�@X;��<�os�ൢ}�[�%.R/Z��}����y{�R/��A��L�U���c���a+�4á��ny�B��D�+,�|�..h��;����ŧ�
"	(����ßp�|��:��Ii���������gn��dώ���>L�v�h<QpOg�/i�=��R���D��ZΏ1�B)z3��O�~��BȐ$ƝP<����	�š��1s&-���6��� � ���7H�B�WwL�Eˁ)שԠa�fw9�ZvRGSBVb��h�\�T����u�K��������	F27�`�"y��n�J|��x������ V��SB,����d��M��}�R_r��c�	Iͬ��u�L�0�Y�}���(�P��gV�ޣ����>E���\���}�n�b�!c��u�&R��:f�{Z�J~�-��}�ց�ja��6~��&�Ir �_xWW���Gf�BB(�C�����l88B���?4�..ʐr�f�9R����C�+:�MiAgQ
�T�o=���D�*ȩB�w���M]tU6]��$[c��Tk�0~��_�-i`11ݟ�d�/x+�k*�x��1�c�Ȇo��8<�sq��-9#�?u�$�	|Y	��m`��ʱ<�)��D���a��B�+�H*l��g�r��j_���+��C�*MI�м����� �\�[많�X����?Z��V3�Vn=���ݩ��+�`�G���D��ٷ�d����'rk��H[t5��R�_e���th�Vm9�3�.�|�]�s�~��IDL��8�����<���7y֋b�ߕ�����=fe�N�t'��ŵ��R���s���]Ù d�6)�i+	-��h$�������ںn%|}~;~6��
���9�1�E�ωk�(VI	�/�/L܈���`�2��y��Qbe�צ �qo���|��98�z�9�ɘ1��1/1��7������Y��j�鎪���r�I�<���
-�E:�nNUQ�v�Twͳ���p�q�p	�����Ч�"�F8u=��o�CQ��xWyXIbe�?�d�S�=ל���z��$־/�6�f�.E�����v��&i⓯�6��ˠ����(�Kw$~�����9��=r`t�JHז��ƮY�*5QwGR7�ǰ&��P���w�,��1�4��`�7cC�����bo]���R�
:zҠ@�#"#���-�upU� B��rٙ�����O4+��r:�a������=�|�����c�\(eAF6��^�\����:k�0���l�Ӹ��2Ǝ9F8E�¨�}�w�N`}���6�g�gcš�j�V�Di;_���V�J��ae����x#�L�Jغ�*�����v�\�����6��~4�wD6ƚ���P7׉�a�R<g��ߐz&n4�C�g�9���#��H�~Z�S�X���N��ћ��K��1ۀ�Dy)���*_Pƪ�gi�ʾ��B4n��M����&��(Z&�%�v��c�FE�\���rkj�����}����v�.�Ki�^�;�hҰK��+�S��:������ui$���N`�	b�Nli�4�}�(��/�i��7$�{�xJ�c|l]p9�����i#���^��L�2���-����8*'�n��bNж���1
K�s51S�'��+��ۅX��_��cL������_%�:%>�C�p���Q��Ap���Mм0g��`0Ɏ��Oѓܯ�^<�bP��hFP&����Z��NUh�[�_�-�*�6����2����YZ>��xҚ9X��.�ј�6esA�0&��4� ��Q��]H%����# �MPL�J��\�N�!�v�]x�=o�$�2}n��^��{ 1r��3<]�7�F8r�e^i��j�~Kv��̑�^-d�=���Ón�O�q�8��jE���^����g���/|�n%J�E��o�4*#X9��_}Ж���"I��;F��8���GA�	c'wA�W��b�@�{`|@��9���A2�^٠9���
����?���1�1��mU��Y+9��wvR�k��-h�@l�[z@٪�w㠘��I��/GdZ+�MV�8k�	K��i=�Xc�$�_-�������o�|ޏ���?�����4��x��7�� <��<���ZR�"��LLr�R�21ˡ�Y��ʽԺЕ���������TH��ҮtNĝ�W�������_{�9#�w���7}ih�\ވ�`�
܊.`������u�����,�:�����]���� H����s$�b���@�bu�3vP��&�<��D�jߥZ�v��V���r���|�v��1��_�޸K�ܖ���N!h�2W���F���\��GM\쳔;O��5���a�vM����X~��[�$P�X�r|.q%���q5��W0����qzeڧț��۽�DXR�-AC#���[b������k��9�d�RF4�jI�Aêd����LH�pu˸��:e��OT���ރų��_��M��u�f-��1�V"5u��&n��s�k�<���|g&���de�C�H��sȷ�d�-�٦*+�R�"��[�*�z����h�����.��{�] QP��
�I��:�;m����엉������b{e����"�D�-W�z�_�6GRR�IB�I��j��%�c̈́����!��E�a����it�\��jeKzs�� j�Yق`NT��v5�k���ȪuR�NX�+�%�r��)4٤?�\bɻ災^%� ;�-[t�R��~j�{��)5l��#��AB�"��?F� {��+e���Up�&�o�(pۉ��y���k�M��֌{8M*�]������DĶ��	�Gj\B�E�I%�1�T��2�bz�4��p0y!�]����A������+#EG'���~6����ư!��dZ|����Q��*oj�V��y�����2�oNN����ԁ1xƴ���T�~�4 ���'�04����@�G���FSGWz-(w��y�%����lu�7t��><;��a	�l�/�=
ȵom��~��S���A)�E���$t_,����k7&a<k�Ï�e=K��[�����:�>m=��>�p�R@z��;��u�0]P�ϴݓ3w��UM�θ�Жj�iz��C����q�#P�z�_#<��i��2�]A���.��:� �������'�G��D6�W	r4e�ö��K���&�6+��a|�,M�dNJ���&4�뺳�K�G�:���|m��ԧ"�,��s�ʗ��j4)�~f�x�δ8y�ث�������dv\�!�ǑE�{B������a�BZO�����Q�k��bb�k�ik�:ҝ;����N��:SltLsȞ�HxJ�8�#���hEI��۔ઉ������}7) B��ӟ�c2��W�����ۨ�N�&�a#�$L�q��J24�Y�O�q$Yuz!�욈�t�O���_4���]�7q�
��;S����o�E�9o�X��rp	�B�?��?��wT^���,dU`�=4V�[���]��l�eYW�s~h����(KeWDC���߸����=�$fuߊ��;����
0=/d4`-Q<��J��y��zo�����' ���C-��{1Ee���;��Tơ�%�Q�����6�j���� ����L���Z����锋���Td
��⍘�,�c��)V{jn�G匿cY�X�M!��n/�a�w� �[����lQ��:}��}so�7�y�L:⩒LQ^~/E��t�v�p�2��=�R��q
�Aa�)�	er��;�A\%��A �T�dmf����{�&�&^W]�c������㘾�� b5r
z�[�Ko>��&P�j��EuV��*d㤃O-��Jj��j�wC؆����5n��,�S�M�ydrTvw �7\)��X���*�c_�qi��ձ��ś�D�G���}�k�w�fЕ�}���4DĪ��N��Q D�8� �N���f�Υ�P$]zs�JG�HZ���(>STOj~g�|;qT��p���L~d2l�Z#��\ͳu���"��Bi���@���cHF��H��
6��F����������8�-Nj�����ӫ�i޸D���-��2�GSzw1�=ǽfA+rytA��]�AC�x���'\Y
t�����وI�7{j��h�Kbߝ�:�Jɖqqz���˭��M"2z*�j�/���#a>"��J�����Gv����C BpE����+�TȍwW�j���s'�K1��^��~e�Y���r����ýeɒ�C������[ER]x�	���r^W}3�D	�Qq�J��_���p#5�Am�w�g!�Ԯ�>Q{�����a� L��΄6
�σP����ɴtk^��7x����m�b.�Z�A˿�r$�����/�c�����.!����"����	W����6}�T1�q��Ȱ5�@ A��4�Ȗ��Y�G0�G}�u�� O��4�=0���>�d��&���s�;��U�y�-�/[�΁ϲ^F�yJ��<�z&��Ҙ�,vF���W���,`���xf�<�(sd2�e�y�C���M�B(�$.-����BKq��Q�Ɇ�'��$��giR���~��Q*}Δ�M��1q�3H��h��P���c��(��"Rv���2�� �'bJ�s���}I,�Š�F���+���vn!�/�byK'�Y?��.�_�b(��.����a�	a�1�S��m]��w^���+��1�j��m��[G� ڟ�WF�i�s�d�\���3�ǎ�Q54yNހ�z{76N^�sg{w�!�O|�]�ZA��^LF��Y�F��S|ىX����.����@e���$��\���\k�SM��u~���@oej�ˏۚ��V��߁N~z�dkBf%�:o��
���W(�G@t]�쐗J6x7 ������xwE ��#�]���;�\���j;��&�z��*�zm���|H�%Q�ߑie���Jt�G{����5��f=|G ��<+��o1�t� ��`�i`�M��ОH����,��>AL_��*�f2���@�@����r$fľ�SHNn��6�̃g�^�;=i����Q�z��!@i�A)�d���\�!�d��]j�Q:g[��]X����D�@;{&X�z���]o����-��Fm��	�Tx��ogF$Ͽ��Ś�q-�GE����
a!�������jH�=N.#J�����C�b�����@kvC]��Lt�h�V"��n����*��y�d�ѢX�X��yȡJ�֏)ʡ�Y{���k�V��JPZl�I�W���pL�'�b���_��5紾=�	���ݵ�gBV'U)�_�,��"��x�� Cu�]	C._ b���wn�-.��YJL�8���Il�����ɸ�������
eBr0���,���X`r�k��k�ɔO��~gcA0,z�n��2,ӃcRft���VQ&Ё�Ϋr�M=��	�����(n���68p,T���4�~��Q��{�\����Ī���m��G�Z����9)��n�[}T�3UfnC5a��(�E̵\e��,L�=���Uɩ����t.='y ���NR0��`eW�C_{/�s�e�Y�4�1]����'*��k: ��
6[����x�և��lG�u���}GE1�j̖/���'׈�?r ��$�w:87ڟ�yO<[�ߩ=�(M��4&��e��Ia�r�~�$ "�W��7H��'%�y�(7�O4)C!<��8%b����	fYr�U go��P��p�ɇ�MQ�Hp2�Fm��x��%8����XM,�Y����f5�_/SX�P��<5d�U�E�Gmx?�ɚ��z�u�,����$����]$kk���Q�H?f<��P��i�ܒ�Y����Y6��rD�%���|�wÕ�ݢ�p꤭q���ܫK9�/���n$��@&AB�`/Ut���i���=�&���:�0Tӣ-�������"�pWU�s�p�̛���ɭ!w�A��Ky)��T쵾j�=Y�a\Y�e���=��&gE���K}�٧~̦�b�׃�N��r}ٲrZM��=l*�R�듥��7.� ��WA���ᗋW0�b���2�؟1O'�A^W��$�\AX���/r&JE!)�B�A���qa!D�K��k�'��o���O��z�ӛ۰c�1j`,�5��`���׍����&^GN�k���iT���_X����hi	e+W������_(��#�uS$�s'>i���[�7J-�n�_/��G�8����M�ke�K��y��*|��I�˶r��%x�F<
 2b��*����J�M&/]!%�I��2���������D֡;���]��$м*�t!��Ϡ������u�v_��A�A@�]�Xdxrf:�2ε~�Xx�a}Vz�kϞbŉ��<����SYΗt@�c�`�:��#��e'��jHg��w��Slj)`Y�����R<Z��a��	�V�=�f(6+�yFU}��qL9/���o��ꅪa��I��i��Ym������S��܄+�,>�*����G���L�jЂe�����j�/gЇ\�l1��J%!2a�VpGW?��ϓ՚���#V�4zv4^9��@��_K����֗�r��֔G�ܬ�t6~eh`*c�b��­�^ķ��wd}�_1�r
��'�$�ˀ��M��C���T�Z̏��%=2GT��,��^��Bu�с1�&{1��ufI$v�T������+Z]�Bu5���*�=VIrw`p�h곀r*�1�[S�~j(:�[���s%V9V��\�b�kC7�i���>%jB�� �?"N�@�|�ߢ� 5`Qy�F�\\�G�������5��J3��~
?.w��ǬG��=������ԍJ��vq���5�Π���]HI��������2!���ߺ�����<�J���wRn�������wix�m�x����ZP{�1�ί<���Z�HA��]sON����|l�� �ڧ;;���e������a��Bd87m:���NU~T��ǘ��L`b�������</�J3�\T`����2H,���6��hC@���9�Bm��>���nIV���dH�@���K�N��-�y
g��7�viQ�6�µ����o'���I!�d�l�Ť�>(l� �vJ�X��S6�DߊB�\r!��yM�P��,D���[�a�6[ x9>��>������[Թ�Q\���i�����Q;��¨�SP��.蚿z��T�a_�*Y(�＀�K��������,!`��}����C-��N�
�Tq�t�D�!�~�,�/:��-3���#~�#_A6r��P���A�.|�RnR�x����R���B��@�-�ewRȸw`M�LB�����ixr��&d��M�^����+�sĤ����[�S�p`�c��1�OVCi�fd��H��ӫ
���t���gp%q�8����Rq��̈[ԡ����>�لq�^��:�+���Q�p�m��ìg,`~�G��a������J�iA�A��}����U�2�6E��Q�۞k�UX�$�#�sS�jHF�D̍�x�O�I��,D�N��w�Hi�t��!�v�n
_SMJ��މ�ږ����dW;���Z��I�hk"5Մ�˛H�Կdi<*=^C2j�nʋM�\����x��C'�w�(Փ�!9Z_䑟cġ�D8�I�F+Y8M*paٿ�U��:��]���5n���FQ�uO̴�1KVY��ܵwTn��i����Ǐ��|����8A�+5`r�c��x�dX��\��o�O��?R��L�}��S���+��'�n��m4u�A*��a���9c�	9�I0XlzZ�Q& Xy�¦�c��O�z���%w^m�$r1�'����ny�����=��g�d��fE�F���Z�un�����+̪҃��͊��*𲠯�uE�D(�I�Ө�OaZ��9��̚)���7��ƫ�.��u`����z��{}D�qE$�$O�	�N)����t�\l7x��k�&���^y2�4�ﻒ~�i���0��,��ur�M�q	6����H+�"��/�p i����#�z���0]y��c��������>���;�fXok��p��J젤��Kk���"����+)Խ�N��=����B�Z��¦� Cj����Y^�����Ry<�����f����5U�7��v�s�&X�H�̓�aZݥ���t�\w�9Z:y�3�)��PM��UH�ޢ���/���-�;�؎�>�6ʻ��T�ok-���rVm�ߏ(���}Q�¤$��_;LR\��RR��l���p#�R�u�U�)d���a�d��[��q�u�8��q����Ӭ��n�?�lGd0�:��ts0��s���Ƨd���[C=6���U��y��a�8�`�$3r�C��lDz������ [��mհ9S��^��C�CZ���y1��w���y��^�� ���4�"L�;��1Q�v�+v8棼s��zf��� ���LeS�X��`J*y��4x"#0l�]��b�3�'�\��э���D�R��������}|����f+����u��s9��<� B��V��ҰZۢ�������������fv�"P��L���g$#�WE�hy�N!@������SPޅ3yv�O�%�~I<�ATݚ�M,y��[���i8�nen�5t���T��0-K����[�s�n@�]f�3i��Ji2|O��q�6�ܩ����Bs]n�	`�����(�bI��h�ʾE�eunC+�dQ��ݓM�ѭ���g�N��I3�DfS0�8�C�%�a�C�G\u�s�e�dXB*��MAb�gY��B����:��$� Е�X��{'65���j{Rw.!���JK�}Nci�.�8��P���At<X7>܀)p��6�h��W���#����'���<�u@�V��!Й�3�=q�L�a>��N�<��/���@�O5�$h$���\�ABn>< �/{/)�R�D��;1p�=�%!x��ᎆro���!�#�'x�9	Q���}��8?\f�x6�NT�S��ß���o`��z�����HE������5CJ��nx���n�.2s5�{�������P�dw����՟d�a�#Ob�g�b?�����5ubl�J��1�Ը������>fOR� ���b���}� �6����k�ls!fx8�Y�̪DZjd��%�*ʧ�7�Ţu"�OYx2]�S@[+��H=T����� [��̿`d+Jَ��룘�W���m��1S�%�aθ������PK��4�N�	'�ʐ�h�����D�ȹQ�R�UKt�W)�r��ś
Q�s���C۹�:Z��r�}9�>�Q  4��kЎf*��x9s�ͅ���5ƪ*�c1/ӳ�eCg���!$��CX�YJ������;bT�๐�V26�K�@���M�{��k�f�$�mI�#B��C^� ���L��Y�[�e��&�K�:G�&�����4�Ϩ�s#8pC�Ȃ��)�����A&0j��D��
f�Q����F�cJ���f+�|���#9�̬L�䵱i'Gs3�M���l���ޔB�AK�"Ӎ@�4|�E�I�H���8V��]�Gٗ1���������ɠ��-5��00(��jF�zZ�%m#ݓ0�� ����H�$8Y]U��6xK��ȴ;���e1�{�	�7p�BڔR�H�e��=��]��w
MX�L_��GSL�$�4�4���X9.&����Mڧ�2�����yq�<O���ʜ�w��tr��7�~�u�a� �͡�3��2�bJ�]�EJ⚋��a�����Hsw��4�����zQ�-���۳����p�.�C틗g�&/_���p�PEO������K���_b{ 1��:=)�@�v��[��v0�W
�
m
]U�p�S�����qE	�?&�I>)B��@���Jy@������h�z ��?�;O��?��Q��
&�T��ݢuR)�4�HN����2� Ɂ�jnH�%�ԟ���Sl��dƠ��x{n7�j�I���<�_�E�T0���
�\�ɟ��5�#�8���.�]�2/|uAe޻.��H�D��?����4n�g�`����6�i��Cjwn�iw�n��x2���,`a$[O��7*"W�bC;��17�������K�_Q����!�������!��UV�bP��@�`��5�����&�@N'QWx��W�V#Z���&����f����6���>�bO���tV�#jX�un�$�=�jj-�@j��R��k��c��wZ�a,u|�U��Lb/o��Y5I�.�g��)���sCi�{���҃J��LM���fN#��d�<��(+���b N�y>�HE3$��~ˣ�5F����P�����Y���Z���$��B��D�Հ��4Xej�t�PS��SX�5�P��7��B3�G��P���=L������|G�ku�����wR�h�3�D���Q�-�<�O_�;���CoH!svO�u������i�aPsԭ�	VCV���W��	C֭�ĳ,\�����E�2��b����p����Y��XV�ڎ0m�#�}�C0T{�6cpF���T�n潉Y�L��JG��
�T�cî����x�;Ą����o������g�*���r���0IW�'�f���22��~�6"^i�ו�tX��W�bM��
������X��4�\�qY��5F�%�v7թ	q:����T/��6��3bi��!��A�9!�#`�$KSį�'��~�,�#��]S�Z�O����X <��k�������Z�g�ĽX��ɡ�bi�X��Y���i�0_`(�+�Lē�/���C��Q���Kp�@z�G�8)W��\���a�ɶ�qBQF�re��2Jh)��bS=O�#���-0����@>h����1=���S�!�>?����"j�	������ks�C�S9���t��8M���'��Zw6@ÄTT2��}w`�*z��i�	�%�u��>�7��_A��
�W�jX�Ħ������1YaLG?\��5�rt�L��Q�`����	qW#zg�d��P����Z=��,T��GW�n�U���c�]�.0�6�+<Զ���N�k-"
��nI��j��/$KJV�t�?�B����UǏ��7�:�bѫy�p�ub�M��4�78�b�Od�(�J�4i-n������Xo�+?. $	g4��1j��q��o&Y����q�Ӯ� ��Qq�����!Ha�:m,s����(�͇8kLΐ��j�E	+�S�˙~!Ds\��.ޯ|��G6�	l��{�G#�+��N��k���1��cg�u��J�C�^�T��xS��-]UE�!l<~�y��v�֮����a�aQp$���u&���lN��[�����;C�z�z���c��.s7��1�ib%�x�c����E[��CO,���\�_��b5jqs�)�}}�>�ش��UǳC��1�Y�Mb��|v�R�ݙ��N�4����N[�T��f'߀�?mlG����v��z������:Lh�8�h�3霧W_��P�w��a
l18�h����|��shA) 4��n	d�8L��i��@L� N��MRT�Z5���R��������ޅ�}:�p�
bZ����6���ڑX���S�:�~���ܭ7[�O<!�)1�t����x���l�)�^���+��t���L�����m(����ih�eȲ�R԰J.Zs���h]%��/�<s�_&-�%��$�	b:C��>��6�y�=5��8׉����n�p�%��q+��������\�H)�������}�����I��Q���+RN����J.���x�h�RE���Oo�jH��R�N�]����|�q`I%b��r�/��q���0��q8���Q�c�<�#7���'��;m�,k¥Ѿ������{�9�9��]
1^I�A1���\�C�Y�����n)��4���S%����Q-�Lb|�hW��4� �x�xSt��)��`Q�X�]:?��А�^�Sc�?�S�PF. �Kb�}�H�U�	������{������$s�[>��w�s`�x�E�_Gt�A���$�y��'��xYM��)z�����wk�,N"6Y������r�2ѧ���{EQ],hP��o����h�p�x�	�8��#�������"���o���� ��uF��,ψ�t�4����~bB)]����a���_غ>��<M����� ��0��.�kLVTv�3`~�Ag�J3mt���l$"&��c��"��-P����^ۜ�;���/
�ȉV�tl��������y�U��x�%|ΓbxP�-���ź��,"�WjӅƷ��/��p��Q���/.�W����'�U����ΐ,A��}��Ps����U�vN���$�a���ݲ�������Ax��Q�0.���<�e4_fuO������Zp�_"ٵ�_AG�SC$�W~�cYP�]�@� �����@�緿R��h?�=ɒ|����F�!��C��!g6^���u­c�r�n��4V�44"�ˤ"_ߢ��)G�Wd�:D_�rEZK��ғ ~"�^�(WӬ(�>>�Ms�F����O:�h�[�箓�P��X�hx��.�	�0M䷐gf]6UY�BN�� )��4B#�4rW���t���0"N�	�DR�X����\~�N����\��l*��d��|��˴������6NojFK�G�җ25NsL��/����Jn�9f�G���4�y�~s���.N7�=�|	�:��3Go��������T���x�C�v.2P"�Qp���U,�h�.`�d�%��SWQ1!����.[-���C��=_1��B��Wa �����Ԥ��p��*s<�9���>���>E�,��B����{0��gS�����RaA!̲��G�S��<T/G%R���b��/��dw�m��	|CXe�Z	���@������/��P�?~�����/�����P���>8.I�pԺ�M�
v�v" e%=� Z-��ҖMn���Kt5P�V~MY_���tFM�Ƙ�4�VŦd9�%�^�<w��,W���Qˠ}�VϰƚB�8�:�}y�Ɨ x鉉�� ���^Ñ�	���Nz��b�!��k� �?�u��"��0ۗ�^��Ƭ�
�*�Be����N�N�X�>�mc��SX��G`~��fv��k�1tt�"z��=�\L�vx���=V"������P����v\�/���Ö���&��J�p�@�~"�Z�¯A�y����#���vڠ�Y 7�*,P�۫�J�N��~DJ�t��3�i{���1e�G���?r��-V����2�r?��Ħ��+B�o}��CjBf��.8��ڒy���X+u=I��ݮ�E�S7�H�ܷFm�*v��hʥ�R6@��8��V�s������ }��<����V��)� �ȧIt��I��k����?�t�q՛K�ʦ3	}�v�Ns���1PƋ��k,<��RU���hi	|\��*ʆn��5	�Ԓ�-�U�Be(|�Wy����$�kEg����>짾>Ӽ�,���WҘ�N��:����^��;�ڍWc���:hJN���m�~Xz��x�H�5��e����Jy�~�R�4��Ҁb��q2���������BT���DW����Ԋh��2{հ>�a�	��������oL�h�-g����2��=��<�ci\׽o�?mC:s�~�ep��#<B�\l��3���X��+��Q�{����ݤ�Qo�OR2L���u�\6��t�ڑ=.��H\�_G�2��/:���Չ
��yG��0���Dcm�����1o᡼^v��z6̞3��G9����^�f�wmN�H�f?�avE0��G,�o� G�e���8>���g�Z=E�\��(V]�m>Ĥ�u�h��eBl��Z��w�p�Z��@zr�Ε�3n�.�)�}2�SP�ɱ"Ӎ�R��-D��f͠���77��1ضV��Z�ؙT�G�Y`�9�S<}��P�R�;\[̜��B��r�/Sc�G���~�s�/T/M1ki�E5o����g��E��{f%�����0)�7���������G�z��&���]��^�	������Z����H����<��Krz��CC�(��bW[N��x.[0i��{����M�L��?;�/�'��34�f?.c �i	P>���ÿ߭�(m�@\U`�YCd�#�p�?�J���>W�g,�S��?\X6CFK�{��3Y��
�y�@�Z�c�ӟRs��`%XE3�����`�@:��gH�%�p)u�	�؂S�F�7L�Q��t��=���k�m4�/�j�U����k��y�|��/҆'�icN"���YoX��y/F��h	g�á�o����a���*c���2�p��JU�:�,:Nk���ݧ��(U���ܲL�'���di�L\����%�T�&�٫�5�,@8A7յ	L}��*sd�?�]�7g��ϴJ�jq"�f+�?��XR�#������~ka7Ϛ�MI�|~@I<�<�
��*tn��\E�6=Q��K�y�q����g$[���y�wLMo�r>u�s��27:�c�ä��ߎ�-�S�y��,Y�a�m�?��� �Q�&�?>�� �ɕ.�IcVA�>xyl�97�O��,`�F����܁�r���ܙ�o�S�U��-�S�D����Ą*����J�>�͓��==�u���^X/,�UOF�t�`§_9\���t�
g�A���0
 sK=�J��V�)M,u�7v��	3�%�]:�����!���/�Y�5��VBL��w�xS�
: v�>@�|߭4��!`��c��,"���������#5�B�8^�X*?��[���ť��Y>�7�͓�)r�+#T�Z�.l<]����^0��PZ��!� HK��W.�~O?�H�$�!P�2���.a���.M�9=gV�9%�ď|�Z�L-�Ţf��*����toף%U�՘^jXa�Ey%�D"�̱2����x����XH�䚧�qU���D��4W��o7��H�;�����n���+"4�@�΋:���b�he�2�v����T�G�S᫭���C5螩���~ב�mU.�X�h53ï��U��pZ��8��(�A�W ���s�3�p�=�Uf���vd��*JVa�ԏ@�f�0�ofI�$f��y]\�@\�ع1T�lơk��7Y�	�K����	ƞ�4�HU-f�0ہ�P���Ph�	XR�|��E�z(A�ee�}循���c9�t)��(SRE7�8&@�Td��(b����0��Ɵ)�(4,1���s	D�8�y�[�w^�������d�VfX�Y�69�C�X�������3�VM��������7W���C�,����֢)f��񴊛s ��w��-��Cp쟜���:#�]l�=c�Y��o�b�1�4恨E�0�K��q��
³}�I�Dֱ+ɚ-b����u$m9p>��mc�t�\u�f�/���e�5�I����'���X�j����3���&Xj:��V���I��v"��m��'ߘ4�Az��>��x����f��~g�pv�5f�U�ͦiY�#�U"���Fp��Oqi��4��F��ȃlp|)�V��Cv�b�}�����o���jc9�Xhp�0��Rc7��m-=��zJa��1�(�{#s���:��2P��Sw��Pw�oG[a[h��_�L#=}�ub�&\�oD8 rt�_}����ݟ$��WD��c� �O�K��a�2H��H	S����=.���Hd��ި�TMf���<��;�a�R,MeЙ��ҧ*���g�_+?�����Ȋ�5oϘ���F�5�Xj�
�HI�9���<08�����ZOX�7��d#*�z� l:��V;�.a�V�.6����=Vq���IFq;>����
~$�m7 h��j�X���=�{�G�#�>]��8Ɨ&�x�4W-�����wμ���!AԌ�la"riT�I�l̻���'����)�����h"a�|0��ʩ�A�M-��*�_<�t��Eƌ�=>�<���T���c�d�F��Z�Jp�����
Y3�$��E�߫Tʡ2D��PDPܴ��ǃz2�Cс��$}&N�A�{5_	���y��q�/~U��8���F�dGE���.SRƖ�w�0�z�av����&�Y�eHDg���=8z��`��RX�vA���祇 9������4��ͧ<��;�t��0���(�Ky��� ���U
�%�op��W+MOn;R��-���a�t��N��KDo�m�� 7k�gX���͏�F,����[u�@��Aݰ�A�Ǽ���.�Ԏx�Z�xL"�ת�픤�7��ul/ ���C��ݝW�-��r3ە%��K0mⅈ�ڎ�����p��5<���E���~~I]^3�c`<L���~|-m�����$�Vg71q�;����+��<)jT"��'|��C����E� ���Zy�9MwE���	�ו^��fwQ.�&qʓ��Cer���N��(ھ��ߡ{s�Ń�1�$�c�Z)~�S�㣻���bP�}4�B�B�8T��;��fE�����J7�<��*1T���qR#+c�1w����Z�Ğ67��X��x 2F���$��".��s~�l� ���c7�`��>��7�F8o@_��6��'ވ �P��މ�/��z�c��p�$F��g����9�#o�V��F\l�1�s7b;|��_	W�%�Il���8c\��9c�f*�4G�eՍH4��L4�v"
@�v˨��G��]�p��=�^?ĸ�j��h0�X�8V�uE�r���V�z��8c�}�,?~ʹ ��	!��J�?^l��U�)�++���IEӺ��i�D��c��������$c��v���>�|BL�pp��m=�ȖQ�04�J�Њ�f+�抭�Xq.��+E���#+5�j=��y)@�bs�lRo��8͠�Iu�]ۮUv���˓��Dm��u�C��)ԩQ꺍�s�8���O܁��wδCB�	�٪ϝr]9;�H�ER��O�]���������w����@��#��^N ��s�">�ڗ��@'����*��&o�6n�����WeL�#0�R����hJ$���WHsR?�In�	I"	I�/�Y�]�`��>������c��`�,���A�Ʃ�˂W�W'�(~.~�a*b6R����Xruٱ+OA5N���-9��8�f�!�2���Ä�_����Q(Wc#7H��o�	�}��q~��T���������K�cM�hЎ=�уF��9L�f����μ�v����0��u���~����zl�S�*[��KY7^��Fu/K�L�x4�X��䲼y��	{�j 2a�ў�O�2�Zҗ�묤��2|[{�⃮�|i���Н���b�j���O�!^�r70�98����d
�aNӯ9��S[\8hI@*��H�����be.�)�C�"�B�<G8x�Tk� �p�R�H�c�N��2>�&R�o��io5�.�	a�9�t*�P��t�T�W�r�Ң��y�p�$p�A�LE� �Q�[���T��2! 	���4|��v��a�]��6��k*���5���L�+�z2����Z�뱆@�h2ԡ/�H����jIr����\�Lx��h2�7C��}��_�T�l�ӓc&��^��� �>'����6U������oBo�#�6S'=
��)�[��Z�,�ta�D�Jm����~ڰ��g���]���IF;��Iч]B�̛1�SQ��~M�x�hΪU|I� ��b���;�-3����|O���tq�m���.D�FBِ��t�Y`��!�>FN� �as���y��q�=���!�hY$���-�Pq�\*Ǿ������@���U/e� ���kt�"i�
r��F�P�>���j�z	�ĸ���>�ˢ������aQES��|��,�����Gݥ�(� �-�_���B����g���̟��q~�mX:Σ�������Ud�{��=��'�K��_40/�(%���ӔQ�3��|�$e���m �V�ਲ��홴�H��_�&�� d�r�����Z�4��v}D|'��ݔ)<
�&����ܯ~��Q :zH�t�6��'�{�CI�q<��TL�z�wh*o���K�k�^]'.%�N����b��X�+���U*��>S*�:�K��0K���h�M��
 �����xu�&�Hw�L��_�z���������r�7ҵ兓���I즆�3��A�����V1��s�_����ok�4���/R��^HA�[�����fҿ!��M�p~����K;U�25�Hʺ$7���ƊߦJ&�*w2N�1��lS�O�;d�?�ԭx�t�<iy)���
�F�%���BQ;_A�|��b;��"�e���Ì!6�"�R.�|܉'7�<E�u8!lr[Q�<��O5�M��M+��1��O�����R����(敚�&u�K߲�Sp�	W�y����������R/��3���&�<�6!�����2����>���e O�rB��������ǜO��;�$5�.�k�l;o��(m������zf�n���΋Q��Jkr���9���{~�;��:X�nD�QZ$?
9!��/���#۞�y��}�~����^�OZ�J"ھ�@��d��.c�{J��������R��\.��E��އ�IR5@7� Б�Nd]�X��v��\T�,�'3^�aـTG��F��M�̸S�v��ީ0�a,("3I�1�*̙�T�)�x�h�B��}�=��m݉�W�+k������ ��1�>l��(�W)�lȴ!�S�!��)iQp�l�K�q:�E��u&t��~F�����\3�((F�X�F��*b�%Y$sV�&����]�.�Ʈ���>�INU��9#	.�*�z+<*�v�G0�E2��'P{�h`@S�$ϳ$p�T᜶΂��`��)=a��C淾nL;Ȱ�����H<��,�� ��?�N;S�(��=�b����r5i���놔����#�j����F�jn,U]6�_�V�=�����W���Ī�=�����/��#���zg^�nJ���\�[���S��#Pf���&�ؘL� �A9�H�e<}��W	-���3����yp;��kG���L�J�:"��w3��B�A�t%��4VX�8e�3vU(�^C�!6�p
}V2'��i�}(�qٷ���O4�L��N[00d�l��Ҹ1��b�Z!�X�х[�����������j9j5��يBK��XA����d���j	U~F|0$��ѱ�|�|#ٽ�6�yn����N��(���d���7%hI��kEY��r�:�d�sn0*cC���&�-� ­4_��Ɲy�$Ml.��&Ƴ���8(�QvE�ty�1��_������`y�A}�RZ�N����,�%��"f��>N ������$�8�[<��9�+@@Q�x\�spט��/Uj�*�,R�~a���$�%}�O�ahڒ�K�����fz��/hgț�����8��B�b�p�� Oj+�,�<
 ���Ɔ������\-a"�����y۰�߰�5���^6�|f��q=˞f[4"��-
���#\s	%#_�%u���7�U`��@D7��g����x�	�aO���OA<��Gm�O��J:��s�ռ��׫�X���~�L��!{�Çrc{G��"8b�`��������q���M����3���Э�+`��>٪����g��	��K�g������3{mI�����7	A�H��*�C�!Ժ�`��q2Znt{Hגz6B�w
��s5j�����H�ţz?�H�l����,�d��<
Ca������4L������V?t�i����8x��N�&w��yTo��L��o5�����R�4VWD��C�;ڗR��G����V��\���{b0L#L��	�wq��}�Ϫ���fQ�$kh̵n���r�c�D�z�Y�����M$�zd����E!2I�x�S���M�W�22��� �M���R�ڰwn�[1 f!��k;�X!Tr�H"��L8�I;<� ��(v8�h2��|_Q�&�)���qC�J>zJ�*l��j������l�1,�V�'g�jS.�LֈsBB����e>�g�$�B�mҕ�ܤG�k�����g��O���-�mP��w�z� ;�B�U����iaj�p���������#�3̱����V�6P�U{���,*�mGi���%�$�}2f��s@���8a;���?�3N �'��]���8&��ĳ��<���&�ԩ����gñ͕�t'鬒U	����MR�����,9�*�����@�5���?�4G�a>���x�!Fm[_26�s���������M�8��	+�'"��唉1��8�Ȍ�Y��k��T�#H��"�����H���x�sc J��S���Plތ�g
v�Fm
���ىn$m�k�;)�+(��;�3]�
YȪ�OW���
k-��|w\ixq�.=%Ű�������^{�����	�sx:�Bƍ�DJ|��q�q(u�7�e%=��{�M����|��'���<䴫��_t��� �o�))�9n�<SCmBe��H�_��k�;ub�O�JB?�	�o. ؏wܫ���kUQzgC�t��)�+�W�Y6����I��rM{CP'­`!3r�\� !�K�jx��S��`6M3
�릁V�Ǽ�� `�@[ڕZ����M}���?�yZ�x/�p�
�������Ih�z�&�O�XO��qAw�t�	�k����Y�F=Ǩ�"�[B�4ܝ
���TVz��qQ��N�mDZ~�g�n~���IN���90j�����F;�Q�Ø0�.iM��>�����&ÏO8��"��G��I�&Ϳ���j��ց9�'��q��a����&�"2�5���񬍫0�.�/9��z2���B�_��j��ύ;at�{��,>�moPu%-�3�a�u�k��_��uW�"����.�'����/��N1�ĐQ�]U&G�,f|JQ����lC� }�`<	�s]/ ��|�뵋9}���H���8&o�g�"�Ǝ�M�_ݿ��F�9K�q>����&HX��=M��D��~�_��;s��9����VXD�p?�C�j2:�V�T�³���r�\�SfQ��,6$d"9��J�s8])T��N� v9R�5�#1����@� b����C�B���9?cl��s,c���4,D�gc��Q�z,x��?��\�	,d�[B�Gӂ�{�7��4��*7���,���߭,���)8c��������]��'�#\�k��:ې}�� J��W��#�I3����ɫ��۲�?S	�� �B��� �o)�m�yc쐢�3jY)Jn:yir�,4�-���//��8�)Â����4���|$yx=
�Uc?��q�وy���,��먙�oгK4H�T�.Z&ο~��R.�^��z9��h�׉�u�Ӱ��E7�QK� �		��Y��^�g���� ��  �ͻ��(��t�у?���1��X���m��cz%(!
\'�Q����<��5��N��p�X���g���O�0���y��e�xz˿�J�@W)X��l�nzf�̼!i�/�s�d����
�%����6 "�:$�TT�ܛ�!�!�K!m$F��SN��'��Z��sJOS��|��В@���G�@��@�U=;=�
ncZJ���"P��LH\]#��y���G�xf}J��S�Z��ݸ�EW�)A�t��s2ck/�&�q?�ٛ��m�O�Ro܋Ѹ�������ƭ',zl�]/$)䎜��"������Qȅ;�̭V����Pc ��u���l���vA�k{�F�ҍaRjK�H�h��}m>7Cj�.\�ZjQi]�g��[�cG�s�YVf������=�x��3ѓ�������`��rb�38%�����|��-�w�X%���X�ٗX�sg�\؟��� ���`ۼ��$���vY\*���R�9E��fO����]s'*6�\�e�=AЁ&&��{"��,��^�Q{�X�nӼ��F7�������������d�Rw�B���2H�h�K��}�1Nq	����X������}�¦0�|���z/?�U1!C��~�oZ��X��݆h���Pt�r!��q>��tx� �p��S��s���K5�����q$�>��}?��w�DU��<|x1H�{�9��Kmܔ��i�)a��Z���Y�jP��"Y�2 ��F�/��]�<���~5��7��� �P�Ⱥ6��8��������v�·S!-)b��;������4�ɕX��#Vb�_zz����w4"�-,�}�A	�KXZo)*%3j��eS��P���C4a��}]�Ѓ�BJazA�c��R�_�qQ�˝~�y�����wcT��Y�9C�t����di��r�4���F�J2\+���O�t��Ţ/�K�&�"��bB1�-ln��H�5�s�q!j�B��L%��i"�v;���RX��)|�2U�5�/a�f�,�-��y��y`��(vf�gt���������d����|�K�*�#	�Pu�QN�V�gO��M�ՠ���1Ү;�r~8�NsAګ�l���lpu���1��L^F:�P�>�;�]៚��y�(K��(�-	������Y��;�}��Bs.�0\v�|��̎Oa��Չ�;yV���j?ΰ�h��1���T�Z�����r�<)|�p�!��%�����YZ����?�m�uE��r�����g��,�=mR�au�l���ku� �d\O��;y��8��J�5�Z{��G�N�
]���cE��7{�FI ����ʜ��z��ōqdx� ��Y?�rth�'��<!�R-��k����ތ%��"߬�0��9�ʣX��ߧ��TYf�#Iۈt�>�Za3'�� -���F]Ә³��m7/װ��|E�+Uy�ɔ��G�š�4*Sۂ`l�[b��շ��u���Ĝ�R��_�$�>��yAT�#$��{�t@NbPj��Ga�x�8��U��3��Z���a�2˫�Xezn�Sh���bq 0~��d�J`���h���^{h��c�k2�균��~.�S�6�75{FP��F�?�.�؅^[��y��+���F�J�_��_ݏ��Pt��1L�.<|��C�R��.�4Bۺ����@i���;!D�d�j�.�v��se��6����vyS�s`r&�g�?T*6���ʽ�o�H샓��ĴПE{��16�6^�h��G��F�k�����<��v)��m��\���{'���uT�~�\�g���\D�,���;�WHt"*&q�煐e�(�eh��L��=I�=a�B�X2�A���g��r6�7P1~*��F
=�o������q����`ɩ��b�$������U=�}.�y�Y%��L��ʡ0>���4��C�A�~!_O�ػdZ˟R+����R?v�7����Zx	����`4ׯw���m����Xt�Z��/�ATxa#7�D�JC�����/f�\��>��
�u�M�0G�&ʳ@�0p���oq��E�R�#K"���c6zp)�Q�`��mz��=
'��C�y,�CX�|i������`�WC��c':�NE��(�B�=C��2�o8s��|+<h�oR��J���O|��M�����Y�ݡ�$'�Z�"�`�$]g0>�-.�pȥ�T���w;cC~�S	r������N��@r���́�WH#�1�~aIZO�T��(m��B�qx��=X�B�y�`�/��b�܃�E�Z��bm���� �{�<�W���v��bLƉ`�P���',�*��-�f����+[���w�C41G��n����e�r�V8H	�#>�ל����V��ދ��C�a�x?.f{�y!wu�#�]�qPK;F±��
�r�wi�MNU��k�$�
D���[b��
3��#s�?�� z�
�gp�8�Ns�U�ҏi�h������Ѽ��֣��u�rPU���/}z�����z�V9A҄�;��l�B�%�h�x��6ś[�����l�D��AI�U."�zL��"%"�Ud:h�����D0K�_P�B⡫��� ��~*�~�*���t�̲u�w��|����}ti'G���ރ&��y�8���w�D3D�Ŏ���E����=i�����|�L�}���8�IY$�1nĠx�ݱ��� ��9rsf��W����XŖ��×I�D�ӊ�i�&�4IR}@K���g!/΂��*�x����%|፵�2���j���vP��u��19)��/���-4�9I��D�>>��b�S�^BA�JY�[@g�1Kg�[�P�������X?��>��5P(BX_��u�ćTbh�������x�U���ըΕ�"7T��^�9R6I�1!���^�|��ω����$�	ho���4�*Ҫ�QkU��wKUЇxh5y[�_�Sɗ��(�/Æ@w���b�4�e!0�)j(�BVc(�a���2!�r�l�� ��,���ޓʵ&t��EE�Z_�����(X�4,mr?��Tj����I�Z֗H	|TI�n�&�Pw�Zґ�݉.�%��]��A�"H{\�&�D���r�J8�4����K�A�"�:.�����Q���y��Z��;�7F��u�s��h�r�lQ�� Z �Y�y�	�j�FɁ���oS��Sq
 �TzE��'c<{r���O�I�u�e��F��V�AI�Da3�[e~f��-���%�@�y�hz�� �����.�@�ś��~J;%M����f��z}���}Y���-��	S���W�s�-s��%��SQ�!�*?Fͩ���;�Ĥ��,,y����/R2�L�� �3i^�2M���i���?�ׄ*د�4Е#Bu�;�TK�|�Ut X�����9�F���B����R46pYS����ż$��#/e;(�˗�|���I�ӂz����S�o�j�OOT��d����.%�Oi�|��(��j<���R��?i�CXĭ�>�4��٘8t����	�k� ��1�Bj�?
�Y�PbP	�}4~/���������M����ܒ�)�㠜	��x�MT��aS�1�pz:�}�@�e�#<
�DE�H�u	�/��u������}2(O�%<5�e�-yd�<Q�?&5�7gcl_dD��;eum��ַ?h�^_３¬4H� t[!e�}hz�5J{ޜM�vp�V?�:�hId?(A��,�YS�ݏ>���a��Ch2Bq�9b׹g��9ȟ���q�(�lm�#g#!�7~�)���g߳�����9As��.�]����/jW�8����$D}g���B��.0o3g!d9��H�k7mGR��N�+��P�я
3�LV��~<���	�~qKb�#��M�/Q��5YF;�s��n���z��Ġ$�I���XTcg��N����tg���Y�GL�+�KR��XxC����C�d���"\���HF�Op���2�����?f���7_�%~�^V��_(��2
�f�/L]��ӜL�Kc��C�܇s'U�XЄB��_߶E�[�2��lW�\�ެ�S��_�F����f�q!�ҢT���F�͙�<B�J4o8��q�/�1ޒsI�n���7�y"�s�e'�|���O �*�*1��:���"j���5��pr\���1͹B��s�WQs-UH1��2�,otn? �W�w_����at��;�ȕN�I��`ʮJ$'���`c����u�@O�H�߀M�j�I �0vB0���k��o� 7����O����)�� ��~���v��G'	��;:��Y��~��Ao�p���I:�'��S1X�~��#�gX8�=�T=Wt,�p,cVںG��`�h4b`�5l���!�[#�J ��a���U�\�~��|�G�����2�Ѽ%��"���������;�/��I� �s�t��Kx��,(��ͦK��y��	��.���7+���ꅊgkM�"!���_���#��r�ݔ�*	���.Sv@�K��� _D)�{�8�沨�q�f:�8E*�篽9 F����ꖇ�Pͭ��u~�"+@��S���^6�Y7~��ϧ+W9�<<>xomzb��i�U���?^"X�Ly_Tc��@��o����G�e¦�r1�Y~Fo��T��Xs	���z�h??)�|pj���M�Y��/3�6W�z�s��E@��֕�����dc�M��=��М�3A�i9���s��Tu�zN.�ż	����2��F�>�z߆�Rm��ʛŨ��f�	�ti��\x��9V�7�v�j��J2i� u6����Vg'���t���^�)^o|�����0�s0����h$Ksm
���h<��
������o���e��Z�줼d1� `(�RYh�[�$�=Q���/�_�d�!xsPz�����?uߑ�{�n��mA��
 �J�$(��fM=���y�*档23�P'�[�i�١��x*?�cf�Oɸd?��u�uo	��/P�����wx���G�Y�¨���_������8�G7KZ�=UW�B�3��^�OӭL�ە�5�u�E��縥|v�-�����	m�֘)JD'���8�N��gľ�F�(��q��~Y'��Ě�
C"�s��Y�מ)��kp���}���$��yW&�i
Z��.Խ��k�c��-�ϧJ�s��������s�E�j� ��}��(���w��'���k�ޙ�t�kF�p:�y��E� �57Ӫ5	P�>���e�}��'}X��4���z(����b-���l�s��ý��a����&�#�GI~�2+4	���ˏ�F���\u+��@�?�%f/ت�
����l����"�Db�[(��9��6�?B5���yS�=����}雉E"��VE1T���d*~lP$�FU��|���{��_._��-#���g��w~���t�yPz��'%�s.�AA2Ҫx�����۴��Q��	�X������0�ύD��<eR�
Tf��7ĵ2�UK�4G������)�C����Z��E!��W����PQn�˞o�H�i�9��9��s�,���ܢOgF�(�)/S)f��#��H��.���o�y��b.��P��/ýZ(W��v��Ǧ)O��E�T֘j�{mm�+�
,+G+o����fHC�L��R���>�wP3�$z�H����e:B��c����DH���|������c�W��"�b�Z�""��j��������C3��Bu�B!F�P���G�6�������ӻrvW흞s����tx慇�z�n�'���+-��Ӓ�B�����6!+�@u�ڋ[C�S�]N�ޮl�������<t�;y���?��, Җ�l��q%ț.6�f�9L7W�:��*�� �x=;K`U7�R�#���hE�{�x:�5�(E���G`��j��~*��D�;�̘�)Q~��v�Y�֓J�^nk���R�9�w����9r�K�yb�t�#P���7R�P����:N�5s'Zʙ� Ժ�=a^}�Ilf�VG�VF�cC_��s��g�_Q��KB��0�}c�������m����g��9�a���C���%ؑyN񞵒FFS\��s5^=(��l�����y�įY�[� �c	{9��v1�Pjlڃxi��%|�b������0_TY��;U�JX��Y_V��-��٬��j),n�&� �L���Q�n%����!���>���?v��W���o3��ú����\�
�o���tTg@�JWfNK�n:k���������¿��D���4c�|Vy+b���_O��w�畁�%Yv>�-N&��hl��`ӑ�KM���mrp� [)߄t�)�V[An_Ue�V��%�'��"��2:Mz��@���k!ul�ʿ�3�  �via�b��=�ʃ�/yV/����������?H�z��D����S��z���"��z`+Ce�(�UEʻ���߭S}�6�w�����$@u��ȴ�!3l�e�{�{�_^G���Ns��]6�`}(�(}��+#�8�PS=�Rr!P*P���"��w�Č�8�U�����eG��D��rtt�2х��4*�?w� 74��x�Χڠ�ęb��4���d����ͥd��u�c���ޠ&~ �|���@�I��D��/��V.�u1� ����3ҿ��:�(V��	��J��4!]N�)/�-������h3����"�z+b��(O{X�<��Ѥ�0���t� �ܡ������ng(�Yֺ3�1T��4e낤��Ed�Km<7���#��M&�U�dJ�s
������,Ͽ���R,�r/K��D�me�n4gA�F�2�O��d05,:�*�7(��/�	C��EQþ�ɴnCg'|T՛������偈Н�V}����Q
Q*ߛ�IW�U/���ۿ^9��(�/�{4YFh���8�0�/3�듍��$��`�i�P�͑rIS�B����U��Tb=��V`"���P#[�J[3s�ق�E��HL���,�+j[<���݃R*_�#�6�����M	���Ć��UlIq�����6���d:�����I�Y�'a��l������F�j�/���� ߵO�A�Qϖq�+ԩ��^ɰ���[Л=���nTXU!>5�6�k�_U�8�~��B^zȃ	���������; ���o�wa�x�%Z�%C9�}���
f钮9gvZyg����YX�9�����1�ƞx �� qq�(3��6���mT���`Ė�a��>]��7��9�IV�Z'�01�5v�G5%�a�4��`5a�	�����x��������'N������,q�{3�<_Ơ������W�6:���gvl��+AlE�J~���PgN���������gu��{.�9i �WNE�L륭hbVsB��'B�ڌޜ���ݢ]�WTZ���)1<e3��*�T*�=�.��u}t���u���'�6Je��������Bh��U������U6�s�b����Acl��'K-�^�T��&^E�\o��a��}���/�:�Ӫ��PNɞ�:�ye�N�I ?yD��|�����@��*,�,� �v���=�NY�#��Jol�$���~��=k1��'�S��y����	�1�S{r�9?�)� �[��t�a�E�l�C�2����4��y��|�]r%�����q�^����8CLl78��D���Cn���x�*.���<��"G�؄�R	 �����fLO��i��E��E6�����QT%=z&���t�jh�>ՠ-��Jı�/�hZ�'l)�J�kBޣ��y*��Pu�j[4#�T`?�Z���=l�>0��f?u�?�h̷�b�=��� �w������҆���
S����$�8�dy[d<���=�񴨺���̩��y��,�}�sd'٤<wľ\o	�N.�0(r�h�>����9���B0���COn�'��c]w�	C�
8�ɣ��`�>�H�^&�����5�;-D�W���)z��_V���{�;�`�>жTa5S55�D��(�����I*7*�鉺D�a��A�tS��R�W�6He�W���5�?��Kדq.\���6��be�z��-^:GR�@1Wl���;�b��\/����(���� o�2b����hޜl��짆�FL'�.[�D��[Ǣs+���A��|�KShXq�Pr'��� r�S��E_gG��o����~�"��|KFx��P�v��x��b�d���^�we�er�T[^L��}lp'��m���A
.(�U��N6p`��߿��p�c3Q�:����Cu�f������A"�M����s�5�M�¢��E�|5��<(o�O��(�u����-��Nv�Q�/�ވ͆�uS���Lh��)m&p��*<'r��z��E7���#5~k8w�%<��J�=�֫?��V\H���N�;R޲��} �ɒ��Q����T:|QB�5�ԉ���u5c	���˚�y2��FD!ē"y�T��EJn�Yl#��~�Wo�Ɍ�OWЦ�r4c���ٷ�p��x�E���m˘L��7����4�.҇W��?�qj�,�A|�'�B�%�1_|L�>���=��U��&�\it'�My�b�_&Q�����sH oG(xмq6BjP;5<<�O�� uPB��NPB���Xќ\�~��?A��\q9/Ssr�zn�Ie��B��ĭ}f�k���T�/ZC=������M��SH�/y��3�R�[%����YJ�*1�n�%��1^�k8�E*`� �+�I)���2�Em�5��B>���Ժ�k����J�])���.��gOޔ�f�2����Y�Q���;�s&�t�}��b)�[��"̉Dį��Ԟ��T�FU�0 �4�ʎ�E���9\�%���&<f[Y�i�G�{�[�hd11ҳ�����谠��^�o�b�IW`^��mګNw�f)�9$7�(\H垟���K�n�/��6�l��#`N�oVw�ޏ���@.�M�M�.҂�@������+Hf=�A��su*c��bB�.�]ϐ�����4n�E,Q˨:�mkA1#�`%$�Q֣/�)��b//&v�gگy�|��5)3���!�T���G�^�q/�8�����_j�1Ug��}-��g¶:�0�C�&:J�iވ9�jsU��O�}�h	�Zo�Uԡ$&���,�������0}v�cc���4�1�,q
���5�[���F�r���G.ج~>i���F<�=W��ԫ��Z�l�0!�E�*W��L�9,է/m�������Q��K&z�{+f�����Ǉ	��ޤ�+CcQ�:C@3�a���洧�n����>��~z�m�>�Л6��CoA�F]�8�8&.ޝ:F&��}ؚ(�!����h��f����6�y�gC�UH��{�@y���g�<�tՃ�w1뒣$��}�d�αk+;��8��������t���QZXAj�"�;�N�b�?����"=R9����SG���x���eC N�J��Nq6������@ּ祸Srw����gy���)j�9L��>,�ʬ�@���5xȠ�^(N��>���)��. �d�`(%��'�>k�b�V��kJ�mЍ���=��8��$��j�$@��S��-x��]��aw�Ma��(�	@N�"�^m�H'�)��fٯJ/��F�cK�opu��o{�K�r�8*�>�t_M�ػ�<��nz��A8a����s��1e9!�����-�Cw�	�a��Yy	i�Ss���I�޶�7C���S�'%�hY|�v,C�t$˱����v�}�]���B�9�a�`�Vc����oƑe"���W���?8N�v��[���-p:$l������œX����3��o�ն4�maN���y>]�?O�|u��L����/�A�R�����L�!��(�����F4��p	��Z9�ՙ�6E-3��ߋځ���6zi�.C-3Qq��o�;4���w��p��-��ym@t��Z���8)q��J[�@�)��+0�!�US�f쯂����I��_� u"XN�۴�UB�3�ۇa�0���)�F�G4�#��v�A� ��d�Lދ⦛�����}q(G' jR,3Н�g$Y�t��� �OR���I�K�g�L�'��~�!Σ��kg��i�D�ͽR%X��.�`b���s���g���Rݣ���-/�h�OŤ�Ҕ��҆�Þ����`��xSU;zBxAi�M��������.U��bi�b��;g��{r�X�۠�8I�H�2!��r8�U�r�'�6=�3+����6��� +XM�~�!��|����ņ�y��Z��	.�UG&��ae�4���ѸG60)G禁���$��	s/�-uA�;g�5^}s���.͍�B(#ɢL�:��#阵�\�F���]U˷��ЬO�7@�2&j�|A�w2eܐ���w �����d)L��=��|mu�ܐ��sꂫ�d�Klk��k�6�t�箣��$g:~IqZ�O.ҁbUy�O$��S��zs�=堄�ͯ�Vn�7��U@��I',;-��J��s�w�->��YddP�Ba͑j9[-_��&���[	���{9���7����C�kם�;d�J"K�rOC��'�f�}s���?L���.0��vE�cT���~\����%slM,�|pgy��˖ט%v��8��C�Rܯ �E��Ҡ�)Y���5�� b����N�%j{d��z%�=�G�<��Aa��� `E ����*M�*	��-@� Ylvgl�sF+zF$�m��!#P���e��,Y�5R�$+K;�!����y;����v�|�WU�-��,qJ7X�Hj�I�--�1K�S�\x9�3�'���1��'���#��>�)s��58��&'�;ӝ(hF�C���*�����aF�q�2T�i�~Ī�����[N^��Tj�e�)���s�0�P�$�����@�໷a�Tb����鳉��_�AW��S�-U=Kp^j_��P'���@�+0���{џ�O4�V��7�2b�jv@g�y�&��Phg[�:^��'�@�yY���̯����h�[H��JdI�N�n��������B��_����J�OWK�ѷe[�7q>�0b�$������hJ$~Нv��k�*&Sb���ՀlYqVҲSKs�����ъ�+��ӏ�{�����Bs�@Z�q(��T��G��3�)/��$o��\��F,�	9Y&"5��"9w����j���W��v�j��v��3ə�)��&�m����cXT�{� ��Ug7$�;̓��0�r�s�X[6��s	�\�u��x$�� ��C�>��o��U(� ���5pJ�����v�0�9��a�&"�zb��a��|;z=yX����_t�%)��&N��=�e�S.�����Zf�9���6A��R�� �9H���]����3�@�Pq)d���udd�x'WB�+�w��l��u����"/>"\f�]8��4��|��ؕ�� �"an0*&���e���:3\��;>�1B�9���q�z�cUE]���6��f�L�s������%��	$�dn�D����K;���j��΃�vy	o��\��q������R����T�C�<��Pquie��:��r�3�Z qRܮ��)��p�qq/�� ��ٶ���a���u'�A-R2��;"����C���.=�o%0���/���� Y�,L����E��|��)�Z�N;Q:h;�,�%��l@z!��{+�k2��������]�'�ҋ�wD��؛��U��.;j�~ݯ�9���c�f�I�´����
������|�u!�C	��w�6�r8�ɛ���KJ��ٸd/�֋8D5�~���ZO�E�7r��Q�W��|j�Q!�=H�&����1��&C'oL$��
�P�F�>/R����$��<?��=�a�p���^7�q�f��]<7 F�-��ǟrЕG�SH���x��'C�(�MΝE�1NVt_�`����dZ���v�\܊��T$��#_�)C�X��%�T~?D_�ՙ�ӳ<䠋X����������3��aj��j�-�����_L{��G�����Ư�i�#N&*����Rݭ)��t�e��lnwrE��h>7�t}<���l�����v��`w���>>�}���]��&N*�aͰVs��S�g��."��[���_-]��*�HG����%�h�d�0�*��$:?4���lŬ�ֳ���'�������ѱQ.�E%�?�D��#���A���w��q�,k���q�� }�Yy;�c�\1;GxOg���c�nnt�ħ#�X�d���'4���S�G͒٠�RF�!����~�&S���~��xs�/���!�Į��8�H!QG���>�U��#�����)��)Z]�1�Q��o&.����y�6y:x'^^�oLrl�cU<���ŭ��"�{�<v�ڟ@ [}�=d��.QP�Wz8��]��g�(hv>�1�:3� sr��k���rm�RO?#O>�8Cx� ǝ&3��<��af�}Z@G�7T��*��g�2�0���<��,N��}%�W4���-D�?;��0�w�g�a��[���P���hl�j&^c%U�V�E�8�r���LX�nkB8}!�+�k9q+=q%�s�����Xq}�W)[��mL�d�tbk���lJ�סK��B{�vʮP��e�@٢���mHC¡.ڭ+�nf-�s�X��CBғ@�F){�n�x�ǟ�֌��4Ik�~ ��~8�P�tA���ޑ�7���,��M���k9��P#K^�Ͽ��s����N���VE��8��[�)v|�\T�ر��K����'"�P�����(q���ɹ��r�:ݞ���3fL!�]�꽫a��N�e^?Y�T�hg��`v��}���2�7�Յ���f���V
7ؼ(�� Vu�ȭT�{t�A~����Om�Ճg薽��gH�����U�v�"mu�KC�#v�.����׶��2�U�L�(5��>����</D��n62�3&t/�D��\�(���ݴ����ː��qw��`�y�"�w���Hz�8��~�:�_e�I�a�w�YHt=R$���7��Tz�V5�@ ݡ]�Rhm'��I��EʕltX����3��'�vF��Q"�B�/na`�9���N�^^��X[t~���rO:��C�leM�I����w��hS��?tGJģ�y���<�̛m���ߒ�<�nL;c��_	B�Γ#�6�(@�>��3�H����h:����z"a2�[����ls^��+�"���2v�Ŋ��v�a�'�i����j���,�F�����w�����PS����j�]�e�NA{^(8#�+���퍫�{���~rpu���W��X1\��z�2W���gk�nt|����(3)\��Z�귢C�gө�;���Ս����%W��[j_ 7j�=fU��h]��O~���V�����9T��4�E�^�~u;�t�6�!-�J2�Θ��wG�瘻�
��,<Ў�|���X�����쯋͈�)��k�H��c��֪d��z2���n���C� (�EP	z���U����j� ���N���.F^"��d�Ӱ��gA$�����l��Qg®׼R
 ט����F����C_HZ�ߏ�<�6��GdgL��W�*ڂ����?D+��*�^=W�.���l-9�9�I6�J���5@2���!t�����YC���!RB��-��8o��SH`K�@RjX��
?�%��)]�������DQ?d�B�Vv��uU���Q����w�J�A͍�{��@٢��裒P��)�26h|�0����>��U �	$��_VC�MN�%]��h =�]C�ݛ;n�Ig�02�*̆ˋ�ȷ�;��ۺ��~2����b}�]n4� UK񧃉�ZJ�B~��"��}�}������1~p+�K��t��e��d!,�%<�Z,3��U�8�	�tI�^6�v����c���E��R�f���۴����X�G�da��2R�4ƵH�϶W(��D���E�ZN2�S��ȼlż.������MC�**���]J��da�.�y	��xQ�
�z��+��	i�wG�fi_f�0��qTr�7a�]�G�TF���x�:��s_�N���/f�5��<�����4h��s[���ʔ��f�H� �T5�����!�^�}�ߘ땈�H��ö��"����ѩۤ��OX��t9 ��lӱ`T��%�� %L]ԡ��"�-��M�PjK�ˉJ`�
 ���p�Q�����l���+M�)�$��EVKc�[܋�~1�<�Y8Y�F���J
��#�'�y1���z}����[9����>��p���[��*��ՌM,��I����%��`�Czr�<;[6�cd^oVQ�F �f��!��u(wC���(L/�/ֆ���Pʉ�?�o����-�nC�UA���m�M��͗l��E6��CZ�C�@���b��?l�M�@��Y��m]����3N��fM�����J�h�'�5%
A ��|��/�����+���$�A3��n,�s����U�e�f�B��߸S>�3�$�㯤�sM4�׷h�XҾ��_b) 6���7�)*%Mm1��b�.����=Ȓ?�`��}`���hd���I>c�R���t��U��CS�7��!{(���1�Ѭ�H��)��� GFt!ÖK-lǨ_�
Z��������#���;��U���!��ܒ�Ys���G�Mȋ`T��(Q&S>�';Ke6�pD�"=���.��v$�~۝�/����v�������BɿY숹L���G�h�G.i��TZS�����`I��V?׈+�	,{a�p��?�~��Z�g:c��fC�H,����k�x��V������`M �aZ���q���I> ������i��*��"P�B�O�E8~��p�Y���f^7�	P�6ϫ�v�mu����+����>K.Ay���X�����+������z�����R�G�kЗ�b������<�@�CǗ" �f���6�U����X5BPNC�YCQs�`H�����B�6�C�tP���kMNf��P�1~z�eL�܃��G�Z%
�h�r�S�=2�ĸ��#g�:��ۗ\"-F+�3Ĩ�ƺkU���(G�����4�8hx]��Զ��lW2&&<r�~���B#0����?y�c�gWHo�E<��/�c�N�Ak5����]��)���2��=g;-��SF��7"����}٬\0s�1��S!S�H�g���R��?S
��g��M����p��wFO�t�E��s{~{�5[A,	2!Xu�/.��֢-k�Q�{�r���@���$ҵ�! � J:�=��.�/�L��]�{T� ��C5��f����k���4�~��yR�ٱ�d �>���>��{5�,#���ڡ�Z�֚M��;4޽�l�L)�M�/�q�2n���9Ls��F�N���"����K���.c+�Xy��m�s:|>��!-��3��?�:,g/m�2�8��D��}� ��ԭ����l�T9���H���"x����Y��0���0M��F�q�+w�����I >5�"=}!NȠl�SY��).��ǆ��t�	�5c���":O%oDv�ڇ�ƚ������Z]�Z&��� =�[��ܩJ�*��v>�u�itE��R<��-�j�`2�MƄ������kd~�V�Nt�9>]��+U�0�{L�ϊ`ʍ�,H���'���?DH�0ǵ�2�)TȏK������~>A�3$��t#���w�ʾWl,ۻ��@k�L�y@��*�f&$<P����(���b��n�?��@�i��'����$�����"���H�	�}K��݂-��P[O�_�Z�{�	��>�f�EA�v�lƷڦ���5�'�",��>o�~W�����;���8�}L�����b�r0rR=x'�KC*:o���8��V*��pYp����zX.O�2`���J��lc+2`D��˴s����:Q�L�F��@ҧ͎�n���-�a㉨&��l�/M�Bu�lvo|	�?��)ZF�����a� ݓ/]�XHTN�&蟣���_�.�&E���//���#JaM[J0�숭a�Wy��_Mu�Y_�����X�e�r�Z�U}������ϼ�h���қ���<te!�:oK4�2l����J�� ?��s�=)�ek���(|��|Ԥ,�STC���FJ�� �,�\�0Ɠ����}~?�/�^�>a���T�km*�"�8Ǿ��e�����M��
_�<"�5��D�}�Ȣ<��8�{��ͥy.�,�;G�d�����'tn�+��\86�E�
��<�yI���J���	����̷���Dn���9��5����ET�,��潧0l�/�J�Z�$Lj�	��vޝE�3�w�= 5����G��x���sb�W7C_?���( ���Op����4��'nD���2/���?���6������QN���_P��P@ļa���h^YE��V�߹n�}���`:������
���������f~�m�l�oX�\9���j3]%�@N��D�IF��:q����@͏��XZ��0:b����`Za���@}rm`�L0r���E&�(&{�>�+�Ӥ:��+˸��i�"��?�����-�z�ǶH�H��&��F�cVU�������@,j=��oqw)H����u]~<��7׫�q�EP����A��]}6�6$5���'X��ɳ���>6	V�+O2�Fp'��L+>�ba��k����� ��~P�������TW���Q�7�∲�*�#�
�7@��N%uo�;��Z0���3����.QC���Ƈ��B2���[�� pJ��������V�o=ph��}��hS��_�>Q�0�i:ԅ���X,���ꠍ�}q�Q�jT�N-`9��"�F�_]��UA�w�J(�ɛ�����u�ي�K1�Tw:����1X�%A�}��I9��K�8�?A)��[�9"�����㊑~���˿g$�;LT�~]�����l���
�sx�#L���\�2i��Tsײ�8��ғ�d�[��| J�'A�oa�1��uۘ` ��@�:h�6Q:����<`G9�K��Dɡ�{=ɫ�wn�n��G��m]��}nv%�=oy����� r�����t���o�׉7Hc:F��I9?
�=�*��������sb�iW�N� �I�5&F��6�S�R��s�l�%���t��Y�.�|���aCӤ�Uː�(Ǥ1���ms��s�9k�l�1����|�?���׉���Y�!��$3�o��Xl�4�9Ã��P^�CȮg�\��� ��9�f�lt��0�Bj�j�[�1'u����3�������u_���bD�e���'��ҏ'��	�J����I�<������Us#Ab5<����>;V�^\�^��g�OQ'l��tEa��9�bkkϣ症�j	Kdr ��ؿ�~���> i�Z�J�-�f'�8������W֮H@��ĮE��E�
����l��}��L�S£� g'56�Kk�:j�� X����I�������(WE�4��~�m�j���H�m�;6��v)!��ΐ���Rk�9�/��뫫�at�ͫ��ԘGXkQ2i"E,�=`Ք�^�vZ�fxO=iN�i��*�/-r֕���#M��]����\�W�6f�Ւ�-h?��L�QZn�w�����lr�3�.�ǁ�i��J�Y��|�C���.�l�J
ZI'&��4\�$�a|O?���(H���7W{NP8�ُ�7У��c���ζtjCi��:��e�;[���I��`�/�Ȝ�\��x_���7Ƙ�s�<X���U|yn�.'qJ�¨ ��,��1��Ò�j�f3��=[���R>���U�l�M]�~g�1�+�!�)�GA6�o;���@���
K?��#];�2�X�����ŐZ�E$ai!���!��*�?M��pG�*���v״�<s�S󴦌����.7����Z�4k���X�jk<�w���v�5xvS���(X�!{E��y� ����#�%h�C�Zr��䝛��}��E�dUI�nԄ-��6��'���Ը'L3�F�Ԭ%�������������	�?KH�^!0�0M�)���&����]�g x�k|�8q�F��%���!�i�9��K��kY��Ǡ~� ���W�P�]��px);y�-�WB��~���.G9���}ؓ_�L�ݬ*m�	z�&����&i/��ަp_��,�����A��$Nx�VD���"�lݗ�ѝ���pMz�
��i����)cGp�6�B��}�7~�M+'���23� ͕��J����x�cLl�U�� `O��7�*!��WM�.T�<��d$��V'\��tQPF���ծ�iHk��$ ��kh;":j�zus�\<����	9�|��rے��s��i`���� >&�*;(�n���o!��w������YW���9�;i��r��RBr�%��y��a�Hl�� ��Z(Л��K.x6ErK$�.U���xKA�ᵩ���4��� sf�L@&�yC����hK��N�'r��T�gă�Y��W/4�[���
F'����_b�]�颒�p�7��~�1��	F(�-��ʏ�&�'�ޒp��m�~�m*քH�x� ddf�������\e,�3��VZJd-F3�/n���Ҭ�UU*(n��ָ	7'jI#0��p�9�F/i_�����h�J��H�7���0R�<��bhi���d>�{^O���J#��H�p[�c��XJj�7P!3�<а��gb��6�,�-o��d�y��rZ��9 7^��͇X6)¨�[V4L��P\˭�d�28�yp�+�~Gj�4�EG`�K�fJ��(3�aK'��k8�V��߱)q�p���oR�-�dE���|9��J ��(�9q��`�6Y�i��9�$�n$�=�_�KX�$��p,<@J��y�F9d���cԎ0��sс0HUϐ��l7�]�u� ��VZI _k=�� �d`�U�/�2�?[�B�ܯ"Q���Q_�cʗ쌿&2PE�7�/�j��(�Ih�S�6�� sC�/�.F���(�_�Wj���Ԗ*EIXp Xvv��~������
�H�';2bS�ɰ$i��G`v	���^hI��w��c����s9_B�<RTR��N�	�_^��� ��(��l ?�����j|�I^�x���0�qf4^��"�DϺ[�gꢏ%m�=�lr���و=�`Ro��?b�,�*�r��X���+���<mN�t$J�K"��!��"ϥ�	��EH8�; ~ ��>�����sL���:��^)+\���#�w�a6�QE�Y)�C��]#$��Rd0�z@�Ĩ����W���Ǣ��c�P�݂}|7�'=}��S���T�S�ky�ݖ�(Q��$$7v{fM�v*?0hqc�`�<���L�ͽ��@���˘K�C����{�ۙq_���;My�9���C��V�;s�z���F�))�>I�����#��f6ܻ�� `_�K�W+-�,4��}8���Z�����|�Yqsi�-^.�16������1�I�����7�*3�e�m�r��<��iH]�+�q���~�����d]���� ����/Q�I�\6���;�����.3^�<��@�=�0fȞFf[7\�N䜘4y,
�;�`�\!j��͌B�\���<}�}g�
��k�F�S��ej���+Z~hV�Մ|xB˳~�J5x�Q����'�Ι��W����ר�5�.����P�OD/�ȉ�~sBw���4gJ�v�=�Y���߰�=X	�`<��H�L�ۏՈ%o7W�W�~W&w��������-�+	actZ�qc��m6��iLSV�*���)�-4���UA񏶌*.w ��D��i���Z��R�T��69�
-�D�s�C�]n\a��r�ZpU�0��j%b���~�:���+}���3$�Yͱ�F����U{�+�k�{�1J�r����OVZ~F��Q���I��/�X��p�qc#���A�¸������̷�){���60�F��B�%#\�S��8/X6����6Fޔ}Y�g9J���+�-�K
�nu��A��8�i��Ӑ�kn�`��EҚ�Be�)5�UE>�<5'_	�ˎ��e�"��Sd��z{�Ԝ��Y{C��3ێ��b�C����.zݵP&[�b�0W�: ����0��l����@���M�dk�~-�m_=!K��{�~���O��s�l<�5�]J�^�n�⣝�L�G&��hE�hs8��s�����h�����8��a@a�=މ��%����z|9��n�}�jsg����^aB���PbK=+��d�+�M���>^iW�<3�NyY��a	�U�Ɲ/ئjbG�u�b������ԟ<�V��q���2��V��kC邸�����*&�Z�f�ft�8ɒ��|̩){���x�Zn{9�Ҵ2�<���#0�_]+D�mq��
���߼!r6�1�GMKi��c����AĖ�v@�������8�*���t3��M	���T�w�� ��D? �Du��|c���j@� 3,�AA�й`�YzC�@���v�� I����
W�n R���k�pAي����eɡ+6[?�&�q�@�i���.J�M�Q�ʊMC*'+��kOxn������`�c�9���IV�x��e�Q�r��׀�����t�};��5�0S���uG�luh�����F�g��D��j��@��y�R�;]����d�	!�L��I����>S��8iV�;|�7 �SY���k/%C�o�hT�;��z�e��u�����ұ�L�W?��2�?Kh�ͻA�?2�p�� ���v�g���*�jDD���*k�?�w �������.���o%8>i-}�w�t�(;�!�������z��/ɇ[�|$܎Qs'��z|K����{��%l(��Հqg5��mw����vK䗖�>ƘB4o���3�"F����d9<��	<'Y��
����x{�\�*0�Ex�O�`��Ѓ�-Wg�����cߒ��N1�r��Q���2�b-�`G��х�����)`��.�Pv9�M���i*�D;;�:��t8ݑZ���@B�񖦖(�S���r��#Qr�W)9u����PW|�������&1]���h����wl��F6���@o=��ɯ(w�r����Κ�43�׉ċYb�i_y�Xc?�c�z�21���'˛i����֝OH�=���ߺ*3�`~s���B����!o���y�2�@ޮ�T��%�cAR�]��j�8!ϵ5{�_y��jm��u&־>�J\*e�����74��E�9ʣJ o�To'���{�N�I�%w���Ji`ra{V
D�0*��S9J1{������n,$�����z��X��nQ�uXG��J5f]�fs\����u5�{q�pN ��s�A)NE�)�nm"���oЍ���SeH�P�+����"9@���KR޻a6i����,��e-����n��F	/=S���P'�����Т��/t�����wBȰj"���V���)H�
�9W�!�R�K��f� ���V���b]��F/|s�2B4���R�[����P����U=�*�|Q�a��~�u~�/�Jf_q�e�(ʺL��U�:�R�P��
b)�KG��QZ69�s��ZK�Z����G��O;��?�c!��;�Z����R�j9�H�"#&
�xX���Η3ǭ=�S�%��dސIv�g���c��S��(�Wv�?�o��$�u	�&�T4��#�fq����RK+1r���r\�V�e�=Q�<:�}O�#s	$�?˕j�>��\������� ʇ��n�i��O98�����*}ďZ�h�[���	���YA��d�t���ݣ�[o ��oOJP�[�?�$ ���?=)$���2+����Ptjʶ�@W�?���J�	�i��w�ɴ��vt��? ��ҭ��h<ք��m�� �'�� ��w�W-ʴU�:�4�ա�*)~>�+?�*6L-(,�(�\��+��H�g!�L-��L��9��`��Z��:����G/J�i���'ݖ��p��ፏ��-�*m�S���b,�h�b�����2���H�=Pg�
��=����AJ��N�ke4$�B�7��?�a}�]T�
�P�Đ�g�h���@#6�����|3{͖�/���;q�:��1�7μx��v�>�@��QV��l.+h/�չ4�C�o��_���9`��6ɔ�gB��q� :c�U�/��R���㑩)��b�se �I�=>/<�	%��!ZQ���<� #�"����l����6j!p7	�8�b��Y���<����qȾ�ʑ�&h6�t�B��(��Y��:��v�B�m��7�쫽U�%�ɜ�V�YZ���|�!r*�����HL�Iu�>W�p�)�Ha�F��#���M�O��V�K�$�f4������E�#���#��[b
���&
�����(��A)I֪<\�Y�|�g���#���}8�1b��d���4��rH�PA/��_�R*��6�'��脠�=a,�%Y�#8�2���w[��oݠ�VA���+o�hi��m��&�)fwt�]t�l�?��]�eͮ�8f�BH�%�j�i�=���p`'���R�at��R��&iˉ�j74me�Ew@}�[��^|]���[�ie�9�1��%OOx�ߕ����@��e�xg#��LӴ��Ȇ�����c��3Հ�����V˭�ɱ��lō���6�N��2��U!~>͟�Kb���nMU�<�X_=���K1�p�A�����������>jѴ-�#A߫�I�S
��E��w��3)���e/+�t����B�g9K�pV��4Y��bY�#�1�-Ғͯ�o�˛�*����u�#�ְ$l�n�����Z@5���뇡��vL���5�:Eƙ�������H�6-B�\��Ig��&[P�A�G�l�E�?K>���&fHH^���8�`z!��u�@-$�E�n���]�!]��������kI�uȨ��tX`d7��ľ-�Z�N��?Y­\/�x���
b�� �8�H��e	������:1�����H�;>@�������	�QM'2�ü�BFD�VǢ�0:��Sk�:�����Py�o^Q�)H�z������*c�a�3�O{�6`����������O(�&2���U�Y6�4N�O�d	^�	�YD��V#���l.��YQ�~��{3��6�0�%l���p��&A��eeͳ�����-����|^c\��ϗ�4x;bxu��v�Mq�z2!f�}e���ϻ���Ú~,�0���c@��qz��T�F�xwK[��E�l���H%>G]���iv�d����K�E/��*��T	���caZ���Ŵ����⦓"4K�������*�d��E�|�&<@��
�Y�n6�+�y�A@$`��j(����1�D�:�F��ܬ0l�m�����Z4�q]����MPk���h�MPa�yP�4F^)���Avx���nv�3�u��P�����?��@����U�Y�-/�#�����U��Q��T{U[�j�}����p��t����>�5�GA��n&I'�?h�HC.T�2�����<��"f�E��= ��P��g�������m�^�q�+I��$�6L�v��U�0�	2�y�8�&Y��۔�~� ���hq�`jJ�w�K�y6��5 o�Ȓ*H��Y!sͻ4�l[�i�Ә>��_�y��ݮ�[�5)z§{��;�n��+�C�eFe��?��}��S_�Y��~�?�wಟFt�7��j���*Y�a2z�9EG��.��_�H@S�a�����H�9���Dx����.��|��硴o?��ʶ��ҳ��,ďX0��N�w
� k�ll�:{��J��e�U�
uT��R|��;���WW��l/3�=���uvB�����W��7^#aʧc���IO���`,��h�B��u��'DГ��ˍ�j�kl��q�n��7�)�[FX�4�B��2�Y����z�]�Pߘ&ჩ��0��������Zh�f؏��H���?�ɾ9ξ&|�� =V���1��~)�3�u<��e��$^��5�T���[���q"��H������u�n0�1��o{K2K\(��>y;N�BU��Y��?���Hj}�_}{U��3-Ü.��H9�?j��aђ�S^�B]�^���0n��|	c`��&��	�$ot�q�lY<h��� ����(zG80��g����U>aea] $�
�`����Y�uJ�8^%vAH�OԄ�o���e����)�x��=y��F�����8�� ^�L�V0�*�&�~��-b��
O�jV)�����[��N�la�s���֖jmi�i�L�E��q��CpʖSh��k|u�.��h ��u+-r��h�sܨZ2�0R�`?-��4��Q���I�^J�խ9z#�����JÎ�>�|�,	[�dWx�?N�����	��!�SY�X�?S���C��t�|$#�n8 z}d��h�/
�j�xzt�rOKa�&�c���3��O���9�1Q0h��F��@�~��,b�9<�Ѣh��7�W�T�m�Q��&�)bhL���b�u~sF�MZ�U� _/���q�"ӎ=�p�JX!枯�Ad�3��׃�&��G�Z�$��g+���*04�n�EӖ�����r{�4���0�u\Z��j�r�%ܚ�2�� ����ס��vG�9۶[���qxw7��~R|�$н� Va����l�����(Դ�1�������:����P��o&Ui_�S|�$�����7���i���m�7��v�YI9����U�]v���m��r�#V���e�p,���W���G�|&��g�����q�?Vz���A��6e�L~~����#����u�]8r�G ���g���Þ`�Q���t���>	��bB���ʍ��w��l3�&٠���7[���mY**54��_�����q��Q*�D�j�%� �/���Ǹ+WC7)
�1:<AS�~i�I�1�y�Ë�j�#�lY��~:�(Փ����o����Ţp�{��Ub���}!��KY�vT���dv�@�F�]��6j9z����9'v��.�-q�<��o��u���G4�p#�ﬆ�mQǝ���Ғnt�OL�������+��9�r>���Q���[3�@>��,���L�d����ߍj�o�ã�dA_NFF���T<�,Z^�a�C| ���9=g�eH��~bG�/-5�Ÿˢr� �!l�&�b�%4\}Q���/��c\b�e����%���<N��������4�y�Ʃl�����X�w��M�N��~{<�*#��4(�_"�%��?��%TV�� ��8��{"�R�{�'h�F��Ϗa�1&l0�Q�KPx�(�9��˫S���8�v��8ͱ��im׸}��r�i_E����
���ן�`9���Rkv�V���'U��Ǫ8�.����a��'��.wgo		�"x���,�s�fY`T��|�G��yP>P��󙩬[х��g]�R�wa� |�]g�5({V�ò7��)i��?0D/E/�UQ� ]����@c� ��>qw_}�(EjBλߟA�ԟ�b'� YG��p��Ӎ��t1�_ڼ�alϡ�kY��qcv	���}c }��d@��l�pzh�?�a���s�e\$By3r�� �ޟ`�kOf2����r��>dS�eٰp�����ok�Nl�N<�m�ƣ�E��1t�ä�7»�^�/f���vG�{��h��?o
-x��փN���0c�/��f� �j
��w&6������e�	HP,�6V8�̰}oF1�e��n�E�ʤ�a d6�V�Q��C�W<Y��)Tz����G*�H���=�wkV2���(������bx�MX��(�]�\�~#�D�n�!73#��V�Wp�Az������V�I�M0l)+�&��,f���\��k��A�g5��!�l�P��S���.?WS%;`�./�2�bY!-|o�p�z�S[\f!w�r��3���p�+
4�G�v�,VWh�H����3>ɹp��'�o�Nxq�¶����
���qc�� !��H�|�ȅKP������_ͅ /��}�Zddހ����O�
�BxY��<��O�������p����)7���U{���S��զ���H��f�@�o����@�ӄr8ն���.і���
s�UY�p�y͆͝8�K�w��Q�VQ��o����=�fgv�0�Em��	���9ٓ-%��1�dt�����͘?�L�uԬ\ϗN�A�A%���+����oL<4X4��΢�sL��E0`����!�KA����z����%�x�s"9f.Hh򰿮<���$��A��E�ȸ��2U�mv������� {�<[�Q��g"��Ym��[鲕������#\�k���cW���LK��gZGw`����%��F�� �z�w/G��Tmw��:��#s�f�:eg8þ�#�8ح���H �)��W�7��t\Z���F6}6U��mP�%Ft�G�__͆���i�V����h��S��,�/����a��<쨐�{}��R���&�<�~�Xy��/i�H��{��J��^��v��:�D)J�Ba|��슠f�?KC�h�s��o����JH;#é�%H����9�Ӟ�~�-�����X{$�c)��~H�j�;��?� �pT��eL[�t)����E���2A$_�T�����<���2���3:T�1�5b��O~d�Ls�l��%� ����'�ƨ�F%��|>''��ϑ�1 �Z�É��M�b�b��z�a�A>��t�k�7kf���m�;�R�JRa�۽A�d0)^�_�L��A�$Y}a�ˡ���_k7%{���M̟c$R���K� ]���H����SP���!����MZ*�������F;�������Su���b�^&q��e�<z:t.���ܨ�+�-{�?���$���j����}�����}��	�m�E~�v>B�Z���k�6>;#��TC'���#�5(�0r'9��-8�n������|c�ߎ�N�6�Ӱ�|jJ>����Q���my�j��������MY�K-m.�P(;�Qt����J}�l �����$Pn�p�#k����!\:�>n����ඓ`��b*yP5g�U4�?f`pn��p[�R
�C�9��W=2�c�;z�e_l D�!���$��UUA�
\���ͯGG������h^��+���JH���.��,�~��kolH*3�f!�~9��Ǹ1/�IXf���2��6M~"����F�3x���f-g����ɹ�%Y��!��V�@��7̏��o1Dp`��
+����v.8Q�@�D�r޼`���ӡ@3�6�u�J�e�ӯanGx��s�����'����;� ��gT��$���5z$U��`�s�0�����n��d�Xw���z����?���0ȡ�U�gl��OO[�v;����|��B�8�6��(��o�e&�V�t�	z�þ`VNI��D&�]�n_0ǂ=�~*n���x
ST,
��CS�R҂���i�#��%@#R�j�/��g��$�@�[��H��%�H~�������Eל���������
�`E�k���~���<��l���8�<0����u��;n��%��Є�\�k��(���]5�l�@��$�����`'��y�9�5�� LM�Ýt=�����p����az�nk�U�!`4n<�>�``�t�g��K+�35���u�&ue�]v`�7˔2`��L�RO[G��Gk�D?��#uVh3<.�������
�`��@~kޯ����N�Q�{�[�2p���U_����w�Dv� �C�3���ܺ�UY+'�����Q�# ��%`Xڮ�ancHT��O�eꅮ�jM$��|�b�KQX�� f��)0rN�Kd�]������2��;��k����֑O�-̞�V;7(�'��L���l,�>�Iz�o�$�&���y�;�ons_�]�`�y���#:ɬd
�2��¦�G��!����5";AÝ3& {m���7ǟh�8�����A�p�^igb�m+�S��j2P˰��r�\�
�H�f7�����~D��1�-1��}�"ɓG�5��q�M��vt���ש�u� h��.z���o=�N�t�f�粴k����j���U"_��rE�1̓�n�p�О�+#�>u���B�ɶ��U�@�t*V^�ܓ��3��mf�QB�⅗ߊ�O���"�7rA�G�_j9�+�B�q��a�B)�=
BmN�"��zш[O�`�v�}H!ϗ� ��.,��xҬά�{��0�n�����@����埂�G̺�h�v��=I#C�4��^XF�RKB��OU�}}H9_�������]oS�;r׸�<��eЧ��N��&��| j'T���X�C�CZ.��}�D��0�I%� ����F=k-��k����s�)�]
���R���2,ٻnT�hݞ��-��$x9��e
$O��P.W�y�[0�]�K$��"Xq�޷�#�bw�d��i��(8�$�r/��1qO!�)��T��!���6�'�qڍ����0耿�k����;3�x�~Ԅ��o~_�!}�� \���C5Bُ����ub�F�����s۵�����َ��2t`{!3uf���%:�<�)���k��yP}��48�v[���l�y��Y��&����� �Y����  ` ][����;�`=��-�u`��[C��d�G�]HTYxm�Шݑ��� �C7���P�D`��x�Pv��yE�j5vB��X��u����M`��HV����[�&�L�ԇ>��R��@)�vgK��R��:b���-t*�J����Pk_+_Q[�0��?QKD6̠p#��ޜ��n'���I\�i{a`ͣ&��^�C�GM�����
�A�%��Ή� ��n���"��N��?X�� r�#�_����oB�����	�<
ñ�~��Xt�^~��r�ֽ1#@,gv�#��d���rb,�!U�7�g/�[~��$;��SҾ9� q����wh�#��N��k�4-oX͜E~�8ВZ4�w�a��൮i�Kׇ�T�Uqɥ�s��8�)b���a�U=�򟃽���kM���k��J?��B@gMO��L(=����k$r�y:)�#n#:��w��l1Ӵ{N'?8��U�rL�S��j[�Y��0���x�i!LI�㗵��8<�ׇ{��x&O�+��/�W������5�Vb�KГ{W#`hj�q�c�"�����QW2����E#�/ U{e��9O��@M���0b�G��>��a�c�Cӱ�[3o��k��V�m?�o�&�{���:A�8�+eA"�g@�M�l���}zB��o����`��K	cv`�}>&���ѷ�@4�y b^��Z~f+P�g"�����0L�Ә��YS:��	r� R��(8���辠�j�j
�ZqJ8,���KO��j�}�v���V�X����~0D��a6��E�;�ߡ G��e��7	H�l�a]O��B��M�V�~�#E����W�1���
Z�E���&�f�-�i^��%��m:4u����|�uN��h;kS�	#�Q�wSK\��悢���;LR���!1��o�jZV�`���o!���H��J蠖�kl�P��ƺx	"'�2�E{ӵA�|d���J|ʻ�� &�;���\� zx�ʃ��/��[�~z@N(��Uа�qBTy��iN����d��nv�[1 `74#����u�Rn�(��� R�+�tȯe�%�p���~��%�Ez��<~c�
M��������ܚ��BYMt�8@��d��i�0���@��6�<������!d�6H/���%`���n�~8�8{en#&-��j����c�*�����!&�VT}������mԆ�'�è}���p��կ4����"���byӽ�����h�oúP�����7��e`������#���N43AX2ۅ��/�q��@=����'p��א���Eu�~�����8��D%�w�J߈Q����l`�e��G�zA�q�{�)����Z��H mn�u I�Wñ1TJ_������)��^�x�gk�)�ԗ�K�&��$�j_0����l�8��ބ��)��E�R������	�-Y
t=�Q�k�I��Wy���
�0��Z1�%č���S�^ }���\GE�=��թᩆju�g��o�W�����1��J�Ѯ��N<��wL�a^7�θ7g�L}4���;h:�`�Ҟ�o��mp�nEZ�+�̾E�|���s&�i_J�Ӭ�w�ފ�u*OAB�i�uӵܾ�t��NJ����<o�<Z�)*�:m�M3ȑ��J�TH7�H���5��z9?D�ʏ\i��S�
�o������(۔���^q[C�]�U�� @��I5g�쇰F�,�-���ß�f/��k.rzlP�9�F���U�SZ��}�8ؙ��>��1�s�3:�r����y��.�!�1g�����QwރP/]��1~����N�F!�xf�ؐo\��>`�x�ee���
�9� I�m4}F�����R�9G_>.�F���w����#�5q���pX�KVW.�(�I$b�t޿��ס���#�o���md"
]f��h����6;���by:����#`�a��A�뙛��1�k��i=x�N4���,?�Y��{b0'K�qH��syT&%N#OЈF�]@�*j
����#�����f���Q9�Vq#@&Xo�[�M����	��\�,7���"4�y�h�������FNP*�R��O����b�U�ef�b�5�\L��:�T�\3���_c���iI;�||��Ln�m׻�W��M����ή@v�],�U�'���������
��t�^�Z�l�Vځe>�\"R�mq�m
tfS����)�y"��&إM^�H��h�
�A�\x��m5-K�H�R�����hEeG�X?���z����sPm;�v�G9�!�D�dFX�&5*����;�~�">��u�I"�m�͔r��c���h����Ϙq�?&�*#{�;��j�r̸�A<���{D	���aɒ��c]��28�e�R�h���O �ɩ1󯥛�:zq�碟23~�i�e�����R�����x��}�۲g=���y�7h���|����	�u�?�1e��^S/M4�,���Kh�!\n���)z��Hn.O?�{�2����Vq�U��V:��	L�H$�;̗���!@�smF��q{�|�h=�)����$y��Y���1��w�?�0��.	YՖN�~�{��?CSPȪ����"5��
D劤]c�Z~�{�C����<]�O
O�U�hu�i����c�1�'d�X���ř������ &i8�P�V
��s
�����j�]$��nK1�	ʍ0N��&�����7�����K`���i��u '�����n���D����!)
�j�:��F�g�4��J���]�߳��-��E��jT���m��ɚ����9�A�X�^A�s>V��K�^��?8)fŰ�m�I�z�c�� d��/��^�͒�6����S�M��A���+Rl�`fJ�����zU�Q����f����&]�$,�Pw�ǫǱ`ɭ�ToU7��$#4dj��v^�Jde��	(K�Np���WX�ˮ�9�ǞZpgdĴ� [d܉O���.�O�k�~0e��]{��p$��iFdOA���������G��^,�%����Y:r�3ghE��_������J�d��}!G�O�Bt;g�s(��*y���^@���	#�{Q�^b�1�Y�ޏ�7�5�uj�R��v�T4�$F��wb��9[�r���uDd//��K�f��7�*�XD `Ƌҧ�/G��� o��9H�K�d��Of��+��⽒�kc������;A`�X�뗈���`�g�=Rnc"��f��Kv5��	4�Hk����[�v�=�L.���M�����sQ'Һ�]�:��Ob]�6���k��������gT8�i�*$0�)�&�('�G���s�)1�ͨzFH(� vG9
z����ǫɄK(�7g��τ|H��gv�/�2\�U��ܱC���m$�mR��B*!�^5EG�.�$+���pIdh�s��5m�˪��B��8ѥ�Q0�+;^%����nT�e�.� ^3���z���?~��}����ŀDk>�S���7�����י��-�$ڪ2W�?�4b��R�B�cv�ni��%L#|#�+�3��ӻ�x4sױ}�C����4hg���AƇ/�=n�X��:93����֎�^�;�o!�s����kU����s�"(�ZH�E.�ԖN��z�Zf�
��<��2�����{W �a�0ݺ��V��1��:+����*���;6����Ai�=��tNG�%7��h�o���A�+�S�C�����sQ.e����R`p���b*��fz�"�nw����������ǊG�}��9��<s�T����_��ejg���`���l+#}R���j�JeV����q��gq��Z+��[�C�cV�~M���G7�����Zɡ�o���Ȫ"k����}�i{P[�%��1|Γ���w���`��������w#z9��k���w�uX�f�w/yz����m��E�܆p�B��������&-���e�?jI����Pl#�K��l������?lʶ�U�;ׁb��G=���j�rⵋ�W���OF2Do�&Y�M`��E%P��ٲ���^�\G���6�3D�g)h[�S���|��E@�x�{�#�d����;���f����
���y �i]��7�+��A�Kt�[	2ZQ���7ƒ� ��F＼.r����ެ3;�e��'��y��px��1����S6�ۀ�*έJy��;O2���.�~�J�o�EW*��P�%��I�zV��T-�إ����H��׷���o8����pڴ@x<�:٢��/�"�6�����,�늁G�����܏�ĩ8$|�������/"�X@�!k8�-Ha׾��щ��Fd��L3_?zߜ)��Ӊ������`�멃�s�~�n\)C� �Y��P���"�^3�%ã*�	�}>�fXѩ�������[��\��&⧺�-d�����o�{�P�@*7*qN�X_�S�9��c�����8^�Z�'�����I.�4���c�1���+���V�T���ݶ����������|���>k;j�p�p��(Ѱ���w���p���R,�r��~m�"��)��ˆ@M\��W���Q��5���d��ڙB�Y�����+�K}����q.Tv���%���/D Ӽd����a�C�k���v
��Փ� }�m��t� ���u�/l�P)�=i�l�T��y�0��V�����
�����&����-&s;�q�w�!���p�ZyY���|�Sji,9�E�V�"/�<���΄#qYw�D�#Rl�'M˞�	�t�qH�[��de�7��5̸�H41�$/���d/&(����a6�+�!
r��jt$R8%z���0�5q�g=�1���^x�Q��]'�L �߅ȑI����4�����x�̿S�+��b���Vχ��Q��� �ͦZuyo�/�r�"��L�!TC"O��$�y�پ6�W�s��7|��	��>�|$I8������'��d=D��3��s�������;�=�٫��UfF2�W��?�g���C��p������'��%|6������<��).��Vr4ɢ�ѐ頸�3�a>�����H	t���,�=��`d�-�q]J^3@~f���J���SI��^���A�g�L�?o������aA�q^]���:�0zy��)2mN���	���4?�9ʄm��H�b�R�����B�A�<L�D$�t��5�����	�� �T{c��6�+� 
�`a�E�dѢ=��Wӹ��IK��3��'�%��CH"�mP(�1HNN�@�FR�'hn���`��*EWNQԪ��d��J:0ϭ�倮�	����k�����2�ƕ:4z�Vt��dϹ3n�R�N!�*-A���IǺ�A(��wy
���Xϻ�����_ـ��v�T@{��fم�)���ꮷo�߂�h@��XrN��<�f���'���pK�`�Ec�;�	��-��f!��Q$�.��~C���8!�Q@�4������1g9���3�����%.v,	Y���;���#���d><F���7V�M���@)��J.��� Ҧ��p�+�E7ұ̈́�Q�*7'�+-��5YU���Y$\�z�]�nF�|K
1?+}YAǠ����n������X��y<9�lJ"�Ȑ���#m����zPKV��6G�7w>���MK ��k,���J�W�{��f�,ljM�[����@�}�>%�N�M�(wW��h>�,�٩Q�=��=�"��`��h��1\K� ����X�_E�~�¾��YqܢX��N� �2�&�R���A/��q���Ûe'3�]�V��Q�����}D�t
D�ټ������kD��->���_��\��T��#�!n�J�!���ט��j������W��6gC����;B�6�l��ê2㤠>(�2L��$Kڂ�ث�>���t�Lp�M��K��i$uy���A/�}<t:-���W<�o�OΚܝu�#��`U��6໹���G;��r�:V;;%��%��c�.�1�ý1:0r�,\�-ڷ�
p�z��b�x�l�� "O�OwZS��8������ ?6�t�~\Ny�G�
e��)�4��m�@����A?P��=k�DT[D�e|�஧���\*:�y�k��f՜�|)!����f�Y���?�l�z�H����샂��l;0�!��dX�+*��̯e��4�(ЄZ�S��'P�?vۡш~U�:t�6gc�ɴ|��y��@o^�W�e�y6�����Y���<$�3��"���<���Xl�dE2��kq3{v���
�ܥ��;��1'dݐ�}�PO�B�����y�b�S�}[��Nk��@=6͌gc�^{,ƚ:��nd(���N�wCpw�$�`�'S�fd��d��(j21P�ÿ�;���B�K1�ѵ����W}�np�� ��Y��#�Y߭�P
�\�ӱ?mG���ݵZ���t�(�7Q��õ ]W4G���j/�C���KC�Ck�&8*��mD����x���];$����"��f�M�!�<mS&d��:v�C{����K�a1�����Hޜ�K�����i����@٢�I�f��N�:y�R>K�ݫ��$ᱹ@��$�d�Z�<Ev��;+wO=d��ل��n�7LX1��=�X	7i�����|,�w����-[T��I0����BF���K���(���_�B@!��=*��u�����Ȼ�ή� �$=m.��Z�V�^$���C��BP��Q|�U��,e�d(���U1N{�rJ��?��D�S~f���x�$)#_�&�j�<�ͯ�X������I��g*rwNC��N����o�����l��F`(�8�j�T3�-�	�M���4�4���."��.��)co�Kp^ޥ�i��w\ ����J1�I}̖jMR�cq��`��&L�џ
�`���v��JD�ҒyP��W,T�Ǽv�,���a��jȋxh��3�ϫ�w[�y��f�Y	����^F@[�O���.u�1:S:��7g��3*�x:�'�܂{Ĥ�K��e��,�Ѧ=��}o�=�ج�Ό�¶���}I`�,�5�p�"En���'sO�|IJ�:pQW�x���V��g\��wR4���c�P��],�ߝP�C��lo��v�S�I➞ǯ؄���b����ՠ�p��b�'I.0�������W�ۂ�/�"�������5N�`?�s�|���i��E�]��nV�T$�x�kK5�23p�tŬ�����
Z�*	���I�4��i,
f,h
♒?��%Lf�$���$`�Q�p�nx��d���|�`|��
����s}��1P�V���-䍦�q<��z��$"��/!�.�fu����&}q_0�^�5��-�'|�S��C�u�X����xʛ^��7bn�l[6^4���4W��*8t���9�yD�{e�$@v�I?=��?U��m��v��~�CϨ.a�	y\��q�Ѐ[d��ߚ�,<@�Z�j��x�vB�m�P����2�v;?ʺ�5�]&�օ �>��"��3\�������j�����ʶ긺��g��(�-�I���k�������^�fm>�@r�� 9(����(k6�f�2;���9=���5��i��q���oq�rd�_�e�3]��S�q�J=i��_�$ʟN��j�����s�P���!	෈p�v��B�Nɛ���7�A�?}C��Z��64|r8x���{�����7W�Qp�<m��	��6��u�#ڳ��ڏ,�e��":g�͎k+��|D|w�&7��6)>v,O�`\����o!m��gg����@��Z��m�7�F˦M�-
Z泅���
��r5�4}��@�=�Q������qe��ҽy-ٌv�CU�O��5�X���003�Õ\� ��X���n=��9(,f9�~�r�Պ|��8!����rjz�-�y���k��\�1���s�'8�n,��]�r�*ă���`.��Dj2I��"ժaBE��諾=p�f�G���`#W�\�/�3�:��oI��{�"^��4��FB�7��{v��#��C�������F��ݧ��N~�R�$z�݊��)dc�_������8X��������������mWl���{��+e�Y�����v]JS�z���c&a��K�nk9:�a���lm���}:��*��ҷ��B�+p�p�����vv���K9z̕��9* *�<$T:�;�<���Wv�Û�սy �n�+&���<D[��%�̸H�����Z��� ��ۢԪ5���F��wP�'���B�����v�Z���C����Q�j��G���}"�S���#��{YmZ�.���'�[�A�Ƥ���l�]Y(6uq�Y��r��1�M��$�^��J��1�^q�n�4��	�����OF!�	��T������,����u{�s~uH�z1�@�B)�`Z���El�7zu�Z��+��~�n^��m��]��0b��as>P�q7�E���w�DCA*7��q>��-vm��a�<��ׂ1�8�[ӂz	�.����|�MH��XIOy���n�=@�/������Vp�@�貐�6��	�ۛ/$'+gOtKG�}I�>H[���� �bJy��Ҏ~C�6��	�g<f����a2�Ƃ���l��޶Zk��|�&�@���D���r��t^r�����y�yـ�(p��(��Ĭ��p%�z��)xE9(�݇��J���2��1���q%·i��W}Xx�"s,��8E��O�x���du��W��ҏ~{���+�V�D��e=2���]��)j���F�����M��
��C������Z��(Cq�;:\�E�qIH���]q���p&��:_	J+jw�wi���YD��i�K0�9�R}5�5�������+tJd���Q�Vˬ�}/�0�ş*<i�r�+�u�'.�o�h��A~�ݍ��zƵ��O|a�sb�s���sc`�tq\s��Ӥ�}��4����1���'J������V�m�|C�ǫ�����L�����ҏ�h������R`б�;s�����:����}�q�N�����=� |��? �&��3�����%��̓+�#�]O{�(m�zJ��Fv r���+,���(߯��e��4$�T�)���#�<��+�����4�*.��� �k���A�AcL�u����w�^I�ܴO�A7u�}�ĭ+�I/- y��n8��?�ⷝBb�L���[�=�T�}q���K�v�a��"i
��y�_�u>TSP�J@�����2�R�Ú��bbf�yɔވ�4����d�V�l�հ Q8�n������s+4_�.��.3f��['�v�?�it�G��
]zl��pY��_�P�5*k��=e-��-��6�<�(���P�;����v��X��(@��+�!��SzZ�m�&.:zb1;�ی�>��]�u'b��7�0v�o�=Y��w��vY� �E��z+D���E�	���x��kl��a�G��L����=�����L�y`�y �N�y"�f��D~ڬ���oS<��{�G���|��bxEmx��j�'� zB7
�0�=A$�>�ERH�00�q����?���O�����#�-ھO�������'J9����1g�%f�:A|� P<�i9$}����:��p�S����S�_"�c�Z-�n�b�@�;��
TAUi*h����?�J��B���/�o�N��\l[�p"��Q��w
y;���^�n�
����ۃ{?�o��#�ϱ'Z{W��˟
9ڊrO]��[J��_*h���޿�,�q�u�=,#t��X��-8�/ŝ�ѩ�� ��cf��f�>[�*��gҪҴ�,RFJz9���Q�f���+�}���Ϟ`�z��e����ӂ���>���i�f��Z�` /�J������S��o�����Q��5[���t�����'o<�~���(��p7簄l�y�"����~��+�q����}���(�SA�큸�8{u��O\)��a�+� '*�4c�P�j���~hWQ�'1��-�ͤI�w�Y� &�Q՜�;#��a�r7t@��tݹ;bb�I�_7V֝o�Lّ.}���+m 3�0�^O��*Ě��q�vdJ��2���/���+�z�%��XO|��ў��A���YD?-��)�&nx� �oL�S2rm$�����Z�`���.ym��5�7�}|'@'��,_X=f{��fj�
�l(5�P�OMciih2�����Gb&`��+AW���N����B�}5*>q��D5�E�A��!��|�Ct& w�ޡ���84�^F�y��w�9*y��$>�v
���%gp��<*l�G��Ү�K�W�&q�S1T��R�����&�uV��(ڂ=o�~:���@F-,��
A����K+u��V(t,t��>|�D)��"����� T�R��{�u���B�pѐ��&M���w��_Բ�,>�����nG�����hl����`��KB˯C&yo7s�f(���9ޱ}�v���H�p2���?� �JM���H�`��:橪6�3� ��K7�*4R��=׽��0¬��9��G:',��搲���j3u��簓��I�����~�ڠ�a��O�tϗV}԰���_�P�Ȋ�k���X,�L�Pb�2"�|�Zf�`ޗ��K��N�"��(lp9�P��
7Uh̻
,h�$�ݨ����{v�Ók���/�,����A|�丿�0�5�1��Ha��7����l�r��~"rP�̴�S�3+�e~zc�k��5�3s�
Tnz)rDRj�|��
�I�.�(���Ot��!k�}u�ꡏꩥ;=�������"/�e�b1 G��n�KU�1;�&�����x9 �P|��6�I�xS�5����"z��4.�%�1�6�lo����dp��Z��I{���b?@qC�?]\Nu$&%𾓘\wN�Y�&м]	��U�F �:4��"C��(�8�mD6g~�(�#������$h����a r�%��j�V�?�H��v]~�V�>��4�w�')�|H�n��GT���x����n�	ߺ�ш�B���z8��h�%J�'W^r�[���@e�i�)/�EĦ�6�S�R�h/���C�>e�Π �:��Q��G�<+l+č���6��P�F3)�Y���I{�P3l���._"������;)ϩ Q�z�'��*
J�G������	�á�[PB����!�����
:��ǒJ�&�n{�� �3G���l��ӧ��=���e�03>y���1(%Hj�ŭm2����*Щ�����7�o�W��)N�\�vyK5�$��o���9CW��#;���v!���k~����,���R�����+s>q������Rq�]l�Ә����8�|{�䊡u�U��B�Ͽ��M�H����'w�<΅|��	��K�ېâ"�׃�>����~��7�I.�=��5�pS�L��.�BI�{?J���P��ƶ�+i�P����Cf �3s�D3R�^��ء�a��u��o��1s���-`�}�5�뀡�=��tZ��E�2��u��oΉ�Y�Ƅ�~����ݮ���K�����NF�Y�j�W���@�T��/\���l���[~�J]�A�'�_5�47�;)��sV�Q���f��&�n�Eb�����VqFo��5�����<кIo[�:����$�
d��E�U���8<��cޚɛ=8�E�Q;�P(/��gd 3�^PN82�C��g�Jg�y��h���j0���뻭����n�zѯ���Ȉi�2y)3��1wӃ�,����?ʍN�����e8�Œh��sl/��m�,��Xd,R]��#�qz��۷�[��řç�_��.�8կL�o�h�B+���j���\Dz�Q��T�C�+���=3��W�?ny@�:�m|M����1�q>�KL�Wr\��YjI�T~���*�'����;b��ʥ0);���d������ �"d��RZ�-�R��Ϲ��.�U��W�ؽZ�߆ƶG+��rY���X(n��:zGR5s���"���U���!1I�ZQ����6�#F]�A���q�� �4�
앪^���s'�ZWR~�������4����>�c�M)9ic�/ܪ ���~���ƴ�x�-��_t`I����흥����p4
˵�Ҥ.N��Rl���Lߌ�����d�TqL1)�N��6^��s����ʳ��֮j?K9~������%bM)����)��B��ߥ]h�ň��OL���}l�^�f8����a���{�?�kiӳl��Ğ_>Bc���6?M+��DZ�<#V?n�i)A�؉!~��l�N���rw��z[vA Min?��~�R.<�=���G���w�\
r��ğL�$��`̤��׵T�\y�Jg��zI�)8�颽���R��ل:�<��e�����*jYF������S���|�=�]φ*�w�/=�Vl+�pa�1�#Y��餄��)G�A��,�A�{������	"u|�(
���8��/L�J�]�c�}�e�Wc<�7��{���5M�W��Ď������eY�a;�yӢ�F@�C:�<^���؍��Wؽ�6%�� [�S�$��B?������.�@��}�&s+���v�$���w����d�0!��Y'�`9��M���i*{�({��ڕ����eM&�@B�6��1�z�MEG��S}+@r�l�=��z�;�ð<zf�g�5:W��~9`��2��q�ULM=��7�.ޯ`���R��.y	�^��w��"��3!+dus�ս��	���P���B���{ɞzja`q5��5	�t]�k���P&J�%>@,t�o� �Gm���O���>>s��õ?�To�4�C�\�e����]�L鲇�Jy���we@��ƕ��,lb|,������^�� ieq,�_+�c	gt����I3�1���˽��o�����rh/��Ҿ�W��>X��2�%��4od�9���2��V�=ë�tVǼ�)a��O�E��� �7uaO7�zlS�C�����*q���YO���t��X��5�Aؘ�R\��a��[ʍ��j�P>��ב]��d�w�����Q!G)ȝ�a�媍����jecX�Ǡ�}�K�a�%m*�?��J�-�5&ق�����O�瓻Y�%�{x0<����4s�yah�-4;�2�Zg��|4�0�Z4�.�Z)uV�gT+�Ȭ����ݛ� ���-���Y���i�zz/~��jI~�u[YxTZ$�GhG�q0Ζ|I���KD��)��L�O�[M�jzXp�,�%��:9X���2� �i,7ڗ���O�֓�[k� �~ݙ\�m��9ؚ�t`����tezL��ll_A�n��Fr��͎�yR�aHO�Ò��h_���2��ۈm�(�q�'(=�V��Zd����!�7�y�ǌ�7$�5�Cӯ��B���a�ʰ��悚� ����q5�+r.���1e�x���}�M�'a�a�R�Qb�m�$ 	8�PX~Sq&�곞3UEu�����3�5n`� ׁ�ZH�f�x#�/����rOSm��9aIPCTt���kzV=����;a �bf���3:�I��
��C'���;S`�ާi[�C�1��W^�����U���Z�B�T���p�Dz^��EZ
_�P���E����V12����*
I�^��G��6�uO�>��a6����v���D�-�VȺ��<#1�N��O�)E�N�(����]�^��^�cؘ�m���*�	'����������k��b'
9�mKYX5��AQ^&'�Zw�&��;7�&��\z3���9�?� ���� �a⌕���qۓ�������Zy��Y��h3��]5��o��Sb�a�&QA�kI��ud�^���_r��
��kڙ���m�y#�m)X��T��J��J���3�6��**���bP�^oyG���nC���g6#��I�V�p�5�n��$�L�b�D^�]$�|fp�;����]p�)�I���B!�)�_�?
UE}$m2��u#w����q��*ʵpA�Aˍ���I�@-�=g"�W���o�Y�z�C�CEw����4�����z��\7<��Һ�H%
W!ٽ�:�	��B��{�)"h��@I_um�JO|:C�|�v��f����>d1�����bM�	��O�=B�zh��a|%XI@�W6`R�0e W��ˑC�`A&�Is����T�w|��i�I]�BF�3s6�Mm�:�9�;����5�\�Ȼ�(� MX�:D��}6)���|��/Q�����Ϸ��q������̊�rL��z�@�1���s+r؝.��Q�WZ]3b��:��O�Ҡ�s�t�.Ŭ�h�GqGB��:�	(��(ݵ+!Vڧ��)�U��.E�?)����2��&]��<�&ا�C�ȁ��;�ð��t���R���˰r����i<����A�5@?7h�I�98�h'����~�6�H�X<v�ADR�W�C:����R5h^�E��!�tU���K�w�p��}��{p6)���
wM�SqA��	��#��]�MN*J�-Xs
��?a�>����{!#�ҷ;��/
�NMf�p�2�|j��#�qε�E	���eS�ԜJ�A��J⑥t����/��Ř�ZI��̓4�P��ɉ��XĿ�4o5(�],UI.���/������W5���y꣆ݬ��Ù�����3��v�oF$�\���a��y�b�5G�!g�e(~�}/Hz~�^����Y�Z��8���8��������)FTa�D[���x<�0B$0A&�S�Y��W����ӥ$({c�I%��%(�`�V#y/���lj��O�iW"��+f��ijt�G��p�?"T�,��X��I[Mv�&�_�+�.��0+��n��2�\D��K�y{��6��϶�΍��Bk(쥴�ĥ��"; a;�Z�_��඾�o�
�h�?pMN�f�=�{z:�v��
�A����>��m磸��Gƕ��۠���@'*�\r�����B)�6����2TH�aIh�-�7Ó���S�,�^���v��/��	�}��P�����ʷ�Rc14+|�[�T0}ޓ^��{��VZ�����R�3X�����&\�C��v�'��L�s�܉wax'�m|¸tE��[��&Ɉ�<��f��奭j0<C��{�<Wr�4~�J��N>>��B�	�y��U{��r��ܬ�x�s��5|A��@�9�L�Ā�m��o��o��K�<���*+����DG��Z/d�ƈ-�z��W�٠�.�k�x���>���ڮ����� �� 	3��zV
#C�jF���СR|���﫮��v�G�Eu�����о�{� !�H��ĳ�C:W.��nG�O�	����k!������FÍ�K"\�xHV.'� R�[�H+��]���u'�"�����M�`���>���죙��S{q��C�R{��G��e^@���R�I�(�_rſN(g�u`�?�Y_0�f��+8WZ���s�pZXj�X�Q��+9����B]v�?�Th����XM��^d�m��zϬ��3�;��Ey���" �VOk�cgǎ��v4��+���mB����9���e�]�4'x뮚�]�T��e�Jۆ��P�`p���T6�����tmw\�b ���n�x����Ӑ"b����R^��v�&.���l���q���3/ʇ��2@�<�ԫ�T����$�TN��~r%T{�ᗔ�e��-9���㇠���<��1��P�]迫�˅��['���[��<���ð�#�������;��wGZ���3�Ŀ������s�;_)Q.-$�vO���ou4�#x��{����
�T*5!��Wi�4K�2/Y���\�/���6<��K���|��e���VI�FD�U��Dm�<�t��2G��l����߭��mSrݑ Lr��!�I����g}�*�h��I�ȫ.exP�
!/+p˄��x���1�[���t�O�D�� �$O:y�����`���B��w�R	�YzL���A=�禋ټ2��`��c��Մ�����	�������Hc�-m�=?W����wX[>\E�)Pi4�b�'�=�t�}9��:5�i��4̠���4)�gGg3q?���Kd�Q��K��=��V;l��*��^̐��]�!�N"�W�SӐ�9��Dڞ_�t�臵ml�|�� ����Z�a�u��5&���i�-�G���ebu�wa��6��ǩ��ޛ7Ɏm���ok��� ^�n�Ѿ5*q�[f�A*HU<u������OB��-�j����@d0���H}���.��O�{�M�r ��/�M".aF�e�+������ϒj�&d\�U"uԋ}��:ٵs��NU���,��˵ܽ�.�:��������]S��8��ߛ_1' ��݇��K�]�����iUC��*6�7d��p���<=��+'�S��#��W�L�8���e���O��T6�f m�g�~AqCY	����Q�J�E)af� ��h�����M'���>N�½��a������!^�L���W�jպ��^ɜr�j�V��z�۞��JT����Y�>��Q,=m�ry�%&�X��/ލU���+�{��&�r�Վ��6��l�m����'�(h�`_�͈{|Pǧ��M�J���wyk���n����b���X�=b{�l~X���e3ޭ�*��
�h��^�����!>S?��F�}N޲Gf>[��r�a5���  �00;��Ӏ���q�~}���B!���Q�FW,Ya��_X�������z����=��5Ͷ�r~N7[��v���,ӄ/��d�'Ǩ!��r!��Bh����=��N��yj߅�����gt�I�Cvw	a��t�3Ì����� ԞijO{3p��f��F�$r5�"�l3�vc��'K��o�����$�G�-[,ಭ��t�;0�������@�У�l5���ȝ@�fYp�|4-�{�5���!��*b�!N�:	`�����RYje2�Jl\��:��Ϫ��p�f������:��p��>����� �7K^}X���_��h�YL,��8.���|N-`ǌ�31~Q�g��WʰU���6P�?{%�AI��d���g�g�G��.߂�U��۟/�E��h��A��uC���ꏚ-�Pn�J�:��D�ro�A��Pɵ��n�ؤJ��=N:6�[D���yy7�N}m�0ug���̐�3<�4Ւ>���x���a#A���9��OB�НG��g��������~�b>ꕓ���\��L�j�����3eW5��s�Y{�?1�5�@Yw
�+��#�F��'4+����n�#�\,��?k�H��e]4!���U�_�⷗�����_��I��*dGno˛Y�.�2}/�|E�pb�yd	C#�'9�ꊎm�(���D�Q>����s�q~�S�6!��TV�*c=�mx�ۀ/��:��$$Kp8@˻��`�tBBƱ��l��Y�ۚ{U[3_ٲAO��.G�
��1E�~�:�Ě�뒡"J�eU����{&�S�z�����	3��1~�t�z޵Q��=�݆�l�`���m�`����m*
�a��!��,����u��	b�'g:���^a���!Abe*MÅ~�����1��x�nA1[����O��P�A�i������%E<�9}�#�󳩋��-pJd���e��.gdX�sZC}��8���/�7����S���i:�QD*]!^������@�U�Ĺc����?��AG5��fr�U_QtP����)_�����^��߽"v�e�!INW�Ȑݽq�F]Q�!c���qrp{8<��ғtز���L����,�.ѰK�[�s0�`�߃x1�f�����E8�/ ��㍯kIꛡ%���N��ur� <L��=q�ǒ�h͞�C�X�Q�������v��f�P�9b�q���J��1��qy�9'���;��O�����ZNvF�b��٣�mD�ֈ��	�C_���hk��mV&p�h�gT&��$D��=GY"�g��^<7%+%�����RĠ1z�����aM�����G�h1,s2o�Ə��av�0�$Y�:�����8�:h"�qz�k۴|(�ɣ��"��ɳ��ڣfHU��?��T�K�q	��3�]ʏT�#)l_R���.�Q؍cW�I#�w/j��'��}����ۂ�'����T�l���Z�1���A0/CÛ�K��K9��~��y��I�<�)��~!T�/��d�mRNs$MjnN}�Y���<�{�Ban� ^o��P��6ʀ��J��z��A�aB8Ѱ��ʷ�sW��[�I^<���.#��C���ThO���ی��pT�q(��M�%�)�i�ev^ �u)��"*lv�8��%�y����w��7���$�&8��y��w)q�y\���8�2|ղ�b3�N�E��m®wk�&�U�Au5�'�!���oj4o�D�\ۊq���Ex�H��TrO<Q2w3�ƎM�I���ֿ�_�����:�Qz��h��"�%�*��P�TP�
:���*��s�p]�Ό��$�fL4��k\?��{&JC�w���\�
�r�	��	C��[K:,쪆Z���7.M�/�+6�bV(.�.^!�+�� :�$��o�mb	+�7#�㈜d�+�!b��m-�5��2E��&�5p��H�����֚��T=e�7�v��K��`���C�@�GQ��0|�cK�S�[j� � ╡�6������#�l@�('e�>H+���?3v��z��A�kH�##U��a D,�y~�>}u8��Zr�n/� SȻ?�����3]a�U^�ٮ)���-r�Dh�lQ�ʹIX|���l5����}Z��ʋ���e�)� �w��b �5NUF��mbW.����x#P�#gJ�k�yd���M��l=L�-�s���Ҹ]������Ɖ!�=+9����p<׆��8څ?�1|{�yp���L����W]��_��w�Ίj7*��~�X�J[�������]��� ��>���]����� 'քM% �zmjk�H����m��X�p�����NF��(q��[�!��މ�(3��(��Ri�$�֥z���]6�z��������qɳ��܇����o�FɎ }�l�[�f��H���7�l��Sl�o͸mS̴�3n=�pBl�/o|��X�{��d�&""�z"�ŲQ�.�n;�᥯Z$��i=���(�����%~��{�~T,��]��Y�3w���E�ȼ_ΠT���)g���e���8#����,ZLaQ�i'#v���u�BMV~�Q����Q�pK"o�l�<���U�+��p���y�N�9J~��+r���x�W�R�S[�6�Y�j��b��4C�7��ˬ���|�6��{x�Ic7�G��W��4[4f%�U TW�"2�-Ɖ�T���[P���9^�4u3d� ne��t����j`��si�ت�80�:����)?v�%0����0wIzBdI��J]/;�t2-�as��Gv�����3���Δ��Oi�]7ش�8���r�`��Gn��5��f���
5A�{�;c��;��G���b�h��D�-
xIm���t����5��ˁqیr�s/������s֦ۭwN�Ψ< ��4����� p��������sk%����H4�U�yL$��r=(q#�_���>�	��2���i�E�� ��;��� �-��5�vqDք���Z�eD]�ÁjuY+����w|�t�����9x�:y�m�D��o�y��@դ��y�[�.`�=�Ó�y{�ج�t�"�h�v�&�>�b��>�K�	�A%�z�*F��I��vqD�LKj`�Z�' 6�ou�ug��+��{f�p	�����M�¬�$u��J��|(>�lT����!l|@�x/0��rA�z��:����Sj]�!�L�������|��;��$��s뫿�
C]b����u@�C�赖L�8�$/s�FT	JC/�l�{k��j4�ƪ~ˢ���|i��'��)�/��%����X���չ��q��<�ȘۯED�[������CB���[s:6�Չ�F�*�j��q_2�2|�Ӗ��=V�9�ڪ���3�� (�&����_��m��l��H�^ds+�%
��ºG�����ՙ�-����S�o:+wkڥ�<*�w�D��_�9��p�0�:D<LSz�,�����_O�r� x�����m�s��5䵽��h��
؍ل�Ήr��٤��{�EO/j(Ӱe�Z��o%q��:Ƹ(�MntB�gj�_�Y�D1�\�}c#���6��S�ɦu7ڏS�]l^XQ_ƌ��Jl������m��7��5>�5��~��eI誺X&~A癆�q�H��)�ݪ��cqt�����.���Y�������*:���x0����kr�s��]�\p��;�	y`�"	�a�P0��"E7yhݥ5d�z����nl%v�Au;��ӻ��L��m��/Z�0<W�ef��X\xX��0"�O�!_�Y¥�EQ�K����tP�jN�
��ٍ��ڬ>$s����EI�@9-�ّ������O7g�Ou(���u#t��k����6kL> ڠ'�6�ZZ�?��_�R���^��`䖱JT�FӪo���F3ӗς��?�=[_��"j�9B�|<�X�hR�5~������O��0I�,x��*�Y�������1��β�\�9�a��Ɩ-`�^va'WV"����Q����&ũA3��F�PUh�w�*l�f�)�lW�{��@wJ���k�����J����q�v0�G��kH꿣�%Xhm�pډ����Z�����d�Gdq��e0>��(F�ƜR�ɩ���D >ؼ�b��v���*�?h� �9���fC��f����Գ�Ҡ��6p������`'�E�-1<6��NK�2���&L�͡�K��*(d�CJ�;R�fm����Gֲ_���>pC��!�T?Z�d�}��k
����L��'W��><驶 �*�����������ű�j��V�º�H	� �3�I��~F������$��\�O����T�w0����ܝ *R���ODή�ms�{bo�vg�Áŧ�^����w���$��Hk�;�����NǣQ�}��`#��#$��o��;C.�`^�:���R�6wW��Éh!1 � u�m�J�8D��E�:%{�f�.��@d˵�4��3�,����c.7?��vPCQ��خ*d~�oF��Qz�1$�M��e��@vVF��8�j�u'�i�f���<5��ؤ�H)�ڙ�p3Z��1�l'y� ��5
iH�\�����{�\�"��u�a����ᘟ�dۓӥ��}=�(�`����$�_&Ą��@��s�PR�yI`��$�������$�^���GB_m�����љ�I�"�̑K�E� ҽY�����"�6n�	���wxA��V�?���|���� �|s�)'�����0��{���s�_��"n�)M#)jN�<8���-�U!#FG7`�.�<@l!�T��YӬ�F�N��A5�e��e7�VX'��x��z�j�Ɵ{9
7��Ok�Т�W1ߋ�cD���Fq�c�P�.$�.�J�K��[r��	e�Z��#���k�F���v�B|IY��F�NjA�5�yp�􀘱��!�gO}j��^�v�$��M���{F�j'�Eɟ� ����Us�9E����b9�&�M��5H� �0��l��CR)�·k Һ�$_��C3م��$^ܧu�'dB�-�*�m�:U�A��j��Ȳ�c�iJ��_!εt1� PX�����n��xc�֤�p`l�+,��D��5jׅ1ú�?�jxup|Hg��7`�k��럭Ln�Y��J��b"�$�"?��Þe�s���{v)IĮ�''�V���8-Yڕ�?�:�?p��݃�y��JTw�Y۴mΊ�b�&�Ø��^\Yv�d���F��N�Rm�oUC�&t�G�<�@x��C�0d��\R�D�p��v}�v�ٓ:�RS��Eo�UȩҦ�*�K��TBԱDI���,�$礣�.��#��d"nB�3���V�τ��=,���tI (��	�n�]��F߱�PѾ�����Eb�B�ߑ���Qe���L@�ׄ2\A��xǝO��,�	iʤ�s�T �^OQ�V����ݹL�X���&�)�]i�+o_���a"V}X`��}{�z�����]]V!S>B���O񸽏Xd�ڎ��})WJ�C '�a
��I���2�	n�$���Z�i�5���;�������Ouoϩk,:o�Uuө�����Ⱝ�?��{�L-�9������X�R#�f����媥D�+P��@� H�8�M܇��?���Qcz�n-̌kZr{��
�]v�*�T�&��̷���.�[����b���x���!Y]�Ng
�}DR���H�����)�_��L:	~�� ۊ�A�s7Mv��p��iv�]����5���ܤW�X�#����\sK1>Bϕ�8�aj��>��
�"�X�p��[q|���&���b�߀w_�+���5b��m���6�S�s�w�]�~{?M�`�"{ԝ��S�Y.ϫ��d��,p��*<`�G�k�������O@�	&����94Hϥ����B�A�}���#�t3�}�;ykE����Y���}q m�3(�]GD���æ���0G�
8]b��m2\Ii4��Sg��iO���7?���:�l�(G��W7�*v~Ѿ����aIמ����Ӱ�N{�+��6 ��%F��\������w$܃뒄�W�b�p����Vᥰ!è��ZU� g �܉�z���a)g*����S�4��м��#y��V��2i�H��s'yH��#}�WMsVɭ:י�3��+9hhN�Qlpn������g��������Ake��*T4O���T�=��n%�\5t.�-���M�̗�i��(m���ꅒ��	N֫���{�&�`-'�Q��Y9�}�۴�Tլ9�.��;��q���TZiX��%;W7'#����_�;�(v����3놅�Tq{Dy��#��g֟�w�v�X�x1�!��L����wx��,p�d9�G6� ��!ߚ!ŦU�iSD}�+e��?�T��ua�QeCh�����te ��a��o�ެ,���1�w�Jk��[�}X��՛VL.rM�a�F�à�'ѿ����7���x;>_����ܜ�:�V4�� �V+��6������J��J���C�\/��C�`Gh�s��{z�V��Z�6���&���7F�w�7ͱn�������x�Fw������7r,}I�@l;*�T_e�[,9؇xJ��0���)涥�{�?����}��:�*���vK7H�9	�����Bz��|S�8�/��i�.ax�oCk�Z�̺���iel���*��M���0~˿I�C����� q�zk���\�SH0-�����ò[���T"ћ�r�qmt��:�����\xp��n"H�h.����?��'��靖� ����i�␳� i>�:���M���Q'�P��Dy��c<���U<��8��O�룮(_I����,�.f�n�Lu�WػJ��0�ob_������Љ��_�X�KW�L�]3@[�B"�s]���O�dZ�7���'����5���?'�� �z�r���N8����y�T�m��:V�x�
�H+�3��*�~aY
sq�x=�LX8G�8��ȶ��3:�B��>u��f��"Q�~�ōӱ�?�5���L&����o1�.�Nv�
bu3?ސ �����������5}��}tx�ȴ�M.�
����Uv%���f��DY�kMܣ���Av� � \��w�I��C�m�y%=�5(?f	��O����)��N�ț�ٍ\�q~�6�w���pg�2FX/2���`C9����J(�t1W0�$�Ž���z��WsQ $���(�a~.~is���x����+��G��&�Ӈ$�dOSe��n��B��%w�L�V<%�'��=��7+J�
�N��r�%R���v���C�$Ƒ)S�� ���	P���=��^\h��S�_���e����09ZL��6�Teh®e8'6�Qx>�~PR��!b;X�9A�)�	P ����<9ضr�'��l�b>1�9��Ǽ	8�����#hx��亅���&M�#zY���Nk�Z�/1ۺB��3	�.ׇV���E�3���x����z�k�P��Y ��V�� w�8:v�L��C4���m䮻E(A%���K��.�Ƒ��inJR$��L�YBOd+�<_�z�Z�Q�ڙB��]�#�O���r�ϭ��������x��>d�"CÆ���m�H���Mv��g6yUE�&T�l����@`���QX�%�)���"��ӛP�>rV�58T��B8�b���7�<�?_;zi�gr�W.�`ސ�oWדK*�h'�����4�6<�+$��?�M�n�S��л����Xl�`��tzI0z��	xTVp����v}~y���z�4�E'�Nz�\݈䷓��jS�+(F�E�5�MkOolk��X�a�J��IК[���!B��a��Y�!ml�0GS���`���=�*�1n�E1�܋E���=AaX�L��RI:�Y�o5mՠ,�n���[���<�{ҧ���嘉0v[��˛�+�a	��5�|��i�tǜ��M��#���U�Ѥ�!��z3�	0�VԮ�i�J;�5q��'H7n}��;�SU��孲�b�d˪��Qw;��1@E���o��}��֬=�{@n�3�Q`���}-*��lP����BA��k�v\p+�k=�Eb9���3e��8u�1�J6ft۩nͅI����|�ɔ`X�I��~�Д4���������e�4����5��;��E�BZe�%Ki�$��s�ψ�*D��e����|۹n~��
^l�R+Qp�WwφJ(��������$�/;�Y`?u�3��+�qHxbE��==�C�9n�K��{���)����?#'���E�5G�Ub.�>}��͏xԡg��rHT8~Dr�����K�O*nJ�t�yB�Y�fm/�#f�>֫��	��f4QVioi��7�2���i��)��0�
��cM:k������71n^�Ӿ�W
�o+�ҷD}\�Zb\m�&�N�N�/:����(���T������&�哪����E�(FJ���l����@���*�0N�_K��q��x=��o�q�u��(�Q.�"3�~4AQIj��X0��t�)�_VH'�f�7�/�:궉6ޯ�6S�R_$�P�@k�BLL/���)��^4�i����ϴjԢ6���p����tk��m��a.H\e߈�r[c�h��%�'R�2g��V�J ��)��G �V���̮���bd��:��6��Nr
qN�#����kl&�l9�kXޖ���Q�j
�y��5�A�aQ,S��\eUA�z���¹�G0F�X��\8يEn7M^�����]IK��?�:[q�rG3�O[��:dv����aK��%
︻5����ѧ���Z�A�,�橤�����X)��]f�R��O���4-��j�|j�}A����Zb������=���歅0��/�a�'�V�N��͇Do}�����؋Q��$�OL���rA����R� !h�b/��o�C�bW@���m��K�A�}���}SƉ���?q~؎|�EXe�am@��>E���խj��e'�K����1����j�']�Ô��Ƕ�96|�p�{K�.�����;�w�#])���'�����d����:�$ަWy�)�A0�k����;Ѡ@��x}�T�-kSR~Ru>��	ԧl�=���Az�Rԛ0Kbh�u�_O�8����T'j ��oNX��y�fD������}⼠�LJ��.�@�*=�I'�d���� O�[d�_��������:�8h��j�r]����"����_�|(L��4�*s���]���g��k0\+��]&GD��[�}+�d�@���q����B�1��#��ih���{MzDNU��۱�==G��gj�����Jt�&w~ξp�������wѲǮ�A]4���ݮ����H��-$�S~��d>���"	50�T�z[l��<9�ӄ[�6ڳÆW3�aXd�+���Ȓ���ݒ��hC�!�#@��d�X���w�Y��f{�Ȅui규�O=E�r܁St9�� 6!��U\y/,�,]�-J�58�po�f��͕��n�hT5�:�>�{�D4�
���3����n倨&fMͼ�������e��7/�� ��[����?5�\���lK\�E��';��x�/ȡj�D:MV���@{�4;%�[��kdA�S�6�O)ZsVM���C���	���c�������^�vDK���D�'��b[�>����\|\8퍒��å�{=]���A�oY�W�u��]�͉���0|�M�!m�Nn�
d�?:b��B���,��)Qs� �o�{]��^~H+��w*���?���-���ը�-��j�H�"-u�Ĥ� �����1�a��f�N(�a�G�X�����.�p�,�u���-R�޽j�.�K`��:�,�8��j�ߡώ#W��P��R!� D�bѣ��KwNG���fp�G��%ݙ���,��""�X<��gB�IL��ְ������ ?R{���Ik`M����h�)R! �����Zi�Tnje�W��E66�4y䨿	dD�?Hl�:�s_���[��Y*��c�/��߆���f�+C�������5L�*�s������2J	6;��^��s�ۇ;xv}��Wǥz�W��%��s&uO����2%#��'��U+<�C#�2�[��K��n�@��F|�8:�i�26��U!��\�5<u=˻�s���?ۈ	��SKJ��8@����]Wc�����r���S'�-����!-$����C �k��)�~p<��ΌW�[��a�+����L�fa��Fѯ���B�H�Fz��V���ڑH���4E^�W_F�����?`������^&�����RyC?+M��`IP�;���ߠ]j��)otXl�=�����P�:��!Uv�������b�Q� ��c��
�y����K_�*�F?��rx_45����K;���ޖ��2/�}6Q ���l�ܹ���@���2���X�B�1��	���HѠ������6��89K@;q����W��p����z5[T�dz�R@�(aM���$n��:�wA��Ƀ z��N?�`����y2ZX�#���]�%��^���,�H��SHwwT<l玷�O�>��(����!�
�Z�L�ōM���9�ڿW��X��]�Ě�Cb����n��Mh�_3���0�k@� �$F�,��L�o||�a�l�O� C��gziV3E�$KKT!B֚;�Z���ZZA�F���][c%��;��m�}C�sg���\9� �Jt�R�~�.{���ٵ�.u�XFҦH|���J�֧(� �� h���uT�wf�az�Ɖ�r���%1&�Ϳ� @�ᰦ�<_�y�5�眬���N���ʺ@��,��@�!M��z�4fd�L�K8?�#'8�ik�+;.��rt9�����=w�7G�4��m�K���,!N��zN��c1ۗ��Y��kQ�vQ�61}=�>��{��\��^u�&[��mN�����ɸ[Բ���Fu�t��օ��by���hI|�����طb�1��X�(Jӎ5�� ��r���5������U֣)�S}�q���l�n������n5��8��ɫm%Ǹt����>D��:Z�s[���.�t��l�~G!��KqEM���6�n%ɣ)�r�V(�"2wy�|b4�4����!�T�mb"_QR�(/�.�/�N1����`��dt���W�K�!�`�c"�nt�u���.�����N��Z4�	�sȵ���X�L7�)L���K  ű��R�����XZX*ô��N��	�Ei�-��6�EA�,��3�D�uk��r������l���ǭKEMs/r aLZ`�1�.�M�e�{~�Y��u��&L�_����%d��!�R�%oؠ���@�J��<���G�;�a�G�Cb�,��5&;V�ݸ��x��{����cM>���?b�f/��1�J"l���I�vrM�`���~r|��� +�?�=E&��9Ϥ��R��of�
:�s�� 	ȍ�]�_Y��#Q�Q�������ڮO�"Y�}��MG�_�[\�)]9�P#A`�'w.��M�	�;�+�"4X13����d�+)�^��LY�F��B	;�����Qo�I	��� ��bo�ă����)��7�߻ZE��bx�e��$���4F5�/��B_�g�$��ޟP���Y謶�T��-��m��9�@���6���IF�̈�?�~@��ݲ}V��+h2	7�X!�Ν$S���j����b�2��	)l��1Oi�G�}�"��w� �͓X�m.D����uF?�}���1zR��Ϟ�}��n����+� 4����
8H�Ӳ ꠓ�q�����lݎ\���SC�BXG�7��rW�����}�E���􅦙�q|D�U��j�Dͻw�9��zO���a<ߟ��g�y�缶����3d�i��=�����3x���2���d''sj7��2~�xm�d�Ǧ�E�O�)�{G�6jtj��hA5"��'/��������ykW�(����ҩ�V�g�6��e./�]a�X�9�v��9�c@���P���.]��^t��@��$��(}��]����)����5�cV�����wڠ�n�Q��ig6v1]͊�Kݕ�P78,�����ǔj��p�U<��?�>g�'�4��dn�m���5���.(k�KE�Sئؽ��������s|+Ծ�;�N�V)����3袗a�yYt�ZJ]��b��u9'�����j��B9iA�шI�_z������(�5+hG��Ͳ�T��5K/�Zע�.I|9j'mK��KU�:�h'@^��� �w�._nOOD���@ M�Ĵ���I�c?������R�
@V� �^�"�i�F镳2	���=���tyuj7�h"�@���Vy��i.�P�@�=K�)3[�x�G�L�5Α����Lq� ��^��������W��s5���f�����-0P�ZK/ߪ����}^������0�F��Q�@p�(�trט����8-�&w�|�d9�7xQB.��V�q�Vп�7�G�S�����A�Q�D���]�2k޲n�i��$�Q�2Ě癓�f����D:j�oLG\�jK�뙅f���ƙQq}�(ǨQJG V�h
��z=���h�qs���)���0��q(��83���\7h�#�wWh2�R��犢�$V��A[���
x`�n� ��^G�p�>-{��}�k�"�d�7���+ ���αr���g�pM)l=��I�_�]��dT�g}յ�=&����?<����RQַ�nQ���;�������*���:KO�>�(��������
HjIr���	�$7���*��(6�c�]gB������S����}���;��!��q!��:X����Ke\'�Kb7�
�;�����6㯱^0���so���ه��e*��GC��y�i4n���]^��e
k#�^<�3�2�	r�T�$E��!��#��:.��3NXWI��.�ͦ���Վ�?報�KVz[���
��i�\�<�'�Ť؄ORN*]�7��s+<'���-m	�B��l��ȋa&$�_�A�@��`i�VD�|�M�m�|SJߺ���	��;ۚ�fi~ _�n�S����#1��g��lR���"m46rn	��>D���ų�qʄ��=V�]1U*sho3%
�����J���`�^�~�{�ؠ�X���8�_[ ��\�f&v`��q(k�_����X^H���a��1�xr�[���Ċg��>/^�f���m�	��\Z�9������iZ�φG�'rtb��������f��|Vs
���^����yD�P��� �{�i$����s"������6	���3�}����z�����I>�~�<�{0!���?sr����Q�����{2�_�Uś��j�����}��v�+����LT��Ї^���H&TY2s������yC��*Gi��qH���|
&	mX���#La4���g�ع×W���/zE]� B��(�ә���#LSu{�k���k ������1�G�єԆit��z���
��� ׊���8F����p��V45��{kC�3��y�Imb^�}�/)�lZ�C�r�\��8nɝbf�z����h�dqi M��3��C)����s�y\����u��`n�w�E��%^��m�vgIcIV�h���������q���Xߩ��j�� _k����Bh�<�A}����ð�*"F��_��қ@^R1��-s)�0b�6�	{M��˒>�e+�ϓf¡/,�h!��jLdOp΍�
}%�lς��<
/p��l4m���m�f�P�w��pHE6)��b2����Y3@�����\}��z�}1��]�Q��]����}�-�j��S����oQ�N�ƛ �l**�� �a�m��&@j���B��3Θ��r�L�D�Q�p�D��	F��� !t2pa4w��~�$*�����M�)�=D(]�yo�\�Ԥ�0��8 �D�����+���Y6�@&mN�_x&�ﺽS����&�˩�!*b��q��Υ�_���y&8�G��1`��n��� ���߁�X�h�b�|���x��	�zݎ(���2.�NW���pS��Д-��8�CC ��	:��{��i>G#L�W�d��=d� (��t�
%46�9�v�j�g&�q%l��d��2��a+��)�25�Qq�A��q��-�$��>%h��E��x>!���%���?�Q���t���d�M@��b������B�cV���?N�R"���-�a
����7`;��!D��++F����ݜ/����g��c�']|�+�2����7��g�s-��P��eϪ��ޑ#�$�����k���_��{TNr�?�Av�O��A�*��$����O!�L �L(�Zv�6�ϽR���6#����v�?9�P\i4=M-c�% ���&~5\3�/8�,�O��>Mr̠CF�e�p&��XE��b[7�7����*�+J���a�.j�-m�%+�%�����k�y+���g�]�y>.V�$���O��5�6�5S$pGɿ�lp� �4�7i}Kz��;�>�e$Pb�Y��rگ��b��m4~�P,��_�f���u�"��Ԍ� �rߕ��Ff�y���sj��S���;~I�����^2��ؼB7+,�<R���j�gH���.oN�,~��o&U��ܪ��>��lV������5H��Դ�> U3p,��!�}?ͬP���H��5����fi�6Ы�qĶ��Z�*�R^z�gD���D�Ӟ*�e)	4cκ3�:A!�"�+G�9y��b���,�I�ѐkw�ʰm-j��A�7���4R�=[������3�$��F�e[eԘ�����(ܖ�0������XϮ�a�z��A��]�i��k<��J������M�P'��P�2U��V=�o�\�������^� jF'�5���JU�X	͉��ZK�'Dx�2�� ����^��
��
����I���9Gl_���x�O��B��W����J�g�oV��B�"��i%|n]_N��+����/�����$�Ҿ��g�=؈�i��ǎgE��^3n�{�	��{�j���-A�CA+�`�8i���U���`�fJ��T`�yyF0Ci.�n�U;7|���<��K|ޓ�l�ƾ�}�������Ln\Rkm4g�z��F��d�7�{�<���'��X�� R��vfFd94i��S�]���s�� �������,ޔV����c2sQ�����������6����Al�\��T�1�,!�M��5�C���,�B*.s�_ښ��שZ�� `��)q�!��(]1ǜQ��W�����y�坘��K��`���o��K��1 0_����5�h���K9��`��� #�d��S
�U*7C���p���1-�K!X��c5(3u�	�2	B�X��g.gN���E��!��tb�PLedS;���Ͽ�[(�C�ۜ��D��-J��|���p��➊gA���8y$o��Zh!���e���N�'�@���#�ԟ�^�����DO��3����o�5�ъ�$A���b{ld�]��K�n���;�9ݭ��#,2*h�\4� >�v�3�FN���+���C�0�ɱTЂ�D�P�WhG�7q�A�u��HR�Z,q��~\�`�>؄7��IB'8��D����U7��#T^��=��m�Ȑ�B�/EӀ�7���D�o���#5���>�T�h��K��he-�����j���)���Zq
�ϬDZ�W#�a�O���7��"�"`�h�hk3����̔a&������v���̂�}����IQ�f��={ټۿ)Mc�]2@�G��P�,\H�����O�d!�WBhϹ�]Z&C�W��~�\ss�����h3����"���#�j�#�^������� ������י��b���T�7����*��q���<L�7�w[�� 1Ǹ����洮�羫Ģ}[;��!��֑o�f3��<��4|�F��fs-B�+��j(�R9�f�O��<�=@���K>X���x�u�`�Ƭ�C�{�u�������fqk�$$77R���]jC5����������6��;�6����r�z��(�<:�x�䜡���D����,��1�׾z:T ϊVGV�!k���&�,@Pu�a�| �Ǡb�� �� �h���Z��z��n�~��m�m�s/��-� ������\������?-�ا�q�� ~>5�p|1��MBI�4u�_"���|j���_��V~;6=R���Bm��y��	+YN�-e�F����˶�7���=@|�-q�
K�	y�PU���f�K�����iU:c�����c�=�Ї�R�Ih3����V�0
�<�D����:1�' \��M�D^8�)m��V�ƅa�r��E��9�������:�o�f��q͡���ǐL�{� U�@��NPr�D�-�}xu���$�T<�ю��:�i�Vڠ
	�Aʀ0'���Ճ�p�;�y�o�fҧ!Cs����7ph�W��8����β��c��M�S椈�z|#�.5�WHLW@:��cÃk����^� 7ǘ;�-�|3�P�ձO׃�N\��*����\���b��H�"��p>5f���q��N�b~
���Z�N�T�oK�a�b]ܸ*�ABb*�̛ȏU�]r�DN��e�ۡ[��ӯ68�t_j�@��H6���Ù�X�M�@�Lm:��X��_����k8�ޗ��b�~h����e�5;�9�P�ē0�4{�$忾�-���Tw�3gI�7�j���I�2L�(%d�N�	�öoO�@F��ro�	���^1|����d4�?�؏����K�oqJ��C-���O��( ��S��,����W��i�uy�e��O<Gղ� k�q���6��3�Ai����Z[�O���^�8����+�2ۛ�ͦ�+J�g��$_�h*ʓ<a����t��a�(����K�
�5c�U٬�E��M�F�[�C?F$�^��� ����A�B�����ˀ����Y�F�M��#q>�}}"nxr�.�e~��sK������	��8����L��p����p�T5���V��0
��k�1��{D��bZ�����e��fa]����+�S���1��#�__ab�|X�j�=?���PȜ���9#K�>�*���P�����wd�b��϶�E�9�����nq\m��8�#Py,k�Z��d;�m��r.��)ַ��C�1�`�(L~vY��D_	�Sg����R\�S��_� ��S+�����Cs���J����jOr|�bu�s&�[�́t.\�BX�����/��yن|5.���&o����@���V΂�*�D�����i��v���9�A�U���E��DѸFf�[ՙ���zu��Z��|�-�jx2Eb���࡛iQ����[�o@+�n��RPB�Ρ'���C�7f\j�P,G�U����)�TV�Zg��v�<�f]��}�
�P��E6�0�|Dw�k�t�����1���Z�1i��p�e��0���W�hpW ��Hqrl#�x�A�E�{(�f�m1����}t�SYZ�	�)o9aA�^,�$8����^t>2쟄�3���mkѣDD��\N�q�{a��Ձ���D9�ex1�5�8w��c̸� V���8�O���
���^�[n�؊��0��3���d��2��y���SnWS�kG\��ŭY�Y�d�|�u/��GE4Ŷ��=�?���vp�*�l��58��������nAx.��,�ҡ8�oe��s��j�:�����^�ś֬랠-��!�g��IFZ��Ti��<�E�ݑ�R5���sNT�I����w��gL�e<��F��s�Z5b:��!�� �@W���j-(��?�=ӨT2y6+p���C)"?y��Oˎ�Z� ~'��#�e�W�&?3�.�����)���=AJ�i�������l�^��<cv	�p��[*�75��ӱϗ���f�Cy@�T��Ҷ��d����1���P���k΋�N*��!t�U �'�,HP�Qiy��{R5��U�-�p��~����|bܧ���>1��=4�`��2y������#�ݒ*�%�y�Y�ߣ��1(+�_3��An6��,�Md��ҋL�g8�@^���``�1b��/���%A(�<	\�'h��]V��� �w�:3N���k�a����ߔ.��48|e┸��1I�������m�i��(�?�>gHßlP7dQ���-w��i��Ĥ���{sV���Tt��©�@l&YH�እ�Ұ�.�DN|F�ixp�>���N'СN9����	�-�5�i�(���,��t�x���1��_�s��zZ���^?�+�H�՗$Gm���H޷W�r��c��H=w�r@�$�����LS�<�.l`�gCt7����0�F����#�+[��@��;,��~}���Y�~7�l!�M��;e�T�ʸ_g����窐)��U�Ne��a��8��Є:�?��-���Hu��T��t�-N�M��(s=�����(���UV}lq	�l�>�2��~��2z��G��Q�d���*���))r�������	��k��#�v����'DuO���8�$�G�Q2��M�m�仹��͐�ia�ga�nL/�t���6>%�P2ٺ����Ur�BK�bF\�v���@�#����1�'{?����Z^���NRTh�2xi��V0�sQ�H*(xD���L)OV�C_wo}�^��]?�#���J���֨��z���o����P8b,�:Y�Q�5�va<|���q3h=#���=��g)��������d���N;��K��-�`�N�V����{���M�9V�\R�0�m �H[��mw�"L�q�M���@������Y��Z	�ێ�$$:��~'k��+�6�UQ՘��������Oﲘ��3�a�-3CB_�⸒>� f�	SQ�ns\]c�j�`*Oڮ�-k�= �+�ڒ��qS�ݵ`n��t��>
2`�"v&�n*���5p���n�4ރ����OM��S�S�Z��|���J��R�~� �ss�-9!�'o�����	ζ���{�cHs��&��/���dk$�����B��w��)�&���Ӓ7<�\� ��f f���$^d�hY����c�U) �c�yHإ�=íڟ[#x��G|��yA2D�?4�'�H�Q�ƒX�=�i��ǎՕ�0� W)\�3qj$�>�K�d��\��I�.��4ڨr��K��[�p-��J�çԮc�vcZf�#����(J�=ɔV!�L�2�ϖ �e��rMQ��1MN� �-�]��F���f��G�5Gjj�=�sh�&D3bFG��v��)Ł����Z
���_��fJU��p�/>?IF�r����I�9��� q�1r��3z�̧ q�hLk{a(�ug�}�dЏ�;�@� ��6�����E2�79���S�%��4P8&}@�nD�˥5��8�1�R�7���>���[f[�8�OO�|$��x�݁2^Mw͈y.����������}�O�F̢1�����q+mિ��-�ᦙm����b�+8gE֎�?œ��C.ې���ځX?�
.D�� u�u�6uF�?&$�}������0fX�����L�$t�;5��*EjV���,plm�e21���ƨ���Qz�{RøŐ~��B 7dz���cL��uڋA�J�sP'w� �����4ڱ�L������O�pZ`T$4l��pk�s����3"	�%~��׼�������s��Wdk?<CӸ $$��(<	"�0��w�R3��l^�iʹ����f3*�����Y�@�T�i>�6���	���.�u��r���,������_��V�mlԱ��e4g}#͡��D� ���6�1�$�#&a �Mz��������7�H�aC-�K��˹�"�1�J��Wm fOn&h�C�d�ê�y����{_��!/��zA�>h� �P͑~�E��:f�KK`Tb��|m�;��bh����{K�tXFǓ�ƴX�'�d=LXJ�K�=e��>	G۷�l���C�/+�Zm%-g�t�w��f����?������������5Ɛ�����F��M�2���o�ڳ��ù���u�5ʌ�C�SGb̑[>9Ju쓳�i��+��9�T�<T���5�"U�5����C	;툚`k�L�$֢���@�[-m�d�N�ێ�`�����`��$rcώ3�} ���/�)|E�~a���b�̜�zK�A��0�5���1:(����6���(��#��2���^���~ΰ���|I����{6�l ?��I�?�)��%S������'�D��"4(�2?k
�&mC���e
v��w��F���׮j����h�$��G2QN� ��e�6O7�Y���̋H]#�ҹ;�~ Lr���8��a���E��\`/MW:[	��XvN���=E��ཅd�[�LӇ�}ۀ�+[*Xbs	��N�K��P�-u\�K	$x�| G#%"I�!�E�ٯ��>���5�g��l+U�#u�p���	���iN�y�b�/��bal�x,K_1�6�?\ڔ�˚+�ˢmH�����H�QO"�r;P�q8Mj����y� ��Ԗ�O���YCL�p��\��
G�:6�R�Wc�O��L�{�x��M<ƚ�?*� �c�FPǆi0DF���[�(Đ�9��9zr^��vɇ�1yO� Ȇ�5*D	��搸��{ܗ��T�}�&	1�D'��"[F!��Y���J�tD��G]r@�oA�*TJ욒�}>�2����-��/����_"G��T#s��^�;�x��Yz=x! ��PW���s�C"V�jNI�,Z�vh~�^�#�ȧz�;�z�h��F�&�-�68а�}D
��%^���_nn;���Gɐ͡��v�Z3%㡟Ƃ�6H�.�&�_�1Μ1_��ކs��A��m~,���u�K���j�l��w��O�� �Wc� ���`���^^�F�-0��K�s+ǂQ���(�+��<>��8눓�y�([�d�4�a�雥ɑV&�\��uQ�CK_�(��'m�؈*��4�v���Pt�{���c��
<�Ep�㳨?�̏�CT/�������7��Eog����;�H`7:��Oe�&���#�0��Of�l�y^��e떍$*!f²[]�Á<��ɗ|W��b�N��:��� ݛ��D�NNSߎ�K�P7�W-3�}"p�,���yř"���wx���=�����Y�qߓ���N�,װ1��ő���FJ�!�ֽY�����(r�yׇ��X��@�CCSL�W�{��HU�KoFr�	b����̡+g�!�.�F,��;ۑs�|�{��a��!�砐��?7��:�.�∻�8���E���:�8��c�8��HM��	��Js=���b�h���.��~���m�j�ȥ&�	�yʞV?���^&9ȭ0�;d�H�A������
�Ytu|דuyl_=��&s9�1>��v�Co_�����I�EK�l8u��oN��D�Z����$�N!��,��P��f���D��~6-T�8R���.Iz����T�2J��d.'+)�=�9�F՛���L�X)&�;��v�2/+8��֡&�Vv!�i~�l���9����G>����}���sA--���9�k��>��{,�Y��K$��?�X5����/�������H��e7�8�.�{0�J��xy�8�*η�;��":��b=�|}�g D)��P�]�������ij��cd��4�b����"v�C�h���"w�q��%!���|X�?�ѽ[��B)��	>��!� ���{��r�A�i�'�U�$���h�~�ߵ�X�$�	F�x�ҟ���8V/����r��nM�׌}��j~��-�%��ᐌZ��t��{�Y�N�O�G�}c��G��DQ���0u"���_d�ڝeCc����t_�>/b��:���b�ţ�dce�!���a�3gу�z'T�����9�d1�ӬH�G�Y�S�k*���L\	A{��z�p��v�<�Ϩ�e��Z�J�p
��`��R��#?)DE1�G5�y��� }S-K�m�����47p!>�����	����) x�)����4�eJ�ٰ�DUx��khX�����Ѯz~ı��x|7�J,7%�u&7*gM����	�D�zN�LK/�+q� �/�����O��Ҟȩ�L���op5����NI�;��=���>q��<�g��n�@�le�t�=�e[�V<��mcZ���Q��iEᏱU�f�CET�� �.��,�;�}1�ٝ���J��V=���S��d�nX����P֭uNa.�	Y�*e!�+#� �f�_��4�ܘ��R�;vp~�g��'�G=�R��=�w��Ui��I��P�E�~II�������++x2.��OM9�M�o�}-��is��߅"���8���\��(�3�1����j��=��D����⛕|�Ow綡S~���{�u*O
�E)"�)�Z���Ď���\�mk���D�sTj!q$�Is{yL���2q�bk|�Gu+1��]z����;�Y�R�ğ�K��:b����4�˱�gi���P�.��f�q��&�b�7�
Wg��
�J���Y8CR�A8�e�ץ*&�M䟰���tR�e�è�@4h���J[���m�Ҋ�4���u������������2������g/�����K˰��t���:���VN8�+YyX���?��C���yꢵj��\����L�`^z�_�0����Ef��U��JZ@�#V����(��X�P���3���%�b&��f�Dt�d}�V����}Cu&S�V���$n��)Úq��oٞ�X_�J���O閱��B���C0��l������fK�j����x��dp�La�$eA��#�Y5X<���M8����/��s��!Jt݄c)������2%���o��C��4?��9�?���-�����FG�紪p���aҘ5�>+l��\�e-���@�o-tQ[Զ�_����q��I�Fn}��:��e᥄ *��ܶ� �I��X_��y�t'���!��hDFU��6q���c��"�'lQ���_�HX6�ɪ�pt����H��h��2e��޼�EË
��l2�?����	�����:�Sgc��X7wo���:#�w��D Т�v!-y0�HM�b��࣐l�x����p^)�����Py_KrM�Z�s��l��7h�89(��7���&l�BҙP�7P]�:}�X=�f6Y3^���Ja���
?�_Pc�q!�H��M���\�uV���&B&\8�Ι�l����p��Rb␰:��9D�&�������t�P	@��.�<��Gǵ�6��_���x�Oh����l��8�*��r�x�0��F=g�,Jb9Z���	�z���ʈ��'S���j*5�fI�z���m��h�{>3]�u�2�>���� ��I|�����)��C^�%�,~ߦ�'�p�Z��������?�TI%��dZ�C�F������̗�(vH��0.�|�*y0�C�:�J)����۩b�k����,#ˈ�Wo��>�9(�訰����fi�X��}�T��K���I��t7�QN[��nPN�pE�:nT�|�t��� <����yS:ղ4zE��Swf}Q��k��Jj74�����W:�P<
{�8����v������
-�R	|�F/xИgz��H����HLx���B���;۟{/����H]���<��yM�	�b��Q?�~��� ��ՅA8�B=/RK��x1�cC��ǋ���"�n:#*k>�ۢ�2[��=jܼT/� Ɲ2�`qA6(2���L�h$�'�o{fsB�v��:lZ���͢��5%G�%�&z
�G�VK�p��n������_�&������i��Í��;�Y]Vo�#Pݴ{
d���\]���nM��"�$�A~Y�j�?�
V��']� z�ֈ�"|��"��b�Or��(�EK�Vc�l)<t�9�%��W�TD�=&���W[
��ی-�e3v +BN�J=��ݬo
���y�'�2�H${,�Ib��ҏ�a��b�
`ld(�PE�{��w�^��|��i͐��/i����t��)W�����&�{���o�}^iͷ�m�FTt݂Uܬ5��08[������3���)��u���T"�8���q�:���T�{f����`�UH��r�V�V�:<�m�hxM`t�!+[��g��ٙiB���|�0ϯ��r#j��*����Vn��˻O=ہy�=ڰWA&χ۳���~|vG�jf������L��	�~��5�8�{���Z�*����	�25`Z�g�:�4ӅĘ��"��(�_������C����	#�	�6V�A���!�0�euf��J 0
i� ���c�9����S��`����^�����<�I��C��P��]���>�3#3�6j_��D*���� 8[���'r[��p"��i.�˵B'� +�ڵ������7��x�j��Q�;��ڒ[eZ��ok#(�&YE33��vJ��`�Cfh!�9�Y�I���~q-�YsZ�{\�?���υ[1�\B���o-�R�u�A�:�[�|�^0��E���&~D`�X�n�#1<�2#���zj��i(wGRGY��\��Àyk�et�<��z���H��䪳���P��
�Dq�c�;dFj1#{v��t+6m.��)��͵�L�G�m]S��ol�%���Kk(N��t�'0�)3!x��@+	!y�Y��Ӎ�(g?�ݼ);�Q�&b���X짪�Ġ���b��7���4_t?�!�`8Vk��pYnb���y�3��T?W���I����l��g�Jv���F����%��&��Q������`���$��c�o���<�6_$�A]���'�=t��X>7��3j6W�x��`�ւ�:�@=��9Kn���
C� ���(������8�
YcSi�uq3��r;�3תö뾮f$غ�l�mk5I��F6��z����#Q��]曛k��F>�E�r�0�����|A@�ՠm�L�;�JŻ��H������Z�va�*5(��V�
����O�IH˯,��.ۄx͖Gq��g%I�^��t`w|�/��g�3c��rK'J8N�lQL�]d=����|7������#�T^K�B%Yb|l��jۜ�i��D��#�@./����Wv���f���KHn��(����Y��a�j?�wQ�;�]BK���ti���CB%F_p�N`U�CR�ab���g֨n�f�~�ya:I��3�[��1��+>֨K���m.?����_x�l�Y5-(Ղ���� Y�'�H�n.�����Jk��_��L9N��nr5��'s�B�FJ57H\<?�[���E�gN"��
�6�d�̯s��A��0`4�8Ba<U]v��S�'�ʈdf�*��j(O��=����ժ���c���GcH�97T��&�BI�r�������}Ӗ핖��|�F'=r��~ ����ֹ���/Ms!;z��n/E-�k�k��TL����}�$�
G䴖�{ ��/�C�/6L�a���Gq���0i+���[��i���Oh�)/a8�T7D��\�����[y�1��Dk�U M��k�|����߿	�!�6�<!N/�%��<��B�hjN��
"�{s�0����
&f"��2�-�a,B���΢ ��.*�)�·�ɔ�U]��Ѭ��N���eg�¬@�K%ƶds7>�I��hL[z6_�������C)+X�v Cr'&ϝpW�G&8��a>r�����h�]��U���usC|s�^DI������J��jS ��vD����9/2��(n�2�Zß��N��^�e�����G� ��i����V1�E#׭+��;"��������hpDG;����<l5��<�V�%'n�+6�����9���+��1&�b{K�iV}�֧vx���HH���E Oն��k�=a��ȴ�f�7�4@Ȋ���{M�+���ؕ���o����Ėō�O��$�0�C�t8�jmL�O��[���7#�v@�cB��@��y��-��fH�@�]$t���̼t��cb7�س1ܐ�ĺ�,��Pј.��%zqO�K~�X��l�`��)	M{�W/0��릋	K~�n�HӓR�Eg��Q���2���[�i����<t2��xƚ><���6���#�zRzӇ����vQ����U��2���ץ��Ӊ-�-儾�2Ŵ�l��u!�X��Їe��>�
GC���n�[�N9��C�P��,�Ob|�S��Kŷ�w�R(�M�I *�TS����6��1�Cf�h4�[�䈚|���+�?]t,����=N��]�=�"�!�������tv��u΅{�D�[�?3�;$YTRA���~7�`�[Q3	|�6	{�P�e.�����k��z�B�N�Ow� >�9�PZ�����Q��F�W�E�����)j�߁ܳ9��x[Z�c���	<V� s>��`��_���l��qDR��$p��L��.��	K/��Xw�hM>�����Scޔ��h�l=�'[�^��D�s�Uv�X�D��%���N��O����gl&��(���!���K���̇:K�B��pD��d��I��$7-�sWD�!xQ}x�_�ƣ���#Gg��0�� x�����Ӝ�	'��3k�EF1U���1�g)E��k� �5�UaO�Z۠*|�@��ϵ��m�ʱ�+�L�������K�3S�ʆ�4�~��)����K>��EyH���	�y��3�}w���,q��Z���i�ڞ4h`��u�47�ݪ}������CH�Q"���O��`��Հy���r����?��1���/�����;p6�%:�D���f%��#5��C:��T��;����毋|�e��+�UH���}�r�֗zp	�'���g����1ch��.B��o3L,��2uc��Kʀ�y|"��zI@��>��7
�d��j����y5�mn��7�IW�#��Q�����/=ϋs���4s���EIƔ�ot����\A���<`��� o�r�%y��v6�r�R����.z32G'�W3V4弐_���{�#��������갫�K)F��Q�s~*,�\���Ͼ�m�ɳ�?���
H?�e1L�/�-/�T��~ ���3��@�lzQȧa�<`DFA��e%J����^>?>�$�Ltڇ٫ڐQw�����,�i�V~���Oȴ��J|�IZf�o�:�:iW��gc3&��d���$��IǶ}ˌ��f�Vʹ�r���~g^�d�Tz	�U����hC��& �)-��>[�Ѓb�<�	��A�M�>= ��e��bt����S��I]vΎpP�Ap��P�k)�~�'�x�P���>��?8�,�{����Ψ"����]|ۏ���4�JAV��T�pR~�k�*�R-�p����90#7�q�U����c��� `�J�D��`��?e��3S���������� _S�3B/��^e���b��6^��|��\�v03�z�Z��/dc��-/�7俷^XP8U�_��H`��Nk؛��8�Z(Q壱]OV���&(�+�G�&^k��..�5�O
�������9�r��5_|�w��<�S)�T���
������b6�$3�RZ����W���&�C��Y:�5&&�T�$T���ˣ�C���?w�X�%�#�ж��b�="���d�q޺�~���~6\!�[}f��L�0��KV%�"T�����Yuj�>�kj���
ݛ����q2���#�m�wnt�4�h�q��,�M�g[ ���9V���˹zji������W�&8( ܀Kb��e
n��� m��x�U���|\B�1��g�2$~��m�L	&�F�@�V��`����`����,���f�]H^�wj�4�k\��Q��]�.K W<Gou��g/	�x���j�t�`����g_�z�S�_�H�[1y�^��oދZ���߮�J�2��w��6|ߞ-ƞ�.9LDׯ�þ���t*�H�kL��*0p0#�ix���l����7��@C�W��Rd��������\3�*�GZ:jFqp��C�1�(�
�<�.��E��9ًH%� l1M\J+�]�G%�	ȼJD�A�2�1���S�i(��τY�-s��8JS�d�W��P5*�oI�S֓�n���Z�%�̱��)���M:#�����Ҡ.hʼ�L~N����?Y�q�9���.G��m�0��]-_�������IY�\�n��?��C�a�p7�gratg�ǂ�p:�����uB��[o�{0�o�����)�����}����u�#Eu9�iǎ��'E��Gh3/GB��bxB���%h,�����i�%�Ǽ�����	Ɇ̆C�U���~𩔶�+��7�|�XF0,� �x����,��dDV%�F?��)��U���!�y��B���;Ս���~�i�E�Y�V�z58���C�x�wܪ?����}�ed�v�^F���Þ��� k��#>BT	Lo�@�Ϳzy~*1ˬYp(�Z%D�p&n�e�r ��8�oD����m�l#�F��]��ǰmuxT@C��#�����
���Q8o�{iT2���k�Y0f������b�L�BP��g�{\� iR�FJd1�:�3��\7�vI��[���Q��*�[��w}q���B���l��1$��&ii��׋`X�k���+�I�Y�����:�!~�m���u������QJ����0�U��Še��;I�{�b)�'�ܑqx��Y�֡n��g�&  W���Q��j���xd��!\Z
9a�أ%�tP ڇ;��Ū��]�+̤���_�"(�}��~�cH��8F���ۙGd�F��>�jP���	�FюT	�q���5�FwhiXV��f�8@5{�U�3��=�N�H�5mX�3���������j���M��b�'�_a�͹x���� 8�����.{�
��]V��]���k��^�$��J�u�8r|b�fM��`��9��c�:���X1�,Z��QM��w[�=s����,c*��&7������o��㖡�s�i�[�H'p����n1�9s�ࣥ h��H�s9��jgw���U=����[V�U��S�n��߅��,� �d|[7�{I���ʔ��Ⱦ�'۵��4�e�q�tp��b:���l>��TA������2-/�@gՈ�5��k����� �c��iu��>��DCvu�2Z��8T��m�rѮX(��wmL���nV>§l]i�tx����x�[DuP��3���)H�/Cc~L�_z���v�D����g����5�uA��/V�x�~
��p]����G�C��'~�ڟQ�/3Bv�߱�\�c���ٿy7l����(k���`� ���xDy�~�H����y <i�~�3;�C��*�氥��|jd����bF��ggl'��W�4"�����Y�FTQ�4��B�Mv�+Ҁk�e�Q�J�[0���+��O�M<*����qV���&D��<�#��}��>G�%��
��X^�F���y�VU9����~݆a�,gL� '$r'����dƑ1�r�ҿ�-2�^�fm�J&T:&D�Yz34PN���<c���3B�(�<���y��X �Pu��Z��(U�M�#�n��%����׎����o�����[�&h���=զ�~���-�Dq��u�2d��ͻ��bZ�&&��ly�\��ܜ�Tl�F�y[.�
3��l߬gػ�#��3�T���C�{����6��KI�~��U��&XU1��@6d�!M'E�����\����Lݾ#��r�QMK�F�.T�� �	��S��">���@��Դ7��J�,�'ҜԴ3<�i����~��R��N) �k#@U��q�vZ�a_���)�����\�y�$m���)��Qi���k���b��(�;�J�?�p.JEtP�!��9D�4�
�5+,�;O�(���t[������_Ŵ�P��G�?s�Szs��vݛ;�ڜ
� �B�a�ۅ���ŵ�,��J{�xT��ͅ��u���Xjw�����l��ڳ��򿥆�;'^��ZI��X:�&|/w�I��	߂��IQs�ej�2���y�+	�^��:���(!#�_h0�Z.$���6�aZ�5�f�ej�A��% TC.��m���~u�b�N�lKU�;��� �B���E�k���N`�\��*M��g`LSp>;��F��n�G�y�͠3jB<��[��
1���T;0Lt)�{�z���n����/��^���^ҵ3?c�DZc�j�z�Dt��-�0ެOn���r��(�grF8��D1oE��XI/[8}��0�0B�/&� 9�ы�oCJ�����y>m�Bg�p���zO�t:�Y v��Ҭ'��\����iu�AH���x���Q�ꪧ�t/Uxm��/fê�0�u6Xͫ.�6�%�o���M�Wo����>�i1wO�5�\L�i3�!Z���!���g���葷:��w����F�#���9���u!��ؗ./D-����u1\x���:%��8d))wT��i�\A;�.+�,=