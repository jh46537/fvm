��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�w�\պ}���'d��qx�Ba=��1�@t�lo�ܦY`f9��GU��O����5y�k�wy5� e%�iHF�K~3��Z�������# ��d|��̪�����PAZ:�;� ��Փ�?�}�F��3LY����U!a�N9+
�\�:�-��*����d��W�L�vb��+�Ԋ��r�����WtUItq���E#�N]h���]���m�5��O�B��Ռ�f�i�&ǿ��BO�7�mT<n�	��S�w5��hS_�D�֜���,����޻����
n$
�b�E�ah���_X�'ڇ��)�0R<���X��\���-���dw��rW�$�N;�`)r�o:�Ӿ�o��/eP.�����DI�7t�4��u� X����<%����Ś݉�c�b�?�+���8w��'�,�v8$i��bS{2�XIs^�4�P{Q�Ž`�M���z��l@X���	}����U�~��@�V)=����?e6UeC����]U[��������[�������}bw�z?{:7?���F:�H[c���-�6	�Z��qPψK�c $]5­�����0���!��`��ߜ��8��>���[��GrR�����K�O��q���a�̾O�bl�ہ����uL5�����B�>�U{�'��p�:&�U�RV|�{��4�0��w�	TT���F�d P?e� �D�]�[�U�6��
�*8�FW��e�e�gn��J���(}Ÿ;{Q����7y!([�=�W'����޾%�&Uw�vX�(ȸ��Z���L�R�ߙ5�d�d�F���,k'�2��Jv��-��c�m;?U�H5.Y>j�����暈".
���>���L�v�L^�U����Sh���U�o	C&C7}H���C��W��Z7 �k��Ϙ��/��^q#��'`
g�H�,����ƽ}�pd�6=�=dj�h�e�#��|����-���Ѓծi��O62���b��-���d����T��u�uI��,<���CU���`QW�
���q�5"�%RGW��)�|�J���A?p!�d�����iJϙ>�^Y�!����;H�(.]2���U;p��l�t-]����N8�Rix�2�����x���*I:�������;��7}[�<ܤ/O��t�'��o���y�7:���.*;1h�����,	Z
�|�����2�D�L��1E>c;^�gӿ�HH���4�8ҙ�l-����pP�a,\j�3S���WD8�N�2f�g4E�S�,h�B�L��l����R��Nl�Cf`�;E��%�s���c���z�;@`i���\�c)�TV�F�>�C�0b��]&�
} AZ�R!�2ڴ�����6�q
קTR�ǈ\Y椗i���3a��;S2�i�pl�b��Y����2�f	��խ��8�ṫ�44�ĩy��w�ӑ<Ԯ�Fo��=R$Y�{���XU�>�B[ǵ�0r�/�Z
t�.9�;Da�Z}�ФE��%����Gk����ͯ���	C�J������Ҷ5��;�NqЄ��o�ǾK��˩�]�S�x��㽺���Q6}r�T�B�a/�<勉���p�\���G���Bۥ{�:������	�`�tO�i���o��B�| Ǎ�}WQ�d�Z�7��%&�>�&�;��}��A�Uf�L��h6�#�/�L�w��X�,������8)D���TpN)d�����9�Jމ)��ⅴ��Ws�#**t *��~�U��u)U�Ҩ,®�������0p����z����Y��/}������ƑT91�mܶ�-M�_'y@q��,0�����ӹu�=6�v|�ga�t�a}�?�0������rCy��=:h�O���iG���@#FFenڄ�(H��sx��h	��u���6�����7�N޶9U��a��(�|��¯׽ܐ �fp�m�-��a�\�l�B�J�MB�d�4��Yzp�5e�a�*|��;�j��:�d����Ϩ3�X^"��Z�v��m�~|g�{4����ӛN����B���4�/?'� ��Vhj�,X�SKc����d�()B�^���a#b�����3�c�S*�'�
��M�B����WtgO�b��c�Կ�c��r��0�XG�kK>�����}��~�+;�|�4+�ή�6��=���,N�X��9鸩}�+�Ow)��15���^��)c)Z�&�Ǌ�q������uo�H���*;9�z������<:H��g�����zI�sKP�m�=��2�u�v<V�\��U6�~:�}�f�Ӭ |��BS_8aх��;
Vg��6�� �1E��K��@B�}�v*��C�%%������L�M��Z�dW�-��Ha�Ե2�+C��	POF�)��1�MK����m��_��hP�u����,ص�C�tc������֠'��v�yI{��p��)�5�}��f��PI˚�2U)����|g�`ѭ;���,EpP@�}	�Vr����G�����k�����b�<�t�P�Zmi�a!���eMyM�=�]��*7�2=���11�8��&J{Y�k��a7A��f�yC����eR��u�T��8�N�� ��Ԗ��BV����J\���D~�`E��R�llU(��y�Е'��҂���T��x���w2F��9��#t&�����[��cƮd_d~�.��1�Fٯ֜z�/�Y8 	��:����4*!��h����� ���-b���v>Œ��^�c|KR�Ն�2ⶳ��ݢX�ĕ���z�/�l�V@$��pF_���er�C���4wS�Εf/Fj�m��G�yE;����TF�`���\?S�idR;��Ί�O<��|�kN���`e�>&0���r��e;�׶<(-'�I+�,��~�^s�5�z2�͏nq�����juk���� �?ś��5���N�/;�`���Н��l;���T���̳��f`ў:?@Mg��%3	�Bg�_�g4H��[��w���TTZ9�#C���L�Y��C�An¨!k3�x��Z���-{�
���V�%Q�(�$�psd�WQqS�N_�h��y!%Fe-`�G E�:�I�����w�3_�O	�hmf_g�L�E��N�����*�?��yrs*�'�FmЈ�GU!U/
�H3���dv'?���O��J��@NLI���bƥ���k$"�g.�ۓ�@*�#�4a9�|k(�;C�_�.��댟�@����H�S;�Qq�<�Xgׅ�?���u]�Y�Q�����pBя�s�'q1�$nsh=���eS�z%�`���{����� <���aB�V�V �����>�Ȅ��{эJ�] �>m	��?a�ڰŸ�<kTl�����&�n±�-���&�\A����}49IE͍�?l�DsW#+-�֞�E�f�JC�gê�)`��|?������!mI�1�h�9Z\��j\:�a�����:}eqf���)�P����6	�$2������7��\�,�S���/L�:��!���D6V���Uŷ"%�F���.b��ݗ�����R�*�~o�g@��&���a{yuG���5dv�kǣ�0���Q�����?��\Z��ަ0�A�x۾HPv4�/w\	,3��an����l��c�e�� ;��[6�2<��I���m�3�{�3�c�c��HX�����@�&��E�t�Jg�A@���~�!|��y^�:��Ғ� N���}bZ�_�Y��q����W赹���%�y؞W=c������U�Y���fc]�i��-Amg�#�M:F#�E�vr�0N'���ô���J���I�;iѶE��d�=&o�>��M_������|T��xޮ:TN���-$���;a4�ԎĬz�����_|��7�����u��Z����5E��}q"%n3%�G%�t�,'�kL�t'�ϑ��}-�63����I�Vd:Fǔ�g�,+J��5A�8��TwPq�!�]6�X�6���D�~y>}�C^J6��ݴ@R��i��r�6@�H�f��϶��f�N�Ji�"<�k�-�ばAUl����gÈl ��z�蚚�����}�z���(]ǂ�K̕���R�x��J>_��,�Vf���yw�#���� b���E��Ϛ��!}�;����yV|�	a͠m�{bo0C����r�7Z����[\�yy'�|.QMnQ���!hp+��t ZO<��8m�(���5���O���I?8�Z��$�`�im8�����\(s��Cɭ���x�9?�uI�aP���V(7[��;�pݙ�}Ġ�=Ch�=˹��0���C�!��i!��Er��Z�3i^��rA�r�z⁧���w[�� ��>r��i~lx�b�mv�� 5�TVYl�
�1�B�b��<	$>s�tr�v��0|��]/�_����,�so���������ˬЭƬ��
o\��VO5�0uƟ�m��Hu���q��8��)oLw@�_���!<3ښ+#Wۄ�6$�l_6�� �ҩ�r�>�V[T,6yjT�9`�K�95My�6�p,թ��k��b�oe��v���&zH?ػc�Vp�d]X�������pU�-L����8H�u��@T���\��6��O��]+��53�c�}��@��6�X7�Ax�W5��ֹNu���@��NK=�}�&F�����^V���CQ��J�4ӱ~�ê���ka?3\?��tm��p8[t�\��-yʨ�ހ����(z�D�{���������ȥ��	��ב���t V�w���㞆V��U��a�3�xY�w�U�?�U"#(�&�m��X�|�8D/g�[��щ��w�*
�J�do�4)���/�A��ʙ�����Xd���Y3�����
hJ�wm�TUG��f�9m�J���REp�N��ɠ���TQ)ڠ�/%�u��l-b�J���#	��\ﻛǈ��>0��]�d7F��*6p��<
E�'V�2J��l�pN�S���d�]��o�N��,��[�yz�=�4��c邏��o��3���3^�&T�,-�j�J���s6�рDٛ[�$��i�G�q�u�z�GHN�I��@�]����q�t�7��z'G�~P��|q�N������.�2Y�j�tO8�A��9��<ʷ�������q?�5Xp��~���d����~�[�)%+��>�:�i�&6�0Y+�p�}�fԈ���[���)1_�ށ�$��h=�lf�Qᎊ��x@˵��G&Lh��[������1�-���Q����4�҃�+u��qt�2p�Ș��ϷTG����Ă�q)�Ɔ�T�APûj}��,Q�/'�*N���R¦��$�.y�}�G0�%
>)A(�s�G��.�M4�]����亵HR���#~Q8q���c�#"�Y�@$��s�o =H�Gj�w.MFQ���Ct������D��>��\D�(s#cݴI����/q:S��=Ϫ�C�y�b�Ĺ�m�j��W��}	]�@[�D1/�GV� ]�� 1���2٥��QZ���cIY�u����dN��(����,�O�9��5�#��}(��Eϒ����ڿ?Z�	���Pk����9�%�'���z��t�SQŨ��Q&� رsI����|�C_�!e��A6,����FV�����#���� �x���\���ոfP�p@ф�)W��}H�~��ߗn~%])�0�����CWt�_��~������vCH�ԝ�����N�|�ܨ��9
�~��+�t�2�M�>��/���%yb'B�N B� u����J��`Q ]��*��u�ğ�Ψ2�6-N�kR�9/k��ͼ��se	}����z�< �a7�b/����a�?]�N����,Re�3��5�g:�M�n̅.|F$Z��4�� taE�M�N�G�L�ح�%P�|�7�F�E���Z�Ld|����-H�/ik�C<Ոٮ�7<��ߥU�LB£�9��-�#�H�����0\�r�������e�*�q";j�|'�Q�1|�� =��a�J���Ͼ�10�='V.j�DĪ���+z��I$�w'6;�:�m�"��k:T`���2(U>�J�2�j�L��O�A�E��g�5'��Z������%���������J@�F\�O�Q��a_�s���m�Uwn�z�{�_�1S��R��E�����AE"w(�:�0 �Vi7l���.�����Ǔ�8���վ~9XK�Re7�U�.֚����U�hq�s���m��_��i者V�1�$hM�4j&��z���?�	c��с8���l�)�Q��$��Q�sa簷�E&w7�n�<�aTc��+?��U�U�3�����c���oD���� �5�
Hb^��O��]��85P����c�і�xz�+��S�<�#���T��-W�T�C�0Pa۰ri��5�G���iz�ظSLQ��'�M�Ü0����s�m�D�oݛ�NŞ��&x��S��0;��g�9�F��T���F%�31RT$�r?#8�B�bKn�9��g*��h�x�Z��`t+�ͽ_�G���T�?R�]1�bz��22�sm�0
�5z�{r�Q܎�������r�V���I�<3��/Ϡ&���R�.�@މ�ڰd��r�&��"�2N	���8�e&�}�u���F���e�2���_S�Ω�b̈vr���z'f����m�����T��v �l����ʿ�b�J�_��E�T��3���[���Ҭ��غs��8��M�uC<�)"xU�Gi{�;��<�I
�>
�ika~�(\dPRW�Q̿G�埻��V.ް�(�~���;�����A���Z�>���{7*AQ銃i�dT%��jK��&*ꌴ�U��(��M�Ԏ�%���r�5�Jβ�̏��Ot��y�ƶ��i�3����0���vǙ�hXGFh��&J́e6.b���"de��G����]�������N�12��?C�amBV�)�}E�p|���}DP����鸝�][�ɚ<�[�m��Y-�o��ڊ��,&۴V�&�T��GgϠ�2��	]�����nŎn�Z�Au�t9ʜ2Hx������q�v�)�]_VkH) �5i�i8ͬ�)��*�˪E·���F��8�^n:t�0�0�[jK�J�.ҴcD����ֈ2��+���^��JS���e	�:\tZ=�z�o��V^�Rf����KCAՂXk[ @s�����-�t��A �S��Ƭ��(rIʲ��B��� y�b�4p	�t�n|-��J�� �p��$�'-c�_�����E�!qBߢY��=I|�>������\G�6�ϩW��C�NDX�*%L�۹��[��c �C�9�����ʫ��d��~}2r����c