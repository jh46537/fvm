��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"�.0�у�[�Hd��r�vJ�?��Nv'�׵�|�!y	�n_���/�hSm��U�����X[l�y��ǋ��<�6u\��#��D(������0���?�����(%��^��@�Qڢ�{��xOP� ���cI�qp]���ds*�iFk^�׌A�K�w��)=f��ÿ���S�w)(�l?!�][��Ah�z�({C��!��K�Ԥ���بF�4�`�/#��|��_��wv 9/�6v����a����?���-=�Q�D$f-W���E�u:�&j�����}�����-OO��b�Z����^�
�z��-m9pڭJ����VH.6��Y2՛d�.U���y˧C)�����t�W��	,�����q�QRY�mN�,�)���lh[۽�GN��K.)_��y����ߗf*��F:���j�`�~v�s��8�TKW��S�焱�M�"�Y�&�.�= �0��}�{�m���Ct�1=J���t;�yq�d�5��'�l�e��%�.�Q�A{�,'�1<�'ua�Dr��	<j�{z��&���G8�?��B%I��&	�l�Jp(\o"�M��h�9@�^w�[�kB�ʨ�ɭ�H�g�|���eeN�C	AC�b�9 &�?<�	�W
�h9������택S�Yz:sc2���4��f�td�����d:8�8c�O�9RI��v �����5���:o���_E��̷h7�'�����2�����J�7b��m�Oly6?�lL��iF�W��	0E���ڋ�1�z|6��Ĉ����)Js�:cʄ�H�w�T�w�"vC+5��'�V�����=w?��f#�1J�-Mכ%�op拗-$���lE�#�B�!��y�!������Awcic��eMLw���:�m���&h�Z�H{J�gz)���<����ռ9�O�w��g&�/���0ڕ��lp�����������!"1��9�<��zÞ��K3��?�o�8����s�����.���.��
v���u�DC��`�C>o���d�]��r�vf�@�a��JD�S����9;��Nk�4�da��7�R �2�r�MQp�0��$�(����j����6_74�Kg����m׹J�R4Y��ok%-�2I�-&��X����ф��r�NJ���9�����"�"=���͞n>>����	,+�;Y�=}n�3F_���8 鱶�Ե0V~��)ۉ�"�,x4q�%_��r���&ne+��\8`icN��B���%ٶ���:�=�x^�l�\��y���+�wiT:�f��˰`�E?Q��	/4�/�������½���i=ܮ� %��~��Qg-�(��Ow�	��G�G�!<s�̭h(��ۦ��&!Xը��,b�9�w�.��s+�s%��V`IIKضB��g3�V�3���$t"�2x��s����Gm��$ZF�����Nu�^��k됫O�	�v�^!B����&�؝�ewF��c��#=��Z�'N�cZ��M8���<��0�(������?��Bk��;/´a���K��^|6�;�A�݅����%Zgn��T�+Ҕ\�WFk7�oe�ױ/�Xl �Jh���x}P�l���t���0��<��EP��sb-y���E�&k6j[-\�ݦ�{�]松��%K+�,��t��ʠD�ި0�pb�hi���Ow��1j�k��pQ��}�j����cNi�6��ڲ�D�J���[�.TܧP�M,�k�2q��&�LG������T�ݵl���H�`9��
HM���V��
M ko���� ���H�Csu�o�)J�5��-jl�M�Y���Α3�֔޸��U�#5l'3ζf��O�*�
������5f�i#P�3�O�Tٗ�E���3����`p_7tۀ�_�dR{��G����0*���M�<�
H��L&
~ ��^CX�g/s�K�W�&�g�"Y��u�U��"U�ݮ痷i��)�A52�O�@�iGN {Ĉ��������9T�t���؅�:~��%|N\���d>��������L��T=�-0������`6u��T��:�_б��O��Qm��);��Լ묲���t(�rx������MM���t�%�~rk�6'6�̬�����-�\-���˂��#��M�'����q~ ���B8@�AG�_N��G&�`����ր�c̮���$�a3����R����!������}�)�n1�Xv�u������N+&e`��?r��/ۍ��w��d�� 8�)�C��H='nr�Cr�3�x����Ȅ�į��b�mF�_���FJ���sD��*��y��i���ud��p^��+�mV���@ ]c��S%<2Q�P\�y�Zb��P����c/��OtQ��Q�Ƚ:� �3���\���Gه�һ/U��r�D��W�`
��/�E��I�}�`�]�*mE���"SA'��݌��EH�*���+�����i��Bx�`�9d�I_c�o6u��Q1� ��d�zh�?ք2{�.~@�K�?��y���B8�H'V�Q�`��ѓ�P�K�
O$h���΂�_�z�{U�W]iW����sqٴ?>]b�6�Jݴ*h[Fb���2��/9�[$���3���v�&{2����`󳦎�_�6�a�s�����)���ǧY
ǫe�zl�vgP-�Zgt&p��^�l���|��Q�/'*��#4�3����:��������,~��{��JD����-q.`4�R%IE~�	�/
������6;;W�G��u�U��&���R������A-,�<�S�!ߌ�77�3tHA��4E.����T�]珝#lP~w�{�B�&����"#H����M��;B�*fr�~�VA(�k_>�˷x)�E�������r?T���3��τ^֟O��aoW�נ��������Z���M�q��\MΕ	$
���ֆE�K����j�%��#�9M�/���H�������g,��F�+����e"����84���-k���;KZ��1��Ϲ�(Չ鈆�vr�ub�ܜ�%�l��-ʄ�@�@�`K4Hp�]��v(YY��<���m��h�*R<��PX&P�d	�a��q�Ɍa4-�f�佨,/�G��p�  ���0ꀉ���Ǟ��UcL���6��U��$R��'��eVK� >�$�ÍL��V��<������}0�&p���2����@���?w$~�Z������y��t�$Ʈ�O]mT�uFr��.��+	7�2r�)��PuQ74� ��[��=�m����#�=G2�$,~�Hh+�N+�g�X'�r���]�
r�D��gB����G�	��"�����q��[�1��N-&CH�N;X>0pؽ�6p��K�$%�����TD�w2pL��<�W�|���r�q����*9I��#(�����"����T��&��x����dbv�M��!��$3��`;���A'?D
#<���^_�t[�bͬ�AM�J\���I������T� �*��pA�GgOH&�!}?�BQ�r�ۜA����rˑ��9�q	6hL�B㬓�	�N�5v�O�,�!aKr�3�ZD>�Z��_pո�c�@&��D+9GW4��L��F#�$���A*S*�
j���5V0 YQubl��"����Y!��'3GE�1r\M����̑�kmnO}ƴ�lڝ�m]���1=F��O�kχ�៤����sCA��q8Y��R[iC��T���VP &ݱ�O���.����2��3�Zf�zS{�h k���(�n���2v�u�0@BKO�9G�Q��W,��)������J]$=�~﵇�a���,�Ǎ|�{F�`�P�x2���=z�f�����,e�]��Z::��y��&L��蝶U��E�4�����z��*K����p���*G�ˍ��뒪�w"�D���#7��U���f1%JRwxZ7�v�D�X�F��۱�9�\���s�i�e��� P��6��T�Н��x����0\YK�Sc].������4��dH������a�����2d7�E�y�������{z�^�A:o��]��2�(�W�|��k7���U�)E��${n�	�gfh�&]�>5j��\�뺙�+��m-s��H@/����fm8�����3ν/s��}��=ح�N��J׫��DT�:�`�+8��0@=^�ǝy�w��_�l��|�!EJP�p�~샖�OԪ�w��G8;`x���F;�~ݔQ��f�{� �S[}��WE���["��vj�Y�陸|���f\^�hX8Y�� ���4���<hr'(|jG��ڞ��d�����)���s: ���|��0�x{��VW`��J���qT���S�}���wZd"�+u�L��c���7Pf�6T�ua����m��Q�e��Ws��P@���T��.*D �LQµ��|����F�Fh�|i,��ց������:ϛ(�8rC��X���ص�'�2�E<)�z�d�[�W��m�&��鴥Ѷ7pƓ_�t�ߡ��kײz	P7Jd�@ ^�����������L��Z�Z�U��K����,��W�nY�wǤǳ�L��d�q��Xz=�����~"n�6�s��Ws_s�V��S�Ae�����Y�R���-�|T�w���SU�
@t/�='|(kY���m殖�cb��O�l��U��|�틴8���H@�1��}X��:r�� ٠ټ��!��%_�h�j.u�uP�GQ~0��rV��v���Hmӳ�b���3Y�R��0���&�d�����Ix&�����+3�P��|���v����c�v��l���^=�z��5�<W `�j�JQnBh����v�s�?��a_)"˻�s�����ETi���|I��yyv>S�A�I�,���BS��xa����zB�k�F�~�i&+�+/��ͪb(���3���f7V�L�f��=g���?��|�E�F5�3�� o��
����\��R>��gk��E0���~익#?�H�l_���ӥ�V<�2(�fͷ���o�U��]����B�>��#��A+u��54��_��8.�]���,}%�����Z��U�"k�9Y?�M;可����7r}̵�/C������`ߺ����*�� �c����J��l߰%�d���M��B)��E��VX��u�$T��-}�<��`,{�#�X�mg�2�T�e$ے���2xK���--D�8�3�2�T3��#�&<�EE�Y7	�7�Ũi��æm��-�h���"i{h7�W�w��-��? ���F'�#֯�[G\ǭO�.�/m?���N����$��X�Q�`������S�i������&LI	�n��.]�R[��3��@�E����@֮%|��s�}��ɿ����Q�`3�RoQV����c ]��ʼ�v���=./WA��#�ɜR�a�X�3tS_U3�oW̜�ã�͈�#������%n��#Ƕ�)TLp�)�s��ǉ˓_Ϫr���:'�£�m�|e�vP�y���h���#)�z��ђE�g�I"h�t ��8`#B*J�A�.R�7y�����P��TRQ�v������=��]��AI�1<���S)��ރ:�N��H�}�N��x���=�G�g@X�V>��x��Xp9Qz��v��\�ˍf7�ɸ�]h�K�<)����8��7ⅳ��l�X0��Z�Qӣ�2-}Gy�H�!쉜�}�x��A;B�yq�h�AA���C����� �Xu/7R�����?���Y���*����C�e�u]Z�z�1zmt�7�V�^VT���ȧ/��=R_�$�'\�������e�T㬞���(Z;��G��|����z�	럾K�`�c<��p�r�cV��Ӡ�}8cxA��z�U�>@�j�m����/"ͳ�_����Z�:��Ow+�IN+i`���9�m���C<V}��\4����L�h�J��k����YH����.r���S����Qk"��}E�QkG�����]:�kb�G�<3I3�b�7�SrP���C���PZ����N�iq:�J�崌D�o,��M�Θ�u)-ά���@޷��S��Q1���[UV�$M깚�P��o͒d$�n�ç��)���%������L��i��cw�pol?��+~��Z��0�%L���Mݘ�5f�+�/���ǧګX��I�X�Z7��}����(sk�F���&��@�<C:!3V)�5$�Z;Mq���>-��q� t�gĄc�aq�N,
ݎ�L͜)T����Jн�0��]3.��'�_������(����n��.ȃ@�5Bq!PNo�讹K��D�ywT��ND��\�G�Q�W��5Xp����U5�(e�I@ȑŭ(��\Rct�v=�[�Dbæ
(��7[A�H�0�;�4���?���	<���ػ\��W�#��=�{t��2l�/�?�m�l<1!�h0�:CΊ��c尮'���1��p��d(ٽ����̤0��=J�EF�S�/��V��t�~r�8