��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\�#��t"�9��͇��<��]��翁"�+g�3]Yr�Ǆ*�Y1Q��X�с�̅�z*��,���8��]��#�����d�X�uRK�-��^�W2\���8fN��e��;��X��PM�}��Ǹ\A�2V^b�q���vorfk�U��'�Lꋼ�k��/;�JNZ���bSpPߣ��ɄW�}~^���U���cz|QQi�:Y�?�"4�۽��[zW������
�������!��5.s�q�����v:� ���f*�}_�_���vogg��c8�l@m��at���{�WN�A��������z��ܩQ�Jh�Ա<,E��t��{���u6���u�V==�Y��x�M�n�`gp���o���Z�ry4���h�hˠEQ׫n|Bn�ʠ��+��)�bQ��>iã�Nƛ�����:�J��z�458�N��n��!)Qc���t�8a��w];����0dP���PE�=��3N���>F9��~��Tp�!��f��4�~���I4����"'g/&O�-�4?�V&&�vV+�5�	S%yrҵ[��ӯ����>f�D	Ex{%?Ɛ_Yz����w���1���Kse�2��3(���^%��J:}ITD�y&]�0��)[���ϡx �M��\b��Z�xb�{����5��;̍>gs����ov��3hjr�xR-4�Y�(�]�5LE��}<�"�����1/���JP�X��k1Y��+_iy��t�E%ƞ?�.��㌽.�:EmⅧb��ۡ%z�DE�-��J�h/���O��vc��ZLz�$�	���8�����t�N����<�{(���\���d���}�rk�1��<�����I���ZX�����ݔ����s��u�H��>��
6�S�o�XvLu 9�}�W/[<*<��xjLB����;Q��Jc����9+�pB��ۚ.�1�������=��D��)~}��M0�V�tF�R��K[/������q X�rp��҈��AMKTuE���r%��\���CU7�� �ry�\w���#թ��U(�����F�o�:E�!g��)\��@,�����9H��(J@E&�1$���b�T��@#��p� ����rK���"������H���mz>��p
v�0��i��{F�s�����<���(�_~n�nNۧ"c��ׅ&\YicH��bB�^��pnl�o�̿o#�[���;/�y��Z�⍾G�j��܂�"��=_)l~�P,-Oӊ�n�X`��+���on�.��Y����<�遛�-4xqE�9��q�c���:�r�����x�j!T��mW���9�h˅�2�O�ܨ8fN��S�O��;@X�އ���	���XT�3�ufwvv"�1X�Q]i'T<�f���S_�`���h�mC�U��#�i�7�:��H�Ru��"$M�d&@�v�L�'�s�{9D��fT��`��<�a�?�(u��V;��%9���s�Qݬs2� >���A0�9��J�asu�(�7c�~� �l�$+�g�������~^"�`�و�������/�=|h �f ��	[˹PE��"kr�(���| o�ޱ�ұ���?G]s�O+.�"3P,�ϑ����Wr-kp3�����೬�^�S?���l���;�Y5�4���q��3�\���<�Q�1������C�a6J��|���R�������̋0���Q
�:W��C��4�u0�����o��T��}u��:�sA��3D����$�(T�s��S��ʺ��������Sbɘ����]G����p���Sq
b4�[�MG#l�ZY�	O�Y��M��;�=�^��1����� �?2/d��k���œ��Au� �N�_��18���a7�$�2�$����Z��0P�pإ*4�a�f�D�MU�n� ����`�eOi�xW]g,v��"�=���K�@}�s4ۏ��Ӓ��0</y/��]5��;��#[K��>��:�J��]�Mzo���)��6[�1�㔲S�&��@��P�R�a]�N�Z���\}Ǧ�-��_ �ȹ�MǗ�Wzф�#�lG�F�0eP��z�B}�@W5��oQ�A�{�����ޤ+������$XB�S�z�^����ϰ�%�)��9Od�#�֢2�I��>�a3ӫ�K�`�8V��?Z��e����\?��tŮ�D�֫ɧ�,_�k J~��_�>o������"���և6���Ë���s��:����������Jb�ɴ���jd��}ЁA�[��4��xL��?=^G��#��!�Gov���'���iK���/��P��^��kb��ޚ�'���^r!������"��QL�g�Ἥ�|Xaɍ�j���l�s��&�{.2~}��?&�f-�ad|�N�� ���$	7��a2q�M7�"u�!��BO��~�����z�U��3{�Y�(h��y�6�?-*��V�� :��_5�K�^���8f��_W��Z���q�r߯��ͨұl��`DɊ^ E`��c6��S|���t��Y��̒6����P�����	���~]�&�1�C��5k�b��{���ד5Z9K�G�x�ʓ��W����
��r����%>�*&�ih��{S�T^�}���7�����#8��DJ�T�����8�SOe5,�t�ڷ�f���b�A��S��q��ߙ�y��� b($:Cs�4��'D�; ��� 	Mk[y�����l���/���«fy��߬�:�gsR��GǜTޅ ᵖ�լ���V��3�V2oJ��Bx��h9�_/ȏ�Ґ9�y7�H�Cy���bHV6��:���s);�X��9Lkˊ$~6@�"2�@J`�@&�Jpp�Y���BUO�E�m��i�by8�87���u��dq8�U�a�)I3�6�Blns��$co�<}+j�ɾ{ 	Q�+w韘���?	�,���� �(�w*���1�̛���)1�7H���n]�퓾�iލ�h}�j�k���_�@-�o���F�ˤ�+��������UP&A���"IUW�WL:R:j�0^�v��J��ՁLܥq0�^��~"�$7��}(yqc���mE?���:n�~v�Q�$�;>s#����h묧[9�j�
�h��A�(��~�X'&��7�����?]�p�#��{IY�m����8�b�WE��:E
-��Bf��+�C,�.�\NeJwy����DvC���[vW�$h�"�� ����}�Nbqp�� ���*�$�ZO�Ac��yu���s{���s����8����[�^�Lsy">!w�p[;�p�7�hntE\zw�rҚ�4���r����0oKby��Q�妫���[i�J�O�=�W%�A�?Xt6�7{��r%hB�i(2�8�e�h�Cۤ5nڤ__+�,*������g�:#��h~��<d����Q� ђ�,�E�p.�Դ��a댛g�#�?W��[���DC��U�nB�����%���� R%AQƸfk]ې�9*�aD��觇��c���hX��aEt�-_@�h,�.��< �����ɻ߿�E����{/I��~s���]��\tX���D݁��7r�3_�
���m�킃\%����_�Yo�<1�p�s�������#z�[ƣh_�aGb��ù���UDr�!�kޛ�x=����F�T� W̰P^�vv��͚:ӄ�&P���.bK�e	���=�0��H�E�[�u5D�G�4�Ņ�&���cZ�Xx�(D����U��
�W��D�*\���2�� 1�8�z����]%���gd$�\n���
.�8�i͚S��0%:��cu���d����l8M�YX�����"&��q�1�O�Vju��i��sS>sN��L�O㲢39C�>@꾂�� j�X-hKʤ��>[M���%�3�cs�0�{��k���f/���-#1��	���S�y����o�ȵ�'L׾�`��Qzu����K�V��¢�I0�X�$FEF��ě��������ݐ�X��AlJ_^��b!��΋��w#�~�)�]J������)��~��$q���!�͈�� ��0�DI��>Y�n�_�w:���Vɜ�7σ?�Ē�&���7?�����DZYvRy�I�Mx|���7�ȅ �Y�5�2�,[*BqH5$�ʁ�AOE�Q�ん+�0�x(`��I���5'�#s~&r'���P���sg���q��:�/�i.^�Wև��f��C� �g��j.��+��hx�h���� nnM�}.3�WS�T3��ֶ<SYrZ����71&S�>�$C�:��/au�X�c�{���v@��翘3"icGR�;��"���MI����cx��p4���)��{@}jo�hrI��WSwP)R��HV|W�0
�
/Dk}�n��j�:^t���C��� ՝D�a����Nne
�#WU�cAnR	�V��^;���M��l�y��_8}��f�u����2S}VN���&�z G���#�y�j4�~j"�s�v�:��d�M/�h�N�t3�=��Y�Z��= ���r�
����y���~��W^?�&�h��ڻ�1.������Ŀ-�Z~x�t[�K�7�ş����\@D���/i�|���{{BN�0��ߊka��@�~�}DO`��S~�q9�0w ����wR���#�{LVO�ɽH�F&�Ԃ��ܥ��8���+�n|S������<��GAh	�R{��ka�x��|q�s4�0z7��;�M�5��*�,�L�u�Y���򑿗�vctH��U"��+���e,լ�UR��W\tZe�I�&�,�t���,o��>�JJ]H�ha�5Q��l��N�-�$�;`æ�����Z���g���'s�e"�އ�Ӓ�C{�}ٴ�"���U.���B��K����:���xIݝՒ���N����'}��Ȫ��s[*���� ��]�M��I��[�3�07
g�1n1���œH��:�M�\�p5���K��c:���yV{2�/����h��SĴ�#�|���A��"�(NNh���|