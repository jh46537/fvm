��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@�ԍ! �AoH���;yE\�U�S�r*A�*�脼	�f>ߏ{�Q`�qư;P[��a]1%�Y�f4�ހ��8������]
�F�VϘ�+-�X;��hM�D���ݟ&�"�\����7&L+N7J������mlD�H�+)\��F��������<��,̆��������X.�^��EښW���y�U&�)d/�O������n.\* ��A���Cg�<���\�����q�����{�������!A�'�"Ť��U�vc���S� ���̕��A1����He�S�1wJf/�T��Xi��q_��� ��l��+8~��JH�����>$�\1�������I>k�Y��TS�a�-u#C��_�������EC���n��o���9�y�؏�e�t��]G�
*�����&�L�{H��6:��O7LK��wD��0����0�+�~m� [Y��O��Ҥ��0?��>%�4q��$�b,x��&>ؖ;�u\ i�Fx�Z��CmuM�K�K�y������̠��xe�ǇBο�~j�ć�T+z��e�r�\���~��D(��2�۩Ճݨ�uaܳN�f�K����v��.fm;�<�R����~}�\�����W)_)T��<��ՍF'f�\�Ə���rt�[�42Ox���[���{t�$��.�Z�1��7V�Z�ە /�>�7��=ɟ����Z]�ӪA� y!٣F�bj{�c�g��CF|�?^"j΁���1�������o����gZ�T�)�)�ӛdXx�9`����}yQ�%;�=b�QL{|�t��38U���U�u��90��"ӶY�Z���x���F��m���v=��5�c<�EZc��(DP���P�G�b5�&̧�}�z� ˬ�`�<���f�0�^ז��Ԣ��3�ZSRc�s��g� 7Zz���mw2_�W��d�O7qʲ������y���^��G��&���a��"�y���
a���\�95��������G�.�zKFߓ��W:�,� ]?��$�<hS���5�*�y�n*�R���p].�+���nʀpKv�'ҹ۫^TiW
��+��s+�!95�\��$V<�@9�!{֨ZM��+�����9p��BY<���W
�#Z>&�b����Ȧs ��G�̌���i�E���2��<�O'?S�����{c��ƙ�����G�ɷ��Y0���b�
!Z	NGGF�e�{JO/��Ռ�,���s���J��o��2���v��'�>u�?ʻ��Xs�<��4�Ԯ�m\&��{#��ԃ_O�>��қP�杪�_���ϰ;�w��壾�I���"�k�Yԁ9�<8g0���p�'�=���G�����+m�T_�掴(QKtӽ0ԅ6f��9�aZ�XT!��/s�9e�ն�E�mr�z�`C���˼�b��m�Ӝ��
T��4=By�u{
����74��*�x&�_�d���$y㼃+���?r��i�(I5�����i�X�DɌ>�꿄�-?c4xal�O�'�,���t{;8���֏�+��Q ��pl.d�6�sS���š��A�cHZ��6��RNc)�@�D�yp��}�U���BnO)�"px'��o�ϴ�{��,��Y�3�EhX;�!Ш��ӑݵ[�J� U�h�i����@5�T\+��u5�CK�M���,<����	�0@~��˧���C�Ŗ���@n4*�O�
=[�_������}k�6���@i*�i��͐����7aH�9+gΟ�N3 ����Nq[	�^r�y^e,nΕ65�S�8lE/䘝bP޷��g�3��6�N�Ӂ�J�T�dꕁ�[�u��^4.���Q ���8�\��{G�;i��w��%~+x�6�(�m�MG���x��	���~�����g��y�U韹9Q*�g+
���N�w�Y� 2�Y�s���v��5t�o�A,b�5�rN%9�����z� 䤼�m{��u!�+�M�[��ׂ�%ևȇ����ղ��p�T�b�������j���!��-l%�С��m�K��(�qxg�-��"��
�NL�]9���G,ǥ�E��i�^QD?{hѹX- 8�Dء��?�X���L�hQ������q��s�A��d� Ϙ'ӳ_P��q2]���f�Ҳq��0��ꇋj���09��P��rQ�5