��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	���uYC�т��秤��sy�/�F�5�
��3��X_��͝�G�����	����{e��F����_�������L�d:���y�Wv���y�(r%�'S���v��a��w	wؿ�@;İ�Z��P��B��@�ﭥo��^G�!�ˬY��P�PJ+Kiks�C�EM�	P8c�_��wj	��Ѝ�w��N�r��F�2��V)<���m�:ճ����Q�4ǳ��5�*w��b��L&�M�&5����b�Y6���*��_M\Ɓ���p�>͔v\��miǈMc�.����ZaP�	�#)$|�I�&\�X��uC�YG�&�e�?[>� �ժ�
QXp�?����IT���!�#M�D&�����(c-�=�yZd�K�A��W3���2h.i�8Ae�2j���U=���d��^��3��HL)z��nJ�,�o9�
����P��҃��o�fh"�ƞdKe�ݻA��S��c��(�-���ή�� =\D��V��Nir��i�"��3-�,F��{�k�q��bG����� ����M�>|�����i��H�ߢ��n�]^m"n���c�;CP��ʽ��B��ͱ��Gf[5ŊX�UV�r^��cc~)��Ʋ��2uo�FeiO�-��԰b�D�운f�"N��P�F-��ү%TNA�!l����8�O�*1�_sR(��D
<λ���S�,.R�b��O~��a[�D9���+�j�V$@��gj����u��=��gN�q�*�+�\<��4������SA�d�|�ѽ��h����[,ݒk"�,!�L	��9�G^'N���뻵:02���g_]6�X�}���K$����v�-�O�,�����O}`uO�ꐰ�8�� ��I��B�9%9���r�ѥ3Bx��p���&Qk.��3;�75J�-Y]��n�����v�a����[��A��>�\�`���^�s�e,v�~j��-���>4cgMHh0�2������4���d����WK�£�+��q�("�c1�{�ꐇ���(�_9O���%i`S��#Ct�}{J��EN��2�������^Ƒ�#�K�B��8�d��;�PP�eT�E�}Ys�G^d f�p��a�p]T���ƌ���o+�m\eN��1�"A���nao�Y��R�$a|T%^I��C�^\�T<��DB��R���YBw�`��D��[��ԞV��&����ᥲ��_'��dv��A��c�ak'* �#�z��LɬC�
 j|]U��a������y��@������䎈��/ӭQ���N����8	h^X��K���tc��:�5����/��Σ�G�� t��a��m}kl`�FB�&]k�5ӿ��	�� �j�Ei,�8Y��F9�\Uꔺ�_�+�)�a<�v���S�3s_JP0���k
�l!�X�I��]C�m�P��y��Ľ�I�������̂_�ˊFj��Cv���0�y��b�C]F��c���Yq�?�)�|�_�Et@7kM���<?���;:9��f�*�� R�͓�z���y{/(˴,_{&4�䜋-nv��#�\�$(��
����e+B[ߥ���T�`O�%���
��K� ɚ�W9����9�! �@�����`��M���V�B���=ې`�O`3 �6���VҲR@�v�DHx�M���<@(87�iry�a�:[VBd�GOk%�Q��ׂn�g��&��p����&�	�)}� �5!�M�2�g��8Ս7H>��&�Odj�Qz����	�R9ki�K!�V#^��-�X�����&U]j�x��zO}�2���#u@�����Wu��w��yT/&��
:��ו�B^nG'}0���I�c������s�(ni/v��F���F#����'�7�$�"O49���ώ;o�2aJIFI]�BHi7W\���W�9�7Y������(:B��?�l��Є�2E*��cOp���S����!�ԧ�P4m�~�Z�3�*[A/Oaſ]�C��R��)��I�{bի#�90B9��������r1H.��m�^��K�����|i?,��V�+,�_=oq�'5� ��G�lmr��Y��<A<Q<��C��y!�|��;վ�W�\-�*`a'��#G���_�N�@v��R�4_ьf:�q ��Tn�Թ��z�8Mz)�[ɛm�Ε�K G�P�f0.�4�d�y�u��.� �B�a��DHc����(v��7C������`��˺ ��)ʚ��[q2���|�3�������)}���C���$�Q'��\Qp��V-Eb��\o"8�Y ��ģ��߳���@P-�`S�F+����n�_��?%��"�Y��:F�m�J�i֕�򆇸����2����1.�鹩�U�^�J,��2F�ٜ��Y-d�pf7�t21�>I�l�rh���ד��V7��`m��M[�u�3$	�hE�y`��W���p�&�rC�Ȟ�B��f�a�մ<"�E��֐�1����и0`	Ijm�V��X�X��n|h,�AW(XY���UcL��n
,���\��N��q�4eX��鹜����t1�8�W�H�i�&y���i����Q�藯�Mt%|2=�6$�����S� �1��}��L�ie�*������j��S��R����y��	�����j7��S���E�_��PY$#�-bG�>���|��6��si."f�k���\��0�CR�O�A�f�oĞ�Q	3ļ�#����;�(\��X����%+)�P!���o��H�S��Jc�����#��s:<B���Ӆ�P��V�%���C�0I�t&�5yg�{n(?��]�-�BB-���Ѧ�.y�,K�������Rj�鑝���Qp�ĠWl��jHz}�0����u�f�����2��M�$�KYH�����虙X�3�[H���cyC2�q�����	 ��=��}޾Ĝ'4(����(���1�RQiwTKD~�4n�6P̠�p2M����F��_� 8z�Y��+��&1��t*xM���Ԯr��-C���"��VQ� vg�t಴�#�f���9�e��P��߀��	��w�/-�c)-U��	P�?!�L�����F]�K�h�bpv^W��I�,+�T5��yH�>絩��W��]�����d���E`�=ȫ�+cV���~ۃs��STɹ����)�id��|�!/&��� ��}�En���e�S�1 dw(DpU�����o�Z`� �ۤ�Ь]�e�I��_/D��+���𚥎�X|BV�^�w(�C>�_;���t���n�p�*B�. d�K�q�i�����`�����rɣ���ɡ���勛҉6���UyU�N(,M4��U�f�����P#����:mI�z\a����li�s:?���$��?ĝ)J4��G���q���Uw���g�e�K%�@ I�̛�6�<��}��ݡk��?(9���+'�����$1��f+� a���l�$��wl.��E3�-���]��J��W��zz��g���y�T���������/�&����A�ٮWv��K�
H[�7)b�{���xS�ԓ�DĿ ���o(vN0Ŕ�S���?D�A�j�(O���e@ɤ�r�c�׽֘��o��C�@�?@D�e޲h�-��
��|����Qa)�my��W�g���K��Eaأ,O�A�$�z�w�Ce,t=sr�6�$i�a)��Al>oN?�� |K����p��|`�nl�7���*�W)���+�Ds>�u����gn�XB�	r�����FYO��<�������Yx	Z�9��b� �^���0]؟$�0�{���ܑ>��Yk��4U�$w�I0l��5�k;WNؾZ���=�{��rvx�xt�����'^���\&�)x��Ojث��@�(ל{��4�l�w
�U��v��r�m�nyp@O�0�HR�t#[j���k�KX1�zM�ȡ�W�#O�7�096Q�h�z� �|Q:TF�y���Fj�<�o�\���S��j ԧ�;�8h�*!�tN��;�H�L�NT�����l_�@&&6���֥	+BqXL��b,Pj�E�"�=���p#/�Ŀ�X���*-Ē��JT� �����|�@�����t��]���;��G
���<�g�$��f����_8z�s��t:~�@H�lη ('�t�ɫ�b��q������;�զ�X����b�/��q��yw�R�7�=��9 ��A���?�+v�U� ��޼F�)�j+<�w�:���X�c���b���-i©�2V�jWA�K�iݷ�^dT�4�Ǫ��X�I���4��_򿏅���F�7p3��l�K���Q���O|�����7Z���Ao��:~��#�kR�Z�b� x�+`�)Y�;����k���;�u��$�b�����o��JW�C�@p3��!`��q$K���^���R*�ˁD{I�;������|}�	³5�[����h��ρ�%ZY݈��Rx��C9�g��>({�/��=�:�Z�[K�t��K!�@B��UI�8�2l��Dղ� 䳱t��E��aN-h���:�Tcz���{�����P}�/R�m����>#����F�ά�`�%bG�5;&��o`����=A�ѯ�/	X���.�DT���W?�Q-�eP	,�46�땕���$"�7��5�,�3����Jv����{��3$p{����gA�H0���HZN;��]l~7��O����ZOEL�	�@'`���G����B#s�t0��[A�5Qv֒��Bi�`��[ۙ�&�Kܛ�57c�z���M+�)�Q��H��GF�"k(+�-�]�s���G�[G" 6w�W��S�pz]��>r5�#\�����;���<4{�%%5~�x��0��A+Ҥ(�l��w3x�����W��e+Dߩt(����>ؤn)��dXL�>{�U|���S��~�0��N���%�nG,05KɻN�≅CN�mD\�i���2#_1���n�M ��1z��~�q��=�>�~:kz���k'n�zu�������T ��ܴl�9J��#.�9�S��~�(8Xe�0��a�����ǳ��< �yR�E{�Ա��9p�B�1��,"������lb�X��D��jdہ�h���9��Eys��f	g���r�Z��"8���:��8s�V�����:F���D���P<ݳ��~/�Pe;�ٍ<�tH�jc U;uæ2?��hJH{��?��Ё����p-"S��Ɩ�pT.��Y�N$F2<�P$��޵�����$�:�@�J���r_���A�m(	u���P��z�ػ]+�$�2���ٯF�8H�P܁�5�����r~���Ǔ-`��5�a��⟅o������_��Utr�D� �� ���?\��Ȅ����E�&�L/�����,=.��[o׌�����I�mE
@I�������o���qiA0�#4R�sl@��?� �KK�p�.	�E�& �X�F�'=�,ZY��\OJ�]:&9��P�������и�?l��zKsA�ݻPɏ)޼�:�C bs\��k�aq�~�C-=u��s��~d��%@��{��;K��9�VEZ&\���M�H_��]�#�O��a�����>���=���?;2�NV���S�-�[hU�f��K�<v{��X�e�8���w���z���L�%�iS��H�a�8R���X�
�mqS��;C�bh�����mm�W���Io3��A��'���>�*+� ���E��y���]Bf�/�fm�<��6�����=x*d�������0L�>w����?����]u?��￯��ZVq+�G�wcV��R�V�r�Q&��p�V�Oq7\�r�odT��2W8VF�і��|�L�N�8�P��6�%�`V[���^r��J�*��B.�&F��'�����謢���t&�>��Aek~�S�T�@�Im<�?��	�^��/lv���e*1Y�NN$;$v�ny<EW�y�a]�#9�{�G�he��LY���-��H~m�ȮB̹�85Ǩ�������z�D1��UG]����!��0 �j�[×��x�}]�.Yln�f!\�z�ra闰�a� M/w)$+q�
͕������I�W��!�n��c�����G�.g6���F7E͹q��ڙ>�Qn��Ŋy��5䒭�@�D¹: �˩��N���2��ۇ+2�(	y|a|I٫��
��d?C���y�	�Hzz�s�x�s3
�/��>b���Fg8
�r��{�Bz�B��<<���O���~�iO���4X߼9�߅�ę���R*��:D���TϠQOX4^��~`5^];�àH��v�*&���dY���ů+si�ԫ}�����s�R�|���M������D�|E�/'���S�E�گ�W��Esr�)R�)�4�$���U4�1��\���=�]��j���=�we�\_�q~?��-OD�5	�a'M
c�-�hF�C��F�֟>7���٥y#�[�,o����:م��y��?ސ��Zj�Ż�4b�]��QY@�&��s�©Kg	�>]��]�ӥy��mQ�!s�d)����������)�������@S���&
Eb���Lxns4� w�M{�8�#]���E7-V'�?����"'�u@����[�Z"�%��U٢�[��yZ:k��@k#������F���S
�;�
'��i��eUX�._�������ҘU^�ą�G*�1p��f�:�C0M+�l9Cd�9z]������n6!� 0��Y\:ʹ�PRu�-�Q#�1��É��(����aG{�� �wu�ƚ,~[�#�u�
�!��R��9�q3?�tD7��)���%�f�g׃.d�P ��~��_�A�w�V�޵�w�%�f��t��"�S[�$�i ���R��_��B������?�ܳ�0���K9M~�;Z��� W����h(��/*H�U@.D��"�My�U��:(|��wQ������}��4�C�No]�LB����M�2���o��Gm�]EwB��W`�yVsz��߼��=����DN1-�/�DE�i'��Q�0�h��0������9i=Ag�rMb0@aO�����-#�uPT���>��A�Oʤ�c���È6ӇZQƮZH��ib����ʊ��\POb��ʰ����m�fA�4';a-���P�c.�j�@E_�?���gh�b�k���0U�}2b���ߵ��r�2��טhZy��7Fa��쉼����Y̲��d�l�[@Re@��Qk�=������ȘސڌLĝx���Ԓ�Y���ڂ\s�!�+��Sz#?KfF��s�>#��p�����7���X$�s�C���Jx�b�]���Ǫ�6�z�6�B8���%O�DϺ��l���3wZ�j��dw �;ib���-+����;�=��T�/PĮh�Έ�r���o��j�K�{�Y;9I���t����P��%M�>I��΃�(A�0(��2~b�v�����͙���� :l�c��ef\�D�1������/\a	��es6� �>�/����lY�T5"���K�3���B�ƅ�����A����=x��TjC8����*�4<����6������e��
�z�.��q�������.��[:'Y:F1���u��b����Zٻ��<ݱ�lh�e���|�=j���}�bER<ۢ�j�o�K	jw_���f�Rl��1��s�:�I�ۇ2�}O�2����ʒ������R5�>��_�����bQ��FϕH�<��⺫�� &P��N�^G��,lc A	n�Vk��n|�m�VC���{<�\��󢲑1�҉���Z���D��|�}�1"�����_ |���P-��jMC�:���lݜ�!u�u�1n�:��Ҁ����6d��D�Iŵ²��yTujDta}*9=��o,5yғ�����ږ�� };��:�b �H���UYof�\�v}�b��c"�pYƶ�q�d�����Y�#�������{\x�>��}2G� l�YK��QL�B��̙�e6����T�^�H�	3�_�7/%r���3��B�s+i������${{��5b F��9YS�Tdǯ@Hܺ{~@�
�9,�N���F�o>I��������U��&�.���\��'���ج.!/F��e����s�F�����r�H�Ug���%.Ar�5x�����/U�_{`�c۬��53���dB��p����z�xN}A�����r,�N��M)Ѣ��އ"�
2R;��;����/�W���B(�#�G!�F/>�Y�,-��u[�e�D&������.��/1ݽ��ۯ}����`5� ���\F\+��)��f+��ڃ@P8�:��2�z�a� �JZ
������8'L/���O+���c�%�xID6@��lR�E��q�����:}o�f�Ʈp�{NN@���5�@Vʤ�Q g�o��9*��H�fH[a�o%]���<�s�9Ͱ�68��S�_�G�$"̢58�X��٬R05�c��T-ou�l�;��E��$��:)O�*��c�Rf���|R�e �lnm��W�O�Z*���p)�A��E�ڢ9 �,9���U�U�0��6�Ml�*�V�6�S� �ӷDd�d���uR_L�����{�~:,�mi�� �9�F�|1�<T֝/��?N!�{˶�<���G��)�2\Xd6x���i�U��	�XN[���n�%j�ɝ�l�>���B�X����vU����oE!�' �0p��)T�� 8��]l�QGm��\c΄wnzR����x��_�kk�-8���A�l�b�[Y@�*_Z'=�	š��wb騼6v��~'��xa֜�������}"g�[�}��!Y���rI0���s���)*i��[O�+� GqA���=8���(��hoϠ�7����k�ML�2�f�R�02<��03ݼ��D��tg�:$���ٺ�
�S ��dw�=� ^���OX �p����q�T��ZK�ގ�f��\^\��oP�$*�����y���V*�+cJD�2�N���P�(�q7�z���P��sԗvx��r�*��m\y����~�k�/Ӗ��w:��(��;�:Z$���j�Z��t�b��sD~��DY����ۍk�2�}��ב0ް�2�Cц�rblp�+�=�i�X��&�<��x�������+��f����� ��bR19d�=i�Y445cB�6Qm��Ok(=���0%G>���"G��dM�KA�;K&Fv�6v#���ѽ�Z�jL᳑�T=09��1��ğ���>�?�,�S�x����L2�����y�Pe:��YI�R��g����}jM�A�WZ�BK��*d���I���I��@�ǽM��i�]_v󭪁2WHԮS�<���5�i6���0�S�e�g�G���
��xC>�&���;2@,�/mI��ְE�]�a�.���Tż�lb��K�C:q����c��	e� 3�dVxJ�0c߰-<�iP0%vH�6v�*E�'��j��m�=�q�H���F��?B��޹7h"O�kr*)y�t�!����I�'���6oe/-�攃�_����P@��OD՝��-�O�~�{0x&������ڴ�M�.�^)�)xs_���b������l6��^KY�?r�k�۲�	����s����@�caG�Q�+̮�JD�� GR��S\�ꆝ����i�-��VT��
�0N}��%�1�,bK�X%�Y4h�J�c�)y�%n�8��'c~���tg���Z����m�|5J�o��,)6K�h��ᯁ`��<p�4��CMU#�{M�o�U�L�9y���'dX��T�<e��)၌u����h�gKd+V���Z�	��| M��
+@]��]��bF"43t֦3��>[�}_��U5}�5>]��|�u ����R�=Z��=E�͇7�U��q[���I�7�&W �1���}�a�	-`b��y�޴���^��ݻQR$��B����I1�D�w�x�$Q�@#�Ì��m{��'#E���x�aXm�=�J����)s3�=�2�'�����w��l�h�����T7�!`v���:rhL�y_{8����嵭+2�ps>�BJ/�tlfxYp����]���Tn6'
���`N�f8|���Gx��v�� !��mնZ3����4�B�c��M�J.�Ax\M����<P(-a���Df�#o>���\a���j{�7l=6G(���{�����bf�1�PYJm�9����Y�x>۝�������@cm���ޘ��ݑ+}s;7��%�?M[]ݏ����.U�i��䪔������e-`�T5�{$�uLY�U�"��9>������%���O��`�BUdY��H���m�LN�[��NfєҽI{0�:����U'+��pv;M��SD?m��d~�c���{��^�
�!�!�H��V����yN	�P�^t���*�=�>��A��GP?�@'2���?K>$���,��o��&rj�~��%�!�/'W��<?���7�bg�p���3�ߎ��W�9�\��snsE��}�˘��L<��G�����p��vn����N�Ҏ\f\3ƹ/n�g*��������A���Oy8Y�K+|R�R����������$/�*�}����g�:���eC�F�0�O��R������em�Ji��V}���y�b큝�B��N(�vwo�e�ն�U��lu��p;M���}E���o�hE 5��?�X���6oBT��U����������\�[B��4��6����[���r~{��3��߿#=A����H!���\�b�y�&v�w������2e����t�fr��|}^��~W�>c6���vP�m��ZQ<=�ӪXn�.���;���K�oS�r�O���К��������*(C5��8�{K��ឡ_OE��f����*[~ߒ.���F���u�|��Z���|�P��ہi�v���n�������%�*`ͮ&�E��d�C��y��'�oB�Q�¨�,�vԼ�n��<���#�m�X�Y��żI0���v��!�:_x������8��yw%����Y�����Q~)N��Y���<�=���f���!��%֩�/�~��n�"�߂0�|דi<����s,B�z����H`�W������<�KU�z�T���N��°��g�_WݳwK*�ԓ�g?����������q�@ ef���A�5"�lټ$�t]FsA{Kk��@��ҿ�á���N1kXQ�v�q-v�pg���g����p�eR3J��.�}�����7$�2B� �	�x ���3�U%uH�U��e�v[Q��k3����gR˞س,�t��|/�������_��t2M���F�6^�ysU2����C�ݪ���x�$��T�GC�vfz��}�c�]���)���3���PO� V|�v*�5��g�4&�[9�6݁�XGl?h�m�Ο4�z��Df�>��-�P	��rG;��dT� Km���e|0Zbc[k�2�ʋ����DH}�'u+���d,�@U{M}
�j�(�Z(.St3m�m2�*Ii�c�a#�)��6t�r��Vu�I	�ڱ�姴ý����v�z���K��3)��c9��Lt\4ٔ�>Ic���h��Y��W��O��_�X�ǧ��I)^dެ��������U��k)Tvˠ�qYW�k6�,���9`4�p�.
ڵٌ8D8��-T�1E7��~�{��)zE+���mw�8��l���onڟ�&?I�3J$�8���_��<dM\W��\#�����i9⭗#Ö>�|w2�>V-����7��)��R��b8���/�_3,�����7	!�u�ۄ�8uQis?����X����#�~�A*�|��b��C��8�c�P����L���
��d��C7I����c@^YE�Ol��D�R�.�����ڌ��#`ھ'��TK�d�iMF�MS�(}$����r���NLǬ� ?C���3�hR領��Q<Oh~?l;���tI@ [
+�{D�!�� gɄ�*����}*)7j~ �e�2�q4AI��/���n܏��综�� m'G��7U�O�A�	��
{}�s/Y����@��68O�!X�����35�t*OX��+�F�C��M1K�O��8<J7�6�,�q��I�J����к�h�g��������:��	8�cSk"��	�簅�f,��Ј&�EA��	`fq��5>'W\�Q0��g�P��hG�j�l�7����jB]��gD�}k8iΎQ FA�ӵ�{4�B�j#���X*D*E��F�&�\�uS]��Z�u�Ւx��TPp�q�q���H����M�Va����	��{��vr���d��D�-fNMe�O���ރ��n�P3\^�0q���vr������2��Ʋ�ţ;���f�i)姕�3k�r���	��_#Wp��G�������T �J������oL���&��b�k+ �b��?��?v�i"4wܚU�.�dO��{���Z�0�&Y _��v��Lƶ7��w�*K����/�4��HK�~��Ѱr����0���lL='�+8�cĊ&� �V�hgw�uAWl�t�nu��Yk�j䃐���,�6��Z�\,F?���T���d�ӟ����[�D����w�Yg-��!�sh�@����N{�(u;�>ud���u��I=e֑xW����B��;F+d�Jpɒ:��Y���0غM�:!����Y)�L�h�ኙ�Å�q�}�r�W���RH����Ŋ�t	��2>������.�h?�*���3����rZ ���dO6���p�S��9,�#��b��K0/��Ց�إ!�gbu��|%���L�%�2�d��u`�����M����^
������a_͵@�͕q��	k_~R�пE�/��8�@�BWN��rI�p`S/m���ni�I4t^��i!�T�:�ruL�rj2}9�C���_.�vb�Q�b�3d�\q�v��`e"�Qf6���~�hb1̴���SW%0_�&��L�J���Ex�A�l���-�e���I�~��y��6-��
�^���};�����V8櫾�Sak=c��[z���,�1ǻ�a�����pJ�C��Kٖ�X�&6��2�2�;3N�r��x5���C`��������
yh�#2���tr-ܰ`�(+^8���p�Ͳ��i�p�_��I�#�rʅuA�c���W����9�U�@�E�Y���Э�)�f�g/���̝�oZ\b]jf#�� Q*�4��!< ��)7��P�,����9���֝x�{�R?��\#Gn�~�Y��yJ,5_�"��n�������ugǢ@�1PG����S��_�u��7X��.^X����i�q��QX�1]@ؕ���	�=�9�^��-ޏ���b�]|�������&b�*{D|�q�v>%X�U=.�X�jv�r�:�0ˁ�/D�w�41��������I�h���	��j��^�]N�2˦���e����Ѝ��EE�uD�A�v��t,�Lz?9���G�!1
9���ɜ8!�>v���CƩ���,��8��fiOԯ���QL$��'���x�(�!0]q��ծ����Pz�I�:⡿������DW��~�����W���_��ky	h^���� ��u��J�L\$�6�[Ӻ1�B���M�D�s
�t؜��1�ª�-��E������4����p7!�Ĩ���g�+s�h4gJ��i�����
{iݨ1ܰ���'$�bx���.F���o�W�w7�pcZ�2u{���巣�H7~�vF*���B�iVڽ2q�������C�"��pv~����'�-SN���R��TZ���$0�4]���3]�� �zV��EР��c5�����J��qu��	�t���Kͭ����[�&>�<ڠ.���P�e��S��*������8����\*�3Y Y��^Y�ȁ��OL�B	gUP�5&4ͣ�<�
�uy>s��K]ߑ�g�����-���ym�1���	���\�.d*�M�!^d`�����Yv����сN	�U����qT��6���V���̠�x���;gF�vh³OYr�9�>v���^O��3CR��VSn=�K~V?���E
%��(���m�(�f�1Es�dq���h�8���%���.�O�{�9���oУ�>��kxJ�E��`�W��ڃ��,��mѣ|O��@u�Sԇy�T V�umTa�INw�9��
�Qe��������b�`���Ye�g?��g$���̗x�Fc"�.��8�D�/�5B)�V`��A�K��NXV���y�JF�+g����d��,%���X?�� v�8����E���O���f�b=
�x%�t-?)n�@��vl�r1�k��`�9l�cb*�z�Imv;R]{.��&Ô�)�5��	n ��J�/w���@���MoK�-^~��gK�Y�����}��$w{e���3
�<��ʈ�%*����/5��(���&	��N�8�U�؈�W��!*�P�D����T�$I���	�2�--`��Nw�Q1=i%h�ī�Mvөi�.��%�Mw01�GY?eir�* #��A����Bm�����$h)��^�#
��{4cM4A��?�4T7F|�D2P�zd�g����m����0'x��^.ˆҊ��y�SY���R��t�坔&w�Jm��O���&��^XS(+��u1~��J}���s��/�H���B�2Fß9m�m�A[I���.	c m8 �1�Hm�:�<���Gi�υ���b@l\郎/���Vuv���G��K�����G�tk��v��`���6�ZD�0ը�������U��_��+��Hk���!.�4�g;��3� ��/�Vє��;Z-�h=$�����0^\y���8�	,�W���S'0%9尺�R\+H�9�|��7��y�`A��^u��Fp���"��!�jauNb�kz�y�%��4G�`�����E=�P�\�DG����DE#�����-h���m>m�h�a��Φ�����M�s������k�1	�����Ԭ6up��j��Q_5�"a'X9�'PJI]4��/�����wg�����q���!�������It��ln��f�
'��n��IY�<ck��r+���u�쒓m����5��|��k��L�O>4�P�
ط{�l��%XAR9+F�B�)�= ,3I8&��[D��@,�p,#e ��f��jRf�}�>��7�}uſr�����H6�[�*�a�����d©��z�r�Q�W׾Lg�����.���4�4�/��*Q�s�b�{'ֺ_�����������9VڤT^%V��^�
y{�3$�Ě�,=r�4�װe^���LR~Ɗ��M@�N���Ӵ&h��s]��qZк�P�����d�W�oT�:�u�fO�aj&��hϽA��;ڈ�{���}.W�C����i�K_r���!�������VZ�^��J��`˞%�b�X�8_��6=��<��u1��m� �h�hr��Eڼi[d�"j�ټ�X��*sc5�1t��ʜZ�r�	C��Z啒#| ��ޚ1�����Tf�v�����ao��v��-I�����/�5�&�3��#^p2��iG@A��G��Slv�h��sq�X\�-*��`7�<�&����pmI�$�Vc;�vA.���[k䟸ϸ��)s�#�DV����?'7"F��[|LL�Pq�w<�,�	�2�J�e�&ד�X����f~l ��H�~Ԡ�_� �@����I\pYYA��xJ�<�䭹��:�`��>��&��	m:Q��u�I��}�~�����tv��h�P�mi��Nz�d,^���I�a�O��]�m��c������`vcԀ���ӏ��C��Y�w-���i��� }��T{����N��,:M�-�ulG|A�ox�ۇ�0S���=��>a��y&��/4R�fwX@��|̈6 �@`�ˉ�xKW1���P�+no����]�g����E��Ul��i3��ԣ�0�D2a�od"M�^�r�6ъ��P�X��N��/:�4,n(2��0���;�7�x,���h4��R�C�E��Ј`>��v9/��C��p�|�¢�O[n�9���ζ0;�:অ7�����8���F�JgX��1�N��F8K��ʝ���]��-�,9�����u��%6z�*�S�ifn��