��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�w�\պ}���'d��qx�Ba=��1�@t�lo�ܦY`f9��GU��O����5y�k�wy5� e%�iHF�K~3��Z�������# ��d|��̪�����PAZ:�;� ��Փ�?�}�F�ԙm�-r)��]���m�V[��zA�?�p�,O�?����5���dk�������'�]��i!������&4s�����	�O�^Ȉ�i�pz���j��;¬q��"�޺A��+NT���2o4ƙb��f��>��[.�NE(���?_�uܴ��M`[�B�D�1k�')��B���=�hN~��lA��F�
RE ���̢և�}ԶC����M��;	�Y䜥�o����������
J!MVj����.�:�ϓ��i/��CtluA7ᡮ�}v��L���2�g~3�r^	�ںEac㧆��k���u�`L1:Ҭw
�������R��1������H��z(�P}���J}dw��9M07X�OI�-{�F4�nWj��V�bz�!4!�� ~̳�xM�=^�ތ����D$�h�0z����C�ly��,���b�8�\K��X�"���-1g��j�&�-s��js��Yl�%N[a5�� +����q��0�}�O�1�Ǝ�#� =b%�k���~��I�gD<0Ghy>���h�s>zDM)1րa���7��HxvE��F\�B��r�߆X�T
 Ʃ����,�.aj��7|�(]�84lDk��{x�����Յ�]w9}��>y�Ez?����e�W3�n��ه;eYs�C�.2��!�><�R��`�e8F�VO�T)3�6�ҭ��,1����Ͻp6YE-)�-3�~�f�ea���TO�1NVv ��U�\Z��B�4M��l�dɌ��q�*m\,�^��a�,�`��E�04!�?}�X /GM-��|�;M�Z ���W.��\}�WaTV~f)i��4�H���ʤ*���eQ�}8�2����s�eXM��Ͷ�C��ˋ9!�N0�88p���R�$IH=t���������c��L($Q�6�f���>jk������o��}.R{��v	A��ԋa�&\���އh1a����	��i��`��ȫ��@^^�,�&:�&�P/�7XF� 8�(�{���$\�,��e�%�A9���OA��S�ܨ��?�\m4t��M0�uTS�mؐ��Hi썕�l��t�u�J�8"���ק5j���������<��@�b;�{E�7�B�]�@���K#����:�i�W�����@��n���0���~�1M eV�ށL�EK���;�b�z�W���!�Zl3��:�r��ذ� �������ޤ�����G��`Mb�ў�����' ~���*�ңtR8څ��@i�׏��Pe�]弝d�ϐ�z�E��caD��Fe����N���0�\%�C/"v�

E׫ķ��+��,�b/�4;��y{��*�#dQi��.�hE�W�H�^dg�(�$�������Xb�ŵTWhl�9��^8b�~�0~W���2�F���Y��_��X��il�4����k�\�?��acv�����3.�\����i�����[?鼢��%�4�菳K����&�_��AH��op�F�\�4����K���#�C�w]3��������Zi��PM!"�tZ)�l���/,��3_�Y�*~W?��H��jա�����l��̆�m����e8=�,���G˅�%���"�$��y篨 �P'�:�[����l���P�5МM�I��t���fp������a���)|I�Vf�Ĝ�\u��f脋DUs�Ya��WQ ��t�%;¡�������|u�;��&H�A��Y68�-[��Ѓ	%s�������B�MZ=t�q"*��R�6�� �M�|v��[;�%L�����1#��:�����nd�K�f\ބF�%E��z5�xs�!��\���%�Ď��Z9n�Ts��=�r,��ۓ<���E���'۩�	�3<��H���c����lӒ�v"K\R��B�CE#ա�tA��T��P��䛉���hUd=$�[怲6�y�Y��;4�|��9m��`\�U;�u�����̯�����[&��!B(#��MD�F������Cr�>�VI���wؚ���W^�2�&su$>]��u��pV眊�|pG��.MV�{��I����J凗��b(ͤ�{J3E[l"s=CAj����πt�f�'�_s�uW$Do�%�x�V��Ӟ�W��#�2�rL��*�a9zY����1ֽ�lW�i��(��K{t��bk�#�V�3%�NsBT�܄r:`�J�P��Gt�z�Y6�� �����fڀ��!1$���ɺ��<o�z��Ϊ��QT��9�&���]���jyH����ް�2���7��%��G�m �୸4�9�u���J<`ӄ:�.�>�@,�Hm"�����fX'X�9V���/ܡQ%��AO��H�K��(�d�~R��1�*��F
��"�Sm��,�a��v�ڌ��Y�y�V�x7?�����G��zcL��&��9�Yg���/}׆�DW�LA�;q|�W�Zܱ���tRF]Y����Z�{�+�ݧ�f�Z�ll�t?��s�'U=������O����Bj�\P�����C^�gb^	0iCj,I�.�mPxLp�I����y)�)�����W�F9��^q��w��[�ភ�Ώ:[Yja�����^YԴ��$�U��6x�G^�{û�/�2i0���s�4�ژL����T�s�J��Ӏii6o*��'��UaL>m��=��X�<;�'��_���D�)WvL��l���?w�����i�����-�Ep=���6��^���t�V��B�9M�4���`�����D�ӈ4������ɶ<Oz~z��2y)"�����\���|��*��
y,�[{�o= �JʢhФ7��=sĻ��O�+��zJ��ΏJ���7~?d�;�q��^�T�����t���T���,u<��]9cT
J���Gp��(���ۙDv8Za���u��k�O���ɽo�>���G<�7_B�p�LҲw�N��?ˌ����]:���n�*� "6�n��� �Onq|��j�I� p�%�:/Ϙ���j�NZ���}��3��A�@�0�h�he�V�Tل;ҏ��>��V�?\���Q�4_Ѵ'7���2�R� S=\�q���	�g��8�)������A2�o�9�G�M�h|꩎�h���SD��m1�r��=����&c@����s��Q�QQ-�>����f�`���V�AVVhvB= ����a��4�z|;��k�K*fX��{z�6��`�!>�$I�{�%(F=������F[��q������E�[^����j[���ș���1|��v�S��q
��
M�?D�b}@���ДQhH&7L%��./u��x��n�u�W�Iɒ��U<���b�%E�S�3]6k�f�2��X��ȌDM���Nf��n����(����������D,V-qC��l%�14�s{�n�(��e��s�֒�S�2�������"�B��fwk��Ԛ-d��`R�l�Z"�c?��-��Ĝ����ߏ�d��1ʔ����(�n����&HT3��%�햰}��+���N���gP��i3��0᜾�]�����o��_�&M3r�W�����N:\�8����ؙFF��0�K}�7!E,�8@]k���I{�"��n��s��M��.��O��?�:���*�]t<��聮)Ǽ�{b��]�S�H��"�D4Qq�C�TC�d����}<M�u|�C&Յ�T}YzPk��f6�U؇4������)`�i���h��!S u��|�uƱ��v��l-I�FO308roݝ��E
�X��M�OrP"���A(8e��$�m�@��0���$�Y`��ө�F8>��)v���� ��S��9���>��̘������!�i�  �?o�^@
G�N��ً�q+�O�ϋ4}oSM'.���n	R����+�P�r�L�"/tE�/�F'�N�S�{���we�لݑ�K��	��ys�-1h,�X��]�7�~��vCؖ{�������1�Sc����b=��ew��|X
��B߻�W�uLj��a�H�0�fn��ٵ������K~���
PF/<�;��,�Wr-���o�x��X_�����7��Fr6�P��*�!�z�h(*�b�d�0RՇ���ֺP/��4����Q�&ES3P<����{��%���J�dLq��ɲ�"''5@���h�Y�v���.���z�À���S6-[֟v��g�@��a��?�s���TZy��V_�6P��e�h/���b��
�rKOOX�)aD����ʛ>�j�f���խ	ě�8B�s����q�ցt��x�����7�Z��vD~ܒO�/��?|�F������¥���|x�J�:��u�A_��/���D�5xwu�M�Ȣb��%�쎘O���_��8�Ic�i���Ʈ�|=sO��ɫ�-�s�Ķ�N6�Qٻ���teRq4r���L ~�Q5"q��4
U5c^�6�r5.�2�jxMY���f�i�~�6��@"���4��6ؽ4wk��v>�ʳ1���ǖ<�.�ք1������*�� �G����G�q�]��|�H��o�+������f]n�,SwUrXo�[���,->��%&�-beu�̝�{�,��5v���0�Q:7�8�U����lp�J3ъ�=�����1�l����m �e�����d�A��~�bB��|�e�\_�yMQV�G��ؓd]P�"-j)�|� u����1���] 9�����Fv\�M�ǂ���h�#����16��<N ���:��,�e�)��d/�%S��
�42��[u��[��i���Y
:/���9Գ (� "s=�w�j��/b�b��sOipx��ga�e�`�C��NΫ.n�*�xo�i�QxD�"Ee�<�l8��?�q�+r�K��$��m���9��ҺzD�"ʚ)����sR����ݧ���zl��oRj!6V��O�y���wU�]84^���	�P�qRV��C����Ö�9~��hJ˦� ���*\���P�>n����2]|׭��2)�SV;��}����q�����(���mէ}��!�z���]4'�t��m��p;Q'۵�,�ٳ�e�,�h�������&�p���df'����w�
ꈶ/��&$l��bA���+|��ɢ�5�꼔���m��D2ݺ���B��~��>�g�)��%�h B�u����0��+�P�C'v3��sq���4(e�`E�d��� ��ع����^_2jo:��~�h�q]����t5C��-{��R����#�p��s�H,�1z�"a�r?a3F�úx<7���"̦�Ĉ�w�J�"u3	F�"i(`
y�u5[�z$��4�S$�D�U3��d��^�:%8�T6�J�旵��*�
�����]��,Oꠘm�'fFv5�2Y;|�Ϣ/�l��Ci��l�P�X�C
���69���E ,B�
fӭ���0��̨*c�|����W ��FQ}�/мd��Sm��1�Sٵ~`,�ىY��l�(��3�q��z��f:�S9�A"?'+60럟���dzr�����dt[l�Kt%;��d�M8+)��s�uy<�q���/ґ���[z4�Zu}�%i����h^��ECdi
RP���vHEi�� ϫ~.K��F��o3PMe�K	�o�����H��D=�ZId&�K�&ݴ�7�?�Z�~�~�����K�^���U.��Ѝ���t����ıG|d{&�m	�Z	+�91.Kh�!��t?Qd#��֋��y�h!���MmQ��v,NLҼI[��!H���ã���\
Qߵ�f����h�幫V-s��?,2�L��~9��ލ�Ԩ�%E"�}?=v������M�o!�٥S� z:=|���W�k?V�u�٪#{�`�\�R2��Eg�u$P�f��QR����G�vu�`���9%�Gʴ��G����ӫ�EKޤ���l����B����adȀgh}�@$j^{�eyXX��F�-�'/N�6aq��l+s��^$���(G������Ll��� �h��eUl��o�ov~�� ����zgKc��� xU��;�B��y�v�߅*_ֱ/'S$��y&��]
�a|��v�^�;�y9?��yk�K���3�#�r�!��4��U��Sӌ�]7�ʊ�X�u��-�I��ɷ�� �����<�挅�+��w5��m�T�(�Z
���BU���_��\4&�3�������� �L��m�j�T�#_(�ߐ�Da��k�"��_�[C�{�	rX���wVE�P����|p>�fi���i+�7��WNC�:Ss����jx��c�\~����d5�\0��!M
c 8�ĩkb���j�6@�q�;�Er9���4�j|5��G��ݬ��|b�@��>��M�x�@	V��QC�~K��٦L��2Hqu5��Õ�)����_F�K���:'�o���I�*.���+�Z�JО&D}F�B_0����Sr1{<9@m�Eqa�Aëm�o�G�5K&^�4���/��d��G��T��{B�+��^��2�����`�*;#��O��31j�w��Sp���3��b+s;\�G�X cNуTh���>A�s������֮��S�@����z.t[Q��e�oA�AE؞��#���E�(��=��%T}:�14�B6�����;�
 �k�<�3e�^2W\���7�E��q�% ���&B�,���$�|��b}�tb�~�����\
��<��!��bc=n��y�QwM�]�V^���"���"n��ͻn�S�VV-�BBB�$i�38��fŲ�+{��xS��T꺮�����Y�5�//�3��a��|�I�͇�C���y�V���R��n�[�	B�#�������� ��6Q���;i/�N0�-zB�E�]���|�C��8�	��J*P�fǹ�4�8���e�A��[�n��ƽ��a+"��5�o�,m��ad-����>���k>�3���gRD"�K�K��ށ�y`��xK(Bg^�7S��рֻ�g����.��������q;y�;W^x�V*�Q����R����H0W��s>�y?h��{A��B�R�����Q���PmNx������VZ��Ԓ��㺠�<Ib��9#�P���ai��/	c-ߑ����j��m�q �!�Ǖ	�ע�J�>��"lSvK�eY� �֙����@�x�@@����)� m�Y�����}Q�l��^���]�����yb[��o{z nB�����������+Á�������`H14�B�m��bښ�E���O}7�~�o�^�rj�X�|W�or`@,J�ʚ���%�{���I$��9�"�+��ʗ�
�|w�X�Z��i���t��26�g]pA*5H�p�dᬹګ,�^�2�n�ډ��B]�y��U�����G�UO���j�h229W%�(9��ڶREݫ���J�+6#�q�����M�GQ*.�KW�(��>�,��&8������_��ȓ�1F)�r9=�WS=e�O���`�>f�:��`�?��"N喎$1�];��s��S?݌��!���I��MaBf!	ߍ�ϕ&�yg�0�-�� ���xԎ�O�Í%rR8��AtX<���O������To<b�r����r;F�_����5$DM$YJs����U����m�?!�ɘ��LW=R��
ܩ�#�k� �T!z�óq��V�
H{yT����[�f��1rOh�b4��R 5S&º8�m�[���ģ�>$��?�fd�l�� 2��u���Ո�:�����1r�}�	�+��v�v}?A�㓹q�O��>~5�x�P\�����-Z�"Z��h��o���?��qa��}�����
�6�<8/���\iq,}A�A.��??⡥����֐%*����Ŗ�����e�I!����8qM������U�L�T�SA���d���X�c�N�� XM)��Zo ж���`qݩUZ��*ĕ����g�a�����A�̂�as�+��A��lC��j��83?"��Һ������M�9�-��RI�Ȏ�g�	��>�[�����2�Y�<��e��q����*�{���s״u�ǤpkR�fϳ;g1�����۽8��V�3XY�5%�\".�	kp6�e���y��;(�QB����2xs��� k�8R�rfp�@~����'}ST�'�����!��l�ΐ��mSg�M���w����ǅ���/,�擁�Qb�^=�cF�VZz�@�^��1V)u
 �S�1�5�8��'y�/��p�A���~���Cw��|C*�Q��;E�F��ۮ/[�"����C��.����N R2	�ξ����6���Kj��B����o��zE�r`�O��6�?}���x������g�%�MG�@���R�������s�$��������iԑi1J���~^J�(~����k��J#�xg5�i�*���ذ�w��)񢎭���Y�M��Z<痟>7']1��o&��YH��%w�xߋ���Y�5��z�h�ʪ��K65�y�h�_S���X*��{��D�����Z"C����O��"�e���r���~�.ws���z����m5s�3��a �(��љ�G��P�](�p��љu�X[�����δM�,4!=�v�����m;-�U����W.���ұ��-�Y�W���>)��<�~'a@J?�"��OS�-�M�+�۱`��핋;�'n�3����
h�:��.�������q��ӹ��3<{)����s{P_��e�L^5hf~oi���������Еv�"���~^(#�W�џl>��W~"��I�ȻFݑ�o��FUoM�U��Q+羔sk�l���6TP�	�Ӿ��D\[p':ݒ�4a-�S�'iO�I2X���h��HZ�S��\�3bz��B��E$
�o~�#��w��wA@t�d�x4���,�(1z�=ggJ A'��R�V�CK���A���u��A�3{�C� ���Yٖ��Trѯoy���ؑ�-Ea�iU��m�\��8驶N�Tn'�+��iM��y�qS�)�t�bq�����Cg-�-���\s�@�ґ.u����=Q��u�@���;F�V��-xz�;f�M6��9M+]�ROG.p��h�B{2�z{]Dv >!��Pщw;���N��"~��
�R�l
���9�[i��P���ŁT�=��=��7J��^��]��E����,�ׁ&��%�#���Y�
�ؔx�����o#�Ѝ oT����-����>w9����z�e��s��z��h9(i��������_���Z��zpϘ��Q����͡i䅵2ɎR6��q�Y��L
Q<�6?����$�PVK���Ӝ���6mr�2�ߖ9ߥ���Nk�bMI.�خ���h�8,P�Z��!,�@-O8�s8 ���,����"����(Q��{J�3�,?>~.��n��n93�q�H+��������LW�C�Ɍ	
%�mD9�P|�v��_A��,#/��1�&\?_��`t�N�V#���ƊC�t�
�����鱼U;W����M�_r���1��MS��)/���'eN��'�\B�FW�d�j\X7�W����7�ڔЋ�lF�f��(��e���n]\��N!O�bB�-�=�=�G�,�Dj��˨<��r��_��ײqC�]Jr&�������R]EE\n�X�7uiW b8�H�p$� ��O�3:ץ�0|K�y|�b��u3��y<�o3���n�YV]$� �AP�ku4vF����2��-�xF��?=c7��DW�H��M{m7�� ���M���_�Y��D��*�T��G�W!�ͫa�z�{� ���3��K�Rr�������~�-�L�0��<P�w���{����>��*���u�+�)J8O��%[��X(k&��4�M�yOY܃�3���1������- �p���~u��k��Un�z;��O���u�ձ����ѯ��M�SJ6B-D^Sf�NCo��k���2>: �u�SW2�O���	t;V8�Ef"ؠ�o���� F�Hv�Nc�+�<U�p������jܐF<�Ǔ�$����r�R�9I�ftԐ�h4`b��}w�`?v:-0�����b �3������0F#S�hh������_/��OS �3+���]���R)=5H� �����>Na�5sB�]��2CO#��'۩w41HI�,'#�0'�I��l������&�쀥9(ld��1��O�Yr���y�<�?�6pvn� 8�4ci�������h������^wYt=u�������ŗ��/�MD�������tF�_�ϖm�Q���(�Q':#3�̂�H���-�=��ِ	��5�Դ�s��l�,��!�����u�LPRj���hG�=dFz�y�d�f-L��a�/|֏@$���Ԗ\��J�L��!���7�x�NE�b���D
�Ɛ�<Cf���C%e��Q붠��ٻ�G��	q�X�o��cH˲��N� TƳ��Ŕ.�e|W�."���Få*�y�O$X��ڠ&㖀"?����\�wI�_��|��~�]I�ʷ��4om�Z`k��H3Ut�_��"^{@�Q ]�J՟�z��No�두=⡪ڝw@��*=\,�Ídޏ]�ugr�V�ep~s��ʡ�ý�n�����FXpɟQ� _l��@!5JT�q�������&jQ���-��-h�X�	|�1G�H�U����6��j#vF㫻�����x�	EA���>�*GGW#�.؞���d��SKS��^~%j�e85u�J�I!��%�H��
�Byn�����6|H	�VT/w 9|�6�����L+�Ú��+qe�����0��<�W��΂A���nG���Z��Kx������j^�v����՚��Q��u�:ӆ*�e%�&��b��:&p�w�1���mq\}>�*��a��FGO����
��KҡB����-y�Y��/�"8?��Wa��.y�2p��v�1ꉗ���D�Z1�pE���f� 0#�&���=[���Jl�����GE��L�zV7;��	�fEn	u�kEy�g�,�*S.�y][���}���K`�(�5-E����Vc��"z�/�D_))l�H�7��[����C��]�!Ⱦ��R1��-�߸�u������P��̻PA6SF����x:�;b�g֭�S2�r,��h4&���-��v�S��K�+��.��er^5ۅ�(��w�e#��0z�,�������$r�楋]��3v����U�o�T��v�n��b Y��""�d����� �Yix2	�	'