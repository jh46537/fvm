��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�Gf�`x��*�=��	�����:.�����*��".e�.�X�2@�6 �j�D���\�Y.����kʋ�`�i��T�u	�!�vMO�s\O���6�̅d�86HhU��h�è��)��QsT�E�	���)�(���L�ް��x2�D�r)`�Jf�B�C� �r�K!�[uGP諛�W���g�6$�$`q�k;z���!�� ��;�཈�_���
�>d�-�HFE�R�1��W̜"���<;����fX�bqZ`�>Y����aY\e����s���J)���������IG�ƒ
S�#���u1K~�f絚l�5�BJh��]��D���� =�ם�� ҩZ�@%w/�q�e���ه8!�(3���Q�t�bߓ-�D���2V2o���v}��p֌���sc���9K~�=���!\���k7!�_��AEWm��k���X �>�Bڨ�b��iJ*���������Ҋ�X�f:BVyJ�n����r�����l�I�j���?�Jlk�t�쫭�s���@x)���R���2�)�9��"k�m�R-Dxs����u��rH��3B1���wU�p���Z�n���G�^D�e>~�!�#oc�}
#hsB��r�h�����U�b �1Y��ƒP��z+��BVS��B9򀴹��̟k�p��Ӓ�b�
v�޳�|����wc����eї��k���ق2f��HE��I|���$@��\]!�zr��5�AǞ�V�����V�D����V!�V�^�ɾ�jI{[���_�Fem�0[Y�nY�7Vgf�?��h����W҉�u@���a�'���T=���9-�{��c8�\5�R؏<�����00�� ��(��H'$��!����B.;���5��e��^�dS�ΠӫI�覸g�:�Rʀ��j�B�����8��})K kW��Ë.�e������j�E2X�[��p̙XX�>��x>��ɪ�T�\Rr�Ͼ���ǎ�!n.E�,��`��9���̞��O��K�(=�������^r��Ǫ���B���G���u�V�(��}����;|�苷y��[�d���쪃$b�`V��c�NW~����L���y'E�*V��r^���� }EC�����ͬЕտ�=%�<�Ԙ�Ȣ&�y�n�"�ʹ�bX�A�:9D,�,F� ���#T��³XA�i��s:#�QJ�2y7�G�#2�^��iAR7/rq��/�"<�'���ÿ�d�X�#� ��������S���U���~������M�X�FFnl���.� ��A����$2e�b ����5�B�g���fݏ�cq*J{����k��p�5�!rw$@�J݇U���Im�V�O�V�Fz��Z�s?=�LWjp��C*Gw4�LR��Z�K&-�)9��8�_�Hǯ��_Ĥ�T}����M�M�V����.t@ HG�t�ڸ`:�jl�pz8�j��PkM��ڰ5�Z�u�&_��wI�\���d!��h��3㽎�g6,x9�k��J,�2ݹqj��(`� �uό�A�C�6��[�S*��dsSg�^���C=0̍:���1��&~^/=��g��K�T�<\ۿr��	�]e岅��E�뜯����
��N��9���cعG+R,m�>��,A���8b :�K2Ds����?����q�<��+��;:�X6�T�4l��-h�z�pS��s�v��`!au�Ŝ�ݿ��uP��J������A�`/�Tj�Y��m�e�Zi��N�
��_�*�G��u��˂�M/̼�?����\�޳���+����������Wt
[����=�-�}x�uO�I��� ���f,pt/�cL	U��q�f����M�E���a�C�]E�7�mnqE�Am���
�\¬p��g_�.�!bƟ��-L��c$��齫�q�\�C��������q�����uܳ�Sʢ�����=jK�83U9���ؖ��&Ss�7���y��y6�Tz1ռz�Z��U��Ĥ`ˠ����ܱ���K���𨪲�xಱ]�nw�W����7o� K�di�����G���䵱�Z�N�~d�`����KAG�{)��x�٭��!0v[�<6[��Ơ�y������]s��B���u�3rI��oR�ʼX?���pU����&���e�<^2�J,h�m�T�z���3o�n�eTK�g"@�k�z/ryY纨{�ʚq�8�[;[�~n�������\КR8���r�ԉO-��s8���2�����y�"��iNQ��j=2���uBg��)�~dX�t�Ri����P�C��X�t�>��f�����)1P�Y"�h��������F�|�s,����.H�e!j.��4߮�8	���9{�~Nh�Ho���\����)a@���0�K#���%��M*���Z:��p�pДa�@Xl�������/�i6�:	�{��-+,|�<�>�8^�ʭSb�_��Q��%y���=������f!	c�����q��vF��	�j��㯎�.A|g��|�d��=��c����|�IyOЖ+э5�ֆ[T�2H�Svߖ���[��w��p�s����;%��7�G_�-��>9�}"P�E�;���U�<+{ cCt�iE[t[�0�u˥����+���G)�*�q��Bѹ�-����tHJ�j��?xC<���}L��mGP��E[߶ܨ��@���}j���/�~l���s9#�/����B��)��v���x)��,�R���Gjm��Pc�4�l��=;q9����7ÿ�ܶ��Ȕ�~�H�I�U&�����W`��3��j��/S���':h~$p��v�x��H�dߒ��D�5�%��D<���x�o�H���w���ٮ�.ÊC�*9钵�J�+��;�7a*�x	Px��P{kc�). ��2�+��W�9�{�8��q�����FIt��b"�c�v��O|^���:�z�0R1����5�d�_y7�<����v��"�IP
�q��T�k�N�.�ٷ��� �`Ɍ�SA��醼-ㄙI���B�V�0��~e��ӕ��M�Ɯ[8/.�8"�K7��$_�!�����cD�+!���͎�D������<��ؠ�}�����ͭ���>C2�d�V#�ÎVWy��܀t��<.Y�*�{6y	9	1٭�a��X6�9v��ۍ*����Z�ݏ�)�t�99ր�B��.yw�B�Y 5fb�"U�(�2��8Ҋ�q�wM�6�^$oCe�`Jv|�n0�!���<%&��d��O.��X����Ēxb*j���ڟy�-z�8y.Ksx>Op�K`$�I�6�M�w@�,��	�K@@���
φ��V�����C��Q
 9T`VA��Э	.k��P�101͢'���T���%�oR-E6_*�i�_m_�������� �)��}������s��)N_�&FD�1�Z�U�]GGt˿, �Dw�j �?Ĩ�)���:���o��h���p�h�Q��E:e���$��+@C��ܝD+�0x�X)J?�aӺGs,��w�%`��6o`7I�������u��T�Ԓ�Dnט! ���W�G��T@��������0�B�h3!��6����r�H�&��}�W�TG�R�Co��:3��q ���j~�rهsUm8�]�����r��|�hy�o�ܗ�M��%jӝ�>�ı��%�mE�Σ<���lwG�"m6�9S�x�+�#����*R�TEZXG�љȺ2!�U�Z�)|V��#����C�u�� #u�`��^�M�b������J���4�
����>guË�<d�ٗ�[�7�IfI�FC���o��/�$Ҝ/�3[y쒼������A"��"�f��"��Um7?�&���{N�*�Ga��C�L��%��>Ն�(b5C02w��A[e�GX�$��)f_]�|?7�Hֿ�������C���X�nV7/�B_���x��3��iV9�p�D��_�a�Qw�R�]��Fk0Zl;�?g^�k%ߓ���������w
�⯵hy���V�7����hL��H�J~X�����	r�h��\�
�S2�_;�5�z FIX^ P=��:/��?K��E��z�����`���i/X_<��`�`��q͒�&q��t?�y�3�WP��H��ڻ�+%�+�Zv�j��-і�j^�\��ѽ�b��Mm��s��&9.���S���w��1حڟ�_�f��(?�zz�ST.��X�g3Vچ�� bd
��v\�לh['�XQ��K����w��zr�\�]�k�׋),����ܓ0w��a�\�MwIuR+� /R^sa��bݟ��OǇ�o��!"�:M�GCk�`8��0����I��q�Woa�`ZJSf+�
.�9nJR�$�/��z�����b����^����՛W���C��?����y�ngDs�2�lD�'ʢ�aX�'�X����+G5}�B8����|'R��HL��->'�|	Pi�*�|!�Ej튡��XsNk���#Ҧ2���A.�?�N�Pp���"_K��蠇�.hQ�,�-R:c�m_� !�����#�q����(�*�Kբ�^�	щ~��OQ�Ω-MU�W���v����[6��Vn�i0��(`�>@lD���e�r�~��|�����|�>r+�'���-gOB]��*�t�â">�8��+ErQ/���ŊEg��׌Ӯ���-��V�R~��ȕ���SI����q9y`7��3kG�=�n�U��뫍���y��*�/*� IJ(���8�u�6��U�VxB�y���)��8���$@��hVREEp�5売�������~ho:@YR���(�21^�(�(ɍUȯK��"����*�+|�@vo^���q��5%�}2��6����42|�?�׺�p�A��Ex3�]˗Ͱ���H�K�i���W]�B���=�=@�� �n�~���^��6*-�w��X8���b�/�cQh-A�*�ͥ�nPk�x�[��j�&����p��Ƅ�$�9�Gi~�!��.&�ڜ͆�a!����G�4�����8�F/j�{����u����j��c����dě�ɓ���̷vC/���TNLP��N����]J� �v۞�VY���A���fҗ[¼��{vF�T�2��Hzɫ�K��:��C�y�5�t	DF:����ߖ�bd��J�|~x���"G+�J6$���k��^r2�A?ED	�h4�-�pإ��V�h��K4m��O6Rtm�4p�g���|<H�7����Y,�n��S*�DZ`���5]\]�O%�`?ۣ�G;�7
��|�� �S3J˕�Y�7��0���E~�hc�`88ۏ�D�Z��A�1�ڨ:��I�y�>Ÿ��P��G�yM۽����n���� Wz;���H4�XU!2S	��j#e��r�J�ԅ���D��Dn<�OiF�㫆�Ŕ46ӻ;��ֱS:�C���)��P҂0z��f�v�����Г�A��W%��*}�2M��M��DKY��Ԑ]րA��G|7؁�A��~]�n{�I$��S����<x)�����di>H�,�H �*�j��+h߄�Q��ň��2r_��;�,Ї��>LP�i��3�l�X&�����w���0�{����kh�C�ǳW��|��)6#�\*5�mrW�\�]�ݵ/��Z�KЌ#h&Z^�������<��y�������b���MY��%2���7�`�h��_�7�:��#��kőm��f&R�VFj2�?�ŇAh�e[@��s���[~<������!CH�a�s:��z���FG��^><����ڔ��2��m���Y0��4�� ��tL�W�0$T��1���w�͇Ix��w�H��w�J�T�p! ��:��e'sB}�:$��]�np�����mү����P@{����&\e��� ��������NJ1AX��Ǐ�#��d�)ʣ³��4�!�ߎ1$$��&>�����dʥ~J?2|�Y&���@M�m���SvNR6���^�Ƙas6�[UĤP��t�Փ��|�5��P�n���7�T=����	S����[�9��Z����/2C�^t��m_���*�o���BU�@�5�~�-,�A��d�7n�g,r��2��|�^�>�	�@�ʉtz˓$%H��o�g@kӺ�u��i��2.��y(��r���2a��UM�H�r8�HEX��;5�\�;+�UL��Dx��m��n�ʆ���S�e����0|�}��>�A)��+�ɧ��+7ҫ����<��	�j�+>VӮ�:�h��6W<����8�[d��8��̔�`���cG�R7+�V������]��~�?͟E�����L5q�(��Ak�t���+#�0�K���_���dU��򬒛sK�K��:��1$��OF�"�=G����J��l�:&�lߩ+m�U����L��,a���Z��c�=�E+@�g���J�������S�$��}��; O�4	�{QxR3��+T���8�"=�`� 7{���8#�
���+n��qd��+������Z8��-��g��y�#�>�|��#U�_P2z�^�]��� ��%;a��7���ϗ�h��^O�be$�N�i���f�I�9@�¼8E�5���}�����g'{��>�iaU�
�{���Ǥc
�x�O�4��9bV�O:����I����z�!$�4�$+	ݍ�t v�+�� #O��zL�k���.�4V���00~�3������ZIR�_Z�(�B�
W�>:����g�7<����MadȻ�F3r;�/����ZG�	gK��^�ԤV�)�s��N��F"@>��P2P��n��w��7oc��rۗ���;7���?�'�X?��O��R�ez	�	0,ar�0z������B�[�~_������hc\�`��A��l#�<�M/�h��'�Zhg/��W��gT�\�=��jj�[�hߨ�e+��K�{���6u6�����%%�J��|�32Лe4~���@�O5��"1'�$���mS�!��a���,\x�e`ځ���Ӥm���n�����S���z'�جL����k�)jD��F��_6���%_�S!I�V��{֢���;���n)�� r]���rdĀ&��Q���6���Q*�_��g��{
z�A�_X�w$@Xa �l^�����w�Q>w�.'+`}P�̙69�K���k����i��nJ(��d�s4��?U2ד�=�sٯb��$p������Q���n߅�v�s"�"M�Y�f1��:Ows�57q�r�,�u�9��^�>\¼�s�o��>�|�J.��^T2*
]�k��zk,$6.6T�/�Mԋ�5�4:�m8��}�Y�# ���J˘}������}���k��Cݎ2��g�w)
Y� �]�Cp�Bq��$u�JÚ�w���$�-e���f(��C���=��K�Ӹ"�^��VY�P�u��A�F����������i�CY�P���5'D+z�&?D=Y6�!Q�I����o�w�~'��%u'�it$���_�@;@��i��� �aB��݋.��k��
����䗜m��BZ�i�C���N��XȄ=����X��-�졑(������(eZ:D&������E��cb���Z�($� �
TF3�kz�7��'��冽{�gg�	�ϥ1�Wyg�hđT"��h����\@�P�.ؕፄ-��v�+�ǀ/c��t��{!�6�L�3�����1_�*D` �՘��l4�v Bx��Փ [���h���q��7�����vcp�zcj����#N̺C��W�{"�S��(n�.� �#�Ió�IB1�O�3JI��b@m�)ڢoH���NI[������ ��:,���xVcx���?O�0�E
���7�t�`��a$-������.���sG�����~(���ϦE����E�B�V��vx�$�$x�7���%���3����V���`^����[r�®�o\d44�� �/1F-Z~��@��!��<<�ky���)a��HG�i�¢K��PU�U���ON�?Ǉ;����.�L�������zaڳ~-�dQe�_�W��ȔM[Rc�$�ň�>=��Ჾ�g�1} Īg،�GXȺ�5R��k���՟"J�5 	�����3&��cFP�8�Xw�"D�����K�nY��Z{J�p%8m�*��e�����x�uP���|�1ޛ�_��\��b^Q�:���ϼq�:9 o׃�jR��||b��W�P�c���k]b�]X*��F�zB���5i���e�k%�@�T�OY�1��`���(,�o���yX�u*h��|ř��9��}8MMP5��S�y]e�z�sI���0�[ﾰ����z�$�(#P@r�B��V+�w��D��e6���
�<(���l�Ink>5���y��P���3-25���:["���=���L�$�e��&��f�����V-����A�y%y�$3�?`��~_!�!ݏ�9d��f�OM5�)���#�'�.�4���tdJ��8�����Y��x�:��X��L=��9���P@�S˅�;�k6G�L&�����r�Q�ᰒ��z�>�^	��{}ΑG��M��0,�$WlV��g�VUg/-d�Wc�=3����l�c��Sޢ�6��3}�&xě����S�7��D����ʮ!X�N>�u��˓��"��̑��w�%�f#�ʴF(C���i�qIUo*�ENG�_�b�p���0���3���U��
����Jg���;���`�|0�4Y��u߱oz�ِ�'��=v ����k!MC��P6�#3���54���fIBt�i_1;]��%}��|�l��*�M��"��(/|�YA>z��7J��&���m���EVם�ty��H��V�5Gm��	�9����qBa�����5(_C�6y%婤����H�\Բ"d	3����&�E�|�o��x�15��w\N]���E���Fz��Y� 	�$�b�ذ"��a���S���Pa,2�s����v��ҮH�Q�1s�B�i-�$�ʹ�69OT��¹�B��%�!��zD�tsM-��|GU)�?�v��I���4B�'��l��V��m��DOW�?H����H�����C6x$47��Z^���n��Z��s��-><��^���9p�f����nh�:p���Y�I�ީ��J������0�:�ڄ�W2l��\!�9�u�f�4���L�
lg��ύ����xY.z2�n$.&��s�у��%�xP3��t��CHA; X��w�1�%���,nT���fϕ�mUL�L/��'�X<����J�]<�-����/<�07/�67<��8�*⮸�85;���tF�,BU,?i��Qb����� �3�ϒ�t��39d��{b�~E]�z\5�/�Y���Rp�]P�[�Y�ĆU�c׏L���P�
��gI
x�B�曷x�����<��OW�gy�w�>N�$����Go�{վ��R��E
�(���LH+��я��U_W�s�w�d���ձ�?C��[ �5�(A�Besh�v�JF�2j�¸z�٤�(	��F��Tc�Z��판ڊW!S#��U�0��Yi.����2��