��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQG�.�����=����A�\�r�|Q7�V��Ҷm�pwX<P=P��`VPrT�͙"��1�ʡ�l$�.�E.��yyNz�<,���O��2�aor�ZQJ��Z$6VN�C�(��Xu���a�,�F�g�xJ� LL�) �렭���	/&e����sf������@]/�rn�?�K*�#1� ��>	וɹe���ÒNE�@1��:Z�=�@�h���}7a}m����K���B�z�+a������<�J����U�]H��{�b@�Q�5�Hݰ^�<S��cL�Y���X���%)��5�M��Tf"�	�������Nх<
���3̢�|Ǭ�/i�lcP ^	&�)_�*��x5L��Pq���5׸���&6�w����5@��N��N>���C#��ӗ�ږ�3.M¤��A��^�Kĥg���"+@����.=�PJ�ij���"qq����se��	WH���=�%@�}f*������!Tѭ��$�υ:��P/`ci���[b�p�h_a �K���e��kjq�㑀�F���,�@I	�4ck���m�읙%�wdHP��P�{/��=�h��K/>^�c��� a�E����1�P��˅�ڬ���1����R�B���&��D+85-Den?�������.�����Pg�*r1^�j�+���
�|�'{��v�Ե�Ì ��?�6���ʗi�R���W��5,1�`6���`} �/�ܢ�8�9
1�&8�ĥv���QH���a��А�eU��yM � �9�M�A� �\g%�A*��u�x{&G�o������]I��B�� \<�?����,������/�|�un����1H.A��X�
�J��Y�`|I&#?�2�'L�|�H2��T�PD�}��k!�����rj��?����(@-r�6�UM5뇙���Fg��\=h�+:y�}�L��Zt�	�N�&A�V� �4�J���J�}�\�6��ZE3��m���03X��|��9�b�����^�E���4?T���>�5����-�ՆH��pv*o-�J�s.��_!<D|b�=KF����kpW�[�%|Ʃ�_���?h9r/���P�)�eD�KFխ[|ь�F̈+�uS���7��?�-�k�#Zzg��(Y゜N�9N�㍟{�S�V���j���*S�&�O 
�ͳ������>;��X@ n@�#�B����5x���B��� �T���V�k�*�u���ә�l�����Í�,
��fyѽ�eP�颃9�ނ"�,��.;�n�4V�����Qr?UE��F���Nqȟ��#�p�Q�T����y�'�3b�2F���,urA�Z�~�D��Q�.�)�@�ydnbg:ʪ��iU�� �֫�`ju<=�e�� y�G�9��b�mߗ<����P׷�s�ـ���#?�����J���j�5� [��_+�ĸ������/̀DX#'A�h�����^5�Q2mhl���ؽ0
��e��&�B4�T��;y=�	]s)�B�`����:�Qi��'���a_�����"\�����9i|���L$p�������`8?�]�{�r�_/�6��v"dW5
��;Y��Sm����`t���"����,�=x���kp�I�6̸����q��n|��J���(�u��d��>��0ۛ�X�Lݠ	���� Jl��*͗w�Ynz3������Ͻѱ�
&L�8��*<�,9K$��|�R���ll+X>%V:����i�����S 
�����I`\;�w�+���X�dR7����eq�h�a��i�,��e��W�^�V#4������k��'��(?��1|��/�ږǳ��+�bޯe��q�#5���_�&����js�[�&xɰ�z��k���A��L��t�|q�k:���V�[��h�V�oc�mI�u���,%0�1������܊��!NV�qc�6𧚭�#|�N_ %$����-d@�M�ǫ��7�uC�.f[G�d1���b0��Q:�X�'5.L���<���C��	2舱�Gq������uʴ��c '�R�U�k>f1�8��V净�sP��mT�����I�T+~
CW�ShhuL��v��bS�Otn��Lp��|��wKX� 62�<��j~�v�֫���I��4,ԏ�Ge�HZ��.�Y7˵�׉�/�jeK�s��|��vvs�4�_�����ؘk˪�%ꁀJ2�pN�������z�����FܵM%�~.]�&f�4�2U��]��m��cI�H1qƏ!���Ъ.&�Ir��w��m%�KI�ޛ�^̶�hb�����'�0�=��
������Gq��L�!�1rU��ƞ�=&�Gx�5+�tWL��A&�(X@|8~a?�6Nۉ7+���Bv��3�#B���D/�K÷�h[�[k�t���6�	8��
�F'YMI0��.�ɇfO���ɣuq{���|�'Z8e�0Y�����3�/j����b|n�?.�eNWv����a����%�ԡ��6~y��Dw���p4s �FkY)T�����#eX�+������.�a��J����78FD�_�P�	�=�;�U~Z�G�� ��t0�/�Նj��a�8횸��	*�q����
S���}�iA��I�c���ʛ�N܇xj{p�,�xޑ�Ʉ�$Q�{���ZVԹYN����~��;���C���X'��
侞���\�.2��W�v�0�:��0��83>q����wi�>P�]SJ��v��u,��-� ���kTs��ul��U�f+�TaC� +��#�k�H�E&�.���&B���3y��ҙ��C͖x�j��5�p���t�Ç�G{�1�G>F�H�N�7P	V�Ѩ0*��G!S��_v�� Y�
]�A�(�^cWT�&�*�+��[ڌ�2���"��tҀFr��F����z��`�aD��J3g��]}���H����٩5-��4c�O��5���-��s̩jM��Mn�9�[�u����ɜ.�n��c���mWo��l!$L�맗I7���J�Ud/�2&+&R�!󚿏v�7�jGW� ��ՋZ`@|]Y����Z�R�?��zJ�(HjL�UJ��H	8�qe����2ZZ��t��tu�U���ڜ��2�/;���n�\&6y�|xۓo�`/��ZK�I�<�~��������X��q.)C!����/��
������3Qp=M7���/�s��1�c@*��H�({�ͣ�N�J��ݲ�Q6&%�ɡ��0�hU���ff�s:��B�0v&��T��-<����0��$�JrG�'��/^�.��ݾ�s��A�ד&��l��\�F��K�((?�4Y��{�f��~�
�0�:H�\�}��:�8 e'��Z�d��F�����~ҵ�fi~B9�ԛc����@j$�Ϫ�t�� 0vV�k����S!$E/���.Z�HH{����=�U2-�mo5̒j6*B,�!s;�r��1��a�f�1(|�o۩�D���;��Z`��L��P	����Tl}ʺ:jʑ�);�軱X��p?,I��n^P�iDyWQ�&�+ſ<`& �����c,[+e������$��L[J�lͱ[�Ce��k�5E��烈����R���X��0`"�J��|Ȏ�T:�˛��ھ�+�t��L����H��!�a��oVխ�il~���jsQq��2PT�qԯ��*�� �R&j4-���&E8	�z@�t��Q���σ��W]/۲Ǎ,�YL-�dJs�
�p'�����9�2��ejF\ϭ�`���%ݱH,��p=����.
�5E�ʢ�7��{�V_���,x���ȫ�:J��׋dؤ���Qԭ-d�t�nC�w�6��������,�CB�IṍS���+��E:���κ����!����`���`��7&7��<���>\� '�A�����]���}D	�����s;�ɴ[�%�F;��/<��� ���#>`/���u 5K���&�S1���m�����RaH���e�Ji[뀺~%��4^�)�rC`J�A�w�����	�r��dj�[�e�	 ��h���N�����74�X�ݲ�`vZ���j�M_���.�z�j	dP�M�+�gR|�~j����k�1�v��A�VSb_c���]'d_lV7å\cm�9���xZ.�J�8Y�g\oO&����֜���_��v��0��]�Z]�ʘP��m���6��7m�䲎T_�1����g��iY$uJP�F�'���7�N��k�.}em�O\���y[�q?a����&�w���ep4Z�s�M�_�S�(����aױ�j^� &R�c����D.u3L�BL�qA@6;���M��@�8�on�<gao�� ��@��(XFcʆ�2a[�o���N�M
z���5�����*��0��d���f̪e���ln̵�9����ʝsC���ҝ̋8�����C!5Q�0ʭ�A�W01�8�j���F2���n9�<����3��
�pX��{�և� ��oPG5�N�R�����ʭ�� ,�M�!s�.J�m��a��0	����n��\�Ia��	NͯL�&=tvl @%ɿ�
���-��Yp<��"������/qs똺�|�l�؆������NȐ�CTq���7��4��w�=�7�g�Ϳ���Ɔ��J7�,i��{�1}z��[������t�����vczE_���V��K��hz�B�aME[eOf�Y7V�ס����x�w�T ����I���Ϟ��X�c���fv	��@t|~����bl�'�t�������e�=�i�>%�d�L��Ȇq$��#�U ��!�Q�JT�Q����1G@���K�����s��t�
J�g2��p7&ע����ڪ�8��N6�V!OW� �LN;yQ��-e���f.��FPr�OM#�`ޔ��u���T�(~f���א�{�҅顛�8©�,
�b"�����7Q�ָ������T����Q�>a��$�j�vU<G?�^@1��-!��l)��p�p�V����a�Ω̠P3�JՊ����l��,��+N�
�f�[�ư�L��~-��NT�dAa�k_�jC�1k�S��[� �