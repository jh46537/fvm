��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�	�O���|�Kv�_e�|g�w@?"����W�� Q�#������O^�_����h5]#�w��x��83�OG���ß�G��ȉ��'T]JQgL�Ms�8e�kç�t����铧�/���\��X�V���^���ʹ�r(�cz;`	��},A��Jw	.�Oe2�"Z0�:�Z�[3�����j��e+�J*吰*�R����F`�`�nCr޲�w��h<P�5C�%�4p�ɖ
���8����w"|J�'��(�^k��y_� 8�ܨS��wk�aغ���sX���$E�uٹ��y��[�W�Rw�P�զh�';��
�x<TC��F(�
ۚ�p�Q�jj"W�b�_u�O��S�a�AMNιZ�`��E��VޜI9�	�~�FG�¡�w��{�����١��g���kb��!\���u����;���vh	��<�;��vQ�k�Ӥ��ī�W���>Oy��|=[��qE�܄!B�C?R��9�A������
V���F��<3`6xuA��=T7���A�q8!{ĝ;���m���l����޹BαF���6Ϗyc�X��c"�p�S���Nv���M�-ibA��N]� A�����~n�X���uG^fz�TK��'���\��;�@]N3�SQ��ɞJ���Q�T�&J
�1n�QRV��*Bg�����\�*֪���T@�Xq�#��:���v��*E
���4�_��!���L=�o� "H����P���c"x���vh�>�DRtz3'"�P�e-?l��ZG�#˘N�S#�Ǯ8G�?��mC�Uō��]�"s�m\����h�1��@���9��J����֯3�m�vb�=�)��4`���
��M2�HF��|�-Ӑ N����0�����Q�N����Z^�!�G����Ng~�yU>��Z��ܰ��U�j�S �~z�)�ئ��P����H����&(!5s]��w9�䞟���E���FJ�k��9��'�C,>�`�Ȏ[�nrn=�Jp��@{�W2�Th�Uq�/Ji�D�]�p���u�Tv����F!�4f�a�2��1d�s���'�����ڏ;l���p�Z�:"�A3�_:�!3��Y[>V��l�-�`N�Tڱ��� ��މ�:�;�H���A��85<�E��T)}����\&xM�êu�^~v�lk}l5!>���;��>�N�'���Ʈ�p�R�:(wp�k���@�4N,��g���U���B���oje)-�yt1|�[��v�$�%"Z������(�q�q�omyP�R#�r�/D8utt����UGV}��@�����a������A7�)1�؍�iU�o'�r
1X����,jL@�=�g���Z�t�P7�E�+OM+�&�x�_�U�����6zp��ӊ]w�%�x�F<�MT�(MQW�x4�vML)�����$m�vga�P�04��댼$�ƽ�6���N{�.<�����
.F(�8��Űp�n�D�$ay��O�۝Ty5j$*���6ͳ\�P�5�7�5TZ�y��
mS��sV���13�z����K_�_ �Xq���`��޳�{��[͠��`cM�G��E��4�(������G����N9?�#h��V����!$R��c?�.��<�&��6��-o�l+(���D������u�q����k����ŐA[Ou+a��h0yq�K�wF ?Xj=��2�Y�RL(��N;W�����ot'�y��/���F�����oqT��%sU68��Ag��lY�΄/U��Ұ��ͼĴ�B��d5K�+'��.L�`"-^��'SK��B��v��X}_�4�����̋�UjC�r�Qu�}�3�,���l�Uhi:+_2�q.
�T�T���k�/��c�ka��⒮B!4T5$��GBYG�"A,Yl{(�)GG������G�)� �1;��(6������F�+��x)��L��:|6�s�A�nBI1_�C����l	�}-8=��~#��mC2��;�5�W�&��[u�0PA�x����\���~ �J��ї�^�Z��nf�6gB� |�az �|�>��L���/6<
����HaEq5̇���{~c�<hk�φ���#�^�U�e�a�4�]�v�'�����v��/���Ik](�C)����]W>��zr�S�|%-w��0��<]d��������	�-��&[�A��t�`���y��0�~��W�nR�y�8�7R�F�$+� :ps0%�`��6"V�Ïzf���G71���"��'>���V�]�4jq��Y���"?�|��!��0���K�gy��ov�:*6��,�<1.� �g��b���0�/y'@f�i�S����e؍�`2$m:�AW,U�Ԇ���ȞԦ�r{J�~��c�j��5�C��4�S~�	��By�}>�*"�� �*�t�P�x~�E��{�x)#s(�֌C�v[_�������;$;�>9�1;���an��{l��^VQ|�sS9C��n�v�~J6���_�����$ciT�d�MB�m$�^�@��B�J^gߜ�mkt��p{~k�d:�;���Y$��q��B����糫]G��j&�������n�|�ۥ�|�ʥ�o�h쇼�$F�y'/p����rZ�V{��Qk
UOp��K^ǯ�߅Z�bwVio�7����˰m�W�j���R�V�>RZe����!�U��5]zޫql�V0y�BhO�w8b�� x�r}�k��B�k4bu	Fc�+u�_XC������
똯td9�zq��P`���9q�r"�=��x�C�����U�eKQG���<�"rt|n������ۍV6�(n�/�
8���$f��}NX�h�����C\jY�kHY���\<�	��ഫ5��o2�.e�X��c�ܟ1�����v�\5L��HL�v��^"���b�;A�A���~X��̭ߊڭ�-��J�y>�nbb�=OwkL��8����:b�Ķ��v}B�;�Π�"�� ��G��M���Q)8�`tj�$�����u�+�+�\yX}����f�-[�0;c���I�"1�jc���DU8hk ��&~`
�K���8P��U�3H�ߖ��$�qF��+s�G�5�sɌR�B ��^�^��Urf�N�0����+��C"BF�ǆFgڀu,b��}�$���v��%�>��ʚ�-~�����R[y�T/�%
��Y��{,���Π�%7b$i� \t�@�_����AhL�dϫH=6uR"�2�Dd�c�+�}���d�E��2�d*�"y�E
���g��%�1�Y�|�����,�|\�'��G����ʵxR���vpg�¶����'O4j9�p��0��hh}r�3�9����6}"p�XN@�P�˞���pF2���i�zJR��vK��Ņ�Xw�z�2����g�bœ��M���	R��X>7
��Ӗ��w��~C��џ�.�ޜ���g���p�A�~x��8r+g���*_г�q�Q��d-6���Č��q��W�Θ�s�pje��ވ
@`>���,#�tZwC:0����|Ž ���7�^���s�� +ĨJq�GL��:�Y=�@�r��1�C��K��`1�u**�ML��_�B�f/�H	�N�a1%�g����A��H�8�l{8^����T��`8��a[H��D5Qd�^TJK[���*Ō2 ��D���wQ�OeU�c5��r2P��|�s�`�:}t���o	M����^z�6���|�N⹶������ݪ&GP�)ڜY:>�'��Us�������I�����&2� �"(@��_a�1j���E}VY7�+\�şm2�m��V#�T�G�A�Y�g<
|�0���P����dHk0Nw6�д����0���!$��>�}f��-e���*��?an8������Q�7�g�_�zVrӣ@є̠���������Aօя��� �r2T6B����X�����@rs�,�d�,��)lW�7&"Z�-��0+nL�T�`��EA"Q�:�I�a@^%c=u�˨Ҷ��T�A�3��W��
��wG�ɛ\�P���F��٫��t~��ߍ�h���?��{��1���_�,�l5��4P/$���Ȉ�Etn��h���A���
s;�8m�?N��m��ʏ&����Cn~L�D��c��z���ao*/�5Sx�zr{zk�c'Z����/��ғ/�|ƙ����9�V*���@����TIsׄ4_�m/���'4ĸ־h�m�i�t���h7Zl7��o�����{�o������Vd���t�!J�UVw��g@̱�!��n�Z!Հ#�`q�}�+>�hfz��V��.�l//�;��-�B�K��&�?���м�m����sg�n��&D��|�N�� /��	�T0:~��;a�X���Rol�7x]����@HӜ2��n��U�	.�Nv�O�ʛ��ӧ��0�������w���=��H�ݷ��j	x8�UL<�19OFJ3���i(��!�^U�6(]�;A_x�}{��%���y��Ze������p~�N^E��p�/y�}1�np}� f���GP��'BP�0�>�����Q�jӾ�3-��3�v�˒��6;��"��G�Wq�j���މ���8p!�:��Ic5y�T�����RM��C�
{�0wط��\��Q}y\|^��������;�qT���%Qw�.{�O�^��^Hi��K�6��o��m	��p
�?����S|�4�@�-Ę~��z�F��D�g!�TwJs� �������\�.��w.�Zv#a~E�Ʊ�k�����6��R�����]��B=�6y~���_6��L�t���<��J����_��`������Fo���
G���iO �W�Ơn�.mک�U�-�ə�G�<X�:gd%H���h���d��łf]��jؙ�/N�%��
�>�W-�Wz���d.�X[*�(%cª�D+�іyl���Б���:�������;��=�����uZ;�m����l�ӣ�K�8#<�W/��}Yd��O�y։?'s3K���ɴ�F]��vK����)�F1�6\-�b�T��L�
(�vEK�Cͱ�Z����T	��(E�m�G