// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:30 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ef0C4EqULxHpdvanOW3ipfABICxAOmpeP2VlcV5W/nsq+RgzGY15grIOaSFdehGW
TmYCQAfrQfppudndva5jdkbT+jOPzneLpzd/NJN8CzgNylQfeKOa9/Y5Tnphi8U2
WjJFHDnP7iXUqFmQatO89kdO09Uwz/esLtrP3/4Wzs0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16032)
OfIE9dvR4JcsbA61Lz+iXtFlPzZlqOb468crKXscnRAXCjacmcDlpPEGh8tUPJyC
WdCzI0tsRHFvQYlnMqaJQ0TQMIMpkFfAxZrx07WNco7cFYleZy9XYM1UtTqBpoEV
3TL/a9TL76E4A9EaOaI/8Ay3JxYyEMTfvapaED2VhPXwAtutOxojHd1ZobgLTyvo
FaLh2TxK+6WEARvzs5hnimkeJvAmSADTl8O3Rs4RPaT3uRXCDJrcWCb5UpeD2Kwa
IXTMizi0E8z+SdsBv8Dp8k1JyC4gR7SQCPEqwpHsP5FHP6AiZPIzo11VtULSn2cN
L14YCq9rl+EAZ4o6MJH50djFodVsPCjEKEpOhE4UymEb5WVd+kUpMG54cFsnqcTB
jkdSx1KVeJKRDki5mteXigKba/3osp4pI/5Z7NrOT0mRYlJdaXF781YWhApteAhP
xR5Ke121tLHuLXVK/LuBuJ2Sg5oQUJ0Lv7Ej6XuFAY9AE94twdBSkm7F25aJvvAh
ytcn/2+m8FRLCJYv2HrMCpC6hhhdqJZA7TxaWvGymUu8uJKR2n6w+ZNiAijMkgkl
0BUHizEpNeEDsjzqhVKFtUeExOyXRNG7FBnIcuQyhSQEDs6QUfUbkeaNsnykM6pQ
WudQgGXdAta8RA7rqo+OpI6cq9zgIb6uwikOk4O4ZDmcNLrBGhC4AkONMR11aOZq
pxRYtwwa+qylZb6spFIOvSIYrcny7AdXedAzgVnf/ER0U6mSjKbpTkMTlY22/al/
SCWyTIc2+/+6YrBm2TKS4GqKQY+juGlOvYqoWYd57pDy6raTKap5S7xjUw2/ukoA
BZSidI//mv8feC2ubjow8Bgb4nDQxGvj7bp2GGWPOrTVp7aCLUhJHv+t/MjkZ7vA
dpKawHPTJSzhZzzMkH6uxgwWaLmbIcqU355wqpTWsyrj9tL4UvMw4Gd+m2RWjqWt
9GUzjBZUmgaJG1Znr1H0engisLaITeX9HrQfqNyTGqnU+rBwoH/eBbnmgMeO0eY6
SMYaLtl5B9Gcej8adJM2z2bCP3Pvv3hQu7QjViK5+awCgO/X0V9PhBLwffmHjzdC
33amyXlV7bhQIqDyS9sP3WQ1XnF3LlUjWD/s9SMNf/AaQrL+m9pwJ44cxLtvyM4M
FbEKS7lpLhmpZNLZEhWXykBT6knyhP9REuNPxzpPQSfDOtv7RlEpcvVMq329vvAY
fCjwqml5aDXp+e/YY0HT02m4AMhSnAisWpiPPrxmG3NS4OW7bkCXy36dM4N6aQmG
lYnpK6BAjT5CiW4mYQPHeD9SnZpYQF0KvHCIGtTfi5QvRfhvk0ygM8oSS4NcMKSe
0WWiiC+vy/73Raji9nUlu00emLtNzkxp2r5hdCYd8lKlaxpt3wjBrvEJzC6rtomm
00yAx9kd1WgurlGb9I5o8lYYoHMoAwuG04oa4wz+om/Av9YvZ9VcK5SLZt36CuUJ
2xNfHvrPZ2e7l7B7DeyIWw9Ydjlvlvh4fT71LaqP0vD17Y0V0dXNoDi3J+uS90vn
D7AK6Y7HHsMcKTowxNh93mwrQXTYeS1KrPbQNcFfJ+eErooeOIoJcj6mmDFpHbxo
6AyNXlYUs1C0FFmVG7HqTr/pLlAH51R1YUJBfoy5ciNGYg+5F1SgeZ0JNsOaO9M4
76uvlRfYsyDVm+HugVjXgvwg78c0FTptYWt6tWFanotL0YLMK8MVICpL/U3OpoQe
ya0nypJcxfJ+lihn3VJujNKdmwvE5wU1PjYVTstSKDKDZcZNC80zqLR/qn83Kec1
JCtwbEfXo0ZvMdIjuIDh7oTjTIhlbV5+V2NYVTsc8xaDGhiU5sWyjQbKmV4yDx9u
NO6YO+Ot2lujrf+2aV0kilxkssq0HRssAe8auP6gfDkRQDkgw1PwniixNDfpsGBf
2VRcOm7iWJNKAqbqfCZdVbrmEanXCSmIyMIMB3PujQOYAo4Q98qmRX4IB8cX02Bh
GxwFp1zm/8jTqYXct2djVTMTwHhxvUjiZQkTU/S85UBZus2nWApswRtBaOJv+u/N
RtVGcFDXpIb/WrkuDvcxvbB5CianSi+q1AKyroNC2AHuVjH+Sv5XAHfnydGtKBme
eLCpfT1d3bb0tzXnyBVm+OnXREsiBvJpd0+Fo8uja+Vz9xAjAx3ke5i/WAPseBNz
uiPterrtskJKXIATE76r1pxEjGsRDLz9gtLx5abZdZLZF80kIPkbtSwM/JXrC5o4
rRY4fYvXkol0LULG1aqZEawMx6OxNxgg4Mai27/u5qTTESEuI+eIq/nRuWShSIZ3
RGuFsT5HQmYE2MBDgLfXl5AXUkP0+4QKg4LwJMfBrcz9Zr4ubHLyUCg3iLed6428
bQ8BLfbtCK4tcclod0YQfogibRllDPjWz4t4PHdXxPtxECwJTn5eois7HF/jgwA3
dfz538cAhRstBags8WCpZBc0qqOdHW865/7ory4Mz2HsiUIuZfk+UKH06mFrYQdF
M6ShoRoqGXjr6n0KqjTLW60RsZrTwttZvMCNP4qW4cgFTrwM3KhTPYbWMmfEG7Kc
Hi1MPhj/OGrpgC5Bn40o5x4/hs4DAvkTRHlOcdczoW0eiak9wsCWxQ+9hH7qKOlr
/qAwARhqk68mwTb0qJ20HYbPiMTlASPWsw29XF5HmwZdMBuiVY+2hrFpJpo7KV2v
6kK9+oo/zkTDfnc/v2Q2AKrSQ6H+AOdITDprHI0/u8kZwbouxayjnPOobltjusdk
g9DvcQn+GenP3FQjLJMEP2DWkVBGSi0mt0DLmGtL3bI+EF1OjLqDAcKf+ahj8r5m
AYNKd2CCrZD4QiOtS5KYB77d6LJiHFPBDAQlse9zKrjQj3L2lEJcb/zkKjBhz3hw
MGaT0LMiA6xn5zKot+ti/LlTuQAxVJITrbuSQAEeFk3OX8X7my9i7bCVfOzkBzCv
ZSb4xZ9PUr9KA39nlAk7GYHNx8bqmOX3JolXU0jBYz1KfqB3Kp2vY0YBFe1rYyVV
IU/81d2WMWBEBZgvaOgfnhuFqQWtgn9mapv36/C8Qql+V9mb1T1RortnIMOmvLoD
FMtiLbMZYVM/+h7AtQa8gqCxXq7vrNAvmg8tfzEe3hCxV4AXPnOHw8K6IxkInzz4
tv3JTPbWb/7+8E0GZAttRUv50ZFvgL63Qt00G2EXSx0opT3RXi6LSvtCaUK+AO58
K62tzGLzbvbaXXSDzTzUxUA2mgQYJIxB1UeLui0q2XnZtUNQzWCAm2QVm9oJaoPJ
DckWQVjhOAiuTw4YRdP24XGV+9Lbod7qZ9RLlpPcyeX9FP7NZkfEQz19+gUW7a6M
cqpc8RGirbIowJqhmy1sSy1pjEUAtQWPu4GssXw6aGKOF4Ecw63NrIwNgzG7YHkk
MntgW2qfA3a+k5nZHDq4ShjUMJF3apS/hIiWn/etFeLbETp1oGDWyHYPPqZdb+mG
PLkjohT8MjwjfE9s7Ut/qAaw7Mivikc6plo04twkx+GzmX0zT9kyTVdd+1ho/lNG
cgnIkatRpqREiGV2WDIKZc1LADYUu0yHVgjpfdZOmvrgrzEwOdXwubnCsQ/6AxfH
OiIhGHyTcWqL+MZIyDetwE/txA4Q1oRq1G77dL81V2KNf4oKo4AomxK6EM5dh6hg
QJwavCUUmKnZMtDOPGkWtSk8RjDAq0my/L2zhc36Z+AFWuUg1AwVs2JZVZK7AWH0
kxtBUFSCNlOQzqhwYuOUEXPb8GwOuSZqeyum6jjJrVG2JZ2bzLW9AJdP8DE5oa2r
XJkDIWrC9MgVnjm97Q6QAepdGPtzMFBuPwsSHQw+3Ht+5HybSPhr3cOTyN/pCT3P
ZTdxP0ndqhZCkG2Y0aa2i3LAwg+bHIOiHVTrF7zfk0C2fJ73Br7q4JLXTvSToZxC
asKlYl4Q62VnGEmDslAUkAHlpDDyZpf9R6eXUdn/9Yb+XPlbjzjThnMuxCg71jm4
v1LZijbBbIoBkOQUIkZCaz7gqdgVxIeIFj/N266q2cFDp2/Og6hoZ0kiHpQvBZw+
zAT8jfP72f0J/p4X9GV6DpToKj2BZHZXkHS00WmioQ1XcI8VSFOwxoXszyMAvK6x
AK9Dvx85lyvcZp4YMuwzvAAQM7OOj8Qrfd5/lxlbb0Uw6DP73iBrYjfELXbQ0747
EVsnNEi21Q36g/Sk3SpCnF/s5XNOuaEbSCOp2mOzgKpBESJmapjlF9c5+tPs1WF7
Ya7wPLC5YALuUsd0OiK8leDJ+8q/AOq6OlarvxWo+wQy1jfsYv4WF6UwCXG2rlZs
7tWhxf+utba7x2hI5Hp7QkTtehCf93Ic1OuvfflG2qKVIaYG/hO87aYEB2WlMK5i
3l6j0lJWrZ8radjQ4vkpRuEaB7gL3/yPCO3UGWhAD7n1R8PPfRBv7Wxi75utpKNq
rwGmHQaOFVDltkcXJVbLHE9gzfXyvODwaoDCq4lHjuPmkJfKMJxUK0vri3Mrg+io
JpEh/ZiEB8DE4XSwwK9LKFosdDowtw2tIUJHuJFKi92MYdgBuGrPDkEWenmRiCtd
xxlATotVTZLrAJ7ZVaheXg6F1lXFgVnyg+ymZsJ+DrfNsdfo7fu8v3Oolyf2PDmS
4QVGfDiI2tVrrqjqX95NI6MZMBiEIx3Cagq9K1X9VH+ePRJ3VSmU0pvLehN4FGhZ
F0A9G0DKHbfEW4WWU2R7Pmc0SGdH/VUzo7Y1VDAx6fEqzPrpJobVLXWzQCW6mR7j
5tOkKDyTvyTSs9X2/HTgmt4WA8bUSEFE8NBJh345SORYgr2ildKKSQiMssovWouY
7Q/PLpG/ZNcVKFQaalJioDDFOHH+zaiQ8DD/u1Dn20Zd8KPPQwscwHrdHpB/8TKu
5YZuXXEPo7KsCqeP0zDVzk04oWTYJfNmNPCkm5hbwoC0mYznlKO7XGuqeGAu/9XR
MmvF5BC8/GU5pbso2vNQxsxddDIGjqgyMh+73gqLKpn03eVPMdydjiv0Dq+x17Uc
Vckc3YJApm55pPSy9bM0GYc45zhYey7aU/LwKEdD7n2/9/JZdVe2xxoUT9LpSZj6
eO7ax7qQer0R6cQHgYeVVWD4Z+R8ZzQBrcR5ZrfE/yLhqU2ea5BRgs7YjT/ME8a6
30/Y7p7IdxLk68pjIozVtrGItWslxz2ybaN5O2+VCX9PnHrkQ8T95mIzdoCDH6+5
vo8sH/K9xsnOpmwQoj/m4n/j5VKsqp5ip34BIgUJIixJ6SEifgwjPtjF/j6un2iq
Voq6nF7tGL4XWLUtjtJBXz/SkH0wQFgFyHDUb0V1YDi9/Yo45MVALxiNm6n8rhP4
DEG9HQcW6unR6vwa8bWEcKtohnS107rbXCSsQo0e1z6ZXyhGAfhfvu+2d0iy5LCH
Uwm0AVbQwlYcZccwN8M71/6apwdrCyzacd6ZTr9zkhp/Gbs3vIeLVc3VpENJN658
6ie7WaUAM19HFIW9DoLmX7/cy1PnoDzfidPyCWJGbVjrUAp2itkTYAkZ2OhIzHBX
LuCEKrjzROw4NSqk3Qy64MOFcuAA+yQduB0sWnKuSqV2rNzkH2189cVpdcYwAWwZ
JhSjBaMs+TGA26Vv3pX0F3sy7LqUs5/+DHeoVJTFmDqLtdo5Ej5q1IJ3bS9rLMUZ
DAR+s+myuJn1blBEWc64dcv3intrI8ZC3SDhbFwyoR7SsvW8zMDPCy832+caNUvE
fdBPVfkEzsWjS8Nbc9RQk1eY4etHOlzKHVqWTNELxWx08Ed086tBHC2Ww1wCHaVX
QV2fS3UKKZNRfRC7sx0MI/J+cTAI1dkiJq4Mz5zS8I1JKxx5ZL6Tz8FBqfKCqQ2k
8ht6nZXUfW/Mj47hVlayg/KUNTPZqifKlRN/o1QiPBygaexatggHUbKFDYpUwle4
KY+JRsoOrnur7+w95taj52FpGO2i412QhgbuDFDRURgfMR8KXj41dLCl2WmYPmq9
ktjs64AnI+QZvjHLk3Vc46+C7/BdCbKqgSsuADeW4ON4NgFGJ40JYt/QiRnUtvBJ
jdWBSkKdj2vXnxCNuNUE1yvBkGIcOMnCrmlZfss3CZrRlBVLT95tPmMYoecyyfpl
EGQAqf+R64t1b9xpAdjYLlDJCx+yjZ20mnHiN5Plx/OL7jgQkqigSLg+Chl7eMlE
k9e0n+ytzg9lzjZ8pRfIgbDGJ4rKHfPe2bj34GFLGtKnJv6GavYswoNoFpmhC/V1
RLONjUi/WrHss5zJTR+q7yFbb9Nj0rqjJH8tLJdsZQ2chsnna72T11Ap5nzDeWTT
lYiy7wBmi8mmESIKPI1WVHCpI5FJU1wOhm1efuDf7mmigiylz3IhlVTGT8UzWgWS
nceuOwTPvlwSaS9WA15kO3dWWw8npodUhD/IXBIceKBrUh/Fx4HLVYX66tW2tQaA
SPy/1A+9AqmdRfCLRWMMaVpBVEsRVH18S6R3HcFWB7l20hpGjtYUu5X25rP3v/67
VMk873uYsE+bHLnGyHDeafKLV8LytN+/P/U//v9R8wsf4P6ZbWJr24+RJ0LscYVW
YUn/4tc1b2adfnPv1HjIeXsuYErIPCZE8+cPORQKoSI9nqQYzzGpetJsy0+jLSqg
VjwS2wug0Gq8pkTMBo3FWiWeFxxA5Ltgsz47x8sDae5jkHKW5t94CbuE1DLw0JO6
ZEw6a+yUIpM8arAV1uU7vs8rnytMw4AwBtIqz3F/TTV6S9a+SyLYIsFV4ZZ0lERq
K3HldPg0GKM+/UNfYGwvO0wwlp+KsJkNvevh6QmxqnZ4Sd/d1pVjLk7+zG3gyUIY
8FpvwoU429mrHKpkgQSZXjoUV8+LMGpv5L2OG6rogMK+zqhxcLJKxT85WrHkCFx8
MmYeUuXuNiZulAhm4loc0pWmHDqFBqXife2w0acPJsq6odQpMfI4vQm49g+rVi4P
gx6F8mYLce21zCPyqxuyOmtYg0fZpzW58e15q/vUf45/pjQTFPA8Z/xV5KfAfv7F
0ZSdNW3OdxDPLwTigrK4nGhUdQj/mTQlSr2aO4PB8tZ81hQumVAmMsq9dFpe4nzw
lZBv6bDvEy/QRnrMmbMlVp1LuJTBMaL/XYvSYJb26HyUyjPC41GRnY9bz+T8fr+8
sjukAUro0RNHqsjbiAMJ44tpBHsjt8Uc6LUasaqKEPhebajngjloDoxBbbC6E4lw
um8j+opgWxdP9Q7GJ6nQHV++LVOTeQzRwpLCDInFfMUxo/47vqhQ3FVvlxBCAxM1
Fajb+7f+11q9n3s/kmxHl4cqDlgEhE6Ktnw/HITElCuztscW+CkRmp/UUNCWrk+c
53lmxaRutVL6/0iRBsc1VFBSqzbybHssBHoJkEyYiEsWK1N9Ev+4AGitFyFVcg2o
ZQur8UazWCLsDZmsUR+cesNo3cjztCltBv5R2QDOmQtjAaCFDSr4bH3H0/cBvwgq
rzJQtLKEOA9UheAPoNAiyUlmcq72NXeWt22LbGbuacOo9mMJXP2zmDec1t9L55NZ
fLrlML+OqsNRsSoTDedHcJAUtegIwkxe+1p2eTFG2503yJ37ph5Ys501wSFRTpip
xn4J0k2txfwemAW1sIphiGIigKZVId9Yge3ulN4jsJzOoO080/Ah5IFtip05vXEY
fZ5ewOeMImlp763VSjRdOELuXhY6+vmwe7MHM441UDcIw6sD6DYiev31RHeDYLBi
s3X65FxwT5TczFXyX/ZZe5PB6VkH5jIfoo1FMMdDccOYmEvi6vRFNDbUS54e2Ucc
z44vappdPmPT4ez1bwIWLqD/itTiWxl2kRLQ4lRZ9MPrs6DsHraYr2qg0TuOUDZA
eW4QwzZ9vsJc36I+PnFS2rsvZY/3JtWlDX75fsAICNywEMA42vOY/Q675wsk2YqE
MQ6QhIh5/07hpoTHQgKGPFORC4WD2BP79PszTAu/sYdWjGjoNGmO+Qqr4oCXOQlA
cl4HCmxW6DyW9BtRKAfZ20haYQv9/r0vVpIWi2RbRZlV+pfxfo+ZxNYe7GZaoLi6
VOl0uPl9lXNau+2eIun0BjlxCxGoJVLuwOKZiqmYVUdCwXaYqroEDRf94jolSFJT
qc5DkVdVrtX+5u0R1nLN14JUlKjmitFcsSQNnynnecXDL4mvj7KFOg2t6p1/j7AX
zbUPi1Bj+DgDkmE3XzsxBSEPVJj+CXsu/dkAfKj1/8G/3rsSBcxG0XoXJ009bE5l
fWQecJZzyX0ZuRq7j9igTym1Vzsn9TcPGNRaXXBRCv2gves6fJtOIijmdyvjwhDq
Xx8rdALIs1Smgbu/3r2GXGULAt66vFXM7oj50SwYU7LZkk2UJ30sn6OZcaSeuyQ3
gL3qyWGTj1JxmctoIcrbgyh/rGpuQSaI8Ege9aR5rjr3FooIbUIS+K66oR4CXpVm
v5/H46CN41gl8Raa/tz3vctv67BVss5dMQjlSRgoUlXbTTtOhOvcEK3L6N112S4D
fkgMP2O4EZHuhchV2mFNdM2S9t9gXEDjVdK8rJAksoIvIWAC9Y6NaSyAw+Lyt5dU
vq+de6V15PG6qHQMkkNsrr0YCzJHm3OI5NCGqUjQwgcp/wbYmpDugjbtLQpe2VTq
JkyM0OW2x2iYtlsuc+9AW//1Q8rJ95/e3dTtldRQlv/6THWLe9Z9/BAWpKK0YTdy
O1zEgwTucTsJTfKlib4H501iaAPC6uzkk+VxJFZeICanJsYLP7B/vSa5QmpoA81c
ySqHFMjQj06oaOwYGX+GCw604rKsIHcCYpfYWL+b78Xe9Gm6czEBxBPINbonXWn8
azW9h6xVakFE2T9KPYCbPSlxBwmzJfMMl2MiidY9x1B4h/+69kJCMMzEq8hHe849
xYwsp64hAPXk8P9ZOrD043peHcW4M7QXp+bSdvBwenHSbNy0RTyKHmUa81UqUEHV
fGj5btZ3zRd48T4tCMuI37OUOV0hDe8ClaSTPT06LZVlvo3AsQ72NOKCxWetzpjo
NnPWqn+jpTFnyO8r+wOr3UU7lnLw1wxfiv7fA4KhWfg2uqgvR1Qpwy0KGX2Cfdyy
4ZAKq6eZVDmF8gvlfDTop/vJSw86/UAGdQmOs9Rr5FlEOzspbjvtE16p96d5SipJ
Hzsb+g1w7acnZBEzvkuTy2nMOiC9EDr4e9+3dTm5TMhGSubYHFFVFw5Xwzt5eiCr
W2//HVE1Fuyy7QYdLOxCt3AtINkwWyRaa+BjmA/sf9BoYhM8AxhCMVCFlUqmGykI
fkIbA6ciXB/V39RXjS99jv/KHGDNTMDvuEcYWjxMl+IJma6DBQ6TA/2kREwHbEBm
MBLmlnQYG1VjT6RLXuBgKRwxQZCXqbzDfo4qlG9O+NeU7lb2Gf/vh1I2YMdVN1Z8
+DavX+NWadEnruvtt9Y+dhdN/Y5TKCU3/JpHSvikv+Uwq48EK6+z8xQLy4MPz6gO
pTFxn3aHJSCF04XG/Bh05DDI9bb3lTXbduT9ETud4O40QGSrb+aMitFRJavUhbsk
f81uoLeGuiNV0Znw58sZOKweheVdqyn4BLamGty1iEjmXhFTCxfFMaEcM3h0qrkz
yRYOUpIVIs8i/U4jFzCWvAeF8CYkX58Nrufh5pNRHzQlcvK4buShm0uX1x/MIom9
GuRpA+eok553ZCb3SSMHoHQ6Az23DZ2dfQTO45aV/RZER16IPFIxQpLikUcn+QGh
mePh7Se0ESyQo6i9Ltppk6E9CmFsvyHoKR0Udq1GlrCw9AvF2nOBSlLOdh/Z7OKF
F6UU6NDoNGD2E4vd56VOye5P9O5oc3qzVLoyNU7Rc9jKDIfRFprQbFN67eC5+cN9
fdFFo6e44omlhXvXeQtETPWj8Oa3VTdk/zZZkYNxaBiaDnAFy24J8T3pjio3XbUH
At5W0fIOApLnTdDnMf+WoInP/RV4s8UTaMz0/jlcdo5WZD/8IzQ9DAP/lie8NKM2
2wrKfTEc0biccHC4KUoihd8tnzMwJAH3qLFUeqrE9OJTJ0MaNqOU78FjgDTnlDfU
iLvTY6/J2EuvCEr9pSy0XW/xFBJhPN8dEJ9szDX2gCH4r+uINLHybdRQad1ByMLX
nFwZFkA5eaB6Ofjajw6oTQfIudBJV/feLBVcqXx0XX8kGMH9JVQtg4O98ZS/t+uk
Uus3mBNob7KkHmUW5pZQnxbS6lwr3K3skLJAQz79ZcNXiOSDRD8M0N6Xl+Qiloh4
3wyp3zn52RujI4WCCuw9CxIV8pcClCXQ9k9h8idCEHh7Z7d5L4t8E5T8Yq2wxsCL
VxLQIrmQTeblsM5DGg+/bZpBzFEsGlxxgQdWO8v+ve1YeuUcMhkpS7DHev+p5dqe
NChQOGS+4UB9G2I7jNsuyndu3OQD0BAJo9nNro+XAuiqXqr4fn1LoUn2fIoAdhMB
Ps+sR+07WjH7BRvkq/xAPMFbJYzGNyLOKTMuEOwotx/dDIjMp0/EiHrxmpp8LdJr
TDI1UnTS++kyZv8TBNTwjmJ+WNYspXLZdFbrBLJUM7konoB6MWAv5luzzU3HuTXW
wXszvEtrsJAGXOBXc8CNtRz98yabeELLmh2rbjLQ9rKmqJXDX+PvHsMO7WkTmb9W
3BAHJ+hGnme7gYfonyMOCbd0fbFLkvuY11epJrIzDYxH6AobaolhcdYwj2e0yTEf
zaH3/N40miU6Rtoj1W4yRlpVNDD8l5ZNL0pOMeoIaaGydUmgwxy6UbQc1y3UL3GG
9HdRvuYZV+X0uiXMcWj9/sidGkewapF5GsO5pFbw8RJPT4TJkH2A57/DXrd5fIco
gyG6YzpOxwctvt8q3rcVvKh++nWwBZ+wlQEspjLmTjC+r/XaEnbRUWRfQiOO9Ufn
sBkBbzjqkKdQJymxr2aaLJ4gWWTlJ8Nho1bTt1dEVCZ0le+kGsMsxrj01l0pf21k
VKXr5IAeznCdA+KMdWt0ETcqrp7R5tFNV4eDpwW0DMgG8DqEebPenSQzZXiZh6wh
JHpmrO1JbS4/1CT/GWvRVdhP7DuFoxERWAgfsPWwf+Kos1I+Vi5IocqWmlBcVOiL
eYaRLqSZ2kQvvrPM3u2eSd0BWwmwc1R1elDz1phPfELNP2cFCwXEeYvvM43MIIwC
UEeZsc4F5X0EAedid5zJHSC4nZtnbWdRDZUMI0u+PABgtDD2ywLTpohzRi9Rs70C
+Zf8YIFkbi2Wsb+Gzc8GT/Gv0XXebcq8F/1vpIhYWX7V5wAs9bqx0d58VVMtJnJ0
bWXS3EDkyY0ecFyWzZo1bVt1V9OxCxjMKoWv0mjWc2uN3AUIpDKZfGSabV9Zmyjo
RNbqm/DUPQNtorjFSAV1f1z50ztNuZGkDv5yregJ0Ei7CC6xbPbEkcPUHcqe1ZQn
RKp49PqJNtSE0MLi11BtHeWX5un9WraAmItn1JGkAd1V8ibfHoijRGYlVHqVQLHW
gkP5x09+IptEvq9XnYzXVZ3EY7zZeHgvEJ9bHw5Q/Su6/P0l71NOAJp3ypBYWxKj
iICG3D7w39l1rVbYaLWoHmi4RkPaBqVmQXRAKWSOMt+VE1z30Nsunb9R5ELXhIO0
k5arjXfDFjNlyuAxlz6H6c3RvsrAI/10usGI+Udf7xyS59xnheVgl5vuzE40RWmX
oFA7dlrGFsLYzmGy9WPIGwB5TEAx+1mgfWXeVCvDAmUYxGhGY4FFUszaeIQSM8LG
QeY73tHTH1LfYSNMCGRIStzUwy5k9quOYiMBHAZb/z5H6Vy0NtyDCaweRKEi9b4q
rNu2PqYDOimAywL1W+0VJ6swK5V8JmdtuCK9ZXu3JrCg9wmgOGF6eidgtjBVMyWm
qHzx1lKtlg/Z7ouT8GjAApWWfCmMn0x0g/pRsbeftxQdT5tSLgIxxGUqacC1AdPz
GCG7tVOmNWHb6Gr1gFiWfw4Lv/gd8x0kWKf1Y/ZQHkBCF+YsMV3LibfS7NkZv3q3
WWSB2bbr1u1s6CsddfbiHDnuFwv83sq0RuEYR3/YrT2GAwFLD9chHWkmlHnUjFmf
yNkOwgMIBzpxhCEvQfRLHZDWF2VywZfSviz3DyhpESxQMqW+91Wdnca21E3sQXcH
C3BFjqHagpaKpaLKSAUw6pku395R05Uih6HOSOAApqEyeYVv5Z1p2g9SOab1wDLX
swUWW6CnDLA2lvALIP5rxOT6cfBfcymyrJUV1dPV7ac+FtJ2flTp2SWLWCx28HT0
oxe4sxCTZ/aXnXJ29+jHUd+bBTnseJE/tli1Q0H5/1sW6f7t5Bm35LpQRRBkqxuV
Cz10WWKBzPuhlt0xSAOmJuZxTK3t/4F93CgLUjGTo/MnVr2hv4zMkeapwjgaXIKr
hN91wSa/KxbWkQRPfJqm+XPweCrqYoygpLeViZu+VyTp2gfebcjtb7iNXonlWYpD
J3e73+lgL6XzJ51oa7NPK3Au5IeWaYNPL8hUpKVYXTvVPe5q6fJbjQUA1J2j9Qoo
X/xa0vGC0Na01/OyckWtPX/G1v0p5kypra8GobzYrDVysf7XdK0I551Yi86S2JDp
uLt2DH52GwuICpOFy+1qOe2etQGBA0iStvadfWFi/batO63TaZUftKc9kslG9OSy
nHLYXekqN8DnBrnBeu4CyXRGWgecHTRqlHguUIoSY1mwSnFQg/qN8EAm99Lq/OTl
bNECjgOqj+Q6D/h5+dCg3p/mmT9YXuZx6QAejdbU3tLCKsT/4xJZzLi3i3x7UnmP
801gk23tUAEae6hW+fHUJEJ1ehqRYcGD8xXxdbfGxDVRwwTuNc6pl/7lMnBfrv26
NH9xKozTBLk487kgHJUHuUVJyiLJOrKNVGnDoWobUOW//iADRJNG/NuB//JKhoDa
8oSk4aCW0r8HtNeH1FUoZTA2p0sb0VP5zl1pXF2U3eFpqHxewXOjcNakMoYAhQyP
WsqHozFPJbCHh2AHfuHG24kWFZNmhW5GJkJ5m0cbkzlXQA+XyR8Zye5Wmsw04DBA
fJ03pzcsxFRZgCVhR0Ly0EhYsQObK9RpnWf4Ob3dxwPf/6tucerpkK9G3xqBZ9tC
JFkbi08vcBjUQE7nZNJyOUeqp0u2Y0cHH8AfozTIKQkpTFjOvoFrfYYkDdASxRm2
QPlxQB5pYpdwQ4fzCfDopaRnQGashLMBYi1b2/DJAjsmm6woLrBYpQmYusQNLzOz
S5xMw1zf3weSMDMM0KBLcGsncOZsEw822R1SKHKISz8Aav7Y/J8UOGzdaTmQIpZs
yghvi/ej2hYvPVPv+4Du1f778Ae5ZN6bN3VvAHWGhpaCkacCXxHuB+crxzwPUnD7
dmxabms9L09PWwO0ghLZhgrK5yZLb46vGJ7Nrux9BsUPNbxjoXCo7itl/MrA9FNY
bWa6Ao+y8XdYTQhMQtOfYRdlq4Lg/nW30s+Rybmd9r2qP1RhgHtrbdY+l9zE6TPw
fbUEikunbt6fkUJgzDNf7irLZ/gDKBIuU25d0lOY5NbKEdBkdfOaucqMSGAEiYeO
tn3f0mkIuufNjyIGByeY+PzLQumXzvsephSTbMFiEfdTDnkU4/7tppZAnmyg04eG
NcrPSMr5MJgiBrUlRe4NaphXWsJ7onR/qRxrLBGs1PZqMHqBFEqnd2z891ykRQj4
779Pv5e6QlqrO0zW4fk3VtaZp2KCI+S6H1FfZwQyCitzZvYvmGEbktNIoJ+LL4h+
4kTclIg+MwU9LaRNUz7BmHs3054YDrzPkv78PVa0OnOPbYkX23pzfSH5bJNilREL
9DF9GXkf5H0mUP4ab5xC76zPy+rK+GLwLbXH6uzCkcalKn+71TkWa+aZ9FEOwTB/
StNuylaYLqMiMHw9KIrPw6xbEjbmqWXataJbvoeQXZpbRjnMQu2YaHViEE16ErlV
5VLVmrCs0q08vR8960IR+HlBBfvV/pgJmHEkLkx5YGyHf8kdhz+7kCJWmZYoo5KC
LSQFronZoww+kMXhMHi44CbcTZgbFE59Mo2mH8HYhzqOD7yvKPNCmwmk8WQf2U3g
oCuF1qiF8CD+rJwwDiUotxAywSNf1zhB8CIhw1LbA3U/PGxCvCT3R6ClMYW08m5d
8KIQ5PBIavBgH7N9PshyBSCbvtB85gumMg6w5GKUP+M7d6u39cuUjTCR2ORxVFfu
UcQGiyvsuT+RtucxbvwWZBxqNYcJTQc/UFNwbtnoE9FmyyKWlXtq+DQu3Y5tI8g1
31TSzqz5tYFIP+MChsFM5PSTpM0cMoujLqEqmGcww4ixvVyu52kdPDNI4VePcuUf
Gv0eeu0VphYD3fkG3J5hzP4DVRss+GPIxusBGoQT+4osY+DRpVe/vqAdTEVyyTmx
RDE3W4pIpXLQe9D1x40A8HBMcrIOm8jHS3GHBB0GIodG6eABalXBB1JL1Ab7EHH4
tIbHg6o1d/RfMKW/X9T5jm5n56YxDMrAvIsL+mB19ZpPKsv9xTyCS29C9akZldZS
h8UWteVa/D4gXEzZl2/mB271mmyaMunRc9z9L4BoNHlKowI8I6Q7W1+9dP8uMmHS
lTX64x+VF8vkrwjg1vxFAv/er27Ph9Wk1AWhpX7izQahJInFzhNc9UdNywOBkS8W
37P/lvBrIBZrkF6ir0qKLqeGURvw24ad5NdhiOlgUHJPHSl9Wj4OPEYubDsJbppe
tIqVZP/uJDXPcsmcjPR0HW38t7GH2CUSDaegXsvIYK8VoqCGJaNjs/2NdngOgLgs
gzeXiLxRQfVbEC1yLZpDOaLMRQkA+pgWUeQeM67VAFIMy/apdQOSuPoclv0royhr
w9hxgTJjnrLAZ81+i2rKD6slyHAuirVCx3nAegJZ1zeCQKUZ3gGPJc4r8SIKYRZx
kkfPRo2sBJKCwLV20MO3maiJH+FN9S+AieYTCH+2MeP1KGJNQDnY5fEDFgv7nsNd
TF7Yu/f52b7vZSw+ThJaouHAJbyIBR1jPoTa4xecka35JRh3v6CRv5OyCKWczNhx
/wxyZkcBnd0sQqJaJGHpIt0XBLIms/al5MKAuZuTzowsE1vhFHxSqLw2qXSH0CQs
vYF7mI4ekkHJV0QRvqzp5wsH3cWy/6ckthsk29llpWXleImsVKRfsTqiSNVBntfh
00g8PitiYq3YKPlnh1D6DFEbYoTvmOqNqX4NGYv9UusjJ6bxf++DP524WWB2uBqV
Scvkfj2qqHkW+7H287tphCQjmKZjH0fPoHYZx7aH3RWpTzslh9WT/9X2UIxeVNiK
NESIe+PwEajLuihh1T+08fPSAdZaWpRBIQxEHE0vbYq2TZ7H8rXYSfFjIP45g8Hi
8LfvERMIXzcU9TDePOy+ev/W7TAnhWvpwIQcoo20SdshUf0mgxKmL6pgfLyBxPFj
137dI6wqByvVP+N/1cK4J9Zjp1dScMZQYceqTn+scalxhgg92rVYf63tv4sUuUNW
n3xv/c7bkycDBTMLMaC3Ew12xJqeRWDdBSKcsg5s5W+gULyxxhlUVYaDrgSrUAaD
6DkGn/yNTF4MChexH6oPhFWm3Z5XrWAKOD1UfmAquWr1NUX+mxeeI5tpDgnLuYEW
bJZMvbRxpoPPIM1ytFZBBgaVItYQAdtZCSJpGW2IczFNS0rHuqYxxe3gwd+E/eSI
EbyzKBiFPqI+k4HC/ySpZpbR8kPkHUnFyASPVq+scEUmpNx9WVfQlFDouxalhMdJ
I097d99E0VKv1gvfMvYIR431A98jBc4XCEaBZSs3IuxER3FIi5wzJXdiVIUc2Zh7
Nln6P9JJfRk3aIje4MjjCefGlFLpb0TtfSAiXdcLhlwsvwOfB0QLnJqLAu+WN1N4
qyJdXtACfdl03cBntYp5LzfS4fz2iY3NdvvZR7hE0WtTS8o1r5k0PuOWim7/zu3V
uX/N34gx1e2oo2+LKmKEPLofTz6BD4KLMAnUIHSbkykOujn//BN5USRDMjSlKvQH
8vJ+wAA45mgvm4kjNG+kxCuculGa+lx5bO3w5Qe6zo7yCjoOxuNv4WTzydHmoDdm
CHY/NqmeKiyNWayfy2B6hz0gUF/vlDEVoxnBgOwUMXV/Ph8gmMiX1CPiE4hVlsTZ
8sDfinHgoUP5rE6t1kmQgmeM1YPEwMSypZBMsu+9uPA6/2nf64T/xsGgwyDVfaJx
ey21V/yAeWiM23Bxv5/aTCy6ELZvOBaMKSz4zHOF7v5fQuzd+pxRs5fTub/4X9q0
ieRD5OZf+hDTFi72yphB3zIh4g9x+HmeQFaW6g3x+BQhwKStGLFl/kr6sV4eeAvk
5z25sr7bP+IECSZHfAYRgIpAtZksFB4oXc4qdT2gEtqkDO3owEa2Xn7cztJks1gg
U3XYd9zAB1i2rmB3vRrqIWLQmlBbb+gw5e/mIl9YUz7mX0iQM63ss+6K5vzWlYym
NgpsrP1Oe8+GYmoDhPLTY/2f4+YccjUHok2lw29d3s09CsUOdurbjT+YjcgnSmHA
vUzCFtsuNYIiVTJ126chyoG8lHbf6lPqSeYQOfJpbFkBk/vO64K7qSr1FbhDpYAW
j+wCOmxRhXQvKptD6Ia4Z+aySc4jVLdu5MDDurBdN+VVmbW0FuRh4A0WB30TySk+
x1XSF1PQbOQSNeB23TWtjNpzsiVESyYuhyJ+T6jDe4NiMLb9wiTXvTUajsRCCoax
XqW9THJ8GjvwOMQ0DxFjsp0woGC3+ptSEUenGdXXL7Y4R+VG8LVtq2zg9ln++8c4
mDcjKcGngPIvCuasoNqSDN5RlSANivx6OYfZG68sEOQnuxFdYi6bYoX9ljlIOZxl
jDPntcsA0WPHk6aQlzdiMjFqhtkhs+QiY9Dphmqzn4zDrQexkmZIAXZivsg6KL3Y
1FEpysJ6v3UTy/cnrkJz1Z8DNExLTY3x0AlCHmXMduxl5a6lmWEtdxWYHalbN5tz
RMLh4vevku9MwR7d2PopgTgSwPspwWIiQNJtB1XUuY8/NAD9eGeUVwtmKxk4bcMc
fSPBZQeiTSrd0Yh8ksGMk5AGvGUaySPkgY79A1KBnnjRjB9BXqbiPXHt23NkLJOc
NZ2XlEjJheGsJzhDu0Vli4PQwNyS/lmN9pikp0WtSSDynN0SjiR8J4ZPCOaMKAex
GU4aTbhOr35iW5UO6281a7IsY79+6OG8TWekq+cANp8UJhIZz3gHOEdl+NEhQhSJ
Jx0nVG4gnSbJx77PwjSCtXwz0DFAucbonMJ1GYq/kvFPuHw1AWnM10dOjDcTiKcb
s84UMAzmAwkasFGvYQlCX2RTm2tps6gQrDkRgwogMj+mrKgWqVS21xM9LY2+t7ur
kClJgq+bmXMQVrR+5zliXBiZyeYAhmdSNjt9vrH0QynxCuEj+/kOimAY39zxNYZf
W2/1qnCx1CDrSqVXaR3TyOImuEsBm8qjxqaaXvCrqLEnkZXJlSbW995hBzjc9lob
ZnggtbYbbTvvUJwJMNlJ4ZvxQ0jjiHIeexgMtqxaAJMG5FtvSHNz4uconlpIhYaM
pO+Dfcd3ZCHa9fCKtpOg9X1g9+mfBtS3+VxhXG2MQ0HQBs2e4j6afhIzR7vvITT8
emIGoDI0yqhKL4iM07wcK11kHawK6IFatCUQVUAH7LgLAehjWttj4/sT8ppejZSZ
N0t9jGgM1+HktdCBuy2Cj2oBJFC5bCujTaJWNTcVd86RQgRojqxUTHYBaU3qHE5M
/j3cf6j555A4WOWFgMhX81z2ClL9qNs1dPTXl1IoyDOxVtQ8AxGO43dqdt95qeMk
LLyiuCPpziXMa0KTou0LDGfTST2Fetg2knu6v96rfTEcv4SgXesPYkkAVEBCcWAn
nF1md2g+WI55/D57yVgvHDTh+mvaxGX/1EHpcTurVntAQOdDWOX8xqfTRDj+OogN
pn3vWd+HoCKhnuJ04T7ZOZdpyrwhLkYzdrVfco1vzXbvOvXNfj+88Bea5z7TpHs0
yDCVD8lcppaq4ci/r2hpVtPiBtic1e6ZYtu35Je+FuHaW8Fq994StizzXj8K7uAu
Jlmn9qDCLkKDI6E9DEeIbnG2YkU0uvTy3j6VlsmgD1n8RY9nZHJNBw+6XhzmHxpY
j9WG0Pw6c+huH88jWkOZfUmP06N7IVOeXLqxcU0CbZmIqLkuKmymcTKnOngFfZXQ
qP81eSOg7ToKJY3U8i3TWXZJdjzdwr5Cp+2jX/lUc1+B7vNwMtGInEi/Lar4oxN8
0buO4uDZLQ+olFSSCCJfjJ12BN/5Yzdi4LnLquMOHsDzDhS8BNTIuT8iBDQUYEEY
oL4nCxIY/8mZuDCv7L1hxQ/dDcJLFoSN3teOsUA0mzkbxLAGgCZFejkvEw1S75Wn
WGeiz8q0ZttIocUcWEvMLfiXFxhhyiGYxMVEzq2E8sN/QWkM3wPF4iQMrSSWjVSc
VG1ogzDeFzNWWCN0NzvUtpcC+po9GhWh6txK8yhIF9jRYog7k0I8FHrv3h2YVEVT
KuVj3ZzXSTNT4QCJlzp+Eze4XvxawCYXTjG8Po2ARxvjRLR0Nptl6f6A4dfv4D49
H6iMxJCXdxgBCHp+qAAa2pXcwqiDHmfHKlF0gN+g2QPOJD1zOxcvHeRpXk2ckSD3
WjYx01Ktla+XclFiLNbW/hxrBC4ruKZ2Q5p9DjV2XmLsiKB0Zi48J1ooPtV20F6i
XiIXv2ooXQnDg/Li7bVb0mi6v8IdA3o+hED+8oY2xeCvzT0RCjlSi7xxQiZZIX8Y
56yhYDYbWJexrWmZx3hief94yvr+HCNxJlx655uMp7w5qdJeom9tpvbbkd+d/Ih/
oKnYPfaPTDEto1NNfBUbaEre72T2LqEc+uQHHPaXcLdEybtu7cFaaLs57ar6N/FS
ps3QH2WWgiR+MPAbNJ8bXUG5UvxGc+omYs55+CgqCxzIO9eYRhhWnJyCmIWGL0dK
v9s1/2ubNcAyIaNJzjHvf1ydxORIhKzWZbFKsyZLYN2CGdYH6f4NK8Q4lpBWVkDd
NXmR8W0MVEdyMB/ehDXbcrHIYjIgFTyBEOqEcNeqFVhvnRExjAwJ01Cz1EUCTwxs
lw9P1NObtjVi1sgF+czkJrh1iBxnjlkKi3xyFMH+gwBRe8Ce7k10/xxgAjf70qQk
o4cLbaLcNH5ZmCCsZX0qIAvs2hrqDiXdNOpyXYPtURKrSH5XpEeXFxWXCwm7JwBt
I05UcRyWOThLk3JFyre9BNn5pg5Dzl9A5+m/k0qkQekn4MQuE1hm9PXSPp2FRSbZ
QdKF2pe0kQVeK3Fh1NAbKChZIKwDbfnzdcNtJ4OWTG827aFHdts6RMoicn5u79FS
kblzMkDFcAsLz2AStS/MWVs5klOuNYxw3cYzEVe8lIMalIwLe6IffUpeMM+64Rjc
4w6dQOAOtLK/W5MYBb9keSikM+dt4p4+AbCO+mXudFHLOh0MQj8Ob2HF992ZYr5F
Chq8n3gczDY5hpWkW0IyuH6LlC8nEKfinvW1YNvmuiREZgbDI5dxq6F9PdmDUKPP
ZNUewMZTa2t2GnPEUcHj2SzHW89nGNkggR+bfO25o6H2pfCSCyiA7TdgdALDkvqz
kFSRWdTTIGDtl3pQ6xBjtnc/UykrgvqKUszjM6BxITUH2isGO0ipLZUZ4qYr4z7C
+1bSpUOYR6wwD7VWR0c/Rcg+lXmsFO7GmzDUMxARG5mZ1E2mu4qbeEl4yk7gwdDi
TMGej+DsHiQnhQm435cMNNV5fzFqxKrxlvmQ6b11LTgVUVYmgjobrSUWhk6sGLQE
DiVpy8mDJ/Qhb6m7Bm9Mk3BdnqskHAxQirmVzpRzHeQikuzumxLupFs0etp92P+H
IkvcjbTz4aR16IijdzC4gzRccfZ855EoeDvV5WXPIYk89FBVVGwWYlXAAxf136PR
WfN8R4gMgSZpNVfYPfphMGKxXaeiwyX5m8N2KGHyfBYznnYw0ZHGzS+xUj6nlhJ8
qM77NgREyf62sRl/QDoOfCPbFhQwfrpnzX3HPlMIYGP6mAx05JaRNBSy1O0hV3QN
j6xy3vLj+Vfpz0zHZvhgcUq6c2cSeMmvaaoF1HA0S2nueS4qXdu00HIeo5I1akH8
Ep+yB/V1ZwLM0QQ/ujak6IbE8+NHl1o89+Op9PikIeB5D9jELs2pxh9siTeMsWwB
DbBhlyeN62F6X1uMtZ7to7oeZXjAPRj2SKZsfLCdbqEKaEbIbOU8aayA2xx7bJNL
A1qGm07JlnTx9b3f0/nmMmvq0FLvEd22eIqz1v8njhnLKPoHwop7K4jNik680DDN
7d9vbCM+qfpvVhfT/XB48Ut/TlNWO/Jj1W9neHti0B0spOOr33NH0mycFx+kTd1u
1mrIMWBrBnAL3lO1BiVaCWtI19hX/shIRvcbb4g2aE4bPvrQDek+k9IqBboKK09C
dl1wtgo/SCN73Eof49/0RegmvLSQSW1whrgebWnV9UWTVInpaa68O0ru75w1dxZK
eY7Of7nBSsXD4QrrX2NwHInllvylzpObTdgZfIwU7GLvojtYbRjcQ9Wl/H2EFtLg
HkcJxPBUWRS8j9I9xUnn9t+mQxwD+XUiwOFsDeeoWRmkDrNK+DEhsgfp2sEYeX0P
qj3xHrkmfNqmJnxIJzKDPtf7jYVJaUai8ujLqJJeShr9X/QeJX8BmDvqzQdy7eeg
DXyjbwyr+cO64Jb9mBsCpLb/qCRDAZ3kAcy313Optm2I2T7hZNeDOBQToiIonQdP
Qp1oscULV3d/94sGDthKN5/DtKieofb4kc7Nh5rGhFCO35vK2uuE5qcaWhSOOHyr
dv4GpSPDjy4N51eiDW446aAyQiwpCRmXmDGrr+OWNrYJlTB9lEd/zria0Qg9vANd
5k3FVuWUFM0du0SyKBH/HhVSESpRBABItsf/bN/3JSjxsgWOuD3tq7eYRFvW3Akm
U84ekwABMyZqJT1v0VLdpDUoIqkv6QFjM8r2kOKobTUc+Vh7sTUVAf1c5bml6n14
5IwOST9yMBULGwb0GSnSMtvLlS4gpQhmCiajZsmlP2If7s6msV8Kl/C09tTovj3j
vG8/StsYquX7efhCRk0KmUngogjJ2c5cX+0HxS2QypQ2Jof2DvQYYMAxHVXMyslV
Eha8ro1bXhIKbClz5O9XFUdy0COJrRSk/n+j7YgYwS2Pcl4Ri3MEjYoy7dYs/EoI
h4zDMVdnye7ftw14jpipqqkdXB15pJ3r3h9PzDL0zia3HHELBUhZr+cwiMvK4XTa
5pUmQ42UFS49jEiTWEWY8MoDqDL+3+N0y2/JNDPJPHXSc+VqnwgbO8IzMlxkMABe
Kevd+FDZEPXd5lAEZnKeaPz/eDcXTIZ9MmqAdbXxsq8l3hmE/5lfDj3/cn6AysXi
2bwheJfEuh43uiPLRJgk5UFERWUzBFc3EudFuCP9uPrkkNuT3ep/XnZgu16U8ADn
x4wbqeir4d/aXCiEjzHTS0U1bDi780dzla8aPtVv5j1PJXrP2rZvNk23bbFvQj9l
`pragma protect end_protected
