��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�;O;�n��E�Ę�O���q��~�F�n���\��"5p�h��7�����k⠂�֎.R2��
?�^�1���r�����M�۾���ҦbR;A��X�5�A�i����Q��.���g����e�u��w�v�v��õY9 �Sڭ���H����$zw��0_��0/�Ψ��J�XC+���y��yܓ�,x�������b�!�&~n:��d����U�k#��E����@��%��[z��a�v��2�}hL�q�D��I�<i��ͽ�6��tZ�K��|��M���߽��}>=�Ј���P<w�t��x9EŽ��v�h��_T��̽�xx'�}�蓹�I�17(�2����Bk?��{�v�G�o��ꔲ�E��oQ��Go|�u�$�6���E�������U���]nam����d��U03�ܭ�+a�'-ϝ<�( ���KL�'(Z�ߡ4o�a�D�L:"q��ʠ�VN�Ƹ؀����gdb ��s.!�����5r���'1���6�U K������'������9�(;����i\�5�&Jț���H4���s����ɮ `�ԻAB�ol�}��g멟�T�@yO���׈wf������ɐ:z��� �Nʑ�	)K3N8�^S_&�$O���#��U@S(��������w����{���Ó��ۣ��D4��*�h�r�A��E8o��ZЙ��
�M�T��",e�D3�-M�������̛J;��gY�jjT�nFn"���_�#9wz"Y�a'��,heMǠ��d�q��#(��a���o5�����59�;�_���� %��n�yv��ыF3�"�ǵ��B���0�g�O��J�Б�P�j��K \X�5�P
�յ��,�0��5�o��� f�_��0�B�cy�;�C}ʊ̗�����<�i�p/;oU�w�|��%c����E����ћG �/
S3
�B0N��Y4�B:k���}�)�i�L�CH���(
��-U��uD#�t���n��ޓ��ݎ�(�	kc�U�ٿUL;s"�h�f��%}���hfiPJX�Zۋ1?A����w�F��H�(��ᗚ&���a�0��8�*.�K3!�J���X6�Wj��";�3�)��7B-�A�2"��Y?�*�~��Jxo�ukm�3�*���*G���[M���U>�LD�y���W�Kc�n��>���z���N� ���S�	%o��߮Q���p{Fi�r���I���xLUS�|��=dia��H�kJL-yl��H�����%��L�3�P���2�4��U�5v~�UϨg�R��ļ�t렓�1R���j	'ş��q�^�I;�1�z>�v���(yr�,���TX�P�/j4RI遂 Z7j���L؞2xߌO2�W��-�,��������n!�<�Z���b}�{0yY2�Qh!S@s���7;�@�Jdyp������r�B����}�:D����oS�j7oF�4�Xa�8Tv$��fn��9bey�q��C,v��K�E�I��1J�}]����/I����Īy�6]�C4��/pM3���Z��;��g�pd����V���-�Z��.�)�$JI($��<31���T��]ȳ���qN$h�,fI6�;ʌ����=Y&,=˾+���B��<��}��^�<�'�"�������=����o��s�Jm2�V����F�h�&���)��V�:R��Z\�'�$�F��ԇ���e^Ls@a,ʍ/��	�������Q��d�nn��_�n��������4�U���������^́U�3/�u�s�[�8���b;@����Z#S�U�&��o
�>��\c��!�L�1Q��uԝ�P[����"�����@ί|0�)� CQ	�زh��'m�
cW�Κ�'��撦�4c��
L�+�X��-%��$�d��H��%jX���������}�Ҡ}��A}��D�R��ϥHreļ��Ę��%���P���X�Q����_u[ w	g��9!??�BH���G�q7�����T���?g�W�!�*�����
��3�Q��@��V�3� �!����,�<�Ld�̩o
�QvԐ<;	2��Q���u��B���jI,���TԨ��<A*��>�9�C�(���_�c"Խ��Y!�j���탉UI��ݤvġ�Ck#�W��ߊW H��.k�<k�av$���&�	AH,��"fճlAQŁķ�+�,�������S��s8�|~�f~��`NpT]�A�#��3�Q���H;F�O�%��u��Hč�W�R?����14�-����?G�V ,xC����)Hl&�M:it5�u�r����(�CV�?l׈���o��&��l �ӱ���)�T�F�x�k�/%��YG��ɍ�ܶfeU��D���:#��t�v�3̶O����=���r�'3�h�!��C�V�9�3�И����ɫ�إb��}}�(�s(�4�wL�\x�0��oγP��C�´'���"�ͺ�O�j����;{��ah/��T��a�U�H#P����N��B��hY�p��vqX*�q"S�a��Fep�d��P�4g4Rh��_x2�'��s�?��^��d��K�����P��=�K©D0N�ؿ˨�Cp �3�T[��=�}xۈM2�w�_R�{�׺�8��2�m.G�zb���E�����[ �7B�!FHֶ�4�̅
U�u�frBďp��|�%�g�b��H�kK�"?���mh1:�=��5ݯl�aL2�spV�L%l�W�q���T�&M�r��8�[Rف<�T)CC��E#q�����>m��uy��������S�^x��6���Ԝ"E՚��p �^��8�[�L��?2��Bv�]�������0�r�V[^S����Wq� G�c�d����3�
�����gP�F'��l�q��F	�ɽ�5�bu���sQu6����^&B������O���_U�1i���a��(�����8)�xs�pm6�A��$r^�M��(G���]�ͱ��Q����R�I������MI��Zjl��C���_i?��5��q�(�Τ#��k��u8�/�Ys������29Eul��#)�{��,�dƺ^]��~er�;��>5Sh]�<\m��J
1G_��l-g�E'�� �������J5�\c_V}���I�2��~�