��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""���᤬����[���%r��e.9�=d�����P��?�^c�׃�ƴ$��`TVϺY��Y��8��D��Z��n��S�L�o��M��
��چ�Ə�!��mN�X;A��忬]�5�J�d3���_'ˇ��쁲�v��ӫ\���1��|�(��MrV�*���7X���O�
��O�-i���va�k�RO����N&I5{-��v����`Y��埱��gX�ی�5k�	Ndt�8�#2XE��OL~9ix�`�N�-�&KsuA�*�0 �\'MɓI�?M~���]�P��җ� �G�ѱU�C묻<Vz�r�P~��U��ĻyKێ*'��o�Pl��"�#1�e]N��%��L'n��'��c�]o�u����H�݈~y[��W�bO�v!69%��S��u�wF�Z^�v)�F������$��x%~c�#��oӣ�����Щ�-;(����(nj���,� B�c�������P��:�p+֝���QG��sd��4Y�{��������>�U���YӦ�������wsL&�W�gm��R�|�� �2o�f��ƫ��{��vn5a�j@�o���)�`�*�?ˈ�Z�v�l����q�Uh�O0Wl�`���`_�\0;�����Z��e|·9:Mq=ܼ�\<��N���V���]��Z}��T4U�'{��8ǹe��iu5~&9>7Yj����F�C1�+�/�v��'�1�$�kI7���!	��@�0�G�f(.xlt��U|�,�%��8�Z�^۳�?�3� �ఖᯌ��1x҈�VE��Á���8ϸ�T���C���R^�Ϣ��QH�?�'O�!kd*-���=e�U��T Wn
�Ugÿ7	/��^R�bybf�w�����%�a70����Z�:Jػ�wLLlf�� >8��Jg�'�c���*Ա�\�[��V�,#Pde~�ds^3$�Cl�{��%y���OY1>��������Qr�X;���3�0t���V`m(u��$� v������~x�T������ގ���UMN�+?Ճ�N�k8���"����6������/'���2��V��ڗ���X]Ϊa=��o,{�4?^jP=		��o4�b���(�..������踬ëV�Xu� #��������t��� ]yQP�.�����7���[�L�T����n �0NǀFo�Q<�0��`��jCJ��y��$�+�@R�0X����'��D��*~
&����L�j�����h'�"7��T#�U֞��u5Re��ﮘg����YS��g��}(�����fM��FZg7���� z[q� � \�Pwcڞ���F�ц�44` ib\+���'ɑ$�D��M�O�d%��e��>���� dܴMo\����C}�N6<��)N`���Ӹ?�&>O�r뛥�
��_�� �UZ�77��E�"h%�^}��|^���uٹ����/9��� �|}���o����p�T���68ؚcR�J}BOn�c����[���[��t���"B�\��-�tM�A�C�ڍ�[��4��"�E�_�� t��[���x��Q�3� �������*���V���d���^��aeIc_O[8g� ��j��nݩ�f�@�G���9q�$U)���a�<� ��u�ljG����Ct�A�/�YGҟ,��ZQ�q�W��/5k��Ac���z,>t��("E?���ɴH�cd'����c&m�MQ�*'0]���͉ͬޏr�D:i�7W������`B��q[zr�}{E6�Ī������}���A}�O��NQ�~ΫÒ]fitfq΀�'���(uZ�Qġ`��}��R��'�7]�+�8��o�.�
H-^.E�k�D��66Ob��i)ο٠�.�)�[lq�6B�O���%[K˪���U#L����`b>5-��{�w^�CU6e���5��wN\`�^d�h������\:��LXB�`w�:������I<�֫ж�;�װ��D[:�1��Ű�%I&<�la�Ɛ��6V��T�ZhY�������dk��'�s��J���Md��8Kf`̠�i	~TL�#b�O�מ~�W��j�P�Ó��$������үX�hxdL�����ZA)�ț��pH={���,h>w�4��3��_O������!��G�^7s%:f�[�;�\l�\�Z��"����+�nG%dff>���r\ng�
GW�?�*��~$�'�4\X+jk���E�ĥ#%Za^ʷ������%�sn@��LP�i�4.�US-�SC����Z�Z��9�*�$h��4���]�5�{�j+�������l�nw$��	#�Q�����OZ^	E/��ř���pIm�`�*t���M/�z�;���;Ĺ}	�X�M.oMZ���ƚ��]mg��[	#ma��`t�s�Z�1�~0�:�T:Ü��lZ@Q���4�7W>�O�@���}��E�(��Į��d�*�3{��ea��~:`d��x
�b�T�C��e���T�|Nёy{�i�����Zj��{��_5��\� *��[*Y%�`]'��
7���z�ԡ�ڡ>:�W�m� �
��8���ˆA@\���D=�{����o���c���gv�yZiqŪ`k8Q���j�|/�(徹4��:�����j����8�ǽ�HnAz��50L�y��y��7���V�͕� w�����~l�4|3�f��%�M��K�M���Q��A:R���x�aZwV�FXI2��Mg��6aos��\���ɿy��J���6?�`����c��@=@���$�UY� �xϐzly�8��t���dƢO�)�����ɧ* �v���WFN��/���ڱ
e�WLP���:�M���y$��qCi��Q�$l�lZ�{8����^SŤ���N�@W�ͽZ�W�$�W1�M�_BII>�|Ԯ&�Ь����_'�����k�_d*_�;Z�\@�Fy4�8/?�ٟ{����#��t�g�����/����\1%P�����&��O�;ԓn%l��l#���q\Xwz�nn:�8V��v.ye的����-g����R��u2�|	z*c즵�ߜB�sN�~�.u+l_���Rm�;�.�~=
.g�X�\��uk��_���e�%S�@�X������ �D��mFEyi��L�I��쑅�0pxV?%���a��K�)�:���d�3��|eU�;ϭP�>n[���Z֞�a��X�n����D]o�J�5JzyV�n`��%Z>��la�	�2�ҍ�|%�isK�1��R��z���{�֔%�&9W�Y�Y����[�M�!e�ccS�X�֕���IxO�Ҏ�/zpGl,�q]��Λ��������/Cc������%�ڔ��K�iR�B�������ȣ��5{�k$>r/a�d7Z������C��8/~��)^��w^�[�JP�wa��Pӧ2���b�L8H峋7b. d��[
�U�NRX�"���~� ֝4�r�Dz��p��ʰ�J��'Ѽ�[&e4	T����ص�!�J�d�a���4�_<��p.����HD1^h�����X��:���1��9p���U��%�ծ�&냨3T�nYf"�>�
�����Lup'
{�TP9Q� ���`vΉ��P�]��,��I��;X
s{JD��{���A��)�P�!��&��6mO��;���9�RzC*S˻����ݟV#xa2��$[�����}?Ɩ��,R�ج@����V�����	��*�Ȫ��ٗ/w��4:=�)5���*�[e͌�R:�<!�������n��ʭ	&����g(��W��>�Rp�#��$+iq�ί�]T�wL�����A����[e��pZ��,�b�j���Q�%��\o�b�or�p�,]i>��.�gm/�:(ث�Nn9yU�/����q[+l���7�(n�_\>��L�@���aͿ��V�5�%�;5N���H����C��5��ox@�utU��:���k
ȟ/�|�|1I�}�'ذ(,U*H6Lh� �(��@�}9X��k*�JV����d^%�8/�h�z<�N��Ngǥ]�s���y��ڏ
��-+���c��qf�����k��ϖQ=O�5ScH���h{� P�}p#�2buw��~mTW�e�-��2<L �C�[��7݉�7clwE�=����9��۞r�6��y��ӂKL���	zI���f�Mł��/�h%�Vr�D�KyTl0�]�����o������R��QKӱ
��o�r���yɭ����Pg�y$楗���X�j�%�#��~���q�}�׺�[�r�	�������"�!Ӭ&��=� �*�`���+�j«â�/	�e�[���A�K�����
GU3z}D�c�=�N�ܵd~Mx}���<8i���AHA!�}<�m����=1(y>W�-E�!� Xtk}_[xO��n����	η����7y�t��EjJ�j(rz���)"����'ĊI CJ9�xm1����"��WĚ�~�I���t��=�9�����Z:T��~�FC7�"nPP���#ex���Z��uj�$�R�:�>>��<�362=�;��������(�C��]���}�7���,&�d������X�P��^��I+ ���:����;Y�[0N ��x������m3��W3T0����N���~	�B(���>ܣ&����3G��S��V��{pC'<oLK@u
�.��1���	��_i�T�J��bE�;�fY��8��W��v9��1� f�,B�o\:�ɢq�d�>����08�D�A��}u |���Ġ!���uwZeu4�+Z�1@,B�	mT����9:�؇n"���hd;�n��2�KFRV�Z�~Ɔ@y�em˺ӽFe�{�[���gd�-���31ta��	�tGy���kK
��A�u� X(����}�C�����Y}]P����]^c^�J��#�!���5�v`K$��X�x^����H�XN1� ����&��x�.�o+���R��]N_bҭZp�hH����l�R?��e��I�O{�Ӡ��Kʒ��dsn4�#�F���y���sb�� ���U�H:��<�[ r8C�8��v�]�k��K��|�en�R�ّ�;��?;����Yk�}��}�CX��	 5�� :�
G�U���a��#�t�M����8�ayn�b��ە
e�U��e���=f)ERO}y��-`�s�7�ڗ�=0��/����eHSѦU�/ƫM���K��w��q�:O9���+�[��c)�$2�{`�aUr>�vį�<ب�t�
�Q��* ��!ϸw2j7���+��k�jh�S��Zfu���ÿ���v�xxۏ(�c�����s��_���V���D��*\V}��YE�h����(��@60aeJw�7��*��Z�Pcj;A$2,�����|c�e:I�̺����&�V\�@V"~e�����Q>N���+�$IȨ��!��P�*\�_43������Q�)�-���̇��R�>�(C��G3Su$%g2�������;�%'���ݝ�>���/o�#=��V!euEiЕG���|}��M���7q�P	ד���$Vڇ�TfŖ��lrp�c��85�b���Vfc�F�lb�����H���50Q�cb�[X��y^�~*���Y���B==;�q�2��g���`ϻ\Sy8�羻?�|�)Rp��		�����r����@��
�Yc��R�U�z�����
U-�]Y���t���r@�K�_�5a�9֭g��em�:�	FY{q5���MF�,�%�(��u�-e��{&� �3�M� {���ԑ��4ɋʹi\DO�aL�qm�r��hE����.��)�m��c���H�q�u�vu�c�q���b�oQ��t�8m+�oT<�t�
���}��%��[�j�:�lr~�P�z�o�E����T�q�[i��+��R~�֐h�Q#�c)���
߶Vƾ}<ٻ���C�}:fsr�6tm�5-u�,��6�2�/���7P�mZ�V@w���[��Fʽ��7r�XW#�?��O�@esi<gָ�v~-�H״Y�×6����yj�#�|ⷺ�w*a�5�dN�4L�"��)`����f��x٣��^I-ޑ�6ڤ�6�)��d� @��
�t�n�|Uݯ0��`-e�J��%V�=������;8λJ�t'C���k��ɚ���lu�ܗNN
j��ֻ���~�m�(�A��BD�E�'��o~Um�� ���Sr2�F3���ܛ�[m�h#�����E3����pvOI��0ׅ��g��;1w�'	��N}b��/,���M�`zp����W���ٓ��D���c��dup��v��w�;�S[��Q h~<K����c_�]ȗ��p�^���f�(��\g�Ԭ܊e�l�
Y�`X��̖!�jФUN\	�u�1|���h�@�$��r�Z2��HEqx��|�14q'V{�d�8��?�Z�)�1$�ED��@��қȓ������?,��kjc���N޲#��c���A�9$4��a�Z}�hM�n��*bC��Zd���k	|ɱ���#C�d�L���0eXe�s�.�Z3g�bq�P��v���l7�GK���oE��+�O�%�h>�{ǧ�ۈp���(UX��z�]H3�RQ�SO��t	�s(��r�Y�7�����L�z:x!����|#�7����f��q��#�J�l
��Щ�
��X��%��Ǘ�^� ����X1UR�T�2
���+;{����Эq<���S�!��2����|�p5L��}o�%5Tx�4�i�T"2�5�G�k���qb<h�n�_��aA��{g��������"HQ�����]\
 hJ��t��Am�vae�áŕE�v�[� pp�,멓�pL�goA���>�p��娾-z+��7�e<�4�ڳ@䔢qh	��P< ��̹�	LR�?���n�M�[ R�*��r���Xy�v� ��]�{�u�EP��^�c�0�4�z���[��7_T;.:�q(��Kt�7�{���>���ط��­cB͇Qg\��I��q�3`�}��gW����&�9)��*/�0;=�Mݺ��P�Okv��^���o���܂;町y�W��$��A��奱�/����I?^d-ëB�;Y���/�ޏ�L�2�t��X��"0�Z0F�Ē�&�1����f�|���dY�؎ņY��m��$HC�Ĭ�\�LP����cqg�\�m�ʿ��w�K�v��<�z/��V�\�Vα׍��T���S��>�)��K_^�� @�jY�D���OO����R/�(���M}�ދƀ=HãӮ"�����l�ͣM�VJA��=��>4*@P̹�1$u����{>�a]�P�.]�>����������k��23����b��8�������5 ��6�[�B;|�]`D�k�w�(eg�P�Ֆ�p��h�Q�T��r�q�E�]R r85�f�@�vǰ$�5�v�B+�1�_�h���ړ���
r����ۜy�E z���P����a�~��u�62˄�6l�gN�L�2~�J�aa�F�/���#�x�&�7i��9e1a������|
r|*�mo���ٔb��{���^��e�{��+�\#Oe���` t�_CU�։\f_c�X�k	`T���~�Ӕ/�Cg�$��Z[�ԧq��.��H(�FJ/?h��:G1Q��9�́+M��
�$)�0�ky�b��8j���̺0 6Q����ʵ@*�J'��~�H�+�K&V:>?"RNh[r��pnT"��䠸�R�����1SP��_�%y@T��� �&&/�Nk��m����2fMʈ�"x7��,��г�E��}���gZm��P��q,�|rv�k�Ś�~�ڿ���]_��J&�'��4�Zd4���im5<��Y8k���������T�/���Њ�ű��%���[��#J�E ��m@������d��l�%Pr�A�Q�6KG����I~��
���Y��o#�rU�2�@�����*�ss�#��e
�-������U�'�'r���3^����R��.;�p�LrǱ5L{ˠ#���V>''��Pt���_ͬ3,\��(4F�Y��#���QW��:�/����35p��~�W��k��}�(����L�6�|�|��ZSS��o��;����m��atZz^�C��(q�z�oR�(3g!�f�,)�2y4:���o1���������6�'�����'!Qm~�e���v]�n	fۈZ�՟���Xڲs:	P]Χ�����y#ī���R���ؓ͝�s����p�L1��}B_0ڀ OF�����D>� ���6��X/�-��1ԧ�����e����2D���OwT���l����̉��9��6�<�{��Ɉh���V�D
�'1�VJW�y� ���o�XY-�]h���*�r߾�*�\I�-f�<kO�H�=oI%S����Dɲ��T�0a�sv���#�t-����'G��{�s���qZ	�_K�����F�L!����*y��#ca� ƙm���oWD�?O��w�Yͺ�Kٵ''����S+�=��>�R� M�.
�V��to�$2�E�c3�DUt,�u�CJ𶈁2��f�����e^��\��0�<Ҫ���Fy���t�bI���x5׃n��"Ju0���3�M���=/���P7�r�_+�R@���z��k�8��Z{�l�73��fm��X���ͼ�Aqr�� I���丱I6,�����x�0��K�;�W��jh�K��$��ǰ��l,O�L��Q��qG��g�����-���X�6�|q\2�=%-������b��dr�֕Y �����ԼhKݹB����߸�L��~d���F�1�݊9Q�ES\ӎ��h��L/ƳS�a��+n���!��DP!%L��%A�_��"�Ԣ�W�V��~z��hX�z��3e�ҧ���-P��_`:�cs�o�.�Yf} �칦���K�#������l$������@�!)?��M�+���M���c�}eG+l1�d �~uL
��� �ȷhZQ����@�b�G�j��"�c�[�V��;r\�5.�k5�m�{�R���.Ө� ̀�,�X���ʯ�=%���E�˶-0���4�cSO���r�Z2�Cֵ�<����D���e�؏�r���z��V��K�Ҿ�jު���K�(荗�e��M���A��/��C�8�� �X�\��q�]9����",
H^Gfv"��]WIQ�֡`p��wK:B
��'���׫�{�i+_j��D�s�dG�z�h���w�������M�����]7��������w�D �eHl�Bʵ�5`SQdR�ќ>��t\`��H�P��tW�������b�jXZGb������Ţ}�m�m��Ov���~��r�Gu�����IE�y�v�8���!��\�x\��7���RC����Y s�%e׸�B�����ˆ��A;���d����ȥ>���'��k�6v��N�8!��s�Q�sMa`�͗oR�HS��f�γ�ʽ�Qoo��r�?e�Ńn��vG��`����		�*Xj��a�c7a ��p�{��VUOG�Ւy:]�-�9突_B�ǕKB
z7����x�V�qC-�k�#N��i�yb�2y��L2�0�Et`��Cن}^͘ix�~�}�%�