// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:37 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JDtLnf+nmTy1In8tkKbWg0MepXt9haFjm735cD5FgAm41oQQrX7QwziSFvcMWhMx
1/MJNJ4Zs4K5cMg6b9RKy2+y/QfwpiE0AuOWkMMfExz+Cjqor2P81gBwDkzZ7iYn
UpqDGqxbvX4H5BWACzgHwjGK3ZoZibyXyeOy9T65La4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
G9/YVpyVhFlUc3Cr2irzOVyd4I01Qj047Dygr2EjGdosuJZ943WpvUpRSwuSgR+J
haOkmMpm42Ju2mcMgWAlyt2sCwz0MlhT12LVQUoeDWY5joOF8HFRYQ1GtGld2sAB
72Ld+5pMEj3kwwyluOIk1P+E90n5zSlVqi73gujyN1ZoKVvUSpKtTDqClDj1pl/7
Mk1cjs09J1Y750vA8UeBqEkzU3LmiFxtoILyWXyXgylj6E3dNmjhDJaBvrrVu0qo
TUel7xW9AA6s0QZ7ytmQoP9i9by86KlaKSmBL+aDBFNvzRMhuqjXDlRjNBwv1Xo0
o2XfXvFc4vV+eKk1yXKL5N+Y1sZ2H3H2oQOdQJg5CjEPe1ooh5/xOPVbDKFjrU9E
VSjjTAoqO9YYdNpdOD0gzXCnDAwpbm/JTgYQTLsQMrDDc10ckAYPYVhpT3p5FhL/
W9tgULn0DKEoE+XF7+AmI6C+vOwgrFi+bBSoexTrevBlyKvQpzlYnbIS1rXxoHiu
0NosT5arrpPqNAwXWSfGqOhpwllHcC38bUBPBvcgww+wzE1NaDUTC6rB7v1cTN+0
ItxrzIge4R/tVx2SSspXXgIPs9I21uXtoDmWLve+o/MYV2YMVf3/S4hHHlPKpx1e
H4tMkDxW3dbgj/s+2+vg0mwt0CHGQL2/E0B/oKRXu1nBLf/OFVKKPr4zmGBJIPZ6
ypE1Itej5P1MRSHUfr2VVdicJ+YQwfEuJuT6UV8tavFnA1nLuopJnP5ttjOl1C3f
QGcYrOtxvKd8AB28Qw8fttjGbQadEmYPRiZDbs7KKbjzWDK6/7W2YX5T9wuSSgYJ
n6LuuOqpKfs/0IaqkGpZdrFGlQkZ5BoJOC02XvrdB7B1iT65Gid12n1oiK0ZAt2g
wtZpgrlQXSnkeK3xrVEpX7zFSOrvEA65VpXz5//oyrVAHXHcgQq3nkWKHq4Kz8zZ
g/lq9gp1UAgYyY4UKdun36m+PwcQcnhUeXQZ7SlU/5zw5+6oU1YhvSOQsfOjgmjM
9r4AUfVqHS2yiMRhViP9hn0End3YDTWI70+ZWK4aIq/oJOlj6oKQb2RaCtokkY0W
sCkuItBQo8IKTIdGtBwvDcoZFdDp4TySrR71am9YI/3AisdrMYUiqBEiW36NqP8v
UVXFZCyu9Sv8lGgiWyhtPntt5pIhwVz6FluHv+ys8Y0BrrTm1tONVF7e9lTkO1dt
++P3z0jX80K3oC2BYb0vo43IL1JAqwYIHzCQZ1N9CgOzaxG/Lps3F5S4w1gN79w6
y1x9BzNj5fLJ40PAs7rxJslwjAiY7E997AJQy0nIZjf/lIIZGoG1Ivw6Z5Sq/hOP
Uqe/IOWzGHABeyfX3bo4pGORhtUr8CpenKIxSBdkjE45L6I7wR+3MtZYMkgsLlIo
6ElNZ9b96ZwFiHJ9ebbRUS0QB9qLaC3ptbYD9tDu85EgKAmlXjQHh9rTRuxBTkhx
7Dj/1pXrTfVHgp7Ev53YDigcV+KSo7+lwIBx2CJXak7IYSRWMLDcLOkxQ0e06TKH
3LLa9RDOWnuH8hVRY/2HCmSpf/kBQsPQt2X9xggAbW/htDPqoFOBO7OOrm/1MzYm
UqCRk/QeCLkEDjPv3LinnOrdkmJwNsNUb/04t31y0Elo7Zev5ZkwSPwSNuxsKUzV
ZTZ5/PeXMuLkQvrs1nCiXkr3BrgeQsQzqDJVfvUc4xZEXgvO9Ice9k+oYNO4kzfy
5kNEw+AtyVALoytp1p9/yQxRjPMNDI0fHdTLD6d2SJVg+J10lbssBN8zTI2fQ987
piY8Y4MxpUiR5NG2/eQjLHPe4+m7LrzSULaq/GnCz3OMsoznI14+e03hjH6WJH9j
vuMfyvz9lQxxtAsXAtMrAAUdOWfq3mZ7KY6UgDwDx90GRCUd5dPgHRvKesIxjRH5
xUEKjMtfJVCJwy19c4vtLPkET33Gi0jT29KJ9426bzz89Qg6QJeOskZQOCjTvXYV
zk46repYCJA5xVFzOyFcKdKtlFGuPvC9Uhu/lESgk5neBwOHhAIMve+SxEJtbz94
78DDr0P4wRFCfv/eR6dD/s/mCyrBHFJsvG+y5WuGo2AoDbeOcqHNhzITuNY/P6dO
zz29FfOsfYnZRla1dcu7G+e71r9v87FteP8gNcgO/xL05DJv4HzYADvWEPwGSRYL
8gDbB4B/3q7mQChkP6hQOAdAU09O8MsAYE1+V+UB9IUTW5ldHP7SroVLTqfofzU4
WQq7ZaXZL9QfshXptIAAmXs7McGUzhRPgRNGKzIiobMtpMgSWjYxN8LB1ndtw8hr
6AT/I/KhrBikyjLsrE9+ZIaE6J9S0oZYlCQWFEMpba8G8S9bR8k5thWVV8L0URSH
I8YAgMMuzMrbKN29HKO18bMJldmagg8Rj3orPE3guE9EDqz3mpWBYJ8ytGVY1Uhw
PawQr9sIanQdpbYPh2KVT5qmsDvDF0XgYL0udKqRXS3JAJobCtF4Ra/mpH8us0f4
1VdXNoiZweJZiXQeAryXlkKPGmkDv0kqU8m5h11rQ9j2EnMIBFuOTE6BJxpUN3Dw
XeGmD5SsO2v4iqVXzqX1tn7owhj70LLNSkFwa+1VT72eE8cqyVjl2ZshQqfeQtBK
CQDfX2hmAarl2aDmPwvon/YcsgRsu2ZURQRjVoNGmb3ekLJWdnrZmwD6f+pJ1u6Q
COD34V+fyDemKJkL+basHGwMlxPgrbcY6FBwWqrXKRQM0lxQqoKKKBq2RooQLlwg
rfF7wBvPZxcYIaz4oE7aIXQQsqtHyYOm9XMghSVbrR0t0/860CZyeQxVVoVHo2HR
4iSiUUkLr7LNED1FOc2VJruPnR8av7H7Sm1yalovWjWAMe89N2dMoCWaUpPEjz25
N1QjrZbHizG07egBkvqIz4L8Rii3EukiIxFoH8lX7P7eiIvp1i18ole/NWy0d9JV
m/YbSta8R4NQzh0ws8Vloe2iC3wCW+w7Ouo/AENyaTAarFRExwlzTvx1gj+5OBuR
LmDKkKSiUVlHJSbytb46bSL6gcxymhMQ6DTpVMTHwDHP82hPL8deEjkiqDfbCa/q
d5KhnIMxVYiLTaJuyuunYGbFFBzuKGqGh6+e2YTBXao9OjPO8aZUdz9xfT0GKX1W
i5h79gu/JyaGCo2HETYvoPbYWBmxQ7nc13wIkbZFocPAjKgGoiUhObRA/agqAYAO
KWbOQOW3W5eOA+o/p3a+Za2hq8PrW0O1MRPGC9bXail29Tikya5sjyHzR+YxaJgq
rfD27bPDsyi1wgMbS4OBwlZg8GJGaId2gDQcAzot6pQG5yXNFIL1I5uqYdYpOg5b
sHOh68Qfvp8mHtBY9Bz+e8w8xXeEovCk10CYQN0xHHMCAOn6nG/HeziAUEIb9l8b
UdaX6WhUYOu788p+mHKJOg2mq3LtTesvEZy/d4Pod1FtNm0qrxuPj9sVhxfAj+76
4+fjjWRU/EueYzBMLQHCdKRKwqdzytV/w+yzxnwAjxLCY5M7vd2YyceMdsGTr46L
QbN7tcKBfBG+FFPQU2N99sKZMhtgc1i/5K5dxqWMAUD3/wohlcGVK99WuiL1AaNU
kcstHbMzBFDhAHDehOLKYm2iuNf+EUg/uwX8dHMh37F8o6ZN1SIYgq6uzvJzkQh9
SPaWuXTs7w5XF2QlpJz0xZr5Y4q5oBTLbWc3SgaBBOjTmrIj6aaT+KERLWHXiISx
SXxablbZpObP3qvl11EFG0M6/pbIG5EXOsjsT5VaZVk3Urd+NLsjEtrANNnm0mkL
0AjovToAZBnjk0hn+gxz9cfzLdyNaAiyyZ7XLxS/McgUKycPyVdrtkEuMir0gWaB
0cwW/zG+a4L9E8H0Rk7VTxTTUAbvuMxMG5nhvYj6zFFMn6qkqlQhU7G0pMM9bia3
2qeAWZESl8r/k1q6PoFgxC0ptRjGVKF/Nmc766MXvwchKmDafeDbnp0fe93DO8Aj
4nJTSJAiNgQIYYdKpRsREBr95NtMz2WsqRP7DUq5bOhiKh6d6l6R9gTM83XXVNSd
FX8oKDAJFcVzGgNdJ/Xwux/muGvnmgYJK4njoyAD4RTVGqqjeWCtuT/dO/ph9lWW
bTK4Bcqcnyf+2XdVXZdZ7Hrm2I7G5AX+rGkwd5d3MF+q2fVrryeAeu8+PgtYVT7y
iB5XvDL8aK6sS6vL/jwOAMXhlz4VysNt+939jSf+3TNIIk+LUlMT/hQLf27uEk+l
Y8lm2mwrYv9VaDImW7lVZOmQrDS+GG6710fZUABGeU8wXv0+oVUHV5DwZ02GKpm0
ydb4MSXJDbd+yDUBZk6mGwtcJ3VIRKeB1FKNXAFI2buW5U97P0CRhaAbO+zFjJo6
MPou7ihPT+TmNpGZHI93nfZ1ZMP9R+7TAjM9Z61EvHzq0cy+6wzjZP4KB62Fs/PF
5DO9jr1dKw7somj0xH0bcdi3g56dt6draK+wKdukZAcK0g9LwAVkgn+qFjGgbwtH
uINA9koCIpNRb8eRUuQzSKaJjblgOyjE+/YFs8Hhm7QBqe4P+vdbMJzIR8rBfJZj
IH+N42GHQFJXP9fQKKqf7LuTEVtVl2CmaST47GO7P36lLsLmQjaUMqE3dazS5tvD
HvoWwV9dww03jmeApmeLAD5s80TSL/mJHB3XvQh8Hc4W5zMKq+rf9moDK64J9j0K
Az8mEp2BpDWqql8lGZLiQOqLLNa7YmWABMg0a5O3oAEarkJOR5zdL/+cfa01pvqb
HzXdaG/uYKo9CWBbI87CeNTZBzFzbzO+a+kj/oM0t64XjJpafFfH6gIw5M5Xzh8h
UgLw6o01WMxZBaO4kf9pnzD4OaeClU105r0gs8poH7H9sihVucqsk1ArZBQxHfeZ
xZ+KqElidrsKJiuyegm34Idy1f6LnC2JtyGKUH3A+tveCTM7GXRTdNx+s3NUAq3K
EEQceKTs4mpxUHd3QuKfO1OvCXjM/rEe09IbXMDTNmgeM9UBrnd7IHwDYFBFFm8x
d2O7Nn3rBC8WjO5sLrjjdo5CUMNOZmJkelyvAmJqfMGUU6LNPqdhsGzTZyHpMG6d
P45JeXueLE0jcgfsVsM4u0IcQwpx7NRUEYzlGDSD2erRKQtv0Gfts+Orto67ukTu
DF94kGtpbkc9+jDbbDZ5Kvxh1BMZDwSgB4Eu+NLRDxDj3bowsAR5nvhYvH2ypB/y
nc+gmJG7qaDZ0NKUlxNIDYlPbiEcrnodzYt+VRNxjBX0OFd6edSBR8014aJ2je70
OVw3CJhZVx95aM9RLDXfU7mMgjumoLCaVtF4fjGf1Ac8lAqTQ9VpXopbEaVkYT1t
IUKXzmFv504XTVJJKUPQwRYISzUhHu8gPLVpWKv7uLsqvFnZRege6NQ/HqPs8h+K
qS8oeytw5r0a2XHtgeagpkb0XgNiHMUN+VgnZJ6OyihradtRk6kZ2eqOOG7M2+BP
fmysn/wq4QN4nhWTv3rAIyAYIuwtke7UhtkHVTqSbFveminnVTySW9xe7n9H/QoP
uGo7sAA7w+ubOAa013ReAWUEwIfj0yOVFxZuT+JDH4z41MQrbHcP76IOgKN3Jbfh
8GakaUXPUVTfJrfc2GFEZmAC/VgG1wLHBkOFa3ZENSXBC+6AQGpSP5+aw+pEcnFp
pGtNa9V4x3Zahsibcrv00Bf1aeWrZqKd0FZXBgaE545RnG2F5o3iMCocMDIbhWAP
VBnavQENl0ESr+m3WQ11BArB12SGmAfLdAN8O1PHeuNlAn7gUWC7Vo0wWf8afeLc
8dvR5HdvPNGwUXxj2bG4XiDVZHdTM6dP8r62TL62Of8p3Br+kkFrgJKKprjr3Kq8
FskDDuXgJje4wMK5SjCcnXmx/IQNehfeqw77WdiOcDpQAnUcMezcG6QOoSew1tYO
C+ogIMb3VG/R1xwRHhW1oMgOowGoXf62eKsSDrG6tzHvsTbhurQ3EvN/hIW+6/HU
tHjmWhzz8ih1tHKhqJ6RWrB5IXOI/rlVz5PrSSehLc0ljbj5GN676UPDUBlEIUCS
yylzaHNc/awFi4tUZyWiO0Q/H/jgeO5cdFZNnr4ob5O3G+lxvMxcqC+4nrFBIA/g
uC4zfB4VApdx5bnWp1PKvUcujohEozuL+B4z3d9EyvYSQc1B/OnuGXHQtAEZBRSb
HrWWgawHJNUqArFe9NPi0c+/Z3LE8Shs1oHP4Wa9+vj7UsCJvasCoXETPqDKtUry
lPki6lV6OkhIsiffkWyGx0OX2E1eFvlQM5U6KPibIjsto7l1SREDAixu+edsm8kv
8xyCa/LIAPKEIA95MKDnPluuD8U4vC2qSahH7+bzdA+cDQQMiT1mAcszelffK/LJ
9lHDIrbAL3/rFu0Mz+BoML05Rd3M6mAY8KRVb4IQOLzfOxM3TxlCUSo7m6+cpxiG
Nxqba2b8VAnie6gw1NuYY8uiJXDfjZoNrnvDT1ZWvV++TBI5dBtteFLfyOonKhgJ
YL7RG60mpXidgkWnBgaA6v8qNRmEAfc6PK7Zs7nps0SA1a/xWR66Q2/v+qEPvrg6
3pRyBmXGGyLd8BCh6QO7nonVOq0UU9IRYwu0AcFEvB2ykgRJUAiNV3bxUX/lk4yC
osCOCNf/SfNm8X37BiBwf2k1ZWSdLeiCPf0cD/HqIr2V96vOwXrbq+7JTMqSsNSw
YPsfYmbmFfQGlvZS31pOms0jRdX6biLJYPKK+MCyTM0Ec+DcP8y5t8LKY9xvkN5W
ChhACYtHhjkwUy7/FElOz2pnpPxvQHfuk2OI4D8Tydd3mZsdgTPy3r6XKAc6sKoV
m2uNg0ZjLp74Rk2eut+amwYyUBzZNIpNFGxzyWAHoHQBpMZ5zMLS3Y0H3138gTWV
lT9WV02Ei+DPgbyWc+E5tkef3MWBCza1ED/K/Xg7mJB/vYSRYyOsXVYzgCzlr909
nKqlY2jq/lRRQyGoQ+sYJeCer9kuoW+hzkbpdUb1DFLGD6wOJQ02kYyEiCxeZcPn
6k7UGXm0tgsr6nH+/JEB3ODiM2hKoYZBEpHpPiw98A/0b+BcHuycxkdDLgrCBXuP
yxxg+Bb2Hju7uPCatIs7lZhRGl/gAsbxxJCg1j0CnKehovLKUEt+7jS2NXylwr6o
brSiNei/2RD9+AF30HUqjD9r0M51BmjltNxBlhsRkkPenytseODPDm40WytP65J9
ANF1XIielu9yrBXRxpcxKiiuaAneypq4VfwwrOcMJd/lJfOE457dCdndkWIPbwRt
vxJuIvE9PBmUjnEl6UxsEB0iiVi1kzDNNpjsoVJWYiR7R9lsVfFW3wKPggLvuf+b
2k93ZHj+YPuqiWYdxMlcU4CZyn5FiSFe75YamOEtq+BLuEdlg92X2aLgCrfHsZQX
GkyO4ZTYRJDN1J1dwxF9F/llWC8ko2zIPe6g5HYZscQ3MagjlN+w/tDjs0l8c4Q0
J63j/lHWMP1y3h1GQGOqkN0tP3QijgXtnjaRJnEc12D2BJ1bfFOLoYOmgq0+OCgf
M1QRZqelOsGXqMTlED6Tfg6w3fCwRn9ZEaRcPMUfKm38gz9ppDO2sjna2dRtCa/B
zu+Sl/K5wGYygYLazFwTIXccFVQHn6Y8eHbE6Z8UI1FfRi+ahTM7uoN+sO5k7Dve
dXrTR1ToijiW4Tso90XcXQ==
`pragma protect end_protected
