��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ� g�I��Jw=���c#hN�j(r��Ҹ�@��\D���˶I5U�q��֋�[q�z��t�KJ/X�C���D%Վ�����p�s�m%u�5YX*w��e3��N���@�CȄ���/�7|�@�GuP�El>9���CDF%��v�Aj"�_X�m�O�}�QL�3�hٝ.�Qe/p�)5�{�vr��șa�5�*�D������:�{�pm��j��
I3:*��-(s�@ٺ��YT-��.�$�$�fu���?��I���tdc��϶��#��q+�=���,��V=�s���L�L�WI���X!��}��l��)ZW��J);45`����ffe�i����щ��@l��L������LgT�F����6j�qr��)q�u�JnLM^j{f���>p�����|-���>���ku���O�R��xr�5�
f�LRC$p�/������|����x�.�?����w1�܄��C)��O�gڣ%Mep2��Zѹ]�A7�[���9�i�����V��V(N�z�������t�/�������!\�<CRZ�~h^<N���y�n%S��#�և���֞,��i�����m>x�k��Q�y�t�#[���.�;G��/��dSH��'$�K{.rn�x��K�B��໌^P���$"��IH�;���R٬n������.=��EL����{�JE��UM%��J�9�Dֈ-���a-��)�i��ѫ�]j���� ���ݙ�a{^�}I���d��!TJ�w#���l���t���w������F��(-.�8�f��Հ.�,$��ʥ-�E?ʙ�)w��9JsɅ��"�2�'��qA�ƨJb#��S(��+l��I8�'��gh�&�{>h!�G"�5D��!��g-.�p\�.�˘����邖'�cMK.��5���0���qn[3�6l�4��n�%;˷�;f"��љ����^eV3���Ɂ��yrǻ�����X2�F� ����cj��v��d��=$�������{��_l�f��	Ȃ� u�#
`�x���cnڝ��V*���	�2��-�C�P^�S^DS��^@�g��r�k��%,�'�-_��8��w`�2� 7����@9t0_�Fk�����z/ ��s"���$��%bA���4�+ԙ���B�¾�`^���rF�^��$6=�B�?��;�+Ҿ�v�C|��.�d�vs��"_gc%����)��Q�$�Ms�$j��Qqq�揕0��Wzec*���H��� �b��Z�D���M���2�>�?j�K�
Ldì�V��s�$Αv���$~e@��^>Q����-�܃�,-+}K3tf �z�X����&�$�v�Ww�h6b��0���5�|3���<�ԍ��ڀS%/�˩�V�����.��1rA�N��D 53r�:�0��
�3�Sd�<�S����x:��O����L§Ӻ�l�M�n㩆D��	�V��Vڎ7vYʡ��}�������_�l܏�k�C���_����N�7׬q�o}X�)���u�Q�>rC�{��,�/u2V,��4F��n�2�.���.e��o���%;i�zf��j�k���b%�w�{u�!�^8���UzW^�=���f>� I!�����g�����w�e�N̏�AۋD��aK-��h{�ǈ*a�|@x
�K԰?��X�HX�:A[���T��q��cC��,�_�ė��|�E�q���IW�X�ӻǱ<�mb*p�����_��� �d	;����M�C���'�ٓr���L��HKC�+����Sγ[��ו$d_=�=JQN�-h�@������ �{����	>�n�ʢ���� ��@�o�9�;���,l��r?Y��WF�����se���f�C�i��G�he6W��ւ�����g�m�AO��(���R����Q�p���U+ْ!��ŉ�nN�'9h�i�Ƞ�FS�L�8�?�������nx{c�c�I�QY��������}��ڇ�H����z��<�:fpOmf��� �����_�Fz-W<qx�wg���p���:����T�Tr��q�$%5Y8�è��*it��v2��;�~�4۠.�E(6RtH���I�Q0̯�F��Ф��9� ����r�%+�Lg�T	R�.t��(� �L���.�E�Ka��T�!d�k<n�g|"�B�"J�r>��}���N��X���T?rgibM,���L�B�?\��N�o�3��ъ	�5���4v��I�����fr�����`(����T��������©b[�v|x�X����DMr���
��[�|�{e�G�洱
�-�^�U����ϭ#aT�0���"��F��9���I�1�S���1��B��E�{�5*Υn5�A�w�]oܡ�����Cu9&M��l\��nt���h~.�n���¨��p��,9\'+f_:����C�8����VϿEx*��'_���Y(�4�3�4`�q^T�3xg(d�6��O:�b�|�l�N��b����$N3�I3I9�$8��B�fL��'������+v[� m�ۍ��_�\JЎgHG|���� �\��B�^��x�G�� Jw
k/O�Q1�D8�]�#
G���Te�7�qmSOh_�[O��	�,��j�?Q�OI�؀���B%(��7ٱt������Nڦrv�\h�a���(1���m9��mgX�� �-lK�n_QÔ0'�+�CK��?nqL��gE�J�>yB��&*H8ЀM����	��V�""f�Ґ�E�}_h6i��r�v�2F����g���x���0�����yI�
�O���V}k�"��\�6bx���2hBr��M��|���f�1����/Oװ�V��N�&jS�_�%ɗ�� �����$�X"�H�ִ`1-��%�� �x[e;�Ǐ�cq�u�ɁD�/��֗�%ϖH}����XN*���iE�EE]�y��֗t������W��؆|G��'#�=9*�︜�k�>"�yu���`sD8�7��ׄN!T�X��Μk�yO;&L�H��>qt�fa�Fr�s�+�'��L I�_�V��zf\MXykw'�)��變
`�=����%3�=����λ��ټ:74��Ⲗ�W%�)#ܐ33��t�M�i�l��G� �\b������A|L�Z��O��5e��[ش�_���jM�D���;̳۠�O��6A�^@~�C�C�����|��IB v�CWSV�� �����Ik�� <7?ׁV���Ah^�h��.�
G�3��NC��	b��,����޸dH��R�؜+�k󲼁���uh����C�0�\�c��;�~��q�J��7�T�r�ҕ�'���˨���
���4������Z�)�q��"�qx�60{�2G���^nu����9Co|?y;�#'�!/�Cw���צ�p�~m���Ukeo�1��SL�*�a�uV�C� d�	1�"&�ʧ�p�u���Zԛe�1��� �K�׵\��2s�t�iWf����r ɩL��Q��W�RMN/`����蒴��x���3m����KX,@,R�"[R�d�E@\y ��Qp��
g�e*W#E��U�|� ��9�|b��y�-�'	M)��Tx�<p۰�g�6�Fh���t�I� ʼj��H�{� ���#v9O�m���Db�	>�. S�i��,*�U���|7b�oZ�so���9���ji�����cS��!y/N��3�q�K��I����b��7���_5=��t��d���9D���x�}3y�z5��3�ET�o��e]��n�Ɓ�4��|o��(�􀘩�#�*ћ`X� K�̘f���h
�o.�B�M���ښ)-bm=7i�=���b��B8�@R�02�E���a�-�Ӥ��ل(�4$x�7�?��8ȭ|u�������,v}�K��e��>V3�T���"dC-ʽT_����'î�����Qew%�wzd��g<+��˂�0R�2ҡ�Y?�!.p���N"	����P�}L�ws��S>ji<K�]�s��{ɾiڷvĜ(�M�y Q@"�@?0�����,���|D�=d��+a���0�SżE�?_<y�����,�qs,J�!�h�L`��~�B�q�Ã����5^�&��?���ؙ�̈R��*�!^$�\��Su��������&r znH�,;��Tbv塅8�!�a2o�A���>bAKp����I	��8��c3{�o��K#�f�#d˩�ET=�0����f�ڹB��w�}��Du]x1�%Bșc˞��>#/xi��]!$y�
��7D_t�>Xq�A�C���J{#�V|�0j��K\p`T�撋�㧹���0�n�?�~H-�-f�)W9������Ua��G����ybJX��=ɉ�W�5��pW���$S\8N�8Q��-W\d�����Q.���]�ĄtD�p���e���=��Fi�q[i���;(��ƞknk0�A�Lx��H$�K�ዸ�&�i�ig���j'D�)���N P�jx������h�(nb2*f �PZ����� ���5$��L���]S>Y�MF�HU���d�
�B���~����R��X@D�#�p�� K��N:�gtZrL+��N�Q���Kw���cy-l���U��AXp��`T��8��Q�IZ��2�����R0�徚2�;ݶ�ѨGK�,p�i_�߻F&1��������4�`Ż�r������깞�$/�#�u	KːO�S�a���t/b���)�&�{O����̛�I�mԪ�����EMSF�V����>������&xAc��� �T%�ڎ�0e�Dl������ Y��K�vδ���n����v�"2�:8�˄��<���eN����H��W��N�#����E��k�]�[���1�|��	���X���$���8��������:+�V��zi�Lq�mȟ����cA�ڨR�B3�s`�T)�s��Z��ҧ&v�DX��5TQ@��4`�R�m��$Uw5�/�1���5�Y՘m??nd�AlU�����Q�}%Ix>W9�|~$�%gv�����*xo9m����ɵu�����g�U�tV���+x=/����?�gI��/�]�D��V�����*o*��`��J������'N4��u�d�����4��#7�c�V9�T�BPC�ٌC���.��y��И�����cBH�
�@4��.�>�;�C}�N�qs#��߈�q�B���By�I���7����������:�c�m@9҇%�B~��&���7�8�ڈk����$���������nԛo�����i�te]2]��q-5c�Ǣ
+�n�B���e';!���U����+�"U��9OM��7q3XuQ��25eP����X�>�Yc�xq.BFk}]�>����5d:���ݺ�)���7E̱՝��b أ�kH/��sJE���Ev�EߐoR�	0�|p4 ��bR�sp���V���z��n��7S������s�ql]|l����r������R�������0'��^��Q��#Rb�=(㑸�S��L&1����D��6��8�2�c��3&��Ğh�E�I�����3���?�سJ,�"�t�W��'�ՠ��Vo�����-D-e����((�L�a�Tު[�=|Uu5#g���εJ����pc�����A�IH�]�� �֓�aӌ�[�`҇$R
���?4D�P�ru.n�vi�B��������.2��� }��!@�u��S=P��1=3����;��=���)�h�r��Fr6��ғf�-�f��"�D�*�����pE�~����|�}��k�qDg����-��$�?�q�L}Y+�d6�8���K$bfFąr1�w�j��Rd���c�}��ƹ~�J��2G�+�G�����h�TH��-�S�Ns�&kt�����o6cF��K��d�({��$E�w���R�ȫ=���qe��;n��'n�堦^D���� ^���@7J#�ī/��Q$d?Q��,���6� ��p���U{Vah>�t:�c�N�?O�K��|�I3�z�*�,
��[�|]<��Oo�(�?i�%�$l�H_�Ap��7��l�w��u�
Q8	7ڪ�5�*�U�"&D�X�k�B���g��?���O�		���·@�מ�~{b���
�#
��8��OJh�Y��̛�:M�-�����M"PN[�",9s�C�uB����l�AL�TnQ߲�F�1ߨc��vմ��<;iv��M�-U�T��b��,�����o/$������`�gr�]U��O�Zq������U�(Ʃ�=�����,��:[UY�@�za
磎�H��,�
�IY��qrP���
�zL+��ԬIH���Sr�j�?A]�p(-Q)��՗�6���9C���	�+ޙ�i�H�p�LE�ɬ�;WC{�ϛBԀF����]G��;u^*������.�W-Ԟ�<<IF�J-�%�N���Kd��m��]���:��� B��ǲ�#��O�(�z�܌��JH�����ܟ���ц2I�F*�i��rS霃pD~9ej�/�1D[�����e >c� ���%p򧞕F���'a��\�<��(�$�Q/��<oF��"4E����2�iO
o���`vZZ�M;z9�̛T�dt�0xc�h{Aﳵ�\��l��5�$������tL�3>a�d�o��?��t�ԧ�.5��qZmli�:�2�8".�`�Y#�J�7�s5݆���9a�{���J�4��-╙TZR��������H�7vlڌ�K��Ĺzc�	s_��DS����,�|
)�hm
f���$.���g����Q��SJ���bI�[�ʃX^+@�VN���TW��z��>Q�y&M#.�t��8��.����~ݲ���w'�b��!3FR+&��+A�"DsW7I�	+��qNQ��&v�ӫPp���}fw�}#1i-��G'�����q.4��i�^m��1-��dn;o�xIa���i0��u�Ϭ�t�~2|®جV6`�нQ��G��jԯ��so#����ioƉs�+��)�1�E,σe[a�K���ߛ�I,������Q��'�zU':]�V.s��(͎%\(��E���Ka⿎a���T�9q͚?dw�\��\DR��$N���_n@G�I�P�<ל��oX"������E�B(���*G|y)E����oV���Z쁫Aj�;�ZN�k���{��?���L��孵��/v>���a~� ��w��B��X��::g��|:砟��Ksv��⁇���&�T'i�Mzz��8��E\����#�jTE�A�^��w����(@�_�Q���,
��YPi1����T��i��ɤ��!ܶ��q
$���.��m�5
aCe�
������,-N�.�`���@Ei�_k�_���$���g�촯{9kC2���}�w����H�]MQw��v�:/*�H�-�p=��{�����("e��r�W8���p����M����RA�"��9�_��!(����)[��}޾�w� Qcn�D=���0�kP�=E\Bbh�%}�ķn<�T��X���t��Y���H�SV"�^?���mgPS��t��+���
�`��4��5E �(#Gƈ��B(qS�#�m1�L���)����J�	������g�VPLu���a
���[ׯ��~v�N8v��U΍	~u����R�� j3��p���b���^K�����!Ec���u���]��;�R�_3�� �$��@�L����X�9�@ޝ�`F�$-T�����Z����#3���R�R[G���<ta��wIc���:Z�x6�s�-<-�Y �+�W��"�ǧM2�B��ڜ�2;ضs�2��v����H-�đ@-O�^0�ڿ�y���]?xT�ےƎ��4l�C��XfDe�p�uZ��>5��k�"���;?������a���Eq�d�p+��(�yj~�~�_m� U��H���ħ�V�5o�-��3���v��Q��|�����'��a�_���{,�����372}������0O��d�������=�[�?}O�+���ߊp�:�L���ĩ�T��Ș=�a�uo@E�S�o��*v+4NF�Μ��LZ���>-[�y9b%S���gM-��+)�N!�q�s�u�K-�ZK�*�<�5}MY�5����Zc��`��6���9[{F���ߑ_�^LNX���k�Zx�@q�^%+�ǽD��žy�gd�0X�ÐJ�I�Y��3B���ccK8;G�S�s�:vN_ϸ���C�{V�x�b�Ñ0���
�4	�S0	��Vbr�̈́J�]�7F7���{�@�oN�"�R��LZ��+�^[)y{�^�e�x��,�~�,D���jc_��D؅�0��S]���b���q�ԉ7���Z����og%T��������c����j�+�3���ˊ�S<�N3�D7
����Ά������ �)/�}�d8�
�]A��!��$�Wt�ˁ�0�7�g6bD#��z�}��O�� �a؂��Yǂ�{y��C�W�C��&��nH��^ �C�*y��ޔ=�*���C+6����pf�8ƻc{���,}����ov0u�V8 �7<�������nӺ�Ç3�*����!��X|�����BU�[Km5m�F>�dJ�1��]�{5����Ex:��	�R��W��B�/���W�GN���k���<G�Z7��1�ؚ~5"$U$=v���� ������Tԟ?����7�)�x�^�S�)
C�����f�XAq�Z�������hz.T3�4P�AW��(���c;
8}���^��鹱�cry ��j@���g�%:8ra���  x"�Ӝ�x��D�\t�����p}V���#xLJ�&n1"|g�ǲ�MK霜s#���Υ4�kA-�:��Wt�b��T�M.l4�6%���z���=C�ppj
�Pq��֬�g�U����'4��`��:��p�>�<>�ß���;����8s����'^���}p���.<����/܍?����� _Hނ�Ĕ���.�^[���tJ���#�������ZȨl:1����>��e�@o���%ǭ���u�X��|�_5gV�"s@w'j1e��k�j�VU��A@1��W�hy�v^f�&I��%�6�y�<�=z�!���V�~dVk�Řx�&���@�a�%�����[��ۦI���0��p�>��g:��G�&��(���f��������Ej���L��e���O(�Z�Ud�W��- �A��y��0 8m�Ńg9	^�����ʩ����0�.\w�"��x��$����M��*�����"#Ő}嘣42\�K)bp=p�����9Dq�/g�BsLm�@>V����HÇ��ᶚj�g�w����HIX�s��ಕOiV>�n[����5�/�7F��ItĄ{>��f�x�¸te:a�0W	 �Iۘ7���)1�qSE,�Y4��0^H�&"��߉i���-a�\�p���f6�u�H�<���Ҙc����v��'d
��U~X�k������J���ׄSL�n���m�8�q�#���rߣ�:�����J A�64�H	&�9�C�.��q�U��Q���JC3L�M�c�Gi��+�e�Ϯ+�:#�����i����������P���A�|j�:��tZ�t�����w��G�V��KP��²�"p%Q�I���!�rA��c����g���v)#w�eĎ�I�J��@a��{vR��f���r��v\Yo������x��K|f�G���,�R̛��Q�1����ߛ��x�\iI��W)*�a0�>����G��&���D�������⫁Z֌~6��n�'x�BM2�Xb)_�W�6;��:N>ś��wa�p��tz6ח�-��c�l�95� ���^T�I��N ��Jc�:L�{-݌��kDT�|�ŗ�;�����t��b�s�X�Wu�'����c�������9\�iv就=�"</�o"�Etmtz7*g�Ls��륭ݛe�16FP�G��<���TqP#�}������1V�<�]\+"N��m,�aX&�����
Np��\֒�R�/�ߢ��A�������(WK�:���&��X�~Msq��M�.^���7_g6@ g}��E���'�,z#���saYc;�^k10����Ŕ0۰���Z�b�?
��9��qV���=X2��T�{��	�^b�G�$�ZY�[�?c���	O��F��c(��^Y���g1