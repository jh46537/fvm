��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���9�{RԱ[ж�8�����������/a��:��#Շrb�,��Y�)n��M��Ӡ�5H�������w�� �Gx� �Vg~�r�5�t���5�Ш>@�t���57�s�f}U�������2'�k�l�E�g�ܒL�������(B`#�%��ǩ��b�y�ّ��o�ka�0��4�~u���͸c"�x���3_�XlB���J\f��E�W����	�]��8� HI{�s�zq ���s,=�G�:F�V����Y�e>�V4e�i��_�F`�mg�_}j��&���\���B�꼗5�%_����^��Q��q�o
|�zyFB	�9{i������ag�rʲ5Fe��Eó?T6��}��K����JN>Cgc��Ӛ�cH�`��(B�� �l��j�*���gjdų���\fٙG�%���$�����tXS)�N�����f�td���kt��*ؽ3��t�����-w��^XY���L��K@�Y<&��F���F7=��g���=�p41�z�Y~��%dh~��5���$/_,���\d���b�J�Jc�i)vs�L��]�U�Z4~,��7E,�~�<�bЄ��
c�B�(/��kЇ�6+���?'��X-%��,*Cd\�H�QJw��Y��)�>d*5Jy/�����֌��%�G(�^`��R0hL�U����v�A�k�3uNh��V�3SIK9�X2D+�����ٟ�`3ѝ�6&�
*��G�ӗBLc ��0n���m�:Ҵ|�Srv��?�Ь��P�[-�?��MW>!Oq�#���gXݤ����k#[.+A)�Y�+�� �tt����8ϻ<�i$�T�(a�Z�i	���9N��@�\~��aP�wQ�Wr�BW��V4a�s| �]28[A�%�������Ju�V�ɸ-�`�,��ɐYc3	��� 7Nȋ}ۭX��5����GܼgN�d k���:A�F3����g�qδ���
�QT�;J掓��Ͽ���Sw.L1����b��}��߇��wzq0�N� ��7����h��a��!�6nO����lW��RSz���7�M�+����
 Qh�?]]1�t�`P]��f
��:F�݋�c�8n�jt��,N^�D�`�o�*E�P }A�l�@�+A;
�[{��� �5!��?�ľ\9�X�D��Yny�Qw�=��q���a��LᯬQ�F���N�@`|�GG`_Ɩ1M8>��<��Q1��}v��]ӛ�i�=����0s2�l���gE���X#��^�ԕ�!SK��z��)վ� 3�����T���a��gK���C ����?���X:\�z'�e�5��[��r���p��������h�έ�>E#dH�9SO�'9T��v2�M��58�:4��2�����0�����c���*Y�ǎ��fJ<����3�FO�<�?��*�* T���<���rP�DR�N�Z�@�Hx�J�X��Yn���_��X��|�Ȗw��j�������I��Y�Y�|�0c��s�?� F�J�Z����j�[�U����������e
��D�i:9�~-P�~6�ޭs�W��c��J�]�� i#�YJ͜,���.�z��F�)��)�3٣��m�'�v�K����
�>�Zr>�/<��ѻ���vU�dGPgB���P�]*�o�Ǜ�c`�3�eb_��\'C��đ�y�5b�ȯ��i���jY����_�[m�R����;�NN�1��3{������JvC�ƀ6��Q �����b;����-���4�������pf�k�����+)�*��ķc��$�H��/�+��u��݆0Q��"�p,s<�
EF�b���[�G�p�]��{Op���#u����F�4�c щ�lG�I�F�s�pQޖ2u�X�&�/�V�:�C:����q���t�B��=�'��z�: ������)���Âđ����A��������URz7*0R�_~��Ώ"������V^����`�Y�������۩A�W��ׯ>������@X��oX'�R�%|d�)Z��tU���S��Z�����)��P}j�j�qRn�hK�BW�1$:�Bx�W��A��]�ܸ�y�E�0	%��ĩ!:�Ƶ5���<v<�,$YT�֛9nA��@q���ߤ10rĄ!z��������F:�:�Z�wFlY���k��k ,-��_��Z�Gm^��ݹ%��%�ۅ[�F_`��a��?���0~Ƶ��ڿ���w��a�=��}��,�}���*�D� s-bx�B�y�G���Q!0��K����-����7��	|ڶ��Ly$����UB!���1>��:�q��� ��uT�^�p>\O�(K�1M& j�&S��4�q����5�X�L�V�v�ÉE����u D���Q&�d�E#���_��-r{���b'�T3XY����64�i�+V��`�,k~�es,}��#�^��v,�	{9U� �oN bd�X]x�c*�Ô�o�<���p<�w̔��*
7׆�-�BA)�W���i�!����q��o�B]dza�v�v�fU�2#% ����8����4��<ۧ����q�P�S���'�s�\�-ͣ<`L��5Uz*T�8�%��٘����`w6�%��g{��ks$?0~������/Gu�99�?än��P��n��6��1ן+}�%h����� u���#9]�Vf�,�љ�ʡ2���`wbfj	'j?_��a�l@		��_�K��.a^��w�
�q������mr:ޤ�A!4WO�8 A~s9B�-*W�κ����vT���E�̜tm�c�a�ⳳ��J�"�~�A�ɭN���V�ˣ��چ��9��o���ѿ�`ʃz�x�HITvA���	�IȖ�����O����4x�k��:ZU0iɧ��1 �]M��dp�t���`zN���Q�u�.�=r�Wwg�9���15���-�V��ڎ��b�E����:�v]a�P�R����1�<����ZKǚ6n��v�]M�.�q��uF�����F�:.���)Gb/)�M�sXbM <6m��M��_ӕ�դ��I���bp������c���T�K+9�|y[������Ÿ$.S=r$�k�Z>VP��v�|E�W��ȷ�q⩙wX
	��!1p]/�kV%�����"o%˹B��z�,-�O�}��ѥ������(��i�0{��8�$�B�r�����؁6`(�)�|�����EοqQg��Mwƭ�~.�X��ߥB��$���J�tg=w�'����>��̏���C`���Q�2�v�P���3j�&��;�'I�\�os��(��8�<�������`L����Ɂ�8�n�?����5[1K�Y�:���>\>�z�ܖ5W��"��˶~=��!(��+��t]��'W�Ed�T�÷|
��@�$I!YH�27�aYo��F�*��=-�@��?X�,�`��U�������ӒT=�Qu��H�g	v+��+���	�`S��5y
�
?�\W�'L	���c�ډ^ڲ�W���M��Qf�K���ͣR L�w�aE��uyO�` ��#�cDE�fC!�9�8~ǩ���3��`1�D�}���i�K
�첗�+Vܙ������y�+����k��=M0����� sy�X)m�&;(E�������k]�������i��+�n灅0��D�*�K�%��ҧJ�]�\�T�)o�cIvAX�͢30[/29���n���H�OW��[,���cgY럹J�cd�=i�*SX�u2O��a��S�O=�wT?�ie�8���Z(�))�+�Z��&�;�!o�Ym�fM�x	�CK��e��G��x�B$N�	�	��w/�H��	s��P�~k����=�N�7e�O��*<(ҷu6�d"�T0��]Эjݨ�v��s=nu��(*�a�I�/-݆\ā���l�?s���f�ב��ӏG��ש��Mϣ���0X�	F�τ<�mM�3�;����Sw��3㹝�?���������l��P��;٤h1�3�v=2߃+c'ͻ؍l�MjԠ��2�4<J��X��Lq�����l��������� �?�M��4*���W��6ڨtXc)����n�se\t���{޿o4����7-I��*PAz#���a�����Ht��T��Tŧ?��B������V�2Y�Z���I�yo���.��3�_j��a%жr�,*�|�)��~��(1Fs<��e�@��?�����H�*ې�Ik*1����� ��p#UI��4k��|Ɖ���!"�퐏�od�剈��KUmE9j&b���%��`����ϚM��u�ЖU��-�0�4Z�HU���𤃷�?���+I���*��M۴�2,o{�L��i�z! V�k�L�]������M�l�+��%�X�t~h��\
O�W:�-y�1$=u	i�c��K��!D�����bm}W�I�O�Q��;k��"ՐԂ`;�4�������k�B����O��h�v �(��x�W�Vi,~��ĳ�V��6U�N+Pm��q̌wsɳ�����s�*s�D�č$_��7����b�ft����d?O�[E1��e�\�Z#9�:�M&Hhe�AG�8KNm�Z����^��by��e��*�A\y�x��%|�z,��
+����a�ߒ��ak�,"�i@�(�}�[����̷]l�r�\U�\ʐ�NiM6�k#�ż�������]��ň��x$<�-��w�WU�����+N|�_F�p3Y>��%�������Lx�}%0�0�_�́�J˴܍�]x?��z� ;�Y���W�7���h�,��p���>D2�g��r�Bmv�����&��P��Xx^��&�,�	�H��
@����U\�qdL��a���1�srn��A-S)	ph�HP�����K�CL�zx�����.�و)0�ǉl���ߟ�I,�XicoT-�F�T�� c���f &C�����8z��[��D7��b �D�f>���3J���;./�<N��ǪH
c[d��)�Iuӓp�|X��p��+��𚤀��ɿ�L4L"����n[�}�$���,nj�tɯ0Z�vI/�c��<�~��v��X#[ڒrU�m����!�T7'��l5ID��n)�-���S����ׯ��C^���$�8�7a`Ze��Q՞}ծ ��"����r_O<e�¸��<)��:��E��2�Kή�,{90ۅ�� @«�392�0[JS� 5Be~z{n�Ԗ����� ꈲ�,�$��_�A�,��]&T�-x3���!��Ɖ=	Mcr��l2@Kw9]��o|H�g�3��,�m3��$x`f���5uhu:��#�ZfC�|�g'?{6g��BȯK!˪�n��9R��^�/�;r?�
���,}կ��ŪϾ=*1��@�΂[R%�3������ ��2��lY)}.�NAGhL���������%2'�h� �d:� �\��P�#�K��|��O�%8��Id�� پ���/t�q��p�= �f���B^�9�C��x�˲f�^f�1(K�!"U���J�U���a��4h!k�f�|=ƾQ��i=Ƭ��Y����W����l�dr��r	x�o�Z��N�����`1b��n۸��غ�!��zO5�"��`J|��I��Qip�HpC��ʺ\Rcǅ�OO��3S�)�=1��6q�nx+�����ީB��m�K�w�bJ�B?���B�����y�L��;c�׬M��Jf���lN�S^H�5i��9����(ap"�9]ff��)�( Qڷ����S[���|E/��bf�2�|J�؝p;��أ��yt�M���EG��3ߟ��ݘ�����~�U�������?���"V�p��S�
�sAOP�en�sR��	'�$N Q��=D�l�����ą0H��p�MǾ��s@T�Jl�ps�����>v~B�ò�~�c��ٰ�2#8�DI�.�6�B
�L�mg����/�(�+tܭ��������0f���<?��@i1���X�S��|����a�ß&���W�s�q�Bd�� ��	ųR�[+C��]*3T'�X_��}�P��jK�[ʥD&��h>F��/�ffK�|����!���s➕vF���;I��BoX �d���zE�敔O�`��P�,��1��U�Ä�}pu����$@���E�zX9�+O�{�J���2u�ou���|� N���O�<n�6�[ɂ�5;�:%b�}K���,�����F]k-�)�	Q��n�����Gv u�8�	�	]��@}�PJ�&���J*��)�����2c�&� ��컶$�pς��i�Wۿ�%�1*RM�_ϳs#��3:�����<_i@烡��1Á%���0�<t܅9�ْ�6�BiE'o��/c���P����c���Ķ14���E�n������|Կ��({��(�}2�'�&�ʥ����"^�K^�����Ż~@�F���wꉎR�ןZ'���q�����Ҵ"�i#k�o�X`�RW��24� �f%�F�vtpF��5h*���S�4X���"�UX�3+ �R��va1�����^��;r��Jlm��߱E�ؑ�Z�kvVDA	�l�L_�\�� ro�[w�AQ�5]d�_��E���k�($M��BSi6A�o)2 o��B�
��s�������\0Jý�U�<�����&k��:��m�ٗ ��ԛ�*�B}�d2XR��K,ݚ�(~Q���P��y��������z;j�m"�z�͡�=A�>A����E1,�8n'�ye��cÁ�{a�� �A*������ſ�Km���X1 �y�IL��}�l���f_�(b�kS[�˘��m�������Y���K�$#q��Ua����|u//����Xq�Po���+��CP[`zZ�+pp��M7�$*Q�¡�ھD֖���W�2G�