��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""���᤬����[���%r�H��Nx����,��l�#��"p�(a�\�����}�t��R�c��Ya�^��ӑ[�L�
�VF
����&�Z����Swd-�Wb�4�+q�Ġ㽃�tȘ�C�<拣��	����s?屺a^���1V�zg�ws�l����ᆶ�����J���һU���m�f�"~j�S�F���xW|6�x�"6*��ĥdm�h�l�����Ic�O�C���{�<͍��D������/=��Tz��n��rp��L����l���D�)Edm�/�7�Kߎ��ux0x�ڬ��������g걏R�3���n>��w$L�хP���\Q� L�
�2g=3/������F��гW���U! Fᣘ�@����4������C4�>�m�/�q�QD!p�IlZ��/�Mħ��Ih�1�
&�0S	[݅���d���F�d�wVÁ0��<Ĥ/b1���Y�c���8v\ϻ����[�gWd?e�^τגk��b�Ds�T i��� V��������m�s�`DV_���g��	;��� CΨo�����.k�H��&g|���x�J�S>@J�&dO����ӡ�m�5���(�^9ɭE�(�sݚz��r���a�^N~���-��O\�<�X�3��.�H_��L�<P�J��>+�(��p�2�j��-o�sp{��S�mř@�S;_�1(�\�.+=��F�F�r>�恊%� 9>(e�9����v��ݰ.=	K"�k/ �*;P޿�Q`�xH1�f�P^԰��R�)������yW綉ԣ�:�G��қ�C1�Ƥ�����=�Н�ȽG�E"����U�u����������mbV,X����3���Ho�Y$@.���b|�I,KP�˫�����[4���_?� �]������S�}�
��-�wOʂ=�5�1�-�����#��{h0�|ټ�y��L$�<X��2Zy�;���fT����2Ϲo9p���C"om�[�s�g�)��s�QI`�H(�{�0!l�tN��!�𗆒P�W�5��;'B���a<�$)�kj�1o�xz�^~�o�nz�:J�mh݂ۛL=��ĝPZW���x�p�w{��_H�1�dYt�bl������z�R���m���Ь c�:�;;I�G�`	���ð����ak� �+�HMı\ ۋ��g�����i���yߥܗ�xeQ��z�fRP0+?�<�v�t�S��%:��g����B�¢�*f�,��%+��(���EZ���0Q+��Tr��e���!�L�uDH�v?c�l�c��A�w�m��.���̕$�>NϥS�8�/�*�}��ǝ��Iq�ً��O	�I�K�<+[�����崕׀�7��7e��u>e�N���suu�,�D��)�O�Wl$�J�Vw�oSc�$5+��d�MX�FMC8Ҷ)��Kw�]l��M�ĺe����g�E��+m(�6��W5!�B4�ʹ�x��y�\�P�<T�B�@HT��-���������`�=֊��Փ��)&J�U���B�.���(�Ɋ��7��4W�1�j�����LB��o�%_�O['WxZm.��''��FpM|Y�v8r/��B�foLh��5o�{�� ��{x���0���e8����>���d�.���#"�z��U~��D6(��7x��G{�7W��x�[FAd���ܠq5��=�i?�D�U+� ��?h��"��U�j[$���[���
�lCF'{wy(�w����޾�
Qc'���)��y�B�t�����	&r�I�~�ŢQ��>Z\1��K�?6Z��l7�o�%�{t3ؖ��=a|i��Yq��x[P`y�cS��Z����]Gh�ڌ��^�wM[UKf�����S�ؤp�Q;�a��V$1� �]��h׆��,4Mb��A�vFWh*�~��0��7��}<��#{��縈x�j$��f��%C���L=�	���TZ���)��n�I:`>�k�3�?�)Z�Vۺ�;Q��3�����b�:c8p�b��)�4��f�m�\D�:��>K�y�->���f�!;�=ә��w!Ml���H멉g[V�8>M�!�w���G�i'7f�?��Ԟ�$RBz��� �,�m��釗�"x�-�� ��h/	�<@Rt��Hǆ[&% ��=Asr6�!�O�5u4��_��j+���z(��$K�����|�N��F՟� w�tVčW@Z�B��sk� ����'��rJ���|�'v�rLB�y��5���5:�DG�u��-A����ˆL�u�*0�!����1�3��{/n���3�	�U�k�D_x�Ֆ,����߸�J/�x��� �3���\^=���UӰ���Pf(>�}g:������j�+A�N�KNħ�Z-��ʩFjn�ў	E��f[�������rXc��ڷ7��럵z�����7�'��t,k>M�	�I��վ5���C�,㽹 Җ:S4��#`� Oƈ�VSb��8��>�x&5)5$��Ŧ��uU���zt�HJH�Ya�~gʠ�����G���fmq��k�DS�:`�t�W�S�|�.�U������L�����<0t���
>����9��R5=!���8o�"�/��~�J�"S��.f)�m|ٱ�=��Ŗ�����b���E'�Tg�!��th�~��+�{5�]B>��N�ޒ"�W��<.���}*��͘1?�e_���vX� �.x�y�P��QS"�+^z�\�`���-���ڈ�Ca���E�2��2�zRKey�?����R9�d"R/�E�)�� �]�/�nb"A�̊��)q��x=3��GsO�'G���r.Q8��~�UK$+��4�y{�fn3wB�cd��
A[���9��G��p��C���a��UTu�70;���(_X�<zĄ�3��%G�����/:����� ��&�u��_6e������QLZ����E.3t�q��gy&��C2�������mU����iH5ދR;L 
��6)�/4e�"��j3�	��6�)P �%F�!���
 c˾��B��;����cT9=;�q)d�j�ǫ�d9v�<K����]4[�.7��p�)���J��v�Qj7n�����-�D[.fƔ��z�7�t�<e!�-��I}5��6�ڰʈ����z��l���n�)�rN�$��F�A%c��HJ��u$�*O�L6�x)|!߳�D��~S�F��[�I��Q_����e�(��єkZ#TG�U�2����@A�ӕ�07_ٜ���̂4	~��;K��s�,YnA�(�s�4����2U�ȱ�I�O��P�#!H���y<�wJ�j|k���6ٞ���s����k^�%���jґp�9�s���&�kh+���`NM?��N�\�w�jyRAhi% ti�\yX������c;�_=��~\*YU�6����J��O�-���V2�Uh/z«�8;�W9Kh�o�B<�<�����lvk��4�	�$-��,�j��,	�/������Z�z��+ {��)@x	5�k��a�H��5LR�X8!?ѷ&�*S\�nA�#��@�1ŝ�"^���]Z�G���NXWkΉ��[r-=��6����v��{��Pg����4��;��]�o@�%�wu���<��h9��K1m��pĮh��	�6�x�{�o�凡��h�R/�$ts�;?	���zI��2uX�uǡ�/����s�a�i�a*�t}5���ep�tי�-�C���]�Ba�n���]�'%%��TY���V۵�RSS��� R�l$�I3aV�F��΅!�.F���P��,4(��x��b"�����L���JeJ+����'�t|8~�D�������G����i�"{��{{���(c��M�$�F���u������K�;��MХDQ_">�����yKB�\e:�Q���;b�#�Ҝd�C|��I'��s��'>Fƥ~��-Ce����'V���Qv���ɤs��~��9��#Sd4ј��2�s����\�!� R�	�k�w&aMv$�
tm*��y1W�	֊i��Kvj�\8ъ��{<�a���![���B�S��dغ���,6ds�� �^WW��ʨ���
�i��dA�ӧ�|�X�И��kD��迸,��a���v�0�=�zZ��;l'-�d���?��>��8��#a�=����a�g�J"�H�+����I�쇡�{��PkX�ޥ��<3�hJ��� �4���ޯ���u"��~��t�HNJ���1�e Fz++Al!�G0U�P��l^�2��DK�'�e[j����w)�{�1��-�)��$�����]���cv�#$�DA`�H����S�S��Jw�)��V���`�N��_�O�rJ�EF�j�u��<�e����ޕUawг�� sP�+����"���y_�
�����:�n� �v�{�>5�JP`q��O�o�<CO~� ����M��(;j��,wd�h
|3<2"�E�
ݶBo!��@��RQ���I.px����\�Cn9��]��?� �Ee=��N-���hu
��;&Vߐ�Vs��}ܲ=N�#��������s���^�'�S��g��N8zW>��~WDy���_�"�#J����9�:�E��`�|��ҵ���(�_\��rd4լ��S��՟ A��{�+��ę�3�f;k^���?G�]̪2���l�ZYRX�fC�+���}}r@}�>d��6�L�s��9���0�԰6�w�Pt1�Ħq݌�w��8�|���(ޯ#!$㚽�o���ԯ���T@B;?aiH����!�5��W�ךfٙ ��Q��HF撘�wQ|��A����~-�Q>����P	�MlpY@�a�X�G��T/�B�y:2+���
Ԇ?�u*�wҘ�gv�Vs����I���p���i+�� ˼�-�^� �������/��CSv{"��M=^��*���i¤3�/��GZUs
^.�l���NX����@r*>LXh�8����4D����ع��J)>�A� �ykՒ�Z�W��;(�`�*+���C��BC�����3k�ߓ��Ki��p����ɩ(���3G�l���Z��g� T���FB��3 ӯn<)���yd���)9e�^n�I��{>����@$Xf��vzLV9̟��e����^��U���8\һ�=�xf�5��׃q��ًuBw��*��m�8������>���t5ۣ�8�E!I\�B�j?;
"x����GN��O|Z��5N8I�g��"&�og����ԝ3Ҁ��CJ{�\����#�_���<�p|P!�Y�b�'rj��l��-��9���f�r,�o�Fz�#��G���9 ��K(��N�s��8�ΓC)��s(w��V�	�s�T�UUL�`Vt�6*n�6H:������'?>:
��m.�X1X��)��X��o�%G�Wq���Kȏ����pُS/@%�G���b�P:("}�\E��%�?�����2 n�=�,Ŕ2+�;�a>��Gx����ĵ�>䤛�b�rL��Wj�pf<m��^�{^meX�X�p+���S�^���0� POa]8����2Gt(�Z�s�Z��J�eT,��^�;$�⯫d,#�V�W����R�� |���*����CE����F.�qq�_G(}r,��k����0�o]����w-����	�8uFh^�@#��A1����EPN��^�Ҽ9{�Pj)�=��e�.vZ�
�ĈSr�Ymv��`Q%�/ d��?j]�}	`1�.��.�w�r��Q*T�}���/=��2=j��a�����Q�ǖ)�n�9mF�l
�{�m��@%h�)�T�Vhx*���-9�%�����2a~�9������T�:ۑh�Z�G_{��Zֈ����zA�H'{�s�1�b�w�xB��Ox�y3���i/0k$�_�s����V�p�{+"JEo~�Y�S%r�L�^��0}�������ǡ�ϋ-(I�6.ex���n|��'�$7*/�R��b�z*���=D�{����D�O�O��CjId����Iw8^����q#Xt��w�0���?TFY�����U�I��b��%�����o������w���w_+tm��/��{�A���X��*]�9p��v��QVĉ8���}@^iU��,-�f����\x�a�^��`�4�%������С��p%�j�������;�e����,B��9�S�֡{���
�{���1Js�5b���L�1�>�KI����p88�/4T��g��e���Xk�3ʧf��6FU�=G�cH�V��o�=���׬6��C{�bӏ�V6�u<����E7+{��[5A�C�w�s��]s㨗%�`\Lt�7_.�=P����V������e�_Pڳ�sPqY�k�3�V�f?�����X�3tO���y3BG�~VI�D�;�P�';S�񭪗�/ԇ縤�l�3�*��8_���}��o��Ţ���kAބw�3��:��)'+߬�|�MaT���^7�s�p)�@�I���nV�N�ʰ+L�����A�k�&Os\�F�b���4��&;���#�����'~�,9��_h�h�]���g���I��怽O�4�� ���t*�7G�)ed�y8Y��n�PB�Ʌn�q��ec0��B�B��r"�֡�lB���i���p{0r�"��rܡ�1*���
Ed~�i��!���-�B���F(
��#�Q%�[%��ؼ74fP�>�V��Yb����Kx��޼��1&Zo�H^]co#^�t�]"����l�%�b f%�|�1[Ϸԋe��Z�Ki��>�g�D;>Uz�em|P�k�M�˱{PF�#��۾�/�	H��n������(o�T_����W�X]���^�)P��I�=��;+�z�{��g�s�ġ���fG�-%�pl�-%�#d�>�y|zSa�'��N��[�q�5���^mmw(E�'��"'�":�l�\�cb_DŨ�.K����>2.{���5�m���+�ƹ�otұT����Ǽg������8��,ʇ�mը��wr��\���(:�x�����螃�GiDІ!KPl���uk��l���0��)�R�`��u�=ʒb~����zV�ߥD?e��?I�(lN�;�H]�]qz݅�V﬙Is�{C��|$�Y��T�9�C�/���e�Z9�d��J��8�D�d]4���T{L��rް�5�c�&;�r�Ô7?�� ��'����k�6�9���v��V�4�<_��@=;�0�M>�A�t�Qb�n���S��`����>yy����O��3�G�L�0�'`�:~��shu,t�f?̜��у����ؼ��&g_��:n��.}�c�FxGP)x����?��T9f��֞����j�>S�.�o��ftTc��I�Z,E��[kv�vjJV��C�p��"U9	����Q>�4��?�ڽ�����q��F��g����yԮ�CÈv�ۤu���I���Ր�����v� Ґ21Rz�P)nl<���l�6k8��L��k��ɩy?J����*��Oq�~`���]����3�sq0�4D*S���M?�5e����cĂ�t�$������Y��X'<iw0������"~ɧ��˟�.폧�8m煊C�����op��u́�YŇ� ���D�T����nK��%����@���r�p�jG]��r	Tيt���Y�T��,M����z�%�P�[��PF�w����t]N�A�{Bp��������Dυ�,3�������'f9T�X�:ģa���P�q�tV�&��x�P1�X��N����7��D+���ru��w�ٗ
�8��V!���"��!Y��MQ�l��J`TR��-�&�%���/#��2���￉�-���ҾQ�!JC.�!IL$�HO��X�r�����"��Ԫj$��3��e�"鳵����i��Pus�)0e0�j�2s7,7��Ve���KC
���#��j�F������y ~�̜�F�ٰ�~�eVǼ>����s�Z�c��\f�/��KUܞ#v�v��%CY
�7,�c��.��*�ݭN��XK�Cܘ ;��5��0��rDӿo>[˳���\6�X�`!�#N:s�m�����3��5÷�H�r���r��!��n�ڰz-�7U����r�I�^?�����L���wM���N�.�Ŭk��e��C��^q0�����u�z�g�'y�U)Y{�J�+az��>s�7��^��j��L0 45�O��i���P��A�V3;��%��-����YxǄ]:5�p�.q���#����̒��$�-��7'���o"s�=n\@=��Q��[���£xc�֤�����LJ�b���Tܵ(�OCݳ���k[�������t���ޒi_]�|�en��粆��n�̎�OYv)�I�@O�S:B�m�+����H���G2�:����j�G�����>2�f�g0L�h���b��]Ĥ��R ��#xTr.ZC|�V��c9�����'"��'���<��<)	eo\��j��ȧ�������L��ɟG]=��#��t�9�&�m��(����GZ�S�d�������]=5��>���a"&��f-�;:�lb�Ց{ޙ����\o�	2O��&��ZTۨ�ݣ)�Z�H�}�G#		��X:��U�4t��.������6d���z�3���K>V��Kސl9�tQ��Yv�]Q8�R��8s��	u>w�i������/v�b;1Th݅"����<������vh�GH��Z����cKߢ����2���c���-�k.�	2��W�-!�3��[\��x�H�hcFg��Nau_֧la��9���n[`��,��mk5����Y��֝�ş���Le� f������վ+ O����l�!�
{c+^"?s-��K�M#�4\=��Z�SΜ�%Y51��x��	�P'�V��.�a}����4����oB����c�QaG^lF���A���H���T,�^A).r��G :Ҡ�����C+83� ގ-@F��\zףD�D�ȋ����#l�1g�������a"�'��Km���+�^����N�$����2�0��ocr�l0�v��( X-�����r�8Dl�C������@�+���a	EY�}(�'���R�i�0��3��]<+o�������LQlk"��'|��w�� �%�6�P8����yб�n=G�,���?_���ν��JZa��'<GW�5]��%6���%�kF�u\.d��ȭ?�XZ�K��)��6=�D��3���Qj�, ۞yT5ݺw��w�Ro)[�e����O�)db{�i�_���C�({�
M��Ѷ�I��!C�,���T%����G��)�En��-�h�t6�*���f��y�%���d0)���Km+����ů���"�(2��3�g� �C���V�ytFiݒHh��Z�K+����!<��F@12[����y����!U�3�����?��2�E*�����-r�S��0��)y\�8_k4sL�ҏD�'I��j�AR)kR����H]~�����yJ��1M�2-�w���豁�vg�0N.���헷��_U�|J��H~�k�;]��JE�~�(r8nV�	��2���~�-��շ&D��T��7��!�F��*�dhW��Lz,3��-��D���M�D��OnZ�	�g�ˬ���h%R�U��O[t�����]F��)�~T�<*�7;U��V

�&�7K��t�Py�ɉ�IP>T+��z����h����%9�jT�����E]���0h���l��pb �":{��D.��a��R��u�
PB���N��CM�������6����,bB�Dt�Ć�O�ʜUE�q3�����&����D��N��OU�<Z�j��m��hP=���'��x}�ԾȾK@�lzXڧVO*��3h�ↆ����Ӟiu~B����3�:8�Pâ�h�	�i1�uN���X�iN�����/=��D�����J����9�m�T�}�F}�D��S����il73�&+K��K����Lg�|��c,!Z��=��Cc6��l���u*�@�NE� C�?�1��D�'O�gR_�ė�v�9��?{��X���d|��"qn�R��e������Q(��d)zF.�Z��
$�W;ʰ�J�<$2���怷H�̖�t��Y4�օ�a��|7ߘ��P��YHN�6����3�q���������~K���������N'�m�w�t�m�|$ɼ2]�*l