��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0�����(�_?V~��
�r�-����)�b�?Hj�N�9=ḵ�����~x�#�5{��a� ���L��y�-T ��G�+���n{g��v���nk�W1��.�%��:��W\�]("9aЋ3	�.�~��9����i����TkG�pa��~Կǈ��
��Ҍ�{������I�OylCA�@!~?�z9��|���_� L�Ku���9�M��I~��;�"+#.���#�^�A;y�,�\�0!s��WsT��ߕ��r��b��a���'�ϕ�&�u8N�@P��P�p,�e]��.�*�3/�"ޤ�*�u���7>I:}�T�zɟwJj���1k2��vҲMW�s�ٱ�;O�u��zuށ�ZAEi�`q�ӛ�5�4R�+@h�\1B���ŧ�$���[����o`���N+���Ս�K�-�����_L)��O>ؤ����J�U����?��j��Ɍ�o���(!u(63/`�S���������o��v�~�n:MJ���;����_J�@h���I!`�W\�=�v�q}���e��h ��MG�:-O�KwZR�� ��{p�A�\�W�t�x.D8���R5{D��\�j8�N/������˷mY#��L�mQ~&�h=IT>�/c����N��b!U�:w���4tv��7qypZI{Ajd��w�މ��̡�`�Y���u[�]�qi@	z��EȒq�A�J��3C�[�ly����H�;}��}��+�:W�KCmc� B%c��� �����w5|�����u�YO�,��zҘa��QM[�F+pq��:e�E�ӳ�{r��)�{j���ُ��W<���y?_ѣ� �Xi�B�k���T�M�WTU|���u�*���M>�%��I�'fab�7��L(}B��8�vp�7m����r�k��QznGM���ބjA٫)��/���1ۼ�����_�b&j���H�+
6�wQ�k�qG�O7�4�*��=d9�՚�P�DE�
S���Nd$�ΥF�D���e,��5<1��6�%�0�Ǣ?X�	4���v]a(R?q���z�:H
��_����?�g�AҞ�v�s�t5M��BT3�[�A�<��p+�
bM=�pj�?�i�f��pJ�q��hѼ�0G3�4n�l�N��kF�z0��{F˺���V[�g[-��2S=�)�j���g�Y��[�(�wr�#0�B �!@+����QS�G/j�������zGՇ���鲌���CO�]w-s7��-{:��e�[91������Y���$?�u5WQ�b�Z��w�^/�W����L�,�����S]_s�������\@�S܉A${9.�/�$�Ϊp�O���|.��3ppw�hԞ��o!�\%)=���Z�l:���{��_�Ӫ���t8��Ap��.&e^����f�U��1i�I�O.��ܝ��~�ϐ^(�~
fK���u+8���$�X�?k�����iX��FP�$�c<�r�N>6x3���S��N�����u�M&�*�w�j}�Q^࣪�z�2X������o-�pv���/hu��v�d��|Q5�g�y	>��.^�cG[��~ѕ�[���W��x@�
���}jAc)
�Z�F��v��E�~-�5���\�ާȫ�r�|TYCM��, �[��<{�Q���_ z�.�2���#��&����pb���X�G8��1w�b�/ Z}����~K@��H'�)�t��>��o��R��._>C�Ĵ�&"[��gh�۾�M�?diڄǫ�0�tH��Ry��*�������I< ���-3�2��d��mI�L�O�G�zm\�J�D�?(�E��i����<�r���y��yH�xė�0��4��8���G<A�Z�P�fu��/���q��Σ�$�
�T�j���̣��&<��	� �ɩ$��J�4�r����7�0lNV!J�wو|M��٥	�5�W�8�RI_�,e�B�Qur���j틢�dIE�)���ϴ�=�讛�&��'�7)����|俬��hmŜ9�;��;��a��M��\���ԃ�F[��;Yg�G��z��/t�x��N��)�V���rq�I�^C0����t��P�L���{�oF[�:.�EM.�sxXG����ߊ(��%"r$LH����`y