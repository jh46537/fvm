// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nVCffoJy/5frwuzI1yqiQ7Cg0i1bTO26+d4iSpMv9xloORGwUBwzsGhKUwc0/eVe
A+eyeHEwEKOidnAxAOhIDg0Veyg+lZwm+G3/FzJjorKvx1A8zeA4t5DMVpbcBk+L
Seu4IIFaFy1pR1C+07qeZloi2ojy13eX8cru4r1CCIQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25424)
gbxbgFWvvu4knEmc8mPVITJAjn+8sHhbT05QVmDALwpFMLpNY1TJACmc1vocopxv
usSiETbPDaXJNocahM0PcvX43dkvEGBHtst/Dm3SJ+J6QUmKn+oe8rI+c4cSwtAp
9KPBJjT+mNLeW4oX1TfXQ0JI9h22ESeM4Ov0+lODF1TgOd8rKyaEo4jsU4r7LQRW
kJ29Hnot73Z8F/QfN8+wGaAFFFnm3sjPK6YbYFX8O5OOIv0ItVQJJ8YS6JWra45n
bj5QRd8fm884ChucwdZLVxu9lDFcTdAgdIbXZSoWIGh6ZkLmX9FjUdfRuspmJd76
Rjbm/88Rr3SQ2l6OdHJXwQ1vHQeySAu+GOObf8kx52ImFBLKNylmpuqSuQgJ73BE
9cpq76zVfihBhOOyoeULpxbcaWlFrHuLcn5Hvo6LIc56xZxKlIWDAjxfB7XtLsN8
8S/YGkawown7/Z5EmtkIW+NUFXj4j6yJ24Hu2qbXB85xUndCzVBpJkeVQbs1drXv
10s4F0br9iJvVK2PxJVUtcP9JL6ArKQKtisqZ0dzOK0itcse/7GGyz4IQ3MhAWpi
aHerFmFVuhkl5i9XPQLTTB3oEaS1GwciYh1nHZ0Nf81TkfSpRir5BoPsOkj4SAWj
qqHa4jNRisr8BWVJ14DYWd7abYYQlb8ROU3ZsgESWwqqrNdA0txBXK07MqYmNOwG
82tOCspPQdDd1KUtLLGfGMAedXeOUVlXKzDfKg9fXyqhkOMEbGWddZ8IJcsZt05n
5G0aZiUi6gzDQWxj9VUZVMRtPcgeOfPV66HcEe0rk7JfP2NAmtR5P08oO2JwYWvz
Ytb5JUxLLyWGwb23Rv36sLtntiEhrVwo0hhuE5XfTo5HhXovA5gVXq4UN7Y74Tu2
6BNlcOEjmABr8XkXk1te4grySmHJ88SGGgzC/RR5Wn+6EHiBIGg6Bp5C0HOJPkDh
RbMd2cIXfIO8JZ/eWb5UfJEMjt9xBeUhQNf0tOAFwXGX+uu8XXauhSCBPMQN8Wsz
HUyHRQV5gIUuCavWZKqySSooUvShrgh4bj+To0XWfXcH3kyYJ8Td+DZKdDJP9SMx
lxHo0aBWTcG/uKvdrCq36pII7OMGiIURjowcx3EB0qRh42lCq8+2QUJBu2z+XmJo
QaxMtgYM3XZb89/3ryfsQQtKrYA7po1M/5pQPLoZ+zBIWLrmim5g1syM2isoEYBy
39Rr9aDjCfumuJ2vROO/9Ro5wLun5gEQRcQgR+SFD3171TTO1V70SSUcfdFNYv5j
9DceWgkGIv5sfZPenqiajsK/IzrYyj1eqByJuNfoFSNNI6grYNKY59V1hrLknn94
DTBXE5wuOoiW8uPyv4+ak4crhOAKOGVl7zaxpMY6yC/ZAD6GbVsspavLIdAHr2Jq
hq4m+M3we5tj2+Fzni8LOTHpN8cIcaq4puf5P0BVhZmgk2wANJM0bu5bLoI0rwiU
bWB2WgryzkSaZ86Lk3SkU6F+TRtx9s8cOUyu1xSx/j8fCKczik9x0Tsk3XST6/UJ
x9Qc86J0d56zeeQBb8kdDwN9OG7D5AN5KDse6sZ3mGfwW7jYxuff1lhG5PypKEQr
KB7R+h0iJxJQKotU6ejt59+DmWww5OlZGQt3YV1ZUcLN7AHNKJJ0ozUYfZPVElyy
YCRTynqg+gc/LAKiAHGfB3vAXYlKtZmTjfKkwhl6ZaC83h9An0rjtCG0bCztLSKV
L+w/VG0lSq+Vy5LbX3KBarAExi0RScLMDn91QKfGUEUv5lCMPEhpeQb6gCQzdcKb
7WjegCZgNgmkVZE8bQiwDh7ZftB1ftDtD058OQEP3GMctb7radrRFjNk/kXUlBfl
ZGm38X/dPsuGdykEyvpRz0gEqUzrRd5D5QOaLFxAZCMfyUBk+8ljCrk3/oZjKyC4
WlGo0WKYUiETREroGIhO6P2HC6QGuKbLVqBXUX1VEQ4RdCm8T7ZBlptL/16xkcMs
BmZnODnQc0NuESh99BR2d6ASVx7sgAiGKxUsBQ8EkKkk4m5MU8gbT1okxyEbJu1g
clyO7g1ReHijw+lXSN5oZ1x7zO/Dd53j/jVjV91IaLjpqp/bb4/NMhncvMSZL/rP
2phKUaIptrgbb/H2yhO4odhEvsicyTto/o1X83WIXv08CtB1r7cMi1fQ+PxDSDcl
a9s6804g5zYiV4QJvqQc4OtaWQ15A2qLU3J15vRX8ve4RjhPSnLNgEIvSZ4jHGxS
mnNMCx3XXxrKOrrsiYFX5iVJiERIhOEDOY5vTANFC4P/ndJilL+mHNpgREjND0Cd
3QOHJ5TL15ibuOV8UBRhhBRNwiI/cdSVpEDcoSyPymzQ4CCF0XO7v+TAjTSYY7AL
xsoZsSImDBpWGuxEBwvOhMjyXmfs9N+4Tizdc332TqfBqnJzLNqyAI45M0ob810a
v5iAM2SMpS6Zh5EV6+6qkcZRLpPejvk70HjvtXC4/nmO+ljUd2OL2qm6xPhuKQ3N
9emGx//AJAlCcm4d+vQ9Ctg2Dc2vqbiE45CLIdkUmoe06bKA274hjCfQKPuosX3o
qHcS5NGJ8gVqwPb17xlUSTT7QYZIxbtSzn8/lcmcdDh+QR5Xwr4YeBQf6kl/qY09
s+eyzv3ENCO0JMpl8wocMPEPkwjeKTN5FLlIG9WXiG+6RfpLvKX5V+ewJUQYLcVn
qzp58hcTlSfVHDjctial2ZB/wZ95ocBFDVhWZy2a+LBQtDpECGryb6t/MJkT2tkO
rw6pzG35XpGqDjJhaxTtzjPcpHM9jR0bketStJs3eOFYmKXWh8COnVbRz0Nm1gvd
Rwot1nykCPWhkm5xfLTV23lybsugD58N+MwPpbG5+9aqj2qWBQAGDy34rJYZnU+j
TyOEfDX13H5otJFqwVfEAo36q33Neg1KxE3f94MjXbEaB5eZTkntgbOrm3I946UP
6L6aq/tvK03a36+nNjYjQty+9fdC3r8e4FmRWRow0Oj/a7pf/GXRewD3Wfbb+EwT
nNfu1+slMhF1Xgnd55YjQdybJurk8VlzW8Z2cuIqREPsczBeAEKZxI5tZBGcv9Hy
xXkICCKGVy2vRp3aEtYrHK6siOwO/dmcKOZTDZDQp6odRt3qq6IWlKn9q+iL67/s
de1dbc8ucoI0RemV4X8Gdn/HJPImx4xn3pFiMVetkaoAqg7fS6kuoDV9SzT1D8Ic
Ucnwb2b9xZ5f5huBw5uwAESl/OMKlg1W52RheXTmOoYlM7TXH7kRsGJTsqnkTPpU
4m9W8q5obw/9yydndm1YGIM3Y+wc2i4rjperkD3YSB2gJpDIq9RuyOJedkCQYjLG
Klcxk+3oKKadn1LGOoMKL1jJHMt7cJaeohaGnCpRsT+CABKFPfPi4utEgKKJEuob
B9AvIJ7naVCMKzz+vCoWU9igtHs22BEVKz4PIqmIarKayOrzXbHBbqRvBhkWBFDn
krE2iRiJpFTwv3e1dIU0jqcSc3GD/HsUG0a7ONQHKbLfwXXP7YZiRJWepg91BPaY
c2yMAoTQ3+hn4WFIZr4L4Q2SaMOvKFwvx3d86+NsOf/ggc0nHkIghunJ41B7t87w
vBIVuvi8FRuihhW4zCgvsDbR32VWbKOPxpqBOaytRY2IsE9sTN6MT324+f+X5Zop
RXyLKYA7cx1MW8xZ5YlYXGLYk7oaZrFx+ZSWA0AiPDnq3KUIUkos56U+o6FbZbY8
Sdu81FpHKOXk+6d3UqbB4OPhD6JBD/mbUaeIpkTmRAR9idNo6iVy48nHzCL8MdhN
mRFg0xvTvp/7sMuF8sBiSbCUJcNZW9J9sMRiLrGfIM5S9wV1tuUjlCGYtWnw8xUm
liRMDSP6QMDldoAf8pKroFiNxQH1u3ReeI22/t3dyYUgx6YyRLU6B3yWIHOn/KjK
wZdHh+l9702GpVHoAjuA50hOeKzMtRDGeeSqB9r5e3wmCtwAireixtmY6dAUXc/m
e7Is9YSNx3HUQn2KVj7DYZNroZwNtY1+HgC40LqWXkDiPissOTYRJ5UNS93zJOaD
Crfi4OJXHgprrgrej9TskmgVri7jbbX9eyQ/nez2i4LYZYjfZzrIR+NIf3CyH+PE
kWXwY0raT8RY4LI3eIKLkD1leIa2ayR4twhmWEGny/3Hgmsbm7VgrN28cU2/B4Md
9318ZKqWF8b3i6u7sa6X/nSJ8tci5q/0tsDCjElTTN6IaS6mAFQdRIzjAr/RDDNJ
rCJftCeyPFSkxwS/XcC1cr0H+MLboE9tcGVZdXkwFkqyNdIOacgj08Ym4vRtxRsl
4kayxbLF2U8UFrMKk4UDN5ab4N8qM7r9Z/HU8yGnRPGOsX3/cRxIJtrTNvvRCG1Q
u4AukmVNWJTlCMfXOHT6XzJF94lNSRp4Nz4vQlyjOmqSqBmLhSjLUISL9p+5oOxM
SVHQ7KXVIsImcn8bxmp66Lv0lI7Z+W5KTBTSCXdtW+bmu/H39wLbkHRtuz970Gax
7PYLhpEGE3yA63y4ZcCTZja+LMOmb0BeQpRhQlOBnO8HW70GkOTUEFlqAeeVou1s
PkPP8n0M76/SkSDO9lqCu2WR0h1gkAFkmmFRJfqdbmtQvf5N4nKtgDIMPq75x7On
eGzyDce7mn7Jkp4Phr9hUGRHzVCRMOxSDwbeqb2XEQFu2r/67xaHCoagAyFUPZne
xoCOnkqF1A3k5vL8WOb6ixmh5WN6ayn3Nv+rvt6Vv1hqs8Cx0F0HMUseZfqQ7QQf
0HezR+yBlCHpDDz0pcJLL3MfYZoHKwnsRO5ERiZ/m5RpZeK9BTGXBnNQ+zrZDDLx
S2VbDWQhlyVDaaMpI1q/T+gbx/3F+l7mu48pEiW8M8fo8jBqtdbCloIlSXY9hLZ5
MmgNSRV2j69exZoeIbWNwMw3nxdbyeetV7qwVoWE/FR6zDMCxMan0eZ4lUYi3oIw
14k6A+QUsJvhQYAIaunqyyy/f4buhsszdwK4lv2i6xnzXiQoxHeM2FJNOM4wdL3i
AubS9BVeUY+4XirXIEfS2FBJ1u5+vMB/0q+QzVe5RmNzJJeP6tCckK57FvEE1pp3
lVjmpFhebPsMjkcpU29Rphm50FIfzCZASt8gBdQTRjbrE89FgkUn0mUUGE7htGbX
XeXt+Qpylt7Fq3hkhiDb82O8FU6g8dZDkB0lc6yt9opFdI18n3hgAv2RZ8XvPjAe
7zGte4AV8uL/SrGgUDOKOgDjYXN5hlgLPGpHz5uiMOL9xrc4UIZ82VqlLU6cRc0o
fFgideWSfyb3fucjIyAnfG+/QoTwyxPJaNySeXgw3+XqqS5bSHrYbf/lLLhrrMn5
ImDYRMAcrBHq2Pf3h+oXGE2OPf1WimiCSX+wcF9NRB7eF5tsDfSL/gna5G0WJBEO
m/PrW2Ek8y3pDUdGa3pe6Zqwid2NYB/Cjw57qjSssHG56U7oWeXtu62DZaO5JIVe
V9ltxAAvj3lc+sJg5F4Aqw0+1I6y0tL4LCkjoioE3t0ADkyBf9y3cN1YVaeM6hkR
4K35y+CSnTjQg95J2qewp/29rsFRIbrzvBvH7bU/mdDSsbjCKtxV6tDFA9hMKgeR
KCIJ+441dfP3/4D9/Csa94geH9LyDUJVdKbr6P5nfUi5BMNZm4VZ6x49tdpjJ6oq
25uftufp+BIZcuiXyE7PkPXcNs6uHf8rfBAI/ufbEFjbXp8cP5lHn/MF1nHyLQEL
XpdNos6FN79ePmSLoc7aLXsnou6Xk9tX79iNldfFHeJj0PVIGWA1FkW7Gkjrt4xY
M3LY9p9wXEv94nj5gTvP+lUpFyeGijv+iehq+cfkzZ8xBTfy08oWqdG/k+6jwoeA
5Oqg4xgi5fFpDw1Lk/puiyggNUqB6Qrt3Iozj4pi/oLikAIPkTdkVWreaNWUXJpt
MpxhD3hVFQ7in7gzlrYeBBGJg0gkAkhA3m0WtRvmNTigyrog/uWTbkkemG48T7sH
e64K0R09IZngm+vHuVxN022HZ8o+osfqR29lh+Q4IRwgJgna9iS8u9Y6liCqCbYb
C7ye4IlTLIU5lXV03xRWeirmCDiKFJh9oFCkR972I9fzf/7rE31Wy05+awGOJlDS
rvzZOzipy+IQVYhR+sxaUwuqzS8vX9ac+CYTOaD5PYCD/nqsJqG1mwFdoCjugf+N
9O7sdre8zQXGtVozYjIPQmP4nCXm5jZMc72PO7NVLePLni7HjBVZLJN2t9x9Mo9K
eHPuXGV6IZ28YWDsppBrN/g9o2GxwSgowWgbDvwj5gjnfQhVjSPPS2pqLAA5dRDb
73+d3nqC/2+cfKOi7GxE5GcrYeGQ0bayJJu6QXpZstR0kf2w6XO1dRIOmbjU5LA0
AZy/jkbbJB/UCRR6yOSvg0/TZeVTReR1WVLCMjSrKvV1RnBp+0K6fnFxsskhzSYu
Nt/4a7REZlZSpRJ/4SktPbVrDzoSUwTxDJMZ4DL6yWSPRNzuBI14U6v4hx5gG/Rt
K2/lMVLsIg+OSwOpdb94fQVc83XjuO+2HojuO3EIMK5dU2YwwgZC3pny5w+V7e1e
eVxmAu3Cf0ARi8ifagoF6DSkleoALF7ru5chkZ8aUJlRHmPOYpkL8ZknxWaMyKzC
DATwDwOBtv0etBBDp2pionhqagrqdh07mA2MFr1G986IiQeJcxmXrfw107ZNhm6v
bubZZUmE1R9VrMUrHMF5eu2TFTw73eoOP7haNFpm4XbZhwkk5+JRKWLOoO52WUnW
kMWCm9syd76VIPjtEIwTpTkDvA0/tUKNLFlem+ZTDnUXF+zeFEt2j3dC9zuDSwGo
uOzgmcGKhqZvNztbmUtEpCLscjZvRJ6FdVHS0xfEJX192uS+55hZ7p8/v3/Spn3r
0BKGPwzrV5gfeV2VszwO3ucAIgDcpXgZdSQfzPT98cUELwJTpSHRdo36N0GyzjSr
JEAy+Xeo3odfEFDKDMGhku85i+IYKGOhEl1+k3cCR8KhwBLUmUrXKap/uGBZSpt5
R8JWAmuZdoYUWPyQhRkJEZLpOZc+UOYY8SmQV4Ka/j0w4OwkoB2YSm4r3t0ZZVom
WWZ47fJvUeU8+zjmO/0t7OPcdFtBPjyGoWo6WkhtSjXfVYlSFhlb1m5OzNgwAtyI
/vYS5s6/U5/tsKOOxt00VKg05PUp6wwLyFjfEEElYxZbAh9LKopLxb08ptBVVN5T
wDataSPSwOa5+EgvOs6h/20kqQ2PXHsHlVa3WLPs/rVikuoMKWDgllE1ZmxwUtja
40L2nHVuexRhIV+aIms0BQbD42P9X2pKcjhEHTErNNcFkGGd8M8WF1ZE7wangLnD
0R5/qaFqdthM1WRBJ27OYQmlUr4ZhKniG6EOBbtjtWpvRqiSe1YCpuPm5Zs7YcUF
Ix05il9tbnTbJggHbgJ05cuRHcCr1XorVdwNvY9XPbe4hwTRNzy9xmolESsBXKbL
oEl+R1DFd74MICXFhvanh4W0VS5BRMDzeueWhxWB54nQKM2ZzuFVg/S6DG+Qy3I8
enqbynyDXMle0eXC5d3ywk7DMW6CIpsWB6Ggc51sVhJ/v9NWIpb7mq+S5sf7ggv2
6iAhwBAaU+yiRmKJiJ44bXFBWHxtjJP+Lr8Jk394y1eaatnUay3Q5+vfRiFHBwao
OWLrIDAaAr1Nj/rCsryaLhCj/+e/o8VOBH27bcmk/LFWwQD4kjpK33G7nnoWA/g+
GTqqdJZFaGMPuOVVYbCTMsvIWF7xH41ooGjaiZ86ATl0p6UDXopD+xyROmE3qnlm
4OvzfanvzOGkQiLKL+nG0dgB2uGqnAgTjEexbfq8EnvLvEQjXMJA7cUvR7DgzWzm
JNxU421AmBZqbpOngoFluAzPDDCuBGVFf/z7kGsrVBN0fkut4uNKB30+vXcMsC1n
xF1PRg353p1dcfSrj8dpjZCA/K5AxzvCkFvThFOOKYwoP+FMg6fohxMf4V6fL6ZU
p1Knli1U/JlhbD/+7Urc+dz1q69BjV4YbLMFDlVLgt7LasfzML6jkzfFs62po9fr
gVv1vBFZEeFhrtsyQYFehiWP5shtby8yA0eS//m7dmRNEba2MSDhkeNj2C0NovPy
0ShxMhlY1Ztuty9vepxbiHDwAOYad5CVebxZYgIz/b8t39UwjvxVvrbyyND9xAen
06BBm4BeYJt95z3yMFFJ+Ighse+eQ7zUQHgPB2mgqp/8LOmQMZQ5Kx7OR4p42ZCL
/r6vxGDjjOJRECCSsLo0dUhsQFILryaoE574S6fkoAV4joIuzeeopK7js+deW/mt
MUO4i3wBQIab19pJU8xn9gp1ls2xPVzxNPE5FXSMeg40fCrxshPQGfUumpvPF8fJ
xK1V89GnaHi8VvUOUTh79XrbdG+wNhlpEvlLRVTgh00sv3e5upuRIZJTolu2N5se
v4HgOkSrhYnfPZbWsbKHLXkckB+B8aRzLiLqIP9IuI6ffZkam54TNy45vqF1Gl8d
P2yTkG+508xDSHKImuPbfj4qo2kdOpGV8OZSWK2J4JjKVcWvk8jDTU4IJNdec33z
eWVOHfLNsJL7kzWbgaYuDjUy+9WPfPtNy4VKgwIjav8rd9fIuz9Arnfm/C02aHEP
jPFWJt/t1uKo9ocfSrkbBA5eEjwZIjs1iZFhkzdm8Ux0dBJYE9giijhBqAZH7uUd
1tks+NyQ89K671gpnJhIJxTpMfHdQMz1gwJmb1I1+lwHUJHt9ATOB2zi++oMJuZC
7dnZIqOTkIjamg78FusM9yhoiEtXIS52epobT0I8t5byew5lpEech4ijlYgaYtyt
UX77p5Bt4e3yzuS8y8RDq128SdbtSUkuXCOIFA5Tx/XFFB1fUTW343/PCS8h7Qe9
CxpiJBjg1ETie4JkjdXFM0QjQQycvXHgMvWypptnTOEdvY4wyuFG6uMcNgcTt+ww
uxKVVAQ8yTIknurpAldLKa+AI27/F84s3OlY0DweHzfw+AHlRZ6VwhqDa7Fb7C/L
edtnH4ojqMcy3gGzTqM7h+kK/oC0FhoanlrAbkEKNx4TKYrLDfFZYN39soNR/Dlt
ONDbjKqHE6BewYhFIIeaZdg2aCQlW9WFRey3xW/HBVxQS4tduG0v91CNPmjlLXJn
E4vPTzU7lRKYyAsNfVylAGRWffu9e4D2uUDSaNz8adrTwV2VIb6OW2ILo7HvqpZ4
+w7i3iXxmYFNOvwxvIzKfUXyKcGTGL/AakSXdMlkmv8EFRt/nz133SFHCTbUDO3f
n3DOezjD1N9eF3Un6BoiG2/+3qUEQ3TLX46Vu6dlV+gaUtVk1Qg4zRJmCt2sRpFW
VZxsVfj86wy7lqrguagLr+K8L/p4jKAeJ+KwkGgiVxqjtjsY6PsQqqrcRjzXSnKz
NqPqSlkEJ8c3fTDA6Yy9oxdU4ESR1f/TyvyZDQE5yupn6vmKoN90Ml16U5QN+O2k
nccg3Hv952xX6jRWjI+Wjg1xIUu3GwMqpYPp/0nqDPV7Zf1HU9w9QkS+7pH9Fa8y
1O1+gMvgwp4tGs866vYu9r9YghtlgjWB+ujRoP/p1nhTLmQB0OunUNZtA513wOai
aP8HwvvgJBIhiP+rsXWW5HM0unsva32fz9n7xs/fG2RsxwgAq1BLicuEJ6GSi4At
moYQJF/jFdk7bouopqdZzaK3Urfg9BWb3Oi2CqRNY+ciWFUvcZ491uUa9DwKS+9r
7GBA+Shj5nSYH2CCXPmtFiDPRJ424ZY2q8Z8ufH+7chhX7qqOnTQXkNFKu8ApjTb
vJb3+2uTUYIyEwwuHsQq6UXzLo6sw8a29wUBemItWUhPHJTgaM1xG5fHkseMU5oT
86VDGkMivnLd6q8416SZtxg6xWEGvGMOlATslfsF8TuhnjYuFkLxnHRzBkPh6lM+
IFmg7LO0NOoB9wutuOsJutPgA4CDo42Tc3v1+ShtDqjiNnL913q+ky8s8fWoxBqt
jZsiuwlTQXPbeRCNk7PlXPIflpqJyF8MBAuMuhg+aYYqtqZCwWHennSb+In8/8yT
Xay6nWwOelGEIoeFGTe8E+Ry5iNftFJiRPTOCpirTS//Et6eHEQ8hUl6aD2UzX97
S6s688HI5V2IiE7wJQiMz2Lok2HXCNJW0pK9G1R6dfXLUcLP33smcYZ7Gm27S79T
OhcnUCEM7nhfkB1ITpA+3tX+TzDkD7RbpFXeHwQAAKdLBGKj3Ga9IszWzGRDmQVR
h+vM/UTo1wKTY4D5+LNm1Vo2KBif29iiQrRGbOlVVOWWXKnx8MVOtyeyRSf9u0I/
7uUOrNaWqAG9CHSQ7a/u0tLvoT7A/FGbyfmsQzHg6VPFgrsHmuYphqD6TCqQtgSI
zQsVLsGje94J2wBbRip/FYtmjfOAUJK78pj4Eqdw7RVrsGl4ITY9Sm/kRNxZYU7L
S4LT44S8LlAjJlfbDUX+C1gHxGqNW6W9psXh+Q8SR9Jghqd9Lnk+gXA930rrlsrV
T8sWJmDwW9iHzjWNj1I66OmB1L5lJUHsGVU66fDITcTWDDw4QZWyOVmP7isdcOVv
f2XswMoATrbb+AEcxi2tbIu8cmPou1qVvBnm1bvJjFyee5o6Z2MFQjtQ/Xn0gv9E
YGcA24Sq+et3am9FGS1zVKgUE4f6mc8WhUXyoZ0oyM9m7yBgCxpoDO7drZ5Twe6d
etvTDoDoWflfjOZ0EMGq74T4WcUFbQcUD2INs0PJEYw+F6ZcfMKOjYuUoFkk1tY6
/Rxl6Jd9LN8hlV5ATxryOkSxx1R8S75f5T9M0NnGEYdZZ2cKEyUMELDxqlvbCR8Y
/K55d5nWXac1NLcExSO3ojqEgMbVl0S1acCZbEMdfOy/Fz6RcupSFNjEWfpnJ/EB
ILGQa7Pc0tG9HLxDKWymxBUyhRgo4TV9Soq47iLGu8CUIwtyX3KxD35DoDJ9k2bi
qbT+RC+Z7+TDTT2wQW1IDS+ECtTuepli0HL0OFS3lqzlv6WQxyTGUpHP8YblRqRN
23at02EviJN2BmuAjTQRzY1hy1H7i5X05gYSblYg4IJchc/4elSE/NOmLe9SS41Z
spYneODopOWdDDPEI7gW7v4fhJMYZg0lH8uIMYPRe1nozFgT5dJJiBK0XIOyhlYs
dxrbOqL3pFLUYcanyaV0hH4/RKRDDdN6dNhvHCJInaMEIi93qTjTdv8+RFqeF5yS
Wqfq4VOTvG/ebHMOJRZQqRH1exVoqC8pbFbsWyzPADPg3Rl9fVDC+1r88Rk5z6vG
+M/FoD+qjBQwZqrRywNhVWyWhNcT/RuREhttnyuZa9EAXgaGGqmqB4kRJVmP4TmE
/Qh8j+GbKYtlmZaL1HV7CgZRfXnWoRZfuJ7Iprwm4ycY4Rlc54I9fuhy6AEtICrs
778TbJia6p6Y6C+wWfOHRRsmPnJBI7OCkv2uhD92xz7wMFbFy+fEp/ozamelyHJT
RBMWMZ0XKP4yQw3j4+WLK3XGjEIudHNMlP8wy33vcBNX6ekvob8o6lx2f1z0bgaR
omZ29y8r8e8/m9iX5aNtPfnO0VCs/3bKEe6MraCcdxVJUplf+4AIPe3gTI/faqX7
wXRsz/NGOzeizvvOUltMn+nDxnJIWsxUethNwNe0y+OWlLznh4iSmb9NA+Uj07P/
pCCve0cRaudXh3NqcShM5alLo1/XPuX6zcUjnz/Ujp7VMO07Gu6P0DqcJ9a0Dd7n
24f/tdGmZIpycWiH0BO4OZfk7zRyGOwFygaM9hEbZXJ6WNxatHbY7AKI1J0Dq5ou
223EC2Q31e6XU5LIvEjB44hwna/fmmCaFLLoxKJFjxfGUcimwGaOpxQH4KmLU9e1
iEbUcWhZsIbZjgfASYxTBFN4klR6gS55/O7PfI+S0KqTygoqf1WZOnTeGnfhXU7r
+esiB9VdZMlv+4p+ws/9IkAdsCn1DbOnmUfw4IP0X1QR2eljEl5kESKyGPXtoRzv
HPJosBp53L9avbDCdCICcZAsxGjcSOoCO1uDsOCaCh90wqtHS7tn8qGOhidnkJMu
bCgaVmEpon6k61FKxGPCa7GonqTZGPsej/Jxkgch8dgYYq6QCtt/ZxRiqU8XQz8U
7UTde+I7pSpZrUZAYSP4tLhYwVLym0lFmjtNOYn8TKkoJZ6AiZfHTP6tkGzphNDS
S24kzYD9/wsFqi8h4lp6hjJlMUKwBipbfJGOfRCr47zmd7HolEmMQ0gTgkkMUoAA
KIEjGmEIyW2KwjGfiVBbItIiMc9jL1nPVkkyTwfsYU8+T3FAG42W7YNl+rHhrbcI
P65Q7K9ARzcjwuUSNVpnMtSJfXKQYFN2qemrFw6TIn5N3Umq/tloIjac4vUN6X5j
92Rs/NJNwLMz0hQ/8BfUfekZe6aDrPaov8xmbeoVgQn2DARj9eQZTkWGoXwmxQPQ
RbrR5QOk5aQPDbjrP1MJHS+//0Z//ZYhrRxtKZ5qIKmXimawDP8vob7AbGXxb6pM
x/faXutuZuIlj3+ZWI1KAptLMGfa2XcSSOiKL6s5EAh/42e5ncaFfdirhzye+xil
N3x1TdwPJaNfX7XbOiSpBI7wz9dbb0JTgwdNRMH2T2DGpmkKVK3kq++G+0tc2Ze0
ipeTaYSG/M1CA7pZY9+3YAe3pU2W85oNWGsQ7+gLouAxKpplcEs0xw3T1CdHFqG5
QkIJYewPRSoKOYBfk8ncYxaSc6BTEC4cVgPwXltepri6XTFr6+/IWmUxRGztC1hz
WKnAvlHFxrYsbMZsLckDTZrqxBJDXH/FrfaKscIHMbPucEHLfIYhGw7pX5YugjzB
eGTEAFz8eZPAjw4EIk0+iXXPgmsr0n8J0ies1rJXUgIqyPzacopmkeaQ8TXRO+i1
c7zvkI7E9Nabwd8hiXIvD01F4hU0mzRmpp3Q6DUqCiryIalfobACZOu7hS1Gio/t
wyCE6sjTeYyK3RXm5/FCld3gdDOqhkrwkGYAk/C/BM5wB38DjUyw5nOFE346NyD5
hEhP823FBwKlgiC/tdnDO/3H4scsysIsOfO2yO9MePtVlrD2ZxZ+6kjH/srYBc8C
U/mPldEgGtEalfSeMQcc4lxb8FqVfStDATaOtrxL4KKcJEj/GZzQZ1gpcQccU1hw
AMpzGH4XNCys5ZuUix3yJbDy+nbyC8USdBaNI8ZCEHcdcABrgpgkVQrk1yiq2kiR
sjiMZ6sCXOcc4OGPeZVgb+PlTNtj1hwB0Newj//HCrdHSAWG+DbzHRtBdLGSVJ0u
CP1snLnH7ffooriRyD+w7ybtUnrfXlrcDP+tR9AL/S7YMbyTkwpT9zEvv5F1Q99m
tFP1DQ9mKL2DWK/a6AZB7yBq740Sr6Omg+ZkPMGfiSqnpsNQS9BvD2HZNqC+u6+e
ywlH+6cWc6+Fh5G4kQAv3HfeL36E9GVa7BPNtY+xtOqROYL7J5uEXHPDz7T0OX23
KeZTPZrBUAWH3+BKGRnQG8A6SCsMvKt9KwnjOY8ANR9qtHUyr+7Hxie4fxti1C8m
PjJ6bD4IGwtMT+89+tW/iXVS2Qm/hmIIPS6vDWU4hiyRWQsSkGD4Jmvw/G/dy+gP
j09ko2dz9S5LQ1mmVpovaYulggQ7cea0c0Wy2NTsIv8voAlkrVhzWiJT4glfuUj7
1So29YviIu3L6ETjWhSR8tY6XGEi0BfuHA2eqF0RjBiIAG083VERdIEMar+62Ym+
or6eKE+tWEv5e18wf6qaRiba9/+XYCBLnR39SgBiwO2NcbTVkM02aP7sYP3yUwla
f4Znqcn2+NdpzFkueEFD2HKuy95Tqy/o81gIGgGNfqBgu7qyomE0n75YOXKfvwmx
T2SUUk0vEboA7Q0nyc+5cwEZqEnANhDxGGDuDnjFZkBG2FfTTDDoUqb+tx/Y1pKR
4pca4tZEd+ZvjaB23V5+aR0mSr0RYvpFR/rNyleuOksREx7YfBOgoptfbMQSHGxV
NUvHejrGKYqFwngRi7qYG4qtXw7zyuPOPOq0WDhqhTPL5TXCQiT5FQwXmwqCxJOi
5bphZy+QXdgAFci7EfL/fdswLRqguuH7bUMNv9PysJoA0IBuK5sPn6FgzM/FNFy0
A4pbH7IhgslTwb9m3D34Xyinpp+jstV7Hf5dTFx4WAh5+1vXQXbkDgWDR99KDCqJ
v1iQxl1YUM7J0EhT9rSLeeZq86X15vRxmBFlJ3j3ahGtpI00qjpXe1G1KI9uZr1l
O0tZK3OZJbDUJcNL1Eq9AIhxvVH9s9cLepy9OGJrBQeC7eagI/Omb9dbLwtvAKE4
R1vBlBL4lonGjOduiEufYHhTD5UvZvsiQCV/ic6XwWIi7txQnkxGSmI6pw68Iy29
9vkIGZIUmKIoTU4lOTd08L1l0SKTMqWIXKgSAMJg/PtwbLApAEWMQ5q82QgWSX7d
wgETCKJnT9AeLXsVBk+M2/66ZQ5psylXE2gyEBgJFtJoU14/iJNaNrb/+pWBnU3W
Yjbl8UXAfG/cMH5m1cIX4WoC87LEclJNBGjPNhZ/+rASfvW9t6/ZgW0zQBXWI1eE
MN55bHFxdMub8wyP/jY5CH5+Bnzq9MkQ/qmu/B2aLlYwLkszafgNwZyC+uHcR2Bj
En/pIBoTPvpYC/cPbicUa4902zHJtFNUQulDpviBtY9Mri7L+reoDBxVIth6hJxT
+uDyJJScXhmrzNqwzfIF0Em31xFKIIROcpGJt4vb0t7fSQBg/vWcOyzp0A9JUq9F
P0zIC6uKEJw6JmLJTZK9pTlqd2wTNlCYSbPw2iLMzionAhCqnHAWALCmq1z4sXhO
xCDdJMciJWy+UIScfc/y9UNVP8D8xgbtZVhLD/fB/TCX/6Peoe7J32rACycCFTwr
3QAmAfYltTh594IyDkUZH/YXiSLH7dEmtzHFOrlQXzPI3pDvk5C3ExHyWx27AO5U
yaywCLA1QQuQGDujhUjFrZojpMGcoEjfctaaGcEx0xnQEN3JvhyRJjzs+GBK3P4W
h1RP+ApdQtBpLHueB7zQp12pJWbxZ+ZhkwU34mY3IdjubARjFUNy3p2btZp5EgwR
FhaVTgOTJB5NBJeRtAqWqzROezk7irfQmq4g4w3kergBBz7ZCNxsNDL+bNG3dzPU
B/dfNdURki9ng9/q0yfdIYFRTsrih5ROUretouZDqikq0czhYNFmkxSGeiNcQK2u
NUI02orZOzGOssSvlx/+X2ZYAVKvMgz4i+PfQsigQSaD3NHp2J5l3TzqLag04T66
r1mez8lM7n3ZeOP0ugzkrMBxJK84pNiy0dpTHF7FV07wCeDKIvRSbzw82Qshpz5V
+I2Dpqrf2ZJErQ6ydMwEjZi1zHZwFCE+qEsoG/2JyQIQNTcgnYL4II4C5UKwoMT5
ZIPh9pEj5Ez652KaDQfdACR+ZOEp9qrhRVih/gWebjBJ9dYQdx48DGSpq3Vxbsyh
WZ3bcChxbTVKeD01UmYOt9Xeh6Hd7COSR2ekIH8cC1lwQ4WzJxMuWDU5AcAd5tUi
g6yX+Ys8vMYtIsKZlo9CvLfLBxWmVPvmhf48PguDxp0dIr/+xONS5qL9UU2iUTXH
J4rdKRSoUsXBou2o9imMzqUCPuv5iqVIMDUC3LUW9dpex3YaD9JvGl7uSZgTsERu
oWbTIY4f/G9MmXHL1QeszaoS2iNSc2zCbmxt0KvDFbn+btjO+RWxOMHXUC1UfeJZ
Ao+ZbuK6EbTpaMjoxu3nxS98x8CNpuj677iTrv1oqLznBIM6Xx+fsT97amV/99Td
mFf/TiQ/LnQqUm1bNtX/NZW2WspeNvjiNdUFuzbLOxPAPwKGORrA/6mnGIG3/LEc
Gl+vYUJpE6qemiDKOe6ktnzLbY1l50zPfeukM7UDOYlukvnihTk4JkkbZXc3ikqj
ADhUL+ljkn1n207KDpj9EFHjA6WoEUufB75lbn5hbcukcle+dDH2ixeOvOou4CHO
auQobY41uXnFVIyc6BHTPGefIb16H2UDumXlmiWLYxavcgM1Fnvry3gT0O8O+dXi
+3Q/Hhn8CPvEE42b1pD0xHMwjdsi2H3o5NF82XFAELBM3fq/LEY5GCgQt0aNNUNJ
9qPtlDQllLM841hrgWGHjyvat6/p9xj4ZfBP0DEIbh+zUACe6Olj7L9z7TNZZn9p
SkZv9VWWbiV2M9cN+Nth592QEg447aO+T5K3vmdEagBVduLkN13d8A1wVhUeTiHs
lHfN8JcKQ/COlinPzh0bEsLCQofF8rm0eeSy6znd/UJvfehBBsoCTJEe6gBTmBP3
2+FcJvI9cEEmT0At6Ogg1w8qhVWRb5r3nkTBznwl82K0UtgMIWy0upLO2DpbnPel
WpsD64GUH290CxvuDQnK+YJu4UFueGoKPjwxFeGjrqKZQTjBli1WY0/4L5m8eXr6
VFo6pWV3qVA496LF9yulWu0cL+7+Ev6JGCHm8+T1/0xwkqHwgosbB6CfB0G4HlCM
4oB3+PAS+o2SjRh9X8dADXjPZXWEodyFL3dg/uIE7A2WTE0iHIhobhsY/HzU5Q7i
C83P1V8L5rqsDH417lqAVQff4VOmWQovf76eIv2bAOZjlMT9zSBQxuoMUdpHL/J0
rIyEUq+YiFI6jMjYDAUlnf15Y6z/PL6xocPtVIJkA8Y0OxycQTES9JxRurhF1aCX
Gh9BGSyGCTzVPNgItgTCga7hN35c4dNgyeOk4lCLNP8C0LtHkhmrYIoqBb/nUsES
0AvzMpZKWg0jKxAe2p6rskj+SsJhVGSt1Zzyvjo2gUZTs8HHiUcG4b61W63iV/1G
QxrT0Z2dGpCg4KfkfMlKN3NP53h3oqjnibbYd2rDce/jdHZ9mHUZKo0bAHJVKjlc
WluFkbxKOiMm7HBpHxH5sQS/+fqTkjXlnWBoJHH0DCFwTdUWn5o8xqD3oI+hasU7
di7+T6+jIliVcxIOC0lvn1B10kNJePzwrklPzePwm3o99kC71kT/p7nUuslkUVfx
6cwbHrqaUUwrrIsJ1Ju0dluyXx1L/ziGELMR1wI/grdYm0sVj9jQmUscI+4vAvZD
BHOhPebhUt8oyDP9LLpKwX6CD0WvU9lBaWxqXePt2r2uyIbfkfebphpIxIryzdoZ
sJsFzKmulaHGSmqEsJ0xpSLfuFaBjdyUa5ITYA10TTXXEb3kf1uLCvlXHeyTfMgu
ym9gMJIlzipitwYZNPHbvBCS6DkBVN1AvX/Tz79ISS41nFG6iW3WTO0TqIcn3CEe
CQ1c7K098n2lx1D5TZ/u05ee+f74wrwo7gHiWl4sjHEhhNvw4jfM2jt/BH6RfB3o
C6JVYT2SlyJHbBoPmZ5Oc/4/6Z53r8gjUSb0boAgdJ3tVBHVNgmAOn+LymmF6l+q
MSTIrRpIBSKVrePq1Yb55wPJFA/0ZHKFaQ28LTBO751R00wp7gOkZ7C+FhPPS7zo
gbXszFf4pb5NvcJiag0p7AHhBFiSWpwU10BPFnFQpHIfN9IMmki3SaQhiwdSCMwl
NC8r9fyZMUzsWmBFBh7CIM5+ouKft/FU8S7NRepX0IGRf4h424pLep0pD7YVs3eX
jDy1noTJWG5FySZ5uzTl8CDRN8Skz2AFNWodfRYvcsrUtglPoBkX5lDA+SQqTUnZ
jjE6Jl/YpDrTQ5NoJGSfr9wLXbC6kjR6eerynW6bNukFaDAcnhAa/dQ4OJi+sK0i
Z1q/l48QrzejuH3Jos6hZgJEv0+4OgOp2mTYq6iiCc9o48Apk4Mcr2tjSYqabXkg
pvZvKUgwInaVDKQj8vObpV0EbnJs3kJtkaYCWhZMSPswo7VTzyhVOUrvXCPuOAUH
8deDBTGkR6MpMBGrNloAmV9Ww3Ots5qCH/pxdIl/FGjvS5aYsQrXKhF6waZvBpVB
gLiPoQJ3YzOzL0/7fe6QxcUzx61P0oGJIFrr8IpsZWKRo5ceMJOsmdPgAEG/Vb4+
5g1bzdAZYCVHFA++vX7521g0pNESn3TOWsQyhvdESL2CdCjsplUOHUYiVn5qK/sn
awuU54Q/ax7jLuRJHgwQCoXTITVnsvVHx1ZUXWr+esfnmrZLnXYi75HJX8lqapDc
13jI2qS9J2dbNBW+3u6b9x1PJa6BLbh9WyrZc8bZArd6sWjkzRlHX9RITITOxtOZ
mRXp2+LiJmETZlN4/oytIQ5RFqpJnds0ITfJ4SOf7JTVmW1Sj3AuAXJwjcvvLR2l
aoBTF2lL7uCRLQzuQVf2CfH55oXzNeYTZV2rI/4wLtVX3OLDeJsAcq04lHPRH0Xn
+BXKYshGN+l5DiqfoyR7WuZmFrczkZuKPSxgsHHAvI5v0sDJmp2KA0oUVhwZaoy3
qUpzxOlDZFXZeVSpHIXBx6rtVxEi0Pp3g3EsxFKfQiHOw0/RLLJPKrNRJ16bdGNi
FH4NBZFbJJV27mjdDeVSsAjdToskGPvHR77WE8nPNzJnTnK5V8gdfyeJYPwk3Wtg
XLqnWJ5uZf3kutFJ5x9ykCoOhkWGmZFHbLBjY/zmeRU5xJbxDx7guTc3OAHkb4fc
BV+Slqoysf3qU2To+VeNuW/7FO8ZdgLd/a2XFkULTOyQAD9dfapxETglxT3/yJDp
DMaucy6OPXwvugFO59kCamPu6OiVX9HjD67G6az5lTR1xF9sdfSsdeAyKbiKuRCg
n0z/83u5EqrljVMHWtx0C03+IQxe017SpaiwxMQAJNyUFgl2Kw722jSNztwgk8oM
mIoQhZJqNyroFpKiOYI/bDQlGyNDL9HgBv0OynaZ/N5rKURTQi/DHi+xvOOgX+g8
DLFidbO0SabyEXqK1ieXLdcN9XRc9Xpgq4bVz5/BxYLiKgU8DiKujgJjOH46cqjI
T7HkXzvt1qnvoBS2xtQy6e/Aq29evbijhKtvZ6GdzJOT93h/0tsxI0ZnzdCeHDkx
OFkvLVZtlsXTHGKKA3o6SZ6zpLxYXXeIwEf3BUw2GPlh23NI+71Y7r9qmu2qZnSm
0TK915HnxhrvCp4BP3RHoNlg85yKppnyw2tkqdkSM9ec+yE7/kcHSHstL5vLwwMC
LOM/TwUk2voW6ds5nrzHCTpVIgCAlwZ1OImJrGbQbP2PhEdXkvcyGd/cjvE/33C2
HFNVwVwC4TrfU7OtFTw238OzQJdGvJ9n2Wycta9/h+sF76eUl0ylAbuE/Mig1iUX
SZXi/ZbXBuxtPs7HjC8T09B2XYffLFvFP/uRrdq+cN/JTacLllqyY9T+7nzljK5+
jb+ik7c9DTvX2qdv1uVfUA0l1W7pySl85gW3XTb1BUzB5P9rF0pOK+f5vUyZe1TC
SG0yIffQNN/0fq0zsJud/lxGN2KdtYJm8PYOlEQkvuBSPFa66m9tB32Damg3GQba
tps5F5GJvK9igydPRxcsWKCm+fUQUcgb34ttKGdI/N0p1G0nduBRUw/0Z1lkG7bG
uaxEYkTXoVxnQQfFP3QGpl8vRbh/vufCKTvRMxVbEZ2HeEsiXli6KQFAHtau1r09
tm7yYaSDFYa+fbljRe9qYI/f1pcQa3IglPXzw+dhabJ2NEeO1qoeyA/YtbwBVh7m
Xv4n4eOEW8sxvVAq1/Fv9OwISEODUQcD4PTBQyNqmjxozuS3SvL8cdcWHcAuVE7k
7pu9ktbEZ5LHC3y59ALpMSLUi7kKYOIFhZYrHdZXJuYk5+8/18QjXBmSoGIyc4De
Cfm8tL+xY5uegOEHctSVvcCiJSfQ9inGVZmCKvYGZ9oc1k8ONsGCtV5Jr1ByoGJU
g8p5eV3NTT9CH51XFm9uARTuUnELQDOZvwAMaZE5wfutB9xyauSW9/egv+vJhFLa
QZiVxYFw/JtbQR9/ZZC71PoCi79fEJQekkvBLQ920tk+fTPQ3rvPr2T6cwufHhsx
kL0Gt5kzc9TG8Uk7oxbumUWk308YBPj1EfhANSu+08dVlVOB0nLp56mzdf78Ek8E
A8RD5SjlwNvIinUkfC1iD4J0KZ2BMcuFQgrgTCdRd0TRL2hwHmJEkx3A/S0djTOJ
abDddl5q4iKZxzvKFCqwPhvPfc8MnhzkdzTq8cWhQefh0Ep05C4S0BYOTeuA3b40
psLAQzkLXnIZY9RppkMJ8cF8qvzItbHlzBJOXlEoI4AiKfNjtthcBFKECr/hCF2D
RaiqYvWoBi8jG9LZXCDj/2YXQauPqfJiv155/Inl+Vh7zwihnYNVIvTJBwfOGBK8
WaGNr4NS3xosK9cmXy8GUPQYs0x1ONMq+om7V2aWDSMlcP3vK9Ezc1+mPO3dDccy
yyt4GOjGAEu5WUtOA/KPFisCGsj9LBXiGUDUugeply08fWeKB45cVVhtp7RUIuLv
2F2pJWwOms4M7WFTjH6JfL609Xn8DBJIwihEcFH+IWszBtMCgae3ywHldwScapwK
X/ujs+ahxdsfxThx1H4zMFveGb78txQgJRrImc5rv/yJpF/gxnVNBh7fOUNCY4/e
eyEwQF5sZkBl2d3k5egXEP6X17D5eCw3EYvbyOjVDE7PbAOR4zJluPcXf7/ZN2Th
7bEIWYyO7PxB3Kk3mEDIN552DMKObxqn8K6DRZvp50H96y6oAqH3Be/ElolCtpmf
2dawsk4zphiOPYnkx33fju9SrOqfmrLzxA8JvWb6gbDo/ov6mMAp61ZsH6AFmZVT
lDIheIrqGMQT3WiteENLa5k0V69T2/a5lM/d5tLRHpFfZkNOaJMy+FxltTE/sctH
gZGfTcV5i8IdI1AYEb2rMzV9KRhKLjM7TU5uOiSV+cLCaXExPrKY9CA/ZXIUFeP5
hgjlmljC2YITf3jQ33FAOAF6P/ao2UsbQaaPg5Flj6na+xNXTLFNxG7U7yGwr5Sx
4m5T88qh56CJu37KX24y9WBMSfdRnYLFtYkz7yUipprowAW0mbJSGv8Ws5UJqEip
NTCCEZD9pxwfzer+y8drBRAMhza5QAilQwrUUzwzA54IuByRoL+Ugxd0NHnEZ7DT
tO1FNfMb90m92VogFZquAdpCfKf1GvHSr+Rr1q2Bl2EfvHFrNkROqsj4tewEfHk+
kAP/BPhkMkqbWu35CMXu41J5N+/RZ4N5ulIv+uMGs8aOb2HEKDUrdrVdJqyzkbI4
bbd486MWPAFfYlnbT+qsazGq0sMU+8VPjlzerltqZBMyFyIhWw0gAoa3Ny2JC4Ki
j9sYW18m6QRPVLW8z6jWMYO7QuZ1ZSEYWQWLvsWJTXfDx306wTd4DzyzRI8dFiCP
6Qf/HD9Hc44Fc/CJZRLkEixzP22SkERToJhyamqG6WlJgk2i1rAi7ywBtJmLsX4K
QU5rubw/qj0+Wp1RTYe/A1CZIc42+Y4lehKKQWpdR26t5Aw89aEYdT7o5V37gHTI
Vfb4zD16WqYCgrWxjLyC108E+rlv0FNZZi6IoNHXewT0j3Q0Jfjm7jZNt4gNyZos
fe/oE6+wv6MjyY1o4pdsVUxS8nhYg/KH+oBV1om9cPMWIKiAyT8X7l+37CYOegQM
u9K2gxH301kAv/rxCugDysnyMinoCfwFIdBnX2mAdsnxofz+ZeFPw/brCfzrWQZk
ZEWeWV371Vzb/Y47ael6//Euw7AfzYyJvixOz8I3L/HMcldUgsMPtg9UXlunky1P
4AIl9aiyNDoN8S+qhAjNHRRvQ24GrLxsXi/J6RYUG/TTZS7QuXOQYF0W2+k4ywvf
NdOpRh8Swt3+TpnijVkmpZfIBu9ona5EagynWJdrsuSZCClPs9E3WZ426s51QbL2
om5GGrh3U1FquVApculAS9EQ+634rOlZsrpC4XXqrMJd/efABSQ/Li3dt8l4kkDc
Lwz1eu77OKDNrXe9WuJdlLL/bU8Pi4x3wXkKDUhIS/xRyUFJ4XAtq8I9VSAlucfp
I2J+Fn7oF0rzGRBUYe2mmZ2jj1uzFhz9JXzRTdU32RTBiRv2koK5k9YYDmlEgJCU
9u69UA2jZu+vpLizBks29bUiK1pqwS6YTl+BnHIuNdk9f9i2YU1Z33QMaksciqWh
OnavQb6Sd2XILgO8gtqU6ndVIwkY/Xq4GQUtCJN9SDIs+K1V08Coh6tcnRvcaatL
mMj65JsLOIux+nlN6kRDJRLQh3aQepNY+3qwTltJAq6TG31XXTMoJP542hyYrwpS
5XVXYeizTj6bcLnFH3ST7PP7xIl6id4HYQrn9WZoUvVsUVIk/rIfldimQHRZHcnm
eDp1hO9CegM4HcPAvWaMGhEA+voJBXBPGAXF/phy+dmJSDLEUYy0/WQsBfW+lhqu
rt92fbgVJ1tgko2VHGdVGOnZOlrIGc+6RK0ZEZjErSWYSe5o8vzoi+iIPdPsdNyD
e27CuAjOPMxeeqMkfIEBRFkd4xMgW/AW0kEXEDGza7zaeCP3gaVjhZHqOmPsnmrE
YQdiKFIlJf78JVFHtIycJK+IKsBRH7F3XmHDGDT2XX1AAYxp/MB7TZxWiuojimni
Q2EePxeZ9wxWXZNpwbDEfzfuGlFv97foBZSDn2jdqLmVvQxZBloSLW6gk22aeMDw
Ak5YwJgof8bzrCjzkaLzeu2FiGXWRGleIiK0p4PVYFaOgzCKh+8Bd8ECcVa+aXrG
3NPbf6hJH5SjsJuKJjmxCVWw3Nl6qYZZC6E+sNhZARTcYrAxVtvrd/j6YkCnPG5F
PINHPqN/tlFdd6+LTOnlVerRe+cpPM8AemJ/8qD6mSHfSJQjH5jCJZyYnmwKV7W9
G/+kVNKcZKr9YG4tFY5KSqFGeA9FyzBuX3iQY2SrrIX81YeU5yZL10HgjAKav3qY
6rhK6AT7pDV/ipakrtBue6CGvzBYhVACi6TvwAjkK5+X15qDfv6Q2LdHLNyqfNon
1yqAcWxsDn90ojZ7wI3JIF7WvyeJ4gu4gM1iSN2VfS9H866fT+LvW5YrUCXWrLa4
mv/62qgxImX/WdUc6Rgg39S6VR8pEubg9z+i8kBNLnRtdptvN4Q8tcfaEc9h8dDC
zEji6hfqZdxePFtN8aGcfn+Lsk7TmenUbtTveQ/bsnVOS0YyZH8ZLf7YOyX7Z4nF
3EzWlnBHZZyP+W34zEmlKNtfISFRvHxoQ0k5MqV2zu1IYbUpHxR36o6jU0VcV3ic
Nw00CLcJFdqbOxjzZctOKnFCioM4wYgR4iuJd9vJqJmobmK6FHW3Iupr8703Ask0
VAvxeXiBnKL7IY0wcbFbNadjJRKmqx+zd7XuZcCqquu4kiTCM/NgPSMsUWB4vXmJ
ehWFdZcPJq24MBxVMR6MZs0s9x+akgJ3f+9bknmpOe4pVqLrf0bqHymAWDAVNlMh
vp+gdD+Jt6+aoti1Wwkq+1gV3NXrkX84FunixQFfr7nd9O/KwKCureQd0zUQvntb
9cjKT140mhWEdbLpk0CzaB5YkXEWmxYgq1cAXbNELxavXovVTUunLnSSckolB/6X
MkwPcSB5KM+6QB7b1U+Psht6BVlA5YAzlyAO8kAuFELl11TtuN8YnVt8UqThzIWO
q0ZMRzdTF128xCqzz1raYndlpIo51ixCy7sL4b69NGA9n/oLS/0epMvd0BE0D0fx
kkHpLtCehN3nayJTHCYsVmyxxDYR55iqOhSEEzY853Sy2YtGvHuNjYOjcIi09Wu2
KvHss5N4vpDXeTr/JyVPZIJI639M17FpNlLJs2GyNpF8nvSDGtmiIJ3QTTKNYcoo
hBsBLJ1M5AF69DgFQltVAR/QlVzAE1HOwgRCt0vRIOcfKZ98a9oF4Qkklha3k2vt
S97ThHxmcqwNMLw5D55hoEwXFvgj7fj4Zuh62xJVppo3adyviRuDckLhPoaekDMs
nVU/4VVZzU2Ds3rQPnz1bP2eZOD69b77ZvazLoTADjgu47AhfqS3yfIUsaocFP7X
Vmt7dorQlKdgZ2pJ6wh8n6V2ZYnaBXlCTXnHi0mqRqvjE54ftPMRO8nUQWVxkhZ8
ix95xVDAT0GOAQm7FodmylTO6cqC5/8MNQN1pkiMM9OaVKgOGUmS/qWPNUSGCo5E
Z/mvKpGAVbTOrz2X4L3jyRzgCEgtL4dmqTrd3fexhR2Xtr9VDTc4stICkPVvGq5v
Zvwi0s0i0TyDFChgY99kWN4MQLkA/fYbtpKH5le5VJjB66Fe0pgPawo+PRWgCCxQ
Cx8Dp1tZD71zE6NZ6q7rZ6X8GZU/11kJiHfKv2IQdDHH2Vn3vkKHNrYflbr+AZi0
VYTWhDo207C0PevUtsaHoiPqHZxYGwqkOC0UlIpGQHUDc3SKW6BnKACXa1fuQlfe
vizazhf+RFpYzM9jHlG4k0IrJCk2RjhnfKO4lPpsXfvXzuxho4UXnNE8b7XPW4Wa
TIxULAK/67tk5fnFaat5ahE5I4ugyC0Tz7JBGJ0RPXbYaKt+tI55/6GoPomwKm0Z
zhbg8vtIcsqQ7M8JUdJBfJYdkY9dieGZI4rypY2wqRFx96iCOVZMp7aapbJuXii+
fr50z01h2EXXF2yRw6QUpNyjkpNIUacGK7Vt0KHOpyNeKTCxl+s2IwBuXx1iO4fz
HJg6zKBSXoFQNIfKSxWWMC28aLLhcFpKY6Xk9gtfNLBfYo8WtFHkTXf4nqs1myii
cgXOEP8aNEdsEGAPQQH2pjOVwN8LINAP4sy9MSzl/RFZd5nGXfeqcIrjQ+w7n6LC
2CuCPgUMi8EDaC4qrmGExRORvG9D0mBrRNDV5mlTkVU0cgncwWkAvjf4sGZ2K3we
WHQ2aX25BqwuZAxugGXKGeXnJB/0pnSGex3GHFmQ0L8AEnU7097fdlbNPffm1quE
i6K9zlNC4pw+vNQxxupGdFsrFQV2eJnPTPX9OY+NViFOolfBI7MPnvP4TUVZ/Bze
OFo5UvzPBssvjTJsQaElGCA8ePVCKuouKM/Nq/nSXXrPRNSfqg8E1SonE1HLvetb
jZfuitnlLLitjw97I/YtyesupW9RFO2YTvwSAqhyqFCTqGs4hy2vHDF/zWI1BAPw
ZCb54DF2KbAG3aoduwtUwPskZDOmwKpM5SGt7mARmoYDfw2SiSqrPDWlVuUHw1g4
V26/wsYH5Fzkj4QYIKahL83JSIMzi5d6eF3G/H9SGDsBNyLssy2dR3R4Budhao11
gJyG+4pTZPYAC5duAccYfyVmE2m08BTBK5og1G8yVr7rEPxhuMT7HEAxLNJvYhsH
LcJrVlqVfIMTZoxb7IS4rIK+p7FDQImtgKP57phT07Algo2ssBRTNJx1Cl+D8FgP
dxunPXicFenj9sRb58ZEs2jkbtLm7RgWiPH751lqBvt1PsUtergCNCUot6SDrbYK
RLZnJ3XdCBx2AAVRu1L+3zZNvWTm4otqSKUw5IvppJAA9Dhm7hDK+hRSPzA4Bebz
s5vvGHY3p7suSgEig1TGIWiKxrqVgbsU/bgJGdQxbKfmHFaWp9bvajICg29RiNc/
rgTMmJeHVH6PRr3PzJ5UHMHzD2D/H4AI3vbrR+HwTeSiICWLdSdRDajNjiLuPdow
Ozw6qdFBTL0GWI9lmsWRg4RonKMKnd8HGG10eknCRAYCEjDH9wzNT3KzIb2C0SP2
eLi96W7OkZUf2klxXhOc5CpUMP6yfrC6Qxf3L4TZ+E3RbVEElVus4xevaskF24sN
6YNVFwCjZ/83NkIs2eZEQniztGn86JG5C9X1jpyqQJnMYHRGHVlxfXBHR3NtQ6Rx
/OX2gtV95CtUQJl3D/xm/GiBIwOsBA4gjP8T5ocf6JQT7FNv0CB6Kfqc695zPUU2
yHRpousWE4lopOEwFOPY5kqtocK7VdqrGtm03f23MO/fduGPgsID7C4xgQMonbD8
Bf2yDYAn03dVFw0acUzLkvQxqmH/Lh8WvXT16ApeGPClSNAYFjqYTSDf92jTQ4Z6
OFkS19cZsd8SDjbPq+4oC2+kVGy1CGjq49t2vbJHCN/GkvdD4hA/RebxgD4emyiE
KgM7nzcuYigQgx5DIGB/x0DbK5VmEQCszb7VFt6VhP0mQ46tQL7TYxJHr7xTo36O
f92G1FyMdG7YOP8JDVH59Ey5+x4XtPXMbTIqhIDU493H23J8wSDhvmSmhpFB15rX
2BopK7yh9WyKjq+xgi1pvd3VuAeDDSgvJCfCOsXizU5+n40w4EpU/1cGOEspBDlQ
3qfeGZnx+9XN6xRMN2qa5O7tU1t33aTLs9KUPov9BbFTpnK80gibjhydJNVJhr2q
2RkyBeTRnn1GNM5HRs2aEjZJ/CnEtx2JrwF809rrNoild/b5HLctI7X+X1esrVaR
6V25gbdqUzj7jWt532FYoQQ4NFXtCHfg9sYsarfvO5xHkVzV2JhIfYfhU025cQkC
TljOh3VLO6gw50KSLcLtMVQZafCQ6HOvKxfoucwGz3JsMtIikpIx7Zj+1kpnBrvm
d4fJy2Me0vrg+Dw5pPVi3zaLNSRb9F2fhc4JRI+gv+p46QS+3W2y6vDYOd6C+Dmc
qVeU2P4DWxXDkaBji+qcT6AGNMJz43jPgt8QyhgR1hfmFw5KLtlDbCSH4E5OoYO3
IKur19JuZOXg0r21CLtPrterT7K5YY9sZa/FM4QF6gS1zPG7KA6LdzcqSy7LTTUf
Xb7qTtpmlyar+M6BaM9CRkh+hR0l5Wif/9yKkg5O25p5pBwjewW5+aaTN++jHPZj
/UZfALvBxWidL1Dq52rFzSwvOWiptfKumwb95i7FyFc3w7PpHuHVzU/lrDxwh9sk
+OVNc5ElLXq4CygZgMt2ohChHIgMzFB3cIvrO0thFnctn+V/wTFx/qAtCsy14uKz
u1ru7Y2TrJ8GvIkO4rwuYcVoZGubYQ24AU6HsrGdMrCHIbwPgmsPzykhEL/evr+J
E+CSOCin8ABzwUAeY9u1foYKsDuNyZXyIJsDyEt3Bw2V3RuLD72/AxVnxLujwAeC
Bl9nug/SuJaq1RLr5qn8zE4r08j/QBhx9zpDTaKmlEpbtxvZhDoN7O8F6ZjG62rP
ab2/rxaJ6gWQMt0x6zb19FvjvS65hCdh23h74xWP+XNWdMW3P4Kgxq9s9QGUnmWT
Xto3+HYFOqTd78ZRX/5SJ6JANfjSjy8R4k27k1LacxJQzsn5o5vEKDsx74Fxngs/
J5EBxI/TfW1iROdXtNR+9fp9U0v1+Impzj7cxWcgzva+4SfPz6cqf4iMNHiy8bmC
8XplYC5SAmId35C2hlRoOXrHnhhenGl9q14w6tceS2vmYvZbJheabK1mZFpLIWmH
l8ucnQveAsgmcTr+50dhUD3oB35pl6rPsxnFWSEFP7TlMf+H/dHphTnCqhBUso3J
AGwSAOGa8nw/TGh2hOclIpFn94Swzd4s5xLDpchO9+h1edI97tc56oYkPkBhy6rQ
85t9m39dXBdDAVwWmI9WQC7T3UM3+fU+4U9X4C9xR9E+ZDdxeab1CgjvoweXKR8z
6VnALI0BzZ32sQycc5hRnNZl/Q65o/tztOW7gjsIvjCA8K1VlenW1GCMqIKlVtJt
hZyxgCyjzBbjnRnb4Cq+4UOacNz+Pbz1Ko915Hu7JLLEOD2EmmTEzMaHO0vk7NpE
Deen26caMqPYpz6DxLRf2qwc9A1DaQRRhHNPOdx5xJV3zYP94O+CDPfqWD3os5M3
Yq1yBHm5LbI87LpQeZ1D9vRwtYAJgVHdSUgRXay3xq2kn3Qx9QCmKoPYLmCVAue1
OLRgYH7uULyYSBCZSlX9iqj89tup4NXU0DrM3PAofeW52Uzo/Nk2hNtkVLeK2Is+
Bsx1MtsROrIhvcSrAnhIIuOoCFSxyr4h1Azb50IxwMoVmWYw6g1w2kVCChRqY8ox
ELVlodS+TcBvE9ewkNMEAvRQWCN+n6+gvo5vNgKi2VnezXJt9SAesU0RIpHsiNze
BQQ/c+7By/78NMXRud4JLlHlJE4uiRZL5uwnW/Ik6lBncSYEHVhhLj1imkSb/7HR
bx89V+Gzx7+iMkXeRau73kAgz6gbMSO8HjvLK+vEn4BOqtFtooxWCVCZKVUXCHMS
F4VR98aStHdbDfN50qrOX2f8ILhjcY4J3+rhdSXdaltvurzJa+4r34JL8+K4QB1H
udWu5g4IaFCxF1MjZOFbGBbMSnJId204jZEKWIeXo+9rFHFP/J04agJCeAIwwukK
PPibbqsyajPs5LQiIiLVGcKDF6vOxx0I98Q9wxSKnN4zaYRD+tAvj474lg9f8VEg
soo07b7gXOkpW/voYZicKB2YXtwi7cQSKcWazmUUDCoIsD5KorQz1b768eXYuqdJ
A5fA/djet6cmH6aVpG11krnUCeb9JcF/inL7kl+I8uYpZnKLM+Fdl+iQj4i79pMg
Ou6RghjRDxmuyEYojAfrgj0eV3hVfJ5VfEjLxTy050ciBbDY0PUeLneF0oswERkr
rLDfEUdn9b6yFp+/8i66DLUrJnvQkHJotvebSYKEfouwD86jEsfj2CyhHDAxVrMK
cbYcK1sauBBiu2Tx61qTZScalPLg7hW72ZuxpsMsQP7/KUVMpj5bZ5Qd5L5HVriJ
Pu3hudKDfYx0bLBT3Z25hpyJ8NinokHrtCvkxMYFHDlRTOBbAZ4Lj6hInKSJETgf
Ko/isYny1act8R6qgI3y7Vlru634eM3nG9hrGGWiBbL3QYA8JoOusOEdP0evbbZC
nE5WldAkk/+Q4DkiLvL5zzuhZk1BldbBNpATx0Jq/FBGb5IyO51CLV+MSPZJ2ubG
0wVwLGZBz3bBZ4lWjkuNXokEAf9tltvSFjyO4C0OVT1XeFRQC2ysa5Eyy5UEmqMG
/axFX7ioehfSVF530aynPyQTtQvLRJHzYK2Aygx8wclO/Cfd8v5f+FD61k1ab5yO
GjTG1a9v/Po+dYzjJ1RbplSqmx+Dqofppxpr5NVMQQdBMrmiuawaqI+9UB5F+T2F
BdREFcecgSgvw5IAIGb5WZyOB10Gqk1itRq5TxpoZgxsaLLnfSQJr1VNpCPFp20I
4/rzSW2LQNdLNnMw2LcXukAe6iRlIVifTBwahmgg1+wrxR8mxCf6RkBoRsmjyosC
VLwNNHsdTtPNmywfzQHN2a6BIAjtwuqX1mXiARpkHrreJ//eSsiFO3iuqWok1YMz
2gidAa/i/yuG0e5QgsdOvxwIQONl2MzMi9zQm2TBCCOWPqF7m0Q8cmLDbwPWVMK8
HOycwP9xm9bPFs49cJkWgj+TksAGjFHNjYgzQfAwxpPfOdm63z9fjXA1CfMlvn6F
vhu/u0bxVbPJVjNM0sgj96NcRlHor1cDce8slwSxOZgDyE5PgES3XQjRBc9dNslX
CvAKGZMGjlzW9H5rXu392s4mIxGwgtqwQvHp+/oE10/cigKyocNql/7G8Eli9l53
c9MO9S5xczam+iHftDj36y7Z0gEqG/qsl5h0c/3n0s1De0LtSxEbNo5QlAvVUTQ6
b/wRMRcpeO/tzGndS2zeB8akNzhEJajq4x32WLUNjF67P4n2m0kvLZVTgWzrWq0e
NVehsoWd6VZ22Bww+CJnXvsrER5gq4ZwHj49lLhoPZgJAfegfLWhJkfmF/SF3S9g
Cxu5e50gY3vohQ63WYZOa9h2alDJ1znNQsY+gPkbgKmVGx+efyI7i7eETA3zdFAr
nXe3/WKZHxZYWCzZqT9Y2bkzucsaR7gYr3Y/VOWjjHb7hJ4RBoB2rFtU1dZKnLD3
OLOtSVaAHOe7PSurAgijN6CoIaa+/eQW6Q1ctAmaKiqKyGUUOkQ7exQ4ygar0ltr
L2e6N7N0s6QT4jWGiFwNg3wQiSrqF24XKYXkk9Occ5neO7gFGEBwhx71rnS7eAdW
FS1EbiXcrcz6UO46P3gW3Hix3FYjbl5WduAK6oabYJaarMcj2NQ5tiNsNlBHlXKu
X5/r1N+dAtAmPPE7K2UCX/vcNwlRuzNFl5TjBT4ObbnsplIVK/E0KSI2ms1nY/lM
2Otx8+ryXfM4KAqNyVnSEJspYI2sYBDMel7qOLg1zhIM/3ul2TzrovBJZVxkQfbY
ntZwA1j0u7CKnyEgWYRXnrNsW9rMsiLzUoq0dL0tcYAeAplzSOQ9s7VwO1UIT4bb
S8nln0QGQ4m6Ll4hYTHpH4bLSi/G8aT2VPuVtMI9gJ6J1tJrk7iO2tjS4Ke4q/lu
lOAJPl9BdmFPAgXDWccOedP8D4Om3WV+D6/HpQZlOgS6RF1xYae8K6SpGWx17u7g
VJryPr6A8FoH/q7xtq9Ut3ScyqiWQmii8p8rHjIwU+aowtiI7dEvsMM5yIdgKlzM
Bwbw0fPrcLlWAswKM+EioLsroh2vPw1uudxjNM3pus/Fx2PSmL618iD8rnNGcoko
7omKzd4G/T1FtUKufelFbpcKkvVEYSKsPabdkwPNrpZifJmQthyC+7+TzL4STg/y
uooSHbZ1xfaCGJMvx0rAETw1KSHYdQo136haOsz6nkMNS/kRkkJ4BcdD09eCzuJy
wrVbmDw2HZM+mh9oRkbt0Ntce1FHVONsLvdxjFsfbS6W8Zd2CfHFnUmib5iJK8NA
xn2LPwKS1636IduGfTQiB6dtuZKN1SJPmu5/zPY4RyznBJ2mTqFbZ3J3J+0YugIc
wvZC7b0zqzvGi5y9yU3vsB3XWyr8+KKhbxhMcigKYgIpKfMRGg9bVAcXWBi8RIhr
MIje1AtwhZxRmERJPGt/qgJnsP15ya78j2Vpi2Jmxpb3zBm718VJalxenssVR11u
Zx2MacGqeqkAZz3nRwhzuVpcfgoFkpxYu1fEospiuAN1ets5gAeL4dj5J7W3qj/y
GEIDXnb6O3PA/2mgfmCaf75njoUi3A6alMGtlJ804cF4oLlWt72I1EsETr2nPEol
SK4bzq8NsuK25+hLHQqIvX8zpChRNgdcMTYMtJpqk7Z2wbotsh538R861bMQswYh
lZAm5GoghTHGVhfYJw14tQy/AKPdBEIyM/InExkMQ4oAgTwI0JaWCJ5lDY9mqk8E
yK6tJsnSWWsbz0rr3sUCV59oPaSc4dBruFpzLm/Ze6XLek0p83OPqySCGU1KwTVT
M7a7z3H+LSPVYa+cf/m2ALZCPln+3twZjkFxAVLjx3qJjknb0OZXE9fZoAacG2Pt
eFJzWmDtgUCIJFm0rGJWLEpw0Nf3FwVOBlPVqCJRtwuAR0os1GNHHJOLcwsUmyIW
muJuEGD8QEJ3EuWXOGdPulD0PuQfJEK6vK6W+yhVkon5uv3MBdEdWU1Hz0VfBWSF
UNGongS16C5Tpo6/XNsFCQPSl0ysnb5Ytam6XlIpE8+mxXDh0C/rEmXcMtmskqoH
i+MRib8N2FeNbdz1Kdvgckf4WkSfzFDxXtmh2tu5vbf3cFR9njmqOzku0W8s47a5
GUrk/m+CRlOuLr21phQKx8k6y8K+pNq12xZJzDuyu6SAS2tnlTJbqOUXu209QGXC
GxP580URidsML8IfdHZClIp7CGJNiA98Fb6KrR3rloxoHON7gKrmQrpPClip+PeX
R2k15dnUxyvAlGfSq1Sz/wBmWEMhQdNndk67CCxJnLMlruo84AgEVHrVs7wANwRo
Fl6zhm5s2TSrd5j6uYySkvQTeiGFUBHUIXhyoTNYGsCZZf92UFlK3tYgbVQ3HMXf
pLbOYCccwO6FdqcJVIdejtBAIahxJgFmQjsU3T2j+ltddPmEZabqHiMV8nw5KL44
uUdKirVSlnJbrMDY4pS/DAnapRJFyicIttNyARvtlMcPy64ujK33/PXsKT9UnaiL
suMYuX2EYC8E022y5bvma+0s01Dh4datOheM7NX5nVEPIzU4ljpBDteAaW2MeBHJ
MgmtsPwvNeHkAHUb9Ry00yEeyzxxwc8WS1b0XIPLh9WmKe/JIm2PTdf7ZoOJGFNX
21qie9O7vwuY3zpiANsYPTFI2LFSUNOI5dkso9stFheqT9mhu3Xk7Dzls0/Pzarr
Y0B0MexxEAjiXdPxGajlVg138MG6gnehcWo3MrdhECx/+L0fDheQ7zeJbjTyX+f5
BZoDnbO7pcQ+PNZZXlpsZV9rdRYhReKNgX5+2+P+uWhKohLgT+DqyBTOzrZLiwUH
Ki5O+LIzNHYJpbclX4+x0GSYHQSZTjfU0zzBpIDaRgchfS5Ii1yOz66b+JHuXr9b
b5fmBkbElca7KHNQWCQevCrYuLVpstPj7wd7UhwoXWjNviCWb8NJ+umBg53oTLAd
1q6QFPZ9F4Yf+DkE5dkM66gvBVapHy5kjihkqB1vtYt5LAkKEcsjwEJ0sQFwvGsK
htX6Gh7HnzRRWrnp4dGG9p2XVDTkXaaHk1Y/7Vyn+lckegSTxYECUo+Cx/gpiXWK
2KkcakUXyGaAyEG9L6FTK4ElB2ELEjdZJzzzYB2PRkf/ruHGYSRFozz9tfB8YYa/
bzojfxumdTY68UUJevZL9hQqo+Z5zx+TWwOoabLywOy4DJmfo8CcdPh8/1REMjvo
R6xktqvtVTA6jEexa/zxLWKjdTYGgHz0+ksEEpY5duRyhypSA7ChT0aSIUo18P4S
ZUPCpxRDpGdZelJ+INPtrGt83l+V8JRBpcJqUVK2s9KpaHU0DaFbJX0uwJkb578A
MVVko17DqVeQHpnXK4nbHqyr9ev+YszPSt5tcdEChkw9YgBnZtkPlz2qVf+AagCx
Nb5d6D66RZL7cDLlTwAcquMf8RPx6g49/u8yomSRsYhBuEyGRVBdLmFf/IjM++kw
zEkt8BHmZXPGWlrpkHXii8ehh9mWyGREwlJ9SmoXHDqhrzyZQggrJILoKE8F9nMG
juqGNqc6lX72sTpPbQvxja0Id02uE9JFJ7FSld3yreFGp5ALO7ua/h7fJaNDSjiD
VOtBpHP4hjqSW5ZOFhKlWooRG0y6iQg3AZMDb5bJwHEFHRPxUv/VitMp9kGkg1Fi
MfEVOKUISaRCV3yBjvQ1gm5eC5qo6pd43/SOcTgaF/vYmwWsgeCm1wvAkIHeMhiM
SguTnpPXYKnl8DeCM/tLeXSwxWXY/r0zSBElPpqt8e0P0JGZbYW6k/QM/r7LuKYD
9dfkrxDHnDU27iGaxjZKuUCeWfyB7iMkBpINYQz6Pk8hHRQEicxtLQCXQO0sm3UI
7eIF18/sr7GQ3jsUJ3rchZLuzhPhV4uzRqkVjslKUTsNm/baC7rp7KefgXyJhLf3
HDU9/re/v+pivtZvoDLYuHOmB/p/XoUorB6MgPRpFQYelnJQOncJlm//Pn9Lthmy
xNETwmF5egbgNodkWjO3006gOul9D+MKXcDyaxuMA42SXEuccAx8iVm96q/jQ8nX
svXM1iWPDs3Wjo3fQYe4nLvkCQfE0iHbtHQw3RUf11DrX9ETgrazvcVsnrx/UrS4
UzDHtnduQ4aiLcBKYKRA46h+VyqKhIIdW6Kbc8GL/cqpGGBdy47tXftnrVU7vlyW
xHjFzftujEZjMMXTitPMti1oJ2IqJGdLutNvHXD2/TIeOOvxTqHuwlEUBmTeVfoh
qu4VV6cuIh38oRuhP2epnuV38cV8oMaycwPacH3sPzIiv8XotWOWvYX6WFjnHMxL
GnloLk1RyPfl5TAEDcRYQvbyNDd523u6DMExUnkASAqKJ7PhN9czm0YpzWPlepFv
x4QyfdteSgwuyK9PNF41jGZwwzUCsUFRKSS0gBmIxj3IEqkMSuxoglKaV+ua84Cg
QOwXd4eEU3TLWU3r76CgcwbifbWRZ065UiEv7Yn/ayeBCZeS/4PmJ02lQ6nMSyDw
BqAmnbu6KNoAcb+D4EenS1lu52ExI3xct4Jsl7IgBcI2Psq8SBdiU6kmVkrN62xw
fKIdSazi7lAkBdCPPzG/KWSLcyCOg06BxeL7SWh0SEm2w2KXjcJBFExFDTApckAI
5HyDD/HIzCQ/nhtTeVxPNoAbZjEhtBPvolqyzCCrQjKmnkvdvnygTl/nz4CWBGb4
jftE0EjE8YLvlYZ45RQ+lz7/LX4LLn2vdCy/5AxsKbuUM/BBrVVf7Rm4CVPisOLc
mX7sWg4rlbC7LlvblG7sP5NEzOW2fX4wfvQXTh1XUvNDpS9HbxPEu7SFjIooe8tC
qfu69/oPx825msxCPgBlGyrXRa+imeXBhhUSSN6B1ig=
`pragma protect end_protected
