// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ggQpt5LTxRT/oh8rO1TrAxGgz/zJ/DUIjvOD0Ot6OWWwe3IZGIMAlBW57tXxRbaL
lqjhlS4pV3EFwdEN/OcxV1I8qL0apgeqRwQXz+O7Khg03wEWkJJhgcrkNF+VdciF
lodxVBZ28fd+OUp5JpH5Gmu889KzZe4+AFTUlg81RdM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43968)
Md2e6sn6FUhQxBn4vqyAachv07p6j3M+93HOhVLwZM9Z3cFBGJNnMCyBmF6Qnn4S
dPgexlE6jLc506zHnAPkoilrl2fFtZcPCsTxcObm2SQ1/M2lBRvCjw3dFusVpR8W
G+OWozBt3TnSbME9C22kWGbBIrPPunKYA6rdeIP4qVAnrKMllcl/GtiO+i9TJKeo
O718QpCnSiFJEKECjpUpULpPGZ2G2J+bU8L1mf/FyeEzGVowsOh4OU+OtcSoDbES
vxqBN/KRo8S+k+2i2ciMvHy3pWZlO25i8SRftQOkMZv5aoOl1p57TxE17QLDI6r/
qmkKoMKCqpPCcskAaXGg8S9F6NYYr83KAV3zMXllTipQbNqWg/E0opjHBOf5OGZN
yFIIFj1rwIAasYu4WExlfI/DVRsNQMQOVC0pZ7PKhLnWYixZfClzw6/U/0YrdurU
5lTffQOXOfdeRY1fHpvLsxSHCKegWL8k/bxCqme4JTjHvHVkNDIb2P7uQka/zYQz
1tz2fiYE3DkERpTV3MUCRVh/QaedvLhJZHrD2+VVF9TLnlMhD/MY6SBVbkp1BzgC
rq0lDeDBjCTM/Zb8egyNtp7WK7wrIuhuVewCCGowbU7DA47KxZZDbIahoT4gxLpQ
um3N9X8PYnI8CULKLo25cAEJnIL4WrNDW5K73EGDG6dW7ndFx+92bEQKCeBzta3j
Jq2phewS0BGI4zgqKJe0fPVeqHkv+6cWxVMonLm80T9dpts9chQtk6d/twOWGPtV
UzFLuvaYSFLDGdwhrCi2blnUQGjoeihTNHypAIPDfc478pi9w6EqJzznRqjK9Mac
DZ+QRaebP6XNRPQKQReNxW3NtswZ5bNTFCcOaDY19mJl+T3ezbANzbfRXlz7ze8w
Y+HyirFzKlG2iOM85TWCeSRUnAfO+l9P8HehvBivJLnLaUbFnM//Sg3BNTZdpDsl
tsHnn2N05emmHfLyPLcZ9yNWxNBuFiW28UZuP8q0T6qug8t5dhNabkZw0OOryE2R
JP8wWcWbuck5eZ5Ign02ijC+vBB2VKeZr+T2cQ5b4OXDBDff4YRb6sJBGZ9NEiz9
sYCtw5j/6ZHKotFOaZ9SFTZVi1n5pT8gXVQP5SW3sP39vaDDzb89WFI0cNYsMuBZ
USenCr1ScPtZF8TXAFEL8/vN+fQuMq2PeKB+W7nU/8OlIzaBLutjfbLTiflR5JB1
2JlH1Nv5QJaPc/eNNjfXWh6mrL3K9VEPRt3pe4qjTrLro0Vveltzmi1gUkNHWUgj
h5wTSHOeI41Jw82Ly4furYR9PFjb+tie4s+mlnFPl+pRaDqN0BXG7eH06OtoPg+v
PXeaBog6WGAVw4Qu3mGK03qRDf1SFhurmBD630Bg8QKcYTYY/VW9WY+2qfo+supK
MZH202ptA69h144zX7TXQH/RHEuElB/Jf2s8SVAz7X+zfeEm0OD4z5VFlIXy/FxA
tUfZgrdCmcazIHOF964YRAmVzziS/4tTi89oGCq19nlwv69kUooSR5hD/Ph4YN2e
guifhrHrEOpdSctnjztfWekJELSVJV8OQHdv0EJoOsitlSta9EklqPEkuZNvd/lj
RhX/DU/s9qiCY/m7z4rEFcAYzuFR2zQyHY/xoVs1cttZGGRtJPuz1sYXx2WUUgJX
b7600futt7EC3RilGvj9xJwbP+zIaqzLNf79yCuYPDHrBc8qqbO6D2ai/mS70VR5
/GhNy8O2S1ADxGFZXIW9z95LKFRtUv09QVeykRC7YEuKy2ptEeL/Z0XSy34BYkK9
65t5IuQ0InHz+4oWnXQ9seJ3BBazx+GQZMTxpqNaEf2DD4f9mhjZv2SjX4vgpTIa
r+dWPfrQmNIHIQf0yeU7APyfDkJ0ZvezGVyTXdF5bh2y+18zq1cUbaiqxt7tM31Q
pB+GayOCbBzv/wh9483wRyf7HAseIgKF+LY10m9JQoJ4e+ER1Ef2LtwuZxCm19jr
/2cUm5ikjoBa4zC9ZGvlFY6ylDa7mXZAMkANIiSbjMI4RXt9N4mDBnzYU5PQHpui
puyU0PWfZoD5toXZYLmGNewynJIqlwAOSk443BGUW5ulhurEBgQ+jS5QqWeTv+uS
OAHuv9ksVfknpFmQeaxvtn2aKIq4xBYzr+m8zM2+KqkdF2HVtkbSSPgEekEcdIOy
oyuiPx5aXpiuyBpc47Dni42+ihgu9d104HXjOoLSnd5FiJdyfUHRH1OLh8LwrNi2
2YZo8i1qXf/ebtooOmO/JDlzPFAa+dwVL4BQqPi/vwSo43pygGiQC2oyCTMdj4e+
SbldosCtoc9tKAYtmFOr4ksHT7BxLH1X0ChwKHD9E/AyoJsdEESqtdvFTt+1G8In
erRjRY1EjCiGzojb8n9t9HLEk+++av35Orj8hf/f846/5IfSPq7tp8nIGW7J4Hou
4fnPbktPacwhYs3DdWKaUe2fzr4Cz6beyK7X5Dphq2dlMBrI0mN7hqc3FTjhstPj
ays3rzNljb1amFim/FDslNOYgRB+yAk5AqG7bmj8We/UaKgo/LO83wZR7Vk0qw0R
kg/CDE9X2ky9dae31r2IGyxNBpIqsroyelDKj/XhnG5oHo6L54pomU5cnHv2x/vQ
5nEoNLR9ZGzh85rm5G75Sw8TyUzWc7/gcD2d2u01L+kQGfH6WmWWz0BgyuDzWIll
bRvtIvgHzD0SnmkcO7uYHsPERkhBLN7ievRktOaJ+GKJHnkGifU7VWfN0QZOk/DC
Ovd8j+UclZuR3m5ZtgdDe4TFlprk528gF7/1ifCTynGI6WpSNEdqE4dAsM0GzPiQ
1P0J4GzFCdc9Rx29saGgVuSTufdz+8DwYFbycwNasfghGVqP9pKh65x95ohDqBCU
laK9m827Fa3k494CpB9qe5J8X63jXIaq6TK+LvbBFouQhRr7zbd/gXdTEW3vExmn
Gtqqs9F/6gc1aXePh1sDaFMHOkYJG+gho38EJkTId4slp2edGX6Yy5ag5oao1/fa
e+34iae2lntp7QIwGWL8miobtj00WqeCZ337itdbzf7gNMWTPHk9W9QhCXB5tioF
iWIiO2DImKPcNwPNVG/HtBcByNKse3PtRDgcox33k6OtE4K+fkfGFqVA+MG9xzuD
j6YsgXmGCFUVnCF3lJg9P2zKlsSWPvdmHRQzzn4SZhCxCGIyBHCwWoDVUNgBFlR4
ZA6k9jybq71WgQgeWEl/Z/On25sDh8wDn+/LNNfzw6MEgxg0Ul+plc62gCMm7x6q
IVdKM8BEwGk+omKiyetRQfM+SUUWASdDKj1ANYgd9Le/ikpZhvtfISOJM9iVDtWT
UgUXkMo1n67DPAhJygKlPQqP3OBbdde9jYgA2Ztc1R+SI+FAeChIpHJCkliIROA8
Znt8sFJSBSyCl+RUuRQ/NfAxqncuV5eJA11cJLDYlS92YucmwyJIooU4w5KFRUBm
oJH50zuh1XDsZHvB+jqAKW89ORo+hmSQ1w9TXvpABE1XLZsvpWu3uj2GgFRFMawA
ZkfjIS/0QMy8GlyaN3MKRmHcGgqHG1qJsAhuGdNQFMtJoIv7fL3GcbGb6mILjwut
jKJfjrlWRNz9iSICwiHFjGTUona3zwWu5AcuIiiq+Bg44yMW8ngPCFMuJOdsVgwo
jrsu0noUfaDFrmXX0XbpBUFHCxCNxHGhZmYlA9/MtxOpuM1t2uD9Q9CDnuO0MJBx
Axx76Em0ZvSLwRj4fI3bRiYD5ITHCjg6f5a6/ZcSnbpt93qJup7o4k9PrviPlfdU
+5hrp5xRRHHJZo/tPbKybZndcPavFV0kEJudKOOBhIGYjrsyzpR0AvMPkdlrzwaf
iZgt4v3njqS7E9JRjVnY6sDBFDCnIFUDVY4UfVTWhu8eNXutxLYeJy+Ki3Bx6ex5
gZmIoKAsPe1Fr94qQzA8VwEvOW3Ekqz6s7oD8q2FyhJ2hlvOIuamNbQ0XSiAdbcZ
10ltqst+S3JsHod5KJ2LqSs2ca++XrvnMbOkcTQjgh2LSobzlkzzU8+fc2Vt+MUI
NAA5of7fyyg+NGvRrI0krvwGvMDbRLDlPEBDq8l3DpMtJO68oKyuAvU1ISX61q2e
62n/fUv8eZ4dMAkHK9rlOlVBeEXiyVIsefAXUYZayLCpj69uKmYyzs0kYP1YutZu
usc80eckTN3P+kIZ1Mj2W5SQwgKolRGoQensubm5xQbtzhCCm1kjLofA+1YRLa5W
f3lsQzGXfcDMuokUVaFf2v5x25mjNq1Pu6kDIamvtXBG4PTgm08oKChRHvdJz5IF
pNfYIhWf+PL7QW7lJBdSAXdeXv9JzX2QXu6DCDAwGC5dmSRYCi3MWHMrJKCYmbj7
dpxEUjmUr2dGGDaBaNbNyGMKd8MABj648cNZbi7GX2whFjgix83ijzDjkiZj9FJA
2fhnwyEjRjCrHIXG/tVBbYUDWy154O5BylOyebvQmUK129iZvhXVMZsYrjP2KF2d
cTajNelw+0C4zxG/ZL30zoRUUcGGSRrdS9EecPOR0wBbGksKmvyuIxgKGpf1mSQJ
B49soJkhaGW6pYTsPpxNY1KQtw3lk8E1gufEtlGBFnoUmPQ3KbCQBMGP1ac/Yl/l
RpOxAq84oD5fz6rrTVw1TEFhe0dh7TFF3i1zO6FY1HnbkImHjrN1tjg6ml7leTkk
4jgkIV7U64bkmgDvE1MZTyItD87W5f1VS+DZBSUG2pa9L5fA+Zj0sJwWKlUNIIYB
9sESx7HEPfZR28y5QYOm+3s1QzwLAUSSoUoy8v6B5HMLGApZ2P/dGCnDo+hGviMP
kM35+YtPK0OguYiH1jzX19weHcOOzQ/wgKZ6+PxoS48Mp+72EP5XL/GL6skx9/Gn
eJD/HacAzMuLxrzswb/WxCDOHoivIetlFnXg1lCfghpJZeFcVhSoy5pYlb7qT9gT
MRhue2HPzcLeLmCXXaEWtcjkUfbVMavaQM7xY3908lItRSdUQbaj2pc/BPZD0rl+
9lgEOXZWJdMmXoTJMGOkpeozlenZZKp0dTlDMSQQ5WTtkuu9Wy9/AVDEDrqXStC0
CktRnkHtHCRAemJzK02E4T5J+JFi22vJLBXGqEQobKkLdTzkVkqQZmcH5yY4e3Ze
hirDW135dv+eJ77nti9xYoawIiv4vggfgwA+txenm2EF1M4HYuyeuIpcFW5Bd/LX
7WOh7UjNMBtd3odfEL6Th61z9vej64gwNv6l1rS49R8y1l/6zURzz92FSrWdQgJp
653pFOlFJIU3DNVzCvnCNMPAOfDDGq/8+//7Rbm6Jb1+dw7m6y12cM4dtWjzeu15
T2qtlYASWDg50RRjVX8D4tCSi+dzduIULf0CvBb/1ALN0p9b2tUJOnrWcY8cw5I3
EVIbCXwVp6fUWFKzqIGBQBg5jCW6nyY7F81PMgizfPSMQozxc7GOGdFrFExvHNNw
FmmJmhL9dgAAmiQqGCTnoHiMz5mrL+aWgp9PLjj3Z1X+j7Lt/U+9b7ODVr0dx/ke
s1Pq7vrPhJuWw2q5UPbVjs+JGa4O8sVumyAA0jekijEqjA6XUg1lO0ZjTrP3NYwo
52PvxOo2C4TU361vV+08RiChFB3ogitpHI7XeTqYvDk0y7R0yKcCtOau2dCwPHgD
CkAprlpyktBEXEY19xPek2ROeuOE0Fxaw7AizaknMPdDS1K4iQy/kLdXlLtHibii
bcUXlBADpbGVnNz+K+Ktx4SFNW0jOzgOXrBUpZz930zLpRBdQYiznSjMUoKNb4C3
+A5blr8K81+U3zWcW6GC2/jjtYmfeqxbDng1bFFqSo3dmPdoTUo/+f7EXAJxuNfv
e5c0/11ArOXmcR1dbn2p/ngqfSyJ/5PT+rHuImL+a7XmYAVYVrb9GCjAUKnf13kI
eWu0JZDLVwXoF0lT4n5BCdXD2eKtLivx+/TZEXSx+6fA43UrGfCYREKUGK0N14Er
r4jfcSEFgCmGGI8kZ/Z7/0p8c483qMIe5AiLAU4cqXnLkmq+XBwSd0PnrcyeKCEX
n9yfFoFhpsIy48MIrkMezhS468lOyPo+C/TKbZwVo2kJrrZV4UKEbX+VGO5/YzER
UEeGNvbcP8Xjv1qUSUly7MDeBGeZje2vzT4kXnKnSV3hPATkAnCAE145RO8N6QZx
jV+Jyuhc/ZqapnN8sPYEFt6BCnOTJRYU/WLVo6HSXKvrhHjlUldGfwVt8zGnuNrI
niIvvDYvedLpV0Y8m5jggfafXP0shEOBR/SSDriQ6iA7VjGrni0wEGXZiOrixY6K
Xktg2qOy19pxEhPTYW0ptogologny7i65jJc6G5v+55u28fJo1tNd2s7K3W7rjBq
SlXWzZqLyyZ07gLgVCplfm7GMEBJbUTVInwiGstxRQRf1Do+CJWBF/iKWwIlkWvq
Zg/jHh6fEC/G2sPxrAxsuIDtgkHubtVGcjvutqahCeyKfRw9cbZU7DURw74UBqRM
eBmiRMrQjH+SUOV3Oc2XLMJsPWQGoIaqhtLKCDO93H8Vmo3YYtog7N4HMHnvDaDU
K5sllqWIUZSQXwCL9id7FWF5igMImj8MsX+0X0hRe/ziJgXybrLedK1gTAv21l8P
OxqHhoV0EuuKdKYGd3choFFtCyLPxOO/wp0w9nk+J9HwBLd7t5QCiNbetMp5YNuw
qKbvGwYy3kOmzrdpDpKHO+li50YOXkTXF0KkM4JN1lF5l0K/vogO/nqY9EkPXmKf
+TG3e1FZ4AeAKtpcHzJmIBX/XhPzGIHTREbaj2/m7HG8vDIB3aTuRtXom7InpiSZ
U6wmRkfCkz3E2SHNAIGiL5lORdTzzYKX6EYwxnO4uZqoQa6MJmfW5U4ONO+s7TwE
Iin0hNlD9s2O+YwiaqB4AY9UIJoXNr0ANxx082RXBSCeUd6tjET2IcavaGPe7cTa
h48LsvvJnY/JBSgP2OMkL2VYks11qoLRo3sBFwoBybXVEopcrs2WrkQO3LEYBeKn
684RkdaZr8z0yXD7ErEwIfKOjGAO4ufvTca580XXXfLWQgtxKTX8DQmH0ngBoEAr
x1cOBMpQYz7K2jRKgDrrXERrr8h1oZw6GR+JLLYYmS5gp6DboE1nxqWe0QCLkZs4
7w6eeXcVlSh8oFbEtl/p09XlMv0F26vQoQ+zTnSYWf1V+1PT9CkJ/I1rwhtrzFOU
9ThlNIQz4r0H9RAjHjaUd3YR80r2OZWAvZ3Xo98h+LucCoTc5pzO97Nfl6kotsKi
+L70cDN5CXQLIM3Cm/IcmpZuwUz88XGZgHe+kA2MYaQ5IidFycsZ84Tjh7pGIBvP
F3Wvln4c9hSmi1Z2zy6zyQGxcHKbvU7kzS+fbXDC7/Wa/x9yZ+/9rky/MjDticZx
lqq3ZaT/9m2VUq3YTAVimtBTgE/SQ7RLQE5HqUp5/QyXz+u0zPAMQvkn6KNtIuRp
ZE/hxutQppL5YDwISu9HJPvKfdVL9Qz+qb1NM1WXCuUr40DuWRiM6J5zEJNnLw2K
zQpyAKAq0byEq3TyYuNv3HB5UiRHsUqm59ucXI5ohNRkjW6Jo1cRJfPL885YKzHf
xzH24/VjU0kN1ZmNz+PJZyB8VYWT5rvXhRHbe9llXlAlb676Ety+Jyg24Fc4jZ/g
uU6oKJLDu+5OxmER/idHElXSlWJKejLt2sW10aMUOs4pWEo1P6GRMzwVPpJVPlWb
dAzzVYyimoJ6bXEnqI3HDpTdHJ/eI9VM0koghyOq1+uGzEV2+QU4CY/+qqLAiTcs
m0tDyqirfbhVLGoJICz3rniwrzacvPT9PaZRFyXXwWirqfyPytt2zO+eDdbQgOdV
oR7Y7QlQkiZHZx4YqcYqeU+4bs7proFC8rUxqPd67O4gGymywfx8v+9+kAYrBhfF
zxQ+doYt911WuMXIyfc4y/MryyT3Q9k5H4voPl+KsI4Bw+LWhTRNRMl2DyB5Qjtp
R9JIxd/B80W6xQh8YuZSSocV7LBpT16YxITx8A326iUt6wOpFm6G8D0gjZymlF20
ulnoY7XOBLOue1v+NZvl3myrFbOs0bA2nvCkb7HQgwRj6Wgx+dIr2r8z29E1xjrw
TI7FU86klxnD5koRlW/AKNncmpZfFWp0XUg9I7PzsGIbXH5PXpBYJL6KYPgtbNnJ
HAqr9nPLteNtnfpcKGCX7jRFbqCsZOHystrCT96TtiqkGy1iAd5SXO+iqtHMyDrW
WlfGQczZWI7QLmr3Gt4MYJCzvq8X1hqPZaIIcptiEx3EAX9GWFq0+ZfmbNIPW0JO
mggR7h+FdNMs9TvpUEhZNzG2ZcL1W+cSl1+WTQ557VEKY1+tKAgfd1GPzROMldXa
+tk8stj6s/pLKl70djXLqHL/z3WmoHkRvlnDVRDCL+qMdcC7LPvLN9ejmxZpoYHJ
T1T+MEnK2chAhkwzc2Owg6ZLNVZgpcR4WAAqGPcQRqEva5gpP3LHG+eigcIaS5/0
45cv3jnIR0nj2gkt8yLMSjdPlLV30SVpprVizT60SkSmMRWpZ2AfpAaSijafqEg/
AzNJ3Lim3tZj2OD5EZrA9UqHg1X8jZJz1XRxjC2gq0i6psJQGgJJPDxMPMoWg7Sk
DUs8+Ez24NX+tfyxm5eNo+nAO8ASQyVCsxNe/AZgNbueewoLesBGsuxrgrXXfdC9
z99mSx6zlL9TR/KzrD2ENwSrixjEsQGeIG+r3GFTCidy+7EsjTq0CU/KnB4vl6TY
m4g6liJkE/LEJilv/aNc7eZtqWPHBD9Y0U7PCFhXNoZbd/uPb7+4fI0qhREXDG0E
6h39mLz5ytJukjcgKZx0an9vNjvM2eQIpJenqOMDl3B3QhzXa379JrkpwaN3I6Ei
QrfbnNHK+6fDHULzISshzsRWL+De39iepSaMBfBMI40SCOGQyOxOALgOnxPuaCKI
1r2hQQ82F4amgXiT2D/1drCOsb6/5buZEMG//+AT3v3onWB5LOfIgNowOYkUaZa7
PbWZFvE9k+XewX6yKULskvjs9mvMru0hg3/CHu2NODqgib2/vkMiaHCpfHhhREnI
oW+IEMjQnsR4H9VlQJOohe9hphGvRfoVNhtwVKZalQxq6igy8KUGix3v/WBK4IGd
/nnmB9TG56lGRLAlsBq4G0f1jSZje55UneI5u0oDqBNkKcDnti3sHJrhCS48lsLm
wqED/lXEvNfh5qmc2uFuJ37CuLsIV692nKmsslgd4NhzVZ/blRrld5k1g/4Nw3gl
v2NLovvHyxXjwP0upSeoB5v65Kqvq/MI2EJB4O0OZIvjZsS7kRVYjruHYA22xQzQ
pvkXnLOuAgV0NNPKezO9VxR6m1033cSu7hvmLx6DbfwkSH8NapiW7Y8s9F5xNZO5
nVvnDRumENEgM3I6xxITvka6WuWPqsISzvqZFIrNp/dxRKEQf/nRT4Je3VpB73/F
onXrfGvCfRXey8rFyZdq1Zly/NqPcmwmS0/8BCgOyDTlqMS/poAKgcdMf6q2Dalc
uSM7BWDfcFaaygzS1VEjsDZ2BR9mngLpiD7Om0dI6bSZwdZIYUVbga2FXd94IPnZ
u7NBndeX3+4rQYeyLhm9KO7Pq6odeP9Wock2QZaW3DPNo8VKLFL9F+UKQ5lNFicS
m4rWXBJWpWogH1iKL3da+6/sa7I+H1Usj7GQMYApU5hfgHpcYHeRhI9HU8+pcEOc
I2su/DhbrMPKoCj2uS/JyX1+aUmyv8zpxR8ajS70FNwkI4iKaePUERBbLJGuWdOm
Svi9C2GsY3URr/8faxpSbN+COY7nhdMV1//jTmvNxur/P8oHsNg45U/Q/x+CRNRU
o46T6Zau+uvRTa+uQ2TZ+kScCp2yk8qBSNFHMMkhdKPP2gRHH7XRufOp43gWlhc6
poY5KZOFUxFJBl2H2rRDn990RgQhfGQSh7w0cJ/MWlM6KpK2rs6PxpdJd1N1Qwnw
+yPa0D7yIf4FHiGIVApiuwlgeAtiaDZTUR0Db+r+H/e71qWaIi7YNfcPYdux9O1a
911jD6GbJMsb4yS7H3I37GvHjVs7IeqEGbBHduxkWT2V5kUghpSovuI57wraX+tz
lyxqLFvA96xtLAV+8JWDdOhPAxS64CicudnvPtte9hZ3WxC6iFYG3Ywfc1SXgjyy
U1+BISEldcVguyid58Puy5OB306bwnU0Wy1FG12jIC2GnFV9cM/si8wBsCvPUif5
qh+g8i3UP3I8YTcOIcSTrZEnQ2HOOeMQzTESOzHHeSTCbtOTmpGOn1sk4lWs5S8t
O48PbV4NtcavPqz4TqMAcV13DNm8JNMwTktTttGOH1lssE/ZyI+b4usgYq0UYyz4
G4YotxOAgPda/Gzs3UgupigDYpEjCsO10qKdBb40NkranwQqmA2ucr6eo+1xRly/
I3Hl9yUbuegdCz20sRLpl5ZxEblKMzJPVwxU/b9EyqaTUlul30uGIYV5PSarCmqX
ZGzXPKca+at9KP9RyEe6vG1r1B1vOOh+P5EZeU2kZ/RksaaOaMl8eQMuxcwPGtxC
IHCIaah/2sfjmhqblm7/hukN6DjEd3df4ARLTG6rrrLDybKnFD4laAcJ2w1Z6Fb7
sZ0TQcvz0oFbtp6NEpShftxxbLm0hJ5/SMJrUT2IqqTl3F876jxZ+vHYnJVOHTin
MzZudGHNN1t985tsELtgK2zmJkioyJ31GC8hCvpJEY+E9IASMxtn40JvpF1iFLk/
Djz6geXlZaYNJlVmOuMo1l4RJ+3X91jHJum53k+dfP1b4x+TrXBxv5Vi0g+CM7cg
A0Umv12lId9BlWrwQP73RKty/B/nW9SdGsUcKMpRv1ogliIwMpOevIhQziw4NI3E
VtQlOU8PoTa38lOwqRPlPeXvN+lnYm8nHUMd0vUcbyyA0IvFVAOYM6k2Ie7YA7pL
K5RitCETf4Qz9NY++6RLtc8l6xqqNuq8WDdWqCfzIeX67w2yr/QcsLvXhSaaGNIm
xIjQPEh7KUio+ZaBgDEXJ/fIYooGEs2feyN5g0zXmmSQcLm4xn+ASeCJumbRRgx7
WAJiQoRI9pfMb4pTHi0EICbFp8Qc2Tjh7iFQbCaPr3BPn3r3HcYBX5ojVSKN2gvv
8pvRQFyU2r86koUslZQIzJFfzi3zH0K8p+2GD78kKf+LQiwxlNJydmD4muGhOjYA
Wa4j3K1IrjCfFtxUpmTwP/fE8v7N0Hr8iE9FozEa+amSlpVYg+07TU8GF5izJyRS
YprpSKVc5iD3p7YK0oSJ0nAhPX7RaG+JrG0iSb+yc6MG6ahuNmfkV+53tnKbx73D
n9gmaH0hqe/mGVJXfkoqmb5o8cJSUpAus0kBLvpOWFfKrKzR+oc64JQ4tTb1RU0B
oV+sksFzFzOGpfqFiBdgLxHNQ8MCXVcnR9nHvnElr/lXCUwochRhg3U5T6fxHClJ
fU0w1ZAQIvG+0XwXt+7NQR+IvwZFu0XXGvgUHgUSr6o5of8Gkvyc6YurkK89Y5PZ
HqWdOj5KMQWW5lhyCOLtXOKa9lwVo7OKiwnEu8oXSGzcHDv8HRbqGalHce8/azPa
5AtWYlbkHDPbE6zSVooFOMzNhcsB6Goi25d6IZQEt7MwktnyKn6ZZdB26DJhV4Cx
L6CRRHllvIlCRepKckEh4CuqOeahh3f1JN1V/KMuSnLVx8OM2MQXsUkdC60jX69J
UlV3ghtGA8iW3OwO3uVaD8a3FtZW9VbEXjlsI6BBav5Lrxpsv6Vx1yijJpjEIfTt
4QN1i94A0RYPfoA/acNvaojV2m3LSRX731VOdGkzR6Jix4PgpLJVUgk/CVuBtsjF
U5KT6y7liM8UWohPKMe3Yy04C0Z2dDtYylhl2XZJjxMa/tuTdmuHpQ0nTyrczMcZ
IlbpwhN3PwRa2tGotrAhLY7eutQyFRLDHRkj15Je8zedHyzeiQTEtrdqxVFaf/12
M3pXsviOIRQLafcOucBhi3XhtDfdvD3qAuI99z/y6YYKMg1+n9+7kOsFYsxNDipp
4pK0z59XNHKAohVrG1dyTB4/Hi02udyl9Jxk8vUe68h71UeEn48t7pMyoAouY6b3
V+kpGkdPMELHeoId21C9A69tlqHRZtFwVliHqe7GcGH9rkwt/BYV0Qsh1FB2j0CB
0Rh80FGxbzA90vlLBg2vEiXULV9cxCyb8lvk+qB4ywC8jrStXzXn0nBBh0WzFFdo
nkQy8NDsfZlr/VIBmMYxCPGczb71YR7BCny1N0apdgNTWE7jb51+O9NgmNy4heu4
RJ1GsvKCNqHWSdhWrcFfZWyh/RJUvfC4ugzo6mnNYL8DAhsWEZxq1jtZv4wLTm28
kG784eQMozZCJICkWib7/zkJ68M2/h/wmRoqTmmSfcxVzOc+rnJb+nsqnHyB55Uc
lFA/HoY0OxGm0iTL6vdlS6UwumLzNVwDBdQhE6XJCsY3coFTgzWUbTHwGW/fORPy
IzwAbfqx4SEHnQaju3MezPYXYJsEVEZ/4X1EhAe/XRPHcvkPnYC0yDrogvsNN2L5
szzuRRCXRCosn64zOz5mJo/Iu48iCmXLJ10ZFY5tDOINwc/2q462Yzxm/mqX6yVH
z8sqdn5NYhyaAN3wCINUhpTalUSluZUEypA7gwkkVE/3ZWSvFf/ASR28KKjWo8Sd
cZ1WOiCHSZNBvtklXCE8d6M46B8zEjf66plCSkpvLehKthfM9n4lGVeWqMInV7hk
SxoSjbQHtyqWTlOt6pwx5cW//xp2eAXDm1i7fIGAmLmOnGYihoElMx1TEXfjTEek
3GS/dC2zzPf0C4KzU5iqf015qpSkW03WqIr6mSuO3ouzu+xErpbHbwBRIwL3c19u
24HA8aFqR6pmhomaFxDh3FmafQv5dXyXcpvYh6Qhy0rfeQgnFcyFGhV2TS1ZYeix
90TaYHV3GB/BUs9ByUJmikom+thX6iR9g53qAg8ERIHy4fiMsSfFfoTF03IB0mBy
mYO+xymezUELBODwUA81eaj5Z45aMqU44XFjwaKm+UESWQmbi2gJmkS1uYLYOcm+
JQai2DDcC4wS9xjzRCuCrusXHM4kgAz3U0bqD8Z9zl/4y1c9gV/e5cpRMXVuVFto
syqhw5VA2hgDzVSdqDiyRhJhfPgF/NSPkFaRFXzjICR50Z1Pmw6FFeNaDgWbPC8D
fN8YtlE3Z1M9fXEf/jEuxuLlowFOjFcAJvwHWBuUAEAheQGq8QFt9nS0kIF7LSev
7Re9W+t5drD2sTmepRuxOEZjcezFacd9CQ3PaJo8N4NNumwnpeOdNwLCBU2ZHioW
A5sVTcouXKUby+hHQErugcHTnm+jyougnEIzz8E4gsgT2xg/Nka5X8bpvPTS+c6U
XhrP33eoHjFwfTecCDdG2B9VnRLvm7BsKj11dAvLb8mPzJr2DkEkip00MuSlOH2d
bhyc+lN9mPXxUtlQa+8yZj/OVF039P9QLQ+xww7igpYMV4HNiXjguVjuDM08cSkU
dlE2opTM3iuVV9w1+0E4EBcYzlsW8ipFtd3LVxJOpXzRrjYyjxEzjfyfnJaEDdlN
HJUoM0bjifVCLKWwr3eMD6fwpDckUmQ2tFY8nzqBx4BQnKiFJzqsGnpBNSFnLBRX
q2y12lLayptvzQKe7sTpOx7AmmNlI8IBFlhL253RdrTnCn+rzQj/xwXE//o3zA3K
GKfMP0ZHzN4fst6495FZ6QxgCGw8EMTIUTwiHDziRhniE2cpOB5OShOZwYO1tTMz
nAZc8KL2xMaB7Mmw3+AtITqvCzgevyzy6gMSadP4CmLv/HpNWsHfeNoU1SR7xQaR
/RqL2ep6ma8SI6iZ49oyqmD4qFzTES1Q2sqnjM65naEwUWiJOxiGAv+8m4Ew6QEy
SGGJJp2wH8jqg1a5hJkpJomZ14g2+wC7m8ktTrW6Bs/lyswb7fK95JJ/9iDbKNiG
kP2+l8Y4Nci74XY6TjbEPcvsLRT9+5ZAdoz9Oh3TtHN6xOpdoe74zo/QYD0MXecE
h1PoTEm8tE0rPiUQUkpzibU6UuvpXCuWiY4gf9/5zDIIeCUGY0L3qH5iJD+CWDMK
v3K0Z9zd2m2Lh7bT3yT8XCG2zfM9d0+DacLjqXppZ0GnX/eMjlT4mOShQT2Tdm+e
xqrduEX7E0uYh/0eWbMH2MrTTwIv2+aw18O2zRNE42BILvReJOExe6eKdza17Aql
UN0s0DgxvvaaQy5u/MM0SjWOZmFZUymI/fUU7Ta97gBMqbit9mUVLJYQddp8pWgM
ktfJia++WHMoXJax6W945ygMYGnvqVYu9Ft/bHCNh/YRCpcWgg/wrPYspmSjtCdQ
RcVIhYylYSKpKPAu/E85cHDHdKiJ0W+6wG+uII3EGstj2i8pyNUZPDLAw9b4gTNz
XH65g33dN2IkubA761rpLuArTZeM0sDqcrmTcD7igfzDsrZJE9HqY/BVXHnlAjiK
If7Na5V9S6Zt0zshwk40DwXba0oTZDr9PPtgnuMfgi/oUgAxOIswJsxdWfJfkFYw
7xessm6uFl5OkHNtkiS0/PzrEkbhyBgh1HHlf7REL7g2X6YuXlbUTAGBghw8bCOk
kkzCIrSdrjQjCAelPy2qYdAGV28ap9wRvVSW8tMh9/x/D+paBi+/N61FchkGyzCn
JetE2zgqqwgC97jN6CdQnmewQqvtME3XXylvbQQosVr9uIPGQ2mHNNUZ0LYZGxUV
45ueE7aqUPvAvQzhNaoxpGMCy+XxjBza43wKLX9F3Tm8ottoMJ89a6oPvbyXl1mQ
z6mjWHPJwKt+xA+b7C1L/b/+STqEN22D6pceaXTmXPe/ixGDNS+RTDcXlUTmExMA
DQVXKZsI0s/+y2c7jBKEiP0fnGe4bCPqhZHtuK1RKgiQiR6AOKE3mOtKMtIEKcZI
CEhrd53iTXInH2kctK3KOS2xGvT+hPKBvPYuZl1IBvom7eKXO6q7wjsyTO5fr4r9
PwjJNisvUmsDoYSD1SzipuGThpD+kmj+nW0RXdi7lEDdnlVkGMBLyH27jcSn8c8s
wVGj+QqHVIG3UtO5AGUy+UXvZvlIt4V/JdMww6mcI5pgyw8UvhLa4kdut8hWuIB/
kErFANwSxcIucxJvVD0s1/q7hX9rdqIAJOq4msHfteey+NfL6MsJwuZRS1bpxPqR
l8DPAySytE3nGnPJ9cVOv6+yZQwEBxKQtZWG/7RLoLt46nRnfK2PnCzvuJlttcsp
eEyXBj4+d7UTtMHr+slNwTc7OpzBeynyqg7f6ZU34BNotVd8Q/cE7ZeYYQSZY9dY
hWZihbwtAYyCTFoIlk/gPKj9pAiXBU0EouW+mpeHhoAjF+08ltCmfaPZjFJHuKXJ
y3XLADTG5bNQ//EXQ8/FITqoX6kkeYX/NXAIBp/LGdKrFONC+f8RgjBt9GTFvfvq
Hnr6nDmtO5VraKiaO2m8cpmXZxf1Ej8UJN3O0zWXu5BFcYEeAzTs6yMglYYMnlzX
tG/6D/e6+USJrxdNLQvbcvI8/c+5MV1NieYQPylUwW0+2zQ8L8ZVmZljnfOjVSWd
njUbSj30WvL8Yu8S9hebAnU0HwP1Qk0bktugsu5SLRqsd8rJcN0t4JPjQHgyzVJB
J9IiOZRBr9+yjxGJnBIDVWObyJ+FJLvxGt/jLlrHliDS4RJPP60v7f56B+MwNETB
jivxu64yuThwGzg+AzynAryQ5rJAMQPSz677Xxjlsx70lgpK5JFpDtdfNAWQ7fkO
MexdjjUqpz8Y1vXMrb+8fo1pGawCFC18dCf1xR7NGPSdWWqMsGjwuEw3kq8HCObe
atRM0JyFRgfC8k9GsXv0xOgxxu3DIBniy7k5t2MjS9CMxllaVkX56WBxK48cA6Co
Lwi3AEfbVXxYyNKKy7RSI8Q4j9vIthSd1k2sEYA/UhgLY6qZlxXYLyFvGkakK4pM
0FgX+bbqTJS/Z3fmyrY1/mEjj5MNyKBfivH3n2iKkLbLEuc9Fn1tfIGjEVI1Ztdh
T28ilAVw3/58FEX0BbjyvDPuamvS7CS6//ln3QTKhDr0lSGPwGGqRqSLJWtOW7cS
8oqNyy4FqLyw0lAtaGpaie4zLaJ4NBLP3lW+8rFhTDO/82Oa8URnfIqnmS0OJdXq
SP/j4NPQXioaYoshOlGOBqI9m3g+tECiW1KfpA7Jgh/4DQC752qbqD8IO1CDMqK5
hWxa/ngKG4ZvXatyY+FV9kKdMJKSLeB3tvDMA+2SDkS0wGan31HlRG6pCg0T4XBq
8CuYd9pDl47mH1W7ogUbVU2BX+6PYpKQt3d0plgt/TqBxIrX1Q2LRI615+3dopcN
xUFmbnHhCuK18J6HhqX2aFrP5us3YXn5FMhDBf/XYT3iiLYb9tv6Hnd2N0tnNnvJ
Vs4EoZfnurNoSoNkFdMlf3h4jYjOyEwORX2ihoRIcFFRfqe7LTqFhzDAKtpVhuCt
1M+I6LYy6cUQvQCBhNw7mdGOmVb5zlsWv5jjN92qBYfgqp4L1fzSVugyBUwAhoc4
4tQ05ga7unTr3ECfjn9BumLxbZP6VN2RbXZFkGP9xIszgdV/gSrDU5GTB5JLE03I
U5pPlG4ogSnVG9ULGTaMlSJMF5RXtOPuT9v4AmMu74K6aq+/9gBKnLSV62LZwIFD
N0/59Nh0FJaalStRmQl8oHjWW2V7UMCp5hVar+T8Us2ka7Gts3O+JiZbu18/U+05
etBLzOGiNiXRGbnLIyGjns9rHr8xwCkVSJY8j7gZ67GDX1c4b4a1nIPiTr6JebQs
iNZyY2Z0fZTbbSAnASEhLpeLm4d1Fr6g7/kBjjbrcxJaDlVTWNaGARRw/Lfhv3A7
yxrwXSx+THty/37RjFN87n5aoidwj0svYba1oRpdKSBDuG03qHLH0sM4EKDh0SwD
Wq/4ER+bvXYFNf0TWHnx5rbWk5j8G4C6iVUD1ZPS0RulnbrpKhZu2O/pmPVad2gg
xA7uhF7Lk2WWG4fjfH/OJ9tpfXA+TFbqsm6S+gpCbS37XnMe41laMXuC6/jru80O
uSaHQlEIJhG8d/6PP5JPnSaZBMH896IXUk1Pvsx2BzSsOsOYBn6y97/HJKNboCWS
XlMKGoQPzFlJ2ny/8+14OU2vYwteM5SIATwqEVBFR643yqjaZ+nl/ZQ9IwOlXpng
z/dPLG+cRbfjx4MkdGZRy5v/IDuXi4wHZo9HWb2FdOi6he9QhsDDYBAR46QYwM38
1lNLSst5w+dmjtT9NKNLe33RNT6RkK738JKbLZZnAINVMjaJHyChWKTXQ/qZfCOf
O4VHCVnhBp8Au6Kqb/W+WMOusTGxF/KRo2AnpiH8Pg68IM3N0ItTe/Dr178or+jt
+HKXXUh+tsDtDrFI3/ocUvsnKvuOT9rhIn25chEuOIcYvy7pX3L+fxvazxhC4SIv
AHaoRS2rdCCUgfEiT6/P3UaLcnLVtTDmFJhGK2IjHoZMBtgQCXlsikAbQeVj08Cv
nQAfEXBmNpWnl+Ogu7Bx0GmkfAOz/ActWWQvMAZHCq/0wyRR/uh8By6tPqCLgKIM
/Vnszd1M2O7/iUZz9kk6ITFEeXKA++6r/7IhuBUZz06GbL+0kcHPZJDy12l/8g8l
cusFB5ULalMUd0Qd+Ve+xLVNd6j0Rc3iLf0+PdPCYRASeDSPVByRztE7N6O2edum
bgF60x8RRR4KzmqBPsGbs1HOUQARz2NPKD2WMQEsTOw2F+iKeb1/79uJuK5qNOpm
5gEqc8t/q2XdvMAnwWwyRDxNHGuEIY1AWdHs2/Y9XJRwt/Db/mQSTREhMuCVhZBa
WLTAWUISXJM7C0pe5dVTlYnXi8z8BDpFxAZ/6PgTR6ykdpkz3JoCyPxnKH6IIE86
pfAp5+EWnui3Onmig9p/F39ZlITWErueEAJ+oHUX9dDJhFvqMYeRtyus8L8ZgAZs
comPeM2h9W9Zb3NibdCe5G0G8gNL10QDoy98VK8OfJ2CbJZkwrJibBhH067OTgIV
ApvnHLTQE5Z4DScYb7evsC6HCoQ+gEN1AuMIeD0VJmzkwcQmHaSYMq3l9TM1lr2U
Jn1XyMbH/YLW49MTPF+FyxHflH4hCKOIwu1LiEhXsf2hqGmEWh8C4rYki4bXCeQq
uf758tKYOou/uKeaMSVTgbu06AP0yS7sDHZr/hnIZLOIIr+1G4j8/tcq5x6nSN/r
rL8FHkJp3zMVuphazeAlD4D7POkdso+YuncBiEmQa8Fh4MQo6KSfXazfU5e/ZBEL
4Gm86EfkJJogmPPa3X4qs08lpO53v3p2GfZdMoSZuncRdIqbEAxR29hzpgSlptbM
rFqDY9XrK11hpv7n4YxPsGOrb/eqDkIBkQ1Pu6Dztx4QnEcOaT9vgJaSpYyjT24G
1ousyb2q5ZqBQ8PH8K1cvqVTkXDNZid+MxJutmpytts+8rTLblcH61N4PNLc4Y1H
WT9+ANVL1C/AqZgLmWsW+N/UVhXbD3zLkO0Z+yMxHsRZ7TIBVBbXkDk3x2UGJerJ
tvmQqVOK02RLvf0TjCWN1LK8Bbhd9r6SJmwV1IOMuJ+b4JCPV4itnxtLvvXGTQxH
rNBysECGiwR2s349bZvPJubIAeOXk5Q75ZifQJuEC30ttpkpaF9A8WV9QdnAQTxS
V/i+E3MTNLXv1jteTarwjsYkkvavoYQxDnA0UqY03rULU+aBUxD6N1+8lR4FX6Al
afihFw3rJEmbj7fyGmz1W2qfx5EQrdfsWzCVDqNwDhNZE73Hc0z1KUbVgodT+TlC
R4cUif5gir6zMSNONLaBSJpffOvW8R52zLQVk+07q0mPtF0RRlJV07jivQQoIlr2
jrwf2YLnciHNyYQCby9uHzcEWzXC2pB2/9zDGfquqvEqMYy8R7aJ5PSvg1O5u/4R
gfNyU3T+Qfc6GLfhW9wcF5CU2qFsr/3CxMeirfzdGphuqoxniXJkS7NwpxReY3WI
sjXzowu6j2Psg1kNxJOuVStpH3cXREZnffvv6WKC9ycqp4xDxBfXTS86sWTK7xLx
7vKI7ilsfCt2J9mzXXn/zPX2tue+DN1Qi3V7QLggcKsR21xN6zP9wsLvHAN+wkGN
qxM/B/+cUrJ+0AcAWgbw4RnWP/tYRAvNC5+egz+q8A3T8eXoOsNwQEUcuaxxwkbR
lJd4jGiuodD1RF9q+Gz0Y+ia1w/7mThZAXT1K/SIo/+n4dSKjM3Ibg8i9WUQ46Hr
SUSFMnQKYYxxEqx9PJE9/5CdMcDtmHuN18HaqKu9pKorBaVqDaoAuziE4n4ptPk0
ES8mjYyzYcmkkMr6RKmUbPfWHJturV7VQgJPDaCBjE2VqyL84yJZ0sukmwGwppd0
yUuSpRowgz5wK92mxNH9MuciPmvfOEHc9U9Ia2QQ3rQHxoeeL7SFKdfgjLtSwgR2
ZRla7qVvlZz7oV05+NGNVqzC7Um3kZk+MR/jTCtdJTbJOgWA6bwNuiCmH5iNfYWW
C6lwwpoOYklQN4akzuGPqdc4cdmtfQKIuCVs2Ar6dPPUanCSha8GY5ZgRcWNs6dB
fxewyqWJnHX8N3WM+fShKuCg/QY+lA66WGuiZZ7gycAG4bnfkyTi0eg0DklgjdNS
Pjclx5n0gXzOtFc5NAt/p9vE5cDaIsH1E27IHTKtwTkf9WIv9DZ6hLQT9zU1v6Mt
DIlA90bxKiOM4usBwPVBOa1Ogdjn6IJCXcRrIPADlhMEfeqZKczPFs3d1yEB0N9A
AXdDFmOT6DkD2i+X0RpgzBQ8evHeYwnu/IiMVwB0ueodJSavimugyLQuvyIfRY+8
tlM2BXUSmKeIOZO+3fISlFcpFR4h5nYU57V083DmmZp+ZdTY5jB017qU/8pnmJBy
3FWjXYC7phsnSOij+io0yS0uBogVi/OwnI/Z4boomfM68Hj+N5DbG7UbvfyuCwGo
FdlNkHq9VE5nziIrrHqTdOMmHtD+SgSmw1hknkbdiMca1sF41Fh64QE7cACAlBz1
X2KxeFQHcuDNOmLxM8aVHrUScFxGskBn7oqLSW5AZ5dDCAAsqvonHIltA3apNRXg
zmmu/7Sd9L/plDwROISsRFtXEFYobafha3yMjpd5PAnn5a3Uk5BiQMVYTC0TGYzf
I0RspDdtgSY1WgkOMgSbLM47+xLWhDOX94jW1E9PTc7cBj4JBe+MTIpPLAAK46BU
gAR8ku7uDM2SapVbSNu05Xe4JosxxUA5oM6rAjvAlkT1W9cxRb+RGiTWcYYLHOVy
YVyi60zWb1tb87bSYwfA+ao0z2/KbMGWI3WBzYDTbbGGudsybTS4G6MrlSbhwh7z
DD/8Yq4r+8OP/q/WpVXTIH5zRmJz69Io0l4EWa3D16tJcdF3kWRknQPhikufAKxC
RIfCBLpg7RNSEjUSCKVfl/tf9n7taT4MAf9vs3draffQhJwirWkfxL0hcPrSrA0C
inZqTr6taWfWD8WNI14+J1SbTQRlJfGk40JoMHJRGYvb9KhmPxIv5IoJTRYhmF4j
WOlJfTjzyKqvBmylH2nNUqmOsPpNoJPLXFtCL+t5/6YeF56hlHe2nT7TGrGU8CjL
F8ctrnHrQFgwiAGShwwOzQmzc330tv5PnNeEyvI0Gc4PHTI6NQCvj9rlV6B3br+2
dM2emydYnFORZbFHyLbTnlTGKpTdVKHJlUuI+ksxOa6eLd8Oled1usT7Xnrbbsud
PG0useHf86CCMSS8Qcqq2gHjtuGYsyHDWYPfIhKCrjyunNJjILIlb80fQI9Ss1yQ
9B99/NH7pDqaOXEPkEXnlnq2YkeJWUH72j71CC+cKDhm6VBCWtfwhhAuZulIl2sw
oWmELPFxRjtdZUitDAzpi1NzBA7zJU4ES1NBjEJDd+ylcB/tgARaY+ZhH/3j06ZC
VPGsDOYxTPQhq6dtlgPZka+Y5oFjFJ0f9ETwAhv/AqRIGCLYAOxhWybhHDSurVwj
N7QEQVOI4+ST7f6AZ1y92pKtGO4LJTwCnWS7YFWkigulTseus9wv+UhHMJWzUbql
AiJ33wUnLUF8gRKLXF9tm2CHYOfvc1y0ZORuRFuDFH53WJGQMQic/m86OeFL2Lq9
o8ixGsZPKGObDAscgehlKl5MDwMGOnK6wRMm9LpTMR46WPsj8dzZ69gN0RRgUn1b
4KuN7EkRYTkMHeiBO2XJMzbaD+m59s1DhEEft7mFRtnOgW1hmVWocJn/x4IuTStL
r79wUxQQvDUc6oOVBzxNyOkssyHSZJLZjM92IUqSNxpfJowNO17uCZiWB6gET/jO
geSFRr4mryT9v4Ax4MMh8OS1v+9vnMnZ99OFDPVI5grUzxrIl/dQCHWBj/Tt3b9e
hcZ+V3ZRwVuUFL4s4McvRX/opZ9QdxQqBXa5o8GhmyAIyttfOGdW2MVJJYwaJ6f9
Uayfu4pYWF5OUoHh0eYHyVvg5ZDiU7TOahDIXjur6h8y8X6yyyTYrfiVozZa/uMC
N/Y4TXCYLWyMKuDZm/2CVhcznZWC23lByKx9DwqSNXQgZtpPom5ZEnXFNXZY9FUG
jTarHb25jnnyWWurBEaoWszPvGyJ3Lf6tAKc8sUFxRyBULzxHF/JePG6nm51B9MP
fgAo0QWBHvrMp2m5Ettsri3grzUSGfpWzzTd3Oaqen/J31T1MoFG9i7sLHK0s0MG
+jXLWEVZDWyKeoo0XLzQnCTRBgN51tAkVZnCVNjsl0BrvZng1O2d0GkyD8Pdd29T
IRKVhVzH57/fqRtVm9MLojMauiAspxq38sjjZzxO4fQAt82r7sbGwk34MnotATwa
i4aKnsjRPGufbES2JQxcPjmjziZfihg9WvUV2aiqXjde+z4mtJy+Sw0j0S8wt+wb
LdwaqDfyM3rdlC7aRuYTfUY7xz5a2HLRkTaKgd2XJAqCc9w12Qp4wmDGpW6WwEEl
V1dKSTyUOliH4zSI/U4hcHNYLcDEJudghTtW+OTuMEcJmy5Igd/UuUWWCQ1iKgvw
yyrYvDkE/fFJy+8kRFCq5rFb0AEamJnqaM7nJ/eemx+UOmknEWbr/6DO9uoRHzJw
8f0s4QzXGZvxMegYh3/GZAbC8m8GJvzVEPkvXyFSXb5/wN8eZaNEU1NAtdC2Ok/t
cv5g0HCz1cm5eg8LGGb0LIhXeojLYpxk0QV1gx1YF4bwwtjU3AsRqf0fQA1FHXkE
QQLGzKiLFgzTaSzAREoCjGlU6RByFrQzf3R+Rw6UFrYtknBaQn+ZfJsixAHRJZ93
/LI5Ol1NcpSOYuqiR9HZvHKq2HojO0nk7D983cmQiKf3DVazLu+ZXxy3TK7xi8vT
OyH4aPBp/PZ/QoMAoR35ORSMG4kQsscZOv1Ad5Ry59X/2uZPQqfFY/611HZoHcJo
Q2g9plz2Y0orgTYZygbN2NKoLkCSZY5t2cg46Fi+/684c9M1LTXcaftrypXm66V6
xBVk/0/Q11ynBLTTMLM5Hyg+P5ubQOjHcNnYE9TVhGnCTzx83GsXnqj2Zv7C/9sO
gy/MxxuBB/vzGAPAzeygTSMb7Kev97nUslufZ0QW9NUfV/Va4BifPLMTIR60gCOn
TNbkF7nm9f1pi5ZQRUOmZFnhGsUz7Nn5FBOKplzPmAnjvdNLI9ilEi91TEJ1gSMp
02C0HE/EmUfT6VuvAlPKSgrVKx0MIG/NUPxtk1ZSvCliFvlgYlBC0dkWj9xnHsPT
GEf7kOsudQaumWtYI7O2PpkNuisIvD76C2NTOFXJ4nAm7TQV4ixOB4Tbg6JPZ70O
shS2iafLjkiqW5h3dr4j6eDaTTZEVX55TbYZV5Pj3fMNY9KGaNnc7oggnOoW281s
lNciIiX/HZvTcFelPYjl0/EW8pHyx1gXWUvkkWnlFfRMsVW81pOuw2ytlSaYgbu/
Mg1fAb8Kb+z6Fk2hnq1E+bPwKjAnQRZgtImflNZ2ncRL3g+5P7YmOxLIDHP+4QAg
iAoxlWFSy5mhGASu6KrHNxz546YBYMSEMscfhBlbcoABJxw5t78oOo+APZQHc6LJ
xAY3eDUlId4yU/v6RY0rj+BmzynLdhSfqsLHSFMrQNYA47kaitZ3HopXBIUDiI2W
U4UzwY5G/UbGV8cm07oyO2ifwS5M/XlSuNmL2nxYQjOu+PG7zJHXhI6j/r2jfDUK
lv4W6Ts7vLZt8+hqHCp0bOHkfWYOoijnBCUM2Ymg0FdBwVQBUfEyFNyINd0MnMV2
uU+1NSj/bIQcJx48wEReCBW4pHjHgNfcF4BSX0Cb75AsX0X+rj1YYrX8lB7yf/ZN
Qb4yON0ykK1UfOWyPYxLQEVlk4UrWD+Kx4HYiVFT7L+dYyPXGWzohXPQlyRmozmc
wADyyMdUh1YIrKvC6cjisGliLC5HWPNRImlrhrBNKvcV27AkSWgpzq6MWXWQ7KVO
wdRbavu2jVI6aM828ayGiqoGZi/WuPLhQEMK5hrf964B2mH3sPTxd2ooLD/MhHXE
3KiHHHBdDzL3W63EHM0zXK4cnlodDfeVa3VJ4GGTmVLoblK+S6LjcT3UcFo9g45l
ZXOGjJvFjM/AqkWdk3g/kTESuCPQdoUApmo1WISAPCdH+LaeLn61N801Mvsk2teL
cIBFOilBpW7illr0RRBfcTUmqCGCds7uHw4GtBPd/cHGwDBSBfk8CtjHNA+V/KxM
2cuVCsrLPLzG2lT026BTe6r/Cu9qqGWuLckv5Cxi3c1BSqwCJfh25QKlHdMOvoAW
RaFhhBo8MNSm/3kmfl7569pi6EUzfvkxtXHfP8RRw28wgn6s+CFqiIK29WzUjbiF
+U0qxUFwV4hjmriG/Hzp74Xf6q0OGPY8KhUny7SbzwzpIlRmuk1h/CDtUS/7PWbZ
A1ZPBHJFOe2wn1mGXljbndx3Fa5cTCu62ElD496oLkdH9epWqboeWztJOF5ON1iw
HHAnzpTaBBkLrHmOUEqQMRTpF/F0rf4mompVQq0pWua3r3D8hhJn05sYQgmL9jFh
wGKYImpLKMoePU1X5VpcE8UuOoTfH83buPWLZ+ujTivi+RaXTH6s0ixxs8Z8QKU5
vnQTgM7WGwGJu38cQgWziq6t0WWMY6hHiaoWI3Jynh7taHuQ2B/FwuxcuyIb6hqN
hMmA+tqkLtS3G+HGBhj4v9sr3D886LWfJnF3E7H7S0opZ5Lo70svADy9PoX5W9pG
7+eJjdpjZofwVe7fh5a+Xq6Hx10xPJiuYMo6y/ZLhXG0EXvPptz2qhQPn5kbA0Za
GtFGt4jvttyM9TLj7mDGoEsu/3AKpYfhaEMMDHydTgY9phZ2e1gFO8IXcpy5//uE
SemoHS+4tPqoBiQwa8lNN/ZcOAFRCL0gASNJimFWmgbi/o2GK86qYwV0xpK7exXs
ojEwDmFVQd2mB0uej3q//k+MbhbEVRJ4dfMwTCK6OS2dHJdlVKVmwLNoTSxcACra
ypTmv4FTXR1DcgZSlU+pRownWr8EvHjtD0E3DaUKNDezIn2Q1bFZBgz4tYB3VFDs
Gz0VIPxQfZw08j7qS/G21PGnYHk7ews4TDYcYBI/fhtwugMwz+LeTy3pLDa4xzph
D8+NWTxhkv5knsXRvSbDaZzUBGY/6TbKWyXAFC/Pp19clMhh4xQGWE26tl3ql1H1
uDUZY7TnLSynVfJjqnHs/lGlPYAmWb4qbXm623x9Q4XeOACrTbeCWy2lrNzMVh2V
6KT2rGO6hkoja5r7A1Ec1Fk97K4UU36v8OzN5evGYlA7zkqlvb1POveGZnjG/s1w
egfnND4IR2spg7kcoqfZU5w1wKaMzQjtqgy1C0OprK6kdThzPYaXh/l9epsRpUM1
4jyPwNSJ73fIKh37gL9xGf4cNFXrkGMLLQW1OUHpu77BAOzCXwoLOCUjaVlnwHQQ
hf5GEu3jVZGMIwWlQPdJGZ53NscOE/LwxvWGM5QVU2HiOWv68QJ2n7Z14wB6cZmV
EUJKLE4Shn1rSW8IAv4yv0YN7lJixns9BtKl+JNzk5TyRk+2Exjua5T5GBfmsEF+
RSoWxqSu0yVr+htWTWBWH3ptPLl/XampTm6HRV6Wbymx5xt75hiEis4w15ALIGVA
2V6yHKPqOFgIkqfT/1VrAr/gPocW4bqmburkvcd9ql53+UDQ9ohFArF+NtoVtuoM
KyY+wCWJ7z6ygoLJ3Favr7d0+iFyLSr0QpqtNMO28zUHcuWn0fDFui7g82PgzLUb
AfkZYb1XM7+4wdI7/aaWwP82SIvnWbxUtj/Rn9FteEyF6l5qUVQo0Xi5f9lOsJpb
MtpxIIdA5hdl4lMr/oc0JyzwN5ZED6+8NhZ9CpbWEYPOJnS9vJjHaVVDHy25N+TL
60qgdtgyH2C6r7enUPCCFjWbW37SNonQO5FmOhBfyat/M8AbdKj+AMmSbG08lKcb
ymsRU9fBF73bBwq4NiLUzlzzWrYYuH1/ITGH2jLyS9cbCIizAu1UNjGyLR81IFuI
wNBwsXB1ttClbcMY9cbekfLJ5rT+XM+4m0bjYg6I4Gu6MvaUE0TvO6ghNjKhPdHp
f0hfaFS2ambWHFtC0S3ZiTM0GIc3cMz3XahftY28afFbwCxTn5IT1xI+gZXiJRjj
0s3kIKIA0+qB6PJ3KKeyH67/X/HA4GBDDtrbzhg5z/KUeKpfM51NI8A3ISVStESq
CHC0kkzvE3mf+CUvpwCJQaS13PTywz4Mzbityjhnarz0ORwh/vhnuOAMgbyamDT9
6eDo5HOaeRewbTflJ4jGbQSjGUiA5pQY9Es9p3DIDZXQ4yZlH5e35k+idolnz3Fk
/ylbR38TAV7ArR9n2T+tyJawoGCtKK5TuUuqAYXWIUEpnXuxtLkTLc1cEnxv6ZJm
MDgC/Y3gKNQBjYd1uwwhBAWWFaUN2QC21tvF2OjszojAW79JSViXstj+3gPyVuAs
OVbASLCBDDm4qOgGL2s2frbDnjDQ4z1HRxGvSWRgoGAg8rphq4qW72l6wISW0S4+
ctgS5IJeXyoxDK9Xn5fR+/WUl8xHeqZHQ3yjEgYozP9+Y1l8+am7MsKZsbw6kB4n
LcV5Nme9Wn9EHmIesKqKIjqJ7LcXRt7xzuTs+km4TlVzAXR+U96PtoYJ0++O7QUa
eOJWbhDzRTuWqOgjgIn9eykqbmQJ+I9F6CIMf7DqJTi7DnyLjWdhoZ4vPW79HEM/
bKFwanI+9Ce/i6HJDqTAakUD/SrOL3+2+kQCXYrSegHGUnnLoCcqKoz3A6U6LYBI
AZ0FflmP/5suQAQNXMs68EnbKQmyAWRq/4O3tpEX/TajjkGs+021M82J6IQpZJUg
lpUl9UzlzC5tcnfBPcccV7hFS5rcMKaQ3Jb9MAaTr2zHELgQ3git9yNS+dNJ1ZbZ
rWyXZOi3a8KRDsz/VufBOJfMIHZy81QOgYScnAzSh7LrRU1W0xUesmDoyWeyPUjN
6RqezB8nh+1k+VDuEARbfBSLNKX6TigbRm256mjRaYg58zwp5cGJo5QOhhbkDZDF
LpEfWFC85Qt3HQXpuB2MgcBZTmhMUhKHiaWCFw8J8rSgeTQrLsNTag88ZP1KMfGp
ywt/V+JZYso02mMJ39LY4VZGG7DPx2fM95LfdTdEPL5fe0N5WZzHnwcmqW8QgDg3
4cFseD4FkBAGklICH4gRCAupxtobOceQ7KXM0rPtoXAN/rgqs8PDWREa2+rw8syY
GFIXSLjFPeCEysLV7VK2vLtau95dyFbsgizfyobJFN3dH67g0lcdhUw5+VQ3dlb9
txjNZXeJ0g9qOKZ9mJVQMdW7SqMIaBnL7tUF8OBNFbYanzoV1vQQ6qROU6/2cNas
5QRsChU11pJjOlFK+0+tTcvEuKHVW46ExC1sRcwJGMfhhSFiSg03TqqOv+J5etBG
smRkmrn9xVBPEWjaMOoSpsMcH9n2HcZks4K7WVPM+X/O7dfwdPXOVJd50NDqXyf8
xU+Hw1uMOVNRNA+PI+YKMLNbUCBovM4dzK5vtbnOYasrVqyHswO29aJnkFI/0buw
M0TgTZD7zVynGcdE9wu6g5S11myoAWvowYqhTkYUp1WIXmKeysRPRliDk6HP8X+I
fq8paS86kspPT4mwS0E1OZaSGJKH7sLo0rpnSfWNeEHqPVs5QKRlvMglTvaWEzXQ
sjSbULRnQz7vBUcpM5JxVt3on+sYmtJB7F4Xik1HS5t8aRBxKyr4AxAvUjq67KiX
BRqEQqRIsRZzFt7om2kmvg0BsDYsdP+ETjov+oexL/OXreK/nrtPEUvYfZVZP/LF
WC4XSDgGpfEr3qatzByq24g7V+/+mIZD8i9HrbEg2xHah/+xvhUGR2NYw4dYE1Tf
gaQxG23/dYJJQdg0GbpJIG6TcWsEZ2dP9DRbn2zKntv9sQxEf2GyyBabgOydsp3N
CY61v4yfZFvXzjoVUhxfOGJgPq5UyR5HzxrJsBAg9/ankxofLP82howGt0Pknvht
FFkuXLsKH1+I7s72jnIxNCs0aP7yOK6gv1PpYwgbdkESur74bhlo5bZWyKbOcc9I
+s/eN4kFaU2z6cCSiVnfDnlzuc0LYxhpy87S7JG4SKAeemAfxQFDto83ICG7tP+7
Qfyac3S9z9XZmEoWBoiUQ7L7XwMiatkTLt1Fa8s36sOxEiJnSZVWvwhbnhsYAs+w
gcQCWU+p7SrI16SqdZNAw29HZtI4Za7QsMW0oZW7wUxNJZQBBG0fwtYG6XlZPwc0
T6KnJ2JfJ/J+3c4qo5W7Q3Ye8udNqp/O682PmrvjP5psnC9d+0xYSEPmSvbqfDWA
OKPq8SYy59ePeDY8Z+nAR4J2FNVMZ6t3wzc65AJjLqRv5RG2VV4Z+JUH1QmJoBPs
D3OFxNoAbqX8rNe8QCHLDul83sJbTIZGOxHnY8DuaFnuq0T4GqFNAqKBtoKHKtGH
Vl50cQr/XCmLiCJWDfych2MaTBR1oIeAHldfgh6T7b+uIJ1izf1tB/9MZtzeBkxI
ezG1DEjNcbD8s+Js297P0aFKZuSHyJxAAtuc6JNmgYi6V0Uo1n9e0Q9pQymwmqJn
cbRaLadlC0KV+qvXBI1G/uvNpj1FXoJRPvh/Yi+vGIseJyXucldticsGxe+/i0Xg
v26Z/ExWBGj9gjoC8Scy54T+yxpgf9JKkIS+u0jxc++62qSSpBordqQ37cL243Nk
GA2Luy9mdHbGpOKSxc5WCn7U2Di4PQfdeWvFvbigcQm48CS8mRXiheogQB7goYC1
JT0FeUlgJDd4m3POHQKclLaCUdrIvz+sWxio5qZhbv46kebbYGTj9oKMnfzFANII
F166leFXKV4HGDlIh2qIrqm3AKv4qK8QI9VPQradudUCi9msa8CSz1oxZ2BOiYAE
1s4NDDF6pDONXM8yqpbGtsZAcI+NIqjp6Z7vFN1zaK1DCDNVr1fDHhVG4DFFWMV7
vfEgqKEXP74JgTWqCKWMX5mX4i/sJvfoS34Q4lnbOTIAPGPNRcKcl4Q+ZY6VHAgc
7dD/dL1q4JEwCVyhIgKEOTzWuVfmDXKG/a4mppwhptt4jj9FE4uIrue+tLAIZ+m6
QgX1oWqT5z9Dd09Oe35tyKet8RtwVh92mImoLD3Q0q8Fnwy12VrvQkjoIyPKw06P
7Z2Cs0kkfutHPAhVgWMCyDp13aq4q2OiVy0LzsU2D3sz9yNbNeD1IxC+EZJ/pvBJ
a8RYZrNSCYnMB+c0ieCyOfhL73tpiRY/M6gOBujrJcJZfJ3peCLH23VoySWNAtXd
xZwl/AhbeJFUIY6J/C2+hqbRATFczl8qYsTP0yu+1NQmg3pTvKr127gyYTne7uKB
IMb9xd1fglCQ6+HB2PEYl+lncIWsm93R2ibj0OCbs88ngIjgvrfW64PqZm+jgGCF
l/baaB8A8MJAJzZi2Op1r76QWFNT/epx0/c0SezDwuyWiNN5gOoEOJhD/9vMdGTX
uuxlOrJZnZu/1liOAHQ+uoEw18gV6YUznzEGAj/9F4YExa8WgSFo5TRWRq3SiRIE
omee2+0MemdQ9fB6yV/XlWAhIEP+16u68XlCd6QQ+kzfom4cn7TXInYTmSeTrncb
stMDP6fn44/tTpnLexyhBbR7fDsvhATFbqiie/k8M7e3Md28ddwGSgjrnYW++M7w
/JY9VCSF+DHn3uNmjvkFCCQgrV/ud26DfQP+F7SIMYWkjEoh8j7+b0jXaFVNAIXl
4PQpGy5WrkF7eqxu83Lqpu+CvM3PzwpKWnvwxa2RiA+ipJUsTEMGaEPWp3S42DPr
+mIDFaCQj44dbrHqC/wBWuwXkAROSDBPaXA/6oOinTwN5LXVzVWcqM54RmyMNnXG
wZEquXfF1rUsV6X7TJgudgnT7WbmqlfKrrG+1NGZbvQJJ8YL0T+j0DZbdZcODYAB
pecg74uw1hux6E1AjlHbOHMa7IXLwcIyDn9eoAQ8XeOT2oQ1eKaaEwsdmkWogK04
BQ6A0ioFzVOoBSDR1V8NDoMuWuTtgwy3LmgTJqpq55gTRNEABvsVebzKmlF8LtN0
qX2W0yX0ZBuIrQxAAB5F3aX6IbRp94+oe+tLZGG3eZz5W/+95HRppHF4zWuSUE9w
jcNnU6+ZyuZoo0XJsjW7ovIsL9ZG9TXmmj0sqYLPKPqvnHHJz9KLPndFYc+2eODC
T56AP5cG48n9Tz9KxH4kP4p5xnGTEhYbLHO+MU11UNlyUs/7UWKnkwlQ2A8wS+7z
unRY0j3SJ1UflyFHV3YqslfHxnqBjMDB6hYCHds3cplZSyx1CN4PVZWbAy7Sj2fy
zFkDA/2NRqlLtrsE0WbiduS9UYGefRkZK7Ygrq2KyU331VAlU/i8SJrapvRhZl9+
oxaj5B4T0akd9k+/qdGkIdR2gAyWF7RJovKJ1Kf/vZO3ffn53odqIVOfLSX4SyKM
M1+oG0JAvdUsRindVAL9oXuebTq7z7N8yd/0PzRdCogak5Ncx9hNtB1vCuVxWtSA
5eNW5JXgtWHVPex8cjb3lR3I/ielef+etTvwyDRb8jJA+TVPk1/z7137feproU+o
4HUq4iEVb/fDHBGn94QFJHj87+nCxlog0sp5WSjcjFh3dW9f3ptaROh1mY9QLw4M
ZjQWJ2INspjF6juzpqjqVVbApSnpePssq3M/3kCsZXDSYa37Dpq/qHPW9W1OV3vR
AYUO3yltWW1p2LEuf7SeBEamtoOMozZYT3wRn10pOhGGeqI8jY1p2+FaMGtUEyPT
/fBxZypQN9+CbldztCmV6R7HR3g7lCt5QkIjOsGZT5WjZRb2xSUKtQdftUxYGvxJ
USqJyCGix2JWvaAp5frryUFJBPUsQGl2L/1AJXHd4r5bbtJa9cod9AcghyUXJ51v
tIazQL5akQH4WylLMIxoBPCGaC2zUj3s47glxgF5cPYyS6BtRH28JVuqI+v+c4vX
R+kohaFmx4554R92mcN5H3dmKlUhVlcEQMK4w5CsEDf27tIabnygJUrGnCd8oSQa
azFu5vKA/GMscNmYHttpB0qFpyc8HR0IUGb1iXlh8yrqdFd+I11RB6kLplLYlHjS
cdXGrbs4iKf/NlRyUZ20Rb17/mV0+z0YgtxgBGXV8mHClaA0sVggOKCD2PRT/W6I
2JGR/gIPKrQSNZW+eDIddEKBZJ8b5pJc2DpmMszvbj+lmaKVqxS0xuhgILR+VLDg
WGvLVfLtU+q1zFtA6gYouJB8YOnEHyPK2eqr9/OdZWHmnNiqSEj5K2BvpFhdPa0T
o6rx5by1cZCeQn5GQzgkkGduqsrXaxFzQaVH8QzwOuPZGC6A+LM12LpUzHoKGqls
FHZN6VGFYOm/Oq2IJzfhNkrbZuMbLiWOPoKix2Bl+0fV8xAL61PNvaHF2GvsoZvV
dwYPq1WdVg/xWq9Cy16phT1aJ50/XpeGvtc51hC3SYCHb0cDElNwVwuOm+2w2aWZ
nU4gX2ZftkJRp78mRB3GrMuqhybueHj4P7BW6PSB+EsVkuIhflBFP6HIV9DGWX6S
0ZqFQcFAn0/X1s3J0Je9y7FleAnmCy1rWlWWgUhp3qf+7Q3LGCQrJTaNInFBNqLF
dYvZZur8T+Sp4QmYooASNFmCmHtJXMm5QG5TFJKzuV+BlkDO+eb8kkFLVdK/+fak
FMp8Cf2vIceDR5GlPDoFLtVY+7sJZWZdyi/Bgy/ipAya2as2PEvBnHCf68aPuSUI
MekZTanF7CateSCh+eKN2ULX2JZ/x9QbTHVBE8vEOSgEiJXHhNiwtrw/aiE7fepY
Ab5O98c/Li4XIARYHYM8hq+IwFl0pgUr5zqE+PfVsU2JPoC5YFt8Ugy3LiZ9s+Bf
5R9icNozQpzAtnunV3Tpefokt2kkynHUEMj1wGOvZpNjY4pnXuXo8jR4UVTZa9Sd
y0QTk8LvzN4aYSut7Wo57gP+vEWT8xADzKw3TcSODgY5MSIB7fDqeP0hfMi3ZiBs
mEUIQddMzVzPG1KNbrLA/IKz1ZJGyQ2+W3C0bVTryk2tZmm03s/klsqrEAblz9vm
xFISLeM4CWG6JPPiygi4+K7w/a3sfJpjyMHY6DGRVt7jowzU42Bxoupmc9vnQ+CF
zLiSwilnfSpArkv8bjhqKyM6SslNQjY977mLoniApp0bZUsENjFmqplXa7lalrBL
vweIho2+ajVC4+ZN5WSfC4xFe/xaQ17bPjfWBzN9XKUMtRmAf7hLMSnD+mCBZwPU
coMAZZ5dWWO/8GjFQxh8e/57QQv5rqywS+0zK5FFvyac4mw5ckDmst11uYi1rdoS
A0RHFO8Ox9tP9SR3TesWbSSRWmnkNG9RHip/4kvViSWNQdfp+gIPIPFeIc5/nY3t
A0UnT91BzQ/RLxuxR2GrNJdnN2iWQBOx8zJVc7GkE1DiBjJPztBw5oLGnzdBDDVH
vWBxGqzObrY+XMOLC73Toxt6RwlH51amFxt4egNlsiPLKVd3ymLrm+QUEedbOMBW
4zMN9TRJzeQcTJkaWCeBX1LKX+9RPBbVdG8uBBEGZe+s1EdV9NV6C6NdTWuc09PK
h40onuX3LZkFirln9Xd04h+63aK8Lp0e+RrFAXOPx6YfOyDLkygZdagKdw7R0slP
pC9GHZRfImdrdtunOPsW1LwDi7aCLDlFIVFcM7sryrFlm09Zegs2g/f5Cbs6SNRM
iKXN9+0K5fbK+T4Yk8jI/KCngosdtqwkoGlTMXJZis9TB6BxZDa1M+ZwBAaph/kP
s0rLPvEEKcQfnBivqw3Y0x7dF4JcOGCZvpFVMKGZTMsI4PJzkHRPPRA0t+HtHOab
sEc+2mQodQfKZLh92HUslvq2HK4PW6BdVtBnoRNY+yxHhVzs1ASiobyPTAdpr3cN
fcoJjWM4NlZT9JMhosxyrCYL+jurYGxjGtU6n6rxYWbdkEalXBcNpNs51Zc7YyTs
KkEY6Tc+eSqf9bTx5J78YNY20pp84KmuC+RTB2MUZ8I+l0i9psFwp7hekWIAvGtN
Vu6IS0IUA/05ZFOulsutUc6mwPqzOju7rjuwjR8ptygYH6S3y238HwLb2584dA8A
LB28YI1D1Em6XDsCnD1Fm0jx41viAcxaLOOFbzlGMX3AWVqQbVwjtHiJ9BUfH6EV
3x3Eb/HywGsHCDhzKRQoMfAoXLWr92xriWMVnVAS1mwKexJz6y52QAGYBfg/66SK
cSVVNr8LjWVrH4MsCjSYlnlKP1q80++ovXBA94YiDOjtchlADs1RcelJudZIzFL1
alwtYEI4XFQCcYtu8808dgWobKx2cHXTYI6so1xsnDk8FSDDag/Nly0K1pPd94GU
P9AW0mw3OU9yBSoJEY37fMp8Fh2q4gtaQHoJzlxmi6RyybknEsbDPbUlbUwcLELd
VSFl2RkyjtvqaOCdgsWgZLBR+0WdM7kd2C5WGKe4x44mYGZYpF8jSPZmDd7PDQ74
6EFYHDQRJqzReLKKfU1I/27oyb85aYq4uvXsuPqwOUfGb/GMvgBigADdduk2+Sef
ZtENg+0mNg87Oy6d2Ykw+RoReV/3dL1NlMeg1GA3/CLV0PhrksVRb5MCFCR1q7h6
bxWM3A6EtBDCetDtwzk0ZljbAz7Eu7luwBohxsNntKTs4zVRQ/FF3MknHq26WORY
sDGzeSZHQ6XhubBrzJpfCPDKKAwdrnwq7XLQFo9JLgPxTFoui8UHujMBwQI6tqaY
lIePZ99DSq71ste0P/nOWx1i/WOHVdF8rclsTWaDrHx34BmLTwAJ2RspRZZAX8Cb
FgNbhBgA6sRIv+MI3cUOl+kBGKyWhtc8I0yRQlnkR0itvrDPOy80qTmoVBZIAweo
ZeEPcKYfsW1cmTkq9wQTzN5RlNvTOihf+4tEKPo1lZMvy1nl/PoCPVSMI/HX1sK5
zoJUfeqxer3IqkdyvauZ0LO85Kl20Pljl6ZI1QqZhY6YNxQJG1fF4Z0b5JIoG6n1
PMYDjwh9fB2oWBU8De+KKToTrHCk8NzYbLO2IprwplXneNPxRX8beH5zLclsujVx
svLvntz4vFWJDFf0b7LSfpQK2xSEXvZ4xcHg7gXQUIPFIK8GtB73iLZ80m3yfavc
uezVaNv/c0yDcHHf4BjLswL6YjlNaafy+0rJwZbP8xbULwaYe1CO8sn10T7iuf2K
SpOsPCQReEVBBrS0lpRZkTDhWdWu+mKWfjab52Ef7hB/vS6DPf+dUfoI1syzfceB
IP8+hsvRk3qs4+4dgmiKCShpJWpvifZTjCZMDqSOaRfifMVyR6whRHB7dD3rY/VS
+TszGSTcEqUR8p6U+kFg3g8j0U+7mXeoKOUrlYGToyotM1z7dIu3KOoXw8fSRmzn
98DGpZA7x/1OGrb/oJyo4bfqRbpg3UfH2EFqmpUuOj8mToOzxIdVjODGDmZUC6hu
U9+vXYRiAS2/RkLh5hHaJrkfcv/PEcJNkYoVimHWDy0Fl+uIZ6UWVJKJcG3sDX0l
Qd0K9DlyH5iJwG+1GYrUvfvy3M2IOP5Z0XcZ5WyjMCLBPXPgTNIIgwjyclxPnKPi
XISD2JREtIdv7YqXEUH4QcZZbMiPlQ/DuGpF1iLYTMPX+a2v+Vn62eshWxi6Bia4
A/1bIBilpPpmqKjeQxdGoVfEZNnuTBEGW3ucM0rQSo5Z6ApEM5Tb56sxuyq+GnOG
oM4NUUvAvwHavyx1Ti8blaob90xoROxwimxZJwazFy7Uc8TU3fL8plxEDCQZiqhW
AkWJdd3rNCRVBL/ffKR1RXTTskbw5PoHx+u9ePLLjPyUwrScGXnSNECJV9koJayq
iR9zvfaN4MyANh0GErqbmSdKFARhATmyxB0Y+vwA0cZn6DVSiuNjAN2REkP1jkqm
EbtKaYXD47pu4PpWvcaMrrV2El9GQTWjd3eBDDa8dj3j2Su3oGi8jcOVztXfiWqD
qWS6Oc1za2dnL+tkwWeV4blWtk2Ce+o1gJVTme1nkL5DjerRJ2f8k77SkNc4Qlnr
UgH33uV7YiIo6azvSAKE4WmzCuuoG9voYzLsIklpx9B9Sq+IkPuP/tr0GtoaZbXX
P0WDx+PhTUyFjS4z3VoxyfEzOxCier9raXChxosOzYSUPzocKRtgDDBHjIegyPnE
3SPq6HzavuonwWheLvNNCxoBYc6wW+/UqN4JS9QEOb77f2zF5FwhPNqtNbtZyUxK
tdaWn0WhoOLUPAm9u4OLGLmHRJfklkCs3TMZOeOruz056E4TcGeqZxrzxyfFxV3a
qZvqbAszUtkrWqM9VtxLOaAA7sHbmIvyWeCJMb9r2epP930p1x3/bjqWXlpcwwHB
vyRTiE0IoMBEqMQcZ1cd7AeSWdf0u7DG7yNO7+K/msTglFsnyJlLdovsoqUwwnWY
aELaabkShQFZ3xuGnhy9uT+iy64MhIETPw3M53OzQKGubdS/IMfVYqSePzKJkVfl
uLtspFUaspEbuRyZ/dJ3iMsqEwdzfQb1lSM8mueTQ85VH+hQqpzg3D07TNUEGcKM
B7pzWfS6U8LD1pCFIuLBmwYjbWhLeIUV/Tga6rbObS7rU1tq8HkmfsUCxwdc/fGE
SOvk2IGCnrmPpLpxCbVCp04NmphkX25rA/R1LdCLRXaE/M57Q1OVgdrhItCBiOc9
ag8B6I/7BN5OcDyZ1crLTTZKROcqxM/ago5gRwJ0cUra7B+H8Mg3Ui9SFqXe1Toq
YMhQjpQYHQi20h/uOjI9LJJCxp+eqoXExA4+VFWaCWsh7M37fWAevUc8C0E3G9f/
rvTrQaPqLNYcO1+GhU/Tp/kqh0t4mlLHspAJej/DGEbZ4oO2d6giY3awpUxLvYlA
aoye3MJjwqzMsgC2TRNMvLFiEbN3ygACaDEL2+2hEE1eZoseDr/olofcFTu7Jgfl
0UaEo/ObLvMNm3vnj1qx9+oJFvGGUR0QuBMMBlje3sMcJMF0Fzo/SLjC6+JOqKWd
8CUJuvrbZsprVBE9oclwF27KAA5cKEBnvSK+eSKgP6dMVfpSvqKkPN1qLRk7VI3h
45ObDB14ZMHlQANudAtl+fmQuJ3M49ARKmRhE35X3O1GC02t9g5JGbnoXITZQ/Ek
Dh3CAuThcSEpd6A+xb6SiYQN5nGWi5z7umByb4wcjhtKL+4I0VrsUjjGAZzzAY1m
Ryp5gELF5jmZ9a4+uQgz7+KxJGcWb7cJegw9/4cRTE5BOFHCkl7fO+Qb6G0X+6Qh
7XUHpvn1pTunq20vJ16BwnFEHbVmM0x4GUyCpy1PIVNNiErvvA3fiWjA1GNh6FIw
RXLabD06FJizPCHC+w8ZxGlXbuat8kkr2mJ+cj1vJcfvjyeh5fewqIGoVZsZzeFO
Wnf3O2Xh2o+xFJ1+tEjLszqTn9n2uff14giZ6sTIuywes61LiIEfVYXpmsc9K+gs
s+9XcOB3p6/btWRI2rhW8H28VR4RyGjHpl5zEBfg0fAExU9/PRt8VM9Fwmw6bdtu
S8dufjsf46Cpn8IDOTzNqKH3tOBgZIeHB6moJkQtui93C8X3Rc/DZRj+mk5rQnDn
GcJnVTN3mWA1IJ0eSAdgy7vg6iwCArPgPC9YQHD10r5+7lHABC3/wQC6Rj/dmz0A
VieLqKvjhk8JbZMvl0jo5WwTLdFkEfsg33JelHOY7CO4iwa4/vlBGG4jBLRVDtlV
yrSSbjUgFfo8aBHiq7NHMSMyQaHyEzPeciSFvNZCn9OQ8jUQ7v/S4DyOexYjHs6g
UQdI/UC3R1JCEZti7I1VoeTuBVVH+PtX2BqxaIWRZZ1dodInPeH+mU++ShCJ3Asw
L3L0p+DcPn+ZCA3zkzrkxgQ4s670B+DUZ2D0f8xylyz3ykltrtyepyh/NIYsUHyc
YRRorOMueg6n+roXEkym2vuJkNN/C7YiqKi0HuuY8kMaw87CReo+18KiiEa9SC1l
33wNF/9tV6QOivrZDsDXWWSry6GRM9rQnR85c/0zzMCMuywqGpzKssLIYFedoVG2
IwROsJLrpqze8uwcnIY63FCB6+UnehscOGPpxw+RonZtAIa9NU9bnLpl3NOpZ3kA
B/WtLtL2ywE3TgYQlB5WrboK1xrRxVHPOCIA9UeRD6HmA6OU357hvqeSoGEj34aB
wlmf+KDN/lgJH+Bvzcp78Bn/Hy5K2UtyMSC9gYdv+jfQJBea6fiGxQU3vSY+WWut
WPpzP30iTQj5bV3r8/BpX37Ygv8YhIr8jQ9wGVih/mrBfVz3c9W2SU5+aJgNAB8Z
hmBSZpG2i4fLQolVCw0nnAwYVry7oVzIIySWaY83i1UB9j3sIbupXORAK6epsEuq
4u0B9w+al5s0pZSfj33Q4M+SKLc9eCBKPjWvAKRR9NeBThW4WevTR0UqTy4sQZX9
cF2wBHOg/w10MeyYpJ7tRPOIXq7XZErZVrg6G1ujgkk2vkdA+TwWOMpG3RzjU5lm
MpoddStZMpLzfQdfkTVJY2Fvm9D+UifzhComDand1l2xSDId22vAuFmRTQ8b2jIk
/pzQqtpsydLM2XcXwfhlCMHw2kpdDPrXpw9Jo1l9sPRy2vOVwh7Ro8t47vUkqZbY
opm7gqCKmlKMirtin6UzZxjuJV+shMgkMxlEJoduEiVvv1U7HUN5plBzJQfevwyT
t0MrAtCNdfRe+Ryt9QXeQppLZtBRmwJ4zerx0beUP1nP+TNx7uYbmh+wNEipU+bb
M3JdpYc+p1ixwBFe/f/8Yns+jkUXg0C9zn2vXoHz/L1odjyxNQgQ64eYeTxYy8jx
f3OO6FEvfywq8gmDtid1LO1czU/5dc3yT0edgwGedjabvMv7uPorsWNOfyVdAcDF
EtI2L7qBXc4Ww/n08pmT5+gmTs8v5doe/XvcTCYx9qbIcGZ7KxdL54L3yp3I9Tpu
BEPnID01uAtOuiej8ATZzTgMi9FAuUHpTReGoGHpFOxIPd5PniZy2v6bc/bt36uB
YU3ayQaZVw9y1pD+tSX7A+a/qPjfsSHwXfpvC3udxz4Zlt/brBo5Lpbg15XLt68/
IZBvHQxbbyfp+Bg6K5HSURdgszBayNQXZGA/j3UInetz2RgQKiFio0Oos2i4E5P2
m78W5QTiUs1QfHe/D2yKPZ8NbNQofrhbvofGjN2he4fE3NsHeGyz+lt42aE3DYpr
FnTBnUc+VeUONXtK8gflGmHzGieB6maSmBsc8ppV5MR2R0I1nvr+MuCwJIs3fqEC
y12eBGQCaESj25XiwgRTd0bdHs8mchX4QNCDt4J3DMzLim2jhV1DwuMel3nlj0iw
nBzR2P85dJVvstU0nDEKgWWQhXQ+AcKvvrdvTQ+NCfkugQSyOcxcecoC7+Pniodt
gFNZtz53tsZHD0FG61UPH6jnoNYwabQsZWeYLnUIVTLpinRVJCNTNCRYVfZKLwvR
Q0ybKaJK0z0nstixDlTevNeo1yRJrORBBDkGwNAaLpxsNkun3zlSX0CLIIqEKYLu
Kzo2QCsP5sxlENklSnxzsCiPFUoOdUMDjk2lhMrQZf//XxYDgv2XyGIOFT/slP35
q12bkvat2Rcg2aVVGkBOkr3GheIpiCZN+fcsio2GbvX9BS4Po/DC3NZOxS+7luzK
BcL/JDZd6LRBcXK4RvEF9j6mr4wg5lP+p0htpew3iHvblx3Qj14+KLNAidFigJlp
Nr+/VqsHiN7GW8FKELcYVvC5Sq+S9X4oY/5/w9KmCNCxfxzNW3qDXbUqU5KUL9Lo
xqGgHyUYYJgytJWvMBW2akYy8k1CCWx3QXBvJYZRa/R6V5jNQGwwdxIqwK+oxiGt
rff2wrZ9u/Uwr0nQKEDZdlh5o6u9O2VLCrmwFqYU2nTPvFXoVhyC+Dfe7WPHLuP5
u+WaXcDmzNo3VQQapcfGZrheDa87Ld7rGbAs/WQhgJRfaaDGi/QsxjVZuOixZ0Ie
9BeRlaF5hjHgOcWDJZu922uU5bgMHtUXQ/rJW01pzDrgncP3XJStW+bLIOQEVnTt
xGEBFkHTxAUc8P4CN3kO3F/q7Uq3oKdHFVu/Q+YUx9f9MkZqHel1xTYABeRCBHQr
S8RV7BXSNM33HDS0DuVRhyc10UlxsFqYz3gjB1fMx/jEHxawt9oibPg4/9ToCG5N
kTgzRq4Yz3jcyfjuTy7n4hxLj7dZBdxjvUB5dE5OTWldoXEsalAyuxHgB+/w4EGh
yx8DyhEGdycZpwcXXGI72iIjqATFY9Sul4OuMyFel3OvzXddO2zuim11qu3Te7G8
G8k7Md0/u1TA/enuNjv2t/pVXAlsNQTbBBYLNyHfXmMh/1uC4KS0ZaeldGEoSCAs
mVD6wV2V3CDYY861lT/hF8jASk66WnF0tDdzQw2PnMsKDIFivRheMIgO0K2o1RpE
LprkAhluIdyOZlGO0G5BheZERIa2Ys9o/KBC9l45gEdRVf/OGGQHPuYoh4RCYqqR
YptXdbix+YzGM8CvXHB9yEZMJ2NYuLlgOBZ/z6PAjXugLZtcXCQqpM2RPZgIEktb
mtdivJuo9hlxWREzQUKEeoZhCNnQZHRgO3QzhSqs2gqscpOijYnq8Sj8syeKZmLM
Zq0bQjJ3BhDi9jHKgCEdRWe8d8/fPeTte1msoFSItjJbR+2L/6yrmvrVuqO8oZdE
Ue6Qlj5KEuoahm4g0tjfz+wmq5+oZpyK+tOFouc9CbplEJuc5WaDBvcE0c64VEtr
aRlEH5eKiq6GFtZuuDNyvIgFu+KOeSbzqanRaGKJu0Ff8gvh00C7rD6+Chu15B74
Atid52bkSu2CvL8G9wzb0GjqI3zh3xOrJriYKdKrqaWyLJ9K3vds7QC5lCitzvju
0s2+fsxamclILaZYVL/MTUof6pvhfSt3nvzJSmHWVjUbJTZe6hiMLLcxLxe0XFwm
shWf8Mivq4mKUkNsMUXMgi7DshXyiB+JYm7qgSnwAs9zL+8iHMQcdl2sMIyr8+cs
ME2yzUbfYS3+gbVYq+WAwL6v2+LUQPy7eMYpN+r5gwDIuZwVbp4s/EWGyOrJMzL1
q8ZqTOvWg+3xs+pLhTMNEvVnrWfGuncIYZESe78F236r9jrQv/jPz2mFiA0kLjz1
4PnYfvmjYFskwrRWPOFm46vud6HJlRAMK8cubjEZmudwmdHFVQKDuKDfdGMZc/+M
Kj7EIMqWrjISxNzDuXj4DSamHmn6mqzIq1MIMkcayOyehqleH3vI8sn2JMj3XKzx
n2UoltS3530EBRXjcNK9PylbyQO+XU1RXE8ohqx1D59fOMF8uto5ZDtBcedWgbxq
IiPU+bb7PUldQ3KLZTRr+5Co1H5+iRd1e6CnhgE3TU8Y0EB/jdVtOxaArTbVzF55
wcrQBPm2BJoMGM7pGYxEvAz6TBowGZI1QIZK7b7QSn/8TFb+n/fDw+Nmzhfhqw3q
gURJVgRLLuW52mGO63IltOjiwAs8ApxvVJwlOZbHZs7+Le/e7YqlTnTeG8rAKyrn
Qi9/mAXnI2gO49DYPSGxRUi/M7r2saAiXek0/f/TRGlxZLwaVUeS495aoVKSFDHI
dY/hFYQHt3S/LPQ4Cob6aYjpUtybF6cm0e79kpIN3PTld4nGFIM+NvV7xKY5QvZj
12nPyMtBWHp0VcyMt98vUey/+Sht+L9f6xSWDwr7AKKc+n3P1+YYM3gkklGQZ7NH
Hdd3rb4XmEIKZFqu6pXwZ4Sdvjrgl5BWUhyTxjrMQ5JxT58XpZzMO/9fr5OGqTv7
CH0eefNcJu38aTNlQjQie0WkHA/U6IIv2KimOXGpq0hZ/zD779XjMcJPrr+nEe5r
SJhFQg3YZ/215n5g0ssuNpJ9S+25lwlJ9JhXNA4ZoarEn+JctWlzatOVchV7PDYD
itf2hlLK5f5xbqVZB1i88WpDc1eVdHgTh3bFQyUlWY9E5rm8VE0D18rhVu7up+vC
3Nu+d7ZJaHbcvuK4EP6ObuWbIZjgnZzT855E+Nu+/QVOBUEBiz02d/9VqehMB57i
srMtl2k/9eEALoLqwI0jWNTKwYmtkYRFj/IDqqWAWC5dhPsb0boR+VYJ6fOled+F
uaP8YiQbDwonkWXbs4h8irWAeRB6gCD3418uo5HlcCHzeZRzwJ4zpGWdX9UQAK41
qfitXcZiYk2oovq/2McInLXh654zMCa3J8p6vz7iqonPwpxVUqQNaIKP5Y9HFsW2
sqaOktD/NYDqiTpX5YQs2GaVSa2lR7XgDs/gPVfJ7/CATW+iFksrl45NaO8vl1dS
omqdhm2cQKNMyAFVVoxhgE+rGh7E7kiw9xDLPplYJLPyPa0yT2fA3FEeBT8B7TT5
IQ4IvHqGRafUhM80wGv1N6/qNrpWf/0NsB3/SAxGe5/+/GWeybRgESFhlnEw1mP2
Z03uQUdLaOYIiEkiaxbvnZ6V0PjBhYBoFfSgvCyFZxBBDUIEMQyivsJU2otcuEYX
ceH2VQvyRGqZ/J92Oh24A0V+3kUr6lBytgVXjH4KbK5rBGiDORm7VnteKTPIm11J
CmPmDEJp7Di4TyrC0WD4MnvgMrNYLnPfLXkdB8esWYriXUr4A2P+GlIkd3TDWuvW
oKC2kXpnM2F9So2Ai8G3Jm6yGAlsaEAjpguGC6Qhw01pagrfxt+A6Q+IO8z4iuR0
jR6+b/qW8cIFWDF5HtwgY+mQqp1BKbaHezsW13Xr9nee8cOpaVvt8kOqhp3/+Za0
ln1ZrOlG7Yh4LZjNZpEJ5WvMRlt+mkqFt7FKJAM5baX836v3An/LmtrBIF6NGHJn
BYtpDmF34jowDW7eTYZ2Dys8GcAE/WTHbXSAizKkAKKhUYRineoNr25GP7EI6jGv
vo+tVTB9uX+x3qLDL1SD90Bo0q1JcPB9O+XiS6d3oHh6YB2YxFYU3h79Pe1ukaU2
LJofGm7kNYYl9dhKKb4aDShdkfGwlWMIb6D3Vqw0uBMsFO0SM+iiaDHpbfjVFeWm
WatytMbf+qxC4ABrI4SAurm9o+fhBz8Z6T23jdC8sg3KwirJ7Fxg7AY1ir/Fq3vo
pPTbBjCN7Bpm2heLItf5oZLnGFEDqpP5CsbW6wkj6XZlAkERP26+R6aCXX+E05oE
mQOxWmg5MmYbcdeJfgVO7rlDKZ0AeGTwM1mtTA4J87ezKRKAyFwy4m2ZJaQdTZ4t
1iR29iHoo4uBPrfEmOc8AuVIEAj7/i4o5MRYe2X6ddUqtq7YAwmFGLzXEQLZJHXM
/matd/VmHUeOiMfClSh6ozPJ2Xos6SZO+REbfPurZ4DdLWa5L0RzJUbVpruv7AWu
k5hNF1e8RnXn4mg+wydSh1wW+M/wIGm+QG1gL0KvbisROQVlrgTNE6KmEtL+Ev22
fgji2JEfroT5EdwXdncprlLduheGQF9tQk+fksTuhxC9veVOkemZ4Tq4RZh2x51D
tOPxPj6TWlBKFSYwLtSvbO0d6MhD2eS1GfxoZbkTAXYPnCeTVYjw5VWQOB8D47W/
AiZ/719XQTXd7OEy+0qEhM+/lxvqs3/H5McbL90u+PevDYnl10yimx+gq06DAqW8
SSYktW95DaitNuoHZa69MganA6kFqPeBx3IUFufzzZatYWv6i3PefbfAq26uDzyK
bMoX8bzh1PKRvh7bAFsRS9mNMG1hZC9dU1wbiT/zCWWDQ+2GmlaXSCEK7JUqZSAs
bYuh0RSeu8xkB/pQLaGzDPhU2L3osSb0wpviVIelJq5U871eqfc54D/kMldZoWnC
bQEuGchpO/jBhGQfUsGLoUoWWXPJCfOsKc8CYokabfP14lPBY+nDLSBmxC+9L18h
eTg3U8qr2WziilziG722O46vTRHKBZiN3WWytHMAW8+JdIUR2PWmMmDiPJG9xM/+
PWJfdLZpBqsjThmVYYpXRzx80YXvsxgZd5iwaC1cISrdDlkKiic6eVrCWgb7hDRJ
cLJoqAJNdSo4ouaD3ZWCUpnsGoonzu+GwWB+z+W4E/bQgFGKRV7AltaZpXKEWFGG
25ICzY4boU3nKHHbH7F8jMc/pBKjCd1hPWpG+Pk5GPFDAIeeKshI+0z/D54qfYdQ
frjYLc19OnsMbgVCsB+mMyLSj72KI8DYbPgTZOzm2VsXh7WFUUwzWL/pzyNzOdgD
Q+Y4dKapCPvc0hc/42qgvmm0nEtG5HzTbLOCFgDwXa0LFFn0uYEkmeZw6RqT3jhX
h638CzsBCEibmuqq3Tf8rA35eNcb8ylCayOQ6t/CXNcUP+viOd/JlDq1+oTx9TgE
1xu+NqBWNNcvCqoPJQ7k7zIC9jWFrr5iCKBtnoEAfmaTe9BU4z2J/cs4fruJI0bx
Bq/tEtVNlimf0nIsdjGssg/pAdyZ5vRNh43JqoIDCTdqPFyTjefn5tIbZU+mcajg
IqL28vEz4HMOWkDMHQYOLl1r4CBVSIuwTSU+AIG3XPgeemP2zUqfNIFebaf2k4PY
kmQAhRDkGzVnIJdMqv792lYWmzxiYoOMjByu/1jIs/wdjmpmUrcPZQlpIBYikO6W
J0iDqbun2bdhk16otppTT42l1M0ZBFtoFTCyGyRQ2p5u1ZPtNdLzvhCYjKPe4QvT
FSxVbfHkcVS37SLZJ2MsF2ciSAyBlncdZ1X9FVP7ND4nDl5KVct8ogNwOjbZsgNK
m9VclA0Tt70NGmx54/1/K+MvArx4G2azosowM8CrpXamvHftRjbD21DXti3lxMra
MuOYdE2m9X36LCyu+4audNRt6b+nG5s40flf3TZ6Lq82kFn736y4KnfnPa4kOdVZ
q2YLCc3UPYO6bVh1L9KwUchkloCV8IIUPl0uE4yVzcw9VsNePCSuDtY22Guaw/9+
3mP85R09SG3yb+m/1wH4t26Mb7OXiB8kVWdfMddVNk67ykfnuSZ6ORvCaGQupTse
DEcvNBKNftJ07ZQFJcUWaALroAZe6EZoHJsUHBFudOV1ZbGGmwRvkPIYWySByS1m
Hh3++6ZTd7DdtlMTIqO7ublz6197iTLtUNmjhzSqr+b7KDYDRs76YUh1KFJyEffC
Grys500CdvbFi1OcjSLek5N275PiBh7nHnKn3OcWjb3tYVahutlQ3+42rid/J6y5
7OAYszqUkBmuIwcK0IU50QRxPyfS+YUanrrjG3jKMOGbzuH+Ysx1WCtPAE5TtXMS
i1RrP9pk6p18iRGNOD0p5FPqi8RvWxvSjMdfPtIxrm2mb/WBweUruV1VPfYWd02L
Tb3KZo3nfJhHeyKnqd+Mxn1OIv/5YGdzW3TDnJsOE7GtRovI61ntXxpGgnNQIzv1
JE5X9SlmXILb8nVUdSTDLAzJKEAoVKL7Vwpi4kSTypWa12hjIb3uSVEt57OxHNWO
uE/Af9CMsJzgYOsJznHRV1FGCt3qWtvoVdH+C7KoV2NqFgrCIcUXdlc32+T2tlOK
e/N2Yi57xgcevIw5/+8M6XzNibenKRnE8UOBWitXESuInMf43IkWRfzgW/4iLdAE
oXdrzctHUmjj8zu96JVzhAQgpmsNFy/fe8qCMFmQfSY5MrXZhVSVl/t2kcCgsJkY
qihUpbZ2VH+OIagyQEnq4je5XHjt0SdH/mWUSDz9ribkcJl99z97e71UAQazDYgv
zht47Yvcg+tgskG51ctnR9G3csk/3UwTZCw/SYuO4UcjQD8J/ND2LbXC3xuw29zm
xDXQhGoAXMZYoDthxsxcKudf0XDileulD1q15xJp72SeFPFs3OYb00QBzjXtdQJn
Wn6sCpAQ57oFGLghItTjX8zAVkkOyJnwF9+PeFO1flKOcajejFSq+1dNI5CxDpqz
V9o9OvRPaSb15524ZunJKW3ajhRaXJCZVcQE23VtonX/gISceN4+vLVWniC7zO+e
wzvAREu4yHM5siND2ZEsuO3ttmM137Uvle5/XiQr1XP60ZBvs7ooFHhodm4QUnxs
6UPbPY3kMhYjfVLeoBd76D+a7LlnhhoaQ3kKWHYAF03mFfCk4EF6YcYjSbBq6iAD
qYNa7e/0WJ8gVAyoOztf16lwjr/xKew3olrmMTVpRb2M8rb+T2sK0yI3hws1wbWN
IXtP+zt8Pu5eXm63gkqbMBZvtNbgrSE8ojm1tUCHfosOpBm4xCdzUFHmG+1U6gK4
3C5rTsNnG6+unjsTUksgZKI3w4ulv65L07oJmVOdcmcXK8ghIWw7mrpm2UJJ8KAY
fevevphl685D60KmqBeRW/yxbvrS25u3botmdC+ruPLwnaUAgEPiUlGT8K3OeDj0
AeOH1kG7wgLG4DZ//wlCxVFtD+Pn7qTcYm5TrCDQOT5AIlBsfeXuteeNNd59QsZf
3DXGRudm+fWmfLQYwRyMV8aL37Ytsd7Q5cUNdZza6RA+ffW7t4f6CJDwHwX94X3H
2564GN+AZlprNgdQd0Im5r3SPWjKRRCSrnlfuB9oNCcDJQec/YiXaca9QhnMJE7K
aViXRwEMnxyanC8/ADoDqJ07M1FMZeenub2K82SVXBcZtQi+VLg8hQko7Co2lSsS
q3tCv2d2dzAd5wF1EUV6sOKTzcMv+eT/sdYf5YVBI0sS6v9OnKVjf/2MxmI9g63c
HKIik3M6Mf5hy2mai6epVe1m39//VXz0K+IVXjRQCaOwIFpAvgYVV70YID+5KkMO
kM2PByZk0CL7Jxui4pNcZqIPSYm0P8TaW+Bn0erKL2jTg+AUWldBBz8gOtrYIENm
X/Moxerx7aHvd7GgfVEFC/DhXz1rboiCAJuV3wZkeGzN9QtZ/C3UznxiIsCeFQhl
+V36ljTmayjMqPw0fplpv8zSWUhBSb1Ff4i28tOm/bcZLPzxEvu3OqD2nKeVV/5j
gqFuJHo1ReZOkX7JOC3xO6GBFV9stpKWQSD5/VpbD0JlTuPoeLSHNxaNwKwo3JrQ
bxMEi2HH4KyslePqcOUviKseaNktItjpst6LuUBGNpTDjJADACTxtp0SwoeDKmDu
5T3AbjBLeBslm5l1P+A7GyhTrnh4miId0M+Q8RIuCLeGUvOxe7ax+mlkYrM0Gn8M
qO/jgOWvBNS5KK70HztDDrtZpA+Vew6POwjlO1I/AA+nOcebbnHan/cjBnpDnLVv
J752H5i5aX5YxCtgaXZfBVV3YqZiwjt3VbvY0vJNYq6YosnsIWHNGVPrQ36/qHy0
LpXLG4yvvM5fWJkjB8Zsjy+ov4pXTGKjZLVfzwWT9ioc60CC5SPoZc7PKFub2txD
5qIV9A/uHy23yM0udq/jD8Mm787/AHXVSZnzCOrzZ8ya9KlL4w1r/ME/2NPtmazj
WF18wG8BupXHZI2NwqY/It+20cuWSdE2nz6ZI5TeYzaF88/3tuP/3vK1KonUV3y2
6Zs4JPpuG/l8QoB8TuP55zSetnTTT41nFi1rmJDpY/kefq8zh5CBs0d8v/D4+THt
EO2lVIeU/fgAENnJOzX/ZUn1V1vj298/+v2XyPaYNfGlflDUGc0iKC3EPe+xhMyD
2TIGZTznlpUdT35Z1WZLNOyB4itRMxrerWbiXxfzz0AoKnZE7SH4BhNT/SPqcw0a
DbdWUybiXlR/jd6huxa/FxkMDilTfk9BTjYr0Sw9OzAtOvNHU8QBXPdDYr58goUj
3N43VdoTQw8d8Yf1brZ/T0C71dpSpjKo1polJDA+XnwHNSiwKHoOPP0Hysr0V+ve
pjcPkeMsYqeaxVPiS8jGF+eaPukgFiISse6kccP4uDWYkT6LO1Owrlao8kblQ+FA
YnM8AYm+MAbPBcF61gP2mACNvNbGqjxnM7ToSxODHUB+h60FyPF0HhxsTMxyMqXJ
51scyCOjQSxJW5HvKsQGyi8D46SotmLAMjWEF+0CRpQFb8q2N+UBSpdrGBlHApNu
RxomOpunQJ7hUJ856iiDcyn+Yhqy6V9PRtYRwlXNh8Q7m8cu0eh/pzy+7gRYIGSF
gyH/KbBua1If5DQgo4gzzSlIOpinRCVY8QG9e4q8pxWLrw30FKFnDmc4WqIqUP4A
FVotBMpJnTtfKNB7rE9+JSD7WXWMwbwDSzVMOpbwNdWypdgjaf5IwdhU40xNxTAt
kyPWa8WO633hUX/Qb6QqXzt5ieVYvngmFHSjTVz6ixyJhAwYJiXA+oozm12EG8ae
X2Di8CDXCbd1kSfZzVQQesmV70meYt3ORvYT7HslueuZEzdk+i+/npTCCNavjemy
xzrnIAAZUH4Bjwy3F8FARAgV414dOuK1/7VqdbJl0ohoHwqxWkpHIWNnEDzuX+jT
cPjAyLzuFw7beSWCKfJ2uRq1viHVY4r8VUJRyMx82mPIIOoF8Ro0utaEu9HKWocq
HQ0gOM/+40ghCckmnkBF4NGiwYf8EcKi0D5/fU7L6ySCQX6MAmgQ9wRZzkOoWT+N
6HlovM48ALY+gVNI5QvPrgfSDAMRYajcPcGS/7j1kSVixaMBYgItsuMhMTc+BvWg
W2uSavhOWsfNhKhcampVpOB75C+D9d0j4bcY1U29Eek98Tvg6JIb6cdzv27tpBAk
q2YOHDJKRSrRa9Tnbx33a2J3xrCtT/UwfT2lREZ/aBeNA1WQAv/sFsUhXGcylqC+
cnjiO7bTAlwqxrbCUhnmouTm/2zeRs++l/gz/kQtoT9Zukyfywg8eslUE2vR+dOX
ScgxGjmbFHzweqlYvlbHwWtuk4xz6zE1LFBB2oJ19XLe2kERmV8RHCSt7JMANWG+
GUHbCrGQVYuRavTeH7cwUUtutHt4Kfco+rbDe2nd5qtHUHW2q+ZAOMqXpSZau6me
A6h3xNLrlhizz8LcwE+0wfhv3+IyDQ1Hv1KFGa45mPlAyMuslKwhO44ybe+Ub9Ba
GjdpQagdu3v6He118RY+m/Dw/T5z4srz5vRBpZOa444Meu/dUTWCZBUz6wbjsjb9
PwuOuMq2Wiy3fUz8S65w7EJeWAICxwuxYZw4HFZcs7mE4OjhVJlIcpfiEURgMZWU
xWYJwHRDEBR5YpL02J8Uh8cG6PnpaBIDVbqSofJScou+MLExDuKq1GXXPvMO+dH0
L8DekxJM9ckG0zH/ZXUNdY7i0ue3B7wjPow3bAVpqC55WXaoXmNc8Ut/zxBqm7Ny
G+6k0hoYpU4Nb+6iGt7t95NCBw/oyaMiCaz9nAZ2hN4+Udq/c3WA97RAc6Vr0+7u
Bs3ZZ5faHGz3zHsWBYPDyeMF+NJeI4p8AC7zdHy+WI9mu6/bhxR1x+31FqMAOEFC
vg82TBb+hbTuvcdq1OyfE3WIFaR/+auE6on1iUacIa1afkoadsltE7FteRYH1ph/
ODjUe9uMEpSZjLlW+DvUv1tIncGvYkkpbSnKUKUkZIK/7saakmZ5LX0wZ/X32K8z
2iypHIXiw20p6FUOqLpMkWMvplE+63Bkr4+UJ5QfK0fhK7KLMHFjuWYYnlG85VXX
aClUYFG2o/0C+57TPCF8LV4zyfGxnSKaFKrsN9i2tXZJubq+unZPCs3yHApOSYhs
rvTsy616goEFvK5eOH8X4zYpXtbr7V/1YxXI/ogp0HBPEKxfeppPsO4wtu/XOYBb
67uoqOQjnMchXkdlul0+Nvvwa9aELz+lLk5ck/W9zGCayVOt+RWaHySb6P0Cp/R4
gl97VQPvpT3pHkVSEXJE9GW7s/gGqC5rsii1t52qy5F0SaH+xKuavJaWgtG/X4wM
eb51g4z08SZhcNc909pWYL0UJuOjHbuJ6x53KcdKZwpklnTq5/8kyT18nmvspwB5
ky3UEamGkF7CEGJetzZEQfNoHYnZCyTYChSxo89tIqrYgu/0IpJEFdXt/8BujJjL
+Ct+Tp+p5hS6TKQWVs3GWizWYdDMHyteCYZeRplmOQr1RKZJ2o7bCX4wX98/iuKg
6jMCIs0bEPRIwJMc6wWnIT8wIq2Zyw3c0R7M76sIZdKAwv1snI3qDHwa5F7SZyt/
eE1dMpQ3vv8BwBVUzH22vWasLKxnBAXBQgMKAIpNYaq5odqxuE7DviQ3eRuxb7J+
yIPtsGXOT8f/Btt8Cx2VlvnQvs1DgP2K9iPq9h+H7E4NgGzeif3U3eWWqyUEHVc1
wuUgHvQn/J2N2Sao6nivEOOdBPzFeuvG5PSJixOTN5Anjr0ETLCegCk6g2A9BJHb
BeILLdYf5q5DsfWuFAfi17RfKwTEN/Uza6B/Zs4lR8Aabd5izV/G2+vjlhfbv2aK
u08VGsQOZkFmCBjCUxG9RIdEi4ylp81vmtxlqR8WwpJD/LUmNwh7kfdxysWyiTS4
/X28avE0mOi0CuCD0IANsg7aNBMX2XwosfuE2aamS+HhGS5jWcjgC5Ci9We4rQYI
Kv3Wb5s/6sfpc3G7UGbhWtYMrTD6X7n2S+Xy7bltXqFuGg00ZDNKTB7IUzxGE9eR
fQc3h9iSH0lsu8PizYBvtpYfNv8r4bVitNDZXMVHoiCDYPu4gnfybqe5mg8T67te
ZmuVtbWyMMHdlstE1JkR3lPxVUon8q8iIkPfjCeShpicgopcOWojtnOxG2mNMlwk
rkqdzxzmFwN96byQGQvovFXPPAVCkFuHp3KbkevSVyZ/FJVBhe5L60FYSCEPzJrQ
I+zkKDgFwqFYmUC1KqOmsowBtjyBBFvq1dbExKVJJlGgQy5He2h9mjUzFiyai2q7
InQkjrN8lohGkLVqKkNJ6McXKYmhrqmMGjOfj7pfMcj6WZd5JMgeRIxKCTH5TiRc
MBBRzUwoxc+r757quvM/6YjNH/lnmXVjLY3gE9aM8GyMdK8UNIcKcAhNXGlah8yM
UwOf0JLeoyVoa0+GMZcnIOfybYzeOdcQDRYTzoTfS5weU+wakCn2qnLUlz5gbVAH
acRjz5tVg6CeaILtKPcZY6SGlsPVI50054HUGGIKc+epCR5+sU4VO/926/cfI4Cx
1NQtOY2kuvmi60tQUgnhaCPouEugTrhgbw6qyep/vxVSuayk9TFMOAkgKKny0e6d
1gKcXDIHWOfAxJVdekpmH2jcE248KMjCREpUTpX90hTlOjbsKdaSGUwh23k2iWgB
7MBNyyrXj8eIWoyH4ZHIJ/qSs1VuwPnUjIP29YWpxLrVYlJCxv2QuB6uBzKPmRjl
4VYVmsLLSY8j/cuRVxh7C2W0FJmxoFywKBO8GPUgWUaMCrLMLie+A0FV+hlQQYdf
Q10Bz6pza7W1Ax6v1EGaYLqHzVS4EX+CKe00wgmsDjaa1vZQHy+b0UNsDN/n+My5
//ZDRZyanM47AaNApdPLZ/C63GnrAF89S5ZnSLKkwlrJQj8PBZRIzZP7JwIiGeQR
KAm01tgO46Xv0HG3sg8eVv9JUTS5mcidbmVq9xI3tCKWGFr7Tj4w905GpDqgFMm4
dYe3CLWy3JCMQrXFSuxR5biKhODgO+HmFwerxoAd7iQxSWWoUh/4jvDIsl6QijWs
7LXHmIjUFJhSo/6LdLej+7ix3nUMcIqjyzaNbL+12TKgUQmi3f+12HbozEKE2dAA
jGLLZffnSFBBwh6XnVUjh1wZhMuWiCr8MemGAOpDL5xklzxte3kNUARBjOkNkJdV
UKENUmZmUJjeb3Ifx5MriGTHM21yKJWEQ4tlHQzUq7Pt5QIuwMxfUFCAv6qhXknq
ntXE+vh3qC4iTISwjiOFtir5UcwFS0cb0nUalbuP6DcR5gKtMCYiUTr1ZC0at0lt
OFN5E3VjAM+EOQb2fPpRwumemdXUqPdfB1CCTxurn7v39okuKqB/dPTqPi+zYZ04
m6a1PP8gMeghqaA3ZxdBxF8BjP4IbK0Xz25fHxbPDyFxujYeAIzhaVfBBVFbl99T
AAuTlGd4i+cWX4zoMot+IY+CrMEg1Tp04hk3p3DzrY4I0gKIBWa9BzFnOvzY82hc
EU1E7tiyDCV70E7l+IDKzazW/FlkjxpfGJ5a2fjyEl0rTy5xYmmt5Yvc4PIZPMZX
Qj6nWsdnY9hAUWeo8ZOqRwgP19o16r8/HXde9opc55sTkNdjpIx/Jeih3pQWvy4X
NJ6cj5GDc8VkYaz/M3XhbgroNFBdJx7CJaRQd1hiId3bWscWizMbn30e76IBx+Bp
jO65IedGEoBhdp62QZF9fD5g2ouK2M5OGe4N0gwtgB52sCSbrb9JdI5TCJrsNXp1
a0Z1k/pZ01gOHt7S5NcnCYXne0r11zPhLglQKZOd8v3h8jqvt+5BwB2Qm5WtEWjz
wbAdCeAvV7gi5OhQQyZMCWV2TgCUR7L+YcFmCoXnpk9JXNq7aMC3qbFcs+haPoKA
9sdI/UscUqAZayocEFbIgXYU/q+6jRHDiFtAihuRP0grPLvrQq+iwlAw+FRBTJjI
qY8OpZkdsdpHV/+mVsrCOyd+3bOrf84fT31lL7/RqEdZ69G53hn/barlxFqNTRhA
T9q0frI/HPJJZFdrRUwEjOUAPbNs9HyKNa4C6i0K4RiQofENZcBwdE6ZDRxg1ug3
F+IG8MVQDO80rJmuqZ8DXBkojcul686J2Q2EjKGniqMgF+K0Muavg/K4M8hkDtji
pxYx8eePVWMKixJv/IxjWx9FHcJTztxaI2LRa7oBxWhrnIxJTFR8N6Ix3W3TG45/
u5wau25fn4F7y9iSgdiVVQOP8/KKN9WRpYs14uMnCvQx4ObXsCj8JHUgzSfbJIf4
zT05/adUl1m0kRQr2EPXMG8u+CW/PkGvMV00xqBF5Cv11N0j79FtYbaaLVbsaclu
jcjSicNOtslngM7b907GBvGaDDFQaDVPXT1sxxS+E8/qJjMh3ICMHAFTzrVL6g0J
ZSrqZDtZxVEw3OppZ077Du1JpSZXUtfzuTLbu6aCCqtVQj/TYR8gw6Am1rHnDvji
fm3HqAuK4A9GEUG4AtJ0QmcvbZxmitm8turEcgeMW6UPcnLN+p7DSdaIC5g8c0V/
gQImJPF9IAy/8CBmJGVUQytbtmdj0n7U1cyVo6pkKSTbXs7Y6upbWtC9QRziKq4F
HAe45FnSPsnbJYV9VucOMjPVNfGX6a8v2f+DL5y4Cq8M8JcaDoY1d1zJT57s1Ko4
Ou3i0GXQa4CsqIMrKJb7X8SXg4/5mVfv8hi8CqiWfzozpKsWRscfXqluLiWetBCe
m5E7f4nf8vZRX97wfa8LVDTSPwzzIqMup166rs4YsOVVM219Z7/Flc1diFJRLoB8
bkwka71yqLRCCGQlPkcGluHwgD5X3+xBru/VwxgRfjc+4iz2nnitj4lVT0cfIRvg
xL+coECGOFJj8/zh5dp1XHP75OX5WQqJGyVbFpiTi7J4Tm9C+kEdGMLWfo0jXv5y
hcQmBIVofsCOEgj5PV+wC7bc/LF3ReAttAq9OE/jvsy2hhoFr7PlO3fnqrR1AmgX
/eWTDwJXxUzFM5oI3XBqpmnTY3+LKez0Fi866ByzHc8eymF4GWTYXD4VVirDInon
uKjlVOeDjaEA/fC7QdlnWPDTp3LBk5d4n6rT9Q2QM8Q+G0KnyI4fLP8LVxO70jC8
5TiaPq3T/jHcF+ExpB7lslc9lF/1sgAgB95ey55iQrZAL8Il/uowLXXg3Ae2/x4P
p1PkSsJdY4elWulzOGz3HpVvtt5ALYuPER+MtdBDUcz4GpnuUzRjzKNan5bswqrw
5Hwb6oS50qcbg6mu6NpgGBIH7NnYqWfeHQXOzA73pbVQIbNGYYBRkk/epzGFDYVR
w9FTxoii+DDl6EwE/NJhsYkzTMjCuDrzb1bA5U3eK29FnPnd8jkataXun23gQaLZ
GdZod+S9MkG7U1l6Y7JcIB0PANojnPLorYvr5NBITK0ZCaqxxohTs73Lo0pMS3Nb
odrFH3E2xSoqlFcjZ5uBCfkPYDs5u+URFRNcZq/5jUCDZY4IjlnVoqRgQI/5NEWG
lLMrkbH9FIqqBWmfjSV79xp2uKwZzQQbwdWkmL9ltyljO9FFiW8t6FLvAARGTnbK
LCiaSlJN7kl/7Es+xlp3Dxhjbuu/cY3YeSGXdOYlMr9SuadzMMMlg2rpQPEWfrqw
wQXOSSgYS5Lj20Alz0JurAmh7Z0NQZzfwYjxpeS+ezy13D91d4L7+jmxSPkg7sgv
zRPVJKzCDCFVP9m+bheubxlc3HEGfps68+1FEmd/bf0JMcVVZLUrW2pjdfE52jfQ
HvUoIorxeZnT9hnvpltiCIuOpeIrguzMOHwk1GeTy9zSzDb6N/977s1yLGhDAVfB
gtqQ/KP0uXs/dNVxdwTk3kKJ04DV7UcSMTF/XwM5ugPfH8sW55HwrwkXeOtempwa
8roopRkKanQDUG3BgFzgc0SNDQKdiSYrNM/KUxicFKl5sbD5mJx/RT0iEiHlggfs
aF2iEISnNaeoFm7pspZaNjxj1x7YAR6CwVws0lulaPMPmKk7qrVxJmiz3Gef24VY
b0bTsNHUhlYQN/CKyFJ5OMpc9/ZMOBM2M/bmwYQ25qhJYVKkZt4vYxAR4c6UrrgJ
gF1YdKGVkEyjoTGlGAn9C2XKEu/GkGS16PO/ZF8cSaIvh4YBleqoRESxUphniRG+
VBe33zkLCsCA8hscl4msD2km5pQTs1iZWqKZ+oBp/NHb6o6pTexh0eTND7xNIPXW
4rxmOaKEMvs9Vzabsa0zRcZS6edYBec3FzTsupx1c3Iry+E4IQMAq0YN7E/7vgEh
2WXurhMB/i6pB0PXTQXmhsk38KTjE45UEvAOYVwVwu5H5uQc9VO8zaLEWq0SxfsP
F+3kvDOD7uFGLDk+hdoSPww8RQlf02WVeSkGB3e6LmSIBgR+K0fNAf4+WM5ud2CD
/jMTTfTt1BXk5fNB8ifOhjJyy4Pl2GlNh2kmpq1IEvK0/qAb+u9VujV3hk2tNkzL
GCdwxAPxGVrEBmX2g40ue/RgrkECiXHjOqutS4jstoHxCu2TYQy3YNJIQCuDYJGL
bWaLxXjsoNAE4gOYD96IW7P7QBX2747MW1Z3YsQZzW+MHi9e1gi9BYwoNG1KAUGR
bBiyDsyF/QguJwFmd3WJKZliKyz5PQimNTthh1A/QAMrnxoB3IMGMPysVE1yjoJd
ZWmNDiITppHL3CgmtwSR/pLmioghHrkigIGbXcAZkFz9IDzMfEh73hkWy/pW0G0s
zcwYAc6+BTBb9D8pP+3mU/4NjZYCuqQzqWC504gnzQ+9Apl0KCh1Pccoc2HfXc9a
6sy3Wy8hEMExrqY0PVx4NKn7Yci+HgfB5aPJ+/n9nfvu/u0ncpiTYS7rOdRI4Jf+
VPH1XXwFzXTn85IDUX9d1MvFZG4OJRThnr/7KbyuorT56t9GiqYW7o31jnRfZw5q
b8N1qqpgZfBTJkhualZODUPbZD6JVx4wKjhZ+IySDfAHm2Pa6kU2irnhBr8I33bT
zm/6DQCU2jt51/qKaXNOVjUjYNL8u5wA+bjI+aWFmJaeray+5zR3+0f053tmrWZR
czRoY8jzfmPm5RRvnksyz97gB5cwMzPxMJp3/4ktkXOxoIQXcMyT3j1waXGqelH+
F9YapkKcR1oQ1AybV0IA40UzKeYXvSrO5z8us2rBTJVM6DpaGSSLTDxZtN/lcWL0
e5jlJdCPbpuAvC2T0d+LkFyc0iwPseqw2zH/jsF7lHln2aJBI6UkySxvBKcls/Lr
Jby5UTbPhre8LxucXuVBRsVM19ef5TP/KGduRXj6J+CRojTQCyLj6MrLQLGpXE7Z
41p0UTqvZ+fDU9ZgQVcnUZGxxy2VeXL+Wg/hz63lTYz+FpDd9T7C6oWb4kKeEMCX
IFaF7QdG34urj3EqIQ8OHnLtK+0KHoa/vqBuSVzPc12J5N07GJvuil/b4xFa1IsN
umFpnlsbn8VVTHLOldGgfyYKscnfi9ntVfa5Otw96nxqTKvGGQsqzsYaMjGmr04s
JQLt38xKbhLjsXtPV+e0DgsU+pXRSiqViDxRfLqyfLLiq7W+Hh9uG9KRY3NT1mtQ
/hUBLKCEC2gmTMlP+8QW7lYqWAUIt4BjhIO0YuxQfBUWeYPiGo1Eoxi5WTRja7g3
KmvHyMieDb7x63ub19RHhBw0CYt5UehmbrwxhP7E8wufnfEB6ONug+zTzx4HVbgt
eSpSBBYYRHqZX4HquCV2qxE68v5RwWYQOZcyHPSKUJDg/Xxi+JdY7X6HhjAZU2s7
GlhiryhLwMlHrXoFtRdS8ZLAvkJNlwNdYgzKq+kvVhkAQIvG0P6ww/5cFMVdL+GH
+/x04qLrVaEXIwxU2qbh7q8mOUYCJ+SyzfhHnDT6IdZsvlLpmM9gmPdWFZEbaJmF
r/nEQ4XxOUSfZ5Dt49syF1Cl7Tho5hdBFU0RcPodT40pGBbO/jGOiE1obgIDziln
Leg7pPX1BnvNB07FrMBTVC8yNJUqqDyRP0OU255AdW2XUbwutPexH6dipPZZ+10+
bLNAIONuQLAnDbAyiRDzy2YOTmqWEgAjMm77nS3QvVSvjJdMppgEpx82BJlkGX8X
dkQl+6jose2MsGjLj8zkYxzcciPHqcmAhFHS3p4c+71wJjto6Umq+G0El07foKum
qGYxnqTzuoogm7gj6lHEEsoObVUonGjt5acUCi+K5ODZYZiaDlpMX17PILo5RCQ2
JoW2YQhyusmdD5BmlfQQFuNa3q8s68+obiUdfOt+Y1FSYBv288t2fPT6XtVVZJmG
WQpAwqYkPfphwSL/jI27jd1Lo2uVDc7Vn0/cIT2R0AaKtcuEZxvGLH4xlK9GDkNC
UKI1zTRS6Sl8YwGIH8qsvkaPSsqW8d+FoijrrsDFcfgDgHnbgSzAHJmKl7w1z56l
xQDvkVYIryfXaZeb0Kj0QJ827IDdK3aT+XT4jbvbuxpduH9GUKWiJPagWudnloZu
uDTdXxlt8zg/fMQuvze0UaKTXucYUv6MjDBQCs9eS9FE1doCJCWQryWxOe6JvL/5
dX6gMR1GrOpdIhxKeFpAOMLOhyGjaEA8uvgLrlnFbBLJFrdZ9ibxmby6hNixrQlS
v35Z5+qzW0TfE/qIGKX+rlZE8/rQOuZCc0DwLge6zvJTyDd3xa6ZPEf/Vq9lH306
UsJlqcqZOieYeIp6DjlDHzzKliuZUtUhuHzt1UYdHS/SS4wREWIRRaFLZqEUqloK
z+NzA1Hl0Eifc3HYsh99FhlZXVEVAhsFDWUYRfugsjyyFhXNC/y5MEE5aWvlUTZc
K9MVoVewJXx0PU/5ttmj1mqfZ9y9CwUf/ZS5CDUK535fDcZWj5fF6Z1o2ysnEbgc
IbiSqkKVW3RRteTr3XHxo5oXxvB7uF+9OeR0rBpxLkXN0U3D4LOTNUH/AG9sMMBW
194Ah0qqk3vjkDrVGEoMNrb5rgU6LyK20bfA5KnNQAUHw5Mz5/yej1PZnzpliflW
GaegQsVrvrT5jjPZ9AMrC1AYITvKpJdLyAsyy1tl8nF/mdjKw2Tw14qOgFEnSAxN
qs7gtlPbXcuRiZ4BJ7qMK0vnzFRusUniWfU8AFj//YwaEhDs/GUzQCAuSdDDPmUW
Ns7CdMhvBSOSQyxwYmHL4NFlR+5yKqgvvph87w159q7ZXLj0gm51TqdajzPrTLf4
sZYX8IKY7qChJ5S2n96hhcO/weatDcCGNIyvSu+EtntS9zEcf2QegA7vz/kbUlm0
sCyqHNGdGG8m35Qo9Mzik4DVSsJud8JEB0mc8iUp7opzF+gSi6wyuaAE3N4Hnse/
HJvg7xYeMhwoAtVEgRCL1HlLxMfSoPD0f77NNj42oxpd2aN/yLjPAeZL40ySXOfS
U3v3upV8CvegGtpwaRHmBai5a5t/mDYhrptcXc+T0rK5eRwDj/PXfeJMbWImD96p
AKYEiUU88/osRRHd/ypTxbNMF3Be7RW+4pjOtjUVPfN+5b/We1BGVEBaENKGjSW8
A86A2HCVhUSj7uuA4aSHXmTuB5UylhDsN6Q0J9DvGSBym2sTEREXVy3cxTc/gXvD
9/36IBplaefjT9zzOczHp4eofdCb9yCuKIn1il/ZrYW6nfX8p8tnLBf2rF93vFyg
8LTgXYaMFjZtoZiDlKBps9K0tHOEhTRQ5K+nF3tWV7GThC4PNaBNv6REvqoXNm2c
5VCAciygvWAhtsnW1VAsk995za7gMZRKn+ADJdJsnkL7wF8odqNznetsKRE6/QGv
5KYSp2ds2On7vPrJ+WSzhC16IJFOJse2XBuNuB4ngIe15RNeN5N91PccWtwFTj6n
59FIgq88H8ymbRjWRv0WbHFRmSfLAsucKNUWfO1si4lmuiXmSwKlaELNMph5mzoD
pZoVPLVrvpOMhudc+llLYuiKujJg5EdNcoM7ocySL8smmR/g6Jazzale4FJLypgw
fpX7C79/cCwZSOxzs6FHkiLr1Rj5b43GwlfNUnz4c7I+qz3G+s55SyiqXPI4smq+
tgT1vcE+mCueMGu1NkexKbyLo72+jQ/AOWZpuYfofppluTo/+sDpiGZFAJzv96JS
qy79FLDbZmKSSRegu94u6nXKZ5BNB57KX75Ci2AUYJM8OO1EKDTSh4FnV/Z+0PVp
Tfsiy5JTyGvcft36KqroT+o+k7DMLPVQkQR3XqCVg3fUZfGler4LngV43uMI0KFo
IYbnnMgHunwzB0XZ1ER4o2BJ+yYos8HlaYG6FTt9AM4n5LQYPKvkwqlg2yVjPFEX
OvgLfkbnIeH2u6M2Yf8H423weMrShlMgijHuU/dnH1ulFRRho0PhGPoU6eRPrtXG
IQjehvYSYLsTPQxIJB4+LEQ3QHHaK4sytEXalz+2pfliqwxXSIwbY3DsTgNXMQV+
OH2YlAVG9GbSZ7cdvv81+l671Ha+bwWskffPxEUe4A6SZ/8dPcBi54ACESne7phk
BMitXVdT1K8Jw3aVJtFwJFoGDGaX/3cWGs+V/gekhFf9z6MVFA2hyZoXFRkixPOu
ZNf6QfjlGdQMfjqUGeQJxhsVWJonHkxu6Nap5Ai/bORj13Uxxvny8pukyrYvSWMv
JAspML+3SVNO8cRxEjMLULWEoUlYGApeiCV2mBo8kYMKTegQFka0ArtRmV/mg/4Y
W9QQAO0k+rZ4Yni4p+zshON5kPCDarDlqVNRxM/knpOK/M6mxeA9FGQ56KgMl++t
5kL5rRbeMNmw50MZNcYLyej73KDESBkKSCs85ymnb828+1o8fnegK3nCoE/HUy6B
VB4O9PWtBgw2/tUcojDCixRYuF3v+z00kk5zEPM1QwGudeKY3O3CF2V01zPjd0n1
h0+2nzJhhmtgbBAJxLnaAr8SQ7Xws1P0IQ/JpqNqK4SsoECTb7MFigNnmFFCUOjn
9tQODAjry9iv+kfAz2JZRImAaCi/PeSaKjUqpxHrcaIET2ED0DW+2LvXrTZCA59x
mHLDNiGFIjGk8WjlHSLFPq0Tlei4EqoV1gPRFG98Q85qhCjaXRb9DmAHDA9KAWV1
7sKOZurhuJbPMbSg6s1Frtk3RduAF6ggTw3odZfPM/qv2+gVMMlFqSv5jnQGFa6+
oCvqfnoMLALZ/R7f5VkekJ5rkkSPwyZtyYyxlTm43DU3+QbYbInW/3VTMyFUgwUS
blnvrq67IiRdqexNXal+UwhrfcLxnk0Cu7CjrHqlWA3CVGCUxgLRNXSqNgX5cZLg
gAVVJePOzVoLb8gkVFS2J6SC5b7s9mg0hNth7EeLHq1eN7ZmxUZjggVb6BUuR1bv
VlKbK3xyCUsmpo4qDQEOwq99qPz9FhxUVIRALRZJhAHBwROYtyW+YtzHNC64ejZh
qQAgmeo+fLdsGQdzzQgRF181VtR1IxZaB62Bx7juaxGfZ29uil+/uTm3eUP26I0d
wfjAvoUII3ZC1OV45DMX+9Pa7cQjZ4Qd1Zy33gA/Ww9ooRKx1qfPOzV2JeD1hJJY
rx+kOz8bFRec8t73O9514j1A72YoqXqHkI6k/aAHyY7nPHYdMTW9QSkUaqwvv6gq
0+hrnlhd9eALSCbv/xoaRc+6yC3sGsppotRfCCvo6EU1mJh3EJ3KSCyXAfikr9qu
crNlLv0BzAuy3I98hURh+dR6un2huaFzCP19f0ghK7FX9HT3DznL2+zFiVv2wXmR
v0HvGnJF0TVZW6WScj6oxCj2IHffHVZ0mSs56dcCJw765NUfFYSxF66R9920joqb
XqBrXJcF9TPLHXp0QDMVG9eITANCDbx7TqU33ljOHskxVjbELLkVQ+Rv2nO/5vO7
SPoy5dQ0RRPjGuZ9N+KpmOtQmkXsT4CVCdHAi0U4Q1XVaQOTySHjT9busw3lrwjW
z9Q5RzVHH6k4nmoVQM3GbtRdO5a4EESaWLrlOHNIBotSv3bCNg+lLbE3sUP+0zwP
PLTWZOqh7frX5gVF0u7NAk1seWcWze3CLGa+Ltwvp+5+c7f6FX8Nl3SYHICWZWjv
LHokX70LPZDUaE3JDWHjkxTBrV3Lupnp4ujLqbmfJ85GTBAcrGbWqZvP2dz9+ohB
/uroYcHc7UhjLk4lwKH17wnr463Bd0cjEMPx25oU95Hkuuno8Tzq2wQeQAL5JPqN
`pragma protect end_protected
