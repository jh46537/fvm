��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�0�w׍��SΪ]�����E��>��顗���="�Ct�QJW�����j��I�����1��5\W�(����a$�Ή����F�#�jT��h	�,9�������H�O�;��̄���L��^�t��zm�s�o+��lb�Ze/?�8օ�V��6����:��c� �Þ=fy�t&[v'w���̿
�k9@�Nv:��I��9�}sUIĤ@��A�e�|��%G,7�Ȟ��;��O��=�R~�u�B
��6f��K+|���� s��O`�����A��m�a���R�1��)Z=[����;X��8�����E},���瑏�B�`6R�6=����Z)�1p"A���K�u����_�#�/KQ��
`^�!LV��k��\�e1��?�k<�}}�ė��ma+*ZC$���sM4`c��p��Ӫ�YE?�tL�EfPGX�yr`\l�W��彥 �h�90/
�Js��K�@待�	�P��q}V�n,C�1n������r��d�n���������&'�HV-wv�[_��V�n���@�>/�	s���<c7�(�������%��s��u�����Vt���+�$2��5`��r`�ċ��KOK�ՎM|닥K��6�g}�S,�	Ka�!�������O�g=���Y�"۵4�= �����9�m$<ߛW���+`��{�2��n=?��zYQ����
����'���sn�WT뎯��եL`�>��"/����Q�[�Y�5�vCXMj��}���ܿ%��/x2f�+_�jA#4��k�?$�^7�a�kW6p��ض$5 �U<LQ���x�=�&7E
�9��	d�"��H��͂�[�--���]A�"Zz��piDv�Y^�^O��Asq��y��ϩb����s� m� sMG���jo��H��+|�Y��ܑK>�d�4ܫ5��φ��_��hתƇ0"����/	�b�ٔ�Ƶ�O����<�����~`�������*�Z�h*���������F8#��v�����v��T��!�NGڰd�h�&�z([1
Pa�q^�4r�x�_��KtY���@�!�˘��ʄy�F-�f��w%��Qh��4T�	�,h�D<X>�6 Y0��}eD�;�Hr���K��7nʌw�v�Y���ߐG
 ��3vqk�����$U_h7������8��~���;z��{F =ۮ<�=d��o�sxU�\�| <:tY���P����u��������b�qT��F8�7g0�n����cL)���*����tQ����g^�-�D���Qwcd��b��l�n��NYhJ��.�G�����Dd�;����P�-A�#vrz�I'�b_�u�~��V9Nf�p��� <~nMa�p^��F,�m�&��͐:��Y�Fۦy���s�G-A��&�!���Y����E��)�F޻o&�O�qE�Jς>�G�{��dX���bB����DTN�3j|o�
ޱຊ(kT�;K'Q��'�@�=�/�Y�S�HN83z�IS'(�fkf��y��i�����->(��IO��3o%�zN,����0�F�0��i�Y�82�є�#'o�å��E����L��F9BςB�����T�l��d�%RUx�R\���%���J���ˬw�g��i�s5�Ʃ�ULt$Y(H+��84Y�q3����בT�~%���(�e����-�P#$%L�<HZ�yH#�K �\������/\�M��7��o0sVR����
��N	���J�?f���)uX��c��}�k�#|//�I�ZQc�^�b�C�����R�㞦�e
̔�\�:��sٌ� Rdy�!����J#�Z���B�x��5X��4tq����&�6!�(�MBil��)��eUƖ�b�ڹ��w"��8��������Y.�V�G5�������Z��Z�����n��2�����KQ��B\潞��t��~D7T/�b��u|�X�Z��.�S.���e�y�TA'PG��Ä��g��Z�#�!�W�j�����S�X��_�lQ`ff�#?�*z���C�!�6�dPwlͬ (1�"U4nn���׿&�� �\�3/�0�V��?������n^�ȫ��7����P��|9��&�(�c����Lϼ|��	��gZ�.�\7���(`�5�X̗FzS:fށ���M�м:y'�4R��8=�E�I{�kv��<;x��*�%w��R�+��Q��ߪ���I"Ja!O��@�^0�	�ԭj��'x2c�
�=�� �\6�wA{)T*�Y��v��^����w��7܎�~� ݹEz!T�S�yo����.�X���H�2�[
��1)� :���ChR߆�.�y��n�[U�&C�"6�������
�a�N�{;�{�Fo���L��<�׿��쾌K-Y1�Ϡ�t�[��q�Kul��&�yQ&r�U�7X
�x�
��![�O���+]}