��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���Ⓞ,B�$t�{����c�,�-��� k�4�	��[%��B�?���4��\������y�0ֻ4M��'��&[�A�2��~P �i�)Ԧ�%'A�R�t�t �*�?��v���Pu��G�� m��C�I3�_DF��(l��EO���Y��*��=�S�-W�Q����Ge�E+�>�ěz\����>s9��!�M!���m���ne�&()3�N| /׾r�ƙ��Sr9�`b�	���J�O¡B�J��WaK���2�����(��_C���q#g�sr>�@cF�S�]�"���qpRC�u]9�Q6�)_-Kҿ�3��6q�沿�E�<�����b�����  f�@{;ʰgLZ��x;r���
 �P��\B��"2�yP�#�]0w���
�%
�fE����=i�|�c]T�@l����Ẁ�N�/�(��Ѱy �
B��ќ��è��ā�/���g9x�!C/��P�U4���qł/��0ߢ���.����<��s�:QD����e��,KB��C��W|"n��\ӣ��]
z}7��K�|�)�	F�&!���e*8���f��'�� �fD'9%�5wk:�/j��q�?�/�̩�e���	�u���X�=��B�W5t������i�^�`���.����%�v�@�*��> �^9�kI��f�M߄2.e1�u�e��8ҸY��xw���>N��*w}N_�x{��V���=��9�J���]!	����(�o2����YBl���� �������KT`�#To�Gv��]�f��5%������P
u\Uk�m�چs-��EO�w�H�����Z�V�,���}gnخ���" �%���3&V�
]��]r��zt�b_(z��j/X��>Ϩ7D��Q�P����j��`sS���0Sl�U����d׵R��P�C�:O�<v�IF�b���]�R���bO���s�W�����m�>70
o���;_ǝ�L֟�2z���W�}���";	���� m\՛Ïu#*�:\��X|1u&�7���㝐ק�P���-)g���0x!��6l�EB��.�	/�I詏���L�v�ڂ\�i��z�}*�.U~�fa.�jdHn��Ր�� "aa�W�	AՃ�Z��S��Z��9���V�����))�o,3A�HF�Վh�^(��D".#�G�����A�0��p�T���x�|u_����񚤇�\�](��ؖE���$��h�b��~���S����;�K4A���Ӣ��N�*� �ulFs�B�L�E�g-���uT��c��!���D�����L�ʾ���j+�RĤ[��j�8��5�=���>^�J�=�,�6&�!��Y����Mj��׀���з�͞e���[k���$x�V�C���<{�b���c=-)&M𕹇�����
^�n;�5���\�oR������L�X�6���)܅�P\�%]\��q����  Aq�IKp��;��N���^�c�֌go��q��D"$��������+;�X,Q�@�4��X<�i����Q��
Щ�X�x��p�\��O;��5"�DQ��*���~*(�w`��JF��(Λu�a�<L��o�3�*rb�$^\$F\]�+����l���ҥ������@W�9�R;�w���3IyP��.W�җ�U~f US�g���yQ7�v`�zI�-����e#�v\ݐ��0O[��s2�u]��������g2���.Z{G��1CS�%@hI	׼ͮ��W.�P��{Jz��2���ں`�[o����ֹ�{sǠ{�%N�����ٿ{d����y�T��B�7��2��hQ&�)����;.t�ߘZ���a��|(��3ݧD��ܭ6P�@ꠓ��q�2nG����'�@	J����`u���⩚JNS"�T��xM �(h�ܱ�@�R�:�I�w]e�0Ѱ5���(z|��Bs�	�������9���i�z�}dmM��Eh˱�^�,}�&�(u_��_mGJ+���,'\h�9�۾�N#k�j�{L�kvS�a� �����+�Ĕ��Cjl�-Gh���8������F7M�V��^nW^�xD�B��x������D�,Z�Z�S�#�y\n��T�����$
^z�Ci�b�emnj�6Ay�#~��F���w�w���p�#R�v�*����n�v	���dY��S�֢��f�����6e8�y�	���(����6`�#޻/� z�����E����w�Y�"��4Iz)�3a O�����*��G��a6���������os��"��Ԓ��uB�W���&qEE��������Ԥ6�:�J��Y�q'VCueT3���e���1t�R� [��P��D��"�mu7n�I�o-2Phw'�<��fF��� w�5���]o����)����+��Bj�l�TY�x�_扔2w�:��2J�z��Q������b@��]7DY���W, rv
[�i�Q�'��5�X`Xe�����D�ŬQ�$�D��C�H|��j�S]u���3���ղ�p�����Su{Ɗ{tg�<�]�苘
����"�ĳꞷ:h� ����2�?̛r.	P�T���PlP���ڶf��ن��eR��5d��/C:�q�܁J��a	d#�_*��b �VB^�}{x/�*��.0�?�D�<'+�-�|��w����Ua,��D���:ҭ%�,����
����&����B���c,���O���t��Sgh<Z2Q͐uP��"Wk����p6!�X�?d�
A�00ê5���>�ga�I=�U"àpD�qVM,j6+��zȒ��/c��:��=�����x��v��7}k��q�wp��l&�a���P���<��˕Tgv;�JS��=�XϬ��BF��O���h��|���̟(���c�̋S-TԾI'0oΡY)�,N�L��ÀfQK�~q��:%�k[$�9���hTH�D�߅ԿP�콃K_^�h��� ����'h�V�L��Z�]nҫxK�e1� �+k~�/�P���Y��o�3���+�װ���	y!�5Q��(;)Ds��"�׷�����T�n����kO:/�Jݴ��i����6�n�]��M�P�x?;_U�0r��N��.1P޻vR�G�t�* �	R����W�'x��d����9�-�[`i��0�6�%4%�)M���w��SeZg.*~������Iy�E�/�i��ҹ>��r�J�\���J�4��S����<�;T�|� �P�\0�1o���M��I�s����ذ65��\i�)n�*B�}�D� ��;�#��c�-�
|�؍J����A�0ʾ1�AJ����)��%Fy
5n��� �f���h�P +�����:0:��s�1qY���1���d��<`���m�����gN�	����K�H�
q�n�~4�aj���� ��d���!����/T�2=@ӤI��q q/H�Y��]�˟t�6E$�5R����}@[�M��"A�޹�8�� mA,):�*T>
��V����0���"o���l��/N�4<�c#I8
�p�\�<�������#5 LB��y��j܍[�ɮi�{�kIk2:i�º.��JB��S-1�C]�0���cy
���~ǽ��r�q��,��i�q?y��"#}U2Ǐn�EY���O�A�rǴ���$�JBg�j�1�O$�6�נ_Ө��uY��2�G���9G�^�2q	��؎���f�YuD�Xzl��V�4I7�^�M�z����:�;����mQ�A���G:t�8lԉq��}��'����Um�[��r�SWN"�Mq�� �j��,nQ�p�b-���=hd �˛�<��fӞ�冘l'U�p�V� ��U��l0��V�c�����m��{$�7���v��n?�z>4�WA�M�Ro�p*U�̰P���V����i4�bICl��f|5��p��T��M��A���no�z%.����J��61��d�4��k�Kp!q����MO(/|�v�G���[� ,AKe�r��f�X͞*�d	����/)�+3�u����&��n�[K ���2uh~C�C���
�uu~|N:M,��y�b��Z�������rX(wF�˒m)�0�Q�s�%3�U�7�1n�T \@���|k�0��tՂz�D&���u�k͑q�p��)e-u^��m�r�	A[��F�t5�N�&.F4L8ͰQTe'`���e6�g#�H&���q`050E��VʅL�u�etg~�^�(gV2���&/x^�yR}�q� ���i�3[���z2 H��6���b��򾞁/�P1��0�R���x��`$Ͷ��n���	��?F�U�uk���^�Ji毸;�b�f��>q�[6y���]���ZS{5���p��lK����}w�d���MS�Y&D�k��:+���v�� ��n@op!𺽔�UM���������Š��aS���ѕ5�obV5�4ڲ@����E�{��q�Ԅvt��a�����IF?/&�G���=��4o��m����'W2�G&��˾�CHh��/��HF^º���߼�-J
t��6x� 1Ram�b
M�ٓ9Z�fH����
k�@.z�2g௝
�7�_x�
��I�ÂwE"��!����ŵ�c�x_st��*LU��)[����'f���WۂX��&���0*��dBL�!'���<E�È�㡪y�ê���I�K�_��{�UlgL�+G�1���,�]A��4��Z�tՔ��dlgUz��՟�	����h��b̮��P���9G���Z8k�x�������>��l>]g������g츩��/�GAMl��"��<�u@��U��C9w��|�r2�;�-��#U���h,�,��d� �=qo���Z�����k.k0=�����>�W[�fl-�'�x�,w�.oT�9JeP�Ĳ���@b��^��=Y���t�=E������M|�";#�ҟ�j ��:�I�_q�#���=�a��`)o�ADCG@�7Q���U�Q�z��x�O �Ӧ���$(@�SZ��6�ipA�ƙ�x~H"@�G�r��U@y�(`����+�24=>�X�x�` �e�H~��͔A"��Yi�q,(6C�%�� �҆W�pq�$�)�p�V��=Q�`]p��K�������Z�cmP�K듃�c�@:��c �̨��i�+�]F	[�-%$3I~���R�U)��X!WF)Q�E>>�_m��N�W �T��:w#i�Lg��q�ej�7O��*.B�G*�&���+���T:�����"79[��t���#>�iMP�Xc��'Fi���w9��j����3�qf<N�����w ���ɕo�r�J%F�g*woi���?wډ���xuV��ޮ_X/�Φo"�$lQ��~bF�ȌV{���P�ʴ���;*!K����U{�I04*�fG��!\x�����iT(����5S��	R<4��kD�72��8F��Z��B�Te]��&��Յ�!�fԣ��ˠc�����A�`{�s:zt�Mu���(��S�'� ��&*����H��"¼��@�uHUN%�jo�|��G��=H�Ψ���hg�?����܁�f�&�y���J�˔����3�/��=i*c	���Г��>���K���@�q|#������npu���#R�&��۬(6�6aLq���� �-��MPD�5���v�w(��R%�}��u��֎0��Hk��=�rf�]�uĦ��D�u����f�ɴ��Gd��-I���({�K7�*��ܮsy-�GEQ@�쮪\0f5O#f�pC@ɉ�j=Я�ˍ(���:�* -<u(DP*0)s���$c_��-��42����!�]ܱ!:�$������;F��t�?L�����0�9C�����%ϡ��O�><6��>e/�P8�p��C,"���|ŕ?�����Q�� ��.�_(%@FQZ-߲��xe��ĵS>5U�2S���uvk=�A�_|Ѧî��eƺ��t�iKshZ7c؅ nY�7��(W�h󎱻盨P&鎠>)�]ōy��߹f��o��p\(_p�I@�a��u��=��Ba-1g�=�|��V��2:��C�h�Ӯ��ߗ�o�]<��fb�|;�y�w$3/8�C�l�O׏��J��NnO��7��l�@ڵ�K}[��,�DHl�"�	l�2���s��E�۽)J��w8�f�%D*�Gy����7
�@�b'�^7h��eޟ�o� �8u�	�Ma�A�֣��V+5����N�/�)����<l
������6�����
�=�Pb�ViA#�ڔ���I>�4�V���P��-����T-0�n+J�;>3��H�>�#h��N�y�eT_)Ms��A��O���@���t���AP=z�y�BLn�7�{i�K7�e�+e�������(r��~ԫ����r6%���x[�_xĭh;��t�AF=�p�=�]v�~;����~���INZWAþ��4TP�Fq3k�j'vk�7(H��k��9���vb�T��������r-�x��=�	~�2�G�Ҷ��Dm�4��\H����h�*�*%`r4Fvm��< ����n�9�ω��c����p2m?a���~o�ɲ�̄Ikĵ�|!������S�`���K�i#SN��3�}������b<��^6k�qAS�ET+yg� �\l�O؎/�d�_��[�+��I'C�Դ�C��ޗ�x�#��D6I7[��)��զ���h�����������|B���c�4�P�UY�y��K�#��oաy;��8��u�x8JM���&x(O��ʞ,M8�<&�k�V'�b�MM�H�YI��ͅv|ہ

[!�:���+Vr���,���J�輂5㰏4)��d�Tӑ�`�s����vN���\�{�W����s�Lʴ��o���kA�kPF�w�9�xs�<슚���b6�kV"�Ĳ�z	�xu�^KtnI�tI?��!4Qʅ3KQ�������9C1@��(��Rhc��e�z$�w�e�F�<K;��wU}�gC?a��Ɲ��h����f�>\�
�*�ݓq~?�Q�z�	�c�8��4@6X0�x�Gt�+�@�E��G�q�������^O}T����P0qѓ�o1��|�8[����(2���z�e�%򫹖v�q$ @�>���2�0u��Z*����j�����&k3�*~*�G��?�����,�Ɵ��$w~���E�ǩ.��f�ۍ�e�2����80�E~s�+j}F���/��&�yŨ�'���W��Ը��xd���x+sx�A=u�w���w�e_a���V��"M��)�ђk�*��"Ҙ+:^w޳��p��\����Þ��.q9���4���sn6��cj���i�	�(O>on�	�l'y�GѢ�'C�5eޱ�g9��$Eu��S,�i_���Ί�ɁhXN�;fkU1k^�Se�*͘q�ZOA���b8	�U{������R���Qz��1�Q����� ��pp�����Q�
骸��`C�������d��'bU��C5���CP��l64pE���&��߮D�fI'KnP����P��Q���Ro�$�f��H�����OL�@�ü��&<��}:�#~1r���D�Xn3#�#5���T������T۵�AX�u6�ϲ"#��W�o��W۾I]�k�n}�E�(�(�������z[�)ٴ�U`)n��#�ǌ�o��x6	fܕg5�����J��S�1\��?3j!dl�*;��fmz�g��*�ci��T��9�+F	ŭmAq��n�qm���	�D��h�lr 5����D��T��U". fz\��q��K�K�d3�-QPJҢQ�d��W���fF�.[��?>�e��$���w001jY��}���'_�Xcg@F�+"2�C݁��K���������"zm�R���U����UHJ��$E����rϋ�S�lT�88b�<��s��vg�	�@Q�q=�ze:���Ziu�e�OO�  ����B�E�L��)�qz|/YO�/k�^gu#�J�˩���}0�/��	�.&^��Q��(۟���Ƴ��`��=�s�x)�X;�e�����v��e���V��T�ϱd٪QEs���6c���Ȃ�o�������"=����&����f1��7�g1�˶7ϣD#����J����9�������o����_��updۉB�@/M�r�mM[������P��q�m�٠Ѭ�GcG����f-���S��K"��}\����LJ��g1����Z]����N�����b�瓒dm��p����S���� �?|)FJ������E.��_���Z2�lˮ��V��������������mh�������T�`AἩ5���X��!�&;N��h�ğ��L�]���_��{V8,�� �/r��;3;��!�Y�S7�iߛ+���ock�)�9���/+\��9l���s�0�j�������!n�mN���Hʎ�[��Hn�hg�6���ԩHj�!Y�ޖ(i��ܲ�ɼ��RQ}���3�����l'ͺ�t�����|�?�s�9�f  �v��P0SJ��z����Ie��2z��k�ƥٗ�Qt@��/G�������F��J:��C6�ߤ/
�	N�c,Lu���9`Nx��!A�S�Nxm�i��Q���"�^4������4�>�}����,��QsW��\�J6�4����
9t�i�1�%�ƶ�i�/1��$�.��c�L�����;�n�d��ÊP-6��S��?t���P.�C�5x�q^,U��
��L!�/�9�q�u���>_��X��|�L��I␌!_����]�m�-��e�G[������I��]���U��O�6��걁~kB�0�ٶ���쎘��D�
��'ym�\�����n`p��&U.�jċ��e�Q��e����x p.4�S�m�(R��8mQ`��Q��j#	���|+��������m��3�3����z,��	��]{�t6�{��KOw)�в0 [��*o��U��.��z��UȀ=
�kj��/�n����Q5]�
xr�	S��C����ȷ�eb`_��� 6�Ϥ�K�Z��_4}����N!K�*��ߑĥ+����I���%e��]*�\n)�i.��a�ӿ��d��%��bFR���4��Qf��]������9���;�ˍ�zY�9V�����x��.	���������?G�7ʯ�{z�����A�ș$P��1�G_�����Z-��
�M8h�<�!M8H���l�.%\�Ƅwm,��P�7�:ch������c��Q��y�ItQV�3GEn�u�Q���/��	��W����ȎD_�F�7�2�v�L[C	��K���x�)(�T�����I]Ju�-����A�o��W8I>�4�=��qY�t_�d
Ʒ��~]�p���H���i���O�.�%ǋ��k�d��D,�v--91���f&���
IL6��Cq���(䄥���=��ݳ�d��"<ͷ+$�g���Ѵ[�zmw;Md�L���Jز�V��ܽ�	���.���e� �h�|+�W��5��U��b5�%OrM�ICG<r�$I��
��ZEU~�~�`�<2��]0F��#����CcOd���La�^��lGi�BSy���fs���ط�]�՟����!��FQ�Ih��K���5�8�Z�`f�yׇ��Z�9��:�"�nɌ}f�K*��"W������ﭹ5��W��n4.��B�֧Bò�q֠Z�AK�cDi���b0��n��Aul��_�?���Y�l����Q،CC?43y�|n�)�O��$`�'�7��Q�ٱ��<t7Xd.����a!q�����4{�U��4�����CM�u*�aҴsN��c�V
kS"�Dt�[�u�G)� K����ؕ�Z����4hO�a�M"W��KRtk
�*�eZ����Ƒ_<�|):e����q>�W�F��8�>іu1/M���mIx�7K����9�:���L�H��
��<���!�o�`}���g8���`��)8F/�L�9�Oӫ">(��c(Li�C֜�0J��}z�6��)��7����1��3�ѠV���TuQ��m"�pS����u���9��(rU^��eEuƟ��*M���*pb!�E��-�ԝM/��۾G�@�A���w��)�U�N��I��uE�U�Z��)��j��Wp��^��z�.�w��6��-�0C+;q�i�\C��.,�������_T��*�xg�O�5����w���+o�\E�z3�~�h-�\�g������ُb�젃F��r��@�^:�-�Z��l�
���|AI��H�0�tp�S�+{Y7� ��r���u`��9w��HY�^6&��,�{�#��
~}3]n�ӭ��5`%��x�"�:��V�:��\fj&�L�mS�̱z��%]S� ��� �OŰ��3w� q{Y��`�%��hc��i^�Í��T���5��O�F��դ'xpU�l�V���,��o���T�@�B�'���Չ)�������ۥ����ްQ��=��t��;��G�J�Ok��L�����:\�Z�6��Rrl�HU>�>�@�B|Yӛ��ۅ��lQPu�ʆwP�X�0��^ܱ,Ad=a?�	�#2f�뢜x5lmQ7�磽��1��E�"�Z���#tX֙������vߠ��<u�ǵ��?��$֚����<9�v&V�}��tZ�D�>��A��/\��z��Aqθ9�;I�
�����B�g�'T`%_��em�Oʼ+Gc�����~�
�*��α�=��2,2~�c����,M1��3�-�Ŵ�2����5�' ��&����KJ;�D�C�J�t�!MX�p�����CJi��b�ힺ|��spT��ԃ�x�/���f�lN����=R���*LT8�K]\���ߏ�^q�J����n���C���*#��	M�gn�%�0(I6Z�}�s�S�ZU1���+xݳ��]��{O��d�Uh����j��t�&#*���L�����՜��T�BaC�$�v�^��X:���vw"�G;�׉���ժ�W��� �Iٿh����]�`	�*Z<(�lOI�+5��=���G=3���S�y�Q|g�٪�,b��j�Ԡ���ȷ���\d(ێr鴭y7'�t�D1�O��1�R;7ZUW�9[����Bm���I
l�3�˞I��ͬ�F����)�ݣ� ��:hs�����#�p�2W� i��α<�"D��a1ܑLҀ!TaO�J�%�J�J����n#���a"�ұ����]%��n,�Q��/�*P\L��iy�|޽~j�{!�F�z<��p�dv��t��w<9�=!�e)0�a�I�&w~�C�%!��J#��)n��$����&���T<���$��d�(CO�{�W��Ɏ����|�ޮeӎ6��V���{�O5�%��7�3���Vp=k7������1�s�����<Ӽ�A��ϚL�c�z����n�PJ�c�GN���ҹr�}����������26Ҹ��{8��qZ��OV���9b
�l� a�=��LU���Y�Lz�I%�<�t�����|�T��i��S�������$����I���J�� Kvl�E$�B	�d[�u��4�ck&�FV�k�?3� 6�T�ռQ~ѫ�g�-�Io���ۿ�dL{�Wg�h���/8s#Bݪ(�vs�K�gIq��a�uҤ�B�u��l9������ɡ�1�=0j~#K�8��=ql\��Ӓ��.	����f ��{SԒj�Z	m�+�`jnK=|�۰�]�#� �RA>N�	�G�a��"'k��r[�7
0�[m��%~ޔoZ�����x�v2�ӆ��y�L>��'=��� �sw
L��|5��t¢�q�?v���9%�hA���WBF�!B���]Ou<.���%W�Y_jӪ�g7�W�f�q/�H�:'ޗ4�T�+�>���C���o��ڕ�]賩r,�,�����!E�u	�N	,����X��J��qȽ�V�6Y��ӗ�.���� �b�h����C��E*u�sb���@�y����	`�����&z�S�W:�������Ǳ��k��<J�w�[�Yk7���`¤i5U��/�m�;�
��>����<k#���:��N
9�AF�˂2�pM��K<7j���xn����=�DAj�֧,U��ȟ�:k���\��CGxM �K��<��;:���-d?4Ս�`�>V&��b\[�p׮<Oȉ��ɉ/mݎ^p
dR9��y���:�aq�-�l6�����J���x顇���]J�V8R�ȳIꝜ"-z���TZ} M���lz4M��Cl��Ű =��O$�Uw���4�Cl��(��f!$/��̃<42��W3}SA��Q��nk8Edm��y��/:�	��;L"Ե�$	[`R��ӹ=���M�/},�&L�
��A��X
�_��h�&��fJ/�t).��Z�+��QP`�s��7�6V���sM����-�o��/�~~a�ف::�M7�H�wy��h<0�F÷qS�a���� �{���_Y��9Ƚ�x��L~��h��̾E���ݥu�t�1;�Ź/x�{Z,���~|�&Y?�ZA���ymp�%h�h��J"�����'��t����͋>���BmZb_���ޣ�X���%��ȋ"��44�1s8���^��7�u7���T7f�膁r7�v[n����Q79�w���2[�@�T��jp�NN]SD6M���H#l��4�CH�KkC���(7��n��
��:N��х�|i�;mu�m����S���'&��������I>�u����
զ��'c"Cw4�(�Ҫ�3�o�;�H�l����
Ҵ+Jiba���19~� ���N�\�r*'�T�	���!��͌p�𤌇P�=3�c]�	���W��,oz��5O@BS��\,j�߻����¥ޥ˰H^p�6�v<	�E ϖPD�U��ck��ֹ@P4�'B��m�i�:<�dND5i??��ZOM`,l<͍!��D cۙ�m��|���y,׬^-�i��U�d����2�n�d���}mU楳!��Z�~�YW�"-:�誘v� ��CŔW2��Fϒt��Sp4�j~?p�����K<s���6��+I�H��(rA����{�M���y��ŕ��¬2�"�͕�w�6�×Vl��V���-�V�z8bp+;b���a�̭���!��>��^���L�,��h�L�;%�����VS$�(��)Kw�-��A|���5�����ΡӲ*�c� h�@��,1va���;x/��2��H��?��L���-��!���c��xj�+G(�n�5�:���;��D����Q�`0%��ƪ���sH�+ư�gi <�T�۪ I#�/����@��4����-l�[�
ڒq��-nl��pZa$O�#CE��.Ρs�d�I��$/Ai��P�Q9�-��?���(7���݌�D=J�����5�Y�j�x�5MZR��N��>�3��3-/@�BIs��!
=CT�BB������x�e?dz���w����=M����.������)I	���G�&�^��B��}� �y�X'��.d�����5�f~1УN�`�b?��X�_���B��Ag��'�=����Zg��	L
�c����մ���i�7$g���ɰӕ�;!C5��kwytq�(=�/D�@<4c� :��;�T�$���Oa(׌��w�p���!�sl�d|�w̍g����ְ����ڰO����웬`BN�r��r$�1���xb����6I�B��|V`�'�����R�F%B:����+ƞs�
B�r���L�	ٜ���I���x?����J�HB���tަ�Κ���L������w���ͦߌG�眣*��^�+�\]�+E?!Z�Mi��{�k)�⏋u�U��]���q�C^�#Q�j1���)���a�O2�8�I�|���$�W�@�����T�#{�)���X��G>N~gҭ/U�I_�y�[�:��B�lM&��@��K�j�0&1E���N��n����/��Y�SfB�~L��w)_%�������'4 �;�7?��t�5��<C}j�a�'__Tzu7w��M�x#�8�F74�x���o[��(�X[��9�A�!H�^�ռ �U5y��j��]���08A���5F��D��4�&="/�(�J��zD��u�Yr��F�&C4��� ]�ł�	;��wk�'�xKZa��Dy��2"�7?+j�}[-X���XD|��{c-&�H"Z������p���@RFki,+т�Oﴆ�g�R#�^Zn�f*ww�ɇ����C���%s˱�oKp�Tv�	�2M���e�\4�+G=��	Bsc=����G�Lߜi�؞h���OW@OY�
��z=fre�f�Չ�=�
 u�����M$�z`���u��5�O�$��y�q��K ��ᙳ�,���R|M:@L�|R�|�p���(DcAjVvǔ�Q{$��ß��v��ss��c�������Z��6�J �n�DN������Yqu��� NڒS�z1f H�'|�a�� K�K��ʣ�����/�9�%,�z��i���2�0AJ�^�>M_�l��O-���7s7�tkg���c�l��C�sx �i!�8�xg[��N��D��j��nR�̜�D�K�Z�p���A��Itu��@���yBq��'/���A�K����R1��֛���!*IFhI��&����f<�����~E!
�.J7��'�xP{&��ra1g)\�K*zV�=U���Hg�C�B�D�;|��N�vL\U;���:M|l�1�T{8k2����x��&��?�����:,}�? 3�zU�y�m� jK:?s�S�q�����v׃�4ÿ�](9��E'ֱ0XkBT�J�fy>(e��VW�f���O#��j�6$�2Ѳ��v���I����C�t���?*���h��X�n�Z"�|�@f��X�gM��ךW��%���$n\�W P�E�����5,��R�9����o�P-z��54�U���3�AJ�x���.-�5�/�NTJ��Q��y�ξ5�Ib����*S�5LK=z21�����B���p�n�����7��jFF�u/gB����^��^��o��^'���Cw��0�ʟ3U]��B�>Y/;���*�]��+��'�wݢ����~��T�o�O���	�DE�l�ՕjP�h���L+�տ$���Ԥ6���bL`��7��'�v��Yc��â�nu��*�����T��bAݵ��ݽwQV��>9n[��џ�'_��4���t�i��S��숃��[%uN(o��ew�ڭ���|��jEr�
c<��쮢���&C1�����9�6̥�~�}z�Y/�Ћ|稟	Jl���k��駷m�)�̅��t�M��$��ބy!��u7�^3�>�Gԃ�����^�1����`#8�+��q���o�U��@ ޒ�TB��.�C�e��]���{�՟��@]��5A?Y�zhͯ77��uN��3�p�< Z���-YP ��ْ ��^h+�\J�L�a��)����75
ǲɷG�5��Ȱ���>}6�0L�"=�Cq\^a�G�{�OX��D��$C�=�/y�C3vӘ����8��9,&���@��E�#�'���d{z�yP�\W���M����Z��젽Q���D�S�z�:*��i��,Z�S�k捿t2�H���G��uﻁ!Eh3Q7�<g	:�{d;\�o]$�]���uy0K�[B�Lgv%~����N	ߘ�>��ܿv�=.z���޳�h�}듧��?=0���,�f��k��r3�$=� �S<�)������5wbO���0��d��F��$!�ӳ��QQ.X^�y�y��%-��~�\����sB뢰I�x�ܛ�3��vNE��-Z]�{x�6���@���ƪ����.T���KI�L��,�D�3�kT}c���N;�h�������XĒ�6�>��(���K�{��K���է��Bv7x�q-�%���O1#�Mɿ���Ky�(���r��a6�NF��YZh�r���z鋸�
f$2��û��f���.|�ak�̞#IiӸ<��ү�g���x:y�����x��T�P��.-�Q����Lî20��7�y�>/�N�ޅ����ȝ�!��>5cA�ܘ��ݪ�y�=b�ۃ����dO�e�[�m_AY :'������9��_%��K�G��^w�* �g�xuG_��b�m�=ps����90�~z���>�|@�a\��7uթ�*�����FtAϓ��~<y�E��X72	�uF%r�����D�i��L��~��'[�����b;�q�ťIZ�9��݀;.Q�_�^VP�ڬ_���7�Ol�a3��gmvjz�#D7FEc���J�ktr�_~Pz�J1�H���zdz�\~?j\��}�+|���L�"���"�9ֺ��*�p�����%*=�͐-WҮl'i@B�G�����ǼJ.�U��O�8�ɘl��h[#ȵ:o� �?�1l��1ۨ��C{��1]��1�[�[�Pi�$ĩغ ���r��r����C;�y������"q�_���3��J[�RG���Hy�,��VCV��0К�;8+	Uc7ϡGhk�6���%'I�R#��Y���Ebj-׽�w�O�Bot�3�?U����7]t�n��_��~d�G�ɹ�!�R�߻�D�ܠ�ɲ�S"	d9r��b� ��R��b��̚�c[U܂���&�N�2_�ؐ�)L��s��k���\>��k)�US�5�5k�  2[�<|p�Dh��H��vQ��ś���י�A=��?oy�� ��zW����
X�Ǔ��D��޷A����C�ߍ���� �VT#���?����^�)&-���a�9�g&K�D����5���[�T�d�ȏ�0�������\E�帀�6���+갏J��U7��]�%��j�������6��{�N�m�����[!�1��aj��&�1ҍ�~�����M�Z��=H�����	�\gY�O*��Ѧ4�}��	'Uw�	�~'��9?����S��>]F�2%o)֡@�^E\��F7o��3Ia��${��&�̟�rQu�@Yx��:�����~ �[<sJ�7��2��j[9�Y��a\�ֆ�th}��EܰX,j!���ҋ��͈A�-���s�40U>wl�C�m��
&�t=ё�	��a��>��ӹ~B�>L8pC��7���Jl(׆ΗKX����tkl�[�K
!����]��ח�Hӝ�4D�b��m�������vHj�� �LB]�O��6�n��;ԡ�	������	�}���
�g�U���?�%�^C�r*w���A�2���)R�����Ch��h��!�0m!W����B!�܇Y��q����s�33���Ӎ��A�´]7;�̼�l>�"�{�i�����R6U|��m�T^�b����S+2�3����T���0�C���v��ߨS3#G�})��v���s��#���Y��L�\7J]|'&tLx�8�����zK�(�7�h��\��Z�L汢 ��>�>���V&�I�SYR��{L����T���(@�����^r�8�w����ұ<��qv$�;wüm�._�$��Mi��'r~��K�����,#yU�������3���{i�@�C�~���M%�l�R8�|��aJ4(��T�[��6���ϖ��/��W��S����ΘC�ٚ5��e�vn�4�Q[b(�=f���a�	��c�:_Ɵ�)�TIm/�/��-z]����+�hg�t���4[P㊲�������U�Wo���Uk*�j*vQ�h}�?��O[��uߍ��
�:�+U�����,�ti��}Qd4&`<�;�Ny�H�X^(��'UZ�aFK�^�5\ cW��E����5�����e�W���}�T���{�V�`-�����:e�ɥ@
��ƽ�\B��OS��~�u�ˊ��f�����\�)z7����O�"�C�ˋֲ�"U�����|���$������E�6�H�2�ۙ͂�ΜO4��8\����v82���Fz���M����8�Upi�r]�C�O䞒����b��T< u;'��+�_��8c�VI�t<~�d�S�ܰ;41�t��v�<o�.Քg�M\���r<4lB�}:�pn����v�����&����t+��R#�q��9�V�5!�Iwq�w}h��]�c*�I�2~�K��yU�`5��մA�l"~4��t���*�|���z�P�A�oX3`�Â�Ú������g�]=���3���ː#�/�4N�M�g$4釅A{#�:��=�m�Q�qX39?2~1H�l<z=���:㬴Wi۰.5/O��-\,��b.i������l��u+gJ 3�!�>)�֘$ d�aS;�ʛ��ί636�=������ky.��T)F)�(@�,=޿z�R2�we���ٲB�6���R��D������t��r1~A�EV�c�`����Q%�kه���l�(�-�h���/)4����H0�3�P%�4�C��c�-�/B��� ��kf��~�,Q����A��P87A�>�r?b��d���}n<���6^�XY�gI�D#k�)EV�Dɯ�RZ x�w?��5Ԯ����R�A������5�G��el�+��ke:��h_k��w-H��1�/�
H��܃��fjXD���w-�hD��ٰ���&f������IːP�@��@��hk���˜I�W���
���B.����F`�IO�|���\��
)��^�x�)� ���8[�@��,�����?!,A�3ֶMn�H��C�]�k�q�,-.�]Y_y%�a�K�<,Uek��9r⅘�L�J]��D8"�bJ��[�?�F��x+5q�`Q.�^����< ��<��Uc��72Ywl!�:>�ܠ"�i�4̈́Pʚ�W[<<�_���~��`�,�+7��7�ޘу�t*�,S
�tB%�@�lyxɩ�d�
�mY4��s�ȼ�ӎ��'{�Szؠ��B��Î�*�8/���V�!�/Ñ��e�-���m�P����T��j�KYm�@�� f(�˘�^� �c��� �d2�.}����Q�\�z��;�,�|��;@k�|_uN���M�Y�����m��R82����%9l,�hq���Y�tYF<KO1M�q��z��'mE���ܣ�Z$�n�SɁ�q��ݺ>�	��J���3֞ �v��GrsM���Bv���������Gv��$�˞���_�Z��I��lq��[�ߔ�1�^���wJ�g��)�ߡ��К#"J�x�dh����b(16�q���3���[�2D��I �y�+(�p��H)_Fv�H�&�ZR1�F1/rk�����&�+��g��|N�s!d�ʴ��<�r1Aw�4��^~v,����{�1n�2��S֥K.Q�aS+��B:}�s�X�x�7��٣�#�ޢ�"�K�n�a�� !U93S���SWS.���?o^.��Xv��į�'8��*�f
~�KnFB}�.�h YJ�P#�X]\X�v�A���4s[ﴹ��h=C�C��?O1����n��;�V&�,��bth�~I��֧���f����(���(ɳMV�_�l���x�S�|���!���7��c�7m�<�6��8{�VpSL�Qx��;j���(�H�v7m��H4��#^��8���OI��,�1��ۢ[����2���n�}���A�_P���b�9����s��<~�1d"�*.hs��$)@뀷�h�@�QV�k��'��j�,*�1�[�G.��M'���)�̧�:Q��g�_nTNe������#w���Y�g��
�4�S
����X&_4IU��JƇ�ǔU3<VN����ܼ�e�.�|��|��DN�$�6\EC�]��Pg�E���� 3`8�z0�J�&�r.�}���ͫ��G	����A 3�����4��R`��o3G�<G%8iZF4Q|��围q��q��u�U�Ń�c�4tNM�K�`P���%�	r�;xr�yآ�|#���d4��[��>|[�B��i��8�!�v0�8WѹF,/�j�:�$�)P:|��^���E��[!�d4��CJRK| �g>�@���ܜ�d>�I�yg.L�<*ǁb�m�������P��9�鷾�ݣ����KD�����>2{��?���]�KC����ff~i{''^3�
J�}���� �K�%�ҙ���`z�>j�����#�`~wv��[�"������4�b�),�1��M�D/�_�4d�>�ɤ�\�Q��JA
�	�H��E0�麞�u�	
8)�� 	�K[��R�L�RM'�j��RS�Ϡ`�8�-��1�y{�a2(]����F=P��፪�e�jY/.�3���o��z!��iV��X~���@$KK2�`%����`�v��)��S���O�o&��ם����'g�~'|����p1�0 ;�k̟xok\�&F��m�\VL؈��E=o�n����@��Rc[ƕv=1�=��Z
ٹz����O98�h���i��jF��P���D����pVn��(�`�!.�B��Y��SO��w��X�l��������)��|yxʎ�|��8BHI�"&���7���@7�(k�~�㫢u�*���'��<�ld�a�����j/�r�]�3!�l�)zl��X/�g�[?'�OT��9`�n`�=�J�p$��Z��K�n�t��C�����|,��#�.�/n=*��
P�;�2�����_��f0�Q�tq	n(����R��H#����F.|�U�	�zb"��Qi�=[^Ⱥ�ψU�@�Y�O�(�%U��;��C�S XFe3��a=f-���Ԅ�"�O�ʊʹ��������UÔ>�T,�(|�9�_nO���o��`HLJ�͎i�_0향���6�3���ť��3l
g�L�����3�ES����8�� �3 �p1�T���}G�
��S���AB����`��
YU�HjZLI�-V���z�c)+L%��gb����K1�n*�IlH����#A`[���uF�ZS���B�z6���[�n�β�i�l
�G
��n=&�o����ұȧ��o�S���ȨqS�o�z��n[�:f!��G���P ��g�}��~�ЁR��I���V�jb��c���z�W�cS����!�L��h5��d�g0��j�r�]µ���AXY�;c�����s�uX_��;l�$��2��=u�6�g�����%xc��	�W�0�_.c9�i� X�6K4�i_H4&"�Z�
09��\7�]6V�=Kq2[b5���,����;d�i)��N�
���&wԯQ\���5&�@Qӫ!鲣�Y����3�d��B���`��ͨZ`D�����\�>�־�.�ߔ{Ȑgg�z&����5��檻�;��b�F���c���s�w"Nչ��jP�-�D��w�c]�����wg���_kq�
&rD6ץ���u7��.D��jL&N�G@���?+ߔԁօ�nݾsؤ��z�h5��冩�#,����GBS�3$qVx<�SH������oԺ�[�5���a�\���� .��� ��͠�9�C.֏�q�"yD����[:Yccꉑ�w�Z%�r�훙�1��#n{�G����&���m�OB�Sc�V{c�E~�!�D@�6��u<&�F�����y�G��TX�SL�H&g��,3F���;��7�hG��EM��FGr�_Iӓ�@+I�~�P&���c-ʘ
��=���M�ً*ٛ�E�:_���3�6ĉ�p�[n/�<?��b�F���Ѡ{Zx%P��ƣr)�,EK�.������a�x9��^�O}���v{%ӗt���*2�;�cCL5t�e=��w�
��QN��e�>p<Օ�Ĕ8�q��B� 7��I����>���ī���xX�����7�\��D�8-Y}o�Y��ҧ��QD�o��f)�cd�y��� ���Sǻ�ʍ�b�]/_a!L�?slU�b,�,�d��i�7�c��j�a����t�Q(�<��7K�A�#S`?�o���%=������:����?O�Tjg�{�m�M#�V����l#%��!"ũ�5���݉�R�Al1!J[8�ztD�S8�(i�߰����$s�hLiŽ������&��(�]�cz�յu�j�5��>�dj�(u��¦e��6�h��9=�;7��m{�O��D.͏k���S�Z�������>��EKO�14�QZ�o�<AP2���}8'"9��@�q75�}�f�j�W��3�4�{j���>��c����7D�p�.���5R���oN��� c�}F?$����\UU���8�݄�(�cf����\��Ԇ+pb���t�K����BK��{�qp�m��ǱK�!(�z�_�uIe�*�RDz5��m6E����-x������mx���8.�uߩ:Gs2v$�!�������F�H,�\��p��g}
&=�fS\��fc�[��rxå���v�-�
(��a���w�_�������۩,*��Ā Z�P�<��Tc��w�-����_�b��^L�X��9t<-~REn�۷mB���0[�����\��c�O._	|�9�v|���~z;4@�-��u�X����Y�n��$qك�	�>�M�ca��?���?7����4&U��]x\L/g=Q��{r��b�yڼX6N���P���g�����.�F�\>���>���d���#��$#Rv��2	�"!2�����ɞ���8�I<BZ�/����&|�]�s,���1p�K�7��I�'I+\���d�z�
cB������
�hk�cq-���;2�v�χ���c�+���.
�ӗtE� �~�Y��~^�GH��L�vJ���`4�$r���&G7���,�[F��7*�~�����h\Ģ���]WU�NO��X�[R��g�+��qϻP;0�޲�57�|����)?�~�oJU!�ͪ�r ;��N
e�"�MU�.�a��VvH��9��sSc��⋾�߳���N��	�0����HO���ST��3�)����|�_�ˏ��� P�wk.Fcʚ��:7�w�H�p-�B���-K�����`����侵{��
o�+�=b/���f�,T�R[����#s�dI� D��h:�πu:p%�E+��4�S��z�����O�����#�$m����~�]�Ce�P�Dوi%={�;�|���GLis���'ǛC�?5�C��JQ�����@�������X@LѮx?%���Ϗ�ϫ���H`�q�隲Ԇ4��]��������'8�B!��PaH��^k���A\(��q����:1��]��J�ZB	�"`<���5��l^bk1�@�]A�`��0��69���j6�t�s߼[�����!HK :1��Jռ��4B��AQqZ�s���֑��kW�v��d�2�x��Y1�����:�YK�yU���H ��]*`�zd�����l�W��AzŌ'}/b��P� G�t�}3E�c� ��cщ���Fp.ʆ]#`�#���O�h���ש����;WSp'M zV����B�-��ؤu�%�:��*.}���{��=a��@sx�Ӗ�x��0UL[���'l���tI�oH�s�M��?Wĵ�~'���drtDp�{��Fu�1g2���K	�7�M�:�^A0�Ԗ���{����ShK6<�	�-���Ԟ^�o5Rֱ��j��!���HX�`�5�&�b��|aK�'p'<��>_M�/��ӌ���Dn�Gkg���s`��5���;ڽJ���Χf��'�P�7��_��\D�-8E2��w��������
{r�f��7�4�!^'<W+���	�o�|�������}mv2��=�⋿�r���L�(�5���H�o�����%$�݅����� }��^�)����)�����O(�[�%�a�#��>P�����
$�u�C��q�h �s��_�y������?��=�~�?D�jGH�.��\�w�5�*�� vv&����YX0H�i l.��2��9��c�
&q�Z�P����p��Zp��� S��G���Q�+����TaF*�hu�(���FB�M���b$�2�FKE~�x�0��Bw�����u���5���ݒ!{h�Rȫ�dT�޺�7VXkt��ӊ�
H�p���Ȟ~5A�C�$`��K�������!�$�(�s���~�!���q�?k�͸�"�EޏN�7�i�*��� <�������]�؛�o.���aʂt˔�G3��T�	��6
��(�"-b��2L�*6�f2:i�*2���`��)�,���ú�|�g��}���$aA��0R�X���KK�ڒɞ���Qh��{�̎)n-�,����D6��#�����3�*�c/��=�i�ݏY� d�_�>�^� N�;{��)4+�|1�qC�o 3�v3/:��j\�Q� ��@�V�Z$�gi'ɸA��.�p��Gd��a����_6�^Z6��`�Z��$�ןY�>���|�ZEa^ڳ^�V�_���D�I���"�]_<[[r��W�y����My�	9h-���:՗8�9��}m4] 4�	�����
��J��Fcu�3*d'��ނDQ��?-`��i�g��s�;V���)L<�s��uU�t&�XW[H�B��@AB���-M�#�v�uCq6�L���e�����$j��146k�8�ݮ��:<m2p����d�(��.R����ݞ=����m]��(�D^5�O?mۂMH��D<��&o�p������G�)�����M�J�/����d��.�=5��+��\�#Gg���]��Ɉ��>�bk��ۺ_k��F����W!�O�{5��'���u;�o�V]�z<ٟ�}��zΈ&���W���t=ԭ�BTЦ�Y,��av��P�k�u=}��+�[�cQaNo�c���s�/
v# ��ǥ��D7��J��~ηSH�:�����8��pA6��,L5���l�RW�iĲ���=�Q�îW;��#��Չ�d��^}���f�)?{�ʝ�X��0������t��)	Qڞ�UNy�x����6�!|8〘���at?9hP�{_o�/�;󪆉 !zT���L��~$	��������e��c�gs�L��X��&�"��3ތ8�p�2�W�&<�q�ƀr��[�Ɣ���?��U��Ԑ�.2�U�?�MkE2���$�]�qZg�C���r[U���ɯ�7�d�E�Б' ��BN!<�!�K��BN������v��F7*���:	��>���%!_:#f��b�i��z�D���*X�vPs7�"ւ+������ަ��y\�g�f���6���k!�"\̥;��f���_k���[B�hx-���3��r y<�C�Å{�QV]��!)/%x��v�jOL����Ï����L>���T��<�A���N/��T���\
���r5~����h`���Ձ��%�⇉mu:?*2�i5���6�>�= ��5)���D
�?zc��FNF���#hQ,�f��-��[�mR�#�|(��<�R�UGZB�u5f�pldK��<v���������v1:���0��6�	W��?��`����<�oɓ\��J/렧�e�PDα_�wW,	��v�7�W�D�|9��\�U�r�h�ř^% &pH_�+U��+=b���T���6��)Ů5���C{@�^w	�bM��A��#k7B7?��E����P5,�x���A�ی\���(c���FEe���xZL��K������2�<�TlB�U�
H��q�)�ڋ�>7Q��M`j��e��޹��m�G�"�"`g�r�w�|%���p�	�6�j�9,{��

z�7��3��\]�c>*��i���'��z<6^U{��� �jz5��cf�R�^��h�ar��o�}8�%5�D�+,kJ�c\>��%�މ=M�e��S}*?��C�u��X�?+�N� �j��r�J���C���W������=��ʥ;
��P��5v������\A��4�~v�D��Z�)rD �ZG��?F���`�W��a�BB0�8l)M��0�;��4�p�%��� CCe�&�F���ıa!�ԃ�Πj��e�:U�l�t8�3t��h��xs	�͝�b�"�o�(�@�U�_�sb��8����B �:��+�<�ވ�|�Q��H�z��X$���D1�!��㷳��h
�@R�v<O�u��I+`��!u����m���ɡ��2�5�t�"��9$�wR807,fc���CIpOUpi�����ꂳ�ծF�.g]�y ���W��K���������QS�I�X�J��R~-ሜ���ԙ�\x�g�L��G��8���i:"R8%�A��t��'��O7k�<}G� �:@�2�<����K`�2��>�k"��vp7��#y���ݹt=M8�
S���MDYš�*n3��6m�lE�F���v�Cd�/.C6q�d<;sZv���V:��o��V�u�� ���/8�ъL�����4�<nHzN1�GZ�=�@^��M�$��l�����*�R���]yQ�B���Ӑ��;�&���ޟ^��ا
ҒE{��8!��+�]L��Ŗ}
��@uì�5>y�횀a�����W��6�����g�Dx��)L�����Z4r����X��= ���|�ld�N��N�ʎ&��c��mB1F���q��;�z�,^�%�xk�}�n�e(y��4o��ЇB���$�i�s@�k豴�R,3a��/�4V��}��-#U��m���k� 5D�L��9��.?�]M;��cN�LK�a�%)��ݏ>֬4Y��	!���f���WEݪ����CC�,�J.[ �:1�Y*���	B�Z2&��87�KbQW'x�D)��.��2��f�_��E^!�"V6Sk�*>��>���� ��\�_F�ha�<�"q�M@�����ʀS�����?3^.h���l3���p�1
��E�\�������xr^+�@!�KJ[�*��bj�+q�������[��}�c..p	O��91���JbݹHG=�g	�M��y�v~<Y����P���#@�ծx��.SޡO�7��<�A���9Bw���j��z�[8;@\��
f~�@_�zs�:L~�D�91KKZJ]��D��؛YPb7�ߣ��&�oL�aOz:&�4��rW�g�ƻ:��ЩsJ�Q�4����ԙk\��h�M�1C0q%���£z{����Lfgؕ%/S!Ȯ>��0M�7�n�7��"�1pP�*/��֊���ֵ�G@<;PUB��Q��!\������F�5�%k>Ŭ0���e�`4ɶM߅��P�E���V��Z�zx{�dH����%�>=�Lg�.����,�k0�w��J7�mk�Tx�7�|l&HJ�OUg�i�D�������#>E����(:�6�N0f��e �1��g�S�;9M� b���ӆ�2�LIo�E|A�ԝ�׺��/���YPZ���7����
| �)&�x�+��eR�kw]��]��e�S��d�'�3���@C�����Y�/k=dd�՘S�#��u�Y.�.
�ZE��d��V�����K%*�W�Di��3A�ͅ�x�Q�lm�8�}"���=�r[`Y"���M��b���_�/��im��kd' �M��yG�?�~�&���j���Ba�h*��%wޤ����� 'F�Ker��R�Hr>������5�>I��ދQ!��qM#���h�*����;10Ra�<5,0}�ŰO�(L����3�C�g8"�+0<��<����R�ɷx(�"Qr��6_�uKN ��Nm�'�O�K]������-�n<��Uo����tфsw�L�0=B�Q�^�U� �. �/�V���1���CxмCm���'l�_%S�jj�.́��xY+4�=�
5	,d���r�%����96��LT��Y�k��I; %���z|���-W)5�\�KU�$=�~TE�O�EN����1�ց����F�C�h���7���=�'�B�����(��m,���T�4���ʇ��x��Ӥw,��2�*\�^���-n��<㑆�X�|(��ު��@�5��}R�\�S��ہj]��gvqgG,,%I]���YE��G{ap����������Ü'��(�,ܤ)�s�ћ����>~�D�.OX�z������bP�s��EBÎ�؉����%��v|��#�q���0�|�rN	C�~7�h)t*6g��Q톪ȵگ�+X@r��=ѤcHΦs��NfM�a��I�#*d�Ӊ�&�	}+����4��-U��Qi�	8#v7�:�'�zL-���!�w��<�����ت܂��؈+�~���|��Q���E���%�)
������WI�D�\8p3]���v�@Zg�G�m��GH��b0f�z�?k�N�[�QVMH�j�_�E�MA��|���Ā��%zpXm�4�C�O�r|��Y��L�	��lN1�qA��Bm/�����Wd���\)�$}����j��VZi�y��,C*��q�~Rg�H���M��)��� ��c���+0>pH�Mz�U��oe^��@�s�r\�2�����L�Ιv�<��͡�"&���5a��7Zi�"U�(Y'ise��'k�_q��� �Y��:�̲���,gKD��}g'$k���1RV_�մ����9�htGƩ�+�E��ހ&B�X�fD`iE��(�⽴�(���n�/�f)�;��������H�{��\�|���r��N�Z�Y�<Ӣ�15q���i���fKWN�`8��֚Y�'�I2���@$�9�Ĳ�CN�}�����?q�lH�#��x�$"2��bm8�5��ǵuj�ُ��
>���Ŵ��ֶ��2�e�P{��~���E?ݪ)��Xq} �]B(߆؈��C���jjQD�rJ�!�-�0<�'4+�� ����0��P#��鸆�7"m�~�T2J&3������8� �NHnP�D�cn$\���]�##�����ɻk o5�h�{8��p�E�ǐHN�l�^�s�9�0�wJ��=euO[�ָ������r�p��S�׿.qH:�*�O3��R	�O{�vb<����@;.�ʢU��R�0'Cx���q���o ���cS�Z�О��_(�z뼎��l����7!��g��Xn+���ax ��Y����ѡ�ʅ�B�+N�U��$��sQ��l�}=�H���F�0f߱��LU��<���:�DY�!5�̒���0E�\���B��8�]m	�o��{���G*�,v���Y�L�E.�?u��rHHF*}G����j�m��3��aV:�-
l��'�;�N�^I+�͕n����<�U������������ś��t�_ͨj��b�b�Z��"��>N]P��^��9�-�{���QZ�sP� ��:����x�Ǔ�y
�r��o(�CR=Z
X-�n�3?�F���0�/"
�����C�cߡ=�FA�J�~hz83gӠ�>M�dCCB"�{}s��"	��:~�au=�Wo���p�d�El�:S����Ybf��[)*/�"��g�5��ZB%�TL��X!r�#��a�_��3�D���:�y`���85��<ρUN\$�ŇJ�{��4�W��k�GA~J�O��q��8+E
C�[2���9�U7�Ǿ^]���7fT+�`�{���J����J1�y��	T�`�[Xs�"Hㆩ���Y\!�w���� #
�ⴤ5Z�Ak��jL���~��\�]2��p���{?\��@�����w_���i��mEח�+kj�f����X6�r`����|h8bAc�M�*�+��S�2�Ъ"~����9�$��V*���D!���C5ˋ�z����X��*\���sX*Y���8�7�/����gg��-�Jq24��VUS*��G��֐,#���t��h��cF_����sc��
�B�!~�0e�H9�07���b�*_˟�B�!���Bo���oך�h�|2��D���&��8�	�</�~���A���A���<�o�a��!b�'���@�;M�=��4"�n`>J�d1�%q^灟��)R�8?wB��\b6`�F�h�������.m��{�_(���/������>+)a:�5#���H�!.�E���V��q�d70.;.��K�w(Y9�福���}o
Fy�X"X&���gԸ)�4>