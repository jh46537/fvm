��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨס�>�6a�
�Ys����'Gc�$��@	[��%�1<����J�I�$��O1������9O�(��/mui�L�'���)J	�p;����ݬ�ת��Ud�����I�G�b��[
X�yc��2g
k�4?�Vs��A�D���`�� �*z��}�໮c��ԉ�@/��\�M[#i�2�Ǔ:�{uqЙS���w�vnFOT�<�O��a�\�	u ڗ��7:�x����1jPቂ^�*l��c#�p�m�ߴt0@Dlr��i�i���[�J��t���2�P�. �l�&�扂�ړu�3���B���g"�K�c�E�%���E�%��0�q���_Ď
�#����H5���1B�@�1�Ɛ�f�����
;�q������Z�ˏK �tC,�A7������,�̩���rL�@�+,��9"kO(��A�!�;��UhX���"��ԅ��h�l�.�פ��(�EV=���N2������ԇg�羋��
�k΅��m�|�>��g��y��o_�i֫Y�V�|a�$�\�S+t}����1��ó�C,7A�j��Vj�,�8�$Äϧ�^W1�V۟\h�D7S��LsM0��_<�?kp��S���ѻ 	=Nk;��p��CP����GH���xiV�z`DĖ�ӹw�K$�?�O�:>�!��6@I��B\v�'��٭��]��oQ?a�ZF�N<[0po<�õ��Ju�G�'�G�H��vZ�#�e�
���M("��r�jwȂL�ȡ���e[B�����&3N���(3ߏ������fn�� u��u�ա�4�'|xY�QOQ��Ƕ�}.�F�5�H�����RO@+���~�#�%�F�ef�z2S����ʉov~��uN�ι��]Ǣ�V�Y趦����/>��P�\J�9B�>��k�e�ǉ�)2w�>0sq�1��E������0l�i��{�eG�w
�i9>��i3�sx���(��x��CS)���W��E]�
���q�����]��:Et�ѷzqF$LOLy�wE= ]�DՒ)���
d�w���"��9V*CMJ�ge�f	A�����w�eǱ��K��E�ndg|B3*>���;O$Z��3YX��l͇u6��,��?��n u-����ߎ�y��΁��TZO�(�Sh���
���
Y�\W�Z��������T����@�����|f�~s9��g���}=#e4�ُܻ�/���0>1|ED�$�sj9�%�ԁ�<����#�ׁ�N����HMsK�<n$�0Z3���L�fPY����"[��sQ��$��N6B��XXS`�a"Y��r�.� +�L�M߬����cX�v��{�;�A���Sܦ�� 	?�e�5�N{p'B�6
y�m>Jt��r��r����gP��C4s���6oS��%6f�*q�5�o�w)�t�]V�7u6%
�0�)1���l��3�$+r#���eA�VG�V��nW7A+�K���>�����@��$����7�<���[�v�H��u�#�V�1��������b&k�:xi�c|M���ẞ9�R����+"#Wb�P1Js};��WH�m�	 ���;�����<�r�[�]Cy�ۛPJt��v!'{�(�J����l���ʟm��0�a6�����}�r3Ǯ��3�(cT�|!�0ğ�}V�~v��cL��j���.�8���~_� ��C&�DFЧ@"i��}��!�O{z�q��^c�W�n	J������S�E1���鱝dc�ӓ���h�*]��^�j�>E��kh���W���]��_;��ey<]\�Y\J�a�M3�C1��X�����;�����#�EI�ֲ`��rc�kJϑу*X��V��u=㐤�m�j��($Ց�o���q�Nrc�OE���?��"�t�/T�E�im0�>imu�]���:�}��K�p�Q��N���Ra�xՃ��-C���~z�t������L�<�}m�X�/�4�_{�:�@��
��n�P��x������-,G�<��WPJ�k��ZC����+=[;;�r�v��i�)4�a�6:��:��*T�K�Cf��re�=�V���;ӂn��Yʍ�iA���m)����*��^���Vv���]����������9~ G�1�"dnۼ; �|n��z��9��#��
�F���Ĉx�^���bymR��?QH ����'{{*�$
�RN�=��D�O������.�ԽW]P�!g#�+��W.qEE*�$�\#1W���/���v,��$­wJY������������w���@�2�5@��'E��k��8�sx"�D���u�Cb�K�q�Z?ظ�FmQ� a�r{%�(���{7��b�Z��F�̀��6�m$�~��.1�(�]M"'�n�?$Z2
�0�$����P�\���[m����$-��b&,qt��y��b�W77�V�o<ڈ��,ʫ��n#��Diƽ�[~�23~r�g����ҁ}l&d�P����x%b��*��Ip*�G��:�+O��jj�1�3i���5�O7u�ΈH0&Bϳ�R2.	����,L\�����k��09F2�gP<����O	��RR2�/��Z��7S�T����Fa�&֩�0�hH�W�V��sV�J "�?�����sV��B-fs�.d�x�!fo��CS��#���;�|f�G��
�qK의�>L��	}N&�M��j�IxR�0�}��!�j�g�S�8����c ��K����ۺO*XË��M�>I�l���p���灦L��/������v?������'�Ԁ�[�]4����^}ȱ���<���F|�8-���������F��e3Xh�K{�Ĺ����F�=]]R��A����-`���P�9R����$(Z0zC�=���.Q����{��{�@b=�T�R��zL���f�R�%�Jy;Oq��x�?��g�K��}C	����V�Bu/y��[��nD���u�^W�mOJ4�qn���1�ձg�"�e}n��!�&�	(���r�v���z9/�G��)���l�b�Lmw�Y��J{���1�����}������Ajl�IǤr,��vDV����k���[���O�����P��� R�pB����A_S�~�]�6�봴�������ϟ��T�
F䐒k�1>�t �jI���3�D&"@�!Qʵ��z�͘���Tj�j�G�'R��m���~�B�^h�^ (����"M�ڟD��c� s{�!���cF�0&��嫮�j���їrM��tB�	����Ne��3!��@�yՋF��g9K�~ ���7t��_�`&Ǹ	Z50��	@�{;���\%�0�Q�$�jy	�r�M#�5�u�7��A �{\�w���u$�B��2X��%(�<��$��R��v���fu8-��1��$L �_��n6w�QO��5&L,������,u�����\�.�I��mW2=ك�/&%1�{c��V��0�x^�](�Ku#Z���T��$�=b6(H�U�h7��N|���dn]?iX�sp�Y/1Qv}P
V��H��e�l$��}�F`7�I/���tL��VW�2*�|�����>�p���2�#m��7���$~O��yP+/�|(��m;î��T*���.%���S�%���O���%����\ �C����p�&�wS)�ψ?�% \�`�V=���<�����^>rM�.}#t��U��y,O�(Ǧ�����]��"�w ��H=���0�o�űX�?YSn��f�yX�d�y&�IuL��3D�}K3A�1�� 2��X˘��i�}�@ZE��Rf*ʝ4������
�D;߷!��D˺�y���ِč �dݶ��gA}*���/�x�(`7l����m~LL�;69��a]��J%=�w]�Ԧ�T)g�A1u�۪1�O��<��V��1�?�Q�vQ��$�����U���X�C1�,�P��~��;1<[B$	K'<��˯�`�%�}F�)%���vHl�f9!o� �E�����a�P��H��=�5�r�1����Ep�sz.�������ۮ��yw�Q֝��P@fj�M^���f��%ď4@�{���*�׶�^���^��5��3�sv�O���$R>>a����(O@����>&"�m�K�*�����X2�4��d3}k��y��S*灚˕S�^D�sm㓖�L�����ޝ�����C�D_���ݕ��(j�3B�P���� e>w���U;����oY�M��Y�}��5��))xu���mYd�k�X����g��>��n;�<�;��pf��JB�+XHQ�e������~���j�{�~9j�U�V��^��|E}7! XD�1���{f�lY#,�^���Vҭ,a�vՐ?u�nכz��"��0<K,o�Y��\Es�f�%�d��"�S���L��e�ʫ�N�nE�C?+��馉SK��š�[NG6� -�J
�2��$���U���e:u��[m�椶��-�1/��bd�D����~�Z��!e�^5X���c~V�"�����������+甘�肜p��榠I
�|#�A���R_�P�k|�6
�e^�/x�}(HM�IR.����fF19Ƿ�X�
�����U����/A�]9��u� K����PW��������R��E���n���'n1�.FfA�FaVƈ1�]��pW�g�bE�1c���f 5��Ҟw�q��$�,��Y���X�Ȍ�d�Y
lհϗhѠ����0��?�]�NU .3�;)_<�ER�X�4(]}˰��,�[`f�B�}P*��6�u�S�+���Z�c3�*��Rh/ֻCP��uʳ��G��GK��C*���2e���")1��ob��slC�0q��������q��Y��䵁�
D�A �$eC;P�s�co�[���A�%�6�盆ngsJ�ONs�Y�T2�(��S0��s�i^5+L��a�Ƽ���x0}�9b��2��LZ����N0���鍗9��Ol�'�Ǎ��`2+M6'��R^�mH����}�Dzm�F��� �{m\lx8� 0�T��׷�"ֽ��o��5ڳC���5�}i�	#�|��zzO
�
c���}e>�A�����0��]���p��i��'�Q:�����4�#�ft����&"�rG��A�X��5z?О*v��Dc���E:�����v�����Z(��*�{o����+t�