��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���c���|�Ɠ��B��P�b@t����EO;�g9��_E��Ybf�Hf�%���KPZ��T��-//�,W���$\�!��I�:�=��x�IL�߄���s����c��o�/��t�n�OXwb���Q�ME�n�t��ӹa�4UZ���g��?d�pf��B�b�E2O�֞h����/7�0x�Ku��fY�\��`�O7jO��u��#&d5�X�3�}y��Ǻ&�j�И�$U���I��Xvԏb� =���p?U(��(��N"�%�0�-�;���CF�햫qM&4IE�ZHI��; P����b�;&�V \Y��!EA�m�����l�{Y������"8��g%w�]��� ��/�#C`��g��;�/L���ݒ �B��i	�w��&�C]ܐ>�F���X���L�������x��{��K�����b���*a������`T�z��{�	)8w��7����d?���������X	�5B����4_����X\�^7-�9��K���!����jC��4��E	�q<TN����A����֯���c��3]���B�J���W��W}�g�=��-�$��M�~���e����u��nR�H���5����:W%{٬�f%�n���~B~���w�m>ņ�p2�i���g��;?�tz�OAm-8�Ƞ�l`Ȁf�lQ�ؓ�G��!G�/�^������gæ���l~g
LE�>;I��%���H�$�TL���	3�Z~D7Ēd�%"�hy2�Xt=I���,%8_g��\;��b��ʁ�$OY���X5��!�.�S�wX��o\�q"9�����钅$+��Y��ɩ��j�`���~�<9
�6�O@�;[F9X��?�'+�@/���;�tqi���YFC����{R���z��ִGT�I$q�k?,J3u�Zz�rTjE'2�n6�7S(�7���7a��3�5�& 8��"��RG�;�5��<��9n|��3����W�����.~t�ָx�)!#�Lţ��&./���<���Bt-�W�ҧ��f�����C*���er�!&��b'�d`��L�[)T��i�5
���{%����&��(-��2l"��0C���wЖ�R=���:��V�o1�n����b��� �������K��e�-^W�X