// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IiDHl3r3W7Y/3gfqqfg/A//lTsaSn5z2jeNTgHmplTeR/n+3t8qKm6BX7YIFvFUG
dPa7ScgeSSSnElflI/JlYYSxnvHifVvVfjpOQf8ICbhyWDKG/MSAe5Kq+u/UThIS
5MM2lqhE/CEL7Gn3HbPWS80zBQCmw0WYZ7xqMnDVjLY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 181152)
It6xc/rNDLdiosDlfhsvZ5IBUT24kiJ0jXzxEBiVw92eWc0xhti8pYSUEsjZkP5Q
wcW59aFpM2v8+pbTIL9GIbDEFRlL088SsKIXoHUfYEyaIDs++e+PKTX10YTzKeXu
nvkKwGSzBPrKwdtsxYYDRDnZih1Tb1PbNqpOzmdLandunte6MM9C9IsiLtnteU4J
8IQyntcGKVP8wggo4pUbPht3bBNPCw25ofcguFlGyntodgNlp2Fi9D568QFYZHVs
MuRO+ifK8Mx1mU/8761v1gFkoVymAeWy5nBfQiOTFqX2XeEWCm0lePwFlKWN2tb+
zE2J5mCxAKjliWRQuvuOveAuJ9ykVH3ZK3ZB9HmEPv47QYm38XEG5fqfvx2wDBUf
01ZfOM2fMW7pro0dHzeM7zclcO6/E50Ck3/IxCHu/crRwF339pz97W+G+0+5ZLFz
ocsV/IAT5dDS/YyQiRC5zmLiBoEWQXMZjs6rXAzBavY2PJ8CZt7kzN7mJ7B5ImqR
APSTo+7VTB5YqTi/p+bX/+1lCXryQ+kY+yigHK6mP1vzbQWYgq/nOs9+sE9HQ3id
SCTk8EGURO9vTyS2mUhHigKbnhJLsKGvPnhQqF1ANxFRThaA5BXwHSE1ACl4LUo8
lmHsEL6duMAFSUgKxzEc/WlGHZrei+j+X0Mwc9rf3ohxiBTRVJ4z2wezQLh+0HoL
1ID8CJuEFMcBFqMlhjP24vRebRIuEjhq+8y1d4Bkjg6o7PydiD2RStw2zRljTtx1
RrsfNft6zklDXQ1ffS5WkvKDLTUT9oPHeKkffCccpplt6jx4ebPJ0U8SuoPfQyW1
yRxEaX7kgA0zuTmxDYqr6LbjaB6Gqo5+eLj/2sS8WC3RBfsiwPmTm38SMCc8eDQj
46xUIQ0kOplhoUsgoduc4H5EnaBWvDreHS5rsvNClqEFUABYCEH9EZjBmjSCr/qU
CfnPxkMC5w6np6688ZdCjjt2wE7oI/f6jPf7ziSaL0OOkGGCB0VgJvIWjJ5fERxo
yYw5DhYNx69uzh8UEjZAarAD2q3EQjod1XgUtzwqtqX6WPH2oVewRdT44AItL+TQ
/wLKbFysbmTftQRvWvnMuNWq6HQC7T3Vb9dU8AfQY9zBXCxOpAPZBgY+IeOErjlz
0uqHuc3c5SXzVKL5AAN8peJtc02etdOFI64N3856m+ol3/P+Dw5CdQu1od1tmFdA
qIpEUcwBfS0huAGLh3Og9mDKDSM/DMIqAjkVigauz4QYMz+YESZtRZsHkuxdpvPa
VJ3S1u4mXEgbI0V+BxIfv4BaPJDyNF35OoFO5/HKJr/Y/ExeGImzXrAGB4EQM1l2
LU3wZUtrKreVzOVcw7jwlGQqs8Yky1brw5dOYxJhkmozvtMoou3vewbU1Spwk0ah
Xj/3bmS3L4mvwmIctv20V8CVK6GijvSugdDzMjaD+uo4zIXVVGaa7gbJVlrRY4aa
nrlkHPPI8+GE1sp7QsELQI+k8yxyM2f+qE6Iq+1S/dVnfocSBfwRRdSFQIZ1aZ0I
3Lr8ksjHJgSMTa7n7KaIt5d3MRT718xhdaLz4/+p12cKYPIGabCC/eQ9KQq7kJro
jgyWK5Id8sf78cBX5O5VqPJQxlpYVEm/oAnB+PWo0OddAoQFwXIkVM7RLQcV+Hkz
SNKEw6NHJa3CcZTKyxm05ph4DIzVeVAXeHJaYvWAtqLFLNLzjcN8rWxzifPouyuM
VihgDouvLQM29zNl0hdtXTrkos1ChVfPzo2GX5Dk3Qey3LJJFavtjM9ioVbheKBQ
p52gs55GpA5XRxbNRuS3PoezE6wSUyZIYMwClest5QbZCZGjg1FAlEbISUCKWzsz
jKWPqmiCaMBkQ9iRzIrlR4NKYa+mf5fPCQ4MUi1vStnerMOdsD0QdmZNxnwlceB3
UsmdcxLi23E579aiXS7Bkw6TxZ8IT+jPEfJOXH76iVIemivLaD6C5OHER6Dw4mgY
scpcjBCZAA7CR+6/c/T0p7puEHQPyPEkptQXP8/E9yhFQGSCAMwy7GVdJKgmfNiF
k5ztSDNjvREYNuktAg54ay9GRtktzP/0D8yIwfbEld+PQmCSM91FNeNia7oD9FSz
ZNhBqVk884Sty4x+XdTsMoKDqTvhrS9i1oFWsF04Dij3bJ4dLFVWnq5UHt43GxSU
Kz3Yi7qU+nHM/GjYTqmx+XVBIKzHqqfYJPvYpBT0cemmSuDwi+09z3iiTL3yIEec
RtR25cx68PTBNdvkQypAYNqCvYmuPIVPjst/9GqpOhkn1/Cf73QXZHT/c8JO9wZC
dnXR3kVavvKEMG3J4mrUQmHbtR7guhEErjdtajoCXoDuvoEza8aIh5/JR1oQewbb
htOH3UxIl8UJJhZ1lmZkRAfDFhmCNOql2RA3221nw4dPv3RpUQseXHG+Lo8c2Hsv
Mm6QwaU+8PO17llI3OwFM55UrmLAchvWJ5Xl5I5lQ/kV72sDHKyo+t2IuStA5xXG
48x6ce/kZXnXfNA+lVz6QqGSAFgUZvhDMNi65F+o10OnXu1RKfj8kVYtc5abxKKk
NzKMSW56LUib4mUbKgL5jL0M42aZt2+Fp3SGEoh73+D36TIQ1q6Zis8VwS5Giu6/
zWJEjQaPovNsiVW05H1cGUT5/0rVvoToyCywJou9l1qcPYtJmkIMSlctUEbZ79aF
3lqVikkX3mr2Sel9WPFr5UtrNIMfWYyA5wchvNqnwB4D7cUiOrAitmzE9V8PXcq8
sob/XtV+0zFzU2QDWiwwdBPjI/WPzZnzyLLM/wM6e502+5Yxx48qiSrM3BXC4tq4
MhoGo8bGcoXD8HjJ2b+jO1hE3LwugtqR9n7mYYuJGP/0F8CvmUduWIfySE4iyDiK
91mzziAXe/w3IEpBBzDYNSLtUdo88Q4NVs9KdcCUTkq/V8ZolGbwCtkOkfPtUpP6
G8fs8zo/o+DQyNZvHd7DLw4Xs/s43YvIfQ1QoBydxCZLxmrX+OgaYYs/MwHs9vHw
voY57kNMy6macnN52VgC0T1oX6x6xFNKakcMZFPVXuxF5rHP7av9iasZU3tkWaFn
p2IH+RjUnmnX3Q21FkcKoP7vZ3zr6x+Fx4TpxgvxFXY9Q0KBMHfAll27MRBsaQTJ
pVWHVsZs9oCAAqEa+3dadA5RW3Tk+DtaZGJDr5bWZA54y6NClqBB9MJb0tywt7Hw
PkjwXAaF/T+tD39yqrWkIuYDiCrfgxqzZkKpPsIzRn+5naMEnmp0OcfTsdIHPXnG
tXE4JSiPm87rLJQzBZwhoDyK5IGp9ngMABPlntAO3qsvmQvgU87LaYY2oyr/YnmA
JArvauRZXVQvByF8swwQfllA6uhsdBp4WWOzMiMnLMrJyr3YRgmr8Nw0X3bmVN1t
IsnFtdXcfJHBW+21zZw5SH8HAqmdnUOhxXLksEzZ87Q61z7HxBAz6KASSBoWUKCc
ZE6z1458sPBalkiokFJ4hNMSt9/6roz2l1jxvBT7frliG+SUrvM1lGgetPNrXCvq
wuDtd5HTI55QxOIxuGvnDPnFCZ7yE9BkPrGdrbAt+uf3q+0XpzKvqlFxik/7HpNP
Du6vVqnAF9ADEDYL0vRq9vCRyZf7TQ7o8fnizORRV9/x+7mqeuRCbzh97JtoPuyt
MVJXf2DGAvKT3owQbGLuMVrCQlq06GxomAJGJJKNFLUzi43KqmtrXMrxrxCzj+Bi
lgTNjxoYBQD1E0fplV38PtHkIyLMk55dibmAkVMIdkpvvrmb2iEiPD4ftvxTyf8i
3VdtD0Z529KSWUz29i87yQcEyR33grbSkT8aRA5J2QjT1eU9CpoWbYFuLcLqeyWa
/kxd6U+LcPPvVUjI4n4T58Svg2T1hD2A0bdncaAhBK52V76vygcAOQPp/Zr9YcLe
8ppMnYJl7V6EPVpJLI4yhLi/fXEGbHY3X3sFlwF8A8DN/bxfD9A5ZdW4X6yhNUFK
qQ6ESTlZ3cR2OfyYFS9iHCAxediO9qHKU56/qGbdAiseDcLdvSzMXVYX++4cZyah
c+/3NAxlT6FEF3lo0/Qz/mRXjHDiiZHyIJCXxe7jstw2mTsFGa5wuNUjuNIbuovS
Nf+PRpmy/zt//w3Kf3ZyNKLkCou2MVY8a0Zx7QUenAc8q11n6wQq2v3hbRxxcDZv
UOvfZ12kCGzRL5+cCK6GVZp0xgD/fUaeRwaeKytl7slqiJjMhTQ8S91F4QznWz5r
2b+PFTxK2zjW7JQeZhlSa7iZ9jgygNdC9ocdFZteNN3ZY/gr/MBcnHeZnVCm3Skm
7mhoN3CgzwYVgYC+a/auUv0C60YokmuKLvH8o2FvjRlMHzrx3uYcanei84fpksK8
Zu6CKDDzZC/4w18nkKnMdg7uRk2GVzHJ4rZfkHxnopqeXtXRE1i+q0d49/BxrRJj
kNbLHd6JckUXYZKJQH2T/U7jkJF0i2JXJzIxY1ODMSSdlC4IvCUXFMZCCQ7nXNa7
yDrAQ6pX1LCWW+uoR8TlJ4XT85JdneyP74gnoHCN5RzXG5vKmYZBE5WeCnCzGHcR
wt8heKiJN0WJsFAqN879p5XlLvXMBTdgSZb4mfUwcegvO+mHMhbRGbIL7hyCxlEe
Let2fGEJjGwQLRnknAu69TIe28jzcR20AIsbE9M995idUAmmk6yzIEgADt/2NFrT
U2oO8t+BIqMm/0tPIekHOLvb6afrStS74rHTvnVDcc+gxuGyzZpq7SZskMHuslIZ
lZyfqpJRjc4zuLaPy0YOqZ+A8EYcLd7fmIsG6fSAR73Sl8msXVPmsJXl1VNxY9d7
sXdfCNz6pgNRhmQWS4F3OC1lGuJGMJnMe63wiTFT+q/zlna/OPFAiyyiKELk+I6q
W+W/tayKomJiZyi0RbsG71mAhzK+5pjvUu6UJp6B902snUVEAjWJr2bfD6jGwuL/
3c4vTetXnEBW83cTfui6/Wu2Q1xgscVT/5fCFKMkwcOFd8f9Gj60SaJihDsj23oX
ibeIAdvidQUw9AE+FZhd/TJUX6XKwBA2Fg60u2rcCtlTdjB440lBz4LXmd3skWsh
aN5LVuHf6AIYk4Oqcjja5AgHQAmTx/X9E/UJBAFYyFTCL+2i5QrKnipUuOIdJ7LL
1KRnRdK9h7ciobzO0KNHz0bQ+rhi8ppou2F78zaEZvGa9rxbMBlRdaLPr92ZW7kD
9Qm8cavo2j5I4FmCo2I3VvhzBwuO/DEJsrEOCCWoTAEuD9EMKROKlGUtiOKYaynC
9HDfWQZdnjJf8ZVkB3kmN8kEu0bGDHPUhN47oMdTXnyIA/6Nt8a6mJ+2vWo2OljL
tKoq+67sVSOikZ9AnkoXyLPpfnbt96t9cHpWCCTAeWJwltdFrjbvXiNQqDa1x3yW
WwwJJ6pMmDqw1kfm9hrHN0zFeg6oBgOu5PCiJNWPFzvpYLZv44ksxvuzA2hFSIbY
kkkat/0lNu96Uvc6odex5ljXptMCXZQ9CqYGkeR22zNDOYxAtKiI1NBd1drQxzi2
xnEokvLnz3bm3FY3c7pyN5N10wxPv+qBDw/5xqZsM3Zb9MscwgftgWxtjMtvUL13
/wDPvXTGxf/dMsc0+djDvUR5wKPShWy3LOrTDwQP9FOjeiPie6/h6BWFOIWN8aCI
vltd5mXFCEtBNOTMP2rCYNXXRC8L7xXdpauUuX4yq5RWdYQ5UOqxJD6W3COtix19
ux4h1OWeC5kFQyF4DLhXNqaEIBuGIWJzQ/N3jRMOPAZhV3mDJgm+Jo2/LclOTrsl
WJMSYHs0Dsc97emA/mJWWB/7Jh79JSFuMInpgTNX8aT91edp47az0kPOZA03uXSE
WpqB6j0k8FwK6D4Ae4UR9q+CVOQKgyBZOcwjbRD/Z0xCGPKYD/XyQrrs8fI1YbPL
oqHE9DHfexeiRa0bt7tzlXLlzTwQoOTAB5bbhbJeMX659T5cV2CkOcBngU8elr7G
oSpbRnpZTKHPBOgFwrWL8973PuOP2NAcGBjYkbH61Rd1H00SrqDY5lezm85S7jgM
c/GYfXTl00Q+c2wMdTNaElqTcM79BCCzNzwXTpaOwMVOZUgHzbejHkQUZnNz/GzF
fd/4nNWtfbDb64/L6QrV7z57En4QaSKxU3p6AI15FqnCVLUC40Uk3tpSs0SZT2bu
yQ6U7+3q+Kh2OuECz+s67Xql/KuiFsIdWptIDxHfX2O0Y9N5UU5Y8msimnyzK/sw
P8/m6abxHKURV5IhuajCgV/D7x0epBtF4OZbQdYVfY83qkKO7corGr8a26IhZxWR
BqAxgW4XmOH5CgOuXAwkn7hv6B4e553COHO09QBhbgypSL1vAoNRyXZ5s5EXtxmD
v++wBkxJ0zq/Mjg8r+4E0vs9KZVBhlN1WVide/2mHk8LK15VxQenppwyOfnGUx6b
DZgAtElPgo+y2yROQJdYYKYcCaoXvlfq1AprtKp2uZu3koH1gJSRBjkxQzOvVAML
ipmFLJxC0lRIs9A4aOA5ueCVlBS0hsDfy2B4Eit0C0P8+1I/o2P7325A6vdR2FZT
dnSk1XzF3uUiUrGWjA4/RVOtFq+nvaI6KTpA1r6NJ8aveKq72pGZsyGBkkeWU0Qg
UNJrHYqWEb1llJJAQfzrlF0oYP94Eed0zkGG5UPH8DJzcmNLzRcmQeZyGA0lzEKb
s2g3AFIBhxJxKZxzswGJq8SnyQy5TPjU1qYGPb4EHTKdnvrwAMblvkITpBZaghFZ
/wqjhxwwUUcE+Vs9FoqbMX27ZpsyOXU4g9wPJ/gMqRws5RYpbCuq+8270OYgsjBJ
8w2OvjYherlcj5r/hBRG55w25jKiGvyAO69sSOjV9yg66CfaTewUDGDs27ZyZsRE
T90ezzFJP5luh1WQ7FMQRq/mn0Y2DqyNX2zfz25ZDU2Vv+z5HEblyX//4p7EfehF
hLjEPfqc2ZHmIinbTdDIIh2k1f4fVbqZyRvtgzww5sq4wyTlRhj2+IZc0DEqR3Lv
8L5BFRdXHmkMDRxPuQCpya+SF6S4iffQ8H8x6rq44R0+aVdLzna2op2w9fT2DpGj
P7r6zLLZlY1yLAgc3gmLQaqBSH5JCp3xpcegadHs0WzsZLz30o5GMHWDpor7hQyL
gpR9S08ylfkw0ZHM1yD13l+Go0YcBbp2/va9UoION9NjgGl67IvwrqQ5qLN84CAb
vgpAA8VScx15+/Xwz+3cZKDV22c93XkND3KOqCgV0dzAbkuPY55RcLllWXF0lNFQ
ZxgHnimYmZi3DsSOprjHzoOaONHP7guDU7THoHj2Kk1QxeUrGFwlDVRpJxe8hUtS
XdF0Kzo6CsLgnCoccGfU6dclDqOc8/bcRm/TRERCkoGghtbOADQr43Plik0jFJuw
XcbvejwsjDoEEUJIqRXR8BD3ILfcqmupKi7X+j83cj9lR/BcSEGhqQN6xlfDDH+z
WBbjveS4PV2LYmtR5HNcDa8gwbhHaiTpbhI0sb/oJBoaVF7f71zifSGJLw8TnVbM
BjbYbGJaxqk8/tMKwKRw0xXS7qtr1TRwJNhhUfQZ4v90E1TG68nQsDH9KaPS+JIM
YoUCXNcwZZ9fnf+28H266ADBn2VOewBC7fdEI1HGVqq0xj6oRQFotOdK7TR48QcT
JHQtlT1jbY+F1AToZRWWan04L9KRbkrjWt+h4T1SVTV+ThreI7Y76nYd3SsdoCWv
SRMw2h5NIukevdaAxN0Ei3SLg7GRmEn8sUjrWlns/QFF4POnWfp43YkXTjjIRPyl
xp5P0eP+UMd6QN3N84X/SLxrxqM9/BNVX3jAWIMWtWPfbMVo5YTMHTXx6Z7m0mgo
qR/RNSxBWhso+aW/q1PBebM+Jw/RkcdqAZwysbWFNOLzHg5JERiPNkivSdlcbtu2
M42z9AkLbVQDQ8ghC3zFcsqWFgn3P/OyqTsK77LmIxakQfmaGLKIH83dIP18SIVG
zo17NomNbAjGi4Mf4eT6SG2CYP4Qi3gKMbCZsN8Yz6RE6F83MEhO9taYNgZLfJB/
ohl51sm+AUNyDCABM7kM+OqoV8ijCKVELOhQLmzm3wIMev8YeyTRHZZqy8Tanp2F
p6YRtNvixYnQ+jX+j01cUgMAlqP1pNtzgUo22IQL2nhbZH5O5nt8g2jGermN5xme
pH49hiIny1708Pb2orDrX8lS/eVrHcTNz7rQbo5ak26JP3rh6OduWfeIXiC+4uH7
k+04wd3vOXSoMTKw8VQ7AaAb3alUF1OUWAmZMs8GVEOj2QrchYwtNzO23DZVK8Wp
UCkiny0jsGDhm4TuElvwUhlt2ALVH2KDSO2PLH96eA7TLCefaF/Ng5rMC9aqonrW
nOHoKIt01ZXjPE/Dig+4LRMCfIH/+GV0+BaMeDG0Ne8umT/KxmSEWOB2r7+0twyB
t8f5p3NAjqt1XEeozVsSkKrHF4aFI01FJQc2b/ky9DnhWBrZkiaDHLfdO1m93+2A
vviZlFwG3WFgMAunH6nRU32nYCXSLzCnnYhr+LM0+0A1G8fB1FDsLafW3YoUD3bm
s3vUQjQLMSEbnJWOwfbpp9zymOlToRf+rc5FahirG7ZGhCGSEz7ccOlrsD3SczlU
U2VZP0ydnR0L+TG4uMq5TxdxzJ8APr5rXUtw+0OSxZcn43moZdzocwJdpBpTMHmV
wDPdID1wPSxfDwEKyG2+dayjPCxxaK+PYjJq2cWLdTSGY1kr9lrQSowedzZAmqUU
Mgh1RNRTz0L8C3/H92zaax8RcErnnX0s0SWg5eU/GhhD+bGt8ZmkSHYJ6h9QV/kM
u6bMQUqlC9C9gQplqb6l9DHvRRQ9uX4ldfkx/st3NyMr0WaH6JOhc5+GZM3hjbCb
DuP97G4xRLtRfLAgHPSjtTkD9tuFHcM/0KI059cYZkZM2Y++YfIZnT1hGpNJi8bd
x1PGpIHGgcJH/EzI8rJwS28SAbxyocE17hZvoQdZXGJDpDxH/sTkEG5ZyAl52IFq
j/QOIi9ydTorl9rOgJfmmvvmnW8gflNLa80Q5AeZY2Fjfgzs5mPeQsRsC5c98WEB
LhD9VWt23bV5K7p+dOw9d6ODMOMDd4/Y0VgCuVnS/dhi430B4lw7aYzPD9xrF1bA
TWubf4yYKzFRzZ1yVkzg45RMONTZqMAUc60ryq3fLDtcZR+rlyxiGYNLXeBcUJM+
yaj4bR0533ptgogzZjVLADdDNV13pzxKC3G0YB1POOPjFkMveYj45v9n/LaG7MZs
DC+VBEqoPxOhKRi3Z+Pzm1pcyJ555fOrPxT5kRoKVG7gjNIG+6ECNDJVXCcyWKve
vEpZ7m7QgXSlhjADLdDvYPhlq1bJe65ISjVAekRFVtbqIWpbziaunIYYaBNLXDuw
r48/beXNP0sPwztZ5e/GKicJp3AbXXLGRRGR7u0X+Etu5VjCqHIENj+vkA4mEGUN
eTRYqDQJL4VBv5Z9ocAadtJFtjaweVum9AywYWGAsfxS83Tlp3zMd10CX0ZJjVbI
+b5MrEMn9SX6rzQHnea6C4paIMCU3sKQ1UAmHkumz+Qb5F13cgx9Lq4it4TXH6D1
aWCNFjWwiHzqBf6iO8qymWzIRlI5u/KlnruQQ0vEe/0oHo4PUCM2cuu61H6vMAup
FTsxN7Vh/OERFI5L7yhmCuvpd5WOrbFy1veRy9KphLay/xNP7OcDxwig5Ugm78TK
evv9n0YYSRZomwD+bKg44mKHzO7wCKCfogk15+SiQnJwlF3OS4mPuyhSWVFWPCAt
QZjlrboRTmNNHM92OLWFuOewhbmHIjg6Nm4JKPYiHJJDTzQWDCd8Ux4RgDDhDeYW
03JSUKuBJ6jGS+EWYYW1yA0m4+zn5nerE20+N6fbSzbY9iUpq/4j8STo133Y8pvL
+PIBJnWOVXp2HVPPxILxfJCngDn4lmPffGaqRyiUjrxyIfU7DGEYQcXdgr+Xfgd8
x1CqJB4JOMkIt1tJJUwbfBy+yh8XNWXeXtvFY4kTi0tDYQQIZsm99/I6026DOiJB
8XOG3C2RRGmsTW7wyAd1gcJnoV7zDLxGRqLQn8K8TG2dvJX/ygNHHPyqsllKLdXl
UBr14UCMobjv2TdXldmy7gQEDDxZs6dCTQOJY75ZK7R6OONG2Jov6e6BKvH8vg7s
QVEfbiCiy/Jv0zRePsF/E7DYJls+A+mDHzTivqpd99XQVbHGwDltxw0jMr4qUdZY
bvxFT/cpNzrzvLgH/rjGPBXsBWZZu2JcBEvhFJgrqvE8IlNOExD7ZYIkPPY/eOFY
sgiBzv+BpI51eRBgoGnde71UN65alOTdTYDZ1ObD2riyqMjjwktVfAN3KJVOWsAl
U+NIklEAhUt8u2x7tYsTzl1BChLRBJT/nWl5tTdnXFlIlt5vLdYplpzIGGmCwE2q
Qd7ePeKwG/IBD5d/Jjv70mJqY6QavwJhraaZvpvyOk8/ZspXuSrCpCR/8KYBLQdB
3aWkOd2NoVq58ehwyE2AOp9O+25OQnBlsyHCExBZjOByje34VqJmIQKsbd5ioh27
aEbf7Ak6zZM2YlBGVMXDLzoJOZzYc2yM4MRIcVqFTw0ms8GOJDiwrWDbd1cp9C8x
JnQToOS4GPia8e+vUgslyeFb1YtfPoM2++O7nuWcCpvRDxraBYCxEKRzhFAk0sXu
zH4yxTN+PMUY0H/Zr5EGrdYYh3C4ILBfCQmKOtyusP4cDG3kZIonFYeuum7l2E0Q
VZcirsomi2KxOOBDEz40Oj9xcIuwxeWKlsOtI6vfW3zAppdrCCb1nxCIVZiPctmM
4JzHxVpBfiYC7gQu2V8oLS2Jj4UqmrG/Y1j4XFXGba91mEf0LLxbVAu81utkNxun
OFqi4NfSI2pt/GTjp7I8jvig5RMX7wtgtXdd9rq4h1KrGVbUtmLyNHKZOc3HqsJ4
5/OrknvFQZFfKDb3WGfY3PlJdV8ZSUQ8Zb86c/C8SpLxLWTZ/YsGfcAl842JRRQ9
DQtZdPhFXzEwTNq0RBXpF3+AXA9Mf2pkyCcBic+nQWz/hc3kstEJvy5MmSzb17oJ
EMSbM1cLeVWaO7N0Kg8lJYgKvfp6otM6Y6kH9Z7oFTvs0fzkbqaVFdFBwIBSo1Wo
w1dmta96N+xIzbXc4UiXhLRytibJ8hrpmClzhB+PiBJfhZPLjuKf3bZslALJ27hC
qaTnfAIoN6Vdir0DRyb3B8urtcwi5laboAaUtjAZIa2OXg2oAfHU/eXMRHR/b4QG
1BttmG9b84yoVssT9COS/s+fkr1RlC4x6sHDrB1yfIUXyC3JlxjOBDTA8L1jV/ld
6h4EsHjAwpnWRYKW3NTgo7PyoBzfupczvyTazc08SHtuBLPswG/gfzGuNei6cCtH
GfSOa7Hj/Ya3vlc7xv4SBGCgHjsWfCaVE/7j28pfgQQFV4cfqYcyqzypjg44smi/
RvnYTSlsw26eysnSEFOWNY7Rc+EjQH/UAvt1rzO54ahnnm7Vc6YuqfaWq6LEbRHV
gUjZEBe0TMuUzupYk3ty65EgnZV4rQht9W7HL9qjS3Qlsoi/zz2G3Tvkyu5TapDK
acYa0K96BEga/YUEl26PcWOB47bXB1tdWJ7bsq1panAFSQbZtPw4L/7dwZMK/YS4
xQYxTCi07fuBwJqk5uH/gMRiSX3sWRiReRE6+gseYsRfgGZbbhYtwsxPttCWDhrk
ZgllLDkzKvjmzB0t/DzfJflk2SPLD8wgx5bmCqeAT7dJFEEbLe7SisHFqW7fzLUq
Qfqlp/wccFoMw91/el6/TsXvgHa9Dm2gptQddyWUa5NkVAIcP9cEEsubWLioPML9
D8CcF8fSlL/R+0FjOaKAp+bCA3TMslr9zrHA1jbfRcmPfnySFjpCV63LF9/P6xnK
fACo41tbOJDBthpMuyZWnHWOoeGgThLTDOeDtD+m8lBA+VzMbhLppxSJ+ffJLTQn
nlb5jVo4GYgBk3buykqQNoJhgCGfWgfq+P/YtjkSJcfyhOK1uCxCRd8Ncgje4IEw
xwYckk7sIJGkQhlso13r9U1V4oTxNcS/uczbGTs/vs4s2a+SjGwUn6f+x42U2qSf
WcUzz1IvT6EYy8ue4SIYIRgWSiT3XaazqqX4glYtZnv5i7o8USA3aCx4ggaqgPvg
OzZTMMKfqI+f1bjcUcEDZeiwXYkUgFqbqgtCfBbUGX9nYKDL1nOoeKRIWJFv3iaN
bssAlXlDfYP7rCkpW8mHc74Vgg6eMq7qliQkYHowTpkacqFnjE9+ZmniNMdoOfst
VKe7EYSdanTS/MKeVKcKrutY4GyVLqpGYsZSjcqCdEBphcq72OHwZra5Ml+KSefQ
Ff9uANpWn8Fz5CRBuyAZxsuoheX2k9HYiJgWQ4JP8Mk1fKFELgK/lZsaFqu3ElHv
HNFRKMu6Le0MjFxcCazOHI1j/lKjIHpYli4Us3dD9qexXWNDVKZfATglKazWStVO
UWY9nii6PWP4LRZcBlVX4qI5DEx/7+2kCDNQ8DT7uViO5E4FJGoENvzpWaKwyKzE
obO8RVqSMa0/DH4HZ9u71ST6FiEzIVjyRPd7cfI/UksXN869upmp+3Taog3fl+BI
FfYq5p2jFPMTxqB5AuZ3gRZDmtIdfaZHGKtO1TV+p+JRWsjCEtfcaQHTCLwrOnuo
99obf1G1niIs7Y4ec+i3YLVjeOlf8gw7y03qIfdrij/5c1Ze2axFUlAud8LaN7FX
CePu4GULXV18mZAPBDq98EyKG5OZbgpdKKf/8EKTre4BHuFvQYS6oNrh78+PP2ip
enF1NdWzNc3UORcunVKmMzEqFA4tRbrd/RxkOqR6b1MjktZmmZTmVQwsmuhnWIMu
VXawDzBWPqBnkptUoPByI4hQ01ljNa2vTI3WY5hpV2XUkX3FDeukjUW76ZycEHyq
gM9yNwKjbqhnB9lSfz1NBEd3a2E6ZCyO7BvV3C21If2jqwN9z2MHHcm4thNYb0an
Ni5niFgpYpgNvftRl/+x7g55p6Mqq7dOlqvKgNoRfdVpCEJi0UFxpIMqSPE8WQxA
01K3QB3lYJ+r4A2Y6HgFXtIhnHv6BAK0aUEyBeJ+8j6wtfTrLjQDmiSuVs3XQoD1
nEp4vOBej+JcHtAEtUxjO21bQKxI/eb/4Cfdx9l4gMBs7LvVMg8aj2f/rr0hQckr
Sy/keRSqdjvadgP24Ip8ofIyKdmq4q3Y9GHzdWtXteww713/AKk8d5ffsh6widtM
zSq4t57YxlW6LS4Kk2qxtDkDW7yCRJocZABu4bBSv+aILDNyxKrGo7Wx0dzgOK36
2qMWoplvbQUpr+qc9GnVwi4z30vRl+v+p7l8gwL8ThPzEV/ot58vpjy1NB42w/6n
WwiJTYhAhBA6H8C8XjWONIy6HL8Q59dfYA2bbak96KwNUySORfKMFKfwoJ01UAvq
s1YmCPZ3l2CapDZqYYP23mZakkYBLJpWyGdbUfYyo5tP5Q9l2p/qSmmn78d0wRk6
mfVWRoFSWTEQVZUaQETHMrz8/TFVNsjEMVAcJi+NWGhQQ0O3nlm4SWmnG69prSqD
UrMPHNbu6jkRg/sp5N8XR/nLdaA+dEpPjdHrHmYi+sQ+R8GF7e9My78bp+eKTq5c
llB+GWCCzct0JaZHzIr+JpqbypDkwmmg2kN423obgz+j2N1/etE90EfgQtCGg+sy
1mbmkKop8IoX4OiygCcOAYgIQ0WSW4GvAk3v+aYWmzNstnFiPCNnYbYGXsLm6Rzx
iGqBxKOAq5ZRpR6kIn3pdR3fr2OccuJ3P24esP6eD9MTZzmngBMglnQrAhut9bqX
m06ZtxSA3GiXxY8AvYpm7KdtW3QpdNCTZiUczSY+65W5hpEv0lUkRaizWlaO3tRy
6k/HG1fkLMG3m1ee9rGYupN7CeHpK7EFnVtepx0A1HXHUXiCAK57KrhPHFJH/cQE
oVnP46YuXgXpuVeSfdMh0wQm2jewnn2J0HAUZx3hpwjed3u6H4fksbhdKvJVbUoc
n/UCtJfs9YVBLXsUvYPwbz5s/PD0NvjdMOMg00LyhCwUc4bJ1h+Jnq4Dz61DoqFr
0iHvisqCao6ekZff5p6Xnvw7KtJEedRUYqg6OaaIWjdhqcV4sVTiQy2mqmla2aTG
/59SlFglpz7QBehhBoeg31YfQsG6fBLS2EHUkJ9ufoEIszCnLKcnuRDzAf+RdbSR
IlMf/xFW3KDRgNi6d4mernTgKrCEXpc3iL+1ccMfRXet7VT5m9mNbhqB6OT2YVo9
hG2jjHuIkCfW7W9oNv4It9dAewKIxOIGBhSkSZ/vaD7+ow6bFeH4I+svoQEmiTwB
BIM/5bNKqlvQ47qfIRDv5oPdzZKag8T0+pAasa5EOSE3vN+Bpp3yb3YbbIxsWYQh
xPFJZzeFHJ46a3obNTahP3tE+4KgCssANPblEZwAUJwVaq3o+qsaWKhup7YypOhf
ll187U7pY0Mc+Rm04axhWCqPk9YljLeBzLqypBv60smo9sIgSJk7Ijk6owfMuI99
Iu7ju4Kl0KEF+GmioHtHigxHwj3rV3Tq/cW0mxGZOKLIiueBGNmvxLudjuJx/HBZ
/uYat+B0Web3/64P+x7NSlGdMytjRAL5HhlYMsWsYbDmzsdHJteU5/9kNCXow3++
Yq293y3k0YIVr7iK67dEoWd2yXBYvqdZDCJVCB6vs961wOgfLAk6b5Y0X+qDFbgv
ekU+6kY3CjthBobFJpx8mIs6vCtHX00MYH6stCTzznQHhENXDYQp77+iVHEuVHlJ
OutqMP0FZ1Mc2OZNALiAGQd+JNgK6c+sCaOHK2LSPgBG6OnN5VU2snGQCtPchl6Z
PV25Ujko6AO31fRG6qxXTgHc/nMuVrqaMZIxJ3Hel7y1uKvPxez8RJSFx76ePEZ+
fQVq8tc4lDu7YM1MAFjUdvdrDtdynMelk6r6jE5XiXz5FglSW6Eiko6NiW6ez0D7
uEqtxSnRwZu7VjyVFh9ogqqLQx6L4VUAqssEAq7tRG5+dDyyTN/NiNZggY/+CE5W
A6Rc6v5VxU5BaiPPox8AdYy0arHXJQM1kRdJzazBmnosjOtDMCPhAGhUhNKyqyxf
cBvOXs+TAXKCOUjD//STf3d7Bn2bqAzA0dOtsoT1x7htiHWsuOhABJesoVOS3YEs
CRnK597CKh3xoj1IHHY/xSQtyoqYSU2He+tFg3RajrjQkbUXaDQSLBqki2wUCEwH
ZvvEPRo5dUb6HkMtXCHb3O4rDVJMnI5UJuBFejLpzkPGgEnhl81M1u/ap6jEN/G+
xRf72aL8UdQcXvbinvwx8FZ8opJ2wxvMe/O/gfvIlue1+GkWaGdc597yBta/jlK8
vXMYT0Ug9Zt0q3rEXwmKS99JjQFVTqzAKOddE8tm4sQuJcviIGSsQ/8CL61pp+79
c1HbYAwhsWU+qk9XaylgYvMMaV4K9+otwAMvyOzlkvCG/4VbG6b36p/AUbi9UQRN
yxY0fIFAdTOApkwJ7egPt/ozb16kPHh+/5CEcBgW2h/ptN9aqtebBMBdQDqKO+ah
9CfZU9u97s3kak+hpoUqGQ9R7xVxYVs57KNCH0rdYjTkCW9KNOMcHXJTO8lFqzcj
M1UJ2Si5NIoh+D5T+H9EUcI06X4waGZ4GjHm4/uFcuRSKGFZ2pRz4+uPxb5atFuT
rAdVsR16OfPVwuTl0Xuf/PufPemAnID6PU+iaBPEu7Wk/1JfjFNvdkCSO5Uyakq1
6e3mi3x8ysonSFqcsBpBd2hGeeTrcFz90wThpqbXPHOs0/Hk5EuoJiLKoFNGsCrX
m7nCHShyI+r5nH+IwfzinBxMU7BtXINikXE9Wi2mpdNVQJV6qu73dHYtUqWj0JO3
U9FDn/AMBHk9+3mtOd0dWi1dtzoDWVpIF0Dz0EJreNJ1MfsIdATZ6tbmCbttzxxX
DbSihKpHSzq3PrptfhA+uLogyuI5k4cl3HcjH915h10Obp07ATEuhTnrbnABvHuO
f0wB2uzb2zYtUQDenuW8iJA4bvnOrq4YyeSZQDibMLWn5Epzi7shi+i3DT13g4uA
/fHmfV7M/fETZG0MiWo1+KxY5r8OeP2sN5zrV+bZiruvoRiqJxWAVZilMGBfdAD7
1zFxtcMv/qvgCK9B9J7ayWbpL+Kl/2QyjzNaVRDHRKw40EIqPBK8Y/afvoRMi1Jn
izDPga3IeKc95j4r9+INWT4BVPV7xE6kc5Kq+gsZG6kvKyBtgYdR7LF+eYLZE9XY
GPr45INS8nCbN5dJfOMOP42Eyfu0Cs2jWtcq70TBPgi/+faECJYOXWbMTsDu6QXO
SYktPjJ/PivFvBr1Jf0Eh7ky2k9VQb0+QHg/bO5FpmZS/mqS0S8wMHQdh9bfMoF0
67VI52nHH7b3FpAQcLViSSWxSMChKDGTt5XR3CS4pQg2ijP4c//jRUF7tdif+rLB
KLkC0+F9zfemK59h0P7LnyX0DviqBRO0R9pN40ijZEM01o0pUAx06D0HLXK78yt9
ubMjnUoaJ5jcv4dmvk0YelHcBfBZMQWkVxQpwu61lUr6Q/MlUkgt9PHwGGDXqPnk
PK8rxivorKfCw1vf0/kYyl3zyphtf2yDqpax9IPF9hYjkQ6zRTHFJ5hpvovfWysq
kZvLuVsChGeEnU9SYxPb8oTOW4/7va/6Hbkog9Xn2pbmiVkQwiKGskmNfOfsCvHG
h+H9qdnxF3/b6Q/bakYeExgDQxhPMapoBJUadUBoKFgfPSKfAYUqwaupBy7m5uJe
6p6CS5a7QhttCNpIh0L5ivjg6RU2/g0+AyrbJfcz68DvfQ0eSE+TAhrK0Osxmt2f
h/8bUkEciQU0O0OzVD/MXe0WALqqYLE+zoJ9UNaAwpHOTntyGWX3AOlG1MEf+i/G
iiCU1q9k96IFHm71MP7UlrTIzAXqbwW8s4wtVUcQ0wAqEvi+1G5oFokf2S05HeZv
F3oPqQ+uGopwYPdOZbx9UWU29P2GZVi5zbnzNgWQnSkakOkHHTkM/RBJyirmzj2L
FGvFE7zjpRxwLt3NP8K7kvIyr/PyDO0dTzG09BHp8GySkiy51bAmvf/NNQ4S8mja
wsiWs9iPGByallJwWMuISxodqHkg69fCrXHNRPsu6z00jpWTE/ZhIeks+gOwRV10
w7RahlkyHwn6fCwK6DP5b39JWFCs2rOwgU3/vVx95rF/sR1OMUZyPmmGBP3+LEKo
liFFXVhnpWADbBfRIM6PNTGsn10M40Igp2LFpoTUUs4HQ7ilZmcf9eZJ1Pl30PUd
mm1bJGaY6Mb9F4rLBZtZEOfPTCggnysSR00ZcFx4xITtvNSc9YpvdCJfulnKaLIb
vTtaLUDlx3cxmDwVNFnD7ZVG7L6Z6k0oMRvsvtSR0qzWnRdEfY6/PdGVY2XMpz0F
cwhqz5HI1KKCXSicPTdjKLivzV6QBFRH3VMfWocLJaAScVFFT6ZRzDI+/Rd+0YAe
93OCcByNC3qNhjkkrdw9Dt+bySizOWDQKZSNTUOw+IT7bXGSXCObftREGbad3fES
WJp/iSXD3z+sBP8WT4p1C+qar46WpIcxGh6SYRGhacmibyhr1BHqCPyreSXEVKcS
eKINevklPCHVIkCV6MqBNt486eYfmOIbKj9yU9woUlQ47bWBBGn968GCJrbGpbtM
35wYKpi0fjVkOPt2amdKwSq12bKdGE5rSxNEplBYilkhpFV/ErIRgLvwevBqGJGZ
BPZYvQoTL+M3VDla5SPpspEGuobvC3YRng8ztA/dTQkMT9UsRJ/xWwbxUIizeTsu
aAFjZFt/Gba1dJUuhjxBz25+ksDXeospWWpX2dcaC9hMMWaWLUgVCg1SVz0M8/dh
ryq+h1IjFG8ZkvJ+Y5kMYahAf51qNHltjT9TRCz4Lz0cS3P4re+qV6pZnuWi/4xx
Dj6Ftwqv63NuPaQUN+w4kEwhPu2DuvEtRL+IDSHKXl6i0Wl0wv0kCfWkB5v4LFwL
Myd4jXbeChuQzHQb3oUQCgwHVIhBflSEMCGD5bfC3kAS5rddfEEzl4Ww4JikcwA1
aWwnZZOS+k1RCGD7QNti2jyriYEM2LZDyu2jP8uuTdj/UC7UZyK7eYhv7hRlZ5XL
m4KwTCQhwx/ioXhAKeOVTQQlI9rzEo189Exdy9ESwwCHFCLTK01JUHbd44zM/Adw
Whkg/pMOx6miVaJ9eft3+uEhVno5Fljcbi07mjf84eSBzQJURZVpdY/tEyfbWBCc
xONej/ZMA+1FJa9aqfCfTgoqXWyCHHDpQXWu5BQ/OgsRBsryrrqYUZ3RF/L7sHyl
UqwvzAfj0dxHRZ9wLYATHxnY/UPK3ufoWY5QziYdAtxuvqpFM7pZt3eRW4EbCNDH
gsMndkMcwGZgS/LOFeeZCxVVbDGYyJyQiL44vyXU23bhEJtNcFITDWtnNS6xENf9
F+0Rvs2GAF45+I1xZjf15AymzT+LSe9p/OwAH/K9wPDCstiw1deYBFPouQO6RR1o
3GfEJ8jsDjmlGWk185DitwW/f7hfNRpsztS1uo0BWJctFpHIhnJT8RzxToY1Ip2e
OgEdmNHpjZLZ8Ocshi1lz/7SL0Ea3OFKEJiUYyXnK7THjQoY1HCEjQOgolhgBZ3N
+JgqSQn/njndtmQKxzGIs2NQuA9fYbeqKQ67vF6BTg2mkj5F4LhhKUEqcPCIMH1d
+xK6+jKe+0nocToVvHazcmz/qw29dXHubIaxS6BJ8JZP7XZjg7zH/SDMHla5pS/r
U8/E3uwaJnAVT6YfQJ9vByi4VD9Z7PDOYGduBHl5E6brKdt8TWphGzywfj1NqMH6
8TgodLZssgluNT57DQGjbnF2sIDddrQs0slR9GRGHTapxJ1UsoWhOcUP2j1EPYwO
2z1n0vH8Px9ESUmrqmZCbVdyUdxevbWgulD5ihiF5sq+e+jEIAAXGikST//uQdpC
2W7hAi+biCJVjy+yCPLWaVbT4AJAHWgtFC/PDs9djnf1Fh8BZ6m3q4Y56lZ68i48
M4zhmEAl2VCjnimzOUqjKC8j1OLVluxdRhB+CzPtwaQ/O4B1XDIlc31Tm3P9sQEF
k57Uf69f7C298w6kU0iNP6F1dB0/hZb5WKnrhbGPva/GpnotC5nA7X/7IeFKVxyB
B9morLrAghMdQBvirT4bK0GvqLax+FoL0NefivKsSHZxqCcBR0817yulxWlVg7XH
3xWdwC1x2nnXQ4VRQgG5F4bW2RBJhFu3t6HT+OIAQeSFKWAZLn1sAUpIlNiQ3mn0
QD0iDDyE1xDLpyppnZwJ3xdVwXOfGcqvYwYoVhvRk6uiodlVLO+IT9ucY8dAqIJq
QPQpvoCj84qSFcNPxxbRWzKQUpVEaSWqhJjXnUaPNAED8n32ASmXXc9KkD7hAUx+
/KKK7kmAv8sHQB1v60GEOJ6KJ99XVE4d5R/qiapaun0VI6oqaqz9a/qzruKfLnWU
8mu/VXj/0LaJh/K+g/F9JuT11rOJ07mYJQrdzXwpW4mBvpSME+sqwCjsdrvirSK7
HbnOutPmeClU1ltF6dZ3GqnbbvLL8OcMO6lTyeW8tfpgDdhZRLUpB1kM28n6D66x
1mEI6LDlfUHoXasXCSbTpDHkmeDRzi+XDCdkSIUAqYy948j52qKwZ5e1hzvLdND+
c+qJNM8OoS5IozXkmoAmuRwFvPpxzcZ6o3RCr3j9Es4umW/uVYweDQC/FCjTeDhk
Q+5CnZDRYdyHULZnRw/lz5pSfpvpSTsFlh5yEjeJhs2s3LQMH67X28xiBJXWUew4
z0AF3fDrB9GmranUsZhZ9s3nk1Y9+yqPv8SxIq3DmPreTnS7Ii1QAdvnlD733Gz+
SG3yV0MKpY04nWX3siKUULAM0BJ1+b0h+EkV/1BJDj/SDCidAgC8LL6xaAihOH9p
xezIFnvNA4mWNk5yWS1N0ZplFOqewi7QWSKer81Il84UYbeTBCWGdPDpK3QZ6Xxg
I0Eq7pP8n6M9aMW6pfjfIa/DOBL+WBsCkCDIkXd81MXfP7AGanc2ut9cHlB+3lBG
ZnEyL+yWuntQPotg2z/r+SSB46wVJJWEejuKnw8z/y4HTV+G+O+lZJ//1uuHN/6y
jl5/vcHseZSj/GgpACoyUv0YNHs7hefHB7Ytv//5vnMYWPkNC/62Hcl+ONG0/Kz9
hksXeMaJPeo8OC2zV9JiE07LR/fPWVBHOBKQJrF6DqA22vdlxZ2OqGG+JmKWCBSj
5S8FDg2/jykokB4iEgwTpBjt7VEKCl0kTiTKK8B1mL56OEMzi3EMTdvCRfXjY3ff
YQywul9cOKrnqlp66Ns/zh+E/BH/GVlmgo8kd50E0TyXmLNMMd3aimBCfKL/FC05
m17jGqM5kYuk8KW9vfaL1EaX6+UMfdmMjDxFCLjKZvxZjXd/g7c1dhQLmBCVQ8pG
yKBHvJ/ssmqT1gCXAMB1qVqpCdaJjBM65pZFn+Mjt6pd8klj7iuQmlGm+9UUzXve
3kQ5iP/LdUHkwEdIK0eJxKGPA7sh8aOn6GptKgR2LBUxg1B/y0s47IbE/V7iZDNV
QywwQZEFrd6DBvyi8sRjRv0aHDOI1qlzt+1dScb4hgbAwvULUYg7OS6qnT/II52Z
BKv9QscIkRCXi9LJnTdJADusce6zfm44TRmBZBDwgOJTUjm1PkTDwKIKeikm0eX4
hXlYqge06xy8mTDlobSsaYbr0y27TxGstIPOKhtqJYrFQxRYGN7vreKh8pKT4fwC
39x/xBrkcRENZvl8xZQ5pIrZlu6BQAeZyUoQNht+PjTEz49wSYVfSitlheMGLt4x
59LxFx9O2U5BfqPFwPHvjonaWQkbEXJV94BW7AmBNbyi2jH71zfiivyGM6gcwRzW
AdcJgHEMGH4DhJHNXPj+v0VTzoeFd5dRTc3x0+5lmeu0qsvisCwoH16HRhVQ4OO0
9fyrA3pMVPdhymCl34EZKUeygn12JZtC3yGBBXmvdopvdlQYD820AGAtU5Of2gE9
tvUmo3hfmmsxzmVWpzlwLAVgpO7sfDWD7mji2f0ENK1LM1lFzCzSLTOZZLczrdJg
lfn9E+DpCYVnjKV7ijwJqODXYGxng9C3cf2IXNAjL27uK5SC6ITYadzNH7kt1kpR
QPRayLiqJ9ByOS9byEiWVu1j3leynNH5hv4OBgBjZuDDMSlwrea4+KVOAyLOOh//
/fZ3hrsq+E7L0pC0qlDjvcgQ5gPGpfZyhC1pTTGn+6jrHp0rc3AT6fXOV5jwPQ/5
8r89rVEVwnMmpHZSM4JczhoQLJ/8scalTkMDZV47TCjkMHLomHV0Sdmkfvs/vM9k
r8KlBt1iDe/0HsN54qVQxV2X9SlkzzbcWv+N2rw59nZHm+dGVyGSV0U3jD/qNed8
rNMsdfO6nnuqceFgI0kZSwUpY4rcihfRSwYKd+9p0FMssHasZxMXVuhd4sIFPP8p
d6M4jH+TU71KgTG6Qv45OloRyKihkzqCSo9nDMXZF1CDJUvb+sno5D10nXiZ9+cc
ofBiqk9qjSbUBoJ014QYKx40m7BFUNc79t2ArjCNZKAlUSZ2sKpSeycLXRFgchb1
2jNEfoXwXtcUXgVxjbBlnd3LiV8JY9GACsTDYB6S8+NU3HiQHAfieK2BrIR9wCEz
k2K7twi9soYbQuaZQXzXgNa8n311i1ysTz75qJvOrb7/193Cx3sgMeYjEtb5TEiy
EHaMauX+54yva8jl+yIKMMDjjCai8Mx+S07NtIEa3GgTyZPW5FZtQXpbY6fMVK24
WBc9AhEFmGdyLSWmNo69LkGKkPiBMCiM0wE3TprTLX5DinLcuFbUfnr+bipqQlTa
BptFw89uGF1yzCIhPbNJwEGo6/b0KL142YLLIog3ghoqZgb6nXFN7oouNGHBpLZi
euEW6B40QNIcf+TbADs/sbo2j9OxX3NKI8hb+WVl9Guun+TsaA4RmF1ax95xcCx5
dRV2vencyEpjoBdHjChS5vhobnEBVU20mS+nKyXLxJ9O3lVVF9FfTiCNrSapzh4w
XoBQZULYwKfrLJ2Bv+uXVylrsIvQ51AJiDxXDw1cmu0ppMphhD/HVtYVGS8Ky58C
ZwHUUdaX3KJ1LlmzktBMWVnRNEvJykJx5me+gSJT7mXMxc8DpO6xghwkD8gSjt1c
VKgfQummZNS5xk87tjl0lkl0rAt4mZtVGgmEkG2ilegIXOuHuoDrYdT83g+KRG5v
mnwsHJ1Lp8BWKiiehQQ7/OeFR/23PrSPhvj7XVp4fW49NBseZB8RG4qVwuAHtME/
OCxbtxJgWsmwz5BdD/i5xHWycDwyqp/t1yjqphwF7twmponpMoUc4SfiwDkz1pLT
q4gFiyLilXOqHmqGZITFMM7UNoKCskonfqDLwdSLFHmDwk8aODNxAZu/mA8zYE5O
0KWKtVrjUJy47lFaRrO33QpfOJ4QnaRksTl5cZyL+bkm4cMjJcrgWyRGb7esEgtq
TfnCMucVApLZgMchBikgyL+Ld9IO7EiT3ixikej7BheCqNjqxb8jEL1Uhd1KdyIA
uNYGIejVzTbp1RbluZKPeZ80mMIJ8EgM+7HC6qqK7nofYmhaqnVaSYfkNH9t0r4i
9Okjujsq8txM/A79a3dlpakBWQmd32qsBx2J+2LU6AuK1iVr5BPJ426XmYU2H0hF
TO1oCDl8P2Rl+MuOUnRgK/i1fEjyt0prX7oT9OkLb2pyqo/ikk7ysgMq6fr9sGoV
ZKbSlTrBHprXx6guGiHQW826KxQo6Lth2jv7Ok0XU7f1vtWeZImFDnVG38mTJVY2
/qaBNjn1EJFVU6BwCy6tHJYzLuLv5H3srbu5oXfFiNDQ2vx2lPHI8V67pUPFBxC5
gZ/3bAhXshAtBTYAPBqUVJdjGWgtG8Gm+HBU+yOZDINMg/vjQ6bMuWXU7BwUfATA
AfbpH4fEaOxRLBp1Xor781hkMh3gEvI6S/Ks7p1A16hD8nWcx2YQX6QRzakeRQIn
jYcOOYGt4iBd5Qbur6PEm2+1EvHWrmqeDYZUT5E1cr1QcuB3v4ZTzURllzFy2EnA
TqcwMap0vRYQ9GeFvMYsYFxPMEd9X5jAx98XULhvKiCHiiKRL4ewjxCgTZophG+e
Ryi94Ae9FDhGHhVdXL5W/casmrewrcFgHrmeCH1HIgSPwXYEP3+c4vh6r+9NVitg
5LuDSw1t7OzY8/aF6jT32N0i+q8XJ3yX38W9aRjIfMmeZgms9+0d1k3B24XaN5XQ
+ZZrtvu39fSqGBpLErSKT29/YutJvmt8Lvp77vWdZy347vit4jiYlhh3o10LR2Ca
yoD3ioz9L846qPPNJC0Y7TEg5TBsBxwrCa16/+e0OEuQYMnpdmS+wPE7ezF1Z9sM
KV+G2Vvx68iHFiIdze6XAzt9TU+eK/N2A+nkgeRN3J2pFarahqx7943nsimAG73S
MXa4nc1EcxLz/20VIpCT+1np9eIy+XlFqor6X9xs1FsDvaLk/ndrv+XbCWvMKPq3
2GpzXXr7UL3wvvZj2mMNyNOx1LX49MEjhhl1EKaRxk71l/r9eiA8jVgbSNHL3Aj2
io19YT0eaNzE7/hLbT5rcfhgOP7d5dSXeq4urZbQi7moDy7/A0bRbC+1Lm9vuSSs
mGI8owXlXfo8cfc9P5ogb6LeO4CJRTCyKAzqgbda9sssEDXQBxR64wtu+nWjwe2D
/IRhandWO8/EbLmDoauG9pxq6ArSFX0Fye80E817uKf0i6SZKotmJhR5RHvOUZKi
0daeWtyVd6D47Tj5P9sV3KFpXOiqGI9h3ChcHrjbeUUBA+7hfnlzS1HmZ2poqoze
WWykLxGjp/I2hsQquEjTzxB4FTOmCytps2BAoCFPC3sS4VyX2utsPbbNcYeoMcye
7myJeRefHTVb7wzEuFjnsBEfEpYJ8Ejgm01mXOoRbZ+jnBaCenOyQIg1uLgMzIbE
4z7qi+YvD1LFKjD1ao3Ti+wp3+AQ65zmLCchutyH92ePXHPnXM1GUEY6p6uDgENQ
jGcw0tRp+2QL9fYFd6erTmEBTYE+t68aok+0KGJq+KzP42dtcIIKlepcx56NKBgm
5PHUaS2lXm6M+FM741F0L0VPTV+EsXW7iXAcP7RWWeagZEQW/Yox/wkxrAS0i0UF
ZMAzkn/8sYv78Sy6LC7QLgYw5TyxH6mCQP5E4DISBgS0nREcjvZu3Zl9xUsQ4vtc
+Y79eXOKR8X+A1d3p0fydiI5XEskQAOLx4tGk2iX8Qy0eq7Wj2YFJIYMSbiCYVsB
HZHhgc2euTdc1svjAj9EQRiEi5BRovnDtt+/LFNJ4Uf6ki0JZoW6E5iGVw/gYqfy
QqXMq30xZ9W/taq88bVkiETATmpFfzGN4gsYYHD+4GoPQfKlHN2Q3jLKeERuMCl+
/z45gWVel/t8c1HNnlYHWakVIHrBAstqhvYEI0scRrP6mPdqS0agxayXbCH7YLdE
2JQkrfnviicf1IRtXZ0c4Dl/KLAhGR0a0wUMV+ejTjtEjrXbnh0BGe2EfDuXFNVk
BNQPPb8UDAf8LWwnievGttNoWRWorDO6ffpcRnCgRMoqBOjAm2ijiFE0PLu7B73E
aRLpCvDJe7wxwlQhNDVMsOSejP7TvWGOv2xC8CBx1e0d5UiMFGIOu18z9WRWc7Z+
73E/0/Df0hlndMvDtMY8gzmHBhaKvjXiSpeKQ4YstJ6P+C1D/eA2IoBGHc1pku5q
DY8GUeY2Ba86BOUtS1H8N3t7CCcdact3wY4uVYeSLHUc7gcMOdMu5mHot+G/GVo0
psjmr2muoNSyYt83p7o2EGSelCTyiOvKl6VEtwW1PcZhZ8D9cNhFW4q4gPYcfDfV
MFLpLyLfzIlSEmPmpefJVn98nTqJDDWnXksq4m6+t+ivD6JuFGPILy/ZYzbdeBoe
wRuwGMeuwFUhiSf0pyCjiQzihw5VgPrnhxvL6tkJvgb4IHkZfIQb2u702Sc0ty5j
QX7b/VHvRCyR/Lf5oFz3YEoV4Dj9mtGkdMfWHCuaxb/ZllZ2psWIMGMOE50Pz0H6
eCn/DWsZW7SOonx2MVHG8i0KfbakD3ENznDTmceDbzuOk0WwKDBdPOaM+11w41Mi
cD42/j4fyn5ZKZl9MTRFpM2rzMrBQIrL3t/hGQuG1E8KJqzlEvt1SU0HLvtVln+I
gCa+MpT4QTjAbJYldm1eC86ZAF/G3wlLKpNzbYtxem/5i1LoERqENelDYrYpAvLm
VX8B0wUaIiRRCl9nC8SeUYJpcX+Bu5zw5oU0pKyr0eTL4YyF4/g2yURiceh4mkAR
iHPrdPRsSe3jGLAcNdO0nyvCvoXwdCsQpzA7jk31d6iY00qNuqbRT9DPWRpLOuY4
/tSgbKNoaiEsf1tvWDKKkSXmAc2ujjMYyBr5qPjJwk+0RikFDRUhtGC+fvvyGtnL
P1WerBO93NXIzWwxc3EMaL9CVYG/ouSGdD5ERyaE+5DpFsoq5dsDHsLezPvxCDS5
DDfMff58GmEVUBHf535P/OPRfnsBudGoCn1+dLs97+OkKRdIoyh1TSN2QMeEZhkT
ByJnk3Xs0SYMO9KgLGIMB6QxaUI6mw3+Nw4CSt2Jhh61OiydkIq59obSusNrmpdY
9cd1HBq9egNR9xQfBPFzHKD4WMgB/ScwevBX6Z3QH8HqaV1tvao1a5BZOywsbHzE
GJyuQlfIQk1q2SPi8QqbT3hVi+iZkiAF/7KIVA/a+pY75gOY2kvA6Ran9GeEoBdg
M3Q8Pk4LgaI6w5//TIwBiHuC+n0S+A9hNPlPKE9qeNc31T0kqDjOAGWZfOopnpjk
WY6y3KbP/yAU8rEF965C2+YoZrv5BRbeIBcWgFPPX0ScKB7kQjtNyHkEmLwmQ5Z3
k17Bew5bV9OZqJ3P8aEy+TmLU6h4RQnVnId2xhmcG5LRuIozud4itTWPHxTj0p5O
Lh7Y6XJTABrTJREllhkQYRVjeNvkbEZU8nYnIGlPSKzvsba3NLCoYSxMw49Qn3C6
wlO0XdR/liZrp9qx7gwqwXDOo6zmjr4h3gwDDJe+G8zXo6P8QLTxejfSBOsZOI65
k9YmLuqkoYtWUFIJ/0P/HypV5jRVuRLRjqGu4DYIC1//IDEhXte7EAGDqbPajJX8
VQSULQr3US/i6yPv3OTgJ9MHFxidg2DDX0a0lb3nnuucGK1aTvKe6WaR4tHBcHx0
Qmk9tEPEBdeoCTEF323fkIM7LgcU1MWLuzocwESMIm63MiDtasI1fB6up01mbVW8
bDDlcZKL2Q4kLJLVFhtNFK+FSbx0vV8jkacOeJ/ud1Xnsc56By2Kjzeca24RnXQV
Y9BRKHqvpOFnR5+ZOdIY3AlbN/HgZo7Iv7vvK4oaiOqd7YcL+TM3lNuhWswYjN+e
DxWFgWBRKoQYiPB2FzSPmiA3ob3PiQjcyw0G4TLFLl7JkSWkDS6G2DtMyReDcN+N
xogwY5K0taOn6/a+knf1OPzs78sd5Mdp7OF07afQaNDgp1GC8oev3yk6gglMc/PN
mg6YaN8+qjwAqzKrpTetgqAgb+0yLHA5HvxBwLSDXyNRgAJ87eXfgT3z9eBVaT49
jEXiuQswo0SE/T+tbUNYqrF3E5V+nqJjno82mgG51o3QTE0DjDDSQ23krTACb+VD
y9b+O2gq3lJPm1kUxy14lVHDILO8ESkrMHHc9CLiyCqUZ1RgmXdATLV/ZLmFnCyf
2ivnFCVZsjDVO0Yp2U4/aag7QztcqfFCd33tCTimArMs2gDU2TWs0/w2joYX28pE
z53y1wraDK0LmJswaZplQ4m5wvbfiNMHRpmlwUHZVanU9O+3TZ6RgBA9n1D6MQwz
iqPPy5bLeuLLh/56sh/mCiHSgGZBFEorn59XjYmdltiA9tpmrdPsNf3cVxHEtM9W
8WVDXZVGAGUaNtJZesi3C7t8ka60GF8i8Pcf3RncZYiDCga4xd18eJ7hTsvSbiWO
fQlcpSbxw+L60JbDP4d3VbecfCUq2Vcuo4XLPhwra+nu0q6l8aQ6ntN2u/Ivt+WF
8tgsTb0Md6Thc3YEC7fs8sejWAP2MnxmaIIgXiNKhSjvpQOBHG1Yr7yQ1tDyU3jI
0HQys1nZzzBFVNCDBilA6uZYnFpFRiYpskmW03Oakwfgx8YY64tkdmzuB1c2++7s
Bp+1b14JOtPRxmD4J4icM+zhfNXnNaVLW5v2Ko4EaBLsEKs/HvMLXGF4+pQaqIE1
zDY63BNKm+0uVCd9cs4PfGLsjQ3isVJcpiDDRIDCCbFGzAlsxnjt4TQbA+EcmKyg
X8tlr8aXllD2zWiKR71odnbtAhXr6nGDd/eKN3ajQXIylqFI9kbXLCYceWFA9gmt
G2R9Q/7npu1WZQac+r1rPKKmXLpHxwA5y0bnMk37iBHT+2IgeTDr7RyqcHhoIUqI
YLBXH1HWOlADuNwQ022t0Gh6dwoPHcar5G1S5I9rLK+Ra2oi90YJM69RV5ivSRZc
Td6OGSFMdnrGKywnRqygFdBcD7C4Mag3HyBDoK3MiIL9AP2zlOsI21xzEm3KXadT
X0x1ibPEhiRE/e5KE2/9BspPRzM+0DYx2ldNylo41q2YTgE6vZQLH89FVXIb5cSA
VZfgjAdl9747cD7escfQPzesxt5bLAkbqyWMY9+gr4m/qHdkCFVAtQb/0t7421xY
DXa9tOh6OlI+D7dop2tucw9QYjmdWkz9ARRDc4tXZ4nYIxvfaPYYEnHH6lLV9Dx1
8IxA+Mij0w17Jrfj8kq3G90TwvLvd3nF4nS0KhAX2r7gbGcqrgepe96Z4rvauBUo
EvWl5Q7h3oFvStjAod9LejIkYIZI7TVoalTzIXGfuTWvpc66zPw7TyfdGdw7ROIp
L4IxZH9Jgoy/xj3Wqv/VwbHaxOKBGM+hYNjr1jPec91kxnGGTVnjAWGQNa2Aghkw
T04ExGfkyaZb5CT4SSE5N86swtOkTM6tbaMpuh+A7m6jpJ6SZ2rD34tu8oyCd0Aj
5yrIfilPrGMhAP75fvgUwiwCw0prfwCtfN8UPM1JreVb06bzv8iyWcXIB3HNThuN
Pk6cF2yfCj/4u6TDQumZ2brgwAmpM15wFTxE/GawV5yvwXcQXERAS+c1kzqGQ1NQ
g8Z3AiiR3x/w64rXcv0mltgjb65sxCdoLAdWwr0a/OaV4uulekUpOL70Z1FsdRbA
I9phY6D5vrol10KIjvG1HBG7hUfwJ0JXbCW/P98DwMyepFCBNG/h2vRHIEji1dEi
DmIzs9PSJ9W/QXHQaMRDxH4ri1LBy9L4o4yTDv0ZHP/NA5UnQpsX2uHaAXhGAtII
qxTPr/xRtq0myxBoAZPHQVDdBO6eGPpv41OHM1LSSVZg50C7g2ogqcjS44/DYu0i
f/0+dwzoIihBzaLYQw9vqos+FysKRvNFeKK8NbZiB+5pD3DpZn6bjYLNn6CjpxPX
2QL/UJO/wko5QQcC/U8Rz7OgYyPjPRtMuN2zykI3weLLfTfw6L0VjdpNKb9SlIfh
2JpFvqyMW/8ei29TUrKZv/tEAA+mhBsQrKJ6SZC5zO19bN76UuEXjw9cr3WLqCSJ
W/sk6JVFLL63LzU8sJD7FWwTfpLZIGcDbAZXcufTDKJbzTZUCLJHvUbTy/iJKBPx
FLWQEpuyrygIN+I5Rm/TaVuUt0+gfq/LOKM3op8iIj9/BCpxqwPuSfPpEkapF+08
Uck9Ui7mlzIjYwcBVi7uTwdxafpzFyChdSjVA6Yvq6C2E6X4NateTnADwixtB1vp
ucmMg+5KaovxRCgkABtO5n2gX+RvAjFrhXVTe/6Dm6yl5zm62r1kL+MhNZ6oLMJ4
t9lO5ARYTXNNsWtPt0WMkwrh+VUtQY8bTwDxs0n26MB0XvW7uMCn8WAH0UBPG9Zg
rD9VJ+rsf9H1BXwpWn2oQAOiI6yhDK86g8/bMRKmElVZFTtPHnIoGcN/kvh/N1kP
0g/opPBWtAu3YHXr1GD4CF3QjePJVmWW+MOH/a6R/KxoMGKCNuuPdgLXtk3cWc32
vLXR5C6hQoq3Tde7DrLueHMRBu/cGkIxIxc27eequckYqvJCwDGY4NUzwcTIUvWh
v7WxQV8nV4ysh5V7ykpzhbTtyIzkLog1LMMCJ0O/IPUSS50glaPk8hqVL00d/DEF
Ls6Pwzz2ljBTD2dVR6Xi3Dg2i+Xc5yUa28yTqSW9anTfn92QDb/ldDT9Fs6wn/e2
Sj3YY9qX4S4iVfZjbiZCdr81dW2lCZP0UwSL61Uv7wDpC3/TclsTW6gs9wnUUJ1i
tPYyFt5ac6LN7Dc03XFE5l26W5CWBqXwo5LSt51wmbiLRn8IwNBGiex1Bv68xAw0
aXRwz4Fvwsjr+vAHyfsr4WdleeeCdhS+w9M/W20PLeftzg0KwJoCj6Rb7hlpxPIR
zE5Y4v0rQwhAVIg6IsZbObXJzNviPagfFdX1ru6kxoMBvaW47SOte4GmhC3AIhaz
UOK7HeRdNJEKYjGyTrj5jSkI6tCSCWOHA6FRAHpYVTZPIgW+/qjz8l9S/snZ4hb1
22CI/XllHvsNDkekb8VzIQ46VBZpqYgci/6zso1N13lrExmv1lUBXuODwWEkfG2P
PPYGZ1UBxkTYIyLJZtzEjCszCTIM2Oo0b5oqRuAS50QIH4lMqrr149cuLHX5uyhr
4iWmk02FZBSAyhKJE3BfNwu7ZNc6/kMSfIXQQ4MZb/2NEioDTXnrNiPg02cOKscV
yu5sJOMDU3VOnu4y5dxHO6lSJWRYTmlFaw+K1JXDsIgG52X/XXDs2XrP1KiqmMwZ
8HuyF2zAeXsAvMXwjt/xCgRZPdQrIryi3oP9heZP43bX/CLlG1VHNkEBg4H2Q82M
uMrEJXE5rrr5mifn75TiYLEb60M/w0uaWzcQ7pmn4OsHU1EO5QO6rXYHs5bEzIpD
WlA8oV27U0Rh4iHc5nYtXPLn6I29jrOvuq55IO4Dts9Su7TBPwQAzujhEd/6sSe7
+r9IPYXFkgU8RtZCnB0RvEzcVpsGWQZtvD90nxxeuUpF2IcYOVxkogcpvjqqY9y4
cYWX8oJDxH+nc/xGEBSsKQKoilEWx5Tks4z44Ozs0Lf78nh0q/NVHrdgouyWLMa+
TesagCwVCCSAQ5PJYyKtczNJdjQlYbrQH0XohCz7XAh1CJnjAwBkEAqN6eqDY4WI
6CQNH/fJuiXseLcg52aoddSdrsjI5lwr4Z549USNEqH62elnHO5I9wQxt+ahQmIE
TxMFADzH93oB9zfzT7q+IL7NSsHn79HEVADpLRhNAvI6wQH8/3IVvvJfC3jTZFkt
9TGGI414U/NtO4RqVFcE7uCx3ho9XsFio/UvGHcB+ZVHlV+vPUprKWDvUG7YwVdI
SQQl/47YLKLDiNhiegj6o0pLMAvTTuoL3fwaYkdg1IjcDM8C3zgEVh1Oea0nJaJY
FtCXdQ/javGAfyTpY+k3uW0x0plPTsSCbKqm/VZJGUKpxZAHZQNK9XbsMsZXoCMz
9kHspf9eLIEFPGHzruhwPLe9BDPcxk2a9ZwiK35HxemFr26HNYp4DUPkYjbPjWcv
HcaHLs07gh9CeyY1pLYDlJeaG/ldGQCtGiZuZktIKkBLlJoSd39aZgocDoXnEs1f
8Ti62FSnEDpzQPoEofnc1LV/CI89v2A3Szc1ytY5ycabI+fyb+lGJ5iKy3DsU8Mt
b7JNOizVZiyptEYwKz+lZgICuoGziiEyUNp4OkKh1TmN2CYH7VadUCnjJyg9YzHv
y5dtK8ndVXngeSKiMWd3IPK6BgzOW1lwHV8qIRfD9dYBvzp4wmHeExT3d0vx5m/l
qg0pI42br15r5wAO8I/9VGstU6dEg1w+Ft4JSnWEleKPROBFu8j8DCM47R+k8MTG
+CyieXUBkv107ZhmB/ovQ8BSMwg1DMHGpatG29+IN31l0QNXg/Kji6yqjVhgz40V
mT+Nq/c7QX+C0oF1ozrrAdxxPTx/ru5OrUtYU2sq1TOLhUqwOvyXy0vAWyK45hHX
ve/sOsKwiW7gRanOJssQhFTH+nMcseqNClSn1MBCJ+A5zG9dQhvPQwGF+UqPBMBj
MSEFI8w0v/iTWz5Tfgb51vFt2jLqDCB0A4z1cmxVitiLSWA2BGDnMj9d0kdrRoIs
b9DWYqp6oueDfUvq1RzW9oQpr81PfNzqnBcRg5kR7+5/dXMdJyTYP1YUcaB5bDFH
/48k8sVy5JuzvhEwiNn9TIy+X86SfjbdcHceR0QuL5GrK3L9iun9RdErJ52WIYtC
penqJgU9NiUDQihKKVgQvjdMfshlq7qy2F2tu2Pf9LoHvo0UQiUfvTqAl8O7KT6N
N93aXe8XMhbSH9yZh39hnS2sK7gX5qxmqLul+HjziR7ZnYcKTIj89PYyBsq592cr
hTrMX2GBlt1K+0S52HWXdi4Oj+mHK5dTgFEu8zIug9asLl5JcWnqVYD1Hh+6VqbY
jdZRgUhK/+4Ts+ZZqDFUFreusd+P13jaP280hwUBhnl8GNGWgNcpBScHyNSLHXJC
eNvZ6FGB7AmiTvH+jFue0cF413JGe9XQgwGw9ctalphv9uACvAcUblAPdiSyoCl2
aLId+kb7hYZTvrDUI+JGWp6bQp+aoylwOKm0gUozv3GmNqBEZOlF4nIeHaUb3egx
FYLXYrsiYjXAzCVhOr1wL6Wu6sqSie83uxJQ+s9seIple85pUYwhn7yWqru/4dXW
7+ZS96oOIcoLTIO0ob2nEa/NEEdU38zaJ9PzfnNY3w3IKYncdhSRQvfAzMCTwPEd
IMcu2gp0qYkLWnwEu0UeOaB32FckMXs7ziK79868Ki4maFeowHdxFjiaHGK6vkb3
2QuT2D1zqCXCDxyRvRu2cfsKHq/K2+pqPIozqOMLC3Mk5YP3EbXCe38fCmh4DdWC
uk06RKwie9nYxH3AZ/xaPWzbdiE6eURXV7uBqpgLZoBZSMfQDkor51RUYeVA9/eJ
4uRcVtFKao3WGNqFQ3pedTFrhks1b/PpWbRcZwDsYss2Mcd5BYAxrh/iZ7TWQH94
yXzvrfDs9S1ESc3G32KKzxvDvupI+vaMo9UHG3znbMDs3rXY/5+UqgLV/rZvpL0B
o9rlMmT6zfnsULNhqdOrQ1WZBMmkz4swVbao7z7X87GafsHH7i7xuu/S+dkqkhED
0usQWrYQ3g45tUIl2Zlgg6KF60Bi1JWiPMsWSeLm7tvZx2izWePoBRyV5pUEXJ/q
q3UvPNQJRZi6rtC0DQ1EzKjQ8dWvarPz0i0Q2eWh4sX6dxZuxQkzXF2RRjcI9y7Q
w/PELqavmZBIpb8CzwihRyBQZ3u1Tee0li0f2eu1sgMpYmwH/S5k06DiZ34fIIro
aIb/K3PjAVTSO1r6Hixx1mqyOcMo6qa+z+BeM/lYRQMqWVJEgp/M/x80NEQBRxw9
+CET+RH/F+sVcVEWj52quEdTHczYoB2IBLH32SvP//5E77Z+ybMBaBuegVXxTj/7
eCyuzCxPuNb8iKiSICLRXCHoi0fVbI7JCh8XpvVT+LDjtXqw47jwqdMe5QoMxtWr
K8L16fU4KwAAkjVtfektWlVEWMt/FPX3hbpAoUFTQsF403dL1QMRnz5nTMiAjc64
nd0U3z56SHTqjEXpBkd680DtXBUArg1D5sW2x+5HCn1rgO87X+tRcu5XQg0AIG70
m3OotXGMhSx5jgjyvfWnN1I7Zijrvo2rgvF4AJqwL0LpccEtsIv2NmFmcbRxhNol
6H89QZm/IH2imJWgIOklTqc7Z2Gu99+FRxD5TVOd/4HWwNRkExEM6ifc/MAMb457
d6J9ovqgadzqBJwyWczSn86QMoRONOsW7a8cMOfWTTM41/TGLNy/dCO9/jd7Wnnd
Mksc7T6Rko30S9hedSpIxWwSkSCSxXOJUfA9YXZoRhFsjE8gVOc3GhZRVvoFCi+A
bhS6uEQQWP+ersfX2xSBKrkIPRZIrzOc8gdbA9YNUE+uHVk0L6f1K4ioczYg13qm
0H0+8lN6pC3rJBb3WJR8DfZu1yFoAV8VQI12HvYDr6uvijzP2xfXlJYxJQLuPTJk
qqPGeugg3fbp7JTAfE7y4SY518WvL3zlsJoExrob34hz9TrqH/QxXoWT8gD4vysT
bujgr44XgYiCcQvaFUwvpQjKdOPhgGRq7F3M1Dekuy7p8vpWait34Dp9Rum6M+ku
ZP3F30/McN9NPhi/fRzqCeqQVNgssE8nwq4zlzfG0du6+mhPjjasrpo5CeAdSdXv
VkiAAr05kwJD7vhG79oz9t0knWFUdZnkJruQ0TL5LGTOu9RwYKSabyqnHqt5U+dS
PERxDU5fq1CwauW1zaIuHpBQYoO3iXo0z/7bRVJQ+w5oDgRfhWhZvCH74o7BesNP
Jz7UBnY6jfS+RBVNlqGNvdYpb/au0VB5HYxUH0pPsl3I9nDWdzgkaZKTCMBLBM9N
yZkzwLY5DQqsbK9lVKBR1/ZVV5iCVMlsAuIspBK3tdlW2zLZosMJOKsuH2I4dd7/
JdujRLEobNtTqDju/AonN32D1JTnSgbPuvXC5j2Q9uCYzOE7j32qmHX1edXWGtYr
E/8ker/slplfg+cwYeYLFJz/35+weyu3tFyqCuBMpI1t+bznXGWE3nItDBVT/9+/
I/8mqjMCBu5jNNwAEhCgsT7LL2mGuStJLqPmduNrgThOGNrYvYI/XMB5wHjpaLb7
XUUX04FjWIYdGZlFSZMrhRiU9v5Ejxpptsb+IoK74uKPvBGbMQEOpDxGGzCMAUlv
J3FsNJmSaL3AdR9abjYdAQ3oHPoZRb/1lnRScn1oXI5Wi/LIeTNjgTS/GRt8c7uF
i6OLQOonrBfrYIFOF536Nfv6EMPHTqES8/Y/FMXGoNrfgLU90VzQVKDnyNhh0bU+
UCqE1tJK/hIpmriLGZusYxrTMC4ZDYZV1CqEeCDf24vzUVCYmOS0meq+jkU/Xknx
yGn0suUL6kp3hvwvk5sb1VpXkpC96Bv3RFgG6+GOxbX9hCCcbu+94VQg0i9vJ463
7FLPyMDK4uUZoIqwdH37U6+cf2ekvUimcxwCqdUSppa90PzTWPIebHOGkzN2SyGd
2PkGXEFxEsDqlUy5A2htHT3/V4Jg6QsbXjULYwhPTQrxUhwEFuLDAYbln9OeksaV
z6L5tHPVRySHcWzeRA8gaEM+u6nGziTildFxLl7YZu7zyFDgMzwWT6JWmknxK2Vt
8k6ZUMjhpju6JqyobuJTTETjbxTgko+hwzjeAguAVqtT9IUOmZ/5hmzmKlbNXGUK
FQzx1LBmiiVvGk4B/QMaHdsl2XMaFCvTzYL6Chrv0LOxCWPNv1iyWbUrToXXjYow
pNBrFs3THwhxVkvG5b1h91EIvz0UdGU64VRC6aP6pWLqZpAeB/gRgKZ2Oum1hiDW
bDLrA2bXSKkmiYPNBMusFKZqlfDKZC5HJtHBwcURa9Dopv6Pw+vx9IMgN+e7Zo34
EEh8We3H0B82Gepqoxai/aEUzn5PK/VRCTts5DbctXi8oUzYhlv7ueGAa4UgW1QE
Bo8NKIXbbAeEYAQmZ1VJwKWWgSD1NpcKaCHbXyvM5eTV4pM9VxCLW0UCvDP4RaH3
7LqLmxJJXyd4PQYo5ORGixQbz7scK6f2rL1/DQfxr+I/vpYvFLtAoS3EkfKGK4JW
kn+dx6/dCMoCGUXQQQ7Ithmb9+Ggl+OyTzSxsh6/WQcRjKFWnXNU1PBOjvrB3nGm
A7SLFTcCE0NM8kJtwIaSWmubSFi4HPOJ9ofEyZ3Z31Ql/o+khIxX0vUt8Ojb7FxK
mw/JNrhbx29yG0DvSS5U9fDGHqzPa3OS2ztp7NrYuSyGDJBZYiv7cd9y1fVIVDDi
h4EdQRU3+yGKqonicZqKwdlkVxz4W/Y8yfGXbCO0y0wkSkpvnCapf1/h4BsUqYwZ
iFTKlxZuxXn0aJQRSZC1VcjkNBLX8ql/7/lZpiEUsuZJHF0VljI5d0sNzc0Elay2
pvjuA1ABRG9HAL5DU16/ea9CKZMkdPXdID7eZfu9DWHdgBSy+ORgRaZRW1BLizUB
GZAljDGq0H+26SFxxmxIPSipPoD4H3yo23f9MpJwFnjAV1nTOjV66Tjgr6IAILWc
oOYDw3tBZBFW6ohuaN/uGKss8KTSGpS/ITsuWnor32NfV0nf7WgJ/I60RBnJvnjU
/2vieOGMHLdGHk3qVSJvCuKn1lsO/Wi/s7H3py2UrTdhjJG9vZX6D6PPwzYs8R+o
2Hs6abteIzg5Cw/Jd/j+NuPZstyoyX4c1bftzbE5Ahzznejw+4kihRRquK1HHAhA
eCx3cpP6XFkseTscBFW0pBboQq1BOYLNetKZY+UqJ3+a/R1ZhkHkx3kkD3+8z0L8
xX/JO0Oj4I02LcQ/CPCvphALeJts723IpSLfhIRIFv9NDmUPchpXMTWMt4xAgiXr
wnZyehyoluyoGvOzbsOD24qE09y05sNQBNj+NtKy1962OLfoxxwFb2OMahtDXml3
BsuAahjgX/GeMsJVA6S8YFbHc8qMo+sLlNKrmvS0eZl5lqu90Tlk+rVkyrcY1+cy
pPkAKfJxpM4sZmg7txggzmfUQOUCIdT8DgsPxsDY4qVekwT/VuVysdmdFi30kcRl
g3tapwxuleOYGo8GWdZeBDgL/6rZtPFHluQ6wV5UoLbm450xuutUC3mBJAJ7yse4
iHWI+IAqDa6CPk/GSKEixk4mbEq1V/wGcca9I1eh6XCq4yQ0KUcfUQnEOIVqA7mF
Rl+rVjQSafBSF8v3SATchFlVxDyzrTSb37WCI53ZhT1sW9vysIHcIFb/f0X5tP6y
wGf+4KMSMrS2gKiq2ID3BOVhYFq4YvIRd1bWpaxQ4VIwWHpkVZPaTaeqarPTq+ir
oFCSnqc1IQFUNQf3ItMfcb64M/AOBuRDDxmbq5y8ZhgYNYW/8r3Ur90BOWVkRBQ9
4TDwUP6g/IWPhF7zFU+EgNzXq5hTcd0o7+3mNxe94lNgZ5v2iie/bTeflC2En8n6
mMqYGMBJXA+c5DJ34jMK/Od0CEn9SNcN2nw5MV079kzd8VHEVoGnnPOGe+/Bfd9o
fYGNxmpv9w+qY/tzZnJTMP2vnW3dWbPC8nnfxe1QQo9INNl8dwNgaXj+iRITPEfA
pZ0mjECl6Py1ZEIXvwVtVNXpWyNpbwNFxcz19LYb7pMAZ+kR5RoibRvDeDeZYMbi
UTPaBLn+1S5X70furnfaVHKznno1uj+gaPip3tgvL+OKofWtzriyEMjOd1RA3pMp
oI0hUDftBvMaPnkMzf4kiAw+eD2G9kk7/rNrkOCLPxYxQW0CduGc8VAcAH20LWez
2oVbmx+jdGmzWr1NcJl/6LfMwwd1Fz+ectLDA3Ehh7hrjJ59sFhBrhMDirEunrFS
G15vhZUl2zAptgIXlpu75DwA9loPAWRKD7Q9fp8Btq3zTonmI/u4YU940NBk1RkX
hk+x2i9uOFepQAMuyDssjLrFo40mwm5dzw/eOtimx18Gv4TwuCXYQmX8hUXDIzw+
haZ/sx01LXsAby617t4SXokLOkLZSWnvaOOpQ8TTwgGEmmGPEPYU71GLep5Ya20h
cCcUvBbGsMYvvzcGV6RF6olMpf2MxuIlpfvmr++wfBEc8UUAlMWI99lUKk42M83j
AMbngpPH4x8c2HKeEEyko2R/F9uHaZW+VKjaLrvPmNp4Uy6TXYDI2K4lLAs4+bYR
Ul8UNzDF+rgH/mzKdkJb+flWie95OfN+2/ksNKLTb3ioRVEONGUCaltUHkTAnaPf
ezuPFdG9Xliuou80XjXLOX0bd+qvEOvmsWhXL61qj2yNEe+M0oQnigKNvp/knLYm
txdm+KVy74cqwRRjpZ7WYKDsLepgQsOzB+xx2AsVQDE+fCPOLbl4Wxw6Qjq12bMg
AndYtjYX7vFxlVtjJ3iBXw9x9vAaX9hdJthBm5Be/aMkfWSr8i3rhUMIc+USl3m+
M9O69P4PDDhcoTETZ09UYw10lNHGrzOLzymTnVyUbvRWOXkPs4PZweXmqclFCuzf
QQvq4cfEIbtw3K7YLFOe6L7Kug0U5y40i0DR7APgtwai7MIBBGIKMUWXyDj7aILK
LcpTYMRrmqcl6SZR3fvuSIc2spKOYi0irnCbyUnGuhNXWYrl7vrhEMOlsOmv6wOZ
IP+thuIq7iJUWIsmPIM92asb0xvpoozNhDzUc98MwJbRa3j4eVzMkbFulEaFXi1v
XBkMxLE0JxBi/I+EFfDwIU0nwH0B77T1bf02JEyfLotLrJcNvkYWlPGztqC/oEyN
1KWPiI8gpGkwM6kTdQUSuSp1popWDCbuJ+cKjnQo3IycjBpYGSecN0CxdnNQg+ri
O7YV/T6VQW6ZjqBN/BNWuobQIY3jPIcK5B3MliZEET9FdmOFyKtyU7GkN0sBvtcz
sRG7kvylzQCyZNqa1iZnOaijPVhxLhFO7WStNtPvfN2pemHqjoqidnMTXHPQN1Y0
JSYBCUqdlOTKcrXUT3S5nEJRHVFcnM7HTagmFBIFNjCy4URrn4/+3r1T5Lg0wjtg
1VPR4SRzsx/tYqg88jHkYZz++SaPhgEpAhzd0JNOb/GCrKY1CiRMu4SugHlXTjZm
Pm7YZsEcAbgPH8ljK6YQFdbkZ4LbDEej7gjES9spjW3Ud8tzJN2lFf8NdGZ9+6M6
SFj5IQtNe8wyDdVmErnjTf+i5GKXGH2zy67aI2qriUVEgTSYQcNyoTfM4U/B63O0
jutM15TWfPCzHJNro2lLKcbFu3CwIz6v4u1Aq45hlVLndGt9K2kLBbs5mNrB/ymw
ErDoDejT6Bhs7KyoxSy6Bg3WY1KUX51SjBFiQvvW0sKEhINbwmvV2MOccK8JkJ16
a4/A2jSu7xURQNzL9wISeJtjYTXOa5R31drddN0YyM9cDjBg8mhCycQoWRIZO90B
vIj340Azp8ANS+JR+KxB+0VF+ayK6tz2V0l4JYg853fuzI4AtIfIaKLEM9rEAkpO
3Xo3WkI8tSSvRBfVzjN/tGfpgkXyz5w5SueOe9h7wE23NvGKHMqhwX7ScoUGWWEU
2C3pqRKpXHm0xII/eRUaN8aZEtBZeDFQcOAUK6al9bC5iUbkK0vB3hgf+NBy9PXN
PfbAQuK3K+eRFR/dLgC9eyNYUPOeWN2outtZxpgWLF5FZGF1HeYXtQJV/I6qsqPa
esmpQq3QoLKEU9Y5Hgqvk6o7FDICcV4cr/BPfSXWG2WztKBfV6cG8yBCQVE0BhqT
PV2DHRPBLc/5gYlGDjZ+3mn4qHJb7qnPMyaT3guoiZsOC4qvMYIpPadzgKovcfqw
YyYFJ2jCZoXnyn4tzfjELTmiJge4lout14Hub3M4ySpHZgHnLNeHOOIJp0XCe/d3
R4ydGyA204DrW4PGl+RcxmuBBhRlCn7Mfmo9uHaFW+XWinjLCUCNwhcIcDQJw+sZ
2j0yVDSgwqHX9l3uFEOQv5yz4YxLGr2nna8NCHaqKhVNxBqRKfP4uDC8Qd26Ob52
dlYpGZF+UXbwK0oQPaDB17Mj03mpTuhDkRAAw14gfgKRbqKPNjos7VTa1GQxO9mI
qj0e/X+x+BkjJwq/5Q1USxx6ZhvHGFuDSYmLVAn8ioQ/sgUgRrrGYoVSM8A+nFyY
ElSzwWgsQ9+5NQ4MEhY+/u5W/rfiruDssGXYO6PpTjJI6GJMsoKnIXtNTToiVgaD
HnNCK4DDG45hZ++j8ocULKyVqqUxEU7F69KPGlWokpvZokPGsdary8zhNlVWCkX9
jczviqiTpbCOL8ogaNa2J3UuLGdzUUPK+TlJPOsw+XN6nP4m2YTIHo2i9Rzr8Olz
FcuyuO2SkRVzYxI62te0Y85R0Rn8rqRm7qoOkWwpn0dO6VaKzGiz98fFhBiBR7Kz
MPI9RVH2ncsg6TF/HW48W5HAylox1zMsE1GTDFmqtesDT8nhi6nKbNYtb20rMWU5
mvxqCmelYivnhgIMnWMCn8QnvIDDG8X8HhU1KESZFSm/cXVkRNE9c0JpUDgRlQOg
MWgzkJEJf4DUaD2HX2PjtnSEZcteqWQQ77k4R+4YL/+55Qw32T46RXjDj1BEnYOc
gGByNs7bXM5jLMlfcePC0strkL8tRMMLcG6FHawWPPZCEcnbw5VIYCWiAXoQlOqY
ceIIr6wywAJdgSoXdt1NB37u1XbXpuIogD9LRpWi4JzqLc3pN60P+lS+mrJlxsgk
EwZHvUyyPR+SR+sBlYODomSC3vMQ/mSuIcRfwe0ynZftyfeyLwQuL0N9/wvJfD7f
TkdSCdQMAb78VQJAyvdbcBtcEGYFfX7PV/b9xJR/+42LHhxhuoIFBd1z9Gfk11aD
HLJGZIZzTmsKEuQOnXR0Ab712zBQLdb6ygdICGS0N5iFRWKl1bcd7nD6ul3Zp+qa
+wsph4lo/OsgfBU3aH5XXypi3H2BtuvtGhaSdXm1e3L9ctJ+ESFLG5mOJUTSiSQL
R//oth1UgTcHdTVz5BUWZnIIZVAHg2aCAEYagoj6T4+KfMTmE9YMC+Dal2lr+roH
F/OWnYPilFbjpqnTLe8X7IW5cv4CTpwlrGAV/1ZKqLaMoMhve4IueCWLy8PY7PpV
op1Je9DvRQ6IJcBCy0OCqMSnVKrDlNlbtKhIWDdM2RRVftiWLQN6lS1P5uwzTwnf
VrQLiVZ/POeqRnJvQhMkGnWgRM0Z6A/2tJguXg37AFEYnSl1yBskp5cD0c8KL84o
HBFH6pRP6cEAEeutFb+f+8L3HlY9Clh8JMbHYyP+mo1Lqzp/mnLfuCE8jiL5g66J
a9xEKv93gIL18Rllb8pT6FeK/sibJ1+GEmMZdy77/9rSUo6/4pAjvxdiYvJvDWWo
Zu1wQW4DT4BYG8zkx583+4P2UNLEyiEIoDUIHhlGnZe+Q8DuCgiHyLcjCGFadmws
ZTsrlrEp0VnOAJxsPhZmkJ+E1hfuwApeY9EHmimKosvMXlaRNjxZMt9YLMKoApJT
8TDtWSoeddK6p45c6PmfBH+RyKMF8YYpCc7CDWjATAyPiCPI36jQs60MhTobTMgm
w2NiRr7OGrXbkrYBKUHPSSORVuKADUDNErWuPASeCAgkuDi4IAOnVCp6OV+whIbW
r4l8zI+w9XvTlPo/s/ZQu6EJTyi92fRk5SkBu7/YFgh5n2qM0EEnUTPCKjIL9u0W
v04vrt6Xw4py/hTr6mPU3k6c21redonvDdUWZpxSHcYngAw2Q0YqrsGIZewYPgCC
37DhBnCXjdPXXCC/OXXvKFiadbpMXCV1BCYvR7BFEX1lbu3MTyBKDJFgJ7r8WqYQ
faOohOEl45Gz+wBENujQ8ZVlenAAzpFwBKXFyPMVflZSgEcKyVUdC3C9TiuJoyJU
OUmDpFDekZCmEFMTtgTE3gLlqOLeldzQYGlUTzyBHKhdMOk0L1Sud8flRFdZgaf3
LvzLNSSb7nOwqJV+42VWR2qd1iFQRXUb/oWQdaJZHh0V92d3I/IAo7C+6A4oxtA5
KBaO4ldRoVo4fR2yesjNbh18X7ZbVGXt/tExwDR2EQlQhIQOAU6OdXu1rB41HUBM
ynIdiIAHUJMsBm8to6uix2ORsKkY/SLZUeYSqsm9ivZ7B7Md5XZgtQvtLipPIvP5
NpkLYFZ61cNDvhSRQo+Wk0NNZE5JJPGtTt8Lfz4EQjf+bNalJyHZOVwFc3GJ5nUc
M+u3ZMODm2GBr+kJXjjDnNKUQXR7lKagKaRt2eyDuJXvIMje2aMbOxqp6R4TTB4+
N3JATaJ6dEZccn0GT/hQ2OpOoQJ1GwVPVA3iEovWDalcZGnTug4O53K1AIehS4Nx
cLaoWLXr+/8fV7iSnABleGIenLo8qhy0fw6WORRHyuxfyDDDRadsf5MTHCqDruwv
0CywZoSSL1iR/IlZlX7tIksCMGhEydwYsMRbY9j5m2BpY5VYjp60AskZXrMDNqgP
7iN1VijPfI20YXWexbe7JOZzB+xPjoSKdBbPlzUqGbuzESDTdbv09uQnPLEXck11
RDa9+uqxPz+LaNrLFYq8uc/LWgQYJMBqZLPLU9bYmX05V0nHuX75s5CqVXwehWbr
BywpVAHlpliAxTqn7k43k0MZCOu99IEH0MbiGeW6sqSB0Aa9/eEzixxwrUmGsXXD
9nmE+91WZq6WchZ41gn7Zj+EwHip/Kw4gkk5KNJR9SV7wS+Rdl6PqR2AoUdhmFhw
KOZZQREMpYt5ytQxZOJe9aliwmKDGpY5XUC3/SQaEXI6jKvA32Eh7ntq5Lt5NU5Z
CgN/oJu/lDIf7GcJyqgZ4Yp6pgaDnVRKV8a9eu5V83W595EdorK9E+ONTQ07BV+e
wDqz+gvhKnx69EANFha/JsATha6BP1CjcSn1wVj2W2l0tMYNFKKtDz8H4vC0TO2F
4JOmNIZxHNdGnlQJW2wPj4BhgfW2NLscqNeDMQN9M4vv1IKNo2Q3tk7t6E76L/BC
2Jndis5xlSMfsoQpiFiYG004BgttOd5qF8sRSLLrNQLRrwivfuLkyV5hz5Hbc8AI
v+XPFCYa6SnwDs8CJQWzqnZk9QjCVlgUe84gvnR8AcHc7tMHS+Va6S4Wg3z2IA67
bGntxc87QF52wPT8sPA0JDxV4ROmbVLPONOHWj9Py5r4PgAwxs2nsHlVG46H2ppd
eRUGlEl74UvvoHv2sxid410RaeSbXdFcNzCwMhO8zXWYxa1qVMD7/R4++ztXsm5t
a5Y98HsIvHxLQyoctw4ExZ4hxppnGgLGb3rmPxgNMAfm1pg3ZHB5r1O5+FSJFgPL
li7yyEqqF223J8OpRcYiLbkR0X5EIpYige3fvlAEZfmGQxZoOUoahg5FYuxjgq8F
OvBOeZ/XjDp/gnZ39q69K4tksTh7Ht2vXdD3AeLCm97atDEdbQEQeucM0anB0VwJ
/yi1FiRgLLgVfcKi/C3Z8px6ChDSzNzLLBEIH0Xel8eh7zjHNERC4XPO3bUJDJMk
vefy5G+dR5ePI9mIniUIl2RjtlAmY5V1sgz0g8acFplCFYiWZIsQRhAz/TYFtrn5
I122GYaxIVM4z/WySbkaVSvLoDIj7rIjNFCrlNh/nB7AIMf9QREkTE5jehjylVmZ
GYpSiflafu3hWw+E4K5gSzjyZHGztaFOIeQP6G6g0f8doJq9AyQ7nRhVdRdV/Was
LLVthm1aADntalEGgOa0Q7LxMMpOfJ+eFTJ825V3ENj4eMNwO3Vp3RhulmpkyTeX
A1gps8kjs1JHiZ7npJLuv33hc3+dXfJAZveNFGiLOHhxK4YYkEaAOWevM0UxS0iN
ZeaJKqOseQqro4+fXe2E/Q2qWd/k04BKJjG2hIW3yL/8sKqe6bzsabK9xwpwZQk4
+4AdMEmAbWAGaAkNUpJAX6+WD/D4v4Y2yS897L/ry34Qa20Qa+ZFb9dUtJD5j0EY
pKPpNAVejunQB1HH+0LmHwAJF01aT+Z+bSwUn9AHyVHZu77WqGGX+88sZjdZRAJt
Q/m10ERFDjGr1SxMOK5OX1tLjEyRxl3Uy5Rp3F08tLZyQuZfbJmd/ctU9TllJwrR
5YIzSNU8qaGDtadWBj4ROd7Ung8cuBgOh9wr1BfMX+SwDT3r0b12nijnGkDMAcX1
hbOz1KosCS3DWJCDP5fh27NKV6Pi1czt9AmaK6HLvZuE7durwRyLZ5xZPR5M26Qy
RkQUq/CiacXLqpTPpyIeLY57HdGsORK0r7FphZQ05G7Cyc/Pr5K4eBHOPwBT+f86
OwI+GrRkjw8qRfSbjOUQC/nkkwKHzquPiKxJxfovykNo7Xcz2jx3wbnMRQ/a/QUs
3lC1ykxKOi3fp+13A6WACZxRYvC86zGsxXvDZLC4jmmc6ldmAi0+jKHr2op5Di2a
9hEKsPrLabfoV5KjHnj9uURuBtJhrGHtyxpwUUyy32k8SqIjUdDkIPz+9/3Ag+BL
NDW8PrXtL8+vDaGFdqt+C8lO0/3TA5i2FBawWNzn+XtSvO+vh0te8/XrxyCf1GGC
sp4Xs5tShKhrh2SPlmLvk7TaufRObRktUg+xpFqbFk5cdCqAHmOejsFoZaxK1WNb
QrUHtSf7JNbYGa1d3/A+vsLReEbjtHgw2x0rvJDfmUe2vCJrlCUe59x6tcjIwOP5
S3nnHQiQS12fKBH1pWrEy68/xnOQmg16Zbk3J+kvE4CFnEigmICsNG6TgELW4xb7
VrI8u0ttZKPQfhX1vGYcHRAk0Ws1bVEN3loSoI7aP8lU3T8rDoJM+Ya/KXDhGx19
OxkubJYbZWvA+cMEmrm64tKvOaPX5EJemKqioWETqEaZve65ioHljGSmvV838w+V
dPzrmff/MPc1uEPm0En5OfgiQDIKqTNz+F/V18eaKiyQEU8Q1RPMbEW+LV1Kv3or
Grr5YITc16T4b7lDDKGGOHxASZREFtXS5n5WhvdQNlv9o8bUSRijjwEgvwt7fiCM
YSjF1WUajvlYm03RGy+NW3uiK8ee8I6CD1Ds2YeuEAfm3LVToHAQ/5AjnD5ceZ5f
FglFPMaPoMmQcLtJ52ig4gVTQo/Q+JNePWBHfhfTTivw5CsnfYles1DHX5k3W8Ww
w84mzbAjb8MAV+iyqigyafqxGNHUfy2RYKEot6YGeUoFAiKAN7z7zSgacP+K7iup
UkZdkVQbmN+okD/a2yeJL2SDPoHUOX3bB+AkHiYmOPWCSA0+aCWaJy+7lVYxHhxh
Unq1F3mlc/q0Sx6E1S2hwv2h/+fxSqk1BdxGHKXBQqvr5fjmYmwiGrNuDFhNgrnU
FIVJZxAkHkrcSK3Z66oiGjt6FKaoTgtBSMWr7U1TZHTAZoZwJ9X418A9Ky05vsvq
xuLFB+pp0kB4Ot/yH067Ngfidx9G1OgaRjQUYCkMBJylRBDwTCQ07F741nkd737g
oco0+ccE7sJnKZyNusRREqlczjeatjlyxUZq+VDD3pa69AckADYpX+3pAC+jRC1T
vbNc8MWG0rnCkbMdMkN49oYa0LSNC2wg9H4QXXTgystvsHWgoB2MRRoIGFM7xMlM
k+2/2aZFwlrKmfBdrcGPa/BGItQrksj8IYjrgLMrNauEnECs/6eRVZgiHDkvovx3
DL2i8JznnadaGHqMVO1FcOIpb51ykHnRPOlB++xPcTFHISSihsMrbXNUYwH3IPGy
1KjLTWQDoJGSyA0e/peHI4Dc1xAVMwrCvGeIkledZOBanQoCDDWvXascVgk5W3KN
ViXv1uOOoKHLjsoVHg413tI+YQH3k/fsaGvZznkO6/PO4+F6a2bmLUrdQCYR0uco
usQ24+yp1IW9WTigid+NNXXGeuH7bB21iAAXm2dKKzqd7FpUWhHj+07vHYU6uAYh
Oou+haPxHhLzHIJ0Cw9kCKcV8SWFcfhRef78jDA+eLDGlnDwofCiivSBLr0XfHFH
4+BgmbeuwTUD4RDB3Wvm0YP9kx2FR95Fgbe5d6cr9ze3qqO9JY06HOqgDuClq7Jo
ZDFiqaGLtKUbpLlCPW0Okr2k2H8sAa2HnF1g/Kyogmg+ebhZndxawvpeg/sRVlgk
MDXFN0MjzabWLUEEX/lOz01gY8uNsRrHz72QLdBLNcIJNfuYuCSw+iRKHyS+szKW
FHkBvSl3bxYn7vKbSjKN9dbBbfZsAjVDa1r8N09IZBZ9Z/UcrjlXpMlDBE5WSRMc
x7WKulkpROSUnh9LMlcL/NcjoU3ChagbWFtyh+ft7ipKPCwXYGG1tqjeBeHGCeUi
GrPuvlcSmC73lk7s7KkifAVsvEp08MiL2VmrIFgE6CqefwzQIqjy4OF/gjW42Rz2
ihLWAbuOak+zTcBs2WdkP99MLAM7/RxdFb3xZMt3RJrqI2gmJiyRhTyh8TvcB2BL
f+xcbVxKvz5JeECDUHM3/9K+H9qtk/Ewz4vB8HBaVfGk4b+KZBUUbrWcYs6m7/1Y
071WLlErVrcXFHZbdoSXMAKaAmhGYpFGhjlU0OPsV1Ubz7x8aQ7+Wtzs3uAP5aWj
/c65eL0KSOSDb6+Ix8aqXiKzRGkbaYBba7yPPZXXR10ODVcnMymJaL7gQb1OFeVc
paQHSLJTMj5lcqxbRswKY7aJKutXDPh7SgNfZSFZRH/6fgRWVETaiawZedG5Z/YX
2CqNLCjqsPB0BYlVAd4h2/RqD3DjSqiCrQzNhAcevFElZwKuZz3yKhrLvh3HKjwR
MVOLrMvgmkhVjGW+e1o9EkGte7yhu594XXlaY134z6KiATPWWpjdXivSIcM8/VW1
iEn/VyNo8zkQ4vSTv30l4RQ2L2O8qmglH2O0AfdJ+FnCA9gqFpAsWFiqg56Y+Kbn
3WIB++9j5XLgadO5ZLc61wGpADcjrh+YjA+r+QRGoX/6/oEW36ZwFKqvJde4BgQ/
MiJNOZR5iBZ8MTvTn+8hPqmoY0GFf/CbpNwDD2S2Ds9ogZObi/4h/Z/ovW69BVAp
0zzP37BtzfWvs3pV70OI/RdBKk9sHrQMxaF40DdGw0fVcO9N34Pb8TjOzGuca/vU
LOdSj+wDiehRKXj5hMAUpMtmli6I2p9cU21cB3r002GuYnQUxnfEACMndxrhq69O
uRnNLP2uy4YN+aPF8hb9qo5HcI/tlTjaqM+jfzQO5lnWojMsvL6EPRHc7DJg5FC4
0aeHjy0Bktpw5cIohbqPRiLxz7PcxhBbgePQKpxve95MwBZRQkEbq3F8mNlaUvAY
CBemKCaI5oKE9al8cZawy550OtB4KzIUNluGYXGTzdaCLZjSIVi5lQ1oGqzSWpyE
FMCpzrUulqsVXpu/Tk3DA/PWMYKMyDMY8NpHf2D0f6z7L8vE0OHaSzDnuOMD5N4L
pi3jCw/bG1ZGvUqYaV0mSFEVf3Hoj0zqWl3cpUihcuhQMjp90Kph4ZBRLqiRItUn
GS6oie6Ftsdtde5RFm/hU2DG+uZ1F/+RKJF4sB7d6WJ2HgwB/hKFgW+qOuATPxJ3
SvKNTm1B0+kQ2/EK4V3NCcUHTgBMDT4YIdVRbVWr1mGowe6J2BPcMVOD5fDVUxt3
COzE68TETgd01rQ/xViwmfWdA3+w8rPCqTXKpZQYMf7g9SyqN4PlAi2lOrJ1rP4/
55S7wxO313006XfCIkmAZxaRY8aNOc/uR3SqEP4i22sx+aycfYGbrWkvfX7VA3qo
NS+40CiMT6EQNLvJ3Tzw9geOYLHC0rkFFGzM8dViLYw6C85QAz0rtq0+e4d3KlrB
uN7fYqrO4x9/iUrH4Ohbiih/eK4KcTvM/bNyHm4WK+RnargK34PjqmESw34ql/cl
Yyat6gLISFpZtZfpSs6FWjNGg0qOAV/FOZCF/RoXCNY15/uzJBgVT8nfs7EQf6wT
qCWPbOI4ITU7q9aEx9chcTgIVrIsqAtKxWtD3kzDwRdIhJqkGl9YdfmRq4yrWxdj
NpE5QAPoqEmxUBg0Tb2KtEbuowh8EqbHGAGydlpfseHJDgaVBxqXvqk8WJ7IXsrd
8/rQGCbCAdYwjhs/JGuuEPqDqDqVAXNeKU4lNp10yMWBGSR6fyNl3UuugtxkkpSy
vS2fVGkY2r0R9LPUKcsBg1fggxJhVCh7OCSUankLlDHXENJrjjQSKjfZl7689Z+c
1/SthYNt3EeUsZgv1HLZd5PgpKZD1JKUy3PiXxnTTOR7V8PJLVZyw2n8vhb3hAgL
cc1rgvjwn1y50e+WclGSRQKwQWbI1faZOPm/nHSnFpkyAeFxTbONOFt4hUmCNE+y
hfDewOEHoaTIhd+CXRzeq5i+t/ALD498XU5CYWL93/LJ0XnIN8VxkTo9kxdtFBkH
yPr2+iALv/GSljvAwJf5yjNDk5g8o3mTQZl9aSr8lpGM6aCAN5IIzXH/wiP3g4iD
ot6/DOvUDaYDSYFbrRfCIK9cHcUnhkwiQUoZ0Rgo0Ny2B/wo6cEMKWyatuiEUJaG
mTea7BebjQv4+uMibzosCyMmxskAkNZPF4wnAV+QOXFTuq/0ZTDchTlrczQs0akm
vu/LoJHUvI93s/qphLFgAJCXcz9YLXHYe84FAhwHL0LHl/IPVbIuOZVppqUfJ2be
QjaLXCvGG4bsgUYzeFuOhyh6zzu9y6Z3DSaULcbR1CKzTpjD8tgW9eUUN0Tn2Rec
OgQG+5BSyoygWOrrwPA5Yrb4eGoqqDFhWG9GTtNVi08VkMkYXRDuGc61TnDQba+v
cwDbV7XlutRcZjAO5d/6MwXJpQGdGp3dqwPmM7DwKytcjhi82cm62WXrQWd/Rahk
Gz2CZ9gMkMDps0e952rxJpbVF9Cq+vBJoxL8B+ePfXGNQ1Lsvywe2JhdBQTV/+z7
Mx+hPLPiJvjcg0wiA0H7ZpCUhHHGhmlogtRJNOKtM6j5MJ+UfsT6MU+YBUIZ/qMJ
xsu5/hHVzJS1CsxBz5S/7pDFWBSyU+zYygpBm9KMHoFbm9CGMHU/glnjuoQwRwTo
EEYYhNYKLcsNegZ4Y8Dm7HHwVt6davVhwkk5HWcAVf1ndShxPIVYXR8sT/KO8GUd
DjuATiIK1Z9zi7T4AAJmfDK3BpdNWW9aSVH6uofV4VvCQkm0ewFxNeX5/deuD2Up
n7p4/n0CrXxqctNjqvm+WJ1MQDxtB8nx0dbSMHsYRWy37JBCGLK7d/G4dK4cKwvg
wJAS1QrpGclDGeDJWWYtPNz4CcYezo1RhZ/tSX7qnBZi8asjK0URPybirRaNlUQc
2XDKbsVC9FtKeyPnAfS00cAfBil8BMAwwpLD44vyY0SdTt8F3l3D5uHM0zK7gMx6
odeXmD1Nx3+r0MjkccbGrrYZYSWL3dWhELQ936ZMMA3Ew/u3NPTqZDmM8OZHuAuT
RHFkq2vCTRCngkFsfxuFGfMDi5z5S5xBaRmorW5YldtZMWdqujLBk2um7qzBFSQo
H/JDwJA3SPRyti8akYQQh3bosuUXEG8ft7oghrm8qWprnBh+yVRVeYXZignhhAjE
TNskTjj+lh8rglrsigXnne1cfOA23FxpBmyXguGa+dfU2tAlkQUFepO+VgNRJJ+7
0YO+aV2Thy6PvGbP68t/LxgZbq69M6xbX4CvK/1tSA481gV3QVBvRxSxTppcrSqK
PwJeko77eNZwZcfuZYO/btFrCVsyTWrQCLprRQU8hMtoXla3JzrUcvDUO0uUaiHn
qqNa+a1HP8TKkn/KeCn0Y6DywdwhegtrP6kxTbk7yWFGFNVVtve2JpiMdeBNSqo0
S/b4bnhG0BAuLf2UnLi6GC8F/XjRB46yjebBwVwQp/EYUQTsOKAowyO02IRfE9kk
tcGgOyKy8+o6bg/eo1MLhTSopheFYcafVv9HHKkviTk5XL0HHwawVTAEMcsHUBby
39YYqtb0uO4bRs51g4dmfO1eMBAsU1mftwFKwbV7Ygw22hORgsGFl6K5RHBhsteD
9oOK7te83ux+xvNq7FtQsBiKnu55di8Wz1sDDkvL5xlBfkjJ9Pu4kI4RS6s0I0/C
/oDprUnuAGU4TtuLUvmnqP+1g4fQi8rzXt1QQGlv9KXdY2oe/cU4Zarz3/4iXgsz
ermgdsGw8u6OG6CvXTXg9WsCKD3AI4GBiww1xBz8jRhBiF2icLSHpYHXHVM8A1JG
i+2ib17zGtq5okx9ZUJSnquuXtR2IpduR2kGFmvAsEhI7S2jqmXmxIPyrkKlKlBN
LWrx9ybFAwPvZeq2ndd9NUgUwPAZ2H9v9zJuchtIKt6zX/2QbXTKCBmJFlcKEQAJ
A4K1unx26gK+dqlqpNejwYcq/kOBNfxCl1zQn09KlxergGQlHZUk1ziQu/WiDHZl
Mb6m3BXRaVa+YvCl+yXMB9/qljFh85U6xoTxQTgKQHXNgcHAh42LrAEztzpB1bSl
akGoeC3KTwAYBmQpoYbv7psAXN8KiZGFyyWPtpOZAcjKjC2IDHB9eR7p1xYSoyAN
iJPg1C07O6ruJ7whZ3U4Fc+/RkR0dOc/T52M7/Ow/DVLnLmvUVVLjE6VSF2Iml40
2K+JA3+hiG53RhxmpGPQ4ewfIiRMsLivJV4I3yAgWUNgD6tsG2Ia4z0O4VRoFPsA
w8ck4uXTq7E9tPJq2eK0RIwcNfMo8evBAtteSPXeIx2ejGWGFBCbevzhB4+albCc
F4RGHodXw9y6PLuFyma152kAmDNE3v5UiIdnUXEK1T9YOtV/8vZUoxpAtM9QvEKl
Odk1XzCZ9O8W2nyxnWl/hwcJTzcWeYtdSQXYO+L+xavCr6ggQ1hAb1BVF59CVOim
ryGXwQozAsO2Jp/YVGJ5ZpOdwC102TzdTgH4Xa9JfzMrT+P19OOLzDHVky7V/1QU
UWyMZbHezsaLFwGl3G+x2j7mCOY0+858LEgD/0O+7UjQy235QKF27fr9i1dQV79D
/1nENcqbydotagLrFVvN3DplK/1n7pHcfwUcRC8BNDkmwSKalC97wiBUJj533Nmu
YRYXKZx2sm9dttrEEDkwyUomP4OndC4mKlvFkr1QMBG2Im74EehR2GK9KGAKy4UO
UOQAj/KV8Psg/hYA6+WDoKNvls2z7/WYDT3BLuYcLgcxfPXwu6vpmNRGRrSA9RMg
cfk1K6EqLrJAEJ9KWcYCADKR5tvvwq5kU9Z/qzm//rwBMUK6roBwym9V8Y6lCDQE
0bkRlvDW85h/xscDWsLU8t7iGKiO+4S0Fdj7KQRUo96nJvhYrbG5uG1gDwVbwhCR
N58C1Wz+S7kypspGUtaNW3YYRizwu9YGNNYEuvzzXn3R8Utf9jWUlV6HmtvjIthg
TwMJfdjaNU5qAgujvB27301T/1IOBOnjtdEwGb0WxvtPSt45J+8LcBMlwSVSQkDm
wHUZPXz4TBfxuMU7MnpiiQDD9c6FUlsPGVbepGLNtkpdsBUPnBnOWy/Kl2Bv4uLm
gOEqooXMY8pthKroTKzcjLjJpEfIHL9Kep1Snql13gsf0fnxy+PLZXHSdgGzdFbg
6N3IOaEkuZr2PP2qr8HZsDaLf2qiP3LVDAdbOLXImq0/uguLSi0wGEghoUOyRowD
zS3yzvkYsUgj5dXzsUtwNWEd/Gj5EX6DIzryDX1bOV6kDpJ3s9N2mEvYkc2ittb3
AvbOZ8l9aaOutTbPrsFV2qphQnuI9tlMZ7/M5m+Oa1aPUpLEv+i+uMSASXP5gTEi
lAvrRaivhyWHARAZZp6BY7/T7Wj+iVyQsxL54jDzoXXI7whs4ORQDZrTdyy9gUFi
JeQHc1Ph3FmV3jcrIOudFcAi0wfebR5bp0YXI71A+L4S1Hs4CwpK+s8IMahkU1O7
63DuFs5AtQv1niE8WdGFg6TBb8uWyriw5suq8XnAxYwkGJ5HAAAqe0xeD/QxYkP/
5TkoesAkWtoYZcvGr+vveLQSEFVmlEAt9ca4B/ci/yRZeAXNa6KIO1A2+9Nk+eNo
1c2OCZCGlp1OgJevjwIJuC7lMOoBw1ea0BtzDxPb+p2KTZvpQ0wHquKbyHDXxinf
dF7Dj1RwQPRHBGUCK7gs7hV7IO0O0LoNNAgzgPy1x+U/+awMR6HloV2iNjY5V3T+
grfK1HzCFp1g5J9aGT1aaQ6g1xwdaGvRSc8VGAmzANH5LIV6bsZp6AmgUrXQiOIt
ViqwlV0uyNv5q/7XHlrnI1OdTdMdD5ftM5bhDK6vR6V0IBNGhwcTQAQXPeF1AHzg
HwJNNe83BDKtko6xtcqzul65nO9IpqqGnJ+U93g4MyijfJBY7lpcRZb2HT/0OzYP
4kOF2kUc8qyam7VdzW/AI1AytHWaJmUMFoCvBTKNHKRGp/0B9L16xmdk+1kZapLX
2mJzyAjzWYIJ1aQq2+xdRkQjeL6GQhNF5gDcYdf32VYRqq3w6IKVzHybctC6YF+z
NzofzpGGwNGFuwtQcG8BJZdTOP9U0ZmxnSebflqtiaU1MJYhTL/Yve9SGC/BXWGs
7b2I6/lQdyC3FJyfwyeh2we0zTxwPqM6t9OFFXkE6e6DMIeak2mXCuzdfa65H4QM
hBuprw0KckjfFTpPy8/73XaT8GIKATtO7oJ+Oe3+O0293IWUxE6PjXOtUQJm7TJc
euPhuEMOFisBfA0vL1uQlG6zEKT2kxWU9nOqrW00AqhTA/vOaOHfCmWTxogPG1ac
gnpjtB1cgDNs8kCMYUN34NjWhbxblj33wieGQGfoRBq5eRS18XzQUc5mNcRoaCgf
Ng5olrdUw1+rRGWeOyWl1cYbdbsX+wD1KebTVEdlNx9WRXjKipynJ1RHmX8+zUyR
NHRmJ6AkmitPgJyKsi/7emcVWfW/GYBZmnpAxYyI4275+aU65TeTGDL6RYqhllat
4db6oZUY+nPvFiBTN1Sf5y0TF9mbiiUmlngaVkVlWYyFlukUaDgDYrsrsCMGB9RI
bnBLAym1L4CvjFcob6ldwoNfBseKvpezDkJhwEsHWMvV9ViDnC9liRDenat7erLi
w3O8yNiyqPCZ+WevtEW2vRNw3GU/PPxYp4Up1bYwmFwJRc6ZyvaksQhiMRTBYoPq
ZiJQoAZfiLbY0KFQRdyuywH4JTdcVaDys4J4T0ZX2ujnts2/9dkP8PcLK3VePGC2
nDRNTYaycSFgRPnwyXLnzrcE8qjXnKRypUxq8CvalwqC40Gt0uEdIqGPCVR0P5QT
+CUoY+oojAIiH1e1F1pJePlfzqlQ3AO+wP5GiFGNzJ7xn1v7tvJpllLYmtsZWSYW
0UjkJ8bb8XDYvdZPNYUQExGbsDo/T5dKEIBfWSJS98z4l3JKEGEL5XgdhDxPgOWD
HvyG+CimGFqwZXn73u5NTT+XTO15mWa1qOTFN1yk0cGPok6cPGSoGRY+ZllOfJll
H5G+3n0uUl4a9MvZdOTaS/EKGleVDcohR17aEkDXgJcgzn9Q9tL+8zCf+sNib9FA
mdZtUqtTlWa/dvIQFdVCMTF+xEAkZwTDFR9fgubreFj8oHLb+mB2O6lbIsTZ2CWt
m1jLhS6LEZDMDZxj7z1SIZrwuD1V3tI6TPY0Y2O6gNTBAnPF4ICPiQHo/aLKL48z
PDhZ8g+ornSIkfFvz/Ufl+k2foXl/8pLbSDSJCr0C6E/H4J7jy2XapThm75Judj/
NxYSteBtqGeAOoZWUhaXczRNth4E4PNorAC5+TR6rdjuQigrFenBorA+st1mCRIw
Xr2+ZcTDaVuDl4Tg5CgaaftfO+qkw/uuA5LuLwRlt3E01zJHc6XAL4/W624sfw9i
tdf++yVeyF54JtcOhUITghlynIcUcuLJLqeUBV35uMVV7cfyq8B716dfXf6uADHY
H3QzUtk1T6sJeChDp7HHEx/UlR6zuYZfXE+6ggp2VIJgsngiAxa1rhq6q+A68rDx
C3gCRhusMphH4MKDJ7UuW25eTivp9o1YK7RIjlmbiJJPklNtItXjB2/SjKfeZ7EG
9Q0jhPlUrWXODcJZKaj34kJqrrgXm761Uq+qy61Q9IDDu/vk7F++WT5s2TEsJirI
qGTtWk04+2Zdzh6cB/64bdLn4hizO2IGT69u5ObgC8rf/WfamYUviZKVECO6KnNy
vaND0R9INtHzulTbIWabZlNDxydzM8E2TbxyleOgHjp9G/EM//RQ6mgRo9gTAAcE
IoUV92peEHtZDwYIwJB3R2id/6nkNCms/H3Q3YG2motbOqK7S3JZAHCIWJylLqMM
7ckr6915J94Yqvh4PvHC6IY9nlBphmzuj0IZYs6Ij5Oa6vEacokPTJ6ihsDJe3F9
jabZPi+l/2Y86OGTcVHgY3OHLbcC3wDdbf16vJZvx+ApmyC8sFf/SP3Ch4Blrf1n
LajsaDypQyIoNzxM1QY8exENJmxwBHHdw7eNJ8n0vMgXRK+CSh+FTWKf8Wu8G0HV
lx351XiGHN9dSsoyxk7+t95qfexEQiPwRkMfESS0Aul0QvG7yiUWWDmR8k56tVYw
kErifAq0cxFs5g8QN1JCLIZ5T482hdEqTmvmTK/K0mzgR7IcJusIKnijPpvyuPRH
2uZV2m+cTz+eZqXnH6nZ7ui2C3vE1tgc27WcAmQS9Sim3NNkMi+wxNpEUQu6S5OG
7kUgw1VFctDRZRi1QxBteThAaJt6mxnF5XSP39D9s/t9SvbM/WGxEmy5NY2gSu5C
2FCpRrap8Xtk0Wk/yYrUB7yNi5FFCqaPUgvifg7V54w0fpBSKNCdK9obTt/IxVlY
ounHjCPOTHw1Sswfc3tB2WyO6qdR6fJ+/TW/lpnEHMqbosyRGv/qa5kSLPFyB9lR
bE5/K2l9hTWo6af6ksA+MN6BBLflSywT0jqw4GoOvBlTkG85rB2BagLnHOOLeeCZ
qERI22Ti706MEYMRLsKrPEQo4zh14P/IzJApH4e9G8R0b+gquHDfl0araNjuesln
RhxOHrUpaG1wkf4YuB+eOXyn5HJyIwvEBljEponogtVofRcxaUV3TaS7NBjp2Wp2
yke/ZXHap+yGW5syxEbphona9Eb3GAvdPG/fbnfsLhKl21KDYRFtmE2QQEVRj6n3
cGhYuAxb6syggRXtVRz6HwQdQSlNsD+x7spRAOyBOwnRkZsEhIoMvBHO+kKXTcdj
Iy4w85q/zeBtW09Q2+EKCBOK/ssLXBbmKaFeOAmC7oqWwGW3hgwhbb/KEcnoGW1N
0HHNzkDLvUfLoIq2mRAb7HARQyMTJ7Tm8w/HGWzW3EmZn7ZALU1s80FzRt+dhdi1
XYWFv+YLahB4uBBmckkWnCix68KTwzj2KPGF651AGjyu2R+8e2ks7ffa3il56IFo
asHXBFrBZNzw+yI105vXxUMv7Uf0/CGnTsMmbIDBo3r3XgBXZKfqg3oGJQUZPZan
saFvBJzjwm0hOZURzGldDb3/Z+ckGoaYVxo6/bpYxV9HkmevKcUb3K8+BINPyrzo
fVZpNTCs6VdACMeNOcfaJXi+8/s/SR+AYlAPAeTA398fHFfdITGUeyVCHCpxNtkS
CYANhqQQPVmYzeJmK1utI/O7O9EFH0WVvlNfblJfwQir+CUzCa6HqvL7qsg7qSiA
uvKno732TYndMUdoYHgZoxpRpIUUfRiqG9gcfssxOiylcwF26F2wHxEU6FyQQiFg
AJBpffvBbCvGR3ZhsEOE+JkY/Vt4xWsvjti5Pum6vR3dBTjVbDUoehh430HQ0zX7
EnU8mkXOFkfOY1wNaHxeU7A84YXrMoz6GhK+PjrFOc//upQXSwiMJ88cHKpN5ckD
FxDdEuz5oKAqA5gI2q/x7vSncq7N6qqU9yf6c4of29XMRZXysXGX835hGrXDF2Z3
pbHuuNZqal404bWl8P5U8QX8VSMf/z/n5PhHqj/LwhMRGC9VS7FJ7lYHJAtms840
W3EEpIJc5m0jLloxqX6Sq9kcztIe/mrMylJwYHBEu+nVj0Vu+B4MK/8EouC2rta6
8xioXvgamkVkojvKe3xEA9T9GO5SFNGvKggRHIiYQD2dR29DfrAsjYdP1evta3wg
ebnSi8gs5f8/Xi1orRqnnczPXuIdxdfSGlh3HvrUQuyz/czbzTZFs/S2Esquukub
y26ZB2qYijHc0nknCDaupqOFTcJfJOVPrxi9xDhB4pv5xf9RYbIek9PIqwbVwQV6
GGKLbAjILtnRjFUBe1cBPXpS4hWEaKIglSxjPRkwTSlZVVr6q1oqBqzGVAIP6FLt
VvXffF4RwWADYVgjQFMj4TOl4n5GE1cHPaBjjdevar8MBKkLAFfhnn7MHOzMQHcO
WRe+9z330iWEoaz96VfEiCxss2nyBk8HQauW5dXEjGod8WruLx0uHRiGsfcujpjT
7qEFgDn8e7RKCVvMS1cRbVIffso/32BK3HupluB/mmEPvC2UpSuiyIlU/yQZZpAq
P12MUQc1ytnfON6SmBJCpxpplZXR21Hm35r1LTOeXHviAXpA1DCD3hHmM31qxxOf
nEdBJDyn2EL+9Lo1/QQ2p9lUXtFCxxmHN5ux40yD3bTzzwwT4RaLDatn+GLN1aGW
Me5yQVKTqa3oKlzGcPuMvhYrYWlOEvm8Bis5sczv19EXEDw9QChuZxfJKrqpH/DD
r0q8O4xBDwkqAIGoy/qA1UJmBj5EDLx2uOrFZ9Ez5qjoyq8t3+VBUIVLaElsHBjW
K3zfwqZ9XJl+F1ApI/zQPsaVs+2Ov1EbbRSGugPLcyJM/VijUCmgUt5FYCYtapeg
p/ZNvdJDGJ+HtgQPR1kilE/7ocTipwsESi7EtEJMFJmHOSw9+q+oJI073Q6n1O1U
K/cfsZcY1ErloOurgdeJw/l/XrBXah2rgIQ0P9IbPbNBB4Y8DBcgOeAaze3w5q73
rh3da07JFHr6boRiabRsosT1YRKVSXNmQbd5D1wvxiUhOBpNOgIpKXauK8NII5Ob
DsHMBnx3LTzVyIrhpaiyNvu1+hVNvXOX6dpzNBPk+P85jhlkcIE3oER8s8kmEfPJ
UwAhPKlJ9eFEVeG1LAjEp8BB75ZwlOwUrugNoZNKtBq3sjKZ8raAmX26BdWOQ2PB
J7nsNpKu77YgCfcDTru+GnlYJRO6mWSjdlw8HEQsqR/WpXJlpT4ZTIPEQeqlhpWt
CDoLqMwGCkpnZI3EcTe9azY2EtsalfW+/ZjPn6MxtvfvqkB3XfoK3iC0G3Q3TLba
SGSlwy+IBTYu4NZ6y3BcoCLl+8FqGIttENwuIyRK8C42P/DZVsCOs0u3b7kLmmKw
5fmL9sGFSWVY6kVmJmzC/fYe2KhGl3zCTs/p8THjig8ekjcr243hstg3Xn6XjvAn
BZRPex6hQ1z3yasyJ4k5SmDWcQiGmckzDByAgcJW3z/5DyuuIw+i+5XZMEzqHUHd
WVh+q7YdRJEvG8uBGZMAtsuumdq2l4IVAAFQidmi771iK7Zs00Az8ImJIPtxTCgy
gdieSTNboQ/PC0iAV3AW/MMouovqWWurHGn6KP3B4OLP36bWPXleULUmU/89wjCd
rLjSxYWEWegGrcCnVRIWgJYJsEa9oWEtGtgJvVzBWpBHwvTt7jJ7nvR30RZ82yH1
MdHmnTIpMg+AI/EBWdZEEoUoxLX94kF/QHkRgVVYBb0vsRidT7skp5tjsm++1eQ5
ov7v1UqqnLbQBWC5WKk+jm/JRFbyOnS0N4wwwX/Aw1cS53c4t3GPsmJvUaWQqJ5r
PVfdLH7PEx3exqzhmVNL/cpatcg67TQ0x3XwEBuNU/zL62ubenHef5qO3IBtRAp9
ysde6dmKc+/FGStVZsAUXwsmnuQaQVjBefywnVBd1EnPQXuxwSuz1EdztOQyggSq
q2IevwUXMtmHEDqCSO3PgtKucZ/T8noxvWPoYC7t1CAvrFqchFcabCi8qcsAfVFo
dS5Sipj8w7kMx9RGmu0YBl/OnuBoAaoNDAPKSiu5XbC9LU7so5mRAcjDr/oMfcKA
SdYA/NdCvb0qn/Tvr7SDk9jQRNm7ShBsQP90Gjexdqz4adjZB2x2bUkTJylE9QtI
OuFwLK7DAPBK+FL6mNM+w1lt8bENltJ3I1UxmBu/ouXMgmKturu9BPh72AvAVM97
Rcaoq6QxQczQGmST1NyFMRDWMlC8yd5wcAdJhUTfhyk/24hpCB7StWzoeyUt/wj7
Y72nfl/OH0gP7RUcYrMQblu/+P+o63k0lSelLS7N3cAIg5fhL+0CScSk5C7IR0/r
ok3gV1jTgt3zoEEBO3CX1sR9q9vumyy8fsau4o0tkA1PHQGsg7kA/T8mouyQgZvc
mA++H6HJQv+7JMufG9cLv8pkxQ/A4DwudCX3jbj2d3/71xT7lWMoAIgk5qRGJhbz
/giImyPoSIuSR0LWndA/qLeFGaBwWuObYqt3bCt9psjhnLu6+3Lvutv3ZtynXPOP
crooT5eNliRRr3M5LH11PDVn1EYvkHYdWneBHfq4aVHhRTQm2FCJHYXaHestysJi
HjPIpFVAgRguXa7zoR/ACun8bvKM2x9iAIeqiS1zZEX8WEAwkzTLYUKr0BRSPisl
TLXH5Yx0IscjWoHA1uofRgl/nutak6a4D2HvTt4X0N1A12vPSuu2R2R8ssQ28U1C
ckuezobOvKAGvb5F1t9hr4JpZxyzlkgBVr3TMOzxUDEQX4MG/X6juLM7mAWyfifl
n6RxVP09AT1rO82y6EgjsE6Gj98rQ04SDhg/C+UEM/wOYuh1sfEYq9RNdlVJIcnO
mrjpZ9FyHRisPzWQXlqSqG7xJO9yDUbLnHqkBFEilc9w/EkXrjHxm0fwOq/H7lkN
PPiu1nBEeSA39c101H6jG45NHbWB03zGiN6uGx5QD+vkP0bZUKWFBQFALl1cLM1h
KFmRTyLYvcQ300vjPX6Ld3tGhgusIYF7t4K6+WxLn/xYB/TykPChoPcTj+UsjaSk
YJR+NvSvQTLW8v00uvp+wfzrDZ8jep/ATf/ZEGNX8rYXYXQ+luJ3q8hychEKRUol
bwRbMxD8K/T6fBX92GZ4cRFk0fz2H4G9mjFo90OP+lchWY7VjEGUMjmOADrE4R60
D7wwvb9yA7deibX6jIGpAkyQMsIMAmNS+G8ih4NUb8BGVvnFCwwpRcYlBXKOxTDf
rg86aJm6qKdXwdvo7EdTTV9q8v2Sw/AvcaU1FudPGrjlijvUqPQ17OzylE6N+LUp
GDh1AOP0llRbUlUrDPLOn9R6etW2hI2wyHk7dt2UkVF4fiden66Hvl0qfwi0m92j
VzldpeF8SGFp1MURyoRSGORb9UIsChBsJ7k4I1aGaCb7tdQt7v1uF6GgfqvJdWr7
2kkmJecrWcAi3+QXSagfwwP8qsvfr+rpsWS134Px2wKwWauWXFogiUxCT8XkGo9d
FpgglbDDz+wfV8CFlqS9tB0LUJbM9ovGYPkdxpXn/l6iC9I5XVMjSG0UIODnf7YE
Vjk5Jl/RgF7IMQ94Xi5M8SyErWoaerZ7QHF99DgYutsIVjtGKYSjnYEWNVioaF7T
XDlLfNB2gww4DuI9AurCKIntNMNmKQ/VeM829c1B2fDgrNkUnA4SKDfPMrbM69NO
Ve31Bq/z5w86aBEG0PI8OpTLT3lgxImCruthKiQCAHT11oQovgzL7X1C1qRAS9A/
BJvrnDW7HBphtlwLFo5f9i1cu5W+eFR2pE5Uy+rB9Jg4Q8WGDVvyWpylMJymdvE6
1hQg6qDmzEe9wNJxW/+PlnhlsoOSJGYmivr/P3Wx2iAPycPJKknnefZ2jIfi/NHY
dnTmBmyhki00HcD/Ze+9NA3HuTFw5qjWb3f/XSSe44Fh532f057bOzhrOaUUw66Z
GExJsa60a+pDQgadEVd4AlynAbG6yy54XxSAJAmOg4Y5KyG5Jn/3nh0cnB6kHNqL
L+UQQ1uH+KnjzOzMBlPf6vyGd1cv+jQK16MPm6spIm2LxuoiORZkBP6r+gCHxxPI
QXYObHKLNDOuBZdjwvtpLZgPT0n2KiG9tVxItPnu097FBKuUkVhQsiA+Y+CWk42p
jWgDsrhqVoPXg2W9Ga3wyzF2vQWJUM/02EvqtwDgqLVX72BApVpyjdqJlPCB8vTP
CB9bFnrk6f3LAAh7b/185IAV1KmdJR919vmbF1SkPfB72D3/RqQFfWYzT9tT2wEU
mlqe5Eaxwr+wswRu7qpKvXVri+4W8Vxxyz4c/RG2HpW7fXm2edQJoftIVFVzz6ns
J6azKbSsI+6Oo9Coi81WhjXOAUDKH4mlBAzXHFHd3aF0e1jv3eugudy+JoYYZe0N
7wnPAkgOVYGea+xZorUFTqjycx1jb8K8AAHXZhM+QXftlWrF6LV3G6cLP7HptzEu
1OgGTKhXXOK4G47DuZ9udaohmXq1CmzNWQjYAw8hRqFGMfBvgFSQHtdnx8k44Saz
OTtBNAUam6KPaxlqHRlidjSQRluIM2xXPUA69SDM8fu2gb1NlgPoun7slliWvZc1
EaMxdv18oohX76+L5yE6EZpvl2yGwtdxRqBusNWA7slqsNBqveNTRv8FIab34sUc
QjYonXboYN7jaLbm0ZTabE8F7yn4VSUE6iPF+Yx9AitsiGJAxoPFNmOmUqZ7dAG2
RLaAhsWRVL3h+SDfs0Iek000R6Z8V1MoHsnREdHHWHOGmm7Npqvz2i+jcV7HuI3D
ZJ4Og9AnFrN/t1QEjyRh0DEjO4oR9Wf5ntpuCCWMVBt7+fjNZ+rkSQDt81zYs4ad
TSwHk3imwt2aME+cnSpc6snldu3Zk0rLBFeQ2wUuAt1xl+3Wbo4lV73WmDNqD/to
zJUSZS+CrdsC5xL01b+AGIbiX/LJTh0rNXb5abO2BYOcTgI3cDz6wBHZvFXIHtWa
Nxpy/b/2buOAyQHU0zOgqK1BLEW5Z4AtGeBwimQlunFwfTpPAtCN/wn4IBTkRL5c
n2T8aztGc9UAoeHnBz5BIoMo3pEqZdyURVt1cQwiuF2Xf8XRoj4r6thUweTGqsg2
Gio0oXWojXocGGeIGgLMAcnIkLJp9PKIPwu72vuYa+9CDszNWnlCLHWobmIvk19x
VGTPcN07+9NO5e+5SgKmhh1hUf176dTMryZ5iG9i/VpbVbUPFrnrlvengTQ+xkFj
ZzJUWfuLxNMjypNb/k/vnYKbGl1SCmCewkHG0f3yQtJRkcgoPt2MxfrpvYwt2Jd6
X4ksnDfNiXdJ9s7s/3xzCxhLDh4Dp5oiZN6DhOvlLA6U7U0NoI3YOX/QVTulSwDg
FdBJdQvpI5ERBfVgH0U8nhdFNnquQyMQmUkjyWseHR7/kL/4mZja4SqIOwDrbq0P
1uOtVQ09aU6vI4DjhsHBhZ5HGvZbC+ozwlA9uGqZBWBEZ7XxKe29CPfjHnJPEcNb
/H9sVgwF3oEPcp1oGpnI6PT3aIrLoNpAA0Jy/VPz0L/Z1onbWHUfHa1ZZZPHpnFK
VFR5SLvoRxLEw97LlJjnbQvhEAtuiBNsjuIN2GqIP4ADQwGzeEgyJT6pkPE9V8Ny
0GUaa3Lw5TWGKHKIBrpD7wLIXb334GwTZ1Jxz/+vSB+lVNEDS7pncJc9fab+q0r7
FGlDbPWpU8sJOAXkNc922GK4El1L/pbznaaqyjuCiCB85uUYsA0JwiOXdITzdfeP
8ctVN7lf6/Cbam3wyxI8IDUpi3Frptc59me6vorKSEiYSNtMq9aBwdRRde1zUr5C
RBDGPqY8fPFIKCq48Wp55DBB6N9rZRTI0l/rS1FiIHuZuH3XjcvNnmbroeh1K9Yz
cbQ5BFcNiCjuaDWW19YunvVOcrs0uCAv1PpS9O/jYWAHq5gTsh3PI/yOpCnzdxea
e8B0tHGbH1KIbJbeIAGcPAgbDeWNPcSYPelbD6lNkU/Vwn2tvZvuAkZ+iHfEYvfW
J5KsQZBJjN7vB01x0ct7p+e2Yt2KU+aPKVZ/r9wBHpjSeLN+MjAWkjTMMm22sBOL
Cp6lHuoveTgGIEEZqj6efUgUgMUcl+Dx76/ETzP2LIG8PKewpXBaXRghYqCP2hgs
RAtg2FON9fr3AGzLVWnWhGRJbv+dL+jOV0L9dzDqdfbVQblmBXVnWa5cq+moZ82f
+nFOmHE3SXqnzYu4ZN66nAZG0ISImlZbo+iqLnIXzlcJPqNnBTkFGEkM0C3Pk4cs
WN/5IMaVRFqzZjOKop0ihQ8bUPqfmZhZ2kBav98tGiieESRN8yexlGaKeMiUuoOI
Q0z1yz59zGxZo8eJ1AnU3f3YL8Zqma4cE8/el/1FNT3NB82FQdMBwoXB/+iYgINA
HFTWea05zs7D6jenD+Ev7WktA5xhirSe+Lh7JcNRm/cLC7Aa54wPzeSmKZHDTPaD
OalSbPPzt1XnGFixIBVbmQi6EjnVRwfGnHUs7hHMVssi9CSKRFZlRTQjqNUF58QI
qq++XvuH19r+dcQ8zCR3qtaiIQKMbYxKqGYRu+ksEGTh9Ja/jssa+8w0h55DQzVS
NrNRDpHbhUii45wxER+r7A2Ox4kwbcunHWwmr+29EfCLY4+hBJ4TdCuC0I0uJ5Sa
wa7sBMSgwfpgjJ64MGKeGUU0zbtJDRDupkGX75B537BXR9NK0lSOUKYKJXR+BLAu
F7fomoYkNy9/WD174iZSgK84ydG9mh+jt122xNpqC77d0JyY+jeTIwzyuR3Y5QEH
q8y+/pNYa3RnPot46/sBuaheApjW8Dmsn7YrFdPVVSgBjZ5uOmPVqRVNzCl6EF5Y
r6GlQeJdFu3u7OHtqSUqU5btCr/PZtnOvTcpAzj8lyuvcEOB+6qkmtmkIrPgkygf
o8Jzw4zSKwP8pjOkcgclpHVk47AWsYMTXb9giZGSBYCdDvB2ZnVX+Nbg5Fx3QRTh
whpwqpma3KpKTcMYFIKaxeoOT4iu7jw0ZPT/PLrQSx7KkFcfBFkGDiU4DC5HsXGv
EW412Yr5PM/cd0oL/7qbN2I4iVDXFCJoZURZh5SkbLkZCWKmwVPT7BKGghGBL9m1
XpADMaOjK1n0+zCBC3IR7oxhsyjcFirRmpFFqz2lutwdbOlvWtWAecm82h4RydOc
xEwBlDMODRJAJqa6yUS+8WtoDZB3RagjbxzbwU3bZoTQMX2rMEmgn/2H5knN3yaY
IrxzCpaVgACDSJkneu6ef0AXYrrpJspNj9aAu1xdwH5FCbUXxNfv1cECUc3xedjb
5kxRh3zY88d03E21M1qlHwWBBmn2F8Jm2LPltRiiXGoxpd3AJdyuwQ8o0czYTAd3
2tY/NqOS3MUSuaa6qqq9qwzF7QiE7/PBtLTxJGm5yvPa4/LumgL62lggwDGdFgeL
eg5AdQGgXZmWxrjXhRaymAFzE9m8pW6pzKhoJ0KnuaeE6SoX2WNsnyD82CWSetJ+
9Q22rgeeQjNCHdE9PEdH5K3UB2q+BYpXsNcE4wSyA6hnfSWJW1s9uDMg/yZkpQoi
s2/PfqNmJgY0Y8ZL0UKoeGgdWiWbXXh2tkXTzZ1olBJRzgtoBKr4vXjH6iI5vAOY
5bif/4xaCOZWQhUTKnBtvItDyLM9hOP04e3pPnUIpISfe+wgMQLjKpTpQqf4MOku
Wc29GLJlX8Nx7X4XX8YccvxZ6zd3GvpbFfQTKhTpyvW7TnFsn/7c+2l+Fcy2tCgn
v/mYPUgVABelxTsjoqAIO5x9OX/FNpOJOyv+iBzPOUpTFpMA5Rez5ru/0ehcnl2u
mecxLOK9BafqRyjm19jmRQlYEE+u158i27545x8oUEgoKri61vVv/TDPxw2/lDH/
hH/EsLawadb/8aF+t1v07/jJythjtDIChMh/UzoyiasihhyP5D/8wBw1v1wHxjz0
D77Rsi6g9R8Cvd5WQ7ehVdJxJXehEwq5BBkW6CPB5kz5qb2GjD9UfkgqK7HUD2X9
0QXkrZoE7ixtDcmi7ZMO9wxL4JZQHZPEDTAdJzq+HHoYtsxFizbLOqwcuSE1XAk5
bYSeSbOYanBXJR4zajXBV90edT1oZ4VWo59TE92TXjVm9LVxRrJOrM3DiW9y0OqE
Z3BaAnzgJ7sWnuo7XQVY7Y9YlzX2216lbvvaaIOGKq4uMSXBJTuO2SXc6YLjCCQZ
jAd6UkR5MRH8+uqNQ3eqE50mo9sdCgj1TFN7ueuEkEpgxzzQ6SfnHa0SKEY1zraa
OBa1uO6VFrVVN0xrUqt/Gb9XZlxq+pRYNW3zzWiMwqvYy4qPOKXLmLWJEAR9P0jY
B3LUR7gKx5J0O75ihZ9H8valo2zBVp854ygiuDhl2kQYxxj+nNN83fuTgPZLseuP
tVoNrl9QPzTayruRS7VHgnmgMkrTX/xrh8aZLFQWDV81fsnMD1Oa0tDovPhGFNip
fQaK3dk1AjFzh5qoQn5shXOE3NVYcBpmDzrA14x3mvUEIn1I/gZ4W686BjmN8tuL
tS50ybfz7SCzmXhxDqovsW7xbVjvgJUxy36Rkrc6MhY1ZyfUn4GBjH1W8jRB4UF9
zgph+uE+voyTMuVikkSJ/hCUpCBPqhP4JiybbJSWUvkzFYTp5d4KLFN6Afs3tNuf
FBMWKh8J3fneOkGTw2ufQv7MvUelwsy7LJZxHaZ4KVzSNLkWDqocf6zJ8d0eJbeA
zJ9HCRmwVWEppLZ1J4pfUmaBCg+yJDK+r1DkOH3hkGQduD0sdrYt9GgI6npbDJmK
Kf7x9xfzVS+l99stxRvu9sIRTtv1zVqGvm89shua2/TcRiotJntkRNbF2XWWpx4L
Zb/SGx58ysL1b6Tds/D3lMzWWb2MdPfANRkmXxjjKPFOKygDVbi8/MEKnS1AxhC9
RgfRaKc5g6ucOF1s5XhA23RdJjdYXz+3gKyNTpn5bzqPR08n72zao5LiRHwYSyp4
0fosUvRYHvt8rDKLi3F2Fc/4BhLr3XYT1D4UgaCSeM22OHR9veBh2gfQjPOZyzcs
jPfInzfmEWpz7HVM1CeVskwOu3foDVaohFyJFJgpD7gHP+3oNjmscq25F3P61unc
MAqutMtWVpJxPgi1GE8uXRQjjw+YwCPNhYu9YOCsa5A7fzObf+gLPtNIj5c2Dswa
fLUVsKaDEFIhsiSc3bFg5x+EK8ZnOoDXi1bZ0zk+u8Ur1p7IFcvCtjqQ/o2oE+sM
RVvR3ZoZMUy81cGFdGy9unpkntuWXKrI5FUzG5N2s3wlJGauU9gCuHJXJ5a5Ag0C
bxgYxZRSq+yZ6RLM/4UhLthOH358Xv9jiYE42r+s/r5iwqi9ynRbBwHUpNeeeyXl
Qfdf5ydfBiFOZ1yFr7qqNW8C/pEhz7OFBGvmEYvIbVqPvB/uQ7gVdBYRvwYlUjgB
EXXrQb7yunwT13cSXYDXcNwyDn9fgj01ELlq9yGZZdnyb97Kh9TNFGB9k6dYD/Rh
xIYpNLP3URteFN/umwjbE4JCJSPHnvjK7D3wea3rbMSE1oNIdtF8juc1LIbmqHIS
98z3jymQWHshU5e9KKcaIgFgrvudGZ/yQJ3PDBwuu6r5kbFmbbsb1wWUeZWA3A9s
dEm00cKeOTh04luTgutk7jQdaQzY1itcYqRn3yzXK0y/0/qu988+tv0FmIbYSSPD
jLkRvwYOBs1L6Ms8Y2UUWTI0qMZnHFZL+/L5l3YX2KRAJVU/Lo7hKAIKgqLq7bLA
z9Bfm8Otnp+1LIcj3oyGaBoYv4G/dcg2fO5xpo65++lQZKNHwY3NNClz6O8Tu2DO
rAQol5MkKDDhRI5vXRXFI3c8SO6/vJ8PV5VbhVUuXqFql1+qmJuRruME1HW4Q5Hy
+XjeyWhqCtZGmLPhfQ9Xg/SCQxbFLFVcsrMog+Xdc/+W3YoH3fQ4OJOAU9ucwX6u
g5mgByFGtxEwuUj9cRzeF8d9+DOTO9ODATadk9eD9jX/f7tg3QOSzfiL2gRrZnc0
4/iCYUQW5bG3to1A8pxbbaqFscGKK7Eflx/xCPwVr5OlVGRTk64itXzmeNwtrqjs
vJHBkeJRfLGWmgFiYd7MPOIRN/c93WaVAOTgxaQcHmf/q94tBKuxpOy9MaVDc0Nc
mRYRhlM+xsMFODWgp9SUuYjVKGsel+CI1KoFcAHLwh+/f9U4NAaICn4zoJ/bLPMg
hn71u4nSp4b52vQxl52vtlkswSTzypqNoNfeStYehng2+BJyP2yPR1VZdTTwJpgY
aArz5lkeBdQGbKEm2SHXL0S/sPkB2OuKuvRAydw0NzngkwYDxZQwMLDfQDmyW6wW
GPcPLiyMgjFbTrtGtAny6Z1smYx/0w/5Vvb5Ll1o7/FsAcVd1EPioNsATdj2Y4wi
WWKFJzb6Vrpsap97CfV2PIdCaXHe11rQsU0MdMNf2I/OBXHk2Y2VCoza6j9V338B
fkVUXZ1PmNcaJpBkuHELvJaAyFg6RdDMAwgjpJKBmeR0Fb//6ZNSOuqrvTrt1F4u
KeY/1v1btggZ6eAfqFXoN31grSfuSzfjFzK9ArJqEttEDFHQTagzUSeRu2GfgnME
wWvLttgcLXQqunjHqgfdeqhaykJEM+8h3PvI4tszUOqzn6YkL3WLoeChGOO2lC8h
VOi/5XjlYGdvCx9nHYt7unFu6sZtTP15FQVI3WjUPtMHeQQsDAiT1m+QdDqYMqEo
SJjZKfosOBvUUvvJFX/9uDbVvfBuaLNUUwFI4mdBkBhJtaSUi4a36+zwLO6Oi3vB
OqADGRT9/mpqywsabgMHSfGZ+Cxbicbkhw9EPSOfPurbAuzc0+kAK4UqQ7kHpd6q
P0sh9whPiiJAimiWOPErjgeaCeefE6RoJ8VG5cvbyu+tJmBh+hnkshcCQdROFUtx
XzD86vOWfhUfzess2OJhCsnogle0IfnSkI8msHBt4XsdjuvNgdkIkUpu7bZukldh
6Pzb3BpsjtLDQdpFm7hIYNEK/HNUUZSO7gE4mvRoTTAIM4Hy1f24vXB3uTE87fRM
lxUPN4cXbcayLaNYxZQDQaLdBxCZaMLz2Rd3zoJ/dXZSy+r/2Ah9nAI+63I8Yauo
gisPZh75RKbs4IE0aZkFuWBc/YoTef+jrXuQlNMIWZigTqKV72tBG74IrGJPwJcT
vX3Avm1sBrSItbe95fDM79w/Q1Yh66asy731Snr5EgSka7D1ds+SjSfzvH+c6GgL
UxH1P5fr0IUKmiXFVvTds+rEu05bJACriYOyPJjZ0B0rKKc5ABLj/Pa/m7rguliu
4eDCzmdsfwvBpihH7UVDEVV4TR9rf2TUZVuPN42b8sXAzVkWsyUkXm4zlrcCgJIG
ZTHs5tWN1hVbErVkNv9bQ1w1Gz5DjP/CkZmHs3Urd+ULBkwwAAr6ccjsLYPUcO97
c4vq94eWYjE4OosM5+Sbla3cDspsmGFSJ0kTMGL0IbISXFi4hfzN3Ap6Ytxwgwkf
xyEvk5KNd5t8EZyJYiiIXZm7wI8aRU0Gh2uv1GUfacb4+65Chy9YmlFExkC2xOvd
aSR1wRG/RG8STVQo6Kt2w9taKSqx/mR7moq9UmsPzEzBBLqfSyXqY2fKk3MpSraK
TfTQkTXqKLLKR0Myshw4PS4+f4m0WQ4QhkeRrYesBeWmIG4uTlo3PpMmLi8vwwHl
Khf/+BCdp6zHLjJUhXByDjnsXHXo5nSCzZkZE99esykzgSEZDX2gT4jClLH7LQA8
TPl/DC7G/3RKhYYGbbvo4gCC2pt47nIfb1Bl5/TktHi2bNedpvPqXnj/2wjl1H5L
Fev0kQaHIUKUmENhWCp5toEjMHC5TrjxwkcKLW453FfGtugk+ddS1bmXQuzlQJmV
m4Z53CvfMn1BbMoyWpeYrOOPRr87AZBYYy9FhREyKiGTpwfhxueYYIDkdttgNCfN
ZVVODdNrDMiyRLVjXVjjVr7LOy13t2KNSV2VsNCu+ObZIWHjdqK1m5cclrGCLZk3
ThKIK8v+zH8j3pchSPfaKXGt0koUk1UNiiWE/d3RpIjQlnGi9JjXSwq0+Ttir34F
FO3F/rexy2BwvxgvH8Glr2NRBS7CvfZklfnh5FlGlcdqNf4wfRWM4K8cxhGpDdmh
5v8UtwU29nHz7RbKRyJ+uQ5Tk7bmU2uY+6iKEqXmFEKmKuDg6gXD+vtVzLDCjI71
ygoOdlDQxX0oheXFdA121dBhbrHGmoJeOFb4qsIGDeWpnf+Zjxj4eSRbusQrcl7J
t1A3zIBUxAdoJMb8xixgFKec9BDC4bq40xT/863hQ/uwhVGFlsuNYZ/rdkJIBKs7
tS8kx+Pa1nFGJQIwPMBLBn+sqXJfiS8fnTXzwcnBwVCYkmxhQxjcE7pWhB4U8fKJ
C529+xtC8112hkxVeFpOjkpK7KScv6H7p02nEE2mZKe/13QWr9MhUSW8WoFc38OS
a4iGRHkspsgFrVef1VYDV3vvpEyFB6e0RjZouvpYYzxfNmrmgNd6CLLfp9ZLcip4
lXkTpTnsYWcyfftMM4rVZi8plcYynNfdwQbaSdjz0rJGtPIM2maqsPt2DgWatIH3
utQjbq5GlZd2EX37loMNFJYh8ot9WWhZirJLFdavQd2ZDExrk0NCDV5NJsmF7O3z
3cho8HVXwAs3wY7mT/ppMCZrlG1Xt48tiGQ0xd4ecid5SGvuBRuPZn+Dfdlvgb5o
WvMQjDsMXUY0rSHTxpqP4nlbZS+FHcRCgAx3r6MvZS22pip1edZvyPX5iXmi+Kbx
VHgvXTmLnyDAdIWNkjpYFm4BOugIJQHi/2NVe1zfA80VnMsDuR8Z+mC4d+iI5CJZ
TAXejbhfcbGyTwIFYVMCPqbSEtFbqAPeFC12lqJkHp43akmLqa2KNve+GtxzTtuB
F+04Hs+/CuOBjK+sReisUpl8QYOdDueR+vOpemLJnG5THfDzcE0s7cmbPqOjH9Mt
7lyoppfrZI+J9MClkQfXexstu3ZHcuzya4ywRFMe9f+/dvd+uiVU1IxnlgwsNDYg
nG6oKzN+xguZuNs7DB0XhauFVBrkJce98V0SfYh0zt54rDMA5rU/zyyW+rL2iPFy
OHeucE971O+zszFwyU8SjS8orYHvD2lE4lKrdMIqWN7id9lZGFYp3ktMUSE/i6QY
+WWBgoIQyxo5O9RhsM/ChWVZXhzCTDPyxHemlvog5gVijyfsR4BExYbBS1T2nD2w
qvxCmdZo7DIEK+AKInBnWystcH/p6Jc9mQ17VfWQHVDZlZeQkgdFLMyv+mOQ9n+k
s14ssyXFhuI5vk2X70E3FYSbfAW/GMi5Mxsuj3+Qx7h7dKUPxSvnA2/L+27FfJj8
sEavnkl4jYoQ4cmp52Pe/8m5/a7b0nnoOA7f//QhLhybGSJgkHls8PHPvYHhP4GN
z4zHB16kAqQubLVJuVcmj6f7YrwIxN28YeW1v59MwMOz8NY/xGiet880D3OP8UiA
delj/pZpBW70DLIWAX03wc1BMwsRvX4WQCMMJZpshGmtjHvj5kUmDt66MQllVTeE
Dfk6+fRDfY3aYyqUSIIeVT9nEpDkz8XZh32ed3Q4v3ygDTLnqkjaUsTB5Q2eFc29
P5id6MGRo9lL9+qVGytZOq6PORGdkzKTMCw1xLNv2xyEVYq17G7Ah3mXuaFH0BN9
bkK3wdLDlURh19YxoooAK9xGqekRjVUrQYzijS/IQkpYMiOtyZMKhNEjHeSW/FPk
o/ifhuHi8DVM/WBgWfWqXyF1airu8YCuCIEmerEl2/M8r2HJ1KBtlhtvAl9a9jQj
FVIHxBD2hUJSdK/Wzuu0xkSXgyqDdotEcSDQST1rH09yUdDPihsIX9l5n7N3P5B8
pE9RsXoCApU7F0HF0EIQy5DGmKb99YMjjpfZVykJm4s1CYutsLgePUKo3NmIzWyc
U93vcqy5kYXKBmkE1Ek2p5Q+gJeKXu+8HtY4AO3LvLxN60So6l+qU4TWdXNCQQeK
DRSIQrvUPqsmR0xNlbvX6lg7gUNw+Wz+kBMN2MkGAXVauOPIg1Q8wMsY4JHgyaf2
7kcWW2S+5pr+nphInnXcTS6CE1on/sp8fgljYymV9/pJYVuZ6GmeFdNr/GGdhFCI
GK+EiNq8xUFsATSIedYZ7J5DoyfptkTI/kXErFfVF5ZBiYmdne9GF4itusFhNZRt
bIOW5BPFI9EPx6aNMvDjuRtz8XcygagYOSDv1EasUA3iurGbM4x/xlX6IkngUiQl
sE9pcF5r6DreJuPG81Tcriop89cXN2zehP6AAlCL/z4v2DTmfZ0RgplMflC7htVb
QKw14XPDDaNWEVYMVoBBHXfeb7jDJkejVZJ0Bznnenv2lnGBV/envHNedso+6E6p
vcnTslpK6Nw5ZtEWkEFM2oQN68VyTyN0Hq4mizIQwPWw1IZD8XG2YgQGgbARJZuA
9l/72+RGrfW1Vr6ZrPD43vVjIFpWt55j6/zin266jDfYC4PDOOPDR2Su/pAfd1tb
4QjOkIBOQOZGsORN7wcv1kjY0go7JMPf99wpNwONrmqEUEDeqIuYj9oNiR59PvoT
SSe8H6rwq9ID1B/ve4OwG0h2z2Bwr3xBOLITn+xC3T/btCI/rUS3E0w9SMw1jxKU
bamRjvliK866GjrDuaJIlWo1voWWFACNIOHrnuZfh+B0x/O8QNpFaLkmIR7aO8US
MIH4YTBPbiFzZojhLuQgXblaEsp7p7paZdSlkFrD0gd1eJLbykrVW0BQFhuZchom
8GW+ddMW4GJwvTo7q5AZcBDu6fb8UmQr8yfYOsyPBFzkANHcUakNKL35uAaKkOxc
jVDTI0uS1Yg02XRGI6UDQWMiCkqzxMMHuLkVHJwGsFZOOslJ2BL6C/V+CYgscUN2
TpMJS7Tg/HvF28nMFiFo1vuPTpta+x1JvULeIPUBwqwAFoMnd+sfjTbbGhcw48l5
0RfNhvZRwJcpt2w+iE7ssMBkbXPOs7og6NDVwOUDOlHaKij2l2auBuNBNDq5RHKe
Yds3qmCncy+m2zcfrTVu05eKjp66nKAM3ZaAA462c8ezfm9NhmpDTAcILuRnPbMO
C/EmvN/QPxCXuyBM7ZkvrbjenpzgvLFy77Yb6FNBhS37nC68OKaf885+PZEjE/yS
3Szr9fGDW+2+jWZmJzK31Xbw5RKGowuv4Rc69op8jHDVIT//9ec+OdAPsWZda0XA
XxKDn1O41oXCAanlR1ZnKWe+akeGe/PIsYaus3rKyHLVMotwETjRSXyylvUVz0oR
nCxgNR08IQYJUNbaZCQ5ONKmMx3S/BuEoHVZoZ8XbC/1ESipkk9UY0G9s+1HJs6X
DXwtJc2ozkj7J/hh8MlqiJVG+GqjS+DeQ1iFduwm0ZnzZMr31lSVdmcnWKUciCO/
5FHDbUf+97bmoXh7LJmUhSNKhBOm+hlCbg9pMJOR/Qwf61ZQPsap3lJJ9ScAhv/T
1GslrczETHR/l8RiQIObFPHfIiMftX0o91aGyV8yke4MVto9SjwvYeUaIdnK3Zhb
F8aEsrXrYIOdfsfAm+65rKH/4+EkDryeSFPG22qgotrkwv5h+Bm3moMMMH8LuN/E
qaLXgfaexi1hRX6HMbtScTrTNWHwuHv40wrW/YKdQnPDO6Lx9NTEMJ4q4+vmyNfj
1Veby6Mf4paaQroeuw9TXmNmdKqC+1YAvejeQVmE7RomLQ+itbFedzlRBDuKXSPO
rSbMj6s2fiw90YxBuQ2dW/2KrKZhOEHlqld5ajhl/2CxNWKuBj0Z5opc0HhQKEnI
9wT+0enDq3SvDk5vcVrsYl1f7OvsOvdBm2FOVKxpCrOnLUq0ShRkWtbzXuKOYczK
phSNyTtIPz8ym8z6DzJxxfrHvQqeoMDmDEVR0WBIDABTBjGIWskkCT8gZfkzaNtc
JKznk8s+85CtMSHfan1l6zpf3qXUi7f/k6KCmw6fAlpj8r73XBZVyq9VgcNvOj6P
18ViYowWgCAEARJbk/e5GB5WhBXJtILO/id9e9L3iWmqrK/oVGzqQ54attlFS11H
cAeicceEwei3/OwQPI0bAZ+udjPrRCfdzlOkN4Z3BHROXajT1SGPXVCdpx/0WuNa
hDjH7moBqmVloroULdvq2cfYabDyKlD9uv37t8Rdz3Q9tSgH3JBiMun6+OkLhkR8
PJcUNzlbLsWQ7P3rkrTSM7pcecilLfxNFPSCQErk4NIwvfwHb0y0aOdCBEje47I+
8tIzH5krRprNB8bNDX6/8J3oYGAeORv+IYU+hnG5sKdE26fx/VWbMMIH3PzZo6dv
BAau3GGnuUPXVAJQrCc+AnVDNdqJ9NodYCCAheDSo6Z4hkUXeagBssY49F/jEYhk
rLmPHbJaGpfZAr0DpHw9Q/pg2oVn7n3XtRruPMFTPmx5APVNsfXSEWJovcvt3QFn
WM7yo6JtkicsSBmUzDgeg389AUJmup2APuiLNK6Qng04boR9m3IS/LY3qkeXzxyF
awygPA/XZFpwuqAI4duO4erL4pl8RBm0byGwKdhboz+LuCsVzhQ+lg4F4TjzgIG/
yZSM+bnb+gkEfIlCPycwhsL/O0ZipzRuWY+ons0bnyfRFOLr6a7iSWW9o0KsePwU
3GO77VK9zAaI6M7ozX6y2ygjpYIjhxe0DrlYBt71lGtwDxH5A7kK78uA4aOdROtF
sfdLp0GdbhTJHFz+zqdzq+LUKChVzpK9EbdczCdMFVM4o0+CXaMe8i45iR/ckQ8v
FygmnAgBilpODqbAiBp6vWDbmKN392lcZjEalBTrtSYPPrQWxHmGtH5QipUAYh1y
6Vz9Z5I4SxUL4Uo5AX9WUsJM9bAAZYo4dksTPJaJBNxIYtH+pbMnbdl0ehJ1u0c4
P5j1Ht2reMmUHMf1NyEzCaMz2IpCa/ekijyQ0YDyWFyrfb5JqocjkrgI/mhsL021
S194gKbDYWxG1oDi1iO2TrKZVf/y41N81BH81QQp27yC0p3Br2ipBW46ii2wHqLG
cuv1qyVt0eTUHVv3HG7VcQ1K2uQIDh355S7G1HsUqJjjmulT/clbOwjx6RUzQoVV
a0iLtwKNdjUbCUGACgNTgzikRRyQ6nJr3aN9HQUaXDOzPpcAMhswk2wSlKWOcJuF
Gjsbb/bnYZ6moJXvo79eKRlqcuyKuQH6DlTnFmo4t3Ox3g9/6eGWTnpI/BfSEkzn
+AgxhH1E83IFI8cGmPanMAOCEpQjk1OISgo2GdqvLKwPlfg0G2yG3bJoiLZaYiQr
fTSKfBSH8kh9nPyq7a3eFBVuhfeyvNSctIQI8v0HKw6FPsPhINdPCrhsyAm6Aee0
f8wvP+mcCyeJslb04X5iH7mf2e6jUVzh7ffqXZgXn0Nl69zyZqZkfpxTttxAntZy
vr6Ib0aluEngUCM4KxwoBkCGTWQjgI8Pe3wHPQ0Uckp4zeiyku1LmXDxxSQ6WP5w
bayTkDltFkD+BLjwnasGnD8pIF7ncOQ6WAmgDiIMkT4H61/5sGSwXBvHms0jDkmF
C/NBITcHd2iLa0lRnyyvwi4WJD2FBkpegey2QmMu6hApAJSOk+UrmVy/JbQ4yOyN
6WHb85w/X1NTVgzC4zKeQqtZj5ej3oj/E3Ph2lo6Qg5Td5oQX/VLyrN1MoI5wEzb
rAKlDnPwYc7x311d8d/aw2sffIvVBq3kS/2s6k+r2t68d7+qoIqnZN5Q0yYn3o26
18akLSqnceaBzwaTujAgfFCovRK8MZDUoPuQh1k31QBhBqLop9LmtpTcY6iHa17P
9wTJCmQKl1p6kVUqcKmPa3NsCCO5zfuXtVwQtF6ZyWOMvHo1rsICs32megMGATOC
N8oSlc+n78fbbeYqxORSoUdyszvYSh6O5F5gKRUcvJvwb37tj+06DPem3fwsiuc4
HR3wrnhMs2uL88z2IqieQyQm/ddFMxX86toiDXay1SQPLD0jhi30Oru32SAVxSAR
4ByLRJ0SormQXh4rp6EqdVQVDNgecyCUkvPnUvY5V6xJbYKLTT3jabDbQS4uyy7p
XhEk6UAq6RCmNyWLdKSryDmRCQlKOaEdIvD+QoPrt5YhMELtcqhsSYLOtRA2Uqyu
RJk0OPFi54ETtDTGEElxSMkMJzcG5qlQEDDPvN++N7grBYKqZCOh2tfeZaDDYXYn
9bGXA0fjvN5m5lMldIVLBjkqiZot9RaclpTPHZD7IkmKWP3mxaSI7JQ+CvBOgGQF
48HDTG7yhdTFZpDMU0E2Q1NJzXZt8EjX/cI7uKpWRPqzPyzCGX8JVXyva9k/7WJl
fPcI5LpBsJsdIRB6Lk9W5ON3xa4z3u8+WHqGJZSiI194KBruQwwKjF52hOxaWXPv
HtQTldcIFcon1hY+5MckRr5uBclf+Xxs2porZQJjA5+wl9sRx1VaC0h3+V3PUCcf
FIgFnQ2FtYDatQJDY0DwE30FqICH8yXNF1zOs1JDNeu1lVG0IdUxNPd9HwrvPazb
xpjJcO15EFqDirMxiOMm51XG3HyqasFyp1u7RkBrvcQWlOKaVkmacZxbWr60Wan7
fbcL9oSqbogfctNSvGEzHmoZQ+JVd2BvzjpT0W05cFYh3klL4tUI25pJqopI7XfD
n2VhKK7to/ZUGKIUPnSeMwSIhjd6wTT0Mn6JDQemZVM+OsxPUw23wsgEMeHhuu4s
C4BGtTuC9ztAOHbEa8knsGybsZa6G6+Yxzy2+tT8AMc2le60fILZ2MinjTdTb+42
+8H141HCFacOu6vCpCBu4c6Y2gUXDzxP+0pkkfbOj1RiHq9xr3ZGBmv7tLS9/c/R
u5wfjShHFegLoGoXYpiUNiVj92fflde0HInVIATir5RjGZ10DDR/ld2KX2Y5u9kQ
QOG07n+m7VpleHzsvszmUP9PSkY+qUIu8NBrhIVh2cSZFj/OlcFU44pQqUzwiJH1
vJ0Mq8XGyLB1AsHGsW3Vfu5YMFWEaQZsBBgEF97QGHmchgVxRKRLcAn1fGZ2yrce
IHLaEaYMSD2jAbR3ypZkz/N4uZnLa9GLhFAeNZFcAKAy3ivvTkw+ZEWXW10weRa3
Pqzb41siZPSzRHRVObDpVL3ZzrlW5cXqfbT4XtlqMM+FtkT5lpEFxZnYWa9pqiH6
krzUg8ozhq3GzQybTFjyot6Nv0hdLDCw8BFtruTbu3figAHs0fyJ/Su071Bp0Qri
ynayUrLEaOjjtE8Or9sCZhGIcZJef5BMHSWcyjIrDvUyH2yKYZzgS+oDc1dpotTD
MyJjiYngvaH+0kPw5pPUcDFMK/Gf+ZnNMMyDGDtigET6B1zSvn2UoIdqR5zyDrLE
76XJcwiaKo91k3PQC0TO2SbO5e/DKtnRngweu4d+nyj29X3UBXhQ1UnVNukI2rgC
iiZjpEW4IuZvxfeMDAmutNx8YBwntGPYiUcDapolHU2LxmaikJIAXJZBxfbK3jMl
1uE5/NbsPDYP9BFeEu8is6xMJd64KjtoY2TlIsp/T8+GWH+5B2dvvvjP0ojsjfgN
e6+QgEAVB8B6ngMBk/2ZDAOFmvMd00AqEzkdOBWn6PdxdGiAol1iYKOK8hm5lOdz
AY1OeMzb8ACwoiTxhkJA/VBPesPAAvGKUjHv6cLkWE3vmywbbn9aeVpPAOVmGB6k
yNe9//q9FXgurBs0nvvG9TaxtQgJZ11nEy76CPU8ePa0AAoSYyxJUdXlzE2b+itO
5OElvk8kaKfWPTXmU7xs6tp+tD40LHcltb/1K7orabbRqGnogD2+V/Mcc61oturs
KQW5/U1hdnBq2qaHaSWF3xtFBcqVI3hbNGAS0z0LxsqmNt3Cm2YC8qu/7KvJxlx3
Pg1LALKzsctYbEO2XWCtoh1P2H+ng/Qa+I/IzlaE/bx0zaRXmOtJHH1rBmggMmYm
63DeoZsanSq7/QA7XxBus95s2l6rqBy8z88z+67sjK7rXS7ST/cv3xV0Ypu7UGBW
jzzvFFjaf9SK6XjJEkBK46e5ticYGqFIRgFiJnrb/mlbK8UD3gmx7HEhE92o7df7
1HKCjx57eGzRSxeJ0mPpYFKUyO2K+W6dAvJzLza572YcMd4WYR44azq/GoOpKhMy
pGjxTQLvYtL0+ejDJ9LVM/hTpAKbYGNX4IPu7iFDj27Alh/KfTx7rdAylJRBpip8
8sK2Ubth/vkQwcPAz2a0dz0HW+1s8Ow0v5qWJbc5hdjiMsBkATuq4gUl/vDCjGTg
d5L40tGFSwpruFe4ayTmItROCiHhSfcB/HHS5JHj7PmXJKjMforg3mWPOhMTf9YP
1ICAT1vD7i0A71Znz2TLK7qEDK8jGn7D0JnQ64H08DMXCo0YMHVm8nnj+guVmpR6
A8e2sS6NSyFev3dJmH7+uRRhXghqVEZBkodsTViPIxMdaeNIxEIAmY0/aJykL1Um
JD3jxdiao0KeJGY3dILQ6E+wc0JNEPbDkYXVO4K9jBy5nNL+L+fCzTSJtzGB9Nf2
iieWOZWQkJeSzqYq184WutqC7sUvpwSW4aJgK7Tn7alulX26zG+q6owpqmoTMzxc
ma4CVflwbF43+J4GXYswd/yeHDH4gWm5mhweRAwAxR7gxs+yvRqtzEH0Q6t33YZe
QwO0goxi3ZxhY8PdNvRFLoEUVEZ4T2AABxY7TbfXr/ZwGwVIoVg52LmvlAHmGTGI
HK4hzB32ZxLCtbmLsfRA+/QEwiYlHxc3jVSUX7ddnGYMN2C+wSLO69yI0s1ML3Ri
Z2P8DRK09MK7sosoPJaenDKKU+X/KWl3k4DYrNKxtRy2NVnjFsJr7DugvCpJSSlL
SuvWoUEeI6eGVW1mIy7snX4ctuE1CiK/GsPLktm0A5Fxk8n22ylnxkBrdX/7KSZG
7V4cyZIOGRR/51GPHjyh7Yuq1Zxrxan1by2uVyQixJc7uQabdSoBXXlDIlqJEHoc
iKTTUwIllAf2mPE4kntiffrmL+OnBqjHa1niOttoF1QQkBPkZtwx7A4720oySi2V
MKEjZsB29q3cI0I4YemQXB8XKOQ2udYb5QschpFXDQ+YUUF/u4ScgMNioN/cCOZe
1Yul/mQrLwQVBv3KU4gOSN7hc6hPrZcSv6cDvu5SvA0qb01Pccdrq+uGi8RSfb9V
R5U6WOPjnJkwKJCo5FzKeytvuto/aZjNQhOUejpHIY4RZr1h9BdBB1qsI6jz9SE9
0vmQghwV4DZlc8Sv5DM9Zmn2TL4lAWeNwCXpCW8tnN4SZ1lHyfxAm91iXFT19GBg
yFc3xVBPBnJCjZOHvRxIpdnrGjpuaZU2zFqYklvhtL9C9fB/EpHFHvHDSYhn3rkP
hQxcnDm/Y5n8bCXaJ5FJuMZp8CpaOLJ3MLyc1PjG0Fewt1HiugQ4SExKA6YKAy//
+26VyGNqhcIHgkNxAkTpQmaIF1EEhGPWh88bTmEznFfOKKIgqskaN2evN4nRD06A
vH8Jfx/xPeLAJ6JlarhZbHFBO2NyV3oUxCgNqrzd94eZXBsjFZwiRo17AN/T0NL0
pPnBFXK9o+8UxWtxLxYhDZI1eg8fo4lMJpUD+0ne89yRpamx3D4rhv54bX3xAolj
tM53XAjFH9OcYRH4Hiw5JO5qVXBsMi3/HjFSO1oz56UgURE/jxMQlLr3uBwy37sD
wfYBybVPLva962fGf99lqEDCeKiZ8+nU0iTH8iXTSdpuhTAm7gcO5mMt0op9Wv0G
ocgHskpkMAfI9OJb6W+UcGw+WG1JCG3jDk5YVkY0j35WBP+Zbg8X9IsKpGRQbuTG
aZzPujNE/hXYtesWLhc7GPmzjVzZW2otctyRSJhvn7NUoQYT7d/20V02G/6mGVOk
n22p8ErQytF+SXsUO126pdbSHLOfNgxVRtf49OKPebQl4PojFu2ArPBUxjxcV+Aw
Odmu9K81scKhl0St1Cq4F/dw8UwNpMZR1Er31ksihS34pDpbv8UoVy5U5Ht5T60S
o7nrh0PrndGzmIA3WZnZD7tcAl3okjzwokeRnBRn8wiDbnjatwPkcfel9ceVk/lM
CAcCA0PfQ9ELR1dNn4vEVi2VAEYM3HoncFMMC8V1n8P+yTtiBO/8Vb6Tpo2oYj96
NHN9E8uBYXr+YKNB9E1KIXo13/ZznZEFQ3RMSAJGFipYIu+X8/swzvua6+HKBEnj
qKgFdlQU2sRV0bGuSbRI4qyJyx1ZmnZ4vpyVqCRD4IrKumbpQU816t8jNxIwcjXZ
AenH8Xc2Pj13eC6QyYNo170zD7EzEkhEM5nbblytX9+fN5DknHx8pp2ezazWBkYy
ZRIWgSk4oXGLAHZsaxZnYxQErPpm4uNldAbO2YJAUJBpofk4ijo+4Z086sUsRxVA
muH6nRXG7sIRJ88GzDIWGCAWu5bg1rsSMqmgkgEBsFcFAXc5JB3rNcvYUQiCgqAt
FpGmRw/IDHQ+55qd0q1chCD3aezzmRfjQSohgIQrYgAy8J4fG51edjBQ60ZknKVq
2HjtTGKVv1tUoO/SXpCuL/YNSodYpfOIICMrV9YtKgF4xMPCimZ7ZGivSpNwhMa+
c4G++1KB7t1IPoML3N1jP+i1epkLq5aYVl1Bp/uGORrdWqh48NTaRZLC+JSEJYdV
TY4sNIgl4AWh3DW2P0D86OYl8wnxzfEtZ4zlkho++xko0eAbNOELfi06+8XQOrNf
x/fVG9KpwJXLqzc5rDS0v4ZSxa9Sz4od1CeL97T6DhaHSP7zMNBJDEt8505AdUCY
vmprMa6wttF4v4zkbreYbUoy01v8EXdVcb/PsBJlHvVQDuOyuPiOX7MxBISB+JLL
3FQyQRUtJHIJSVpPtTszdC7lvwaJ8AlkDuGo0/Vm4u8qyI22aL9MlMQAXm+NqUKv
1MT6SG47wMgqhftvztdQ9bpzPGrjaDrWy3f4j8vtX07pY//MNF1icY+LxIAIND7W
kD6coNEcQjN4YoHyRzVP2k1D8dZ99rAu/ZTLmJQ8NvapYEivYgLVMD5vrgQtxSWu
Ct/MOAugSfF6yuHaMB+RhYKwVZeeuJB/GG7/1T2gtHDRQu/MbG8elaN6XMKAebBs
acQFV1CJYCHMZX79DF0uGa8uhZvANOCvqKmNGkbm5qMGP3OoKIA9Cic22+BR38p3
CxumNi5mVuYWj8bWT3H4LQHffOyCbAfY4VBs6vn6HU3BPnsnQNxgt6wip8vicSZh
wNe2QVGc6xRSChs/U5DACe9QztvprbtdY+L1QZj/gyWwxQRsGcqPPf4FpEyUJgnu
oTsvV+iJR4xD1LtPedv1PUm5qTMso5J0+gazfyZIzXxLKuUKY9vghhUDUqgrFqHC
kgA/qaly7CRmag6DmX3Hzt7/cgXb9u8GjxVTpJ2BAaNbFvb2257K0JDOzKqNcCtW
mf36l5Z8tfRSNCpTn1cBkWHiQCAoPvLmf0vITSftzWM0YwWdCzCJxsmaSQ4MJGAF
T9qyrfmEpNjTaKHfEdk2L5UA6kUUXGErVAGDN4e9CcYxL+hJ8E9TRxtBcsAdCa3r
JkjZhriI4KhaWVL797ViPz37/mT5ENhKv5U3n7pkBeyTlqwWhn0vIndNXNYS6UxO
Iv0haF89XPlf0mFwMt90HHe6YdfdHcuf6IAJvcp1jlC/IGxJBuTlo0JwZjsCmqw/
j9CeEekoW9tpxDZuKmzZpdfuecpz0s1F01WdMg8awrp0n5WLRz2pHUKaXY6ZPO60
vN5juTKkUVIP5C+Es37qCj39NCK8l6+0k+GHpyIGUYEBU3SGaOBBKahzsxmWh486
DcTMrqEjMxrc6YgWiHsOqurm/HcvV4orOea5eqb//v+KG8Zew4ekcMqk+/6v2Yyx
VIOcpnCtEPQHoYJ6IeF4GHGphC95kuVqQ+LpJIE2N/mx2wJu0Hz3KHzMqS7t/kAW
8ujIrrHEQTt3XIa2yE2cPdMmjIvEHjUbgmckIxMK8dJKbiokDhI48UWmQC+jAIQB
HPgnMEm3uDAq9JVSa2nMCu9ecECv5yQZZNt8xl7NGzd1WWkDiXNKGAGVpPaExL1p
hcw0CPNPWu6Jq7+asP/N9xRvxCpXVwjg1Tdrt294LfO2IG2zC6QohoXTcdyAvXwG
oZeFyIK0ayb1NAHHrF1UmlnrGRRYGOwZ62hDcJcGTbRDMZGbIySgNu1l9Kn/1qwg
rntTxFZuJn7q+JjdT+dTEGdqltdZYWiKvdWrrLKfdqzpB17ETAPgYIt14IfuAmxu
iHjI9esC4ErDAbUSpzcX5eTjfjNjxGjUw3zroo7RmvGj8LBfJFtiv9op1ZE0wexe
MKbM6O9So6b+N2NUgk359U8CsC9oloU0WA+GTt8Gj0+u18YVszLdzgSTn3zJZLMZ
uggwfxPSv8riKNMOMB9fCckMzyiZzBAlSfJ1YaD+6Bj8m8dfpg5RSnOp8Ffh59vx
OAbiJGiE6Y7CU28ct5YAdEhOr6/JmUj7aYwIZ5ie0yNSGB1950zUYtmYkKvX8XCJ
SActpmLbHpqLzMHnExLX8NcdJ53kO3GlM5RcFEJR3FeGmlzG7SQudnX+HpC9q10u
NQb88aI5X7Jp33zBOlFFIFfVtUQyOuquKIbwE4DjMHORhPV4/LQaWBt4pLYIGIj6
WVopJ8m6Z7Y2oX6+YA/9FnH5NCiHYMK2/BXW879sjzC6vk1He2oWZZdDunzSSc8f
l9kplpLIqyRIiWJsIcv/Oxh0eV+KuXJC0JJC0+rkWOJQ1wve3cw5EFAxJ+T1PRM7
76vnyJF3go4BR2A/iHLn8KLnYEO5x+03ZM6mFPFOkRF7F1norIog0YDsCZfjfCZs
G8BVb+EyCsmr18r8JxwUv25AgTP+nJtcMwcwG++ssShfNNPBploaBKGNyuqliK64
0QkRlA0Vr7cbbL4P2jj9DfewjfI8LpaLJEnDAPkmBVvD1pU82v3LFZShrkjE87sK
lpKnIUF0M1H+8ZXXdiMqtCV8MlKvOooeK1EFqXAJz6UnMCTWEBQN+oNvarkUhOhb
csLZZarxSHUARpeUToGcUW8yIjngYLqAHwe0ksLj6e1gp420Xiy+bG/2nk5OBdP6
gVWkbBWYYdPnUNcgG4RB+F/6ZscXd9HQso0SNBbONDhlWhQVI7ynQREQPFNPd+SC
LQ6wJtQGdgJW2o00Cqq4K0yUeXZ3vlpDb/wFFzPu4xe+2dUoovdfatKh7V7fp4sB
zJVC1Ropqoj4HNH6MoFpugzIp/F9Tfcr6vypUEt0+bRoCQKMtqSeE7jR80vgBOuM
3fVp5AwFhaEOl1FcDJ323nnvP4y1zzmv/AuvTbP8iHUhJ19piUe5MHQs/2fAdPwI
LEISRF6Ff6lUX4YhrBZdHRMTXK+cnexAbR58+v4aG79BU+AxYaeWrRFPxCU4Kq3e
ZXeO0iXZtfjB556+9OosfBpwpSXlBOWW+EBKIPc1WKeIHrfjCoVmlPTwtiNmlRjp
UURhtFMDLH5jJ+fcqhW4TSG3p/pdX+p5r9H0gy1rclfLn0yak5AgiysbT8ySQ3bo
LaCRyCLHP4W11QJUh6tmKzw8TSaGLs/BI3qDgQ6oOz/Ro9NrFtRiOhJNktrx5z0K
VX9euVOVAK0kF9puwF7xNpv8oBDprply9HWBTrkSPn166ezU3iIuJnMTcxkimVUr
k8hfMUci66B3efb353EYMQpQh0V+f/7G8X4ZQ7qQ/NqFFHmevKaE1WVlMxswiVnv
zwz+MKJZnhSyFGq3yd28lH15Sm0wlyEm5LqnE32iPKM21ew1n+8QKRJiRT/TTVDQ
r2LDcZVhyorV1SC+y/QK/S5vALdnoYSrqpp5Bq41QMMeIlXdNpF1TDsX10jrdxNk
CsWO8tJ4Mo103zvXb6cZ/kOqn4GbsLkkXtFQpAFqnju3mlz2qxIWba3AuLjswGGS
yMTAZ4eQ2M56fXwQay+XOBfMTdTQf1WZqdN9IszJqwbhQ1TekwAyWr0hnzLt5sAg
542qs7DvVxeBcuGt51yRXoke3NArevE/XUHuhFENnAzQco6NzGeRnz883oCH2PsC
O6sB4if/TnBrOTl/RhfIgRcXSRYd46E8yuFqWHdga0/VMad15uAVZtHPsPbZ6eS2
+xFOBPTYQe7nIPnCW7Sr31+tPKm0i0n7eQb7645EhQ6fCwY8FKi8Ur/kcrjjQ6zn
ldG86wfsQXKVAUdzlBEtT4jXBIOjtiL5iiyXSO3vw93Dhs2W8mYth7pgAK0q34Tq
vxDbxzP8zMlEJ8n/rIOuM2xIPPBGKidrSEYrtX1ZdBxiaoAG1F81xnrHl4K6w4k3
MKQmZHhwTrM3ytbeFngW+hWSJCiCiJyffGcLTuIaUrdnX/LPDNzVRGvQY4wl0vAJ
na4SUQttapwsA8mwh3InBJUJarEs85qROcLFQ4dQE0SFSJmCX46KQp4G/g66grZc
ITuGPIAX6WvhiDZvDRpaSp7usui8u9lxdXB0vhyysy8TDOBxwTXrSZfbaI0q8rQ1
yeI1z2Fw8FeXjSDEOXD6ftY3mEyQm42aD7cJlToOM6ciYVJKR/fGhyWBnIdtyI+I
jw1U9cMV68JNv87OdzHDbrHniJ5LD59ro2Pn+khjDG2wlOHTOsfI9Tsximdglite
2j9XUb4js3N0BlUsql2O8qMzvp0SPfCt2qDyDdC2q8lr9QhPJDlryWC8z4CTqX2M
+TzcQFN9aRG8kJwDQi3cNRCrslXDUExcV+O1yUbLU4JFOrDsSgQkiIQvjeseOnQt
iyO5Tn3wYzmf/66eOZTD4WBYFWHdXAWmJCVLZjA74qxmVHe8rvJ2clVd4xO4bEuP
9QJFu7gRCGcS+Mdnu5QRLrY6zrJC66I9dBWovRZdVq486CmzMD8sSx8VcN4HKlWl
dITJjfhl0faiO5ADXcrlbUFXWkV0bWU2ZJ2ilRfblx1iMStr02RboSfpzePy2bBg
D9AdMn4QPjgrXO2kw5JVy4u/oNic/etyhJKeYp3ZEX4LaGtqkFCgZzNB/cifEnOJ
wtA88cDN+eetd0nzM+8hk2OclnW9fzE1KTsVPG/XbzssTMQy5DBn0GzQ2HSh6pHv
wYTNw/VzXKPesSfUThhVIpOOzxs9XiuxUyd+VzNpb/msl14+pcT4QYEoqn2XX28r
FIUqU/UKtldgCrqLP7tuWiZJ+0M7ZD91PBmHJCL+lvi4dIU8VFkR0z3NPHBQ8r1t
k7l0M+mDU8OnuN5quG9KV5x74uDiAMf3Hgpw9r1kG9MdHAAr4MGSYBOwkIbf2r4i
AziQrd5Gia1nZ653BrdDGMZ2FvZXRTWN3/cC9AVmKC55rdafdGw64Iryoj4BpKpu
Oebbg3MygoJx6bvbr6ahjiLEuevnIdzMtfhvFTGVHkVVXcfzOauLGbrp1Qs1GOgq
BRxutVj8z5WHwOFUXboYhW+H2r9n/uT6MpYWGhKjpKVc7VpGSWBwtnHhk/XuY4F6
QZfxaZzELAWVTthiKi/Llqk3AjNGSrVw+GTAcw1gmIt/JRHYFB+OU81D+L2TgUIN
9Dd1a7D+5sbq+6dGNYx3jN5mIk++j6T8HVJ2XiHqKms0tIOEWMYFJluU5l77fdOf
t91zcvuUxX67SRlzZ0PrZUoIyf8ouVIRRik7pBaYgVNbGkKJzgUhhhyE1pbJvH85
wPIcYN27/Fp9rhtftjGGyzeCf/Ncpyq4i/LIx3hdT4y5p2E5mK4JREtbBj2PgNbD
yqqaCjM6X34fop1XvBVL3RMOA8DtHZSVdjAezD/3qFNERn2FFoyMG9YK4i9g/Wx6
9JQTEvcvRsLrhVWK3Q37xGXWkcWOYdsldidJT9RUQPwNXNly529vgHplgLZbQ35z
fB49TIZSfW0bWBWPgQ3As0AWtAyusCveD6hY03pn4nVj1ZOImf/x5LhzaX1BQrE7
z8ACRXZ/PwmtxQ51r5yi0K1M5/d7nXT4ThV7+4QS3RKP6zQ1BwguGujxQHfSkxIH
Ch6+OKI/n516d+L2GQEUAgozgZbp7nPDdEHZXToP7wT/rhAP2Rt4bb1CwLIuvDVa
pPUX0kZtB3XG0V8Wt7+Ux87782AEpYT1inA+qTfJnlczkuhID4KlQGt82ssOt7NH
HzZN+kGmM2S1yK2/v2gODxFQsoudFpTkNFmeMvNtMBOlylSezrHo0TO0TPAyFsRD
7zdkcxpHIUFKZV0yetGObfQZ/fraH9NR3XTazFUu1qoLa1gIc5cET2xPFFZCeHZW
JRK/F1lcRmBcRlGPN5YFYInuWTockLwpkx9Y02pOKkvbBlP5r5Fz7npXg/d7eFNk
DoFC7i0erPqsVJxe+dmlwCn9zC7HV8AudZVoPBsysq+bxl90/QLAchA6LotsqZo1
HmFGC5Q5PRSYfeOsEQ6wnGZJtcdOjITnKvrK//WLLdRR/Onwdlxhp2VcjfhRxWFm
CyKp4iqaG2nROlKBCZ4oNDMthEw9WnePJlyq0fhsDjz+Rs3eCqjNasGgSBCZ3oXx
ngoPaqzJghF3mHJgrdb0bKEoZkRvU2BWcQ/Zx7D4c0e91pYOe4bctYJRCw0/oDlN
xH01Ync1qbmtHD2CcjgjynVSG1W2H7HiYyNt+haMT8b+taSoJXSo6sY0tnsHMtK1
WE0vcyJnCZIMBiS/fncGRZ+bC9BPdAm7j62gs6m7q2jvovQEJFum2SEZxcFOBRmR
HvhJZ+5HZul9qCIrhJrV3zK3WAlxWRYC/HAYHG33pGYy/NnJXHgESiUHpbpBUud+
4tZqFiXNssKwvBqf9s2pKW5kk+bCmV3EyTPBP6Xh4CZEgGonJicH/XikjNqYYSev
niIqm3bAMEGAtacOtGsS6iVx/R2337Ms87X1N9c1aoxNdGXcCfgzrGBDfHqFzujm
+/+sXP4nWYGO+IFF9aYVndO1xaphIwTiFe3MPdpNWHhIU/1loVgznHEr5n63eibx
gzy3G2nDamuj+8ax6Rjyz0+aothpfYdoYohFciVN308fJe1Zj3AiINFN74EPgmwF
aKhSzAnVaKs8gVd0R4/XszUVhs+ZOJ/PfbeqA3IqamwcEP+F2qvV4YaYWHUcH89c
N7RGvQy5ilsXZqh3pkuOvcsnIwoBeF87vluJwjiasgBxWimQWl9gk/v/7rKOC6xo
DzLqS/P2X4qo75YKBiD4ygPgW4uyk2flxmFl7ik8ugUsR1oLEAYFvv0Gcfdqm0DH
la50ZAwJB9RjnlMHIRJ8DwAuL1qhmekeYQfh0DMd1DWvOlQB9guO21IaoSo/2/Uh
O72CTJNLGO8ikYxC5S4rizjxPgpBG+AXXme4aBW3qACmkNYc5bVXxkoBlpl8AhZG
glizSSTBzIGF3gP0Dddq4tno0C5ld5hHkGxtyDo+FDZ/IAisEBUuITN0oP5DQPpu
ba3ypji8uQxQ7Ag7ttlW1ySi6c+JirTZVdSObpCQDZkC4H2r1hmod6po4s1iDPP8
D/3/JV2jVPLIAuRsFMLRDY1JEfYP4UiDAmf9l6fcNKT646uIG7CvI1gRQZVmJatQ
dygrKTJGp3WdreJUdg4E9MoRWILOJ5S1yzac5WyGObVRpQi5P47sv4soYHbaou/Y
soU1aQHOXgEQGtV3NX8TCu/I7bjLg7o98n//MHlE6ir2ejbMjmHPPUsozZlez7PT
ArxSyj3YyqCi/PRzu22+8QHuxZjue5t6BdMfCA4y2fxkzUiIMgS9LIkmBhvQ8zbR
rj1Gv+UF0lx/EROnPqp7dQQVfBPaFVw9lYyyj2k/5vya0YbQqM0pIFYahM/Su0Tv
s0t8C0znIPWTLPWP4DJ94+bjiJqF+1m5iVgkWCGVMDN+DUj/D/NkG/Nd3YCrmgQ5
29e+BPTh+rJreFrb3bcEFqI3KkmyXaw/n3FtuAv06R7IQ38kAnKvY1Aq4OvUyvs2
jQxl1Jn+FXpOxEoyCeRWJ5Oo4vYh54lipsAaQcjDxHRRxEn0JjliF/t7or+dI6Ju
7VyT8r4aI3rgh5Z1KPqMnSGpJ2QqMyktHf0CRFERjz7MFFf129rD6QhxfNXUsSnQ
POxor+RW0uM/UxoPFHpfcBgpHq990wj/LYGHD/2T9s90U0ZaxQgUHLwi0bziJZrM
tne0ZDKxNDKat7rhKoXccaoPe2vscQaPn8THJPlMkBULoc+H0JgppKgByFUbpIQA
wNa3ex8BRTbMikelNMcdmS3NEJSsFAkz5b5GWU7keXLVjFsz14TBslhoZyyltVzs
EfrcTGYe6odxYT3W+HP+aO3uyQZfs/G0gmLxYHjUh7EuJQGI70shFyxEYtTZOUtt
oFdPyCBZ646nITCYFrTE9gdUG4BR3ECBJfN7jXAZ1xTHdXxEQ9pcIbXJqhzmu9ic
6gox0Ca9NJHuAkcs2GZ0FR0lt4yZzYelf4viuY70p/Efmdz5wxVsH0pOjKMElWyn
H3kbSXoL4RAG4AYN9RazG1G9XfuQFddeohIaiNgvzflx8j42Tby96CZTL8IDWQoo
ISR9e6QfPBtN8KTdQ1j7Y4qhDzcPyiPWuov63fH4+cKRXvjaHsOrcR3gvIO+xvhX
l8hAauoK6amsvS3KCsZ/Neou290Mx2ArOYxC4/a3MRzavP+S51XQEzQBZk09oMoY
DyXWrSrq4bprODmF+DbhtFRf7SdAU49Iw7KKGRbggqrR6ZHPZqgfbqKN2wCYU+RK
fSGhaimcJ9l+AXOdOEkCGNHXGoYmWwZ5WHCzYP4MTXjGN+1CNEu/vHcWOoSgfI9b
y+lcYYNPCyDn1AjtIstq7bYU5cAQFvGUUtBkD4ocYMUHN9YR5J1I6tdBdWPn721j
/JccKYGufMl2ob4kGWOBangZyNmXQHiexrnScSg1KCCUHlOCOdhX17zIMeiSkrcA
9x4mJo6rhqUOVsZ6IHnzcEWQsNVGG7ijaS57lh+GtvKg/nlvT7/Xc3IUg3tEVMit
Nb3e6hE2RoK82x8m0m34dF8XjYRiOX1BzfH+63a8TdRDy6sq+/6iR9zZ3ZubyjIx
mC21x0+nQlB+N5qcNnOm+1izBHKUFzsnTzoCrH0UMkTVWSXvV6eFNIPGrDQbZf2v
pf5oKwlLv+HLIOsNyByAhVhG7i7rk7hC7VUnLLQ7IkTkPR/B4bq6gsIkbGYitcfO
qYF9wGXxa5VwCbHExuc7It5x+deIsUcGqkmgOcsW1Lmt1lpBwJ12Hy6WUmU70kCM
yPdu0i2FTaJ1Fa0T9QQQCKWrqlh6+uvT5YvLNhGZ2t5TmsLbvtRD9IBnKSI+JuTX
C5PpLexFxMFKhLk4NlvXA8kACQz5Rv0LFQnQcjIfrFBQUSnWHNz6gpCHK5WDMqtc
TBCPVdBhtBtBMYIrKrC13HbtBBY7ynf/Dk7nlrVdfa0HMK1cz0UvXgiAM7yjlv/q
wyAei4lhliuG5v8To/2PAa1gVlu6s4oIJ8ysHy2oktsjplP7jijhYhVJp4QjEj9H
goPbMlhtbVaKDSuRG8NEK1s0JRVtT1YN5nQdmS+WwlJjymr8e2JIgcdRfl5auW2R
ox+J6WRHA6QOE42w8wDZpIOXryNxPdKnAPBYXrU28ypTz1ADZKZ+Qo0FtfjoxvI7
dXFw2+uRBBPbx6wCLAe68NK3lrOx9Gqd0nuf4z2Gv8dkb38WmC95FmvCSzUeNjKW
9k7e8OPOTRFzrEdC2da5c4+4lnyFEpR8LZ6apjy9si3M82WmfHDJvgDUrRxsopfB
Pex0SotDnTXi2K4j+julCGyHPFeN1WSrefcZ5XGB5l3naV2gE6n7yYeGebmDfLlS
Uy+JNqjiWgfcjUHXhcp5Z8Ze8rLm+LMoVWtDyMiQd9omDHHdhJAzFdIZG17NF0pG
DGaTi9mWinhj0AIQX91X4CFRqZF4djl2MSm3E6kX6+ODe50afRl52lYdPW6qejuG
nXQAKJ0/dR6xUAhIRM+eu/wud3s2s9Z9fCW5rm4SwFXGsUaoCWnmEOXi26AtWl97
9v/+ZxEgD0h7rpSioGX6OgkgLmfX2Q6Lmo1AsCOZIItzt5s4OzFyu6JNmNkf6ZmF
GeksjLw0Tu/JhTXK+95IGHvw9GjtNUJdmXkhOFegl0sWdeczBFjPN3idQXHYqD09
7vdks81BhT+Jm/UsBMugwxOPQMmp8735ySS5iTkcN/KMOFGSwLNpq+dZtRaEaZEp
GPv8XqJ6OA7LalioR9AQCJjHJJgy4nBeZIvUx0uwlI4cuQie5uYdx/1jN1PMB6z/
pZkjgg4N/UbYbvzqSK1o+n8+8axIlNQDyWUM4rOzx8BcJKIFpaH5EZV9F3D7wVgr
KOvvCs50PGtiMsohKNkWwyobqq1yvE7yA+Glf7rvMF+feVoxqeA+i5Qa9jyZLOZz
ouL7lSnTtnK0Fc4IlI4dDdUQkEGf3Aw7GnWwNCQ7cj6ii4qO4izCSnQ7hyq4AnP6
dF9CDhZ9Vnqb74e9pTAWUNzXUcmQidKpZ9awxi3pLN6ulCt3z6env8HhqUoKjvPS
aaQUNhizm3fuIvbfo7UxnZKPzHDWcMO7meieGhXndaRHK5tW/nwlnbBrR9Jmullm
jL+QBpfBId3OOjRMp9Qp17cEMNiPcByjy46e3WBX36cVnT8E4OvBdlxW0J58NxCh
BwKIAEx3XySM0153UqnvbpDJA5BsiEzSpBRrczGMN1k2kf6kkKz6LFdYp2+h2vfI
FwuaVBi3B57LZC59wefbdmpD44EMjBVcvsYhtMaZn0w6ckEJyyHn0a0FaSxREOcL
qFNIt1n5xRmZee+Vu/p9RRDHF/6p4+Oz865eyRTRrFiohz8Ew8RQGX3rbN8gmCAF
ZxT2niV/kCF4L1kH35NCNUdiB85sPqMYuaRWxpO48pVa3Bu5MYRenPeCgiIJF7nZ
eFYjxNMnJcm2Hv+KEy+D0zmKLS4p0R7XBGcWG41GnqDCBgifa4vj0k0JeU4/sX6/
tvj5iye9OHRWCu41aEf+Bmb6atAHR8kgLEP/0oLlfO5vVI8gWKHKebQVz3FESWGM
kqzUVpo6DG71jUi6eCBWLZqWQ6Gl6fhWi07JXIfG4oqVfRVMuwIU9WcGnZzq2XFl
eUC3ty4EkWSH4C9h4Ng0P32U0dF0tnQWIuB98iZL2PZ3XR5ecnGiRZgEk/UcEcEZ
qLU2RiG61YMfiWGYD91bGGQN3yYI6bnWnyI690gPQwwtSJRvS/URm1M5falcV+XT
5JuvBmZn0LIxaqWzfv5W1UG2ilbhA9SjAJq+ECuqzCjIS8uHWS2nfIipVFvOcfiC
HG1zV7I1MNgtYF8f6j1QtQfACELpppp1DgzDenDDedLdPFTOs4lb259d9dOXzmSz
SN21MYcDLdjMhjHMw5p77EHSm2bESNah+RABGM2JWR0E37j2/+6VXgfDUk1AtiME
yXd/NxfF31xDRT/T8wblA5Day8sOS064fVwd4sFszYF7eI50M4lf5Kll5vYotc3u
N9PKSU7lw/Vq6qq6HQojgjKq5pyMxHqf5UDOVpl1I/TG5Si1WC1OvKa4piyN+rNc
jFaopaXKrWf+W02xsLg5xl1N3sqLRo3ctzL60hqerS/OZKAPCYcdLqi0uiOOxTQA
AOfl+OyjeoSCWRMojuAnMWOvseiEDFNBsAxX2DQbf1n9FiNsSUMaKpWvjdc2Fuds
0LA3v+So5pssezgEZiD2gdkYpvnUYELSO03gc609HDlGmXk3sqhv+09uv6mfWdcH
k8WNupduK3MfU5zbEGDhGqUjJshiCLCAvtXJ0Ac8HD8f2wiLA/hG7IltxJNWHhYo
MS92mY9Vz4z+DjqvHK85VFZDirz2h55BIE6SzK61GdbqC5fTsx14hdkrpDsuXjpI
0MCr4n/zrld772GkHfigJG75wA/ZVldsx8rkvTs9kO1p/zyEaZTkhHlYk9tPAaSj
tNoWXZfP4OSfJZxi7i9dbMgGTTqaWCzeQDYdSoEg4QOc7f18VTBkTdlp3+4geU/h
pVgAWjTKmtFlORhwsfku7Yf2leGo8Iznelg26UWOx59SPJbDeCnkzPrQNCZQE+lf
/9s21gT1eHd+iYWBHxoUtheZdq5FQLHZs9bibUYEquQtI6GeloYVYhWD6BslFAc/
t6qYZawYYJRVrLGF2tXqiJI6hhuK7hLYaqy5azU+zOe3nJP432xqQpqA5HP//RKk
tYor4G6D83tjLH6mwBOMUqEk86F3pd/kTsI9M1e3MtbzVmje2V8W/PpUOFwJVJQa
5TEnICepWONlbDM6tg0JMH1tK2j7gWQ5mzq4nQm77QbQ8VAqLEXfqHsz6UAHLbR5
ZGCowCDK37WnfGzVid/5hlQEaAj3+y0JFk8LUQuvSyTaDUmDYrYbDy1kSWG2+2Q3
10y83NwJmludO+mXMl1sV9pF2R1KrafRGw2Xx5agbhXBD/TkI4WZ3IHmSWnQmb+7
KvD3wlcyEUyOlTtJlGyaimBhYLlNxim1RX/AtY/nvV20qcAJMLQV8UNchj+NyDJJ
P9kGC6ZR86F5dLbj47ejKqtl+wTRMwHVznRimjqbcHIfoO+ZXDujCDzOaIgDQYgv
7B+TbZnbOsk89p9quHSj/kOnmeE7hzcm8LUFpSOBYGef4JDZl+hwQuRGP/jtLuPq
VlfZ5ySLbC2E7XGyhrMPw2Fqp7u7HIBTpqVFUWe608Ou02h/KM75CHY9Xn2iRZ2F
LMCe466bdB1j1qx+gOGnJ6jt41mzsvZjp8HvZKPTmuBa7qXKpJLFgpM8D9CRpRZC
f0sus5UxYdMbHZpyoCD/sGX2n2U9plbplSixVjQwLPihm6Lz06fbf9jwbFHMVEQk
CNzrBzFLGwb9GTZ0NgsZpXGYcTB5kTw6Xr5Q5GerZmseKujJhSn69zoIShWrefWF
d+Kp5yXSZH7raNpzaAhJDWdxalsjvBMClxi+am1NQuq9et5c3+0lMqj+74nNNdyc
BHi9OacNnqK3iYAxsKaSETLizIDiK79Yzst8cRBC0P9QbqynpCUax3sOLuF+/MrC
1mtQjO3TD2/t2t4pHefW9/b+lrYs8tGKVUweYGWVFCGzduOdDU5qSPNtnKNDt4H5
/nkNv9oVWrAcbqc5le/YCOHuG0pdjLDr2Sb3WwwkiaA3pn8jXui8fmNctPRleV0w
sd3A/I9JNPpauy+I3hzSG2trJFlxiaSOmh4kVXeuvEKuzQCYeE3q1CCJi1Bjtc9t
iIob8poh+s4ZFxENP6gIuaRcdrkiz4FDKculeShR1XA0t5wTywOEwKG/XA7W/H5B
9wo3T+bPn20sBTGV60vYgAeh9VtHqP00fwyDfZo007mC60jDSpxV19wi8RfnvdA/
hWJJw90PBV2TpOAD1iIqLklEN7Wkfl8Mj2q+tp23bRGI+/R1G9bwKFRWapxQKJga
HsmPrTk5KlITj1tBa+nPY2Fmmt8ZDpdr5Ee4hQA63z6J0dUswGjVyYbaMy8RGE56
eAIIcOsa+jB07k/L/ovTQqppdoWGovVrYkPqT1gGM2O2nzv6O+ls+2rcL1ePuRgh
wVJrJX4owRAqOiYQb++Hz+hH6wz6cvjeZv0Y+tkkqOoNwfBdQCpZE6tUqZsSOryD
Ui8QByE60OhgyYuwVYEqX38tVDHxYro5Xzkmkepyr1rxs/yzldtXSRllxBCKtLl7
wgfL9Lj7KUEodLsdUJjBd4cUAP1bgq+rtyJ/9FfTT3wvBL5nPvC5nC3lvVdX1r6u
Ejg80gfuFvXVt++EpJZWqhhpvIU3lffbcPAfp+GsYXPhp28asn+GdzlE0HEetDiH
cf2QDq0nxg2JPb4e7JEYevtRII/qAv/rSBd/k7YGlWrzwlaV/vYcRqO0gmo8Btic
kF18bAAwWrJ5qPyjSIMiX+uRVD7z2rolyOS/dRaZw0uze670rkQtyteWwqxfXLCk
dZLX/Zc/gYCht7OIAuFI5DPBua9lwhDHxUHwip9OgWy4o+lmrYdYcjKMhyHrOxY4
K6bwpNDhrG3eNHGeqBkllZe/j0A3X83x15qNvCdQQPVo81xBq9MDLXA4eJmTnnEA
lW9uBKCZTkvCB5VILRSVvxj9wolWKt61D1ZmCHd0M/FnnQcRM4XT1x19XaxX02Zr
Jbf08dUo3MZJFgee4i8bS8Yk7Fdw1NwqLa6iuD5RIXE5iLZvflA4vPmz9ALnvmc8
uTQP+L2jWvE7oPnHPauuAtuM+dKz9X4x6eTDOFqLAT26g/laEEJTpQH/P4BGYZqT
rZ7E0Mlc+0xBfSL0OEx1USaOYCFze6hKMHRoMnsgYxxF21vytBjwa6wzJBHBmC4m
ogCgv8C81oeRYTpuihfRNlKRpHkLU8dAFfAZxaiErduMN3KsUHT78FsIifgzEGyS
znUlY7Taezh28ss65QSSNSz/alrlTRglyXclEfbewbnSBPzwdlctpQnBvigBOsfo
gS0mF3KYT1MoXJ7tRr9DX1mFAZl3daDcV4KyfzU5hYyhP9sxSBZ+m3hkIKUfiKm0
FOTf3//GN1yAm+uWca1/+lBcTNKmw3p91h08zpCcLmc0YxAj6Y2pe90MhmMtr3Fb
wa0F5Qoj0nERh06stfx1TaB57VlDimDr4XM0PJZ5Bev8GZwgUnNzmo9MkIkKEQIV
m6yglR+zvn+PSkbWF/93I8r9UKruxOsL3tKwgeHBIW81SotzVQImhGuuIRBc33vu
tk84NUPyYUldVkFvgr7VWK72x3Gqngv3I7vYmwlcwC/X1RxDS9orqLEYAh/ZFtBa
8xrQ6niqu3FDZBLJXaaaJuW/TzcBNq2VSlQRBfpEIgpwviZR4cKNBRMo2nQg47L1
3C/xyhJQliMhr+lMAHG5t0ltRnZYtCS6eGn9geQFzO5Pj1h//mvpeypCcf+78edB
pPh9Ye0fKeitWKJHM5qJziDi/VBD2afVGWccyky2ijL8yoLAGoTNdLcGiwotZRAg
vdO0Fv4RD7TPFwz7Hv9vlhuGGsMQhHwaN75HcX8+TAxe0HCmZh/reTWZBZPbzh5i
vLFnggEM3BGO25NHO2+0TMuhKcEN2KE4kq/ujsUiRZUmPqDxeGWRdp7uOmgEHCHU
6frXlZyfX6lrV+SjwbgjGclrU74tlgoGrKGb3ORRMHW8R0SNJMDljwN2OdAzI0ZS
qRUTp9IP+ouVG69LvpqgkQ5SLr/zqrHUjipIAu3yA33mbwX5HrQlrS0ghHSf+oAl
IC6WOmCOzo4memHwj52r5Z3XBxqJM0SVtFbLwxdVlqhaKfmsZyGjlyp0jpy/v80l
1YTBXwJgLADMbGe+yLfkJqKM1mzDIZBY0fWMFk6btzQthDYBInxGkoSy/oAQxLny
P6585KOrMLZonF558d2HLyE2oZzmHkyhr3z/q33NZlHwHrtUuPCfuIB9/JL5cJ2o
ygqnixyg4MkXfDz5pO5Gfyet1tF2lAIilFqKEo9vr55H56t+8BMGeJ66a11Lkl2J
yR8mk1xfxANTgY1+kZeULO8Et/O9Ms8RJFepS6/Q+7I5xQtGH50xHIcX1f5hPrl3
cusZYf8dvXcPP2H3m1aENJbO7X3ZDZYS7LK14WaAXEFEcSrnQ9Cg19zN154i34B+
FuavQNs3MwiNW9hnCdKF9OLhP34feKpQR3tO0nPpEKhenr+mtdnlUbwF9z4LgpwO
mdvUEje0HjLBF1sGEGMY1gHZ1KXH2lTLVKMmWjE07IU6g5klfs2/yhTX9JNvUwd8
8Auifj30V4/Tt912D2YxMvzO/YvnmKt7VTyWnAJc3Ymzwx1Ys0NnXB/DMBiWbTJD
Wn0RKgaDxkwwOu5Q15rvwH8+MZEwYwjyMXGrVXPqgDxhUNgs7PyrwcTc5/2SWyPB
wB8mrXY6asYue++nSK8JZeV7htguLSV+e6A9mWjJHdGh2a71bQFJ2YCC/6JXnNJX
ceIzrKqck/xnI7MTMbLVxufXlt+9zR97oKC76SoizmBjUPZn0VQmL2h7xewf48wy
/Ns+qPfvtAzqWYWzKz/DOwESROaLfw7ihhP3EOEwpfx1/AIT75aj7uUs/1ho498Q
60mmGFpfu9MOd6rcUbABHyuoMaO841DwItqXFZgVy/pk+mUdYlObqqVbRbQ4j+Fh
lPu1cjPRl3Q1dU8kFg5xvYHloLcXqkf3Gm85cPHsNZriCjIZsJ9fFQe1dXAiIQ66
zN/JOBtfNC/XYvJTZg4BVwUeW7+ouotKPuWfMlYPp+AnZ693BRRvBdiumR2pyNdU
fKd3rMt1Y2UMKM2OfKnTEU5FsiNlbIyL/kZG2dWv5/+kQmX0GYP4XqDmrZO337Ct
8iOW+migFKqckqz10osHKAN1CWgidWPc70BYwJzPB0xn+vSygbDEoonTde7shH1Z
snSO6EMLG9d1M4OCrlbxbbfdi551o7MH5sV5YushjA2Lqb6hMfeuInjWTpttlf4g
JbnXxBtRF9wlBu6vBm8lqQ1hOA2eoFsHUAyN36qJQJNkI82DH5czu7eNccQEUA71
rLJabGcCn8fsY69/3OvpBmGsAg0n4yiQat0JOgIEOoemuLcILbfGXoH4FJSxD+o0
fWa7uNvGuRGU0yVcHQcJ7MffraL7knB7613yLQlVwZ4rOe/W5JgzgjZ8m2MIQz6o
77BRiDwIsPimQBiFukwUH5GfbEiLoRmDGrYOuDOymdwltIF3JH+AmfM04WlJD5Tq
L21tTacwAMVVw/MnTdJ2VxrVfo9Iw9fi/A0KgJgZbpQv82N3b0xWl9073GNXGMLn
JUefNiqIuljzhpN9eR41zpzbqYYNSvZlsy3KvZBlQBh+0y8xAZB+eEhWyqcqQ3ki
+fbFY6FYhs9J1W0r9XbKNK7ilPb2YWzq6EgUBOv7dxe8sfuyw+e46vofwKJEI491
CBlu7s1dqR9E2WQ87G3tIS17F85qYiFxkJoaDZGBIAJ37lwq4HmqA+NG7Og9VutK
SsdDKgBJjYv+a7jRjajIIvi2DDNTQbSzfOq0RACxzkHuza9PDTWCQ7PnRUlRZeKw
zqOo3abTiO3jXUZvOgowo9bst0u1n6RdL0Gm2Vgpqj8S5qomtgGM2QP6w1Ed5jSZ
VmVH6GzUfkZa1x3CA7NZqtg9wOrIoNVWM9sM1DD4T9W06vg04uHGeo4oFVO6+9cs
EUzG3tn1Hg7ghk6PRdkCNn+H9p5qJFXJDx16tbqjYkbtracqLHAuKVKCbWC4X5Hc
6p9b4CZTpi+z6XeaHuAyM5/Qei0VgM2aIe2on22G0LyH3XY41mJoA/lExdBzUOqm
Opiae6lQY6frDd6ImCFXGiIsxbbIre9DAxPxAEX/cTIq8NnKQR4417FBuf3vB487
9/SZhlvbpN12Ti/C5GTb8uHcGe5x2mdlCo2H9BekWHUJJKJ4ypZNF2glLYOXzdoE
OtgrWJSTiiEEoPlVriHDMB8eMYjEGfypkKLFE8hEc1fex5DMo7Us+qzEsRHceDgM
+oAoP12Uw/ZWsNDFeIzdHm2N0m8CWX7HqoBrmoO492PFaNcdBrumlIPhWELb0D3n
6SNwErXcrgRs5phupwSFsbm0cimVVL2hMrZGb4wojcgjbftUqMCz5Oh7XgMHKe7s
784ojV2UcdqBLtGOLP1VB3wqF6gz0Lp0Yxd+GnwRXhFuD8XXj6o0qoOnMALgOcDW
OlZn+fXoC9Iq9sh+6dZkuWAcZZRIwf0cHPWJAoR6sp/Z48MHX8SjPR8TCAgiKioV
a6KqMX/ue+4WCdmCr+tR+x80bDoqE3AxekIbYliBHA4dHyhFNal0fmmvdhwsXf0A
702E7Rp9AomaZD8rTrIekkbhoAMUV3xUCq72jwU4yuC39oeoqPgETjmNLKa2TXzT
xCxnl9qneeaVQOG/qI20yA4j/gGXssS4/kXEsVG4RPS3WFBYsNhi3SVHnViPhLa9
Ljk9TETuX3nms0wT0URIbr2EFfe1CerXPB00mXUz+aJnhee0Y6u/4ukexREG8V8g
xkzuCOUexK5tmyTsejt434wprB639qU0bBlAi8uQU02ZkeohlHJ7/Nzof/FWIGY1
f+EMbW/luMh4Dp2h77512SA4UzYhCjaR53yBgoERmUBoWxglpFPiIFjpFY1jcI4Q
zXvnykwaJcKgmZWeHcE8r7aOlCeWg2nYKRizIJ4WWIXj5jTOeITkI93pbrf985/K
L66rLpYMzzxhO1x1mRMGMsBA7MuyQQe+Fz3mT5+83WsPZWJlmEOQDs0hyTC40rAu
UPnnbWJPR1t3Mj3xLURyNoCD0ZM1qdMAmNOSApbpxQUOJvMFFQbxE8Ho5eu4XcTf
RcRl4dM1YCwDF0WjbPd6NzF/OJ72HkwxwcbkvI5S1ZJf/5CgK8ArYJ9hXH12rycp
yUITbZD/Yt5zSG6RCVu7dufdVOeDdWf7aSjZjwRPgzPCaY7skx9lyIFuf/7qa4d/
XwngjxnYDSm0KuUA6hnAQNs098t5F0fC4NrMADU5bunT3VaMkOlqDyGk6Y63X5AV
OtBbV/Bo/vq/quqWXE5lwYJeZDJIwwhimDwxRqzcaxYG4ECEMJ9p2VH/dAGsxrMD
crt+zGz7WWHk94IJbnBfULOHUR0D9VHntzQdopzKFeYI53PjDL/FbM7J22sBbp3f
ZNnxYo4Pl21gFvWF7ty9cNifov3hDs9HZ2zlFHTCFaNCqetvQ1TXIzDgHD20f0Nf
Z4uarCclaeDARueokETuEIAFENsEhoLK6jzj6J1PuOzVo7kFNtSfSUUbHjppYkwQ
PPnh0HpSkSOyyfp9V3Rmjy/9uPDXyrlTVmHnyUZx1bQqzFiQBPeSEXoolkzkIdNi
kmujkFI7KdwvvUlT4ELpyVj8gNE2kzo0ASXnqpP8t189Y8PPdKKqHMtXbRoVYDLx
vk+xVst6BOQK+HBtuLa4rjgEeRktkRL8wtBd587vySdl+Db2HKt4vq3pCHidSgqq
EluiYkG+9VE1q3by9VgA/1ody4IfjVQA9/X5yMOxBjBWof7JkNfMkA7wQhi9MkNL
XfCMiTXz9q9qAVvAgzpYxoDF/bo9aEPXkgytjH8HuHnktabilDvsJ/7FI1Mruhkz
t6UI0K51OLLDuB4IodrHWXG54kcxytHoiBgHzMp2GRuAl5bZQeXIeYvzenJfzYpa
0kMcT2AmfTxs5OydPcOPE+kzU0mG/bfw1KraTFqnmi9lUyedk4+CeMsz0RJtbMu+
1GdQG4oaKNmZbItc1skMcrByFYX7emOYUK8nGRuuPz0yS+M7Scp7/6JM+j7OuBrM
u49nWELyOd6t4OdisyzOGlS1rycgGYayFUihXq1eX0OoGOqLCHZ6JLntp+0kqemY
t3Dyk7xJOHiTeIJVslDswdg/moAMy2Y/Ii8gY+tB48ezZqXLyZX/+Y4cmRQ5I0xR
Dctm7AFEB06S8lYhgKsI3XrvvP49gUFBVW9dKeERQY3zU9KJBlWNy5y3Y/x9exd8
0weoPx43kvseuK09bh5QSmtJOcToHaB6QteuTXtfObwItxawTRTXS3I1xlk3vKvF
UOze4GkKL6U+sQ9BpJrCUSYm4omqsQoybwiRAn7/5Y9YoG/QxAdmR0ccDF/fHQup
u1RkGD9xD0nFVhd3k1oL2vgSnc+cuehFeipxBEi2dHRzEm7d5Ykip4pOCzusWzXD
1X9GdhxTZiLQ8t/QWdXaovQcPxc4pw0L9Q3OZXBHHwLG3KknJRzso5nB/Sk16oYM
9OVGUMZQYHAyQsFAYe7hwOwc2tLu8EABiLIs3BVxtDUrSNjexn9iDTQzk02UsIHw
Ol4UhQJXrHeEJPirgK7HvQz3X1nkJoydIYuyD6TpXiHTzRAb76XpSh4Wjj8Rschk
7hxqoHsGoYdeQZZcdFNzIo4PE5LqeLf1qJT6u1jUixZEyuvEE6NsElmxLbiYt0bF
PGg4Km/jSTwIuERflWN7kRYsP6Bg0CGOO/2mOf3onShdyom9RvBuAN8d4ogXk6d8
cj06AiQcbtrnJ5Z/OnFQ11RXBHRUBTe4xtziXRIrTVey+ZWYOH+Pmqe/7Qb2/rx/
Dx2Op3hhWWZ8ItBax274kpKTCjcL8TcHJzDmc8lePMug5khiUO6JxGW/owZjQhKE
3RCOglk4v7UGN7U2UXHdG1oWb5I/UcEe78gJokOvre+o2M4MinjVCIu7igKeoOQB
AbcdxiWSQVwlpEbXrqlT35vW4sGlS6NkJ7e1XfzJnO49CCmgQBPT5q6PHa/n9Kuf
4GNl8Tw1clmNMt3sHoAco1pyWNnIGCYQ9EjaDOp9Z9NZyJU3BnqEMnJv/SvnMaCr
+PsjIKflD/8U3rjiqThdLcRJt9cSNmAhPlINm1e2YaKuGot0KHIvyHwp4zmL3LjZ
Y2sjQLZky8mqihescytb6LhLOk/jZhe0MHgkFluzHcgC2pt+WlLXWZN0pnYUoSpb
BjUdonREjw3+Xrmtye2ROEmCE4N8W2W1T13hiJ53fEJVGXrqramrNjgLWRSRxTcT
ceUYs7tgH6FQiiBqPazhLLSD3W521dWITk0peNMqgaMb65THhKjyItqMdLTSW9X+
v8GIjmWgPSdmd2rzCypPVeIFUhxYuwgYO6NLstE6u245D1xoQY1pfuYzS+s46aWx
a9yOT2kXlA6eXPDy4Dl7xZfX7KwuCv4QzqnQ9t8l23BcdVXjCY7BzioDlvm06CSB
6yhnWofMgRW4UyIAgxbACGCDA9vx/1s59bLU6b++WD32Q78Lk1UB6xtbMTG5K6FF
2Sm6Wse9Y4TKE8DipmpVesAKRcf2Zuswo3ULUzpbf1fXmPoqTRW/u89sV3SMwDeY
ViFjnMPwd8LpbheH9tnIQ6nbhZs/cs8gs3/ctRPQPULQ25AJknsuekbQr5O/hkCq
MxfpIIjvvCDI/i/JmAbFQdtbMefqhC8wJ1mMGD7uhwJoDBeEpZK5vx/63oDrFVpz
2bsf/p6YL4rxIJYNWV/HnFX3kAbnZaQ+3I6n9qDGxy/mBDeL2u+y+a/gFN46whIB
GqviKXb0BOpnE0jwUts7YILxtQdmYqeOKbpOLzuyJvvLhuwnkcNA3wUemc6GrVSv
vdDyX2AUniSgqHCi6vaA54XqAeb2oImB696SkpeSNKXmOREBec7uOMnoYIWKcZMc
7RVg/qxF8JE+gv3+4RVRfKfpXMgj5GCpx7+Wj5rZqL0ExDmp+g1PtS7zvGqjBYiT
2Fv5Wkp5BTIFwpLS148sF4TkPDEzxMYND3bq3uJH+ig3m3HSOyorl6ci6CAnS4aT
gUyQTNEWAF28GTP9BXCThRjRLoi+uRnP15BlLStsDOSRilmHaM6qWLcZahhhtAtg
HmrdANdNZRNg1Q21BdYD9GPNc4RSJi1qJuzEQZl07MOtrXsQ2ucLwoHdFzPXlBmJ
j0wKtOx+r9JRuMpe94So+Gywawa3l/08l2nLGKWZpNq+VRmQCyEZHPUHaPNDWIqA
cDt5TCkfD1tFudE0Ihf0kqHr2z1FkXd5MoDyEXMDTW+zS+IvL6aDHhXqLtIGie27
XA91uq6atiehSd39pJ0Qy3geQtA94elgJWJYn4HpwK5eBuBnfXKO2M+3MUz+oIKI
s0UbaDPMEH/IqTlq3Aov7UFStNyFd+jLTkPsXN1a7Sw2q/9JO1QDcTisX20vabLp
/Cs4AN4v7B4tkZ5Z1UOrqyym2+gwfM2QVq18VVdx5CaNjACZSE3lwHBXP/nnZFQJ
MufN74qCKWKkvU1WnZpybqMVJhdYjrbAgfLk3Bje0UfdqvMG2L/poT5VWJLMuJFW
jFP3HghEC0OjoRAXV+Z6cN9lb0R/PP9jG7Qc+8wGE/uKKcuAwPN/Qc+obAYyfM6W
T2VdM+IeBO6/WG8gPvCwE4Vn2lgBQytqZ2H0/9LtNHpIHBP6Ni2AJn/vFDry495m
ayqTcLcLooEPA8EzdlUqCupAfnIa7HODX5bWONsEOni3o8qQQVnYqRcZnFyjmebZ
E5V5ZJOoB0H7XbPU0Qwu75Fj5gn5j6bfMt2GHV8j9UKTFdL+GW57AAKCK3wm7yV8
Ssu8ita7i1TpxBjNtfrKVb1D8fo0Bl+u2c5SWHVKy83b+mNmfhm0dETJgJ51aGhl
CzA+SG74nY6MYbpVClN+sRE1b+rTG1PPIcYZaIT9h4yk7TUcBJiyx3iIeeFS908R
Q4RSe4Q5BZqdnN3UqqOPT7VehIs1KRkACzb1tv/fk4Y/jlcaElft4BDE/jSKRMYW
FZpnUvrG1dCrD776/ajJXA8KTSeFgPiPXVjoc7GzZVqJCP14uKk/TFnfoLLuCgxJ
vZ9ODrPD+lYi8at7SyaeAxhXTBjAASsqSNYROUITC4k5Dmw5FBGHiJXVNNDJz4B8
LJOWfpvCoUdxnapW+fP2hXEK1ErtTMZW1ze+ccsbwBLAMbyQdslYetNEIVY/SEuc
GfMbrJmx4V+6UJpMxOpYFeIXw57VEPWhfDchJPsj1u8b56ZilfkCcxfBkggYOcI5
U0ZLvTtC133glCcvwbqwYxnFTivQfTBpbjUv3VZBdl9cT0HwmDua/+xZRWo9cEWz
gioUlZUOn1pRiL2WHvpzkXbx7LCeQBv8z8AnHaY6iNcHwXHP95olHcvo862Xc7tF
ShVJfutoDQTVehHe0ci4j04PtmfQb8ARa4uYiYCgT//ltssa0HcksIBxwpgKG5U+
tcmLQIhOI2RMI1QpR4qe7g1pK2i2ggYBDzszf5wjI7p7f5PEQ3fyMUiOf1x4fwFg
n2LylsDtKlnuAKrOTwjz0NJNvCJ0fzW6+cws/L1vu6xBsvlOMFWSFLODD9SyjrjT
h8mwKqd0zzCZMAuvbMSiiNQ3TfWTlIWipdp10Yg4DrDs46rnecPzjc97cHOHp16a
rDkzjWICllPygNlnzGCTom3KYLoiRjzMR3/39cBaAediByqqKKvyXRyT+c4e7soS
/GkiuXPsPwns4oNmEO8h/40Pi7AvqaxeuwhIYzZ0UCLkIXMgtQCMZMbrLXMWYWWw
vayIPQ87FcSgh9pJ8UXdhsbef1kTI/p0DqRpGb5yxNvcHT/qfkcsTKsJhuAROeUj
0BdCxbY3DyO4din9hEanqn1teNR803sRHyvF2Yhq/mq8lcK/RsrMxEq81P+zWBKV
bBlL03QHFTQfbZPruySDSHQvdolS/5TnL1csq52k8K6zPahoIi/VAg6jZcNIGcmB
N0mpHpt1Kcfdj0DH40tz4HIpw4Bx8UmATVI8B0JLWo+q8LhhbZGpJDQeKdZNRugg
pY7u8UUDeI9CYXbrAdSTflNB4RNBYHWjf1X1FlKvSkSIvyrrX57Hgm8EiupiZeYD
ZATH1zOhEJKS1KWkGvZ0pY38wqUyflEBFyFQDuMwNZ8txRh7f/Uxszv7UEfGYchi
vfGFqnc0qrbUGprVBAfRzGgbY1P/FiIE1anM9dHw5FXDWnJ4V6syY7JR7rJX9G00
nCrKxRSRmVixusB8BtO9A5U9J0tedoIqSqIpiKR/sQdArZuNhJKI7ARl4XDRuCYi
6i7BvmRWbcTbImMewHd/qLShxNczmHS4qPDnfcBeNYy71byJuGRp5d1pGDgDONFk
C0rGS+radLiya2J1XpFtqsWTMzmE0V1ixj5+ei0V/0TsrbclXOuUQNfUjV1UK/yC
NQD7qqSmvffUy34ZW2urRzekRgoALgd19hPyC8cgJyzP7mXutclcXrtbYJ5hqJIG
DilYo76Nug3mT17stcDbBugrLaj8l5MmuK5ieIwSJ4dYYKsO5gt/v/EKPjYnG040
Wf0W8fw8SSoLnAP21o1378mcutbYgLshoeQ/tdYQV2r/10ikQj6Y2j1SVqoEl0vS
2AsWkr8rvNI1xWArq5ewLWyBUaWkK/oAMNcdx5IcO+24nqPNXkWHr5RVquwnWY1G
qZdrxQKeW/d8j+ohKcDZ29ODt1C9fJp5FCTdHKMU1a1j9X0HZlGsw/IbdzPU8YXy
2oqRcTmVoPxfPLraaUyMUqkowvVILA7qguXQHip6LbvrWakpd5iQj4meFdvvl2D/
QyeJXT/6X9aZYHA5+HS5wQZtOj7aHy7CJmHhK3uzvGHPTTgH6KEn5w279A6/qymH
efLe3s0b61u5l7wImB1NbCSbbP6K5sr3rbHUBRo15XghbCAXAUhTbZnriv8O6MiE
w/BJ9C7Gtd1iZwQL06GPWt/2o9zaQsHzjVOU6tnFAAaktUmEEMNholQW5cbtRS9E
7z/SUveJ0u1pWaK0LQfuhAaV+wXV/03f+R6TL1saVrQAgSYXZi51fNzuXH09WBvA
2RNQ3lgoGNqHhJftpZ4U+ZZ+OLiP5MvtaECfXV1fPY6BZG3gkRHaq4KWZMz7QgKa
gmsfQ8NXplUSNNSDamfM/+2JLFY8RMEYAbQujZHmT6yOEY2cQWvpVgBgO3J2GMt8
BK+YFE1Q29SbKx8ZC0ARNIagE3unOVQoKlaqF/rweUUbaJgYC/a9YwQQDgO9xefX
/Gqe8RPu4jd2V6Q8KiD6e6tKi+2DnbhKLHAZEVhe1dRib1/V/4c76OZiRktpx2/J
VjqJHWFqTlgU2UxmKdsZVfH+2b36eWt/mjdD86I2HnRX+ydRio1yV/hCJdrYhjI1
y72qFmu7n/Vlg6u7GMAA8gligLTOSA3E217gIAXHW3r4+1EivqYDfPgMAtcHlfHe
SNGGd0JbLsTVmN28itfJ8Fb93zAvtqFX9CMah6RW1h5YpSQYhi6DSvoieGkAw4PI
4zVGa9wbveUB4MdLtvkZF4zRWAO+Ziq2aPOaRfxPmGwcRknEIJG+YV7vmiTMgdIz
zdrKpOcp0Ro5qX0oD3mkB/WSXY2oRqD99sp97Xla4hsaKCXWjeF3zK6j+msTt51n
HjNFdPp4x9S5AT4X6I11V7i88zy0Ucx5Ej0PO2iSytHgGShF2ZFlmPLtVqMPFDC9
Bpl2fe9pNgKNv34NMh3CdsnO2ccSH1s1te3i5Ud2XtJzg4Te8CQqswRwfhKZmoR2
qduJ/2MI1ecyYm/wzGnMKXTcWoyuIYxCiugy/T8rqHYAKRqz/qBrqRMI0kVrmjPR
uKTgItaUVmEamsB+Hc05gMj9mJHaUiZoXdrzdicTmNzsSubEIh59R8Ysw5UoRxa+
gFUZTfg/0iCYC9baQ6rXvguTgbNF0bcRmvVVuq3rKuKrDYofuv2fXZlkPlgJjHVj
iL/csccD7iAPtJnFrH4EPZeqfTo1nBNFyRzZXxXKGYepYijbZGJGLM6vlzkgbEXo
uvpWNuA74k1Hg3CNLlR3kudN/pez82fXesZYHXWaeSB7vpJevYT+9TlcCUAJKgwk
ZUNDI8rNtvkiMpLrKYSP4le5O4HbSdYFq74rRI8Y5ZoSEPJHcH1mrJ2Dj/MPjSEO
+UctHbE5uvsHAwnCDAwJTxaGAH4IY+6+sTZ36XXjKGDHYJuTWsj6xh17MfCqK9bV
aAA21iET2AfEBlU6YCVVm9U3e9Rkov8nR27MLx8dDbo5yismU2dMO+xqpxPdRnQB
xe+Tc2KM3VH7CHdojlPBtkJHqvOwg8LENHQ4d2VBwrbN20P8Sk5rprJI2cgJO6eN
7apa+okHVKkASNiP2C0Y3yf9p3ZW1ITEtqQP7QoF7inenYpJmD3NHVGanpGGkUh/
/Wov2iIG8rAJXmNbSgfiJeyCm8cf04kkkYojoXuP7TODT77Mn3BnwXYW8SGugEHF
Iry/iROeVeBlfoVTCDz6ZK0OwBUUe3juUYOiSccxjOhAIvyDgZmIAb3SOAbTpxwk
Yl2/+VCtZ2izhdej8VD0WQDwhan43s10AwrKnHeyAd6fCaOa1Ufh+Yg8WqgcEZ8z
XHtCDwOzBoirMC42vOsObw+c+F8xCPCAI8YSSTpN0gk5p09xQI+H4+fXu+BFHPwm
BDQt8j4ifCB3esnxEQEciPkTaJRaSt9RvCNNUl4hvtCj4Z8qHubzMCsu+TTE9Qyn
Az5zCQyRx3SEDHS6wnSlC8FGFq0pbC38hunp61C82NC2UBgai01vto+t/v9nR/UW
4JygGF5AsiKhGF9U50EomJrvdwRCHqTu4AAEPfqBjpMDFGkTiYSLM3jaSRrB3TbZ
hlT5NqfF013NgPSQOKnhqHztz1KGJhqWytQcrltmLdQTVSVzPphCWGRvGN2v0lOE
VgllTD4aVZbLmVW1Y4ICRoRF7m1hqiZvKCfrftZauSOS7WgXb6MdvIqLjzvdaoYD
AnIMHKW3nnyNuzl5oOfOA606i0E+wbviqa1J/dpH/u2fNUbFXZ+zX2NEfaupvlrv
Pfrj1ELToFud6RK7iS8FhJjqJLFyuF1sRAHzLnEz7fF2rUf160WiFKZ+aM+u94tB
LKGCuur14RTVKfWRu4fCl7h4E2k62h2927a7u04F8j192DBeXJlzp+VBpBL46gI8
R3PHEJ0roMs2OS5Pd9gvt8NMTNSXeaplqBrcAVCy6oeeu+Kf5TVMSM8t8oNf1iyZ
zFgVxI+W6v+OBcPKr6nwHF8vdWirYlvbmNsbnrmRazT5M5MBo/Ez5745iypdv7D6
NsYx67CmhzV5OnGNVKmuRRCfX1WkSf8s51MMSgMC4UK3cTVa9FJqkiRFwh8K4SI1
+GYunrTz+A1fVE3s+xsvS0FqlZPLk337lbrbxn6Ag9bQHMQ2IrG2F8ysynJ657Bo
g8yJQAusMDhKE1elb/nNELxGlptNIP3e375VmkQ3vTkR54DSy+qrJ8iaRpFrh4vY
hiAN6EKkEXgcX1z405b/w+WoznG7wJwW6T7UOYqgTW9arF6JxxGMuWzlqzjsPy04
IMi6ITgkiiDl9Gwcp7c+jvltpuMtcX+q+axEjQubXJrFoOgoCUwuEApENKdW9kVG
Dmxqoi0MkfibTO7aGhbiSDBBHhliRzhl5oNllLrlumSlkQV/JhxkUKmf68d5ZKdi
qxSsYpT4o9w1LWDyr7kussjoXWybraZw90ALZMueH22I0Yq7Z/NZtuE77wQ3z/dI
SnZYDmBNh5l4Oo293KrpsSZ8pIUg9ThO42xlBfjCm4WP2aGElS6JrTAmGcGYDT9x
feSdrDCuiCzh2HO9jQknzVH7wG3WgsRAbTG9AVZTcK5SpTGjb52YiVcLHV14poGJ
NaENGJzQSe93Y2cz8wkcdo4qf6FOawkcJb/vNZ2x5jTnW1jE/q857iJBG+cd/BLQ
JNrIgyCq6tdb1x4/2l50n+pC4QixzvwaujdwyRpVBxfHZL/TOB8JeMr/+ZGdtfIT
sVmN3jRgQhtDtEXpELEj8/L1QFb199aAuWe1kxCsMLWsel5RHmB0BRtxmhBGq4+K
O7yP7aSfO/Gjigy8pYyauJB/dAdx9EcPbDf+8UruZCHFox8jV6eCVs+4aQKBpbnv
6zM64oHv+aGu7Sb1BTRq9Iyrs8Enhg7/KPkWoAIC2FBsCTipO3ghyE09DLht+KzJ
sFas3kou4MEBdwof6rLHfRjBk0utKP3lXQiWln71mxM8TF7tvG88gmJw1Nz09khm
m5pFyR29zfe/4zooTrTc1U8nH8JDl6e5vk++1BKHTuoXAJWJfz7fGCswiRjQKf3b
aFb8BuIjNpjOgLXu0Q+yHJtpAj3/kYnV6Q0UrjgKQhCDn6ROwvpPOjcK0Wh5WTRM
50LC5+bIieJocRuLpDGhc+NHLaT08ksRJ0hhguw7VvvnjVNVkn0CUPce2XQ08xSV
UnZ4BdhUg4qHpJ1BH0ekkxJWqIbg6PR3gIRvdSfnNISgzVNE09z3np9npOt6OPIa
5UDxDT5kgfGUOkWbkHkGQv0Az2EO8/T9mc2wKpjhR3LTVBZYsVsmUZl+t1HeW8C3
6gD1nxynIv+o8D0FbubNn2ZeoHPZxBxLQ7JrYEVBIRHVwFj/jIAwFResCSpEnkbT
aKeH6KBz5Xr/7eE4DrHg9Q4zuwN97N5b4HwwmppJ/wY5QUneDhtnPoVkJ6glOkWX
5WLeUr79KhmHrr7D8cmfRC1NIEh8ZjP1yOUZAhNi7DkiVXkWwdGJLtANtt4Xk2r4
kD87qMqsLlv5zpiI8ld4uZk7o0nAlhPBEjCyocQ5d/BlFOVApxHqqtjDVhwRGtb8
NckhQJY0LnzfBp7oJVGFzAy6n4RR30VwCe324WU3lp6GueJVnc2QSRXqg9Q9eS3B
hdiQzNx78rccqs7g7dE+fc77wmdWGs+AU9cwO+sRC0te4kPnpc5qzQRdmIkzGH+6
swgeVLRSc5cMDQnj3+w40fXakZULQARjfNVVqJzYFJZSiYVFoIyuxL99YCn+oTcB
W5A01RfrLXsefv/Ai5CZaSv9g9AAH0IxQRHMlwoUUhUtVx/o4wX/uXhb6ZwnMyZI
yBZChBmOy4MhkbeRevsbYFSfh6HV3MaZBTxmC/rw4KIbG3liX0ePx9428QPBpZ/Y
/4pXe0bOvgf9SSHSr5K0a/gI5YVO0xxlUYfbQsch9C1VtYA6VLiBa3E9Cs4y1c5U
j8xtQdV9oEaFwqlDmmR94CU47GYbbA/tdGUTe9w1Mk6ehfnB5cOoI6d8OgVn/26k
J91Y+2BMT7QKGv0U9BF1BCdef33bZ95lXDJZ13chx9ZGl9UgG8YbYERnPpSrRvCT
oPFmik8cMewUSnihi4CrrqPMbF/oUT7ULBFhZkZGuCSLiVk8C7Lxay65BKpuC1mS
O1mvm+uAXpe5Fd1ELDjQWUXKjgZElZoWYFqjAhOyqEPDiYZP8S2CRrCBa8rzeqtn
2vDpA/UP9DIBSjMvzGmKoAYtUcDKyHBWhaeFCWYA2PKWUruHIcVY6oS3ALwuZQXe
EHt3UcqvRE2sFLNgyfpEA1qSrk+9zmaVkNIUi53E611Al54ckMKAKDnNSTZlHpND
/3K/p3/CBQuMeZFjR43AVIkojw7EB6ZyKcDiD1MPcsnIPVtvqX4nBPwrCNvDOvjB
Mj1LE+anoHvlj3ixI6Ipa0GWA+HZeQwCJX7gAG5st2YZbGSUpQtl1ppwx903hWJ9
gIhdET5Kg5KJxai7BoDO63HyX+LUb4MGfn46Ep0g3GMCritF2g1jV6O/dN1KgGCA
ge7EnkeCVSq1khFa2uooKgRkTfCX93aDgiIirDbgBteb/tTnr5PWsTGUgnkLF2Fo
HFTtIaAlRZpP3BSOldUFQWgPmrKPn01qDFIqTciksv3M6u80MwjV3lwwLDwOmYR/
cXpaeaFy9xjhvAnuUPPP9wZDV5vfGqtLT6j0PhbgMb6EdY6QmD6ykrF+d74jOGwb
9e7j11PE+WD1sKOkR4EzFF2Eun7PGyP5ti2iJD4g6/rkjVR1SPzn3QVtjMrlnJrR
CrFWyUjSRCbd7eVsY33cNUfIE8GQpkviHXobThvvafZsQQ0RkHHy3+7kQfx/EyeF
b4NDwYOTUc64+bYL9GBxzLZcrkzfVnwCLOkUSMJzigxGhx8Il0HLdu+j57aHrtXQ
9q3NSpFHzXl9/C4eWCdS00p4wbJWobUrGvoXal0HzfL5UFS0F4dFgsw92E5PWAbH
tqBWSd2wrWFN1MyWLrBiIdcJowovDF/JL9gCV3ISgFvFPK3MvfRF3g34n+jmyTIw
eyfnkKNDwFh3JnXIypGrlOjWhrt262Zdx4Z8XHV2n2RNREcFszqdjWO1XBc37Rf5
rfh8i8uCDNAnQBTijkhJhOjLWMS6ZB3ccSiU0dNdFGnSHUw6Tqtbz3UJqvVg0pdr
Dgq5ZIIAs1VYUOrIuu5h+f2VsFX/pHEaiwiT/Xw+x6pP7u/VibkvkJNkNb58nPwv
yqijIYj4XjsAMQQFnqcme9PQPFCpIdSP+9cqY4IoilDOw61vhIXJJMTK8R6SVFYq
lxXXAOgbEd2NyFpSTBmUZrRjmtJg79tRPhFgLL9so9hVnpLwiwNb6oSQI6S7bq4X
yBkxPHBAn+OXI6RcsW5N4qlCMA47ge8fGRYxve/QthQIB9ztx1TMtB+jxcu73byh
ehL3e9laOAqjSGcReNqiM6I2W2oixqsutYQ4Fodn7GrMGniuFlPWI+7N1nVoWiIv
sLBLV4Uz2My3XQdXIej0jd/KJqRO247q9JD8TQMlIGhljzjrUH0Y1KrzzUeyPE5/
vmehVhpqP4ppx26Eta+/tUUAtTfzvvu/Eyi3Szd4kvdHWG0eHEtuibMET2SQK7E2
4yZofIwh4mTkk/zZM6CHeJkxuINnEGHjlshcso2xB6EiEu/IhiTNsCawxbjPdn0K
qdVL91dQPtLQP9kfpaJU5dit9LwmSV1+pk3rat3p6Jd1ortS+mLPviDsPK0Rr1tQ
5JNTUYzmVYxWYcpAP5cRoVE4FvDVmRAqc10GO8OOxbi6QrAvd0/L/eZQdh8XI1ZD
Qc16eH0Sp8zB8tepRKWL9QhWlEDqyt65PPFVQv4w/doUumX59zJ5F4KIN3pcLYAT
CXKhZy5dyd+8JgxI8Sfd+1uK802taroQt7aOGG1M3emOsNt6NsLgcpE4pl7BS/Xl
nwzsLG2iiLLJy2NQRn/Ywlqg4Jxf7XcOnhulcRnuERFMPZCrEktqOteiXbmZmjqV
82dHQGJtEvXGtFoZYcqiMtc+p765HEMajje61e1Qj2Dk11cdMrw9Z/fBUOVfZ65X
l6HbRFv3MXgIJ2PhjoF9cr5wJFjSnaUNUcD1PJMHGDP9QF2NIngaKKLQJKHx/Uog
Q7JJlQZvON3rM/D4mI4cK/ZMa0CT+od7y1a8FO7fCIOsHNtsiWXCWWh1wFYVG7MU
EMcfDZpo/U31G79alhYYViC55r4UZNewBezPXlAJXYc6p/q3vuyrZXehUxWFF3o3
1570S40a+WlbR2gVP+fz7pmR0I1elOMO5EHCzOt6yuwwJQ/AZeP/SSrExIkk8ZMJ
QRdCq16F2naJsEj/oCcpVG0ODzK/icWs/F4bTMRs2L2mWIzZo1BDbwlIoxEXzXKc
XJqaIroM69EeK82xw9m0KF3zqwKVuTnGr+l1GYJFxCrSnsSo6NfvwRGyTo1HSQRK
8G+PrrtsW7mUoTlW2ROiC2MBa+DKvoglbJ2gEMntBdrQdEgjrIkhXiGwUCY3IOis
wKTbbtRMPg6Bvi9NPi+oWgXn3kdIuoufO3gwH0WRhC/5ONIErXeK7BSp/gL/0OAV
1YJtbjuGFj5YzDTL1z+4/O7vn/t8j/QGEl548dB3fGTn4ceD0xivgR8/La60U2sY
wF4rNeNoR3jkWAZMk+mX7WTt1xC4fMuSfWZUHgQBYZAlfRKM+RRD3Fv+XdyYDUCv
AuBZlGYdaoH0x21GtPnVoHJA+tFqv9P456UQe7jtgfwg1TjIlj14KCtWtrzphJas
oIWOeeq8cD7OUm12LRdWhVMKdmX3sDBRwW4t1F1VlACZ9GKfR5/GKxExYgMCBstA
26gRHZMGaWQR7h6VgOjGV5cbH3M9I6mt55NSIpg7nEBbPaGs/RsGeIZ9/NIVben9
FGQiZEPP1iBxE3oqBGCpUAp+xUXCDfQFuJ9e4uJe70A5c1+0CZYKgNXZlH3WliGl
tlvU1ZjG25m5qRFbSbqFYh3kJPsqZY6vY8QMLpr+VPjfH7pPgDJyk/2jBA0tK11A
FNGKSAZkq1+LE8cyKrHwIVMKUdDTFLhDWdb2uB1575Yy6yr6Q1C0OF2gAVkc9BSH
TgQnK3aYkr+0oEBe3788cOTlJj8yfbQOf/d6IQyQX+JOaA89uohw/vXa6q/eMIzL
Dsczm7eguRrR00/Bp8Ug4tkXynUxAG6+9mjdM7mQldjrWtiY7Avosy2CjvjF2FPt
D/Hvz7CODiEP3ox4hshTVv1P3AdkifLj0YKPfzPlyJILO96EUhD1a9tf7crVN2JH
e7dInRQKWEolNooNNgqZ3qOdIRi0hSOFYIBlLX8faYiOqKPZqkBWt3dQmQPPBZqD
CZhOIrr/zJ86pLiIP/nXeR7ezYbHLPe9iws7kMEllb9pOg7qc+8qlTwsz3ipHTZV
hcg2sBLzp7qEKzGsn+aLHGQNIpWJ5L6HmDveXiqX4h9sgFciGjGmFPmveI86f6T2
luSDYNyWr0aZVd3/S/5fQE47Uw5+BbdYJyd0C0PPih8GLUMhVuGhiJcLaTKHrgUB
yhBmWUKegyFP9Z8E3T7lrkIVtm8sNJaE5v8u0HfsfOB1qU8RDCpmvk855OeWSTVZ
OuZALh9Ayml2SjIA9dCgUv+ukyi+rg/gWetOZIjgi/sshy8Qq34P9tdtxz98e/no
pmxnWL26W+m+t2+jqPuFKcYmxLzSO3G6PcGO/BINnjvEqWuPCQbSkIHXAHIhHPjm
mCl9EmFZBdJJvETGoljqLKXoilPpSL7WkQe5AxD5jFEQFOs2XAuju5f6lFNwXUQe
WuB47DljcRaPL6J7lesQlpCY04JbgVe6cCIRw0IK3w+Z2bj2K1e3EK9f5BcmMQES
kKwGVSoWZVPFZ5mokd0wB5Q2nytqNQ6lIE9p+R8ZhTYUC72lTueNLYLht/PyjHGn
TNzo+5rQq3R1HjBzMpPo3ZDrkWdHFhM6iKV/Y4F8D78FqzTNfAKtCkUAlUi9+dfd
Xs0MB17DAhQfXAqSVS8xd1WM0chCiPwoj+8B9k3NTPRTvKb9f9Hft39Pmn+DTAoA
d19QJMOa3DAxCznaXA1ceP/JR9vylsGxRcJsNmYJl6H0xE+5Tm89Mxlomw1OTg8L
t72yczGNDgx5HtswwYdHUjfn1ddnUIaEcNqMBx6IpzQPn0CIMAvmUhxXWxT3CART
lyU+kscbnF9Kca41ZSacNKGhFdvsmDoCArlvDOJEur0k6lfQsQwpsKzM7XXB7CeH
KNlfEIrpNIFV1Z7yIUA6rLotKo7QdzWR1Wv58/ystUN1dJoJh+QCrBWAGnImg1SH
wQ8NRw72Yd6j2q1kwmYbE9AjiTw/0FFje1JqbE6pDICYKjE1zKDacNKgPR6GYRRL
JzFxUcZZhFA/rVdI/71BSslYKcJk7N6zX2OMlwkFGw7dL9k4236unb8uEzevfUFc
ADPvzu+B69CSwp+KWomZMizES4jtdDkm5aq/Eogo5Uwqr23o9XVoaEvEYEbj0Dxo
GY9t6dQi8xwsxESYjj/KgKRFWduMhBnFYu/5Is5fnyFUANVZ+YuzzdHdwZVa1ZW8
KHEkGGluDjnFIO0noescO0H7Xu9LGEOCtA1+OUqkiBI8dX9g8l4pSs8d0uin5u6B
P63x0wVXcxQ/AYqu27GoZGX69VMhaFRk/2jMciemsnli/vzi2t16nvsc6PFifplx
6i008rFzCF4FfuWOPrGNze5fKK8awn918+rF4NQbI/bZxOgwLi1f/0VI77pUO/ir
pj+D6UmkIzOHsWlTBwqowc8bY1ECEqDFJznQUpLvP9Y3ITl3KXj7+l6/1+lTDoe0
A3SidF8+FMsloFbH99K8KhAM5+RRdoHDvV7EDJxpAeyvS1D5KtclMPSiKtN/9LK0
hfdc7zCOhRWp1tlUJo/xuwLs4CzADbqaTCrYtAM7qYH/lCS3jj87D4VG6B4h0fJ/
WpOnErykNqPCEfpB0p4RWFmdug04GxUdq0oZCXzi7P0DDuJolJTf7u0B8XSFpCpe
ijKsVPvO/F/Qoa6q5jLlQL3bxXQW5sT78w2gUiyZAwWyujIdii+MJcxsSU0dKVVP
n4IMQrS4NF8LAo61Z0KFfsf7XqD+OBg44d0apn023uwgwkX/bOLyZWMAOK93hw4H
aHtn67f1KMfgz5/46xInBo8nrO90Hsj+z7QuenyEdADzj4fkpeFhNBjXqeugSuAX
1waH2efzvKt5LElCZ1we8dP6lw//AVhfRm9O/OjRndvCs8/O21fTMdAK4Eyk2drD
8wmPknBEg+EbNP4+2FI1A412CJQk/E5KpSVhhPP+sMYYGtpTN+7YV9MCQUc85boN
0we8epfztpQomLSzxJYo6F91etsRC1AG3e32UoRmeTSCopTi1Du4fpQntxWPVsCa
hcJDnRK/E/4C3coEpq/dbhKIGCnVANOtmrAdJxovE0Y8XwuyoHJPYjcTpOE5vD0L
C4uHbfPgpoSBk3KZGWba7ehx9rQMlMUnbruNj9xUNx//iiBBGnIaeMENILI52+T1
lAmmqmmuBovM2mfjCO3+tWV1fcmjnzXptTx8dESPqbaap42Cvu0e7rqhKuAhdr0H
v+L4PXRL6I/JPw4gt9v2Tg0fqA2UFGIhn7MysoU4Pp2wKh2Rj0SMEfI8TId3Z5f+
Kmk7AmIvU6pzUfr+j1Gvv0v6+/Ku/xHvydzPAbZFmAmI+ONfF3ea7VzTYv6LSsCc
a2Ocq7bALZgoNtUn52v3oQiNthk5C0niTNjxnta4Yh2pqnCtM1I5zoxNtFgFSqws
SqELaMbikX/l4yJZ3uzWhJv3FkXiWk1xi/0kpmnBVOFzj6etXlxjf6vTjrVsqI5l
0sBQlrBwYNRyW1VHPudjq3B4SstB9QBO5/kaBREKCa1tBYtePPkLoOBYOj53kDud
cm9cRtpXLhHBBCePkVD330A3Rami5yrv1EkQ4nz1TVM3Tl+ChH5NnQFL2ir6xksa
LSUb8kahCcZd2QR9O8zGosJjuSRaRHjwaix0h2bxWv/t6NFxXdWChZJusIWMolUk
PCLm8MvGzzMDHPtGhgaOeZlzCQz7KbegrNZM+3PwX1OSCXjXqA1xlrL42O0zXHE9
8jKkp7mfW5mScKFKCW+aLix9sH8zCh4qKmsQNlJVT7TE0b0KIWoS/Y4YkHD6pYjR
rKn01hb3zJp+ndDDbyk/c25C30eFhdG5XgE0Z3qwCU1V5E5H1tYUHCzaHJaDGN28
7vRrv6q3sgm2RqwtuL0rxoJMtCse+lanuagcUS1SHPw2+eYJM98L/nlMDhU/UqPG
YKAddPLw3rU4lyzpml5au27ZK1hpToNFWJb6EEbKTbQije5FD6eSWq0QrCNLLjkB
xP0JUlc80rw4ZFp9A6XLTI89iLTT8oTEe1G2U7mGWGlh/XANH2U6LDMHw1Er6bSE
KHKgYlFpYiCP44CBBRQcfaVlNUXvJ9PA9SH429ULyBMxm+fiVXCrsT6OWJp6l0Y7
uZ2RGsn1dvBvGL16j6+rAP2cyRMlXB1UgD/ZgTu94dpd7q3w8JpirS6AqOHYXeYB
8Zl91xKcGoUOXK1i4eQ/rWoBQAysv3PwI15JNEw4t4OBvrKQ1M5iWm84mVLUZs9J
WQN3cSOlRpywD94C8xxHaO9gvI4eU87q3msncGjBx0q/CWSdVgiNffeBJToZd5Yt
PKqGz1tCk3ypGNRGyNSR8NDkDgQN8iOcm5e7gyJMFDl4vOUqYFpzXphODYGAvNvQ
PzpDJafM6CJmVCpzplgfr0Ks1TyLBBdemHz27Y4x7xUHztPWojC4CaN3WeBk2V9j
fTuJXVoBr8WpBcza73k0dIRXxZAAIMS16ur4blgW/iJM50oA4gZX8JYxCTLtrNSb
aQ5bv9ha/xJrvy9fLka6INOUmRdoVp+yILBzYaPewr3Wi1sY3gDkZ4JfDYMO3Xkb
Fv4aZdW4jSOOhRmcYhvGAlqou/jtHClgEFYxXcnBwv/3xHnNABQ/OVPHYnXQ0ZzI
plymhJ7tEJcbm8QqpLa+nElX7RjRCmTs8M9MkFKNFOLZ2Nsdv0TfKLr/ebSjnrF5
kNh6XzJODRZlJnjvNF3SCDv01B0mwMAuubhOuk2ul527v0Eo3t//KNTG0JoPUSPH
d66SY6hR1Yvs+oFOyTAvLBR2zNKvWiWsKxSvg8GABT4yc4bJTii4afQBTpH4hDoz
QUElePNWd7tRhTpeB9UUgkwJoMrujep28/zfwfC8TBNsMlGeHFJ00TyPZ2oyvjpI
eVVIYIFsK2b0HhkEe+S4ZThI+oIylXsdmh/UFOYL+L+FHwpbzHwWnvmKx1ETNZLz
i98wEVuXvVbFHemhYkzAaa8dIESp580tZVOwApD3ymHnkR7bMb7MWID8tFDHHGy+
wcNTt6ATBWVtwwa7G2bKGM2NZjaUyWHVxiTLRG/1GFXfcoeBHpKhHfBlJFcjXZX6
gnGvgaj/MzDp6eJNcKvvYGGrh3FddepAFGcZs5+IliPisdKWqE7to3FdhBX3spXy
LcVyOwGMCQ24SbK3RCpzBmbtGsSMUM+Y6pg5CWLivjnAjJ1DfJruNcMUcsZ83usB
Flzs2Eavkp3tkngNOAxcwmgcX9H0bDL2qF8YMk4Y2mOcaftzr//8ZwxoxdbkNqX3
u8ihQe0AMovCUomvcqARLiB4j4EijA8GugJY5O5AYiSCgZm1N11EPXoEenT5icEp
rbUhzYCb6ar3e3h0oLUI/CKWg03Z0OpUuDmRpwfT3pJTiGIXPUov3HSsGrQ2l6mY
ZitmJShDA3N7+LqbFFUxCT29RoqUG3sHvUgrvGxhaTDIsVJiV8ywILGh4mMleE/m
U0nWaokf2HL9ZmAavAjkb8VSEKOo3lW9t1WaeAUyGyaj4RV4eGXQIfaaKoZxJNGr
4FVy3uwnwZKiuJ01HtNUVKhqGIT00daJmBawwIr6dtz9cRlvLBoY4JCAnKweyVUh
Tt1rreXi6uPhYvBN0Lxtv6kRaBQ44aAocruupYMBfy77IPVGJ57ogde2R14JYBrq
1JVRzljJ36Va1lqy9UdxN7KdHhRjQfHlQstGgzluQteDXpRiv6OBvhCVk5yvRKEb
smaSh6SEEeVlJZPaDYmn8fB7zRqOpfT0UwJvdwoi5ULmeEJMLuIjUkRYNZoRdxg8
PXoL5XnW4rUwAQorMCkjPofPhbX243yMPUMWEP/zDN9HPeDxnTJLMAs/hF2cqi00
LDNr4VORFe3fqCByNKn7/Z4Mu1ezvcDNNCrzOUQnLgzSFKFQRMG96e05gDPN8Su7
Mu9TlBQviUPMjqEAs9pLggy17gAZFMYucKp6TU+EkpkrkjQrlvhzY07w7jKN/+d5
BFGv8Gs+DIhMYikC6HQOKXtnW/kPlNFnS61H5fhYFUQUe5G8i7LbhhdHXPmgJCiD
EkWEP7zZEbbVHDfhuUOrTYhvl18j01w0wC1CMSXyfa2mwhRpSsIuTXa9f6VFYdtB
uzCQrLf/jT0HIkrTwZdo9sjBki01UnUzUaPrraEtrRMjGs62OOm08azW6o06zJSc
pd4lF+pn7AES0vHjsBEJXiHq959q6dX9no0YHzvx6UxlNO6aHa9nbh+UiFWcGLz1
X3nF3MU9fMiIKoPeNK9+Fs4UZ/jdqqBAjgPc7gXfrMtFS0lvRwwsiPrKzml7gwfS
2t3vKqhRq5WpHtlUgJQrXWLFy55/wGBlZT6pnIZquGuzNU9BNRffzjaAxCEEqcov
r01vhicMUAyKf3Nl7r9952aqKoL9OuxaHzBqJCPyx3aGaVrhEG9LnuxdcstsiXe5
Soca9BCFbM90YVv+1QHwykwMO3IH4YgK0DpzmiCCTURONemg4KBGddZwheHfb1N3
CQ3fedPvyQ5gpivsSRuJF/XGifAh66WJdJeKnCuBdZ8MZIWRkQ8ZdW4mG2tRaNH2
g5/IHwGEbF3abPcYfyYGIB1tkrtkmBPyP6ZLuJO1Z1kxKPsv8GmIrs46XxO9O7Z8
RHVxBbqh3mVYcj9cF4vvpNxiAQ6OPVrk6c/wpdjP2CF+v1B+8yRlXlrmPTkeetOb
2DrtldEYhowEGECJ6RljtMkkY3blrTO/0WXheybQJO+tb8Br47izs/t76mqSmlud
cMvUx9bP+UgSat1VTzM90TiSHM8RtD3UzqaXH+jpX8jh7VH0+mL02qCdN/Qge6pK
7RbBg1FGxaxqHLVhXYLoaKsrwC8KwfYay+Xj4mw2t2vBtMUJnbIrn4yK2evg+xeZ
9hrtbXBapkLiPgv/OYQyOg8ZNvGtLtpB84lralZsj6Aaaoou5tgwl2OxGCOFRCnf
ll4FIoc9dnUmO8GEwPbi0ISIOq0Jh6oX3GgBJiMzO9dD/Z0DQSguo0o9XIhkep29
hQV9BpVQ7IOutIwAfNIhVnpz3cHgrzQleVz1TezQWSbgq/jfULHYcd+GZVTgkozh
dHy+joJ53zyxUqlQbQ2w+suFAJ8yUE3JhPL5hKxetB5mgHHUvB0KE6E0FMJn8Sgh
MnuLC/PunPOjFYEBjibZg88lVIimtUz+rx54bhACkXTT8pFOMw2aPTnHkwMXq2FL
xBfXVn+TuShCRJymhdDeGh3hOG7I9yFd1jsXdsidhh69K/KnRsdJ7/ouVrHlPaPv
ntZaBHEjaFYNmajx6Bh9NsNvhbtci+sB8cIJGZ24cRN20JTMy4ZKxZpp+t98/zY1
ue3Vu+x9s3HiC44kk5pZM12XgHKp51efJQB71jY25SUJAhMqQ65nYdVSZbu+HDh1
RJsSyLIDvLVWTVP8FXTW1oCIq5qp+SGkvssBBnGvwmI/zpMKsRPFP8Syu1ZTQZaq
lFsXsfwGo+bbwhmQxRLc6sXdZmei1RFGg6/DB2D2p4VY3fsB2wyTZUXqoZ3S5i3S
XOxjTG5xqumq15g8PMC+Fa0u3rQjsffh1MCNxPJ1q+0hWFo/d+2qLZwCfd/4wEaa
EMN5c9aHvv4A8K8HeN569GKBgoGznUCleABhq59d0fYfjYExC8fF/oFppqbNJesw
8tbr7qvo2nEMQBaxbkLr8EIoJrauKpmhUzYANTLs1RRLwg25i5nG6CfNfcu9RUDf
6wY0krTniqZnBStbUWaSJF6M39cnQdE4SYyR29TMX1aOBklv8kwPJZDFQKhcxVYe
uKGnvMFMUeHMDOrFuvN0IpZuatX/N0Ev8M4Z4Dj6vTitg4Pc5q+xqmcTAvP3eDMb
Gmqbwc32nHBTyHYl6gjETHDYkU/eDT500RzE3WEQD1pC0zi4fZ7gA9nWV+9drZJ8
CDOk0d1oHSSaD3prVGLJj0FYC3r4XJimX27yd485hSdKANfS2GJi3aMnow6IoMfC
Q816YFyLtiAI0/NdKGsicGgrPz/FUdzD1S3jd/RD48lSaKANfMN2G8GuHK+ZLBw7
GUBmECsaG54FoaOqiqgFmxhSlXenNIswCzwF0Gh7yK3dcj0SEETwJieQbxpOoBeU
M2zLTwpHTLX5dXkh3e3fCT9tANLZ/fPnSrtfLMAsHPkav+HtYXKq7iPx+EM3n7gg
mRNMtSVQrVKBz116O6c2G3GZJC7WKqCCPo0ErOs2kGDKP1Ni84tmOW5khTymge1r
hAelIJSfs7EoN7gCOc2wFFDw+C5NfR25Y/1YbSceOcqCvXomv4cFWD0wkeqCshrt
fgb8Mo39xy5pYiFyjtc+ApQVI6NpBBtAsD/2tmh1KKzcbTktIQo8s/JkhBY2hyCC
nj532RmAkPWvTBVj3VyUFWuP9MN3pxqWtct449XIFSH+NPotXcUfFsWH+WWVi1tq
vuqEfRVZqj5hRVk64rOzCiSDXpdIMb51Dr2c+DehEqE58NnPcVQz/YAyOKbIWk36
w+PeLp4FXFXo+I99bvPprz4FRnhC07A4EbTlKSiryd3ytK6YvXVXrgWqaIwqGP9z
iLnqY1hDspm4y/Nyi8iTR7eBJOAQmbxFt7SoQxqsTL8Vaz/it77gtvO5eC92fZ/M
WYzTPnF8sMfXPRYhHJUjgjgJ3PtyAGPK95t63bcG7o0qX2NwdR7NIt+jw+gbxnDP
xiweQePlxviXb4vm6yJRP8fPyzRxCiYUAX1+mKf7I0Gu7i+YyeMLC/OjKT//RWPW
shyBZua99Y/DiQx2jbhiPPkOeNqSuCSHEHnJY38smbQObP6SkRaPpAIUGsjAR+O6
qjrrvfgpL93XZq8yubouGIeV0Qng9zqHIHdQVz6HUuxR+SL59+VJU83qdGCdp5qg
e+XS58hTJ2A7d3RobW1pFZDteId7SIIbvq0+7OJZ619iIqh7T7QUFE72fv0fjQf6
P//nRObRxBfBg+qYVJZwkUHZMoSt4fWBOQ0mlU773r+jA8XifuLjzA9kJS4K9xzv
NG2q0o1EyDT/ph5DhKslpQDXfq36pur4Tbdq1JiQ+tjj6L5NnBtV1qlOghRkFh7k
HQCrWgMmzSA/RskFo/j741AJhL0D0b1Bdvwp9dkl44+a0/g03HjO74niGQ+XAnWQ
rA8dEzQbs07vcCQBiDUFqosQsGVpBosni5ISrPka/UW5NXJjJEkzcbX661tyndmz
wed2wQxRNHsdzE9TBN98emnEiJBOgyD/rNx3sbEc4qAYJls3ZfZZs1MzL5EPJTwg
Qm7rAXhbCSAXqRoK2SyErVIto2iP+gs7Qmsm+W9aXmmunSHSzaHWnZHBJxu/Ezg+
RHKNA8Q/lnVvTrLIGpaXSUPsjUm8ei/5XEpeYHrx6Jsj7AZuaSN2EZ3ggn7KnGhe
4KTa3hYHGUaDOf8E7LXcAcCRTIIbElbdfA2FfyM2UmTYQWAE3ur3UI19b5BBvU+/
QUpO0MZGyEP0DrmTkXCAqe51X4yUNDIevnDvuWYgyc3MXtIOdO1zpEWrrIvx4gcr
HYmlanx6iRGdynlIItOqDHfl6IrMS027315LN7QSUw4AdCTki2+RRfbXHxzU21hx
neLX/WwK4N8UOPawc33qd5pJSFRBo+gCSYmApGJHVFF6IPtbgPMSlYAkb0rNv/vW
v9vFoIQHe1u7gHYTrxynL76F/LZfY8kt6jk8bI4H5HOwlYCWa1byRBUZ6KbTbTpX
el7OUi2Ef9acAk6CGyYYLy9h9KTcB567uNAUdebkWxCf5DjYE/8ugkKpN8nIOvSz
mZAI+WvrFF0ZRlUwe4v47m+2NsfapmtJT9fH/rsp5HV06zs6kxXHukITOAiV0WjH
Z5rMsFg6771xs2G3CEKL1o1gcsXjNjHDXEZycPaE1PUT8k04Wv9eJ1eTIi/+0MbU
FVZBhJyXgD+2VAVzOnqXlzKue3MXj47M1bT/W+cwbawOpRaKNGNZIXrdrGCvb+1N
sJJ/+jVa9kmHJQ4jnn44Wq2QRBodnICXx8OENrmKJ8xR7LvpMtzMl5Sc5iwZMO/m
7SZJJzmDyBDG1JpljN5WymDQLqAUcgju2zYq70qN+pma0KVy8eQsQnGO1R2VHtuk
rXKLqFwuCzOMGy+UlrBA8V+B/ly5fFT/OUHHeCBHE3tp199iiynuWxH+85H5A5L+
na0P0uVWFmFrZB0+hmGqVL3977A+JfYrqa1xy0uTXxJva32jRsWXiH49zkt+G50E
/CZKQMQk2VsgmnjZ6pgMeb5GDw8cEElszuVsz2nwP+4q8jid8maZegA/kCgFoghm
bwNnhurzWHSxx75yxcM0xFVvH3fJlaqghxlFpUMG6sccKP30Jkdq8rmIWIxj7qaY
sphUmQJuYTp9JRtonOENIgMJaGvZZoDE0qNA+oqfadI2aiRg01jwg6vp/X/pEeK1
spkk884UHizD5mnlpDaOZHZhaQ1xEwRrn49fjzXqCkJV1EdJuQ+k7ocxgTQrwE2v
0MsdWmza8wf6bKHOz/gjnlBP5Xws9xYkfD/1dkE3qoca+5y7K9bc2Snk91IJc4wa
ubRI6I5dy31A8v1grlKjMM79wdB5COGJest126/c0gb0wm+t6Wa2yw2U1Jv3qzLr
ni1Dk9A6ISQkObnyy/zfxoq48audbr2zwZXf7VRsB3dvf30MMEGpZphjkE6utvJx
sIP00bkBy9ZoDvVeQC33Fl0gqtM/F/Ois48/vCkWZY54H3hgk1k1wGzBPXpa8rLh
48coTG3hHtaipEee93SQMyKPEAQV/20seARpMwnWKByB4Qa4wXJzE9dQZ6imAMHP
GOa4L83cneWPGUDxWTuThuFgTuOHf9f+GdPIUeJsAVAYWKzzdMAWk88aW6oWiAkv
cDGeD3pe3NdQKdMpivwcFTLRx84+vA2k88XHrxwutUzOXX1ehEKv9NluIg0WDc46
mkouRxQbai+YFaAsyRAzXjomSgCj/ImmFzu83I8kzH4wdqqmuPbMINKA124wYav+
2WTPgi6AttflS36+37iLbuYWWejraep2u8Hxj2EnXYzLPFLhr9f4hru9eVeV/89+
zl+K1RmJjK7OL/LIHFqbLjIUBCQ9NXwBoNBOf8vcEhQfhtFHkFq0UXtAzqw5Ykni
/I17wTa1O+5oQoGsMQxk5dLI0S9hv6i6S2qF+baGwBjKO+OGeTWXIF6GX9SXqk77
27G2gLctJHlHu0JlbMlsPhFCi6Elq6F5wZjR4T97dMJzxYqhnLH5CFwEPBaYePMv
Ss0k4PnQbX172fvxZBiOQf1nUPGhZf4lG5y1PUz5Xoeboz6Ir9pHjMc8ySl/lYEI
8F1G/5lLcQFAq2tGN1deWsb7ejB0Ojht+og3tA9k91ineo3i3HLNm0RKI9gdn9YT
HJnN5r0nTbk9iQpZJi5KyO95seoa48iS1W1QyiCgKHCRWRwBSMM+zVKjuIYSbM09
NNxjCJP3QjrtXWeVXryJiLev6AQ1SGcF7vRk6fsbixuQeh6ke7DhHM6FyGlc/e3/
1MhVFFsq4rymywKmwVI728YYo9q7fn1o6Dw2npc4j+7QKgvz4sSc/RpAohaSQIqw
HY+i2UnFcg/7FIsFMtDb/dAp6zTsW+WVZJo/kXWf/kylJqNmGnbEyITJjLA9njRg
bpbOsRz1N8WPVi47JCvd0ihC/4IB1VBR5gdI4cfNk+wYA72G4SrJk3I6Da4soKje
eBFRPCZTHubikvbmiHFuOJpNa51q2seNITkC+70DGXrlvx4mu3JuO2b8ndtgDQH2
xhHSZ2QvJ2GeeQLSW05aq2udSAr9cb7HP6OGOw2OaetZlR9uRoHle34WE4R6736A
729vZNfccZ0mAv2iP5SuVJCMa2Tkpzd2tUrgHOepiR1rlnsvpiOmRE79uUZX144P
7VmhAeSbUlK+IfWEG3wPKTN+wtEX4oC5CFytmXqCptqQXSh8GFGadKBrh4aSFnlG
bNBBNT7I0wQysL7CbG9uBC5c6liFDHQ/Dw890dRweLXFBNV/jxTLS6CFwzvOnwmQ
j3IBoUr+3MTL70iLsclo5Px/uTR8WFpysE3sWh0/oRZJCY5BIY0jqz7l3H7hNiGt
Zlr9DLky87Ullt64tm3TaRRR0AvAvPIEOC65sxc1+3RzzBIg3DzFi5y3ng99jUjK
dhDeP9Jr4zeeCGt+/f4d9ry0PAKSgIiJ3Ay6U5jZbsPXI72QbBkB1o+WmXdx9W6I
S/Tl07z5/BvptsJgOK5uuU3bOZ68w3fhED22U5qQjFiHI4owi7BeXGCyQ9ezDeyC
K5kiCRVQlJN3FSLeokVOVhyGsLo4eEpR51eBgoYY84Rj6vF2Qi03l5F5sNMXzrYL
GS91spM5p2zxQYfpd3thST6BVKBKOOAgT1Itw23EEH5ozV3vvylB9CAEBNcOG2X2
Qb984+0q9DG2ND3UC4ZV18uhwpsy2yngN9XXIn3MgE+R9ODloEtpUA/jodggeHPT
9ci4PZ/5beA0fzmS9TeRgNREORkqQ1LxnK3bZfdUcaP0AENY8IL3ow3L8HW+uuZ4
T5Fx200Ceeh/lwzIU40JaGXjzVNNE3pDQRuiTghBvSAB7KvqXa91lnMYlMxHEKgI
3YZ9G3RpTRLDxlww2Bt7Ltwm+fO+UHb4xhMguMqATVT2CGrsNFlQh4FLQEvTGsl0
WVqTpDBzJIBkGQfpGxp959Pa0ezZRL0X6RBTb75AqQd8u8faE6ptHa9XuUiilNkP
rb+uldnmoT4VhLCJLfkcn2yun9d8XnBJBeUB0sQqIpW9eI0wIDYNLqQVoiwidSjw
cdaJpa3ZUpmb3Ht3M8jvEXa4uJE7Oco1BfeogeqjMVxG5DAmpXMn1A/Qa5Cd5fdB
W86bUJFro8insVvKxbYp8gbl6rp4lRSWOICH0c2dBVHLYlD5u+ots4pIdhupaVHC
rE/LNwCgu945HtCB1gWf1gJgb4TQ5EzA8y61XyEpPe1LZYToREw2FpN0IYAGDhFP
xWxqIwL6TU9nSuLrvuiqqJE7cNNqvvoys6y7erILbLPk188iVD8DWE6qVG2l1Zt6
9MSaPdzQ1HSc6HVvA0KlUGxF6lHrFD4AvtvHU+7STbMtVgFP3ait0C1hOV51YCdi
A2EPwFI7vhgCc57EuZTjqF3ojja9cSsBv9L73mutMu+hubct/oKkr1AFFINQqWRg
EkmkJJk44j2T3J/3QQlYSqQ8sSrSB3avR+UBdu6wioGLFe5XFg4G/aXF9ncI5J5h
09+EgSUIpDW+rm42FYVE1hBPTXRgnWxpT7zDGcFpZOBjf7NqG274zICzxAIgi9HP
j8hY8StKKEd9+sA67VSv+xMWwKUMGBBErAWz4lfmHWJbU6I7uvyS8YQk9p9fYKd6
ivEYHQxhMK0KCJ89fsBOGiVs3BCayM8sbleHmI4smFER0nmC10/4citnvzKKh2MG
2qT8Vrd5fT3cFSLN4VkuPQpuLuaGuZKja67MJjKd4J1Zlb5aH/6RZBP//MrhxiMv
6FF4VcOrpzEQtC/M9V6fYbwH24tyUGlSEzsxh1a76QkaOvMeUGdqt9z7swbY0KnO
frOq4IKp67eX4Vnk1CZBda5isRXPKhrOGyi5ROB97Nm2wEUuvjsyRFnuBSZmebd9
l5csrcYCvfu7UJ40L8UdNUcFKMkikyYbDHP9jthGxH1Ktmq2OzUBT6m6+gz+jGhk
dii7p7tBuo/8B2M+Hlgvj3B7SamxKHS0pZWmCES6v4aTpQkqzgjr1DCFJ9Lg0M3O
gDiTzgVYCZNTIv2coGdljrXV/fsrmhQBUwzz6InCzQFEUtahjJw3f21xi9xkL75N
L1/t3/qI07Zng1TnfOUKw05Accy+SXQ1LsM+RAjX9wmNA52df09ETUNmPoM/FYj+
GNrOViEIPX9u5pyjrwoWwmNguT2CqPFm1heFUZuuPVh4PqgO9SYyPqP4m9cphxYx
8UBmssitJAj0vMnifSASpSTykn95keeVcnf7Us1YYTUstrmPWaLVKxleJhtQUo7h
3vwxeG3RSSP4JJ0TSgQ7g1188HJE2oe+SIhvB/+2SDNRFSyp4OZkX2yMLhGRsgQ7
wsqR3lXvHxOlb3rDg0Z8VE9r0y9y6BbIolvEjNubYXl2BvlzfYgQeV9+smknXG5n
CVFthEvv82bGRlf3XAaTki7PTL1kn6PeNWmpudTXvZi2lXZdVO0K2FvpIns0VNEy
VplVZ2zzvU9sgdIMVLFlqw3AyRtNOdWijqvIFqqs7OjMHvDWRWbRQy7arWSfWqCn
F6nO3yXi3qKHMAJhm/G6buvojNt7czwAOzod4VhPZtXA8qlgDz1vuvrGzehVtRux
UhFdlF0tO8ZdXATueDPVJGS1o9ldHmrAp0Fh1xHSHVN15kUxS4EBgzSKqPNKTGLE
Wgrbu+SIZi99XioHSZp9/kyKyG8quYlj3O+JKy2U3iA80H8Q7Ovua1Chy1mYn9A4
+Fy5rCbCvL8vglfjLPTbUZOj4rFnPUSYEBi6KwcfRznBeassZiibvbaSEyo0Z/Nl
j9yquvRAIf7kYhuC7l5Kw+k5UZCn5Dnydo4vlxrUa1byhlbnbXXR5yx53Js33zyv
FkcROZ8QKezcP89TsOVBm71ioXZ25uusZUrD18W1vWlF6LsP2LnMZFIhLm3FGgDN
Mk/5NB6rRV42YYqGv8r0cDzNFT/T+T8hwn2faEU4ea9kPMoSrThweFxIivR774IU
nRVpk/qlAy9VvKdAGTQnukFhSFs5gYiu6LLj/jOBOWgrd7rafU1LW/iTPRhPHr/A
ADYm2dhcGeCNVauAxBmW3Q7X+wix9jC3AQ/6Yy6tMZ3cwA9dTA0WEjYUqIUQ4g0N
bd8QDUhErKV8MRbkZYHkSMgAIuKIiA3U9Q5KTIAHu6JMeg5CwxlUlCC7q75kDNn4
FMxQvpa+bL2PqKl2Bd8+pdeVcTvkwHvwD1OUXis0oI+fIcVylAZadTf8EdKXt2Z/
lFWmwDfSuv2TSxWU9fudrdn73qlA9I61marQWB8QEq9gZMwIevmjn9FagJWTrJt2
TKk/RtorITBK32Il459CEd4wrdcZA8lksWYuKpE69uQVJuhBQ3hNnlGTwldvzyfF
LqkFrkapSKEM5Bey8kfNq8qlLNPHUue1bg5iW0GXYqMkKrHb0TF4jmRryXVGmwRj
zjECAranb1f19K6OzGDkEFHffl5EPpS5YqAJYl4EDQfUg94oTRYGr0y7GN/XHmVM
JHzT5m4oD2ESbkW43QDvqyxtjF1EQcQiqA8+Z29q2xTqz0jWN7tLMZpFmqImidGV
E43FNkxX6Tg6OlSFMezGwxID4a+fR0/8rHg8EQ0GtdhCnkUUqfQ3wmX8627mRWCq
tAE6P0D82DoQeXrB5AX8P4BZWXdXkvb6yLoEUqKyiRx/i9Uh9ZJQ+4o5OMdCUo9d
gF++9Y3EDTsFVPKcWJmAWQsalVg01VKMopCboxsFPy42st4bt9yVMFmP/8yv8nDU
OFcEbIf3XYlkq1eQ8Hk2Nsz4L2zEKQc+jVabEICPBfObuKVoi1JNgXCD2i7QIIkV
hK/7thMEvy47UwxzLp4aD/77PJXMq1GSA2WlERTqn4w/crVpc0QD47uNwGde8H2a
0P6RU9HPQ8speqmPIgmuLKrAX8FbVIkRBvTcfllcIdyv3XQqurecmQ04OvLa3BYX
A3vaYT/d4opER/cnsSTsp8N2ytBh3mB7qs19u2+ZunPVDeCXwikA6l/E93RRh9ei
E71jg0lH4bLAESkl53p2nkDm+Ar8ZE+Ls721G7Dv/3nBA41jGWjPgsyh8nDI8GLM
+uH9CC1MTvIJ6VxIDyzBGBl9nhWcfWoN1lbPO43/tijfx3RnYltBRkerFFdqtRCY
AMr+kvlFMAyQJLUkh5+G2vta14Bt68ymi/hlAmNfHOzJDfF2T6nS2syW0HoqSz57
5NDeYDaJmWtVDWsbYr3UUHKBaY4cJY076tGoNNN1nGcTkICidYaB/oL+7GUXFo3V
I8dQ/HlzJkjnN5rVvzOjQaTsJaz7KehZHofrj//ZdXImevoyxSuLxVkM7XyKzM6N
Rv4xGStKu6kRuIUKFvUPWKspSEpLGiZy43wdg/SoP5FZ3qcS9ISh8drGlE4UB7Me
ERnd4ITjpixSxlr/TzcyytsaxtHXwtg7DPywlF5RRJSvrGGAcpzw7YPVEJCyRit3
T/OAQP3yXHQeVMXDCLGP46gbSjM2y7oUPGkbZcTHJh2iIswWfZdYaZ31Ec38uRqR
fxQCXrC9Du4TJKhdUVexlrTsjdDaK5o6fI8s8gMYGeymDQU1+Jw6/vmwE0jnQxC/
2YtT2+M/V5nDXV7a2ZZuVLS1TSM8WfnPWCRwuzympgRtWjRARVszdnL1n1Iis3Hn
asjVf7JQvhDVns6NL+Rg2QoCZgwRLtEw3FpzGD4A+ekimxXRWG5taPgV9akDiKqG
XMbuDxyN1Rk+c7sn0nGIGPr6VbhxkM/SDhy5dnd+fsYcJo8MwqY2jZhmqKp7R5HZ
DedEQBlh70Ve/tDrWgo5rGOjSthWYjVwg9074h8q+B97mdYdBMh02rtiA0bWy034
u6h0se8rlKjdHKUxSZ6YRpcHhSNU39sobFB6cCly9zfHM/NhUY+0kYkofxb4O8OK
hN+1tZ+OOGYdBISea7F80DN3XbL/E1SJ+niv72v+JaeCYj95mHS7312PlPW/dmEw
UFQAhyLRi570w+VKuKJ8E7nLEegiZ+ocMqtzwaXrvFU9RZG8goc0MyM/fUzfHgJX
VtEnbKc/uUH987V9wRUnGFGiG1UBOzw9qmKeBwxqhWly42xmNhm5HAhpW6331p3j
zBafHQXrNm0fMfFnFFOn0spA0UBKFgizbs+UjNKvsM1nTXBxS3PYc6YhVmzCQhni
Np4wWre6xDpN3krAqLOyw/lZYr+6dlDfLO2LZvG6UD0Tj/Wa0+hedRxK1G7m6AhV
r8yGlL5nR54o1rhUeXFsa5r+98cPf2/PH9o3npSItMPLKjXWTl/70jG2fwV5A2uN
JzJmXBNo83S7cuKzyJ2v1xxYBnTV9QzUfrBSijIOQu+lK7/nmdyGP7epYasaQSAL
aJ88Z+esptM0H+TGtmVN8ceX8hiWVbIRQEf2Vrxivy6wJMXAr2PaHoJwG3Bxv4gc
N5hnF1Ll8cX8PW8cqLjTR7g0YD2Gjq58HZgt3Wwufl4g1PJurQFQdRfeEkXr5SXi
UxKIGYiF9xUZRq6Y6Iz6Y5CUy4iA3jG0jfh8QfFj334tFB7duh/WGfxlFA0mpSF0
WC7jBlODDG2LXkS1kmu0HySCHYC+wU1k8sIEFgH49abGCyAbCnEuVoR83wiEE52w
+Uv0JPt6U3MWBv7Z73q6mP48dPYruq0Sb95QpN7iLs24rBI4VdbRbQzr/4TpmX1/
MUgZa3gtH2JO8KVkLv2i9aTP06pmpNIDC9Xwk5wNYMbPIW6zFRr4qYn3StZpEnq9
EDzMSDKj+7YYfMifegqrfN+KX4p/YZA8FthqTBKbc03RB2R2IdcVOn7bpNmrPZOO
OIwh/tiCNKe9DnGAVh8tQF+f6SXW/lLKbEuc4JPnOCvYu0dmm9wZMrMyjda/grYe
62tZ/eGVLuLKLIFM16mU6iGAdNc6cOsJgHpx9y3v3eEu4jzrX3euXZBucrTA846g
gb/AH740SU0uR0VZCH9Dxox+LWPhOWPZzxX4cOdKBFsmJgxrRSl1ce11XqPZHkqY
n/uwk2jnuJ8v2fz8AJch6TxMNdRhPzxmYKXk6as+pFz5gA2TrHYyAlv5T3HhKsed
lj77Pn24m4nh0I8BluUqu7jYBonUB+nrju0G5VaDmqS9ya1Cv6hcMpTW08N/V9yt
OUQ/KM6tpNf5AwDoO4CVO5HVmPHDnUqzYhYgN1bmFQUzfBCmx3b6WmSgvd8OZz3X
tnrvkD9IKF8VWuyh2tpVuYrctmrQ0SrZxNP9ym+KcDm2xj+p9GXmNr6VVhWhPTop
Iq2wT9Z3x2cyQCrAIggbPmLxSS9fPXLIJceuPQBykBH4O2gBsVOcxMcSTPs61NZ4
EM51ocSgCxLGOW0JTJNwqK58JgYREIZyB2QQXzPDd7ed6kh1U0t9r3ZRSx/q5R1T
Qo/ZlM14p/tcuvB1+Mg5zSuTF/bqTG166coX/qSS7bk7OYBk+YAqQEnHaBHDNYhh
YTwHCtRdLHGcqxSKJJPOzfajGFKesZ/55CggW6weTv8w4Bueh4Ae5DAxLiFw14zp
GF2Tvto8LbXO2XKKhv01vtegSmtR+yfWjZyzEclaZ9zOcsce6JmptB6M/fAAdA/N
HjHSIJlkg7AOHE14WOS6c3H4BulzARmBwyzLuwxI2polRq2Fi+jVlUjlqj7AjozA
Pq24zDQ4HQqbXDPZfRhwE9dTXzlyOgFCz5EcShmZmOnu/FAP8bZAf4JIjtMEat4G
n4W8ZtlUr38gSFDU+0YcbFtGerxedXHmZSgDU1vX7qUHaQMg03yeyiHJwWz2I0Ll
Mz/T1tslozeWYd4+dnTekOYrWGoxaiU681VPnw+A+uEPMplmQuqgk+Gp9+X8rgqt
JVwqEQUtR0Ir6kQ9Oep2MGMwnDu+T95YnPPh5F8NONJM8V+X5wg5MzfbWFOPVkOk
ln+nZ/mfeRj6z/NiRfspJnZUoA/9Xq78W9GKzkZ1Zs/q2CcTfZOvCvWZxu0Kf58Z
zyPxItQwuzBCz/H0N1VJNRg2x7BgTtlXxKjEMGduR+jMHoQWEb1dpNUp1iFpbl7q
mhQJymufFE+SHjwkxAVAgsiAeLDvo6O4Dnxg/yfQSggWvtXloO5ItdaXNmDTHZfA
2XxW9qNPCzPbrQj/hz07KxWInSskR1iNVXiDzFfhLAuudPCqQy6nXUPY3GPoSQBX
I3dO42hldbU1RuSAu0haru7I9Q278xx2SoK5N4GmwGH4Le1jzVOSw5sMB2FFrdo3
E2uYnDio7ZAD4u9EyJuRQPGPxCtnaO3Om00dDVcCC0CiliJu4Kt3Sa9i9SJISBlQ
KzngqDcQmUK6c/NY/m6hlzpV4hXCtgrXYQn3zEzZUEcV2m+DrBwE2mS9XY4nXah9
aEaZ8Xfn2zPjF9pvBLfG3cIUYhtD+2DkIDQsXH4FobP+tVSW68Wy1tRu4odmi/6Q
kApGQnjdyMas735EwviQGl9etInyBO6+dY3wl44+vIITIRmRPTwA6gMrWtncYolz
4ZILXgdqS1DU9h9x8SuwKx062DuLse16Jmv0L/yhlMpfSpjCJnl3H++peIT2sYz2
LvfDPsgIQuHK7EeunhTXdBwqbXPXs2v47waomZv28YF9nZLDzzh1PZ91x7VK7ZUC
pAvOWY4Aea3KwaLWPVneIWMw/Qe7SBD3YjauJV8YC6XILN1SYSARd/WsST4LM55G
oQgYOnUr2D9S1uzU/ZnV3VO1YZaKbCUraJLbOPRsrEK8mqoYVRziF8++nLpatvDf
KR10fVsjuJtw7r+EMZyhTKwhMajeXnnp7muesXqL4r5u+k3k5rruw3ZZhlV5sJ7C
Chq4gJ3iaADk83znIYGr3JQaHZ2h4GXwSahR6TMpv7uAC8Xsuuwqzc4goHzMibEq
SzC5LQmuiuhhqDvwrwAm7aR8ajr4bl3XmKJfnN4gu/KLbikQzf+s42FHqJiARTGw
JTi2J62HON7QrXbCXRpy+jOdgL24PGn0GPbrB0iqegiQMWxiHMml5V+leW52q2ba
ECdboDn1SEGKJgj3ANqUuizeE9HBsJyKgPugFDHcbTmXHjXR0Ua/6jgXUwpGW8Gz
vyKC/sRWx7D4nHKhVxLX4V5rxuCJlvTW7kWnxW0sCdyzSDPnUAINmd6Hj8hrjPtb
GjSEBMEmvSqJl9hIR/BFOr0ZamkLrn7CPyTPEiImFKDJmhkf3SVWly8I+2DDKxnY
wVeBig0pIvtooGmp8ka4iP9/PUfYed+sprE8blPFGQOEYxrmgtb2BAwUxhGi9akS
7VXCeiEBo/EyF9hKS5pv0TeYQ4sY6EukG54I3uDLnp4EEJSh7awnZIaU41wmkoJ0
mWGPkw6XahzQ2WxnDXiM1HWwxtRs8iPnVV5pucdsGRJRrWtGycY6FnLZ9rhiKl64
GEbejE3mdHORsPOKu5KXf1OrQ7x8/CK0MmTzVfPT5Wm4ZpHpJCzcgV6K+nmYhMnn
YFRzqwRNADYZrP1n2aqhTLhqci7ovGuld6eGmdp1GG/3IgcIVFutji5cKssbi8+e
Nq9vmi3eIcdvbMx6Smg3w+VGjrSxPISZjI1b2P4njdJU2r/ATDnvdCbi20Qp7gEt
klDDZgFw7md/iexP4Q7VBRgd9JZngUCnAcDw75PTaWu1TTX+0iyx9Cp33+9ysYMd
b2lsXm2w+o1NvUT/6Q8VQ4i/GTlVk2DAF4XQxFSKjxf4NptDq3QGThwVY6tmmEKg
tvzsbzhYHoDWzReslHUEfq4fWdQqgee2tZQVI0PNkx64KNwVADe+vqv7k2CsBbob
RvUbrekQGFgTfYzDl2RTg7lluhdHqtSeL1zVjCJDhJfJwIoTeplxQ4a6XYiGfj4Y
e3qW2l35WyVAcXfkkOChTEGcBoinRKkFcRP8tQbO4vZrYJ/KKpMzsyGTmAMJ2SR3
103081TBlDJ9VOGYrZrKNIntPVY4inruj+BiSAB07WO4FOCngzejFas4EA5b7mTw
vjPUUuqdBTUAPcgJRWOpvAJtwJNaUcjVn5sbrx97nzGWWdc1r7XAFfx3zMZo/R/s
Z8L+wIZ4uarfZKF9jBA7gbgwd6mZVtzNL2Lgn9iJqbgbq+DHPdFF4BGv2N3iwZeR
tO7brtNoxwued2sW2reD8RcNySrroSkZwnXwGSkKIHx86vPXv8CQzrXzHwM5muR9
ntYGOVzaGXOOA0hCpPWG9HVJ7fIM1alVcJX3Z1NqM/INrTbkXNoyBW31i7Xx0YYU
Pq78IJv3qT65UZoISp+/0/gyV6mVnoRpRYYZ+h7OHtkGt3NZavk57t/Q6NkKsojg
kllO9B/j45qKyTfdXf5zBkkaSRyhh5G+7H4Pg4/9pW2fwYtuRY63QQr26vPevonX
kjnWKNbnTDl/+JpmkaOL2WYwmA3/pWH+sLreXOxZNbWC88RhGwxZoJVmFfOqD1y2
FAex82BJ8NR9k6qqsgxbA3dJIq2HMMe9VuBAAHvUm2kttTAwUMtOTM8pB5sGWFbD
aiZLG4c8VQUHx4Q5Df9E/aGplkCtC/IhfoZFdNQg3ziqTRVuk5uy+WQCnnj5EfVY
WGZ1+/EgqTOhKaStntWYnGe85eJz/1vh6bM+Y69sPjsce/gvZbNCgw0fxKZnHzYz
89+lD+gwxsDLUHNXTxFOlCoEPcjDYv1HERTMOlkPcZK8jnSm9QJDBNTRIuKA5i6R
3No5vlGKnbAjE0DtSYLE1W3KPN/gfB5Ms6uaV52/DI0EUzsPszshsCQRo26Pesou
0r5e5rHrcO/K2mIQarYH9IFZEEFxKPDh6/KlaBabRHN3fSMqS161lV9eMixdIF+M
+cBo2dQ35DrYci+TMGaLXVKZfKOEek3FH3ZSMfmdqjcs94GkE+hirfBI0NPIazHu
DMLIe7lm7C6ydEuFhEoARWlmLLhUk04rB4UmiZyUxEUKUF7lCjAVNvT5F7Vz2X8K
KeY7y/0I+BIZlqDAlYpFmKER1D2gO8g6dn/kkg63VF1CiifkQASCxIMVJYEPbSZu
1y8h41WA/N6n6SL5yih9Nkw6nscyPMqKwkz2iaMiZyQmn2oNhwems5BZjkhXluaZ
4duS2uDnd7ECCjR9uWK1JoG0G+wJ6SPF033sTIe4MWSmlVjvCHOByhe6UBufWcpo
kahZudUBcL5jMccvJJlU5xy96ByhFMfZMuhYzu6lWDUDvefzfvZO/F6+BCAOGLaI
QzWczA2T1T/nkGis9KNlidNHLhpGlpxxtSgFXG1KXmzKcCqruygIjcXWN6RRRdbk
OG9pwLUXmR0IcZCYlH98x9gVYD85jPiWBsDNiuhXo0Rb93sM4q6Tc47wwZd3caAL
6QXvLBQ1nOXiINGnyHLp5Smf6Nn20ZBqg3EYp71xaoodWu2iHRmL76QBS28uYrkj
RY71u7SClJ5nK7CJY59UeYB18bfFO8J3M2QUJD4En+gb+kZJtNShxCxg/Oja8hH/
0Jx4YQhrJi+H1C/iRbTcuwj+UvGB9sgeLVNm0UGnHv52RdZov77p/zZxOCey/Nc5
HVxrXdzu6ohUR6xkZoH7jh4SmkmQ9XHNpYT0ZO6gmwuPZONKeqjyoI7k2/TD2OmE
a2QiteAPXd3vBd7hko1Q2LZOEck4tCldcl/XJiw8CGqmwMkhSNkmK1ZQcg6VaEfB
OQGlOJtvfTJt2WJIEVv0v4IAwqAXvFYKTCo4AjFlchqMr3D9lhhd+ADdblAb7pcw
oNkVosYC3KnlssRxuMMgCBbwQ9tNYyrZwQQ4wIlGSJUlvP6I9OSbRF/FwEOBsmYI
93iGI+UwuKS4etUc6d5b8J+vn2Z/4cd0lQJW3VwHBOrx3NMr2DsuJG9dR98uDLfa
J+sZb0Vji9UK7OOonxLDfBigmelfIq3gFui2Da53Oh7iMRvWc+dgM3cMZOB6WtCv
ISq8DU8/y1JytNLN8+BYz0q9abdzn5cHKvhGnOv1ilOYhMnQIUPuE4raqa8xBWNz
uwcPPqXrnOgp3+Ymwif+9bSIPZaxDaq8UkDwPaMxi+khk3zWuZwWuE+DUbu+cnp7
kR/nTiqbVW57x3vBc4XaN6kG9jNKQARBZUWM/HPAkiCKZd1xZdns/PE+kR2uLgy8
tNPtYj6SGsI4iwiteXoRH/uly0sHSLVqKJhtnfXSLwD3NiTXAEChvkwwTm68dWY9
lk6ZNt8QUnhQJ22YKVtsnYb0PrNBekiYceVIrGc6vsZq1wL4BlPZN9U5Z8183SSs
ZyW3tQcuspMcDyTZW5lLO3yYyPwnAVpv/CLwUomFi2CZ+T+L/aAt9jGwNn9bd0L+
DVUMcW9+fPmNo1QeXnx0Z/MFk+XCNSVq2cffLchKBNFkDhL8ZhFfbNx/p3a78zwX
dOKBZopeTbcJ9k8Ze98knldCEiqpP0ejvgyLiEbesIxJArgRX/EWw4uMXNMSRRBx
2W0xFAo79Pl4MzFclOn136POL+9GWUPLVw2/34uJdhSXSaU3dR3iDy9mS7f+IvYu
tgxNC2FIQ16APMTNeZJg5v7tbJjUez9GCb/2ifo490LUTVdPxXy7hamQVzjlLrYb
FTmuyq0t/MsQeck48hJ1FcYtuH66mg1j05FgU4hUgrlvU6l+5ClqFT42n9oJjcBK
7cXQv8Z6r0ntxmTL3+xDjLpM9H7qbeU9RUnfjUrwYQpWBHvBTtzzZd3Bn3Ss4qP+
I1SLe9lSliQYgD86yZXRIP8hypfLrPaGn+CK21p3FH8Uo7DYs9vGhsDAx3UrSH8L
qIpx2u2L4JPPnGGJbtY4ZU1/rdxYaw1vvMhwpL9Z+C0W2vA0JqwlTTLYuUCPbY/o
WxOsXAH140CFb87b7mhcgoRP/hqeu9GK2gjppesqym4OiAfKW+7kdi1wsWqV6nox
y2nATUHnQ02HIOJY1BFHHkmg0qn2aPu/OW+l+Y4yKrEIGUYCZ7HmmWEqi76FXZaN
BuuG1kwfsCiMEuKatyGgbJ2FoVaxeuJsEBGhfcgh7ElVbAyFGc+6QT/rUtpFK153
X9z18716EsKio+WGtavcnoQSBdLw2FYRJCOhTfGs1dEGiQm33Lo5DGb3ZMqsJc5q
mDIaNkngZiNIGUFj/iu2/Ec+IGntz0mCRNcP3yAo9qzvtT1TPuDkVAfLl8mgPXpH
XqEbvzOQv/GrsDNPNb1XX4KQW5InUz8DI/5ZmPfD9vQKPQzoD74ti1fbylYWfFYT
C7bO6EO0uBeRsi/HpqyG0QFEZTySxSxG0vUEx/UN6v3xQMscf2uEH14a1aKndiWE
YcQ69PNQ7LPGWIv/vU0wE2aDNcFNcAgpHf+wP7e5fB3Ygja55HTI21SAjQabpVzO
wx/TQ1jp/DeCRIhc2LFRAoVNnuys1DlnT59UCpdd9/vljSCoZmavzVwPfoFBI4Z9
yQswqzZZnO9aLBHOJbLkLFvnJC5AZxKf1mG7OgrAxIaGNnhfrbCzKAj8xEiB4q5w
Nx9vOK+87pjVdHSDIM0ALoEFB6jSOFESinlsIA3blU1Opchb1tdW/RMTQ7xCDCBP
rwXRbEXUstGvTSDZgSXM4/cgnqLZ6/6IvEhKDa2c1OpibX6qIZceFi/O5bMRd8aX
vLR/S0Po8qzWDYlKOB1osieYZ8viDg2VnEtjstX2K4ecHHy4NEONdXTm8s7/PLhT
BzpoBnavPSPvEf9ymXDAYGppFa3q+61yiK4XeUzEPvGNq2X2mw3ToAqYcBrZ8P3W
zn4FcWqk/qgIVyyhlEGfedzS8Gz9MAaIWKcvQCIYHvJiYouDHDvkGRhsWDMN+gAR
qLZ19bCm55jz0s0SmbpcmkH7smeherZEDys736CGHoM47MRSeSuZSCZ4mM7bEeEX
ktizFqWjWfb3DCt++Jue13Cr75840MMEEqUs8js4mMnE3OaJ+KH1BKRqlho6P0Rq
Jn2olUJQk+iosaGMFVvE6wWKTXmK/G6h5XRlvBvefFc2VK5oV7py4VJdLEHW1lHN
3SsPSayrQDXBMT6421Obof817fLK7v7V58AVkoBIyJGW6Pf28F2nn58OUocEsPmn
rlbR7MF6nZD43BrAA2YXdgZwfxL+ZXl/Rh63+5lVnfN6Y6cGykN+CBYbs0A+nqCs
fcpMib255PQxpzPMAstpNZlxWB7RCbvXN6Bc8d2D/aPzZExiS183GRxMF/9SXz6x
V9jnZiIUmoTffUljjlkP3Qn0xU5rB/yzLE+CCzL0pdbOoMVdk0w8hlkqaSoEHQlC
hG95BW65sM80vQGPhVPtwuiGSGYLidQjaS9H90gql1xvF1DJXRLdCN1sorAd8a2G
yVmg4wsM+EXX54e4gcNCSafTU3h+lb5WwJaJphwLK1GKDFezdbXBEDfrE7xmfz+f
5g2OTdJ5verCsTKggSDzfTMBqCQICRUVEe+SmM18tHK8U+XST1R+p1Gj9QGs1zj4
rfjOKWF3/vAddXCh5JNvJglGD8wxKZcW7m2c++P00k6Kt4wK9CFLJDKmPBBVqBX+
NiqsXSOyJxl7hg9b23EXd/w6ZwpNbjmkwz2NMca9ljqo8N+XOgp9X+Vq/v834kt6
dY3x1YfUpfirtdMlYr+aNt6cxA+OYjIj1vYU9KBnl4p/GCPdhSV3E/arIICIYADn
qborB7sl7U13S/uzSx0P30Tnl6dYv8gLt8mmoOt0OQ28Dor3nvdrvtzdGWQxlce7
mxKImWv30cyEux9Rc9bWu22W7wF67R2naOeHZmDMhtpNlIf8UppYpnSZ7cxJlZYF
B/2omAOn61pG7ZEvCXXAKRE2H17ipv09YVYPW5o1HK+wxBtts4ZdmNKXKZVxGlQe
oVDnkI2iUiQ9QTIctZjC2PUsnsLx6ZkIA55lZbsY/HTynm2AhghM+NqGygr78zwU
gtNviQkb2luTLnoc6QP3aFbkoWBfy53nbd9ApZWXlEOjjcsf4TBkXYAGaGW75iFq
NJ7nGPN9feBsujMG3dMuYwSKgN60yX9+1cz/5PQmL9xvIzrxEarw2O3i+60MLALC
ihAtsZhBPbNS7vggwwx9aQtiPGE1sZjQGchq9U3OAtcZIJCdExm99Wm4lnj1XWxd
m7Tg23MAB4jKFtVsc/J7Q1gpRFgccJw2nyJSv5BliZY8cGy0yOHYu5jkXQGsHsCM
AAVTravowDrwHK/q4WjNIefs6UWo1GwWnyieereXoOrtEZz4rgJsZki6Tf4mp1w6
N2DBO5Bu9xJXef9lNTlNO2Ixsl0JjBI5x2ciC7teQbFykgGR39lqWa9dmJ1NpZz7
u3buOKHggyXfUIyu7i8mXZWqUNLEmQt4lkGPja9zd6CY71Ihr0tYKoSvKtBcTGZ7
8XklPdu6jw6goqdXPAfYEe2me0q5EPp39FHHkQ784HTIB+J8nYGxEf7f9GU8GO3W
quTSbK0GpE50I38QTaufjPfKd3ShrYEkrXlqcukJOjiPrGdUoCo3oH0LgGIfZcZk
cgioauD9wN6DhfyrYaU3EnTVdtpxJ+8S373y8x2PtCHQi4RUAVW0OdC1n5E9Q4mG
7Eiialz0Km7S7OUYKeyyoNd/LRYlv9vw/++AL/erMaaol3a36IYnjrX0eOK2AUsc
gegV5VaIMCvseF1ck4uGw2wKNdVwi5TN77g9Z0IoFqhMVc2pFd1qYBWL9/xoSr2M
QfkJJfrc3HVUZD60QWL5WaXAKicvYryqRptJBXBzf8J/jCVBDJgixcfWf5Ht6Rn9
aEm7UQ6SpsEUa4CnM40kSbLfNfjwn/B/TRCybU8k8Twhkz1nTQfjQQq6pfeAom7e
HJyeIQz/VK/DU0wUak85XG0Yh1T8hp0uSKq/m7R14P/LAInqjJS3EGNJuODQBk5D
ZLeRtwM6FiT7j9rfbPWfSf/kACvns11J/f0cVRReRhfti8M578GVyYhWaDMkc9a2
46R7uylhb8owNXz2IT4Sv8fk/Po+uAqRSxdga8iphOj3riR6WhMfp2TtRTd61zLC
B+hBEivF0yeLIvCzMB0MbkjI3KWRv2adybz/z1Ik6CBEu66QBkTz6hnaLuPECEk1
iJ9wc8JTQXA/jQB7EVXCm750cfRHKDq5yR+Kz6jSozJteS3Wt4YO92TDJCPiC/Qf
lqENmZqaAvBLMdhb5bnqsC85PBndpZNHN1zy+Z1o4iaJ2ojX76RmAmKndRKpbvME
GfT3yvR8SaavgfruPsVL4C9i5xJJV1vm4g1xHu8OcOXyYbY8zLw8WobBJYDfSBce
rahjSNewtC9wIyIm0PDJkqKxKXzjkZbVypOacNcVAYN2yGK+SxGscovXLX0x/wxc
fdO3YmPCrZlFcNSXm9bqZFhRSMaR/xIoyP73qTlX1W5t8sG2XiJsLRfBiIIYafaN
uA85oU2bgVRHLaqklYLWC1Br0dTA+4TrCJsMnBpNlLFRjYnQ76UECuD+XhbKLR+N
vebdZa/0pLG1avD9Wb2AhXMqSyB4QjxDjaSTTLjjOgkQdiR9LjivmahewyT+MLN1
Ji02Ns3h4Kwru8Uu1qYtB5pV5xjTnf04YEGk0kJIL0PCYP8xNoyIzIdA2rmx1Xkv
xRnMlZZGV33+IfRqrXrN0HOAsfnUGN705MG50piCG+Iy+PqNVr2uI9Pc23EekJMS
h+WXoXcp7ZOCaR+3tgSRiq6er+XWx6T+LhHHblAyvvq8S9VsseNapxXkGP/fXgfx
ucgi2hq7SX9U/HzbvDNS9DdzVY9mKOdpgNv5LCIujP3uPT2sKpoR2FNs7Qssx388
Mj2RTQuD9SxI7QHRHZqSbeonxak1oIHPGtoEf4No/jZaTUonWmkzYuHHzCVaNuCC
xv9uag3LrzPJ+IPzKjOXJAnkroBfXXIZ9Y6lSsAOcPB/e0azHDYmDloONM8QuPJf
Rm01IZTbnbup+Te6bb7474sKRKmxdGZgd2TkI+1SMmaSc1Cug4vxZfi+0YhtdpjD
STSa+UICrJJmqe3bBw25HoRvm+eBZH1E+3wobHWCNJXJrIqTw2TZv0bKvSQybZEs
nUyQFICwSB16clrKhvNpkeJ9j8sjT8sxfpAIwpg/ZRoUwPA1GyylrIkfvR0ChDnB
fbwLBtk7FVzBZg5CC5Ei7uYazTPTZgoKVdfuOCXR1mKpoZR4hPEbvMIKeGYRORMA
U1Q3GlFfYS0sTshRRvZz2KGtWfAeHluWCWnXBcjU19iZ8GURJGzvbTmk+L+XELWZ
CTBD6mrqJH3ioTPSNwvqBGDXT+aZtvYniKXdZC/b2yYTlq2h9WnvTk2loe9sajcZ
yrBRIYYF0Y3iaYBgVScq0AomCEIETXUI29tMOW4jtvPWd1xDzcXrkQmA/mxDOOzV
ICTcLJ3TDL8J0BJCW/YlxxqPD6svou/OZDJx1RhIeZrGufsTFiVY9782Ghb5v2I8
aRRz6vju8tJeWvsnIqZr/Y72xVpJ31Kpx71vkeIaUo3cbUiN9FpUpS0HLRKs2vIP
t6xecWEoghtOAWt8HJzfTy1Ch4a5+pVoLC5eB73fIjE6oixukSH0vAsQMNvyg2Vb
mKpFNOiWuCSb+UY8TguoHo89DtDqqXVHNxbfpMfkEpw47L0Vsv/pGTUo56vat3qt
a+/yjlZ3rFyVt1DIsyvVwRfbI5zHirf0s/2TQe7pXBh4xXezNFylNpvCxNQs+qgg
EbCa8R6co14jgpSdbwgv0ON+AwTdvM9LT+OXYjsL6zrrrUJ+LB6HOfSorv1G/Xa9
oRHAjsS8GoCm4P9tb47E6yBIjF/pq+xkGgCYOo9CZ5HLXzGvcSsNRAJN4t74lpQO
TqBuvBQmB5T8+Cdz+zphYbT1hn9egoeFQtt80x3eTyNeyLn2WvG+I4+IOBBGzrYd
BgkhuL4kqnbmEdy1wl3tJWD4CAyV7nnZx/SZ0W2hM/Swt9z6hmPwfmksVWZJjREk
btcZJP15CzdqkngvMRq0ac06P8QTTW6NJKOSvJEnoe6hDcoSXE3KiucUwQrFRujN
6kNTIldokgCNXqWlhu0h6CLNMWvhKyNSh6OVH+0PMnKS3F7WmPYgB1otQO3A967t
7PuMKAkvLNm/3KZ6oizwkL84u6ALGu6QCamKbbfKp6kX29oUNvktTYDu3gUCnZlp
KmDTg70lhECStgzsSuy8+3cPRsNocTixa6kzT8j/lrl8E4x1jhn97Z/Qs4uKJKKm
NIcPzNbg0ktxWNzxrKlPYC7QZBvkxDJ2z1/fEAi0HBycwJsQsyVf7Iw+P4xRNYvz
zO6jYWPaC9pHSKKOgYa9uwnuIXq05JselHUAq1NGH9Rfgll39NqHuti9yUaVy8gl
EfGvMon4PzxNO4IMuuzJmDq7bhzoE4e1dnw3ztAu2zf0Vm+NdnYGYzvXqQ7M1qq3
NZGnpUUZEFSxqH5gjSTDmxRT3XyCjOsDntOW2z6w56BcfOWnOBWgp4Zwko5yhWLp
b7LY3LJIpXr8F4RvQ0Z2fUtJ+ZI9LuarMweMpJxt8nETalBrRAdz7wbq/cagME1T
45bWLa2aMqpBbbD2NB4Bbr3IEUQb6PFNK6usDqU9hrrHukgVDGgIG+yKl51Mmuwp
NK/nQ+9b4Efrf9RyvzTtUYnsBuFYpizjQqns0Me55z10sUqSAuBj5FrH0L4xWqLX
xau7UpecLs8n5FoyzT40hJxclJ5k0D+aXevoX3RdiOwkBervnlALs0urlCiotc6j
tJfPaF7RPqWuJ5q2b2+3dQqlAiB0WVYNWd+TsW3g9zLf2RlnDl/YXpcbvHSF7Uxl
FjmAlumhFgNQCdg+nI7uwe79GmEoy4lMsvQPbmOh6cjyymLujQFZSGOoHa2bXwPv
l5At8X3k1Lzwkv7utnh9CMc8GCu40Hf5akZlNp4eOarIZ5ehrro6zM0Y+9SyVm/K
maeW+X/ajkRTgdxW5iGebbYRQScSEbddVBN3CoGJVkW6djWOBFI+UHaQhKM/ay/G
PGpQDLa87MBPGToNI/z2p9IR52CEVJpFXrYwyS8yASgtswO/bfs9We8LG9qSxRSv
61rjtjmZJm73JSVUiE6lcquj1whpLPSYbDWtGOOEXsQ6ESRqVkXGMoAct+O2pwHc
g070+w8gvi703Vt9H3yofBabSLen3kMWAwSjCdzCMf4HKtI9RYdNvOQIsBR7q2k8
IDxU0g9TUgsnYFw1h0NNwz2b7SIPm6+pRc0C4B9sb9uIqXw/ysVALOcQSPsEFPgj
v+rzOC6/ykeZHzIOQbF6TiUGyMSS9POmfvPV7B9d9FB4u8weqYt+bkGjRIB10I7J
8llHC66bsAyZ5d66n4UrbcDuhgUNl5j303DkWK1xxJXdhenZvtfWs6ca9BKMhOh/
cyoRfmkIjHGwY040fFHL+d7I9ehxew0Tdwf0jjvT+tRRTRyJUKF6JJb7F1z5w6or
7I3xMiKKyLi4qTr1Lt62FJBFzS887RQnDnxGyabR1+K0u/n9qXzCmNPWGvtwAVfw
FEFp1nJ1/RVs9OZidT6U/lBWN5UL0iVsmiDHl16AU7UpMTLY07w+EIh1SRbHZ5xU
1b8+2yIbN1ewBSnPTP4kuGaZHP9zfwr0R59h/RBIjDhxGqw8etLFs2GHHAmzZ/RK
81K/LGmpJYOIzFsW9wi+f123civYmlu1XIU62gI+sahXOaOYtrYO91Jo5eKtOWch
sSeaj1TV1zN4uHj0cPBJSv8zfxA+/+c23cijO3KPDpI2z5W3BM1zIBCSNrCFicPC
Jdx8Zwld/KAJa/R7IguWsWyKOOLnsugPLgGNbGLASlGomhrTUcIoBLCRfaa1XagD
b3f45XD6n389MxvQPCWuFp7k0mGQw7gdWfzOKimlRnGxa7nU0ogyaG5M6bIamRvZ
aYGhDhl++gD7rHGJ4+4f2VbID6iMwxSXewt8FLQr0bp7ZyTlUJXGfJOcwaz/ZV47
KjsI3oMMRIPs2XTtL9ivpxCV+3GOlquq5amq+EXmVYv6Y5Eh+oZPA4em3s+JM8Hl
l79/fP6KVoKDmUAJu7J9dbcQGBYay/o74/ZwOw8m3ry2774LZG8dqxDm/wlJSykc
U0jfGSdjehMffiJ6RPbQiOu2WZpPC91PDabeLWx160W0Ye/v8ZBrNetpjDPLlsHA
nQ/yt9dKhqR+iv6IjHQGSskMc9UlAXagLtCGfpEKZlrpEZc1aXtQnaux6oOAk3Ch
X5jBzFBz0fKMmtaWhpjo/3FHRkx75H+cqmQMbr+YixhQjtnrsnrAYLukDZ1DSHd8
D2JMe2a3s+ZvEHv9SGOLRAeE5K8bnR5zXc1/dRL5AVvwJ57eAnJouHMIDqLi4umb
3LoMXijGks3QNlIlPdaUOBjC2Y+zzECJOXbIzTU0xqhTuSdygMv1mgw2d14XD2HS
LtFsfwwLeaN+04+udCjzieXs8QHXp4qxZ2mNfPK9oGTMYXLcTDuRH7NgJaLQSlBd
6OXqji7uGFlZZIMMPwCsCEuIfyCeId1mo7tARHYdOhIKoGV9NKQDQQSEcJm3vKda
BooG56DZaZJFj3wCKV9qR3nGuwP2Pew9MfcHBoxZrmpE24BykftBsXVvHkk9kSgo
E6R9DBSjQ8ZheQA4L7uZ4ZGZZe9kFJAslyP6BAa+3RuMX8SdPlXEK8I2llp2E3fO
8zTo7ErOyM02IBKDWDNV3N1UPeIGhSSvIQ1EgM+eYoPCla+meChF6JtFIi67sPzy
5oZCzeJOGbi7I/u2cyrBUQvJ5Hcq3LzUUYQ6Ss5AkH0AEFizTuL9qjEuR3yqfssp
LJlbnXzABVtvd1NB9qvjJIU+E62mmAP5RnEGCIjgpsNHGbvLAt8qQ/z/uPke+w21
FDibYmZBOv76IPuxXJRJ/MoJZkDMsdNRP4Ev3SJq0AfeXlpYFnuYwNc1On48ZdvC
FGpDYlXKa/LH2+8GXXZlLQmwxXmVSMBw87mQy0SyAgU8PA56DMoF+ZogNJSwOZb1
a5q+quFIwj5KaI3iejVBZk1NTT0kb+DVAvvcbGYgrGv3Lxq7mwyFhEaOvq7q9T9z
gSTsaZ39CpKRnA6ZyFpdaaaSpBbs6m2nvivdqG72n202fROcPRXIanhc8CGExe75
+Q/4sB8tobHF3A1sARh8fnJPfXwOYGfcakBBxGwAeJgkimrrCSMfPZzY2qLmWn8H
s7Wzy2ChreGSRGB/8DLCqUSoPKP3GexGJoKsrZ0v8Gch3zdS3q5/+qyhivfhfxj4
x6COUhVBBrbH7ow3TqidpjV83AXNfN40otApewg6r91KWHKXdmRDuPUSO6lycPS0
N0GdOdVGIJKHfMAKdE8PoxMtV1XRLBqhC5DvEL9fGOSCO35z/6GDZm/7GYobzgUq
sx/EmopNJaXtDoiuv4385w9ol9E1vNaee8ZTsRa8VBE5T3EYXs5tJ9XW0SbZKg9i
oPZ5mI0jTc2mmELBS5i1kf+hWG6QaX3r/ULVs6hDb84wKLRgiClJUwRXfzO4ZGxO
kGFIlcOUikFy9QZNBmtx94J1XFABGwJ/hRYuEAguddu4sGguEQvGBEw7H2f+P/hY
luR2t78AOEMGhpBctbodfExD9Jk5K11UJtBM+Ku5REgXXY0yBOpG+zP4yZ+4j61Z
MhAHlaubN2VDAJuf7WoX7/Q+PNz3uKDPFPgaiUiCaqOUIm4kGPsRQr6lhmyq217L
FFlq7UQEvBLeQ42QBgjFs705xApLzHfHqr1eNL6NYKcD1i3OVdhPA65TE37QeSkw
kxlVbCvivW/yXWjdgU3/ldtlAYIF3OCbgr0B4CHVxDGpMzcpR5QWyiEVTJ+hlWAp
X9uj1PpNDEyZ9MzPX1udKx9UPbMjTbgYAOlHiNU2q5TUdOlh2JyWJMX7w80plBII
7vHLQascAFQxgYf4oz7VC0nCPqshTySLLV/XBzUt2NKeQ+HbnLHukoR6L2xfwS0z
xCuPT1tdQ3d+a6B4IaLF093cAb3V8sUk5mca2BVfr2QPo7Cz1ZN6ne6L525JYs9R
KJKJP83BulCo0wl5hnd1x+GpakRmwctAxH+WsCGFtoKrdTwFZuiX2MY4cNkLdD5Q
UI12Iiqri8kKN+WrmmgK0/vH57Z0Flvy5ZLBdZRTXmFLq7yCuoCf6U0y2hzXeS3z
xJdpNBluK+/gbP10OaAegtj5MY3F6rWG/dIBtqjBs5Z4CGeYU8WG0ylzbjmpAUsS
Re3iAylUc47iIITshQnC1c8UjfUHE4ATOBi6eeQbEQxUc20tpel5p2uPaDHTGVgg
VxzGEKqrdT3TVxhixlRHnsf+G+rvLVgyUJcyahPETA+dZWc98BZNTyxNMe/qe7rp
9s6aammAOmxCm71zXXQNKRhhaPcVwevB2BGSwg8zX3BqPaJVOQPpU8ZdEFNnsjbG
nig73oHbTLc7KKOBrFbr/bQwsma3MDFtvTtlIkpo8OAsYwaYRsqMmuwQzSlCL+jv
j9CR+wuj97zfV8khvX469qxryB3W5AJYFhLvGy1rktlw68V7IhJu1yylPv6pwR8p
CKwynhD8yMFtbN0JnE74olUsE62yLNrTnOIMW/NCLb9KJ56/pPmWgnSUeJTBhXiZ
PLZSh51TtsbaHWdRUaZekgg5aAYMx/2A/lkG8ZO0ysa7KXF0YYDQuIArpZVcDh8A
95yJhtyBOjQc9Lwo/3GDezNcoWqUVfML2wO/aCrVpfX+eBKjpg+j4fwKdTH7ormi
98u9qcfh1au1vGX9rt8vllOSEVuHotR/U6VRF8hGoDzP6TYmu2eIh+A7UCTGw919
xRHMdPUP4OWb8BkMSV12NT7UMgaqLhsX2jSFRgBd4jeLCnDbjZv5MMMeB13dAvnj
nGOn5NL7u6EJeqf3ySAZdkZcIvQlxxaXVruroAXYkjrRxnF2Ql8o/uDO6qgXMN1L
ln1ThyufBH3MmxNieKO+5Uw8o0xI/hAueoMHWXf5HXjrIRQRZosdIiOlRbWOzTW8
+jLkMN5yBSSZ4mZQT0o7FcLqSLEnSHr9I4i+KxSvI8gPnqel1jx2/mhgqWuJI5Na
sOBBs33eNzvyKyXJfu4L8VVorTJ1h9EMhMW5GaW85aHhDZLXDki6o7ZXF0Jmm5RP
MCGgOdyTDYidIHLTRsOeihk71FKsYJKwyQblCUUmgwUcsFWqaSxPDne9MT4CMqGp
rqjpzv2D5iyqfqc++GQZ4SIrUnRtN5AM0h0Ihar32VibOZn7RMUA1C+eL4RY63ZW
LX3QEf1/RwLWXEvWzNWbsjW+XfVq87FXOB2C3tVBXxAFFZw6LI9IFHsriWbeZWD8
gMsPbv6MpnneXQmZinbg1m1JqIY0y2LNs71kAZsmPTPIg7BV2nBC4NP6msJcmdv/
TqQ2Fh84vY2981OxBLIeZHp5flHqv0ed6hzzrCo8ZBT275WoderYg7mQEI9AF+fL
GHs6M5/DLJQxzNJCdnXh1Yietk6+0hD09Ok56FLLj2sBTchqbDsiksrPLtoVNHln
WFWO0x8YZOjWNsJrwu4+11J0vI0+3zb/t33hDQQPkCnh/JTm0ptM4dcKB9hElZ9F
MHk5odVcpi95kw4fWxynFQcufgLYOB2LrbXDfL2IcQYGdY1wNEWl74nxGN2nh49S
YZvD6eoiWGd22Hx4UNcaZzV7EG8DavP6Ycc6RQ4qmvLde/X4VNIgzWLFbTvFcsnM
2XdpgDVAkIRutJjfM79uwkaLeUciW+/+0EAkRjlOMez36Hx9JIX+/oMpNMJ2V6CW
0bXfhbQYc8WZtAgHJwAOUj6cwzL0JMGZaKWvKaNoLvIzr7z1A2y0rspIkbF1R/6l
/cOkR0HWBabscCHSg9Bh21l64wFwVGUPoBgM7PDcamfNzjQSDmeyCVU5rN4iPM9k
/fRqymYQ+3POy/lV6eHM2TlgmnTgbUeNzV2gbMruL3URJkpNtNzY81yYYt8tV/xj
rDEr9SIIdVXgl4nv6Trv+wrOS3UA8N71oa+OOMqoh/7wMTfJJ7XBZMOKrgdBJiLN
BnfsazDGX1zHg5zWfpcq/+6BYokKaPY+NwFH+Bc5woIToSYgyRFcqoy49SldE2JX
Wa25ZWhNKy5sQksBgmyolgIuntPGYcPjNBegeEpsiSQwtnEyrzO2reWNBbN0v9cG
ZFX5c10nqgIwu0iX9qMGG414mfRBgrmqzd4AMzcLuCYSiknhWFBsrZgphHCOuNfb
5CvHxBIPzhQxbHC4iqSH/B6Xou1DJiLns7jAIyBSTbiKIBNVDTUDXpiyRLSJBv6z
1IehUemo2d2EwZIVszNN8Htyo9eOAZAX8jd+vkYOANbO4EoxrhDjYnw4yYCa8eLO
eb8gez6y/1YHhk7RgahClzhSjOV2dKGYFPv3ZUkfqMlBy75bqkywb6P3w5BOEZAm
gQANAou8qHswWAPFB7ubdobrO8k3xRWDbju3I6Skc7wXWGi3BdK/NNnZIjfGSn6b
rJC3XyXQvqWFqz035Mg6r0VphoyrNIueOGgInk/dHwuEi/tuFLbx2eqXkekZYgZn
0g5B14/TmZVB2amvxMEoGiK9fAMc5qk6zPFrpvzgllmhM0MJqcaZuXM+XuaePf6X
nMaEq+wD/lgs0tK2dX1fqvCQ9CC5+F6msbUkAUtbjiVgGNMzizitOw/Y7mn8m2us
3brvpGOYxG+JG0QCgi/Q2dyGmnH1TuOMqEYcjWUyjyww7IaVmnQy8b9RHwfOfnU/
aPB9nkBeETRDujOkGoUjRGleF2gXoPwwigZD5MbpZds6vbSYwrQ6XVbZuR9GOG/k
LrtLPE+biIh9euS5FDLsl20g4eCJJzN6xK9wDG8kSXzQm31vOR9ATbrB8VskmxFE
DX33QoFu4qiOOmI8oofvstjChOiEWIbHdgjXEfq9U/y9WICYM/n/OWn5bX6JGGr1
7KtMggNUx8IWoUssdf39YKBvUft92WfLu5QK0V6NmlDI79+Xr6jQtSXWQo4nqtoe
oS9Hb/lS8f+vZqBx1MPG+ddzxENcqwDjqbzKntyx7ytWJkjZtck7c7TGqrHuEZiT
psJHO4GqycLR+4hiYCUHlVcphc/WIGdMFYQ9rs7dMR9HEcURbM31Iv0iXziOp5Ep
0K+DDedjKuIWAa5ZqSiMZNatFRk19fMoN2hHmRb8/VMB7OtRbWbxgpbgeIi8eE6D
0mkr5AXY869G5qotToxNxGF1z+cK8mRmLlTzeOMotkrkyH8RIFZdWLp2N6kUDxnU
StpPwmvKNXTZilWm/QYv2i/Zc5oerOhPuZCBB2H4YvNye4D/KtT6XlpkE5ALW92U
hkyJqJeErQ1BmbXrM0BIYTs5etQmqIEDakyYGcqoBFv4nBH7ldCnl8CN88KMrMDF
upCcVIDMgIFdHkolexxwTNQfBeb+w5dX+cZmlVKBny631YomchR97E/NpyZjYGlP
/uXuYdEoKN8w3J9L0ty7k8q4p1NebWXN/+JTCZ0qx4tirphvfJbZpbU+ClzB0OOz
/VqAgdAnnHMSV+wh5sUmpjE6ur69TlM2+MTQ+dRn1bdVZwUyZOvph/CkNRnHhY0J
affAuUsCzbUEquJcNIqvGR6gIvGLuL5PsEOX8Oj9v3QLjv1ZQO/TE8dpRUoyyGQn
llAhtkFE1JR2S6PqoKaMZGLqaUPAapC4TVu2QpLnE9s6Q4edSK3IUlGtn9GffoaW
WJePLoHF2GZPvkY9+PdIUSaiw8EGybL/WqLDN6yuNdjjVBWDHnrK8afa8Lgf59Zx
5V81PVdP+bz7DnP9QyKt6i+kWmwTOs0MuonXW1iqtWBYWP3n3zHpBorkE/WTIOnx
7Oun0q6+kfxEUB5S7BrFgT3Uq5RYA/vLKiiF5rzI2JT5mDZuTQTPwWhAUZkZhi03
b8DWTR0ke6nvxbbAdsg1o7f7j+ILeapb78LqGLUl6eK0eON/sI9KuTj7qeR6eoz3
+u14itcybY3ApCnDPkgTzgBJGd+ek5Iry2BQyYDnMl3PWltpwRnaR3mc9AczyQeF
V/JLFS5Zs7bsz8nDFUZztTQ2HiL5Oal+gawZBtX0NU+FWUKa7B3WsTLxXqsTcQlD
D2yXMCqQkSq2k8cnYw4qEJj8f4y2eWWtYMixWIyTmf3AR2Kc4w9K5ABdeilNMSj0
HQF3oEDseKJddRJD67T7dIhEr+Rw2RUf/2gdWGVjmuvV3xCdRD/eJYqGnezn6C3k
ltZhIOQwv8pdEcb5uMNzk7s9OXdOiS76hYoUHIZdC8cWLY9gRMRnJ4fvWDjDvnjt
WL9iwjQI7KibIgHyUV5yDoVKNwyHvsu9u4zc8AxSCB/6EsH4WKs3eymHbNK/p5Tf
qII0ouXse4D14XD6DZFbq4lYKjljYLP9d0nR38qgNwAP/GsMAVhhDb1m/2/csME8
fx4a+QH/VoCrQ0jB4rMXPJirb2Su7tyLim2er3otLAIXfbkBXglCiNzLIX6deODY
I35YAC5uKSU951aDenrH4XnvlMugXKVeGpD1RHcm9Nz7X8x6hN14mX9GY/XBj2VC
VEvSFKUOySUuJlmrDOUxMqnl30X/D46M+PemP7YZIv+18BxhDObrYyAB4LIJHAyr
oKBH6s0pfLUR6fsKl4iok9ZvrgaRzu5Z4VMUvXCDQosg9Px6Pi0NESNa/zyY5cE2
U1ZQRtNLPe7AKScgDn2HSOyP67sRRHM8YZnxj3F9gYiL1PUGz00fc4JjvuwouUfB
efRJqkM+xYYFtPcdjAXWsunxL4ao+KyTDY3llTw5JWO1zVsFgo3yo0oSCqbVjCfA
PpJcmNBhwbzc2HA6VLxkj71XHpoikvW+qBsIWAXr07/DytbbiZ0Igx4HaA+nrHvO
hJc960rXPYc6pC2hng17KTgnPjjnepIghxCPhET+pePcHSldZ7CyfGgqfH8sHYTs
2iV7Qv2/bJfdiz4sW2JFaQg32oPoXpNoRLkPe8n3M4DJdrgMbH5JQ8PFY7WKhKHJ
41ut5TdaqJao25ls6xv3AIYfIoeUqbZVRblsJe8LpbWjirJDK4ZXqRh0eDJGsvOB
DT93uz5p9AM1jpdbEHU7K3Tfi/k6+HJrZ9cJcqS6T34HV8pgTiAd2i9SZdzhZEu8
1rrEOxNLQsJbrYA7+v+gxxXNIWuyluwRUW0k9u+RCRREjo2vB46+7jQdyMGjJtJS
w2ToDXWgC8IDqk0wyGIBsd2y9ycylgolxLB0yZhNv7c/7AXsdnX2KH785wHfLi5y
Pn341m+nyZPzvKQs59rObIriS2+h19DEbKqGjT2uVO/431uIZmuoTi+LhYba7UpR
bRj6dQUgI8JzzqxxOpbNUnSXZ5ZIvpYry2+1KrbRPxsFQk+tO7vNvSacysfuDk0l
2RrZphDDuhZIgZ4V7H4ZVSENDJ+DqqVhzZgox6xkym6PMVVxsEmzNY72fDP4vJgd
WjS/hKy4ZbRuz1kpWsBZLZvnpyfFtv91RK27xyiaBBLF0lbKszrj9Ul4aRj5RJtp
xSNJjkeHABtHKH0mafdZHOsqaaU50ZYiKMKaDyVzYXCacjydKsWGu0dFNSIP6hOU
nx+CTyVzrU9i6M73L302iIv4etzFdJLxRCSdL6Wg3dOpRqFxArE7c8LrFrSfKGGP
MqZeeFbwkTy9eWScJxHiRo+efJFPxYXw8QpypROp/6lyosAmRAz+6Qjr5JSKZ0YM
kJKIud3EBOBCmHJJ49pmIqXB8zJaNfA1qQeUnXe8PDFwsTyY9c2T0EJolZmfxzXy
VCM8pO1Bf0aSPqJFoZcUm0yHLtpveIh4vipZhY0Y08xtdrf6vtDaaUaCxJIjY8G0
/mgBliIkeW+mafqm6zZQ4mvPp68t+PCgLOQFykit4k6ijqN9p40yi3oK+cmxZosk
Vp//RPvtCFyYjlYE8y3yEsTZL/Ta0hs1536q91Rulq2LK5WuSfehWYR7K5blsV0e
09cAYkQT+fpdIkI/4x3wQj8R+BUCrYFCTU6LYesJjuXwY59QoKyX686922PyQQRT
UERp5+w0lYXArNJ1tUPqGrnRf+U/rIN9bmKGPBbO/fJC7amiDWQT/Jhoqvs6s/ul
GFZnKBTtHM5yc8YCJ4k7//czkRGRnlR/CFfnFgi14gonAq5xbkFKInSOEAmRc1Qv
5N88S9cWq2CAjWpZefpg4M6QQLI69Zgm9W+MAfHD+bXRNCScg384YsY058nD7Gmf
qrR7T1ERgEM6YJOyHf/R4ENAUct3i9hJYF9gwFO9qfcHPFxDr4Y64bzc4mZ3YIn/
Hg/KCUoWENW/XV0N3iWkMSXBE67uFjJQikChxYdehQpi/yfinPNVzEFGuN0bBUxA
69SmsQr5y9z/wxUeBCFxEVVanh9Q8GM/K9MDAMiXdTJqI1/bp3WvBQmyfDHuc6wH
tGF5WCJAbQQN13pwizwhAYBYQVwAznaq5T2ioHGMhmpEo3hb30mxhzNl6uFlNEnR
dsAktj74P6C1PgzN1mysi5a4xiONFQagFkSRYTlwhK/Wt0kxXR9GOyr/NlTAo8jX
mcCzjiPssEDaW5ibmI25ZTqavrsp8bgWIC1rTEqeNzWKZqelLKzrnmA7ZkEOSirR
F87EQNlSkI/YEwnTwq5ODvvVQATAGt3ijV/hLWTCouKsOdjRgA2IUobey2wRngU8
LmnZ61TFuZVPi0Wx18vpyxPVL2pqHMVM4FnQwaXBi/MSnCXiHREuT5BhjWlemBxj
+eDorT/vlqNxcRli2nm5xk0Wlp23+nof9ueTpVV0AaFG+xcMgk4T9Q6U8333aZzi
pTrZUnsZM5ADw/KRq6udLxYtVDxmWnrxLkFAXc9GNzps6MRr9jN+xByfeea7h3qf
wCTJqoZQZwJZETXiwGGlrHDUL+9yDv2LmD/9qp+a+ASgOgvLDRX6Sg+Qz9YNFhmM
T+iw5gsJBYtpULJuqZrGE7GNNUMBEpH9wO/X5k0oE3XNfMLx9z8RKyfglydG4kg5
gI2+7LxYkTy+ct7ETYOe/kI4NrWQx9U1IFfhW0UklmpFsXAA/LmGwv+WMukwpQU1
bMzFCpQZmLcRKSBS1zDG5W6YZioY6Nt+YBwPntl3xToQIjLpAZWxpwT4f0/V6gt6
CIJy9+KLiHjrK4XUNR3RFUY9miSykjlcjUJbHVz+O+ea3URfuOtA0rbREWRgBHpr
HfZElzGROsngDdBdGtHSwOFiWinVXwHavmhn5Il/th8zL/SBUWQ8OmEL7a1ywDF0
WusFzEHEiy5Jw0SOB9zg2m/SesPU1jfmnYb3kR4k3c5JRa2dApflngxgM94ji+O1
gJxKDACKugvM6TrIf9gqI2btekmY+TVX/zz5zvOWS/JjKnENlzSCAmT9XSVXCbpD
oMCG+LcL3nQy4TZxYSLK68nN3wdBBVJvdscE1YFcC0UAu2hcVt79wCr2orsuI9SH
CoKhh0WQLjQdmtV9ImoZQy7ZAY+xhXDy3EEUKphVAPG0cR5dSBLAhaire6nqnV2m
7agCVfk+wPN2OM8ACmwxCNK3lUhLNfOCzJyDNHfjGHP946BNleaYG+43KHdsisCf
UKDbLBLamDW06CRTAZq5RlTCkoJL+hJqrpYIqxUXn9L4L181y9gJ+FQg0Td/vgY8
Bw+aQyM0ISIWwFR7eRe6/DKSmood6x+bktl15UhJazU8uJdnPKkvlDAuEvku7SFN
UrSevNDfA1z80cQpWU1gHJc2ri0ruozvW7z7OTZ66ToeNhljtpytmQvXoFoWAP0+
78EBLEU7ldcjFBnGHkiqr1qK+87cbBagYDu1QVBFyDKRAxbNN9DPOJj1YfevVEIF
22G3MA4r4seA23JdPZ4b/QHF46EJG7eRnN2zZgOA5WNtR/lXfwAlOE0wStyVpROr
Epix764enewwHaJ2SgD2lSYr3+pkDuncrCQswPYpdwOAIl8YMhcf7Q4FTPjEvgAW
i6vyCjr369h1zRLDT45F2QWWs1P8crPbk9Dj8LfYRazIWzTBCvNqR4XKsWXOG9pi
gyQHfDRPLCJq5wAMeOmyEFSd0CwmsY5klWBLJC68AeenIKpfzOfS4PwxZv8RUSyP
Q3az5SStpOgiz4zrXxvEkab79qXi8Lu5DuRiHh5fQ/DHIzbaaRgUrYhIh8DlYzvX
gFL5xOib6mo21bK5MtP5T5goGqcx27afVn/wIKJ/tXCQxI9bIbY8w+SuyzaqiBLJ
FeuNfMFqUsZ6ZTwGF3rBKQGjTSvRoMvWu+KjY6i56nv2JcP6ls+iUmD45u/BeuxE
tVyMjvfaQspfkvC6KzQ+jCCsojAQgiL2DihUHqRuR9WMRT8Sf85+McQu2x2XybCt
76Z8VxJ/A2JetJ8Q7VUl+MPVnF14m3W+xsVQG0ea16Jcnz2gBRKnHGnT/IPhdMvl
eb/S4V+ClC/rdBlMM5ONPZQFG60rrco2hGQnUwM1Owx7w1uIvB9bRTZ2CbHDx3RW
d5m8fpH8v0SCEH7jHNJMoDHS5LoXJAaO6zHTbOl2JobURcO1n6sxPhnNF4l1SN/N
7kiazOdQEOSYgKljyJNJibrO08ZGvObpAQ/EoiajV9vPBmAn0wENntU/+hAWSaap
vEzf6OX02A4Af2OpZetVrUoRBVIAyqz5CLLKdtr1tYbxrDUVx/0h2odrDP7cDOfJ
gAZj/yh6io4Jij43mQPv5edGYjoYJwrr3PZYf9UqMlEngGeYnfwtd/xYRM7S+LM/
XwN5u5E/DZ9x2NSJ4UEOUVd7abeYH+jXPeL8t6IAJhngYz8Ognc9NTx7zDbMbLyU
QJlD6ScUc5u1B4k0eaVnmiiDntPr2DSmX4c9/Wd8iXjRxqByjBrRciPqxBfCKePe
khqCXuqiF3FPe7Louij8iRlRW0nBkMDxreYZ3oeFwwduTX0JHHwyC9cHGtLbI6BI
qLU8ZXp6wgQU837YNwD97n5EJTrQZkSJqkYR43KQqLAJFBJGjd2tjrlr2by4o/PV
2GDdWxqEb4mLjCznfrPOlCDgQVeqXBagYq2zbd5J45S8ztMkj8iVa7uJt9Skf4j9
lW9s8vPiNjwMKMCLckGHp3/xaV0ku63UYJICSdPJl4t5y0VNBAqzL7zbzD5nSfUk
3GvQ7YiqdGFi2N88kmK1/mHdoS0+SrfzCWmPDDdGd5smZUuMIvl4xv+TTwCkmf+W
63q7ETUOFQdT22nwzfDj/X7So9J3uLN4JRGh+xJo2uZmlapH/xeav4Ct8hRsnQiU
GG/PUSLCFkFn4or1VY+BAoP/IpK1mMMHoutA93TuHHV65M/XD12mkJmm9n4GobnP
tQFyvkxiNLS3UwDcS1u2sSp+S8AIyWDnB1hV5uKxlepyh3hNhifmVnHVJfZPTZdT
kFBeyJD3I3UbX3w5CeTmNbcb/QWsUeue7BotCbbDwgOzmRglZ3LmQ30fyAaDfnys
QKEYHs+o6TQqtkAqiyDtUrdnoLUFPLNDwgeEv+upaq/ycLuKbvDSPphXNmfTLjhS
N8t/PVgnIbhvP2CMUh2+3PvNVt0CXCNcp8NJF0+tVaOzMGgkvle6GTy9aAbhVBiZ
/AME8V6zhAQVMdi5cKAM8xpIBphjJ76/N5tquTv3ti4ZTTc4d7uSHylLYjgbU64c
3yeVaxkvBQKBSZGyiLnNP7KVbKkGVtR7tGZ8ZlX/MuOP4RGA+7i6Og7fnTXwNsO/
eJURwuMqBZhOgGGZ8yiAOjV8zDViJmGkDeNnztBqjL1Z0p8CGfD7GNXBtyxYPKI9
ldHmo2DNQcv16lbWBKeZIltuPlQYSd1R5Pvhjqd2GtX6vZUSAbSCbtK4XuHdSKXz
V0NnMG899Yy5G7zpIPioh+o1LDqRaGCjG+lnyYhdPaB2m6qDyyBEOFEW3TXd20vO
+aNoCPt3lbMLnOR8xpKIQyZVyR4clEyfwS45UaAkW1DCIBF4uDrmGYgNPpNI3QkP
l9jHZoos4OYQL4NaOecaRfRjTttU+wTTq1CcSTL8V6x7RJPyznRkpzaYAStr/ahs
H34iFbT7THOa1RiJiLekGtuA+CL48ARDzztrQ7bK+GUAn77ubJTs+e/Y0flO5tcY
baUYY8NyrfThleOSvw30E9SRgwEr8TJ0LvVqk4DdS57Jm7fyKSEMve0uyhVJqDdi
ogKpu8YviINY/TUEfaJEhJsv2h2zyOvtwqGo3WSs3i46PERDw9yOclwK1bdkdNik
De9BBd3mnPdTm5b24Bf0s/ksCClc2qo05vEl/BCRZMHlR5XZlU1yTU3BhisaH3n5
HIBawGT6rtM4mfV1CYlYT8KPURIypegSfYjw7k38BicHfk6JXKtyLAiPpKLVhMl2
tr/8lcBOaJQ6kseTYquksY3LwBuAEYE4RrLV3nxqBuePMIVV/zP/v6vvaKHcPmPK
1wQuAxB5nVX4i5aoAX6f0z6UCIGGW0MRhzwnheFvfUyN+F+ckObWLSPAaSewL5Wj
rYCAcyLhTsFI7R0Db1hzJxgH58IRUDkUbh7gj2EI2NAZy18jr5l0UM0I33aByZ15
QGPeNP9gzppRTNen9ALGxNVUz9+kOC37ILfcJQL8eEieLHEYdIbBJ7RDoGa5q8vq
pk/wO1/UdPybhEUqpfEpgOyjb7GmP2VPmmJvdxPxEY+QME2RPswC9PtopiD09jRH
FgtRRO5D77obFO7haLH//Uuow0f1gX8ybXWxjDDNaWQV32l4z4k8OqzyxbXoZDQB
KEvm3Umsk2oTK1vDPQNYz2s1MhInKcsqwFwJ6VdyamXbdB7MLyEdfEdx4N+X2QoN
bfjek+UU+gRKJoVtPNS55kiHM8RCDD0FnVX6MwhcctadZpFWz1LH8EU9juBpTYiC
rbpziCI/XZpnME8W/0FwrytWXrOYlqSi7Ntg8XWQYz71PD8upNFRRBV5LKDDJyOw
Ovs6UXdU/mhHSCnqEe1acWaw4pN9WTDIzbhWt4dhRx7kBzy3lYpv06fcy6a5Rc+6
fPZSKWSc2DL/h2kGJ6NhrDBTlB9fAlHNh8qQS4g18mvv+O5yoeeGVXy3vNwTF6SY
vBSk8Jj5GdpSrTyOmAhrj7A0o8M15UDCRkYzCxnZ3+oIoFON2RK+ctdi0Q/gDWNg
Vg+toj3U40yXwOq1xuirhWe7Ea5dlMpjxPdo4wcxtKr5kVvAjQ4My1bqTU7Ic2S5
TjTXuVAinTud9osP5onASKOOukrrpBVdCRDJVRdIhT1BmsgDGXcbSz1uWgQG/WmZ
tFNcV2lU/7tI0WwMrtxwj8QkDBv0e5rJqn8+SeqjHCtwROpwMGW7GFn4RALp3dOS
ywo1XTdAMB59nBt6bzIZJvdWLfsnEPkrp0UEpcSve7+P6uhbQ9sTxAZmq7u1R4PB
O5ionQKqpU37/XJtRzEVElZ/XsT0jNOnSzgOmNKGv8vxFo2jZ3MWwDJCYaWGMssQ
TwEiiCW8AuGg78/SGH/6g+81RpNpCYm86qfWW29NiZ19bKlVsEJUtlcD/8vcXCoI
s8XdZ2VEJ5VFvQ0rn4gKFQmr0nzeUJd2dTUN9Ed/TL3ZakrhWBxMYteSFNvkCiTY
UhKg6WrCocwOBRiE69Gm8i+LQpirX+HF0AVYWGYTOpB8zHL5VcCfTWu40sPt6hf2
gecHdg4nra2Qp6Vkuvt5YTtNjJ6iBU4acXqF+klT9SUA6njm8QRCWE7ysKkw7Xsq
wuuOKLclRIWJxSU2aTPY4uJwDdRqiegS01Ri15OIaNdjAMi6PxMrHZSlZuzWZkrf
V9rF/eNoJI16SS/9UufS7Tt4XVcJghkw1602ncljl3xeaJ5gkoYAGLg0UM4hJCxr
UwxrThodNq6goxpx7482M9NaTvrBcPEOOXUMk6l4643sPIikLoQEc+ImsyGUDiZK
mDPnn5ikGzyRyGGo2SFOtkeGXDz8C3qiZICa0xdGUHDq7OANpVeM+uBSu8tV79xq
kITjFlkJWBDvYNPn4d6dRmTEMwWJsvHEJiANrsMRq2fVSPQEJFpdztM6pSDBbS0F
5Uf0kTvFO/rQmwjEBlEPr9dC9plcFSEg14YyBSkfH+uA1q8SXHfhWaS4NbY5q1aB
Nf4u3TgtZUdUevw2sLyl/Bnc2EaKOrR8VS3Xml7c478TulGzT6nZOBWccIluiUZr
zjv0xzza1eAQo52CYju4FkeKou6w68wOkDZ6wZachFJRmoLi/ffb8BcabzkFrGkT
1o7+4KQW8KErA82l5FVwinR/gT3Z3cRq+6BxPYwCmrHDdJ3Bam+ZRqtq+1b0Jw18
dVrNjup9ERl7+MB6tjjPEULq485HFewvFmjpRyDYYTx2uWyYoeqYVwAe2E9CVrLn
Q/hqz7idL/+cgCLDuloU7jBdVty8duZk92lfkCtSc6VaXSuHzvl7jcR39Ygzs7Ll
3gyDvWCxwEia8UA3PNfe4Kod90zE64cnxtA30BYaSZXC5HiqeOpihjMS/rNhZgzi
4gO6R42e2AUTaxxHQUVLlwlohVo7nOscBJj+j0ZxLZvTVmgRDLcgcUFB1cYhmg2L
9441vDeO4XQ6YyJV9r3U155bQjAfuMciOoOBjQD2JwhzzkLjU1DiHWb4KJdV+xhM
rdEFMUHDqKcCTiYCs0h7ay4hvyu/faR0V7xRFPiNdjUq0ZdyzsH4kDMMdg+OInJG
nvCvaQddBamofwDfEVc8aw7Ac+4nmy2gtODwoV8DmvlUWHtF6P1mv6MUdRcl/4Du
hbSMdNV1au8dhf3IdlKLHGcGYTxcZJamyD5M3hYj31XiaEPMCQtoW5XcOaGdzzYN
PIL5b5GxWnUNFTMRxZwzte1HGJ6X+aJ4N2L+QoHGzoPcWzceJFJlP4xGmtIMDyOH
tPIyoHXqFJ3wsvN3Kwyr2w15a2v/ukgfQxoeNC4FuugMIyTpQIWF8oE92tTNN5xR
2KR8XJfeucUKHEpZPimghGtTfwUGd10NtRhlIlTRagRSXMV7vslVrHqKAQ6nElOC
Dt0S2K8ZG29sSeIHVAvJv7H746InwtqS3M3gWq0DUmwNWzFjSMR2Om6UEDAl3Yg4
ipoVqo7QB2M1RDxHfr1JhcEHCnanA8WXhVw2Jak09iVo+V0XlDl+TiYex3F1UcDj
8DjsBNwSVjV8zgYA4liDSDmiFO28fUeKrjFAwdj30USzJ3aluI2BudnAH6duS7vs
TaYPSTxpQ6ujgxZNoNuE+KyzWaHafUfVj8WF0XnNdLV05wurTYJVQPnd2Ci+i3gE
DGYhDJ7I2sEWURvv+WpVs1VzsiqG/R5Koc4zytfMzhm+6qlVB0tadFsLyTM32msr
5NLOKA23Bhh7uybda+v8X85bL9nm2+VXYGus9b7QjIAdnnRBo63XUY3nmV+Os03+
z7TnWvl9fCkvU6KlPuP6O9sBJwtEN4NdeKL4OxGSWs8VhIgzo9mbnPt5jwZdMfWQ
2z9DbitetcX6MKLWzXG1RocBIxKTJUzt0Lx0LmGoF2px6j/YjgKqCBSR7SaQaVBS
+uIPQv1TuIMYiQLjQtpkoXkSr7Af8dOeE/seMpDlD7htxNJhSyBa8518en0nhUV7
AWCCC3le5rZRREahoqWNVhD3tW4iJtx7/oW3AE/ArqZaj44bwEmI97tK8LxMJtW0
aHMXpacszMx3/NmuIotAeW6ptcjQlaset3RAFfcYuv0FTsHzhtNS2ISIyYducjSQ
rUeZwV9NHlElZFQflJO9vMbpU23sIDhluphSnlqPo7u3vfc+BTf4Wj+9jU6WftGn
voZ1qNMuq/8hcxZUHv9PAyOPeUd5jpG8CqJTpuxodiCz46d/YZlzXo9m1di+UtQm
HSmFQqv73ozPCOnswe+MsvUs9syNiu3k/Pa/s+Z86/BTRona6TtHRS83ge7v140j
ZC+6nNrt+MupfCGTRhfUayzICfk8/C0/b+XvdTkCT9sos5LyKAV9Pyw0BWytOfTz
VTSLQdVPcpThMpnspR8t91jux/myis2gB/8A8vgC1Kf176DtdqknC4MoIKcClkwd
YTIkurwZKVjwR3t784YjpflHGkrBCUPOoXaoiVKMSF2mSzH8vqmbD5tvCS2ST6eD
6FsBK+dpFd9k9guhD9mCgOEuq71oCbasWShvEd+c0WnkR7Nw9OPa/FiriZrernl+
TJXLKh2upbIS4/ElrltEjWtd/prP9OQThmSuh8iksZKSBSHW7RNn31Ao5nwwAP9V
Iql7rzZKRldG9CqSlf2syPzf7KojVi6DMNpELt4HEIiDFl9wBncGYD84XbjlqYx2
Mc/xgZzUr9KWjpaBi/LCmIIX8YIxzvhCIWg6lRE+OwCexWzkYwvKrmJZ6m3yPmB/
T/az+vM1sK+YQnMrJ0Ge24Qjd/XZO03dMsab0YsErURm+fR2XCZAfoWB7zqTey7J
1PPzKyM/YeJrMQNrFS6Ie8xSl+KjBEOfRxQCs+v4uJG+22RNqQMf/4N0zcdQSacc
u/l6ZLkGP9PFeKW52Y6ldaRXi+RABaGFrMc2pJOepJd6dYJeVDOGwvxxZSwMjUwk
f3RgET6TJHUdHJMJhs4SFERK4hnzD6a7KavDj4iX9GjOz/kvgxOEDArqrKLqwzlz
HLaVTPJXvQWdS5fonVUhV6aGaI/Yrwxs1lHpeN/8auRy2Hnsge77TRmKXQmxAZN1
2TQym2FMQBXwIe/e4cZgrClrDMWxwGWm0qGEVGZwV96mMFcEcdLkM8YFrVERL5Qx
KcL1E0IOntUCjTf1M4ZmO/5PvPHVZXhNMpeXFrwWxiGYQcaJLWiShomoBJ41xasR
EhHrl1RjGBpR+/Y0I/8hrkrLj3nZ0yeGy5e6KFS0yh1SuT2zxyrMdVFNCHYEomsW
lXAlqZpKiPk2I45rtOc/Uj69Ygw/R1m0YSuLPNZ9oTVW23n732q1Hu5/sFo4rfJZ
XuYBZZrjEo0j3IWeud/zIMnBc1WYlzIf3JnxjgvmDFvlmYpBSoYdNsj1KLZhIrPA
oMCUzabJIPEPqaLwldTIFUn6GrlJWMwOf+7kNCq/4tZ8q/5iX0Z0Nefv8uczcBgY
UVvTQjoi7gje75ghmPXzQQ5yUB25tFkrVl1hZV6MoMavYce4QM2rKOzVC+MZKWN2
Ly/hZoE/IgMCHSI1OKwg4jZAw2Lr6NPGv0qvyftn4efmW4jNAAUNGnUW8n7JSehg
GymZjtREERprp8Q1OkIzAKvTod89SbKDWYZZ3OcDHjfPyxQR5HkQZbZQvVfpl632
aFL36M6R+Gt+KXbJYwOOWmrC3viR2Bbp6TPxSPJMy98gipXVQGMtXJqFHnGYVBAC
PCkp8TipiP6zCvH63Q4C7ABrjEp0jjpcSfkwD36rO+wa9+1LQutzWcOavuD+/Q/T
0tPiExkUm/crT8md/wnejqlykhWa6673g+GNHKtxzjuyCxkaq/Fzq756WtK5AlqH
jvjYYJbmbI7Xd2UrYY+IvuPIwdR4ARRmxu3u4KUuuPEfXikkNaPuvuNR52T3J3Pn
ts5MbUE1jSfvs+W4D99M6tMi2lnBNyGJIfCVO2YKqqu4EENQC9yuBiQiC86bPBMP
z07axo8/8SS6xhcrBun6AZglV6OpJWC7wIlxHHNOMqkKFR2nBN0UIRwyvqs95GUr
fuFfB2IMhQqCorNn5YivoZw2bALCOuZMxTgFhVj0pRRFv9snIpWr9hg2dCgJnVnt
HHMkQzl+l6D6XPXQUdfs02itqHEk3Qi535uSSzyjvHzf+iCqVioXiOFmnb79xtd8
10fQ712+0NLpQcAB3MPNAy03FQ8Tr3F+ef5ztBkuJWADHeDBe6GeE7MgNZyIp4IO
wE+6R0TLoqv08QtxI5tIdhKTL0ACNMLh5bV+RohxkE/xkMf2/pmIDHIh7y37kEX3
wmJtTToHYGI4EqrLoVYzxrdbpNcSN6XV8BsyT32g0LRBGhDisw/CrkhbgvckeYwm
fbuxGZhmqBKU3OnJQWeV6JAWgvJmUpCnxELflpg4fbUwToAZOs5YxZrPY/xUlwJg
YsHaH3TYpeXr2p3PMUE1W6nl7XbBlc7+oeL0+pAh78fF8+1SBMUxp/6ky6tATPlj
bHWnig56NKa8YbzkZAx/eOx5xAmdR23ckuQBXzQWOqCqKPCP0NEOiQKUKwEBSABS
OzUIGs7+5gJ0UdOfqUn2BwaeHLj97hRg2zBmx+yESL5XZD5uOhccB84JkHccPGH8
XzjchV+u04krBplgyxv8XLfdVCXEPcfJJ0fe1JbyeBLHAS+QPFxbvozX4qKa77rn
q8N7tWgVW2KRb6y3HOMsY76y9/YoDWyosry9mxYh2JLeNxEscbNM8KtgHgV+386D
2nVMpnCafTcXnsaf/Jc6mFY2z76rEXJbWOJaqawdv5Z3+Q+G5ZcU0WUVdkhofQb2
PwHo+6WnpXWdbH2Prt5lPq18LwtHovSAmIgcpZs8BvD6xh9wVLJSz0YRyn/Q3gXA
uuGtG+uwIOSaea61zNn3VDthiXIHYws4f94Ne6W2biWwAyIbJJoMh0wO9GO2R4U8
SKOFciat+JhV44amj0l1IKKyQZB27KIWqJYJE3VNvYpmaR66VDZjfrGjv934lkXF
hD7TOulQlDIN+0DIsSlPGYA6mZw0uagDgOV+OSBlG5FWnLlZOhO1QMYGimKNgdbb
IfgCGmBFcRCaIl1an42XHTMcf/MQGkGdUIEVa8AVc1gbd93AzLBaAl/oFB05JHXP
20e6YRGq0SVnxyDeuBYQRYNSb7EOmt/PDREJ9XJU/jwlneb8lMRWDULl1EBObl5m
YD9iZnSi64beRaRK3Tq/GvAM7IRrIGIJeWJ4mh3YCf2VLYBdf4I0ismlHzp6EX4i
6Gik6iNik+wrD3UdG2JNo0gRS0os3ueZEjDg2Sjo7hsRJwqUCksWjQd2dxB1ni0D
VkkCs6YuFfoebC6FK7CiI8ljfIqXaCP8tCub2ki60OWOft976zsGON9wHdud1ZRS
kllipYujyZkypdKYIVK8t7CL1VrLkDfcYYhkU7OX30tvLo8FyaoQrkrmxW1SNAYt
0C3zFEyG8mEHu/KXD8yOAa453Fqtr13Q4p74PSU29aVtZrUshyhWFzV7xjw+bYw/
Zo6EpPdFCCLifBEK/mibfRj+NdNC8gFlZB74Ih1qds//aVWj1sb0FokXwFUytI+6
teNhZx2bW4DHvGvU/LztxJetvhLRXG3y4FpJHZTzY9tP8yAPxinJAOyRuzh81gwz
YPXjRfbtE13DOOhZC8Rra7c1Ziv02IlORlJJyxWk/CkPrHXrbryyjNuWfaTDHtMC
qKunip9P+iZQzIktaa6KGiqKY48d6MMnoFdGByUMJWmYvyk7m/GHzjR11EMQ3Ay5
bYz1DJmrkMit6UvGsyxaz7HkW9tL94cfADAaj2DutGOxeFiF+ivGi7DT45HYcLLY
NWlFpVHuTI9YAEqc4leZbK4qcZOKuLoSqUoc3qLJ5MKdgC6ploUxP6CqjUXn6y64
hV+7wu7T7/nuwKaF1QQ3saXAwG7qVcgdlSftiyVI82cWcolgzeF+qp+53ZBxTpiU
hyI9o/p+WX7QnuaJG1jMXag0nKsDUW9fci4jL/6gPgchpXmEtjUTvvIhsnbJEaJS
uUU7UsieGjKLC00DffV+4OP1yb1dm6Vzq72rikemRbk8Br18HHOc9KChneuo5meq
YAczZy92ga6i6GN6vsqalcx9MD9jqf5+09m/jOTLp7bVgMbqzsoMPiE5usxrX5XD
El0CXK5TcWtKusG3pLak3FBVc8NxgCVqr+wa2K60UrhvtyXKm4n+KZLMrdk/QFr+
SiR56WByla5j9SSMwx806CPxYE0Uj7vynj0oZjtIhPN5fs99BXgddr3LjPYgDB3O
V//ZzeB0mvCwuljbhJKfO+6+dNZ++eLhI+SLJ9TUezEAgiY3pfkvn3VWfrZfEADe
cRKXhy5aZXBCeNJRAofNbTJmT4vXHZnt/vqIz0FDnernipF/dnjHwPirTjhu0o7w
PuKg3IXMP5ZD0z1rs7GNob2Zw5VooWUUGRnYWyMKkptGqlhh92QiQHV/K3XLbQQW
8HueTGOQFKVcClnkub+FwkG5ZJgPVqkgyYaIo6v/rY0/hlDUr4zarnxkSDaigf1T
jYSucQYtJ5cTy8yOPVdiDo/Zv9pruS6VljnGVQnHvj6G/iFMwG87v73euPr/tZSk
9lrLsMy3ge+EyhILGrHUs46UN2EDTRgjE1ZCTPzDyLxA8q/Rfmp2PleY2jbXO8RT
4AzNPm+pSVRwVCx2ef1M7OqfKBQqzXD1BXIgt3KJiSO4wRrlsTJqcSVMs6t2avv5
lXtWU2GJWBgK45g1KiONHFcpQDynCGxiGJbYWTck/nOiiSGKVaO/4FLwyqGaTCnR
DbmBZTiI0JA3YTlIVsfnQ/DfNSrv+0Ss4xDJI6dXMPnVg5Sr+NHLBQvOoPtyOEfV
rW+6GzGM0jEeDgt1jSqWWFloKajqqRKuJeJxmBDQMvuDdb53NOajQHVlNgkxGgh4
U6/w2zRXB6FMhfiDte50Nbeyl1A3gcpHfmgpw51u4KaECdLbVc+aKmHNWXnFmwSl
oeFHzphm/GyZUxm9i8efsvcGsUW7nj+raJo2IMidxtzIJnl1wmSVjrnxa91MBOq7
xerWaVOTGKWXCcfs2YyUmMTeT60OwoGBYpPo6ihPx4fxOFLACsrP2enLtO4v4O7m
GXUf4QihVAmXtP0/pQMIiqXtuYwuD5qomCuU0U5kAuUC8dw6j7Ni9MT+trJgS+ra
Y8IXBDXHnXcn9FtCdHFp1oQ9MaMZGc9ZlCqDYqf6A3PRQEDRni3QQCXWJRxHiEsr
EkwKpDEN0EVtZQ8LJIrGITHokvQjQPiEiUHxvClhbFW9FLAHdfcsj9NuG23IE0nY
j4LBfhA/ZuK1+G1fqxSmPF11sxHSJ76DXR970j4/ipq2snBcUc6zZrnOHaQfPTDp
Wnyt8dzJWq+I2D+z0rGHpK510jCOC0zCYDPG+Jr9fjTGZR21tBu1Btwc3gZshzHt
zHUEwOZGEoph2sPlA+fDPJ+cozRZwfpyOVTio042sF+nbKUBvnH9NmKHJqkiW0AS
0vxycLTxqPqxQN1uoZZX16gkoo9eh+TYh6hyYJI9rS93heHDEdvvUcMittASYkrn
10rUHZGqymzfLQObLfAMa6e35Fmj5Lt6aJ/CmYMUcmTCTmzufFSYHvbV11XLgKfl
31QbTWo1hAftAVa3z1dz3iCzV3XqplQJoqMapRItjQ+tmCZqXaTVLuJna3NfNzLS
xme3xg7HWJ4b8El1lcrcvazTdf35u/5Wpxw5F8HzI38Nw0BawDIqzFEtkJ/oltni
BNQX3x+XkJF5izofXA0Y3Xg8+YRjRexyE9baNU/dox7WlcGTLkOBVPyu94uqSydj
2Rsvi5T3HY8OzoHJhlUtkia7qL46idp1BMPu9rSoN0JYLFQzk2p/QMX42LueHD9T
8+QjTPzF16CxYbXFYNPVDqgtNsXXY1KJI3CyMyFBDv+cOkoZN5SdQURiJUFAU8Aj
Y+3T/tOPwNegGfEoaJsawg390XUHuLQKJOmwD7XxRpZTb2BQdjP210Z943qJyi+L
QhSLV0H4GaKeh+DH1mT15GqwVCLU+BArmXGub3P84QCSKcm0mIOYL0+Z1AdFSsh3
pT8S4S2oNzNPiybfOYjzqhg0MGrn7tRA6X5OVzMm0sP4i9kenNLAl0zUWigNLn4u
F9Ohw7V1N+8cT8Yg8JnujTKOnIyAvcL3SWl+OI+QDoOtdrO18ZLX7XRU0C0PE41L
iDhl44laH2WmwEbSMNgZ+ELhCPL2zPpcGoSYYLI58TJoWEWSmIAullgDM6XHst1t
Bqe9pTAghIJOGQvFYeewkujv70K4jhKHi56i4KRd7vhDJsXhlC1F4yo9eiCIKpAM
r/fo7BQcdur+Dv7Jsfc36Qhy1KNoiwxbEApEm1MQ6xwU3QBHFgJhacqY+UI3jaE0
6AHtgPVYPUBfwwuAZBz8pz6BWGIqKi0m0imY9SECgSqw1jdwByuWWlWXn1qvI7wB
s5qgndj/nbqRuh0sXF6qeI7unQbIixwmseE0UJnEQBWGCBqMbDPAHVPA/2Vt4CG5
nREuQZ6lsASEe6LscN5xZHpFjBCh0YG7sznlknakOn8MNlQgyMoFr+s5aykZHQQc
tQk5lPPwNXuny1dtCcGmI6jFD3qSB0TdP9cRBRz/TXcisROzFI4Uc/UiLH3KBSyF
2JUlKDf9i5ZdHHG3S3TAAf/nPYXuAu9Pp0+ULfE+Mgedkrvjr8YeqxrQBB70TaIk
4TP8u11XRaWx8egZQonuWfL3PxxsVWpekTqCFMDv1DS/Zhc5kLSWg7krD0cb0VI2
KmlcDbk9OG0T3A33gLlm/ubFGgZ6V7gegn22NJ/hthltfG7Q4JRtTOzEhmZE9b86
zVxRUfFHT+svKeyormyRAkykBBTJZIzL1/IlWkhu429Ywh5CZVtIPDoH+jjVhqSP
h3YBAbzlM8k4llP0EX5lyEat9yu8ObTw6R5wbOeYKOphLNYCuTWNx7la+u3V2uH3
6AP5oAQt63gnbsCyV3NaYtSUV8ud+Rabjbj+iv0NFncAz1xE4MGuNKQw0oTbqzEI
RF+TXptY27suAH8uYgLPp4Fp+FAcK+ceTo2JS8pepJ4OBvE1txpy37rpgYFJXKU5
t7SIANyWoxRrlyU4JVG2vM1l8V7s1AqQ8jnmt0kjasdatMXR6B0alNF1t9wM79WC
UtWeMNKCXUkDXl0vFHQSeBkHKgv0M2DT3ZorM3WG+6ZLK6c2prNX6Jb7bOOLKz5c
vf5pf6XBp92j1RWJhYIkm7fhcdnfU8waAaRuNi7rKdC8nJa8bDs+yt+TifvZZe/1
oA2VPRq3+qfkZbzMvZEfnBx+OC9rFHa54ErUp/+lsW0X4bVkToE4uksfyqh05uqJ
Z2OA2FFqiUlHz5ZL7Yhe+kqmHcd3qIyQhZ0R0XYs5dhy0NiMeuu28wY6BnsqHR/I
POwR4sMiPQ4Ynr5Mx47qmqsqwnBGAgpexBcLewsNpcFsyyPIBWdv7SXDz1NiBPrV
KtVtPpjoPqsbuUU8zl93MVuVTpQummX93aWbzr5t3XgUNM3XTAMMwKalawS8KXpX
xEo/RRTTZ6/pHOW7hV1L+jeuGnErypc7SoWfkWqCXTAbB9vkhL8i4EtLTvvbFSiz
p1smzNRd7K/TophN/NPONPCg8eVMKscBFQe78jjdlah6YNZ8dECZFH8R7pWJTfmF
6Leokyb9LkVuSkxhMJpX2aKQa3DIJhIOnWyF7XXC3XKXNXK1N3EOoDmFAC1eC55D
whji4NqOTDZUYdp0XaxmjkvmdanIoHxYvT8aGFZRd43ywBlw2HgFyg3j2cu66kl6
VHIKyYGu+1+VLF4RCehqrE8566Yzng3UazjKPJNj7ssc1tj7sW+O7lZi27JHwWQM
gfVgYM3ntnu5qUUar6c7weK8jY1kNWIsHZUaNvHvldU8f/PckZe+JNQkjAGOAetU
2ppXer42BkzX7HAufjXUF3jNsMzdXfM0PB0zJCPHI2uDBaa7ORYBWNAF8sgiQdY2
Qr3+fAqbGlKIBGFICTepxPYFCoYsItYthecvqcq2B4syyU4f9YGHx3XPfkBgMMjQ
Yg5CAnG+SOnFaT8Ohz+L+0JZno4xW0HTaFhcOJIo6FpmMF1NLGsR34zXo/xoNIQM
9cZwj1yitl/1kkvmKhTCC/dALnQcVNEF0yNNQf8zc4CMLZj4ZPtcxLrj7CRNtZbS
NbhDIGYm+PLTTShUxLahaLP/41sVrpLgjCGVYZTzG17vinzI44QmYItAYUGBqlk7
K859En/ni7Ufx3g0HxE7CCjwEpYEgcEEvvcqg+Iw3jUsjed5B+0Rd8x6s9dS5MjU
qDklaMX23CkQLGfAQ0WQxQz7OwbXa6fvPHFiZUrFAHzK/rYEs6EZj+Ju9ocP8br1
1gse73znOvYtZR/BPa1lbaOaHvXfdPnfI1xrw/RBi3DRTzlWfvJtLpia1i//Ku61
erWkGPLQTAh2tjo1USlfsqBNrp2ZDlEyHr7+DKQb4dYOxmwyJcpmcCQrtxZ5hFfT
w3IxZTgYTxR0nPUGc6XqeJLHsX99x+xaiYcGjW9wGeMaaY0bIk+628wclT6pBlej
1i5NXWeaAfEQFvErRvZech7n+eE8TPuH1FhAnRsmoZS4lKPuGV2zMSlOwd7mIJQM
j7CEGjfnvxmKcflCF0T8Uk4Ek5zgVmqRqf2SGdKcI594HCR4QvVxgiTbJ9tUTwpf
wet2DpGLi4UiW/tbfFktEplwo5aDhyxQf6Ih8wLlQFu2tMiIvEfFmrc0pA6qZ7z3
Idco9NKSaJJz26ehygf3iCGK9ZZ3ZkIVk7p9tTH4RBP5f7HhwUPqDCGCaLVCOrp8
OAz9u22F3MueBJTYFPk3pAfICUBYKjoVN8Gfjz1qNpOUkje8CuV3zhmG+byRUWZB
CJw09O1Hn9cejXj65JJ28QImNFb3mpXsp/33nbz0I8IPRcX9obbr0nv0JxP9sOlS
mYMEbu5F+656f5WK5swGNIIwTtx9I35AHcyNSVZWRD0csEZPl3KJkUR6LYMIbzTs
BgLn0w4DzBw/3phueYV9qup+/XhUkqnZxs0azvglfzmjiGWwjEH2f83cTA9mX4wB
LzasV6KoUPlUJJAAY1kkknjAG29rXHHI6UXc4CUuszi0twfnMYiNqkdUWBGzrjVm
l9CKNu+CBX9sNED6C/ihTCeV+JDJiDxoMb0FfXDjYhjDbf9RIw6c/exHDA600Krb
mvLr5jU4/uVWACpift/12KZiXP9dphUTp34u8wuv++YkSRhYBFaqrPREK0HQxORC
0fJy8HCJm/FdXR5oHCtMqd/wlVUv9LB39VJ9mkTZbNVEAIgpk8jSdGsWX7d4MMkw
ouYgJgHO/dfAzsuQ+vXpl9N2PD195U8601i4e2ntz6CbPvQKk5OvBbzqvW+rSSMi
9t2/KBT1SX2B1AdaBvzBPAwk8IRckRydNVhPI0sUUmn1QD8GBaO1NmhVg/ef1HAa
F1Aqd4FOWu6Y1QoMVh1JETaAwomsAciyJL1LlQ7uvzwWee2tXFOUzqLXs6s3mJX2
b58Xx1TjZejdKjXkiQIzqE6IxCSYayDT+Wdy1DMLVjeTD/PVT9thFRgxl98YDNo2
surnKyoiURtV+377vuN+e5q5SMbrSdg3ZAIsJO66TFBzwdX9mWxaE2DMyEd2y4Pm
sO5ZsmW+/up3StfLRxqs/n46PJ+frn8VbHYe/l43V16Htgg0MRBZ/rA8/kTVpBof
SvPyOVOv2v0oQAzc2NllvmViJDEu3pnGfM7wKFNaEB1xuzvlfcEfGM2ikIZ/XX4E
gS7suD9CKKeH74ECyWRH8i//VBS5v8Qyum3pa9/ddORdteLiL0Je+2vg3oujbbCp
Cd396VigROuOKoIByrZuSLfqDl7NkxKlLA7VNmVneL/xMKKjuWOuKJXuHemRPqKf
ni3DXFMFUJ9ip1DzIwGX5l6rwqgHwGT6O2k79q3Kuc+G3RA7XTSjE5/xfonHqqO6
okYchsjFwX/YRGCS3L8+ujyb5blbvVX7/5N04bOMMvehUSgr+Gxmnr740TNhRVCJ
rDtWNtbA3t3GBjmmoqAE50n0KK884ic9wL4JoCvFr0VX8rrRrSpeZ6T5Okqcyz8G
CZsFEl583fKvNpJzQOAOR/bTXmzg07G5/0qx8dyT+YE2aKtun3373fSgmZ9Ed9eU
FEs/Y30YgO4BiyhYJRgQs9AKYqa5lEgnaKMzDQTXkWnALu6fWR6+z3ySU4jRDS+r
S8AXqInODsUTvfqgnl51IHbAuzotMP0RESJoZli5bMDoN/zEZBK3byyZ7FzzmDrj
0cLx5G3VfWNMmzMUjU6f4/1bpFwVHef744cLTgp+yOpr/BHFt1YiJLyDNcGrjM28
m2/DRjPZ2lJWvX/qZer+HZgZycpZlE2qNbhBhYZrDF+Cb/3zDe1AJO80oJEGuT+S
2itEhUSxYLfO+ItuqxQZGaxUk+f+9FWkGqmKKtpdB6EVbmFMCQneHm21qIxA2NiI
laHYpvHR/pHHAZc4K01HU93+sJl5IKdIec9ac7jX+pR49dOc9dWCVLiSTxxVUdqH
4jaHuENI9xROhn+F44K6fALHq6Fc4gF9e6QW6U5/Emay8XozNKFHt4DKUJFQe5ka
SjqmCykqnfiV0xAM9voWXe+bz1szKKvNlBLkI+gtb9IZ/Qx4wNhq+Uc7oG2pCH/5
XeBDetBqFReM2SC5AfrIaNTOmNpRAuBUXBTLTpb8AUzQCtm0O64Lql1GOUn3lh08
+if0PSGXfRiMQnQNz3G5uUo2Nx1yCBy1FQXdSJXyosS+i8AXjlExjX/2ghxC5CVv
v2mYHR4jqAs4CcZnTnWUthb4SRH5vBnGb45t61Y4kGJlDaERMw5ek+zcW3wCM55X
FMXDwGUtGUjf5a4MTAdJ2eFRQ8iRdEzTQWdJs2fVvQDUUyDOCeLG6o5gAX+uroOB
UWYag0US9hRtcMa/v8NBbx1abxqisNLwphnG90Sz4dV8MMpResA8P4QbyAx0aF+Q
BpTllUfN5oxsCoKGHKCUKa9uNWsEFa4QlhFd3aLSJDthVZDSZ9O+ZkItKZVZM8/g
9npVZ/yU6FWyJa1u7vlQzqpu8k5v69J0S9WPW+G4gCn9LWdm5967Ae4A7rWJ4dpF
+Frpu2Kdso9EzV2NdwmH5Djzqu1moX0kcSnj3IbSRiqq1Hu/L4ObF653Jp3JXH72
naZO6zaQkKNMNz2iGeP0BJxi3xePtqk8BahUhfuMaCh93CzgLy6afBt1IGNQXWpL
RVryzuTp2raPNgCngmaB0vZpMI4LoPh1wTvW9QNk+YOHH2423YQohcpK9yMIDLwP
Al1+8Gje5jeiTXZywtbIu4ocZjDbe6KbSMB/Xiry1+qoG7YRf5XjtFXQ8Yr24aIs
2AFK7JRLeqNGWnXciIdadHMbWXngdv663wi/je6O6mLBaMaFx2WoruO7nxfm8lSv
s6ZbyeyfcJPiRmJ2SKMc/tnNsPKbjIhiPQWBydwlj6Yulsn/xaFTQwcUAkEM2pXf
OZ/w/evjVu95g+/GYkioUNUabSI/6wM+R/ulgu6y6cwwcflcNhhcVpqfMdSZjWbT
l1/16vJL9T8Pjlct+aRVYk9ZByPcTFHmMnzJJAGfaidWy9qEgwzu2lk2xAlfmaRz
C+ZdkE/OfvIg2cPVnaevbqWNBiJQJSPM/4bmKc1ontCl4nJvuBOjRVpVONz5aNW0
ppVMuANalfiBj4KamjE06vmJ2OcBHUEZo5abemVjtMEgeuXP6XdluffiivBivuPv
DB7K+Y34GgPxD3UD7c7PkLc56enxhvxFDa2vnfpDmNHxbrivmN8CmZMiZtMCbqMm
fMkzq2WiUPKm95hamlyhjY6j69vkXwpTh42izo34V8CdyyzjHTKE/Gbu8Y5LjI+k
FABmt7u2cU2AsZFQZPWmdeW/VH7ZR1QYRsuLB/EZo+DmH+J33NEitoxO79lAne/v
cy1x4lCwDLPnL4WvpiwCSuP/S+nFlVZhg60FL8PXmPwdYap4VmTps7q6WhrIfW7E
eILhryN1A+WfRPBHRj7KV3r6D+4HEr5FJqohHHC6Gu4+Ondhh5ZVr51FYWzVKrgA
gQFKURuvB9cAVVS269nXzpdFX9YQqgjUMFg8T46sG6ktlAWOuJXVkH5oR2jtvkRD
pLW+r1ObRfRYIMRb5mTKOti8n+e+4piv2jSsYWnH5NsikjwzYGqwuPNBVX2Wq/9M
mzL5neQWiu8xjaTUiuPH47kiHjWQ4IBmMR2kDfLp7h+E6xJJs9MJF9Whs8kaPPMn
C4ofqfj2fm/AZScJ/H3qh4JBPiL7sshvRrOOT+OBiy99aV8CT1pqkFDaCt4iNk7N
nnBEd423igUd+FtqDzcvlZUJuTIoMVXfXlmd67EZAbJAZH5pVzbNnK9wyrySKt+N
t85brzpTDnIji7YQ91MHx/g9J3rM80OE7K8Rph6tjX/C8MkXS4zvrdQkNSgDdOpK
8Y5kVNSoMGbrIX6au/sPeESumQ4b190et+6v8VPilKiPhZOHs6F0ATpxmHGBzd5N
2HM7CTB9B60uA85SSrQfs2qfs67XF3FoHufyfa+oBWkdlF82jHH8hHo/ZW9E/qa/
oMM0waNco7RlWnJ+UAnDB/s1qTHfR1BxslPD2Grq6FBrBLInDMWyoJJXHsA5S4Xv
W6lNWYTBRulvr1nmCyKz526xqzcJNa0ESY8TiKBURj1IuiMmCffGqzcfykVqQyG0
9ET/yAlRhd55SFTza8rQJQGarzGVFu8Rnsk0YxO9KKklo0Yj4mlLQpFquF+pzgJ8
ncz12JMchllqkb8ttdheyrjjl86WqjfmkgCt3VIOJghQizAO+nETTIirxWt8Atnx
5aq/sd8Vexuh0BssFH13PQccvFYW45ClIE/rsnSH6rk/mMlM50B2aOaJoW+P4rVT
IsGPdE6pK1/sGGTkRb4X19AvBDXhGF+r8v7EnUmdBcqFtQjrGGFIG78To1xX9M9S
8t988lBenazL/u1lI+qU544mFws69IbAkGT2xHv+vW2+Evbvy2RlTnsevn/scdxU
apa1mGR5uckEmxAJhOJOspNjsylgsZvh6JAS/Td8W2va7AjURiiaCp9rU1wwoMDM
2HG9dD3/J5d4d/xZjtnWnAo43/VPTVk9Cdun2dyhlgG7x3uk9H04qvT7dDrpi6HN
G2rY9A9tZqsZJVKnKuggjhMcfRZqpVFBSk7P9YQOIgFUlZvNer1cT6UHynuPc45f
te1z8BkvWfnhXFcFVx20DdqeHyiOVrmntQoi22igZQmF0MxzhozHdARuaPu7OgE8
niAv5S9SMwxBJZYEj3A9QilHJvs30zR0UIeIm63+A7NZyXbzxnlb8TqehdtF+TjG
7p31x8ynj62u0ScBw9Uf0NhxotLVgZ+Ptp7OMrYWS6ZQDkSBEu/pgXDm8aWoW6K0
Do0JTuy5B+tBTOJnkAj/gJ+bzl2ZGRo6lMA2noc7fK5ZNOF5YTZxO5VXAZY5B2j6
rQDDrFm1M2yZ1nkzy0OHclasrUBALYu3bCCzQSROkXPMNeN/+ZbAZx4nkYGmxKCC
DLFeUa0SVgcryuh8Y414hwQMSd3DSbIGPl7RGgmn97l9syXHd93DaGijSCfyYXMf
KFTsxElcyyaF8mAadp87RVRAmqzJCju0vA8mF2RBubAPU1Frr9F1uan0dRN9vJb9
n2Meey2B41KS56mhVhM3VYydezLeHFYv+zfgiGnNBwST0KTlwKefqGuhD6QKhGEo
N+J3KfEhQTa+XpgCGD3iE4O3nGUWWzznYkk8li7aYy9duLvLZfzGc8LBKf0U5Znr
kOPd12JOL6XrTosqtGvbbOqtDKvNnNl2549DUr5sNhKuyqQbPrHMNrNTzxyXjjKd
mgBW16lDNBp4eHogCUD0riS9+LcSuMcL7UvQQstPCqwa8+UVe6TeocjwKqCsYuCS
ps9ZomlsKFuM9iAVTqNpZWL3m1JNX6nqVocPUnPP1ggjtOq284LzaKFGotQYYsZc
HFPbpNxss/ilDL4Ju4H6ANOv9fQo4sfSiyeQ6riEJO4D2g9xqAQlrU9MAKsnbPgj
HAaa1bW10yc6NJx5VdesKd1zB1CgGSATwDITR8IrrHAd26RPIP4w42AXglWo7r8Z
yklgfT/vjQA+z4eaW3TPRt8bDrfdGBhfKX9qCvl+7IZLPbVBqEmXA+D5FbOq1asf
VQTGCE/H+oIrNQKjg6PAzYzEUtALmfxFuT0xMpZU7AAaj2vrm4e2m7pD0BgYoCfa
l2apcSrMlx6ZFq7LPeEHcQi1eB2NLjB+SXtD+EgzC0gMLzYaoRw7734dMq9qAmMN
OmGMeKQhechmO7d/GMBatBL2Yq83ssCuPSTKxo5XDIEH2lMlq3slwR/hz7DRhXOQ
8umTXfhsGO4XHyaYfkGxIc/sGRiW/+JrSUaQgkkibevyDX1TAI/BZBJ37XgIwXAY
v/04sSs8zdOATAmEQCuB35osBpU3n2CWmyJ/rvlSuIaTgG98m6c/rNFVeiKvFakS
O4xJ0a+hJFfJlwsqCcrSn2w5/QRaCGlTXOL1XvU4WwXwVdXjeUtCAwmobDUXIumK
hegNMRo84jcLnF2abbYJFqj5f8A+ADD7Wox6cZP09GNkBoh/jaOWHWWuc3eo647B
dOUZtwV6sPAijdrXwadKeQmorodHvnrkxzo5jtjoWTTlDPtujuppb+Ppux08dLRr
NHg9BWu9WsMJ8UXcsxBbu1INOyV+bYSTVyf9mC2vPq7w5ze+7cEa/21+2HPaiJl2
vjZ0GRRm/QSCTfLFuc39cQV6oU0V8Ij+24zgTO4VmgBeeLGCsMRrejnKRfYdRThm
tTHN5awNLNZrzIPO2SYThdi6Y1a8M39RuYOc5/AWaVdP2yHIS4jaM0P7sSVxIsPf
/VzpJWCtk5EDr0PxBTasCxtDy4MHcRsbIQiwOg+1DrBto0w5nG9TugxYUYVeeMjj
ztzbedJlcsgSFtV3bFNjKMudffsgVng+3I5U3gZhgPf+ENWAQHJpiVDHHlU0bdIE
YYPE53jH8xkYcQ5ToYFqoWXwn8FeugYXGpkt8PicUtGiIhviNcUmhm4DiYK+ZfEd
DijgxnLHp86dxt1dcgbi713EtwM1j2n3xy3yaq5Ntfct9v2mQ6HD//r1RpOmERUm
9pwwfPdrX9yBRMt0XoEM0Bmbe9l/oti1t1bkpI6If7srPJ3nGjqw45nIcXLBApdK
FumGUkmddygLB+Vx9gx4QWddKLQL2D6gDWLbvTqrZIx6jL9Xi6xJsJXHGGHM6oLq
oef3O9KqGmw4MvSkenl8Cs8R9jDd92UYzyqnqFM5pEbHkr5QxZJOBfdvdqd5TYal
qfKKwv305u/M7kMVCdXmWpGrki8Q8OM5DTFvUQhrOOgCqnkJx26+cJfbm69NkS2P
uhgcoLSMUVfvONbRjRElqWFZblVLrbt5kTcRLWXWLl6tOwyoRek12TQAu2tAn3hi
qCjiQkZtsmAYKZlqK5U8lbMcap+1ZZsUfwMoUbjSlSAT/lRvrUn0iNAj0tOroIQi
3ltCNh7MIUaigZzLeut6AI96QGdQfDA2dOl3SYwKUk9LX2EalgytbPcw1heIy8lX
Z2j7r49MM/r/f9ggQ6w12MOMV1ZLMSZW5TqTkQjWi37wrHa/TAIWaJZNGUxkLl8M
R//os8YwrCCrn04oO3cRuMJ8BKBSXMZnRF8AC3CdYRAbwBd/V5YsGgziecM7ML2o
9TX6Qm8bx74BiLx6Ct/tDogvR7E4tpARN3HcIbcnPjSKq0Bb1JHQwAogtPGGoZUa
bLNxjFtADz8gBaA4H496AM6WDdiObVnrPWbTpxQVdJPnkJm4vE6scrC4I4VARH/a
f6OoCbhfOAjY+Ew5Kk7/+u0gG9bZX45HkKxF8ESa2Ay8jVp1AbSFmeJTZOVAihWl
BqoXxEJWKUfWJ1q0tj1rLLZAbx6ebjVfpt+ESN1u3PqTsSxMadJD9orZo2+Nv4/X
I88W9IHdOMIF3ZI3U3rfLjubOPWQlh1rG1pkByFShchp7loYyD8Y0p6as0TECH4e
Xd9Dw8ie43WAJJfY/2sg8ZZj56q47dSmJe1YcSOYiBcc1eXJYHIb7x/1HG0vWtuH
AAW5IhEEZ3CiZiV+st4jHQN2J7i4yB9XNuVUL6ZDVATrNa5Y0tYJEz4TQbThX+ND
+QCXhzFbNXa+O70Yd0jlj84CSLagROeeaWILYLiaAm/cUv8WDWbMsk00x+A/SURZ
bUZ1ivtyGFIYyHiVY/qi0bgN/HJR5U5GKd82hi6izfv8mp/DKLAPsS4JuFiEai6R
o1Hdj1Mu+M9zuAbT+AuDAT8JEt1S7myOk5ZATAKRf2UofonPKdpR3sDl/QtkMnXH
6O+38spktSWebSOaAP5Wx3BHRXAf6nGDgJa6eAxgFLinQ1156EPDDKh/pd+/wenT
+SZzogRLO+4VMZN6RUBub+1s791bMZ6luej83u+EUWxVXH8NRMKr2YbN8qwK/9Zq
8UJpmdih6bg+kXOv2Lsg+EKp9oI/OFURlau71IFa9ONH7zXiS1Nppc5o4fOb+M7e
JSwIEkUBq3caqtispDOCgRjstzMwRYJoo60bt3PcGlYFM+0NkoUnWoUZfJ22dydQ
kfhsbIMqnpBMbek5F5bQF0tZZkZcgimBxfF04eh3h4fNtOYYT80fjErB2I9yt37N
2YeQ1Fo+r4DgxXYncDhVkSoP1TCzeX79rDvO8IvoGaM5wneRMSV4QL+lAN6WhPA5
sy2ygeMxlqUgHtxv61jsXx6IZzWgPmIXI/jc8Hq80+rPYmpSqVLWfwbwldpe0kRK
vIVvtwWvVht1oHDy44rE0t8fX/cK0Gdth+PZZnB02c11KlMyJ1RaeBqhMzJc6lSN
iAkhLaF2b9MUpQ5oTrdx+Q7p+yNiz4mybEs41KBjMByHcrklhA20GZ/woy0Ca80y
2YIg7LfCfq+fI6V0b4o6fGnddeGLcqtbL47A2EaidkwsYNvuPiYMR0GtZ7Tb7iDN
G7ze3n2VBF1bEsMlkcSid6qITrf9H2pYy1tjRqIJKud4TeLlqFnHxmH8ACypsA0t
vkdkECCxMIgSaoGjbuSkAYrnM1PUl7n5qJMx/KehoaBf9quzVyOmTXFr7FmtPizN
eWvk3X0cwDXIo1X0kDRU+A1NS0RTbSXtCWEV9mECmmHsm9koh7+qYwSE/458xyxw
XPHwDo5Mq3qaju60rOG+HgJRzVLJGlrBi+1k7LjZ0ywkyNoQ44H01paItiGcEN6n
LRNelpn6PDM6UvcbN4UjLzMMDxKXbT/uiNvbNdd9lH6XT7HqjptNQXH5oqdfx48a
x7Lpxa7OnS8JAxOq0xE41q9P4HqH3F2TUV39GMqrBWobVgr1rJJBSvlgO29BGh4v
GkKjj2jAgeqp6Ozacv4udmdhl6WLJOPokbaOZxJ+Soz6JS4557g2Tf74FJb9roGH
sj+KGp42g5+uroUSl4VMdJ/SZe+YuKX0rttcIs/IcOcM2oWR8lQJ6tuLLMvu5/bN
jYtn9jsuZdLP/RRDM4d3F0KEIysP+LNAihHc43o8C0AHavd+NMSFsO1G0v5JOMGz
56/rDRyYyO5LBQIS0uoxN0m6y8y8CCAmcP/awRBZjNHQOc9e7Iz7QQ1w1jLkhpuv
+N/3d49BZB1FLpsjQN9QKR1D5yBRbmm6nHuQCM4Q/PcdZlvN017GHZ+sIigSBVHp
nv4MjCJFmsqQ/KU4PpgXiJX9uklsK0fgQLEyYUzn3CvsYsFlhhcfrry2rm05ZoJk
s1bm2UW/QClZ6rvqt76S2aS6B+1fLPzCAKzLZbjAA3akBJEdFRG4wk3epUjf+NOx
iIbd7Wd+oUN4O5NZUhOPr8uFFXAc2aENFxEN9QnW18zoPDqv/p+AqQFLVP1Yz83F
85bSzGBlCjBhDNDmFSliGy2f+JDxByN8farwH1+3gosfbLLn7eu6UthIFx0Xrdbe
3zi8lod7mpKtr4j4F2E1SJqeMtv5B4DX2VR8Xz7obxE2g935/bkiOAgjEmUjbvbM
KXB/Fx0NYEU2yWyK4AkBfk7VGvutqZdLsBl+lmAQnJ1sK7fO/qDEr/ZxexiI15h/
ApYldAJPBO58xNr1pUdiVk0jBWOHv+0ZAXfprbOYCCPnBMb+iubcy1n9O1OB6T/2
vkISTMLz/hYh6+VGwugUrcw2FuwSqD5autZ2siO7vWIQvbrCetiTEM0ofRbm3of5
41iMeebviQBnOKqmJVxiiMZ60ABedXd6eK5mtkRss1gT1KeW3KqkfMzWSgpjCvWt
3hR05YHJy8etDaGN7HTDD+oISSfZPDWTTKnhs8B3xYsB+qxDaoA1Siec3bDnHnaY
BDVCNt9b9llc+gKN1HaZSvgdq8+P8Z5RB19r3Xu2eMOzhx/4VrBwTeOTB1XWpWPR
KMZk7zM/y5V3jP3LAU63Z+bTUIyYDYOa4KlBLYg2/KNudD+94gh1wjetzDNXGKK/
Srv8pnRiZaUPfdosuY5+PIR+bqokft2ijDMPL88iep2vIAlceHyRxlRE0JjvFPzD
RS+62SE4HGWpIYFasITWONfpkPDFauWxw8MiNG/yoie6MHQWvgHgWGVW0/x3ABlL
rc6se4XkbBCeILC2URiCP06MVLP24+ua76SN3q96d7O8mEQ3r5h/JY0g7QVXGBbF
ZwDs5lR65X1SyR4oJcngPJ3zRKXsqMd4/DqvoWneAGwRKhUtrefNUoBLhh16r+iM
267VQaYrM4NYfbNpnm9t0XCj4H5ND8fXRfABkcnzpxGjCFGv5zzs5wINHOyPMEbG
X0kVsKm1PcttjpkFIlzDHgsAMZ5gPwMHVlTmRdBqPsTSW9Xsq2J+4EFctdxKJ18n
/d4HyCeZ0PivdnSZYIfa8JVgTaIr1WzTCSjvqHiJNX2qpVi3geTnqbQLMhe0lN7c
125Vcmb/t79/JUAsJnw28/DpHx1vgqGSkb1o6Mvbqlniw+rPzSow44AlfreHF9Vj
z6OSE7kg6ecK6JtLoxKFtnwoxcoSP9rqOLDCBS7c4563hTYh3wN2UfaMzzdTH67X
TVmw8ygU5Ozej9fmUPYex/yVNwuf7ve2l3L2PkU22zdETM8baBAwm7BkCToslJBI
26EV8kmEAEn/OTAplbz0tFtCHLel+uVPg1HfATg8ZfKOKKxF3WdkpTSRr/cxyx5T
HCXknfCNc0v5Z9xHGnfFa4BhQfmDyy9pz2B/Zpcmhv2nS4/xk9HpdrdH183iDJaV
FDWpW9A8iPvZ2jGlR+dlyRUd4UZF/NryqytqUKX7r9UqfbLss6LkKsu07ghiBx1/
ydV1vnNS2Hok9sVU6M/GfYqFqU0QBnAv2BzOFJUapmepFN1cdUFCjQTWZ3FrRyPB
qEAoYLUemVmlBwzfNiNiPtjQvNc8OgpQZ4/bifbiDbkiy67eFMKCFASrAaklcVaM
XrbYZS0+WfXMwpm3mz4ysUrB80LoI+UM0A2WNofXgbvBjWfW3atwXeidGGDJTy3S
yrkD9Ffy0DFvftMYlJQS/QIHhyGyOZqM0p5npzRK8f+9sz1aZFZZTEnJV45DlhnY
J/QnIjKDkoXonZsmY78kyDGfV5NFTgP7N9fkPfhjbRq0DWq2LSwSCwAYbgQaDxuM
iVTuYUTnnnaRSqdLDR6B+8/9fA1kULW5Z934rEyAl2YmRTqWgZn83c928h0OSZQ5
G98omyg0eVhDn5PcZPuSCu+XLWWD3LYgFRurxMVBc4dkXTfSbCD3ZaCaTeT1ICDo
48KerCrCC5zABDyeveZNVBFap5Xvgwnh+i8LgF2kpIDiyrGgwMNfUl/o9TCAvu/1
91U6G0UdtBqHaLwYt9i6d5zRSZmP6r8NNUS0xyuswRxB/Hb7MXd+VEkcKDc4P54r
r9udOjLrea/s/xlKydVIXKDwgGMOIFouKNEbECfkSJQz+f+SglTy4C0IoY6yvjDU
89JzAs2rMVjCj922FKA5AzLrtnAadjD3SAbmPa0t7V9NaKDu4N/S3mD+FYvYg3Kb
SOGzsDO22kGKNs+IqmuSGINvv/LkGWeiwvSvmO5HKWqVkU9ZPZmYM5rsoNEtdVON
BqTbgnDi18t9ApAsIlbjc8So1RsFtSsu5KCrVKDtHz3HVX2rz0Tg0Ri2NrKEJdxE
j/iLyqEKxrvEsq6I2ejnLs3heb+xWv6Rhxqn2xsIvkAeo5/x2NdOy+wjP4j6WDsv
I2W9wLYBZv7U+/JZgYmAyxTNATfRJsKldBi1hL7G/vLNMnJCyqwS28xTtlDI93VH
RWcxmkvfS9Jhpak5BQaeDmzZEaAykwIEqF9SKfPcyC8ZUdOx3GStshdzOu0wXcM/
LqEt131RWfigz9mMBJc49L0zXXlRz2i5suGKFswSbtyDLfhxkai/SvtYFROezNUP
E+SKBAuO8U26HsmIWwlOJjiJthaadZQyjYc/zw9NZLc0kA6HUaL3UVT6lC4WeBhy
1LIfBST+JR2jLL9aI7VaWpD3A+JheRnLlXm3lyL2mt72TouJZjrjVJmcTAJd5fbl
x1Y3H9Ui42vf0dHVqSAkTf5dNz1EYKQf2YeB1G05LzZGgHgfKuAbIBuk6F4UmAd7
B5jlgdu5EEb2W3qRfH4sSYaq76nYuLbXVkAsvtG1SnzIWLxEj0aqK7pB8OcRP8Nh
R/3tDP3e7W13zsHhKDfmo69OHKED00joQgrrX82lo0612R+ErZK+JswvE89krTPO
lZl/l6adRo6LaKSe0cj10rSaPB+jE7A7/r0zcJEtJ1yWbh8QRO2nim1I/xTGz+iZ
J0zczK90H35mSgaMJNPbcqMQN0unKlVJdW6ZZW8KTVfGMCMrNmNvMWsiNIAvTKq8
gMiAsieoA2IhEmWuVpyvRyTcD51NGuTPQRQC9Ba7hFHFQMiz4KQAIAeoJQTPhBCO
lx50e2MRhLKlcW97uvmX/ZZcsFb+AV+Nh4xiAyUSB0+3Gb0oYCrMmXm3DznydGdn
ZX1m6hS4PaDIYPzPRCvLXOLmaVOt/lGaVt6Xeafi6P61M62NhDP2c9OB43ndxxLD
EeOxDq+5jzVyeSjLYriqA7+6qhJygAOQcRBbm4n27Vtb5ONOcdNn0EiJ3NKYsJyJ
Ly5XTwb6OR2t+SDsnvbWd0/l8oYBLusf6n+cwe4Dg/Dj/1S5KpU1Rg/oVL7HjkLp
4mQGAeOmetlFKvgIku2C7KsF9FEUesguIoGGE8t/881M9jQZZU2Q/OhiCU/dFXMQ
ycf7nj8FNEU+cW6yLVy9Ya9mUO8csPXti3OsBu+oL1/u29RcUzcSD4gPGvMheu4F
a6dfloNGZnHRNP8Q1SkPNNe978ZJ1fh4ILPA3l4USeFZBKCBrOlJYe0K6SQvYmaX
uhjtgGlPr6bLg3T7zXPAOvzp/E98s3cYMsbCgyo1wLK+HCyjUS4eGSGRFvP1eNcs
UE4v7GkXIYiAH2QmS5QmaKI4B2eQiAGhdaqmBKfYIeyLdSEZ3g5szK3tHdpYbyGP
npx9NoMVPVblj0IOaZsa0yhC7BbPTIHfpyf/XT02kdHa152b1ZMwaDU5fDXlWUCm
5QI/wjmgwCVR5ehICj0SD1PNX23PH4qIekjKlU5oEza2/9XtOhh3f46QJoB6HER6
eM6Qhrmzxjj3pWr4BTpce/8udYMXzagLy+vKR8sP72SUDoE3XbUwqMliIKJkPe2l
ysUihX7klfFS+98PMWLZa72Mjp2xo8eBIdf/d0xOg36jGpxkFqoV+MUAbtNeuFrD
orWekKSfKCzEOzTNNQdUmE+IRAKtc9xlBOMWbYFpdbYpt/akku2TeAmYzjBFMsxS
AF1h2rXijCbQrNQUGuxp0yUlbjKOUfVh4yRzU9wWgzNHx+ZTJJ5DICs8JxUPD0J3
FvBR9/b08+bd1wEcZZmD1sHcsuclg1IL5gtmcb4NwyGhhG+d5CRv8tKdSjScgHQc
GbF0IE1BhSi8t/6wqZsRXdCUeAaq+KVTknB13wKKHYt37BL1bXQ8Hvb4GwyI+Va9
riQ6gZ/mBravTh3/GRZL2b5T6WgpJYSnzj+gXYSYeBcNlCyLZhGfR7buxQMAE/+A
WtyRv0T032FMSIpJGTGxo/XkCYp1zhr3Og9DfTgVsGIDDR8ZIHzQ61Bl2nGmDrP2
8xD6cwIoOi45plW46mUEYilHmXTKtCKUEusoQyfIypSKOoRHmwdKefITDgFAqbFU
UCmbSOFnfj0ft0esreVryBHmcJTJgcDv0RYXpiVv1vJZnXAdp/NEuC2939olAS47
ozLtO5n4Psw7bZUqMCukPJOuH8UorqNfp/WpCACoNcs/v187i9hY5CCcLDZQl+Fx
i4NnBECKdqUzS1XD9ZEcEI+aOmTRWYl+mIE6aUZ9damLXHIqB2J+UFXcs7QH6kx8
jiuYXUN4ey/XHODEhufAu50N3zNsYogU/kyIte1yAjjVb4IrYiPITCDDfhsrT0DG
yjOoaaumKpFsFEDaGVzogS4USoR5PJqbOKUvNQwBUlu5CWQF0nluhWHLgBOpdo5P
Q5I8x/BgrITajvWMnNeDAiKvzTJfg5beZfYhhi4/L5Rj44AaH15YJaJy4MxvX9PS
JXcRnT8Mjgnqhf+9jDLBB5QmgkShf9Okq4V1FB0gukOeMUV+bb5YCiphOueYKi1R
JetkRfIhpBgA8roAnnrEkSulBQhrnqv6gZRFL6dyw1N6quf+6vE5+hLng5A7sqw5
IqZubmk+yv3jItOCenwnaPRa0VjYkYPfLV7Gf5a+oPrnsRQj5h3pgubbCGOacb7x
+r/ETyT9xHEk/E1fIecAOMnKpuJGMogCWYuLacCKNLKJKbu9FT1sVC8j6ah+8rkl
ONGuwtt5d5ocBbJ4G/YqrMWlkjKQ1ox5U2OK1j4PdWEytiej7tR78u+cdz3tWMP7
XI/zx4Vx6Ay4WFfNcAw37KcL5kIJw1M0IVaFm56m6OtaY9vG9xinUfuN8rDzYxYJ
myFv/GoxQFxaFAWTRDg6THtHd9Bx3XCr0OS+yq1+iiUTM/7DSMOYE+sQ9CsTfsXm
payJk+HquKOeAl8qDuFQ5eSfZGQGKXCZIPKZP5GRIgzNp8qhwnCvsmSxxFIBLns9
EmDSN7hwlBYmyOKb9TtUL3vP0dQGEi7Q9m3/bcNnV2iOGs8qipsjaD7knIB/Cjg1
1/8Lr/2RMtgi7dAkCLAVtaomio1E1BlsBYsSaa6yN9AFl6EYD2Bo3ZcHNpcAWVU+
jP6EIFR3mvhHuJZMOe3uKd3X12N4iq2WzYlB386y6YcaJQTaV+o+5lb3rUjaKluO
BWgGwg+KPtzSAf+w3N9tK5Gb8J9Zh8sW8i/SPJB5XNz/2O/L84ADuJOfR6LhbMHf
N4MH7fctpaNYw1rJWugLz1jz/LvF688b+DShQh97PmHwIaSzm42v8/d1/9fNAP+g
krvNlvjC6/sOxGostV+un9ngVbP/0n+UMl+xpfRBbDKtqXU7ddVkFpLc75qWjmkv
MSgGpZvOjQUJ9rBXvF51kE2P11mEwSEJTgU7zjvSZZi+5RUMUlJU0qgsTyoKtzWd
QWFVqwiO2EVVVwWyHAleGaO39QrGASymNFk+1i7v+kK4iiSO4kX+wJ2OgithdIJH
F5jTi51N4y5tpq9Z3Fm8gsLCqV+YSRif0i/Od/yx/wXll1gLtrC7VSagcEtsPace
Gxc14pTLM52TdeOoo8voWQODV6IFrS3iDke/PnW8EyOl1gM2MG3iX+sCMCdCa0uS
UvFiOkcH6ZxJUv37yrt0kUuwuuQQTPXz1DRqfwKX7VG3yemCzzK7+tgqJg4YbaVm
Ft3HYWiw/zDIUYagM5FMHpYhPP9w5H+5CaZzXQn/Y4AbokqRH2EHhMktTjlmX1uV
33P/PsnLAsqMDK1pPWsZ/vyflkg+8AyxfEBBkL8EQgphwkETErjdlYyPtYCAk80B
an1GnMKzOMpkLGjQ7sGReBlxxLw5zVw35ZhkE8L2So7Z+/oxpGuc4MOCSRR6AObT
/dlcKtnk7GYdafW4FV/5AiFGExCjxT5GvZ65AYjArQvSOoxwElgar75NvFOL03TF
l8yGyd+TnTT09xYUeEOZlKg1xJqaFDhtMBOl+F7JgAcvs/JDlbQz64Zej5TIy1ZM
R0k3Rym+6TotLmTHIIQXKiwTsPgTkQzFAGvmrsfI6SFtUCPFCCTTZ7uwy2QSP0tT
L4jro9Qlzj/QYz+JyJ6M3vce01h6J2kyZShrzFjP1hAlSc0f+5CQv7Bf+hFgAhDb
Tf371Lc95mFngZLmjiRfspVIEB/ORSw1EUaXwkqkyb2dwEfxrHL6+WFCN0U4QH0/
4rtK2LiA4Kbp1Mbt8i3C9C29y5O7N1ECXFDm7ni27qGBTm5DHVErPzlR45uraM0F
RV3llh1IppFXvZjimWXv05cT8mjiFWVwoM9TfndHvnsLmpq5sikipw05i5FCuvEg
LYvtfZDl/tulPnIOPEpMT8DO3AUzdxJJDliws1XjnJ5uVAZybtl/djbJGh/Xzy7N
S6QX73Fd2Gh1/IDNiIXhwf6I/EgwJZ/LTnH9ERRb9tlOj/UgKy4oTfVBf2GAyH+9
XQQwBm3gaEbUvMhokPQ0cOQtgHOZJUOgvGDdbQYprwble5Uf+KCBwwpbz2mYScYc
F9HpoMXcjCErK4l66ZRfpT83ojwk9zcicY0dfr4AGT+1J4yDblj5UYfPWmN0g0I1
E4OHeMJutnXmmhbPVHiFkbBp1b2rhB2MpcOaYYFFajYuAGePia38JipN2spuOIYP
ijCDy43SqrsFp0nXOFUG8Z8AWZ5mvyxpZuYGrUAjY1e4iZkFb/N1AJaFL48csgCC
Ldj+CMNlb48EJpnVqte9FDI9LZhkO3K86DzdhzWcIWknMTb/zg5mSK5qiEalx+pQ
O1fuAx6eDBf8wvID0OGGQ5Z5d9yP2jVlgKyGht+dRdvvtAQrYzPHqJnHt4vvIjUE
cRh7zZVFxJ6UH9oZ8TFnzKuhXmB3UGN5ypGy2L595VV0EwYz5fjw3ROzU8agpQs/
NgsqU8NtBNiOFqBhkJOCsoIuJ4eJCfbSmL1nsvnLpWYMl8kCoLZdzyIA5dAjbOZH
5kQ3996k/wFfcYNh4CVyNUFsnAE9m1dO0B64xlnMLA4S7Q50XTa+wZhlnr+tIFO6
XUGcCmKB4p5p6IiGi0vMDf2rkrxjM0PDYYINw5eYdAEY06aUMQbM/W0CSQnBpak6
zzYqlQ9AxNG+6KhGEL0GSw9FxriGL5mjacRpA6Q1tW104I9A8RCkCRRaPlMAa48W
wOUIRKj4AZnDO5RnGJlGsw2fZlkcF0Pw9ITgs0hv3VwJrfBt4Vb4Z8y0URTDa9pa
YnXhJIk+aTKddy57ragizYJKpZVRh786IzvnMQSeYiVjshJS+sSPg1TtUOcp3bFv
zBYBXjjj//d76bhZW0bbqfAUzXAZUn3xAXTMwcc7hXEuEfG2ptL6YsN+RK3IRRVG
+jmHjXwW9KoL8fXO1nYHH5wd2vG2wfiFn4er4eYcLzTRzbnMp8ZOlVe4TBUoy37L
Rm6Cb9v5ysEnCkQ8HgTQktlPGsp4RVul8cKONsEXt9WUl7aA+avQIt0OZ9W6UAIt
uB5NRPc8J1g7VXNYmoykIUZvWF+ar5SciymIUj0ZQPTlZKcil+sAap2/K28uu5hy
m6HQpiSNJs1UMKZ2hy1C8LhnrGH6AMjwewZzvLmypYNOuVV4fCZqQaOMmKsHLqxk
k+nyT0U7d9PHqqi1WtXDVBYubq/XDy4lUwIl1K9NTYegvOpaAB2dVaPap8Kl4wv/
W1oPa3a1OSlzlJnHLdzMc/mAbeqZxmoCfXKan4JnnmkdSUaBbhScekvnOcUeBITM
QikNh8/0+3pYII813ykNBGuglpzBHh5lowFPcYOd8HyY95hGTAtmJR2Fj1wHHuQu
9jyXNM5siGKQ8k0MwdH1BrpXzUuQ3XYFUo8iFqoTW1JQ6LHgI5xI/FRcLD8Kh+n0
kL2VN95/2pzou1//scp9XI3NTTq44bkGtKV4jDvMtxP5MoGjbN1Lgv5ddHiz9Rkn
fBiiDZ1By2ok2TFmXFD543FPKyX1JSKFEPvrVYpbLt1X9jZZUWiLNXESTFi0iMvN
XWhbSGuEY4jmaNXGvgklYO3v+kGKvovLjJt7vsDOX1Dckl3qgi0J45ePaHrxPz2J
ujhN4WVZZ/dpPiYp3ObEtN7prOJ8i6r0CEXyAXPoiZJgLq0IrDeMPW3DJ4jt7YwM
ScCfhsCgePz+KqtMGHuW9uufU+QThz1hv48FRcZOgM4j8cqKS5Somu8d9HTW+OmF
VB5ArooV5+qmtLVjHSb8iip9DAHcgdVmUPRzJ+ixBqTyOyMRNta4QUV0P+PI5cQ0
oWLtE16TR4PS5uVLDvvuqsN2wwhq7BUv02P+H4QreS2DN2UnVCt0LeIhh/TDwgWL
R+Hg43cDM5ogxlC5ju4Rud+PKXI36ZGmBLpjP17t93zluET5sPchH7BdkKcP3Kyd
zbf5QsOrTKBa3FqHpzl9tGNCTGN/jXBd89EZO3KeJ4KvG/DpYoWHhJ1d1rOJNObF
OJfBeIVp+5A02gU2q+dAwIsdizfmCj4sHKBPHgBeE8LG09tp9V6bUApI66/SiP5I
VaovUaWFIxSm22XCMPIxvzN6NRgKDlYm0MtB1Nfvbo580NnwcUq1QfPmxmeJSzGD
qP9mVmBgtmWJWkeMZA/dBBFZq8jJStOweXtdNB5CeqjTx3ZiYSXOYWFv+4l7fYcM
oeCT0LmCfOgmoGYqNloT6o0L/nWeLGjcIZ3zv3LoSCfOkokSYZKBRPSaOCAddph+
wgpuwxEV1IabQB/kLHpA09wbRDkjOOT68qOVkjKJQNOtLteFf6+3H7m56vtvOHEo
xHJJWacln1lf91osJYHfSEl0dT+xkPJ+L1/mU38Cub++Fhca3gPXMvJ7j+QB/Yj6
CNuo7jwEA79TNjmf3cSup4kLu2G+4IJBTY3LKz2z0/gB1gIL+rUAuiiDN8YQCuCY
J9GLS52K93G7h0AwzcCqo2R8/DHrQTXCGB3gby9Znml+c4LgJm+VBV4BvsaF4gG+
uj1s7wFMfRM2IwXWy0srRDd+clpzhZgUJSbSUdYWolm3NGtUSXbvLuV2sPx3dK3W
PPflmQ+T2yffYpbOEgDHzAy21DpzJIfkuso41Od5etsYKCWDvNI4ZiWJV3Y/7CGN
oSsYGznwlj+Q2ZFkFJpIVdMVPGsOLsSGG3ckieBa0cuDIxSxZgwBnZQHYj/cZ9Qu
/u56ZrpbztDi2kEE+EUoAMJE0RAc478soYDRW7Oy36/rM8IdLPzdDe/r8DeJFC0r
quJAuLys/r5thKt8U7CjlXomw1U3yJeTlLDbI5i7IRzjxt8Hdz9hGKXXOOY3RBAG
S47bk6vRLjAbbj0oIfEikrEXl3cfBcfkJiDMrE+Q/BStjJk4Hzu7ttQx5EYRlg1b
E3vb9Z/JYQG86SteCe0DIrxkPvyLskpvbFLbq5ssBWTO7fgcXOgiajQ3dpeCV/hC
wqZrClJex5QT2AhPt83RAvMWB3Aq14qofzPPMaRJaOvF2WWBJL2XAlay313VOXX3
ixDdGAxfFUzpSbZYsmVlowrr/QNw1CUE6HSaB6FvaT5jZDWb51mVN0Cg03DJ891F
y+S6J/pkk+1KXN/RvxWvt86O9ieXQDvGqrv3K+iIrmo+Rskxt2F9XVgTEZoO2mwh
a3wtsKpMZdlHrD4IzQV2FAPtmkFscbB1EuNafWkf/FohUypfN6UvMcXf697XThmR
LVkUGO4jwPozNl7ntHFP1ESC0z/Wutr34uG8LgxSiV+575MDFI+r/39lCjZ+7/xs
NqUYorWN6Dwc/ESaTsnBWxAKuZYGhZsiVTJ4R4Dpo22VsJdNhb7PlEksjXVJvxUq
yZVWC4ZThR+5FzhLCQKjqLHKaSGudJK2W9XaSrUKO7Tj1tQKDGIURw5kimfEZKVH
AYIBszlm16Um9leEmkVwwwFEiUQuJr/j0a5/RhCVNirlqGYfT2adLxCObrMwpbTQ
7bksGTOF3o1yQIe3AbEptmBRvyatij7mRw6gjmzJQnwTKf3mYzrwu04PXBLgxZBE
/WSnBscEAmwRQyqvSlx3r8e2+XhWBZ8PAEIlc0Xs0Lnf774Bjnq/0SsN7A09E1wa
U7pQdhwsAEYpDE0Dt0XyXyICJcdbya4fGTbEyIzR9Xg2uXpdIdUTvLCqEK+7F4RS
Dqtl2/q0ZZYaJmf/CjZBNdGXaxLyjBXuT6Eu60163gxj7RZrsz9Ks+G+1mhviN8i
aT3be02qzqvFuS2Qsw5LuUICI/9v2M1kmlD3um0ulqn7z+agDlWEmu2pj0zsnfMr
TQbe4OlIQUQ4OT9Dg9MDMFyV+TGxqet/lNRI7J+Vobww2ARahX2VMF0S7XMwb9US
UXvsIbZVfBpejG4WHv+E45g+HlZAmTpc8CBrat646EzBi4ASumRzJ/pQFytJYHak
UD/b+kZP5Rni3DCepGaSzI8+d3GdXlhxglPeQRpQ0W1ujjcjWvF4BwdYGK9DYhLB
+TLeKGtPPS3fIsyoL7cW5Mf7zOEjMK8zCRsHaVV4yZKHp+QnFqn43xFW0Fxuth2m
Q9YwOPyZWcVLJa0bzVT2GnbVYc2P36+1gieD0JoTW24FW/ghEHZGOrOUeAXQT2hI
InbmPRXZndHzvTBSLG7l/O+yX4BZCPZlYrOdcqg4dz4rhvI6T06z2eau/Stwvo4J
c8HApISatXB2e9nOLjJfliDxHHUpGCqFsDz1nF5lZby7b9j0N4i4YplNAY9GBusN
IiD9Y0W2uX6Gg70WtSdaG1APyS4wCPDkG/c0I7zf+gRnMkqnGKc7Uxf20aYEBLOT
NOr3lEZpdG2CJvy4sfLX2yI+mN5nHqRfl4RuzyYTtURGxW7vDPOzchsG+FrwjUm3
1n6Scvx83kh+Nn2qdw89JyqrBHYWko4TrG7wXLhOk54JdYOS/lFTBmvU2ccUxiOk
72ozTn0Z7lpGFF9yNc9kDaV2h6s9D6m4zH/+Tg0LrsqgO5Tv+iRes4boPEZ+t6+Y
P2NfeVOAeIPXvp5o1/4DHjpKS/22g9MW6Vi0n3L3TX5OJ7phbr/VWIfOMJdS4cRl
8/vh6tkJfISAY1Vr3YZ9T+v8enaVAWpJLylyKJqp43ZUqmWdQOfANVqPq7YqYgDX
2jAqv9UPSW2a39FepmF8uPVL1AKUznJoFgxALrZ26yConFXx5uR6gB/ko5jggmvv
bT/Gt8GIOjJOk7MxPV9CCNlC0JobMyapIK39jhrE7r5nOXFJ1uTg04O/a4/sJDZ8
ciHWJcCmd6/32U+Ut3Xs8ynrljO4PfySfLP8PvyF0xsjkiiGtXmWisQ/Nq0fLX59
nyvWg7HqSShXrq2c1pBGWEU/L3bl/6k28aWEkGCcsQQt8h3R0QErHej3TvF9UA49
ZEcuBKu+hqq+P+D3HaCIvXOr1hZDajixocnRo78Zzf+ildK2vNv/Dym+kfVjU28a
/hzQE2ZkRQ2R4YDyx8BHqBx+3mgQmQf7AXAQWWuS1p7M7d6NX6IIA2dVK10lb7Ll
e/s9nuUQBM1wFHXzDGQWInUAyMQQd3tcPfPAsPSmi7HvRf0kNs52NOO2yMLqlCXn
xQ7CPWnRoCTWhGqn0dPM7K1wKTBk+vlgvryBZYGUocCXJGxm/PO74HODYxD9ITBr
FxVqBPpULSC3GmuIVUt/Yf1VBQoiGljsr0dc9mo+wEyFf97jyO/MgUuP5J31H2Ej
V9RqI+oUCvbxQWzT1GGDKnMIxxGsiY3Mkkjhmrwkum8H41zMspwe9HyQV+WhdqIA
67s2E99PtcIgz5g1yIrze7Kmxup/0pZAJbSgsS7XmXiEDYyzOLn7etiLx3nf4Vur
eSdDfZNcTj3/KT8uDRE2yRsdl6p7//cSc6CoGkpAWaFQamai5s4jscoLSzgTFC9R
/DWFrPgk88O5NuTelJNWDGW8m4cgHDFIdf0XZZ+axpE+nmIWIaRTYaoMIK+g2Xjm
MarLx+NhyvtVHMm+jZNVZUC5Gu8/LBUGreS/KjoZFC0sQQRsl29a92xU5lE9qESn
u6nldwHrpechGJkwdPcVwrMUwE0l+WP3pRbrJo8OTBmhsSLXG8l+qV/Z10pb1o50
zw6exZsuypwl4BbBwzW2rXe/MgngNmTvXmzlPjDvslLdID3xC5Uy3aI5OyvdujSN
mnsuC1UK3rTHcPaxcxahATx3UX9X8ajtHBHFWGxNMo7l4yE2sCJCL05ibKL3kNs2
MUMNIayZs3nBtKXmvzb33C3PCiI/+ZqV364Lnm/9ezSuPb06SDgC6qxWhteSvTe/
1Amb3Zza2C8MWwPNk4gVVyt/MqfJHRmKZWOS3OwREZdj7roJCfp2qO29LSOKCpV9
+pb4KAaowBqZ9ZnAEM2kZZDs1uAgVCR/ebJQWWYS9lpMqF9HGr3bghYXQQ6YAZ3Y
mOvQLcdWXjoA3vIcF5C6mYLjQ754Vtv4f9kJs558PiHyRHAMES2TTojtb8TFs8p2
woJZ6BzG+i+QpjCbcnOgxHufSseTSgYNmfED2v12tIUkadYM8svItKdsR9nll0BZ
0bIoTSPBc8eVkwG49nvKab3Y5LY7jmllLp9I+2raD91aY6J9tnP70Af2PfbPeQHH
dJsbawXm3YQFF/WjzsE1JLh0sjb2lUVBpXH7uG+GOZfCOkbWnNyRMftk9utKUWJe
gpR8BnsKCn2dcn+XEKLXVhymo+aa+nTX5/jWvAOvo22NIDkgI7R66JDLbMK20851
kjff26cXB6vMI0KwKL0x7HGQ+NF6kFxtvGnP+/zRYksK29DzvaXmRI8Iy8bCpR4O
mXprNAmDgI/cKpqio5GSWmwI2py47/gGgQ3KI7eAfLdJ78crYL70TvHf8385DZFI
3MRJzi6iDe8/YLvbJ/kpqAYQkKuD/y+N8i+/eI9lrPPa3C8qbAyRaxfzoL5Omhea
luHGzjLt7ezmbkAuR8VMBgeyBxtrwoEwzHEodYqOzhh7GqjFS9G/6x1DxFchFzub
brBotBXgEMLwvprEKOrxSvkEdoVW5rYtIQyINKHUTaY6rX3REeuAAmkSYCjky2zr
Pw0Erc6mkIoD3O4vZ6NDlZVM1Gfq5VlscDoYeita+Nnfbfu474RiI03i/+vSKr6X
P00wWthRZyB+r9yGVr3XQvU7OYb18ll3yiIfmbQKrQ/sD0Tpp1fvS4zw2i7P+qJ8
1/qd0KxX7f/JyctQrwgc1Fj2UNnbzqnhGyjv4N9xt3zy2rE70jwR/jo9XDJ4F/9l
stuicQjCLSlgqCpGd/UNeTq0Z3RhU3aKPdr6RIg02KakxblO8H2qqadYoFiBfZYm
MSDV3uWD5marPOQTFNtXU7pB5VTwFcPFdb/gu0GD2OsThB5hosu5xxruIPfYNfwj
7L9TaC3xNxYhF7ffwo0WSn7zYAng19m8AOn56kZK29DkpFV+3ZGes5VgyjjKZoa7
VnNdcAIAKymV/pLdbeQfBTEUkg5pxH55CHBSiC8vJVw29yRZRCLgEbZm5X9yDm26
x9FuuEwM07E6l8KNLnRLg9KUDCCmfwYs82q1IOZYstpP+ar0XixnpSjIn8PIRv6R
s6QVFeNSvP3T78BreeYpxPajSM5y9AU/YYC8vYJNaz3YyLe4Q3p0YDnk2JIhaPre
+ncJdcuofOcYAURxBtJ85d7ALeQYLLiMbYStot3JNWA6nwRGMplaocW5Yv4noYUG
paPdEBYC5SF4kh0Lvck7NRV0fvXFB/AmfakR/gKkHk47WP94XCxIfMqvjwMYxqSQ
Eb0bhlNqC/lKUJBcr1dYZCC8aqL91b6ZtCr8uPCu0qOCqy5F1LLkGE7CBx8j0LFJ
u1xBEjBULeC9r+mbgzA8L20k3VEorkJu34D99vzvUlZRmY4zj63kO5hle20h/HHx
Dm6TEoQx+Ciavo4eF3WQWD4Bsl9KrVkLk2TdFHcHR4kRqZ4WDhvzXlZ1qPq5hWka
PWUc8QBYdpUOfQfdheuzkaTTwPJkCzOMG1X3pRDhehr65ldzG3owjv2oLAqndjd/
H3QG3CLfj5aYLeN6kP6ZLwRwW78HEgjYlQfnJ+ZjFBVjChuyXFLBfixkHMZxeHLz
8tM/TFwezXQmaYlUDBD0tyUjVSxdASTsa7WTgWGLPaiM0Vy8dxt/wEpp+Os6vhhe
5sLf/fLCM+6axlUb+O/AdhdmHPsElEUKEaogJJBNDF5pxAwkZPUaSzNcNzewbQCv
n8b1toV3gp8sU13OUk0qwcIYOEVS4POV2R7UEz4Q0jWhIh8C+xe9wtmoIKI2TNKm
BpI0obORf5q/nMwessppeC3t9YB73QN1/vyvruV7n7kZxESkaTZKJ8WJ33jeyJgh
BLAe8SjCVWVXrN9vNkcbx2KYgFxfbcFLhmmBflOuKzxHEnG6LnQudjaUeSw2hqN1
fMNeXLC1n7k+aj/gJOgMbYebLkB6othSuKeyFLyi4CzAR/1k2Db2Djx/B/tI70Lv
+EEHaJ9DLi76JtZbRmdqrENgPQ7B4S/pUhs1Ds/FyMiuS1EAUW13zIhROJIKIRZZ
DuWUitBJBgPgTXa7j9YFHb51YOqZX4FiY7t6oAfuWQPatRSV2kt5ooc0We2PJbVs
01tQXGFx8gCMQFyCF14juyIH8p6XznMAPBI7/gCXkxGx1glaksdXN/n1oHbdaZKA
weRXV0x6UvbdfanUjZMAn+6RbU06xEcqzpu+mUZjtfu+BorfOOuh1JoyqGMedTxR
rO3ToF4aObgJruWIALD9EqzCAevAFSuyEh2T1qW3rkMwLatmRalFMHI/2Rn72l+E
BpiKmTx29vRoUajBouLfw9Y6sWDelP1K2WLF+29RTP2ZubzON0CvipV28DsRh2+f
1VlfpKWGqJ1Id5KfzwNEykNUWf2CnwrQ0901SsmDTBAU7L2CZ1NtirE4ByKiTLlu
rj8wylgGc/0AoA76nbNXpbAy2gzmIDOTnfh01a3pY8HFrJ3k0/gn+YdzfOl8yF7B
GRmGu13U/w5peNhp6tExAfMXUbOglLFs/JiBOh5Z44As/hF4FtDXWfMVyUmNGkyH
cTzEaqWw8XgVB5qO1HhQO+36WlVJBfm68+fh1iVQoY9NOjYOso8qhFihxF0ZNKRJ
mPNZPfRpZ2K49zu7HSxPRZkFsi/ZgMxwHlZhtjAzNSSDuLzp4C0lm14dZN+tYItk
NGoY1vfiLnq8c35Wjw67a+eoyCPDK8a/4YBqYsbAIRMlxo6KwmVUdXVwNVSi6rIt
zMWZA7GWGIXRfWntIo31pd+LJuzI4MBspRjV+fymOPyfcj9Fjrp7aXo8SsZMrWB/
XDJCpQ1ZSaGS+I5zP+QeGUzcyBAEmgzkbgk2kj1ELD+bBP6MXzl/Mc98xUU6warE
tQDWLVQ9m8dSsst627te7Fyr8H2yeQttwlWYKiCBEN9DzAqkSIhHMLs2mg1N0Pwh
nCLLXn8MnXktlPVZybWJnNLbauxZKFQR6rORG6tno+pfNmOrlifvQTyRHVh5Jv9q
k4p+XLNQwXtECVZ6Je2YYPweKN+vgZNmZRkq6FUPhSxlEjH1f7uDC7hie7SRgdHJ
OE/P3fKQVOpjVd2UF3q1GwKbuk5laUPaqC9VzTw1Vl0XG0S76U9HfKbUR8QXzzbP
/JgIoUZ98E0/ssDW4ApeZ/puYTKVN73z6AgtcE/8YBWlZTGA1jfLCeJJ7cQoQtsI
srjO2hng09gmti3Ipp6XuQ6cdzC772QvcLxIk9sj8ijxr4w1zVV7KY5zKFCKpj4H
BZkCh4phqo9iDDQm193ujomGWfTa79BiGTtDS193RYQxy799vfqOyALdWoYpeaVR
idQDEB2ucZd2cjscskh5K9VybUcX7xwrfOGWoHBs2EbIeQMB77Uo4HXB162xXX/d
SHpHLV1Bict5kOgULE4eu36YbBXy7x7vmDBA64cTsrlwbjl6lrSxh3/bbkTsbSz8
Ff8DkJIz9f4u28leoofrOQ87JPxKddSpZLKZCuLQOT35bF5/2tvRi4NlFIhHgytG
ERGHcIkULfUFQMxJ78DfBcKqZM1L8kzUn0qaYAFuJJAGL8k5f5smV/0t8S9btGRc
HVfDkvFtvF8iG9zXgRA/RT7dwaLe0Qbm1BAVGD5ZS7C8sqAuqgq+278rJBOON/0L
ldEEiE62lb3LSTrCLoCNPb1gsA/EeyvLuNXBoVXMtLhvxHYKpMaedBAXSK0sqW9t
LmGU+uvpW9zse10MNDjjYltMKBiqNLh+Hr0vhiI7bUC37sD0tEXw1G4g2UH8MqXn
ZDo9/xCf6ghswuix+BlapQEHhqtkjIyOvVf4vfDhiIuVaTg1cU6LDONKL315uTQ0
T4zd/b42AIRjRTrDbNgtOTpnGcne8xnousYi+lmUkwOamhyZXiOv5adA24/HmJVp
r+u2XE3qKGZi4BgL/y+Obi3GylhRhSOoMSoMS9Mu6ww8XeW5t/dSzK4ZEZiY1GU2
p+VDiRZiN1WXNW/tu2S6+6uQV/jg5+z4P5Va8/zs6CgHwBnzabmZpsGClu3pK/Q6
Eka6ikBZCrvvaggkt7/kcwmcF4mkfri14IkKiH8RRcAvX7oB8JofDegTxhedAS77
/IPCAuwegKS8SgDDusT/6bmMXuKV3oYS7e+WyWYIu1ShviRKfcBAG7ZPokefw0gF
hKwmL3hA0UlQoeONND8arUeQT1iHYRbTxuLiD6Kwkq/DQ2eh3rr5zhZnYAeB5/kj
kmusa2hwD7a51VJuAa9N6tputoZoXOdycl+ytjlCsNbuTMAYFWfJt4jiP069Cm7e
b3gC+P0HuhtUL8yJAMaeg2TkYjoWp63dLgIzf4xkYxd6hzoC2rIxb/X5LnTG/fAH
PtmRgwf0hrFoZwjaa85Eqnq/V8GQHIgL6C8HhN5ipamdV0xM4FBX8mllqvwKo3sX
zy6MrYzHBFRVrA12FZrDLhxCg40mfMtajcQGViWdN0cEMPbUW1762eBomETaAdKK
d5v8FUHDB3X70MPGUx4ou/P9LAwORXd3Mda95YF0PRGytZ+MY/ZqlMpMptiCCU2q
ZkEn64yAf1J4iG0YPcPu8QJUDLlvwutb+ySnXZUlsksD9XlfVtol/q2G44/qJS5t
qHvGFu3XbFal1CCKHgY6Cj9oxujBrQzmuO1bfScdx5RvqWrwo1onDyQWbJLN1N4y
UbpnTIYuPEDu/R1gIS7w9a+oXtNtf3nWX493OtFdVUAG9ggoaylXlPiVjT4DJuuz
b4YCZR31piGdI29/5qa/AAaRmdTwYubu+T5s/7QFTK9ei2aYrG0zWmVpmx3a5P0d
w0BXgRAw4ly2SZG09nLuZPPQ1FUsLjtn5AkFTQJu49XB6OLTLm1Y58rmC0Avh+Ze
Y1BylOazhxbe5uoCqzFhvtC7GZSxoDiJ+Qvt+a6cyNzaCVIGCOrfXY2NZ23g2mwO
u+4UxLLV81rYvGX6XF+USWlBZvLbWLpyc9b9KfJ8xmGdApjUrlotIaLke2NP5CsJ
9ThmlR7L6s/58wvejQ0mSfQqOvbHirHJLoWmAXYKToREU/ejDVdGdx6Nt+HDhpn1
UK9e95xH7hle5btP1izUfrT9L+aByY6L203J8SXSCx07iPT8FlanvzbkfO+CP/Dl
KTUkGuDVwN1NvyAk21Kv0ptcaC2v2tIKtB9Z56Rf/tsGOvCIWlMHh0iAv/nSBZKg
APU/PArxjJLznAf7+Cd2OVDOv/eGvmQDQz4La6RjsxgDSeuoN0Ms6xkUz6k+2e1W
Ix9cTt1STvrvYmOGPQiapEdRlxJzfPOOI2llqABHfBWCJkSIrj36F6wBD6QN/b9H
/p72T2f9uVKomH/1foctL0tpMPnnR/G1yzQYhpTAZZ08jG0M1rYH7Rly6EgHdU5L
NMvwizKngcmCVP/k1IOUICztrwxj7Cg2ETwBScD56Qz3Kx7+n9YgoYa+cXOeTWfy
d3n3+4QbhNSvLvVWtA6hiOkA/Av6iAiVQ0Yl3PagEkh7+G7Ma1TLaE0uXjvKrdNp
/1Qx7xMx7badI76AANEYBlQDDiEGJ3f720g2ZEk2sEVtY0wzeLE9dKzupLJooiGr
EV9fJbqL4QThY6xHBh9qBXmjRvQ9hLvxfTy0GjB7Fab433VWQgM+45Tn9qbitEfx
HHpu/uHEtZPocYPtRfAK9YfX/pD/zFgfhyJe3IDGW+aiM9vkXvl7oxasy7Zjqlh4
NIV7DA+Y0XOPXzKYG9n5IJp/tVlB5kzNYQ6RkligzF5BvPUkkPvvOSZz4061iIEV
F2zbOQUvFYgqcJr9eSlS+s10eT1GBVgVLZFWzkBWRXGCo4aIPYz8iDeYQ7ZtIoDE
Z2etr9Svm4PH+nTEiyvxlo9gPzWtx9DC7VUiLeoFZHngXKYVXsmY9zgBw7WKXq9C
wu0q9gIn3iaxed54yTFkyU7+wwBio6nXogiH8tzF2tZ6U37dcE+lOVtjBqbsVxyE
FikysZx7/ikns5soRDY9Aie9CSH5wYeyxgwbKKjnSQwfN1hFIvkLcbt0XU0eFiVj
jAbDoqobmOhGCF57RvR+TTfJGkXbNDNT7C7KrdPeNk0TWR6XNNIf40BDluL6SIFX
opnzsFzbK47joy3Aq5KRQUFlrWLpxdT2eMn5Td3mt1uz+qyPs1d/7xC0dbVaiNgv
PPXpd63Epw5lvg/k39laPjLKnz7zCcBPxWfgHDrjdLnFcsBMbtUbUj00Kmwp4X7J
u2QFvcInRhXvGF9FSKYcVRMjgxvWtRRI6V7RBHMwjRwBc03yGUtd6s2rvYUAbZVc
1EhxaGDKJPE25T2xcjSXJ/nNPVlrv9IPYIu9qGHL/+v7+U5D3O93cbeHh+4iNsI4
P4FE0I/oyNNwE7lMPDRjl50V/mTRcDDMnmGFii9Aazs9d/eBkuiOa00vU8Tc8p4N
m//IjxG2RwTbJofcSOARgrI8IJSlZ7EvsjTccqJiZuSHIcB9Zf/KazeywVCdnaWa
I4A/ppUmnnHEKYbDDboRVu7s8nz/WZAblETxy6VgP/Gg2FITzTmcChfIx3+krjpp
70WR1uNkEG4BplfmUX+xfOToPXXIA5hPwUw5OUq+7UTAvi290txF4h6yxta1A+PO
L0fk2dBlFxyGYt+xR8EMKdsXa5B/wU8lBO2C61xN+iUQ5uNbbU0UR+/vApUsFAd5
cArNWAfq8Xzl4o5dSK4dVcnnLwLNZYCTnlGPlYZHk4W1U98ITWf2qOZQGFlGtVFQ
dU0Vz12DgNAuzTxDdLsGSvF8B152tg6gtravN5FH5kH72dipCUMguJDi5pbAeV6U
N2JIJvMq23JenlZQ10NoMM7Yj7aZU/ksNkmLl61QnzJ82P1MOorHSqYxcsblCcDZ
yhNXGcZqZBfgpob/Kx6zDVAgzJu/8n4mUMrpbHmI/9XvLhI+N6a6h9RG5/rZWei0
V5dhYokKnc9flDMrAtIRBTFeYEhf/7k70Z5pXZakkdplvUw408gLmvB2AP3jhIIL
laADpUwVor+t7TPOteoJ5zgVhSLpxaT6Nfn1WRiFpy8bXgOwSTMuHycwFwq/LQCL
3fTz4yHlnAz8fjgiwJzGBOpo0UrCI7SEG21iFaegnR1d8cYS+aByfIpHIEplJzNn
iOn55a6SMXtPCNlxr7pTOk3UWyyXqwUUeNjdJbfbUmNawyh9DN8JSoijE3DjWM9N
ZBq2L3iRGc/K0AGFhT6qv30zbx28SyV02hcPKZ66dt8hO1v1Ci+bwRee3VYJ6CMk
MWnpTsqMr38GBoMEm03xLG4hxoW5n9L8tVcqeME38rDv46pTExA7QaJ4ddaH/Ov0
HTZWBDQEwgRSjqYz3mobkcxhQzF027h4wSrzq0Xf2seA0ID6q3vIztU0ztJ2rVmp
rNQvi8bdWRnV3Uz+CIXg4kLfaGwh2jqdGzNFnvfhMCBSPIZxQWw37mWT3BEhVr0k
GLGBw8ohZ2rbA79zDmjMMLwtHw6pQIvrQhE5A9/CHM1vggOri/7WPB6rxlcElW2P
huwt685W7As+Vmhy9Oq1TI+Ra1FQ64FGJ6QM3r3VDFF7vC82El4VagNFUMcJUfys
CwOg4fJM5ZxPI3NuCwk9T3+VttW2nwssLMOjeyvibKCbmhhyUESJxIPIpv5C45/f
FbpJi9EtBpJ+SrwSEkE7nj/iKfej3Eq9xeg3sB0xEBLkugM65cBBfc1P2ZfLSzhS
ABjGBJAj684B6hkqAE15NyeE0EPTo9Imn0lwcf0GQt9wTqpIzvZF5j8LGqlE7NxK
yJjaIi+0ONo5JpssGK0O2/Dbm4zxEHCdPPoP6l3zkhyles0Ox9OnVLV4DGYpksQC
iCCBuKyaeRKYaiuurSKGFs1UEuCbkiN+ajeHhGrWITMn6JBff31dzBlzr/rhn4Xu
gQrXKG8HaUxf55P67N/CtvGpKIzpL4BtEJg3KANJLuk+r7EJUgDytuWv/+wGbt/T
AMFjp8CFbDp35RmXF0w94VnuROzf/PBwRCGXvC1UPQlxpzxDDe1hhA3wvelRaIhl
cQQ3a2S+Gy7rdTslCfS8XbrjgNclZ3JPE41VrLHSEB9VRAOI77FwBNolS9R7g6sh
cbH4XdvhsHQz1XnHRbTYWz83I76UjXt+ORw0QewUdaILEWvYWoPpRlP3979badYb
uNFr0/OlFmYRk92AV5wy00AltTcOF34xZqklkgFEpSogL+dyyNcsBqGi2pIivQ24
+zKWkCNegzshFdjKDzIGRCswgnIOuKmk+S3IplDKbq7uO6oCoOVCejwVWDO0TRKW
LFd8yvVoUOpEckTodJ16p1lsnDDsVee0tZYqM+rfqUIcNgacByWEeLMhqs701hNV
sjVNrWiq4T1gwo00Q+M5+TuhnY8rOvHx3tiqggQ57IwWSqdmoEjipA7Y8hY7kb7W
iKxjMGmXcV0OOGCGDB4QS8RfwKBfRIr5hu8Q3h4GBGrfDv17jW2StuFhbIWU3jPz
7hlTOnjeA2MiFWwLDJ2A4o0KAVSO6xqsl6jG7aE1ewjDDK146V5ddckgAR2zUlTa
GbjZb0uuJDEDdH/JxRifHmEytADYJD4IE+NhofDTY9kniJtuje/my6nR2CSYXbHr
vjnxF4ENM+u4U2Ds05eV8MCOD8Pg2Ctp38dsn0aNwGuxnIY8pOTzobUSChJI8exH
t3iHHAIZq4GmDCqrB3ktEgkshHDsm2OhbO8n+yODfNWziPgkvIN5b7HelArMST6K
huIVnVXoDtS0cld9VrgYe4mkFO8vS8s77AjokhR1iKHfu7Bd8++jHL3XA8GIZ05G
zf05Yoo99JqxuD9A5rLEAZ8TgDQoEaE0p7YsvdHuOnAoDU2Aw/99EeoJkzI84BKU
2yqef47PExFALyHUqJZwOUv/q39cKITYuXVBtYOWxO8krBTlsaqglRkC149YXvJO
t/7RKHauYkkxkAVnsn0+eiPJJam5YrI42OizbIcRYS2d83OQEdNXSSYrK6sq43qv
PdvPkRJdyu8dCdNvuUD7DihTSXFtc4reRFZUZd/OILeR74sVposm4x5o1iTAqXPL
c8FFfyctWNfj3ZCj7leadOU3CP8v7Q+lMcckBoqNQjuMIu8Dwpt0z6HH6Xh+ZiZm
+7atG/63T6RXo189r9WhIASctX6EOzCnxDSdtPdio8hWG/BcSoZxqpnHiXnBxLbg
Nq/Z8dn0WoD/5KqFsCxF6lCVln05fAdaZDtqJZV9b0hgk4Wn1nMQYMHxYSJcOw8B
HHpGzKzmeZjiWT93QHQgyRd6s8H5VaipqkFDHsKbfkwFs3X9s0UAt+/bByYJm+1U
Tq8g7wqIxfrj3LQXeO1sfYSoxsctCdqPMoNZrt6iMuzCEpcANKHMgoEI60GzQ9pr
tzdHo5Fsipn+b7HsQXdgyH0IzCLYezT42KzXOXbTfumzOlxj2ABGfaWdBkOwnQGn
SM1RkAliFFTdKOWDQq+HPtKGbZ1P+NG6wqBV7MBGlteyztJyzHADpRwD3mupiUc+
I8aqXTpMveelAXtBFq5jYfhOXBRgqnZxe6q2oOQuzBGgYOmZqzQmMbbavB4lD8Pw
9PXlMoSRJ0u38KsNSqGZdBaxHccXRcffLhAmjanArsPuycnEjnHwqUXtlUTwGKs4
komv4nanro3fSyd922tgEYGuSettZqDxVaZWsBnvVCqCnCR4GPZFmXlLeHuY0Z/9
4pl4f0EtUF7lXXszhPZZRc7+yi+7DOyplv94YtzspjJTWhlOOisyi/lN77ppmCm+
VUVN3O8c4KD7kE5O88+0EaUxRGzGKluGOxoeRgg5+rznHTMEuyvYmGetBnQ5b3NR
pfAz7BcZ/h81w9ovh9Q7akRBrWNztwZ6SJiiG9l9Tn4mZlNEGv2miXWJf+FBAizm
+mqs/BZEQCqPS+7VLGMjGIUs56n7XQsEYLSPRUYS5wjrptJUvfnOiSQ0vLjP0WJP
tvsmIeAKUgvAE5+n+Li3rTGSRck5v5+bjl60a7mhOAweltdy03Frv5I6/OXnmnal
qo53EeI4hGyj3oagjaIpr9to8ax1BU6AnDb+SPKMxb4/Dxc5j6qNI6UH31DA+Z49
1npEHvCSy4UbrWKBMsQw2FQg50SXAzccQ4S/tD/geoIhWmbkzxs449IEm16VMkGv
ZP9QGuHpPlPErxtLK5hrpN3gkghsjYPNDn6tlk8e/34Wko+k8Z14xxpM0R6XkI7A
EJ1EPc/41XURRR7b9CCoCRC/OGaIhdQEij3v6fBI7uZXuNXki0GNJW5ZHWWFORIs
w87QKhVL66qgXQy0s5G2dJkgINkYNF3mNsyL1df+/wds5Q/Vsn9X0e9H6o8OwA0N
XBj1DY0pbyQzXvAH1ddJzgbCXelLYoxdPz4oCQHygfSHIwAZnV75ZXpig5vODYJg
8mpxO3M1gfBV0lRzNu5jot5k6FzIa/PBGY8EFOAKZ03Sm1y0Q/qho5fpshalKo0/
BLLrQ7r4Y8eZL9rdwJkuZ+cSgon6qdjMPPh0XFmTFQsS6PhXUcO/TNezBx8pI7uE
XfQF0i9tIfFZ9ZR84c9u5cMih8HPjmrNIVow428RlDd3YA43wHhJ/ZXnidx5bzyg
2e6dInHB+ktc5OElZ223U1aU6VOpTv5zC1xc41GhwQ8O024qUe6ZcnS6kCPSWVms
kZw1uMuKQ48nzT1ChiLmXuwjrf5YOQ2a1XmAY9/nIIb8a5SNMs93VgMC3b+aUJlp
uco2fGaLwOFF/s+CUrkst+WObsucNOcAsHaV1J8FDn/f6jx9E7hYkCl6WxrnSnY/
LLDRmU2pw6WMR5SwAlOrNXKwedr+yTiDNXPcDTIowBaUhc16etZJ1trxMUuGSzcC
zoJdQ7W/EAV+0Kn5ACswl7qErh8bwfCxyswTcDffZLWq6cPRuPFtFj5qmz1+7z6/
L23ZrRlVIzdlp5Z6y7yZDyXUuOvJDQG0e1dq/+SYonrAJH24nYzC3bP/3BXq8QOM
dNqCYbcwyi9ipYgnDbhsWVwWIbqAI36BK+mAuHPfit1OjCzEpN898i/1fp1jm2he
WEEYpaUxMN68a+izs9wQVvJnToFZwUXqsc4/DmD7iBD5CuT8ap9cfLfe4r5IWYzW
rxcOXcelO63zMrY4Flxx5RoYuIOiWuIzyl3TlYfOMxIK8rji/86Zq3gzirh1Khe5
qZ6Y6XMu7+xaqbjOk6AXeWJXNtjgHi9MBaFYRNvuJTAjso3hTb9WqCY+QSaZ7yYw
VgvTw+jdUbBq8UDrKCUZS/XKgvmNNNn02pQUPRFeyBrZcOE7xVqeYG4nAO9QtBNX
vE2JBKe9/1p2Mi7txbX9xKFBBJue9gXSQnAW843sx7nb4xUXsG58sYy2nqiU2lfU
p8RdE3fRIWzfo1MrfBWBxj4FjnZerOiNMz2inmQJlrIGSE2AOBkwSZVtkSj66Z5G
qUcxuRSj5P03SkeujXcRRGkWOhKlhfpPYbKvsmnsVsRWwvi47pa4YCEFs29gMIuI
zbFuiOgPnkFqanaH1N3OuGAOsqxBdTEQLSvX3T95p14vcf2xwdwzGPYUp7+Bb6Wr
sVfH/K/mZrxduU9C7CtstNi5xASC1c7pNi1ySxpqA7J0H0R+KecmG/wcCbNdNsLV
A/7bB17XZoCbmkkopa1smbmdUEabcdoN+ic3VMHt5uzu1DTpg0Pr8qyta8etrFgt
l+Nbk5SA49ozoakKPHTphgImRBa7zubDzU7XtD7OEcgH2MAqhvkQI/0rZtjW6Sak
CZZ5iBGE/BzRJDcVW5oujKuE0uJ147sqTclBY4d5Dtj3BVMXy0GetKjKd9gCL9p3
kGzuFrrMo6iE6ds81x4Rehb+fbcZ3/n5x5OOdb2Ht/NVzdVDrwI0KeFzsfDzDa0V
Vn4Wdx+roXtleVw52sOuMX8a38rY2+R9dYlT5UDSrB14YtGQT1djZi1q38wUxnZI
0tMSfA9/U2mtOaSwhvTxGNJMPeAFVq9kDKg/q+ZVJ2Kj5B8+NtDuCuGIPqePmYMY
wa/0lSs2uxuswAvlIfeYVPfSsaCyG3iZBCItzVEO2j/AV5snYQzf5wfZqTrlW3r2
3iy9Qk1N3YNkJ2b00u9Wf7Sn2i+x31pGABG64VruK6m3idYqUMLa6kg/C+xNUUYR
U38GFn5lSmChEGSBEVPLZkAGOjpbsoEVFf1dXIfscbnN0pdx3QTCjSMzp6VnH8z8
GVNERy0gbNyDbU3ubxpARQxx5zdGB6BFxDNc5UJAwfgXAUhPTtcvOuT7HkDc5kbr
NwVjusr5L8iuE9lWMWaWXh4I7Gi7mbvmBisVxybvgsmEuGgDBp3YI0238aOW7Xfn
EEeo6rmtLCTpoyW2GawIu/EQpLzmKqYdjniDBlq6MjKhgH5+uWRoK/f9D43uO+0F
o+fraURAyy3Wz9W2ZYkmc372x3PzEDB0uwOh4FvgtpQPdLv3n+2AmxiMJyJcAZ0I
8JC9Z1JOUkNra3yylEMNzypMvdIfw4Lvjww5HCCMxENumuJegVZmh8o7ZM4kKX1s
hIpUY22raX25kOmbpfI/LOhM8y2vzjcb/VZf5XpKCJ2rj/c3h8ZRIEVZ0Qh9rqxM
xRAu93dEW+7XfRO5F4mz4yZLBkw9LPhEV6CBYrviMXnO4fZf1TfzISQYVEJFWSst
tNm7GUu+DaimGhWQouAp60REo6dAYGYZzyQCnHVJCubWIJdKEquSE6/XKSYJmIBg
ftG2WcBwz8LBLqlpCpjoUTmzWMdrjZ/5GvVN9i24BC+ISD4T7RrwlysmlP4iU3dF
Q1sEJA6V+TX0iOM4OYBq3UqDcdTLA3HL7ioi8ILOjq0KLHSzZ0gmCsG8HTNf7E49
kJOvPBBtO9bKb2WvRL6U7gEEQKHBoEq/BGgS6VFgTkRKpEaW+1N490ruIm8AXFaN
aVtCAkdnU5JtxEv5As+y/npXuMicNtMshe0Ha/ba6vs5V2+sYPa+VilbyQbOPFac
nr60xyH0Avlroah9Qf+sBo7IEElxCBz81lJPdeHUQiVTbwn1f3SO6BtcFLGoxDnS
QzE9wC5qa1RrNVFLEqH54f4ZCV4+rWFCnLt/XeIQujRUOfyel6MquhyD8KKqLxCX
KCoD6ktItJGz8Y+ecPRRjjgFRmF+6dmS0QkMisryYX3M1/ylS8MVDYpq0Myha7jA
ogcJjpzD8Mkc4d28JIq4iW28cN8J3Loc5o1sJK//7FC7IGH+57XBJB7aNb8ykESw
pZZy/dCKEy2K4Xuyju7x4jqWmRBVyn7UIjTCQuZYWiiSWx8LfBjLpoSyCP2Ihpdd
L/+FPT2+Qgnmakx/VS5EEwHzcLhVZ934VxcY/6XzcURiZ3xqy9SUtHi1EFMjvhvz
vQRP1R6Rc3DVrvkKX/n5RKqMvOlQqQl90hFkziBOyPLfRzNC/QrW9Bn3xn5uKa5V
pc92nC84JAyID269Q4XxbEDNOHuDEhGwqE7Aa6Mp/N5QUnisUAqSr5EQ3DclQtr9
fBhrVL69c96zNCeZU/hZQKpB9R2JAkOWdT6b7JS1+3gXdA3aZzG2glcx8m7hgU8k
aafOsilVixGqVWTQ2wmbA+CyhBSGfVZ9dz3i3T0KyMr9WwNf5bYwvDIonWZJTUo8
8LsFhaZmMtrt22vroHUnZHqQLq8QeEs+xedTfbMElrMUGkyIIsCr3+MfVAWVBiK+
FhZOlW8FNfbOtTtcULn0+YDKbjzE7+WvUVpbcfRe2Q0Ce47KLmmbgWcf/wknqefw
1fwgCLJHCTt1UcPXdVbeHMCfZwfUFbcDqrPSzFQMPsDEAlqMz6Wj88TJcUUYiiOj
gluSX1811B3CxlJuWBfu7Y4xcKp1nmMs9fhe+/ftxYVorcTTtlReeklIQwtyaAQT
EnTWEP5a003erS7PSB18TpPMtGxkBI5CBoOItMjcbRijkl4kpqaxpU1cVexFdhl2
YWG+cU1UL+wn9OOfJE5RSgnD3HWaWurWD+Aa/2LZGFBS1H1qCwD51CuuTbwcfb2d
1GCTjy3Ndttth2Ow+5uz6b5/fH607covZO+G84XNOsH6UnpVFPs815B3cp/3eHzp
VHjjVARN1eTdp4iFxC+D4/06pSAcpS97yguSIc/vNQNMrL8QKGAaOYP60LmrEqUw
3d7LTXHexU4Un58aZMdk2MIVGOVgQI3yv4yzVs8g4Op7dT/EGBO2WYEZ7semOHls
siIpkziPyzOZyg9DkuyPVjgcokufvnaE98lOzsVY1xf0WaDFvUudqaeuSUfMD1AM
Z4W2zqTpJOMvpYFKmDNGISnwUAw369VmXme39pTaZtwit6rkQ0todjSwUtoSZlOZ
Z2EDopgJm6e3707jE2HiAfOFCjIcrCO+tOkpTJbLVY5rwGx3o5Wsye0SdBLWkdpY
8dKHNY4lD1gjIS0O56MDLIRhiq27Dl6Q8ZKM6rqq4fK2XlQifLpBmwv1FVndiPda
ERC+xxRL1GY/ovv1jkuaBM89D38vEhZNNOHMO8DUhYkWt10dXROjxFv2DhScq8JV
3+tY+qZ/XhG4CfYXsCQWYk5qBWEWIM1TT9Vcf8yO29I92RzfnNHU4jp4i7leOo3v
ULR6iB4qaTW+M9YaplAFaDR71sSaphpIxnYEq0s37EdXVcwKarVHg4IVa+qakO2C
ozBJ//aKftrYClfqkR87Njv/F5futNV+64cyVqLU+8gXlLwJchP3hqXtStkcC6pJ
nqQfnYusmqTvvwhHuF45Cy0H+dVVCjhtpVIMyH6AVmtLg2aANdleMwUO0bn+/dbw
DsX0WblMFtFgggh5NZY09np95djvO9ThzGSJwv+b0tt0voIc8HM+znBseniKgKrL
gtpSNOWDjO/RcLKW/oj/eJbPk3mdA0ChsnjdmREwCdJmoR39wUVqL45Ti8QsTrqh
rqqOhk6QP6HBVNU4XnVyOeGMP+IoHPh/OFZpXhV1rPmXzcvDuHent3dF7P5ZEXuH
3swPCdi+mN1cA4tiOhYh5XHYHMeRTS7vzFW7KaZKsJkehzvIcxbookGUwTbi2E8J
u9NgADJe+lFQv1J/M5Ip0NA/UGTyVWp9+ra18m8voGJInyQsBJnQ+UFU5tlZ4Gkm
U3yzTOaKGBewlAjre1iIyfSmKfRoDfaj70/ESX/Wb8rRyuqIcuwOS2NJyDz/KxVI
i1OZyP7VokowTcfZaMhocJ0zpM5MyShZ17kah9kRcnFgZXIuuPF2dkJvbBKg30hU
rN2mYkljWCndAA0ZhyyEvTxFMUqL9vjLUAwmz50XLdzjvSWqabrZL2KBB4+8o7pc
e0pDMkSOxjEX1RE05cWkqkIWyEN4yDYJwBAHgUHgPV9e0sdujYpt6DzuWfuo+RCS
GHZpvE7MSfS3nfh458cRpCcuTeHfNoPm0jtcvFI6jY4ue+OC6Ycbn0XUjb6nTU78
mU9MmwoQB2r0v6PFmazLh75lUn5yQ7fotKKbyCcVzVzkwT+dTXsdz7CEJvEH+Qw1
j1C94jCCTHKeY8d4s/ZDnxSL6aTg+1iFcEi2yzAy3h7DcI4NbuBV70kMnXTeFosZ
njL64qdLxrb29kTmggT+i5jhpY7OqkxJo5XYQsZTJrVvh1EY0CvCfOPz2PBnkDxH
Sw4xN8YFWujrQKk6m0i/d7ihB5UUxhR/ihh05K1kAnjWiFh3rY3D6oziuuQSwv+p
IFpiJ+OnF92k9hBGAOBVbCrn6cK5tJEWvQGL82XZ2NEpvZ5l1guy4HmP9WB8+Bxr
BU/x3n407/THrsyX6Gus9wRH5k+Y38H21K9zrp6Vh+lc3A/17oadIxzU412ypXay
TRsHH5AHSjIvaa6GA8+BhPC65TvmKzqAdAwVYyvIczQhFRLcdfAmxc/hBll6TGEl
WQNtJxXRVEm5t4fy9HwrdIU2o0QMEy/k2IMkE0GhG7yaDLAn7+tpsQV8r86s9xhp
YY6e1yn/PDieNuHb7IYgrqUl0OPgk31HtPtFmjaVDmpaJ8FfFgEzmJ1NiPINiK2V
g92L7qt/2pSTcFh33n+4gkLYjlXXOXyZx6TbOjYFRaw1zcfNw5+RGgF7FkodeXCa
p810ofaCrxKlLaXbwyXqJRXlztYlbMGLOD8Ha5ca6sv7hFmNxyDrmKUJTc40wW0z
FVozERuDGuB5aUFn62YOeN2f5d8UmVXHonePgJ3Kq0T8rnpFs/qGFyN/ybWLf7/F
y4suMUwGNQpXBNyh0n5xzMqATGO3cw2XYGB7ti3AdMPJtQj8o7QudeUJ6BRfqEOf
Z/b34N5KetqvEhJPh7GBgSm01Y9NXpKm76MS9+/IRTSObAYesBeTFzJa9eu3jsH/
YYfhqB/MNyrqeAFWHgak3KvoVy/b772YixqFOVEg5QJ+ALaupG/Z9383SO/yiz0j
v0BIFuF87zCeQlK6ZeHkA+9jTsC9RBwbQBpehF1/RWK0XamKAsLCfTGfhdX8XmBw
sceNfNoEvykEdXtNpA4gujrMlRqn/U3hdAzn5zu1mKwpAaDQWzAtQHdDg9p2WAx8
rXjjw8RgBvC7tHLK5QNCMr3KO79tQsv0PDaGJIyAX65zA9JpK/Pp6jbOApsNQJfL
ZeZREbqCjF55MpElt4RYwB7SheSqSS/6H05OJaX3qFypxm84qv2LP7/1DeJOoAhF
6b/TEbQGg4YCjOlJz3FemZd6/+e9mlc3SGRsTX1LnuXE6Zo6/+Hjgy+79/431Tph
phkZS06ww1g8TOZJI4aLJkrQjCGFhtpFRKoJ1nqO2/zFmgqY+c666WIiRzkTLMFG
8T4L65R+j3BpLnNiYt53emGzUCMoysLbPYElca2IxhydDnDyy7tCjp/Us7yZjPBX
HDEgoM5pYmA0QPZR4Nc0lYvKXeRqo+yxtEp+QLmVTPHPOznRFrMDItTsjafkWU2J
S3tOTz4Hyo54AEl9Zv+7FeWWOAJIcyxyOQXZQNRAjeoTb49ZAf9cKOtcpcNAHwxs
Z4R7Em7a7hWDpCONfEjgeecnC1vAWhhb2Sh1d0a7zorL/5twOrt308Aqz1r/sgeq
FH2uRGB/SrlqRVjlO+xJTKxuLhs7drwrBeGC4Qe+xwFrvcWloRUY+0jbGB9KA1CN
ugHOT8+u0JFif5/405vWHzGi/LL0HxD3frVBNSUwR3I+ryJaPiYoPkwVrP+tYNrs
E4ASzyO5vrjNhl7KAa3QIVBQBfUYJJNSGeOm4OoEnbfIlYbyq5woQZ3RHeYDuFUS
WSw5Juve78JP38nLeKVuJfKfcZY10hwKe/e0VUcNf0xt2+KGWNY1aQzr9MjgJcus
2HVf5Kz8bPUZ4YWsyD6rljaJcpSHja03Zyz9kcQcNALahU3xkpML7NzxcNkNIeLT
p3yIwtLmIyB3/Q8Gv+w148dvG8qb7q98FLCygqHKrFa5DQ4/cip2JTYQqq3q50bL
iViHA5HAwh5Sz4RAingl7oMm77CBn1M2Uk9jqGCGaA7k/Txqi3RQoRoy6LFqBDCL
qHiIOGVkCw2uStoNg9UEZ7+0FeZi2s9QKhrnEhU8AQbMc8Ver9F6Qq6McfFL5PDx
lkqTbEfYNuHR8Y6oS7COA3gNxFEO+osZAmYq97dk4+vevpVLQ2YBQMjEwW4YL2Ow
V9tSIcdHTVE4vCyoJ+xauKK+xbCjhCn1Bc56pKooZQ/uspguDMxdJwgVJRU63a+Q
i0esaSyPPluEYhVX1jJr64xIBSINQ+BdKN94TNa5CKE5sz6YDbNl483AjZNF56XH
NiPkWD4BD51sebJp46zOXzPgw9wgYEMgdPveXdbNfzqWKzoaZeJCNlNZfzBTQDhR
k54K98W0sPxebad4C14OwAhWo26D92uo4WrJez4L/WCIdQ/MItASatqXTgKLD7HP
9VgIoxmlyjUA8RHLnTFLQsbVqbR5ammZkCjfLlYZ9lhx7IKkJii22hV1PrBP3GSq
Sp2ltlPVz7N8A8wMZs9iaHwd92Sb826pYa3niEKmX0BLpCPx/p8sNEIGxWKT4WyW
LZE/lYCAhE9+GQy2ILOfJWaNe4byrnaIf5YIe3I54in6yAlFJUnlBnMvyXuQyruO
b8R0YnrA5X20/NSiGc93tdtLnpxqkkwaGiyiwJKJaeAVSpBdVMIDkQDrGD+XQpZr
sEHJkizkvcN4lynjRUvlLqTCmtFB48QkVJk+39oJ5u0KCju2zyu8HLUS6+a4pHlP
GZZfEWHdLz046/ODrKOZq2WSEGk6GXxP/NNAW/4DFunAEONtH+bTDGJV66BTbO2j
0CCe4VVcXi2hg9BxiFYimGmterysG0BEuFXn7K/SnEyqMFzV9OFg1FSMreWugcko
jfS2YQ36nXB64Ar//L00qxU+ERu5ht6vLMD1L7gRcOZkbbJCrxZ90kvbTZzubEXr
hYUtIWn/S3S2CtrmYagbrgELMIDwl19A2p80uNyZg+EantF/0YVM2o5apOLqCDvn
JI5QApcf7jMCROd0jmImIMDjtZ/V6hGt1Wzyze3fa58gedK2WU8vd2GkrSweYCBD
k9gicu7Qo0sawZJebtvnGVtHIu172I0IU7pLspp/I4hbrT0T1nSBv5BaWWAeKmHI
KcoRIvP64CBnIjQhBl95dZy2DnLCGhdEDOgDugeeddr5wCZt80gTOZHJiBV09V74
Z0Sy9+128ggH/4JyVLTGz4a6UacslQ9n5cz5uiLdeTHhb3PCos0QV4TsxhhrpIqe
92h5FizmSwzdCFVy5GC3motuon3sumT00URAax1FqP+0mSxsSGoDTkRvZSoP5cTw
LJuync3ruYlK0BOKQsLE0WifsdDrQx6RRbFi5656KtY8FOIy79H3+5wJhKpJgGj2
Jc7alFIBSgmW9JZ/gKhr4rRVth5Ua2mS99pRJ6OrVhPH0C4XbV+Tu6zxKEUR4e4V
LHt/+9y/ZQRE0hXA3Lkbi4GL44jSgVVr3n0dwnoEZJ8H+SACOzE3isOAhOkWq9bK
8BMsIyvVY3jzY0cxFEPAU1F3469I8g1nR5qRQx53vVNRa6uXmtL4GdUwKsQJA7OJ
eC+iBJOxgLCq7KR3xREWMolU44cu52gsc1OmgmFl+83pUaLL/dKN/UipVQh8mhGo
KSeZv+FDBHpJ5PvBEqT84+Ow8FlBKujA8YOz8PuxPjgqmcngYrf6wRAhlxdHK3WT
9Phn5YZNVr5d0W6gRP/X7rUH3Hal4RJ9JKKYb7nIvy42ecXqtRFh2QmB6guZUOrw
UfUDVqGuDoFiQ/X5TcEHmeW1fpIrs6wSq5mAP35gUr4ip53YlycY2z2MqM0Bt7p2
urEZZ0hqIaIJXLX7gM5AzhpRoFzBr/wY9NzknzR+eTMxDQm13PenyrsJuzfnwIJ/
Yc73Jz7gYDabhUhKy0sJe/8x7PNtvpqc+aKcA9CTOLcGjMFRY8cGvx9d9s/J2aLH
ofoiGybe/MwtVt4d65eIAFCN3uudzGkMWAOArSnmbgSHFxuVRXfRTamx4q+c+kYI
ZP5/TBuY1ajA4FNbvk2ilg0MNWnoqI7R/DJ0d+y1PuPT7jazEItzoNYcAlQxT3ub
aF/aC0wjOXw/9xEg3zjM8KVYRIlv9+VAqW6UafBuRT+y2IcWufLgB9qHQWTbINDo
rCC5JzaNWSg2ymskMYNXWdxS4nhqFh4zAyDB1laHYjGDgnz9DiGxVWtT3+1SEg+u
hUdQ2ODtPI7Y8PcKgNqBi50HchOidVMDcvkl/0HW39otZt/10AR3BqWQYqYTF0AB
5P8kWlaAm3WE+a5urHziSGRx2oQ4rhDCij0UBSqWm6yjXHhD7wQWWO2tdzNIK87M
+81i76sJZ6tDJtHyuYdtiKdjFKtGJhkgj1XDVSkxcybWPp6JGX0mQx0eGlF2NzzS
gbfJUkGnWOZgcVezpA776WC0JlUN3v4XgFOgIRLUnhkgHVVu9JYkPoyBXNcbZUhg
9DjucfbgqECiY3+bo8P9Zh/3UtJVJO2IEqukD+Z81BxIX0MJldjnVrhlDd3RdSGQ
mX8p5b7GxNLKzjzDwq+0nkh9hQDtAS/MI9BdhnFdwjehZBaQiwxPq/uayoEJQg6+
n29YwOciirVaOZh/SdcV0LpQ54DaJ062Ap6gyG/H7jPiTLfEH/Ms04iYE0vQ5w5W
wIwNMW+JkbiAk/UG4vP+Zse3jduoL9hCxliv90irJAk7UJZ/AvTLTczYvTRZ+Edz
0gV0qMDeaFz2ChWq9CLa0CdqUwlurbC1wjpnKBp1wXCZCrrWOOQeB9jI90ofQU/1
UVRBlTVgQbKbVbJTf9PgRtLpHWNfJYfLoohAXvsn8E40dJwUHzxIKwkvLmd+vHPR
4iovPSxAEayu0aD8zgEmp+Bzoa5IHGnZhnOJiCvh7iCZLgDxIb1+X/OsMoHgGFTc
Tj6Bk4tmeZRERtzspqSpMp6xRyBDZQ90YTOx2mef2Y7rsemgqJXY9md88c1Di9g0
J+Zcs8HQI9PA9CTs1a+y/qFfH4MBQwJo34DkjIX6Z/jjHNIP6KHpcHyvFmsHDMRc
RfL+yrpAWKXNaMmhQp1Lyd8elJoMDnZKERVGOUZfmUuMQuci7dHGy51UXlNUVLe3
3N6tKEOPezX6oPTkIsm/RInndtxP4Eyq3borzgV5xSzInDo4XG3II9wGavwXTkwH
F4GdmZZ/rX20HaPrxMghIat7/v5pdUgKkasXucROhPv2cQYD5FVhX7eHLd6R0NA9
gLKkTYD2MUQJXQJaQyyTIWutuanLZI0zNJajF6ee2hj8hO2gPAtkBPDUPQll22Il
ZWjoTZ4u80nGhkrlrn5y9SneshTvxB0vGF35E7z9bJsc92+zIoh7UaHb8QV90c+A
a5MHvtQnXX0pwKYqihTDEkj0v47awgkyWBUdY3FBrflVEDFMrH9VKMlSOBCyIFuY
tL7aQPQtfivdlI+zJFalS8GWWbII9SI8CPUGGODtCCJMfZr1/WU7h/LiC7RiTekJ
WPdQMa9rm16oeISSjy/7AiHIFRoU8rE74JAF+4HnWfOhziX2hOF7lJyvkCiqXp8N
ju8QG1HB2727S/+vczeAwwLCR+uZJYZtZQxib/LDcz+L726yn79nopzRZvmcdEWt
gz4lftrP3z70z+KmcsDdsblbG8o/a16hMR3yveTJDm4v1gcqVd0A45vvqTWVs93s
3QjRdjMV95j5kMPiO5oGqA/weFqjR5a47lmN5nwcrQEN3TfjVlZfyVfjSo59Yxty
1rLahewZR/DF1D3eyt4lUXrd5LC0cYWCDJ7pw59eSke8Q3Q9jxbnLlqpRYCAqSjf
Wis0ef+2a7tzdH9Y6Iz82p0U/suWzYjYer5ZJaBbt8yiPxRCaWUujYfWMlo1IoHG
+cKS56rdrPGHLH3xlxYUITNj/ofeHfaZvSGzPgne8O3OOaDyOLtsMoCKnVrNRQjy
IuzMXKQtZQE2Nw3ICVLaHu8Bgdrh5RzTSgrbbiqX/ahvzD7b+rNiJLFv10SoMwqB
aayk/Ulcbtlt02n7lRPLziOJ4bMS2yXscgzIQSgLM/ssMuJzeOu35BK5mfJVmFdA
EE+mZLw5SSjeGWjFrch5TDkbXsKVbwMGUJOLXHKKL3tZ3KjdMYB/Tkb3Jj8oftB9
wdLpWSYYSswy2gZXlCRR7JHNX6lTrPnidFARBKhaRU8QMetmdaRxLYS89pGhGmg/
UxJTi6DgNPI9m8Fsl7cRkUOnEiYm5bVWLkhzHpFPYI2sP/WuRDl7YQa0ZRUqr2qQ
MYhJM4tNWQ3rD9xyi9YF6VTqJj7ngKSjGm7Iki536jzkV0TmD1JKUq23dwj1eVkR
yRneI0ytBO7rYYUihILelctZtkSLmdckGPvxsLKrHzFlDO/YlkOD6mKBanBHAdZA
CbY9uH86kLt1d/KkYSbd2bF+VSwT04cXoMfzIWOJuwnQIBLG59vmogtUJyG1uUMN
hJEX8EH1YxyzFI7gs//QEYAVlcm2pklQuZxrfE0KvrPqLNirNwXuYdWksAX4dFk3
SJh0tj+6e1ky2OjEq5vmB4KzH5IRRWlS10P77oChu6Dbf6B/eDTi2P8c0JD2mB6+
/eSeaOKT2qiCRrjUMkcmaZvRUcvKSah0TVeYk7SZcZMDNfLl2S9pSOQSkajOXNC3
0SH8hiJd37mv9+eRE7jcxSx4hm5Simnq+prwPr9/0uIUNTKIwlvVDCT3p1xwnAcd
qgif9B6KgHQG3ZXQ7PLAz7nXPqpswJ2Edrgc+J3HmIwwlEhjWPMXqXEdMRnXQ/0H
K7gClejZSfencx/1mZf2wdToWT7M7CByZ7hFg3TB1LlETH1rb/qyBzrQIEBgwOR1
avyyK2gkQeYPty6icSPnu/GSlNGVKwlJSzzf4oTZLwcPH1ozPQW5WDz1t9dcDpej
Stv6zhDNRxLndUzuLme1Hx7PGA+wBdy6Xz1eV7ED4OfkXa6hthP/kgblRINNaCEe
kOcSgebzKoZBNz9ZhN4LuSzCyU9BsyxmRJmCkpzVcQJWIBH/m/F7r/ldZ6bawtHk
1widMRprlmjQOPH84Vh9b8OIzOPYkjzGOMu0hYlbJML+vyS7xH5fd/4yo0zzSkPT
/CGD0HHnEzJDAr3TMFmEx+XU3ocHsIedzGrn1KphEDeGbzS6CpJT1ia2naiq+6Jv
RHmGNeQh2W1axQVQ/RgmAgaEnya0uGcLccE6lQ2Djr8n+ElRJKO392glpticq8i1
j9TTaJkJY1mqXns7M3YseA6ZG3cZtbiS1lb77dUtCr4XENLwj7u55iG6n1FRyIx4
OITzq+WEL/mzWKJ1DoVAxkXg232bwQ9/bcClOH3Ws2i5VK0GXF/8dTqnpjTuXTcd
1IAP/rZiEdPegKQkdddbkw8ep6ZG+rJ68ehTFh5/xRJXxFj6uMdd8AYXSGxr74qj
Tz4sj7V9NAUkGdQG4/6sVaZqsd6520h6UO66ycWwn2exMEUtiFYBFc1MdzJiECNy
JIc+WWNx1QdG6HlXXzgt/MDI2cQCPV3Vp95zjfqDoItmYi8bSMmDeRXfi3HfhERA
cLtpOvvJvVwT+ljF57WRCocYnsOpWrbo/Z4JjzjQ+/EsVFlRLGka6O/+LvHoG8pD
w/YRlR15SekyReSl4yQLlNAHYphiuWuNJHsrGL1JdNkm2u1eiz5uUDfmxOEYzr0G
d38wgQzIsYC55Li6Yg3GpGC3NI/ktCm4ygrOLjZm+905zxG2Z3bqqZt2ky7n9WkK
4ubBNtrIFutqiOZUafvloR8UenE1Gnsk5+dP1vqQ5QN48kEks+ogHgdYg4XIHE7R
HkNHx8HKBWdgs+N2E2FlQSIrf1YN1VyokyKGPQ4KXsFwyAR0GlUC4DK9vT6dTt+n
YgwxxNz/qXM4Sj8wCDFp52OUWnqKPDBNukCEG2ejJ6VnFmv5BCiAGvhonE0pHzkw
2TiQJgzE8RmFmaafY7Ycw0iePr50/DZC5ERmoJueK0QgHNXQY3yTcOZDv5Rf/UOu
4osjzAMNqIjoSFD5wtfQBdbhECXtOM3eqaJRCFPYdBsCD3w74Becqpm7AfwbwLH5
J3VnHFI1HIsceOY2tEsc9sUuPUTaftSyZSjkaB+DzIlq1nNHB2gWpONJ5o5joREX
I8en9cWhBD4OAf5FPXIJitzgQSeNo3h/4mzJNaCVmXkpkkdm2o5XYI/W+Mfge6X5
hHWro0EZU24HC+EsAcChx7dabhgh5o3WBn5xoTCq4x6GpXXqCZIhPcVn+qpm+wXn
TCfE1WZSX3LtiDmwH0JsDq+btwgRcbEI603wiCS/t71ITCmTLnq8Mt7RMeCnD4Cb
vvARyxFQgHcpcpepMUkmWPGrQHewoE89Um4U4DKEUMtJNC7LoZ8YLLziQk47p0Kf
qVymSapKf+xj/VprFAmNdPpt4i0KfW0Sef0sKXOg/OC333mrk076LZoWHgOKbHDM
bUDuHzkuY6KwqjwDojJbs5Grvr1+GP0kbQNnNMhG5NL2jEGzD/hndet5TKsuLZ4X
d/u7/t6Aq/H9lSwnSUko2gVaQQJRztzxHiID5hLYX5sa/WbbxivO0SubZo2yrQEW
b9CDwGwAHUdjc8QZEZsl9jR2v8tHYEoL6W2qXlutmJh1ZiWvhPJ664lv2e8wYC2V
nRwnFAODUg0dYkBiaIlb6EIC/yK2iwgpC4FlftTYdOiMD2vG/FG0YnwhkXZYwbuP
HDr8cFmL8vgDtXuC/wWO3+tyePfshwbzNGiGq7RSf0DYwXnzisp46hSdknnrmp/F
9t+k/UPaJzUeqD/Gp5EPeAXoMVRklSuPZ+Q9WXAo/5FbQTZxfOQTuM+5d1GJwL/z
ms63CYBVgXBJF74/AITa7nhwdWyUJxJFAj1WLrJIEpzf0o5Obos07nO7l7j0Np+n
XrBw93lAgIa81dodmKlR26wr4/JeU3QAMq04X5QQRZIXpLebtqd3q3DLl9uEYmFB
z+FW4Dah1barS7EFa/qQi0dxgjyVAQPj7Pwav+7LLHlOtnQEehAEEUxKXFw1R5mC
Kn+OS+2de1hnDXwV/wSAPm/RTC3fOkRMBlcmWlMAOWJRsfFGu4WjJJzqOjVYC3Ns
eF8KHd2IrX7LXDG1jvf7MKJocXwDowdLL/sLeTHLk76ygYRSCWHKT7FYKGYDz2te
9QzasEsXQyaXZSzbrVdieNj5RLgtYwNKArJoXpVO3Fpsjosamk/oMMW8Rh+ReIlZ
GfNbJiWB4VcKKoi1MaWyB36vz9kQnETx/2dpCU6aUKK5mLd+wHguNMYoKBeZQuaZ
wURnGqjEI9/cAiyOyUXxe14TBc6oMU+fxO89T/YwGCvZydNjVoztX/ou1xchPLlT
XAsqCZJsgPfqY7ANIcDlPt0gL40IB+yR7L1ITXp/d+/LgvL2EML3Odl+F7I2S+eX
oN5GMSJ89R3dJG6GrNU6J/LktO/EeofUglp/UqFi5VRjX8cgea4lL/8bb2QRRu+m
ME6lfE6FwkhpscECT+rP9c3Ju1ZX+USDVVK7zkHoXEeMR1WA9ofmm4LfQ+hNNMEW
aUikoslUhyIGYs83zSILMgLIUF8fQ2dqs3xpWm/nUrq1S9Pj4hnDJ1JRhpbq+84H
M8lKWz4ja8/f1D82KBZuQnTVzO8yDW+7gfu7pzGu4BzdJORyon+YIy5fLqfCtmqj
PcJtTGSCrEhR5HLge2/gLMysc9FnkMF3SMW4g1Ow8a4fV+mkHx7aUwQg+hAHvI69
rJCrsDDtRYHUr+jao87W5374ZG0dFmb1AFC2dTGSayXVz9KGKfKRWf6kOF0Ej8wU
YGIoUTStcDDV+0XSAxvSA0aW4YJimc47ObDBwnyRMJQu3R3Ux7fopn7gpxtVdP18
U12m1mfBWLJ9oCJXHt1GVh6aFiH5QFoyPGRJyT+BPs2/4uoVxAy5/zgPeP892a+F
LghExDgPOcVHSvBIgxf7mNWk0cjOS77a2hTdqF0BniFIlbXfmKpgBD5rg8+9L2Ov
n4sxc80vc6iALg1mrXqU9N1C07NLgAr/mxlUByZQStQgRKF0PsGasSqgjNOjrkxg
OXWgWey0tgLqYfvZ55RDkliv5UzIsQY0QD9dCUNXqHli9Dj9/773kaP3Mh0bb44T
Fo9PI9rNZN+NETQgRIM/pK9xX6aMMAEiTiBoYH4hRUc8Fryveu/U8WRla+mzU8+u
4YgHdr0hTXtAz12E3XgnhPxvGOMg/y4ftTYN1PxUpP5unjdQX1DbgTIT/LG8jFVS
ahHJ5/1u/1yniWXi1nYiNcEuWfEbHeEJ5ANYQnT2qHF5t87qBFYIVHU4Y+IFkykJ
9QJoGIIx8sdJg4xnUOMKZJW2e08eDW8MMe1ZiSuewk70JzfWJCNfbhmwjia4t1fV
ZdRxPFuBFWuJaIUnDS+KL6DNBXxSoq4fBtEMjZKZe+ZI70+fB6m6IdIcHwQuLXct
HarH1FULhxuINicBfzEUZqZHJhwZpIaUE6zCStseKb3IURW9amV3p7mDfzzCPZBT
g3FAHNQot1RshHt2lqP19yTAIQbPfns+9pmPezYlSerVDALR+F6gapUklxZeUmsS
zViiTQ9tJ0ff73XRkbE9LOzHbxHhySZmg4YKLg1cnyvxJnxFQYkll6yVh0RnkXXT
AOfqSd6BNldo6YzRxwdxQn5/ktsFKpOR6lg0OWYB8/hw7E6acbdQY/ST6uKho0MT
A7AE5G2VEWlHTD3Az9E86y9Zs+Qcd2L0/y2QT5+FXBtOZkfacB6F5/LdMd0USJH8
EeOMVUhJs8S2YhHMZJFBBNEjPzNBU1S2zOyq9Mr9Rri7GTjdPHVCUKb68UtckUUF
B//peoXe3tatQdVU8sd984qvGXTm7PP/c61RxFP+7Gh8TEq5c3Dv6n+/klj//5eR
SfdkDAQK/ri75E6+pNbEyy28ifnPnC9ms7v/dT9IKKV9vCdiuRj7GUszT3D4LNzd
nesd7f5B6Wlka4n+nxJ3x7uuR3SQ+5VKkRP005h1teUn5GOXX8LWwWwEhxI+pMLx
YwZ/2s8/4dPsz1UOJnUvRXGkGvaCq0tvXfeMTryKwlDV7EPL7lDhNwFNMIFJkCLf
PCK5+LdObyF3gFKsWR7D8M/9b+g4ONEd9NHhfKX0QHuofvOE3Pozgb2VUTnv3m9I
OcHpGJJrJY4WDDo5ESDBpAuXv5zGcbzIyPG1JjbwgGV19D3KlpEFQcD00JmNOYIR
wtlw2ajpjabhvqXaQN4j5s/jZfLDSZzRrc04be4zt42KhgVa8/Ss9OHsxCyG1lE9
DAhXx4sIQMkrVoqjnIRF/6CEz24Y2GfxNPLIJrismB8OtwneTD8vJhyajA3BVc+b
SSlC4Xzjf/IyRBqGBBxpqhRegB1IUQ6MOXxaTcxYGJzavqZIWsHRz3qUsdus9S5K
3HEBqdn7iNuIrtwpSNw3Ga/DYQ3d7vGxPJ3+NTGyIDF1XPZ3jMv1QKP6z9puiIrM
qvl0ctIQIY//zFSQdsIVq7AQdMk1s6EakvgU1vSSeqvSDktn5SVOQCPdj0oPm90w
QidiOOK9DyUS1qmL3ehD3vWAnfkTq1r9A5J0I5pbejH10wam/4BsxRYEr42GOz/Z
f+RsRsHZNsGD0cIUZO67G7Chq9CNKXXqkpFmdtkHNNyscuhSjU1mJxrQaVTMe0oe
zKWhvwYPbM8dzXxWUH/HrvuYrsfiYgMlyIGC0UDpkbaOEG9OlrosqjH2ELcCTn8o
yqQBF6eH/+K6fMHUZ6zlbnpwMd2BuGniORVvIXVe42KjxM6qQuUCJX93BVmsJln4
rak/ZSc7zXfIlRg1zNcIj5m+OmtOnzj/UoDx4TzV/dhlWK1xAnZ42VBjvQLKwaEv
hhg4kEuuIpsPImcqxvIMkFEHlh0uKGo60mtB2lcSGBmY7nl5sjdCuWYIXIo22wkd
4ZiooIw9PLJN7j+Z52McJiRNcK1ZNfGO6fp6md8ONxyipxVJZimNmPmlTogfqtIv
KVFmMDFeIec3dMjttHOOSjBwFIp6neWuOhSxvt2kLApdZidQUqd2YwtSP2hL+YQy
mlb+TasnPl9g5DQ286cfXVFBELoNJQ8cCTqvkkEAft46EvDOAG4iSGUohC6s6wwI
N2qkx6LF3DwRhjxFc0jGFRGdCnVSDD4ho9xG/ljkAgYgqRrcLb67f6eTHbW5gQUe
RIxswKUZeC9ROKY0+8GeZK1I0bloFDGPQqjbpCm3Y0Qxr3Py1RP6vljhogNGY6VR
XSRWx+6/JljyGdpi5uzO1Isbi3OpSQRwqrb3dMX4Mjk/wB/89JfUhB8Z+kbiUMpr
5xW+s15bOqPSbN5UkESFyl96RoYSF3i6GasBdkR0RSSZ8oH1B02BEFSeW5VYOnXy
mofew1ahPILbKcsmnwonMUkapVBo296YmrpWDw/0Rg2A/3oyCvhYSmA5ZZ1mag6g
CuGwsVFH59LuS9s50E1HQaGiIcxoDK1UlM+UOf6B1gGYC4aS1jpyXtV4WJxxykWy
m4ET0lVjuFbBNO8OdZh4gbMeh0le/9UKtrq/gXUjEjjst+1wGwMI6tbZ7DXtgYam
XZWwikk9n9Sfz+uj7idESV5XtrYoHHveJXDN3z8JFn2AtAelBTzW8ayZ6fx/323M
Fa6227LBmgyDtweJQ//jLebHNgEYChrFvUHNrouVTAIQ/1khsZn/ZUo1d8/4qIJ0
B8R5wtN53ZmBSVZDqFkRKIzjWVQSmMDOfz0bV3rxpLpwNi9XmZMyxKkAn1cbVPUu
kAy4+rVywMXYEHmeC31iZZCzrzvpIRCXOaXnZjSJYQLjxsrPQ29ccbVavetlS7Vx
NZKU/IwssnEKLzZcUTxN8+NnceVTkb2kHErdoa4k+bxbxTjIfuAApR7+W2Xf0Hqe
zf4R4rqdQEc30rVgWOPVMwyX7vinRavsEaRAKO4Nt8dLTvUG9sp9VyzhSkSByMEa
Z4cR5JKU+/d4E8zSTai7djvimZJYbY+hoqzCaqbWe7FQRFGPg8eXJJkVfcrv1vOS
o1T05tKuCUawddSDHRj/b+Rov+do4N6pWrELTfqf/3x6d5EZCWS2i1Xw7j8zr1Lh
/RPjMytcHz3aZVvd2BAnCloRHTLU6EfB90veTz7nG7RP3LwFrXcDpug906Nwy3rN
AHGzfXvzgeUPX3JEOFuuU5nKgjKlOSdLNDXGw9z6ds1Vz5QheK1crqUXEG/hPv74
Jt29k710WtvE7hEBxvfnf+tSu382EcRltKIf91cVg6e1ORY1ha6vH2acXyvrDR++
t1TnRyMQ0f/r03m0PW3pmo8waDsvtAA2a/dOs79HD0cOyaGWXYbChPVY+nMrrVA3
t/8ybXmEZalDM2d7f/cNEQSDWRiJDXX4n9uC9J1DQoWRmJ+P9/T0R/8CdxZ5x6DM
+uPlntOHseSSseB16hJPF+c+EjTcpGdHidq6YEUhiSvRAsSYqmw/j+kk9TopTn/E
8iKgzPHCc2dvsBpMkzpD68bAzVJLQfEEoQPbv5oUhBP+K3aCZAT/zefIplmDVOeu
p06u2GPJeUQbfI675Hy+mh60h9t96VyePFNZvC64OVdpt5wr8vK8byUGl5X2F0Bk
WvcpjY9f0iadPTyscnMXT1jtGwPv/YfX5/QLGVm2IDk9WDryPrpTppe3HDLex4H2
NZVAq3//u3GVkkN6pSWI60HLd3ZEyaO69zBOC4tlXjgWLAoBbpKH4ivL+9BA/mab
uZ9eTZxUIYwattQoOUCjhFIJHicU15WgLiTS8IqCWbIQ5Q5w0v4E3u5ckx0km5Zy
LZIgrhvaWRMS4eiPFwyvJyTcjkIHdEbfEJk66pDYbh+Ft27uu82xsjj5n89sojbd
3Pvg951Hsw3NvvbIIzeW1n72BzbfGqiRX0JeDTAC5AYO9s9fFUtXFjOcnCbUm1jU
tv4JYH79fbfmNPOxaIdAeXQFtwLWOVTnUpmW1+hsCz/qjSY6iojLPs4JsSgok4+3
GNgai1pnoRE1ktL1ODJaGDcKO11O6JhJLOLr2OvTnic3hRR5jg8mGKV4j4QY+ECa
k/RpgWlJjJh4A9rDhJApo1TyewszHoujr9E6rdt1xzqM7pajG+oNegnMJaOJq96a
lhxycXORXg8SroPIuyY0TjoakmxjlL2EmG+1Vcrb9CLt+83VXjS68Bessj7yaA4p
axJ3VYfsRcCz+rL7sc8+lrZdGWgtlawwWOB0HPPVfVBq4fmhcqGpQzQ/qWkA+TIv
7+vQ8D9wEPRfalBoiOuyl6ZDJCUvJ23PLJl3aqDn1I5T8kIp7enNVxgejHHedhhY
fs2ELZtjYnBXEmucFyGO3sQCQ2wXDtRSnItgcMla248gXPs12gRp0S/Bqa6s7mgz
7GZj/M3dDXnz3Szafh9z50zcI4Jygnz2+jLMh8f1A5sE7zyUhBKaXJNEWzazjn83
MRlorYcg5wU8l/LduFer5EVvQl5TPrSTXGUzYgTK8376TsXI6n6e9PcVdvgHSH1O
m6ce2bJaibZLlbXTa9hv0Wb/pR/0bBVLr5wyCeji2cHdDkgzaSUKdzAAgIJyAuVS
U/Uw6fkxox5N2LVBq1875i59e3xs/O2hvrr+NcCpTgPRTHjJ+0jDufdc3pVktN6c
p22rdiOEWGaU9akZ7XwVn5TdcnEK03FSsnjFuUGn2MNSZrdCDuItqR/T9hyvR49D
wZEVFassvRew84ldvm2g0teGAdsXGXXnxlK/+CFzBQqfstCeI6xLIBpZt8AvwYp+
70QaeA8u4PAAGNFyw7jTdOXzJjOC265JbCkpWU37aGO1AzUHsFH0+bO3+8gNYe69
/TRCKzIY6zD8dzJVXL8B+Ga7BSlXV8FPGnREkNi7RjthNmIS3651IsmSXTaYgtru
3tzz9wdlD0XOZT9ZUj+eUc9MLVNiUXyEkRNB7eGzTih4fx8EBclneskZLGapY9Yv
pvrZqRsRHWzg4YEeAGt0LVzfhTz+YAkvZqp34fo532dz3EoP6ivVAHSjgvfxHyfP
dThvCwo4orOYq6wjlFifdHuTvTVtHywNYXSKK+SrZJccWRjpJ84THGqqk75b9rCc
3qAY6ZLLnBHiMIi1a/ovOkPpcx5jDrG+bnSVW78esrIcAZNZqf80beM6OO8wSvWc
dB56/hFN4IOFUoem0tK/o6IetG0xE6/rR64LKHDY+5GDOxELxGXDpngJPhk34vPH
6FqD23Aq3ddsvpmE1O1y6SU/4sEwNKbWiAEXO26gYyUVOb4ce1CLmRXU9+iGSKoV
mMOKADLzTCcqFLVMk5jFxlXXX8h42J9gYFdQPBmvLQRraB0/Qw7O2XQhrIPVoHHf
Kji/3ZpThedp1W/bkKCsMkRPapw2geY8NziIdIl6Ib3ViVJRi7P7wiKflk8kzgVl
NfNl0+vnSlVRLSpiZw2Hv7JUEydZzVLvJXR+hWXxItPHbZl2FtJ7q4er25tlHQQk
hWuVsnJ14xzumcQRgSTRu6Cf/IT6Lmb9HqCak8DgVP7DrTqfScu6woo9VES1iEy8
KYBmbNNw+jivsHg1U4QJD8goZ4Bie+spelOFLrPF/IQLOsM5w3n5bqrZoIPtrPl/
lG0Z4PcocxGIScpfkpZKbwApi+CkWRvZK2ESK9+61VSsLJe6O2m9m+9gYHrTOUYg
HF6ozvmHvoudgkqIeRxksXeTVt7wcsVVCuYRLE0efjQZXd5+vzJ56JB0J29LTWt4
OeMNhGHXLDGtGhvzbqS5UIefIky4TZdKsqbgpBJtabpB/nR7uSN7cBVi80xoljBq
FeO6F5fv+ApArePrar3H7NcdH/XYNg+BmNDwtS8nxfX2M4dvnKCLpkJeYXb+F77L
FAVuvZc7Ccp+rQlWrSRbZpCCkR0U4RkMW8nvn2TAqaupDIdXJ4/TOVlxDulOTukI
QHqpjZBOfs6AbTo6GmnRoI3cT3yIinrHDMWFULKYALzpoWKW240M5Qo87gQ/Tw6m
cv628PaiAryMBaJwfZq9rLlEkHQjdZNomi9IH0f5UYigQslpdykgFhlzstCn4P8r
cMk+I2BuCwALwz2fWHIQH7IhZCIrMFfGkXu5WhZ/tY4K2O2kv264oYcDYQfzzRjE
ORwr9F+jzt4CMXEfKFH4I1QJ7oCadNNUK1+qtv6ki00jqCwwI7NfBKdI7cA7X7s/
I+TNkHMg6eeDtAqkqlgJtIXLYQawx/BkIkG2cK0EqzgIjs+FRije3o8rYbUl6n8U
9CN85DqChdY/NuMwIL0C+c7HZT9YNBZWfyLbqDUWjyq4Wc48TBxNy50P3omOWg1T
6m+J7q56yrYZbLu4BiaSYMuKyF3emwU18EKFlLoC4suTDIP/+Twzxl5n+X9IyMnq
dk4jjSKrcHWl4l2hGfCidLdwKa7NrnXkh2rcCVsSwwzZ7M7X5DVL5uTF0Xc5lg2o
+GQFoxt726pDGUK9TZX8S5sV2cvoGRkcyK6y9RxKtSGH163xyEpwjnm3swLdasbp
0GFuMZUmo+k86yPIn/dpfew+w55bNMEqcw7lUUHyGiIVxdic4d/NNcHdSiMCwHta
rZlKCsfj5xIqn3JZCLX9HojpBCZHKtRjBiWawqqjCl071pUxAL85R4oIR9q3aREp
ZsTaB32vUWqXRE2BGQzQyngo1zgE5krhBD11hIBwtyVuM4VdyifVF/YfZ2OR6+J/
0MeIOI0p5hMAVHypSLpapSMPC7ionIJNjFYJSYyTy4EdCn5YFttStLnhuYAKQacm
jwJKLl8wXE206abBwVPhwvsuiEMgTGbupciZQcrWadzRmmeluRn3VeBFZCt89BD7
R0kzBf0yiDnYukBfJo7VRudL6KD84yibEnhxdzOJmPQoggO8DHCXNYbxrTu9HVcK
8NzQUQTkZon7KylZ8aNkDODt6CgZfOpqEpFVn0Rg+kUb7tVPXy5fJ8dHinJWcySv
qMMTvc9pvn6LTMOw/bEWYWhu+6VXXY251YeGfx3diMxSbdzbav6VcOgNGyZJq2kv
d89bDeggS4ZgHQxZEInTTW+9wEZfITqG9LcxKFJR2nulTnFsHARmXNhdgrBXSvWy
9jcDKgY0xeSAJhhSWA9X9UZk91StEmCksZJi8hMu35g4LJv8I/C83uj3UuATv+yn
y23b+5ffFqJOl0Qj6qfWYYe2FxKb4e+Rp3RyZoaZeLd4cN92YzmgS5+MH8sblSAg
BMobPajbvbVY+xvqYlx58WxermmsBz3sT2kQsClrpowcoSYywVn+BFFhMFBNGUWh
lXqDLdnWY6KPO2hN77/iKdUNLRQIieFraesYj/aT9tfEpcoPgPMaQyEwGSGzHl58
UiwyGpcgvEOLJtCzJro0qRq/9CJ6jJZriCz0nGOKDlvib89ymp5TQFAC9Sx5M3Lx
zjJIl5IwK3eRKK6+RRqNfTQNR160TKIoXNuGKsE/7nVRCxX69fWNuiCixnynTeXr
Vtqo4tos7u/poFRaldnY0fnmxUKZOVOeTi2Gp0MqgqWXehJJsdzkzn22QMhCLG0V
U5HXLIRHqTC+uy7gmBB6o8JwSZTc7I5jhSJ3KN27hK92PtSRu73Msb/2riSIUODd
dJQ6+yjPiGu9evSgmNnRALhcdt5wqqZKRCPZmTWm5UpnsNu2dlCPlpXPeB6HJn1V
PyCyModtn2snPVCRGYWkyX7GyKGbW5rVIPsah9GxOBPS1Y3T00az3zJUqvTDo1FN
qBmcl/m+DQewNhhCU8tvOiJoEQizFLLzjNwg6RzwHjAYSnrLJGMHeJ6wtEtYnk+d
466ob95pvt3BlB33p9pMm19KO4fpShLojY6boA36GYdldmNVT3BVQ6+PRyXoSZsS
eoPCT+RmNQALqD/PlYKAZ+Q1VFD+f3HDbcQQMFI4vuYMjIFWJbMRzQuHY1LStBkO
kWaHjb1ER1Y1WJ8mflIKrigFigIa+VvlfoOJPSIYafgxglFw04dg20jr/Lly9XIp
sJhh2166AWQKrdT9mzC+oTt0Gc+LTVfDv7ra7Zfbvo1dn1S4roxsS7cf38c9wd9f
JQSGvmEQJp0o/AfzxL3IHcZTPgz9lYwbEuLyqU58xYRs4OID5gILQayS52ILDMFW
pWdjG7Z0zmTSJa39d86Rr55QRkqjgRRZW597pntrWs4E9VIZuIdnMM+OdGfFUZT+
5LrhIHoJCxc8jxqWxJpHDySbnmbpFA/leDjvPAAOV2Q7FObxPNXHO/oeaKn2nt80
IWEUBqeUHwilskT/ZDaVNfrv5BKAzohcZxPjCtiWmA/cyN1jFWpbbRVzkW66AMvX
x86KovOgVG3IFEtfJktJ4tUXqGwuaRaMwKLSeQPJKzojn8rGZOW5K6xDy/2DL1Mh
1cJ/TIEJraEKqPi8M/loh9Ihs+ny3Lj65Ycq91jlbngAM2RYwBXVLJ+QYMpB3Hzc
0qDdgBl6jF8altDxo9IHpUkiURMcair2X+l/GY9WHVajynE1hILVKm/6Pbr8URWW
4m4VRdVzoLssp8HsQqmrLLCU7dQVd55yLPNXJlX6RMHqe+7BYNv7lMVEX1JIumhc
tqCbi/9pj3rnlFzkmotjJ/icVox4/6HTe5XP+UIZiZOPLSu/THCdKCaM/q1yWjQK
SIuOSL6MhWYX/3E51HHpuFdC1bJ6V5GvI0KWK7HLGmXzE7TW2ps5URS6FeQa86lJ
Uia57n/ADLhtPfbFlr2CpwMXVrEq+0urU32pIqJBn3JxV5Nrbu47GUpBAcX+BtnV
Us+KJbFshdEie0HPDoURXv7cJ3TP3nKn5NMK5ivxEYTQYaq94BRxg0B/xjjGJvNh
h52OBk2vaFYUToA8sYlkzeGkOWLuBMDnnAVfpea65LNgl/RLu1wc0xUZzMzYJUGg
st/3S2T/3HfQDF9rIhAYZsULxGIV4JLfahUD/FqPZ/e4N5p3rq18ZYJ0nD4tgHqM
FFWMsdVJC+SjPzbqAKGFmd3nQ54AEybflNhtxfmOs8mHQQzy2HMwhWc4h7csAUE/
aBKNYjb0e12zGXshhZjEck2/n8K6oySQ3DILRxDg2uiv7EHHQvEvq5ZpfVr/ttBA
aldiwBZy6hJ9UHZ78S9Od5axLxq9pK9B43D+jy9/MXJHEbyka1NLFehesISRajNw
MjCOBgtusd5iszjpg6WC/9VKQPdAZ2/+W4tm3iqB0aAnULW/X6ZZpnn/8R5qTGAG
Te5lXWB9NmS2gfwLfbiqWbMeaYnuN93SdUScA6nhTt0rYzaoUbbbR9LXhXcHh8U3
XdQ543jh+V9/PecIAmZTJAvEXYJLYEzrixbn60Hpm5EgtFUoqn1ob8HfkSEoWTGn
Zc27WDfBHCpa28wsL32zm2bZ1dWMXW1cdTRyHMs0+QpwlDSkaz45Riakb98HvXS4
4HLCaIDRnMrkDBItQ+YeylCyDh4/Hh7kwOEhglDKP+CqDjKcmc+AkHCMf6vlYlbj
UNapkSOuA5+A3Mbfn+9JlYE+UaJn293vJTqT65Z+7n300j6MnOnh4qjymujxc5qf
79Q6K/BAYBVXUtB9x8XMgZjr9dbh/Pl4W84OvSWeSxit/yHtiTlWLgXS3FzcoLPr
DbYBHdbtT4h+nBCgMOk3cD4Zud+XfIl/mkcPWB+I/gvSMuuUSLW4NZjOZSRAMDoK
bBqXDAYUYIm3CDDq7BqB9dMtcFhB+2Tx4ZmP9ovWNg9+ny5xyPqdfiHGmlBZ4bvh
+wBPOT1q/seMC3BmRlooPy93qQ0iy1Alb1a4UXoC5KqVPBNdxeUfWlvJBCFipkPh
f2w3AhQnna7h3aMTiFp0Q568w97DMrphBDBr7ypHe22Qur/vShYTqU8Zd3LgqbyD
309W56QMrRCBw2lT7JQjVW3/FhpZ1cJXG7YLVp6eNLny3QGQXTRXNqgDnOoSWNuE
kUvV/uCkK6Hv7QTVp5huzLd4Z7WPKhkdeVw7Cqx645bgljEqIjL4sKMOIdjPnUNZ
A5ISZ2TaB9hb9/9aNjBt0T0QuLWXB8FH0U9yoVPita5nBXQsGsOxwCpjrjiT9ItN
2K9GRwdsvYk7EOHQ/c1st2Yp+/2tjJBmTzZA74njbFLwu0HhtIwGas+8DeEdpnkP
e7XQCovy3Wt0+vCGTXrYEycNbrxNkXQCxCbBOO0MzvEPrEbLoFYagzPMaO+yd55R
LvzTIhkM7E5d9eEJbI9T7XrhVwrUdlD9YHv5ukkbJPZNtfg+XZOy19qOM35740sc
Osg/qTWPFUNnWNMWn5NuL8k+IbbqAqjk9LZU0GafkadCmyFCoIoW2iCHES1YoW9k
g9/YOgN/8Cl/M29D/DIopYS8kDGpVPH4BIxpQ9DKvJimaJisk2mKJV4++9HE4Xtf
LOv14PGm2boKu3ttxT52OcTmHURpbFpOiX2G9UuAPZsFxFCxBVupUasznQQwV0gD
siFym/N6RlypVi/DcKeW3ynjwvV3B+7E5dK3+8mUTlzfPwhv1GqMPI5/O5P/9HZh
w6tUTHSvjvjk9ZLH8z7HiCeA+9pFS/XvbH7nEgYMIIHfD/lYtDQ5I7xY68KrY9MW
sh6VeiUiu6mP6zeca8bZqQsvFORgqqgpA/5ei5JF7q8c83KktDNv8VQFAdYwi+PI
2h1OhYV9QXgrmSjk8gYDUUG/LiRPpdRfS1CP5y2eUgyNlbGeYH8vstXs95bHjXV7
TWjhfVqS0Yjv4OyOzYvH37/A4Eesu5hSyv2wsSFiVQY8W/umfcGHa8Vt/Z4fEGq9
/v1wU4DHcoaftChejle2MEh8Eb8LUGMcUMPhx7sb/EZsAo1JKsAkyFwT4o/z1UY+
qu2zvmFXyksbuSspnoSuc0aOi6Pc3KqNDWr/r/1hS3h/LEliwAxbgWi+0GZZUB9L
lzm4jbS8OwcrkUAeBuLppTZpgd1TAuKRKgE6kM3qIPD8tVyhjHisk7Fyb2MDOqJL
hwFvG7OHVPx1FMnHC4gqtuVDe32KxeNapjgXLvH6qIe6UHJEcXlhewrNyl0NNss7
7YG917QrxGkfmtOISTLnaqruxj+9/C2LRNt44GlnAfTg3BOHFf6ZT2OHl6u81AHb
bYgXZ5jkN41wbVBgl/7GNuWfM4PyiTHg/jLq1OSuSCSCylGuXN3QFzTUFF4jkzco
NWm8C9lIv+RMzd2mLX9xDeHvA3txLjYW6RwQXJ2tpnr4B0XTYQSBdUIaDYyhGKZT
B1xa5E8LfJCZ89L3ufZ18Y/GyBGN9I7RcKNdp7cgGiCe+1VipnEJkWsb2BgsuFn6
aJOC5J2cOvpRd4oMS/BnCJUjeQHOn3RNM28howTdWa4Cw5wwKQpsn9/YB57RAh/G
oNruitzUd8O4zOs2Tc6OFYmHvGxyzvfsh7H36FwcCQGMGPL32S/UspTXKgvVEEbe
aoqhfpz+OJUaTYz5I1FZJmpYOL9xCif0no0rZOaIr/5+CcTswkwhDjlx/1boAdid
eKmRLY+AVpaaVBuJx/DPPy6h1MV9tUcwguZjXZBtFqahegVc+2LtKL9jsw4HEK4c
qidUqp4eNWqVGApmDQG+zY9HMOkU00yGZu2aMGqyfo8qQBSjyIgD8Tb/YyVmjLU1
oMwNZoEzOPGsKi1j/LACMqRD5UKjgCrSXIpcfHX6ccxGICoYkQXi3e3BD+v7fTA0
qgg7QIlbM65gwVYp8TQ1IhKllciDLaFNNE5dY8CE+L6j35bG+K0a7QEc9aBDkJrM
ILAJSv3kJiEsbN8LsJZlJ64R7W+0WDA0HTL7zoH/eEOs0Ygrx51DpHXMnzq9ZDUx
+NCe2b49w2SVul0BqLL8aJ8VER0GE81jBgqG6Rf5EABI5pR+eCevvvh3V3frAzdU
H3NzuQRoqW7/TIwhJCmY9eHhKKKgzvHrocOig0rlzBwihQron7HDhIJsCSGJuhai
z3QgjFlxOvTxdcix2bWCl/OcEFHIPMPzjGsp98tcBQ3dKAxvHHuAWikXBuFhbCni
vvX6JwisOUByhaNkLBWxctjnIpBwkRHpagvvraaIqp5uqt093zTR4ca7F7RIMRDd
CLxVgP4iIKwyy/HeQWemBBftTkDGTNMhzMiqysb5SOA0H4f/MWjKgltsR5rWqlHy
a0GFLJGVg8eDmK6htBBCW+FUQVzf4ozyVgY9rEKbChjRUF33uci0cAgnPPJLZ4pH
ChjMu56r1c3ri7CeOQv/M3SWHUEAveq+pJP4gJ2s3YEqaFTEzy8QXck7cfvtQxkQ
8nhCxHL1R+W2VQpFbVQAc+O1eq8YL5TeAhrICIRSoAlRomJz/NNOJLTvUrDKmthZ
L+R+ud0VbS32hV/9NI+RyWUROgTuqCpahf7NbgWipbV04rZ0Gr1vci41AFdW9/Ks
pxjBPDB9W3ZhePsjK7nPOPXxRQFFHW0rwZ59IslF3klQjbVs9vW0xotl6Jj6GlkS
QmJdWcPy4xccA+wC3jT0ndIx1TrCx6fyL5z8yOaJV0d3rbIwjNAXHc2jjvApjbLy
mTODFJyZZOlxAaVytGt/ajtcds2fu0tlDmvs1rn5kHe81LWZmAm7xuZTzQb24UdV
vmWRl7R6RMLx1D5gDd19DdUMlSv/VREEkJVfGqiujpBbwokVI8w4mdHXc1UJtUGT
pUmrnoaouLH7neuxaEP7iLxzCuuSBYfZ/uCCDg0EsIwaLa+zhZECDHlnAxZOusNG
0phhP5w56BFPnDZMUqn8TdAj6oR84QRaT8/XfEW0pLK4MmeJHPuPzvysKAilAzmf
xsf4Vx5d+yDLQQfVOsUKAsUk8dh+8VnjxckqFqGupNmjeLFbvwGpGnam0Fgirmlm
vjabdGkqN89J6A0y8VnK4ziu934kEXI/pwC7+FuUp0j2jjsm5TbbSHO+Ty5ZAZwS
7vbaMZQnT5ADkTvg8FTvEcE6W6PBF71HwsojW1DoTmY1SfyUqlukHCweDO2NObv9
PEeowYTNAsrvaS6efVHcA9h6W9ar+29gUZSfpMM7v/eZc/j1yPcAGDTQR8F71HKO
bHyjHls7yErsKkp29PU4d9NpIaqjzWA96i0xfJ+Jielt26ivi7QpGZqrU9yPM4CL
SwHiNtmtgql74NchkV7jHxkmVDuJqhdZeFe56XvSRNHytzUGL7DYZ3F3JqD+BVfH
WxP2w5VP1PLDPNoubaDaGYpfiRSkyfJhwrzLNEak1jKvw/bHb7NSwQjszNO+5HHg
6m0CGw/Ot6Cd5BQFkdhuw5fZciU8unjEFIYyDDYylg5YmiZr1vEsvWL+9fB4VHrE
AQegx2rWqt9XswERMucdh6NTxxe4lXel5AOMeIGDboaO1MbZKaH0SSOCIwvK22Ys
0lpic82XesUeWavTRRkJbChaG8fK9sqt53EIJk/3o7aiRoqhMngmZvPsZ3Fb9491
p8unTcue1+OlD/A5HybCMUZd4hMapxD8+sYKy6b+ucQ/4Ju1SQIPQlcZvr8nuOCE
SeyEY3xY7/PtrKvM++PH3yUxw3w//vKxNdwnx4pGsOywdf8s/mrAV/d+3nWX0xzu
rEPL9lKF6JWBGIW891Tg5k5xqmaJGt1PNLR7W8PJlvJDY+Gr0vRC0vYO+7EipWhT
+TUC3/k/fM5FBRmtFXLdxH9U4JFPRC58/9/VeRpkkAYnYbiqHQHMZaZKZy6M5t5M
rXrtDqdXH9bcrTVO1LA90+UxJK7c6Rnzp9nD3BqfSNvoCxlKTiaKLf7AOzDp87Xv
JYcMMxAUEGfGMHWNuB9AyWJVQ/MbJNl3uHimjD0268Pz/OrWKj5Q1QFILdQddj6n
I0hXjgdbZwkYLcoHk6KLJOBdzsgMJQhd49Vg+eYVU8VbrxvQtpMNhvdv91hZgU+b
K4/KRxLof0L+1LGcdn4Z/tshds45tiZVlBf6/97ei/6Zsg5z+9v+HXBQahOSA6Gh
x1t/e5w07ZXvzDHUG2Hu4f3rFSytX7mYb6PBnJUyOjmvL8iPmnrv97hk52nLi4Mx
qqyYcqcxjIYv59mRGdqJi1/A6HA1TuWP/SnbTBIcjZQXHqv9bf2PmOFCHHgnj3t3
OTTmhPLHfwiodoWu3EjbJ4gKhoJj4LHRK3G/VhhGaXrGrse7+5C3JwlxC0vt+j6O
1xXlgMNlA+h/ygdBOhPwIqFVSjQ9ewtUvpG8N8LzPVDZwjByx/sxYyw0m33ZelXV
eS0Vg8cffpohW1RTAM29B3gUmBcniPzWKUd85ugMkbRysE5ElVb9cQj3Y7CJC1mt
efTQCPoqd1WRdMLdfCx+zOnHs9hHhTzW+ciMDhvfkpTcyHWr6fYYheRhlmg+OMWV
AsbOpTrVNYO5RoHPsv/8ePgUAVbmj46nNTCyvLl9LKq3uVxtxEmvQKo1ukrBwX5h
c77Y8LpxRemTSauMRduTiU+2BV4NRyddYeJMKt+hLAPu036U7HxLZuIYE49xR+eJ
0IFuA6En6ynJIVI7XJyksHOI8c6Cd5NPy+T9x0bHapts5kpt3IxVhrIeGy5W+GSx
2D/sbCBq235JJrAoPPi8J3IyRyrfoETKtyytjVUu9CaQvwCekITgGJJfsl916lTU
7HK0dMeFz9+1JvYfFraZN6MaofI3neKolXmPqs4FgGukjmMJV6oE32ooRQaE5Qii
JeUghWGeZCnOaR6F9qjGgqaTBg6GxWRV1jZB2E0udI6YB614TXfDmsrRpRs2NZAQ
9KdNoN52e3ahDVEVyTPQ0FhXl77l5+7wqy/AkpG+vdK5G7HHtjyqhL9Pw6huTqPN
vXodVf0tmjeONQC27Udw2X10+tM4Ya6TyNLhWy4MzA3FefbNlWUNfIny7ZB77oti
Nv4KZSZuUcNg+3mGD5uQIyteVAyqOddF0YeJN/51jhPhKDNJEpWVdNDJ+5drZ/tM
Nq4YJsG34OmQzHMH7fH54ZRugg8x6gGgnVboBmLa5ywcDMSlUqL9RK+dxL32sd0i
aehpmdRNrUTbAc1RZiiEocH7SPhYklKn6syl7ZlN56re45j3c60nEBCZoehfrVoZ
Qm+Ro20ijOmD6CkcqQT12y/duGWx07K8cx7ICMTDJFH7v/mJp11vajHU5wws2sle
TDHKajpzIluUVYenZTroaZ362Dlohe7SZ+K+NQjymNKWz1IQLbpPnZFKuVwsZSl/
8UjAyLCG0t6ewLOsth1Afow4oXHUFIaxk9+cnDza7IDdJd6gH7ISJsE2EB2i6Vtd
ICzcC+snatkFC25N4QkPC9npp0NSnvd0NJa3tIiplHNydFcpfy3A4kwiy/y13jQ7
T21d2AGlbYZAeWTTnXMvgfzh3iIeq1gAUb+MGuMNIlkxVSxU2SoFhZdGB8x3nG6B
mV32d2wZoobm9zAcixfVqnMPK3SOPRp3qb4uGaD526ryap4dlzNrOOdLIPxZ924v
rx5n1w+5rrNP+YxMbQQS63RVWGU2cq9MOBEuA1mCPPsn87vv43L17bcvuerjam1K
fUKhsFjAl5RIbrDvXZDBrDceVv137VX7Rk3XvGO16VyOhP6aqlsXbffMI481XdXx
bNxZYsJTpVvvNt0fsF6FMqcVwhWYJTW1TD0+IE/dhB4vGEwydAyOVApAKKO2PdCt
Gp2SgBtcm+LUGPJRpe60BtJe+f5bsEnNo3dPWKsNA0j6IuFY+wcRTnQn9MaO/ckh
5HCTsW8h8k58cYMtz7GuvUZLUClbttBC8uU5DKKI1eZPbVq80icH1ogZULPTeg7k
UftMo3bcAcuk/mFY92am3qgVGX98cbC32hz5CzYf7T/KzGJF9F2f74TlRIIIgOM3
QrVLdFEsbFvgj609m9FZMkYSDsgM0MRLiMrNl3XufvHh1woxi8iWMFpHB5KoHPfB
N7B+tGgZtD3HKiRth4nHBtwpdFms/qmxprx9M9NTfpAP1Ys2s3iUjtdcouU5Ff/b
PAWdB1550Qguh5SZ4VA30jJ8aVEhaQrq0c1xgo5INBxW4+jrUn+NTsOq9HsNvY47
tiBd7dk7GU8Cdz8z/NEnL8zDjlgNcmsZqmC4AdSlxAv706owECHV/I8H2d8uW2v2
OzBnBjiOE6adzrS5BpPsQLMIpTC8+Ph/BCDgz0HB1qjbBIvXD/y0C+i/QNAEtRG6
RNwq0npv+12wjWFg/TATXFvtaqJMlEfg22reF+GPrpprRWtXm9zz/8MRpgHwnnnM
+OBZoxF7L8XlGBMoXEBC3K7cpkDo9rjKYTngGD8nLdntDo814vAuQzZjJ8R3VRdu
5uD5K23H9EIPcgt+TOFcjQ/xBLqvloA8EEzJPqqyIakQbne1i+P8qEGAlu2a1GAY
+fSWaS8T0ExRdt+PUbFgwf1JoUw3K3CnOiODMM8L7w7fG2qh3xJUg537ByAsAclp
54AkIABVQhxzgwRZSk0N6UAW4ttrzhVPa4yWnX2eQDjiFIuVxoCS/Hf2PjbAMCAS
gGUPyjoxfS1XULSMjhmUW2OvpJqWdFfU3gLVn/J2fT3vzDtTLTrDvE0sI4xHHeqK
pW9vpnFoyQEgLVmIGTyiorBOC0YRZk3cjkyjHv/Zacxolq1rsaIxJ2j9msoE9jHw
AfqORK+w6nCcTPbqTjpBs3nxUAQWEIFWfdKL98Dpg5qwd+PgWqrJYGK3f7HBo8tB
KW5kwwEQgX6kpj8LRar4q7W3qxVpPI7oKD0/y7HbCrDhG01T4POXY+iTEkyKb6Jb
NhJvjVaAs5v2SUY1LTbXvR82KGUA08eyegF5Ac2gi5T+1GnCdNMxDwXCmaQYPqmq
QIgF9FBtdDWRVQlFvOTJorYGGkgLkl9gjsbPNi6oTf+MD/PGQU82jUfWlmVI6R1r
yrouzityisr+tMCAkdaXCY34CebkJ+PqxFKN0DZI4rgdNhPSya89yZYvRlMq+xDb
F7Cf2HDv3PWVTgUhS1YvIUonYuBu3IjgXxdhJwSohtz+P12XE7IvtKyPHamRwgLM
ZAkonlCqIg/ZAp6VsUmQ2GEgHRDgHC6WPZt6uYtdgEnKpEVOftl7CG2EvuhKnX/T
QYBfl1m4zrd3eILCwR/CJscPPUgq17X/g2AjOSgU1rFp3EG34PJZ+Z+CkpcLuYnv
OXagwxzAPMYhoPU9/IiJRAjSrgr/gJnZArd7l6rQjNbk2PvGfEUBGtjr/4AF4beb
ilmkKnCF0HcVQHcu+21Qw1JzOwXzbh5Fdz7MXsbUL7DiHDNxfouIRUhnNx9XCHKc
njdmOM4cfb2eDZ3UWSSZGz3Xf5OSV7Qy5hFUFnf0mFvO7+iHlvLXqVozUaQ22dCe
NtqtUrVZxIAUSS/nZV9+3q2DptV6EN8tQuTQl7FNr0Fisb8OjbyWV44Sz6LLIc1b
AHYgmRPtmGxKwxiSS5qmV51OaBrDHQ/l3l+25oIjlbs+zUBbBOkoOY3R7roiQAYB
8W6HNt9Y82e1t4yz3OWfnjPSfRAfiZDTxfRDQ5f0W1R6vGHPHencNFIFZvergVK0
L2NvIk/SEJLDNSghbq3ICRhJAGShDg3DXINHfzu2FACpHfkqju2i+xZvwovNc0+u
tc//ANGoaHqSKBZLYN0Q22DLLA4LPAoJFksqlvTvhEXRfovhRVYzhb3pW0+zy2tr
0440J7p6K9JBgwHj3WVZdZc8utTbU27My4WjQp+vmDsmjtO3FqwX1iG7u+ZXi0AJ
cVng4LDQal1P10rgRUirLMwxtC+UrUA7UZV1GgCFt/BV/EQQmGbENpB+V5zLl1B6
0P32De5iV625QHKB6egc8fNZnEKGscvLhVUsn5F1QED68GjMA96fH4tndrT0XxoB
cKb4FxhFroNpPStsz+33MnWMVz/GEmbgAslJtohtIKP3+VN6L1uRRR2WFkHo+7AI
gQ94EdIJNeghl20fYp5zk+uGA6tgkkbmkWK5on9lcX8lKpSQ3M5e/LvUbVR6sc/e
ocuUuperem8qenMJa2EBBuEkLPgKQlPqzJhXMtlh7bcUov+2yVWiVgH1fd+CNPq5
gN1RvnUqlmkOT2bgfh+mB6m5uS2ELALai5xCywow6ieN1HghuSTOrGlG8ut7ipbT
BU43B0D0kCN0dJ6Fj/s2aUrCGEkqWlbwge4sT/vo/V9bv5mGYwa2qDlDUAca0n3O
E/bBEC2ThknlpQewXLNGQbxl0QgU6v/cu385fBRNsVhyTE2f2fRSRRGiAXM4AnEo
GFgGH52VRIBdv3oG1zJETbP0Psc/Z5Wh0jEtTgK96rusBnL+N2QqGbFJV5v9Wav2
GduCzSBIqlI4GeMp8rFj0UriRwkLpv42fvpqGZWYOHkN70ypVqHTQyEyDXI+s4tO
pUIAIJg3U3u9t0H1Cye0UN0Gas0ukud+WP1fQDEgpXkxe6jA2KjDkDVf+Rb/bAvm
P/5zqhgc1rshdZ+Snpof8Rt8JF+8pyBuVLHTZOnaddM8VbelJAt/N0I5jdvG6me7
TRq3EvSWjZphFG7lp1dZHxn0HNAJKXDAIN0Y/lQXJjuwB+qFD2goL1GN9tlQucE+
IredtR1sZdESDJttML2As0RB3Dyb2+oaauPGUi7V5maONPgFCSsde0zvs/s/iZK8
CYX4JxeGP4Gnth7VWxOazjZFY4sh9iVS06BQsg2NTIuvbCm9tSNSGjsM8ITddavA
1qKOGKglQc+bLRHbuFVSm0bNKE2ZBfWlsCi8aMd8boUf+KF9RvJvfZ3GN3y2458t
3V5KrfyQJL6t6WiEkRvfgIXkOF/8ea69BY7Z96Hoa6mIRS/dcapxdXUWRo7uxwd0
vj9qklXjT0pfxa8uVtrBuTkt90BOjfYoZT/SJVtIZUB7d3DwUmWVdhpfviOMuhmB
4t9UBjTL5eeuAr65bmSpViyxNx/77mIfrncoJMxrJNIS6Xl9Lklm5RoeQbIvWBP6
uLkE19c651SfDtO/Aq1ezN6ug0hPqF8HFsuYNgJ3gajAnwuEVofBhJBo8+LxE1ZS
kXKf9j9MyBlL2m42i8FjqW2Dgeaxm9dJ56C7HB6WWHHAHCieMD6BxCrGXFYQbvj/
GGdYkcdOOcS+HNaE4M4SpHMP2POO4/NBBS/FcH2RHKP8mAzA2qTDV9gKeWlc+1VO
TqOGE9gUHsAk9S2cLm82HyuSK2shj3eDLe6cNTa2CZrJuNVDjJtLTFjXMLBl1oQL
HWPVn6836wdOwKQjUuofe8nnq90jCmU2GMGoaYVxs0tYpPna8H1BkAKzlXcqakIq
o9Q7hBCHPndeYqSxQWe0Rk+G+Paegabw09d/f51spWxNaEPffbqC8xQP0tjHFz7Z
zzlrAq7DKN2BVY8DucsouJmwFDT9ei68o58e8up7g4GooAOD7wKz715JyvS9Bl7f
wa35Mqkc7EofFuWid3urOaLdqOb9R66NVBMkaW1FQ1jFdBu0CjjQRWb3i162PoHK
jmX3GBsjn1sbJc0OBd+l0YN1JsvHoRY4qLYS/J60Kj5MzxisK8CsBIRcwBvuH1f+
0HVy+/qINY2rthu1gfPLTVMBxNyOxcmCn5po6vauJapU6cJyL3o8zwXhdP6uXS7U
ScwH0oVrE0VizwnM6fC6S6j7eeevLIdFxA8rG6XzKrdoffW7FvojdIUJA+gz5J43
VW0l/sf3upYwuKSqgVIo4EjAwEaD027imGnrK38l7AIN5JnJVCRVfTtHxglHQZsN
xSl4GBAZLamKsCA25gElU54isJsIgCaXjWkX7EapFLmWDEEiqOS4Ij7M1XQBoWgJ
aICvSEjprHlOlNgreN7VSKinlCKPJjUdbdVnQzi3b/622IL+crVimTe3e5+dGCH0
NkTCCuhpMiunhvKgxNNDHKhCb4QD9YBA5o0U1HUfO/3mPQ6Iu7LUhzoPBvmxFdnv
4WpJFWjipEBQhaZwWBygayDiZxMSHv7CG80SVXY1l2pi5s/c+jYLojDq+UNHzpe1
xIAxlwMbyfPduW8eUZgYGHU0hK8LP2Tz6D9zie3TScM9HJOgm5wrYmtJmiBKMAtl
dhn25oyPQCti7hB/itkOsh6zInS0tI0X1w79z96cMqpTA7AzF1Gr4z2BPluxsiNh
TqP9k3w4SN3f1r+cQwBf2ZJRiuu2Q7DLHVgWzPmdhIVaCrNioz1exikPWkNoukS6
5VJK8ZieoxBv5CGjoq0JUBsAKJ4An2XkXclSsVUP/Y4MfqQqj9RLZNXqEiD2SXWg
f8T/n5V5B8T4fmw0Gl5WpDg8gziTJmlM5jQuedHrvH5bKIFIqzXl47sZsCG+iyVd
GTD7mnpEOJa+oEr258HAsFbCMnaon995wlQB+2vZhFpssnERn0pjoc49Lr7cx7m/
5wZLKKjLDn1ULrEXv7wWmmfKdq9YxnxiOUMcwhQgYCPVoTMvfOMhDn6HK3w6pqpk
1H2cQsZKOb9zuETs7nE2DXE23EwV5DXszJk3jmsVGj3iyen5t7Ldc82Zq6ewI+2j
rDbnj9YcB/oVF5UvV7KKUHGbkRTOiu3u+82BmRnB7ZVF2152aTe73lN2HpoweW70
nHwa8IrhV/ZQCRADIm6+PF/CAnAQ6AX258FI4D/XzE8Lv/stUtTMu4swMgpvRJGL
4XQ/kYGPwq/9CNuY4OwM+vBa9OTrbVpFqP4+68JbjU3TIvsuFVL9UctgVPAbUgeu
K2q3/jgqj8OXL5n4O5e7Wr0+VzeEvVTYQ0RQvt0l/38C7POagELHB5fNMSItaSQb
RCF129H/+MkKKqSBDoFzHFsf3IsE+axm5Hi/rC+hrIwMN91MD0vP+rJT5gHbOmgL
YyAXDfPqxDuc1ZoLou3yHntUrnczSXOJY3PUIoQe/KLRtjFF8aidJxTu7qa1ElQQ
WG31JfuxAPlnppY7co6tYgTkDgFIARFSm2jbwbyHeh33UIlZcwKetcRQvgeSKr8p
JkAtIvpn0kC3kvLGHmyAqzG1sCoOWTSEMAhCh+WY6Mg1kbiXzyEIzubBurNJ/r+i
ldE9xnp9Qjguf/jG/oLLgpPAyJO61xMFgjrfonQXpFEWfKzsXVl0mtMm4pzvOTqA
wLjF+p1ciAp+6cktOXasSBfnFghevSSlh9tYhbBXI0ZCqrkgYPdpLl64pFVgwvmN
n/hzaqrTPMXBaI47ahd96/mnseE3xgTbtgNec95vwdGWToN/yAl3irCHgwMy42qy
Ssu8VJeRR+r9SmkdmMmndtx65dpjqbLUU4JxuMCQRTzMDCOrAxStbBrZ6QObSGzu
LwsOtcUEJ8r4Yk1b6kKE0++TnFf9kQUnc8ndDhejl8+e8Od26m5tmmR7lxtQVRF9
1SderrcfG3cVvVGB+0EmS+p4l/9HlO3h0us1pgI0gNr8Rqbp00tnC5gu+L2rFOzF
COB0RN6nKa9b2VncmP6LIR0Y6p2A7GzrUXQDC2bQpAXipD1dO5Odhbwt3TTm1K28
TmF2cUoBtLBHB/EURRjwXGcqJm1mQZKFjqBwC6LM6yxzrUiiuoUxhsC+sYFsX23a
M8DW4XlqqzT0ViJws/cQPpa/UMZ3ov3Tot3FPak9nN/20qzXpdW99BI9pcQZddb1
zvQoPfMiqOLmpnpn3wKM4fkHVxSoSziSvNNjg4jXUlw7AYe1X97OgFFHQBRpfYRk
qTpG3dYhzP4P+D2UdTRHHLbWvNsnmmvWcT61mBtK8Y+TKflKUdRq8mV8T60g1/Xy
cVT/04yiNKnUClW8a0gXfRanEcWufC+uEDUHefqkAltoeZmh5Q4QOekCEfcfVJdg
lsRNHBK6kchYL8BGrfTopE6u3QyNbV2jB3NAYcQkqkLM2/we50ocK+64YL4C7J+k
ClihnVV8FM4wEpWk7DphtOlmz0t5v72pIEYrKgBy2NEDWDZtY7UX/6dYxwFy7Biy
9mdfUoBY243aNJu9oAPwoQ5SkdupIhNLX2/CglAmhqD82ZkjxR7b3uYh1El26dgu
Hu5e/yeis0/kobVMrOULqcoYeeL3iFrm9WeZiAANEFnyvt7PkalE3tGXbjjIDfdm
D+V5VFOMg+EkImMeaYBaXsYQgogvhdTnsUxkjnPKUQ3vaRUQclZ29lsiFAbfB3pE
rDW4OeUVmC3Fx0djlr9eUlBVGF4Sx+Wk/x1h/BXUFk1pS3PIGtLEZvgGFWH8o3t+
aJkt7RnDBNVn6R5T3DFRH2gskmDlR+b3MV+4A+f6WEgBvdqtg4E9fh4cDhimfFWZ
tw10dYn6rC6ZwSycO/c7kupkXzwUW/ZxuVKu8N9ouOUFDkdBSCl5d9aWb5sZIV3E
yf0S4aeww00BPnd6Q5z/PRjtcIsf0U43dH3UjPXbS6Nemm1WNyzKzZKMRpf91iB8
nzadV2sl4IuM08DCAQ94OqNLOQvT5WgdHyV4ZHh/x54jbYg8ioDhCxkfcBG/8LV2
AKAhdfUjAtiKa8stGYqGrpeMTvVNaoMMS7YwYfz3qnBBbHXr2bgaghyJgL+Bu9VX
kG4SYuMl3W3TN4FesV9Pr/Mxy1PbXbzvUZbuBzd2kDdfmGoHOw8StAEQtDQ9e5UN
gdOX6c9WJMrIHL/nKWYWF+EvVswY0yNhe/UBVDVETJqYB//q3Z/6uBaiKuf0zVU5
DMey7rN9alfOBVXSAxe9Nv6lVAgb2dZSoTMgGrZhVfBrJ4oGSG+9zezTtp82iBm6
Oefnn0teMTlOLdQj+Y8/T8U9K1XovanteomfQW3dNoI80SSqz7aSOZaOTiHoHPwQ
I7aAGWwqlZrZkt+KnKPnBXfDPUOQrRe53nBlSKS1nKzl3HC6jiqu/TqDB30vSiEh
1KS5uoh13VlwyFzhEjCPSsYmtVT5q/vIaQbP/1mO3Ee+PpK7cpQgBBKP4fKjl2/p
oUOXm7/cjcg5ZLswlxzzpqPiktYFKDdcWC/dkZdGeE7K3NhqpJFCowSDuAGfPWe+
xkF8rgz5SGGK+zCJ+FSMJo0RuQ10hupKgKXuNaKZTb7/WQ2CfcICUYblNBl7Szn9
0ez0unuyv1A0SiTGmI8kld2mkXPXuZ27NUlIaugkjHsn993vB+xJaenvnk9VMyo+
GrhYhZjNkQ7zOTNoU/ZVIqkTsSUxuWvBC6mxniea+RZzzDN+cm0V0FLjASsxgQ4I
z/u+EWr5tzkrCXkqGAbFwv7p4Yoys7PCIyKJlm0MU3FLlsHD+nnhuHg8mJAgxUaj
S0PXX286BrwKxM7voUtgoMLCTjfhQy1Ch4xFNFI1kPYNuIjWmjeVoy6sxQ38XwoV
URehgt11RX/uOZhVjkvcysHPd0xUUnjk8umFNw2DM7xMEZcWLmB1q3patmm9OYp4
4F+T6yhV47j9pEeLtLWqq2s7zt/ITibg4VvC2j3JrU0hPqctuyfeUXBma9xPArHv
btvFTTHk4asggRUEtGodL7t8/ukLNOf+tZu2zlUr61lg+mBvf7kNY1ryNLYXA8mu
ZQjb5hnhA1MT56iQ4JDRGsg2EBGjXgP9jq53n3FAu/MAqbcirY7Yp5K8VJfXCyzW
IP0zVmbI0mIVik76EApNHe7CwfF1ZI4Q12d/WcPKdrjcSOXoBRfHOqEPzWfiTGc3
MsQZf1s4O1Pz31iVWZMQgL9c8ta+1U3Bk2oYFOuXh31ko1xNHLzBHqmOJdwCKzuE
CiGU1AOllopBGNXf9CkFwRSNjc8IdTX2EcIyFQ2KBkB24WakxEz1i9jpmFk1C0uj
NU5mhAKnyuAvifQA/H2RQJek6fsNZnoPg9Tc6PuZjl22gVQCWU+gUTa8toA9NhF5
0MZbRPNhjrO+mcjArnCk2oTFRO1Tm1fkV48kBVAneEoQCfJv7RbYbbdHbjBGChNk
REiX92FocknELGOZTOQL8vNuhGsZ9YmMmPmm5GcY06QfKJgjmNR9DhADxrZ8OclI
zHYHg/EVwCBEjrR7rQhKQcUSP0yPto5oJ3kZHHln32G+ON7W1Dnc6gbct/6xzgQo
LFIkQYhYMOWnU4fX81oS25TWQ/zK04W/wqHsCSQujP4nfPZUti0qTdFECrM4cEMU
jIlt1WxtuhUqYMZ1gDZrcNenxtRo4cutucyS5Jv7EGzNdF2pkAi1TxQa8MCuuCz8
pWWjWo1wNa7arWbS7rijGkm+E2Kjvuj7VBF1LLA0zhiU8cQVtPOmZ48zwGb4H6bo
c9QZjrQvjtzuzfn1W2bVPee9+RyoSz0ERtfChRE/XL/MyecPQqiuNFtGQ9X6+fib
WjFDCoSU7fknzQR2w3yPp5thQQP8Vuwrc7D3PGqDwX1cnt8MrjOezi6qQCf0FPvf
6bVm+7RCaA1ijYRo21a3nVknMmA6V0nRqqbTjANcpB12GRGDY7AnYqPD5GupJqj2
vt70du4Q7p9kt+af6HCNx+5mM6kUxO0xjAvkhUjpSfBSTXS4BzFwoctoojATezOW
YlDZxpi0rRSkwsNWpDASqGrqtEyxCmDfl80l9YmecyDz1Fg9r6Gyr376CejGlUcE
HJlCJBEnqV0lt3sBquXAYc9V5sgSlyy3+dMaTOhFv1ZVh1XGLlkiBj9vM9GCsI/I
XcHDiHJ4dJ0tzNBvpjyJHi4/HFOoyEl1YPWayE+8wW2BCQuOTzSCB80iVfOf+oAT
iknrRM7K0UrFcYDAnEC+gfR0ZJRNOrHe6zLv4rRfKRzgEAdMnKUI0pea1NZjh6Uk
oI6mUWCl63UVspuKS6+9pclEnr2kdKY1UBYPapOiLEMudhFCVamkzbRcgoAjKYWT
xIOi053nT6nSKI9KRRhQihaL0vuE+X4iPuIIi9V/PFKVvFVVjo3xKiTJE6SEj0nr
fM7zXmju+53H0u8QhHl/AtgARuoijcpxWM1uxNxHNXEKwc+m5psS/ebI6vQ+7MMl
mJZ4/6Hu5qjP0eBp3yQ9d2rKogEmjyUzhWdEWLf/5oiQSXt4Ggm9gtii9nCNQtgL
WpGS2x4fYahRFnDpHcz65A3I/8aHdqlA4M5YZNG/NLL01TbGkWAsTDYD+KVF7Ofy
+jXuNGoF7YQBDYhin7KlYgLBXA4higFNnqUH0BNeHD5qwAfV4vL29bDlHMcjapKn
IlNqViBF//b3iXA57Rxqak3BUaNWBwqEDyKOjGiXMcT0rvillrOmOUot8prwXOob
r9DLJE6SO9lrH+k1Fa8dLScP6ttXTGzalJE5L3Ocn3jJ86yUTWwDCtQnNF9ybe2M
yCrRsXdXxKJKBUpRER+nA/FMLlB99O9Zm1G6c1pnVku0zysYYrjUyp5nkZ1q2Xbj
L3AZsSfkaukbUjns2Q0lzXNKLtuNXM+4tnKxKbJyCbSkGgvWB37w/sZFJYmW6Y9T
kdVc/2QL4VghWq8pyqnDceXD1t020qnHzkCON2t++tkQ9ILEC9QIFs2EDVlNOfz4
mRpiZUnn1yQMnBvq8lxpIT+Pr37ewbSnyfIR00+yZK+EexWFF5s+dQ3oDHqq80b0
s51s87oZIXxfwgOtAPHuYDRozDijmvbxkBab6mvRk1qhy41UqYcQ3F02CtZV8B7o
rjvha1rUKn74/eUH7yzqSJisdZZAXn99/9zxTmQP8PJUZpQsp7PBS1jEjODyqf2X
XvbtMHGtsM0ZDvlrwQJI9iWSQfuIZ3YcbKeZ/UgfCLHhmfRRdpPJvypdF/wQrU3Z
IpNkZF7Oo24zFg1uRAbo00Xg2KtnNl3MgbhIn8r7QxiQZAZXDWu6dCAmV5XbIIma
MufFCLpbPyURfEKktTkUXBKDOzrZgH6EBiOBQTTYgh9RPTTTj6/JYgJ7V3XYOr/F
KBIyli5ADA+ncCeF+hl1wYIa+nqXg/4c0NEhkBwM36+Pt9lcuiSNOPabOUJG+wFs
Y78zAGJw0s0qC3U2fh1Ov0HAcRUDbKI1tvs/hylQHQOJOw7rU/XhRvwjhxyIugJj
bSniyU64uIlelzba14aMBvOsgYBXvEXdbKLtOqklEElg6IajW/D0gwBKn004JVIQ
N38aP9W+JakPVEq0dS0yzAwrhaGhBeOmCOLe7XnTo38eSZIJWpnoZpwGbzuATBX/
s9GD+fZYITPixM18FDGbjqfh1erjpE2vd27+XwfqU+r9La/Ab5CnKa7mnqMuTHK7
ubkKmxV8wP13FVKaxk9tlpJ0mcnaItkI2YcqbmL14tNxluMucChFH5PlsAQzNrIA
4qo5AUw1rlHcB2y+UXeUL38wAged6fdzKAKy8W69+xkhMhrm8crM2z0IPe3XVrVY
8PkROWnCJxAIVGIft0Dc1H+2P4QX2uVvAbYBvkMbVYjdPCD5H6+Z5B+DVNGAwver
wZU99LsvdYYktJ9mlglNPDMozt3iknbUK9S7V5YpCWIpuKILFDmhpU3p4fy6IamK
yiADpuvzCw5fkfJELeh9gFQgk5pMXWLWny4zwU464zrS09PXCSAPf2ugeIHxFOB7
Z7L6VBrUxzPsXNO0bRaKMrG0XsTxeSdUAe5TQw57MY1eq4QiCyB1GUn+DsyHZApA
uP6zJtcPCINyISOqrFa7x4AnlDWd/0Fki0CEvn7yah2CsF2qDA9GykVII+QkMPAI
ESyZdQpMgcuD7Rb3fufcKXNhVxTA1Pu9Anb9rEs6TLaNe6Ed+AV+A8uhoH0i+goT
TTQwzkK6g+MZ+98Ui/It2Wv+6n4cH5VLSNk7H4uWpveZa5mvz+z5Fjpgp4uqUncS
AB4JpWAwwXoa9/gGhc1/tTd4FXVV8VJAO2T1ChBGreJXMcR12jwHD3aMyYYEPA7V
C7pdaZN6mEWm4dEVTRpgugPoW5Yqdt0DtA9ZoJfAqb6/YX4f/tQBNrvfhKQ0zK34
V36j4kftL0y/rQDRtkjPxAGESulXJZMYPdtKD21FloVdI1dY6C/7oVU90RAkFZK5
BxxTG6KTX9uIOfvSUhgB7kU1cjnMwHU7SrEoFW+9DRJjEGXgtNFcUYmL2lbh98Oj
XsJTwGhU2pJo0pYMJT/L9XR6efZvAVZdNICvlgOOwOGRVewC2KgPrxCM2MFON6Oq
SAOCUVAvEptn0aZYFiURmUyPfXunph9JzdbgFGfoJJRSTRFoMd0jhJ8lLzzF0vv2
xii+3f+rJsg78eqvBlkgr0tSaadExz/ecGgoPm0x6PalzxglBzTsWFamfUeMhohf
jhwxU8PYxNeISsgfV4El/lCET9SCt33EIBpN/46Ykw4GXT/+7F/BbqMHKkMahgKf
ZDHqSSvLD9M8JNWf+CGSJEL9+5giHygf7lcdbPRhEjiQEJHwEqLwZu2g8w2lMePj
zqdhQdCAY0lIX1BmCJI9gBC2byYnJH3iXUcRUctvKlw6xVthe4ChvUHD/jIwEGRJ
w9nmuYd0vmiBTPMV8s/T1OvPO9A/liiZidYLQPW+73CAI5/V+uUpS0Pr15KczuMA
gy9KdpW2WRQRcoQLRh4/QpLkv2QrDSZhADC4JTGf2aXfEVBn3IuLwFzZryBiINce
eegU5BrDkyAqWR5Qa8ugXeaU7HZtAWfcRSGDRUBYwzGcnd4W3dBNwH8l0mK79AS7
p7xsHdWX0SqMaHR7Op2impQfsYk0fFSjwGzzbNzu7cVXEbEQHKm9PT6YohXGoNFK
kKfTfz/bD3neHaUnTOcAZ/BKJFyFQL3bY1rA6py0xW4BA2h6DkLfsD0uNwl2au5H
Wk4kQ3soH0NdM3d8fwMuXiuiZOplGmRR/qP7NrJm9buXElykgrhSpNytr4ukGtxH
OAkn4p++6bi9Qjb25gumnI0EdPcf6Meys4mn4SBcL4QaJuXtcdJ2lvsuzV/W4bsH
o3AJ2+A2O18XvbpS0F4/HFnChnpRO3eLeqqj2KtqDr1YqH3qv/0+GJxy7QDEDbKZ
BC09aXkEV7y+al6Kl1UIdCWlfFHub3+2eV6Tdo+b9J2ItS6Z8PI6dil89MtxU9Ly
H+rwV9TlErev8sPk9a0D5+edbKBgB8EnawR7Ir466MLOLtYROX0Keg/1V4783zs6
bOK8020lXyciF6oTVIgn+RoUDJo5o38tc8dPMq/9yQQABE/ELeo0aEVtY0ady5Sa
Zh6Lwc/v7bz8UGS/CxIoob6X3+OGlBLVgpSbK2JS3WG8ueW6l3IXWYqkhqEmos6/
6sqbWqjUjStBHC/DHOPov6+dHEB0DR5aH7B1xx+N7p/x9s/AwuY4XjkhqD6wYYZn
/XdK2w8qiMsBpmP018MKImIqPuYpdmWAposXwsk+T3cGQzCFDME37ZjYLysFOV+o
OEuQAgVww0JOr7Rcjif2GUj2ONp49kLV3kakc4aZrGmWNuYWdJHHjAxeBUI1FZ6h
F2zJ9tRmcvereSp8Co0fRnRPLDgxbUPZUejfr+9F8gkxHKGMyhZzLLuOFot8AQY7
yyswpLzC/WQEdcRiUE+lMhR9RfMYU2bcwDRZL/e3gQ4aOsQRUJ5IJgjFatyGbLk+
R0XYNKuG8iBQtu5D4OaKX1GmCdrSul1wcA//CcgNfXAuqvhctETCkRU0KkgMONmZ
bngOVmJepYE64Cl5OL6DwI6Pe+9GRx9j7EB6WjsQkV2nB5n4e43lvzQO488QSDK9
MQ0X8Nn554hpWILiGJv2lQsXp0I7eXi4+e+f0Vwm1hIDrKC/6dpiSx2oyYtsUrwe
QmP+ehVpUfGUb6UiT15oD/UYuMWIw4T/iD1R6PwkYbHqTnaJHRfaMwBCnD/TQ+iI
HAawrzR0HixdqTMjwT20auD1h9TrpOAzf3WCiumGUIMbUZkHfk+e19slaquHLKOi
uVmbpf/X+uh8Naeed+V45k1Tfzr9n5Vb4B9yj4kggI2PArGBOayQbZ13R614K6Hg
tWPLfJN+lQMGedaxrsjOQYwB3KmJXvoVwO6rpnHGN0ivsdW0ORDrIaDrLl11DFXj
rap1jg8mPUTgOHBhxeiyLGEWFDV+zzwF8o6SJJolg9jTpGl/G7SynLj5J6dzrOHY
NR/HjJz6/9y7Oi/jz76H+M2s/gGVrLb1AJXT3mWnaBFWzXQd+iTKl5ISZ/IrI6rp
MbIBHS+Vb7Z4G+1XbIHW3O1vc4r642tyrHt6Wy0dmL+goJPx01YUBh/4BOB1kT8g
TR40TNmz0ssD5CbKDlwKoNbe1Bh87/pMqgK/6Yj2czZLSHaMehPaU5i2LBdQwZVJ
IixbIJln5EnObiAt6rhKECQlSZ3Uqw8Yym1bLbqFfnykOBsaoV0EFWfgGOjNuUM/
mUtDW9jhMK29vMFkUOnNMPgsF2rSplndd7M1RibJCq66zIfcanjuJBJUjMDAaAjt
7kD3eRSKvphwgJBFyo0RzIPGUhtjUrlVLWA6NE4KFJNQXqb0rw6KndyfLe67ARHt
4wZM0cXFErJyrfb4hZfFKFE0N2NK4DwazVV3g5327ckXrtf0PYZIV9bsQgdv1Drb
943OgI/QyHTJAWsxGWw9dK/0l1s7Kc1abaG6xXISHWfCJFzaMz0ZzWhUOT/D0myY
FmbNqAs9iNJ3Eqj8aX4gTxXJkwwIoSie41eEQ42ZuAsw2JF6J+D8nvqvNMeqhpQs
8wMKcl9Gz1hE0kXM6Hsfbkq8xBTjmPXdaG22nqDsgEZ/5a5D1/v5c4MaAUAoILOG
XX1sfl4r/PJb9p9i7lp/knihXsx3nEs5w0TGbGZFrMfywuwcTVhh+vnQrFxl2gSA
/WzMFxD3INOCKjdSo3HZOMnQg68gTinJtf4K4FxCW48biKnOL5ws76Es4Z6hwUYj
Rwh5wGCo9RPVkt0/cvZk4Dkm/ORL1npFuljUf81MI6nlBIU5YNSLCCdlERdTOj7I
ifq9pP366jdqKJAv4gpApbaIFY+yfY1E/Xli9cYa9P/AZ2K6envjnvyVTq29xlDl
s2ABJYv7aMm1zS4CfN/JebXuwA6GpVnpwh66pbs04SukwGU5XnqJs+NVb0vvVspe
jloe2qc3h2pHPbWv83flk5SPm7h0J0LgUAlRd3Du2xPTak5+jtvq+J0PMy1XYRuI
l1vP7rQsysjfL2jGB9zvMbJEkz+lReed4WQrnlBandmn35l2TDunj5PGq90EmD9t
MvCkrTSCaQReN3xy2y5F9lC+3rH5k0n2vnECfJGKRMW9JrAJQhil9u3P7GrjtOH7
4GH7Qg2JHMJYcZt0CFI0kGnglifookg9+KpSJz3aWPVVS5rslHhJW0JaSUlCVZCL
RFyK1UVntbtvxtOpxd2We+OLBJTR4Wnw/zn6H6O0m2iyuUMy2Pr81vXN0Hgxa9OB
kN1Z01pDH5EYTknSihOieycoTYL7KAPE0+c+iN+/2gPJd4NeI/QL335TewMEjNeD
o7zI4FU5Z0Ze94Gh37WO4k49lHPUA3Dwy4IOM5As7Fi5SPW1gXtYnQxWEuTE+zAg
rs4tzEY2gayruy3i3Zur5Nksn5sdeGn2Lnk0D6G2+XO9XWLiPHKzGSkErv5YxOX+
pOH2QqxQ1lKGUUy2H3sDLqGBMn/FMIakn3fw1R342NCZszRHj6JcLUKu02Z8QTb+
yHER69oJwMBsT/GMxbHt6eJjQEhKRNdjViYU8lCB6Qglpc1BwKEuZP8UY+bjA3P0
CvB9SxHbXHdbyG4fEIJ5jxUUA2suI/l4zXx8nuKSo7k1sKmy9C5OzhazidIIA0oL
NzycyW7cBAOT9BNJ1A/u7wcE9h2zBI9p9QwsSHFPFVY6mQSxVFTQVrxBCEfn1iHB
wk4T2wuC0PoCivHkLb1ajXi6zgxzhs0NeS62sV82CzKESpxNCMCwi2mNtjAgrxCI
JlFC4NpM4tu02g9Gxp13iufCGpwVaaNtkQoyIsZyEogw/qbEijIvukmigEx50KbV
5MjYjeCCIuxWRSFh81PssG38fCgbiIz1wf5qdx9FcPVKfo0GcXdSpImtfWjnFWlb
glX9qQ4rsEk8RIlwca2/HM9V2K2K/2uNmEuxymvnuuoDPiuySssFCMa76VQzI3Y2
WgS3GyZ5CMBnzQuOa1SndRkGRrWV/psWfamcr5ygvID/4FaOUo1ovklUfOXzwLEb
NDcYJO5YKHcj5mRWKGG7vck205WSllJ4C7Yj1HGPRy1GeS0vJYbq1xYSqa3oBmQo
DCBpDukaobsgWUseBPDHbuGmaWRZEGorCUC2yhucbtdzaFOGQkosoZVo1c9hQ0xh
eC2VAXQTL4h6WMJk0bEBRPPKhr3PbPlRErKr3Qdo1Xt/Ukm7x3gztS/wCagGMeH2
PRRvGm8Zp7LRV+PkzKasnHIceLEHMtPGumDOblNmLCVSZa+t7J0MOpGJp0dtv3nD
tdZPRHk81Iz7+qwhNLeiJkjzdYEiyx9/HhYrrqjLbr2GqppUlAiVGvBNhL1wTSME
+MA4Jo7ok03GBDpnjDwwpaQ+Ht5aV1DzbsCASjvei4X0mSbF35jw2UpTVFLe3HDk
hgl6UIP4kJlO8jzgAJsMrqVFBUGzogAbvwYfPeDCoxewUYsV2G377BucGrJ6FSpW
m6mieD97ujXl08AknqdaEqDkvGlwV46H3yKgFRNf0acTx4/dB/tY32wqbx2/bJ8T
Io6j5JAFmciFqPLrhyQKm00GdtyNd3q4u7vZUm/OELlXjVBYlwXQOhAAonAaeszL
bGQNuQyyJmi5YwbY/TKqS9EnHOKu5Ap14+/ipc/HG6cCmoatTeV5f9QvYtXMoUHd
Jne3t0P6F4wjdmNfrvs/NGm09Cm1W92ya3recAosM7I9GBMDPKqePxZa5HHnpM5R
KvqXbhUobH+bobOgRGavxDeu7Qv4SdEw/4c+yBDU8UIKYlp9dGPatDxJNG4pikLA
07Sp4bg4aEL2Cgv3f7oSg6Bqg9wdAtVSugBOiC0ZgTKcP647jpX1d72bPF7QdKTq
+9j7b4fZBfLfzfw5WEiVbz04Bos/YET/8RaETPnkIOYRkrJctdHfWstcFt/vE29o
W5pag/SEWhNPM9NlTaw+3yrkHeVzXeOnzr2lBnT0mIQWCn80/p/rzaviYn7RjB5U
g8LZy9IiP8AJf52YZ3MDIpDmxQPe5L8SIiWMkBnyOGsGvuUqL+TxNTczQqOv1doJ
HDnegMoYcVEaIdlFtOFyYX8DcBQ5Ndbnq9SxGICKeAchVL0uDuBCw7tZj7AQe1MA
SydhP8ok99+6jdU9b094LXsW4O690+gXoGKkpZ1wA2Mj/6lpQVZO/9xpjVprSpkg
VfNadqvbGY8YySiF608TPrP9Z4qyFZcyc+EsunkLC4niThaSFn4LJxwFaE2td534
dtTeQ96MYORtol12GRIj3tEfoP99MucE3dFo2lLuZgPqEvGput7azktzF3Yi2IPJ
gMaYBeVXMSFtpwv6MOOgajyvSXYcjZgrd7f/y71pZJOhQf4qgTGwfXZ8wDicEjV4
r3ZHwBuJnv8wS1u+IJavjaKzvnuTl59dsPwRSQWj8DBkNDGVf496ZBX5LN2byri0
jKKPkmNK+n06rgOp7d9qt/09zrI0OiRxAbA7hLstMNrOtWkM3LrPJYsXnoyhiGaT
bJ02Uzmy64FWnxLCvUYm7+RKdya87aiLgoRXRprze0B65XWUaw1XMtpKI/lAebeY
EJx2Kuin8EHKQWGIv38XgW/w1Ow65IzqRn5IdcMvwfrkQ+fJ8BKVxp9q8DbENyNO
TEpQHpsWsXPKtA3qXXNmNJy/dooqI5GbLoFY/bBt1t9VUov2lRdeCQCmVtpHccFK
EQdr//0PrrfakrAL9lRLVLPr80XuAlEHBkGG7ZH4gHBAMydNKgJ6gn8yT/5fDjHx
am/hIAZI86f/xA/mlIRoeBVWML2bdDGzZxSwxBATRDSbLdm4+kIyYCaPIEjq8wbS
OEHLWz14FPnTgTA8+bCIz9GZmg4ITK1TJsEtLZCZI8647zolW4oBfpdbF/SXOTQ6
dCi2afHWrguXFQ/8FFCAh4WnTREDdE45bPeJhcLy7aCiAitbeEEBMiTAvAihmWBG
kDIatInjQuqqVRlWZ2DUNcLDc5b2ce443eoS7xVBU80W7nr1BG9iBxnBqL5YgPPA
PRSjeja8ufoQqT6VQOHvDMHz1EYKG4aob2vM+DJsjeoybnI1CMZ24OUARJr8FMvj
O1x1aEkF5GBZOWoT+kWGQ+q3tgOENKM1F1CqTW3kKdNbSu/eXH3hKzvp8xxwnO0z
tlCIV9XeSByBqt5JxZEUWWYS10disfjtxysnva7BUIpNmY4O0uvyid2Sn7n4X5k8
7erTbOtVTVEaCelH0pA22ahst/I/d9EBVoYSWwH0vfV0eHcn4YIvKcfhCWbdJwu7
lulAhrTMGUtSHk6xo/TdXEJ7ylwvZC+qgZdlScrm7pYD6iZEoBpGvOpcoxZfyM26
`pragma protect end_protected
