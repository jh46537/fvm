��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK�Q���L�OX]B�Ј���}DO���!"$
0���l�Zy�@�Q�䎁�1�;7gF�%}�����Z���MI'l|&��Vߪ�^\�Q��EsGF��	�M�|��Ӗ���'��T5^�] ��S�3����':���gm���k�R�Fo�m����>S���xvS����#��T;"�4���ů���]�٭<?��߃�����Q�hw�y�|p���F�_�re^�i�������m�;<�1J\%`2�y"���
��:DN��x��m5���v]�f�VD�E�6�����1w�ſ�@�
5�2�:�n�� ���)v��4��Z'm)����u�2t3���;F�h~%dľv�X3�-iKg)����0N����J�̂#�ا��ӽ��{`�נ�<],��ޒ(�4L��%H��ؐ#�g���
�#�L����Q���Zu����<��틀΃hfW<�WQ�;~�w���jD��NYҘ(a�� d1�x_�����b���=,��3�����]������}��!Dt	o�Z��h;���\�qO���pb_�͒x�o*O�Ъ��(eV�kJ�X��򰷥4/�h�O͖����`"��vq��9����J����s>�5�$�Я�Dy�j�8�oz
��nEVM��etR�M�&�O3�ȃ	<5t7�q��+��G�Qabw�ߒ^�am��׬�j2H��"L3䤪Ý@�}���q�j���	�n���3�%�K9bS�~R�}Z ��D��T{
Yq'/��z<⥄%HqE[P�]j�7�zW�?�<æ^�)c�l_�<C�ɒ���Pi���{�PY+�HN6��a�Zء��a֨T��+�� ��}��ѫ�>;�8��I�Ȭ�9��|F�&�"��}LG�}��Ow��饻�Qt���[.zY������������G�]��N)A�kE����ݢ����դi�N���~�%R���Jf�?O�.��_S�QӴ\���m�	gH�;)�>)��̧=���s�(+n�s뗿���B�?CB�8�=&ݜ��*FY�dШ~�	�W���X��?�)e�rε�I�NC�s�I٘ ���Uq0EXy�Z*�+���U����hmk��;1�a��[�&\�#U����Z�c���`��沉��Q\ɇu����:J�W�t[�V�g1�p���h�������U�Ԝ���)���e���Fvn�1�]mse85�.	��lF��c��U�5�r`Y	�E�С�#)�"������@δs-�=T�E���^ ��7Þ+ؼ�t ���
���94&Ɛ�!N�*:i�}4������X�YC��;j�9���3:c\U���%l�>�������٤��&.��򮶪"M��)W
QK5/�<�-H|�z�)<9�vO�cЩC���'��7-�3���(�w4A;���_%Çd�a8]�����G��	�	�X��>n�/�\mݻu�+�
Z�ğ`��W�^Ht��> ����ε�Y��[^7&�=	J��iZK���n�����ȫ�3<���r��.|��!l�L2�L�\�!%��[�F��噙
���d�x�&^�Uk�'�L֟^�C���煗��巸P6.T	]��2�v�T��P@��hW��n$���g�}ip2��V�5=��?��i�.�5���g��(֯��s�z�)�������9��Jx#�ݗ�W*;�5Bh^/}�㥙�nWȵG�=���<��֧4\�,^�{�/����{s��~S�~Z[Gl\��i��Y���~��'�wE ͊���	f�^�!�+sH����Q+:�M@0[V��� �X�LjI��t��
�ry��/9�������}+X����f��J���n?��P-�p'j<���1ӵ��W$Y1��UA�$@�%���*���d�7�3����&m.�:�D�VIC�B<k˄c����\�s�GV�a�%�oi.��V{�l��v`ڏ���z0��W�v������n��X0P�6�4g�	��3m5%DS� ��j�'�ؕ�L��%j2��>���X�/��m�Ỻɮ�N�sR�K/M�:��_���/�-�v6z��
JL(z8kjK�ER|�rG7�8�yMV�T�+�������١�z�L�Cq��E�ێU�ޱ����S�	;��E���U�"˽:S�>A�oV��]&L��B�O.U�8t�o��dF���.����\����u�=H�L�8��q�U�f���@���������{��1 ���Yϐ��x�Q��W%�pC��,���)!�L��s؍n�ب`p�V�B���B��#�=����^�d�	tr�����h������Z�?XE��nZb��O2����R�
e�.s� �]� Ǌ�
�n��%�����G����y{�?u��:�w�6�j����+Ig稀Z��m'�㏆TsSϓ�ɬ�C��I�1�f��_��+��� �x[>�w:# X��"�5�>�e8�O��ZFj!����\�ͬ��9�+!��_�Rw۠4R�#E�h7M�@L�a ���c��ˤ�(�]Y$�b��K19�g�����^�(�RS����B˝�U^�@#�-�#
��Ղ�a.6N���ٕT��$�a���,}܊��э��x�L\�����6�&�¿�oRe'���Q��@.��#�ۢ�y�Oֱ\/�欝뵃;F�0y�{�>�q����+�o��]ms��Jb�����]k��
T��89KH
���ǅAk�秔PIN�y�;��Ɉ�xn�/M[����TK:�wA��rUG�0�>d(K�mM�P(���o�Sӗq��ҽ:vȝ̥V�=U�����+���K#�Atgwm($V�B��5��{KK����)�f�]"ȖzDX��@42OM�py!M���/$���u���`����k�pGxғ�(���D�t���󡬉h�0��;�*D�]��~�8����O6cV�'��x�]�ł�Q��٭o\��)g�n�+�NyP�!͟8�C'?R�j�:�ʨj+[< \|^(ťQZ��f��j1Y�J��Y�ݝsQ��}�ܶ��p=�m�/~e� ]-��D��C�(0T#��/�z�X�k��Qpw>.��v4 0�(8��Uj�3��5QЁ�qq�9�](A�+�a=e�����BfT:� A�EM1���Q���ғ&騱�|L䛵��g_���_�i��z�ϋ�>�9����I;�,ۣ|1)mߕ%-�mݶ��[�+0P��� V��%h�]����w|���A>�)�{�t�b��oT�d�%�#+o_�urF��/B�'��A���{�#�z�5;�/���S!��)����H�5����\4� �>��$��Iu���� ��i�=݋�wNJ�t\���~�M��O%G�ɡU �N�s���Ta6ٱUE��q�3��k�#\2���=[��1��V�gБ�LWK�ͅ'p����	����7GO[��C��Vͬ^3:�$:C��p7]H��������s�֩l!�۠;xQ��۸�.F����Q��ba�p`n�ͺ#ƶl蘿�n��êR���Ḓgg䥉���ƕ�w'd�8�yzԇ˴��̰ʛ�]�b�����+|�G��m'��>�*f�gK�����_��; Z	/�h|�t�q����|��yf-;���?���!�0}|���ldg��1 5�/T(�|�����?��x��ɚӗ����~'ӡP�'���'y凢%�17d]X�_9N���m��>@튫��wYprssB�H㏂��(%���-o֪�\�U�^p��/c�ie�"���)�5��Eu3ad,Dq̃-��0���${9f�/�+�_�A�9_�6Se����h�t���wؖ�>pF�#\P���%�)D�
;��H)�*;�2Aؒ9"�e�_8�n�h'c�.��Ɂ���2/tj�6X�0�PQȐ���$����t��U�M�}�/�7m �Y�����4���S����ψ��t�0e@h	zK�����.K|�E����=�C5; ?�