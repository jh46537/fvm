��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��J��Ǯy{{͂�[��N��������]m�ˈ=g$k�n^v�{.��ʠ,�{������ld|N�u��v$�R�i�f�,Y���v��w@H�o�v�w[OC���UQI���&����RF�-�5_spU8��Ʊ���������k+�(��P�{e݅3�S��0��醆�a�p��ڧ{3�n	��?m*��uuTB���1����r-sG"ة��oE�P�pO����N��;woїc�	����aћ����#��,��O�����Vg��= v�ﴌo�ǭ/���9N�[��Xsr���%(Xy� C:>��o��*�c1x�͠�҈����������x1:���C��ɂ�a��ܱ�\���I���M����A �eNY#|d���������e�j'��k�X{�h�Eʐ��Fmg���b��p߲t5Y-輮�>�����c\Ӓ��=g�*1�1�"M��I�Bv}(�~(���6{�Y+JN�0���G��7��k���hY�p���� 8��)��"ڹ��}�-\��sd�e0^�G��Z>���2�q�4�=m���ђr�s��9���͏Q�"���ޟ��<�+.�����}\9���ޖ0Љ@���L����5z
��˱DO31�}�ri?��W��ꝑ�C��Yd\j��I�j�eT� '����`�~<���A� R�5u]�,����oz@�m���秜����;���|5�GJ�_E/�)��y�4���v���g%R�*�-gĥN��'n	��.ȋ/��.|$��z�&�J.���a�2ճGs�w�x�p������فS���ܰt����+fڅ�,��.XD$���\�J�Ҧ}l,w�:1Ze�A�^�y��t���M�A�dG9�F�|�O�PT�̩�Þ(�<����$�1��������٧Ȟ�	��3#zv��v��tz~���r���:xM aF!�Bk+��5Z��T�����,m����ֻl��Z��mj�i�3� $u��pT,1o�s�϶���T|.J�3�\�v,�q|k�mO�q{�h�U���!������0��i>�:�MW��Y�S��A�XgIk�i�c���%cc���::2�%=�D���\Q$Z���5��(5x�5��������m{�xziU��М8���xo?�
���o�=4��[���k���FP�^~o�ڑaU+B�)�TЖ��]T��������j�m�GYJ�х�8&h�c�������2�Omɢ�5�/Pj��k�S|��X[E7y� Q^�q��m'Eb��u�:P��/�?ц��X�l�/�!����tֶ�_�W��#��PU^��W_ʫy��*��1�5*p����q�{���X�x6x��1u�0��As�A��t���0��dӏ�$?C�g�ظ7���1u�����mT[N�X&z�S�G	�����/M�;޲La�Xp�)��׏�!nm;f/��:FE�u��_��c�v΂��s�ˇjf,[�������R0ؐ>�P 1( �����	���F�������"WyE虧LE$�V�o��#*�����w��b�9P�Q"���Ӂ�Bzi�B4�]�vrI��R�X���r�=�s��2䈡̃��9�x���|e��}e����+{�W�-�5����"��%m~�u�s&<Ӭ��$�vtF��Ġ������%���⸫�4�����×���t-�"���L�9�nt�XŽq�� r�"�8�pc��,PZt<2�����S�Cmhk'�SUyB$\����U:�����t�5��b��2����>r�:F^*²�(񨽀��ryE"��Yc�e@v]1��5���8�[E�d$�y]4�f)�j����˙��O�� i(����v W��,i�|�l[�BeU���H�u������;,����[zͩ��mE@ق�Oޝ�PÈ%i\P�bZ�0�`xg��pb�Ƹ�z
+��irI=���%�/�o%�"�lB�⡀��@�_�p���������JT��Rud���N��h��_�y�
'��`odd.e�x"�S����f���?��R|d�U(��Ϧ-|��?���x�K����fP��z�"ߗ��\˚���]N� �Ӫ���WaZ�7P��#�Ev��mj�.x�����<<���)*�@� ;U����}d��f��-���Z�1K��frEi7|v\�ҋ���� �I g��6_���=U��p:�A�蒮��Q�M�;���|�L����f��K�������pvmØX��z�X�S.,��iST�/�,��qC���/���>�\�N�R�1�M��.�u��-o���a�	�f)��L���G6a;+�-�i2�Fث�?a�k�EE]4N�'jܺ��F==���i/��E�l���ӫ$%��=�_�A��b���n���;�����t��vowJ9��gmd�7�OF�J���+���K��+FwE/��뇮9��!�p���t1Qv��x46�2���L�p&*�tdl�6�&Q)�Mj#�W��m���ۣ� ����a�Q�Q�Y$��#1��0}q�a=R���B�}k�'��:X �Zu��^3>�l��|��M~�4C�e)V3~����'m*%4�P���3g�jj]ФĄ@�4�Y����6cj��3cG��N�0T3��3�9�zu8�VO��!s���aL�q�S�r�p���u���2¸��:;7������#BH��]�|�jp�����ФB���C]C�x�ϕm�Ձ,E˶i\$��P�j���q�#(bQ�Kxf �ӹ:��EkS{�'�F�E|q�2C���	U�t�ٯC�9�$��`�dr?0���e�b�q�
�����P,T���`��+i{?idw@a�㐖����� j���N�M_
j��8YP�)B�/tc{�����;u��/�I�UQ��h܈K�_D]#Y|�7�	C�Hh��{��i;�'���VM��<���̃�ss�z���������9��E��u�F��d
y�٥�ZO�~���U��8�ʨ5UeLe؟V���5O�P�(=���ʵ��K����׶�oWn��j�Ec��r}�3+eD���S�,��M|v1�F?�d��+с�jk�]��9��G�r#��?��vIhfS��L��ʪ�t!�r8�r�Q��/��B��3C���r�.��l�c�+�;vB��W�c�O��[�|�+5���$��Tٷu�[���F����%������`E�cƵR����r2zZ	���8e�����F�i+�V5�N~[m�|���N.�/�7f6_j�#/*�e��|R)F+�u`�~W)cy�P��Q.��{��SZ�t��}�mP�qZC�O�o=]��*�ȗ`*H��O@�Rʳhbf�V�I����S,������}ږ.����ѳ*��k��6n�����$��h��,z��#��<�]�B�W?�뎁�;qSZ֍�f).��0H�LE6�t�,�7�?��l�09��Kl�w\in��u�A��e5\E�+�ա0�^!��tYR�Z*K��#m�"��-!2�X��3�j~O���盂?��>�=#`�H�����AA�{w+�vVd\rPڷ�
<�,������������'S�6�Z=�d"��x�R}���S4�Nd��]4�d�S�N��(q""c�Pb�ٲ���jq�Ε@\�5�xOʣ�Н�����) �U�"��[Cc3�s	��A�����@{��坠��ѥ���Q�(ߐ����I�v���t~�^�%��t�a]3m����80[��k�c.�>\��t]66/�<�	�f��C#��H��<7b0.Q�:G��4���\��C]�P �J��ۍ�����p�.��mV{��
��_�L6�؃<:��62O��&��'ٚ*@������Ti�E���EKY��ưAwԭ ���`���6�<h���A�k��)�	I�OS�� ��?� h���~3��Tpx!����/P@�@��=2�}�`W�sZ��箐.׃�!�{<�`�����,�rySI�?0�w"\�0�3lڃ��$s��G0�̞sX]'�ত� ����T[�jz��U������A���~Vcu�X����uJ��B8��H"Q��D���I�}{�񬒖��	��fr2�SA^@·j�tQ$�V�\�'��T4����a8��^ ��9�4��1��=cp�H1�����l�ȷd�x&���-�e/��p,?�q�o�ݶ�"��?ۖW��2���p7_��c_Q�d�9����Eg�0\������՗�܇��@�׳A(�U%H��3�:5����[̿a�O��>�ƌ}"��F���_V��[�3ܳ��VK\�P��_���rV�+��faV@��N*���g�[���!�Xǣ���r�ID`iW���eF��Я[��]����Z����m�4QQ���(���qu���xK��H��sC猩(2�a�i�6�j� �S52�h�]�ځ����|�z^�L���=+V�պ֕}%K�+}�v�nb�m8nW��C����E�:VF�6��C���Y6�lF�[t����_e�8�L��
S�ko��^4��Y]I��'O5�7�y�O�v�d��YEf'H��˺dⷘ�Q�����X�@��^�fؽˉ��#D�.�a�{���(��&�r��4�l�U�˾�30��e`{K٧7�b��U�拉Ţ��T���t:�وX��R��t��:����A�#�9��@:P��-�t̷%m)���+k}Ѓ�G��GUڜ�~D�����6	��_h2�_;P��s�X��\u5{ ���.����=�(��L8"�����]��^uUX�N\��[�)�=���0���/����>3���0q��Q����`*`ڥ���)�?,�t��\�_�y3rR�����-w�Ι����6-�,0=|yS��R�����W &��[�2m�߾<�"j�B���7*}Cy��xz�� �I	����"ϔ��7�R��oK� ~�����Ȑ1��X�;r�����@��yލͫL�8����sЍ�Bnf���즪OM�����FP�����K7Oס��Ǘ:-֧8���Pi�Y�K��J��V�w�ֻ$?�� 3���d�VX����$H6��(sE@��q�s��ǥ���p�,jF4A��YwMI�S�FQi�p����|2,�����t����!8�%��L��܊ g���@T�Y�J��Hˊ(���J�#A��������HSgM�Lİx�=n��MvV�{�2K`����34pʶ��|G���5.��[�{@����	X.Z��b9��U-��	�����n!_XKq�[}�-����TP�M�s�����̒�^=P~��m���X+,���֩���|���3td�l�±8h�3�H����Z0��Aą�ዜ�w?ۋ�u&��+h�eOۋD�/�Fp}�UW$$xYu姶�s�РDr���/�]�]]u�ŧ��&m"D�S�V�Ԡ��K���T��"��A�AΡ�\dg"dsq����2�xR�$�8��yo!Ϲ
�"Gɲ�_iBӑ�&O��Z��Fo�mi�jz�~p� ��j�
`PY��Q��Y�^�F|Wt{�ՃL�"�^Ȱ�L����+nW�<����| �J��Q��TzBE�<k?�a�~Ѓ��Y�hp�	0�lC��|�2n@8�?�6%����E�.��o:�D���-��Q�
�T�0��zkY�I�� �^���a�a1�jABb�	�y���YP���A��0t�7�ˡ?�8�g��e8��ut:`?�������A{������|tZ�	E�^���1(���m��(��f�yE_s���M�pi섨b^5��aT��������hJ^����R1s�����������9i�c��������.���Tb�dy��:������cz�����6������|?����]�D~���ܔ*�7�Q��P�`DZ7�1P�B;�V�r��Ig�;��ӌ[��@�_����+�E >�u�o�	)1�M�i�;L��#u�<T����u�ժ�n�D"Lj����]�� y헹#�*���LF4��B>@���M��i��BE�4տǑwi����o�T�alu�,��y��@�0��˚��8�=ڲM³��E�+�`J�W+]�AE|�0_�.���8�WN��H�m�	&s�)>>
dܨ���X3V�8IqM��H4�hGj�Fw��"���$l�h��B4��Sx��}�;6�9��A��E"f>�΄��۱��k�����������F�K3��Γ�?u������V!L������4�����?6Y%u� *��#'pF���=�ڠʻ��f�K]��FL��=�[{/9S�t����_P��Ԫ���Y��?�ib?����B/����"y��K��_����3.푰�F�e�d�G�R ��D'�@�����Fm�+���|��0]H��'�ޱ>�ar���I��rH�hpf�^�܅\�֚>��E���5�`l�#�`�iZІ{�>����LZO��� �Z�OZ��#^倴ʒ�6�����Q�1J̤v���5�I/�x����:�.	'��z>�����VQE��2�l��Сuu2�6��0���չɨ�K
sF:�_���C=a��w���&�RN�j�^Tk��%�M��K�%~Au��q� ��¹CE����/�t���n;��	�׆��pr&Ӌ��UN�BJ��Fs]�׭T#�S��%1GL�3��sI���������L��\�Y�������&f|`�Y~�w�a��;�h[�.����]�T$������zp�����-DȚ���#	g'�ȉ���6ݚ��?�
̎���l�aH�p����������0td��錁X�� ���'O�挌����2A�q�go���#�����;I[�kG�Xq!�qL6͞'����T��/.�u%'nN�,�2���KM�&>��ƅ.�򄙺x0+����_�C���L�Q;(���f���]`,n{����Tn�.t�Э��~�j�pkga��Z�xp�ᄛi���&\����6��K��ڞG�fҠ�{�s��IuΒ��ii��la�c���[%^��H���cX�}�zaL�S{�zS�T'�5{O����f3(	�$�ؗ'�<����<Ľ{:D�m�~&���1\��6�o��OW�M%I��f��c�n��B�(ى��p9uUw0��h]���.�\�WgFQ��]ۏY�	K���}�A���,:��D�ӧ:����9r����D�TøZ-�F��`U����u� ��#��!��Y����H�@P�P6��jxs"�����a�Z���%� �t�h�0b�ټ���t��	*ci��I.�G���k훔��v3k�AA�;��x��F�/�*1�^8�S��{P�-B�aFr��.'�)j���9`��o����uB=�Ht7�Yʺ�m(��#=]�"��~Џ�t'%�Xۍr����¹�w�ҹ��2��I j&T�,�f �=vtse3^0��X �r8g@5�J��Zch��ہ�11�V-}�x��-��Qג�6�V��ѝ$Ʀ�HRh�]�'�@Z� 
X�W�q�+�KAn/��	���a3�]���9h������o�0���H�>�Y��"���A��d|I�՟�>���s�^��b?�!�[�#�N��.�8ƅ�f��NQC>@ݥg�f
o���|A	��󡾻���=�Ӱ�kFtD9&3^�%�_��M�W�\��Ԙ��򱑜��L~�%�������aj�"�����l�oC%��-���GШ���3���<����ĕ������VS�ry��c�c��8���9~�t|8�4��~�H�d^/���gT�4w�>ޙ��3*�)��o�sp�c,���3@����hO�Bv���+D�<'�=��M��:�K��j��� �*|��)"����"Zr�Zni�KU�r���(�Hg3��˭����5���R5����W�/��%O�H�Y�Z�cuV(�R�aJx�x�ࡦ{P|�������w�F�GL\������tjS%��n�_u��з���[&KN?�xg�S��)V�����5�Lw<-.�M�"��G�T�rv��?��_b���D�<�=��_
�Q*;Ng�;f�����@�����~m�ω�c��W.�l4E;;����U�L�{,�X��^��o�N��tLg\�d֠�]Sn����;�ٻ�+���\I۝�=Ap��n}-��EE\ľBa����C{�)�KT�!}P�c ��?X�xS��;.x����\�8�W��ҋT�`����D��ׅ*��Cc�2$��2�z��+��K�F�����N03y�t�sY^�1����#ജ��u(�M%��arq}P����`'������mi��,����V���5��E�S���j���g���y�<MZ	]�>�PҀL�^N/]ƽ	-�FP�U s������ ˭����鐎���A;���*��5�g"���k�(�ۆ�8!z���X��Ee���;!��D������LQ.`~�hCI����}7M?�v�ʽ4��j\�+eғ%�=ıC}4���m+
#�܅��
�]ФM�Z3����ɚ�ࡧ��4��︁ `���2f�Ɔ�!���}Yj#0<vR���i����z�mM,��7_���Sa���:?���B������8ÛWo��N�3/���s�S`x�.؍I�"��^���b� 4eO��~5�\R��v��7Ĩ{��杻�KJ���1e����A�\�sH~M�*E�xI����v�V���n�� v#������3A[���g)��$�;�O�&쉈�Pٵ��-���kJ]��&d��5 ;��=g��<��b�9YB�ћtsnl�Uz_όߏ��e�mv�@ �W�hÈc��?�W��[B��-)�_ګ�ׯ0��̕����������tJi$WO��S�j�HVU��نЫ��.�EA'�K�4D�՞�j9����a��O�c����;�Mh�|j�-l���Z�G��U��뺦��sX�D|�o�M����|?�mI�`ͩ�����c�^�#�`c�t�K�������\���x������	Nʺ����G٢<��D?�%L{w���.Y���.e�L�
A�ĉ�<*����R7��;�!��v��&c�u�J~�V�^�ӈ�c
���)h��r���ќ�7�G��ToF<�!���� +I5 t�l�S�Z�4��
;�3��������cW����='4!4C�>���+t<:��Uo�^m�M�U:j���΄�4\[D֊!�dJ�d1P��ʭ�������M�w���j��ɗ 4_��^΂��=�7�˱yUL�³��2�@L�o+ F�
�#�p��R��:�W�*u���:���;3<�򡿚8¤�I�� �ݙZ���)��)0U��M��7G��v2��j��d	U�׭R�n溞<B�%*S{�&jQN`@3C��Z]��MY�#��%�>�=�󙎋��P���=�����e�7��sO^�b����5�(&�8|L�H|Z���m�<��Ke�A�ǃ%-=�X����+��q�ɍ�|�� 1�[CG��j�]�qm�G#'[[��8B�<������2�󬨂{�_�����A���xD>�_D �mA)&��5��r������|�F�5�a�Z�����i��xIK 7@w��g5�TDI*�'�U�K��}g*	��bըuc���r|$�rBD�����)��V��
e�蚾J����G��XMP��4���ޥ8��/�DT��:�|�P9X��x�,�F���.�(
��4$�/��D9;�Y�:����k�r���σg���m:�D�rXt�H�%��+��0�{��W5�t7��זq6����������I�y���kM~�~�k�˖|�&X�ʹxG���rp8c�ۭ� �TjO�l[����uXIS�Z/��-�V;����I�0��󚇤@Z^� ������|�9L�]�S��C�1�;?�.w���އ9�^��.�)2���N�$�\���v�Z���l5hz8�KM%��N�ʳ{M�)kN�*���!P�W����H�ս��+N)�I����j��C� ۴9D��P���Vɚ�:�
B_����$�Ynh��;��v|�"|�\�s�M�w
�ZT,�K���޶��`�p�c��-W���t�olG)�C��/�8��©�l��y����,|�|=�KkdU�-ҷD�
��j�~*���=�)5=�ֲ,o��w?O�b��"�S��2���	e�>�+G���+���n�c�/׽�67�~��˵r3�A}m8����yܮ�D�u�ȭ���
���WmY<p����c�גQt�	'���X��Y��5�#R�O�qu���}uiJ|fFR�l��/}����ȵ� v�nqn�0Z/��Í������E��փ��� ���]Z�`*���n~�{Mm�x��6��*>9"�r�*���()��}�1�e���F�i�{��p�[���'�ih��OBI�r��R/@�*�Gh�p"�Q8z�+� �%$�O�$�H�� �e��P#�A�4JۭK������d��ڳ|;��\��-+��>?(�-���� s���R�!f���Ni��f�T��*���t5�P쩫������W�]�2�|�9>� +Ȑ�w���D�"|r��������®.�q)�r��$�5�dl��_�Y���-�}[��e[����b�0~�b�4U�l��u��y{r}����򖉖���xV���w x������I�Q����T@�1��90��-���v7��akE�֓w �\sc��#��Gڳ�17�Ы�g�b�]q3^�!)�I�	v���!D��U?!J����]Q� 8�R��&�m�Ls���˱�'����f�.��oe���
G��z�:~(%���$��g�މ�Z���`\u�r��{4m�D���ع���;U�WD�T��v��~pxι�G�0v�U�B'�~��ݓ��U_�J�d��9 �������'r�`�V�r�����X8�*��*�%���\��W����E�<@�����g����~�X��Kw���H��}{�	^^�r���:��s�	M�'~J	.�ސ�����j�=-���섧��B'��Jvt�n⨾�u��_�2����s��3fb�|��[fV�u��7��$�1���҂�P,m��M���j��O��E{�*M:�]�աV7N̎�[��-V���W	�1�P���0�bx�Zږ�7��[��.��29���M����c�H����@A���(�ǳ޺�xÒ;�M���Ws�94)Ns
N�t��־�W���h���h�L��U��uN!��	)͘�t�(J�H�-K	>z5�0h%A��o��u�� 2�bJ���x�m����yPn_kr��j�����mm�T~`�%�3P��E����Uщ���>�5=�Q=��ؘ$Xbc@ݽݭ4�
ǓL�F7�
�L����������G)wp�U�r��M���;������n�_#r1$�,��l
]Iǉq���^�_��	|��F)�?����J��7ع�֢?�jE)>C���X���<�q@��l@���k�p�Yz���Q�"Odد�L��V�5��U�i#,Z���7������?����>�\y�$���q.��.�~Su�wi���T/��gH��Wb��i�Fʋ�m+���Ks�%ޓ,1r��|��_n�jZDY��3s�E�3�@M&V���@)��L6h���Ţ6ur�d;hW&�EG �A�\���S�oe�h�b~�l�tW�(�"��[�J�IJ���Mʻ��}��C-�r��Ӫ�ҫ��l
�	��"˦� ���ϫ�c3�1CI5� �&��Rh���RֻB|-u�[�SB|X:�~iN��%�ԋ	���c�l�0j�0({ �5������kf�c#J��f���3���L���2�P�n�7��V��#��@��S'÷]_�ֲ	��Ҵ��b�V�!�W1�DX�y�դ�n+$��Aqf���>����d\�.}�<�ݸ�"��Y/����d4��':J���9C�B��#<t5[�ױ�(j��p�p=���	;�H���΅���C<�@��4.1Q-d�KS=<�)hQo�Ɛ��������Ujs������r����MGnE��%�N�!���U�'���������?�q��A�|τ����]��%M��L��'̪�=4m?}���o`�ҷ���w�h�{�S��Z��߰q^{�Bjd��P �M�Ń�('��o��kߨ�r�����_��݇*��#@�S����6�$�|�,�i��h��̏C�K\*�h�wgx�AGp��XUj0���޿5��"�eP0��Ns�� X��fϞ���� G�2�����J�u1�v���O��������� A��h1���j	�X\*���eǍ����0��U��i�δ7�D��,[�~r�^%�bA�I�k��ң��C��@`F?�}A]ڟma�C��������U�P#Iԏ� ���]ϭ�ﳪ����'S��Ŕ��)���\�Nn��{�$���'X.t��z����B��O�[|�8=�ҺA,^���a�)�ی�)�VXf�@�d�ƌ5�E@�Ybވ,��$�2Y�-E4�Z�&�`�6.�'FB�:�������{�{.06 �1�w�,�p����:���!�^��{���C�����L�����\�2:�yO�f6gE9/�UN��Glw�7}�����R�.q���+9���,��"�� 5g=P��\��S�R������' ��î��n�e�t!D$!��r��ħ�t�V��=��*����^�rB!����$�V�	-����dm%���@7����-E-K�*��X��������L��k(�K	3k����Ņ���}Zf�1�.%"��R���%�����J^]b����Z�J:� �Gi�ȸ�b�*l��W�n�K�����;�y�te"�)�+��S��[�,�9ss�U3۔����=���G�������	��f����,-e*���X�����L[�&D��� �z�GW�n;�)&��T
�����ʢFM���"m�+aI�P��g=�ԝKAF�Y���#Xz�4���Ȟm�4�=(��ş�ܙ���K/*&�PK,7h<'dQ��T"ife�?�@�r�筚/��D���R���͆U^�J)��ME�cԹ@|Ҩ*HO�^O���#F��R�ړ��<��D��Gц|����Y$e�L��\�#�{��N��_hD��|_�.L�
�?h���>��g���M�V�;E���u��"�3��H`��۾��+�y&��,tW��5�<�N�ʭ��B�CbG��������c��֊�#�Y�Z��xT��䶭���J���aP�K,��7
:�!�;P��i
gO������+R��D�]��۠$�~3�C��>�*�%���³N*�qW]�x�F��,ʊq��ór�����}������k��pG#T�	�Z�r��'!	�ԜF��2Ta���ǥ��Lx��}�'��Ui�����
Ap�OȠX��/�(4~�{���s� �Z��r%A��H�o��Ir~���p�0b���3ګ7�=�`����o����	��!*y�)�Jj.�>fG-��đw�9(|P�28Ȟ�f�"�Qg��c����K�z/|
Te�-]�y�Q�}���?����P�<絍3�Qv�zZ�Z�wn�e�Ȏ�	��9�7�ب�5/�;J�rX
��w��:d�7q"mֵ�ci�%���GCu�٪�9a�@+�Q^<��=@X�����5��xe���KP��2���),I��*���������(e�j�(��T2(q`�_n�>��N������Nmyz�4cvQ�	��=�S
�����>t7��jY~a�qg����>�[�}N]2��Ȋ[�hy�����[
^��
���.��Ñ�[Ubh�6q��rI�*�/���`&\ ��`\0��	Cà�qj���
Im�/��Y9 ���vV�>���M�(U�+} aIY�
�����B.�SNs�~��y��a0Dq*@7%�+���L�x	�ˎ]׀�|.�i�����K���W�"-���C��A�다<�
�����TZ�;ۡS��3Rh󥸗Y�zH��h4O�oIZ1�У曵u�2ѓA[J��3�h�n1l�j�\�{g�1�<Zk�c�2����2����G~��O*i�R*"G���?�a����~LDlj��#,'UTL^�^p'�ӳ�LΒ���YߓK�P˗$yr��f���A>�ea@��§|P��7���\� Ս����J��˺��)��tHh
��鎈6���a�&x���
������G�9%7�� �����C�.����_^5 �����窮\���8���O?P/n?���[l*������J�zA�gm��_[�"jDش�����b� 9e�#h�	Fje&��ud)�ƃ������F�f�ĔcUڮ��:;H�k�ccJ���׆���B@�{���"����~}{WsI����^�����B�8�$�{l�˗����F ݱM�F��R��8qa�����"�h�~�<�q���d��>AI�_��/LM�_�^(���7	�}V�b̀���!����~�e�����c�������*l�Pq<���	�y�'@S\�����g���UW��I�{	b���	Jus��0�����a����-�������f�>رf��;>MC���!3NV��h�X�4òQ���*o�a�Z[[Q�����`��[r��󨄱v��k�Ns�K���bu�\��_�
@;�T��h�"�,�b
��>�)��NτF��☵U��<^DS�����o'ET�P�;��Ϊ���$�q�5�k���xvR��3����	n���?�Bb��1��֢�`qJ�yy��Ɔ��0���SXy��P�m��Ovo3�=]R<t#H+�v�X�z:G��P|�/�ݗ��4���Ŀ�s|�n"ٯL[1EZ6�[;�/SQ��e��39A����xW�!�x�c����
�\� �x���"��p�U��� ��Ea�'Wuf9�cI��Ň����\��� $p��⼎�s��L��G������9++����L�-�>��8����5D�^�B'��F���Xf�(-t����āmFz��PEOf�Φ�-l�c���em�Y�hU$��d9`E�.���:�8���"��}ȉJg�M������6�K�F��r��	�Y�؍���
PO��+�vE[.h��wn�[�����y�Yx�� 03(J ������|~N��9+�|�v�������'��%|��ay�, ��`2�h 
r�-aӍz�Q�zG��D�W;���	���"�؋L����"�%����i�F~�N���M�ț_m��!!q�Y<qNQ�<��� ��H��z��u.��hط�&qd>�����1ew�N�&$�@U��������#G��[��95�t��DOc������o;���AψDɎG2R-�i�1,Ň�ӳik�u�Qqҡ_	�U�C���VƮq1�G�O,��d�Y��huʷ�-򻬣x
mO�S�/��NĽ�;N������5���KG��Q.��r�LR���[�g}I�Ar�������[�x5�\�W��T[C��j���~]�oj1o���"
����^�_�hص3��t�Ma%��%9�L�`�M �2S�;��n]Luzj�S�naCc"(>+�|���m�!���� �V1(����'���,xp�)d̗���Q�"����;���%��g�`���ٜ�*k �S�^覸WYG�o��3��������Zg�`���@Da5�b3��\J�`e��@��ض�W&���~�OD�9�A�^-#�
�Տ��UQ$�,Q�J����H��ice�RF}��l�d��o�$�2�Q�js�����njA���
G)�9y�8h����-�dI��r�����0ᷗ}�/�������v����Q�%�ȕ|fO�"���|X�0}7�8�G'��Pկ���Ӯ�Gg[�b^g��s2�<��i�c�S},"�N1�.���+·�A�����ɸ	+1m�<�4��9��7�3Cٻ��{B�p#շ���uDD�>��RK�o���O��!���Yh%d�װ�c�g�>�M�]�}��"�|����S̒:�SƱ�fQ�6��El}c;W>ZFM|y����N��S���a�2��7��]; _/n�<G3����ͺ4�ƞ�I�!�c0o�bQ�n�n���ָ&�^�`4��E�s���]���V�{d��<w$�f�G�N�+�ű8$F��4���q�a蒬32��3ۜO��fխD!V�4�̬��9hc����.�q�8&��A�p�DM��=A�o�z�9ON@�>����h C�V3e)Pe�~f�l|�đ����Ě�R)�?I�8L34U��Rp�R\)����
��`[f3��R��xG5q�$��� �/��`����4ZgQy%ȯ���T�H�]�p�H�޴�
�jJM�� ����}�(�٩�iu�%Pm���hҏh�pf<(�.Z�4�F���@h�[�	�lg�2湕�y�"��v�5Np���eý���hp�&�ֱ�h�k��7�9^����]{Sͥ1L	r�u>3V��ϴP�z~_&
��f~��0`�tf�e9�y;[ �9���Ud�80��=�.�����j��x����]�k�������sU���������ۼ������H�|i9�n0h68���h�A{��F��6�3/�����ý��֪��l�mA�L�s��U�o���TRW�_li�L��K"��o�=�q�LG�O�a��J��_ ���;%�����kS�vrǜ�0rY\�&\,R�M�f����Ziw~�On�ij��z���y���X���L�����k�Yߕ�Yu���$ܲ:Q"�ۀg�Z��������B��I�%�Ё���V���
�l�	�T��A��p�����]�.�lЊ���w�@z8n�s���)���+���-2%�̹f�0�]�/���b<"7|���q��!c4�r��R����Q��*K�s͉,��ް.��;��9˪�տ)�!F�')�kJ̱1 ����eM%1��V(�ڡ��2���C� �$[����W��g�ju��u!\�P�9P>�q��A��]�X�����}�:���4���}	�%@�N���b��d���{}^x�F�z�T��>Q�wOd�#��Fn���%��� �c��i�{^�b��n�ޕ�`N���{��Bd��=^B8UufP��I4���~s�S4q��!��^�(���Y�p�:���K��3��3op{��(p4��AI��5R��IbaP��������t�=C��O��@����?�`��%[�3���T���W�as?K���C /![��}7oI�s�{ѧI�q��s~.�nF~.R���ͥ�ė-���z��y�e)ᐡ���		�|;�ۉ�7k��'�Ɗq�BؼH��$"h��w�g����dgZ:�1/v�M�@�L��(��^�>8��Q)�'7���3)�H4�R �a���&�z�s���w<w�4#��Ŝ���-���c���jl����S�ÿ��4�`b| ��*�!�r�~�n�e��(
�S8T�9���V�і�7a�*|��r*�Q|mxMD�@'p( �y$��Z�s�&;	�k#�.2'���o�(ho�a���pԞ�6�˽�:�?�IA�W�ʌx�����g��v�d�Z(�dʪN�� ,/u�+٬��QI��9�D�W[�xj� �C���Jj�U��t-inOA����y�إ\��J(�<��h/VxZ�U�S�\0�:P"И���-�x'	$�!^!GW�+ !q��V�T¶�c"�#`:]T��x�<�D���D7W�����b��FP���v�2�C��}�;��=,�D��)�/���}|��@Ԟ��^��1��K$b�������9��7�Vl6�>+��١���+��P�Taη����M^$���s��m>g�TT!�;v��c�-��<�z�s7d�zL�m�OE�mnp�@;��f��8�v��N�?��Њ/BH��#:H垼�K����@�CS�'�D��?���!�3��9�+Y=��w_є������T�D7���v�v�-yI�;Q��[��.�8IIB {��ŔypJhe��LuH��c+�f'�Ʌ�+��������p��|.���O�a3 �s�v4V��:�E���ll��Dr,���R�K����Y�h�f;����W;��b�K�����&�ep���,UU="z�i�3��Y�ۭ�Q7	�f�� �S'{��U��"ezu��a�+���~���
KT�;i��B�9co�fI�
Mʓd�p�X�r%��c���S6�Y]�D=��N���q�}���U�c`q�4z� cy�w_O*q��j��ք*u��@�z�[��F^ꈎD���}��Jr4��~��qf�ce�I�Oz�.�h�@�>̀�3f�¾@A�˴��0��+;,�0��|
�����50UB70P{�-![�__�~~J�)u�"�A�	"�ӂطq�#,���|9�N���I��D"�����6���� d�WJ���'��U�ۙ��chQ���ܪ�N�U����.L'tl+o��P�&诹�-xO�M�PM��A��`.�����h����M�|<��З�,�!��r��h�lc��zF�:�3�L�0�3�$onK-u�t&j�1�8$�ok��;����)4��.0���XQ����֧��������#�o"��_њ�v7#��C������&.ƹ��n��8��<�ڞ�F�҂��17�a] ��F\���)�%�;��'t \;hn�����x22���61�osٮTF����Ơo�PUj��^�8�ㆭ���m�r�Xx�;��*&�u��� ��f���N���{������Od���S!��Z�/��-�h�"�����'��>B���k�K���*$��T	�+����d�Z�H���ڎ�s������o80Q��!זJ��a���R��C5r[B�0��
��86&>� -���_�O���|p�K6�m�E��|q|C����`��dy�!��'A�W�k��,�Ht����*gr�2I�,�߁r����K��9T��"C;tm��d�}*p��9�i/O����
���"u��t��d���ly�V�z�)��߻�N��K�s���ﵨ˼�FH����(a�t�%�=m��N�l�7J����A����kU����,o�W��^��F�G���ٌ�a������Qr���-��V[-��pε�6�A�Ojm+q�<-Lw]��$ӫ�� UN�-!b �U DVx��)�z[n��]���2GH@�8�u�� a���z��7ւ���yDL���"^��A�� ���!S�J4�kY��fʚD�"�Z�V\��;<DYz���4=�>|��o'qOC��i&2�(�k|�ޡ}zo�]yh����x��'�X���- =\:+�UKu�Z�x	3='阰R���� �����qiӱ�rU���T"�e(�|�pN�x2�#�	g-e��\� -�l�S���s3��ՏCۋ6�l���AU*at*l<�ѽVr���~�j+�z?f8�����F�J�.ަ��'���&g;�ީ��.� �C��~C�� ��*v<.��yeg�ճ(7�lt�3�d$�p{�KL��<E����C&��Od[\�g���ė� y 8l�T��"���/�l��ƪ�"
7��?�������y�-���LP_lư�
��a?Wo��$��?��+��@^�GM[rja6�|�`�!Q�^H<��o}�Z*h�b��|��$�\�l���:F��fe�-K����_;�Ot(4�?��(�IVo	-nЀK�3t��g ������Z�R�de,�����*��� �<���z�R5̕
�,����L����Y�Q�4~�ۉTe����Q�E
�m�yß)yc?V/;���4u�nlu�Q��5&o��+�?�#�Ԏ��B���ӱ��-ב�{U"�
<
{�k�l�e��lȸ�1���_�D�V�NGó�ds�w�͊������e�y�'rAXg���@c1X��%��R� iҽ��K.p�U�7��u��h����p�VrV*&��vP(��������/e�m��� V�E��}ρ���I�L��o_�ȣ]���;���Sc��σjV���۠!���	@	>���[�㪅���\�vPԹ�]%�����%�mM���$I��4�K\����Dđ��p�*���
Ud8�p��q#y�wp���e:����z}�s�����&���K�{�o�a�����u#B��Ug��%�bekλq�a�}�KC���5WN̫�x��M�8Q�j
>�Xd�GN+��4���v�ʤ,�
�A��l����X�Hb)��Ɍ�L���0�"C����-?μ��������E�����m�#"���L�Wf]�����
<���;�%��u(Ġ��9�|ˮ��r/�m��9co��j���>��R
�nU�|!�hp�<c@q�_�z1l���u����c/׺�P�S2���>�1jS���~��c������5�+�@zb �<�C0��j�Ӯj��s��:�C�U�!����w���5$�΃|�F���0B׮ ���8�����g�q�����ĵ�R�?�W-l;��f�����r?^u"�'��6:C�7ȏME}���Γ�Ğ%?���F�N�7BM2[�������Dt�|��gq\�:;�vo$���>��:|�Q<��^�"�@���3|��Bq+KC�Y��U��N��G��9^�ڶ�@���>R�VT��	s��V"�<�0s-/��ufśMlt�[Y��E��wB�H����]�TS@�:HhK��F!2s��Dvl��SM=�@T0�((d.�嵸�A�c�;Z�NEh��ʺ�T���m�u�g�����P؉��8��P��<E���>��"�n��t�~�%�u��Zw�T�_nUEզ�x�^y�����f��3���5��"f�T���˂�/sW��Fn���P�6.��vd eE�ǜ/��9{��p�����>����e�Z��GTG⢑.s�<�DP��`mUA0"�'�T�m�#y�*��&
9�����X�^��2@н�K/~vs������3)7̔-��bH�����	�m;�W:��-6M͚����1�wɏR׽A'��r�@葎�hsi��R�k��V �\��%*T�&j��g���8Q0,��<#�%�ʋ�B���x��BT�|7����$7=����B��@j�|��{'E�q��{�]'S�\�$�h���C�Gr��4>~r^_r�ƅP��^�O�?۞�Q@{���`�q^�n\�l���-���(Ѻ�q��ٔ�	��5H�^��2KIl?�At2��-7ؙ�BL]:c�U�<�s��9�:��d )B��������H=��-�f���ׄ�U����dY�L�t;?��o��}�|q N�sD/I{X)�_�ks�k@Bq'W�3\�_�u��Y����}9�k�P��/��k�����D"Wv���Ģܒ��=���J�Q'�E'���;��U�n�J'�dE���Ѱ5h�W�n�� ����Be��c�a��f,�X�~~�-��w����ld��S�T�m}~��A}_��Ph��~��¤�6"e�I����D/S:�0�d�y����g6S��1J}q��b�����bE��wѳK�f���;�nc�X1�",��Lq��h��$s9OY�q�r��P0�ZI�jl���L3>_�* >����O��2&&H�s�2����sϻ>����v�ԠI���өT�+ �`xz_b̦�t m����HR�w�Q%��RĲО^�o�D��L�0 ������߁������ �d�儃��M��E.�bq�Og��f������М�l�Rt~�qRTV"���������Yʙ1�(���P*dv�oN����36}y@�Yj.�رcDȋ��p�H��+�N��=��Y�&<n.m��;ɮ�
aV�p8?j��3��k�m@X��8�Wg�a@�ں��O��6��?	,����0�5�ٸ}�O�L��բ�㑎��y&$G�쪒�`�� n[��Q2��mZd��rB�������>��ˎ�j��$V�Ӕ��v-�OI�g(�v ��L��t<��Am�1}���Ԕb��<�'�����w�g�r��=J���&j�\�����?/%,Um!�ޞHD�.�hB%���X�pk׵R�V���*W�L9y�P�n��=�o�%�^�WPR�G���d(=�"�g[-6�����n�:i�/ļ<�n㚺�5�������X��yP�fu�&e]���5b�$l����ǝ$7���PO��i��;Rn�G�p1��z(�wam%���N+�(����u��Uc�Y���?�r,����(�V�Ɗ��8К-JG1XB���6;�а5���g�(�.�e�'*McG3.��(jt:�2+d)���LI1�c���0���o ΊD'.iG��ID�'@1^Eܮ;�V�A�˜��z�3d:�)S�U#���W3(fAeg�d�+�|@��Ͳ��/�S"��k�]�M�j7�Ul}��Ǹ�n4�y0�G�~���c�&���+CM��	"��ӫL�uP-@k�����h�ߍ���p%&�݄�}�EP��L[u��=B2w�m����2�,�:+\��+qS�F[:@qڢ�~�y���S"��^�Q�[#d��/�Q,���11˸��s����ė�3�m���C�%ypX-M��f ۦU�)�:%5�� �6���f֯�d�ej��d�(��]�H����ނ�CʴNwY��%ޥJ<�cj������f� H�Cı�o��Q0Ag�+v���wӬA_E֊X�~�sb�㟩n=RqX�9L.}�I�lU�����Of��+FM�����7~��w3�L�VBxO=.E�n:����ȃÔ�/υ���_M�i5l�U�4�h�ƴ�͒!r?3�!i����� ]9��]dԤ\Ue��m;�~Zx4���/=��<�3Ӫ|��a�~�LT[�*�,�m�	��w�r�v�k���}/dJ���9D�J����p5�`�'�Lk*��o�&)��ۧ�]�����	���c2[ݕ�~�^�vx�+�]7$��L�AG��e+.�X\��ms�S1�n!鶅�u��]pͤ��(�E����A����ד��Ӫ�s��F+��lI,~��C��FqEҖ��t�����6��s�kD}�#F��ah�x��������l�:��SO�#����ܼ�n@�|�@�j��@�]qoo��]�o
��[�G#P�CPPxP��� !�rs��5�.��%�g�L�)vI���쪋��3"��7�l
��_�)l���OQ�Lޞ�ѣ��M ��@����	:4|�����@?;�;<��i�N<l߬��n̔�=�d���kz�������w �n�W�p/46%P�3��5��ؚ�.���P��X�G��wUs�6�e�}ϹyW��a��m7�;�>���?��<Ss�G��lE�ՙ���sWX�[ >�����XgH��3=L,hH�����b�´!
�1>�ga�J��sQ�$�$��d"׆�I��$v K�mc�%�(_�L+������<����S�$e���=%DT4�Ӝ�n��]��
r7��_�]Ķ�/K�����x�SK1�-
Z�
֚����4A.n,KtI�.h��h��az\q������s�
X���J�ʩh<;xr���V��@.��5������̘��7�6	����*���YVB���KP0�{��1L���/���U��z�$��6L`�� �$O���b	�<�hIqm��_pV/�1�ڻfڭ1�%m����_�q��^�Pr$�[J��h���E$��Ŷ��C�{䵉�KR)��(��6����f_� ?���f�P?��^U����a��؎�D�]��s�/g�F��ll���.�ϯ[e��#L��Xh����%�_��^	�4\ﱜe^����=l�Z��ʋ��	��3��A���D�(R,��կ
�W� v)���"r[��y&���p��.�0i�5s��;C�f6��Ή/|�#��ņ���$��G������zŴ
Z(*Rw����x2~��?�n���JBe�D�oGAvg��;GZ����J�G"�2E |}�D6Ǧ��ꢬ\��Q��]6񮵇8��w;�,(� ��<ohi�s�/�Pcu�ϨC�
@��Wp� -dA��:�q-�|z���i��#C�6%p��\�L���-��Υ�{�Y�r�b3_��ǀ����A�Ǿ��@^�`���
^�}�g1��1����0�%ZT�T'z>Ke�ݩi���	�5`�Q��$��z��TK0�Bt���W|O�="�?��	�I�� ���ȗ����h֣en�^�����x��������;�2�
L�Q! 	O2�.*�9X�D#n��m�RO�J�yJ|.�b��Tt�<�f�������6�h��C�o�Q_��	����Z���⌙��b��5X?(�^����6�^�سK`�l�a!���N4|`���a�~n�!Y�uic!MI��P�f�.\�ț�_E�XY~֖�1�!��=�"C)��Lop_3e;K{ R���=Z�z!!H��V؊�-�@�-
[W�[����	����i�c� +F"+������& \��a�\S{�:�Yy}���SJ������J��q�F*������-AF�?O��%�6w۬�S:���	El(�o�bQuϣf}eV�"���XK d�G�(�m�f��:�["��_�2�0N.7GQ�阀%�k�a�#,�G�zI � ���)ѵ&7ݺU�S��R�φ��bWKC��2�}wxʫ��Ĥ�REYu�tޮĒ�+�P��3u�\��g]��i�ὡܛ�$7���T}�����m�S��VFŲ�&%��j@���E��g���r�=%��+���7j�D1��p�|}@����/ȯ�B?�P��6��<���z��b[]ם��@%���Bʩ�?���d�|ې�H��M�c|�((}g�ݙk^ ���+ Q�y+m��q^r4I4'���^N6�]<�����ꩧG�R��/�P�����Ǒ�8 ��&4� ���i�>���,A�W����{`�>(���+mA��]��4j
`3w����w]^G�ވ��ț�9�/D��;��`n
?0���"zKvHj�=0���_s\P%��f�& �3�%ͤ�Cn͈�i�ȭSC&)�����P�^.6�_(�e���(�V�q�$�v�bں'7]��Z�t:��%E+�u�d`5~/��-�����
R�T�U�C�ψ/�.`�q�@ �<ae�d���P����w�p��k�?l�5WhF5���LC�_V�$�/e콄����΢Y��@'���y�$5	����b/��C�1� ܃���lHF��M+S���c�d05�������2!OP��)ܕ#	Z�{�SD�i�ެ���Wĉu�j)�ač�n��|�I��;\"e0�SU�-|�����]�ٿQJs���N9�ʏ��P�(z�F�(S�_SȰZ�c"H^��=��V�[٪���I�k����T�g�Ff�%QU�A<j5;/�3	���5�=��գs��31��h5��ґYcRx�JF����0#;G�9k��kȱ��r�Oo�Xo>!~��λ̒������:�m��A:+ �|������i"��m&��I@��3[W��m��p���M�M�.���h?�P:�IR�o�6��d����i*�Y�|)ob����fZ�����Y.XeuC*Y?*�x��
�Ѕխ�P���X������4*�l�۹~G8�S�ñ�J�jآ�!�+sȆ��y�&+�,�\��C�"�����/�����W�,��¸;�f�HV0��_�v�y�Qv������������R
Ge�Z�$�@?�)�&�Ǣ�|�^���0�;�Ԇ�9oP��hr
I6�����Z���AP(��8���s_A�y&�RJ�D�!�5��Z8�����q~�\~hf�
v�Gx_� _,�Z��F���^{p�4Oi��nI�-�>N!zSd��jT);��5�ۍ�$�����F��N)]�N��/����w���[p�����M��n�7�m�^B.�l�S�)��P�SUf���k�	���/dQR�F&�U��2+��"kvG����2��
�ޣ�K����֎�G-�S������
(X:Нˡ�Z�+k�LT���,�ι7"`�Y0J�A���١w�D���+|�p�����\�9�&�c�̍,�'Lؠ����F_�T�h1���JFǒ��3�'���*��7�<�J� s�zibI����K �T�=�ϖ����((C�ݴ��;��2P5�N���3�-�x�m�ǃq��%ED�x�ز�o���2M�i��SU=��tN��?��P�����ObNE0�	�K2���΢��uA$b��Q�A��X1�K�R���0��#��b=������Q����ʅFJG"���wM�dO�{j�`v� ��h�s�}V���-�� gY{�<���w��V��"JC|Nk=���2��Gq���!έ�!, �	�*(׍��)X���w�j��SGX-�78�٨JP"����lk�|q.�*<����2�H-w�w��/�fE�(/(���D�3~ܘ��c�kb��4�b��X�E���E����|
�� ǭ'�nh�p"��U7�C�D��Z�!h������'�G���M���5�C[02N���\&�^�޾�8�;}�󙶠?�%�׆���0��3+�p�Oc�P�=�����ᥠ�� x?evnMDr�
��P���dSrn�qA?LR���)fk�\�������q�WSK �v��(�Gc�p8v�`�Uk��^粴����Y	D���q�,aw���ZX���D��G��µ<������ �ST�%
g�]C�*�9�Ms�&Z��o	����`�		6>���s���)^X䱹��On��"쎤N��a��f6�p�������^e�؞�J��,q�>�q�q�lłė�Or���;l�M��Q]Z�ve��:�GaZN�2=���ȶ�2}���4U<ѓW�m~ڴ�CWM�J�P���˅�s�G�2�_7�!H(�/���G��bKxń�9*�j-��u˂Rw�R"<�����-ت\�~v�P��k���Ul��J-E�g�w���y��}g'�cR �kSvl�l}px�8��I�t��i�bu��ϏO��i�)95ax���n�Cy����k'�v�]�#�S)���Dh�A�e��ݐ����t�/>���H���=Vx��ߥxw�*X�v�̗h"p�z��a�F9���G��In�J�w`\fAN�QMfN��_#�l�G�.U��8D��9D~>��V�p"�G�/=���Î�4߫?�u
Ҭ�AɆ `�A{w�f�K�B��s����3\1�]Ɩl@�z���ɮ" ��8ZD-�bY��������s�ܫCh�9�(���{0�_��x�KJ�D���s�yՉ�B�4�hn&��U���z�^Z����s�݉���Q;'W�!������.#,��"r@cQgWF�"���ߦa9I�'��B,���/I��m�]�.��x�#f��1Hu�����wDq���%���� :#���Ԫ��+D���_�Y}8���N�n�u	���x�j�����T���/v�
�\I�f��LN~U����P�Y-XM���=�4����|�	Xc�� �X"B�˪����OW��Kd�u�l��=�8ȥ�ǐG�8&���E`�VD�7��Ơ��!���<@��:�� �_�w�4%ZQ��}I�ԊLx�^��~$M�hזƀ�(��`'�)>�.c�W��8A|�? ���<�C�7�-��+�F�A#)��(�~oi��j��.��)9T�Dj\(�<��!npT��˛�j.�13	�D��W���z�����y�q��8G^^�G�9w{*���c��?�.ۏI^*
�o��d� ���Vl.�5.�,.�[!2��I���2����KZ��vh����/ca��0��6���	����Y��m�&g9�'�kLӴԧ#
��� h�����5-��zΓ �.,^�~�T�<6�6�"�qA���BM�H�;e\C���f���`'\��i�vYg-Q��s2���8�|iq�yO�z�Xe[C�n���E�&���f�E3, ��3�R�	��1���-ꤒ���pr#�����i�(_��,����e�]d� ,4�X-3�t٪L���1�:�<#�I%�S�g3��= ��1��7"�Iү'c����pA�,�{o�!1Ͽ�|x���a=��x��-NDNV!�"��米ۆk���&\�Bv\�)�92d#u� ��FIW���"6����V@'r
R^�y��/��I���t��)��^H�)Ff�����ǣ�+Pz
i���G�k�S�5�C�rX;�F����gn+a�O��_c���=��']K,�uR�CP/�l�C�@4����T��[�"�d�#&��ԗ�kuہ���h���a\Q�9�(U��W)B�}q��_R]�/��h��n.��Il��FE����#RV�������톲�,���ڛi�5 ߘ)w���C�FD���T�e�=���aԜn�C��}�q�jF���y�Y���[�]�]��{f'��Ձ�����iT�}@5o�t�\���u�r����XG{�:z��@Z7�]# ��`�r\k:.B��c�=��?��$/:bY��b�9�D�.p����F�aҽ�X��U�5牚 q��z�X�Kb�=���h�ףS0vW�5�$-�<��9��UjkK����(�Ƽ��Կ�!��� �'K]g>�%;㻪�Q+V3�&'Tl2QYC0Ҝ�����&�C��	���~h�-�*���E2���=~3 ��C75a�_9ն��M�x����a���y��}����4ҹ��T*��Fl�/���Lw�{�3g�wK5����Q��=��#{L]��}c#�f��d����!e��7��4�+鱖���l��a|�+�}�qs�Z|�A��e{>@�h�w?�Ĉ�^��[M��yT���dҡQNإ��Cf�s��2��w*��2�̬E��N���_� iS���?�;���O`�5�vbQ�&��ZMbj�,�QTk�9
Emn�b���e&��s�媑ߑͻ5��f}�)	F�B��g���� ����5��k|�X��=���s�G1���&��]F.f�p�5n��+J�mhW��w��'gɮ���J���mt���}r�i�Ѽ�Dw�R8�!J�^$"@ck��m���i$#�b���j,�M9�.�L�N G3@}�%9> �����x�0���(r5�����5��=փn_t�d��M���Q��-+@�%�H���H�`��ߣb��u
�U��D7W�-��1���V!�u(����[,�$YP3��w��x&�R�ȉt��#rS�q�4:�+ &��ĜQ�k}I;w&�bG��`�<]P*ٛ���Y���l��_�p�
�s�I�ǡ�W�I��E�>���
6,{�8���7�Z:�Ce�bb�&��F\U��6�$f���% �&n���&���O�����dyف�Q_���_�-�2�
�s�']cK_��pr�v���ɝ*�hA	�<�,l��
^��R[�Pa$| ��~��kwR9ɉ�YO
bǭk��!
�(:���%��k�J�x�y���uD�:@��]䞕�Ŀ��^���@�÷��9#���DS@�w�'��C�AP�򅀝�-O?b�q�kܓ
3�����Y4*�\�U-�<����h傇B�>L���;��}����Xs��dU܄NY2ՔRzA�$2צ���f'�l�!�e��`� ��{���K㲼6�����t���9�o�2����k�
�Հ�����q��`6Qs�g��R���Ј�?\�B�����~ҳ�s�)\��R����v��z��66��� A���ծ�H�*yn�� ���Fw��ɘ�E}�f�������� L�