��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�'�I����:��O\Y���QS�;���A�HaWլ�9"����*�V���v�4�)� �f$�S�'O塞����G։��Q�|ݵ���AhQ�Y�:����M�h����8���� L�(��df��H�j����"�fߨ��2˹��w�*�:IYOy�/��6��v�����3T�S�L��6纀dҴ��K0X��v���c���2yބ�{|Q�T����1`1�K��(G�����j�+e�'A��g��[N]K�rE\1���dl���S#՟�w��p�g,��$�Q �h���q,hvԎDF��^9S�Y�x?��6�gzsm1��)9����6���qh(@�X<���E8�'�%�$UC��+�!#��=�>����&��ͻ/;Y!nY6�a����%�`X�9�PaGh�M2�[����?�Ih �c�&_�>e�"�^��,̍ċ�
iwv�k8�����l
�p�ڻ_!#��"yX��i�u)G���^X�����̶�5�nR����	"�F<2�Q�ƪ���*ԸW�T^k����M�jڕ�A��.�\�� ��ks�������--�r��s�!8�o�U5P�`W��I�V��W��ɝ���@7�"���"/i�I5������(/�<��A�ǲK~�\�n�w�(e�+���·� lw�}�s��>���货f����QPo�2JRh��3ހ�����-����(c�+7�tF�rc�T����^���D�pZj5���No�Q�ѵ��ZP�@�2.ɌxX��(��"�!���4|��]n�H��<N9WWr�ʲ��f�C�(*�qM��92�n*��o�����m}*
��]<�k4'x��\�ӧ1N>FS��� (=����%���m�XHdy󚌃HaQE8Ѝ�.-���Fe��ө�%�<��~vHD��W���I$���z����6R�L�#�i�#�)�8\�+W-d��x�hXT*���Dv;W�>��x)WW�(h�k�
�ߌ��1)��K �;����ɭf%�d�õ���q.���2ђ�	v�<��-��@i�t�YD��my7z�SM��p�y�axۯ'��SB�_�����pZz��PM��oP�S��|z=��l��"�]\�R�MU����A�DG���ɯ�3qz�=$��`��x�8)!4r�|� l��>�ݛs1TW�:�Ǻ>��"CP�[��B���b#����jZ��qŋ#�@٦�7vU_���JЖ����gZIui������3���h�c�R�F��5|����Љֳ��Fa��qR"j� 
π�������;�t�%����3���L���َ��m�vH=:TQ�ݖ"��P�a��;��[��k�6SԘV@�!�7��ڠW�|��ßp��K$�������3C
���1r{�9/��_��l>"S^�����{t�O!��m��ظ��sqJ��E" `Y����Nv��1ĕw�8Y��d|(ޝP��q�`rXHÛ�6��JXSx-I~'X�^��$�K%<�0Q�ģ&s:HE�+b�oj�u��b�9�c�����f}0S���M7{��
:�d�R�Z���H�w��V7�?�(�L�6���Ы�q'�W/�*�mk%�����,%���������|Q�J{=���]�v��=dW6ӤbːJ�o������������˵��cY��D2��~B��v86H�"�3��ǯg����B���jw��������
�z�S��$�8�eo6B�w�.���/��g�~Oi���߶(��Ind,#�J� ^���4����K� ��70-�x���}��V��f�ɶ��h"��{OZiN9�����2)z�}�q�|�A��j-\Us��̭�N��&?��O����i�f3�朸BO�l%�=�f��;�ǎ����E[K����&<�il�������^�����$�L4	fVf��m C�`�h���t���)�c���R��+�����b��pz2���24��?�|u�C��Lִ� ����O~G�Ֆ��R���������Z-Hv��<r��q��7`qF�%�'�\D>W��r��Z
!\�ƌ�{��t�u|Ԫ�S�@�� lj�/�Tsg`�+�5�c�\Ƒӕ�,"��WODu�4Y+���f����%��A�|*>!7	�9��ٽH���򛎐c ypA�|�{	h��s7����?�7#�'S���k\����ྱ'�����rRC�(���}��{h1p����:�݋�--��.�2\>6RJS�ʃ�6U��#�5~\���N9	3*& T�y��y@+����}(C�nG���%��t�䏵�o2�)���yz�-<�Ҥ�KR�Q�4}dioO��)�\���&qh{7-}D5� ;>h8�Z��� VgI,��es��"^* �W�t�xE����Ef/3��%�|�F�_̴
렰��V�7,�H���m��ч;��-�s~M/��Y��+Cȼ�C@Yj�nz�X3o�E�T6E�A��XNeE��!�6@?��h���}��h���`��%��~�|�,�YY��3���H�%1�E�I'Ƨ��!�ňԱ̈a��h�hW�Je1�8�(R�Rq	�	H��{�\��r\�|��*z��w,��Σg�=]@�:�T����l`ا�p�z8�	h,Ne�Z>��5V��
Q�w����Fl���jLI:<���*_đ�T���}�k��1�	6S; �yX��5@��&栍6%�#3�a�V����_LG�
_�t}��F[b���T�%��(;���:	y{X}�D����[����nw��G����(���
��yZ��=��8�"�ԅ��Z���Nz��lF�\�;C;�bW)�6Լ����p~�
SV�ɉ��x��gie���@?���֪�X�ٖٓY�󸰻d���q�/�?��A���x`�h�3 ���kc,�s��Kr�ۍ�=/ಝ��SA�w�q	��g�u^�<�p�k4��S8@��s����^�o2�ҫ�
����
�E�O�u��ۥ��O��*>����ڙ����L�b�XB'����G�.�������P�`�[�7>D[��`� p�%C�Q�]q*r�N�z`�k��84"1�)�F��	�9�2���,9�?Z+`46����`��]�����	u:�U� F�֝�)��CK������95$#|(9��,ID��7�Yv�I��k�*'���MQ�]���S��Q6�-����f{�d�nѦ���0dt������ͱ�:� ��Q��T)�T��߿`�?H����z�0s�F� ��"կ�۞(����ð��EdY�bk~^��MXZ{�����Q�α�Uj�ըL���ۣ���쯎�C;�p����9�ꀝs�g�l�{�{qH�퉼��R?<[
�������	����<{ �i%��T�.:��wގS`W�'t�nJ�� �ىHQ�s����kB��3L����4��U���L��Zm�$��(l&)(��h�ʃ֑[8�?G\�D68ژ/�Q�*�D|�l*�Y�kT�8��DO�0t����Q-�pȾ�s\�)�E���k��>M
��Kz;kɰs3��IOX���İB��&�����@����H�c�iV�|�Q,}b���i72�nC0}iU��|�]�*�2�H���b�5p�,�,�"f�Iʴ�2|�t�)��_�:������m�~����C4p���E��8�nہڷڎx	����6��R�ާ����~Y��ƚ*��ߗo�L|E�1K��]�*��$�+���`�rN'�! �oh,�4�:�W�viork���s-�a�	����E̼�j����<q��aF;�������W�)�p���f�̓�����zy�`9�>
� ��9�4�"�N+/L�uk��%�Q(���ةc��Yl�Rh��L�O�0D�Vz�/�����Y�F7��u�ӆ�P ����}��@}O7���a�GOHg-��eO�5Az�%�l��N�
�l�w/\�l����Ž�@X]ɥ��ج�L�)���
�Zy�����O�e6�9&>)���-��U��\��$"!J=ݕd�$��u�Qj지aY��$�~�1l9�e������>F�~}[o.:9-R�8;���=I�n[�_y##E6��J���%q���l���������[��.d@x�_T��nm�Y��*���:�E��'����~+`�����y�H�xL}r�a\�|R���7j1��W�ཻsn��틭�af]�"�O��ı��C	~�8�q�^n�����������#+(�������z���/���YV��Δ��	[؍!�l� ej�4�17�*��:�������:�7z�.��K�m� �Ҧ=K��'�v�xA�/̎n��#[+Z.`��u���R1-���Q'�D�r|�3t������G��ew�FE��_2‘4�Oխ3��`Zbw��z�G�Ǯ�O���v�:Is�D<h%!�sN�������<�(��.��.@SVӚx<.������9��L<)յ٦;���+7Y_�/aoצ[C��1�lQs� �w��L�s��3ɭ��`_ �:5 $��&�S��ǂ����z���Vq���[��������~n��`��,�ݸ��������l,�<L���\� [�O����:��9������q;��F�ݱ-��H52C�K`=��U/v�scc������.GT�2P�A<��Ι@Vw�!"�&��$�<�cZC}������<t��}H9�ш]p4(ʎj���?�s�Nn�jY�ӥ��K��p7Ts$f�C���ب�4����v���:�T��dKA�ŕ��噬�����������͆�
��"�rw ����E��fC�W5Csw�	J����16�c�6�@��j�8^;�X�UA�(Z��ЉjVw���+K���Ny�ǣ��d'��[@o��8�� �ۼ?��k&�vj�U���y~f�VZ�6�Jщ��.�;�?P�_���C��h^`�=��n�T�FtWT��a��"�T{�s�^��8۹#�T^-��*�����E(�1�!�C��y�4l;MMS/\��*����eM�33��O�ڨ��z���if7X�k�O|�K[�,����k�H�h@�L ӗt��좪?����:(.vf��Ga�{���j /`٧��^�������Z0�0��f�ԩ��΁ĵw5M���Mȵ������;(�KR!�T����iV�e\����ޠ?�1^
L��XX����1jX��*����iB�keZ/��sa�1�^vKt��u��s���+@4?H��D)[mSh��xEz���M&�`��hA~0��G�oԫD$ӓ�U�*~��=i|x��-�l$���/g'Ƹ
kM�N�f{��j�&DY�+��%�^�<�$���fB���b�I����RT[�1A�gr����	"���U���� Py]t��H�a�I&r��F ��/���s���Ci�>
�Y�T�<�� D�s�f|^�}l'^��_6q��y������ԝ�X��Ժ���uф�M?ѾϒP׏�R�#�V1��?�����'A��r�l�[�� �C�-ı�(�Ƥ��b��W����o\�< 0�������	"�"H�I��m��}�!�8�	��o�ڪۚ9�r�#2KQR� �ζ��8 �.hr|o����1�'{?���U���p�\��چ&	��at(�տ��9�����g�'�xv֋��I�i���;LW&�Q�V�i5?�8�msme>-ľ���ku�b$��D^�0��?p�1���ݸ����$��_^ek5 %�7"{;�v�]����R�n?Sm���$`׾7K�HC���mҍo<�Eۓ��I3w7��O