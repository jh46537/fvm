// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DJCyWyOUdtFrCGISHCjST2vQcneDzLb1luOEqxw8xrkNfJr/V6Q9WOW+jtnuiUbV
Wa2DR5vmMNg0ic9jOfroUVwfxtb/Nvvtc9A9hqY8eUWtmwlSpokhyi73yCLNoaRT
xh5wdXi1Xsd5R6fXOCbaFJpM3H0XAz8pKnR69etGSug=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 324752)
XxZiF+Mlrdy0/bDChsk2+s3xHEitioU37Sz05vfFZZ9kdrXz4ApTu4Kg9rb9nBNf
CocRzeJpTQLnAd+oxt4oKKTXwwy9BuFYThQd9QQlxBEl8lEuG7tfru+6nnDGuRN4
u8+7/4PBs/Fsz/JMsIEyyo6oGsnpYo7kxmWUynhUIKsfZ3nFmEFWqQcOXCaBf039
zAnY/5YIBHsyEOFGWwX9pwVKYqu8lk0t5Wq0pWm6F4sD/tNNZrjTD3zP22mKEfvi
DDAb4lpZEmWnX69LDYpkwK/i91sy4ZM+U30VvEtpMH9v2aiHA1Ks7Au7KE0zxV3b
UibJj7qHzF2YqVAcURMO4+V00I1oR6/FQ3vPAjnzgS1ugTLe8ldpBSs3ymOrMg5E
ZWK88WfIDCogjUDYfQSbucTKb0NPlHL1Wr6ZCLMZrYmSsoTmy6fkcQdG3bZzbNnp
vCKeoPpvky5zdaiIknXoRBb8/Zh/hgcSUNc+xmv/FLONc4nYk+nA9PZtEebxrwEO
uwfXu8t4NNYIN6v8nMSIKC3QePsOP9t63cEN6hd9/p7Y+8fnGBmU8BJQEwSZFg9s
ERTRIUXuZcbgeouXuRdWIhYFBceKJOTgx3iCV4GSjeC9fnFvU6XznWKIt6fvtN7v
Pldy7ymJLqnXC6+2yl0oWcJB7AIpuaSqJ3Zuhiir8FEjAL2Sqk3+/NNmt70HxbwK
+U8HLzNj3Ln4QNDGb02Gpv46FqrP0ein0wQYPWKhOQartRXcTUtnemxEJEtzIW0e
wnexIhyIzsf7f2UQSotvVkXnaJQsOYYSHf2/z9P9x2x5nxT51Igvke84XDeg2Fbb
wduk0gekL4iSSQXdtXsmton3CFGFVW+7pN4g+4uJDDBZMmZix5li6zYEBs5lXpoB
Qw773Ztj6PvwcOnlQMCiC//JNZtOpeK0S8XtJKoiuivsGBs7Qa2Up2AiCECw+raD
M1h+yN6+bAkQbDHq7utXghiW04NHnJyc26wveApB0HSo7HwVRsTh8YWRYsYL4xs7
6ONnHiLDE7uAfhaF9dwCCq6e+V6K7DJvDbAsaprz0C2Dl42n4vyHxLvd+aNoUfz8
bVwGkSI9rldixPk19B34PxLO6lfYwAvfcbN0JTd5eSjvh3x5reUELSnFxUy/IrUu
IeA/7VkaMxA+ZTeCV2Ef2sUf0i6QFm/hgrQfH/NL6+rJEPCVdzgWmqZCyhdU8dlw
eb5p8m/3jMoHrT0sM9MMtrL1+/a3sSVCGq9W0LowcX8B2+0DjhHNZ8RoRDIDPJ2H
dauDEdl1/MCTdVaIMiWgCdsg5ltpo1opd5WuUD/IJ96EwVmnDoTCRmnKuju4ajaT
oDTf7j9D5oYaEbooA5Fs9bo+MiqV4kN8NDcc8SK3o1T8fGXhJEzdzrWb0196G47Q
emfY3hANRMY1cYvGzylYxHWi2p7AojCs5syxq0k5tH6mfyQI/LMPPkTdV3SfqREg
1aayACP06Eo1nwHnC93Tbs0zImekbhylTpx5Q1qPZasJUb/yqMHPV2LwiJfyjjUX
u/ok0UHlZ0fAIf6MfMeU8CkCKPLHGHKIoQxbWeWB6E620W/xdR/vRByUS9vYKYtt
seg8Ki/P2diiUIbXJzDPyjqubY7uhe81yyTrOjBk0p/xP3A8lJHH3zjyicqQfbvO
h/ONhFMBzvHacb22OVC3RBJ9EqpAO0RmijGpSDQgmK4WdLvW7S04V+IQr8xOv8ZL
5rfKSlk6Td+lpbr0OPylvuorn451GWm8dmIGk6ZwMDJDvbY/BJoY/NgqRdVzgI+Q
WjUogXOlhYac/Fy8YA8X9WFG9zT5PddLBQtvLjgJdAAZ6N6tgLL06XVb7Tw8Zga/
8xIIUkDgiUeTuFpu5HDjyvkYpDrI43W4M6cjM8QGoMuIUtQBO7anFgN/Lm3cPLfP
1h0GR9lEKC6Fr5pLTxUdhAZvFJL68wfRyyzbxHsup9N375C6qyVA3nIAnmdQh/f/
in5uOXDgBdEvEB+cj/B8u/st3WtcFPrW+mhxXIsOiZxom6ExwIec71ZO12Em6Ow6
VWPsfjnHCUNX4rYBoEg61nxWc+4Wnnpn6kI3lLlhUHqRt0gIuLJ48dRgb22XUmXX
nOZqZIqcXgdaY7wly233TbI3rTUZt+yECAehVhqHKif2y674aboAcy+RFIeGaGGO
sUnBO4Ev7xkZNP1d5V/Kyn9eU+8Bqgb99fbXIyBoOT3yWyxhpijFhjiXMCyx7IwI
QHvf7976ErRCvHBd2e1eQOwWHrigYuvD4A+SiXcOVAG2h2nIYlMI89UYYEZBPLrw
Xp2qbI+aRP1xSLQozZD6jWEKYIOHJW5GgnQtsR2cEUDxFRsUYJ6IYcY6tUeO0zpl
Bnc8LfYpr+zK8RzDRtIlmldaGkxMvQcr2KOyOf9U7hZ0loBYDG2D8dCFD/WhCyvJ
h8fjwWyPwD4EeAI/ZEhBM5POTyEJI13VhTqldl9Ze0iv6kL7kawbPPWEWrqlVgC8
bTQzR3Ae6jfyt/Nsn4se2+ZSKb3Kzk3ZRjQ8eI3ernbxD9A8vhwGXs5ykAaGUG84
ZWSfcXANi+KerEv2qeJx7nvhuPBSYFPnH5EzYMIXWB/F0JyHkteSUtZU3JTRRYFm
CF0nxBpQ3tLRhmWLTc3bhhgfzC/H1rkI/QfnbbWBROlmK1rMa4uPliYFKzWPPoFm
wdkdSYGhvXmp29UTHbK9o2JjGlHDhaFL2qSNXf6kQx6iM9rU8eUBKytUWnJiR+eE
HycQSCPP9mExeOEwilGG2ztgVDLz42ahBjmvBZ6ibZutXqBANi8aPZvz6S13IXYg
BXQglLimBl76wNn0zE5LLJS031oxdGYG2Pp+RORvtcj+Tz3IKXHUgS4C6kQtyywu
Eyhf2BVi9PHzhdPWYSzo3WUoo9fSxRzUI7A/RVfqUgkNOgzScrbTLCGXyoapvW1i
U/6w/9fnCBVmlIATjUsnvqa6xcyHli2/zDdErzswgpuh/O9LzFiB3Vp64pDnhmHY
TBXAYSJI1cpu9ULzG70shH0UqouatmwdDJVqsgk7oyjdH+LIjebrIqJsyTH2gn4Y
anGwIZulDLkbBm2G2/f/NIXDhASA5mscvggztZ+LA+7vMJRpQO7xYrXqR+9SD1A7
lPEe21XeWhYZgd2DZBSu/EV5z744iYznc8mr6Z1WeXan6dKTC7NfmRAwy49CJwJi
DDL9gLkimjWY3IbmSytFDM20T3+doLC3lCZ+u6suksyhK/j9wwKi1So7dEmOb3fT
owscukCO4UMPszf6GNVl7eUlqdMmy/Vuh0YoBxcxQOOVmIeYZP4izdgxFB1o+Bur
Xlw31eOp63Czn1I/J2NljI5jArsm1uk5/iO0UBT7YXp9seJc7nWly9D4WEM32Pch
a3oEobH56w/WKWa5MKHGM4ZKCtWd4o42S+hw658u8uCjK0DB5rHYBz6weTT80CSw
luuBxhMpc9zESnMs9tZNPwkpbMTAsp9LTS8/u67psiUgTqzfLEKWQy51j7vveXR9
PskxTfd236zmuMbKKLoM2iZIREtsNuHs3RISXI6Kxcsx/wGQ36p8BvxMRCjO6XuT
P/haCcLWAv4G7Xl9JWVJLoiKPSjrmf4Jxw0pes3NHVbQzbyUQBY2fgnAp6bD+MmE
zndBENigEgZKLE3UEn2dl2rV6BYaCwAO/IY7k1b4Udz1YHIgR3jBHtJREB0eAntC
OtqUdflwwY+giGeQ+Yw+fLJPF8RBPtWaP9aVdMfB2/DurdelK/DrmyJbz1TAsFC7
1lRbuYjiusaetGAyDoi382U5V70VSHk2eKnQxn95T8Aiue3h2qazsTp7ks6jtG8d
MspxKIGmKV0wOwdBS5WhX1GHovW7U1qebE6p1GaEJu8xCJUEvX2R7maszXmL8B48
CHWmzwg8O7huPHQZvhX/W31gGarc/PytByBjHVNRWMQQHPqaGr/DYBa+MFpYIYky
eNHn5GpibroG+O9ErkBQZ03jmqaGOuJeBEFhIJgrmN1SXrfQl7j4lMXFy/BnCybW
CMlxuhEeMHM1zoUv0P0VwWDop7qwfvuyqLnLF1+dTWwlX4fnNv73E6kw0bLxpBKw
/HGcKH5a67twq2V+HIUlDNjGaU2sZ+Z9n8YGtJGM2f6EVeqd1aEel1fJU8TBKwuW
qr3NU4r8JweaZyMpD8l6eOD08hbSZtdEHqabWwK5vL352zZAQH6GO4X0OIU459Kg
PGnF56PoZeRr32MCiaNftxDN0JU2Tr7OfDmvQvOLhrkQXBFWcNL79srmhrYwMcS0
r/BlJhdPwsD43gpH/nCaz2wZAINP7P8p4MEm4YzcHq/xh2Tlc9CIgMHKhD688dQv
9eZabBfT930Fn+U0yHC0xU2E1Dxibrggfct+XQY/9VEos1S0Lg1rszHh/X1LrpeA
FKlIBp0pzqEx9X5gjBtpG9QfENoreSW2AGbWyfe/rIygKryC+EFLrVVON/pbvYAf
7AjiovS/KWNG3s2bP197PFeLD2N8jHexPj2oKJrKt0rVN3pqQxnHfkDdyYvKWOVO
o522mVA3gjWx31f6yDj1HE6d/CW0whBVYZodVGwdcEotHv3ovvTRX0nU4XZLwsGM
a9WfCcKOc+giz1kjszUQCpNd0SyeyulWVkJCaZMZTysxzMVjBbc/itvy5bgTwUoZ
GwUck7opQjD8i3Ws4XdjBjUJF68xEaGP65/OJyQ/XMTpeM1UL6Xux0NfiBTLSVJ5
00E7r/uJuDjp7AYqckxaYXTKf/4Wn6TFWa8xBFLnbC9I34kgqk2W0Cq0WsFuJK49
BheGywo0BGaDJYtGALoYirMRMlPGEGRUArjF99uhDG4FjOfCD9CXnSy4Km666exb
HqZC7xF680h6g8afiPFSsWx6sbHVuIZNQmzYmtNak69aQwS14bCTKk5ywfsEGHeZ
dOYEEztUbzywO14O3yV2lE7LlkQR/StqIuwSB8yXTN/385De6cHRVwZ4+jxiexFc
l/qcSbzJzoLty80dD49bjFJXFgw7s7N25+JyAlFH7oi1EyVkmo7iwwId1v2ra6pf
WIYMssiAzjoByTjHe8tEo9Sj9uhy/jq8d7zU20iAM3mZvfvXINlQodtRXMoRbFn5
oApI3KS7scFAjD4sVk9LtEeZ73XPjijZmm9fLshU9w4x66zUV7t2SAp8JqvzpJe8
nOGYQ4rgPX05TFitY5Z3o45TWhRGFQL0OzH/0QZDdNkLWQc6Ss1r9Ed6jqZbZzRs
uEZFcG5aLipiAgQTXbYe/Kxx0ojc00lA3dszpnJECafGHtt8kq4ipqmOKs5iEWdv
2pV2bwJuqWrITCtZdbV2cNiQAU8DzC1vfWy4opbfbrYRU7xe//ICyR6yQOzkBWBe
lXva0yB+57Sa4R38Eee1vJwBD/oBVwNm4Drgg+eT7CpXGARkIuTpiHPW+xGvR6IJ
XpwYmgzkiJeIgQMEVRob2y76AKVSr0kTedJn8Ifht/jpGMI0dpYTqGoRtHCSJdVw
l6/w5edWZ0P2D3/mq6mVjGzZpIW5dkfflsQGnUS+dO9wX+BnaOP2xYgL3yzOAPP4
pCrC6Vb4CSzb8Zz4I4jw1GcoBfvKfJSlDTi/nY1+bIvP190UTKM3Nt4bhzUCRglM
U9IQweMcW7tt5Drlg2n+tU2PSp4ft3cGVM/JkAe/SInTcmdNrOMDYrYoDjyx2UzD
yEJ++AgibDsxNKeraQ7hQKB3yPoTXekVrd12Xoqarl0ZA9K8cKn1B+XGDPDRcjUS
AYzrs6XemHSQIAFYsgx8XxMT+Z9zIE5grpsWo5iDzqZktprgeuuGYNOBz/owjHt3
H5OK8DbwX4rX8KQnk3J6vuA27pK1SJHk2lx8C1Acv3XNQHJiPYOiUGsk1dt/X6I0
1/kupgvNkOp8NMXzkpliJrVH1VMYsPaMkacAvGX2HOumh77wk7XYbEvaPW/zoTGE
xUZSBgQdT27cRjqP76o14Ya8X4rAcA/RNlHMZoqAaLYZgxVJR0uSOLT61cCWInlH
wkUiuxx2dc5dPGl9qy9VFRueEBIh0MPKyp9G+VAWWxiAbwYfGtPAeuvu9UpExCff
nu5sQ+/0wVowZO+w6y8Ef1XBgJMwd/NQ3kq2SHYJccO8GWtsKkMoorhtb88EbG9h
Aru6jGFsAOH/WN77a/RJmaisEcSdstBA4nEkLK9h11lPBQVKc9aBrcaFgWugwAO7
hmsMKovf5O4lTEULCYFB/8acVQEqmt5fftfYvlbGk8bJ2rSMGD9d0Ak0W2/X69tz
jxcCZjEQxb5CUY9BDHFYUMuUF79e/E6Mzmb7Es4Ja6XZ6kNc6r3bQepXiT+KrL+9
nLzHHOUcS6psTTUxzTQOIHUXk1iYZkxtUkeM2wm5vAvwI+ko1hnwSH0x6ws0CKqU
D+fWPlJaseFY05BdWW7Ob8AxLOmkDcZBxpCp0ix3p876iA/+aRorQESNkenaAYET
HD9x8b+qcr8RzFTPduOeGH/cGjhzOmzwgiowGVtZAurUsd9F9byD7KNziKqPEQvZ
KcJ7NBO6lOAt7hgcV3ebzC7SJfstTNj/QyiGBKz5U1cx/NEnSDJIuq2i8vPkJRJn
JhQDQDUHyrFUXnuS241J5XSaQzviFw8/4lxkEzXBnK+ZgAw6DLkCwljA/VQp6hr2
l5poMJ79m6xsPNEc2lI551XjZxCioRPt3Jl4T4/jTLb9BBIyW61IYN7WghIJ1Dx8
8SlG+dtKEvOiKJiJVonkpAlxNEt7HBL+1J62eLLDqjCTN/6yIZyO8UJVE2E77c8Z
NtTepXct56DtkcjGJIRbphkYdUkTYreU+2M9MDC2iw21xwHTkFuYCUU4WyZJa8o0
CqvK54oNKb0HEXg5gyZ1FlLI5bwCvgp06zYvi2yfZ6ZJLsztj4RPR5sPkv5/AAKP
CtNVT3XcKyUtr/KWrdltg5t+YSDygZNyiYuvkh5meSY/7sZHix2AOtyvBus4napp
eS/Ne/emobPuf7HbC9bDk+RQ9cGnxCz4x0t1Nqgp82wRhWjI+QmplSlN0YZCJT08
9AuzS7FLLGdb83qKLN7hXw6vWF2LD57dqUcAU/Cv0eqRrOsCkPzycw5WzFdpCiZU
iZSrEpDJdbksG/kEIaE+0EziX0ebxS1khAIl344nqLTrARry8pXe0nqRpgiRCRpi
Ea/et+YyGYoKpzlbbbCUaeeheReDciWQt2dsRr18V4zvQvaxWj7S0ZT0UT9UXdWW
lSR+GtqGpcLJo9fk6uxfSiXwc07SwMhqOZwxq8MsVLftzTKYi1ixkSg23jAW1S+C
IP62+4n8fndXzQLfN4ZLI/r1dLpHT91xYoYj+msLiroHxew181tXG6NnIptce/0w
dRJYKRVoCUybpUEj+NumKcPrJoZc4JZuVuegZw012CAF0SD7ud3SjbXxBAYYTHSm
8puaWCUrEk109mcyVvNn9uvBVm79Lf29dpA/0D0QD27jx8ys6i7tMXjbWFNFznKe
aHhWmQls9IjjcuWx7EXLJ+p6d2mxPd26SY9jKWTye2QXZx8LhCQdyyaXQEN3WGzG
ddo3gMlgD20tUTtTOR8ELr/PCNoNheH9++AO6KrVhyJaIWmcb2I5MQpYaiPLW00P
BMGecQ5MMKJ1XBlCGQFkyawc0MwBRE7U93QgqGxWPCi2l5E0Jw9EU+awbE584bcD
XMSvAApCYr72Vc4W3WUba6FikDSSwo5Ij7RGfEB4udZQWlCIPstPJQlQdFY3AWmn
PvlfKVED9wtLjzIgGLPVRgm3w9hrRR7Bwg6Zqc33aS6yf6CCK7CmMfGc6/NZCtvd
ZIIpOaL7AKJuI8HWwCNZIExFOnIwfjQXvGpMVjwa6imDPVMfvaza/TgMOQe3zGwk
FsKyNtY9qOyKyQUyrTXzJikRgbMKFPcCxmCFCRXPcDiE/jpvDp0De+3McKkmM3Qg
7u8bp5fITndXQNARLcrFA/J+XsQvAacXf+LffHgNN+uPlPubF9DPhOhNiYWK6k/e
KPVMT8/Qo61vzGjNgoRsetv4xez3X49YxHlYhXRrl2+M20QhlOnh9uwtlrRDjkXE
/7ajiKKa9ChicCZJKUbMZ60WdZXlIzvzuFZqwqPz2HS4159RCkBLbuCTX3lLAJzV
3zRRG6PcAmoKvUulIObdBw4QPZJykWDC5aJUIy2YlcjGH7tUBbcV7kKBxDn1417F
NazZB+GIGrEvlUCIA9M0+HrCkynbFQTzjAH5OzeXjwGZnRCNb+g09OkIWC5K6iiX
i2+Ut28HS0TqAjHhs8fWY6UW0/pUqV5hHHjclCROu8vbKgYn9S2PNF39OgkmqTVG
Hk2xT+QwfQ7lcFQjQBD/9UJ0PojlUCHDjGCAvJOYl+ms7AIi8Porw2Iezd/EjGl5
kkVEqp6JVRfdynFMAAHvV2JJpNZte/2KI/wDpSBKjnEUc6POAzjP2c6TLraVbHmA
ac2I4991OaD6RNfUEDi7R5A27lyAna+3ph6CBBWBKEsL6MROd5Q+3oJ8yRU8MruG
DufGtpHqSWr5qreleuFgIdA23Ln0WfbeMhPTd980KS5ODr2B32g5QTDSFe047TIn
Mfrmf+1wB9jtBJYTnYLRqs2L8VlVOUYWMMwLW7GYIgblz5I41FcPGALhHEwVaJsc
v9c/VNI2exsIFre7FsviXrBXM/fUaQGQZvSv16k9QYx0rQjoRgIlEbh7df/pI73W
P4JDXqXJ90IW6jEHTXI8KNN5J3mlQkfMtlGHdW2qHaTMxMHyzWo0nPWYc9My7o58
i7o7MIXVZOhy6NOlaxskZONJKlTisZ1PelNOFXtKFXe1YZ6pa2Y/EGA9EkZCfjo/
OPQ/q9geJBHB4PjVRogCmQxn24lsRoAjw1WyxnadRyLoujCsbtoP5E0BSCm8CClq
fqSS3pm/GIcm61vB40mkfmHZuWZ9xlSsW0gtTx0apfRZ3KhgeBfvxFLHMFEqvDA6
khgtjgnXWIj6L4Xk0VrszDFOhvpQTyl+M+rc0AHjfWuVeGcvqk5gHy0rJhegXRAf
4wyzx9xwZY6hzTBGEssQxZ4bXxZj1TsxTdQLa2r2qhXdIo/brYb1wSCSajZv0D05
A3lNhwn3z+zjj0CcJekwDYtjxnhgk3CgX2+GDtmt3ssUBtTrWFUgke4Vwtn42+12
JH+K4rmhy5Lcfa5g6NZjxA8PSMBErk5qAB2TF1+FksLblSasPLtolTxmYcdesZSZ
9vATB+P79/2SeQwOnTSiB/iPsKlY0UBpiKQvCnco74Csvg1BVev/CNQ4XtYc3C70
GvjnGh2lWXUs+eCHIiNvdh6l4p7Q3e8mjibgt31e5O/dB4ErXpIq9DnuN9HYaRDm
0lfCe7qU4AOjX0H8HGe5uEkLff3saWmw9uUvqlBls30+571pDSKuf6u/uvqo+XBK
YDEKszWidQG83/nGR1NslYHjE7qyr7GrtTzmbb8dhfWbfw8IxiieE+6wKjgWpE7+
q/9DCl3xpnZtHAAa+QZqw5d9jmHfX8+NOJ3rs1dZg+DkVSV8MYNJMhzjzhQ3V184
KrDgFnYJskkt6+cMLujp3PH3vSR696qOMARraK85t6fg5TAR9ajf8G+9nuHe7k5y
aFwPEhg1g1P2hhTuo7rtiv6WUvE/PvO6fpTwMZTrxwy/mK3VJ2507hYs4X/I4JvJ
rTCvZUuR0iuQZGuQLNVz/6GZfjiTQ0UI4tg+G64dYZIcbRffgJg+kub8gN277Ci1
6SmAhxQvFFJ/1BnwH9YDzSDWlb9dy9KQ4w8gw/HQ9SMrMplExXTxDGYGF5toY3wQ
VSskBpVY4KXhkaAkBLJXe8DwiG3FO3F7YoFTChSff51Xf+Y4vVRiTWbngsPNAj7a
/HbXmJYNgreGckXjHMb5B6yW850ysYvsMWBVsMZlLWGQCBmRApwmKMI8EXgcyCeF
k0Kr2Fx+ku0dVF7eGI7cccZLtlumQH6dr7Tek0ub3GTw7SlOy1mFHwZMRA4Uu7OT
asf8wWFn9iT2tapyLMN1otBF2Pj/oGJg79Hivqzk0IOdXMPEYca6KE3GJV8Bwwgt
xLrqoQoHOd0ZfutUtGvaHp6xMpbAhvaBVGq5QAZBILYL33mfWaAAFnEdfrWJxLRu
mkH7M8LZw5Cj2yBvgzkwgKr4kSauYQ31a8VOc/cBH7mqZlbn4QFA8N8Xhk0mirkq
sjjzyMuOXsOiJYW63akHw9SDTAsDiGjqA+GA/fsONxWvorxdIX/r9kuCuyTg/Oc6
EWsFqNMDmRxIwoidlI+LY3KqxTMrR6IS/9y48tSg4CNVyXbK1QDyXSJN+8TaB5zG
MABY/xBHI+BeoE9EBHEi2jSVYvWtRG7+m920QgdkW6PENR4jWCbNlzcnbTwT/OSb
GCM74HUppha/rjSmvVUAk9oERMHh2gv/kItuVpt0S9//P6Yli+swm9k9u/EEaWDc
+HoN+YcC3Fc0dFpq874R2CwhKrUAwM6DnoCJd/ND7/Vwm7NFKM9Gj+RyFE7UbVIf
KuWk6a8nWp+fQQwJ/f6n/8o29R/A8aRW/cksm/nciL11JDIfZui079Rrvx5cnnhv
pOPR6j8z+CGJO06rTYPbEWR0lQjcka1Utg2ZxkgRVkzoGuJlLEsZZPOF72tMH/GD
XCaFrwM4+CvaGT65tvFLr5kw3xWZGHPyNi4gOOKyXEhONNCWcrehOfj1hevNa+dT
yimGFptzhs/icjtBu4L9a/PfH4y7OeOadGrm5wUZVEgxyaIjiyEegOK1J+bUFkTU
eEvhbylTrgAiZssVf7WnzvvMJwE2g00w+seVK6A+Pjh517myzWqBXpn8mIktSX+J
/P3U4I+Kiy3Kpo0zOB8T62lu1axxsy+x3mNLlRc47zFKZotwLKmYe+ImLFSVL7W8
kTcsZr5lGterFGzIPzjJXK67lloyXEJOzz6Rx0+FWTm13JkksL864FjgsfipIf4b
VbVltFCySNMTULAElueny5sh72s+7S41xhvlmeM3K/YYANygsLWt4USismEdu0cn
Ifde4BIzCBKlD8m/Igu/13djeFGPCkHATc48x4uaC/mQ3LSYt2+S/lorrqV501kl
eAKLeOrpmtHBm3UUnkCyHNbjxG1IFee3IL8gjJqA/5K2I8o9s4geyVEEa7TXrh8V
P7e3ODHgBOZzvOKVJb3ZvlcvA3vERrHuITDepBu1ZbMDvKtCmlwsM7372fuR4NPJ
2yOxhZ3prCVz+9qddf04EwlQCGtskNOllyiy8UYCtofjLcF3layiZpYRsmUwVCp6
FjHnmbhfj5s5jwa45hgjHjJfqtYgMGadTcB3r9vbW2FaQjJwMuuYDcJjm31Qz8Kh
CDZ4A/XoUDSmUEl82g5rNX8gd/jCea4BNa83Yxt6zLeaftWoWX84n8QRbJp+7suy
RP5TcT6YLfWX2bVRJxZBjjDQU19MhsGKkcYLLiI16fsxn83ovUts/aUxd9SgCnBW
oP5lycrbAJKBBgrj4iDZZ+DuQn1uc0vW7I+oTEuA7XCej+k2vavIPUjHebdhJZJs
M6iIo+8ZJ5moqzLDEnMhyjZB2rmBDIqp7Eo3SjCJsJGQKGIseawiaLeHIyhmcvYu
KwZrQVGoPAhcud0ZR93ir4aK06735lYrLWrpVeaAcsB78kSdbx54V3elLvivIjI3
5tz7zypxlub+Gd03jy0kttjTwn6z2h0XB3Jk3EUxr7bEHl7HBtqLXEEpXTE10Op/
EQKg3NcSHjh+2hlOB75IuF/88DhzMumXtOrypE5Xt4dEEs/bSs+0kBpjzyA/8bE5
wy1tTS47WiptGjshlHbHSsnsS3Z3A0cj7foMhbumqgXjPRqTJnYoqRG9yctbveQV
VMG8CtWO49DDIUwIWsmWBbDJd0xF5/9+4vVGvWGOdwrcATyWS6MOdlxSjxSaO9vE
KxcY5QU3ET9SLTJvjwNrfhiLmahKae5aY8SGD7D6P/CnF53NRf53zRcI1ObdLh+K
s8UgB3o/Bxf/hz+TtS7gBDNEefB9ttqODPTSIBYaxtjq6OXFR6gp6fPQa31Vy+RU
kMWpV7rbHyTojI0eXbXdK1TQzLDHafGkXTTwTOhKQW2WSYuJNBQZ/aud6jlcz6em
sZXeNPFxvrgFktlzHxUffSHsFehxZSsLZPLXzl2PHkh//7MYFK0umLsRHYks7Hig
1zHG7wwkLUoM6oLoTfPbfYmtZTrlu0DypIFXxpUujMZWq9JJPVTV5IQoXMM8nHtV
0t21NiKoYs22We4xxVdYV2u9L9oE5anFHBuocxvOhjkADGg+pZqCo4DhaRofW/XO
8oMGGCt0KO+teNRjpA8EB8+ACRqSEQWzlGTLPZnE5Iyc71Jj7OubnIiLFajR3pAJ
i52KgMN3dFXDnB/KkIaVmXBdvdrWSkNEjbQkVEfhE+VsE6RM2KkYVTKm1yILjPrr
8tbN8jJTC6dkFutjvjmKLxlr9EYIG7UQtnF1HWiLXBikcZbeLL9u0vYv9w0rGfBX
DZaFAMVz/aXHKwJGGEqNeU2vkdztT64eNQqErBv1s3ATEvYP6GVlg4N9UuUWvefJ
WzNr/gPMrkL+UZOsfjJIHGTcu5gVtwNVrMmHRMUzKfZZuBWetfbzP1y2sMrsrQr6
qSr/+EEGkcECJjaw3vY1aC4jH3t2AQUfznA2BKN880yr36ZsenSel3fg/pS8VavX
LtdGWkfQGBACXrLVR1mjQ0J2xyDoaCzNW9Hi+c57k9EZHxaD2P6sSXt7vlHx4pQE
DEKlpNbQAUXy3kWYTPd79/ZgB4pAfPrVZkEHQdMWYxttObX+6bF99WHjM4jv2Ve2
ccHc3blR0qPRocsyncT8wYsFJcpz9Gu2PqbumI61MLj+yAaa93aYuV8gpVgop2lr
OVSooPdPS8SpYX9B2wzrBYyxjEbx9GzA6O7gqPafM8egCrf8fSBfWXbEqXMHxjH5
GtEWdENa4t65+SIEc92WI07JTdiz0cmaimoiPbdCp9V8BwM2ReX3MojCqvGeq7fu
0jokyWz+z+oeLli/X/nix1vKFyfu48pmx5tFjJ7dhxfgGKq6ladARPt43RJJESqL
hhlAEoxE0QSgQo/F75L61/DD8wR58VH3JRrzMDXPLbMnE3d8v9LdhIYeNXbZ2Zee
99/QjTXNWUxQ1PpgvnAWegMmgxAEnG491Kbee6Ad0TibgnmscjBZftmfjmc4w9Gt
KUEYR3KsbvP7p2cVIhVGnVXTp93Oe009w0VuRE6QCgTz88UlhoNkp+oaD3HsU0Mf
YdT8lomeerfFes/gCSeGHbpqNB7ItvM5OrsCC785TeM7HVvAyhe1fJxn3Ew/hw/i
LAeufeDuvRrGfvilq+242335oSgM8PfMqzWNC0YgWKDj+XtWJKfCevgfDo55sgEF
CX8AN6mLCBPJh6kRuZa9ECW31eQVHDp88TS4Mpl99+g9NXhGrGquQF6Gnga3KYma
rGylntXxsAEPxuA3Osz6LLro2k8dtVMU+XWdOr2PZLSSp9OLlooSnkKIk8AbQJ1S
trX3OuwVpLqXyahAV8goHee576w7J7cZ2UWYNw/HQcJqNyHiXWGV9TNsnSAZSPoZ
zcDR3ZspH118IDBP7eTPq98kZ3QKB5uLT8lKBtllfRDJzGjG/KYEFLaiOJkjncm8
jQDgYQuanxyfCD1WHJPw7geJog93wdUtz+fzaMhm2qtPXZ2tkyF9vwCsq4BfCcI4
YBBKdJkArkbCcaBddpz9UAgChGVF9VMs4KdiG0Zn4xBRSFY/8YhUuN/jOYYWltUa
k2waASd50lbA4jjWDDiSKDRFM73E7D+bDD0BEJII1/sl2js1LKSB5bz4aF5pQz4o
y0K9fDLG+DzIFExkae+8x2m03tJlnKFz3RozrFjrZ2FzGLcJnDm493PLc+XYUVYp
l2WHZftT0PtuprHMsAyPsOHmeh4MbDGqJhwv9XHcvVovB0ePNWkSLVxCyYz+Gyc6
cL/Hh/taLaRHJL+refpXRN/wdAc/jwD47OhOHLllf2bRpGKF8BXXxee7dPMvtDmw
FNCS6kdozPSDguyGkf+A7v3ZbvHLZMw66C9d0O7pTE7Wb4XHvg9L4fdpTfC3mz8O
EB5hBzSZ3Eqk7FnXjEDVlkH/ZFjNH4Wan/LXOUNVAFuWqNyHUthQFhj9CbS62p8N
kiUFktt62Q8WbdRUh8RdxNL+7m+valoxt2XfxCm1FDQvnK1wcxh+64Erdmv38Nni
TH0hn8U5xIUvYZo4aXCOJ4Hzj6FCw4D+FeNkTa8CJ4J/U1HzKsXk9HU25xZJmJ+Z
1/xxpmnlKOsj87og79wdoatiZMI1kV0/Joyl3iUDtFf00ShYw+k/Ro1Tnto+e/3u
jmrkMXLrt5U7yKsBosVuNZx4AdnQrthCabXhXg47ZGogaWZ6L6iqtahFPA+dWGEU
9V6aGYNzIocxOTUpgogW+qhlIMMjM24y1ZOWK2EMvN1s9ppPQQUFBecfKlzMFwTP
WM99rwr/3U+tseCqatY+tuJVrDHKWELCeldnTWZF85JnM1p9ZbpDk826IVGfVwtf
74zPq3P4NdaA0waiDXeKDr0R0O+65Cd5ihu1AHd+/bD+bCT04qV28Cn2AhFLTiLr
IGllxEe1b/az3wizjfLng4WnvaNBth1dcMH7XwXIluKJuaXHIZaDK4B0oWMSX16e
1c67lKMGR78pD3TjevA3q1rIsuDEmEG6Id2Pek1l2O68E3VZoprJeRsCuJI3TS9T
msqid322h/Helho4EMdE1OmtTzKCQaHxOdCNmgBDUgQsi/To8g0hQgU8XEPl9mei
gNAsesF009ivV/IUln1nRFMBtFhNMVjs4794Own1NntXAG49dIYg89iEDM7iaVUh
ud9oE+WpfkO6nXcH9ALPsG/azKaAGbcs7Nbqm6GcJs02kic4DcdFbkrOcvUssiSt
8fahof5cWh+iZ4DkmWKuaglLu1/JogICae411Y92CibCNMHwhX+TH+rc/P15hheJ
4DEMZUianab6sar0Sc5Yp8UYxNrAoY6lOnpnNvqeWpXsUBNT1A/BLi4A6TIe4yQu
NNTT+0jlqXa6S9clVrXh32A0VgberOZ0D/OoYYnRQAp9KaRURDP8vvdUpWTqcbG5
eGNUqtSue6yPLXMhF4kuYzwAFj+nwdtWbbKhgqfG/V3HIAvrdn5dVau6P1kw+rKf
tV83oRncEpaHhGrkDCPrIutlPGaNM1t4GPy87iWRStC17ZHvtR25Ssv5Ovu5vVtH
qB6/7T0a6PdowwrsplQ2kEy8bkge4Bj/A5Il6GVN8WRJPa9yYuK83NUUDOqkeNb5
hvgfsiMURx01cZkatM8fdgP+nOQ/fTKVzjj8vXq8Fw1a9H5NNQ+FF67zwAab5zmT
SQm7okRL/wkjnmpGQ4Zlut5gKpCV6hd8zn1dZVBLeUC4R9F93W+UYt7P7PsIgzI2
7dZdcq12Ew3uDM2O/VBIGKboTrIT4R5129blbPFwYK2Ltfqkftv/U0g0Y8PLq79/
aNozKGdM8kKvdzkFBEe5rTh7MIDFQ/ScuQxp4K1KqaYg+PUMPB7rr/KsLzx2lfWz
BNFg9kHEjt9HXGkwFhojpRZyIvFKy4aG4kmyKXBg/TkKTUCb7J7oegExf8rY2b6m
8KUVSUl0ArLmTgUzmCHTEmQJcnGwmqRgCNQpDp61hPEI2A3jjDGAxxoDBW4DO+cL
YSFYNsNUUgYqlYsJjTuT3AHKtBaB1HqGM9J2GsdkLOjZfaPP7+pW7RJxWq0PFyvY
Dfiz57kzLuuM9XDT+mhzRTtRgEuANUKwqgLy7embUG78PFs/Hq88jtnkY1JFFoiK
re9G+hyFqFPSh6lX7P1pyucksIWAy7AyiwSDxjtIZfNCniUEudtvVuZMpaC9LCsi
XGY0/B63qj3c6uC95q/HI0TLXLfldmfp+ezOWj/Vg8axUIpX4Y/PYiQeW7CYPPXw
bC9x6TYo2YSikoASyu7BUwQPQs6vlh2bFAwf3wifdmM5k6CYBnYX/5bcgyuU0/+u
PafbJx+2CdOcCdXEgvsSdV2ZkgpenwBN721J9SlOXIcSE+2b5S8bO9PMR2dCoU1R
YJxr/mBxMCStqyqd09bO+VCwW3/HCH+jrs6wv7ROVeEsMkKhZw3cAX92HYWRENWX
WJeRUOE3FFM3OA7FIZm1k51aUjOWByDMIjlWkn5anVsh2mAUqXwgRStSJH2K5byQ
w2y93pBddflFpu1IWfbME6Wo3z2eJ4XvGQKUZQrP1MA5iWnHkcZDANkSRSDA++Fs
pboACAPiwhtfNehSde221/1K5yBvQC9iKnkcp2omUsZNCgBi2uRPpDjoRp1e5KPH
3uH9Mfx1lVue1SpE0vldcLFX8cipIq1zEnn/XVzJaQAv1tTra8uNPcKD/up1/mkC
kpKVnX7hvJJ8ZjLCHtVXDYi6KkJyBwQ9ops3ZRtksj3+WdeuumboBcbZGXOzJLIR
OiQXcvorFSGDy6N1T6SLBLYEKjU6dY/9CykZj27p6oCu9pVW8vL1+jd41osZ4UPW
h4wWmTwGIHghYFT2ZyIisYIVGFcMEBKSxIagYz0UeTzlNSnVpmm7Uqi7Yv0K6Jf5
xwRp19eg/GPjgzFwX+u8sj2tGofH/ZtAmSMQRUXhyAAI9jzm3Qcz4bkRaE9dOlUT
rvPzVfh7eDaq+HzF3vaA62OlCAYzek3q2SxjMyCLGKzV5cVmfaK4B7BEw6+03/ia
kpJrAlp8g6Dhj+19Y0CSWAtOHYqzUzUI5jjVjFdrPtS35wfCDiL1X9XdQ/Vgi3q/
5QzCdP0JApAB6e/ctSlFNaMeviuXgIosp/QCvkracad5T+Ob4i7OzbE8fQwdurSu
uuyMilXqKPirOJYorbedyPhTAhi5GZw9rg15hOQnbkk8PjTDNtzloljAbvHuEa9Q
jyDzodOBT2JLTEOTlKRaGD1+5HHvpspY2G9DhUDy94DMsbXrAkmbkVr6bgsGzriu
dtq4ImZRFQfYtUkO/Oor6P/6NWZvrH1LleiL2ZgV1fcDEn6OCcsEu5UHAmsW44Un
zyeexw88m1gi7eIgTVAs9SE03GwyMR6vn+3HYYHBhsmC0ZP5ET+4QUOYrEmZqMg+
kFbPApLlkhqQURdt27TKYgrIyKs/zE3itmMBrxRuqluXN3gK0BMlDl0FVbEeP75U
+l6gdtGBOG2sDisqU+ygj5vNKTEvH2E2mdrkjaD7NhQJ7Z5dPyAMZ2hjdFzPrldk
vs2D3w+i/dACbMHVM29S2pXGa/t2rYjYYHHhL43m563Ob5RKJnLcTOv3C6hMAyiv
gmwplJytE9pQunDhexqKO5X4PIvF6u2PFUWH2GtmPBQPxLrtRj5gtlFVcvm1KYda
eHVY7CjGQY9QVBfp8buQSjvcQ8knUwcnK5WgjATszNP3Byz0vyQ8uIL0C+I3OpCa
Cj4OrujA0fSu6TFT2rqB226mYM9SnpbczR02WSScbT+vaKn8I++lboWefnHAC2WH
/efGc9ahs23nacT0KxBdz33me13pKeM6YpEcE1wTfAxD+kj5cfEfPYcfgghqMrAr
eb2L/7rDKMh3+MAmTqEiBpmKOB2ycfigvHJuyPINcXT1AD6FKoaI6RccBZUwuN++
5SHJhd1jPDVIOEjAttiXi+3wVaEoYj5Ptmbq7g20f0/5POifKUxd5Zh07p02vvbR
Z2+xQwfs4nQrFjYapQo/j8DeBQAgM+OE4NI/rf4FT+aulWthdyIKLSt8pgQW7h75
WOZSVqKmt0yMQP/xJry0kEmdY5pjruDiXO01uT75vpIDJkyv16NTFp//cSfPDHJ5
XiyfmTxBiKILwrQq8SwUQOu61v6Jf0tnJaPov+35IdxjqVyL4/jPPiVTaptUGOEt
q8MUvd2Oe5VBp4GU11T62zTXQl4GJ0lpXAYL3nUdlRGDmCrWN3Ip+MOqtF4EDwaT
AAyTERvqFBEFWq8dBKfsGEAjGBe91935xwEz7yQ9vOLhgLw3TbUIW1zW81x3Vg1A
JmImRptMmSi2s2al3K2Tv3R4R9O8UTOETD2XVXclQ/l0bcZVIXPlwzR0OzBmnJi+
ygaix/hTVZJtTB1NUjNX91F0LzRYN0oRtkUTwIhiJ2uZ311F9pXucCenE330oa4m
slvM02co8gfMk3EhVHcwKHZD4DUf219imIvHwv7emhdSkkzqs/WbKrS7pGPdt5g1
eaLyb8wkUb+SpO+WU5wUchx63ThaAX+O0njlaJuFDf9jTSiv8A0POI5M0t0oW3yJ
omhleZPsw16Ro1KhbtBWZlS5PGJTSDjwYnTBltGo7JkgNmdmN9wF6iva9h+CsvOw
DloAQ4hhBwhZvVb0HvjFa+lRDg4htukxyuEMHtjZBeMIiy56/+cc31ua/cPa+7Zr
HhikKuY6tzDq3klgswIF64T+v14dbQ11JFdAxzPN9K5jc0p2zKBgTX0oNCeoMRmJ
ypTcBgxDyv0rzjLaQTx8oq9jhXMq/n/0Vniv7+bwWOLBS7dKIpn9wk75PkrP7Yth
cHh72LI9CpYQD6ORMJXH9j9GdnPwt9abqDvvd8Kxo3DHRBt/2bxoVl9Ns89uMv8H
LnYg4jdRmfSXQiH7Rs0ykRppJ+lNrQgrPorW5p4Rn1lwBkQzJnqm/LVwRJdQGcJu
qtpy3iSI7qax66qsgcSvU7zFRGvKnvlh17tihU+Hx3GRru3ZYeKUry0dhvPVdPBN
HZfzuVJcaWv1pNV57UyMSPW0uCGOJGhp6xr8emfjfRK1k6/R44jBxZG1Yks5hmGJ
oHEH0pbS8KCxUP279gUPiVr8Ou4O0lIgkkl7OVxRT3q1V7mWCdJVWuGXLVRRDmdi
gZQHuDpNvmlXTcATrSDEk4NMVmR9ABsnyTavAtg7JeyHyj5cfmGWdsodi0Cm1Ut/
tKeaHMwsdYH7uII1cSR3vgC3OSZGYcl2Cr3HQE8gH3mcNLwTA2tVtsh2Fg+dyL+g
KdnkliWpWnmhJyRkZH87Kq6eCBmwWHBSzH84j6Wo9Fde9abyabo1qps0qSdyk8dG
hLtGO2g0RqUnMo4KzcpPs9uP/kQpxREEYBvaO1CU5n7LI3LLQuU2/WkVqwE0BLuM
c7/wg8p54junMb4vydaZR5B7xVhgF/yBNZKlP4DdcHL4i8DSNU2noAEbOyQTAi9e
D9vVF2uVY0ZrzmPPj6gj0UTBgIjHJ9RxFMqT5k0BaAsE5mcdmtB6vhmAaKi6EFOr
dTW1nsKaQz3dPjXUb9huR4EZ7qTtkVUAPZc6S8ejunJOBLPK8Tt8eSatSrUSO8LI
ivaqrgTXtex1dnKRizUaxk1i425tCXlvF0AnUBSkaE/VAihjzvmqADel+tjdtUsl
F0rL1l9bwK3SGcWS/XSSHcu4V9bt2BKywpHpjfWS2ITUPhjL45ZBfI+6htjf5j1u
2gVx1QtBdN3USkb1bQPI7yRg1cL1e47uareMw4qmzQYWcQUTUhcGmeyie0iB3ftm
eokZ8ViD6dpmo37UAoSXLgjTEHsrOHcUF5rs62VTasaICkEe0MnjDKx3yXbLe82V
l9iusL4rMsnyxK5pF350XbfIxEJLVll4A+wJLxeUNA64zuOaZv1yJBlXH7XsTf47
OBRCe+1HPSNLFIfex3Mp2kCrR6kgLKpECGRWpaR9xCL3wgwt2lYy+KqeNB5K2Q9N
ESDpaVlvEl9PunFWRW6+W/ogopbgWsJ1XyQxZ1vZY2AyIityloiHbw38cCxl+DdA
9rdZIwB7bj7SPU7x/qOjX03cGa40XZINl91swXXmjTVa+nzNmq6Fl6sBF8b0hGrP
Ze3EzMCGgyPE7f9ZHU0cYfLmtwxlVQST99Vyy6c78RkdG0kHH19uFTULPItZn0+b
M9sD28BGBOlfOoBBHpQk4B9f4ebX8tC/YQ6MMDPnNF/b31CwtJTtf4lk2fF93CYs
uaFDcQBG02hEgzV14SpKaMd3UrQuVRVyPD0q3e3fBKBAVDfvbYWlY4HxF6Z8SrF/
WxrhnCmtjHHxVe/F2zPuXpOpFnn4fFZGDCiXP3kWKFAVzu0qdw+6WZfySgqSxCF/
8kk4J4aZKvwyovjnUW4RoidaVbJTK2ZMRuV8r6Omrn5JM6DIHZmXVPBFqQbOE7XA
NAOXuHOVC2EqmYbC1C2EfhXZw9CO23G+AdCPYg5YwPssjCqQ9l/xlX2zc4FEaeLA
LknyHNaaoOWVRoA8PoEcdv3SmupP8xIdINmgzwK/pgmMRSpDvNV8HwIB66XkGu/a
my+V1x3YDqcX8xmAbM7aMjM4A1rSeR1ZL2EO5zYxHmXJwe1oKW9nP4wgVZpPKaB0
FZF1Xhc53dVsdGH2BAOyBKwHZGpWm+6GrtTfGjj9OK5BC8dRqvxj+KUhoqRLa1UT
QMGqHUrkKB5931YnHzoO2/9tqNQz+ds1a3Q42wJ4Gw67XMdH0jf1W7wsRTVz1QvR
z4QLElMKx+xfl/gRHwk1o7Vd3MxCHOOuLbFuyankYnXOV29Anqv5xaJukZuBbaZL
ym1SR7TaBPzwcxOMw+ftRmWVYtTllzOIzl3yA2YSNgdOYgcIF2i60Za7EOlNWBmo
FoTfhNvlFaELjFgVrayFXMLh+8zlTuZEXhT71KhZ++SV5/4xXytx0AOu9obN28ct
2XCz8X39YmP/z5qVUj224K+SjUlqqW2B6Tg/UL81F2NLS7S0xmw/YA+pnrhM9uU3
aaKYQmNgRXegY7UEhHaRQT4BIfoQBw5Tr2awMaplcrndXsipXZrxJ9GuUxaU5M+C
ZG3oSCWteNN5owNdp+CIHf1k+hmsLDEwo1Mc7TsB93p0nRqHk36EDxXfjayfksfg
5VBJXyPGca0niuEfGIq3aQxKsxPNNxipcAeSvHOP6eT1uwPUKsSsN+bGROI1ie0F
TcWWmqSvebHN+qdBlcq1Eb9YGdB49G4ZO3ZIsDjV3a8e6wdZn1/kVASVaTf7nbke
875OktPSnbkg3qz4oWg0av7MbHnGrsaVdyi9EH41E2RSP4Cy80xJBi7C9LHGmpj7
6MX48StSx5vGRWrU5zxMtPGb8Yg6i7ucj3RHRtRZC0Yl0thl1gfIsC6DtfmeWpmj
CCS5Uy5GaYu9FQbBK83rCxczkFOO+cKVUu7lhSrCzyMyHXjiOm3OHAtST8m3W2Em
bFOT/hNHabeQumctqsDz0YWxr0rtgj6ot2sQ0EEo8sfxXoXzingcEA0WmX0spIVH
QkC/hxSd4SGsRs/IPOfBcPl8fpnkct5/NCSLGehcjCk50tmTVChRnjMV0bg6wzi5
OaNNq52QbitEUAYBa4QkLde7eYfljV88bX50+e3t3JowuxIJLfF4qv1mWIsk5bAl
LgabTx5ZSBNQ0z/YoyhjbBmMP+w2yYajLlEANEWo5YPojFAWYxjDztfAPH+r7WQp
gnAGuNbYy5U6hKOl0fEXfHYXqon79LdyQ/Tei23K70qQSq3MXIbVH2TxNsFERvQP
E4D9mWMJBkcIe5H6PdARbVuqzA2u+gGuZ/Wimu6infxIEVUlg8ztM/fNQuQ4Y3IJ
AmXXcAbhdC7ns7Zm2RYuuF2FPus+xhgw56xFhqzs42eLZYTvjncgqqT5Cc21WZ4P
lFAZFYpeAiiYM0ysUH7EDBe4Tkb0E5HbHYjTtRah+D7M2aGDW42WVwwnS7XIFmn+
vpraPs21iGEeJ1R3uZvyuEjgHVYKMEsNKwLkSynFuRRutOGARMxecaUtmZ9L2iZd
49znkxqmatlHs5xfghYN3RjNYGFghzC1W3IBTXTfyT/S57OPAf1zYAh1rR/tGcps
LVadTzp84bEssDADCvOYD72kx150tnEGXqVfGKYC0hECHNl57eccc+BVU42ozLG2
mRTD7xRCCSav7zh4zrihzaXJNB7uRpAYQVjX6+DJEAK0VlPUPlChBEt5KOT/SMwC
zCjL7fPhRsdl/o1A8UKr2jhh5riy/bcQ8shFOyJrF3Oxl6on2qhCJsyh0kgoxPoy
TX6/1gcB2UDIPphfeRuxhlMeRKqvgurdU0OJTC41uNqRgjh1O6TGVn+SUZEQJB8A
VpV39tCos+J6KKsdfZr1TaTim0sGpFvqg0tQJiFIWmG5H3S3LaHHlS6fYE1v9daP
o7VPeQWYgZfdQYCRPvfoGPEj7UfxWtQj+qdFoUz568nlbCjJqgIF6puggRo5Vq9L
xDE+axDQP1RqOrmBvYKpch9e9PqhNJfvMA67rC1QzGlBAulAlgjxgxvPxMM29hYK
JFJlRhJbaBCiZZiRXGRVyxPUrlZoI8LADr37AW/9HV2YDLbUWucF6f/4lS8++qDp
yW52ZNMf89Buz+QZwsbSyZABM7lVKj18LpsNwtQa79zhQCkxITylwBIeGNZKHPd0
etCQIwpKdDd7Q8tNhAfAM6uDhChmAaJs0n1qVTjHhVHeE/2ny3FqRjsAYkPsttaQ
E0skSk29cgpDnYsG8lAMhbHL+zqdYYVHfMiz28X4KZ03EjahAsOWn7N1DeyPFV+9
CwyY081wr2vIZM0dGgekTTl/tpHvVNxgu0LJFVUoTF4+lXb4W5H+kLAi4jdhuFjK
/CVrIGoAcJVUj6gdJhRRgLYH1L75R+B9krNTloiZNKKxt65DQlGznwyHrFUzljF4
sIW5eIQv8t/l+fZSZO1H6UaVI84ua1S80QXuxS3jvWbkvaibeGvudR12vKY3lf9I
xpjTmwhNPdxRMfbdfeG9lUlMJx7dzJx0wmX0nuLXoQi3nv2nfcLYULKP/aDxW2Px
7TV6p7gcmAbwKR4nNwEffIh+nNwTCuS063d2FTvzv/wgGVcO0/HA1eJH2HW4WH46
R8FpqUM7ZxUJqni5yxSl9WOH4xjqDfF+fx0ErSAAlZwhrSmrAo/ssOxD8Ea5QbsO
6vxqww8ofdZPWKaJIn69UgK0odmJEo2CYhdMELYwq0C8rYrzej+DsMfNmifiMMjh
DIY3DumyKnM4Bel82ucA8+7xjWHUEu/1MEBRmkEC1A7+mPGoJqjcniiOHy3KMKBq
5TeTkeTAyZTg0w0zrtuELMVddH3OnwWcVVtApa+KpogopJEhXyqqYsSyzEuosuV9
5ab16tc/0ATItHTV2ltVVLbMBty3Tt1iDDSREyZSNt+kDQOFvkcYedU7LZftNwzC
tJp426LLMax4AbXXRnDmQuN6EcxVg38eOtGxW0lya3PT2Y4FDQqqhoFdwIZMDRlv
SPI6pW8G+FcTofm69Y6V2k8sBIKkE12wQxItGrd8/BtRuebsBCZW7Jyo7/g3mczK
m78yHb9xjbcjcLhoCxKsf2dxgarnJ36oadk28s5XwVySgudsp1Pnmgoj4nbsocsf
8HNP4sZR08vrkf4xqjkLmNeo5ZcWOOaGELpmbgpY+9Q3UUQzCbFK8ZraD8l+Li1P
UUg2ELi7mmcP8C7gV08oDw2/+smkTCgxlWXo9RgoxFIsFopF+r8SfLgX7KCaLS2B
1WZ/LjUqfi4iG0WeqG8Zd0s4yridFy9fWX8Uuoc8dNUSBNsm8qkHQgiqmkf7eP93
N4F72UugoRzzigF7RQM/rzlHlRkRjGrJw6YXbLaJ7GG3k2jJdGMjjD9Qm2qBmrIu
ZNcpbJhf9ubuoOpeTTP1/pdtaakQNUIFmV6b326/nAAILJd4bt7kzzMBgr/kLDl/
NGNlYp/q+lJmUXG/CY6+Y0QxarcOhPMNRn0Y2KrCIKbMXJPr7vbCtFQ6i8h7+1gb
Gga5PelsYIfAcA0KXBzo/4ZYhQwiCLGY6t3Tnt9AncPYxo2HdJDMFJxbCCgEi4px
0IxOUYH3ACPLdMtfHc03AGq9ZqCdpvFV+NuEGj2Aq2zCT29RpsPFv4hBKt5DfCnE
eGlZJAm2TNZN+FHyduSWpzZOJTB5bh8L6VehFgfQVaIArKSjwie6gFTkRLwfVXP6
cglhELe256Sf1SkDsr/br+QkFn295jLUsywt1w3d6XybACYblkyALl1czk98D189
PKyZug/hajsml2ASS2ZT4f1VxQuSmypMOhp3vwUWjqQc2pCmbIda98M/H3PRQ77k
+oIIBmYDRVGL52s9fqxNzkSVIdZqcx/PpvODb1MmoAUgp+eEwLGhLj/e9kVYZF5t
od0eCg+Bro31M2y2lM53uKRblEkJ9uzsnbm4ahzBzBUcIhWXHWvzGqKOUnJTqSY/
C2RnGoM8uMdFQAZwXiUl0UitPnpPfyrwSyi9g+hHTpov18UqCRpYD5mTi48RJMVM
QofK1ROs2nB8lUyQoPBrn2Zq93+k0uDEwWQfN4qZdqoBeS8RTp2LBi3NOHA4P+Yj
5ZC0iJcR/xIqt5D/tlipLseX+Egqw6v98w3h0hd6CELs1+M2QOxc/HvVYr48ym+v
kWHUYjDxcdUkA9GQkknzApDzMdP7Qbkw6T6AZjKO36aiVM2hVKCelsIEx5tkYJG9
s7OVtPN268tuErb7etr+E+NM2ygHyyn3I1UEnvvjTnlsJpAyAp1jXfTlFbGTJYbR
44Npcl5eYe9haw1HJyD7u+/0atc2kFYwS2Hxdn9hy/rIO0vTztoMOrG8kEu3H1nd
Idz57nBKzZIoHqLx9IDJeZEXXcFXjB+nzzwUBMlkE/PXTb/up7Y4LpcTLA5Qc5vw
mQOvskImBB7E7UBPWQySvgtlhf//TRPF8cxdhj9R/49ko+xKoYYiUI8J3rj+G23F
8pcUAaHmUqVeSzbGaXuahvvLNYCcuEiQfqb4krWy22ILirZXqwiIxNSy8fxj3XEY
Sjz8bzwkOoIQVJv/MrgM1aBrmJL50VhF1Pwx1gg/rJNDuC0w5IPYFERRCcxPIL3h
G6NtsRAEyTqLsPlX61VekQu+wa87SxCQ51XRGeykvfAyqWKxEN1314z+gHL8AdBz
WKHdXQCSJ8CvzlyJD72kZGuG7cdEJ6Xgn4KTjMjIZubFO+NFka8LsLTd58CAnICo
0uaNQhwrjq9lsK1VJrNhPNtoqKojxbSMpuOCxDWuAwBk6syfV1uRfrwmmvIv3q4l
ZfOEWCPYFsKIfeh8t8icEaJ+n9vmrgoPU2xw8LDkzR5R8Cl7Gn67QRRYGefkLzvK
bQOu3qfqUIguvUaJudvz+JWZJcNVNO1a8IX/OPeeDKmBAHcw1knL5cfIC7GlrdO5
w/SzAnHSDf7JUe+qeXnXuUSLMgG1LxSVRKkRyBN/vjBBss8j3mHpNZPWGAjKxIyM
qVtVLkun77UwRdOEn44MlSMP67qbLHjsXxQl5pV4cZuh0X/l2JzMj99poxX8dtsw
8aaOeEwRRFIBhKEJt2NGUBwlCCpemlkuX1HZFxp5LHbER3Uk/kSaUzJ1b1LWgmcO
u+jVjuw/vMDXymfvMP2k9DRye70b99tTowDntfOv8vaYvRjzcksk+T6/lh4YFivE
fLVdme/NYoqo+ZEPisBkfh4g9HhjH47nSbMyS/2ncVQ8XLW6U5HM+woh6/oU9qlw
XOQME7uMgcz+GdccnomiYYBWdfH3jj+MukNbndy5TOLf1p2wXMHpKG8No2oqlGi5
xRSiziXsn1rivciopNjOYGXIJun6F5PfiqbO3k+HVJ/Xy1BWu4HVOMK1aS6sjQ11
nccieluemxPORZOnnLWh2fyfGzD6O5zicc8DnMRJCmxKUk0sGIgnievAXOoXRv3W
WZDpbvMN+mJDkdy2UfoIyaWgnPXz9E/XJzomNOLU3yM4Ww32e0D+GsCZGUvAbSor
D6/eytCKMti0ExiXKQAQ12uzcUC0sCY1FHkNC+YtW5PBntqV4zMZdefG5Udzkh7l
1rW3P2gGl9/QiDJQaqVrUjumtLCgR1lUS5WBpRTggBgZXmqPYFpHXPoue29G9eKX
g8AEVwzsV5gb3jz+8ahSifGFr1ElV2/Xcka1KIvv82WJQdrigpT8vGR0Nzxnem0B
6T+fjhzuQgDcMJVbNVJZEtdxi8jW1U/LxpvBBvLmhG6FGe0DTzSRJrkGD/hZaMHJ
7rfjgJ3AnaiZorvJt12jP8U/ftsaG6ulmL8uxVspa229jqXQ1EYeRmix7dlJxFvO
VdwOgBTcVyQmzj13cqSH5kcxANjVqV1V9X3lsTQt/842tsRSYHUxpcxYcaMaDrZo
//CqJgmjXzJGtI5rxuprr+JXsmKLc2vrtNvLydtVS2FjGpO+Z1UbLiedY9Q/aDM6
HfvaUvHbu+d7qJsMw69ttvEtzeueNcxwh48psAtHJ09h97NveFIsG8mVZEnUapEj
iENINXPSxmzBBZHPU4cdv1SdS+xgXTxF8Ta+MDneF2xOVgBzKGFpRIihW+xhuc/b
3Wc7e64vtw7vJKCkYoF8ABMoxJ3DFOQ/s1zMDXGCg/dyA78av7Wfw1u/S2gFJhhX
jr33Iwnowq/PeKR1uQTEKzVCq5usvhqVPMwtYeZPWUjlxaXPjNpykbjGSrNxB45n
21CHVH5WkZBiu6048utkvxhawjlWaocjlDukWazzQn3GJhZ1C8F0CQXRyysBWUR/
gS8b3q8bIFJH252BUIOl2GXQyv61uBy9eUBwZHLuYUsEdU5ZyRQzW4eRLIPHGoz8
PHK2zz1gq0h/ZH0QbSkdCEtXL/XskVT6S6N5B9DBZG0kPzw0251wCj8sPUXVwoyj
5lMb25cEBX4otx5ZSYu5rx0lKJwHU852FSSP4SAThPLy34RuRfy4G7TTMZYkByBE
0nGFQdaZAHFOFOedtXfSgkryhv/1AMWixM+dYOl6NiNWVLwfyMhR58tKWRtH0nXv
iZmG35WzDY5Mftg2dWRXmkqXNOavIn/MsDr8vr4UZ5cDotL7WHvQzFuzLg1AwTls
wkjoJBdNnLT0sqV1vIXOxaAx6cJYuZQ2RyGWwRzEnT9F305TLf+hPnWEXZ1wFgaW
t3laWIPMJ43EnfZs+qgxcMAYp5XK380MWx30Z4JZb547AvXGZ3LTUbQ8iGNyuNVP
j+MnYV/Q/ypeiBIsuEyhm9Y/G5W2uCk4fA66vzARCg6euJLtA5438JZc6vx2uu4l
RAkRwXQKw1Rgj/o4QkrLHbxF56s5Nsn8Q8zaDKHn96Ym9E/DkX1xNNDLakuTUTXK
6CsSfwLgDoxkh+MDQjbEH8XCoU6/onGKxV6Zy/MjEaDc/ON/94Vcm9UzPwURYB2/
PJfSGJTW8HGcEHvKRfIsBJVuP0iNzR6X8hmruU80XPR9oMsZ/uNP/yOscKLUrUNk
MChfyE2ST3bSNFlnw5gdO2GH7Q2w35xvF65myR5sI5WHOMSTcf/Aa++yO6PXzfvb
QKt52FPV69XW+F9TvPFZgfAOG7BaadZ5ld8fyi6R1Fn1Hnv18I1A3XNU1NiLzZ1l
+YJXU9YXDZGjpTrIg5t1KvzvRmtoJUdjhQ3UAuNN9EGZV1+qshQAmcat5X1i1VCm
MhwSNfrwN4iiQEiL8RUTMNO7xpAl2djV4fdtw9FDUOYb6d2lB3fJWjWuSyyawJ/L
R+KtiITEJ566MGxJZR4duPecwJVw7Sjnsbz1IeahX1teo9TmMLug+jYobOXlbf7F
/Wvad4QGj3IicWQ7CuHR7CugtdmZcwP4cSo5eSixmTguAb4lx4nvc4Seuh8wC9hx
rkMRaHrZWUUyT9oI8E4qCDHkkAc83Bk8tnPmLauhq7n4rnYlDQSciwarLtfEwRC4
+xBB70pOAjJM0VaI8DvsNFWo5yTbsPlZah7LpSpOQ+h+xEdJtEMHlZyIcGX0neBs
+Fj9OYTXOVdro+teGfLyPrSZMeUnIdxAsiXbw9GJMevFLppnk63fM/wuC98lKK33
AZpXv5DtlRYRGSiTp0YFgqh5Hb48PKJfFz+1lS+YqnoSmz+bjsEKnGeKDhNeta84
No0awUIV98RZRwFRy4qJrUW91MeBDIjdLzQs8SItWNr3Idk+5xsLm6956XQzGd3m
cEZJ7QL1fTXt1NIeaZw4IyGMnHbQ2ljZ+NF3Ik8pCx75aqoFODTVPccRltkw3sbt
P1jaRzP09+xVZn4LPjMbqCyVA7XBgea1ijQRCwL/KzBPDX0XFK6VVY9qklTWfTHP
otCCJWLErmzww5oqUUIEMzdqJngr6ENPgBJLFGhboufMkE2VZddFM7WtPl/QbdoC
VmnJNdrAbxN2ThUlDx2DoddClejovMSXj5HusbwF2Uh1Gmt/27jp1qAquyVs21vP
EcmA8bah5yAzqMBzSixvzC09Ypf4c/VmaNaYJbyb/S981sJ7pHomqIyURHK9jRCv
oyJgiIqEEA5toSug2ccYgufYgLwN13fPwetXoTwZi4Ea08s1r8ebFO24aW7ykAkh
kKh0BEqm3wwXaPW8he5ffBK+EVZbF78h9HrHdujdPQEe4YsuJVx/V1xoIGZJrP3c
7z3OzXDYd7LoHPb/pJpJ1QuqtsSjjWsvCwMn1xh9VWoHIm+2dffflSdPERMf2uw+
pXB87Mee/6/kFuY3mBvcAvLBLx+If0ggex6MRv3WYcx5Zz3IWAVTw3aS3B42uvcu
ec7NL17J16FroeQ0hn4QYjS2Ov/CmbJu7f2P9UN7f1o4q+f1WLkEoSb++fDBLVRD
zQRQFW/VO4s8vmThV/Fn9TWtrigVfiWK/MNr5qZey8XZ7JWH8v5zpwDa9mIasouv
XfDq/cWcdW7MsWsnTkQFLNKLJHoW8lgWjTCMrNjBBMutcayn7OIHDwb5JocCkKyz
pwRSPWs0VcyNS/MP0sYnqvXk4CSp/NiwxbqP0+sWkJu3yl4QgXCmhWnNyl8uV0MV
yqf1rn7RCOSR2KXVgnlX8nlEdX/9Kv8b4oZCgX3S06pEK7g/e+beA/N8q2qo5Hds
LmYJ8HU+RvpHMhZCoCCOiPpoN/bc7GfrhL9WH2CrdFevI9PJdMNO8tDducmZHd5W
Lfl5tPxpjtBFCZ2tTCBeetv3NViABNXo16YzRExCGktDoCn9nkXC+j2Vddhkfl9J
cPtjsL7X8T/RhVeWn43HxbRhgS5uiWQlmfABxqx2IsCgs5sbFqFMWvCdPXsVz6X0
zVTZ9xORKN0FPebiB6fZ9AxNdp2s+GxR/3X7Xyy/DN8/BEKAW/A7UKduCsuwK/TF
fmBvORKqqKNOf7oK0sodNCKGtxId8aSke7upSmeCbPsYxABniucdoJzOVMa9fxIZ
JgBrjmruiZvKen8B1bEytQ2nVOK3uQGVKCRI2F0Q6xB6vj9r3c12CKawJCnZS1F0
NJYX28tEz7926H4ndt0h/AWapYNRv24nvq3tlqzG6M/2Iy8UOE6WDGdbi4wtBly3
X8c2SLocxs1J8dEw+Rjbd7S7LQCmFAkkgl1n41TNQfz6MhyIYnIoeWjMz7Dxkm3j
WnjPzbL2ib8vGnnDWHj5m0V68y1MBB9KZr1dNyj/+77iS+8mbRQ1okXTGTmNT0hy
12ASOVQvoTNWyYQpbKICHjEy4hDIUeY7bg9HFaB4gJeqEXBSBODN7bSKa7QXU8o8
XDDQ6VShv9A9gzlAU7x9usk5fdFdq20qLH8gx2/nxH4OT4K1ZP3jEOT86jYSvcwo
44+84/GH7oA9ROWWx0pQPQbMYIozbg6LAOjpDkiIhXI7s8QzWc6VgopZpnqyL+pp
X7o0Sagc2i45ehm1edoCZ5g3B07gZguZG2Nyp2JhYQfBZePmHhsoibKeTBoImNBx
IM1gy5ZOpM0vtjw9KpqOKM+GeibzQwkWTnoVtQJDZUX54+aKY6hFaiBokH8CZ2Ik
oS5vAIgesfHan4gZ3WsK+nI2kRrHj1itrWtX4wDjpog2QuMwUCwI625iC8zRmalR
k7aTr2Xvwj8bcwYhhKGKtfHuivT73kzqYhhYdzUvdLY9bmzxo8h7kX5bM9JIDRMa
61GO25//iSGUYqRTkcIcpP+Fhpe3n8En+qInwT7jjCayazE+msPrOGcfbOy5Zicl
EIOx3xa9bowAGLEpUMF4qPZgcH5Y9O3n/MFJ28BrEa4qOuHJPJWzT0gh5bQVh+kZ
wOFIlrrCRvgrG4UpHmBfgwhIDOpB4ybY6w92KPCGRckA1qDiGP4qT4Qoh75KtYGZ
Y5G7LaIksLYz3ViHDm14iJW7UrlsU4OYD+JmXRtbAowOPXEm5vN5E2reUJQcINSA
mpbGOmMJRVPBRlrLsAj/puBpB+vM9av+yq3zpFxSCWUMT2gQiC2mGJLCLshA+vwD
kNvZTtYp1HKjYfX9RhC0pogOtL1NvSQyaJvtwSujdNicpVA/VZQdGgcktBkAK+3K
e5B9rjVvPXEQCS6r8LIsx8tvjQFjKAu1QWJbF9BoUq3jr6gt2OjXBDYlGWFNdkw8
URGKHzViGPugaBRp3vWhJLr11bKIGK7t4OHszgDwLkYS1TAnGkIgi/l1gDc1tm4m
g10+TFvdD7GWKQxUgeqU4vZVGeK5qxwkCuUi5GYqIKkcA3kt6Q3E4l/ganX7TdCA
vcV/3o6KgCYkBOkX+MopBqpGNLrKUVVC0MBea09GDkluxCPdfq/rX5cRgCYSoH3R
AIN98wLiIw1DW2wzigBEXJTBoZc009CPQX+YRE5VPLFLcPygbgPaFlXGiMkebkHq
cLi8tH7OXYp0vcxuyp0Bykr6vTC7+5buUV8CPjm438q2x6wNHhFsmb0+IZUF6nvO
lDF4xwlZbUz0gsAcGxhaCO0QgZOsYp1ukCqFQcElvu4nsHb0cvn+kXSatTKzK4D9
Fp8/NzbUjuMRLb6F1HztJ9/mCkcbsHKM0gIxXnQVixyarpEzI46joPq29ZCrPSl6
DX8+h3RNTqsZuHCrzVJyqCjofXc6o6eLICrH+pARtXVVlqCmwNaAMPgkOd2SD7g0
1PpjIpdMZ1o1LJYVsxGumWaAbdZcR58cps/NpQmqpKqkhk+aPXB0CEC0MtRWc+Rs
PAPNg/DY7dpcVsU17jBsZqT1Hi3+Gi6TtYnVO9r+fBuq1iiaaxYQWlnARI55Xggs
EffY/9WSdHU5u+9R+4fFcQb1Pj7N92ct3GAA7p4HsGG1fUoC3ravkd5QqfGPZjPW
cC9trQ/f7yGZhrdOnDhT5NOlt1uX9VRUIQp8TvJxemBra8qXizmVkEdK4sA7Gd+x
g6soMiJun7PVsehyhJ6QIlWqaVup9lYJfrsFQVrlLHUrGHge2UJJJ1SqGS2Yd2AS
OlBFL3yWaK8rSbFlVt1xF3xUdz7GMjqK8ix0GKMrOt42CgQ867AU0C0H8a/VVnhy
dk3sMnXF9FlFG4ExKK8ptMkc6cxgB19bZ1DpR8mcHhcxoCNB65HwfWJQfg1TEPDr
VSZIdvTG6CJxDgdHn0p9yM6CaUUg9sMYrJydEiXM5+O72TGF7L8wEPCWkGlgPm9I
Cq35csGRWr20k78V4OrU++lPS5XSzjAjD99LDxWABcghHXzAGCcK80BD9fCROYMD
IFUJWLTjqQHsWmqLWh3o91ENRGELma0227xKxur6vv96+wgT9o6uqhFQk/yGLi+y
Eu0gn9wrVOlyVh4CW+2Ss4pgKYH60znfR9GnHQ73zGREem115keZ3F5vt+vD+cUM
qSteSiKQQbeGz2XEHMxw12ga53kaXfzBsw9OUr4q5QbFzp/Zk2e4LH7wKKjjMCIL
dgciG88Kqj4t2YtcGWgVt2SyYQljXaWxjd9yD/HTFbTQ7yb7vJrAFs6ahrbBvMRK
fZ1SG+U7EP4oL89fVmlW7+IoB7tLmfXUGnXfNAMMAguGMa9xZbX48JG+qolTUhmf
btXT3O++CwHapbbUBCF6TJyOvBe3XRBMC1LXNjVmStEo8pMt85W27GaAvV8iyJF/
NdZG0RhGh5l322HJJgV3eFMIqHs4oabELD4YpAzEY3avuCC3A/OlwZc0pSTCBU8q
gJVS5A7JMjFdVEYpvVIp7lMum4UidC1/FRPiig+sRS+lcYb5ILz9f0thf/gjpdYe
Lc08935/WVhmaeQluu4u883E6cYJPRu3KJHZqmYo/j/3DNqKdGxO9bVQskAsicNU
zTRTV6X1Y0UkuC5mrdOAfN+i0dRuO4xFzxmPtyiEo8N7x8220108XL2dmxn8ycg2
wOhNOD3xcfY63xZm4K1KXgBw4bx5N/42+YJI7XMlhtoVuaWQU7Kl5s87XfshrDVk
ZyBlH4yvs7VlzeIxYyfEqndrOLkDdZtCFL5bAne1gybgrjweS5tUs6FpoPBCcXng
GdLx+1coKZIJrLF9u+livi5acIOi/XygqOMQ6+wKm3uYPRZvJ5RAdrCCRHtDPdp6
h+/djSf4iJGwueZUxHDob2GkZRTYL8mtNMIOGDbLPa+wbkBXofltPz/2dAo/LDLO
MMtheIYzw6wtSslrzzwNxIad4siI9dXoOeQeBl/P85eH0OfA/H6KMz1bEpMCf8wQ
NcgPjx0OlsmxGMBcMcx8CaVclfq7AP5Y1ePCkmIMr8p42dm1QS0v/okX4RlCnirQ
hE2XcKaOWfsszO1YvYth+YMXWZXPCkHKRCOn1YUMfQusGsuKIlhN78tOaoixh+lg
LjsQPu8cEpzzOe0r5rlxBrzGftXc1PGq/memf+yXGQpQAqF9PuP9WPBjPMYL9diy
UgI2Mdx0lRANLVRYWojFCsVrGqQWcWveN/ICX+iaUUoIHEgCxEdeGHyxqusnRIPs
mOHvbzcJlqnXU3dDuYLulBgnAecS+rbFutP7/fRGastJA1ELBTSDxqyotSx8xqgD
TaolRbTsvvGosBFZs38HiZpLy3Hr2SWv585nU1dej4M6bwWiTQWko5mA24OV4QNH
y0DpC0PD6rBBJgTo+y+RQCrAkiv1Eem2zP0pT7CQnGVaO1Dq0HEyhR3zROa8c0w5
dQ88CMJEmB5Aq9qidojW7Eqci6He4ptOw8o05Qbhhk0cDcRYl4N1BATDCKmmunFR
iyDtgX8CLl4cjMaigkqNSwIkGS7Wb0FIhiDCvxUA1AIUk31GLFAUuDVxiKL753Zc
RaM3OamQaBBs79CrKac3bdNJJOCEpaaNf2LrwbNUuRrmgMXGPzLRh9p2+HLpp5ma
3tOTxGb7c83wIHeIx3yKiAOKoKKS1/ORX0PNuN9smlCY2kW3WEytXARW+czrUU0J
WvGb3DzBWtZr+lmw0GUWZLM3lbCpLlGuyMLlfJkgLJayxrsgvZTBQ14BbE+r1xN6
pPvSyMI7mZEOuY8GfqiRlRdYiCKXmE8CiOxhUL1xSwOxz1sp8gJJEsl+n+ubgyoY
bLaMpbaiPPB+VXpmRb6jHv8eAgpzPuCdG9+d4TmzvQJQs6NydbzhrmEKQQ9W0NZt
O4Myv9qkBzi2pRjA6AleIJ5fm2iHAYLG93l7hXAU6ODuGqVyuKeQ+XrZPSl8/+cu
XY/l9EvoijfRrcgiZrw583Bmx7AEgOdZulgZzwAs922NBoe5iOIp1TP8OqMNfm6r
l9IOB4VPqVaBOrnfcuwqSH+gmMQNLoTIVx37+wT/e3TrfucwVX6mhFdt8nXUrziP
QGKOX0B3hpjtvdTX/Dwj59cMo5iRk4BcXsYpTnv0c3BB5ZiryU8/g3XxkCx6DLuV
qBY7Ug3yQteHCdYbGDytxjtS/QkIki2b7ETIS3sbvvMKN91ICFLNd15ibFH02AUL
vWTCZvefnVR4IVz77JX5JzC0QBkQQD1TOdcYiRgEgRoPRVtgzRcWplyh5fBHmvdB
wg1uxrFB0oJWTeHUzPPYOuKpGUs90dcFCRG4c9Q687vNgpNIk5w3QgDoi3B7HWrZ
Rsi5f23/oyeYjQ5HCV2khavgtf/DwoANIcHBTG4tslyRIL4f2eY1XIFgkSwq9tT5
w73ZsIBOxIwpEIpTDjBYP31+CGpy9wIBE3PcDsbf0OObhAU6D6M3y7B3wAVg6Leo
uLRRTP8ltYQvEgxFJ4+0+d5P1IjQmStMQpnYULOsIUh/grDe1/TCPeYTTRvTduvZ
/i7zpfUKFJyGHuQWh6tIBilniwyobbh9/XB4pc09uLvwEVIbV2VgpYXLJenYqU1K
/VoYxN+4Kif1nPQ3ZkK9OQhyIq4Cs108bve4W67X7YIQv3zC5rGQ7YtN6rxajt8z
5OfoyopuYXEYF1vOBBUq/prZWCVESlQ/aYrbuRsT9aKiaPZz1QAB4GLDCbwivX8M
mnmOf3hzveQwjlWxJRMA/9xkhFQcCGDbvJXtv8itskkwmCVH9kGP7qu977S1sFSW
5kR3JBLVgwGSwLmZQaoRtPXGVE6wO8GqysXSHzqtZvHI8hyUuXHHnqqJC60lDbF/
BWFe9zMto2txfR2ZQcLOwzrNmIZpv3ui1/p5RMuAeAfvFs/aDVsc3SC3k4Q/7ZaM
qL2lxt5WjXxiXVYeoQJKkU7ZS5b93GpDIDUCrrbdbdu0siMJIbzt9o7mDtlI4VR6
2LvaKcnsp4f2AOGYVzbL0+JVWK0pf1s7DZNFlmTDrUyBnjB3017qgjHQA1I1gk+M
iFovQ4TLY4B1E4MFnQ5U0Nw3JfmmCWWi1OpbvOOGB2CgxqAPAcvUIxSpNmWsrPT+
5zFHONJW1MO9k87b0WWezea0pnxDDAx87PbaZShBom4AlERMyxB9155u+lvqQGko
0KYaXw2Mlnj1cM29kxFZUxuq0I78tJeGMNWa3tAu3dOcTIAOFdnS9bvpbT1GCd0+
tA4v85gH461LjMbB3BOC2K0fhDdK1emWamj+XlvnsCxr2fLEmhhWGrH/LtNyycDN
WtILJL5ZKhgohQS721Y4ZvJugw79BDoFeoF2w+VFu5+k7vV0fa36ucc16TQOUaTo
a+p2wLXguxPaFLTdoq6tiAllvvxCjn7vf5boKgMJM1/RyoxqtRQnBBlxzDfvAB8K
JQ/jhnKrJ35PyG9ECWMKjrt3AlfZyYuxfuI6MuPVRK8Kmra+PEzxLxuVMf93UTJf
JpmC/TSwIbpEPonMM2zrGmN+gINMK/WP8oGMRMT72qHnL8Wl8TWQHyPWWb3q8vol
omFIKSRwOU/W/c4y1X3eowu0gpQqgVcuZW1ejIQcGEpmNASsY8XUl2SA/Via8jgu
jzcER8AcUh2uuF+HvHNaQH7YQUi7Lry8TAgsPE6A9o3J9Kn70S/gKggHFCiwufpQ
9aAzYUimzDNxcPXxWX/DC/H1DjzH54xhhF/3pkiT+q+kYxlF8PzaTm3ZRh4Ykazi
o8z6ovUQMs4Xbi387tv4zaXndCmS68ViuXL4eKzbScbZBdkoWI9aYH9FHprWGkBz
c/3Hs099FYu1R2QoXSRbCvZD3FBRNoKW9AhAxIdEFmthqprP9JbI+Xlz8hRgY27O
RMp105Z441H0wy3O/wlmb41nXCNLT5wxa9Rsf3hzlr3anU5+UfDm0zv/07ymqMXP
H+EMd62mmwaCrSdOjm0+/8LMLZzQwgCBFU1E+mWxDwwHoyqg1UsgLjvQJtTjbor3
LBLgq388uuSmffHKRXcytpkSWVUmwUMY/wf+2B9wCYsgWt6Hbx9ecLxBH2u7jGOe
+lgTehAipQ8IqdsVm3kPt5+Xuv1sejuA/PZKXWLkzO3jNgok/3Tl1y61FM0Y2/ug
k+pO/XgoZ2uNwG89rjFfxqA29WBf+y0j916UgOQs2JiH+xUHRz8YcOwM+UjZA4O0
lZTScnOr5SdzRy5FBBkEnZZtWkpOYOjsQR4hGZ0q9OGkAYs8+WOFT+gvqq3vbCYk
kWgIrXW+MLdGniOJyzr5b5nGPsbwfeU5rH9s4A2XX67khyFHe4vAyOI7xsDOAgej
a4VBswr/yRTX75MnxtCZ9BoCyrsaDb8uixn3d0gl38KXWkhBSwQHdNoGoxNlFH0O
4ozIw0lEe4lvR0GASOJxaatgd7+I2m3T7e93Jk72v745jvyfsdkL1KtPl1n9/LC1
UA9XyaCSVslBZBWawuT7mtS18bvnx3n1s6eoYi054N/1IXaZWp6ZT0NpwXVhBjLe
AbHai96lwC+FRQs52tg0HsA5a41iYBtCxVEGeHTa3iFxxivzfpHLDf5VgNkiuAdZ
b5xTN642P5l9vwOXoJ58G3XZrIlWpqKdM4wenMh+m1+Xa17gLgCO4EOM0DASY29A
O/4jk5mUd3GUDMyCdWhmsosB9bMZjREfaAqvUVh6J0muvs9ICs5cLY3DTiq4wXjn
bzozadYrhzGD1r9/kzOaj15dguGHWFi3dUCEi3fSrDVMee1w5S/NZE6fUA38lb0V
CeAPF1zH4yxaqyJqwn8Tcau0mNGmh+B02VnZihy+mWQ4ea740S+0fA10COt+EgSX
+spqvkkfmE1h/h7s+Sn66ygjON1iievS26vF/xQ+CSsilaPA/pzF6tzsNk9qpInV
UAPDFwOYPx05q24KdEArLeT0qfMmS+sYc91vOTUotpKEKD8p8EN+Ttsa4SdIW0YJ
FukUbUg9yLckfI5GSrvNK9uLqwHAI0eVO7BNtZo4h8876b+cpri376BVlmoCdH3R
YNwW641dgXwSf2kM6nLrwo5dP4YpbADjsuloCH2CZ9+tCx8P29RasXpAurD+KykB
4iMquRKxfGesDjShc/e+5qPY+Cw9PPyiyiZMBv7zOLcRyPvHVhNSPXKm7mNscdcL
CgDJ3EXaa8VA0D09dDrHvCJw0MkybriNYpsMf2tACn7siZhgzdH35NMeqD29DjiE
xKf1dQxMUKq6Croycj4DD+qth05VzA2+YCwGjeIGtBI25LFI/ikgoCWiCpZyLaA6
WyWuroBiobWcORBWvH3HRWOZN+Cu3vplAFQhKD9Jc1cEOaPFx1Xnm6mJFKqw3icC
YtDsz0cjKyaoVfY/M73WnkwBSMWbdvMZVZBpJMKdc+fQhKHY1XPl8qlC0l8iKJ4Y
dM7Why/Y/BXl2M2pSVOJM9KYsOOWbgSIzGbs5jTUeTLYAPEKbXtyqSIfCYjWzaRN
0SZUqt6Lrta9qtEQ58Bp34cp8SJpJxUNpqZ/p/VDKYfwnLcZzTE1ivn46o43wtpr
0VMYmzIL4ifD7FrSh+eiGnl9d/A16B0dHnmjW70h4dOBJowcXUF+ZeJrMkkx59Ae
oDiF62mhpbx7jQvAie0HUjJmcvfiEOLO/jUlHPx/LhsRSDzUuvogkaF2c8l3DNF+
fVzRfoz3OEE5kWoSsPQYd2kLDLtLUIgERA6764qQNfSToj/fBy4P/LFkxst/SoDZ
Qg70lE11o7sBqLy68yWZFQaqf7fpTBa4YNSJXzjiotNdUvkprIY6cDwS1dKUOiRN
vCWbDH54/TxUMqKkqiQ3kydIZQMX8yu8uY5ptxsmAJfIE4reptMl2NvZmrI2mzly
fzqX2kr/IKdr2Xo0DDc4fmdn5bA+VUDDuO5u8g8QN2C0R7bqwb9jguSk/hPalDcW
SLJMAv4HXHYSiDXBT3mexRpIAdi6RcOzIUmzp/V5B537KRtqdIHGDG62rw2e0vd0
OZDg5s2oR9NWdtS6V/sxUlfLGxdRWj6kyxQyJO9e/42wfZPPe2r9sL7tWvn44F4h
sCJnGBYrQ9fyAelUjrx2gb5G63qafGUyX+uV/54N50gD1ExFkWwYIFsMxN2eo97c
/IsrgEZnoFUgMWs5tbZxcQsUaKde5UXEUfKXalPVdA64P4BUQ1JiCsg5Px4k0G6K
COBguZ8qLkrqBvFb4WFsxjAqViSgJfHVvyoxfp8agprF/15ZCulk5DZCuLIGl8JE
WgZV4cZDHs8/pddZIuQOt4MQErqjxGZfyWRPRR04pEcRO7RwY3cUfWP2MHVM8AZJ
cC7KulzJdKEnzOIpQ3IxJw1UgGD+/oXPApNfkkilhe3GXgz5NB1MtmYtDVmOnUIA
4ZmuMBGrFlga5mAxPJoAntGKq2lqsI936GFhPeqpbUovW+aOvp//CmhSuBYghsy1
zK9Bws6Hzkn7pEXENSVHmUwtoPTQcCdg/oylub6YxdVcFJco+NRtlDltrGggVjTi
aOvTNruXpOJi+QcMFHgT1a4vD1jexa8tykT/UjE/u4vGzm8p2NiPvXjhKPm9ZnKt
AiY+vY45ZjEGhceBbAUyTpOBPkYecRGB837y0mOtOhZqlcwJnRGeyu///tUgk9m1
XpPTVjfwRleT9uFEQXu+qLeN0ws4o75TI89s/q7hiVnbmRQOjAdmFTUR0AggWLle
/YSOMc8sCShiZMPx5a6Q8dvSMjudnqdrIykkV6I697mBeOZ4k2j1jb1J/oFzVYYC
uJD9bEPAv4CXUSrSVqEuQlGbpHTio6fDeUa+kEAeSpln3sy55aHOff5RbThVLEYY
NKwPp1SSdCvVXBxZrHVjI8pZvxeBDklLqGM8cV6vVdEhckyBq8MnUGygKs4vJEs9
Aw2Y04sf6YxF4UWIU+Mv159b0ldSMABbSq6I4XMAObtx8gaqRdnGIzJsWKSBfQv8
vs0LG0+IDZBqW/LB/P8Pt/9JttAtqfNvQEapzq/0n8EpXagIc5D7qPySYowOdYVn
GL4y55ANSuYo9v2UiIVu/0OQ7alN5qkoDVhZdcZCY2WTsoRjcX9uMuSUTU0+RMJ0
cN64F+9YCo1+Iqw0nxci9xR+MKQuLe/pNDvUjpysO1Mp1O6wTH0NIdvOFfOWLoZJ
FEXAsWAI7Wn/9jpHbZAshJRKXpVqfqxsBNRiFsrLPrqtOPdGQtJRmTYQfFqKOmA2
2cNfowBn63hvMbthJsOfnbKoychjAZORTMyw+eTRHo+zecreMRn9R7M1WvAuOQoy
5uTz++J3CxhsYRFhO9XNKnpGK+jXXDNB3jRwxY3I66syR5haKCnBNbE5SS6Drp11
Evh8ODRLOFzebwF7PZf+3hxj8FJFhxKsFEDqdepR0CRtaw4+sc9VYSWPpwX5OpDL
SRLqfxBk++zsb4BQgz+MdS9fv7EH2lhzxq5/dxtMGZMzfoWpCdzVFwpsvNQiSRKg
y4p+F+kcyarvbOekMXW/DvZCk+FRuDkvwxmgsSmK1ftOBJeAqd/RXgAx2C9m1zVu
7mxV7FMDWocwTTWwQuOLicR6CAU34zsauxwWSP6iYLV5a+AYQAlkrcccvaKLpV8Q
qM11wAHcfI/7yBstnTSBuDS+U/cjwRaunAjnWuayXdeQJsr2xeaSkSjaXe31MB1e
34qcm0MTLvU2iU9yLc4tNq2P+AP0pmmpuVh+2E1e0YRn1O/Bl2LbnMAvbWd1FFsy
8AS7q1ZKNVN83maCE6k2mWuIWy9d1Dcn9IHZhvJiRI9hqMnVk8ZmWPOtEgdhb/Bb
njqV/3nzTRw5LdRuPA3kyGem29+naPxp34FfYFgpj/fhoky+D/TdlnIuDa1dKUm1
LVGQQnboFbXefhH9t9XQZsh99BbtDo6M+ltL7vKhItFcIOzrkxhbuta9n5VYk8hQ
KVPPLN5T1opY4CyfHzXpwQ7T8oMfScEcwmJlC1w02MKEfRcEFHTn+yopG4dfk4Cl
DF27NM6Trb7XYDysuUabM2vXu5oeMcn4KciWfCqBvPRFjGFpBQptJKgk80daNHy5
s8hg/W5kW+liFuXFCOyk7muJTGC+uH5PITTM6WULMtqf4Y/eLOA1OU5LSfRTCFrF
djVsFj8WFj+bWmKOGBkZ0Z1nMRjFu/zZJwpfgds9qaM38WcDu3Yn0B1snd0ch9nu
Z89kaOUCgMYWMs8n5rW+LtZKssryZT3q4yMWF57BxoExUnYJlSc0q64vvgmc0leQ
JkL3wtTGc3wm/P9iWar+G8jnW6MUKTQN8I59pOs89cQGbDTVPkSNDUBJ4PbtY31k
mpUGhvJpfXxfP6yvfzsmbulBO+79SYEsKM05R3Dt+dDYEKgn3dE0mQlxDrzsWSgY
gvu1KHtSRHiP8gPukQtIP5gzJJyfWcWf3DS4h6kpqAUk9ruC4Xnd1IXDp++b2Wej
SsPi1bWg1DILYwIqrMlaLsy2Bnz02UVGrs2Il74pVcKUmgo6iUbSbs9+sWfIM9o3
cWD0sx7vC7zRtX9nvWrXv/DF128JNnnjUiLf3n0sMY5et8XH10LN+tkLSVDH6y6y
UQbMWN+J5bWb4t+3ZncSuOYwiPzO616veeYqBqIZyl7XIF4m0opKcYuHPcbavCVh
q5eu2zK73ID8s6Q0EHmXTikyLIHtE/+G3FfSa848Gu5HaX3ktDx5uKdQygOEqlxd
dT6tHelalDAY8bTHUHENn+YeCsLqWP1g7/rWu0GcG4ka6FYv95N2+2Lvr6bnjawy
9KS6otP+Sh8biCRqaZmNRcsd4KDbjJQyZPxxaa8Uztsik6GUuiL90eIdyomSGz7q
BDeaatLfLOswaYp5/Cmia81AjM7B3fXctTDsM5/NfelHs+9WUkzGL4oZAqjxwjfg
I7ifjLJnFjy/GWBkZmBMTjDwpgTZ/FritRpayUiLlektLS7sD8xqCMnMJikyH9XQ
9Jg1weHn/6MZfchwmeS/2L13J9nJ57C8oxiu379WkLDyXROkcfvqoyC7LW3jJzO0
ofHftu50LXf+G/X628Cf67bfJZenj2xOAyyDu3nI4uQwsNTNhhVOoh0OqOHSV0IZ
NKtf1i1rlv240KP863Gry6k5C3dwo0QekKaEH0e4LtymJJLf0xcwN/tAyaUWIew0
ISz8XKzNupMaNJiApt22rC4uRbX0yrJAGOvSD8iBV7e8Hu6y21yy5FIP1vHaPJ4p
k3GJnNMf6lu8iRcudgVyK/TAGXYzaDwy9V59DdNNdGZwgSmOlEbyY8u2JrXvCqOE
/7v7emVinPMZ+q7VPtk7oS1BGjv/Aem8DhbRopDEVkm2nAmEscTiwLZvScqBR6YH
RqwmPT2LoRI1aGs+0QA6af+p4WBEbLQNq8lPgkpP8c4ksZD5pAX/izIDlRUDInXq
j3av+yANKQJ0ywOeoDLeB0ZmzctUJxzV6WATodlXyfeuLnT7//RBUJu8SjbzT76Q
v5swba4H323ro4/qY10J6cQfx3KPbBwpwDR00tq1XN3vjG1otGRj2TIVYJOAW5n3
MKe9d6HS/ojWyBgUlxxXHbrty4ltFrTo+bhYKSdvzLpUWRZ9wT6V3WakMC/2dTPJ
WPafogKZAIeSw4b4o/YC4pldws0vLoC9c2prCX1yLCpKrBpa2UnX9e+LcGj0v69b
5p70el4d57IieqIMiUHejJbmJfyc2QRQafcHjgwaXqlAig04ISdETlt7zWZzeAI0
p607n0nPdqIuUtw3aSX0nVIvYwS4XbmMHtePp5yRhvKiviD531T/NhGlxjDiAC/B
oa7cPdxcMcS7SjROBjqJgPIRofAQIAOptB2MELY/QbdYLdyqlN1YIpbfZYyS0vQ/
XIyGhOkMyUjawQfptdWvvXNsWCO8hQPzWNFK/x8qiDUOY4HVeOhGCL9kW0Ue0r3S
ilJVyMwieYFiBjw161tO3AOBIS3PJFYAkhIUjwilwBf2mBtmcH93SZbRwrDztRkJ
bnUpI2MuqUh3+Gol3mnjUwh+FFKssV7SnZsdYwBpRavJpgEC282pY5lFIY4RXsNu
1UDx0oqEbVeBC8BQKNzwZt6MwIfkviXEHBH/zhZ8Nj14c0r+UdonueV0MfaWwV2y
LcYVXhV/UEhgAF+nj6ju/QSk949JfKEUmzPVI58Hr9xsOFftLMAZeta03Bfo1jZd
SDpKW1fm2mVr9R2a4GWuExJmYdogH0EGMSbaiL7mb2BdHmuxFDgZNRcb+MgS8zUJ
Enuq1e3Rs0y53Z4eudcM/gxnPp/ew6ATYZgRZWx5hbtQma0cf071mVrQrLe+zIX8
wI6GBr/5um1HC2PPCddx18gYDgqahp1nujOPHbHaUO3IEsMjfIh8x3olt0YvLaQj
dDpNRpjS3MEPDNbWnaDUN9zeQBPovF3SsN7F8EwP+9p/8l/Afvg34SryMfR0YJoj
3kNlT6wKbPPY6N8sydmjKSD3DQktOQyXsYp0Vx4VuJJSfF/1ZdkYyXRxzODyB25R
1EPaL3+xVJvCqOMnmrSJ9ygvzXyTBSzBE6/WU1drlXy9mUFqrpY0si7b7T3jRMXZ
bYxq9YgFrbiopaM4zvrf/Uy/EGCl3ehbKDN5w0VL/Xasq79jc/uJVegIgDrL5c6B
g+I7yLRAil6EfkEU3T9pTCDtFre1Qds4jV68xCXpAg2dA35zFxJGr4m3Y9R42VVq
qeM4dmh228bnkg4VPdrxnj1WhJhC7SkbXYcp13A0zBSe1Y9jsCWqF/7a5XAaBZZy
yisa4RUtPtTMNsI53iHSqF1DY3C4RTl76kmk7oDdaK3xxDobSc9Ge1JnWzp5VsfL
BlUVDlqWSFx7Z2P51+NMbxcn3+lyLRPwhYkVolSzqeYbSCauDygrauVLWc/7hjhf
q6u+Rzba+YkrZI4ip3Dp/2FgdLgxoac/ziiHhl2H6FBAEQ/uaLBeKuW3gPa8Qh7W
DbsICX5VoDQQwuZ0U35L85WGIbB5/BnaS8AjX1h87oZvu8rkGltg2eisQs/zvbF9
Ri0w95pme/rf1PKaminlsb1+I0aDS/qQudxMvynbOwEbS5dIz5Fz6ImDWR/yCCLK
S3jz9LJDvv3Nnr3KDpufVg5dhIUtoV6qvymSChJdy8EqOnv9rpiB6RRl7fV5XpsH
qW4Xk3XY5IJX/sL2RbgXF6FMQ69I/nEIc6SMHuPNq010tnygTV+Dp6HmtbMf8fyh
eSGJKBr0s3taZjzSN23VdsDlSkXiul2mQYuAf0ibYDlfDGck3utKmxR8k7IrMXLA
CJoLYQe69c1xgWyPgMrsV/D6UEOzch1fOftFCY9Fz52TCQ7MMhU+0AAeO/PvI/Jj
XQU/8pFntd+p+u/avecDCyDyLuCc7kU9j6cMYm+kWt7xfCSsIcBEWNP7owXI7eI1
G0Dt1Rzh996M4dS62NhEhiuFJ+jW/ZlYPApPwwN/fA7Yb0q++quWMePBbOE+LGWQ
DMm9Xhsj1XnvOOUQE7SHnMhn0kGNdviBb/uhkumxZT4rZG2ZDu05hrEEV1zsEweo
QWCgjFaZ90UfFw02AkFamgZxFWsDU1UTb56PwEkqP2wdXEsRp2cBlXqTfOzyATEa
vJPzFJ46X1Vrfxzazm9cI5CCV6Z5nxrD2NP3u+kbhH9WbkXZt4FljyB/5FRf8wNl
Q6FYerttyarpeKHnHwir/rd7pQD0VZVDFosJ1PRB5R58XZtfYdak9OdgVFtoug1M
8oSmPGaFF4M2bW84ZQMuLWtsFGKMVXLU0EZLDb4EDyZWY35ic3TeKcsya8JkmCCF
iggMcGwAlkRjlXmsnwFUWkym9wq1wm82SDGylmWErUuoQHKAWIorNZdLHqZW3uwC
AOSkF4xhJzioyBv8pD/zNX8QL6AHVAlYSrOv2oqXsGhFriQofezte91NzBEUAqpM
GJkZzf337oGB0xuUbjGCM3ZKBRh3hAB4tBz/yLVYRGiB5nqxuWYVWRhJijookGte
JJMu2h+Gy8J3CFOo7CAkzb2/KFhpwKykTNCIZjAH3OgRn0tvAB4EC31xJUE3HUuO
Fva7VU5feOVjiEdTP4F71ffCFH5OIKP/NraXqQaDuW0xxstDbux5SsU7ROXiBQSF
0WaupfC03LTzE1EcKLX/JBE347XuTU6X0xWzD223kOHMmuot3QuzT5u5IjB407XU
KLaWKReM3lOB6hjzF7XYF+6Ye4Cg3EVDthcK8yB70UzyCRWzptaeVeTLTw51105x
QTEoM2p9r3hk6GGG3oWMEew4Ba9dzDkryDy9leWQFJ1vBfYpmXMCXVyn3HASAPUV
DUoubMOFChlRhMN4R2nJM23gPnqeKEwXQqMdAM8scYRgvqQiWsess3k+lgXGtTEB
PlgjyrvB9dF2mzs+SEgOnh4eE9vcvVmCo8qJQEmeidR/t+xBFxI11/hMRpddUr7i
CAU2VnOYEFox80rl0k9l8OkCYFuf+3U9C84PPR3OP7t6P17DlLNKEF1nBsTS96Hz
utg2QU4YA4m40yGGXUMe7yVT68+kjyybatIGDmPIB+0S7tyjR7w22YdubaaruC1q
9Dm5yDqwvAGxBJsMCxpKeMBzcIjI3ahgVPYJP66e8J3UKorn2o6ywAN9DJ5hGvjR
1MoDbNTCpPgWF3lLjOS/sj9ezFG3GQdpjFI0mryZ7eXWEeV1y9rOtP1xeXjGN73x
TYM8ufPYuPviMkX3NfFGW+uLPT0W9GnxQ33q/dHezhe4mKw9OBZ4ljTySBvQ0EpB
Nv1rGTKMIlwqm9IBVolGrTTGgx5Sasf1uXcqbyzoBuGeYvb8kBqENncJlI175jBj
GPgxmy9kQp7RTL/8z8TkCBMXWYLuhin/oD4GptwJPgLjy+kidXXniugls7pb9jeT
inaJ50ERFBSmzF7L3Mp/+nsz0qHrIAiNsqsVsL6SeN1KHsDfJWSygRLZVGR7U6eu
uwXmAx5kug60jftgYZc0zfRpddK8WmMztyEm/Lx/i8q0aM8nLtMGPD7bVy2Z8jtd
8AnJ9I3rRcS3UsdduqzyQWei6SN4lGYpUZ/2qR7Zt+G1mv8qn0ntKcuDFoMGxEKL
QnYRz6bBiuLB8NwnlHjfVxhp7RTJv/hCFfGSaQxFVyfCGaWSkDWCG0TEXOkqYPlx
YInQu2f06ty5Ocdn2NEYFdygs7CS5/mBYQaQctiB+ePFmXfKlU76kzR2Xc+1Yiks
QkuoXaW3HOLIpkNsJl7nQqFI/vj8BquV6MHNNM8tnm0ZoWZVENhuzYZkRjKCsiH9
QIzONwtBbK/q7jcwQONwXEDeMfYzQ9E5NOhATwii/Z0Hks4mA9mxMxiVsh9/Pysh
OeHWTjfn3yzKbOj5t7xlcmOAFQbfmuJZ8VDlvU4SVIHmfsTw46kIDoodvBIkA6zC
SoAzNGjQzBlnef6OmjEjtrpLDp4EdCWxTyfPMRN4DL1cDflLLZUFiQauULgfAnWX
aIJXGVjoI9xRfxYGs0DYFehz2IUUOqGTndKQ+pQX15Yczr2UfuNsGajZh6wDkrsM
qx3MzGFlEn5w/c/hdNlyPWneiowibO0482g3b7yjxfbDwJLZf5PT4wFkIw3TS8Qu
CDtzg5fHpLno3clSz98wdMhJTIiWTUbMjm/UbI73mmOAVkJIxc6b8gEI6mmH2FBH
wNtIxnwBaEdhVifigLy5MsKAIU76SmAz4vRxa5V225D6QPQPJk13NOhkGou2jN5f
v704mHzBX3NregYE+bsPRqXZdt7hudhAjc9xrXCUsHEJrDVouBWSPKZVPb5GerrB
MIoZIE2hI0xZ+1DQhMtd+AZgtk8PuawtdGUU8tn2hLNBijVJ/6/JSSdBK94zOcRC
rzAOlfieRQLYtwFonn1d6kMUdRg3pwremK5RaMCNbifFlWL62kAEf6/0heKu/fCW
A71Qt1B9G0AfilHxQLt8DxdhGIkdHy1vlF1FDfsbzdKK4mXklMjx0MP7mfzLxEyQ
YuipizqtG/x3eGBdMIDYH5AzIT6WEGMTH6U1/C75LvkiyAIby0egT6CiTwbH6yUX
RNpQKJHQXF0YiVgcmyuJIeUMrVxCuLd5z4HvFMNt1Z3Rm5xsInTOQZbER7r5sf2X
VvhNJdCx3kWdcYZ3/wREtJmy/1TJacY4yeYgZ6AoYzdDmAkVcGMl0fqWI4/UbSWQ
M/Xq/bCyJ56eQ//LgxF8UByVZGYIeRqaOXkniYIVZcHCh9AuVgsNexYl7ymLsGwe
FU91eqn3sLtghPJs/6ikkPUSB71/Hdsn5uKxbkDGbrKFlcC/dYQbA0UwDgxZJVPl
BitAXtyM+K7Nma3ftUPLdTUTcX9P+dmQ2PPLeG4djhynS4EFol5CyB6445Dfi+31
NQuAKJ3jWAbfZc6Sys9r9SHEYSrIoWd5gcDb5MFYgtOjo0timAPq28vh4sbFj0iV
LAYO+XGro/9YPUSi5J+1Uru/r5Frb1RSmIlwD+bgG1AuxV1/VDo03A9/6u/dttsC
294/NgE6iE1IiDDIVD9KItXtywzxwT+hKlOk+7cY5yqJEiA9phVtLghUWmlBOEtv
vdwkkGdzwCTVrZxZ7xx0Vlql0C5CraMziOajmxR7qnAEUKvoYUNmTZw0uGdeuL+G
yJYwT4EqB0G+p9ykUbp+EOuoXAbZvyLeLTo6X561pTA4SqWPCe/YBFkmB9zJzLee
c66iks/fgevOWqkeeThS1wAzEexO9kPM88bTKyG9hfVJjTDtqyMQUmpbLFTLEMk6
j7xYMBakkIzWTZGg+tjwzDC777WwXS/UHj49OYbT9Al2OZ7p3pI6cqAa+IBWUCFw
cE9Y7o5om7fbkNbTpuMxEstY9CKvZhz7c6CRRhMzZNw014aRQFjhu4xNsZGVH8qR
efy/KZ4xnFy2pjq3muvAi+yG935utCnzsda148QKyJRxqOfZuFKKGcnJdPyLUJsw
I5LHESf7cUrBV1PjoxNuYzATOL21zNUxWYQiUSXBom4l1lJz2oF7uzVcxfIgR7b7
NcZXPMSygVWRxzviptjkGC0NbEdrUFBVOQF5JFZQSTQ4YCiAH+VuUZOAVB9Zqauj
DBc+CGgYBlPZIVO604N3cCoICFUxG2yCW8WNPmSEWukKw0aDC9tLRv1b9uFjP0jL
ybPUiSS9FF2HU7CYYmQvw0/NPoDBVBcxD/jD6LY6C3bi628SvMVb7ChWV0FRDbaN
TYKFcxeRymbjR4Q7ORDkvvPXUXRLao1FMLkII+sCiosTltlnZt/887GfFaBuzIMy
H7N8u3l9MI6qZiMVTnVyAyjfqPuxy5OIAY4P+EQB2udvqn0tTPXVmxWFJPjZCdRa
8ixAv0eTOO7pbD4+UHjXPbXWOHDrjyqCd3ZUuDDTkEnhcVMFaCzccXu4wSVSC/ul
PbCicnlHXuM5hjRdGfBk1VrrdAFNamUIHUsp0ipmR6wBBvdpiLWPH2kDD3uXoQUQ
Udd2ItewjA4XBY7TcgDjXWUEGxWkcZ6xDfQNVOX0UCy2V14Im2kUGEl9zpgo93/j
xp06Kr/QKazPANTs9NAWROgXlUSvKthrr4Gc387DzmYXgPRzFcsPi//DAHTy8El5
dbQgxllfe6984lcTDbwn3etGY3y2RKQ0p38+qxxx5vq2LgTm/aVT7Sg1l/VjmA75
tOP5TLpTFAbNQAfZ1fh5Zd/Tq9wNPr2FQxqJSTdr849aMjwaa9YAZOJmZrYYnU1/
R2sLg4ATiKvn3r0+ADTKrX6fpOsNfWMyGRMGeYAlMJ8feO/gXtgjEj89KCmzbtM1
mbRep1kY3ByDvM7ecLCL7rectdcQoGcjkwhFzbA/68UA5zRzBK/tdXlIJbLJ/KxS
7CnIzSdqgCvdc9L4vffNbpfy8AfsIxjCsNDchwccIT7meKIpJz0BSG3PMZztj0pJ
shKmKXPtpQ5EDvvGbNvQaXvNJ7/OeCKpQy32eAffMb8vgTVs7uvRXxrX3jSmIzTD
DWRXQ8vWrGUhJ3iORNhtoX6CSOnsm6FUb3rZFhhEIXqFOS/Z29ducpE3iXMuOTqN
mZdxL/LyB6erJZn45H39NFqcXq3YBBXy7S/h4oQGTZb8h8JKuD/rKUVMMDiDDSFP
r1O6YZsWRNV2LBO2yUI7EyLs0cYz35gQWtfhUQUOMi7FPExTlBQGIoLADWR9lKcK
DexYd8jHdf3pkdiCctppnOd+x3c6oumSgjQRF2Oqvj6Wrn7kM/QfFWjKxB00Nllw
6g9N7Ur+jZ5Z6OfJKOY6Ag287wdMbWLMTaKQxrG3d0hvZyN4um9ln7dUuTdqKv/7
3cLD1ar3Z4uC6iBTeNVqAiJQ4ZMC9bTbGD17gqsVSYfB0oWj5e8sHcx5QvXsH3r9
0sJ+Nf+n70mIs8tNbZ+Iik7RiNSIaoeQd1Gu6czV5p3HMdLt4OUJfWA4SZr1rVFC
CJCZNjbu2zd43TKGJfVnaOwm2mpIoPaVonBPkHRiZWW933cUCT7Gw/8GquURb/Cp
LkBjonIVbw5wTIqmbL8SjT4vmzO3zeKCuiptv+nI6BmF/hM5PT0zummhRjAJWLSi
zGyQh2ejDunCJKhFfoVqwxlFcgIiUGGf7bitTkBCA5KecpPyJjC7E8rk58KgGOHe
pv2VqthTCuPCCUzoQQG7qtZFjskhakrokJqW4V6KV8UgJgEfFpRJuD9OSKfFxk5F
VGBILRwU7mYh5r+n92OScS3IniwlB60j2fW2CT4BruTQzobpAhaajg1i7o7zVcIs
0tu47EEwnLQwYquezG+sKudZxq78BWvkKBKIg0DAXBj/RYx+EYD6i8VgvNkA8iTa
5T/IMrlCTfdvmVyCWp6+vHFMO5qD36t6jcOSce89fSmVaoC5yRvhvYMf3JWVvJYb
3jj4KSc2XaqBIQLfYLrHMjXFboSZBOEA+U9G4sHn6HjKM3qGlx0xnWWJWf6/2ns1
3fvJJg29dMU/+9laNzE893REhxdX+MpsqZq8LnkLxWjulj/3STHd7EKuW79nK92G
2CRjD0xLfzrYivsa+u6nyM2Ony0ftkl9v4ZXQ2tzZcCSuY44otsNEY4/6ixtECli
uS/4aN7uW8cmivRy7PkOd3O4/0qYcQB5SRWYGAulPC5W6Pus11OLmRCF5ao+7pBa
u1BRyDdAA3IIV/O3BuItVBYf8aUrN+0S3thxIhnuTxB2NfvfhPRevmHs351DT8gJ
mOOsPCMJMeoCDio6hRIdKwBRepdLPIRx5LD4gtROovWy0OnSZGEgZHgC5YF3APHR
7tp1OuYZ3c6HtV2hqy9n4B15FrhwuPHeRXMNqnQi9ROma7mAkiAsZ8ofXbHuJk44
oOHV5BLEoL6AzT5EgWKRfdIquxozsFONmv8bzh3l9EXHurVpDGrsDQKNsK447qu9
5mOhwxElO7r96Ebnme03H/lnJIRjCM4UBs846/iyelvDSqyLbjWYizpXhoi4g/e6
x0N7fjKEiWTKzq9bPpHu4HXAXFXXc7M31KX5P7RpuHZPoWaxHIJycRWfZpFWuOml
B/qiZyXyR6x0VacFb6KKqDx+vgNOuez/eVkhTUwd9Kf1oNhIlNCAr5Tn8Ig6cKwi
YZuSl7kkbUObP3AKZqraQoLZ1oaAw1wtXdCYivmmc89j7QFxukkd88PnA1ZSsQYk
CggZq30bqs4gH4VLHov9oIjaqLVO7blV9S5TTIC56tb6Mt+dkbutlMD/u6JG+bIb
f8HbAwoDkz71UzkQPAVUmDjpXfXYifWGa7ybrVAlMaZEdk+mYBvUTGJDszvOLu0x
TtAYaOdYFY/wCDNZRMu1U1wu2WbST8+cOv/kaHXZQXOCA62p8ZaD1yj+gV5Jw/hj
pPs3j66wfJ8SuHkTGeE84kwGfutrcamHR3kruXckMh/h0VQXgEP94P46PNsdyxC4
xQ51Ovkv3Wu/HOD0IPhXHGt7glZLmqnSKS6YL57aADPtu38e9CiAyYD5k4ZL+dp5
Pq5pmX5RIXkMi6W+DKl1g7WoW0pGg9ZogKVVuXhgopTCZuMRa/2Q6ZSmmkQVks/N
6eBGWNhrZ8mlpzpFUR9+z/+6rM36KwhDXPGyfdnd9bJjq9UT7+TE/TvMnY9dpOzf
sKDR9Ugox2K6y90SUz0kOyKCcsDbek8WH0IxRVSZBu0ijFPTW9FaCCRcHhukcRla
0oQuA5w6bPUCmOsr0x3aNcczgaKCnyU88KCIgWGRj3ckUcQJ3a1MK4qvGlOgxBDN
wOd4Cx1PrkbhlcacgVYbHgCKj+fmugBxkyqmFWDq+G1+ap5LyLhv3FgGJXht7v+R
a416o68rijhEI1pQyiybPOs01vMtpRLYmmNr460J9UIkq/5IG2vxfMy0tM0bVxXG
c1SCgAcvZpLSPGxI1W4yZshrAAowT9lJWkwst3XTWSmwuRdMTeCxw7GsRzoDrnVb
xYXj0Kv3rmEld4P9m8Oah1vKFimxFzlCP2b18rX8ZaPnrzMp/sG1X5axNQYD3Xwb
YbTdpcXjPCdLsJx0VkpJRi0RhVYnwVJ7LbDoMPvoDtAtopwz1EgIVenCL23dwoAy
syTeirx581fsug2unyfcUrSHHB315yKFcncfyz32KZKA94FbTrrBM5Ew1MTLHins
92bfmaalzUn63VaZEJHuX7R1dV1SqFqRWD5c2Fij2TLl3nqwJXh7ivc9oUVEr9PT
dwQYGuv5NZ2Lu69YWIV/X7kKqwz4iM0qnGrmTwU5VvfQGNM/j3pdrB2HGmRkni+e
ygcMofA5JlulhsOvBVk9rSE1jlMdAvymyfXedKZRLDtjP8mq1+I6dgnXgCYOabLG
6b9wBwSmHjCFVAfXzOHwjQEpko471udwedirAzigP48nLHatoxoEVnfrxIdgvolU
d2smeJQsuHPU6gYdCOy+dp5ntX1C8kAuvXSkkeawWV3tc3ETRA5EzmRXxrqmhzp/
dQuw1n04n0iDeG3AMjA+luhtJqMHTtWD0sjhzagSPFolQCZfKCDcD6ucWEluSgJy
gPo1o13C0AiAU7wLXDfjO9zraTjMkfxfbuk9iiztrw6DYr62PKhUoo625BhHgYnQ
fv/Gyzvy7q5gb6arYcMmOe1pGaXqlYKtfyiJskcKAftb9xkqmfVw7jwOvWzXGiFn
HIEkFawD/zkl1Xf+RFGsWbK6mJBu7tGVoVSoP9ArR+J+mdpWIg18BTuBuhybR+w5
/YxmGwv6BGocCAt0K56HtTuDvgm0rETOW27NdSMJb2TlpO38O/hPkMdUPeHEYcsI
O41F1D6nEsQaN2r7zjgY4hlgXKR2OrYZOzz0Vc5M4/vql1VktE6Gpsat4IVqkz+l
50M+ZzM/J8/b9Fz6C9d8RJ/0KMjQGjpLLgrWrpixmzovPrygZaa1fjCTGbrycfTS
C/tggpSfQnHzJrT7ZtyTuExLOEIke1UFdUzR43nEdPqHFls8C7HL2xHT4p/KWJMX
SBoWr1Mg97/5bf/u9J7SL2Ype4J6uuNbjknSQjmFK6M87zg1qUcSbglXmfs+SUhd
PYFe/ipfsR6x5tfXRw4zD6D591qO8uVRU0WKKQZID0frgoREUGiMYb6YhdPyOSNH
gBElNxFvm9/79Ejb0En7uR6QVNXxGs0IfOfSl06BSCJhRS+EOpgezXOEWzxG6yIL
VQZeZKyHLu7ECdPzuaJtt5V/iLIB3WO3e1KRJg+wHotnCutlIRUBFD+ZjXIB0FZH
X1iCC3Cjsg8gpYY+IiZU+ITQblbYT3MWJsT1rhlo7H3sZmxB+0amf1cUK6IJy2EK
DOB2sAbdXAoXrZ6qEAqQKVHE3IXJ3A5nc8rLwHDwyiH5GcPOzGgUW2K//xNvQG/k
dpZKTNmkd10p7/dXRAENGL12ZLS3/EvfFtVw1tP56weIcld5e+rtoG8B0c1Ybkw0
VPa4jVuna47h8atg1ZolGlz8Bu5eFGGAV2/O3RJOBDVHhdiZhaoZcs7dA++rHZGw
FDnPmnPdCMQwI5npM0/6jNkAYaRK2/3X3m16OIEJGUsqqdQV2/0M+3vrBu6HlM32
jnGwNMxFDA6SbMAl2yHvXrQi4lqwqbjyeCuEaEk+Aoxs2JtNcBog+RVq5Pa1Gxsp
ytokUqu9U4UkVsqBQNjaZSi8cr8xZdCfJpL7giIQaFS58t5foBm5hleSI8qBqOtk
ziUOhbVbaI58lc0vXRO/aXWZyIZT8jDpb0tar/H3YsNlHHBmDyBbkJ8ZdT9QhxuE
Qqan4nAwh5BD3q2ObppqxFo2Grq4CRX14BurOJDp0TYLrjYMI4x7/eB9bL3ctLAg
EL15xsfMOnqVDP9MM0Pf+j8js7nCgTRmEyBmVP5PC8rqmcEGvjZcxatS/Hbzi99C
oMYzSdPgRCX5siTI9lUOTSp+5AuyhqNViX2q9zRtZ3mahWQcYzgVsrNuv3FjBVAG
doIejbkwVOiiYfLYe38SeFK5my2TXiRohCkGNeuhwQ5J8sovNyPepi+A+cfskiT2
dvm8wV/KQcHqeXm2nsXU7EXmlt2QazajxZtsRGKatyDRpJYoALTlnIPtdZcAc7ad
X6VJsBQjTtzxBQ3Y0MYQ43fSKnDFplipM9ik2TQYRRieoY24DrpJdEwsP7hSPSuW
FXKqkeN0Ykl73WFASaps9IJD4fzwUEZFDBHp6BixuD5q946P5KOb5YXomw2gU0UI
uJt4YB33EZsmAGBeR+haHjBc0U4mvzyXEpkgBjky4R52woXNdFOWhNsijw29HEhh
4uv6hMGUgXkaKMlhSUTzslaZYk+L/wqQFvxgOQ0rmYJNdVmwOEzL0xwbLguR4FqU
aF2LoL+ivPEh7pvPZJ9J/uMFNuufiqUhsRLuloyzk5JNhl+3zJBI5gDqpTzj7862
GfsR9vS4h0fk01oTMl6jsl9KGWsUnjn+gIeLgM8V2jKu1qe4Ccwg0IAMnrSShd/l
FkkhyeD7gzYOYszzPEShUrkiioQXGrqvBTaMvBz9IRjLZkqo7txO5q542jx3A7/m
I2J1jumXdQzXaJBTXXLDKFsNiIb4YFF+XNQzEEnz9TE4sIZrTz288nxafNGd/pVT
W+3iPKoBns2cLF1TmVH7j/PvbSIPAi3kikc0+f3WCUU94adqfZ24JBybZrSl9ycn
rKd5BeksCW916itQ0I8gyGC84RvnMfr9WwCjI+2rWVkQxhEp+ljQvBSV9XdDrE+P
yuo4xLDYoThrVbAv7Hsd6RO8oCx198G0PyC8Fvrt3py2O9SailH1XW++UrDZDpB8
NBsSNlzJ0jer6Sie3kbs7UvVZl6fuP5rRJHvuUIYYUMbSNXZ2Hybw4ZW6oV0UXbg
Gi59gxaV885mRxBiB0xdZ0QR88nUrhztUP36IegUjThmvjSVunFtWSlaZprQSMkC
hrcxxDeRQ26Q7JyKYYgIFVvUPEVmhCGMkwd0xBkRdv8YYesv8IdHDqj/3+bZFeyu
MWT0PuJvCL1COfqXXNvu8wlNPFNL5K5tMd9aD22BGj7Ci2xjZdrwijalPjzb1H8C
BjHQT3KC3lh7tn0e0tOUmmvEv/pqE/rnMTads4s8Mx6cj76vs6LixzCEq9EaQ6yZ
SCSIaSjmV1cwF1Ur+5KAIyiiZNGNVpVXIkff00StZPiT38CeLAwDb+4HNIp43Ymw
snEMpDO2lVwqWdZcQ8O41FbaC90onw4WDcyT9Zptg5bmHZhc76WlsMw81/xHHZTz
0kOWkmeG6kHwGjnd08XRtDqFGqnos0IAdN1PFoPun0aod8qPXSXffgW+4mviCULr
1PlJj73+PzHTZ+R4GL839nIpiFUyikJZn4mqPziwTqTcbBIip1eilYEDLjWkbfLF
YozE1XTVReE+lTNBKeyiO2JgL0kk/bU0AsITlHxnPrSZMIo2mNfF76SSGOAsNTeS
+Wfg2JxNzKrpMiK5mgu03FOzIsmGCRRB1FeVVIq4oUiKaeGPAILF5sE73G+aq0XU
ipZSwl8MsQxQjuVkBVrU3OwozxEPLlD+fTbHyQ7/ICm1t6Ne6Tgu5B95+mB23yCi
3Ho0W1R+2+QsemPFuuN7lcOQeEdU8Sf8lJ+BnI2NR95YJc8n4uR8i5hP6Z3kttm4
d/1oBhWiQqtUA8cd1W3aekg+lWRpkg7NSEcd1cCDCBwKWBzLWM7n6WYfGKcJMSsc
iSQp1DXnHkXBi1927fPAkFDVQfhDvbmk6jQv8eau0qIctbcMS/RBHrAneurpbnh4
I5KyY+1rBwKPK00d1umTCOLCkxDI7Yz1KlvT6uZMS9OTDg8u08nbpe+NvZVcnyt2
ArYgWDhhm6fs3AABXow4XiLpxzj5LsE46+HZT3RNQW7jTJ+zu5FZlUO9evb0I+bt
Uq3r49g5AbBJMoWFx8gRMyf9N+ff8/T+xrRICzOjWMWEs/kW1T44OYXuxdL4e148
ZDRoLpVHTuziHa1l0ZiJtVNVjPtHBSRnY5H1DoVYqhtWpabKhS7HEAxkucLe0z0Z
w4YziCb6ty7kc5rnCqqq1k0x5uxr3Eagj3WhI8lycARF/W215GHKBfEVisMfEuza
XkQ/OA/DEga5S8o1Xg0JV7Gh7zVxuzZ3zR5ZQedMBwRi77vcUWjmBcdBQ2qhynQU
+2lCMyS2hq81x5AX7h4ljFPDb5xFsZsHs8VccB88XTzFoL601Mx5ZdOpL2TS/fbS
FP0G2Rn/2Oxwy8qNzgUwl4oZoN9WS7qeF9EHid4Y33J0HndAQZivoAD9gSQVsfXR
/ssLLwdkTm1002FbIFEo6STj5g0EcY+350sV0YLEY9ZFaiUklt9DCniIcvk6YS0M
AW9yoGUWVo9sAAdKciZs6b5uZ39FI/RpkeyFUaW5NqfVJgo+X0ggWNm7En/6tJBc
wZKhHOUGSCIQffYMvx9Lz5KLuJXV4A0HC5o85rFWQF8HFETrqwfuGw0Gg72fcxuV
GP0F+K3ZYfnOq0nOsktItUWgntyVidlshnMWsx9ra/DFPYfQNvvPT+gDEmGtkxor
+l5ZbWxtaxQl3YuoBONvzJbqWyiBxiEhU/FlzdQcqW2wo0LSKq2OBdmRm2qAXMMO
GlCqdv4xGVKpEGQ0G+tL3TB5MumR5OtOCyvGlPR3I8GM9Wzb5K7W6OH9s0lRqsYe
UalOp6R87k2khW1UXRBSq7rT2pbKAGHQAwvfv6xCKI1NiBZMLCYTvExwLDM4+Gxw
rWIYYBAybcPTeWSWngVJtifMpLqUMKNNPax/3w+mH3PplToG3zSo27uqR2Gxqwn/
2gdPRw/AOYWcKA2NtY19KMDdyXhG+VUilzOuJHDTMQTizSfjisqgRN1euf1oUAKt
oKV2W55TrRsr5KKgredcShH3OlH62uOvG6UQJV80Q4uk7CsWxwxyq0KelPzqZTKF
DNYPIccepzJqPCtZK0UJCnwJO4zSnMwvMZtCBmSCgLh6SCCis6RHenfIT6vbxOmu
xM0ikoIcu7hDSsa/6lX/7i3oEHNaHbjjLGhI48K2SOy67YsXklU3GMuTfxK+2FZD
pxo+rX2qrZBm6l2REW9HXcVk6WSu4xF3lkCL9nmznnansgfI3B4tEemmo1O4KbIR
dzCN/yyxJkVEt4xCjABhuIS0pjDY6wbppauXcPLTiIeixjVAGkNqkwI/KKP0as3G
wogYCHqzobhDap7tiQBMUBqKdIn7Jg6VUljdMQffh8Q2z6ma5EzS2/zJzy6mmlU4
4yxP4WQFz8OM4n/3Hz0zt5mFiIRZ6LOzZZFNNt/M/3ItkTIy/Rk+b28DYFFMPlzb
ySfDp4qLCdQRjiCI3sMa1vWTxRgvx+TVADKNZLK4jCmfrmIxFnnhYP7ZWY8Mpd3q
KmerpWXxqb00AOvJdHSTpQ72ZXijg2ywFKuRWJUtYlZ/GQDnAmo/hVxjropyi+UL
+PNefktbLGUogLPLppOOM3qg9oOkssszpyfrLUipE0AbY2Tt8S1URepJ3ZGsEOtD
wWZHWkXItGy0AWjatL6HAizofzbCEhVcDg18OU/HwDYQ89lyZUQxMbv1OCQY+1PG
exlSIVcqwC1YYEyl+KodJK706G9N5ZBHA129zxt+MbUPkTZbaysHBkB4UM/OBZHS
FIL/b70tlVw8NBYRigAeJWDM5DYBS7uoh5qxZtbwCjDxGL4BM4pLqxkbA6e377Ql
zk8pdBykZoG9Qm/JWicCyU4GMtzPGIX8qgw0vIhgJ660dtuLvj4Vajj90dJgxa8y
BQ319TNVs54O+inJSBTYVGUbWsewTP7wObbqCf1XA1rjEj8rJ0HAAJtqNs2WsT3r
Wnzo/TgD7GbckIhm9nBVo3US+Lc465KhxTQGshSOCYRucDJIJJrVszESOdBI8rTQ
B9zcyjbLEheJ+vrO7JiVb8fY5iGTJYdcGMYjR4N+daFKM9+zRv5+rRd3YJTq5Gd/
oFUj9cn66uRMjddCIvilro23raTJQXC8VpGzpBwTea5ztOE19fj9+n3Rv5HOCemR
/0crd2ncCCE8wKibuPSWn656Me4zk6SS+JKhT1cUYGNfma7nA7oxgf8YPR+aaUsn
56DHJdO0AqOQ8n7wJDz6Qe4u6TJ59/JBhbNLJgMfFWRa9wI3Ai09VvXiax/Xm5+v
eA9c3BkPyzZ/+NrokCfcRNau8ydHC7Q4EdYlBCh5+5+rBqpvtXDkVPV47ZC0wix1
8N7TX9GbK5yfU+g7mCZxqkLQuS1YlYcJuQ7WjzCZmlzLrBgjD/Kwf8U7FMX7YaBT
6Bju0p3LUVbyySfFMnEn6hJuxKspFvmWecKXCOHvg9xbMQCkqeXHEbFejcgZmk3a
qSAiVuirPM56JjQBoVu4nUqFSMXHiXSkSZ/tbl/hEtE8UlRy2OkBfGBKECjroe3V
zv32LtTVQ3+aF38mMG7tKcIcMHLJLh5mP0jw8J9Tz5sNDzSq58EIQkIn/4J56zP6
WeCQi8uavkvJRWAU54WG6M8k7iGHRGKLmC1/X66/wxEcqXXCP2MUwwHHYk9vtWez
iMfYb81xjfwRxJMCkKTTduwJS/d0slTTUx7laTIJEzlvxdMgT0MbjCbNRjwbDAiQ
MQBpOGgXwjDwC/z6qARREmxOCs3JUBDxxoSgAd+jOuLbj0EufVp5DL8fDkTUNLiP
cf3QiONkop5hn5v/4qg+L/pvIwMoDz194BK2+RnMKFZbW9xkQZjv0b0ng+08Njln
gjBmGGgvVzoUygdu23wQHS8IRuJDODEuXv3dcEm1OcSBLldgpSeUJDC3eaPKZqye
WqQne+6x/2DHnfFWd2plk6egFvJ5X4hzP07GiYlPWvFlBAMw7QkFKVXSE9eRzHNr
p+N+rovqnB8j8MHWDcfMkmIhxZZmHSjsVIlWcbcNva0tenNxeSuD2puLJrSaP2QR
XAaJmzq+uu0i/b0FELVL6P5LbLL0qZC3mf3HxCDU9srgkQOZycG8Fh0d11kmpDjF
NrLMTacKVRWzCfeqWNlyebMMOla5Mq3PxhC9KNTl8XUjKFcjSG1AbUjuUXXCaBUR
cp3hkPDd8K7reTOIVwpT8m9vlsyg4zXrvhnw0IwBUni/QFzosorwZf6E0188FXil
nCSoseVINhGxG7QHJV2uDDbcoG5/ek528bkmGBWXWsEu485aAFQfaEH6MJmn1VhB
zclEPuNRW7Kw3Diy86/YePdHyTbgFUiUwtjAMVju5ssGgSz+DMVb2CKmQH3vR5L7
4kpKzJIc+kPUnlvJveP1DV8mwTCi7FaHvCHRX67NZEPMWgK+Pu0VAXLlA5lglkSd
Xr/goFCOPhqSzNT+3X56sA/Mc2D2mz8xOZnIWEPggBz+f6G+s7+8dShp9WzAbJh0
kSKdhuGKr6yi3kcXu2vYHA8OFKqI2gFmyO0kY7EXvS/xSiM9kAnX6UWyOSZMXvsN
EG4X5B6/bQFR2g83M59A8NC2d2MDy9zUkoYdOORwToUSgC7hWGYLUsZHIO0Hb9yi
g9KlQLCF63CR8t19VE9d+zz7xzrGKMgxfZdbyIqhnTWMvCl7x71cdVds5T6rh05a
bglQ2sOsiE6xV2Z7lxURLiRdUP8AdplmwWrH+FWnj3/IPdDQ818DRl5kvY4uwvCu
QAGd8AsBClvqSoq3vhZsTY2Ei0SCgXw1h57m7vbPKruLbFZaARghE72/gSxxDrLH
k2HS9ggePB4UKo7uMuRi0TmeonApDcfcHT3u+YmpHYf3rbQffaC0yLsTQuzflE1+
0X0ypYsQT6bmY8c6hDbmp1FDzYORISUeW2mP/ROy/L3fUNxdWKDwa4nweRqaCtyM
FrpF28BC+krdbMOSsVn1PAiuvXUvTmd+T4tsj8hmUQwmsxQX+rEa1kLZFv+YoPNO
5e5uWT4J3zatWgmFm6Fxb66ujKtStHL8Gmg37kKpTt0lfVuYe2/votlfCy18XvzI
JuoCkWZJEo9gl3JqHt2rIIVarr40CyRzuLn1w9vGB5VdCEHtTVglhGX5FEuWp95S
I/QIsk4OcJuVmbrjKZDdTFLpJRo7FAJT8McYPggmpOs+RuHVIRHObrAAPZvA3+oW
K/iZIuabEviQW0q3VV329GP0yo0WreVgixu5rhydcwVyRBJZaypTL/xQsawHmDeK
0KC4zbdvDrnzqz81IGuZVZ6+jDFFSxFRj39Qk3zn6YRBENWK+HUQHSk9oBuqJbJM
2Ng5tqFZyFe/W3EfmnbyhBIkm3xDAqxsd1Mgih450BCHndqya3gtsFFwp/4Fih5M
8WWi4uHtCJjbD2mrnQW5BAi4SumjK22l50k4v1zaqtTcqUkBEKVbcJDJ8DLsUQni
Ezi5tiry7CxLCQTzPagUEtPYFpGDx0dgzCWojhQDzhHw60LL4wOsRroVxsDkmWlW
Xr8TrEkZhV8m9Q0jNvl1+l0dVgx47V+1KWDFfsLCTQgRtBmCenyZlIJFZ174C+hA
Fx/LOBIu9+gnn0YJcfZ89YLCrlwOpouVkw0q8rHU2z7tnlg/NoSPJTdF6V6cJ7Et
4GqA/FsUaD/0o5F0NmYoM/Re/rhn9Z1CpCeIldkvgtUXmxEZsfxr8vr3uZzITUrf
PMWwOJDksQ8FhGnGf1imUlwc4bLMIz2b8CBzLI0om6Jc5a7O0b8Zg8jG3eGef3zh
j+COcE7CkSI/x/yIMxbwAI46nAoAAm7Glk5ARyK7dO+cbs3Tm7TEh/Y0pPDxLW3K
pZPHH3HB0+yrzw03czNhLpJyc3kQtAQbRBAivBgvbSX/3zSc85pJ6nteDEQk7bVw
wa3iCHEUEmWmrJnQk3V3cilFak3zZbVcwwKd5ks7MvGb3buLdEHL/s2zKirISAvD
nCQTCEdQ/gNDpl/+TlXj8xKwD34Mngj3TeY5cENRSTxj71GvOZEbeYpQk+C8bJo4
+ioRwc2obU4AGEuCO1Uxu/i1+rA2nvjGhQzAapPdfh46nqmx7Y2Srij85inWbb9N
9Pd5X1cPGsdCY/r9eqL9dnuDO3I7dhwTLLtQH1u1PT2XEYMvipTZ5mDj8+EZyC2g
Dr9jMNUqYTTXFpmBeNHcvJKdZXn3C3VNZdQ3lijYaRkHJ/oTLuqCK7ypeIDBdCmV
7lXXQRoupVgNrrHWViSaBcgYlONZgIZs3Cx/1lPZcC4rXyaVJwE90x8aRp2hBiCD
fMurEzQKKBPJZu7/4Rc5h3x+Ps0DiwBJ4P+FI9LUsj/Chm2PLdCLapX2R6AYzOcV
xvTGhepg/Kqb5CjGs3Tn2bp27AdIwh0u8f4UeJJBbKF5XbdhbIIAIxrz/HAklIJN
zZUHP2TxgGlAh50Tjfg554OpUZWJXKcJOBJUDyyUbtD9YG9DRrhfUXmV1Gxsw/2J
kOUbdm9YDpKEuS010ztxrf8QgtLow9/+SBZfCVgb3Dha/rhGvZT/+UhCHDuURamI
Y/WYP0ihejWWjDVqWBAGstIDdQt4aY14+81fZ4uswBQQG/7WWu3aVmSRf/9UFcFm
py6XF2Ttu2O7bP8HCgJMh5aHxEluCR1aNrm/qKk6Zxh9EicgHPFxC3cSWZBw13Bv
N0DdrFDb4djfYn3W+VrQtxXklUmAKN2nY1BCJrQzWqftRGKAm3ncdLEpLkZAiOMg
fFhGOVhYjsA6KiT5kFtbJCfXvDrURJuB/m45qT7qsWCJfsOYk09SxStL30MW5GIU
fS+pRQz9rsqYHEl0UVSPLbWxvMBZrToiPMMQ6BlboqYJaMKj1Uyz9WRWKa4X7leO
lqPV7UFfW5jdU9A2smxB6pPZgUlEVsVl8ETJUxxWTtclXUPIQeINI4K3//bN1Xv9
Mv8ejR+y18eue5U/nGerScEv2/vMhqdliVfEOvmLyTGoRalJWBQyV3pp7WSpG6ps
sMVvDsKfakodSpzwFNLNssxhSStVdNskFP882l5zb3SObBpAR4Wx8QWUsXnBP9je
x2ZcGo0Egf1WicTHepDCLVuNK5alfV8U5oiLrM3OatK0Oip9AzF3m1ROxVIrRsZq
cJ5r/Ch0kMP4w/aFoqOpvMSlfybtakcBENflYRzD8MelXJAOBg4vOBU1gBlynTfQ
PnR8VovFBkDTRacvUNbCM5RwOjAHdUI1AHYBAyOxfX52Lq+jCDgy/nFlRPtIu7ro
TIt76nDrpf1051BSdfkfg0MPNBO2gBS1ZYx/hHJxqUGWEGZI7uMsX7/L+seqAxji
W3OaLGMoWrQf+fyuIyldr/mxWfSUPgsDiuxkXIcpD6LsprJgBLxmtseLau/ZAwrK
cDDu1H75CqtwlxIFL98PN1ImFybJRKiUPqDy2c2RSOm763LlnlD2t6ovfzILwlRI
L+zhWTYRsml7VZ/OL5xsXS7lZ2Yo85eKfHfVe0OIfNj6zoFci0C9kEnNCORo+NIT
OnT6FtnXn0fM6M8K6V6COGffLtRKPEyodywBbCHbiXn/U7bXPDsRkwWUf8d/xJZa
CKExtOZNWg2SMCvejQkyJml51tsChATmbqLCl86lWppvOGJeAEZVhdVUN9R0DJp0
ieytIzP9Ei3mKeVoGP6XLvN1v8K/bnzbkkssvoSf+XwUQuYOVpUxe4ReMoLWClF4
S0Hp6GoeiJIcq4JYUEAo0co7Y0f3AZnweispM6KqPPVJuCBlAIFjWwPC0xTRR8ek
gvxnpTQe3jR/gd0W9XOTS7QCTABQVppdAtdRQYd6PMJJLyInDEteyYFEpaI5Iw1V
+N6TBH1AHDG6slxQv8+OkVhVHT9Ip9d0EfHoTg5eTKOSlgqplabDlOIaGQSubFmJ
68ckslSw7e0Q7fG0V2ZVGdBbxSow0HHuVvi9zAWgn0MK/dTZajhveydMSAqxGaBx
CrIRsJruFklDvJzVVHlrpwCa0MjCV+01tWBVdz73eJHuCWIbIofdV/3aoRL0XoI+
/bfudiKinq+DfRUdLJCCYBFQkno6IhxwL20qdCoL6N6WiNk9uwRDv1av3Z+nUFpe
fTH/CJ7IHtChwc51HyVzRKm0+OO/C2XMAnSp9E8nhlpoQqYd9sgoyvI5Sdu26D1A
zPViJSAo7/ZWDSHc2LAKlMtMD3q4xfffMmg5bbHCMrCjD8hcZOxCHtPoXqoQcfBx
hZ9RyKU8renmxIk7Sfs3fd+0uOKnesgrZ4qUyviVd1gdflK6IiggVlghx7NEKlSw
J2Jp/yzw18n5MaofnYWzX2JBTP4wJkFFJf0uNnipTQ+jI0VFfjHFlAFTH/1R1/6b
os4tYCOdcQxO6KjdDfdHzh159SqccjLLTPJZ5ejOEWusAMcBVD8NPiIYIWb9NKIU
ePpoUETxncNeVTLFX1Of+5luvCUND+QHsl9dZZEZXuxmEgGwHmIW5JGEGXZJKj6/
/7DI8YVNIe2cxnFhfE4rm71irT25pgDuyWxLk7GO2BnjkRT2n+YAsuvKv1naQ8IL
F/T/ZdqcV60BqUK2h9zQu2CLgKlXuWFrfPgv8yo+NQzsuKlDcORyhgikZ3Lf5eq4
u5vRlIZOl7I4lXEy+gh1kO79l5JrPpEjNO7WhKbO3ZBGPzKjvWCx3d4id/xWpdYo
sitjSV7NN0fcXafEGNt8f4jvI3A9Z1Us0j33PpHDAzxhFBU87hItUOa9fS3s+puF
/DyMBjmODMvZk0DeMbAbNsyHQffqq0D516NVrPotSV8CMSRodAT5Vg7RS3DOngeM
ZGNQLcEXCeeYVtCLcYPZTFC5XQentokXAkbrcowt26VtSbbILge2CRgSSuXnbRYA
dNbXY15VGD+qvSEv5E92Sxa+P8rbATKhib25QP6fsdDdCQoHR2XXoxPcu8yKfTFk
MrsHwWJwCbaq8jlR3sW6Sj/iXxM8KW1jFnekE16W+/EVxyjKKv2EsIy+Nlsd9nnV
2/dqZle92bQwsSWMql3GCELc/qn5O6LioAKLb4Q6uaZpyJZvZXH+ynuwijaqL2lg
l/WxSH+J2Y1YrUyz9JT/rKUS0mc4V2pD5aOkPd51a64mrX9B7rCho/ZB8HgjdmZ5
lYUlDQz3iHroaR58+LZhay8J1wdx1CKZkhjFZbAQisOZvd/ZpYkfwymScve9cXSo
wQUPsryeqy2XYlfg72GwemuLoZNn4wGZ+5nSqRHPPbaAk8TkbqRWW/ubmfXkdBGw
CwJ1qlHUYuOAo32Jx7S05ZbvNhP4nnWAw1sf6OyeRA2ShTt4/iQm5qoFHw2pryaW
FgK/fadKNjL+iBN0VSw4ssPXaX1vi9D/+BoBPYKYLu66r6g6DPJ2jWYb21qgrqHN
ZGYx8WHQpmNCg6LklNJjc/Fs07yGPU3rROAZ6T3g30532GDHxjeMah6a6CDcfcMr
WbPMLAB+JC8muS/fRlXiyi6LQdix44d5Qm6+Wfjk5eTqicfTMIb8kD1gtGH26NCl
5AullsCrKdFTrMybxfIpH1eu8ZcJGhkoAIPMrtKMiVmPup5qyjtpPyhC6fsJuOoz
gbJOuNsdAqaHwarDiUh74lJLyxf7dcdGZ2mVxhgdD938kl4Z+5xJugSaHn4w++H3
SktIWCYbPHh/CfaX72FU5rWiFqCbX6bq0ay1OdRB0tx9t257Ecr4y6lKUzNuDlXC
5QdYwjjVFMVv1pfiGmnkNIGKVa/I+tN5D/KSCewRpe4pOVoH3+8AlpSTwlsub25s
gmbKnJZYg3d9ERBH1rwPmWOfrw2rRUovGefX3chMaZ+HS26fM4x9fCXh5o5/ZUOc
sYjsw/iZP891ZFbL4eQF1QD6BTaOf99xWYllfKRN2MmeML/A+UyVieN1Je7MLh8I
Dw9AVcNCLmxz/k4FGKOa8qOw2eTFPy2p2LoiE9tUvmSXwuMFsdVZ1N8RCH3wYreR
Ebbrkn+frIEBj5DPvRr9jYAqWpxqgQDkPwuoVPrcaDYdwTc1YalmfixgpJ/Uoj/V
tMhUeQi9oUfzy5hxYwJo5sDKhScUbk0iDdCkdAh+Q/zR95Qmjt+XBlNTpUHjmbjG
FcJysfii9pNZMMYpTidtj9PfUFDY7N7gyXeq66RpMxddqrs/UKJpvn/m0lnJGbVN
L6XXWtBFvcIoXwwiV8Yp6CYitj/ln/FhQ8BpdFHjumWa1g2TroMKby+KxEQWDyhE
013narifFZfa8jR8Le855roO44YWlGnvOc4ZSb3Qo5ui1scu2mn4ivMmu42EgkyW
nsaLsysUB684XE4mFzthZRENp5WyS//weWErv9v3O2DcxBfluECdscDjSPhyN0hV
Xg00yySGmT1vzdmU+JsSAQA8XRpy2bMkQfXQPkBqzuUrcKdxk/5n4BtkU/WuGXFK
QRs2ouMBjtcFaYQJ33emJs6YvW99xRxXpiDU0c6j6rWzazvxJ2q7zEAV89BMBC81
Plrp+lz8DvV7cjfxhTSgflCWhqup+0PfUCJxJnMR9QrVYlMFbZl0+5zWFOgitMyI
rkDAXVVsvi+d7n+eh/kSHE8/Qr5VI/KcXVvJ/mey+AqWcncXGbaET5O6DGfIxsDL
mH898BhIwitMhPU8+/yfUaKN9g5dnueEyZOLkpTHtbnb5nW9sLBnUN5xeIU+N9GO
KUfekEbUV+NUxqh4mhGoO2qpprXa51BrG9kN0MMk5shpsk5huvQjyyXVUDygsNQV
gkOhroaJ1fE3HcED663p9IxS5V8rpQ8Wo4HwXMyi+fIq6M1jedn1vudyz2sArvaS
EfsRp3q/VvMb/QoasqWKZC/VKzf9wO3en9EUQOEysgzJxsyiMgwcoDOgrhL4ONGS
y/1SwvL9N1WPdU3+Cg55SwP93Gdn6bOgUXJYqtp7rmoVNJlJbMgvDZhUF1q1BWFo
gUjAD/q+IlIiZy6/IwwFEocxX5rnAyo7x+DTa76z9KzJ+y+5d03xGHJVCAaYRQ5T
/nmjFdL4oVGD6TUHFAXfLiFWSxn0fI7dxjAlC3trmjimSs8MWN8tuPI6A/+s5dkO
OPgI9fLF5OwBdefB+F3SpHhCmEg2AQ6sKYAWnFvUF6kDdZ9zaOYPHryg9Hp7ATyd
VcI1Y/CvG2s2mA3dlNTKklqWbxwekOoTAQ4GVwVyCcs/TZN+/snDfMcurcIybMc4
scN9XpIQN/ileSRoixZBjJ01fD+ev7GAb7y/rGeAMedYeTr69yAVa0FOviqNl2q+
fqbjBu8MzqnogFWWH0rGuWurNiWjOp1JrQ4+p1O6kAw3DUGXbz89bLc0wstWT39T
kQczEEZN64sEWthYZnn7wM6z2JYL04hL7otMvKtByLFPL4Q8utH5iDuXWvakBqd4
riGt68OxchL/tnk38a40MozSJy/tIGXYaKEOdYVUCb9pRRnJupZhIx8GWe4SyAnr
/2N3noQSCDZDpYAEue97abeYXnRofF+zC6i7ksto3JVkpQ57ZryM9mWvd2799goD
rdHqx8C7JqrYxb+MByNBSttlVdyJY2DDrd7EbmuNLQuoRY+ul/HaMGb/QJtUCiA+
ltNH7v4vH2TfxwPT6h9sr39N0f9vUM4ykDtLsQ3UuyL4lvhvOU5vEADjouvsxeFZ
5Mvjs1u/FEsEsP9qvNY1m9sKMlhjbLzMumGp5kmY5uJi8i2v/WKNCqHEy6n/XLx8
bDOSxO7naqNkvvySk3xegF1MPeFQrmW6gjx7oJpcwMizkImicole7E0+cKVDMzx/
Cm1Bf4vdLXsXlL+vqbR2wdaDN/TXF/frkO17kB02dj1qTDuDQdgGC8k+dBU3xh1D
44EUZm0YIOLrBceJ36EhOKoeYM+tUCYiaSO4rWlX/eZGzOCzj0voH76X2Jdi1xyo
/xjbl112sEXkD0K3SVID822YyLDvqKwQN6zbKY+VgF88YNIU1VUUsVF0PtLh+6R8
AGsKWoS1zS05kClyW34ljhG4XAlp4+Yme90U5Zw7Ltvbc0AEKN7TG+uIqXnvEBu3
SQvmdA+vIbg2bx1wSDWjUVyO7Jl/pEx4PJdnedcyx05hOq1KqWHxepZNRElvFGaV
fU5YWS0Wij3F0mqN5S2UTSkzY3ec5v6pF4jGjZAvVhiIw/yCiLvvVzh3gy/9+7mn
7vIWT+v3iuYzbPinmg6KbOuDx1QA1O6sOg9uow/wCuwHZ3+KpA8zOOU8JRzA+clQ
KoDcwekKMV8yacJS9E3hDCzeWCodqNOfTnCQJaPMAyR2c0P+aNeOWfzP8Xb227ZI
gN6QH062l0dkGBEAFj73UNWNbywUhYRd/KmsddaJPM4dkDmTXtZMVpdNjyPfjiBG
C05mcnRvHl4RkyMdW3PuX+ivft81P4hWpQnwz8S8PXefUHfMmfEnVXZM7IbeDCGQ
9253jgGApIH0ImevltAZw4hUjgkmEfUBBqxauO7PJa+rqBDSBGW6xeTaNAJ8Cxdu
bBosRnJHppP7DG/fFsMdp6QCsotB5Np5cpb2oC0kX9KsL9f/ubc0lPSDeHD10Jbo
C9r/O0hNxmOzPlm6+mBZcc6ldtn8ZmPp09kriyg21lEaq2SfrmwulhCVKe2RcxVL
PB68MqUvm+9UR5lyjInk4yGj86BLk2XHCuPuCF9cIbfGd2+9/51UJOd/hzwuAIMe
IyFn21N4SYIj0CAuYGcosi/fsMaQH92rjPVXapw+Moefi3Vt8zo5E53hTxL0eDqD
kHSRbdsEwm4gTKz+QoLGWFsoIbpfJiglSfjCZp/8+GSDkMOPJly09l2hCVsLzjtw
DN2oNHhvFTGOLszEspJ8ItC5oNO0O8ueqCqgMrVpj9s/B9dCXwa1F0eYlDBVGaLH
IHch8lj0zITkcQOG35GbXjZDRTZQMqDhJmEMCmMijASGdd3cWyc8llY5GOpEKjqs
9+7oHlcBnAJFE9UpNwEw4FbySp2wjYmjp642mX+WPY754SLUejASQWea8sJ3fgV8
jaB5iuxubb3TVr0yjzNE0mFEOQodAwFlERuLfzARQqSHlretk8ONGV8ky3JHNM6h
ihAO++oO/w9xXfmf54OOoCZQ4G1/V/6x6x0UWsEWI2lw/x3tzm7P/c00YCvWwu5v
1cFUDN5tPzZARxqT7XFdhdt8HXO3rq9BWxHN+Pl0oLNDXfDl0bGby5yNfFkB9JPQ
MflNaC8iopsM12kePTXtnrLusQw1karQbzn23Mx/oj9x8+7+sPX1idFvkj81b6/h
tDccmTTz0W9axma4SN5NJ2SBE2Q0TeeQoOhyDfpq9eb4aw9NJ0BzEds3gQi2CLq7
h+UZ9d6NPoHPkO5RDVYXg654xTwQFoRkP4cEZOW89lHckfF9EM5M92Hk7+suvmw0
x8+mNdyqcf4aP1+O++VQa30NM69azfjxv/jBGLglcdUanVX37qCxl8uMNJJUTYj6
y8wU/Lp0d/MvxLGgkKmZQAFYDsEEWBxHbUTqBB6Jw6b3B2+gAqrs8nCl7A1K9GVq
3KtlmDgW0WaUqLRrF1gt8vOz8SLiYCuVoQLroS/9ZF+O00qUq9IMyxXKBmql/pz1
bSnbLNv4epOj6G5IqENl3wykt1WR+gKixJqeptohr94qOmz5+yNFbdd+F8nS1rWv
uTgCk/AX2lZy1kXm3s3AVl/af2AHNd5BIZIuqDpssOql/j4ZRKTs5G9K7xGY0DuS
R6TESq09jCdE518LnZLvXt2P23krWzIgVwLusYIXOvF1lZw80QKs4YQFyXpOaNAm
HOEDmAzbHohQYcA0sIG5pbBV5NBxZHGk3EWy97xVsoj3lQwb598QTasDPe3RPKUm
VnvbtEHMvc2MLZ2xdC30RG3SRNlPXs6nb67H0DcBzCIouBoqZDfqMOImNYftWcdM
pjDBp4PRIoi7FU9kERa7ycRhcUYNC1aofBmG/xoJ1c4wexSxIW1s184NcrQT2ky9
ZPwYS5y9WVxsXahpDjJEGlSmZN4dHilTjqDKawMrqvx7YlC38W3BpPae9gOLMORn
DK2fO37jxkJk0ufrpGz5YEVFG3aQhSl1BOuQrgJCFNpQagziWFw9F1yh1afUg2au
EN6ExadMdt5lOHbh8EirJBVvlbNMDkDk1x6aYrJkxkj3eILx0XmbVmmLUUxL4TtG
MjDcplp7ytuRQdqrCGm9A7xGhRLrq5Fqn7lg6zQgXUzFY2LPkYe2QCOr4yN2u52R
DIR++jheESAKmGKhxmtz0w3TJgtSOSRBMpao6IU5CaflD3zDq/mgfDVrpHJ1met8
hDfFp6gNRAo9CB/s9h1HIF7+UrVsCj/hE/EjwS47xfiMNYc+lZl4Bh3bPNWnigHY
036b9Tp79wuYVC1Rqew4sYQCYxFVL8Znm1A89OPc4nFHLq6vwF1ig1EeeOE2+e0Z
HH3V062rpwLpC9DeXbAcwMKGCHj2qECIaCyYB2oUAM3R7kUSJXSrr+yy729IHyO/
njjdoMCf94hqnKQLLzhWe4Nl7hCO2EAhD7GW6q0HJwJ9kF/RQ6+QRXT+ftTpwYNc
Wh0ZXXqcImyadZrnKnH8VE3rDhu1+YSdtHdfCRC2FUrtKBMRiw4tYzuanybPzWgM
sD1+xAjojriGwG2m89tfbiJ0+8ooGro6GiVwNNoeSgrm+lOSRdge38bQRcYOWtv6
1eAA52+RvTvoJDpHtAasNj911o5b1u7WopSkmwhJdxRZ+PFUGM7mXyckYvW2k+rJ
rEQehWEkS+QcUwi9kZzCaW13lZJCJTJrdd18nuC4SGJgIY97rfUgcJq/XbQd106R
2suTIaJlORYRy4U2ZEd7ht8if9ZPKbwMk+PwEAxP9Fsuj46to2sh1v9Qzh0Lu64o
VaGOg8Q9dO3x1Ryo8nvKcduPyuvFMK2FfDDAuUnpnAGQZrOzQift5usT6ehck9Td
XnPx6WIEZq7jA3fWvWDPEAjbFvMIEvTcXMhz+p+0YR+3OCFJG2bC+xS3shsL2TzG
ALJmy0qvB4vlhUAKPI1m1thZsRwEZOyqIZGOMfPNTC4qGYwNLjg3p1pAhXosMnUc
1vCd97Apiu8FgPISgHfGyA9iuyv+xUMuKzR/WUmx0luYNQ4wlkqxZAoCxWhxR7+B
XVcoOqnF9OEGgjE4z3+KdC+IQPJniHv7kUhDCd+2wVmxOUPagluJ+I2y58o9iqVZ
2spKVOHsFPwzd5Pk2ARoIEJBb0E6pDLZbWsHLLVsuT6tdb89hZ8s94/9jW1kGuRH
Tp13C+fDJyiZq0OnmkfSRllOLOwuLdQtSleU0JtnSVdNDIVgmCmuK7O7WTlCJuC6
RMz0wGBL/pzVetLLCgEdjvSDkHzlfzytux3awISR37nf6onR7Vh1fN05hcLOhVq1
Shzn2eh99l8J3VkOTDQLbKUOn5MKIAdXPyG0iykxy9YBo7WxjnkOYXN9JHuJVKNo
/RVKDgPM+gmvys0KH4vbef/lJ/4qIGuCszAlpFHlEiL7RErn4BStFNwQKXEpxYpF
jDanfM1d0k+1aWStK+Y/1ZHyMZEnWxoPfv8VxYjpC66ZIEMx+NwluNuz/isMafxW
h+z/fcfNsVNnCosUYUsSX1YcCeYao4yDk6jAsSM0WHPTsCFx6Oe01IT0nL/oWkSB
cJLkISxVz73GYahLtx3R2TXAUbkAFc+ZP9BMITaxDZ8RKZNvNREj62zK3bhAqcDP
rg1bcKrPJMVjqO+yJeH5uyG9Wcw/ReVxLYSGPdxoDCufwWndmTCfyioXMu/XIVaW
TOUmpKk5LBSeUKW25NyT/3VKTYI8ldmhO1BmNJ+H0eEnR8Vx0awGMjHSjLT7IH4S
+BWBPTV88jdoqHzcLlRgWSD5y3+S4A9NNn35PJZZRn+mx422r53OLTSltSxbBquL
RV5WJ1zvZK4JDIQvl0t+h099CPGP4PVDsYvQ+nBD+KNfSjM95Ru9Loc0ACRjXIMb
bvko7YdwfturIu0WeMeI4GLYE0qacwQqVdY7L5hSB0XOMRp0Dy1Z0Hmor0hVw+vq
J5PdU9Tuw/+gFYg9QXY+/rST7TTtx/2Ha8SF07JbFa/t/0Xqjqw9GCLFoYwgvIxD
odq27b4kMSsO3igB0+hnfvGaAYS/SG/n5EvhVn10NVPT/LLY02ONkOSK/JvXdUpG
E9e6YEQBdS0Wkl+DKIyBAlp/ILihGyHzK5HVwFnxb6AuzBYVlxXUNELtJ7GnXZzS
sC95orV1PlVRxBQ3bHzU4bmc2b1Sczg6HgqelYX4mkhuOVn9NmCdLr6y3XI5cwUQ
IahP9OkEHPQJl/7DJwkPxoNcgMOT8zKTWb3e46+vtCGxMXaFzEMCGWSMssDQ8/pI
lbmsNCM6HfSbx3JCHJxOPvU1bZURoVMNkl4Qh4aLc2nQHpiFe85D+4ed8D47Ckg0
fz3XGZ7xES9IHBdhVzPEw1MazsHmpBPzauy506H79YVXh528wFjLoyBKHWqgoInh
qSKqsfyT4IjXSvHZwg5fq3N51VEceSbxaEqbV12saRIU2tptaYtkoKfiIyPrQ+Rm
b3h3w1P/6BaESR/koZK4jmWxiFckXIXdFWSrMRa3Z6TQhwlqGJQc5uxJoVvNHn8a
x17+2Q/laCPcX1PbIEVsq+zXEZKgRYlqhw9G9K20/6bCZT7GtSjrlZZfHxmM8xem
jBFEIRSvfUCVAYP41V4/NhiyRrSdIhkHhhTtXmiaIh4BammuwYW3SrQb+7y0QnVv
cas763iySViIvrom8VmdHOgd0Y6C5J2uyUc2FnNBe6J/w2QaTMUrbhGrfYK4Jji6
B1FM8ri8nw5yewzInY1eGiHIQr51pWrGG2x1zGiDD3iZH20Kkyb12jsjewttydyp
WTfAEpz441+/y8f9Oc5uJFgPxDh8hdNnIn43ULdfOCMH7UIaNIdqB8JwxfOn9XQQ
BeCzmTNi8alO8QbawD+5CGd+8dXuWjbGGTKFwVtlWpfsWMK7H3I2OYR8tmSx8BzR
sFvulcOmHxkLBG9vzM2QKLsBw/zkYDth0lCG1sSsPtwXkJB9W2H9y98tiyFaF128
SYxp+LIEfiHnFktNhNSH47Th4aoAnoY+nZVBiNWv99t8aQHRJGOx1c8ixoEtDam0
qSCJ+lkhaPzKG6YrDHfg1cgDb+yxHLyDgGOUpoluukcwhTyPR3mtHDJVet3VvXwn
fJCBCQE8nuhYX0sXvVBtjcGEEOj2jRneGUAqQzFwFo/AFSKmWNEhLEUfwQrQ21pS
pzLzySOZIrC8zWtZ8AL6sBh272djgHPRuu/Vw0MR38KRyGOZeRL7CKUOnDxndHnU
usZih+HnSuAKGwyoVl3QxWKgtXNPqarmqbhg23y/GjhrpC72ZhhzE0KK4n2R0ooJ
n+GxD0I1T4MC37Ck8WcBT3V6SeoLRUFxLkX6fToFvb2LsC+xsgpGE1X8NA5HJr4o
BEX8ZKKGSW39/li+IJ8KUeUzw6jTsHyrCEmQ9VQa3y95JrMpMYoS8c8RVR4IY2ua
RcZo79vesDlvyZLM2q3mK7WSusROE1aIsgDl0oIotyyFMYYz5IO0GgfrimIgVc6y
Tkicck8j70r6flYp+FQG62EPP5ykNW6ITfzhk752wDnCD1TkB8wM59GxbOq9TWNp
meGuXYRPamlqifKqiZdxbU5hjjVWp5P+lsYUVEqoYfn+DajZH8wSCre3dR1W9vCx
j613+C5NVpNqnbyFUtVcSV/MocxVifAWIzsVEm9iZYOuFMxiVPcN2mM+5PIFVUnc
eL8B9+y/8BOuRcHlaqq8/aLfl/tbbZNqfS+t0VClza5QpREHqm16i6+8VcyaWmy0
4RUbDUoFW7Hz3P6RjZRmi54chqSGM168vaQUhMnA4vYPSfUF1K6Cw20X1DdC8rJm
FACQikqK/COUSldD3JoAg6bEeUkT81KFbo8mZ59udpmTA/ocsXneKC5YOwnbInaO
2IK6kwg5p4CJagJuey/AHDYCmp1iOdcYCxUmntepEWpZ90BCKz3FkaqtVRgTJ+c+
zMbdNCGDXDEXAc+xdvZHV3n052i49BUUiOEUjFGjKZpvx1Bvu3rjlLsh06y0+IGF
+S+GTCitX4Uo5pC5LiUXn/0Ho8xLQdW2rNDVEMZiVeAbe4DVgOGjugMEj4lcPgwT
4+ssXqa2ejfL430bPrPxA04DHy3lLE7kG+a+dhME0GH1qfLYMAzlKkZkhAR/cEBv
iotMXMTPmcP+NEiK6lsBIHNDXG0lXonwUwKlax4dOEv9EDIgp1xJNwq9bSTqLj6w
yOI5o2iUOHZTjxmJv6Vxtzn+uixD6f0ZBEsCDXKs8iFPZiqaIVoCDApbn0EweJXf
zD3BpAUmOfUu7tKBoUuZTa+7O4n6kwnaIe+W/CEE6MHHSC9j/y5B6yUNE2NxynMb
hSOyifcRAA4BYzHVt9KUqHWzG5CZM8BcQRtvI2H7/J9JlWTajkHmIDl7BHMXr13V
4j+eNA+FciaaDdxHoLtlmvu6ZXRKmp4kQLcHHvyb/KakZD2RyZEvDuvMorEpbJcF
dm9wiHaBGhb0F/wb9UbPxwzxtRNDlBO2DzSdjuNfBVqN+fPuTJTCeTARzeJl9qL5
7clSVNnS7bypyqInORt5rATTIO5HMZz5IyamKsEDPKpRF+RaDdT3P6tgvbdvek3R
cxEzBgOQWpwHyUM1jA3DzZcVzt45M1PasU7HmT9sz8DdMXPSPyE84slSQAbQ08bH
ahyD+2uP+PotzHlIVrr2IQ5i5cFZ8AqxSfAzOB2uvJIIebqWulCeDnqYeyhSW+fA
to5aUxeDsc8OcSC12+gvi5J6wlpnLXu+oNhiPxjYQ7ydwPDoiZSI3E81EE3wGB0d
fbkqo5O0H2c5Vkvm4cULEvx+sBKPI68X2XxHysrWumYWUbOV4AmdXHJiVaZA/EYQ
PhkogQPERcOcfBw4Us9SrpOxFhcqRmYOg3M/1/lzQVYGtNWA67n6nyKPKGLY4L3/
iSGkow8o9j8PosfT8OFgtpPqbvhUFHOx0Xc5+6CCuRWciIe+W3pOQ8AaF4DJsppc
kRa5tQCTzyoOf/P3kUVMnSeJYHTmGCJfEikl6RtkeVLoMIih34fGOPCfdDodwxbc
l0ZxHNSs5rJ62jMWmZNdM8cTF/+fygY3PxkecCNYQNBO3UssFzYtgpekY1qs55Rv
9Db8EgqJnqJa8+xa1zJoJdu6IvjqRCXzjtLjixeA+vVh62Tewn733eiXMsKgeMLN
hGuf2gt8yE49CDBavFZbso3Wr15O52qeVtkG8a5Q6HA2DMj9NBp2GG1oTkiek7iA
n3EOp6Q0aWr5B+VyTIYyo8MD2Nh+sYTqt4LQ4AOO3+RWogalqV38fshQpY4NuGX2
prfawO/FD+pnJDlRNFvf81YOLL7Frdk5+l/NMnKaoTCxwRcQnxP9z41niW/9GEo/
CRGyBFabZxM/jZe9J6lcRYTAhRn0ZXLnqpBConOmjd1oEcXHPQZjj0X8bNwy/m9E
F80OPzg0fjYwGowCAuXPenW4hvcw5mxqopZna1v/VV9UUopOLmqyuWr95B13uFZM
HL9S3LFzMT6itfXLPDxoIodQDheSl1L+EoxmWx/vmmvmcAACyA/pYgRd5pAPOKm1
ZCwzHHYzIs7B6z6c/5PvzGdOO1NlJnL1NWBxspNDP6EUXrPGDkdW7YxJ8moLLUI+
SM6IwwLFRDtcGBZs0wu4e7fWu7X2Gy4c6M1bwlPz2W3SU4YTjpsuSWUSwpGjCvWX
e1Xt4NHYg+Fj+ao8dVlC2rbUkBatrD9xKjScjTVV4Mmzs2iGzJFMNdVNUuk/YkYu
J79Ic9RG8U1vhAqIDn2NrvixT1HyYSfUEg5bcEEVqbxzRjjuPv3W/cGG9Cno589y
c7fcdEaWPD0HqBslYn97sDEws0kZ3vVl++CRQB8sVDzPw9rRYEr0Plx8sHvrbqyT
JgXO22QtuXNvPmVSGLYDL0/EvZcMX4g2qIFqQenCvJ9va9/ECkHACmCMpeX8IiSY
D938T6Qer7LzjfvNBcTBxc34/wkqaZL6Tm1/R3tjjQObStgkUnO1gDhPffMXw9hG
IvT3h5qbubGmHd4UcZ7Y9JsIyG6q45mkwI3DiXh0mpJ7QWhUukP/6rM/aLJ2UnTc
7U0kcY0jUvP+TypPsWNbIqoD+9uKn0wNgkUMCUYnhe+ih0wNEPALsPhqmfJruEmo
UONKwd6FxFUjebF2CI8OIUB7Dc0cUDDk7q3xUokVOjLiSnPqC57hvRywdZd8/B2S
cS38C0e+uZdWU1I1YO4elTbA4vpTY4ErieFPziFOUIkMng1hppzRZJuOv1wLgtl/
b6B2i2lHpDV6yI5xhRJpcIO5iWjr6C11j9zIv9qC2DvDI1n2NyrjtpkPste+YUA/
oNpLaxGChoK8kgtoqpy5GHVEz4d2cW4VkRr6xbQDAhy8PtNdARH3UC5qHrbsanYd
At6Zq1fdQW9HbJmV59VPWnjjdhca4c6fUzuBXKUiQevL/kOel2J5IWvf0LvzekyL
S2icbDdpQO8ec3u88KQOtijiL91SmUehR3Id/UAbjzwzIY975ZoYB6xx28ZOx+1w
9ATCwjLUzn/LtyFG0mD8W1JsOZkBnkwriORE9Ly1Ytg4OiIQH30F29Cehasc0j/W
wxt2mFtTo4U4VxVGq4ydJhVO2o9fP+NQWoAZ5zCG72ZYPNZowjRu9KJ5ZKPH8BPE
CWNTUxziWzrZETDFHivriddCK/J2LOCpJ4LvWspqy4h9obst7a5xZ1Y1keq/7PdV
yeb4habARLeD7idEr8DWSPV6GTUhfSTp+zpfDk6SwNxpNA6dYCNsjTtHEuxBXTlY
GWnCMbeDKIT2auuxxMtIMMziSiYHCRMAoDcwipguIldVV/KbyLiz04BUaPiadhoK
8FJ6NzxGEkcEOieyFRrG3QxfaEbFYuw11aLjv412Uv5SmOTAcJp94qCrsyB/jRbc
z0Lly2z/eIWZwk1ubMxn0AQ1+TxXbn2V4u5nugrlI67xlZQSQn3D/fMrA+PweHOB
+ch3jAkR92FtycdB70/QDFFjUyKXAqlelYAc/4fUZz5RI0EZIqa5HNHPSj8+jVoB
RWVm8crkG2tzlVvfDB/6i2FrL47Nj/jofRPywmwFEIEMY5wRlR4neYzXmqFVMeb1
F9Sh/ALlNz7PWJoOk3x4uOi/sfRQgztwvHQDM64fkNgIH4I7hjbwABu+iAhZdLcI
1fSGJwepwXadzVCbOplj6gEPq303p2ytDeXAknQCT2nzzo9JA39VbJbsGyyXNfxI
/j613p4yBNfjLeyfP69DJb3AvaIJ3oC/EaHZc6xvk/bUue2PH+9T3IPr+UYIp/6a
sNSLBUkt7gos12QpYrQ9h+URyPV9ntl5CVyQTa42P7uXhNWKRPXXwb2VLvLzqaQf
036snjlSHd+v5gldp44pzyS4lyHpVxTwQYuRGS0wshN9n+eNTq937jB9sFj0qBUV
ZvrKg03W3UxCKbIVJyjSpt3tsQANq5QfnlooYaraDjihBJ4SwPnPXkbKc11h1j5R
8XYw2JuUo5x1lWfF0tDqAZB1JxN2kPfwUdWThLBNFA5U4PFVjgymWFOpQCfTL1WQ
1uq9FBkE23iJZZ2Nyc4Ey6fBuyy9IIKPRa0Nj/LMCNx8GKAWhhr4kKByRLFdI2ns
cl4c6qlsBpgZYhirZQ/55OWQniJJQCUPg/kI0WFN9t78GM2ajE+oIpqbCElgUKLZ
Mwgu+f8QUy4BnKpAODMz00IXj6CcEUi7BA3YiTFa0LlWnuiBDQSJNl9w1zW4v7o+
xFnoUmv0yKKeKo9WkcV7Kp+QpVbqVHDx4cJuyBGygUg/r7ybr1jh5+0MJ8mZlpWi
AV06xRZQ5ZYHwFmF0djBreQXVaFID3T7zTu4cOsEWorwgXZDmbobQu5GccUBaYIL
afAwAdtQDj14hQ4xabca8IddEC1rIXhig5xXoAo9LTuORt5Wj/TY2ZF6WpIIh5s9
CuMqyJZQ1r0M0e44oDHj0kEokyd5Br+BGDpnlw0m+NpfZyA2fR0scSwnyZa7dpF2
AZgs+H1XT+y2zIbej4ZztN5agKZ78lNlvKcYzMPLW6/hlNk/QsJAkUa5kRzxYWNU
VYMsIiiqQFimoClzVnaTvOnvIdPLaWfxHRHEiD98kg36P5vK5j3g9LIfCSfNszYv
WdZ3XO1dV7RGzdrqaEgbQt6c2BV/7hObkFVbLqxuEOWZRQKgEEBW+Rimmee7HFY/
Ms1Fdr7TfMuPCqeL61MbERSdI8zSfCLqKRdv9iqKHdQC0Ulr/mOUHLqwzHSCmAHZ
DxWd27YuHWLVQjdJAhWQ0tBKds2JMy3dxgF0+aQop2VmlLrFC0fWlNsDI3GBfRA0
1w4mfMrESXwzwiuTE00/9KM/4E4VjEoT2WmmXxdLphjx3NrgMhWTYuvQBE82L/hM
QsY04cHAajapmbQ9e5vgDK6UHXhu2+oBqdc2JFp9Rz7BAbrk7dKOBEGwWbCj2qB4
ScTUXF9A+Vr3auK351ehJX2FGWLvANXGSd0xPUuKxByIYlLQxTuOdplEeinDUPnj
SttVa7EJdPPyNYkhx0esthjxwfWNRruS1kfiTGfMTCFitlC9kLL8+BpnZgFPcyRh
M4XHLQREr79/ZiRoqfUuebomCpHZY9CfcZvmnzqS+uFAty+bc6FSGurcacIeqVWZ
0wGdcE8T1ygmbUeSnxFo+7oHHfpZD3aJnjizOjnPBzWydi7Y3zQVOc796OJlShFP
0g5sdFiOVIL1LnLB03qwvS31bRai+SRLvnALC52Y/tU7DrjwhaY0SabTMutryeGb
RolbxCy7nxqVNH3aAgEwZNYpbFt6KthOmqNJEO9hAt4KS1gF5iJC65lGzJHxTx1w
XfgrrPc8LLN8w4a0yDZd/jpMlea0k8GotNcMpMJXHZX0weYF+PKYQ3rXQAT1XvRa
+onerFGgrrF4046KJiS/FEAo0au1cUujUtmNbNFK/g8BJOxJ5tqaWlIOZ4L9WqIF
7jUg089QFhWr9a23x15m1BHVWlXUO92uCdNgwgPNA3kVB50qYraDa6ezcmPC3vvV
kEKRew6Ceag4mb/ghSkvd3l/0jms03jLiRq5Rdlqdi0eR5Ax8YKjgJNCuVzbFfZo
Y1ycxaY9Hqs3Lhe/JWHiSsYN6L19dJWnW025Y68JcEOfJsGosVVl7tgwziOUSgHj
oZPP+qYegucBPiWkzwIctHHJK+HTqGLhPMgeDJ8PfB0xLWP0TUJXvdDle6DcqS3U
jm5kDMP/NQZB/SCECoiZlXFNKMxC1oViirPkbP2v5BwQjumYxkI0vQZEqZt5eeMV
1M+sBAs76SP8VQ/lP1Ttf1kyhUh1/lGpU6Ey9lvdvCJ4M6c2l4zwec6ObwTeTDzU
JYjFfDG/KHVRtZGDa17s3Eeka/WUJEWJajCQzZxDen87JT6yo0SqVzSwl6ZxXDvg
oaeHd4RR+a3uGriYTf2gzNrgBolC7CdaCh6ANQdKqNsDCqM3JOJwp19tVPDmLmbK
e/tSfRQAw1EXrGDcyxixG+oCNFxixHuOygUBrfOyELp6l8eijNnHCpJHuLPcAGIl
i0wBgqw7QEGsHwI7XcynJC3wmsdkzT/okUlrycnw9Le1PqjJh2OGkT6JnRk/x5c9
ekOu6fXWqBz1516uvcjjlBq7pRQCDIyNBSjXIEKLyLWCMPESGUfI08CtEc3PPCXd
e3z+ky7PW6AoQfTAYW4mOKbhvQqrcMT8yF4lwlbMqmICjk1AVpCSqMXtdBOA7+IZ
5WmnXGNYij227v0AWgixpkh3CW9EMXw9z9xvK+9oDoFDVZ2+9/oDjwbz6TEheC/Y
s5QO5a4zb3+HLB/q7MyP3KpKrNIrStD1dP7JNSuM/Jmv8snN2LzLF0yZ7K3YnyBK
oWz0Go1Z54KB/YgzAkP6Zt031/E3saHQhNs/pCRo92ART7nje0ATar4f8U5ecoJB
oLiGjgCgKEUi2sTOrQ4BEVeP18rMEcoWbtosNudGz468FSixksPm33FIFWARx0XX
Qaw1/AbBlNLztakemQOijW58kM7pWiaMNfbAQJT4RNKtlRyrhHftmd5RLodrfXDE
n/M7z3xTjXCaVAPWQOk7cbwajTbTc/9aI8TzyHwg+reim1qTGfcdlMZLfiNzNWCF
vGJCKomxSys/5kAQVYQg6ykylAbMOWMoBPgkcD8HRiaYXRnGAug1Zh/tGKKQALGP
NLnN+5rAfhqybLmFXRgy9MTsMQ9reiV2YvbhjIF68gHE/58DdSyasBUGNFx7JroE
0+oE/HzyiIiuD0/f809D+/FsNgF7RV2DrN6TKmxEFQvRmBoCHJ2YCZGoGsdo6zLp
g4pUCq7zSJnp/XOaFifjXAiPRnEt7ASuv4KwiA/ySmGOi6FMTj9Ss7UpzeboRvMd
0NNLQMNwnTdTwK5IrwfZiIkNAtV27QKr83BHL+8NYz28x0+34V+mcRAABAPU+piN
OxCrit0TRv7ULNoBj4FzVaMtxe0ITtyCYQDH2d33WoQndszljw7qrsuVYjVcGgV0
G2xkp29ZUuWLb1vPIFxa8cFXGNw8AYfnOgvOegWx+95TFk8BsEEThAI2PNjrJgB2
PkC8DbgGbSaZBV1BKZSEFrop7H1n6Pv2Js2NHBIg00l0X72AMIpOtz6ooRQpJAVy
ah8LACm/lsKWJy0KH0S3eyWHHRTh3joLeniV8WYnf+6ZosDscB5zNnLc+vRyNDOM
JCPrKWEgATY0cHh85JLLZqYP0hUCULn13mc9rK3/eTnkmfWHxezEM2WkgX6q0Rsj
g438X1CL4OijxmfhPs8mW5ON30b+UrLrPmwKcAx7WzQ/bXCTp1kc0o2j1EAMf35Y
owa04ySacTR3MiTm7MmSHNaBEVpdZLa+SsYk0dmR3nWiT6zCbiRpFXzHTYivSC/k
ZdeYhLoMr7k9TuXspmtTND2sEqmQZ/+GtnKqnz8Lu0T9osRE3qdoDi62GbpP+eKD
bWxDA4/WTnMKZHQESIQk3Gn4Am8+uoUDTuaHuLxyiGKJktT0PZrk02HCtrnZhE7F
zX4GGlSLfKhONAojGrtNG2r2e55qQdDVZXC1qZEPVl47IsfTkqgPdZXlAs+xrFwq
D6E9LF8+T3Y32zeLv/KQ32V0k9SMi5Rbbs0bFiO2GaaQuDs+ejox61nQxSQB/3Id
hVYAarjrojTycDOaTiSzgDVZrRPgYepmlKSpGv7149LF4rNckHmGBi0gviXkIhO3
nASQ2q34YdvTnGwwWxd0B5xlP4SiZqXmtoQHYLhhrWHwTvemxH54FPp6PV+YW990
N2rLAn4kpJdRi7kT0prVmoOLWGn0D5aKdg+MBFAudFqibj7TpGoGIaoogAGjNgOr
EF+JOP3AlKq/hiKcHge+39q7GJG52EbVV8sP/eH3rFoHjwrigxQ9oc9TpkjcAVFi
JmElz1LxkcdlHeYtDnS27CoSW60uU5cCyj/sSngq8fP7xDMFnxa/JaOIGzbU4VSt
ePzdB9jN8ZpfayAelXwEp0q3gaB0OiznIGDoJBZqBqadgB6OKe/fdH+Du2wl2xgM
g/Et8b0IOzcJ4uwA52LAMpayMgi2KOdN0dbEskas4bDA8raQYTZfeXcmajh/TYsb
EyvuZNe5A/pEgiTGvkPBAklaOT/rfqbQUKzPMKbZB6LfCU8n5fOm5/vzmYwwd082
PsMy8Z0Hmkg+6GHm3KAQWanpjAKHxJnSye9OwlTaueMunHdiIgoGXk7qAXE86Peo
40zI95XCkGM3UmMSQDFkzUmg0unQ4qqN1Qssf/WnD2p7UjXgaArp5FJtFT7bO4pz
Vo1VQao5A+ZykMdRVeahe/Z9oi5PK77iQK2V4gTosP9f5AjWt4hjWbWB+Tg7orE+
zcsIeiSzGVvdLqGES81zCJM/AD1u/LWEZ2jWgiyuacU+j3ueWmhAby20SHAtLlOd
gf1JDxZTYr8SegkwgMV1C0BwvW7zY3ucDgbMqjntE6VxMIYjfxCtI6+jr7jj4F1A
Uf0P+QkkZLf9S2V7Rd5O+kaqgJLISTpk5ZppUiUb7Ob5wPeCbgQXz9gEuTRYN/7C
vHE18hF07AzWpA+VXNjd8mH+Y4xpZxwaTJHSjb/jfqFx7gUG1OvHzd0NGNQ7UKpw
JtcQrgMjMWS/fRpaWTXLLTuzw0x3NO6prK48E97B2FdIXwhls7J0rYqMhuV9dXlB
RSCi8vk7s7IddokQqYA2bxUC5XcfblyBCEWLABLxbZE+XNuVhyEpQ9Z0/9uNxd/Y
LKOCCuUuNA11qVWDB1b6syjdtz38tmzkgYFhG7rSW3PRhABcvMUDW4ZcT0MysU6u
Ffw5myhAj8rxlFRM9WMruu0W5Tcr4NxF+jxW/wozE+6lthnI8HfJ3dyW0xllKeTz
eLRIiBkHmVVTewlthrJPAtiOR64n0W4VmoFY+nKcHIII2doj1PiccnsOv7x9bnKy
c4CxqNrcazEWfHEINrmCarcGISfY00aTSZsFGG0FOV0801xHUlN0AQ1dVhxOUClP
frPu5CjzlmKYo1stmzNsofaZIwm12FD4csoT/u4Pg59GKaA1SntWvilbonsDVt2w
g9+nJcj2ogZBwrU/IjMpgii9S5LElnGnDWTQ9rvQDo1LmQa1FvHx73s+B8EN6YlJ
OUwyvBntdNfkoyurzRwEdVqBWzEtF+V8/1SPCOad3BmOHFq8AWYma6Ua2OzTTk3f
bRmsQAZec1BoDvPFaBRsX7i5mChBHQLrn+JA4jrQBUicapC/2D7O4IOVUNEYnOnk
/HSpXDWeKG9QmrlMvNLRKa0I/fzehNxJAPUpj4akKxyeOAz5LudEHF49A6XtsaHZ
L4VRV+yEueTJJ5oVvzQgilbPAqHtTqOFt1IGcoPYNaLUZ7XQuGbzAVfR+8nOk35G
sXtPAM0V/O+sD7jswG9cg4GveYLoH11cAz+FcC0jIBHgmXN5mtYp0N/o6bTPgZs/
yhB9Vpk6oeQyuHQAZxqsqnF/SRP32q1iNuoLNfdFcFWghzx9nb/TzUHaXK3bp3Q3
xJmIVcHWydvkY0aCIXd9kafqOD9shyD9ergfIPeWLBmdL0BNKTGTIZfgjxpCbZji
DIefX30tOtzw7zdIxmTb2h+ElwDxdoWkbYk02gj6InmbohQ+MKnW+e0PfA4Dj+zR
gTAYpKbLWthHj9bk9NYcFD1HOGkZXTXrLNnxEj/PnJEhH7xZYMHF9v70VZ6e4H6s
B/7+KFVUwf0s/uQClL7tsvrvqKovKo2l/wNCE2rAocjLqe2L7fZnAgEvMtHYNuLp
oXFClNHMAxjEUvgojeZw37qPjSeaKEKt7AUP8wlBAVNVQlBHUKB8p2klAXnI+Fxk
Q/xp7GuuElBLXQZdQHygTAHqJSKuebLaAprdze+W78ACo+bHkIAbIJeahseTGg89
lLantVNBf83sBrBy8fjKi+6yUz57taN4dLABgLjEQxHAkO/cofimE81Rl9GjE4/H
CKGwKp2UleTOyPDGYk8a4+c20XskVvin6ZnP+wTDANQ3lH4Y2c1djCmuLsaMpN5E
UWvhbDk9gsWHF/b1nw4ZhSIwWZ2vobdyEzr+/mva/mxQdqt6Wy+irjclq+LVt/U/
CveCK+A5N7mKljKbri5pm7HX7gpvgW3qdyJ3Gl2F4GKbji1xHEsn8qS1n/hI7d0l
RGiVtpveEW2tAz5WyFqWNYr4ycKsMXQMD6ks6MekdmlXDRNt74lyI/O5Pke4uYeh
fuV41Ow+KhKAyM5w65J5J3pFmEyGNsPSc1thR1bdy/KtvODaQ5QseCxldyg9VXZf
ClzGOaCClGoDZ43fNph63TpTzAGsK7n/fKcUT7PSLHU7WPzQOLqb2N36LKZZqGuE
suQnU2V1A8/PVq6rCNJYSGETGjiYy+EI3xbqcNedKn11stRGncW/FX/9+cBNP/3J
6oSdP7w7UOftzrIGxB0v/dWXoECF+BplxDtPcBvv9FnHOFv50txJbT/ODnqF6QMq
xmQJuZYPVpv1XX0sV1lbowCrHZ0fat+vMyQONNpPZq4tDKKlFIF5Boaa13XXbSFv
zpEHBp1B6TF9jRw2k9j4fUVJERbEhyMiLnRsOCyinNwhOlEJWQn4LAPXYMdvO/CK
inHiIh5HvbH/4ELZorFu5RayYhPmqxvS3VgpKLD6/J1VAHpaYTJ6XRb35oTlF9FM
TU5WQkuxil9KaLPAz6oRBPlYXSaeee5eYGQ3wUC6qC9fAn/d9RfU38NW0C3bQiLX
C+Mrwha9oO3Nv0GgFL/zWNiSrgfQJENKVPVgj+sfk8RYrR6l+Z2IiRKQJF+daSuO
7rAQRoNTQgJjIb0HxGDeDdgAZE9HOMmjyiViaNKBRWbipZcAIEwTtbsyuHO6yMpf
BR4nWyS/XsqnTH2HwBHsVzmONcXOvPkGI5PoPtWnS0PIJGLGRY1x+9ECcITxrebF
T2mXwuQ+XTjOo55oyZfRmQI5Wnyjc6WaSuBgP5lHmP4P3hd4mkTdsV1ZMWXOpVc6
DER4aj3Nrz9C2JNDuWo6sM2bICmHvgv9EkmxLg+X3Cf/WaulB51tLnY3cCtq3jW5
D4UCDLX7DmI/9h5aUIdmWbPcxFLWyHu1PY90k97+r5PnncqYfGLhevISJhZjUmhL
0ey2lPHxBsqu4E1ivXJQn2Osd8sVfaxYs/T94iAJAo3tDZ49z/SncBCuaEQXb5Ku
WPSX3TciE15P7gB7ZM3K/N81g5nE9I7v03nDjVUetEAqvHdY0NLecGdxfDBeQ0VY
MhUfJSXCA6xu9XiE4LNBMhkF63zb0Nzcub5RCInLsAC0y+dB++bnQzlEFjeEZg1+
VM2LkmVAGg3hFK12MJy27pg4IrnXX186saBOeUNoPl7CIe3khyY5aTG8RA3eKLwR
Wm+BrtalSQ7CDIbDTc/7W8AjhGyWPivTPJbpSp6meBTUn1X8F4e2qmKw7gZn2QJ0
W/T3e+o52dDoqMc2l+DUlB7noj0Q2Tw6nPN7uLHHAVKuDZNXRbvtIhEHaL6i/Nhy
LRsdqkRXGjlqJtp80PXJaSWApVbym6D3fESKSXIxxoVT0oCtSbMmTz12KUt1XIfL
rhWoC+Hy4v/ZOp2B3suwguZegKWbGyykH1l/GFjAhHYzxB7EOPLTySIHr1bfq1wj
AdCIXTSmM/xMjuD/KycQK/g++BYvS4BUqsOL6F3j5y/0pE6lC866cLgtefUMRNch
mCVPjvrovIm4LM1UtSrCu7R9b/vymfsJzY9sExIhQxfAL73DnvNr/FiE6nE4k5IO
RBe10RtHwq+q+nkuTo6idD4fE3fQy1t7vcTTlAAhHe7nt52H+q0pg0PNBWEmcANJ
MP31o/Pu3IGSIm0gJFqjiza3vK3uEjBYQnNGiW/4BweGd0aNQ/mGfi4VPp9wV+rD
AlSB9xeMYT7wBhkcqxbGX18ayBb+nbnAOEKylh+16EGNKHmHixYX/1+HW+XJjpBH
qZMiSaFjth/minotYjGHpwqoxbNxIoQoff5s7jvJKzHLi3zNchTogXx+9Ps6B5c9
W9FuUfLzGGdcCaRzmFPrCAodFhH/w+y85N9lXUtA6RIdmYFR0gewmHERUa05OIgb
pIxfWRFICbySBvhEIPmhY95qe9u7plUmphQsgr8TkCreGIJk4++7boatuFNnToUh
qRWNSt5ZWxYvXkuyNhWhnkUfD5C7VWHvYkdPp5/AQP6prTB1Awrwud1iT696vi6t
/5jauaDQdqLaPA1Sqnr0IO+4TRf6ybPYAJCShVRkuZ2KKXX4Ew1rBbEoVc3QcxBb
Jk1SN0XGl3JXy5KFXa7p9kbrhBhgcUARItgUZo+GGV6UBZD7QE5bRNeVByUw9F+L
bja655sy0rOpEVRTpT/mKv4ephya9mroeJxYXDCSUhcNJIn9O0gfECGcLCJG9BJu
jhL8E1Z29YnTnh8flmh2n+U4jLLVJ6JUdq33acdFogABgNibWSvGEGA/h/NQ528p
awUi556hSBuElY+zhPRJm42BW8e6pv8avmV5AffYARs8GmBoj9/vdw9fgENtdr1b
UUGBtKTGoFhUMzmnEaftzLBO39SOWtVBuC/1rpPeDU/ISTzApZYRYns0iMns6J5A
gjuXYUnmAgkVlURdLSSNql6Cie8jAT5heNFLJRuWSmEAq2eEwFwpbQZa0tuJk+j1
ksRg/uBhyTpQ0OF0t0z25sNyWPIe5bAPnaqharVSKa6cU/27U5SbVnsoaf2r9Jw0
hHqFpLg87yLZOWCA07lAitokB9ip63nPF8VK3U3gaMW/R+9c4HDhV92CkUjro7oU
cq0DPexU6RcxBiT1Tyj8mXYvGdvFRVjfwr/WJrwNwvSGpC1NCplF8kNyHvd7jpKd
JFfzuJZzGjnrD9OW1uQ1hlPbMy8ezGLvo0DImImtTTAf9vaUiNoV+iEsdg5pL5Q/
0xoEFmMez0K3RKAQ86+wid78AdbJF5MD496NHXaFmHvTrrG33wJHXK2k+JYIw6hL
3UZnH55YjU5O+UvVYPVea7mir0+05zLumDt8IGZIVudkoMCtKFstlc7K8wEaR9cg
cIvquYeyzVCY6QTfjrmPDlXi3DJABt6MiHac6sZl425EzFJNw2X5fm3hGiq0zH+4
uyz+KvTphhxmmhkQCOX+5C0muHC5kDZ1z0ayflrmv4mnF/1dW+ndQbwjU/IrSCb0
1Ug21lh4hWac0khihV4KJAZ+nGe6Vyn/s7DrGwehmKp/uEwjeACAwwVeDns+jeXM
Txh6V8b8KNYjPxeQWujsPorQ5HQkIVRRYHwXJi5pRTRDs0TgyBdDdGeSvlmMyDqs
xcWjtJXrOJsJywhwsrgJD9zLWEUN/pYh/kvKjY+5H9HycQNKXEVZiXMDvF7P2jJk
6HUtB2meKPP8yH7WFSXXDjqbNLJXHYdGy7hwIOqI7N+JrI0xsmWow9zMQzVEZSou
g7cjNictQkUlUEtp1ap/Xzf8lnCoGY/Ipo9oX7YIQz8kP9PbMa3b77FSzHkhdhC5
0EnpMad9gUQq/M8TzqpEhSQdUd18lPKPJSnwBuYD3QBkaSHzmY+kZrKkkx7M1f5h
DPPz9PyBPBUkK0vyAe1neBsr3IxrIOTfEhDBGkFGztPEHCaBdpzB2dNpgiNrybwR
ffkwDRpntsB+9BQdCEhy89X/eLA9tmrDXtTB+k+pvXpjVRzZ9rN7vBkbCuJ2qL6i
jWjBmS+UXcDSz0Zq86Qx+l3LWA0CLfpQnHyHQrlPlYTBQKa6F0xurtzFTy39p7YX
T0oDEcVHxXEG6EMgS1ahJqlXg+MuLojteoAHeq0QowdBvzAIEh46KwIT/XmwmSVD
lSGgJDkAW3lYAS4e65lbE3xVIpenLbqfG0D7I+1cJqXroZRiAgbPMZSgK6B7tOVh
LQui1JJYjcRd9BM0/0RVrQRkbd00ZWvRKBrxwngje4kjT93EagmeHS6RG0glMX79
2kl61VsvLF3qGK607wamJZwTQnooJS1DBA+NYa6EyvesjxZFf+NWTbYlLr3BNOV2
NOxIt9p5l/VoNSXGhye0zIl2MeD8JIUAqfqZGe1Ik7dwGCv9ItmyrqwIW5hiBr1Z
F3g7eRjnUG5K1bgvpsvUubArrpldtm5a3oLFRzGH/r9N5rTCLHbbSnbUz+eDP5sW
wDZ9EdmHNltAKVHYaaQxGdwtv4QBT80Oir4wq/VcHjafifPBcdZpUE5G2QPa8SSg
pWsY71WS9pvX4dK+tVbQlfxk/+4y6sigC+Z810WvSWwuu4SwfjLYrFVqWmT8aelf
gmi/1ZiBon4eEYYdtMVUptcz6aKW2n6Rs8tZiK2aH0IyL8NdaWaUqxNHolZSF9Eb
/wLNczM6GiC31J+7Qh90Rs2XBop6l4Y/JI2x2n/WFwkmI8/aPeoFmH4fqiHeSC8o
DjI7afEqGpswmeKdcB5SokBJxtxu/18SHD/6esjjYvdO5qS1rkqt6xEdewBOdjGC
yw/ZKKBYrxWmHYd57dtcKgpxzATlcgvnhLE51PVqHD6z2VsxXi87se/oGNAAPt/n
cUvoB4JuzECDEPmvNo7MidnWjiwKqcQt7FSCA+EmU6Yj7jZmxQbp4Hu0dP1f4bJp
kOqbvyR4l56DuvnlHRraNTyxjP1Em3ksEH64NFI71EmbhuTDbRzso4KS8jPaZhs2
A3wKN1teAkdSR52dS6FrUivc7EzslrZ3jo3szvGB9VgMykGvsIrxWgCl3eeXGBP6
jeDlGSippNmbrRVUCKUstpRtYNPq9d46wAudjUrI29SyvqwVIzkN0nqzj5m1IMkC
YrroP6RuSXjWxkSX0akTANaC8bUU5wXGTsP4Vwef4ZyjZZEyMf/Gik1MiW6zywY3
BqcU7A9lwWC3aBw8wklFl2L9nrXKQp0mKagkU7VRwYL3vR3jAVe3aE7wWxwJ6Zeo
0jRdxa5p06Qd4Y8qFV5S1YZghWmfdiLl75WI/xQ5JBi7SygXJ+0O9QUcYDHRux1T
EoG1qYjGW5tX4DF0T+zxJ+a2yUfc0n8ek/rlTU+JlNvC+h6IyZddAHW+lXZlvz5g
xkNBPGY1gD9Dj+DG+D0aJDm/OeX+M9JjC242fuERjHEXwKBOnnKtf85/4ymxS8tb
3dCSaO/n05cjoQEt5amNLs50fskHDNO8Cxko7k1SQestLLO+NB/uryovHZ0lhZ3q
/rU3u89t84XvQ6t6rRw+yO9YNuY/MSkdMz06uy1j7Mt3zECoxgODRl9Ngh/01Tpt
0MYt6L0QOFX72dmvoPIHA/AuxSQMXRXGodSx97jj8vw2H/9RMFqtZ1Nr3rm5i1zj
0PBOvZB7hobeQPpIVVtGrmdbifFsikanZWqsW/fSvv/bl9KKxpxZGfpXQwHuBYvX
f1JE7+oTaKvgONJlP+m9l0n9CykxH1FbcAag6Gy2FjjnpUTlSm+XdbHOumFs6s1w
py8P5MVCGcFOnss0tz8g7O6dIh0/KrJRsl00weoQKJxggQIFJMnn54nbozw/e5vY
0lY6LvKWn9Sggmtc4azvSMHwysxYAnp5kp+rGy+gKULrG2FoFogBbtSUO1D6WXdH
lRCTulD+SJGNtNxxnLQ5N4fOSgHqNPeuhU2gVuqI6mPHTXrrJl/Xljn2pGVq4uEg
OhaJyaKKGpcYRryVuAbEMLlvhR/5qASPNaLGNOb5NcD2xjXCgXUE2m+qUrdDc8UR
n5kQmnXpv7lbXt8BAgF0RPpttK7lve3ngOCK+BFNo24+2wIhJ3RUHQJrkLXWRoD3
cwzzVs8/S29kUPdTqizMq6eaQNcgw1Joa1iNFyWnW4wPri1IBKE1ZFtj17JWNJDZ
8c195jmaHeT0QZbvbLp33eAAhm6tf71vfm9jtMoN0okwlIbJU4DwF3nMroeCvXEa
wR2sBAsgnseMLttN7Sgy2pEZ39NjT1eJQSAa9La8I+7ZBsGGNIQP7xk6Aag+38pm
saSk4wu+9kltQ6jcEX6D6aHMMpdsZo6y3XMYW6RMkoSqC4SJcs+tx0KYL1SkxcfG
nQVlYXSrIFLBwlvdM+Ew4WAS8CjYpPXTm+dee8yj05KvtSRO6GCkAJoMQf2Fbavd
T1u21AFwDdwLzrWhoG6o4M7eHpcA8IWZeVrQsM+nPGMm4lfA0+RugLElaHKeszRy
b2XuL42wNxzQio0XeEHQgu4kzr7aHBmT0qaenJmtH0OFMnbj+ZDEIYTEHa9EXq1u
pr2rM/o/CSrE2tSnvzxmxwZ4FXkRRgWDODboyrAOdQ5xkYjwk7OGxJwt0RFzVGJS
gfMACQ5McbCue+ZcGvokrXFUxLvrqfqbm89UWIvnHol326oHGoPveKgOJSgkRpSJ
GOUfY1l6bthHH6ppLuSKSuf48OQBDtpWcJKKd0ODFX2GUd/LLgaE1pRej0WAtDCO
y6Ax638DJVZA8L64avQGymlXKrR2NEvDicyvxdee+ep+55+5EKSw7kpf5WWm+Xh3
J/cvEYDZbpUUndYdMHXolbFNTgVbpGWUfBkgjnb/FLBi+CzQxhCGVkmrILOQemm9
e56fAyYMH/nnXgFzNP0IkEA5vzbYUGhUNlnUeE28+6RwCqMnt+4aj0QAJQn3g339
b5av6QhTZm8w/6qTdAYkVoonMP/geOHgQEhVUotoyjh0OcuWNFD/8gWXMrT3FujS
5zDXdifq2wWNyp/6or/psW/1j7ol5y5s6FCnKKS+lqrJLWeByZVHiZf7zJOt1DWZ
XCoukztNvGFbAPO/sAbYDGN9cGTTUpvdq/MNhZFBT5TYmrCrLk6MME7tqXzEJ4Yb
z+K/6+FshLKK07Px5au4LxiSDopZHglZWeE+OjMBoLVWQ6mifA42KUANfNIGFyOs
lu7b34oVYGxAkmXx12MdIdrrzxgviQL/UDUdxvNb3LlGYqmMbZPb2Q8H9Jd1SrI/
+BbD+DSCu5IaW4QKVXSs+zrm/w1G0gkZRcW4BXfqRTfrnri1WzKwAaa6gi2hsmc3
ngF5R+M945ugrmVrDSpSnQQEUR1AZEhKTge8u663xIKbhyk2DsvQx5TeUEq8wNNy
uuNPOiDq5deKebaCxjznOfZLBwQmArbMi7LdWj02LQYlFTzjLlCCInMAbhx7uooz
mwgZevvFHa4T/XSnrHH24ZPHDYTc7poroZYEqvIhkreYakJ6S3I6Amm77urTU3NF
zVSTUg4ngSYiLOn3EXc/aorukCnYKBhJSdWAmxEO5mLwzjszikJYHidKWDIv5nw/
va+Mpo90QKNb1k+7ZuEle3T0+f3bZWTzKFl8TMq8qY18ujFo6HVrq9JmANzpIzv8
Yjj+KOaBtfwNrKYDjGv7dH9sttX/3M/z9gPwgb1G1FS8pz9ksJN/M1UOnlmWDOaD
XpTfa2svXVMgsrT6Zu6uwgL4hwLvWLqk5++5UJe8vcluULCONf7sA1Il6I/k+BTd
65Zhxs/rw+0cSbaIP2X0NCRJ04artIsBJ5vbuXXn8az1/0om7I+uQQ9ZB4vgoxiw
GV6he2kVIXt/v4u8/UNrebzXweblnyBioeNbV7OCsP9ekCT2Yu3abIg1wEv60j0c
Ve4vZFHULMX7Pgz2jdNUIgHy/3UYX8Sh5hAkc3dufCj0Ix5dKgPKl40DhSb5sTLm
Iwo2sbs+N+dk66Ftiif4tiUT30vpRDgHZz5TDhk5hwXe8+IVYSyWDicN01bGg7Ry
FwoZBXwj1OcRpmBln19aegq+5Oym89+Tzux9S3pvrNiU+Rpda3hy/7Pr1PbZTQQd
+5DlGCEv4XazUJvmw9znKT6AeNa+ZivB1UFiLKCsLGbAR8+jrMxQCVtC9F8mUhAE
w/iJ4srOynQBCDqxzML0qJagVU2voLqXG2bHHuf80v3BNl+lxkwHtntWnFYcHOWl
+1P2JX7OtEA3rlgBBLSwNk48sMd8C76o8pTeiInOCmeZ+bWejvqH66JXjtZ0X3Wv
icW0XJacAi29ofzOd0kmDVf/Xf1QoFt9Q8NiMuIATIsf3hXeSq4XvPrnvttDEqYD
F2CZNTCj0xx3kPZy0pD88++73rNaSmmX8ef6Wd8QQSuHgCKgG6zOZqcjBTxJyh/J
3/MNe24PmCh2Tv2MNyCbQapmUb7+jauwEGA+52zNqFPKDrz2q2LVXlaGj2OvPoGe
Pg0Np7xmjhibxb1TU+M1OQ9/IO4qEj075NA7LTHzP0b6WDLsCUcflOZppXXKLX+0
zyabaFSLrup+qDaS/qw1oYN2NDazpfrgYnIvKnzt6qHlRuBmZzLn8fOhAjDEDxmz
0IC6WCe6UOYRq9iyT8QsLQR58D7jO+QAwgXCVLBgTZc8oHne9ZRRkn+BRKM1AKoj
fR0A+G77AUEsgbQ/EaumAiawk85LktmD/m7NojQ3jbbfzLhR22T5VO98Xk5Z116S
I7bJmJGk9SRynmE4aqY92eFfSeND6WgG7yu9Fq0KOguHf8j+tx+YWQsCJQq4rG7U
xla+WE9PSlQFEC/F44moqAIftIkfTzPcLltdEnZDzGg+odtMmsSfjYJOgfs+0lcj
3c5qXYrbSC2K6imIhOzbYWXomN7MBw07k9gK8zsl6KpCQ+M13pmi/PDi9Ktia7az
n5ilipuG2PzVJsP0wX5iQlNerJTQ9ULSO5j9DpiuadCh2aYFMrh0sItlDe/Uh/Jf
0IdsTNtPVZpsV9s/aV/EV2bJqaYm9mplblV51vrk8dXocJnC0jYJ26sTa5OHmVht
N4LFffDYvIbU02uTNrhXaNeq5+YY0d/YOpBoMnyAFcPK0iDKodxdKA8yAhoVbVXh
wT8zTzyXIV+1C591bxb/l0IvE/4H7TR5VcOiNhL6Oiia0RH37z+cpn3N0h2YtHj3
/CWJrCv0pwhKIWXhWG2N/rn94Awmth9z7VPil8rcED+NfQfakl6ErIhL+bbcp3YD
Xd4DfyCBPL8jyTgxNSXasAu5LvkjULNT9T/esux0OSS95+HamkT5hoV6DLBEeEsq
IWbmGpyA5PdcrxKsVoYzgjTbJi5IFo5l2XZptzVJwUJgbUzu5QQr4/QMJogkA7db
dQEA82IL1gRREbO2LNW/TRPKV4rPnMZ0wYrvzcEy2jv5VNopAkmtBJNhi5furoz8
CY/sdUdmFmgTdWocoWcag7sDFYp2qW6sRMwVmOBfce0FpQm8914K0gaq4ARBPHQJ
NvO+2ZhdRshHN3Tt70yHpqzjfg3NinuaIl2hDn1FPgtclzIiTTbcLQFrlPMfbVYz
lmwHmF5COq4aNsr7PjEGCby1xpHTSwLcyOdh9UG12RmQl3hVwaHglHBHGkjkUc0k
4S3Wi8Dgeuz4zqzj82CoUUO8oxxlsCZKlaU6Ev0/HHpwUXNmmf4EkZl/VLBzTNJM
b3ddRQz/VBqJd27HoEAJOrkk2cgw0dRjKK40uE5FYieYbmvB3A9LRYSK1vi84HG/
CjwmfWD7smNCGj9w0wSLFFIhPXchK8VcXspBOMcHzlbaYmIBlcIZ4UEe+dHsWNd8
K14KrwOTCBDBLw/oMMQ50tFph4k5RFiXC8qIQEg/qe772FLO2myosHHO11ltWftz
T9nZd3DSCLINZxCXklO2cQB6v0IoiVPl4Vt+q85Z9JlzFawgDndE1aaXMbUFkYhZ
IOE6T5VQN8Uqs0K8pVn4KFltv3RA+wLd9gYapW75zHHHd0H0SluxiBGj/O9ur9Mk
8LVhNo7nWyb0o8Kb2Ue1JnszbevMwReeeBZAEEr/mlfAuSkVbzvR0P9F2OJ6hGFs
PEgPComLBsyyOzf0T+yg58BRyKbaDtg+udhk6hwnUAHi4Ls7wqSkXw0L31dc67fA
ynocVV23on+/fwp3aE3MekTvE7tKAxyPq6HUUdeTyETpfNUL53kIhPciyOCAkuEZ
8j/+rtUWD/QaQTTrvZfD32kRhhv9d9VZ8tnixW2xbuZZoV7tSbJTUHkFjhVw2jj+
Z2uv9K/c99rztS7ZRS/8yXXevNCCpaYjNOXaWO8VH37ccFalPNNIFkJcGBCorgXE
F6gvyZA1NxSNSNzDNmgDVxT6l0Bs3tdizurCGlWPx7z03uzntbcIMPgPIG+FMGty
EGWscMSeCV5cdScRy551szPHazLO4pOfL8LkczcSS0MxeO4rW+uUp1j4XxHcLxel
PsnKIke28JzvlzWYp5X2H/uUJzv94RJbE6YHU3bdt7+4ksBZ3ddsqVKX2bO+sGpV
5UJGd3vHB2CoOzcBqH/PsQde1eUC1huG6Zc6h+Nk2IfggUUSfNhYfjDpgcxGVoQ5
IYm39KyWgM0Js/xlFFLIdd+3xriydObxQ6+C7WRS0zhWQGJVzuEbaIPWxe8j0oni
+2mCTLjYQNR4vXGFwgskyRY2UBU4qkd55zngAn0AjINjWDxxOk7wuU5qna+KB3+h
C0oNjWRYGnsAqutmG4R5fyxTWj3kN5nVTME+aSGtpr/HgSlKCWAiO4rcEP1KK37y
RzzbsDWc5+vbO/nKcnODCrKE/K6uEk3i1ut5QyoU46lYbu5rBANoKOjW8ScOyD1q
rzxuNjV38bx2wcUgt7HXLVAXTSR1LaE3Sm7kfflImAcJ2Fo/jOpxl+q0ZhK9eAAt
kHQf5G0ZPcic2B0DlWJSvJzbeArW+LjxXOlj1H+hCh15ELxtcTmh5oeyX4RQ29b4
edNKQC9GwN0CPu/LV17i/eSnwwOo0Ls5wsSdTZDra/zczyhvsGJ+bpXJJsEwlSEM
4wGoi5y8Tet05gbWiyqNdmcAVI/gZWmvRW5hxETLc3LZB16RAJJYij4w1yWSVBaM
7jgCCHx1uK4aDZTd+iRnt17SsVweDnSJXsjk8dyM/aAZVEKFkpDf2TDstsibJWaC
bRmRY03OpkzFg0NablMOizGtMNUNlkEvkdoBa6n9ywS9kjTN4UFPXU1wBp8bvxJO
q5q8msOHYxPBr2bAKMI0F0WSsPliJRlD+V4wsBO3eDy//2UaH5QEv+33UmewQ3VY
/znuNLDP7CVN5X1hvS438vtDs0YUi/dPglP3w9jEulwclLpY+plHY3472/nlAaVG
QCmwqUuiTxvFI7FsgleByKCSxGDtgV4iJAscpK7/FbNkyfuWpwQQ69HHlUHK0k84
amyJ64PSQy0Dm6EAeKuEBANQCyw0BWISse9Z6jdpAM+s4L15lCkxvQJ+5zH17ewn
6+spW8oxFFufitP2ARJF6Fc1uv/Zb4VuFmVGhlty2wP8C2jotk8kIMql/8gLDrNV
P2gA2yi+/xgS+uG7JJjdZ9F86At1OSp8QnMXgA/RKkXYvpywqKPrsK2mZQCouFtR
B/yY3pIyw8AXlLPStSNygeu0qSirEFh5KeRIMufbxQnjxA03u6fNP8N+/98p0jti
E30J5xI5l6ByHVhlbAfIiUP8Qm3wMdJo9ODlvJfbkIwJaUDlys8N7JpJ+lja+bSo
wc8nwi+W7Ut7YfxeoYnff+7OtFCZPkq6X79KqA0y9/R3nIcxd+nT2eZs+gOwN0yq
3/AMrwPoocX7YfU+gCB5ASpLaOABZXGrLIT8YilYh7R5DKYobpSWO/p/Um0JC3kc
O6gnH4kMUKnR4SOXIl2SOca4cXWKqOEVOXHhFr2A9Nf8YEsAy6h7qZtp4Zs8AyPs
ytv2FZYro2FA8CJrmqJdwx83RdpbXCuKP9++5vxk0sjppS1/FgUE25e05a9k6lEb
5KKmWoIg0/lxB4CMv7oCUmRRf3QJrdGd7Y4CVPXWEkAQVI4ZCySsW3/7mWivTGLI
d9ecu0EneWF7EIiNKrQi+Mo622ADhLgo7TR4S+XFuac+PQZ+X1dx+zYeVs5W6sQP
lP8OvI2DenebwWi/AoqGT3shmHomwQcm2RTJkpOQ6BvsaLr0nzdoW4GCNcU3LOk1
O+yw3Vq4dFkiJ3R8J5PytVYG/bnwsIOBn0zaud6b5TAJdH1QSj0nFPOkYhzyQBUw
Lq8aerFBycTZXknFX/HDStYdNJVPdKZz2xxJ+JN8uQWAb1oH/578Es2v+6bGsNEj
23OuAWcwr3MBTWxj6HYvkiMic0IW6L9a3F0AjBoFwxW1DL6SbNpxQTMrVlXGnCZJ
9xg/MkH1mfpLPrbpF23Im9M9H8NDDJR3C/g5w/qpY4D/5eNIYcrEJklvDSv0Juhi
k2Q4Kq1xXMYvicD4fs95XUQkOP6ae0ZFQ3CaE5zHNvAIfZGSwapn41TIU/IxQlrj
lFUnXyYzUACSFMX4TBBDRsO432+MWfJP342uZBQGLkih+3pxEzcZtbWErp6R/k8t
e/FnpoTXyzHe3YSBwIrqnCCYmNARA7J9RtE0Z3RrF+Iz9q+Qqw8I3y2LsbJYF/BK
I6q1R8Su9/FNYk7nkKirInPtKmQQfs5o6F9FqdjaxKQB13jucRg+rpn957A86ugl
Gm6SNXBru6/vj8DwJ1x1EONc9tlHJrvr/EChCOalAbJ1nL9aPvsowCrKFNRLioEL
Kpn/WXbnSLuBO0chxLmQAFr4lUwRUUpgO5T75nR7iMRFMG1YuLj2DSSvEk5lq+8P
28uaOdT+IUEUH7PLwWSnWOPCz4vmaz4HHCPKIXE1cWAj3vdxKWE9oea40XezcqGX
sMTjUicYiqBzcbRt+BcmZAMAXJGIb835J+aNkDkYKjr/KMYn1yoaQQ+93ko+0gTS
rAU62JtAwUMacl9v5MImZKC0gJBoD4J9wPx76o9P/NCjR+vggZkXlY7HkZTBOyTT
RbbA3N1usdS3IudcP6ZbldOJ3hdCp0iJNvj6e+9XqNUrcNjclUOECax/kgrSrZc6
RLdAupBdAVTmXODIs/HwgTEui3mA3JWCjnqcj/SVzghn3nBlal0XyCOipEXf5f0Z
RctB0XnJya2xF5uB75AN6tlPM9frorHh3FRMBhQVcL7zau9tBGCY8kj/XXFF9l55
z6/ahRP5V2VlNvJw8TNtxoqUKlJs25dPpJ8aaDTsAMBCSv1PtdsFgX2bineCSGJ4
m35DmmnRgJekHOYfVCegVPkGWNkJk08fKACu7AKHO0Nn715iTUs9G8FWOU6MzuMf
Y0/I4NgUojHjtZdgBwL1QiB7nbnJlxfrRetXq5R2loRKW08r8Z7JpQMfaA47mS7p
BFaBVHg441v4TAnZg1k3Mu6qQPsbaEB7bK52Wwlrul86HJwjtOMrt62rdk4B89uu
EqkoylZtZep1BwWbLcQc24h1V3NitW9MJRUq+RE9m40Zvk2G6dTP2xZX2h/4AbqZ
pdmPfGQKZvR04DvgoYu7BKFhwTaPmVEWteqPl9a7CPywV4RsKdqEqOkn8YlbvC0p
a22UAfDdc3BBf7DdSxfkmURn4qEt/p0+bcY3a90ZTniARTuPmfmlzaRzaU/c3VpW
dh/u/ZKR/jiPrtjGErbUo3etPwGrhtRv11Wj5uxSnMJHU9SmARmF2dOS18v/dMCO
oADo6OX+x9uDwZlU7s0TJxswFgQ/Nuc10x2eoUY4hVy+FyzuJI1L3KpBTBd8/Li7
RccJ4oSnm30RIcZtu16AT+ThP4EBoPYbSi+4BMQpqyaRnwVNhXuYCT6M5ThQY6eW
jI43vrWRcHH3JgK8W/ygibih3d6OiBQFuBLyiBz/k7/ZFUpbJ0yO4DlmPP4QqCvM
6awjHCzJLqUvF9TAU6Uk3XEh6y8DK/54SSD63mPl3u1zD+Ym8A7XkEekblpWf2W+
fLjRLtySFczEzS9J/oxz1NDLoanGfi8dAZnHff6NOHdqC99H+p4JQQThkwgwT+OV
0PMzSkihUkXxnLUysQADkjr6OCusEukhIlFQWhB/8vCfGUzLz/rh6wg+dmmRCqa3
V4fwrkd87s6XYD42CzE4l5xjD2ZwVKMpHJa24Afsy+P55dgIEQqCfoDw+jYcfukI
vdGAm7Egr2IYUfe1L2da3HDYNI5NIioZkRiyNbr+4UmME8UZh2WoyGml4YNSdm8d
It4lPnzanWMsj2JTlAEkC3rkiN3E+k0e1+czbnWa227T0BUzx11/lJ4Lo+CNKb3y
hIo5t+NEjde6t2duqqqXFfACrwv/N2RJFaPDH3QLk4ioFwGkWu4zYAVGbGSljoHI
/Q8UTc0RrL1VPFqgz7Dpf0abVZPB54MzxQf3rcdBHNZQfT119V4eFFQsL2nqwTYR
Yg9Peg3cMAuZ4roZqyWnsTzqFvbghC4vhOJeDhSzoL5ey2ryprDWDZp2KgpYxL2I
38OqMXRpJB/RVRx8AS0vqy+ZgcEuJu8D3s0vJ+9abWuxTiK9SrK+PSTazClUGdHE
FNkvU9trM4Fcc1r45MUs91TBopUyFGgTR2ayepo552HF3AHP5IB06N9eAh23fszE
aH1yj2hqDN+1j4/gTJfpty7hxDjOQ9LUuYzIgGA6X+2qCMjR9sh5M1X1oV+nbnxi
qS5Ioj5yYej2o2UV81EuM2ekDSMpEXB2xkvq3sVDNscLQmh52/AJYp5wa0DZ7GtR
4apVj47DsvryGtnGlpeAvEY+1MF48YQQDhQqg7G41bcswqYBIU+/aWH6/3oEMLlM
zHCqVETS5mInYGnQH8175a+oUE54Y9VJuOKC7DIBgg9T3kH75taM4X5NjHrLmdXG
nvC+0s2hFi3rGyw9bIAAbLVsO2/W1jiwYVT38NAH+mQlyLj56m8ae//aLLVyVGQP
hL3j1/79zk0QNW1mZfbFLVp+qHefxu9e6HE3lCpDwuiBQpLFc/vw9ihLGPGB2yES
hGbEFkw8Y6kMKZxdOfIYoJ+bfqeVFc0g3IDsa0zZrrmuWsqa57KTGOdKOQNZCJtf
rYz8xTKs0vC5Oc7UQ78eMx3BVSLsMSnDnltzvMZPxumtXkfWElVsvpj0lAW+miiY
QysQ5yxvaWPsAsAsSagUeQhIzMpU9xfgA6hOJd8h11LvIgRVpxIbXQt9V3ssmR2g
y38cGucnvQgLpGFHWD0ABciHSqu0yz21gscTjkVDR7NeF5gtz/UeBbznZKAqZo4Q
t9KUd6eTp1XRVXZ/Y41WukGnGAx+6fcLKXsXlycQHiU6HOR3n8cQV/REIBNOR+XU
NplGqxRuBzrB8ZBYJBTVvwPHT3Xo8qR1oy6+TV0X3p0zirN39kmdDUEehPkUY4Qc
YoqNJtCbQw5DN32aI33Acu39Pyk3WObO59GvqnoCf0dAdPaUOYkmTlfTDeJ0zDlj
p1JYKScqn3/REjViupdSWbb66622B2miGFBVZ/4AK7oJrAAjkadzaTlLU27RxGBK
/YllIJHyiOS1DDer8jSjW8n9tnEDoR8fTOtADwYtEzNpQwAdyTPBG7+ujtJFKw8p
ZhGM8AyM2QwXed42r6iYLPXzYD7c4u+VPHZu2aK0aApbQeyVEiGZKEnk0oh2MQK1
2iT3m8nq3nkMzoSd1fmnsdNswnpJxr2vOAnFmJW0U7gdOhY6RugOC4Cy4gqOafwO
TxoYVH0AhD+mPPn0CqYrSGUoIr6+VT1b8NcdA9eSxDDZBR/K3jXob640N2etv7XC
y4L7Dljbt0kxMkQl33rOd9Dpu/WS83fZxqWFlNdpltp6L1j6N6ITAx7N31l6dJzn
Y8WHhPkjj+KjAOHuZ6XNyLjtomokBBZXJUtVuvJA/G2arbhemxDu2LOo4tt6vUHM
gkuzsuSRjB6eVz9yUJbJHVZsBVVPyKPvuQKBgFePJcQWqcw1gzFcGE4eGR5GJ3bZ
tuRVAY8M8SUzoShT1jKIIx3FcIAvC8HxfHmOR21rJp/ijY5f6zOI9+vVl88jmmHn
3WXdtVXIHVA8gDMtd/E0TeoTZFJpLIn99fIKZX/Z3rTAlMv5s+XtvtuEW7+j1KZm
XnD2K10HBpW5aGuCxbE2kMRd5tXO72iDRxUyayaslUffjqBRPP3ufm98DJLa0K3n
IX3PlVHenMGWrcnkPWWG2snrJrZsnSFXJMiwyIgYZ8lwYGuk1vouYB3UTrdnfPpr
A0psIdITQgTZZvmI9R481vdLmfJbaFHMa9EX7XJYGfsd43nsnVCC2tKSyM7CchQT
jqpfURCuIM954lv8sWizJCr/kiX9i0dbGYTLWS7uwZtcgbg9R77O6govXzoIWtI0
1yLLlPLFN0EgUzisFxI56JosgGfucwS6KZ5ZUseE4uauJbW/sqPYxAo9wJGgLVqX
JGBWj7CFsmHYAD48DHYknwwAz8ldF9IMMDtSaFbpOCRZTfkMr55XNHzjhn8ZR+nX
jnbZZ4vmRm9OFuDdyRYzlmvf+3k9mz79owRJpNa0qVjeZt4AubaWzJll4J+yM1sl
iFpS/WERI/Sxu1Ztkvsy6rY2gL5Aym/TmMLU3SvsClqvJg8C4JLGEmCiLXsaaV8R
8QJOZ3K48eME4Rj6I8yuc37vu+NxfdNDTDCSLxs1pWl3ODLWfD54kbud5RP4BOZ/
ZgxNmBYCQzmg5SyjyvE6iYCLhaI+rowuJQrs0JEqbzur4+NrM56GJo1gBKK1gjnN
/3feP55T0FDuA87xEfx8bE10zNcoE5qFHsjXtORmR651o1Pfj+OsE7dqDzD+nGN2
AsWEIN1Cjn1DxcDEZl5TNHDB812bgdrwvDhN8WlJyMSD4e7aVsY6WLUCkcm8MtN8
Vpm+4G9NJ6p8DOswDefm87yZc7I6sqgT1WpdCKaPF/ClwaKtl16EVI2kPphbX2Sx
iIu6JguPWlA6zts6VCBd1kKIMfQSRizaeQniwNjMZzAPL+nf7BFFvXzzFiGTsizR
d9xvOsqGxNO3EGD3MnC1X3m2UyEihxOMtrYoNZztaVox7f4iHmYGvwAYoRcpcWSB
W4Ne9yKTh57zuZQSD2/BoEB+h5VYS7rWBLWq/dwM6itCHrJKe4fZICwsF0rpH4aC
VAG6OtXFAwBPPs6ijRLNt21xH5KcM4/P4wI26WSzkNtatrw0ZD2gWgYTccvI9Jtq
NMbvcDEvzDWgwl5uZmC+S557zICz1dAlch+LoN62X2AenjO9ZIoCDEnKGFta3Lt9
mNHQCy8qpyMUE8Otp3pWZAGQHwTVa1akP534FhOVyYxLwPNGTkQcUYFgDtLOV8TA
ab0bUJfjTx9ypv9tyQi5hfioNElgz8dAUt++p2YkJ+tMKxDl3AwRqru335CpQoS0
PQdoyP/OcfnxLwMLtXkTnDNxrGc2KcLsXZLhu6ZgvBa62aMkJR9pzXTJi9nWjtwN
U/JxwPdD3XJTB1qpCdeRBAKvRHp2sVSNh9sb9A7CnvfK79MUEY5yozTBlqTL+0ks
ce9CowqAFKDDJBeTc9bC5EQKHORgpYR/N2BDB2SLWV4LEsiLUAo5B75TQxKhwUZm
QsW6gw+IhiJTu7kBGdaBVNaj4271qDwiGEdz6XHLuHVsgbyXqGL7Cja3P9kP9LHW
5cLGOpQx9pLrr5fVrOAxzYcC3JGH7F0Xf2zWwHDN6D0ni95+BcwW7VJIcyPmaL4V
SfjSVvIGFj8nbxLr28wOcSk2jy7A/tDBhL21g0SpZQmIMFMiaok39KrjWRwyZ/hw
V+gyMyRYt071mckpTTvrH57LFN3GmByg5Dcfh9oXpfxIHTzRuwSnkM4RuIMiHe56
8RC4vdvwwEIMf2GWq8XS6f8LgdsXDwxlQj/Pr2pj0Zq52RL7FTERdS1DxKMntcEo
54BW6ZAUO+g/HVSnninfqlSXP9iZ7LfWBWWJTEivJAicPqe7V8ts8GM3qgs/QZVY
KH5P90gQfWGvmqJXjY6So2gnQa93nP7O0tDcSA68WEsAwfCPB3MkXpydaO6tZVx2
P7zkvzG+9vpZ1K9YkknlTJdTk74w5gaOrZQpw1W1ktiDUh4hvrBdy/wOiqfj9o5y
rAbRbk1GpHHwNuK0CgzwHwtYJvEF9hAYyXs3vWoFIYSOnPW2xElsgp7o1eEfhnfG
1FpkEE68DCc58jcHnuKuASCc9YS8ru5YnTevHh2bAuxR4EaWlQA5EayPWH7RJqub
hhfFZLhN0yaMyPQzaTnClXEVntwGE+nhzC/1haYj5Mmx4ewRcR3LMiiGYNLJqayo
kCm602/kjyG6ywgjQBZr8SqYal8gGVEaqUus+0BmSecLdKVe78kWhmVumGo6Jx00
/Ku+/6WEcsTmfASXO+4OGdCCBbWeZt7/OON2Pnr7lhH26j2p4rpkzlsVS20305wN
FH+rbmrFiFwv0zZkpXxmRlg2WLsZjmlsqSKmp+CB/1czcDR7d0dnHtWdb00e1jLF
tJcLX2XxJAG5aOB8C2WRCZ4gvFHe4vRAPLc3GqwMM+aEkzbUJWRiRX1ySeC1CLap
LwZjvKqa5Ug+IT4EnMfxM1iLXM3P3VTApxtKJ9Ln41ix+CEq93JaHWE+WCoeArgO
F0i2/LxoX3FbHnyOkyPKSJcF07DlC3MGUG8tMH2FAgkKOD4Yg2bNy1aJbWJMR4RO
UrLVcsOkwBcF8ZYv4TnwjThTFehLA4GzYfJYHKRbVeZ7hfYD+3NyKTvwEEjSNnky
nYQfMgRwnhjKu2pfUJqZFQL2i4DjlGUuK4mgGpNuK+ngFEZpuirw9Z+U7DMarJ78
22NVMUh04VOgAIbasgayQdwnzLV7oHX8dgYx5MMViKiCkQjmWyLv1PbS8sMMKsKY
gnV1Ra189leueaoNd9ZAQgTsWNI4o6pMLbNteIeWslAuDreNL85yCcGAao6ozzwV
H9+X92aFioV6D7a1DygO0l7BpT6iYpunUoQDsAJCkKnh4+j2qwOIq6pLMZR1K4lC
As36BtL+AF6l76Rlm7c08XGjDRuRoxV5py3eEoOA0NMXmueQuumAJYCboIXaOqHU
TV/pLsqcbHVgmfJK16s3lGiGudHt6yf+1flnt3wNCP5iw0yudAkSHDLtcm+4JEJi
J/b+j4KIl/qFvtmim87e9Ybd4EJgq3p2VWZG48YIOzhuVRcULsEABu7wGyugAdVe
jubUUfoWsoR9/ud5X7YcdVfA78oLPwewbfi6JCI6sWEWvbs8RqptAH78dU74/FCV
qmVt0xn4osmraYmBtB0jnW6WwuxsoI1e6ocE5kvKKywyri/8eD+iXfQcNDbtYENe
bCyqq3txeNDnKdNRc5Z5SsJOz9xWGW4ecGLLdkKMO7sgKIDCekMkqCXS3CeVZi8V
0h3AzLa2VFxU8aoUNJQOtlcyajGrLAptqPA/nlWgS95H3URsSarkFo1aMKQEk+I9
MhNvAXF3LRyxC4Y2Qh6xJuZplrW24So20VQDPoDyDmioa1CQJV5Vb3d5w9OlGyZh
QVVD09PyQqylKCFnbEbF/gxADCfGG0QW/Ksyumk2omkp9xZYDtxwCamyBqGJcYJa
/9++6ZOGrjnIfAs54yGC+nLUQSPcMfRrKKVp+RQTDzQ1moLLPvvBBob9/bDswdiX
e863OcF4dC8uODzfahlShC928J9UCFA90wY9d7GLrstOVH4FXFK+36MGRrIsvQ1W
5bnH8Gn/Qh2VeNVwwH9EfLsMgnV8IZrSwV5J+G7smrdd2TxosavpLECoPKD71KwO
YXN3yxqAORhXVqTXsAlJMZqYxGCF2VaJFROpqqOtJ7VD3olCxyxoP1YEF5YIXakV
9Y5WO9zuX+z2k81s9ISpQGxZ/dGRy9wnKjxUhVXleOG+wGRpin0c/3NPXnGuoHQV
PACu7dvfatek3B9bgEG4ZxO09fSMc+6Xo+ms4M/e0nPNE4phz0y+KeM4IWjNbeTu
00ymy7Qlmr8tUCoD20iDHEqswpIyz2cU8AB1IcxUzrheq1HKPBWScZEXb3sG5sgQ
2vXPKPd61e3xwdUgVfVbrCs/knEctTHgLFCrg9d7hakvZ5rnFIhqQdonrTCb2BOq
LryMifKzvB6+c/CrddAkjBism1ngDMeQA+1TnI9G6l9s47i6AiaHnOowrewWITX9
TZkc8dVOsETZIssLk+Wam03o8qI1zOY936xAMHwBiroI7yLpbvzQ9bdyHfHZz74S
f8wYlC4XHJhgdje4+9GeIJQq2tk89NpEjKAoiWaz2K1z7sV5JBnQPkWz0AEERBFi
DD7KTkMvDBQu+mi3uVur3uQztHjB2cfbqO1SftTj2LkEENS74JuHYXaPp3oFRJLs
mBTemI5Solq2tq/GI1Zrbi17iD0korNwecSmc0lVNFyCFJzlNTyCPPeaK6ht2pta
kzR19IHYptidieN7TpJ7vDxgj61f1/zdpGgBUxxhYJ95wzk3wxh8kLKEVMHUdQLN
28D/RRoMKYehTzZYhhSs9+lLuix26MCm9otW+srf6hKAiSZK2piE7I53PxIRpWPF
zuyxIao3BUG9ZGIKjN6UKmYSBocipaAEG2Snex3TwtnopoJAx99zeujZ1fYpu/KX
e3rZM4Xj6vo2t3KzyXUsGpYnqNR2aK9k8Xt9W4rcwDvAG5nNhjgEs3qiZL/sU4zY
BIoLNRqtvTMgV2qwRk5v+y9u3wM4R8ccbtNOVGDO+zpBplBoafzGHm5I4mfImF20
qi2jPylz+fosQWW+rkh2fBmrJFrsOOwjRlo+4pGXU/bBTSvpPaumTPKUuiBIxaZv
KMCieOwNZPXp0L8LtZgdgrpEmrl3eQFOR7Cp+HeRSNn3gv2VvZEGYIjZLiH19xyk
ip+LSyA7XzjGEKPwNBrgoAPpGrbBTkJ6eKV8cPf3Jal6VzeYQnVpsqvUxiV3vHMN
ernyqoNXPILWVV9/ILJmHT3wXeKoyi5fetCodcABXPPLxbyY43iizB596GdG6/l+
JouPwrUQjwDZigyOj6/+eNU2w7c9fCbIhGaEYtqKKthJSifWYm/KXCch27z/vIL2
WhmbJhiGD6HCZ5BA+OFhaoRhZDpO4mbYQXafVgECrVDoUrWi+fdzo9hmeafDh5+J
cbklzm15ih+haZBw4rfkMCHBdTsu3gLb+A8bPVHGVTxTfVudBxu/38OoSNKVDKDh
axL5ey/O93Uyk+i0s7hyevuQprmEAAi8dSB0ci++YG6dk6poo0htz+Ofb4yzM9lj
BpTG9qoQKoaio/8dDJxFhaEMTJ/YNZL2M4hLvZUn9xY0XNVShOupeFeSQrLE8u/S
8a/ZbBHJfZiq9DJzRh3SGRTppTtAEHAZQq40zy81IbMBHPOOxGgopDA9lyt+PCcE
2kaVaefMZRTIYZ9CFdmAAlWp38fkTDzOga/1kirD5ZhCgew70jj+HNmREPUxTAor
1srNyzmNCLGbXbuocOQvde3l4zFJPH5kjJleEtwS1Ra61Z7KWBamNJRdpxcZxsYM
wWpkoHqEX+gSA80OcQVap09RdtJ+9N2R2WK5WNSBSuESc9DR33rCRtTUD0IWR6FC
DVSSghVTkKIms6ePqrLtwI8yTYXaJb723IjSaVh+PGCHWpS19mZZfV7Y0tXEfBjV
C8oXWo3s02XguOBVEwsFPCbZzyQduCITRFR/MBAW9gst6n5JIuME8ER9ZN4quAw2
qxK62oWns4DnOBwYjpCXDHmrQZdRftpRlb4f81hrtdieRVHRoXM6t67cDfVHWWin
o3+08B61u4mKNB09xnz20a4dAD0uEPO7hdt4/3/IhO5uwFurNWW5/19ZivB1FSFD
kRa57TJO5/PBv7axoRTsZukmSAM9vr9ZpKGtyS0tbf6kW1S7n38nTPGVX/NYSmpU
WDZZaDsLRoS3wFgpzQSHMiYC4JxjWukWc6gZeQ8Oj2a9DtTV7hynBt4TNeOS75Ef
w4l7ZQiKjadr0rEJF/jFiLoVRoV71pQPssWjlXhOz6s0EYA71muU9NGNbQkUDEqG
M2PvsbOKMKgB2aBuOYaZRwrbvvnGwZ4B63oWIGyIigufO9V6DkVhpzrDfRksC+O0
sNd8tqIkFbWHOZoMcCySjP9DxZKzcYM9P2X/4UQzldgQb3kaeDRssQGzyeIXn4ex
4q1xMyVq5znI47jtfvbVj94JKoWtvfwGCf3rKCKMcMH8GbJ6D/Y+yL/Ia/mwzObZ
ttbK0FFeMbkmwJmaUZwIkESHxdOgr2uOuPiczfeqTm0NwfBdIqk7OwAy1wGsq7bA
XWfxK/ZnlkAB3koQJION9KF84RJMTCXOY/bxwitw5zdotUvJrr8eYUK28bZ4A0Im
ZHhlY9mz93WUQ5vhuQ956ThifIlWvuUpRYbO9DwVHsjv7uJOJ14MRkZ+zfAjsmTE
Rh8za4KAi/LB632xbyKjNBI9Aj+FBybq+kMZM0X3b9ijPjg1u+5EDu3J3aGXz1ip
gYeOCAuzX1E1SvqzoDX/EDGundONPjLm+wjuJJTJDbdzDe2MvokD/2EKbIX4weQh
ijUYthWqzgyZF3Mjo8TJdIlaMXkKkwlAipqHlVs+TczvV9kqFWcnD3CzQ/4X6Nwg
c1gUF8BTO2mkD9IN4gUN0PkOjQ3RQThHmpzt2wM0Fl/qZud/MZdk3xTUHKH6puc5
CbHr+Hs/ASXRXqO6wDAi3Y3hk4QFA/h1vZYvgACC566S8alac46+A/nfMNdEg9JZ
L7X+0ovBaes3PaPrvvv8srwQ5PLlVJOVMNa12ANYxHslWFY44Y1+rAfY/qA/qt4z
dm3j56in+m+0gC3fOew7kFDCVbVsb0i3h6ATpXStiUZcaQ343Lje44J1btqSVwIr
t5o08bsKh6mHyATtLi8wydqKj9PiiW/Zw9CZuX0FiDnasui4mZFG8j/pmqkwK8pb
s2kzG1xzQFnZLp1klY5sGfwC38XVtRj3frcJtddEffULfIFO5D5ApIvd/JpG0nR9
CAVC+oK0wMpkxfy65yRdgL5pnxH45TU+Cf203ecYI/MwbUfe8ZdsR0yNUuX3nsjw
GoPRS5AkljTfU6H0X9fZ7Vy5hFVELVNJSOZ5ryVdh2jN540DMPeJSITEBlNqDEc6
dDT1Bv1e/HUVcs1kXIvhgQMgZ2NrselToTOwlV4gNWLrIoRsosIMDp1oph5Agkt7
DrRST9HG7vS6obpyqnYzaWTeDYuocOfDZ5xOnlIRlLjNTcc0fQFqYP+C/dJE4BLD
+PuPFmIQigk/LIiuY+eSR1SxLYrYfIoPxfdLXBF+aXR3BpLAGjMJH6BEJm4EZ5io
MEE86sz0Rfm4B+mvVUtBVJ10rehOwzpGxv2EzgykkKtf/6vAyPYI38ZziZYFns3v
vcda9twToDa62c9fEY+6qSdEaXHPRimSPc/p3fw6+HWK5W8Lff2gjQbYjaffjjeA
xc1nz4C8YuNrEPOgEtv1AglbpgAEH5U9p0whOC0s+faDR9A5YAqUQ6A0EzkN62Yr
dN1vW6gtgcXDZnaUj+NEi/xHaFLPFajl3RFhrxAagQJ/+pSqFTR4k9w7Q31XpQCd
VfKvG6LQW0hNp648B0VIypOhEsO7kzeR3Wtc/FTOVTgqybv/fQQRwzx++hOMLcWl
75Bf+fAN9VKW+YcCYajB3qwRIDtYormK6+vt8eeRPfJlMom3NNv82qgvarl+Oa52
ZNENKFymqj1uoBa+Ekc39lCNHSAAOHdxtqj071Y4LX17yR8/XWG1Z1Zlw/VcYRr6
vN1LM4ZL/wwx5EHDbWT5M3elMRK3RhLCrIlWjbtcW5ecQj0yDAyQmu3nofrib7fX
Io/5EAxTvhAGsIrCkKQuGkkDbin8crvI9fCMJ+pFRQf1tNr3lU7Lz1Ewql4I+DKz
l9kKR1mDYTwCyMEOBkD+9RhKLMZGQyD87KutGR0HIQcwLHap/TPOBe8V34GzH5ug
XCfSM13vVuqT14KA22DHw8L+MMmFQBqj/+a9fAz2Z1A2LkHexH5wt63ySzzQLTSX
IKgZtK2D31TqDlPUq4mCa6/SEnG3+7UQ254/CI4mzyWHNaWliJc49qr1POUd9PDX
Vn9DIl/eHEqYATVaeooGo4xzp4eRUcpeqSOH4x7Lw06a4IOQMHh41OQNVEuogVCe
Q7gBPMT0SzXVMxF/La1vsfluy2sJRWyqhmLrK4sQlFex+npB+1H/sMtffqI1X5JO
CziWZlkIjIzxusm0U+ONaUjvH/B9GtZdFgxOPDaKOmwI4z92OtJRaLKH10d7XlUy
aYiCTZrb9jCiX7E5li92lIQ5OOKD0zgvbmd3mpRvKbi71Vs6oAmZMWam0vcaWgL5
BuIHoKzNNw6IT74x0Fm7sOBAdju2rcPKGvRxEIqKYOlMSr80mqJEcOo7xbrtEAVJ
WCgPEJL7loijPzafJM+I/Deyyg3ZsdqsUhqmtjvw8FgiK2ea729XPGrrQLcCStG8
yxdYvkijqKZhj4hhjoro9MxQzqQPML8Nhwd6QrXlhYlElCnqvuSo1VPCvlBmiYXN
ObbcJM3q5iLQ8VGffUwwQJCNCLq96jD+mBX4WlLKLiVZRlE2i0oPen1UC0ju/NXJ
CcVyzcxi3kIZU1UY5bL3rRNxOlzQsXKpmadV9NR9+xWdSSiPdAcqq3AtU1i58GWD
vjXZFGQg+Zd413TWkyb1a3rC7zD9no7KJ+QQ9a22AYpg9s/8m3z1HVziQ0G57MP7
FPP86pZc40R1pVR5i7ctr/wjpFS98GJFcZrHo8SXrR9TmHC1tp2D56pcg16VUkiV
OpH08EKlNM4DgGzRgQo+OjgHahFUxRKpOWo2auTGfj4xkmVWyhavjPg2rl89V0jH
4au1WXSGohiTUoh/y0URMv7paUDM5MWy1XOSHIKiTLUj1wuNXbb0waIB3Egkwelx
Jj4M9FwskjUYj/sCUPOMvDECOlFec66eyixv2f6g+g9x4t8iNDHNSTzBveZAK/Ao
eRo/6SIBUjI6KT+QUZWP7nEDYrLN5r87RYntBXzOxe/dLAdX3HnTzQ4pnviajPE6
lVVZtpYCgGzubKNprP8t/BOt1dfu70RiHYdtg2nGPIPsvU1we41aYMdYHS+Ujfwn
KKdKf79X4U24W7V8mDOKaopkVyr3YZQ9aqebUqZuZQHsuiq+plXvrUdSE7tV+3bn
2LQwWfqi0FsLl1Oruo/83Q2d4yxy+/BkcQogyJMJfqemr6O4HdiQ8VxKw3fQLmkc
/DZLYk+mDqRsH8wJIdfmYyvUbK2tbethiRJxNMkJgoS4Fw67mXLNnmxnyyn8zMy/
bDdheA2EK3qSIPOE9T43EUBxuxmABCMWEPRKeFRkagxhUQFBQh3G5KI+ECewfMDL
rXsg7q1N0FOCtQ9pBIHE1dIEp5kax2C5kuNdE2PgX0EUWJ6D2b/xqvTjs9oxojcq
axy1CG8ucmrTasHGWHLaUZ9tUrNnnA3dhscUrtpMcc3j3z5KF+fU7M7pdqkhkfkB
u9i7VIQTrwX5viAHKvi3G2K/pExZr1fFCntoWDvGPziVTBs7Cn2UXspTVnJhpsge
WwF3mbm2vWaB8l8qkJogh+7vHCBaLumnz7WYl+CGTvEZNerE/sELGp7GpK0tzpQi
wUNnM6js768ZQpO3rTsZANCuJOVuE/nL4AkCYyETMGLL3sW7iSd8yVYMX8E0PDqS
yB74RRHg7+GIOMiXF9zPky1BVAsfsbodjhOD/BTf613NjvzGu9xVKYCgpXYp3E/Q
RwuGRCk7vHkN3nypdWAUH4VEIfx9qQo2rNuKZqg6FUFjFHGddckmsM0UIO8nXNgq
jTa+vuIqNi5onYNBgpNOY8gxVGCypMi0emBpMxvfVtNqpheS5mAwx+a2GC52JlpN
H3QKEyjfcv0jx9Sl8NtFmfCnZ982dn2QBm/TnP7OLackmCmSe3pL8FZgfOg0jcsO
BEjtDRDwpdUtc/nPZ1vXB8WCyh4MLTTsUhfBdCh4TaRK9slDtNAn2BW3sI3jEkeu
IyLRx2/7IOxMMbSgNgiroyLrNrvIHgULKEUDhTKIeiH3plZvKpCZvGcjiOQDyfZM
3zaPkrODJUiX2Fn8hCoFku/OK6f9NMIYpjikRO9HfPWamo3uTIHYlmnkn3QzZkXb
0ZzHPTCWhxvRLyFG+zi8nfSsEIiXrPuxs93TehM6dPtz6vVD5FH+24JpNFxPVWYB
7eoVglNQqRQNE6WgCNaS2/+JYYwpRV7JG8426K/6IUksDIXi+cOIMagqWpfnkRSd
Aa3L/fxNoVKebMz70TTtz+4JxpZV8482PLp26kTR19YaOHTdGy6nAy/+3AZMhba+
NENLOiFI2NP7pCkqd/bnyH5dUVHBS1i61LGQ7FIL18L1l5SZMWwaynbHkX1uBdAi
BPkgVpKB4DMI8Uyd9KRHlrKvtNMBNt955tPkDz4qFma3k9vahdjggB6TYjw5QYpK
gUHIq5TF9Sxq+mTlYbJSz1ngchYJAHzPgGNZianJiykMbuMmDLB06cnourl1gOqX
Q6UKb1k6nPAUwhXFTo7NwqQCTbHNbTBL/O5bEm/qfWOTa8tPAaTwh1THZallpSkX
G/cElZ3JEhRfBA2BBYimj4ZS79eupRW8JqnZ5LvLO7dN9aMsyqQ2nNEljP3MRszs
H5eA5cEl3x2I6SYCnF7ZFybccueyCjgsEjHgabQvgQwwtT+pQGoA6XZovV3TNtXX
euNqFrJlPPbepZ6xCH0QYdRF8Ill80lSrYC38CLPtVLEHdBwGV2HGlOnkqqhEFyr
AXUcjvGWqfXsp4o82FjrI/yugFSBTxeasuWWaKdUw7K0OXqM0dAe2P0I811GS+pF
MmDtCMCMdIG9wsLOLVrtH8UVps6JCaJxJctzCyG72X4hUdfLEihmwCK4j68kTXjN
6RM9CjlcX1DSDLUKnwkoKTqiI+3S9FVFArNCavPPl6NieW/VKN51TZoTpaaKOOv0
hbaok27f3EsoGGyOCG+wbui3UlPfQGc+pe6I2EisNAckwBECjWUkKNpEwKgURZ0M
sBRfi8+6vx+bKNhUyBAPBvAh7V5kg+brFKyzC7b9/PgSwmJmHw06NX71WgpSMiFu
/q4dK6geP1U406apl3P/Lhsx2MvxtVry+jKmt+1+IIiIcBqrH3cdhv4J/8aUKgas
uXFixom+Vs0WGiJ1M/S4Kmm/wPlF1YerT+4jvEsSSHH0IkFF37IPojEoowUUsp9d
UaHGa+FAOTgDB01Svw+QUWfVzgOx3CpNMP/HzqqDdQZaLcfclr+6hjcecLjP86Gu
/bUsWDaGtGEW4cK3kSu5RQOANHLSmCmMMdvP4YDkasdVLnQk38K77kfNvuNDC9JT
oGwQni8QfzsOQegCEIyZfPos22eC194VRTGwDb58ZzaEWMTtoWZ8Z4NLLubLOydk
hlND40amhUbIAjxbWqG7amHhysDuNa6nIA6JmNR5jnQhyi6Kvv8IwvhdNcPnHR3g
xsUoqa6N8rq05NZuGVwo9K2v6ZgOdXWTrpKZxA2DDAPDSSE4c0hQMI6VYQgyA0cI
6wV6USo0ikbxv/h2z1Ok6OC1UivjjOXNFwLtELmyA006YYPFX2Y47DKYfjKZDZjc
tbnoDn3Fyg5mBJXXXjOCW5rh7VydZyxOJZln9O7SDwPOKzND9HEpSc5TZWpsE2BZ
eLuVxs3pVQRU0R5FSiX6YU411KvFM+tvyoFArHJ/4mg/Vek9wUOzl/6SmcAW28DX
hS/AuWvfp17MgbLut1Is6x0fCjujle9mtUTrmwl1e2aCFO7W1vrIfGovQIuJfPnp
hFnTkUadNsHBkY4MJx6oSlYg01YcDcolIUKIPgKtR5nwWdavQqYlrxYxhjL+rpDq
ay80J1DT1qPb/K2RBtD+mT7hzExhhIYkvGYXThoKYfJFmYM9/SUwG6F6U9iYI+pJ
6ZWMejxh0IfdXwA4dyXoURF0lC9S+1zFnj0SvMFzHkhzbdgRSAH6zruUt0dpDQDh
ncCy0JByK5mJLzK21mJAWs41FP3JmHPzFZL/Vjoe0C59k1BlyBL3NmHTP0ykbmFN
hvrety13SJklm0C05GAUh1sMnwWrcVs9DdFaXYdBs0YBqPEdX1H+FxyhdPS3Tzco
61kMl4aPj4IFZEzRPdsMCw4tyVz+XQe2SDvLzyzvkYcFUW1K3+9xrnKzZ9nOhD+/
b74yed9JFsYjXE3MXLJcJGIiUZVXfnxTQFBpPI5sPVlCIhLKId3ruDOHtlsMaQKt
pbpnhSGuX7HnO3ySxViZ1z1GVuhR96VUiU27utIVhxCnJWH6Ppi5N9p6l931cRf5
ruxKGePKpw8L2CTNp422wT1iBG8hlXjmObV87ICaiaqCCe9S0DjMiqlD+TWZqbJK
DdeCJS5933WzAnMuI6pVnqM7Y7zm5qDpj4P0/+B9VPmHlTDb8X6O2HWgTRM6byxP
DfQpJEf2QpgZ2HcLP8j2rJjUaEfEuWeSy8UfBWR5x0QKfl9p4UrEYGCHTdnix246
lL80FiC8yNExrLuB1VW+iNZe6IXQO+zoIs+BavD89RK04n9JdyrBTJQqjEemgE5I
hTdEr6PYUUAYGSPQ/BEdW4JqNLOl8uxW+DKxi0P9kdOyLCz4tgq1neKLWQJzf7GH
6K+mpmbTKZVXB7W9+9ygvIbiG2tj0ZISmC09GXajd3c+1M7TankkP5zE23YzjLG2
4VBs/WPOqe9fuqVAvXCvwIL5+yPoh86EJHa/QIg34oA36vAyrf7mxQh5zH7lEF0Z
EBIt3tyb3r32hptwQTyTYtJcolHAAsLP5XnrX/l3o9fzRRKCRQotRfadG2KQsWWb
y1aBxUxJ0NiY4H2HFUt/fCP0YOSiFNJmMmjCNsV43BnpxA6TZdItngBdqG/9Ppul
SEYHnRw98FOzcng7u/eFN0uk2qKt/IWOAEjpkjzIYEFb4/JSmE4JBZAD33gePArj
U8dUljOUCP542M8Ldc1npLVm8jWFq7jC7XIuw+X8FuLvftbhlzLoPwXYdZthBZ20
e959qi9XEugE5nbUnf0PKieKKJZK8X25ktPmtNuhiN3vZLv0dF1Zc+W9qdpGaKSO
kmNdazTtPyEzf2c9VAZg7b4GmR93EshLnAYkv4SSXE2YxhAA1SrpVnuyB6TtCVRE
cLeUlq3+/QAqAQZ2Vtk/dsb2GEhHz3a9OdIpI//Lx5UYSXSUkCfHJPU7RtPxzLk/
pvofREEtC1+ltTP4VAWLlFqeH9cx7EKQO/DqGMx6NBweFSKeJY4SAzBsKVMjo066
98LN0PbhzrGF1qrfnL+UVfMxgTSun5MMhsKpZ0XoHINwBKMB7qbGHW4oelEUggnH
eutnTinXfVypGVajS8U+A7Z34Lid6f1XTddvlhhmN2swA0svO2H2xNbwUMo/Kpxr
6g3tZmQO5aAXQ9Fsb3qlKJ0UJeul7HoSaJ5ClhEZaQ3nLwRfb2gMjCIEEPIn4Etu
Klbds511aSwkX0ht1JTiAwfzLn97HoABGSFq/KLfrC8EofiB/kSlVqhvcnlb0B+d
2VtJJaMszvj7b9ZnQ8u5ZB6kQmYVkjgwqAJNhDQMWFZNl7u/vXdgGvUvDTg8QGiC
kakp4N1qKOW6NujwZEL2Q+gNshsrCJ9mKX6VzzLrHMUuPvlPWzZBDfkGjfTxlrnA
fH/8NxIZlFc9dDHbsS7v/p7ukJSSvTeZkEjbRwHkPjPv3VFB5d0Sd4syO5FTcuo5
VdmoMltd2c2LMgos4ekPwnUGGCBq1TfrUhtAVvMmoV9GkZJZQCAdVxK9+JPzuF43
EzhLnZJl2gtETCyOYM2JdUzEae4LhsN25KJIn7Fg9fl/SlbqQl8lZacKHOmmLJuv
aoDmZyh6vyzGaA5g2Zu0RtYv9/GMPLVbzlkylUnHlLgpYYdvM3+x+iutzqUCYi4o
ScLYDLC9x8CuQueuy3+8AM++hdhaSHcsl8Ue/cqelQqGAFBb1PWSSapMy5c3jED0
S8WoJEtVGbr0V2lF9wyj8BEhf3lJK6rGfRv4Yx96mDz3jhpFkAAW/8RM48+FNDmg
vfxk6uGLXrlAjJZfUiOZiyQF0lTXUbbHhet2ksQRLVRrZ9oMFVXIBQjPNKZ2XQur
VdP0sYbtTkDuqN/r5M0jLaXWuMWWxFM6mgzpSwhiEa6oW4pvNBvvhoaOWrKqWGvE
lxpkgiodYfNc8q6eWlS/6tRSgzCEszlkwQfG4xTVhp45U943FQnvuP6/7d7YFK49
FlwDN7S7RPELTKEnXrJ+YwrqHK8uTI43Dz/f2NuDKWU6lfdrdxRu8OPjym1b9wWb
I9xz8BsO4ivq9DQ77O8fo0O/vhDdy47rve6hgos5Uf81IcmuPS+13bcHC+iWqCr9
SJiPnYSayZR0nOtuqX8XGKB3rUizHovd2yZDUNKbHqQodlL2r84Hn1hh0TOdeqE6
RRpbYDSDjIVdj5KGp3fe4bNHgbJQuxbScuYpi0deMqXBX6IxhjF3WTnYJREiOqeP
DcxRxWnfZAYPGZFQifiOqFl3x7pOj/+C6H2XQflgywmheqBOQa9yC0mzlTOOSE4F
TK8YOqpLwCQyvEjvCsPLPz+99Ckgzs/4QYBv6rEsMrO0RXGZxYqaxtWnyOz9hwF2
KDAlnZ0oUQ+oh8H5lLt/j4SG8Fpi0jSu9r+M3iPvn5dzV5jVpb9M7esXioiAFu1B
uzbNrfmhanqF9jJ/WwICHCOdcxU2F4QnFP+Iq28M1+so5/KgajliO23WXt0epTGR
Ub39rka5RuLIIUqjbkUrJxnthLKi0p9ozVY/oA6iQGpnFLeDpDZnZlwpdZAj/B8X
99pMI9/+7gliBuQ5zlUbtrhvngckzqQFLzT7yr6J2XFT+nGeaufh57GxXfFkdZ6e
rx3VJ0YTfELdwKVyZs6imqKCriLwyACPR4BTZIZwl+6EjHWkIv9X5PXCJsy57+af
wdAjRJTevG3Yvwh7lDTIud1CTIB86NZEc7E9ZwVsgizZwItWTesnR857h9KvwzEd
2U78+g1fgoqaeErnikrQ3bgpUUFkPrLbSWV/1220Zv91y0wVDyIq019GPHUZBkQx
ofrE39cWtzwvtU1wsk4Bsql8F+oXBrCOhjH6ESAS6KOp2GwPBj8/l31trW0PDcXr
dHZ4NU64/uWk/u+nkVHDh8r2v9eGGhiOsfqhH6bAZOe00J32c9Glr8eRGfg+F3TV
JiPlxYh2KNBiwE5nZvJ12wChgNMRtmuvprReymRlckedPV98WvEYlQfE6Da7MJBF
ZJ3yFeXUgdlUAL6Zt5fF6ddvl36fOcEf9IN2M5/RdqEYov8xP+nXu6Kst99Vm2Uc
nuF4DAaXKXlI/FmRVoNQ5zh7c9RNSjLse7CoV3kNmL0YrvhLXm3s/VoIjC0YuRv5
J5jq1ENIadbY6zTT3CxlAlxfIv048lVd00MDEK4FbQJ3v+Yxs6/vk3UF74w/qK/U
ofZNaOzkw8bLwllTimE4Ccv+BsvCqPvWdF0z+NJbwciML+DtuDXA9g28mfRlvHip
RgADbhF5f5h2HmBjRTkHaG+HWCSdr/GvaAmcWfQ2e8eGRV52f9rKoihLDnqAoh7G
TZuVBo1EP/DBJAgddSO8xC9iwcl1dw7k+zujYM6js1ekGXdsqy2ZLP3QrDe8jEXJ
QHULajLYv40rxvUSsRYnMzEdt6IqWJZzRgULh6p0pJsB7CdbU1ipLrKgDCpIC0fI
6BVA2lL6IRYaYtatyY9Ru0eMVN9zi2nTU7Q2HT3F4SbyneAlDu4MPC3AYplJb4GF
fiEmr13fnE8uBGIOBLOIkA7YVqJtejlw/DZfN2Ec5P0YSKEuTTf3UN6/Co4Sf7Ju
ibO4FNst1p43ZuUiwZUqd2JPinfmID+NonKexIcjKImj+ceZSPy7KSltANYN9LjM
WRh5AHz8YnnnrO/vgt4ovvLuJJSnoIeke1XeWn0KpAklc96gFWBuAN+rXhyoSLwn
o5GM83m7Mge/NkdfArzAwk4oTlrhiCO0dYhsGHPQQfz15XxbbHlDJNgAhVlAHRl9
n9aV/QeS5OM+CaFDR0MyYxjC8NQzwiC4M8Pwg997Ql01VxI+SEn2xovNTgyp/oBA
ni+xyXYXRVzzZCLXTf2S5AgfjfdhDef108HUHSNUrAX9DY5i9aVdka+aAlK2RDRQ
cx2xEaiyLz9u0rVj2aCJ3tnFGinHl4htU5fFX1Kbm597UQKkVZDArHdPPcJyc9lu
Cogs5Pj4cDSVjhiyb65CU9fFotB0TXvMdglqs7nRF7OT/jM5sHtHpD4jAY/9QPdJ
/wR/eDF0ajK6GD85qE0UyLb6QcvmACXwc0MKE6Akvs5FFY287aGtL9dvfrJwgiH4
CVZ7t52QDYGrh8kOwDQuSN2x08PLJTf9eyYA2IzqAERAdJdEBQ/ywimzF8phl4O3
7rsoS+cnkkF1Q972Il4OfoY0qiyRz7wbs/kcwOT3fxJqTZj3CLuDrBMIlJSCfKDm
jJmBlvCQsintNSD8VTB0ZRxgEu7likfD9sKnJV6a0yBJFJhEIQWLDSWdpptTm7No
SOF1TQwvf22Kj1cr/tBJsyNuppjdbJ9h7g+cJM7Hr2/ynBpqsxHdjmwl5F0dCkIL
CI6t2JzPvFHKdJ5z68QLnsTDLsw8hlLBq0AGJuzI40rb3AXVG9z51KgQBHZcpoUc
lFH/TFMsmgI4/fiPAFTLyop1S/N/yhH2CdgLAus1xVpVo5a39GZCtpQrAbBfraiK
hNUyNCG4mTrhswNxLDPq9fEYS9EOOIICnSvWsHTahKENtsQsB2YjvqY0MO2AtXJZ
evJVYudOc3RHLBbasl9YLvBFmRx5TZkpHwL0U725gQqWSBJ9kaPCe/Ys6GxXTeOc
b9RX2lujQ9Ze6wH4ztDVAycvw/dVldwyzuwrxbiIkcE3Y1LuOH4xFs2FloNFngo2
SGgbVe5muFMkdTydlSvECo2U3cwjLnG8750K+NPIiJsxa8TWuYwRv0imK75lkbHV
vpWWgidpK1Bpv0J/U0yXgTWSgpoq8wm5GTH83vnZG9Tat4XX9cow9+Oyw22R36yJ
Gm1hRpMr61/OcsUjsyU+ErOI3dm1Y35Qck8ziFXi8TIXrMI/0hWzXd9tULHKzHnO
ERswNXS0A3lXwCE2GbTQ0+dxJLKgUGPclcJNSme6X2mY5nq4w9k99wxDpnJG0PmJ
dRzZY/JkpOEUncWc3cD8he/aZmReUC/1D0q9WsBIGoHu+Qcw+lUfaKfI+GDiP/o0
m92GEB74ICxoezdXc7CGNApTSom+RsrNI9n8o8RaSy6r+GKroxd8g53ajpJJPZM1
O60/wrkqdx8EsgzBOjuZguglgUullBdy2lE4+siKAUypHQyhZ5FG0GlasBKWJlAv
0x3ib4j2PO9rO0kSzWNTX6H1l8dQtXsYZq90f3Y7sGkVX9VT/ObfgvhLIyPa8aUh
RHWKVCx3lpiBlu71eL8tPURscubYvCRq5iZtK7wxWAslqvv/d7Bn7PjCn0G6iscV
abJkrcN1z1P1kfHQSOIdkj79MumfjnpWn5fcGC5uA7G+9uYxRaGWLsS5Luj10yei
wySyCEwmrtXBbe1LMbOhOiXAKCif1U+3qEZi9usnMzsskRnvmhPW9s0zqIxi0rvC
/8f5GQQUOk9+0l+OGMfeBXMiwh4lyFatI9ckMDdyuQJMd3eHrvSLThKdNqpy8dwD
WLzTHXaOoXOJL+8NWtudFydYdNXuARIkWj0T7yWIzk4Hk3ZoGzBjwIiNcyQ0w1Ee
uBqLKWaE/lbFpTbVoB4fUSa2/5k/SpfcGpC85r5xo8cF/DT0ccwMWIAlTK7JwcTU
ESB0YzUihzvV+/EUF1emsAkczZV+KHKcx5kNXnj68x8027YrlXY3L7Xnk2S80TrC
V6+yZxvJCbih4jjgF88wcdtlUAeTFW0vMAcoqvDD1g51o3jJ6DOPAFTvJpxae+uO
ugbQc1jQ45NWMw74SO6UH8+abYCI2t8Kem5J//rUxP80AeU5Xg+W1/gl7lvW7KyW
ueIGYcGCyck3GN72qiWI7l6eHuriMq16/TMJ5mHtANV9KASLJoVHMCft+VAvRgxJ
7xWN/v8X621ncRtXzEJsE1DVfx8hIclQtrd08YBWKhM4ZgkErBwdvR4TJC1GrCBF
YnORBeuUi/pIyATA36Fjg5jkOCUB7AKY1G5fgZw9SwTPVe90mnAdgX6CAeTpkcI2
46kGKRi92pFUO8EaJH9AojNTLet+g6ZAUQHyCrRym16bR8AkCeCWvGl1Vz28axFl
5PtvMKAbeoRdz6RHeoY0rfo1agTu86m9J5kzG+tZbTbB1p4hCxPbUEtyXPPKGElU
xa8eNPnAmUSmj1up8c7FQpkJbwjwUvEyMYhc1EF0BF+iGVXaxx3MyJiPlF3vS67k
6qcxjBZjgyMoWy1WTewVsRIfKWToXwfw6PD4AnufV2oZept6ZXMr5wSfpFDP+O0E
NOpVjJm7iO1rnJAGhm/RdOXeWhVXPHzzOtmlj5ifCST1Rg3SRL/NK/gYlxJkdZJt
2TR0Fb53xgHHb/SoFsjMThNDPF3dIiELe8Du3xXDN7DxeTfMeySdjWaHdqo9RpzD
nyWQYsIFrMEdIAmA2PtwoTJMoAjmG756ktn6LrpOReczaYprRlEFBt5pe2lAmf2O
8eoJ00vE9lEYN+RbD5A1Uv44WuW8/gFxnczjEeaCX5d4bqMVtz2WoRq6qZuyjpRR
+i79pgzQGu0tC+zomcnMqYBaWOtvZno+2Vce7rJ/Y5At7U5OGk6UzuLFfCb+U8dP
TNvKr+ZesY0QOQ/xOzR1RvDVoxuyUGJM2XaSw887ZkWi5NuSZCj/n8Tl8te3/Ka/
5zD3yw+xeTunq1nNVG+KVQEkg5x+I1ahvaNfrzD1vYx9Lwhb8HY0EM48NmxalXNM
Z1Ub1ipRq3ojnZWjOdHukwtS5yKf3WnZcwJJCOe4g+9tkc/8aeTS8sJ4Rcvj1H/M
rheQVwfAjZJm3uHDfK1GHwQ+UiPhpR1E4+XxFeea8z+fLFWd6YWYaRX9/dTiZSNY
k732iFYZZwcpZTkS6Mn9wZgNRABOfJykeKrE9LcVGp6rnGdEUa2O5ocw40q0cAit
xD06Ft7OfBD35O96Zdanf3E9yux5IWCfQao4NbozIPmgUvS2lDw4FepRTOQUdZae
CKdxJwYvs4plXRkQWxhVFCh9YtWhWmTk3/Z1ZRIP/4v/A+RT3YGIELVYlaTNAayK
cfEXIZEiEJPHcYfTSHYOtXegRMqn9tKoS1CXLfMkndbIVHar0tWR4rsyg9ImHvze
BrSim6BbWNxRQCDRmY8xB0qDCWCMrr363sOi7JWknoQ8LLu8QIb87F1c3yqTY0Fd
ITQ/dD6H9Vrj/sPQ4y1S4bdlDjMutvpuTDdcHMclHo+UNChzH5Wl4lXBple0HsEQ
BnW4hWVXYICUqjo2neKIgFIol+cWj80bdluSAmXipqEgcjKhuRmSb9senVryMaI8
7jDX70XJEO0zxQGAURtoGCilMK3sXC+KznkxNAb4eKVd9bcnL8AO4wwi9oUjS0J0
GZQPhLOUL/H3+2TFc8AG3o4tJWFeq6RmSEY1OjRzhJV2OOvHnJvHSMADhRGTmBZp
Zm88Up8rxcUmfVXS+995S5wv4kP5ZzLubVm/7v5iHUXebpJ4GgKjsxHdAnPSoBkE
3k2f5BEK8Uusi0qT95T9Zp0FrN5EaAMmeSQmrBJDDoNvrW9R9b4Acyh6KYq0X9Nm
Fgc1t8/hOCi+aPbTXLD5g4mbBvGWtdK2qIxvbjCAFmiQaGtFlzD64ep00AOBRgxo
HhJo0v9xy8a1mEDn+5Gv+fjTase9bnPy51n+7ul6miGHSI77BZZzIi9H1Ol/VTU0
v+fkDM0hntyL//XIGcpbP5yRnfIBGtDzbLAYe3bkk2S20I3AXxx1IsspyPnXu+Rm
NwGE5yFOGYM2cZSNs9BwSDj1HresELMINfSWh4HQHC1mYR+dtdP8cuuzmvoEd7Pj
fGNOqp/pAna+pu4DqGmnKgRWEy/+Fvm+FNplfFP7qH2qJOeRLjHUtu3//JkEioFE
dGsOEQnjPi2EmTjcdUHy2D4xtf/Wo1bXZ/J8JJfBqbh8RTSAxg+5lrOum+PlNZ+e
c6w96pUctZ8NQnN7TptIjF4KlAvBDHB1gsJYYZLxKwITyIhxiJyKyEaZLBi68DoB
P9eRpFvrbNSfu3z/C+f4Hbc8uDkfWd+mIs8NUdd9Dquvtb8g9S/hN+8thnU9Hrgz
NixNzrC7RLHx4mcE7UlRl40PvtA5ToiNuDtLq7RXrppuN1qi6vLY4OouywmiK+/R
5QEy3H9mNyopFjqJoUPD3MNXGyMnoiyYVepyxMfGPzEPhGq4Oz617vGNcUWsBvna
3L6XFyZA/SfdnOX3XJyTEwjuiGDppt6/46AQhh29ErmW7mvNyjRd5eRYxwqCu2yj
0JDVbkrsgidjFF2sclRZBcm85TdFkUPRns71RhPmhp9/gDYrb6Y3lKhjjvbK/oPb
8s7ZYYPGHOFcnXCWtbagB8OQuaBDfSPYKKl21wKvrRND+fJF9x/rMnZEa86aL9du
d49iAYW1JAbL0PfdPnfQ0bq7mrigjY9RcY0YjvCAIFvV4Es4FgOUhxHDdzY0ZbUU
k+Zi+rqze1CwWYd8/tAvriHhOw+6miLUr2WRQB+kfpFmUOs80AgfJ5DSwfqrMfvN
oHWjCCFu4Mgcn6y7SLwWzsgNoAELABAbq+U829m+wH6v5AbDAaRn7x6fJk+fHksE
NklG8pohNStTXhA+IrBGOhZedWLwJiat8BIdSB5v/oWe1KSbBKCq8Exn3lFehzMa
Fe66H1JdWEntY36rqUFZMkbIEqQV+ziWKr/RAu/IgJheHzQm+ug7rhlJQM5YmkTn
e/OVpyuSyW8GMRIB2jPvKOXBnQW26W7/1LcN2/L72Oty63qQI/n4WdwG5QAeF0WD
m5Q8R9J3an+w8pDgYFmD+r6GAsCYHGhad4Ue/YuK39e0qBb8v7E53YaKo9inNDVH
GUKZgT+j6sw/EGCL0ltt25O1gqj5fpzfw5+ZeX3ykeU+t+1dUjpXL6KyGgLKT0Xg
5cM5+Cv7Epiw7fv3u0SwHxw2zM7TKTVVgivUTFTAR3tCkmk4ct2HVYgpV9O8fzv3
wOY1x3eF87lsrCumfEBF+AKkrqwxv3TU4720PSI20UgzFv/w4O5P9x/+9LkinMdN
NwrooEp5cJjvXxapi9msneFzGLNSTcfdEYsuteAkANh7/xn95V8VdGWX05w2nSRE
9rCducXrWQvX9REg4GDOGxBYTqGqMZiE9fmZjTOj1wfnqwAUuoNosXEmiQMcij8C
lE/9+4AHb/nJLMsz/pcnEuQ0uJWwE7clDOjEGZVZjb84VtAPjqnKoxhdkiwy1ALb
Retcv+LZ2VDOGie5pGzTa5ZCHpFYIZP7m3Tan2szOjltbsroqr2rhCiTwFhG0OjA
IM8bxFXTmQHTxbldaFk6Juj3Z3SWU5uhoTEnfWMeUI2yFremMuLOp+aS4En4qbsx
23vGOIC/p913RFAVzZ0zggFq4N91IV66g5r4uKdufZL5HCPN1jWgBhmGhFfnfGJA
OKIrcglQ1ietmLP2sKXaBfTlrhai+mmDSUu73pd1fvXEjqjtbyKiz4H+SwUGmYKz
F/BQp4/MoYSnLqkD+WYtp176NxyaNqs+kgrCsaS3WbC3XNt59Hlyq034c3nF2ZoS
SWNuWrPr0S60KdU0vuHggyIrhdQeBuciYDWGTmRxD+wgVrxu0Z0lSbXkPD6a8ram
tLgfdwMR+l7gOd4w9LU+KbAIKliI8kNsleXw/l1g9zgiNNMGHG/7Kh2HMy/EZj6L
W0QRU7NAFCmwU2iYHkHnZKfw4oAaQeUe0AGoqwk6NcwzmXWtZ5D01XMqnq7v373D
RuJLN9doU0gPQ2qMn8ovyXAqkhXgaMBwFiO0+rPcoJ7LAS/wKBZwhjDADIQQ1J6Z
kC8DEsPo9qSL52lV2h9u2fLNDzE7Ee6F+E5WofO+DempiweGkBxVxdbcQAvRUMen
QZXfICQ8LoV8GIBiKFiklzOrPRKBOgXvfKYScaQPyUsDZok+knEE4vHXfDJEFKO8
FNPfvGI5F/6Mjf6jA1powJXJ9zmbBZtDL9wTu4CNAfvDtz9hhSH292bCY1otAWqH
CxeKca2n335J4mdldHe9ntGMeQWt5ACCNIkJ+FOminXn26Ixzbg5y80tVvvM5PEw
wvqkmscEI8ipibUOf+NUCjCxtWINJOX2Sw9g+nqGkDKetKMjG2xGyU6cGYY1Z/4l
fe6gYUjt8plnAZUlg3digxcTX5HaVSfXFCsR5x+ltVI6+RD31lr2YETBdCUhofhM
F5xuoYmk1PYJDeGh5mL2gPaQz6zXTFvF7A+zQJIokuVBamrmK6kIs91sTLjBTfAa
V1uLO7R/O8Jgy/ELQ5f0osuXan4xMZ6P+Aok6WBciXCVK1dcrbkTw2aJQzM88UID
tyzPqLWosKW9jIPAAE4BaO5d2djKsmIt9ki5+XSfbL1ZCZUuKzIqmFrzkRkrDXfD
5uPUP0ZXWKqKa3i5cmqLRo7up/QVjW+qrqZH/7pLqF9q7TsIjAK/G3LPLTBBFpSk
U4ZWyeu78CUo2/pZOsJPIZ3AI6G6GV5OwiX+NC7MAE0E5rgOX3EH/K1gPQGfA27n
bJTKABbs1QWGm7GwbBoa3Lo7q8PGadc6QCuSSiIXPp4LFPv62W3O/l3GmNshFjAA
tEK1esKvHcLk9tx6JF0fTM4YZ5PLUmczhyV1knnkggoayCdiIBeXpWrCWG+1aARL
tZImPO1kfDJ4iAUA2Ae22xUse3v0sYLKrBkSXPvX7UGh+ngE63kMdUryGpT9nlXI
oH94EYVKG1F4BatdcyWHHdIxjpFOx6K0rUPU21SYXfvy0Ty/SQD/QOEQdBHLyxKS
URZp9yVWJ3kl4Dd+g9hyF5iZs1KXEzG5TzbM+Dc0YOY0rmcF2O7TmJvHl8xMzajg
zElR7Vpj43xwUQFu9Vd7A3PdOk12egavxw9NiDiqPylxL8Rzp3fNYf62fqTSIdHi
Nv6wiLDRv/oA9olPjKrBNrhUD6r5qYKjKrfNOIfWkBVXK5Ll970EwYEqnl/nsZCn
EUQIaBTh/hfgHrgu3zNPCWJcYrBXLE2nkgmyw1/MwpiA5yMgremnHPUO+OUVW0rz
XgDCmRq6QZNoDgs059BE0fnuu4OImXQK8ZRkqtbZxyMubyM6sk3tjhnYKmo6lnFP
N8CKxtXxDGbgSDuEIdNQBhkOQ9embjYczzygoj+i/een1aV47TZkNAflqjrCCkcO
ESlbt0MoqIk2KeUjHTAQe8Ic7wuutR051CiyG7ZCc348y65JebujW445d2OUJjoY
X4xF8pTpk34E6fYMkDf1s7pqkRej12kZwETUM1vT9hKJAZAGj5WL3dZ1BRietu1g
gk9G/t7AlyUjZBpp0dl4eW4Sg/WVPE7GGy+XSKPttsJ67d88u7G1yo/H95JXHlcV
sYXIsb/vSuz3+tkGLmgvy+TnaI8Tg9jNqUcSBUtq0WVGEBV//v4cQdBSwElC1DxX
BtfOwCoIOPjZdU9QPskCQX5M5ZFMYVUb/TcLAsGaJUN9ogeD+IOIicatLCl8oNcS
pWGVkH0nFP7tinDaKG8TxKCIEVdju0GUAEfYuWgyjThO0lx1PsnUO+uyHTjJ9eld
uqIjAnJE5Skr8d3fhXU/8vMCun5IfbtkMTyLlhh0Jn2lgxAb2Mq3yEHB+S2Mi8nN
DWoP7Haj+jWtVtG+OvQIbsWqF8kMXKwz799hrkfY5Q5b/UmSDeZfKIVlYFnc2ZIg
ZTQkAkGO283Sji5OzoY/e1T8pscaHnx0Wgjq7IB8cUBqFQV94X7qt7IB6RzDPTeK
Ke63ts3A3VWvzVj2R7zbmu4nkLqJbVwEpj4HuesWQX5lDsIQxVEWMBuHQq9f/UMZ
7VDIWwqXM/KA+DtVNS0nmNTi02yAwY3ibqe+Iyrnmn53IbsvbA0JHzpyKl/0kHzO
mkuvHnbCRyFeqZdlVFVdQNWtHyx+mR+ZN/LXhuqMMsGcZ732aSsHcNfBWy4tQQyn
TvFmTi3CtqG8MvQRWeb/X+UUEyJsEe9X2ka2XfBS48TtT+o1xvdHfG5JSbkFAqRO
eZ3vuG9ZIBgYjkIU336hfP480899dA9tIitQhM3uYeYJ0DSHXnP/mbUNwWCcCiIi
lD9lh2HW8mmdfuP8K7SapJdXH91SmdrfG6/X46asI4j/qjr5SzqIgLRsjwSVjvt8
1eF/KD+97dY3eD6K6FnulhpEDGo+6QWOtC0H3fk0moNvSPnfo2nvZStxlS1kYR8X
SmJth1jgt6C4d3X2szfuzalHFbJOmWW5ZZmujFHmKmw/D+Kfc+sR/GmbidyaGYoA
g/KYewl1cJzSLsOiO4UvwJc0pYsxa1lQzFcyh8KohBXrpEpRMJk8SNc3mS7zuurI
75rBpVkUO22NFzyaEZLtOBBfu3aqsJZtOiYHTmji7DrHBz3HEaVC2i1XRkE4a1+B
+tZz79lzDUt6pKtMcJgHfEvCiF9vjUaQyZqC1ODULzXIAlKb9bnWXImiuCvhd2PX
7qb0yKKgEZW/SMrPVIqfVhB9vXGJGtc0iUPMpCmEZN50SXeHHGf8jOX7Qmzq2eWD
JuuuLjCr4jf/OlpGUPSF1heIBctmR5V4dyCIDFcNgHvpATwzErW/eJUM7/N+XlLh
+X7bld5oMqjjBapFAXuH0ALDXGj7jm/JS6WHUg5seQyXgPEiKZoNSKrVuJsMzqV/
LDAQGpjg1j78ssxtvR45/yfP2PElpHtfbqyIUN/FjS9x94dFGVRPJZutjJyJvS5m
9vxhKOSpMf808JxXxYDYX0LorYabQ7d4yiMVIBmdhWVFimsKop05T03SRpt0X9yN
fL8ilIv/fLDbHWgBYITYRJ7ST8v/XItpYfOsfwuE8/xB0+jkqKwzPvzWaStF+/5g
1WUHxeZrEvaGn+rSeEyNTvMi6wXIZ/VoO3fgpDZzJEcq0u3QZXUx7Ge8E+sF2juw
4BJlFaFMBXYVpqQ3xLEvpJRg0ft6p38j5qWwxAAOam40dNcILz/TFOSEgcJiv+ZP
vaQ6yKVmGFHFJofe/Ye63CuZsyEHACwhT8HPpasc1t0oOO0iSTMjm8Ya0ILK7Ix8
AHNCHfUUF4pnnqaHswwbVSG/4IWnWCBfrOI/UaLiR9+clVqZqRF34zHyiEir7gbl
bjSRTHpXiFrXPLU23lwnlMAZfIhoQu6QFE/sqxKSd+UFyML7s5rNiGGq0b2ld9LB
PpzrlMWUGZ6IT5EOnb3blG5XITuVOijRfa3oen+WUlOoG8nh1W5MBXO0Bk5ysIqQ
9ape+O06DzN154+1MIQHoQFw4VFb1GXHgBUKfSxCtD/shUWY+Rr+6BPn1WXHnmqn
YBGGftoPVrIsl5E8DKggXxnwxBsH8DsS6AGsBWHFu38BgOf50/1upV3Ey9rg1Z7P
24zsrS4l/sOH9NbYZ+c7NIXQ5aeCVRWM+hMZ4h2Wkr4SQP4ErQBymdhzWE/54XA3
wnpO/HyDjoCSJnPaZ6DP8YIf61txlN3fOoqQE2gauv7ILFPADq453vOMrJybsO8B
cDhLTEZzCfVPWo6nz4l2eLfx/UT1JA1EWH4gOgbQEyQEGTX8UPfVlkwQ7h6bzCRU
S8N59WWqLGeDxQmxu89T6yi68/bjjHXWBP1biiVBmmWpdhQ5W8K+oOXsZ60QKXOk
900ez3azS9q1grXqc7HUF43+ZGHlXXPVOQlv2BPxWbLbC0XgUrmxUp2Jzdv58R+g
ELP3WtBhw5dSHRDhFtj8osx2XIm7P/xby1rFY1+OkEjuGR0eUTmLmqEt+yeR6CS/
Pe4arctM6faJ+nf5E4ZlhTKu6sdcVED0RQSTlQiQVQhvWu4QmSj4ByTAuXT6W0ZD
lishlcy9EwtBX9A+uknR37nEpCT0sgwKUOrysis+1IN1eKMgmdD6ZojmMY2cjIh1
nrQji7f53Tbv22dNGw5+r134/xdE3cc4rraVfM++6DCKvCFBX3S7aGUYCFDcVz0C
opCKqzn6GhRyTvIVXjPSeTjjgYwdztp+j1MQc0YR4NlR2xHevwnXlUczXaQhbV25
tnedrs2/Z14Y6Sk2vmfeQKVxjeiLyZV+AbZIh93M9f0Zq06ValG675zorUDdM331
FGAYYhx3YB9vmFMU1GCjgA6PQLXJ08pv50cmuXb/UoLd8DR3e5ewUmqyTj7Tdzp/
jarqfwL+C7fHH7HfzC/RAZjPrHiNCaxrYG2QhaWuqy0m6A940Et1Qae0CURFrakB
wCPXMt6RD25WB7ggON1DmtaFnt0/QMdpU1c/Gdrx4bNk1iUHQnfP3CG8J4uhVSJo
Q8FcS1+ucalZ27stpa83YhSemPklGan6wStGCpZgWDYOecByYrqP4fgNjkhodme/
WzcDKWx3HzFxIuHIF15zpO0Ezp6/Ayrv+F5sASVS2M1qCAk/8nXu0BvjE4e66vPU
LObaRqmem7BMa6tfErsDxz1bL4sU9VgtMy2I6RtsKU54xiJSUeCHrFr4+oQanWVT
02IsmYVjB+Zt0C2siuMSjQONHN+g6zGNKijvZj02KZhdQmvYW/YrAjPQ4K98Os70
901vFqLrOgnnRnNvHbZl28zdtFTUiYkuHFSaFprld8pueExsYPrAPqmK9dRe3wqv
mlL9AEds0MRiv9Zs5hmzp7ODRFmW0amvvjZosOiaZk7+hs8Hok/ZxbBJtAitm/RO
IedCf55IUZHU7Zk9EqDF7pOL4wjDCfhwjVNIpOvnn+fJZmrHR0X2xfVeHp6speVT
gvdXmDvBrnAKN35JRnXV12yv6fXycM0SoQ7RRXnwEpNws6juH+Haevi5PdNSvcPd
T3Ae+KsrXtEfxLtRKfte55n3wnmSm5s1qBd5hPQ/4yn2/0Lw6PfPwp6Hp2JUrL65
QALjWdrxJKY4RYiNW+w9UCA66mtxPS0022at290bqTx2X16rHKNvtlGh6VECvLoQ
+0l5MiDYKh6HDZQThSwOH8rohYiwG97GUo1QC2lOaoaiFWNxDIi+jr89xRFezGZK
H9dtpOPL7nSZwahGvyWL8FKHmLFdL0qai8QlmiTk/wkORxClHbb6mfgwOLFC6X3f
sN6o0n2EtCcMgY4JZpFN6KTnXdo/zdJihAYHD0yWYiiMeqSOAjXAwN7kwrizXoOP
YfawhQDqw4RxgzkmJc8eLmgkzxO4D5Wr3VTkcOhbzoG5Ils+ovtYQdSj8nAlA7b3
YIC4Vt0lRg8Xtb9hTMsxZQAL1tcFXBczkRuVESlw5Kc21fVsJnwdnzCVi92/pGRL
5uSxTvQWE6aLsBfLDgVQL+5tp5x1PZ4hMo1J7kyvRBHQxM4W2bd7IzqzEDUKeLeo
mY4vln607pJsP9FlBLNlme0KlN8HnhVN1qsPtc45KSi9rKAmpagYSNw10tf3CiEo
yQRe/W5Z7sTL32DVhkd2cqPQ/TKtKeNAVGu13zDZLc23gYdP0NmWt5j9qdCAEVLT
ZMxcbjYIEnK/bNnRjZSjGKWDYvYHzNBDjH6qkQA0WIyhPPxasuvxFEaZVE4x4YKX
54L6uqre/zPw4MJBLg/5mlecF/tP7nX4ZT9HWAuNRGbrmQ9ap/YJlPU19lSaPlu6
XzGJoQb4TEgK70jg7Dv+uPU36nb69MxF8cSN/vxEwMoxSDDXJzKCtpYe0WZfpMPs
HGi22reCiVcBFrCHDIvSQBnOPT1dzqodl8fWEkYKed6yqmO8/oJHBcAezIBSAshy
21n3bWkVyWzIOq5oYXhfVjtG2kEsn2xauR3+vWxpm9Z39vGRu3fkGgOFgAS19Ulm
i7mm6LzpKJQ1CoAB9cJFW0PpCb0+F/S4/aFzA1DQqjlZYZuX8eOWtglCTL/t1CgS
FUX+zwCpTq5w2YN9FX9yyxwqPVDRJOHPxMkaSPP7yyBA4N1Vm8GuN9EuPGmSuH9M
fUWhOnPIr5of6/gj9Z8cZcm9JA9A1ZtQZGyCc9UpOhf46MFrEm4jhHZ0sjXbS+Yq
u8BMWTSy08ZxLO1IRtoZvW4uXOkY1szIEUCl3u6yjtQwl76Z6j/bF0CdlIsmFVzn
JVIRWBvwzGrLhvF97etiKGkLOWwHwlK60qBo81Ftj4SZr55QHVn9ojGPO7yGsynt
kDx9W9aTB7z4jzRAR34jAlbXgNXld/OrbTGSc3PFunVIQZMFkDVVh3t+n5I0gtiP
31umn/4Cx8c9hB2ZfSXFGVOUkBl4LbBinOTRcB0ws91n0q3AIX/dHPGNoCN6m4k8
ySa3osjYwgp2H2onSN2jyts93icE34ZGNBID9vvQ1n2EtW9VdNHKGVnRWgViAdRX
tOU+ctWUJ+yBl30bbddaOn59v+FtwD5SpAHdRJrXx/6j9Lg2f3kNptsp7rtntbQZ
XTbom/dCIFMkEdrUocqoVD+8mhe3yDvPYoSNz/oF3VLdvCFiKKSZDbQxvmCuIgXe
fdi3v84A8SAA0n+kjbm0EG1PBU1TLYPoaqU1QuIH8no3Jk2YxyholQCKNtwG3A4z
XOYmBkID7VWfg2TF0Z8qYRyyu5bhOBeLjHbDDrzTlBYVhtA20dDtaFxTc+NMi1pY
5MQ2hv13oGcu2dgJE51YpWpCYJIqdXQAbwgNsUQ4EC16ZaqkjpOeyNAMDv4NJGf9
q0ntQsDrayjFy6hJMYwc/p+d5AE8NfQb4mrrJpT2DWc2D1B+ac0SMnxX4C7d2Ba1
AfvNfhKDTEOy6Z9q7cGSE52r9vS0yrjOCVHwhtdW8SqoTnqGLYJkiIVayn2U/GQZ
gwpQqDM5fGJMrzp7pmB/xIEJAJFyiYBvuLco2g3GOq31vqGHgcrszAE3m0+8uA0+
iFqlrLUHb8JDsk47/TtknQeCDYADxSInPBl1ljHz7x6FXG+avJLPmc1WMfgrNKjR
pBz0ZdyMi4Km1PUYMrD+w5G+6Tj5ByGulClWUGrgs/9zBf8nabphQXQWFYldYIoD
pf43OWIcy1nINlY3mxll/085H8XqI6QcbmA+VS57ip9RGRIBWR8FtqLzIvSIZWpW
n1x/RrUFKBv/qfLMLQlb2Wz8rULccQeUVlWC+MEui7xpEXYULqxcy4aoYSGhcuUT
F3JAWbvbEeUSDSCE9HwTHTmYPDuEkrrtj8jdWL1vsM1y7EDN5GxnGY+wwbADOXne
RVV7c7Y1YQJ/BB+LMu22xolNOQZplvZrwsRq7qiVhtK3iNgnlSuFj9g/88HPLe+v
cUNookHhudnLzOImYK4Z5Z2xwF3lEMGHR12Yb0NcG3CN2I0VTTRd6Bu1Qg/6bliC
Dow4I55dSe2tdBIsY12uEdbWOJ6exHuA6RlIGARr/amIWSNxlxP9QFWWIa48iULn
j0VxHwryz9BmzPI9PutNCtoOgs/irkryRuO2Onn0Ijw3M35suGp4rYJHsYPDRAVG
tGwNFygB6OAtn/QKPQ6IEj3FrdedcdGkKF1pV4UPCRgx7JWShcLAejdI+xjcuFiw
6jTaPir8H2seMsJfT9VQzsdAuDl6IWcHeUeeIcNi9Bw+2C6+F9vFCt+DCxoe3WrT
l6Tt9N573BtheR1AD6TjaTbTrTeHgROSdd4n2YvhCDQ9BFyVNyfX2SNmuooUj8mN
fD+gCuqF8zBKVitJpQK2bSgfDa1iMJM/WOX77ovHC3rKPDrdA4u/zV0ylyAyJsyr
b4Tf//kjk4DGkubNhQRwZmAV0Ys18OVOOSL+3KazL7G9QLX1gr3bR02ggeeL9zBA
9D60qcjOuoKiI/Resku+8pboRZIteiITJlkqc7KlNNBTahE0wsR3OafjW0bPyT+y
HeGyO3vKYxbTQ0ZDgfYtOH3ae3AKwKgIImTVs2Ux4TNdUFn29wzc2ipwrNR9yjvB
gFSd9YsqxrNFzVMFzJYxwVSqNcRLdvDOJGZEmR/GNoyWIdM/e4X8WLxIOsbTX3r2
V+9+CiSfMgtkfCjXYDUpsWjHyUlCfGiO+xb5rqDm9kqIuJiJuMkveTssFkVYrllC
ofg7tfApy8wWzF8hDnLdoMK8Ab/Q0+OVaSJsCd31QF5SsCOgOLdWCjJrPO4vfQYg
k+HKi2n8kUihZhzxDtmsDEL3p1HHdYGwfjvIQhbhCWgXhhH1edl6qXscE7Qg0K/C
8SKI7kRZoyy1KRyllUYJJXfJxBUFqgpwFOrie6cOn3+f/aFXZGcUgFtyEQ3nOPOc
zQUPDZ47khpSm2QxHBQezX9dUsU26aj1leh6dWY9phYt6IgqKi58mPlIGZhoujXd
U9kk9XMjubGjqbaPDrHvtb8DZOsqweBMPurtJkaGDFxvVZDaN7fn5DAdkle/6xLp
KMN/CM31OZmcyqfA+4iY6vI6Esx6cKtT0xC9UA0k0mWK8ipKrm/3OCwe/wTJ22U+
vfKP9S67W85s3jT7aWH5D91ILjzvdg+l5EBLy5Rn315WR+0VHs19kr+h4e8afJRa
hajosJV4lYCTqwtkJBhVDYxMeKiy1+bw6gSASy0p86K86YL79urG2SKNfiAn8TC4
N9hgYTohUZMIULxnTN1B1Y08dIYOmKcNsqa5JXretVdUZLiBFpURH9V+JL48yR2N
jLlgqYSkho9VV6c4HslVoSmv6XR4c1iKCn+9Gw+ZlSqzgJRy1/U+nf0cTdT27o5w
3KWBukGcpjeSEweoq/br/aCP5U/eX1GGQHKZolIbwUxCYTtu7e4Wavu0Hmj8aZ0R
WB4LT9R/Wh1ZKMwKHL7g2iMBkC/ZyHew6svgaIpyBUMho006IHw3lIJKEjME3Jyu
HODDGMgfl5SOWaABS9jk4GojyYNrMAkqo2uAohlWoIMipc9oumuiWsGljyao+c35
oXABYEeGU4n9Mkx9lFoHv04iUTMNonIZNRAaWpkX39rPVz35BuBqL+HoWBHvYbAX
xa6brewnOWg85mO/ZYozE7pBfe5WupEoGtlUAIPIJLrzGf3WLxVmXXynJFd1ATSv
wpk5yN7XxjmQkmcN+sPgaAnJk3xVfToDkPRl7clvAoZT81lxV+TBxV5wpmFSTKjh
fh/l6IDba+5dj6A7Wi9DL8jYouF2Ht0H2KMK+TrS6POaXY4T0zoePGJ37LvL4x8T
hsifv2PqOx0P5gl8YyV7y1aoXluYEsh6hAMmbl0mSBOB3GQw9CIIxuEF1VTVHi2e
x530knugI1oC35U3O12VM/Fwkyv8Znud+emG/uYRhN+THTnLYQa5xBnUhTy9fw1k
jLqgqVxJ0B2b7gOpdGWg9muJ9xKqcroPhebM2AdeviaEvn4L0U2WKpXA5Zf5L/mS
sd3yAljSBdx2A2Gt3Q1yk2KcPQJDO7PRMZTm7Dgy8bAFIGuTr49lNrjDfeGp8xpn
Vm/mRNLFajkX3zgOIZic4tp3W5o4ZzwffQbeylYZxw0CHnAmxmX1OFEufHEouqfc
EInwAZDn4DDZG3E2q2WUZYONiusuuoMMfD4Uf3kWoUahxxdXcnlB15tAZlGjev9H
y4cT3BmgrnfJuVUfYABDvGdGNP+MRpYSJIHgAvqB3lGGpuy0Z80CS/EeJGEwV+lO
gvAi6h9QoUGXxgDfmPuE36bApEUsUEfihV+iG5WL2rQjxHvVG/5RrQ115WakOlIU
kVH8a/DmfV0gA4zRPCdHJqdN63Iy2jBb4+8hdAJFQmHmTK353N3n+mbGGSmiI3ah
o+aque/RdbCnDuD7a62rr2Jn2Pm9Gcr2mBsnmgoB004EAVYvSv+Dsu9ybrcAmfEw
/CJQVhR1BhGSRV/u1D2Dr31phuUQbrOO4j32xb+/GLZfiLzo1tCXuppUS1tERciW
64vfRvf0XxtyM0v7/j+1vFtCjVI1Icutk76hEShS8cyK/6mQpEo1vj7HGynENadz
iB4wle3bJhO5AdfMcAsIFhGSC1ZD6jAl9qVxinejDVoxuPq9wPcYIQBLQUNrk2rc
VCLWRodqnuIDgPBECQeEsCJXehqOT1/eRMLxdUIZeKWoFF1OEMzn3sCy5t0E0YgV
asfBhbBj+Bropy9vZEfcZku595Dw86s1RoosB7eGSm+rT+EcZNmoAMoFPeM4Myy8
hVPKOHtkfTRxZ0Jk99ogytOO3vVC1GivCTWSDwHFsrvGuODzwEF1Imwiz8fG5fr8
sQtulj9sJWlK4e22sbf2m30Bq7trHW8MdWW6zQg2BYO8NElcOLg7pIibQY8yNooB
eO54J813qwpfYPGqhaxxErumdld4PNcWXcmLCsSSl6Bl+UPK7hdzml/u7x5gNdPA
Xi9ObwkKhKLzn6/LRgKAVQBU2U4RPo7jKhFkXmhc/H+DRvUJOidERSonimRBeuW7
6fpxivGYcwBAv2QSZqi5g5VqYh0PabOgcMOd2bqujoAIgWzr8B3XM6IKnFbN5MV7
jX0AXg2Zy9OsAz3nfTy6jEhPcrvUySxGIEoXK4oX/cuiFCKnUV0rRN5Ab1+cIfUQ
i6MR/73/WyPXEwAMTh3jZ+kkij90wxWz8GJTuNkjEcbqScnwFiFbZ1N9f/Y/XWEi
9tho5TeTyksfyjKBGhRxpo1nCrC4qhF1lHohVOkE5wrMam7RUR6dkoYh8/+BYiyn
QOQsfb8hqowJGe/I/fBTAk4NniSKhU7Csgo7F8Bct2YF7F8ETWkoHYtO2nwGvkmS
NExsqldE8vrLZVooA+7TZRcGSe8ChNbpxExzp9OwOT2jU9LaQ2nYzcwCVtgio8B4
3sJwFlwQn0dfkfdXrYOI8dVLkHGlXF2RrbWhHKdz2K4fKIoGsApXq6BrHEaJbl4F
nnr1ahqH+816F6vMKR7BNCKyUtTmyeSbwam52mUurvWyyawiwmbRhucg9PlnH9qY
H14NEhm81sapxMQy7VbVAGX9u/Mfo0xp1wZy4uTiYEj0y8tBQRCdUu8iBhKPUtMT
MLYfnW8g7aYw9oVbwl3efwjaJRNglrGCLjcVTVumbo+rMPqB5l/T5JwmnijbH7xc
Mdc2mOhJKowoQ09xJvZF4kCUeDkXzYfD4XmuWJvbyjFpFEqHeZqM3QItKjkTnqFL
PmkduHiQyvflVgUo1OHFeMT2z1XXrKno7vLQRLY7Qpipm1x7BRhRXOLTPz2vu5Bs
iUr9gp5BCxwcj2cGNt7AWZB0xEqwPkdoAytNl5PNx8za/iDJn8V1zMs/ZKoFQ1PC
Mj7zDua/QMJjLiK/ha+GgcKyh7npPNxXOSL7mNfR886SlBzZ8phT6OwNK1AH8D0T
DNRtqaK1Qmx4Hwzk38HvHx0e6GQRmzrK+WvaFbM39KwAQoB4+Po+OI6Roir57weS
BRPqv1gJLToJipcrE/197czx4QZCIhN4p1cWnv5IzDITW1TfjA70Rqb8vzdsmOic
NguC7yX1KwsS93K7jb1Ianssh0cOSwZGE9SkJAMIzMSG+30LuQZJOwB0m/OzYCcg
V5xY76oMdBbWpTMbcnKuiFtY7h1Cgcu+4nJ2t9j92QUS0s0xKYiS8tikVXu0Ii/W
SjCXMbIIzxACNEszRo3dRfYo3W9P0QUUU8PfilN2KMzRnR656v/s8lDGKUIKDyQJ
Je+InbBIG6rtodRwtOX0VoIct3Adwd3gNMtrA3tBZIfHGoqyxasskUJYKM+1Qmg+
b6vZddNTy+xtRAUDMjtHHIog4Th43sDgq17sBmPfwulpcwtvMNzd53trKNHW5aX+
R/6oFiBLDKH4n28IWUxoY7SC64m3WMj2U0B+yRtzN4HLnXAN9iFivcoQ6RZOZYYu
JvaxVyNXpyKRrmqU2O437cwJTyU1XHWWb6W6/x2qVP15kO/CwdMcDB5jj+ulIwzr
4KvBeHLv4fZZUTC9gwbxtv+wAX6MBBFjlC6+J9xUOVjcKH0CFeKtsLpNjYg9FlWe
SAnY9x7GW5ZlzJSJmeKy1QfbHeq2oqv8XyGBsW0tXyjQnU2xv5Sf0kQ/e00I4ve0
BPtAlJwxLdgVqyWAMtF326ViLAGq/3dHAPj7PZoCVCzpIWPFs46IHmOQXLeyuJYf
Y8BZA+oegvCoHWy/GkjAjHLHowk1FRUSQJVrT7grSN5EZccrYDdDjGCQbnf5lHmW
ztaFJM88hwd3N651Zgqr8iatnu+M2vU3WJ6HQZXhB3MMwyA7Oe6+kLon9vCuoSNM
xjPzjy7As+PSYDscixXYLsr4tXDxOMSnyr6i6YjeC5maNjNOQsOjKV/OsBBzHQbQ
xgzreaUQmtH3EKokfiLBUpk3tuaL9eS+SRwpsUJzF+BgaSSKVYjvxR5AXPlI//kZ
vAFZ39PSNIuUpq5KFoMyv2VLzon1X4Z3tKIxSrY5JqycEOO6Oa/Z/iYS54MEMrTi
nwB5ksvlM4d7hHbyMItSiebkDLTNe/ZrQvUHnAyftxvzUHws85MXePskpg4QJp+e
e7lfCjSP1281jaPV30JztG5h969f7OBKjr5uSj1E3uwBXRzWBXf8Ep5E/xOp0ipB
XNFr/pjPftlKXifjXGybBcI5GDCfojI6dcqa2sSmuNuLMrXw2FRYviT8cZ/8MfRc
fCA1riXLlip/x/fAlgkQ1lIFZoDiPa3vdjdPkdX3J0saXn7Z6xvII6ThS8u24Wam
XySBrAT6QDqBY7JSnCXBxVFWHL/T4fas7ZJ+I11aZRHygGO+JdYuBvEJQJrbRb0W
F/W5qIJjqiQAMjWTsGqkKtc+97O4RNF1fiHzojC9HEnr+q05Wvdq7PcQ7sCXvRBP
JbIj9+vSLglinlNob2/fVZiPrQLrNUsaFCytsaTbMyoA92xzSStIHpR6B2FatKN/
OL6bx1yePbjlO/GUHQkQg1ZoakMOICRJ7GjXCkfEg7fQZVnV5BUUhhmC/Fcx4rJo
p91xslW7C77KI5PiMmHR1M7H5rs6fPLdqsj6DQzGBla5A+l2w4ieceqhpcY0uHoU
+2eZFfjZ8/eOo67Hrzwnn4PrSnlkwkzWt0FWwDBTaAqWua+mJHIveeYu71v6AwOt
5IU4I2nF7tNeFGh7RuLSGjtdnoH5YAqsVbgsbAyGpNyzpKRcpXgk/MoIwx3xJFN0
A9ZOPs9W2e9MpsJ+nij02P2prCBgNZkL8mQ78MV/AgXAx1KIKSfvd0ium4tip0sH
giv8zzrp/1fH7thuorBEIxYjndmBAY7QY0TNqQIhFzKfTeQcD4lWpZm2715EhGK5
mb3W1jVeDhCPX7wZPOd6BuRJYrHmJkqbo+b92b9VoOJQThuZQzYwgxzQ6U8rKtxt
c2BQ7aHRlXGvJ5vK9qVqqq944QdG2Tp1zMPqFXvRXW4FaTPEfYDhkPdgrld/nj5U
YFtZpHQ3dUL6CtkcyzJs+6IuiKYhqzHzv7YvASa9XqZExz/AimDf9jifaWNqVxmx
oemXQebP6580xbIhAjExXvphQCF7gixThJb/pU60fj38r2k9wfIUYtaFqNCKEyHb
VadetUu8kItPn2yBkQ2iQPvqV7aFSZE4+htsC14wuKX+qLA59Mh/aOPdfuImduSR
AsGiCQImbli7ivafGQ8UF6BDO5gZPUrE2e0CoAfGqMcc1vFC464ggMLd38hCUS9C
Ef1E+i61K0G825W7zhsyoD17yPdg5loAxlnUAcR4ZiyDXRaLPYfI1YBDm/P9M3lb
e2PNVg9gsT3SZEmbaXMTi6xXUF3hbOS7DrjEg4PwJuv4IO/O/gOn97X/mb8hx+h+
22vLO9JC07qF9aYZ65kT2CUrObWsVp+CBViZAtr8Er0jWXM2/iJO1HC0KARW5sID
VJT98uQmyjyc9Xns2Dj2noVJR+omgFbpX1XCWe/vO+V6SJK5ASZxwydVaIpG55h1
2QHz7TuIcn1DlS80MUtQwkN7Zd/Go00untoy+im+wcj9GfcvBjfCBssk4XeJBj0A
0KGgPlDSJxzC487tKZanmqXOhkhPysMjcL164D+v9IvpKB6CucK+ime54WS/z5xs
RdSpu9aLyQ5ayxZ8TJ5c8CJu7BXlJ2pDVFYyShWVX5HPHN+grqZdha+7lsCsLb3y
hb1svNzu9P9I2zViV17XGPPUwjHXThl6miwnpQl3BFwQ+lZlEmXpHcIOnKDBzj/W
xNaYkn9kEjhEA4a/nmVh9F6aIYEOZdk3emBGQpNebUA7JJlUo35t5W7I6f8vUGH4
CakO/sJXRmjQcqZC57HL0Vm1NarJK2vnlxdFBbRs1gt7XqC86XU6lv80Ir5po1X9
ihtJoaE1isDmt2owItBS9u+ib3cCzg4ZrfRanwvZV5rN9MiMTarFsZllDMON0bB2
zXmZzrE5Kn0V17KyK0adeDonyAtpXhdL+9a/ZXlZSji4hgHA8CboKs+AEP6sgVuX
lds7EAub3o+ZfV/mJcDpG9TQgHY0K83QhSSgQxy20zcTZ4MChCkpCrIybTGSEvQ3
FIYzNqBlPfT7LQDbwpAMnSgd+V/AkjdF9u0ojjjIahm132O0dOwaLwly+0yYmlgJ
laBRG1fo+BOFSszyQVbyH3uVXj2lH/dsf4oUnY/iEFWBoY58ROzdV9BAJ6/bbKC0
X54Gr4TujlXu0RYDEj1Wn5LXefWgZyVe536nsnkaDqi01jGx61jDxbct/p28zSth
9uDgdZW7QlOjtOAS3bLq/zaWZ/KhtQahM51ToxSW4W1g68vXlJcSC80Tz6EJPA7m
JBA0GPNvonB53RNAFyGO673p1XR70Tu2+ABBH+AQblARGvcjFSiCKSzMi8IvKgE7
mK9iEg645JhTlQltSjYWFXF8uqZsbQqwGHLrbcaeNfg4fMZ3rbYyXZAgmkZowdmT
MqISKHJq6NmAHdKq7lxDZuSOvN2lpeyQOxKcZi7WabgmwM7w41wGSORQuq1nxkf8
qzHl9KYLRcQsYgjAFF1TFMPQbgLeMdieCdISoRxWERK8CSppIXZVEDlKCcswAVfP
f5B6WPazHKAjLO1i9xUMqKqHw1Fe5fSKOu9n9be5XkcAkq3FS7N5jBbt2SVCZkhM
CJXWFg1kmJyRY1AjtxeEeYqsi2Tm5bwdgtDFqQK87tM0xlaXKv4gdQhTmxiWRuQ6
hsCHNIqm1OLrR3R8z/vCIJgF5bC+WmnGJbWQGRR2NwWSTjefcuNvhptymi1nmCDW
04WJVfaaQjvwR3MYslg8oTbHKva0E2V/97PZTv1URSPnUwHMmAuAvRdc+NXoq0ob
RcFs93xerwwDIn9jviq2iWgfiOurE8C5sYv0NoIBYbqDouRukWSLSnVoQSPW7m+2
Iwgva7kF9b/87kGG+GfBebXS3hlnN8dbAJnH1fjPgZKoW3pwtxGI54E3OYak/FF2
yvrg/dAULTYWW27yMwz91Xhqkv1lY4A9DXsJVWBveME71s/0DrpFbKPT195kfQOS
OU0x2hQ2k357ga+WuoALyAItpDDhWELn82xfD3vfpDv0uF1dv+4YLyeL3CnE96fp
zLG/YPRK/khg5BXxfPJKnKLUzm49/eUZekAVvbwdeA4iv/OLBpo9XJiplLaPDIRu
ECyFQH6jQoobvjH+VOeFJIDMmSsdiyNhlsLscfgwGzK8CSKRlOFb1vuWfy+6cy3Y
5ic1cZW9ZIIkznJcy9bHMZUWozNPvVphVnfzQCcVsddP4MIdF1GBBtypx9Gh8eme
1z71u+Ia9xHB0ye7FqRFojwMrEXQF3896NeEfsoNtwKZ9pxBrp53o84KPeOClbwa
uzyisgUt5gQp8eVG3ETFKELwMt9plEYKLlg1tcJgYsKBAaHnUHSh1dBr1WOpvYYM
zdxJ2tb+/YhvD1MFlLPK7CKL3L0GqExEIP0OsMLUAJAZOzZwQPxAOGd9SImbpsD2
1QuHar6BBLQ8JQgqAbn2kpDXjI5Wjz6ckgNcIiMULCTapRlGllurDyAOdwJLS7cO
r0JtgdkAku39XD9JROukwqa4ETB0wEyz2NKU+jPMTIdAb75Xl9hZ0Xnt4pBYUkK8
sUZPldA1wnoI2JQJ5d2eiBwDhjNTwP1ziVUw7Jw7nnZc/HLrdx7JQeSw/P1cmXQI
om/H1/BsmsPMVC4H4YGkT/86XliNC2xcjutGWEukhplh9XRsqxjeQlL5unh8VWNP
lq8KNfi0v6XNhaByUTYoxQNG5cbR1NixEePwDFCHo6V5I2F0Y71ME0c/Ate++KSL
jQZZpJDnJ5LKfUpLxDR8K9oAgnhrtBgA2p/CWTuJDAweg7gUG4xpAIEvh1C44a2u
UGhYjZeoEdmJtH2/SQ15O9mkEDIAZvTTM0z4ce5PUdcqGFpZcpwPL2jp+QpgDbHG
sfcpmt1KOxBmIyGYYAzNXkjt4qGTtNogQbt2WzKIj8RYaNT3JDgXQSPJfbN6Z6Up
85IZGXV1O7Cx0eZcpZA/tfx2e3FR6V25aKFB0SQi8s4y2Q2C83wYyBACkVqgLVIU
u563aRiWbHIuKZCgKWVk3W8IiVohX+BthJlcho15O93tkDvkXQTcEyxJUi1eYzBQ
UrUCcTEOMyOgWBcyNBc7KrBl/5kHMMfX0zG4oPbHB1UhsbC6gCrYNMufJjgiu1ov
yNvtDxdv4OmJRCjfaqRKDRWoiMT8EcicQvZ+4B0ma4pBU7wBtUrahD149cu/OnJ+
OwyWaOzFFD2EmpBI3gNXVSIVuuo8yjSxqA74m5X311Cfltuqj+5AT1KWgNfwU9RD
sUrby8Lb8x7+gqCxImIbjlrdsSSNcGNTplgFzHaynXeneTAq9WJF2RAVi5pOa5VB
xs0igeLOQhG75LQuHO3ZMW4BUzD98gQ053wAbwZJeqz9aDEPwdaVf3xU8xVroLPy
7x12kgrWl07Oi4yLrZw+XRp2RyFD0aHby+MJ4xd4eysq2DRezagpY52E7u/JJ8B+
zJINsNl13dlBphXKLu1s5FoTeXFDgK/V1TQwOddEJ2hWWc0v4Wf6I2jkUb2a9m3S
VGSjvG2Hgu+8cIyLPvJNd9Hrt8hsUpAu5LrkaPlU1uExDuM328xzdyV9Jxk3pR+P
kwWp3XT+VAs/dbpa9dMGbgo5LK6+ECUA22eCwrqOKRtB3+xfBbq57OF5C/SSA6Jf
dXhxpHzQbgbkF6xqOEN7yS2vHh+Yrv9GNwdpNizK4LxrMpp/hQfiINHjaSxaMNYC
NG55IIQm901wcUKXRe6yUeuvviFkBf3r5y8BNAGQ71N0iz+FITNl+NgoaYMliSJ3
WP4goFqoqKoqKU+GqO/fEDEZWxYcHRvaoq6Otw6OodEXIPttTkvi+qSgM1LPj+LH
1kPf7yPXfBgEuPlfrTeDjQYLPibb9+n+F9/lHaN1aAg9iCaDLDOGy7+6RqHd9GMo
BjoWZC6fY+iJ5AgQxpKSl/3QA8f6P2X48R21FPedwAbXJiBikl5jLK2/thXIlR3v
FJ1BCzyt/WXbgcysNOxcQRZOFvGyh3uc84p6+cU8F3KArNaq8ck6ayxR1rqWrhH0
2F8kyKYNmxCVPfQT2tEb8eWqdUwZ/HDW3hwvCybmpaByJ3mDLrPA+K+oCm2qp6WZ
xFhG9Z0VAoDEdiezIXowP0sgTDjF/D/v09W5vkSG6K+9i+7oP/ktdabNMBZpbDDL
bURvXuoaIC8KShOTsmBcSKAwNy6aLuzDzL5C9KF4OIuGUdcC8//OBDJMM24KmpI3
IFzYjw2FP0auneGbMIzrfEQPmi8pZEpiKW2cNrgljv/6o4HK7qBTh6h1aU70K2ZH
zeZwF8OAgk4Lxu6T1JfEzeivsiRzacEjA8IsbrUyVWFulcxzD5zfNmsqWtuuFOKe
IKNig9Igrbbg/N3gTBetSm8/wS6BrrNFZ5n61zq5AqJ63OHypE4mQnDmK+Hzp5T1
ziH2GUZ61XBSjJjFcbOquEUs2iemE0Q+WM4V2SN9eSWzYlksFDHP9U7ZvO/uJFgB
lu69byfHzqNiaTYjALfiI4/DEnwlNU2j3RRzwkOA+5R4hl4t+HvNfSaUeCN9ON5r
KBCH8JEjSQ+JUxe7hOMnpzgPwE1tnnV0h3b9MsKViJKH51KcywMQRm9/lZPh7yEC
gQavKpIG3AWoZQlmQgEwypmovO0VNehvTmLn/N2F1Bkpl6875Rp+jH2devW6D+ro
eX/BZ4VOSbaqHGTDc4BI6jcLqwrvUJPHFIMuWJxaSsR2d5yzaa36W7njYyIGRt6x
BwGjxrqNCGSSarufxU9Rk6Q8n3JJjVPEZ6rDq74Nxy9Fw9B5l9ZUPgxXOXoVrdTY
AVoqh2r0p8EE3PD5c28GM7j7b5memU5v+RoTCTp+rm0frnmec2+gcctzbpOeecs/
eyJ2vbLCgDx8o4arvTSWRQvYriZ6uOtASHX8ZXoe3aaxSNAH/3VaE5XIWytyaHhN
6hS7wECHvwpvmFXnLvhWvdvSyHL3UMlDexW0BpYhZaKXU666PVP5NaR8/maI1Mck
+qGzVNfGZ8VBj9fUBX0buXouH227+Bd6ygfmo8hqwj6L/x2c98GWotZvAPP4KGHq
BzEDJOJNoyYl7ajWJ6mPJqAF7YWaxm4avoBLEZ5fX3tdYRmkJ59mK70qDlfJsJ3r
BMQYVZrc0heX8u4EY1OIbifqAOyrYzeFenfAjoFmW9HBHxf2/AUIublF/LGuKvIg
odZjOoEvoIAuRcJszPPt6ytMJCIjNxx3ojDKoPgekPi83ZXUGtbZ1Z4pJIII8dDA
X72FtOyb9lHVyDGxlZAoLGMixlXftN3JqnGQNKTpSeA3Ax5zEhjCzi83wM+dCh4+
DWcZbte3K42cgMIEPrU03FxhXXYf2EfeSCNuKu8S4jOe2KrbO9zINBQrY7a8qEX/
6o0Wc7nNfFgMk+EnCVZQzUCrqDJIpDwWjEGrY2t2GIFWtWGBHcIzyJEauj6UBLNQ
Gd4MQNFbyeqO6qPLXtYS/fMIqSXU/+eNi6mJ9iNByLi9BTpaw26N9RJdqlW2gI3J
pL41FBQkVyB1EfLeQ3hYxPfkhgF81eJ0mPN2vfprO7aDdABGl/23ahdG4HbRBFZc
wkcJiJ/b0jTgJSIHCXZO8zv5A3SrM0BKX/U9QKBxFev3WEzhkitjuAhhKKXMNNJj
oxsTiT8eX+xxP06QTHizbdtYkuoEtFtEg85/Xz17E5xDN6qcBDue/R6qdzCGKfxA
v2IXsCxyvAw/jcpAPwbbDZT3v/qyNysN1KKaMiQuo5aFapuL+9gXuoc8AfGcc7kt
kYEICUBgrz7vANQ3gbDVTEf7EWqgeUXLSam/Q/vEY4YmKB/iI5gA5DvAlmBzqkzw
ekkcPYzt+Uw9HmUu0g1DsWOjvEBtS2MEn26JChgMNvtDyrh6C/oAVIt+qnaUNPeI
mshQPQqclvFa09gxFekjAlPPV12paCK53DUdxSFytaUF8/3X4znVXky6h7qmmDwa
tHeILSB++Ga7hB63uu4557EFp2u9A2on29MoBXy7dc9vU8OMqOVw7SC40zchyCXJ
IqhjVkWyVTvnWFKI8nigdZ+kif9KMbJwtpUqs5KUIc2McrkmrWi2V02fMNBVfWhD
/1nhL8l92oahLt31Ww3pn9kySJd6LhHYGpAY3w9g3GJ/YT4nLOYYMkRGtxUZj+GI
LOXWo/uE1kCH9WSVtNSzHd5TVD2yTSrZYT97PMon8zqWYjRDQnqBLSHewu7n3Jot
r7pzlU4MaUopms8shnw66ckGbKGY7JUCXfxXUXpAr2AdFZdx2mraj0dNTk6WW/zv
nZsfPOF1s9a8h5aDY5D6khfHQoLqGJRHa/vm9BVh4yVraywTqW7QS7yrQFL5iSqi
dz3rsXyk1UHiBhtMp5Th+L8KfCI9+l0jqzm9bU+mDiRecezvhM8OIHqirYrwf+qW
sBNe0tZKeoaWv06dXE+Jh2+Lw5EWyZNHQKVvzkj7rZlHaSQPj+YrURv0NGs6Ns9Z
TL02gvi69K7jwYOQT9BgzzWn1sgzd0aeOZEu2jqCncSCzy5aaJttVitWWSzgDsMX
bBVlMsbM2rV9NTzCedvWa/oYam/FMkyunvgm+t3hJncISoDB112k2ehGbknH/0FV
lXy3KRjQ4X/QfpqhUe3Clfcv1PuRHLFhfjalLVuFdhQOrTjsD+fxYIRQW1qsfT1I
2tDb2TwduNv+kP6HdVobAiZtZt3EV+oMg8PSvPL70mMtVX0twyQrsB0GXQ2AFHqi
mefZQAyPtg5hJWfyIsCHb1LjZrz3v0okMJiVVXy10X3RmONNwtQVQMLbg8M7HyMW
kzyjvi1lEF1oXiY7aksKsAe8D+ZRKhoRUmu5Ke+nQUqF3V0wz36Ia83bu8OGKDXH
U9GpY0hOaJ4Ffptl8bvhQWQ77rK+L+JRpo3iccurNR1Pw2HuzVyWYgTIoCCRsL35
19ngKhYBFbYmBrY9duGLGUK7cksnWOLFvgUMncNZNad9dlWD8pBYP5T7b0ZC9aCA
n7z+GVP5Sx2dRz7rc2iE5SSJbYxiOeU3afLFNzPQwMCEnxS/N5vuqKqxqGzxaQoJ
oY+KtFHL6YuEiVtoq8I8qFQy9nkUWNOcwKqhBUvTszozfCRjEtCHkxtyJrz6Y4D/
y0zY1akIM45rVS1URBtJPDpaEXHwQPhrawAl9QFVLUl4a5EVyAP/CUxCChXFDhVH
m9pdRUwELI7AJNVyFvpmzVCrlkpDGXEms9BIvBqVij5Yd8ArgaOqJmbUe84hVZip
hdVSWB26B70KiPkB+8oct6p+FONBs9h2eq0b85hVh2qgB8VAZ814CDnRmVc4oL6L
03Ok9liDbC4RNM/AF2b13K/mfpdWZPDjHTRt8EMBm6ibaSMQ5FEqEU22LE2HwM/M
+T7P0jmQJtaHg85s3xEtQBZvx/WIGlMmNFiMyCCFYJvvcDWP46z3jPzNUOQlVcuJ
D3Eds+RosEe+mutki3gO80jqqMqMkLJXUFiuvdhRf6d4YnTuPT4LcB2QQCYxZLNQ
4KePsqysMFE/bnk2AZVXCtZdu1tdEuDcsiSK3V19J9EEjaEE9jV4qJ6STccUw+6Q
3QC0REDfhm5a+JG9AkeNbEMMAwDhG84iofdXorkMkPCalTo0uBMPoyuRKlxn6JCy
KzFZbu5DtWmAueRKOGeP4VeEaOgiHkrpFj0wsTS21TbWsmQ/6C/LClrLcX8rm0qP
J2z1JZkyG71oUZfbD2qvvolDEA5/Psw1JkvNjt+ZbkvlRmaKCysTe68R+X3Y37GP
q1519MMcJYTnVk5VMrR2h6+mrI2EwCATNDkOxxKqs2q9ggqd5IECrLwn9Cx3SDm9
I+O19PxeS+/IDnWQTzOwL9Le8egZ9aGvzA9sBIaRYIcMCCuzpso9+yfnyQQPOwQs
bcciOApTzqb/rf4BxWsutJ59djvlVeelMzevC80vWibFTcGTrKDquSDkbLqLxUbe
b9nmkzZlQfbyavsUH093JhXX/fbPmpZMv2nXminu19rtrciEWIhZR8TYLtxfWRKh
F5yIT32rECW3sCz1tK4iLtYY/KN+/35j8VwpYZz29oik7Pim3YVdTIzVxEAZAzVP
LNc/Yap57uHM5H/u3tmhi/nGtp3tYzGhEN4P027g3wHAFBuDq+0jriLxUieIh/aq
6CPNZK2xP3XD/gM3/zNRZzhn062oHdbW7YMp9uxV70zk/k5U6P+3GqnMk2Bfui74
JArJIVCbMexV8AwDBKHPD/yA8veJOnWWvgBp3uJsa4EpiKx/Yzi/qrgnktzJJeWs
yBtlOBB2oxxSdGowos3nphYnliEXPZynoRqF49FvUm3ggUWupqTcNILFUbg1Exv3
Pm5IfR9a9Gfa2XjGaUlLovKibn/+8AUOnmfZhdtffLb91cYfAkdglhQiQUEAJa3h
uO2z+di1Oor5kG3I4kiqTcG43w1RQ1/7hLBfu3JQoV/7jK9TtNTUZUGp4BfncnpV
HG82CBAF6Q9t+byO7FLNF9BpDJCPWzbz4YXe9S04P0YQNAoHWhROMj6NeEJpir2V
SRzDS4A3T8g21u/tFldyIx/9cHQUPngyG8K/VVU1SY7DatTJZhfilLqdEQye7v3+
39bl3wMhjsGNX8vGR8p92hOJwGMVHbxHA5DBfVcnN1DMAPFTVyYTw6lN0PWDiTPP
QLF5eeZTdEimfB6PtzfsYqT3pRX8P4y/sAFU+dI4L9h66sFGexs52hncc+1A/dYb
KuNl/gFgZibKzYsfCI6d9AwMV00p1l9ntqsrru7U5GIbB00u6Lsm9OiIQhzWpNhn
c100sVHVlYwGtOgKbt2hG7wjw+TKqb4Q+znDsN5L3iUaHvIbaOASTrTYTma+ETQv
FWtg/187gCZELkHU7l54ffBvuGnSCIjptM4ZLrzdi2XwLnhHOUkSctI8Mrd/ui5c
86PYGXF1MydNtU+VAJIF26xVbC61MI6DZ1SLGQqB4DGJZungh7HtvRac1gpKIqkM
y8Zz5wH0aXDk7hdlHWXbrQJqZNGzW/7V3LoA7FaWglfgxthMstKQhD+Qez6EiCbd
58wtncZPjJ7cMj0U/qaZxWcyc6KQdB+MZRK39CoRaibcw9TsXcm4UkoA2Q4i2KI3
EQBP4F7v9ftrouvnKYlxoe3LipeALLKK4VxedeExuWTV4mkU545E2NP5+JuBmjuL
goSwYwTqRW2fhV8r9dIl4x7RFzU8G6OsHYftxZuhV30CqV4+2K/xeRvIDdLN3msm
zKjRZF9fgXrtrAgLR7tcsFT0pJjc4CmiBNMzz7JaRULyjRqfGI9OJsIwz8CD8uwN
KXWG6GjXsLcr75NbtHSqR89WVuuA78qhcnzlxUUjwft09Q3JW89YUeAbssvVk2Hp
V+OO1/6t2L6bIjfF4Ikoand7IAlLbhvpxcBqLe1NlxpdbqyRccPm5c4gsJeYOHn2
SkJ3La+SKM21GYMSEKqMzCl7PPse0frMGt7cAx0Bis1TLvF1wCphlyv5PstIf8cT
Oem50cA+X8zvp+EdfqdZGWytwxra29PeWIOMWP+QcqQaQFso24AJxzm3TY6ZLqiN
lAbX25R1Vd5gi3vv0HksVwleX69OTMpRcO5/JFgtaATWI6l6zPpI0FgNmJa/8f5i
CB38383i6wZW9tDt3KZyd/5PYWGkdgbvRMJa15Vl2k77n2ELtiSANhgd2k/lTdxz
D+oLZ2D7HHNs9IHhDzDc6CsNAELR5XTvUUtHX20OYCBA+sY5fTNtEwxgF4V7q6uT
wXHoD7WoP2F45eRhpamAT/clLfhS45Nehcovmrk+iyQdt+ADkSV0bc0iB17shmbz
HBn7eMGbL9oeR0J0npx91cFhSEtdXj/8Bp3U1XJH75gB2/l7yqHCMpBaoPHbEsID
6rfte6weEUC4J1VZHkWHXt078L23ZROq9nrLrSkYHzd8Uy8LXpT++vTzInptaX0S
hPwJCjGB7zjHJZHdb1mRP/OF/IxBFI6QigDwE5qUCIouR7Vx+viz+vqdDTEL/YJM
t7wZatXlE5LVjinphGiiK1foH+BrpSDogHcS8BznWEYkijdgQBfxuZef4GjuVaOP
QGYwYtJYzvo/lpJjzhc2bohH8tgo8/kjTkk1WcbTGtFsc6wUAut6BvPxb+5TZPDf
6T5RPe79NzovhKPFv8qBAfoeh9PNOwK5qjjsxP49Xcq9VCLzkCMi/eCwoJgd8ARS
5hBjLg+ZR+/U7ewbUFFOU/sg8mKLF5YcXgLa1iZA+cHpmm7lVJVF7nlOwBfQedHJ
9PP0sFt8nb0tC5pH5Hn6gRGuQNzd7wtBg8U97I6UE8TMDksFKC8FZ4k/EdUo3vrJ
Qu4VmNPsg/2v7QWVmFqbXZMLVfFyArYUbBVJ/hByJTeXh6/KMkOOQYVQpKi9m5dP
eEgF+Q+yigXcKnbT6TtaztfSWTtjM7eTsS52So13zOcpkv2lxIHSDHZtLvGwTKx6
6Bfqxre1VgFgq1uropAn2f7cfdu2xU1jD9FXa+fsJsTZW0rW8nVHnqwjVeAyzNXp
rUxCkdGLBWu5+hFjOiMysPaZfa5D0xBmuxq1sanYztFsZqSyIgper2hDgVxAGHfW
E6nHoaF4N+/H0Z8g4W3mFxuXf5OqXbxMeGQ92t3WUdvhGX3cy7zqv1qoBNWPf0Pe
YxkWRiISm2w8Nw46WxlIz6lMrW8MXvcW/eWt7kTynnojTbg2K6+ynM2bzmp3udOp
tG+l0ZrWlwgrFJziA9Rl0Gk0JgAf6nx8x+6AZLsteCcRQav88bA9x53epUNL3rsL
VYg1gQl6P5HyMhBBE/dJSFVjBum3E2XSLUszLUNnLG0w655T4HPUCG1E4Z5cJiR/
Lyi8rK7ce7NZf9g7HKdtPOH6qyn96cq4LxDcDFv/eCeEVo9v/cntfnh2vIWP8+g9
DvwoHLAiZxTR6mwiLRwBFtqCKFZvJS2ii2uVHYVa0o/6XoMggXYoUHqFpcd1fUBO
yU9+xYi9/bNvO0zO8ZII7tgVBgtwjyOHYO8RLb9xw3i3xU8ZEyouvJJaz8Y6VMeO
yDBElDDSHmKIr+tw51MB87YFALufm9C0gPtExkIFlipNOrGI+pQ+9viiNP2NDfuT
bjuAFE+GKIeYkj4PwC5cmduCk8XfsSfn99BkT00f3OCC8b3NuxNIeRoPBHebx/sU
3TOp41ZIyOxn3yz0hfKEAVLuB8FvXxKBrDD0Erb8Aey55AtNgJ2h6D58w0p5pYGE
aA8tCKty3Eu2IKrTxacQEvCeb+8Z0IHIG9nVrM5LpScgVOEXsI21O3wcb8MvNJZz
a6VYzzCHEaU3mfyjocfSNdtsalZgeWx3tKEg0mSmSQuDujz1wanc6lnZX/Bxo+xE
MBqr1/Kt81UoJyxv2pogjzSTsm7dPEWjsBkz4k3FzIvUS5NGLcLQ87rVF+NIDZxa
R0czysgFFYese4im2eN99fLi5y/lY5pSkKv8r23o7lxj2VoYj8kWNJqGxEIuCuSD
LCHugNaqGiARI2LVytE0LCPBlLv/GvNhy2AIIsCv7Ku65iSPa24Bf5C0XoKs+H87
8HDYuL++5gMSZgyCcukyrJu3ovkLoOzryhV/VmsvJtphwYLQMJQrhE92C5M2m4nu
kqY5u7oSVWN91GmV2NrKkFM2wgtu7coqfbRHfJEMsgwH/buq9DpSsuBBvRltiiAq
UQM5OpkSh8Ht+05rR4kFI5tVVxfWMMd4gz512TeeVNT89xGmy23e9d7xS/UCNEYS
w8E0QJJaK13PT/ds0ymkaSJwuUL0F45XUgvFQcLaYOypW5o9kk24RtIT6exxzQwz
0c+rcJuPPhltyvlTygHAnMNLCo+KDZz+QVERiVN5/AY9rRUgIERDWXgO2F/5tAf4
coGzkhWMdaDHRYFX08PVAplvfq5b9elQzJ1nQTPTcT1M0eGbraNngPv1DEI6qnPs
j4FpZkWPr0l6Q3en+AYXcn9dk5ZnWuYWFEMtbY7reQt3EkaKMk7koL1yTRlSjBP9
YzwmCatQVrmfdFFa/Al1uaeNPijjt0r+Sww9os76QWcCoslkOmxN3qbd+kXJ/VzC
JcEUV1uCvPOLijN5Qoj0gYikxY4BT2V0xeGJHGEOtn1zepVqE2XX2UfbeXcgwk6O
pkIWJv1UAv1wqK+prinTLOxri+iYBY0ABiZqTvg4DDWTUjqtwWVIqDQMwRGjPEWV
PoBwWRMxj5tHHAaf2/MdEThmSrg49fRSoGnMSjtdDH2St0Yb3sIA5/efRgl3rdDK
ExnEfcbkM3mvxB7NGGNHtPAUSvVQLGV0wdpD6hCSdylNU7ra0WR0ofjYuOBEqPGJ
ptP26NMvyrM4PkURVrOi0Wh8OU3fxzJATNFnmJ/GX3yCR+Ng7h8uluvIDUUqTwKo
seTRpWUa/9yl4xnPUVX3D3sB0qTYCrBR8Xw1mpnjhrJQ4TJaO6RJE3SR1Bt+FMzo
Hhr1+a3RDkA9oM8oAz/oOubEdO2x0ad/PEwyfDaCQZkvses881Bi5SutkPkL6qmr
zStLexA66zridx7bzvjtZZGdb+1xm/x3wInKBv0M7LkFgHzJSlSQwlS4xKuRkePv
XHL8iqAtGsIM1hUgVSb1avQuaRFqWvIYf83+y64xwrZtRtvyOc2IhWnu2Xq8buco
SjA2Vgs9ng5FYupuCo1TYSHxN6hSjRAxjnBGHtYOsKLXFuk78q7s6MHE7kXf4ZQF
8XI03MW8OTCdTwWlo+3c3n3QtCHOu6qqvOx+n+MsJbysYRcioJWj1NXcNs+QhtPo
tLC3DXTVOJFYFLgTCU4oNQSTYIMmIyePHBtKVu7xarOIlNKD11FO8gD8TL1y+WCr
vCfSCGNhy8OVMuAGTo3EJwK0Il52vNicwGo5Oh4wAgkC494eGIRChLyh8AzlJTCT
OTjnd6mHJx1n3C1ImxI6XHAUwznGSsJJEgWDYg0+IyMGzdoH6pgjoHIkIkjPWTWk
In3jUDX9e7lMdk7YP1CFqb6S8t+mkj/JVN1Iyrwziem+rvKkI4ck2cd74bfok+md
Bj8iCoUf2DJP4rLzJaX8sD3d05Dsdm3ul9kknrldtJVHeOrnRX2sFmlw+z13GJW+
k0iMzbccaVQ8l9e/tvdCG6c2MRXZYCMjyNZf3RxA2ooM/RufLkYkQNu7/g1z7lX5
xYbtGUGHeVZ9C2XwbdkDArUUdu0BJciMr85ORycsuPfOon10GBBg/2RCTw6Jqe4S
HElZCxGNSHu6QhfIkx5008BZmng1AG8vGkV2OEM8WIJ2OD1M/U/+YuDfgld/v9u0
10OdtX6Lx3p5fExqqALso+4KSoImCrQp1wsjJkKk7EeDQrmOVKWEhZq25Itiiphs
dXiIRyT08WCtETEviHaUIehjOyn0DZ9RgZFjaPJK6eN+bG1Ef/Eux0svzrKQ7fgk
TcvC3iOJ9JuDjZ5XNLVQVTvMQcEmjTSITNiw5UfE41zpksKCuinR5RIKMY4AakYy
fDBP/jBLe6nfOXBUEb6n2GPaAl5T0ep6u1KcBXBX0b0aH1GjqNq6PsQq+vipRnRE
S4nd/Xp8zyxACwLg0id8o3uDWduTYyWFbtELGA9tF25lBNvLJ0DRxHEycffig2Lt
1fF7sdef62XEUNBohVcXrUfUMMgdBCgr7Kzq/RoDelJL8T5zY1Jsdus/fpuAe2H9
HhAtUsjydr9JPpSDoNH5ghv0caPyhLfDPCMQV+P5pUugE8BDSuQh545QTKf4g2t5
S6gYOuLakI0Ty2YSkKE4kGpozAtePJmYsI4URrHLqxNLT1JXeGSLw4bR0CjHJCme
dGlul0qQam8QHsdHY3X8Kk7tjOwwrUWATpkm8f/VD8DIegglmvSzYrR0g72pQ+68
yKSfCAbNBKiWpzxr7r2LYNo3XReKZE+qHy37JESdC5nM0KXJlR/N4abK7VgypIV2
WAmPsA6jMLF+v7PhYTgD+e+Jjf1j9DYjzM5NopjTmoMJa40Wdza972yrgnvfvUSr
07cPXi/vlWuULDeLmK6TheH6PYvIi4V0SqalWeTGLonYxzkbED31XdLdWSk1N/hB
fvTujI1tS7w9sE02qBVI38dA/DxHProGKyIuha1pjGDeWr7zf57EOp8wxvmPTMgH
yLkavo5o3/fFSwBftHDhtA7EQ1QXe1JCONL7J8FuPrAYWgtcTUtqlkzFDVZJDie/
LFEJHKRe16/rGu7HXzsN753o7oCXtiRzeRxLM3o1bbiOIMHakb6aRPzGHq2PMsHU
5g6ihCBBhQHoqQUs5fs/BOU3wKZEd3MiL+rZVrGX6xkDEnG/5MfRsKy69uBceEXL
DraTmN/n/JdE4CiuQhSKfOAe5JFrx/MhqsudkGcEopFYlaz604bXhmo/zX5F+nU6
+IKf5cDh0HWaTOpyaI+2W3ejASDpJHiDBGI1AnCqtdpRRLgcpjLyXvu2IRZuOYUO
l0jrhyivljDIgEQUTF4lxotiotmKHkz4BNAOrZT8OY+1dT1aq5WsYzcdSxRjvlSe
FovPyQMOsmRFXRaO/xeaeObuLlgNMpAV2iyJTD7rKim7ZFj0M5Oryids+9mSzPRx
HxVMPHdDYgVM9kGAfviOY9fhCK7N7bIjvlKU9+bQxiQTiOPFqjjdAJ0jPDlCjVUF
/uUO3BjSR27Orm7qJ1L1M+zvQqoXKpj0Br2J71qLTtS5yww1C4Lig0Mmq97cb9fU
qLaubeiTnIxJ0ssEAu+5/+3qT12hZrciYZ46IkTt7egQpP9T6Q5Js8hXHrr1pRlj
IPl136dhYjcHnZf1CFBxdAqCqzpi3+XUH7GZBKqqwuFX25+Fx+JGs3sXky0pFYYS
CxEpCchErJTfobgp/mq2xZ8CjK4qPyd2hFBKOP4dWlSWGeDFwVeTGwI2isoFrgQ+
5/uIDyoxxvmneIvRdYsmBr9zWQQzLYqWwiSiHyvquK6uuSI2hxCgYt5vSRAnGaiM
DoEbBq++DMGQsBQajtvbo7xI5eqfHiTzDwRtMwOzg+2M7V4b4z3gX3okW5YTADvg
a0BBENHIFq9LK3U/vDiU5xLYJvLrMruoNMyh2rCmV1AvzCSvmRlIQ7WjzToMjv5c
lax8dB+r4nvFnDrxsPE+fSkv2b/VeYFNXRVo87dWJ8g+M42VSZcL1jQTSjGG11nM
dIiLM3jyuGV0Ojabtl9zEIXeNm00P6g+lc39QHFj4J24V3EBJWXSRUrWGZo3hcks
r06rkkZ19osz+idJC3INVWzWGusZRjvt4KLHLVCA6qqztki9J/EwuCc/ETY7lktP
ZK0xuuOEWmIFv8fL+GRWLm51X/fAmSRITXzC9p7VITeDlweDN4HFYGUUrnSCOg8e
Q6HVJUGAESTSQfT9qiSpdVIE7jwuJc+q7aAVNqaQSPjzm6fVvEYEMat4wkAMyA1Z
UgYv7P8txhaYqbffXOjG4CmkeNMmBqt9lozpSIWRqBgI4f3Lp0hKe2ru1Truug6b
pux26aNIfHKDiaVwdqaP7MY7kjGZjzYuRgneBJ+NvcXE4HGDT080ikZWrie44Imo
QmuWfgPtZcsg92+B3G+QTA9t70xwB55eRYu9NLsHFG6WkNYyhkYs67a5CCOtgf6z
pBICdfR4jlkW08vopAgvJy/AYZSGXMiQvHZutut7LyqbSm6QpugdXiMZ21QX482y
fR8BRfkgTpWvL4xpxBSkRvhpbHEAEqyfNrPrQEh/SSExXBKdh8kiQoeynsl7GFBv
kbu6P2Ff6rWPmJiCRq648Li/Yktw7hPxYf7gDRDvxCAKxJz19Ix93FkLvgmcQkap
CJT/3lwUG9BvRwNWiNpPR1V77vgkzFjk/SiFsp1sxuMyqVXJ4RUna8ebq/S1IOKA
mQY46QBWcXG8uAzV8C7gIS/SVdHHuialue3CCtqIELuN8XMwtR8V04LSqcrWKJDP
5MQnf//jC2Qa+Asa1IhvkLpIkXuPYdj1yicWfbjTib7XQcfeB9cY3ECM2j9YIowz
QYxLtvPpL2rGom5L2fA/yTWMVDE2+llethtOCgh4Af3SdRQliQNFQasQMrguHe7H
Ruj0Ib7WCOmlWwdN80t5/TMyfkWRQ/U5RjoqneiHPCi45H6UCrS6V4y5gLrhEVQB
aoTBh0oBVUIYkw+/SlNQBb4uIEKxS6MA/R8t5aLPPw1/+gDp4aMs2/gAYP3vQw2X
aggCXVwrBc3HLMH6q6ioYgdSGpizTbVp772Ytt8pnvDvYWRhtZ2OR/Cr+hkDwxdJ
cs+DAsJH/cSBw7p4rM8der6zr3ex6WU5abblXW1DEOB9P3naFn8Vc59ay0fLhnga
eqXRBw1q1lxPefyONT0GqXeX/dYXsQJqgN9YO9ATmY2mA2fDOBaQDShodLiLkPP4
atnS65+IDfuLk/mzood4Un2xoCLeUNkNTay+OppQ21qqWb5AiDblRJtS0dRlz5+A
3XBbW+xF+aQ4gMbCaIHF5NEK7I7q/5ItaLyF8MZ2uGbkI1jGAlDbeKpA8Ck6euQo
CJHlU5LFVQGHpE9Hlc4yf2U/vfjbLDt1eUku7kngWzZWuXbYSTsEjhfef9CxmYUE
PCj+m0GhZ0qxP/DW0dgxYSwUPsWBhugkWlGrdwFUiGIkM3Zr9KQg2UYXiUqSQcI7
IhT8Fg0Xml7OKnm5JUwkCwKHJ5JSrdv6XFrkehiWFbAuN+MNKCEe9NdVqdXK+CsA
j0bmVZqmFzEsJDcPuNs8jn/V0p7JcYG2d5/4WwGm0yKFt0rnvG0iavFVtXShUJpg
FxK/TC4AtAEyvXwipB1KxU4r7wHtBS79Y9dUnIf+IIqt0q1pM/M+CUTml9YepTj7
as7VX0Sl+56M9KAaimp1blQPSrnr9cA+wgjjRZ2SBT4Jpl+0iUzkhrjQV+xmxnUm
BD7mteANp5wLo7ON5BplFq5183OZMeqcIwt5ng1COL4tSpsbQD/XrLFET93h53lt
3jO5HA7XSxgcsTjy8nG9TupJSoE6gVZ6sZpyZvmjiysrFjmSurQJ2FF+HaZMvW7X
RQDitXd7xEkQ8Jmklqz16bq1XD558k0s7NQ8XCo4YEDNrk48J4Zl0DlpEFEVCMWq
fj7OPguPFp+sHwo/n/kdEZfaIg91+eN4Z6UsQKRBoa2COGWbyT+Ea2gg/7S2ACwO
MzVCix7CPuR4LrubwRDU+mjL6y29G+s8Dt8pJPgEowE9t51pD2wmpKvHVBmXWP+W
rLuOGnC0LSFJZfPuHTkSGI2RyvZiTMry2iaJcGc+2ldgR6AJN7XCtUUyGCLrWVI4
zgH+RB1MD8EoNpZezX2I62Ti1UNdTHkn5ah04xrdK3XAR6bq9uE2LCex9HxPdL6m
AUTEDzlFeZdrfUZs6Dgm5Mj0VLxee5zo910spTuXbm0UfFANEbrHT5wM1n9HL67H
lq9RCvyJbNLkqt3yjiPjx2aElJdFXfHQUY6rDT1N4wYMtrLTX2DsJpmG4rDhDQdN
XcI3mwKsVm/a2/rTqDSgNkHS/VbzMOy7zOfOu83tEogxdMUKZoMVcBCQS4e72tCK
6ctxygfxJQphksDN2J1jxOvLzH8eIM+kdtsq9o+gRZVMO1zzsmeKn1IOnt8Ucfz7
PV4KDZ5rGY728/0IqYg7LdRb8Hb+GsJkdZWeI6C2yOIy+uFagT4fews/mJ05nMmU
ey/qnBaIeCZ40WkPFVou8WVIqTEZdygKnSCeK+l8sA1Ca542zo3wD2pHmmMHssoY
QbWqCYj2CZFurhHCRlsspYJWEWPl1rUrJq6l2Pi28///G63xAyeY2xTeeeiIWihC
H/S3BLCmMgPQYsgkE7cTmc4PmUepynzypjS5s6mwTLTZl6iHIUXP9+K6MD53/qTd
7/FjG/SKn6kGqCU5Sjnw5DE/Shv0YnOz3O+W45IiHuHLOamrCRPZKXa6J+fW1sSe
dAp+ej3gSkZdXEP6DqG5HUTaIugUBFN3C2MenNg2WodcpI+NBPW9NDcouLSPT3zd
+HpS1lyRJ8GQIpjOLSToABbAMmSoLBhrOI4cvWgyqm915NBF6HGFVKt9D8obZbNu
FncGk9UOYxh31+1X1KW6GKBAYS+5dcZsKkdunbo+MGZwvvY++/0BVogb6czbP3wv
Tz9arPkFicOWMTmXalIqR4h5vxgYXapf1fs3EEAyqLuHafh7i6OD+QjW8j+JMAf7
jvxj3ZHKPPiFalBdkPwhS8Reb84KSPOOnFJiBhzLKuF9uygXxbGmhIvQqdpeLMt8
PYiF1Rj3nduMVecOqu7c4QV/LVfJp7Z38wMjY3X9yYgDvBoRWjkTF2tjfdwQwVst
oksVN6zKO1AzFUKhX8hcrKIID3JZUlB3mYI6db0au4+p7ndpcBxHIOMAakjPk5r+
e2yujmX7PGe+NEkp3b/Kjst7+QXtVcFbDgxY9WrWVWXz97VFmn1cQ2ox/Ed6r98U
RvjE3msC46nzni/zXOF5Hibup/Asu4cEDYmD9qi6EbHl0nbVydxCXrl1ykF5qchX
TnRHQ27lqN+oLscbrgToZqduXK9igRMEGJmBE1tz3GXAxdZYxG7cpoRIAGWNmPBL
h2pbKrlW3lEzw4w4HVCSpSvooYM82P4OxzNNeA67ZRxlw6lxbu4y+FTXAoNGInT9
qc7MMNXPiY1fcPyhqZTyHppfPtHtdPv4Eh5k28MHt/MavrBENzJ6LDYAPEdUOo6T
hqB0wy+F1tk4sa94+OIVj/kaNeRM08OxMlt7/sXN5FyEcI7tiCo8UeUjV8IWmHg/
sbmz87ygL4QGFe2d3VNc9UOlMLTxOGZmgRifb2GhuC3lXGiiAkXeAC5IGNl5/ydE
IwYNujqdKFm5iFXeFiHpDXm7z9HvT3Zr8bmi6wiqw0irKIyp2H5h1msNlw3CDbpP
vbkRaxk5w2L8c1BhSK1Ra5OWY6zbIpMYOLpvRLHjo9s0hdWs2sCz1CAnq0/rCOlU
B5aRs8uxwnGVTf+cxpd76ThsuI2w2HEqxYJUhVaGV7PBihl+2otDdUG2rXEJn6oi
/swSvpSutuu6S0tS1M3bih3OqjVICtZkPTmooVsMZfgRpGRo77Q9Y4uAIIgwY3R6
p221xBVUh5Teohm+JXqT0xPDcAfTInQxcjjcnSEih8Ps9W+k5K8xFKSMoa2w3znW
HnOm1EcC7qPF+CBaeWlbrwXfe0/3kHLwVwnw+XyoGDCmMYtzuVB8yQVGr1N/MZs9
UVlOF3v+Ykh+nGtkkc6rO+vplPxpViOyKMh+vbL41PPfXMILI9Xg/nouOtcLkoay
PodMhN42EujGmUYi/sfwrGPaaitEc9NfVaTZNYtjo4AEW66+fRX+ROmJkDOO1vcg
9hhV23ppch9XeyKl5Ram3Ziu6PflqOZaaQkp2RHVth+mAqUK3MOcJQxN0SxS+AQN
sXS0UN9rBlm/QRANbDozw31uNsWhTjFoWgS68E5bXr5hftUim2+kwQh7b0TdsA/N
aMjvGoNBHYUdsk17jiU/cGFw++wzD4Mw3oJeCRBFabzca/AcqvoHBL6JMxJr6g+N
LkeK+Vy0Iafojae/dfk4DQajXXTZ8/hddP7yGbhWHwMp4J/tGgRT6pX3O8QdaV6a
wzZpGUpczqpbTBiAeX7E/W6mey3wYivNVvQKFq41/pz3kG5FdWZCLyN/yAYt0mOd
IhbP99zL3C4j9iVO2iBAg8//7ISPnkSkJLV0MWTrHvTjkY1wZzsdioKJcghnCTW+
PRaovjSe6TnTahXwjG5x5xBN5XZUuO2JcncSWGXTuXMKIhHmiQ3wusBoNdX0odwJ
ZAtEFMv6T6y83gHPCq1dtkBEt0Q/1m+yTBxgCWUpHGyPRjIKNpBdGYzBt/0qOQxE
4tWVekvaWG93FerZ4C4O0PGtzBa0jTvCKNvKyH0K0UzbhxWC9sSie2srH73OcdrH
2/jjpLVmURZ4I0NOvIRrK3NbXiTR7AIPtiYAzyD0ukysfslNENJ4E4coV1tnQHXk
jRYBN+Nb40n7TN2nWc77TxvX6tC/u7fWZk3gjVegF8Ax3a2KW/HzvQbXyfqiJMMf
lMb/XtexgbhD/Bqi8c3ckx3lTrqf7WmOuya7n/LG+SfM1RZ7xoUh1ID0mlKSzN2x
jUEKPCPoUvNjA7mLdlt+7yBbEr3tbYJEa+s5wfPSmicf+6kqDQJnrSAtaFlRVFit
vtJ3pJG9GG3SFNkQjeLM+k9uAkIEAfj95JXxhsXP4XOQM8NtjijvHqBQOevWzylk
wivPXW3UruwcG9W9G9MZB+kJfEBaWOq6NqZiJfZXA354ry66ShG1l7sokcNyFl+g
yH9tJXrQWSSbW+ggR5bClHHkNxKFAD8arSMhSUWmzFmpJRwEGX7GlezSYhgIUELg
yAqz3Zez1neCjEIGcbbUMhOckv0UceDFwr4pofPRndL+9BM/wvHuoZjc1hodl0Ik
xPhnfKRAD/6sooi6Z2BcMbjHgWB0OoOs7OyPAbd3BNUe5HOSucxo7jRsritqMOsT
oqTyXH2kQ2eQa1iP2utoFetVkeNr9UuFUlY+VChqzTHYzs2nxZXS56iXH4eO/1bH
NkEXxloMvg796Jo252Vx27J+67uDQ5k1mFwixrwKNu5EiFBCrpZbL8dIszVGz07b
oL12GUHesSrOeyAru6J9xNUQDZzEjuXw4muWCFXGBdkEUtEGUZTV0Pi2aFMdREg1
PhCKUALotvq735Zws2DJPhb7UXMlNHO7Hq2J4CYI7y+5pptKh4xzOhbqO7VsYx+L
+gQHi1pCAU/wJM2e1puHL9WaSgnHAROS46RwRTd4iCDCn2vuRR2N031TmuhDTVoT
cTwQsimY0K6/LaI2Vz4PEVAass5OJjf6e4qo4O565djzdOJj5nSOmQVNbyRm8DeT
iYWvwx604tkOe7YKQWE+sysC1T608/oS8Ap1A5w8lPCrLZAR0qa8A33JMBrTA6ua
m/o1bAHRXs/6J9DOnB2y1hMrJ0JqhcQ2LhOxuhJanOk/Tg2yHSetGEIN3QbrdGjR
YVRojtFygHEUAXr7eIhWG4sCHXhxfezIZvwWNtuCXBA7TbWpdsojDpWgTeKAf86k
OCEJB1u29lcvOiBFDSG8wTfSZ9NsNqMHhNKSDKNB7elZvDJqOpxW/qok4I9oi1ag
b7VKMkpKUlcaTezLbRZjvshBuJKasn7wZbcDvKPwpgp7w8rBQ4ehRipBQhHEerUn
ZTX0bkC6cbyS7N9m+Bi6Rqf7Jnu+5dosAnCtD7267rijb5TIih/6Sgj7Y6xMHjJu
0orOqLzKzewuYENHcobOrF2qXHHasWOFbxQZZEyw5LUWCsvs/kwCGYu7X1FzbH0+
QMLP/twrIZ9fto8vQCa/NvW7lgxk6uFiEy0IGCs+kKXhMkPtLPctCYv93I/vKedx
Olukhxn+txh2ExaE2HwcP8S8OlHj03maDrsXwj6kAi3Q4ukTAlkfAnBFNnO3RM5g
RV5bTYsd8WhDcoCK7RDE5zXYkEQ2xuVsM9QQxToAzz1Npu3nOEkjx3u1x3zCp4+j
xH2s2DsuD1mklyyRPFuMN+OSDiMDvU6PRSN6QfpcTpxi5UzXbohBHkEyYA6D+2yX
gTvG9+pXOO0U5NaFMdBDVFl7urzdq/tRg9pbyjADq1IlCAepy484ZA/z/rqkwRvk
bhoPFycfPP0q0ahXjcSB9LnNpq2CPmxZxj3P7hlv8Bvb9YdcWb5esXbX8L+ZP2pV
jFNJCGkE00ti3WFkpTgXY2rd1pwOKOwiA4Xo9S0AmT0FcVF1luucIQRq6R8ddV6X
LkTNFHL9MWqaTsZPYEZfYtIVcaY/zm/jipk89URhrVZaNTg7lLATq5u1AHzKv2IH
93RPAswANNFwzi9YC8XeN03w0SJhZUoPUAnJJZSYKu2ZOTEmgaL3ZVzFL+TbTv5d
5pNVK48rsUpva34hkybFvOn3Wvjy+TkyAIuPAB2RWHMrEwmEcDmTWLt+scEoiKgI
wtfgOOHlEXs5j0o1P9hbu9AyroHnI38Wo4B8hJdlNZbngDNBslZjuTTKitEeUAhn
B+qW4Zj0CjN7iR5+RTuYMn3R3eX0yEkEt7atUKk45VKlcuATt6FhmHRp16ZTnRSj
alrMH3hJL1lHdWYlZN/THLuKpU0jlpL/KMHBpLCBSFoOMA9UAY+x9w6hL7zWBLSC
FjHQwA3cAHiHP9KwHQYMqbmhqL/2uppPw+RfyPGvz+yaIbama/i8SvQCNCaejdZg
Ys33d47ktdgiI+fAESJvY5dD97l/VeoAjT22lWQacidpc0fyzOQ/Y8o4nARpc7NA
6TyIc0jxZH48RyfMXnLpDSyGFyEA5GOItG/c8GEfq/9ncbaVmkDqoLvEjWMQDbDn
JI+/rZuNJjsjw2syfQR1jkSbrd4tNrJdIJykcRbvTLS8yb5Wd8te7H2FgIAJMliz
JGQtCT3I36BntRLliGhiKe+TBAo3iniJUnziaA8M/B4Vx/N6yhwDEQ1762dI5p8+
vlXW/2pizU7yoBHXMTXhwQFcIgHkLgy8jTwUOOLn26MvYwDEHJdkmSYuu/ySBQ0R
ly9Ao9JndwZGCC/qlKRNL1yLaskfwm27Ee3oZx1A2QrmpunfRWKaPB2WagjE4Jtj
VOTPIAbYOsvkG0xsKlIurmv66uApOvLelx23h7l2Xkgtw0Z4IeVtmhB4aKn6OVpP
F3v6wBM+yu8CPBvnek5hQzg+jIZbSrh6iHsna2msl8QYbpz4IKWfZE5W7QtqFS6N
JKm1von7G7fKaCOCZ3S1/sgv1cTszPGa9fj+4yYSJMGrvti34/fnVIUjwFYB7MKt
h3L9IPg1a1XWJh91fF1wBNFAO/ohJae7Z4V6Yu+1aDiAqtxBcHgqPExOAlb8tsCq
I4BGzT99xvR99GwFt2Bew+yv698JXSzsjRc/nKTQQQmn7qvoKpgqUgAqk1JODpz/
2Wujf03WSyWyjiNexD3kr5eAWoaK8qTi+CFEo6eCpby6nSGj5VCc9wmSpCIS0dd8
6qt3FqbYfmtMbBFCJNIvaFPD3q522FCS2jtrdCceyFsgzHvoL4hWmkfM2xMxpYOS
Mp7ks+cf3XJUbKB5s2b9dBONzZrj0v0TDewXzrV3SypIspb5WhOV51ViWwW1qORO
3mgPmpykG8qMky40xxT/BkBNAhInDIbBXMGzKxlTSeTt2xNIgy7LgdBP4kksU0Ru
mqTTbj1VEV+phWMgoVDcxMxbJlSM/P+zEbn52kc1bwTZV/XRG/ZNMEJzBy/nuAsE
tUvZ5dBt6mCM8Ro/q+IEuWCeCP7rPn9WNXlSgBSSMZOCHK4c/sflF3WH2uaLxHxl
AorW0jyIyaVJQJjqcMatsVRPmCgXTsSjpROBpDxSpFKxmY+jwU6xvMknI6FKbNrQ
ctl/NPjjg2YNm4eZUPrlBvulXlwfBJyT52fcE9MGcv42zFI07J1ayvqftTCVubZU
T+EhNp6fYF9zIITxmz5m7X5C8tni2PwtTfmc36ma8D9U+8geYm5TLn1vqLoOLMD3
hUJ6JktSlD0MmfTHw6wT2Em5+MoD+mBRJdiJkOL7gYBF3IXxuPWRufvXfceoHSYw
zeIc5bHzxsfBzbxSQVnEycBWsjvi/9rMgJ69V3S8Fsj1G4nhWV1/hRPhhj0tm/9C
n04tEDYkylBPj2dn1CbvH2Ank30SgHGBERIpg2DKBzE6BQOlpjUGdMIF5hx22GU/
sVCuRIImXk28ZsWY2cw8CYbvoXy7ifL7Gd0SJTX9eVTqJK8e4WWCDEHm9mf1Ch2f
vb0SuID3IKzkQg/hAPnAL2LV7iFHx7PVtBtpWe5mOUH/OnQHm8VJlTvoN8hhDHvP
bpHippcetEsbN2NMdP/B9cMBpc9WxAll4SiTg8uUIN9ywppQ4hVgDAoMj6CBTIe+
LtEPQlxmb7LRLYvfFWBmxDD3xK+ULW1qBRmM5ITnokxAXFDMv8kjgpasgPSFmzmD
XtBDbpUdsbeXr/VNubAj5hW6u9XleTsCeMlXpG4TJXSZN5FXKINjZ2esoY7KaKZ1
9kfONdNeJ0zA454+6MJ2a3MeqRHFrmwTnvdHlxmzzvSLIS52rfktZHIIdRgRxBtg
u5BU9N/Q3aINWA2Ui0vbbGG6sy0jHipOV8mQY+sB1EzjaF4McUDh7AkRdphEOKGU
X8zfN2CGNEDQnIeF6PyhdRYrjZLDQLMWZPrNTI6pgQWMWk4NHOcEWb01ozWUbIni
upyqRcKEPT2Q3HfzeNgmNAWfj8bC1Fftn/xZMxyH+ZmREw+S3p3yR+vumtmNix0R
GqNc2dNyjHNV9XpJC+O7kPMOJtHGD8G39THFJfB3M4cX0mxLtBhxIHQ+rJuE4luW
6vbILg9op49TcOy5JdB+XyBg2g9cSJnB3Mc7heB0ObNGTsaySqxkUVoX0DjRk0MX
LTn8o0KiHZ4csWjxN8PFMJCC19gXvydLjWjRFT4gWyYvtNjKcH7Y7L9IvZvlycya
9Jod+XYaQlG/LdukLNHLUZA7g9TkLhIHopJiiJlq0iclG9UxecGtyl9M3+RJQBIc
72WTEziLV587rQ9XotvqZPCW8z99v1G2Q+QHCiOVa3d3L0bshGUs2QTAR3BA/AJ0
f2GCFq0pn7Ed40fLr+Y4QBGdMyvbI+vgrSALviNrcOwwD04iaQMJH3Yn6WpkIDUd
60O5yU3BkRcVgEIJiFvrpAkczElv9qIiWDaJVGj7xSeyNGGR5IhnD3T4XT7G7Hfv
wKfBEJy8f6plN7SEKlcTa940C1vnDsl4PB1Se4uI33lXkk18r/sv/G/xgJjBacoT
iB/kQwgFr6xniPMi2sdITsQocEm2fliiWKQwpF+GhlSYjsKbpPIc25BTrsK/5WLX
Xg31kagJgLG87GnllXwGRnsNHXfjvTu6VrMvQl6JKvchdNEY6PCzgCoX1IVs8TeN
7Nwl869Ohtg1EZ06NcDhXXIrJ9ZKoo6ZtZqO2+ocpPShznDkRf5TRepnzzk0ILVp
muWe021MJg/6HMPp57Oct47fith/hIoxUV98kQO3KT7k+Y5sN8Ol7/s1FbRmr4y3
n7vnqaXG3aheorEq6tJuhyLwQ4sGBOiKHQTLMI0H4DVxzhLhoEKNTzpe+4PzHJgc
DsA0GWHs3dr3ZG9UtN5S0N6etjMTLmAZ3CNLm0ri6ryfWcCxXvbXFeQFkufFTda6
N5y/ksJKQDbV+ukXIjH99R9N/4TCO8LoHxpV2xGfKEK9Cf8E5fozNWdeat/UaRGp
iTQiInbCSbwJeFY8VTPN241eq42dWW2Q1N0J1o2gei25zAmFd4msyDwG+222+49Q
cJfvc91M2VdUPVMnD0AkwUWjrRIrRnx+liH4zADX7xWKjCnEsQo/5Xx9FzU95lhp
AShVDHT5rtNum/lM0RsmwyJnAi51rWqTgprjHfpA5G0Ut/eBSyUa61cCz1wehgIG
8oGNAw086JLZZ/HpZ2BmyQPOHHySSighz9HbOwTOGV9RLcjPcmzu67mgu5/IDZMK
TgoJwZtVMi/HueLMDXPv73iQXr6R6IxSKrgI8e9M7LXn0A5uN2n7f02sCpQqQ2nZ
caR1G8Rh7xa8Sh9ilO6mg0k3GVhCdLJrrcSVKaAfrTZSUkw1CBBJgnE2XJ7LJE7g
uhapqCqcuWm0E0LZm8H3M7Vb3fLoFDS9/WSMKcCV69eVZkZJDqd0VL61QmupZPB3
egfcvvodGWoEUcOpsdZTlIDeFXfz+sRluk7cDcz34Tl7Xc8Upy/Hb6t0nN7rVh3G
i9PgcX4b4S/Nx4o7FE8oF/CdY7cm3IRcBfoIFQ23kzV0dytJRTswe53FnfqipClZ
khAYNJkQGRMwze1ulXo1mgtgMytmsEj49TRyYl4iY61lMVjkyatEN1iE76DQw3id
30DG6IA2z5IeNMJegBHkurA1euw3nPQVl/7C6syOdVZknD76ac78OrylTciR0v/W
AdfZ6w+tnKKo6Un+Y+HZJZ/mLLFGGG/m5481uHjY8n3bpFHAQhc7T1otoZogB2Vv
pVJepoIKE0THkmywOr/1MTaAIJEbJs1KPVYsRno3VhkVDqnZgXJ4f1oTOvNt8SSr
7Jp7VJYqo3jOLxiRFoyXP9bZchX9Fdry+uA0oYt7n+CHnu0uI229yb9e3869mib2
vjHQPFW2ChwdWVf0pEkapXw5RNPWlZ8dFMJbw1/qLNItX677vpVvPpGoLbU8T/Ca
rquGtCPUuLA2/WfWVeT1LTehCRsKaDkB38gcv6NuxMsP2s440pT50v9/aSwsNdvt
/lgN7GEwT2kW33scd/JeqAhYnMDe4rIkVW214btMaV0Hd0GWB+0R3wP4lfEKNlpI
TBICw04WMRYVcB9oU3l0g2hq385Jgz5szn59j06dJlvhshRjV1lPLHRy5TzrK0UL
70Yj3wUUgO2IQsCyOMLbiLouaVDqLUrp/3fd3ctw59KBeDDikygOh/6Lnk6MEbaV
n8wCo7DBPjV2GAVXzr6W+aJv5xTdn01yCOi5ikoYeYn8tZxDkmIRd2DPFW7RSslX
5wzlc/bhOxEmiKX0WtXK8mEvhC26VD2gbyyK5h/1etcjfOeOx12mtHbPJDoAmDsG
oQKdg4dw1syLUUoV/WnaqtZ7m0uZwGIrtZFmJN1EXJCqPHkmqy6G5Xj5Sspgl2A2
OCUiW+9jOHLPm1WcibVlBCJYGJE63xZwF3t6S9hF55GtN/nW/kRCGdpT2z9lbVMl
xvGugZZlmNO8MZBSPAKGdXb0iaW94hvoxUowFQhlBsuE6zzDxC7G+c5dPT05tSgk
HVDTvs2FXJP2nJs9V5WO5ijxkPVjSktwzJdpeyLRPhBqGmxt16ZVOSUJ+REZU12t
c7nyYoQl12kJMuyR4CCSBzycOPd+2wevglTwgrRMC/qrmdGpNh9Hb9U6v7drUG45
h0LH1X5nrhucUzB5J88LBXzYIigXJSL867zbMyrQ73ZVwXb+usFKbFrSZ2mYKSwL
BO64WehFBiyRvUouqnwRPCqJXVKBsAiZoPHxEvLgXkVjgLYOA6Sc22qlU1/aJlXw
OkKfnbtbf+6QonQDi60UzL1rQvTYwvMnbzexbFUYqsakE+C4TaHvcYmMq1dkRG7N
B7sgwucwwZzXsfCSj1N8Elf4KqxLWlv5Ej1gPLSbMCKHPKnMrLgaFIbchZXGfHXj
t+YWByrYopAbWbIQfZZ/iOuh2ewqBjoiVqrJ/KjajsKtBJ9+pMEK8ovT2ThFjAPQ
ZbV3fpeB6KvKVaET3NpZ2v1zSVNKZ6l4ZweVAqA7DHiukNYwgPBD9cTfVgwkQICT
/B4EdIIHYtIz0SB/sZatXEDYzjQwnrdcY+LwvC6VOm6lJPnfP8f5tpCPwjchMkFJ
nrH3xrlZvU3/RvUwurGoFQlAKu2JLwQ1n9xhVu64bh7WaFA2Af8uDgcJl7ul+XJb
4Wszq6waqXC9bH8/PSI9aE4aoUZj05VYtoMHdB/liEsLGjl4EON68euvZrvS0b2R
22f7Gcfn6HiafXrlR4bMWH8b/Gi9RtNfU97I0cUrDWnY6g5YgOKb2rj3ToAgP1NW
72VmlZ3HNCBLeTjmC7IO+5rezYgpJiLXZV0/IuGXJZ6eRifV7fD58jfAxJGWARaI
xGstkI43X36RC24H2OiGAQZsLIOSNyoxTQe5rr/zDNKIRycL8bglUl62dg8+gcp1
ZjWrips4a+e9Sc+sYAhIynUeaevcyFuarnTWjsgEaAQoFQvCOSZtdY0bLSphFvYh
83mQLCY1wNmzovUpKpg6JTI2fq59dhjNGPs0vAAAkrQw+SPNxxn2yL6n5MT8FrZA
cGLGeIPOL9DfiaWcaKX0xOJ0kaDnZqEfYm0WjCtCZ9bUZxF5uPsI6W/aUtlhsbti
WiI9mJyBiNeVhEx22OZvVaCVt1OBnVmh/gepV03fKnkOhnrYdr0uzEV+eIJgIvXO
f/jhvzRE+/D+/PC2PFWAF2xmndc/ioy5Bx89W2m2BxqduUe6+1t4kJyXtzssyFTZ
mrWi1h7FjWv1A48aL93Re8eRDH1XaAMFopJiwJBTxdvcFv60t3ov+KyquWyDUKIH
/n+tso3ONbK7h70T0ShFSoJmysB619qY0t6Mm2m5YvhUnIiLryCRKJdK0ptbmki2
1buJyy8ypRHLTCia5nRR3mqfVgQrqoTi39Ho6H9nGJRQp++txBMLAaXFt7yrk6CG
7S74nnnYimapZkPKNzWa6xqRhtSxjgnNj73aI2i354p+dZTG6nAuO3Za9QyeFnE4
y03bRHhVT8UG2Mp1PB1yM/rFpn2kalVVs/ERtHj4l94j4ocmaEO51XCnN+NjlrEz
sp+x9NW3dRLOXFMoWWhagw0/74MPImX3G26o/RQNI/0fXhV9swTn71err/mhHuKx
zWfihgGm/tj2Z12IIXVNIRirhcxOoeR4lkNaf3l97OXB5X2kLKw07aI8ehdNttLl
NWTQfexXxUhdLCRx9m9n5mPSVcZISq03l+VrFkCT1JOo9eTxIzmMWx1LdD7fS29F
b9csImJ7Ycugi44xz71CapSr5Bwhz6Mk3SPPwmgGd7orgYKpBUJ0dPzX24FrHHR1
if+dfy8WYrM7oxKq+NnJKdq2qKASXZQ060JKUtSWb5cM7pzWtwxE7KBTa70jm1xC
Pc27VFSzEOTk4ek3A73q5kMlc+2Rh0UdwzhO1nJhtzFPZhiU+yCnPYU5HDtXMRny
/AnKuZ1zFqKmYp+f2NT5OpJ1U4sI8xwwm+SUuzLgYlSZqqanXCoYsfm0on2Mjc1a
9f9BkcnR6bjtgz/RMLVAwgwyfDtd1kebxr1E8Yr5KAgDv8DYsqlGJEsE5jdV8I+q
/JDQoBKspQjZAGFgN5yE8RsYDGIT/7GWqrzzLafp+GSACJ8V8Wb+vyofeBtxMB9e
/D5D/QoMpQ4Q7fTMZEwPXHJIhKZiAdZp7rcBadzOkJwa3Aj7KrwHJEPBsRevHXbW
4hGiUIQfVK+uBzmBXTVrfDpr85YEXUTDBJzyl3H7q7arWRcIR7oT0NBxcvIpf5zb
8M7rPZTyQFse4hjsdSRPB4IN4GvJjzdfV7H4+STfNq2+qYEjV07Gv72e60gjA39x
YKGWFfB1QI8wxBSv3hVQIaw3BARWjXRshlPvGjlMhwE+KMbckK0UmCkxkfChGV9J
XQSOjCXBZoz/72hYRpukqKxMFGoc5yeWhE7ruu3THijTt01t2b5fZ+zmIDt2tB/f
tRQGB8uFcAzs/f0qIx9cr6vmMszJwE9kcBH1JEi5ep854yDCq4OPnkmKbVEhlQg0
21ovJNmUM9My5qcJwu1eUyfZTxZl6TaZ5vZT55pnTD2ScYgYujhmiwXotf5MCO2R
t1A6SPnbn2GkL52NEG/qXF+lwy6yzb9ZOwz2Ow7rSnPU4xqNp/W9apWBOP0+FKZF
9X9Q9YprPNzqGPLTfQgIA4+vuu4y0pHkkWV/DEYQ/Fve3kkf2DFx4dWD3DL+co+5
xehXlHSDuI2pDjZ2ynfn7UeauI1J8gVrNrPm29Lx9DJDRwV7F+cRxVwe0sHd/577
mClVe6CZ11lzV2rTDYaPDEe+F6MgFN8SVUMyZrSt3sqq3l9mzjkqsTs9eoTWB6SJ
J4U+3STUaIySEFJFcOBDlfUIrQSQmaF+8BwO6vhI3mrg2qDRWPn5SG5X1Q8MzLDk
nUrXBTPGa6a5h0FoxN97IEAWCBy+5a0X1QZsRZn4HWvrTpInEmSz5o4lk8ivDihR
v9Qb6ztI6TZqKzJt91xESRTtqQNMF7cCgJIk0vMPe7L12uMtEqQnUlKtYO45C3ia
U2WLGOWM9ZiqA7nB8tE32pfzivkebGVCcA9aXwAMepy8LMDbMgYIowuepOFX6hIt
yu2Mc5bDmgI916dM+SdOkCibzeSxdlw5gpltF/grJaZL/GL/ypA78pMb9kGWOmdI
Mnejjhp+xO+/5JCg9syZ26CxC7oBbNbFZ3yFtKubZwrkcoLcdECFfnlSl9HWmTDn
QCwoytBCAYbBAgkrH9ceH+FHNxFDCzT7s4cBKJ+R0m07i8EMYTKVx/4jPNtTGFf5
Of/b9FTO8/FN5SSKiOCH4jnvv9lEs2YdFLlAF0MRVYsIEPd+LOzpixyC95teEcys
h4SVuiSdLJifZf3BJGy7cWanNfnkwRIhiveb4TReedYFmvG/IZACj3PIR1QK7F18
JVy0ovSwc9Yyi++Vb56ma0W5NG/9RtWPkLK/mNtfrzKKmxdcmq0fs+YQ9FOXi+h8
mq8umpMa9LyH7zMr4vF8SiOkQ3T7s/c0OmVeofPKCalOi9IB0JsSs74p9rkJL8U9
9zeouc17TdOV3CjteG+RRzx/UWHRi55Rb/CpBJgPoabpqLtSo/J7KM7uZmbvo8ta
rWkVuCDWsW2euogNy0SiimYPYxEPTE4AmgD4+oNXwJhTzyggGWvRp2b3uenCLi4u
fT3KOMGpn8HTnxKfr73wGrAiUExiu5AWpBzM8B3S48L5MUrm1AnOhTjTvNJsVvi1
85r2lxQ3yO4ASwfzVD7oNEkDQlMTlcqBeNKqdL93bdJmhCw/nS/jAvPtAMp1idp/
yBhNt7Ue86xK0qsX+Z/RviIBYaUZpRs48utCsNfhgwJ07Dqct5YuMrWC/LMip2Kq
TVQlJtMqrrxvgw1lB5k565V6IFUJ1veGpQovJIa3cQh3vJK5/Wo/XG1BWGcV2pI1
t0YYzFxNp8JtcIDiYPMluUyK9gOaxeLcJXohAzvtPVG9MMLL4qpl+IBrsVsJS9lq
wQ9mXgv9opbSrNZzMb/pRfF+BH6QK6zVyC94iJvDjkSv4Ejl/Ip8ACxFsFOXfaOf
SLB1pa7yqJYHfv4kHgbZ4LAGaY5zD9Ien9FnHINcuXLdwwmwHxaTPEDps3L/5/ql
PomUcR/Wo0DtcM4M/5L2BPUT0zFPlBguC4nMERFxpCv5lMITa/CZ6+mDi2HA3FhC
JcQFL/XH+sQ8z17weWPFb4OyErbdpIPyt7R9HfhlAahGbV94YnwNHk9zdNo4Bb3k
aTTwfc5JSm7n5b8Q2lwaxXIPeCmBOvIHW9yBV2df23zKEKtyIVOUjodconFUJr04
yg+AqO1ulA3rcfrqnKQEthi0INaRRwk+602+bEG0aRa6AmGpQWsXq44ROWxHB0tQ
G4mXPlmkQiN5f4L4EyYWDtLUSl6LJ5WbY7npl3upw4GI/FF3deWsvIZ6awcIqahZ
IYZYH9Ja1ZUn9hNAsXi6Wyi6PqOHmzx2FauIWtuYJCIJJDvjEJlVhVrsoJgsEkjr
F1hBwAqTeqUuuqidudpnJYZ10pqQxDNLky6AfwzqZkzZVXJubGDOD5f0rwa5V+IN
T4XWjW2YzVTN7/v8c+nG4VuJcorcUCWZyj5bgW3IA0ktcEsNbFTpX7AkAVtIsP4A
ykI31cSijMrJ+Zus0Rd42x9t8toTvOAknyjQXkIDQxYRetIPl3iJ1/W7rqhyq0/F
3CvM0hSgG7aLKfB2JnZP8/G06Nylaj3bis7sNm3BWddroP/N1JzY9d/LkloOH/bI
+vE843At+JzS9Nuu4ZQ4osewFBHi5CcARUPCCIptobXR1ZRgOdt216S07i8QmCZC
ByY+iUGC8sdsRwI950JrDzlEmiwd+j1clvZgyRQloHoPUWqnCXqrz/D78u3JX6U+
3+Vk4MNZJ1cdkWMjDL0BBLZB5btsahoIEa0PaPOCdwcjkfLwijBLAaio6/2W0E0b
tsTUPlFDpBqR0wiGNGHZgyy5DegyPa9GcruTAafrrjgSwBo5nn6us3KApFE3VQFC
bOJZEXsNNRJQxt8YS+sdyDTm8laguXdf0ox/HsQr3jVPv2Iuq/R7/fZoF2CG9MAV
jKz3UQvPl1m54g0JE6knmlIH3Yc22kYY9BH4ng06Uq28ic+0Xi7oF5nd8Mw9Jrl7
NAOSECh9MYjEUbb/28VFRp4a09TCHRux6bAgU0Lj6eGoxDr3TNjuHB2ox/T2zHhK
hNT1tuoIClp/zWpcsAmAQfFbYIP8huYk/KKqfg1VoPBncQJqCPWYLIdbfdTIiLaI
h8ES3jtV/+WjqyR08bfJUv6Cm1Qic/Xy/ggCGxUwza54caGJ7ytsjj3FYQAzmcfb
wkw4NZ9+HfBFQcC++SMRXQtbpFIxWeEAomn4mw7Xq2yQ5IESRa82TwRR17zPGxP1
wfcHzeoqypxopYf5iXjzpVEhHnAq5Vuc6/ao4LPKUVm1Bf1x638i59Lt9G5pttym
vSUErjZ78fc/QuMjWgU/ziOOt1eO7GYvAxA5XDNhVr2dmZ+UWNiAI9gCAwvLd+uG
AeqkVAC4e0aLtMRMzcpLXlJUb5/7VAr9zWWYy52hSacLkfprnLHoBXd6ArKpUjq9
NDMYyCqUpX8nfwkPgt/ZHjbdgPQkwUqvfL8TyuM/sqbk1RiMGfbq/hAW0FaCyNev
oo143H1czDN1lYmtlSo7uBvaSaWgWnF0bAe0SHG54AvPRemj4pMofZHBBvCv5oR7
xXxOi0QkZ+C54n/AZx9hrmgz83GhB3uukVi4GvORHNWLSiXM6xYqCfceitUoqFK+
duBs7lMJ4IRBbEStOeEjtr8Z+7aPZV4bzYMU1MpoVtIQtCmgUErZyk1XDW4hV1zU
6E2GKZ8fEILxrGyrWIrH696zAHPcSRBgDGev39ExGfUvhsxB/kcbxdq9Ut9YwQKm
gi92NQjU4F4i8PyTKRriLLYCv7xD5QjdoXDCSPYrjlgiMlS2mmxUXV8+Sib4hZYH
dQR+Y+/CJM0aGBOjTDwrSCYXxJgUHsqpcvhaY8OsObjIsCVHUomvm0hPmG4qIhSg
AscBN+wCsgAkogoI9VnuYGItQvjTO8ks71VE616GmfRaSc5zrSezC9F4E52hsbHN
OArBbQJF8XSCeCP2wrjuthOQX6tWyjaXF4HnqnC3TvKuL0+knmvglv8Bq7hkbtki
x+PMV+1MPsctM5ELY4IxSa5sBZR4oOrEKdEtnI2b5TiYBlwOL6bp0gxAELYniwJv
aT8yJPKtNZS9nMigezP9liamCioSvhgHrGR/VAZ20artofSTrZXXZ+T/T89h25n3
meOoXD18S5s2uFn1h+rfa24hgpsL+yDgf/Ou9jZkeu/vB3vCu804+Vrbfnnhoxtc
4KlrCYQFJlIaLYElMvU9R1++zzBzw0l4BLheQYGM96Q48i+Eek63KOf3qO+fOrK9
JXm8GxQ3LmgwtGXr/5Vsky012oLyD/+MjfJIdxtMhX2zzV/kvkyQZr3gOmCptVIn
yNA+LbN6u72KwtydB4jq63ZWd0+VGt93uj9mChfyGjURHJ7+cQQOf6cknWzb0T5W
90arMEw63/yLdNAlU4x60B36D0HHfb1lB7f93yovRWyt0sWlbA+kthHQ6jq1Wc/u
pXvsPPKTwI0mc8QTkwEnjymcsLJPHdWG2SMcQiMLwSohoDA7ApwZM0lx3WvWGmN6
RUsWpLEt5AFfVrOXfMG52Czf0POkgJeUxlXhSnwsyjUAO+RD8WMCRYYyza+W/Shq
QRxvRD4/A3t7uW9WSFYhdMKSzaTUlju32FMjBxuIgSIvmSYe5kfS5hFHrxeTZYtj
ioa0Kh1YKRuREf/O8ZjC/VppXuuss3qLnSpiCsbF2AIO8JMkflCjI9XRRfO1bJWO
jFkr02wpsG10wdTOmaOfXNSxavs9sluTR/5+s19+12wEEcvBgDUXBTRpAVD28AhZ
93RqBvhVxrxbd71BtUgAwE2Gnl2bectLjHbKJE0PfAPrHRydDoTxGbU6RJiWBuGX
RnUZPlaCooRD31TH4UX1U1hB0sQiQmpfodxU+OqvtGc9THLPLv2jQlnKOLmUECdp
hmX6ra8exUyzwI6hDGI5nF44lAXnXPobbebfeOItaYQeHp0PvyAsX+wpp+Axu3qP
RLMbqbt3Ucpl/Rkgr75Z2Y8DqJIB6uLaIQ54RyiGd4EIDnti8Rm/WcekMxBnaOPx
mketHw3eo/5tLAN+3iDMtsEKyaEaLsGk4o1e7wT/t+hq/zvSnXDNd3K5L2tCP79q
KjoIhRZici8sXT7JChnfS4iyd7UeOwzisJzHGdw/83CTMM1CacC3Zht3kWIGjL1x
5TkDIb2Ie7RLZ7ay9LwtqJCasI4LUuRsch3K8+sSD+0CRJaFmbMrmmS+gDzKM+G1
6PafHlXXrmQzUOeeRD1gqKzJ40uaLNq5bZ9u+dL8YRi3Y6A1KU9zssr2AeDnEaTF
uWXmfUr0i8C4hygo2L6ScjEhbu7pV/JiXjdusoFvzViRMaMuBdSxzG4EHkJBta0r
kJ4t8uNIjd1hJ9ZA7Yzi9MZAVQHaARL/IrC4uI+a0vcMQhTsRn6xsN674EzQT7Tl
467AIQVRbrT2oZr+PfQbOOX/4glrrgWVebdCd0EfYO8EVzG9Pyy6Zy22gU0B1pqW
sdWvbt53pWEnsHSFV5g8DXws6yuvIwWRbuDYXihstijKZ7N2BF94d94navsAGWoP
vmd9QjZ6ZSHEd8UVR6gHfttn+fRkXo4fhj+HLcGUb4dPw+gWuFoHvN89G0pykSD1
+o/43o6v8fFsUu2Qhg79e6uGRmDr0ka4NdBFsGhlnAjKrfr1uUsJNbZbsGHVYIcK
YIj9KuHh3p9vps7WK8lomNodDqfZmtXJnzdvSBx2KniGutG7G+pMjEqOaSUaRanA
XkaSAqKYH8ZwCgM6caKESmQ1k+YhK90IDGnBYR6JxPo9Vh/HRjVMafNOlX5kLOPg
zrB152gTUAGk6e0TRpIFlQXHfPoqMKDWHL0yXAgLeCfFWZBjXZs/yrBodzTzDXVs
j8oU1lLlONenwzm1pDV/F65vm5A/6e0c7aq2XnwShFZN30jAE7aV2r+3iK52hxPU
DJwqhiEl7mc9q3Z9v0pSghOrfvWCbvcxCvx1JRkrQr2JnFlQz2v1CDUFqEkqXoEc
f8/kGH/a2ynMfj9139HVrp8hh/vA35bL4+klimSfdfTehF5ppgVmuOitvko6aP2v
phCiDJrSdfgppSvb1lwD5JBbBFEtQsj/m3fkRYWlrq0mZ+CqZn1dsUUWUd+6cgSF
S2Zr3yZAi7TLhTbPrm/2hDVyN/HE09xsQ5buc56r8O/1hvs1ml1kgHbhBzs6Irmj
16smN9Kvwzpy5Rd+cvvnlEZL6ZLhtCzIvbFYnZolQN+uLGN4d0YgvilNTiblxS/U
TNfX++NZWqBsq14dWDiQgMiNN5o4zVOxLPk3PPPmvv3odGKjkRasBGurpe6M3I/9
+/IICgFmf6gA7cMbQIpQjf+9f/wj8OJEHL6uxTZXdH1oz1iwBA6ZlDLOnDW9f7Ro
vNkezCawyaE6I81/y2ZuxCo1WsnNjvP59gWZeFY8vaa461GjZFawxsV2I9FTw9Ij
GiOrNUwjtl1j78nyDStjqclh7kK2+biG1Tuso2OipfEfxbVmuPfT5sDlgoQQMJOM
VRr20JFUto3dF0bDmHCx3r+skXr5YTZKhZu+EOxVp/hRII8wglZMqVeHaEUkQqS2
/3FJgwGKDGSdqNOqDlSLujH8HuuotbKD8eIF8Qii/Ry/ORgUQn2h2Z0DSuk2YSQ7
ZsffbtWhxy9lBikw3SMReIlWcwNAfyNhPCw2lUBrwz3sIdQzNriSJvtj/P8VRqx0
sJ+nusNEELdvE0pbU1+w6oKNx4/ioe6v8Tc7/nNpKEBVh20ljbctZMYXiOP/njld
uge3hVCout+sJrrpmht52iDVpiHhSr+PQXFeSA7EDcc7EHLrK4euG2YfMcviA4M6
FzhJNcYBg17FFCHnlp4ksaZX8McsofyczhjZTg6OJC3BRcQgUvio8iVNpOh6OEI/
Zu0AfLsHND3q3CMW9OclLdKoKZNGKGMGYWOKaLtLcATeSaGce50Du+QEmxAhZg5C
JxlZS8UoUB5F7aH23YGb2I1En2OtO2J1XLOt1oC8IWCYy0evK6Qg+PLxg7kGjmui
YSShDWspzv+YiVIoq9wGjdXkb32qCddLMQY8beAhleuHQkDG4DoG+CyecFQpuvCM
rzphL1QWE37mvGyzHCx6QheceUDhFDK7W17vSmB2ERi355bgZi9OH0yx3okHxGGn
D+uHmr/qa/xUGiFm7rPnIwUXsdHVlHC/8jXhU7k7tKNr+YFSmapJa8eOfF6S/sfN
KsCA665CgMqOJ5HC07K0LtLqfBUg3ha8C2y6Eq1Fry8DWOGoYq2vC8+tyE5H1Yvp
tTkFfQXwd+tnj0Eueu9ok47X69kkTCG4VMWPC/hOH2DA6dkmK5B6wjTSCwaBTfBV
26nr42wCFqaxnblo1eWPQWKTSCgIx3ewZaGfPKaTuT1PBbzQzwI4O6in77DBzDmB
XA0XeTdKN2yjumYrhDlG9t4wnyNPwZdXB0aScg5GmkqEzzmMb2ErC1WVz2iIyQO/
OgqU7ZFgOKsm7gceAd7zCbAPHlgW2DG0m0XCT2hGVwRcsRK5W+9LsdY6fbb+eE39
/IEPw4oNSOBajc9n9lqIDnAckN/01B8gHNUwNeqmpbHhTc28K+x9m6Xiq1UTbpC/
FxiPTN5VGOQl//PzxswAf5O91BuFk98wZTxYJD/IWZrDTTZetR4zaJBZaK1+TYT+
aAhIGNBIiYKWQNH2b9ozNbldtSF461GzOZUV2hiYdi6PYpINiqrDw84CMrDdpFR8
ZqXWT1YLjQ5tfw8rinRp9yudTZ/uXjKHy7flkTDG6y+8FYWvCRAsWiURw7egCMyp
ET1tvQuJ3Mdd6EJNCoRwnlZlR+L68Ac1iTjHWijHsoiGw/9XJvcESR5XULvWnprO
3zlWP7C2zUOFqhJznYOtEHjyw+uxWdYkNYjoi1CX74+H7UuUm563hRoqksno9J5K
W2sDE/fb7kvpTsfOpYTWssPMlskD5ygKKXgiZDb3If5bE/ZwdWu/cyFnUXS7XzH1
/th2o0JX8lWRqjQGUVvJjcAbQuE7YcyO1IIlu7FrLStdiSVG9bish72o4e/1fbnv
YEseQy4P6RzuqKNtjjekbNtBWPfjnZQl0fPCUN2zGacJ45XQJx/5DF3TqGvQ4TZV
HroYbTm036P6dzPWAc7ZPPYEH0/Pe0euzN+Y88pqRKC3gMNgJTy05QmTEOiAnFyf
IMvlXj7rdGKN9m0f3oT30bEKEvLJhqMVpk2UQ/gSEe8biT2M5FvUqGkLocP3dif5
ln9mkZdWOlUpxTbFycgG4JKHZXfTqThaI7yrTyKNhZb+Ywyr1opsXXo57hi1JB0T
M/4oxMSVlkvHXLZYQ5Ixp/umtEnV5hRU8+Ihzmk3edJSyCZd700wCuWjNH0/pGOu
+Fck7U5hWK+4bLsGo7mJcLFq9yjR37LpD0vcvCWBuup3uBDAAyEiQXeqIIbjrGI6
CSiHqPmUo/RlCYyM7YwVwi8Me8nodOheI49sFn7XVeWnTRFcJUfQnf/t4c+Y8D8k
j3GnArjg2Itp2iNcPWJLuopiA1ZDNInJrGIfB8k6FD6rCAs+p7kFlZlUR9FZ8jlg
cwW1szPiPSorOGuVReZo25+6C34xIDY+yEzm+mUDWn4GoPOGy/WNZTANzsSaD66S
knhc5Bz1au2ZJRWxgHOzvvtiDKlbvfvhhmzcAh1YyAM98FL9yNg55vAS1wsk5GWw
4wb4lQt+DrPyA8ct5cZOCvdOvAcpBz2IZSYUETL44Y4ygquNDAvgrzSJIUiBkLsX
d5f+mZpj5lzfWf9IG9/jVLskjD+gj9oAuSZz1lE50mqiQZi6rl8tJUdI0O44w+HV
I3wEFtsCNz60WqdBZF+PsXQoEnw6v7+OTPu24yR63mpO1m0morThM6GbzlqtlmHH
DiEIcGktlFwXdZI9+Lm/DmNp9u3gvbpF4xYkNG+HagAYKg5FJaJ++DDY1leCro/9
SCvgVIx1EqxotXs04SfnaOZOxAdjf7QVxkbEBCXTdQs2TIwRnB2PidUDt3XjmQu6
ZIRFSIukVquCMZ269Y4K0a/jjd/wryW1iV7emDH+xOpDV6Trk8HCEQ0LvCy7VcHW
JV0PQ1+2wj0tiy71ufVGBmvmARnwbZ8+SyPaNB1hrWBCHHsTY/hVz67v8B2Ns62D
rrp9eJ44296JVm/hJ76o5NkIhRQiUB/zm7Fs1J36QT3y6j+DZ5UZ4aarRZICMvJ1
9GseWo1F2YWRYoCp49fS/i6JLgwy3gtoV/qQVpyJCRwVqiqnhj6f1DedRt/GHnMM
J/qNrY+M8Rc4DR7U1dVunmLhIa1PvBNoeL22F0rdrJCEES/OaDSIeqVm5cOVYmML
XeOu9kpgSvVE+8H9/hNL1EPxuIne2iK4TW+Eq+by2xALbUkE/QU+B48wXMNrvX8i
MPxHq0mJbHB8QLVx0/QyuE6U//hu9mdGi4GXBNlqsHu2FH7pwoU6lyENnhNbVjUs
Spbvq1jeo+vkgpy54IRG5Aj9eee8kfq9ngA7XposH/ADRL+zX4tas0r7II6AgACt
11LmfpLb/Y5DLeeu88rRt9n1x6JyVVia5BNLXC0a6xmqaHMvHc4dOOiB/zChBABK
012G8ZDc/nXOegBviyTxRZgJds0/+Ryyo5EtvR+9snCPuG5wzT865Nlhnab4whIp
sCZ14hykS4XvMsTMK6X1T9eVbITM9981H8OoeDYvgQrkRq1TAyGwi7Lh43x49VZE
BN1IL6a0ww1Ia/HvyfJ8/7y1FTA85o3bghclGhSJGeg6pcCLWFT79iLEmnjpJQHu
qvDh/rgqpDQGOU2CxDkiJmRx9dC2Wq8h6+TU3JnW4Xd55XEshD4SZgYMuxkG1UYV
wfyyf3CRYY+kgulJV/b16mnNQfl4cVsRMYJRsh18qE6n1VtxrRUDpr1u+SMENz+7
IsvipaOH3VfJalI7UywcW9u6EEYhCkzj0hPVwGXpzBE06Y6VvXm/VxDJlr3CSMWg
6zOCMstYpU+bqgtQiG1QIaawMDDI52VM/Bwts/kjw+I60P5EN6BNFy/9ma3gZoUU
qvAEYwWJS4GSEP6jzDmE36CDrFjm88Y0zF5GKOIu2QcCDgTSQzmvHnsCpuMcpXc5
/OxK+Li1ICWYl8kUvWxu/tzi3LMmXW3FkmFFUgu2CZYCLa9+qIuPLWAwteGensBk
KEpd0prcIoBbpCTEMkAfoE375BrtUnyqBtGoN9kbotr9ODMkNc7FWUiH9ECSVuHZ
/lal9Vd4cC+EB9vSCGWGMV0LKCY73pwg/+gWqzlzYXUV1HAnN75xmc/npBVQdTh4
mHYpzCbEJgjS5Q753f8ZLCZeOPS3JUC3CTSalAu34HH08EuaNPqyzW+9GJeq8sVi
JyHZoV5XIxVJcnPMevh6dGE6dhz9HrBkMmJaBmFMF6WNnU8KKFoxfC0IVqPJM2Wl
V507oiBeU8MBucf11zXrj3MMSxJk0kgZ2PCyyj1nYVmyuyW89j8LcWjfshTayi10
3omqR7Z6okbRVTV6m44iI+PWUWyatORwRpOhi0d/Avv5+ffL6uPeXSkJCf7/lWxM
THxhjeewJoIOQteGCMahAs+IReudi2GHhGqdbMuWk4SoUYDZHowhes5PdSt09x43
9wIChCVVjYD2ZY5SjWILr7tXXSaO2pC0YpKVmpe50+yWRr469MZHLMtHjUobIM3x
sc/KbAnvPbfAheq9oZqlURt4+NTaVQON674O3JKyyaquK/rx1/V9Xcdn7yHJzosy
VcXsPGTAAnRRe4C6fLGec7pIj1HyQFSlDOpAUBM/SLhyfmBKgjZXq9WlCjXTZtEX
vgWyWLoPttOXvZdbrbiuwidPSYhvb4zkXbRQdHKlITm1Ud/lytGSfERWAAo+8sDq
jL0BqjtXVRH32t6CExxc3ze+XI48xR59UGgUdcJdHHo8yRR9LSdNx2pcED8uFVn8
AIWqAwccYu/SdtACYtvIBr7ztS+WWFEe5GcCA0S4q8qoFFjwkxNLxZ9/Kg1WnL0x
72qv/uyicZfEZmKMxb1i9MJwYvNoZ5xMFwmzDqwg1DO4+ydhfojJFCf7IVe6KeeA
xa/sODN6JtlBsKHmi1q+IWaaPGQkT0Dkf7xN+wVD+WBJvBeueJRvL2SLUAlBajMo
oaHTQSmXKajr9yt8uAVDu+HKfst9auODrs4CSIxuCdzp4koBTdvbG/0EvZUL01r0
FKML8N+MUu4Tn+5an8XPsdIlIoPis61K1XoYkdTCCd/WjsMTkIe1hqlUCfO26Hkc
TYrhEYAUxn5yTBstwNKJFkWMjjAO6Shi8iXxZZN7CNw2wl1YSlOeZHpU4huSEerd
YlD9GkX6kdKuIFUm3LVBqxxQZ6YwLeBrQloLabI0ioyjVZIZjOBlA5cq679OPU+1
0xPMwHEhQQyDMeORPxak/IP9nCeL6C0M7MG1Ox306lE0jnuqS679vKn7IuhK1PW5
VjwNsIHXamqBkWQp/NZ0li/OjRMzlsJ5HZeBBcPk1Eo1nVbGiSFc+eGdWbMZkf5o
0e8JPNiwHvVF1jwMdefPEeZdnOyw6H9JrJgZV0rXCam6iJ9hlDFON39SMQGYLEfk
pqIIPpF3QOaSXpmoVuvSLhI28xoILcme+jnDg/4Q4kxb4VLsCAfkLtiWFmLIPzno
3FiDWubYhlirk1qSnupJofrDvVaSsOo0Nj7e4unuACodOmfvFpL1418AcWsLVW83
z/K7KciMf09tKVIw4nYHFVH+4gjRY1TYKZF9mK7iXVj6fuFhtxeCadcDZbUpX8wa
2eEpHX3ZKoppEli/UfJG6XTjO5CXz8sgrxkeqzQkxXlv+lm+rgOjfa3MLUyoYUkl
K/jJDFOzwasDBej5ZU9lfZ4ykLr2x8GlcOgqOUrg1fvGEdKJV3uToj95KxegVV/I
SL5rO1QWfo/jqgsujihlNIZ7DabkrH36RON//ItAVeAkmaI75cLx3W7xXP4+C/+Q
YmvsFY8FEgVaLBlRVlc/0MMOQmlZug8LqcuvNO6zSbrP8cw/ZU2gM0rffRf+4J8u
oUQRJNwKvPEYCieF+yoXWbVdvkbC3fGlfHXq6QT/cK5iDvM7sF06x/PipoBTWgNB
ADygtIED4jJSILLheKKgHlqe0WIDcnTAgs0aAG0D8AxDpWo0g/9YFyunhvg98COu
iB5LkaLMZEd9UzMp+iU8JUNR2G/KEnGkvu1qeJfO6fnTgmj0t4l/361/gxCbi4OU
I567wVoRzdnBiTcec+n+adB0ujINz9k9jVEgMuptgrdMKEAb6mNqOpHVHBPdZjqg
U9mMebwFlE8X2uMhk4DFa+JuOam4VhLu0Bp4p0T/P41X7qWEmcicPvqoAJExSAPm
gsXSxyUdFDc2FrovgBOQ332oxiQMXk/1lArJtJI2TG70jnKap0dbjN/WDPeOwd1Y
stxh8k++4QAv+3hvgEx4ERgAmJNjWA9TGvlFgLrBMUEUSNEXz/Cz91kI73GrMreO
hZKueZAGoW3sKf+6kAXMyTYxadIG54OVk2mH0mE70mC/Pel9hPaakwi+HuG+QfVF
mczWpZJ1rCrGqYQkzm/tqSBqgu+rfBiNSyhXA7/VPw0v2RV6kjcASmjq+v7/UF6z
/dqyi/XjYs7nmgYx7mpTwD/SXid6IDtK00DIcf5t3UXcrRXPwMpVqcdt5PvZyQAd
ef0SVjMMvU6JCs2Rhgv4S5b3hMv6B/wqtKAfemnRpI9IRgE4Gmty8mIXhUI4+Uc5
cDqj6wwMhu7qYk36kstXQ1bDTnKwx2hLGgZ8qpCewu898PrkG2pUSCAfZHLQI/Zw
AFq6dacyFkWU+NkISI9k8tisMP8m18Qu3OeFsf4zZbmDQwp23k+fhlhCGHTIC028
d349m+5hx+M06lm5P0MdFYg8saWAUZjT/NUetTbkGQuqI4vCxjuCc5bxyywWf2tf
GGC3tISZj6wi4PXpO1rtaBgpQ3cpBvf6Xhd8OhPiiA+03f+wJYxOrpqJ16ooS/C5
u2uSz1faKHLHizFp6HYaJmUDhJ/XmGjSwNtjzlO5JB6MKMuro+5W3Rv3YkUG0gdl
KvrElzXIsk5/r8BEvefHFn4RQk9DmrGnxKJcbt5gl+U9dG3bPpCYYoMkV1BvV7oN
bq+xSBU2Gk0iRZ4O8W51ucfVYNhqwDekzTh4Fe5FyK2TPR8WONSF5nQhE/aTQ8k6
E3Tw9qJwFCVYtVuxA9g+zP9t0pgUywkXjPoDWhdwRrywfmHz2QeszUWLZYu5Z5OC
BSRkklqKTjjycOQF8HW/cBY/qQojD+ys2Klrr9epgts9dUa45JEk5EdtO49BZPjR
TkWY8OrQ0vOpgNkAQw9qq6gRyFxdwwFTQ/JCU4PO2PAAzIs9BbEOB6mBfSf8ERJj
IqshrB1P5HdHouPfLx8+21ZG++B8OMmx+LG5j2dfD9gHXQlEWQyg5bJqZodlNlNG
Uyy6hjQ87Dn9BOJa1kd1iBEw+KGxVm9usVgJ4HAAzBs9nFNsN2/+RBED3R5zrDfY
0Nodah/FFCDQqjybuCjJaLRp4FfVK7TE+RHCk2Og2ygAkuArUalacsTZQGhrzzk3
FdgGtgg6OGIFhw6RkJiPfrbcVfkp+FkqRsDGyS5X2IiSkIYJZ8lv9wIHufvTKjdE
QHcuEm7C1pbdfa3SYA1Z92cU3ap2cxQeKU0QtvDv0mYXUwQHSk/WVQ1twV41P59d
ysErZhVOgqQ1de6oxxSynqqigIXbFS0W2yTbVuR7aJKqbYzU8scWXVx/Sj4YkjVQ
HklFXmAKgxPilrggdgHINeY6S1rimjdkB4e8L14aebB66Lcvyw0JeHng8Bz8mtqj
lxgEWHCZRdm34+5uHgmd6V4pXjJ1zjtpZG6aJuREjSMNEyYne3coW1Doel9VqdPu
CJxbxAxe8gqmwzC5MAQ9LjxcgoiUg/oZBbgGKmPVNzuOU/I7B4IGomNvNhaRUhmi
MZ8G0R7fvDbrf5pgn/5IABOPZdQD2pJ+NtELqinzL1BYiycsv4JWFeLEp2Ea60z5
r+WJ+ql4llx2G2QHWx6KD1x6B6yEUpFG0rPaT44xvyrwMGACnmWMzWa/xy88pZ4T
uZjOiNhe27eFd0H393MRoKdI6puzz7/UYT1nYI0JQS/oZBjWl2N2IEk2S8fzAXaz
GxMqyYfdX24/pB3xA0nbkVvetHTlHWIuGobATWzqKoHpfn3AwUN3NrOjTT6KgC0D
XlL23UMJISXJc5abi5rt0MZi0IiE+DAiFXF9o4EO7SDnPh2LpvBYtYfRsB9rvIA1
Zeo7Fb6NKk3K029pxxibRjBy4MjSkjPbaY9wUqa/Niir3Podupqlfnt6UShskhte
/hl+Jw8uNuY2nvKUaE3rsWx6aJTlfC3SYnK1tuDANAT22tsSsTcrwkbVFN0MricO
C7dNduqU5U2bOdnWEcPxciXRzIsxVlnZMdR3ENH5ozWJu3b/t1aAQTPNe3Um6IR8
ITlWT2r6z8DFdXR3oWZ2hPK7qa9454JwynZ97qBbygGprzJvF50afODGUB/Dbu0o
oEgxWSaKYdc0v/+vC3OwzWMai9QNb3VcK2pWt2lmwNB0meFC/DsWRmPGmkavAVEc
bwKOGcuo6bQW1x7i737ATvHkgObmFtjth6gJbnwGiEQHnH1WQRA7wiMgfFQo53PG
TyllooJ11oJ6HwAHTG/rHHo3T7C3m3DjnbDfYM4D0F5+IzhIYdglvfl4dyRteoFp
DQZScC1mdgCgMtQzRmSJIYnQGgScInFUaCoOlrqGNCakKfGgL3g62JXNOPKIrmBk
c2/Kn66Y/K4yo1G2jgUiFrfuBDZN1+A4OxlnQr/5ul6opnz+RjPchLw6celg1IfY
U9+7BRbXwkKpZTVKRBW5tDC78hfsWjUOEgGzchX5DZpjyCt/KdL/mFqGlATE9EIB
RYEs9CV5/0rQtqajsFSWhVdVFJjBSCvgdT1USmIUHL8phJ+cpYw1yZj5MgLypMyf
VJtmp0HIII02gOTJNZvA8cnxXF+iJSjyHZktGa9jbBtVqIC1VegqsTb86EVm7Brn
o0gZfkvIsBC0wR4gWEzjCZf1Eh7FUQARdwRBHls1H9daFSE55+YihlxGbSNttP/E
EF71/1aYEhFp8ameeiptjo5nSyXsv2AZtNCyLDZGLf3Gak3Tno2O5dBnlT5Hf8dw
Eb1RluQHp3/7OYMIlkXtTI2+gwTSWNgkeIS/2hwCoKPG9u1QVuor+lgsoCS/JQNR
11OvMOqAkjg2mvRJIOc2k2DN+m0NPmCUThS9CCsV8FoyszDxl9SlwA9T8+Jd0xkG
8MKppv2239XsoVKHGYV697DCyKVVwDmSL7FA3cV6efhWnLNgTAdXXKeCpAIyjDsz
+JZJuCPVcrr3ALZ3N0MoG12KM2xvu/UQaibAYdVMOKsMpDEEdD6xG8uPcWszBGtb
pRzlA/MvUFR5FLA2BNuuAudi/pXfWhV/wy1ePWFsX7vNhNId5yYxLK4WBtbTF4Qx
tro9i/8iKQg64kC69uEU2A/iWRH/+1BL3gFurwI8B/ZAqGmjAX9HrhKKCVASyMsB
8Jkpm7xU3bodk+6oXi+ZEMUl0foW4V7StpF8MGi9reIzImgpKzs9R2mn0er9gbyT
ye45kibE9jFAYvjtySbOry52p29ly2uaiCDXnQMvM2CvUhT8mFFVQMxgoeHNk5yS
leKpcrX8i8M7Z93nW99gp5KaiSTcm4E3xRRc1VKlxRLVVhVvwbiHvqaGoNZeUOKl
taTfJcKuFnPlpMUhswOHcjtwF3p3OBqxPKgZwW/MMSdSmEvp46TNgr3KSPffNndD
c3Mrqldpns0xKYnb6l9hnxI6uNLlwua0wap/Gh4C6MKCAqQyarBcxcvFvqYfxUoC
2pBolOwHorDv44OTVPHmIba/NdoXfptfzQK1LmToSx/7TyrNS1Q4rokrNbqatlge
LV8NEZofJ3WkvTtRoa9BUi55DM+1hrDuYpbGbfj4kGMi8VzAyMpc37x4RABRPUbU
/JW/JkiASBNLtebf8T2NmhvDunfag/FR0eOw3Pal2Hf6AJ/9zWKdU63FX9E4G8mB
dfE8ngb+7qLpSu/D9HjULnekPa6mW1S2eYuTpKYH8ronGwwUAYdN8ZpZW27WTd5J
Rg4I9GOHuEFEAgrq+K6YaRWqOdyBC+B493Zx7tx+v9xkcbPR0aFHQp9ff733fqyS
F5faE+NgG4v9Qqly1mtWi9n3zFf2OHrSlZSPi/lgv8JZ7Ysw3mQdObJ7Ib5/Dnzu
e8Zju2y4DoikLTRUTrmc7wJfm5zIahoD4WDOg4LTxZaN1R3tXBgg+ESa+KrFY+wo
sH0qp1lFAgIKQmgCmi6ginhaCau6tXtaGl1GsHkGkV6YxpfaSJDEETRKczL/J0KY
lhhDcjMCAgtUs/4iJMdUAk5WitAQqoBTCalKryPGykyRoVmmUXjRn83YKlK5W+X/
UgY+AHiTFDHeh3TDjRpKtZBFgII6kpy3O9Nw94nWx+zXBcyiTdnsuwyYAvhKhCm4
nROmEuzyQDwfXhn5Su0GfAG8EAD+PAWu8heEHgaRLXX+4HFtwrEclrfVV2wtkVwn
b+mBHE65B1yUhqYqS41NmQTdXu5Jx2WOU+4ZXui/uzBokTpBrMDflrSqwCNRy5lp
frlDa+G2XnRIjjn/LytxPM8X9uk+QiIEP6YBMLkUMTu0MnB+7aOM1PVZmb9EAvsW
nxzRgBqZpqEZMQih0GrbE0GDupQuOMX2hJzskiL6gzxOh/bjGWvE9atiQlNbzVEl
7rR/+S7spr/yWtmbAF7dILzGu172dfPweh+edMCh6L9N5H6DEedaYTCjvRwDYaou
S1wkyI+7S6OvqMCHiomIi3swm19TKOShbfji29/kowN6fZai9obhschBmeKW55mh
BJ4CyEs0kHrj4pmYYJSC88I4hwZ62UM5SSJ2FpOGm+LNl/wiW3zfMG+91fPQhg0U
RaxpjN4E4FfsHbNuTqzOk+ba5F+6wqiMxbAf8DXFeFwPVKrdOc0pAx8xY3K69Iyp
I5MrA+AnIvZ7DZvSoLWlkKRG9XgOzz/TX8RZmH8TfYLw+6OpObCg0cjBbycuQXEd
RHoSSgaLDDY1lGsWbBz5WfGkmwOv5yqXtrMOFTI651Zyf8SvhQRhC2S3nQO4lMPF
COxXUZ6Jm5P8/ZtQKYmZZkjqU1MlaGuBWJwwc2BbNwDx+tdHJESLNRVqIhJuKP6l
gO1sY3mKnbNUsr5MQLU+wtzsVWozS5AJaXIdPYNwL2WV0XYyAlTJK9HEYl690LGJ
K5gTZhx811kNZy2Jsq0fLerunwhaW3L17rZo4mO0rWWVmcJIPJwni/tAf+EMPqoz
pSegRJAmYfi563WyYL90P89YbIgyVCQZOfLjV4UGLof7MO44OjktAAH8XZ2LFi6b
oDgqBvmyBk75o50P6XGd0aSy3Mwqyme+AUkSAe2+dB7IdChUUlxQchnlQ4cdbMeE
EeGO4ntL9r9ptttTy9uDfuYwSAfBXemDj/0p+kdeppY9jl6nYFEBJkN7QqGFhuxZ
lVvxWzaF+Wut1eylOQf0Q8EgCMMA38/EdMZFbmRzvXbdwHAQuPqCU0Xku4by8IxB
hrllLiiuZ6TvnEZ/UBebZBHyQxjqSOIxP3+0nSIF0dsoeK389cq4YBca8w8H7ZO7
/EXF9a0sgB4bOn7WZ7ARqMPp1cGY20Z3s2fda3MCQSEYbEdze9hFYvHOiaFoyIyG
mKl6o7hwLUxehDioK/6sXZTy03IKAapbIYPWw48Y66Tns5BSyE2WPMvz+eEZJ1sG
xE9/Xeu7chj68mH050I+3Lpqf1xIdiav4oUWgsBnbyVwDZ++g37M0gz8xw6xWk89
ZxTMwldJSwI4f343k0LNS6jPm7L/b4XQ/StO59roG0p3DcxMX7zqPrnas2AWRNFb
STwzp5Gok48SSpD3zoXLFIt5y216vkvBZNp+I08wKyWdXp41ywnk765edR/bgeCv
Rn1dQpjQNebUGvvH3QRRkkQXMgX7gunP1ZgjSe2PzPQsbrNqyNQpMSFXqAHeMCIe
iHT/Ez9RD3inhtf1mD6QY5iiPz5999ytTTHuzq17LQfO21YF3Chp8QGcKZJDCYFs
Z+fdCEeuWaSyoSkq+HPg2Vt9ld38LyAysLoE6BEZwD3A+Sn1o361r2y+aJMWQ8Y8
a4GLLIT2SWunKzNAyUunXgo3J6+NqlqfLrx07WwTwbk+aM3jUotSzlWovmSo243N
5ioTIG16uu+YvmI/1ePN+/Dvwmt90PgZGOb5Jbja0Hmzzrn5pmItpfR3bxQKu4BN
TfOvxlC1XDRHKAjtgUWRXEVqWSQSxQInz94YrkFYeXWX68olAQR31qe604B2iYK+
yUsf7PtvnHgiaCFvJ6MUsA/ZUFcpu2vOK/nsdqIr+jBVER6xO/sbA6tMm0yOLioD
K+OrNujUgweOyB9QzEcUq9o5vV8QdzbzuHYsP6Pw1Fn5Um4VQcrchwhCkxBycXfQ
6xdhPaPmy+RJiEc8MOWT+wxtKyZ8u9cm2EAxuWT66NPENoZHQ0CcINS69MUu18tp
zpVuyxvPwH2LcGRecbWo5xbQ3/v9RmEg5Y7WcO2UtzmY4Cwx4tKz/F94R7Sm6JtU
zX2d9Up17L9Ew2IxSkNUfV3Mi0S2pyHMpEulQJeAYEDL+PcwOkGIggSKnNtqqllO
iIyz/GLjo1oBuiI/y2Qjz39cMu7rZlkimLoakefHGW6RhP+8ESkamLOJ9pYDaIin
LbTjlfBduWoq1aLjoMn4YrXM63Y08EK9zzeYtnTwoPJkXJrNWsrStQDEFque4mRE
yRFbHNH0WtNfQbnxpnFDoHtTj2nTibkZbW4+NBVb98knMU1AMuskn1gt5bbop4+8
+AR9Sll78wqTU55TqoCKqNBF0aP5nCtx6fVDYA0WorGkX6is/PkSXxq3DN5+tnxH
lr6V44bsmi3m6zBHz7GYTDZbt60fuoWCOW0OQBxZ1dC6yBqNo1Qv3xAh9TayYCeU
FUlfNmtdEANk0F3yROZIqIf0xLL/A2aMrkhP/fFVbSq17qAClbtn1kYkYiGlFIXH
qrbgWnqvfZfyPh8icFHuf/YlSpfT/a2uzKMaStXFqLi+NyPvF6pvOLuVLJLRa4M2
agIlAT5OEvaQjeEORFCtA7rQX9p427JLjjYegMdEDCXX3ET84tKnQClzgneoH+Wn
vN/Vr9COajMh3ZWA5Iq0ytiOGbPdhAgzRbFQ4GEm2eNjRhprb4YFrFx6ufSBOd9X
tlIVDZpZbWIHiCDnFVGRp9O6dzt5czkw+V/vJj93Witrhz4+SLcCqCZPoiDwYjBI
wqgHHdJJa5g2OXbJtEl1CBzFq9J/2y3XKr9DmtizHvgi4cfFZmvLDzQKdYPRC7Mm
k5vB2jE9lURsiQ77/9ktT5/dE008QIDThl6vUNYsyBPQkF/sS4rfSlndmzzWp028
wZz3svkEaCmqzbnZAFfESRTMIPV+tVzYlcRiuWt9ZMcXD5NphwBmwuJm80g/Opuh
N7L27vC5+6QAo4B7B6f3OzerHwYULjp3xlfSjK7SgXjN51iJ5b3sy3oLTk0urwQv
IihdLhC6g9E7/lOiM11tezw9EBpFsoZUTgAgv3ncKO9ntvIyOEcoABaN8yRzx30g
SOqK42vk7E9o0ika/5YfPWXkaWvJnYFLzM5c7u9uCQSuEh9PFk7/UrEMlDSB25Xh
V9PV2ywcCeTDU4UFUt9Xi5oRFGl18jKk6f72B4w31Fz6WX/st6VHFx7NDljNpvd2
P4B+MmUqHVqvpBmAy5HkRpOCEEzYTv81HHgCkzw/0PdMbTmIOOk3T/pjTE8/MCva
X+i+rYRCbAR7nDuXaOAa7J/HEszqB70p+Ts2wIrucq/QYe4CUqk0p6mzRFlLkxjz
4qEO/dV39xfFyjQHQ/+8jr7OUMBT4trw7QYGa2dpY5qmWxQQzCQv3eDqcYa2h6Bi
mbKwbk3wvBYakt+/Gfhmpm0/PZJRKdc335EBfSCwXCfQEImgCgar5IC26cJ7tzFF
3WP/Q5XiQXRBjOg3OhfUZEKGuT1W3kbOOGEDhVjg69+hg0VMA/f0kbQxsXKRZpuI
RsJkBnxzQmHw7zNKtEpQKTRYk3TweVyaf1zGVEuzE7OAN9WAEizp+1pxeaGthSlC
MORb6VylJeH+OAQ6oZf7NXbgEcD6wsU7aL5Fgo26VfI/rHj7q9EOirFkMzxoyAR8
WArmNLa4WY+cPdR7/A4RuOT5/fQ4d6PNEBRDiypdiW3IBjqz3/R+qDrZIcmz3mci
rV5DG11x9T9DQ9h47f2W3jx7Ez8HBfd2Ueuj7FMSqGyNb0CoZ46zBixPP3M3rkM7
bgb6sZjDEgNyekEGuBRFXnq6T8cVD25dOgXW/8kxkKbvVBm+W9PKIndx6Q/1tRVC
rRtv0qVUVFCmIgbLKQv+WLj+B7MSI+4fyjUUPTk1JV0CGaCj56p8uyfkBdz/nCAp
FynPVxcCLnPU3a5yjoIG+sL9+pU3xlrCrVJRs7HzoRPKrFwkb1Abi1cNpMuGRxA0
9bW2M9VKSJmmhE5ecRjpUKN5sXNqoabmroMx3ykYuJrb5A6S1tWiC8ke8wLSjTm2
CSIKw2iuh6yG+DEkPglFlcwfJVyEtwthaG7Y0rVJguhVF/ExwMWT60Z14WfOzA2d
Z0bBlc2twvb1qyoNGcrg8cHt3BXCQK+p576ZzYRKsMEmHUmiwT/047JVsVK7QTbT
Tih6ooarH4yIgId7LCXKwQcHwNOvlMKPlodNSDpgSzv8SpYd2GC0KTs06qgLuX6q
aAsXZBPSLErxH9L3+JxaJcfno92Vif4rrwUM2Gh6NSpaee6eQdO3+GwfLPznTGAg
R3O7Mm+1VMUhXaivsW+fnfp7ZGB5GVGdsaWbeWqNUeaATLjUNh7L+PehjW2MbfUJ
eTA5l4WwGjCwolbDYIIFGxkjqJvTXwpOh3G2XyqO7Vux963af3Bd2q30RTJF0G4H
nhStCZNsR7+Nv0mYPpvHcAPVmgglgDKyKjGbLuxWxlbcavtDKUyhpAhBtVRY1sFV
MRpxLC6MH74f6ktqSblbhCquwajN4F4IdXmkvqZHPpx6rBAj5q9gV344A2C6Anut
s0yaoa6omhKeOlHPHzkw2WRF+LTwf+L38ZCQpG7GR8AKnR1xsiGe8RI3T07Zgw9t
vvkYUBIyIQq1j+yHdMY2x16I1nQsfFJ9PjGJCrEfoj2jjD7/r6/VmMbaT1ws6i7L
2fbUyfNo53nq98CBMRImAsYZAjYcvaOmVz/cySOLSgrzxVQx2QFGQPRQUOUrqDOl
XQxm3eXcV9gWUDkyS+r3Sr2tnoJQB0Y3TU7d2oeiWwNR+Si1ZrZcJv5wIb2+ia/u
Vlx49wz/6SkXyTPaFL5/UziJjnzzT2C5hZXjTlNEjrt/WkAFK1IiPJMch1+YpZ12
Gd13c5F3eefNwNbwYHhMkxfF2EsSM7zxGKyyHB/AsjPvLO6j1c7hQfcSdO7bdFFk
Yt5lIM6lCO/fzllUvbdy6wyBWHJhQ96eVQUAwg6NswPY/Ikmm+H/+ZjPv+2YfjbG
ZX9nsji08IPpyRuhvaQzsG943InJNOKPAtW6kIiXG+K/CcF8kWCRsh1NVlk+byxR
LpL+eedkJMPVzqqBMW9YfGKidD25JBklqbWtjaAdNO3ZMfirpVtAlGbKBNzjoWSF
EcQGOaIn/XaWI54/G4EzK7reuxklG1nOjMmPhdJad8wxeFBBg00bGxH2IHKDFhX0
9Y6U88iaiqk3LdyGy1UaagfN4LSrwdqmgmLUx+81bYf7l+FwgFYIfHwla5AV4vSY
Gce7cHEzhT6stef0R2fxdWjzSYRcXh8+DLx4w9oAsIxmZY87L0nM+iLX40YeqmBY
4emMotBdklWkSPA5H8IOKKdMR692d1B+TVOUxEDi7Y7fFmVVNOr58oHk07yN8tal
SOQ03XvcCLTNK/bmTOtC1EYXH26HPIla3RwtbqepIqL+38cQd7qaTtZgj36Kguj8
pxTuP9+m+OgOcrCemNe+CrzGHRsfWSeo1bl3l/TDc/jNHthDA/cUhjQQNA8/K0sa
YF5lsvkGsdKd7OMeyUHR1odmymWtye9Yd9xjKDIXbYWlE21kdmuTsh1ZRA5KquoX
YPOLGBEQvlPWAnoLQhQ55eiT1qeHxoOQvbHdA5pcwF3rDCrY4AERgdXzQXgffQQ6
GcMgtzGf7EMMD/41mNpV345EyhWwjZsIeuKfjSiGtbLZ12G33KmgcOD3WBdYcGNs
hktb5tEf21JTQG+NSHoIzHMBFLJugBmNiLfX4xOB3642CtznmnbMxArxz5E4ddXo
x2DJ6zQK0r2Fgjjb/iq51nLRHZRwxe9uastJnXVN4dj0r1CflujejMPnrE0P0c5o
8CEpwBKu+Bv4XcNjkxkw4GDzMFXGsW2bPAB056ZzxDK9MNhiKke015VWBh/fDBa0
HwR5UbZkBAdaipDQCMioV8L4F21c4QHLG4/BRYOHEs6ehQgAQQ6dizBpAB4xLQfH
bmSsVk9AvMHEE34szQnRltCFsaS+332tyka+Nr96HHGLn3yqzW6dIm4AhFNU8cFO
7UVdfAUS8NpTwaFB3rrm7g/pn7xC6fw3riOHqijGcuYuoFI/KWG7vox9a4mMrH2y
10nEuFW4ZNiF4AisKq0/Gt4sRZO4nZg6jmt+GtjWIoBUgX1rQHh93IdNRT3DP3b6
QlRlhHAhrYyApRbW5iMZ4hTyTJNbS0nSAwK7JAHaPGJL7WxXlQV1OhbTl/01NiRT
5vPs8Ydmc/XyiP0Zyv6jH/u3JkX1jpHfgTf0k+i/Qv3xpNUHt1zrLBlNjagJoEog
lFjvCf2X9rAcATcJw9JfVccNg67qpaxfQ0PR4u+BdqIJ7+S10gPFAiefBsYB/Z4U
sVBr9uS76KuwVqOdl7Bue6LYPOy6o6DsAWL7J2iNON5DKFR6UaNSPzMocz9V6fO5
l5B7A6mjX1P27nM7l89AUNtVjGrN0TqJPq/ciQNFbOT6Q41mGNcfIVrJtSLH6x/S
PDK6/8bduwL4EMievcwilXHa6I4JsHKQZ2BA7jzyhhE/D/VLfMjuaqaMLTWWzn+O
TcSb6E/eMtMzv9KgiFgyouBDmoJEGKzU/3veG3xLIKC44k7eJcp/2u/rK2oc7Ld4
4SBSPhkFo2RMhgp3vV4A9EHXpIp61Fwl8Dm9B/ti+l2YXGukGW/9O1mp5CVj7UIG
BJtoSDQXoWvfwHyUohNhjvmWEfoodQ7RLZuWlFipLGtR9fo9Oar1pMmDhfbl7Ajw
jz0nKb/1wo8tDFZr+dTZZKPRSXLhGGk2k1DZ0mrYK5aUyJUt7nNfhKlY8sNkdS/n
5cr1kg6qCiGYo/gleITDRvbshhBptLTK+Tix0FUjc2u1nnEwaFFdRwxRMCysaisa
9fI5uyhfnLwYgnib8GKQiW6gr6DWYOuwRo1T4gUaEIz8c0EprG9ikLnApenfyGBF
wGGUhzSj8ToMCVi2Z8GeCsdkOsJusR3wd/IWJNfVcGU34D/7ysZ7Gi7rjCkF2jmx
B73P9K0XXlKk846/He7GSNCh4Nq7veYyqXuWOd8+Ues1XR66nZN5mBmEUVG4wj/1
SYelGuPpE7g3YxQc3MgwDzqJ81R9K1i0e88HvRDmMlBNUqk+08IJPr19U8YpHDIf
lrEVBtOgf9ZZCS4ToUoUMTe/UNEH62DypCXY6O1PlALp7nSHqCeh3EWLg14uVw0o
U+NSCzz7cwnUkSk0ciHYeLa5KitrN13155V2lZpyjj48OTuMApDkPxqadrPSOZx/
imHuj/Hnf/1SrflH+xL06qiMHnP0yTdjJ/G2FpxMaiAe+wNCb9EnXMA4GQyoz6uM
arw4ALDh2tAeRiIetMYE1kh/rcBzF6216PA9xM6Q7XUK/TOoeER776FSYM4wMisy
IGHZiupEmlIdG9ttC6k4OrNmB5D6DlMFYgNL62aeaMuN3DG3GVJJ3f4lS8kFH3jY
hg/OR9251bRXvZSrNUX4MxQrOmhL7aMfGNaWvFFwHJFmjWJD5peTL8j46+3KP6ir
3+DH3Q5FL4NwskbSG+H8xiSVlKXC4DksHZbMMbPRayASNdMwMgH/0Fbq6AHTunWb
3BH8W0x7HJCTa5vXatDP0WKGPe8ZPSvZq0iyeecq/f5onlVISZHo/GvCFTaQf8Md
mklI4YH59WFbCGMqipxkeHFrcMsfhpJrYqaR38WRzPtTY4+JZIGi/Agxs5V1qOTl
nkycpEX1numgb2mWxfmufXbAOLB6VN4mFwuDoSxeIlCK7pUlCNjA4yhieu8XBTMS
FXbjua6ZyMZ/DwShjIo6BWTnR6plBFOXBqQF22Ff4Nz1/WwhwvPGOlDSViU0BDK3
wnISnY6FB6iLdQ7L/J16uhWGllsW9Id8DIp6srCAe+yWi44xJ/7zMNTsd0GH13Sx
XV8KaElJySRfu1k8iEnp6K6YxD9YlW0u9IuCx+0S6hMWLw/ezoewvunryVpQcSFU
lUVTmKwqYcuoyq2g1Tuc71DlOGRcF69On8YPeZVKReuZesPgmpDI9eLw+XKTc6vg
i8BfbtuXL17fvcZliyqAxraUFHSBThjm4p23XTenYXTpQpyNUfHgUSaK2r+NgtCe
zJDRwFDXYuFOwy3JayX5GTGFSfUHrwTMxe3z704ZLgVDtlPh9UeBYEdGItTuZt/p
5AkYGsy+VZeJTXJMh0A2t3bTQdzWZqAKUP5/4JiUNP2/yrgySkikEjo5ZJfJCuwa
8yncLE8MTRq1kn8R4p59TzXl298+ethl6bWOBeNPs/yMiDSANeAktltUZ6SmKnY1
IR/03tZNQ3exSmCYiMBjvW56niXat1bIJ+oynvxcwKKUsr7zysZCLwIRMhLm1wb3
Ty/4O3tJLnx7fwl1YRR+RqVq3pOsfuFTLSxz7JZY20ze0maMwBAr0EuIh4CGGGl9
pMuH5kYY7iGGvoqQ5jh2EVuSFVYfNL5JILFIajStHeX2e4eB/1CqqR6xAIVUhs0j
OeG3EhNqQZ2JcSORbTSg8uKKRTH/9GUQJgz+fjbe4eQ1Uh3k/brNsXCiPoGZdQwf
eV0aESZBsJi876hJyKNRebRUIucmXJt5dDPhqbqzNyJtFLkirmfT40+ioD6kDKpm
mcmkcDnXxzAvCwxfDPP9dLAkRqNGO/c9PIl2e7Btfq9E6CE/YAEgpL8a9ZzFX/nK
r5r2g6TMN9Zta1krM/cAQBsHHKYO9xvAe7OvjLGFCHfomlKiYuV5SOp1NIlE5tVG
Ac4nSZPbsArMYaJxpJp70ImC71baK3w1uwZOM6Z+1B9fqciquNFWOj3Ob/yJIU8s
342JSSSkUILSfrgFtJC7jWaRuXXnC1V6gJlbslDGuIYPsJk8/yzDzeGsVIKhirAC
ALA6Rkdy3bFHA6YffnmS6uzGVik9fVp5Xdm42YiwQlVQim4fejWul0SO64YWLO6V
uY6Ngoz+qbqUpwTf49RK0WdoIyS6lyCEz/DKoczFGMM1glJ2EuA5ure9E/gsmirS
B5DoBTefZB7B0OrqfiUkMll26/LLkCGfMTGAF/aG7TOU33i6QKfxfzO5Y1jmOXpk
AFYPOJ87e9+XviGYcRPB2CsaTeBXXRHmHqQ6lhmK5T64zPXNa1z847Ukpm6gOVfe
b9dJQ9tpxGjcBlmBX+tVggV/zXorEGHq+4ShKL0o+7l57b37zmXJVkv2dIUgLsd4
HD/gVopzDiJp30PqG1c+1EZcj4lf/Gqo69eAG1Kz7AcUn7bjTrrxvJXZS0dtzM8l
0CF4QW3y2fpnSrXE5KU1hOHlpwRfiMR0BzxkMrjGpZxRs+V0tqttru10gM726VAj
YvdH/FhfVodt4KWb2ilGZlZocA50EdVvfmXQ/T0cNxQFwVQS5/v09LDXroFu2IY3
G0R+0+6EO9AoMMzZqUZGQbqC0FzfYk9CnAxt7Tfknayx1kxXyTDGxwgFmYEaOK0X
VhWabJRqKpWZs39uiFWz1AQXRGeHjtjjBeWET4xQHX8seiP/VZORkqDSFytMx4rr
keda4qITPAH4voQM6i9lyZYL52521c4WAFewLoGaB9jJKM66M/5CElpqBD6VkfIU
4u8POSBh0HQJ7nNK5ufCOSnkZcfOvlW5Er5jROhEkN3LjobqnYED7PbY+R3E6eJs
WtpfmOOUQOOqAlyDGK06/uOwnFH0KXd4AxKY1hL3sPSoRxqOsqfSCXBX/gucBbyW
mAotOil0ixMRg9COEQOKUrSS0qAkIgIlVQJoXUmnGlT1x3/NH+cA/AcJBSOHNKuI
H4NiOTmZy2KabJBc/TjwgSwccEnabXlvSmkhuOQqYOoo0afqiClsQ1lHXracdeOz
pB8ZulCavQbByMAmSA4B+0CjjkwPXVVfSsuQfwqsvSOopYQq7awoiBykSSG1fmF0
4Dwoa7GPGK/EoTZpRaFJFLZ8QYyOd08V1GP/U4z5fnqsNlLevfEoi9KhMJXkAwPD
QONSei3Ff2Nir5WkG4f9IrXiy/pXf135Ro5Zoq1mfBO8EaH0i/NBFFhhUO5l5MzV
TZxmY7Bl6vgVtrMHswCZF096BIJtToJSrkA5BAKtkpzUAQOEXyLD3LxVAy7CWDCB
wu5KH0/6ViqU2TDRdrKZN7IL9rqyDhTs9JzX2BJACp8OZ1Z08zdh7YO+sT3ghBFx
qwVttV5+jiUYZfQWVlKt7SFZX73KQfmge12S7nFn2sR3queYfwpAnFP4p/ZjIGO0
uo2ce0Iw+e2Es5C2y1rCyWZsjTniVJC5FeeP5h77RWl1te0a0kbQfMp4ZgyVE9XQ
XFm+eMuAyF/DRz5m4VermwcoFbne/hUlPhGLt49R+3BuB1s4EU+uaiLwV+APv3NY
jnIjJpDNu710IeT2dLncGAedRXE2eoMMg7fuWqk5GlcfbNL23n2msaJKgkAQbxZG
NSX+fi8h9ISbqCPVsNwlMP5jCysLymlRvhYUOR8LBngpBCdWGSdUQdSJvTbpbn1E
Nu0OGRIEbdgmh4irpbx4DU8o1+rqLylDbL/6bn/GCAk1otdYtwZ7CIlfwqEuOKBb
3QndJAnF+n8mmeZHjrZiuaHJtI96ToVlJLHLGsrRtVTSCkWZiUEHlVhT2V6FFHty
9w8Dr8yWMYCIep2vc77ZIxXookQsL7+yGjaVqfXZPZJUliPzso/5/ohVAh/VVTPn
jiQ0E5purxbnCVkSZtSnfj810LQJBR1aVSUtKaSIfkmnxFFJWRo08S9Qkx3ioH6Y
rFF98+8KZRZlyKobvfVa6e759l0yh0nzPkfe5VZIRyhyIs9mjJBW0lGfCl70RFgO
wXVdE2Iv3Isq2oBbN8KkHqaDgmK+pFxAUqBg93UI9Fw0nQulU8ChWfaXErlNru/S
aREyifbLRZqT+N1K5USJLX0HCGEh2TqUnemS/6UORqw5OPIht7LfNLWanKiyHC46
HCGnkTdkSBukK09YawMk0mZqFxU9kFVLZOWK33ljnSoxqKp98Qs1W1zOa0NZi9aN
2IyJusMFLW3kXP2rQumXr92kgBrTIEs7aCD9GOuHlQdQorJG7n7DUM1lrcf2khfB
38MYadDpZzbx8qbNTfoWQgmOaPEQXBUUp5IqVsfMN5hDESGZEBYGNeGRg4J3RYiu
1Kt0UkbCdi4TVUirzCeECJKVAhM/TLdrpfF97rviDIwABuzbBvvzxo+ga1LRgUOq
96k3JC5RgKXlgnh6JJf658viFPc1k/pRz6R5LKui9/+t08BLqaRLc0wr5Qb2ANAm
X9C2ljH0TxtZqRz9XlwmuBak4mM5AbuL/wdwvZHSqsDQoYqA3CCPI1Jwodi4Xrhz
3cYQoQRvZ+K7Yf9sfvUSJHweQDiaSTYSzntADPLc6d+5MwNiONtCX+VCllGeAobL
gcBs2YgGSzwfeC2e8tR5+mvWsNwjImzgnr+MBNivSOyrapXyplYQqVsHijdyEsLt
8lcFqL8eITckAOq2vuDvfbxDahfnRogy21R+mKIN7nY0GXaCJNT0Amo3t3cJaeqR
aQD8zfvgZ+iAPWMnSenDt9Vbc4PU5CJRvBGhOmH3Zl1oF/Xhm67R+hRBnWrT3PqS
ns6W8i4ELZE8y+hPEf4KKF6053ROwCzg/9bLRfG26u6wTgP1CCdzGc9/WxnFEx29
tfXAVDo9uL3erVfievgvgVHIVdW9W7AdGrxgJ+cswK0X42lmFKYSVzEZkczgUTP2
YZMGHnSECmRUee3CA+pBU5JQ5UyuqZ/wl0DZmG4MvH0UIm+EZZ7cn9eMVp2i2tJK
wX+PNnyZKX/mU+tQfisetcRt2rz60vwTkjBi6V3TCreS0swDoRfoTrpgLIY1m5qS
PoAikVgfbFzfpO67IyovCco6tHOyhkdjdKZNikRHerRdJBubn6FtKFJaEy3HqCVd
15x4A5mPJnWhaaJ8JViTIJUW30Nz4MYRW63ay+/P7iRfoyGaN/fYpgjn8E935qvI
3Nu5SoIp91c5e/p2EikrFaZMvQy/NWinfmeVsBZGsg+r/k8+8vmEmBzaWRFo75XY
F3+bOZxrWbgSK7oNVXEsjQZmBCx88CZv7E6UFPy7t6jfpzmUWm/EpUUWL2CNVGeC
yOhXDLgfWntOZAr3U27PV9w7T7hEhTdA1HNUBEP0NAbiORLBui3xhvXinYrz5dvL
dqd6zwRuk8yMhE7/ERjyJcqlYWUsLyYjLpaPVDScar6jP8eBGUtmvu4ZcXmdYBQo
drMNOtK0/btcLZ5BzaiwQD46/i8rZo0vFP7p70HDVaVftzjyzelKK92sI+jAw3nQ
Evu1sewibUsicp6+s6CtEhIvVI/vC24+KGLZbJyC/2UauvV2v9f0r2xgWBo3/vM0
OQrEBkQQ8RNyBo8B7W/R76QyGJcviq/Qjcay3HxAP3D4v7I6I1AyvSrPbLTLVvtJ
zlsLvtiWvtJuyL0QukhO3FjYZGjhdnSPB4rzoDgSwfWMoXBOAxnmm4G0AUr1ZMiV
i0UFsrcEtp7ja5TclMDpRYgqFEQ8sygy/57KkqHFFkHyYuCG17If1D8GaDMufO7b
Z1e4ZxSbqoHL3ZSjT/K/TpgrRCanvqguJjh3wUW4qzwiAN3ff2mbQHEiOns/aLep
uwKr0zFR3tXr1WiE9I1a/200CzFEIM+ZirYR8kCT/7k15l/+xhYzM2Sob0/aiyjc
K/8RFtMvDk7Bc43ZBu2Kejphe7MwW59glwHMlwZHcbJzN1U8hl83WsujCnpASUNY
MSRjhUq8S+ChzPi40fxtnWeHiKjX8ITE/KDD8knDARO/0rYcMQCa/c0EsJ34FTsc
7Pfux+6FvKHsC0kXHdaI6CiVRklheTghkgHCFWR7OL4tMOfqe0wS7/tsR9HnjlwT
dhAAzJ3vYfLuq99V3h7UORy7eAWATNxBRWP+HHo55TRTs/68mMH0tXBLxUMlFKds
5p/3tGlBI/2LsoKKJB5UlFOOWyxVCxYFm5IqkTSMKW+gECAciPTgXqg/hNiLMex2
lfZZLl78kVFfKQ5Dti+gyFklnIxUGZ8PZUTb1xj7nvFFoTjC2ieOpGdwizq79O02
NIaq69+MT5mJxOA3Gsw2yJ8wR9jctK2+BS7lTrEzb4ITqdbnyDl3KFudwijoLHbw
2QChX2DaKvVnyMbYeYWSfEHBG+1Uqp271PXG5LT4ytLWkwxijpUTO3oS5CCmIQ9O
UinxTIZrB2N/8qvC7Kn+IFFenzkdfAW8B2zH5pCXJmPXxruKUY+0FHdKpDuAZR9H
rCAxv1gaW8Rc1gKPNmCkZmlQpQ/NkGrafd7cPlat5lAndrrvBtUKKHscnCQObzIU
xJyFu6uGPn6UwDVQSNtOQHkz0PcX5Bcpzl+yDPxxOz3tQaMRpPmIWPYqZFmGQ+gt
o8nz7IEUpO0ffoOmF6+NAY9HdqPyAoHRVtlR5T+L8u8ZlmlS9LU8aMHsNnHlE5Hg
da9pGAJIkX2NrcoiCjdnkw2XqqnRdU8S6eA++RQVHuHwgytjiPcLCPyU7WEjscnh
S23/FkuHrn+pzDEkVwTaGiZ3nZ1Z4Q91iKCitUZrXom041ddJghbAkNXs9SwKPZ7
bNUpF6fSET3kh7/uRag25ZyXfgu5q0kkbPT6k+Gj8+ESkyB00zEjTN/DTTamDAlF
DTRJw5cojD2m0K+XYoubM11qJjLSa3Kkd5mGmtH/7cIpPQ12oXPm5VFgqIczNyDb
rr6+7Zk3fOqQSPWZXZ776WOFDHLuSblnDNmxU0d1y6+f/4GgPRBBqzSsyAVvpvjB
oagRpMYXojKgzPWJUdk2uCSLHiSh3W43cPpsj4P6IOJeJA2zwz2hnapyAofoRhai
LHkOJ1G2fIsDchpVl09gwo34OSxxLZQLXuOkZH2UZKxxP3QX8DsHLqN7/QjmvvOi
cyYC6Orx/tHJ7u9noL/uElbhrqUhcquWH3dsPyG5gCXKgSxiCVEXx6ci2JBUyFg0
ItvO0HKb9g7LSnTY5r8cx9FLzJEgDEZHYiyXbVu+gaGGyeuhmX59i2Qgx+ZszvQX
uPfJcdXW/erRzqFHVxOyc/bJtZRIii3sLUO1lL4srZ0dXOEX6h6Yu6GyYNqX6O3+
LRXkew2Fv+HEgfvK/fT6VBhEWpq+NXMEF64r2AMbVKFk121W+8OUB24K4vqOH6/f
ZO4vG7P/tr3WNcHgk8hdA8v++54dpjT0ONMWR3x5GgOLACDHzJfq537TY4bYIiZY
I+RaaR0oErCtiPlemWGwo54JzX4eFxTePxuYhpPtTWXGOIgHqlO/ZY92fExiXkXK
cCwgenfw7WwyVQA+gkMNJqna69rTluwF8DFI5nEi4j81fZCIiKLH8r9IiNZOMA6m
JyrQfyXl61ZAS3m0DHRo6y0gGmmF0tARKIh75+y9xGo1W7KMo3nsitbqNKzq5qFM
7gsV519AjBGQHVIW2Tu0XPaWkqq6/7hrcdt5uJGE/MDO54lUYFsl4UuBnszxle9E
xD1DdGiZrwKoie3s7Q6wrW4faE7uO+ypTFqUPh5NhOtODaozT5MLolii01NAa5Vg
zRDt5RPWWGjhV6/eEQWwewkY3hs9fz8Z3DUCMffVT3bX4QdzrI5cOfk2Z0MHyg/L
pSFJOAo/+IsfePZUF02kso2ez6mKAnEFxL5VGTtxCB0zL+K3JFoNWsIz+tGWoV89
dqvQ94Q32bKMwp09r510yFsL93ve2k4yFjr6ZUhxBH2PjmdloVjraIyF1nseiGRc
urz3ABoWAxnW/liGNs1e7sdxclcotKdXrt2vj97zzp/iEZK6G01wXFq5EB3pqYd4
/FcEqhPd1hKT1MenuMBBpLK8H+lijHmQM3gpfX4neOUgzeYTAIL8O+eVAp1KuZTE
TXpvMyk39wpKUc/7DJ8pwLYGNgcdwr2vsYWqCvD+V5zN9IwYEMRwRDlU4g3xDtou
+mrJdHjQNUqdEjId2wXoaoEWTYn+CTpUQ25ZwIeblkmt6u/m95XLUSLvabiUuagn
dfK/E1ENX1vqYm/re549ouJfaIw8WvK0N808WF327Qw2EQEdjajDW30MBVUPsmcp
8q3gGtsbp7/jJmpFInIqfjvW1BEDhLPXgnoajiyE03L9H9ZByk81ABmdgSYCy5lJ
KgrUQ1k771dwn7yDi5lBCZJDv2XOhi20rtdNEJWt05hW6BiKnQP9kmvcozgtaRQK
Ht2LUiqZ+RXwr8loBG7nTDGxiaRxe5EZ/i7P0bhSRD/DIIJtUcyTOGZTV+js8bRn
aEw5E9FPONvwKpjdFiYMNltEfljikyDZ727QAmVIAsZCKQH2I6MGbpBJ8p6u+uB4
/CKLZDksf9KOg1OB7SczUlGaGDl+SoyDopAGeiMOcQvuk5+GBeUpAHqXDPGFeoqY
bLJZgK1Z5kkr/wdud5UQ6LcDxN4Nmw6Vfs+Vd5bcQXNMIS7d9rrBp0qhmI3B8KiN
0MiqVQNkPuQPQTYqSjOCQTZ32lHiHZr3AqAxvtwCdKZ6BPxDWNIN19/gd+LHMtgn
OQTptOcCaQ47B9XgcVfUkUtPa8ww8J90ItpW8cg4wg104JFQEW+sP8T1EuiY4erG
swrLl8yOi0wNwMfifUY9EgytWVVGgOJxcWT/EIdbRH8Ik5cZBVA73pvNPW3ahMDH
s5Go4+e/oMVwSFs9gqVo191IzE7/RnVNjuQPfBCM1dPmRprkbtwdGQ2/cdw8TCyx
Q1I2LwK/zL20XXpG/LSLR3KgM9WFPtJbM/MnUhw1w3QQVfNfMQSIv69TJsxbuO1+
+A7zTRjxgpY/sWPX4qkvIZU4TABxGoustPmfOG7g4Ba0IsgtaSQyNWuW48n+ft14
sFfD3MktsLxemOLN55nzQYM5PiaV3D+nuFiSFpUH8FobfKrqAnHOeKoTfk5XfZvU
m5ybjzh7h/9AnodKYdWyU53Xx8g1JnR+eUvgWl8i5iXeWASwxTFJYKMu+PQu8M3X
qOja6eVXnhMlCdiPGAj0BVUoINojYndnC5xuvhx2alFg6J+rvdECMiJIk1QecBPp
ZnndiQM/+Hlho+yGWkIZdWoHjQJbPBnVcPIB4fn6DBcMLVEp9uZZ8Mm2HWhxjQeI
1FkYOWo8Zo1LjLYLHmCwgx7/ZWdpybitQEtCxdILvYBa+FsRi0S1R28kyhoo1dVw
zgLfPdGnRevgnffM2TSz9NkJGJM+THlLqlTv6DX5LTPiBTzO8+JhfQaTMt20MuoR
sTL99JQvsKES9edsekHyE+RVisdSGlvfcRneq1H4GPMcKXHcYc2z6Zev8hE6zX8Q
+FW1Ad01TROH/TFhfgJ5COtlz7dc+gNr0s9Oz8tWr/Wenl7Zsf31NxHV+kufjEHj
+En/qkU44QAh3nEJrQnTVAfTEiEJ9CV6fMlRuvX7ADarx/FSbce7yzVESh6JUS8c
Pu5aBQs2peALWj1nVMYev8AqCacBrIstC+nNx2r0fMTG9gYqxAMuRZZsVD6dc1vB
qTxhmHrPY6aL8IBzXqUJZ6QpWTjxTEMeO8QAnm2jrXhp30Y9wECc24gfg9Mvm+pv
lN9A78GswE6GYXafg1kjeK2CiBK+/IkzN42bX613LO6Rec9ZsKGuNJuANWTkJrke
0ZEaM6f7QbTUz/IY5hfQCh7bTNHzPE5s8cXuv2fHeSi8hwJGujoVebf0GN5/ub3p
onownNI38Hat/mZvqZvfVDLg8ljdNqkIoLN5JdOvOmPDJXscZ5H9GT3hyWR/eVUs
AZ+WwOcB0OJ0I+y/CJDC6pg/b35RSvo12hWjjIjH7Lwywq0uYNtzB+33q3Uares5
mnZ7WXWxOivk/BO3y2sU4IKHYO459gI4hHnlEN+LP42bFKdfYXcKplWVreV0ojnQ
5SwDXZWsNHNHKICUWnCB2MmbDnKfOmC+iOL3qezZqHtjTd0bVbdR6y9rDdIM6YDx
hB2TpZCP8olJcIn/i7x6kkMgtMt7TCS8hBtbud/FTn4B1pat5k7YjwLFSpOMdF/0
y1RLX8epFIy+opbT+e5gzmjWBq95Mrq+snOnNFaDvrJb3NEcr7UYkANk+oaWc15L
kHZcbOUIDOqIFP3zWN0oKBrf5BiN88ntS4upy9AW9RbuCUD8oqqcZGWUheEEKjLW
enX1AjVoKLdXVxEzeq8kxsEQmgmSl7bJU2x/DNyf+lbymObSxsRrga50skQ47wyb
bZJDZfsNITMza3GDJta3qCmJpANPJpKqVgKvPvg+miM2M9dZGFq5YmY5NXLe/0rY
VCqlcv8CPQkhH0bhSDGeMxvA85nKJHrKvndWlRqvzIwiXnKsoVjHwOg8RgX616Fo
1gCGhvJDMU0qerMIDH48I67OOMVSUZ/2yH14JTA/pheNPJXy1cbP7FJAAe/c+T8U
aFsID8JusAXQpyq2o+ro7Ifwp3MzezgAw5DS7HsvGDawHDNGrqtWtAwTuCcn/3dS
3k31cUcu2B5Ui14NIL/WKkeOfLSWpEGrdqaKFqxE6iNI1iEM2iPvrr0xwcRBLA7g
Rak4D1Z29lq6FOo0WDwI3KB0oYkWIXYztdjfM0UZcRc1OGO4IKx0S2fwtMzrfCBH
E5jyuht9rjqSIixV5vsmthlcUu94zgS30qR+AjSlvDOkEnh1rYboVAMs/rzSutA4
i7viLR1hGCKNyZJZFPbwgNMCOXlhxz3e0S0w9oqDfduiFc+374eP0boRGXlKBWbs
goC0dlJNixu55EQ2P+YWPTOArXB+Bja23eqMvXbAeXG3wHpp9MrgVuIeTp1g/Bvd
Jy7GsQJvk+nyNmdXdfIxVq382nOOM0yzxZVS2nTAtr420WE8odbuO2WferAe4zhV
1S/jpo0zVbzZZb1Y0Ntl83iU6v80jG9AhwahO+1Ijdw+6u/E6mW6P3QZ2fIuvlbH
hhiWOJEJS/0PsH0VoQP27V6IXhr8pCGK0plfHYI8PwopL2NzEdcz0FULw5mtyFfE
NVOkSHW4w2R9zqaig4XgWLEcWUjHo7uKlmatC4fV8tycJ7OJasCX0URUBoQuzKwD
b+T9/aZRMSd6vdR5PD51YukSCiPRjoe3uK4ZKdmjuD4dMDTFCsyweYh4TANskNER
O+n/m3FP9jA+9Xzr6i6JwcHdKMPPajFaWRKSchrwjJ+3ka7Z9jqXde4U062bZUL7
FM+HvKn9GgmMN9pi+REb5Il5YLfc6mKg5MKtztrx44JotTp1jHQg9llIeMYdBxN0
VkCqdiaKZTEYCsvt/aZv/Wm20txYJ5Z6OtFzqfb/ZS0RguqplvAqqXm1a+z/cDTN
GPTfDSCLjY5qZrkwsAKr5VnxOLCgksNGC1ODymJ0Bge6sLXxNxsT1outyhrB8x+l
eo47fJbb6lmyQcjYSgclz+T76CAIaJ0kcd8yAbsnp1AadoAggcxqpw4ABY6vYHz+
U6YIWeU2MuJ84iyNY3Noktt2MYpat9pLVky5eS3CH5UD2yUoV1sloqV1DTbU40w5
z3L+sgopkpnpTFRyDtRtDLpuJpQs4TDUjTnTIvLk7FxCAFDpdpuwJEd6JxMKUByq
Jyxq+oYky0mSSnMQl+vvY8wXfIy8JCaMlkyoCpyxmEtmyFbKzcrd/XTRKKUMEE2f
W/ZgYTuMsWLdRsXG73lsapVzQ8Qj3ON92mZEp3coGkdofdV5zUphFodLkJU0V3iH
NC5dH3gTq9//2fiOh7jAlXTcd4O8k5oZMmAHN3dPyNe51zji2h8m54ZIL9KyHVUP
FHaWyuAOw0n/oA7QBQ39DusPGJ1ns6+0T5rNLiH6/Ny5aOFr2YpIYk3Rl5dHj7eF
c8LNYi0SMP/ml+L4uOJnTh3kJI18oW2dMQjxKdwzZuepSiHzOxrjO03m1lzsXwFC
u30f401J4jb/ujeegKStVXAyqOFT0ZSLa6V2n2fJ2yL9WTGy00pF+KURXLUeAMOJ
Lx54MGjZsHa5cGEEoZNmoPS8gQJBOqjL6PI7XQ5fGXAn8OHObFf1lC9d3c+TzglC
Jm5cDhyf5+3rJznSl9EMSQLzApRjBVJKpIA+XbwYprhpriXLWHOEaCsDMGDnFp+B
kAVJYbf/YgqC/Jpg8e+VqFA7MEKMqgl1X0B+QC2VGJtFL4WtzTWNHvH+7FIQ5zqQ
dnMMDqg7/a+IHRsXjGzxoJJHUjJd3xshFz3falwLBLynscq3/ot/2iEEUahc7gHV
/BjKQm32TxemeLeXJJjCYEQYSIIa+N3adLelSgxYPaYUOa2Q75DTSLlktAXt9wp5
SzWKWsitO2UFJGhdYm1t4Rwpcwl3VR8Vy01rUsIC1JAl/48O26uiCC5LEXLsssPT
tbY9rrNinWWJI3q5agqNJlQnWPlRD40A5eDD3hONxMlXCoJqC/XeADATC91n6Fq0
q97F330ieLQ6GJbY+EqLgK6bLIbMUVZ70h319sS64hIlgfpZ0rTZo5YqfDooYk/Z
hETWq0xJUw7VVAJSS0ZX+BuSTJ9KZ6KuVEmdFzuVlk0axQXoJSpHJWPIR+Be7ivE
5b1zfTBErK6PFIRrUBLyXegq4l6VrRQwF8NgiXCd2tQ4mk8pFTnVK2XSGIxr0y6N
Ab0cTA0ZnfwDeQcqeKWUFO0OwKSU3vo1ELjVVxZQqRn3VKDjiBS/UxXWGrOORwJN
KNuBeExldE0aFxxI8Gngyk/ozH3ychKvddmZaMLoZHkTQ0OH0ouDVhGuvRq1K6Yz
jyGSnYGLHthqxZ0vcfm+vtDjMYQv3ha+Ia7+u18/kVEfyyewERptn31MwAy3C8wQ
F9iMsMSbI0al7NWjEsvbgXkt7wIVdhdxLi/YU+U4gq+3IzfXmsbVPaSOiuPsY5eL
2zKJrIQ2YEJIAnZo8JGUXSbdIYmDWWgEIeap5STbrNEbM3s7txX4+M0hA64xzKxA
cyi8fIrHTRrshXpR0mEUaItJoSyPlmup/CSzo2FqR002G5UkxqIpHtiB4AgMWOjR
G4mYcDS/VL17FoWBVVwlBG2PF3BtBaZ/NsI5kNTwKFv3SvhxkD+7EH7goLoJFWeI
sGpZLYor02xwXd2bIYTfGZu35TIROCWGG8KeHm99UorMqrVrrsd7Zt8W/OTtnusj
0QOWrTFj8GXRyu7K3PQ7Ir7HknK5D7amscajo8+35vkh4zW4ogjLa3jeMj4Wqmj2
VFhOy/Xxs2Z3hsd3lceHQ6sb8Vh2lMr1D259AAFCT0FU/lDYM20f0B3K0n1reE0w
r5FwQuo/LAppPCfEdRiYP0eIBx9pVyM6XVWJfdpSTwtegM3NR4bnKgHdWt/RBiEy
nOQfYSjszo6xiu5yKLZDUmxXr7ZSFFqfEFokd3CQQo5WNyT3asgNxIIEcxSzbiDJ
SnUwGGV/+co25om385G1x5huw1DBUQFt3nUUUqhnSJN0TqVUORDa5unwPcmhFgZR
viAoXsoe+rIAdKWeyXWii/lM/rq4sFqJwZQedvZkD/k/KamB6hPBqm9bCZ+g6fzB
IANJh3fHk4MJYrN0UvGjqIJHeO2+QRM2h6qER/C+1D7p8VxLjrwdxoBjpTbEl/14
+DXJYYzFx49jPnUGsEOPl2Q0tXzq71jcKfBqLwdGeSRgQfyWmNlYelZK+wIpOiW1
2Aw0WQrdQM447oICyCMTYP1qIx8abdimc6K5GxUc6giqX4SsKDGMmHsH8390OIY2
DVEN7O5LDSk55U8LuTA65+whFE7dcx4TK7JoAWhUlEZAjj2E/N+qstiFHRl36Li/
EYA20Kx7G4x+WUdiBE8cKpUKCXGbDJhLud9y0wzijLqLZ4gW92L/At3B23iwheJQ
WrP9vjE8HsbEWK+CCVreZltzMPxx8H8yXOHuOEE3GoqiNCtYE2BOM5A6AmssQb/A
56kWCyzDaoGwGpoeSz6W8blnExU/ZR5jbQVj4evYDEqFv6NqnhbfBPPpTMPetGSe
HUyt5Rw1gCoHJ7tTZpQG6KUxURX2bCk6jL1vLKGW118ZIEitzj5Y0zgzKhb24pTd
Hu3M6e6rfnjDw2uffVwQVDuChT9v2hflD4KQi0TTQnN3+ym0ZsXPdSlb4Hjaf0Aa
LxBqSxTTa8DeqSkjLiiEFiV1aDM4JAntl+uVkP+7CfCETtUKnGBT3O79L48epY9z
a779NAm3uIKqSOrLMWGCTZ/xbgE3w6bRjcWeDgFOBC1i1Ru0vinR4TAqwi4yFYYF
4QS1oLmxyRtGkcLMWfOx7cpGtZTx1zALMb6r8m9TRqVdElhkgS50DncqIf7wGK1Z
4aYyalmYfwYb5ifdRMi292ZxzeHlmddaalb8lAnUcrCl1YXakN0Zxun3CWO1wnI/
iIML8VjQJdNjX9Vddl91cr/IStTPzJkFXh4wDd6EOePxosbNfKr4CC2xhOGM2u06
fZHOFTcZEvwChbQVss6Z7CrBBjGKacpCeumTyeM6y+ZxakYEY+X8CZKy5OtGCEHN
BwXjkySC85QddyT5/a1YpSvK8v+sZ0U1KOKvyO7zZ86V2a6eGPqcQwbVBii5k9Vu
8p66XSZBZP35vwHOJ6IsNL+PX7v/JtIoXH1qXPcnRKk5uSubp63VbkkcZVhkY8vc
l/3sK1ni5TU5Kx5089vXTP5RKP2IapE47DDXIwNPKna1De6BZteJ8JNAXb5AnHa3
ziX/s1Gf5wVcm0df5TyD+FjStweD5jEXV5cJo1Tu+a7dzpJgWMyPh/U12yNW1obq
jJAasH6rfnafrrBmCZ8DU0Ign6DwpnG252VF3/9uU9cGk+5yOE/psA+SpQbouEop
03MYb1mN3bQVuxWURrk7sGRm1HY87XL+RVqVDdBlgPoRcPxI/VzMqsXNTFiESYZb
1q3O7XDkVhXc+w07E/KKI8oCxajLqNSxA7l+mZPeK0O6YwzCnthaU1MwXe8VN3Wq
B4awN36spBGzmZq+ZVKEpvX2qqKCbIGmCQnftbh4CrCVoM8pmOyPyqDbspDOVgdm
VvoUb9aoXKembQTmavmgOWRGze6n/aKHkeUxOUKwvrMlKntQ4TLO/i8aSmMkW4X9
2lIGHGVK4KBUKZhfbNNjBewhVaZSLVd91Gtxs+gbEr0t2kBug5vO8MyRQj7zx2Db
l5TRLOUt5TU3zxjc9thnG8Ni8KHAMe+O0awADdcyrx1gXl7/0KKlkX7LwlBqNTpI
Dl7kJLJD8DFB8EMcW6zXvyZ88KiT8NicF84dhCvEE1H7xEz5P9GQfrDfmqGcAUyq
7oQXWIMRS9jt8U2lTohf8DTjZqxB4qswrpnJ0oM1HhT4O2r4sh0pE4xCz8Cvs6Lg
iVpyicyZKwYkPADCYEXawcB/SULYV1koxP5WdBZ0QnpIGPleWDsK8tzsxid8Jm4A
Id1WqPo3q+QI4XiBF5yEWbZvdnRhzcyKi6Ub40/5LU4iQMuYZ5Jqw/uU0HDJSbG9
Okusbc57xMeJakrlJ5+ghqMJo1Iv8AoMxMGaygFoGX8wcU2hMzPgM9L+rs8+arH1
jEoFFtwjat6v24weC7HxV3relznB9udnSPCOoGMguWbL197gvE/LPVytSufEH4gv
53Aqxzjioib3UEmcv3J5uYFM68r0T0j4z7Vi6iYSIIXqN3dFOhyNEJJpU0fJD4Hx
79bUogi2K2wikYHOKjO/1dNwp+Zm6rSKTsQtH9pinGmeST1qjizc9H7piQNjbZOf
UxNRCHbr24ePQ1NkvFXkTQ3dnhnFDQKS4ul7rncuUXd3sRiADRsvOkYInVkqzUIG
uAiK6Xs0/ukF7COMrJLme54Ym5NdwSjqt9QYAqsCjF2R+CWyJ+Z0URISGJW713so
CnWINqmoX3ZLjQPgDb0qXf1ML5dKw1WsShhaaQ9M9N/ZOexboThFt+8+GRVO4E3j
kgRPgIS+YoALq7Uv0plo6xjnYdxL6qR9LUFOOJ9vxtwnG51EVURXaI8Kd1iSUvB/
ivxPBOhBPBA3qlL1W/1iLDMJe9FymgjuL3NsD/kAQpopHNVp53CkyO2Kcf4XuZND
5UCfHNPR5fb+SkyGkXxE0Bj8jn18K/YxxzCqh5b2jBzqPk1ZXyrVY3H8wbk7fF1I
c2Kp/yz/c//IMVKW2qdHheKHBlSgd/VGMyBO3KSvWsfuUpJVNarIBrXl1Z8CZe8j
RYtYqPuiPZdvSGwivKyzfSbK1w6l2gtr5Ksg9NL5syHltMD14yw/Y9DvJ+GIjz7v
g2aznk2rUSFB70a3ARfh1naheFubZuaBFwJ05fEaaKXOK4MsRdT+oB/LiBE33hQ4
bE9Wj1xAtnVeRjIvyMKlpYi3/V/vD+9Lsfp9+eIymwrWA5axKX0w9a8toA/FPI5A
3Jsuz8YDHZYsT/E9xHtGOV4CMAnmo6ODb3NMbYIrrjFx472yuSj6ghRHEInFb9fT
W2tpvVg4QAMGCOkTjlWPn/0SnTE3G0GLlm56LDukHaxhzERh/pzyFas2HnSZpqk3
byGAPmFy+zNN6L2JG+Js8ISlMUnkltG6dptxFnD3KY9av3Cvj1sHiat7X0nB9nbi
RPEtH5AEOYkVkJ69LtAuy7DVd7nz4Uyo0TQ5UCAtuJLn4YFpRkhpEMNom5o11olQ
itF/6WxkbGad5Z1CxsnmJwPRL2f/+StZcp5m7sMCoeI3390nfVUT+sDy8l4WIah6
fQLm31RpBHbPo5TgH0FaNbKSSaqxUXE/R+ubBgWhYwIyaKZXaHQx6FX/gmDMeVal
f4Apd4HIF1NfgY4xzfFWOeUEBdaOgBfpAZprBqa8I545d1xKrkmkYS/8d5WooqSH
4E1+JJUTvhmltPlRuikKAjkKtmsHvPyGVCSAEryAr0BMu31M5AxqcBpAC5hpnlaq
oc8z2xxcW1F0CSbUajr33vaZRhI+h8JO6WCrQjb45NBlRI/Z35McUv0vnzBvvvNG
fxiLijlSZGDQeK2cY0ajYUd5GYB7Tddjs6lfeS4dsbE9jdADPEz6NLWdgHssd3AZ
pJvRZYgL9pEgMjEhc7UXmQyhlqCUtN1TWPcvCNcrGYuNCqjWunDL4liENQgSWarE
RCB/vfFq0f/kTRNkWJMLAtZXLjMOkOEGKV7EFzY77eFzBr2pbFUUO1tmSL3zLAaj
hEktAkUdbTMC9OwQDe0wOolHKcWtHpbZn2lZlo4TX5BAmVdqRYLyVC2+QSG0MhJR
eBtgWYw0m4T52EZDSv7ZJS5kkoUeldJBjlQqdCIpT0U3kijuPehqkUdaztow/JfO
INrA7PHWCfGj4VrtO2LtblG1PIubWb4bpf1Xj5uP9ozolYpF7bcALkSWp/6coeoV
qdBNE33SNYKdTuvH/OHOy9oHidVz79LD+x/3dXMXDn5aqhXu/p7e8ggASBDk9QWo
7OdUi9r+Zm11jfImzTw3DH98S5XDxBCRROy21vYUQpGq9Fn2hhTRenXjJko0bvu4
Obtdby/87prVFV0MMPKigpTgJAbZv70OqJbInbkzRgYWficMvYzXa5BmqC9ZBXCH
IYIgHtaQ/ERsx0tcV5aWaApkOuED17HaARYKqv1oOpo+7vePutfMCOh1Ldw9hN1b
eYY53Jg17mbm7+sTs42ex6mWS7/K/hiXO4c6LtOgXseso2VSZFPNQM6p1KKHZD29
cXGdhJpw6g+TY/LKlLs/C93AE1w3DAMzYo3dlCLxlz1pwnN2OldpILZR2WBvibvJ
Ghn4daD3J4ZQXeNQy1JVGtJdCB3zF1kq/us0T4JycNE36Ov9GZlkEuc0kxK+QQGN
d+h2XfxV78UnBZJ4Wd4pjfK1IpaWjVQFxw6jUIK2FC4n2BMTvXV5Z95UKKooXf/B
5vObxCpJaa8nY3aV319P/3IqL9gAC0iD+Vva6h6tjwV5+Fd6EkCHZ80YSu2os4Ff
Gi0r/hHapqkwyNNhkoh7BJd+eQwqHtqIQkoFLEciEObeATtv8vFpVPApkKlvDBl6
UqoabOyP57uaegXkTjpMltkX8NGtB5Q2Kvoyr8e0ajOTOq0vV0tph98X1P7/y9SB
T8G8N8WgS9Ra9ExNyIIZApdPiatdxI+FZ02BOISeRgGddvCqcPzftlBY38jqTXID
zSYOpbvRGBzV3+fI4e4MRLCpTB0FEVFPEkcIq7JPJIqcGBqTOiOpaDxoTrobgnus
WoYocWurccB+buyJV/Z0+4OybQkBhITkragUI6IRwOXyEAwasiGIOpISs4AwgDpA
whztm6rYCZxQ1xYeL2AYaiNCR9OYekBNvt2RvN4icnt1y1njiFbFnQrIbm7kBMUH
USBgY/K4c2YAGQYp5PcC5rk9j8qu3/UKFB6J+r9fZCxBb5EmhoQkLqSF1vC9ebnH
Ya72UWpVmh25AF76r81KuTYY9bheKUQFIch7IvpiG4sVBC77hUL06dGhQTkCieJT
kglu57ZdEy0/HC7zbeeZCaE39Bwt7TCKFZwju5X4KQE9Kfzk2HkXB0p7OwX2VXdp
w048UsLwu608YrLGRINKEc+LBxvSogRG8J0Hh/XJa3WhilRlkwjW/JVtZSzKvvPK
vzcGHSwlvIL2le/bcrPL78wfcQw4HeMKVAc8Ak4oi3Hgc+OPWS+mq9WfaVXb04jh
XL5yJJmHbUMwce3ifj4DCC3Wi49YLpEw5V82Nf2lxVAOCUkh6nQsouAhR4djzFcG
G2zh0cZ9fDh248CvRdHgGu43pBDiTWNTFNjcOnh33eRcOyuXRra0qqilKQtRJXpR
VmMmoqtOcBzQEm7Oib1ziRkrTVQ8OJLFHIya+2iOHrTycnA5z7dcAx7ruFUq9gFI
PH4YWm0IGxRvREz1octbDZ7P988G24Oh9D8B/fS2pZuPi3eP4qzVULqV/XpVXreb
VvCfO9nrEsI2imNxNYS27Lt4lcFr5JkaFUjfwUZPsz/YHBLaIh2W9MeFNp31nrDe
WqcnDIX7wIHTMEY2ywvhGh19WfHAVXFXtKTyrXk31pVCG68sG9ECX9MrO48uCrLh
qzqaa/0v61tPQQeXpgqo4IchStLXoUPILFxN2hDgPpDOFpfu+pf9KJYt7Rlm8Qui
TsAmuMh77cqjy+ZBGNaRdT5SqY3rJAZEO+2ZgVTRBS5Bm6wAI03gn/6hs9oyJuNG
h7GGMyZ5Rga/M6c65DkBV2KoFyt9BCrCscEIgk3/oT9yh38sKpwFPpTLiBrFrhjW
LLeGe5axvQWqJr88q8J9DSFJhghl95Za6xnCvOVuHhxCb75abstrkamwDkrHm77G
y4WioEJD57VJMrakZeLNLuJoZfF4VNuv5LsqcY1jeD0rQucojEswx8X3quJFzTSk
V1W0AzLbxaXTeRqTWGHyFNJc2UoFDdIFIeunNNg00Sa/wwlD+xgZU601qs3QFtrQ
2XFjl6/fg7YMOBNzOnvx1L8M9wk+HmWls8kwW2nTE27UyByHO31ELFOgZBiqzQvN
yDw1xuNpfyUeu0IyNZpr02krynCq1YeB+SoifobN8+cV3CH9WhYylvP7B2rxgBDX
D5CPgd5cGG/vcF6hIhbI+rk0qg4CkLQk6y0RGEmpF29OjXFQatwDwbfXkHHNLwvj
DaAAM8aeO6zxMSWF9fk4jpHBU8mw6Hj5w/+JYriNEGcZd+QkCzQgaQ10oFUENkwO
eEz0iP4f4kpt3bduJ4+/SCZdPAkLPIH5g+COlqrE7i8o9v9n8j2qJboE4hOuw7zK
/XNykGtnIn82aF9uv+KDTwI1mok2jiTNI5XQkn6BAFFz2tjTNwAIthXzHvUExaRY
2HK56abpaav6mBPB7oDjR4pMtZrcGzgd099p6RZFEZqs5u2AjZGrCpVET/zV0zsX
lYvjW/KlRQOu8vTTUTest1aucg3rPf/e2XAuZzcLJF173APTxsfFUriRsMPkfg27
2EforEICAJ0xwuxIqt2//UTp+7mzfh31wCUDZlq5IviCq6zL3QTDM6danRthXwvS
NcFXOWtPhkp1NV5RHUpdDEjGI0i1P4AzbQe0yiz6f4E0EuCTARVkHDDwdPqkvnRH
RbAqLzyUZ3DEbiZI9vRyK6/yzqFU1em6UIEDaqP7ngwX09PfiwrPx2AVLIZ6T3Vn
ThYlX3qp5FuAL6cPRbdPvkubfjq0OiO2MM73y3q5eR/dHuo31hadpjX50Jp5nxiU
s5riknkgoh4VvRuFwoRf0wyNIBcLjGLjkMJVjzcBKoQ15O2+db9rY5vKIrGcSe9y
YKkcO2expp2fBw4E59w2HKWfbuKCdpg2N+kCH0x0E1sk/J8CwlsxB8kVtF8SBzNz
s20QtGLinOZHwanZtZ8fUIoxm6QaJb5kcB7kLy6gqGpcegSRUkOBdmtS7+xmn+Ch
NnSnwG3VHqxk5W6As74rLsLyDFuD1UXDnxUp4OYErWEKR/hQ4A3Li+urlbtDLw4w
1ysIIvhgzCbgxBaG/M1iK6Fxhl3n26Tdfe5JtNLyuudHjoiR1uMfHFHYcHNRNd5f
yHWHUvS1OcL/xsubaHrxWyc+576edYbjX+hZZUTnnaUk+nITu3KeGJR4eBBNsriv
RPMkm1nSET78Wqjt5BGujrtYNSLpq2A+Eg8DNvebg2RycjjzL0wXL5OprPvYgm6t
yIC6yQPoXQ5niFjLLOzj4uf2C3MlHKgbG7QZUawXcnwOo6liq2AprYPtXr+416Oa
+C2Tcu2uHE7kfxunF9D81a8dM6vM/qJOfBOaUTtl8hY1IAhA6UjIPNCRoneXVFh0
8aeycTXbdAMY1fS90NVrIgm+TeLmV0GJnvcjsnxUNe9V+0MSh3nH1VvSDARYIxaD
s4PIxh1lhn9V/5BP5AOFIyvM8azeJxNaN0n63GrEn9NaCSuzHGEvcEaVpiGudv6F
IVC57u3uZsWCKwjjp22T/ZelQ1KLe2Rv4CxqhWfXKQCC4H7xA0YNHBJy925zpLTt
crD8zm7sB7Cv6r+NlmLoLQnkpvBbQnLRn7nvJRQpLpXlT0DBS72SQwOHQ7a9tP1g
e7dI71pcrN2jhaaVQ+Xemw0cvrWiVStrfNp7tc8OiWZBniBnboyARmgGO1MQ+3uA
ksSTdXiTLf4itrZA35ckscLXRUi33v0nZMz5rPPyaWn49yUpTltqGCCHMkTpJvS3
QapD4rHVg9JJBISjzg9bDe515iAZTpYoY0mig+wlj9JQNdF272das6Y8pdZiuGHj
ZY4W2SeXVMOmky4n/mADoA4UMjtyi/IkIAVGMS+HoC7qoITwZIAtHd+En3coS6kL
j6ndYNuNaIaJ9FJlC8Y9p1a+RZLaUA3RGUTM0Yr9DhXtmWNf1OdyiG7TWhm0ySSS
CanDgnskItbMe7XcAHPKSzdaG8SohZak4hCL5Q+qCx19pX5YmiLkbDvnT+eRI64z
x246byxldJktHQM4U45gXnhCrtZvx7daoOrBjkLYscryuu6ATsZHpA7wDFBWKhDu
wsak4Do3oB9UmcZJNKJBLjq5JWaC/td9nriNArg9m9B4qT+V0PMwYXyDgIOuHTQg
Rcb1usWhuQ2I/jQRZfkP1BPxupXr06GM0Wr4YK39LuQmpuQmxqMg5FcUoWbdsRj4
x/DOvK9TJEw/AITGB8un36hjNaphzfJ+0E6sjXSHeXorwTmefnnqdd9iF8NbQycf
MkbpeITzH8PBzWXzCKFnEeOyrCU6BQkdOKmgsWHookDDtUG/iADCrR3qCBIVuXn8
xpRqpdyeIudK4T1wNGyUfezMRZzdRIe9CmpXQkPkkB5bIuHXNR1LRqR+1Z15Qdi4
mVYlcmpv5Me3hc9v4DiPHY6qtRfsg8IPy2e34zuVFEKDHnXfPVDa+pzh6Mg6Aesy
VZAovGJFZGNhjEBNfQfZp+G9Nh2sHoGCmX1bLd0os6JEvr99YiWmNe8Wyj2Ds+st
46XkkLvONuy69d3meZnzNU0810Em3cbGw9fPEnCsdeSaI3xuezt55zJpXiwdE0G5
p8gc4KWfGDUimRP9cmQx6WRjK0d9c0X1ugftovifh3SuUrxa8Sv/r8279xcYlQrO
1PziJVv2Vmn2lDkuye6182Ql57mC0Jfk1K0C6SNG1Ok8YG2gXKkEe++42pRC2L/x
am1G1AjGO2ismA983nLaDZbfea7wIT3rcQ9FnsO08Bt2ej60e97ygfK1oXiB6FcL
EFKb/LSeKpPL/SSQOXwVcuUUQM98TMGvmZGtQihRL6rdqOuAvuvQ/RX8j37oL5Gf
6NiIbjaZ5uyVaFq96CvP+Xj9ELiHrx/x+X//Feq9EemXYF7W3QC6Khco4lURUymB
IHIW9IXDqbk89PYicm5gqp0p5O1j5MvoBFmPUdcrM5rmc5Njz4HrKFv10V8bDGH8
mtJ7PC9Hev+JwBb3szo9wfrFeHknmYml+8XN6so3NjzCL0CvAM6gl2icFJOIBiNc
w1GWBjLCuRXZzJeSc3b2kYEdxCVa+fUGyj04ASfwq3lvkoGwMG4MYm1bQraSLzcp
7RuH898uUbycBHeBjaq/3nntq9jCCkG2EdgGkDcg6Uhw4xLJZWS+kI31mzneLAjg
j8rqiNRYdsAhZF8QVZY/Mm41lRqpN7BYVHKVbJFU4IZ3D27bUtxgHJcc2ay9PSIa
QtOeU8GQjIC0C0NZk7YMHKKDfCBJofL1o+MA9znz+u/nvkTgm6nUD4ySa7innmCU
/f0ikBTIkTnlrQjE9Kcb2gRl9IvFznDO09fqcplsVurHYQhy1xmg4hvn4vrLGopS
LOevoegL6CLrOJZN95kUj1vRnMMESiN/aK3VNQMhW/Z6prRJQkaXKk8U8NszYoe9
uZeodneRs8QVAlEA05m/0FfoTE78XQTBMNwwvhXbVFyBEHttZmL4v9G4AuzkxTka
H8fVlrCmTA0KkW1/HsKqgQ+Y8elFyioB7BendZ4R8TDv8zIt9Lw/MIwmUzyJr5DG
J7rFfPPas34f7klnd6sYeI0VZtpOtsTSIymlIi5SId0WN71bkLH6fkZRVG+6SE6Q
8VyI8xGzQdWyZxSaG633p+RJHCpQ/Rt0coE04k3PmP2wr/5VEK3MPUpXKxVeqjJ4
jpUcDLmOmsMpaIQqA5YIDypWV/w/Qad36yUt0elwyxZzENN3qs5qnaSRqI/JBncI
9NFb41sIG4hutsD5BJBh9mr/0vKNxEaLVTBjfC1WMmfswxgTmwcD0sSoxRC3VAuG
94LJLy+/9Go8CdhMDbvqsel4DCmDXk/yrUc6ag9vbTZI6hfh4+9j1ktrThvgJnWk
8F1b7PackQvjUAaKazwHR8yYPEiESIlCx6sUuwGuFXp64FYlss74W+vT9dliXDgj
Dv1bbIkiQ28+ejTClZfnI1yjJeYw67DiYTYA9FgmtPZdepFFL/bk8wAws4P+GBb9
DC/mxrdujEWK0YGQvf6WM2E1dCEt8KEOk03CUf4FUS5Ckn790Vbm36qoX8xVZCGc
Clj6hXiwPHviSLq2yUqV+FwWpaXV0J9KX3kuGwdDOCwYqGLZZLHArrg4yA/pzY0s
BBU7qnACtSkllqqDiNG6jChutAAerJ8ldeMb+u5HIE3PjgjUQjksScq5wVl49GNj
y+f1yhCtu2VF5zk7Tr+XiLuIuBJEEt16hw3V5Ns50joNu0wQD3xA0S9aMPrY4ldY
5y8c6atPhBLlQ3o3C4PldJytAAEOxnbtQ2MPIKfZOkE3LDcaJb3rGywEKd+JoBev
F12O5tB7Z4/3n1Ow+5Fc8DfE8ripHdB5eq9lBuRdcuZ1+AfFDMEpRQhyAOr894pL
wQxCXPfvim35yvCsxqdvf14fu4tYMvuPC0IUCKmtRBhj8HsURW4j7F2lR5ahfXQJ
z4IU2A7pS+c8bQypmuuuFIWPBSnaVhV1ptCmeOxLamZGE+aV6My9KFsj10Zlc476
mVzeYXGiE1tGCaWl3XlgtslvZvb/tvJgRINOZ+kQ6+zBL+6JmbPA7zZQBvMn57ho
tfd//nevwzLeS4hQanVZxzknC8MJQ7x3upIk0hk48m8svkHQGBjgBwGW2LUjlbNw
KuIZvFIddFG/1l90fIgH5IyG9iA/q95MDJ4hqjJ8t2h+SkWOPKv5fcbCaOSZfPv6
xS/EHrie8TkPLj0BQ1/YjeCUmVu1xKS8LJsWdWUJBzucPmRjsWgDyO25UPky6gJw
P86AWHGYl+l8CGUdc+KFODpN2jg+sHNUeIuTcmroIyy+SgDz0nXIHRvwzJ66r/Im
wAaaUHo5LI3HCJaVoL5MH5oK+PAQY443fERF4ydPkzIdm06GwWQ/qLByzRdhaaUe
vxyMCq9WC/7pErKxvDw1VQXyXR8cY2AFwg9jI/m2eN+q6YVCoUHLibSPCDr3akGn
ooTOpWVPZ2SdFuvQeW6c+GieN59m8b5RC1ttK7sZNyBF5Nw6VdLIxpkbanMHhTvD
W22RIDCx6iwqPXVGJBt3Ux41nU35CHAltQ3FM/mnGhzGWcg3RiVF5WDmVpFYbD0e
JkaKQkMYp2Rfc6konHaK1jbz1jEEXIZjXe3kzJM79Jb2w1VsUiKMcdIL8suZjVKW
6XgVL9sb6mTtnq4m3pCv7nVhvDOU2HTvx5SjSzNeznFbU3d4qTvjPRh7PG/dwhGG
hUww/OHtkoIevRShwtpq11LuFQkuFnNbR96tXw6dlMY1l5nxBSBadCtNpXDTMX01
H7u8tEDEhIU0PnMF38T5cWCp8xTT2f2pqOhgGOxdTwFycJMJVj2QQRt+752vIHp9
50FSZeotxNS4n9eo/lp8tGALnWzufvSuxjo2MSFjNyg2wIxicCITQLqYyQ0EO4DN
bcrt83bsKMetFsGSVcsObC9Kdvq6YURagKm9X6WNGGMkrtTJUTVyMLbHInPcaXBr
ezNJycNenZX8IKG4EzHko0qJbee8cdEm68ZkTPj4eY9DJ8AF+s4F7GhP67SaGr62
teaNIvANCLQ63hQyip0crJQV/1PCUa28ThQRSGET7InVPrXFQHmSXENTE1ZMRYZq
PE2Hdd6z+dFfsl5Kka44Ylf4SPTOZvcaaQS6OXULzvUhaVR1x7QLHa+k1XWZ+Qa5
5xLHuEroC9SCWtEQcxtTY/CTf+1oCe178OD2ZqYCd7zMITSeaLJKISn8d1910Zx3
qsc/yIrZgtExZhR16Do7iIG2zGp2jfNxWKIQDNZSJ0D38M2NyYUgx3ANfro2HcCz
DtcILWmvHPVb3EbHKc02PYcEn1D6wv68sU4jtbrVwI78ztPo6gBRFlAD41mqNmu5
jqjaoIQafrdOuVvkJ6IAhCyPEJW8r6vGj/48n8N0BAbupGzjI+H7hTJczE33DIkZ
ZY0QCSYt8LJYtliRXOsUvj6A3ZjBkiFfHZi0OsvMozyvOcus5QS7vm7L+uFyltpf
L+liJ25zFlGLsfoP7by7YJ9blhfYUtoEi5Ucv0yOZOTbfWxXHoll3iKwNOY1GN6k
SLDbGgiaYbdsvCltpKuvWLeM7VyB6bIGJPIobB9HUJLhmmXQjwu1CDDU/buebUwB
E63zl/q8WcqikfENPN0FI86e149HLt2Mq1L1/zxVFxIl/2KxPN0o8pxvOy73Gopa
H6Pqmb6zxSi+Kdxz22n1QFPoIsIi3qUmQzWIDKQotj0LckfZblbbr7bMfARyP9qO
hJFT7iHYRMt6nBStu1BTM5qY4wSiLDInWm6rDpXOhUinrMWTRzPpb9nj4ZU10xzh
S+b7Xt+SHOnz+wzzt5on9xwkTck71Ol9/2NXKWi6Ko7Bwathijt5dgXKVSWBlxsJ
wMKK9q/IBQt8FbnAez9sbfe3DbNeEX9yKgj5wKhc8cH5NHW1s4k64LWESmK2EfHH
PKQUSewGOX1khs4fTcHgIPzhibBBotSwRBi77SWyJZwy/JaMzjkYaRsMj1G/vyQp
9q1+pke9LkaZ+2lNOBOa5mE1C1thWBkkFfTckePMx4aYphC4qBUzTzpq8FYo6iV7
5XUNVGnvrDseqvPCrVaRn6xXW0/aH94K3RpP4DcceSWHCCFwJK14HnDognKbdf3C
P0ufQbWsRPQ9+45sfoSD32T6xf6T8yH2yJ/AjuluacO/QxbjAPCIZ2sJ3n/OLTwD
G2xLfHudhyJp3K7slDWzuMONcbVOrZsPOhXdkxFakw12kMFrshQki+bk/FVN4663
qPI4zbjcnZ5t+QNdWxumaFr3z+c0yHvFOui7hmion8gOyVXpyv8elAO+GVR0mX2X
v7kzwozlZ9krADDqqZShZTZAhCXzDMjTrDugMGLSelxRJcLoLByqIwXa4fUuBKZ9
/8RiNAOTpM8WXEtk0hVXwaJXhnRuIYMtdLCL905trNDG+frBevfQuWRSU48CroQm
g2nuXAQaMnArrvmw/xoKbdTuM2n2VN0m+fn7mRE7cxkjby1ZSchrqRGR+mxsGCxn
UwJ/IAxzeHiC/9S5h9/vVyp+QAoGBjuReKb6Bz5KGuTAzbCsGPfZM/WVpTMGL8qg
xsoXN+IV/UsxlBEzL8JxFL68bg7c8MnCAXyktpiQfcvbqGxZUZT4LTujluRZlh2F
I13adhNvq6TyfIp597Kl77CoxydwShHIeaZnQm3AtIS3KdqeP88A6qohkBsFvQtv
cLeNZhK/mM3K9mM/h6Cid2v7ewDe4Gzr5+EzUB0YScwaOHzT+xguDwo3EnAZTgg7
9w7muXDrdrBGsPSZEbt49ILm7G8oyNw8SiDMXLgGCsK66riMRAFoR0wMOqogfi4b
BC8Qqs8HPWVgAYZuJlddPhUSI+Zo2uB2YccaiX4Vl+QcbY1WZs4SHpenc79L+2hP
D//pf4pc9POIuPACMdcjRqwL0A0mM38JybcytdH3wR3WQvCeG8AkZdDT8ZXzkpTN
ZY3MYgHPFnYq/EfhImkfOXaPL8K00xp4xmzcTRDReAIlAcG4mtHiytfik6HhNcph
vEQ4esOHmk9ZaFv86CRrXP9gUOryOFtczNO0txle/CZkFFsI9DcV5n5I+T6fm4BU
/86NAvYlRa6JNeQKsd3w0CV4JmmmQvHWjiAP7qnBtF9Q9li7KZ7K76HmzI8/UUm+
mA7+nks7zJgaxFE+rKQ6XkolkXedtrybeIhjyOzmu4w3U7pSRp3I5CjmQh58xCVx
YI9E6VDr3497o9uSkoCyEdiZdxtQ4OUtrb3xFYqsd5p1RtIJXUNDpMJs/PQXV9U4
gQeZEdxZoVe2HWfBrBPrZ+FD8wWW9sUdVdDZrCsE7fTECVFEaJEo/neTSVMowaxg
e3FAqzf2M8TDb2yBRmGEj0qIUpAGx8hsnmnnGSBIdLDagSD9ERbm2JI/VRLeyOGE
RvZhRg8vbT3oqAjvdqnMAn57W/Bg6gQlTbhdwUfw+kSBcaBHkNC3T3nd5thR111R
JoF4R8NnO1QQNdSYQYlg4DhJT7YlZyrmEziZeBN9zkSNFQUL8/ksibvaaQ3Gdgjc
sTBKrl0g90o9CBOXGPSLrLCnUKFau2kpQ7aUpAjZJAvhBFvpa6eKLYTSSVYza1qm
+0h7weYaWeQvRfNYbJE8PocCz0ZY/J2hmZd7t7GfbuBN2Q6CkkIMUPoBgRC9gqzD
wPlsOax1+B5PQ2F3HqlcAzOe/+6bOgswpdjTMDa/k4fBu8POxJ4DwYRjMeMD+yvB
bYPlw2oOI/e2A4W0q0kjQemEsJCOVI3YKsJnhwKMt1vu2IWm/B+Evk1z2jlMfjw4
uYNisunFph2MbA5yZJ4tchoKM5UXP+1FbAkOOKCsOFIPSuz2YB39WhuFxOoRDPwa
+46W4Oucn2Bq6KOiQGk223W55xBB+GV9RnqbH7BNKpxkQJyQsOmjk3I7vQt8rIDP
Z40qIZAVl5npgc+fPcDhua2VS4ry/MwB0HmReOWJi30tNwvHfbvSoqpls0kmXEsm
zQV7kzAVaAFGfznoY6LxOGtxzhOK0dse6Z7TW1Z2D7F1qmTKkVNxJdDmqzeYA9YX
vkW8YXWQjMITPC1ReloJ4oF3VFMnj2l3tVpQNOl3/TDNMzf6ztPit2HN4/3qZzfW
2D70DiOhJ/XxAYBQgGqggH5N7VYL3Og/wdfN6FBkK8Qygg4Fo2o4neh6xQTd2jel
Hn1Hd9R4hKfI75/Fov8A4wW+uk3lGI58r3tnMCA6ofIzMDKc94AYLfP0VrLhCqW5
AKi5HlHC5yprLoTq6jexCQfgkzbprZ9Wt9Jo0ZNy3mlZ9WKEyF28ohReIDiDoAh3
xlcCe2J+ja8WYSj15S7oSLOPPJkmeVUkIyB+1f6HmqOohmHQEYIMwcH/Q+tGFdBH
x0ByTPgbqQY7gDXHZqEPeXgN7InjQ92reRRNbWrmsxjhTj3Pbl9jFQl6kGLhplhG
nTtfdxhRIM3xn8xvcFOPedCSGTVDzltiICfv/2rIJdwjDFIFvq8fRIItLl/MGRxq
RH+5CDBz5sJ7h2t0lN3PxNpv5Rl/1yVTIZvjf4EfaepxigyZqVreuGJ4gDPM6cvB
FLPAPJgekjidQ6nhzVAl68heDG5UDSnK1ZWNWZOLmdMFkZSkEPFv0w0Ohj6JZohL
yrGcgmC2DC8tBrN7yE9XwuKQ3MpNiQw+yGYiidJ25vi4+Db4aIiGA+Ciqp+WY8jW
kWW2VXQPbg33ND7xTgddx2c8TBbEgOVFVdldNMQKcrU/E/wsRKyewJ/vjP6/Zl1M
8TfdSodrbY3j/vqmoF2cPYXCTh5e6m0sOZXGjx6bGK6DF1fFep6FeleZI7ojyo6x
d6UzbxnxUMIMgpqMOeh6JPHwmjUNcD9oZ6AEfJbILWYam8IzFmcmiCqEA8IXw8Og
ZYVo1LN7YUmEp3VPzT+5VBPE33vyW/hkTJrck7GxKj29bwPL8sAU2Pau5psaWP3s
KphIaQZXMfSnHDN8nHZK3jMwakP/119ul0aQQ/B8Ffy9wH+bD2b0fJRYPaP6E1Pj
cPzyFFaI1vSNN7GC4MfJNkE3d3+34jVj1mX1alJYPLiXmP2mJnoVC4d3rzp8HvcU
HVPE+DPuo6MRDwjE3qnPumjcPAkVOihp0iQUucOwrw+cyfiiHgK3CmYKlkqQNL/5
ykQUV0nnkYlXBho+VhcfeOi44qqcBp//hsFRlAPs/YTx1Gwlrlj6BT9M6znIbf+o
EhbdLZO+qDndLdifAba7FBCZimRMHB5nbcqr25TvlanyiWGcXdAIzMfEkYaaHZqS
fTbqUFcheLQXa+fLQZP3r39RWAPUC3gjdpJ2Q2YSfZmpt9xnkVzx8TQmKI2gprCr
ubKvzpZShOb6KJdWjw1arJ/4k+Roxnoc1s9y3xtKt4NO8hxNT6b+y4OUo6ZPJt+i
8jhhpa828j5uttxprj4Lwq1apGNb++f1SLw07/BOsF7lFFAC84hO7W/27BismDKb
r17ltY1pFpicdGBSdT/l0tUje0Z2chUVv1Z0ey2lgPI78aph2rLYuoCjL2yAwFCm
vsJf4D7qYSVsrnvfdA479zjDv3Svq1ljPpENzQaq78oN351qP1s9evjuF9idoyqH
hZEDsQr9DgKBMBAYGodUCxDd173wcMXI70dmj6O+1Sex1D4yM6U3YRsk79pdfN2l
M49v4CTgDFulRtFD2hO7HD0GFE0a6IeYPD8K9DXvf/Elo1GdeYfSs8PlEVciEp3V
JMqdW3MPj/SljgJbb4bZOwX8TH4ij7DuJ+lHsSgShU76UY8FPm3jIDeopFZWX0MR
cIZbqsg+25xxBUQS5waHoRuRikwQSOCZYNK77qtyEbSneFqoCSW3q/lr/oK5hizE
TCu3SCQWH6mtMMOpme7y+8CCWlM8vjnIPBDmF5/kX8fBhODWJ8lv6VNCQApw1Xdd
+JGoyIdprj9sJGDW6hEsqFkYeJ/VkDH0/ZChEiO/5kRZmbjr9r2XLSHF7JiZc2bD
0WKTbEVDw/zkIt1tWMFXTXI3FnqBcfom4fopS1HhTypuAZmkwQRkKtyQ0fqS60Hz
M7IlyvDvFyrrc+8FDYbjTi3LdZrGrjwuKTzL4Ffoaekrq7skruF8Mc6RRie8cwPo
/JcXlrnKAuzn2LffbZwAS9Y5IerivP1tCxAoPzYK1nhzFnLhkRfUYnCh2Inb2T44
3yZ+KAVIeXK7ravFwjOV5ItXVe3mXa+ehg//+4pFQJ/aQK03rszFG1Zx69Z+f4ef
9MaC8qdEW8wumRHlKdJaIq+P6/ZUJQqCCjUybwuJiGRwhExbfvGNYpt9zhQlk97N
ZFj61ua53fkLsznpzWFrwHG1rWqBiYvb5RYsCSG6YwdumCdPzj6Yz9pYjuuI7Q9G
o6TJ6mu3qhxS7S9A2whTb3vX3DRUNPWmPEz+9C3CUtzw9BLeFpiF0S1rhrwW37VX
Bl7mYPvgXXu1MGc8hDG/Lrf1NEzfuCPGLhyIgYVbwNGEi2OOj2aqrNXRKZsV1tE/
T0P4J9/kpmd9n6A9+09G7bKol06zCIkyucln7Y4EiN26jMdBSLTW6E5JcUxNq1XY
6GMp4DJx1Ts1y7ouVsJdRNlz+wriwhQJnt5XM0uuZgOUhhskgLOar6T5a+jHXhs+
OvkQZXuspfPr4iU+IBNbWqhQ8/P9qOAe3klgu3GPopZLI7pgo3umNjqWgQlb22gP
meX8XWPBLdj9uURu3ClrP2D9/vcPhEZtK7qKHbRK/13Kyaekmt/g/UaKTiAqiKgf
ToX/Nu5NqBx9Y7CErf7EKA1LhjY3GYyCZOpNcJ08wE3Lx/MP34ZURouqtgoKELBF
ISsuqNsJvL4jzREPzjigdT97yUTryMflIoNrx9KWCTzsiknSFVbkyv4twsX9q5HX
a6JVFsPYZxnamtB0anYVeCyQq395mdkkp2uLdchu0GflTfnBh5uW/FVXXplpnUcD
7Tlxj7WXC0JZyyHPH2GfKMl9TIhAZMkbiZEEeP4SpDrUIVUEdEhgME2VRpEY/Jz0
RYbIH1Vm5mxKb9Y3r8slFmuwobAM5n7GBRWWc81bk+vBZ7t7zKZUtbACHxGGwH8U
Jd0agk8tSyH1H3pDkaAxb8zvkqTkhMp5K/PwyToIaO5FtyPZwloFES5aIp4hpfEq
Emqbwjixo59jEosjqv+sv2hHEXmIcVl4IOGmPO/LNNvFQ4FQ8Ue23fYc8fUOc1uG
hjHz397sYqXCtQ5iYzgIq2lddK/tCt9VNQb4wD2QxsiDF0G0pk0c2U8HU+jrwIvY
EO56LrAmAiwhmyY+OvlxUsGNTtn/756uwdMA/V7zF3vnaH6yt/tqqs0PRj5rI+5D
wSqtrOogTNLoNRVUxJSluoz7oO0TSJ6W8/mEWk/HtKcZ9YhHa7aYrQ06viipbeYe
rZMJYxN99WUkRR3rwEywkg8eDc6N5uSFnvpN2VHLrOllpX7havm6s1oyeluYH8g0
i5nChDrlU2HzIpqfpqTrhxdXmHr9MXWLELcZ0Bo8o3KdnJTmt6nEvDGIpWIf3dqA
yHEaRoLy63+7tKVAr0UXWwdfZ5WIPaUYMxMtiJI0CY/JlzPFlbbMcxyK/hPallNi
i8o9r12cIc8ysoLEMR7CWWymOgpHSreGllKzpBxPJMvZB8+nUZyKPI+y8kITvExP
ODHz4sGQLLtHEsUSHafJTNIhJbGXfuBtXZ+DxVsrLdeOAHNmKal8nsppYowRbEMc
Jy57HZl871GuZOeV0DxB1laFl5iRTBT2Km8x5TZwur7PutlB4q83UlRYvK0szkce
qb0GnZhMcavCIwzS1+65u7K1UlzO5dvC/kuC7pPWzjgiAcfVpfeZ8yU5B0w1yMER
TwV5cWlYTRot9euEOhNIEiEQHcI2bQLpZEaA1YWVgFgYadMGiYi2TVtk+dbI7Oez
msM346nzUFvv4cFGmnTAR/RvnUyEnzX2S8WEtqp/4SETaXbKdOYt2mgqNJU5+hOm
kT2BUi9hjlkfnBoFeaxU8Ym4J4mUtVWuP7ZVrAiuhwQ3BgNVq9ZO2ccN66bjOrLc
Mz8xOdFw1doi3A8O2L2eGLJpsMa5s3x3Lo1tjjICTLVy73FWpSAIlYOsI/8yjCH+
gZjvDdn2H3c6hfb1dIfEppqhkGb1C8UYfXyNcslGMUvPofSADBNo5lx3O/RCa1nz
u8LAohZS+tVrqs8hXyAW8UVayB+z0VUEhLfj5CsYLCzXzoQLj1Mru50xQ6gZfuvO
HbeErwvgOa9DUCJp8Pjcmu0XukA6pEhr7XTkhcQ/rVDTWo2eFvp9xaeKDDphXGNF
dF60WUhvdxqJDBjwSAcW1E9RZzvHG2OpT/efZCaC+A7h1+nJJvP6XNL5xVelv8II
9S8BXb9K/UNF6JXwcDJiYX9GHEHLOJGWV2Sg9LVAQ0vibIeYlVNOGzMlNb7poeFE
kmPvAOdM2lZL7rQJWVcSbJcBkWMx+9udLc4WydrT8puSEMp6iSDadABRIqiFnw8n
yimPJvjxbD/FoSPag6jl0lQRvA515qO0BXOKklAh3qyYGcfmc1hjfTqRWMoRrh2e
y/4oi2w97K2Jx0/5GzEZkWqnQDMjaoVUbx3XBne6h2piLw2V34FA8gfEPF7gRdXd
toZKLTOgpPRzYEmXSfKR2ZX/ZtBt0sOtRvS14qmLH5nDKF8NgFzdfEt2LVuXZmhQ
bq66icYFZZhjyDia126GdiOgYpCXuVbt3kiOxqhrFTPbQiCt3J3aiFdWafXUYLCb
Ln8ekxEyjvrV4FBjG3sX+LYx2LnPLNKyLgmxFyWS0hbviX0JzYCkgIfebPHE928d
+LYPYmyN2g6n9qZ3Z06qNmanp6MejNgFBTHRZSZenW3HVMeUg4JSswGFe8hPyyqt
8/JrFPo5n8aHzUB4zDyF1I/fSBg4De7K0Av+RFA98PTZq9f7f67HvmheVJI5ogYG
94fGtbi6XM0lSC6MCo97EKpBCBEtB0rQSfujvwf73fYcEyBYHwsVQy7xi7Da+SFy
+k3IJdLDxINJOZHMpdOTY2TCqLYsYziScoRKjlUe3SsmVUFrPw28OCuojy3EWnZM
SWcpu2tr/L+4wsAb1GXigeGUdc1fRo12fZvpJJOhDzUexPtDy4n1aADwtV1BznEL
GloEDYxIfLFBWbucB0n9uegl2rT0CWa1cQqpWSY0SoScEqV0ZjdP30qeXcKh7xtH
E2J1GP4w7LieDoHAU047HmDWySXS8szooWy44EwWG8mVWeJ8MGB0H7sjFhzOFEZh
m4n+ESKbv9ij2VwsF9KuZhP41yA3V83sfRCKtfwRHIfQQv4V5u2PtdkUfcPraQD2
hsrkFMsGK/IPY9VRcaPr7zAGi26La1NZ5ANTrHR34KVGNYxMpgrIYvZnuYwXy4jQ
RST/+ckYfjKepzQCUYjMXiyDjzS6sy55cR1eUKew5gCjji6I53NPzUkN7VwtRBJu
vz4gzvzUaHidDIAQlZRn67rl8jr7mS8ehaeQBOeq8gZXQElExt4bSj1U4vdpswZ7
k/SMnlMvIYsSdRO7gJMoiHIC1BKHv9AFCnJluXE/vpSZSKY9LHklbMQR6NtFiLfi
B3iSyZcV7Q0WmQT6H/Ga8cPiqRROOmCORr1WFmokLCUDl/h3xD5k2qqMQLd2nvrJ
ZE/5ZTL28x/dBJT4EFetOFDjOMvfzS8n11VolD+zv3uSwGvxWa/zRKk9HYxi1fJi
7jh1KQ/c6Ipu+IjlWQpPZjHk1BoVgu14bt1uTAJzGu0LwG95acI2dFvX3p97URgC
nIeW7vMEMpGVYjA7Eoke1u74JbhEnigCZJwZnPFj3nIa23FbCtA28tgH9E2L3qIR
40znTRHQ+oFeBTHspO1pw9NJ29EMlrbwPl4u/FFch3eO73odBSAiyV8kFhXFFOJW
Ll8wogsOQT9JwgGVvp5ACP00expD39/BdKCn9EqB3oDSIJOuZB+TQ3TKYN1gws5K
c/sYktb8ZKl02lP0nXPkvVmSVo/eyCLy/NV92bg9jbCvr/pVA7iHS6mR2LdS4M+7
wZZqAI38Xw5jB2Pbi8ezbF9LvQBo7zSSbxDBGmZmHDVf6DXI1r+Ay3RCQ6dZQJVZ
OqpacE9CnHc+X7oCS7LJXPT5F+k5C0VzqzLRCoJFkhxAtihAjTaeUbqtFIcN3GjT
Ow5u6ALB2mwvGQLmr4F+fBMxKqmE7jd/TKgXV/OxHashmtRDZtFU33UefMb5ObJm
qG6TJiUnlsmtlymalAdfOrbh+MVvEOO/AlkyFbFxQlXTLJ1ggU2Su/Mfh0yW/XeX
DfppuoeWstaJBZxBFRyllOg8B2Uq7akBqZSTxn90QfOOE0BJK04gTbNqLvodnNDa
qlIIYHeMyK3S56lYq8d+kzc0NiBy/eWbo9qhpGn7+0npKIMDlYtPkGe75YNhaQBC
1ekZ52fIjVorZu9y+A/ucCHCFl0aFRkvGsjlUKlOBMBGiL5eozEinfWIVALdiDOn
iX6k7Y05ORoCAUlcc2veCpuXKcfFfdi9v8GZNHcGpcHRogzUW7w1LEEHra6//vtq
hwDEqklzkcZP8FUSE597Ky51O8Li0eTC/E+/OrXH9txJIG7LOD9MzXY06aT124J2
PJWINpNo22kNVdx8x9bgaC1F7DpKqN55EkD9MwozkltbPxo/hjniv71qv0K9eQEp
H30rR0j1InmjA9xWH+07h79awhyWKawnGJJisW5T+6M8x024CdMmB3YWS2SQb5P5
zjgyYdGFeHDyZwWlJTBdzoDtjl9NRHLtm6yY04ALJHWlY+LZgr7vYXr5hrTwLqrX
PGgyYSkttRhzpYdz8vwmHmizJiXqwK/xL+Bld6vgtiPHcVTwGi6IHsIxQU17pyKg
3c3GTwkeodHEMIbUJhSD3gdeMHcvsyRLbxlQGVEy8cG75nb1V+pijJtvW/NoTANY
eCcq7bAchT4oz37GEhz39iCViHN6NqXaUAFJ33hENi30rFnGqIXxv0uCj/FLvhEv
SQCa4VJYAtQKY1LM9qgYk/U4AVKmZXDpk3mg2UMGsdXAR8rtNC2tmVWAZgGEol2C
jOmxz2uDZaOd8YCNN4mcF2/9AQMzibgsbxPDvqJxjLR9oywp7GQLp0lfjhpdahmj
OwTgyBKDLklVfqMXm6QQ5nviGSkNouztLC2V2KyfRQ/Tv4XXPFoNfkifyh2ewQix
LaLkDOmqeUWup31Qm1/O4N8Jhm6mTac5Q4LobGZ5QcCdOtU0FIVh0tIchCXAAcfJ
tpGxv01S2+N4YrPfBRcEPLI5hHu0PqMBIog9h47R8SIgOhkp6rsi2MLLqVLcUJsc
fxE6sidr/PPsRbQcemXuP1TtOUv7fu6hhE4BsgUOCxEEqNyTl/pC3CrsGR51Xlhd
EUtFooRruBTKfY9Kd9J7EaLzHd5mSkfU/6UGQEIQLMQ4ztygXfBW2IgboRzNQZdN
chv0tpXW8yEZXtjpv5rSYCJj0BoPlLCe6QQwkWaePZq4FwWwFLNZ+7cFkPnhRBEh
A+5skJlBrN74iztZhPoh43ODFaxErXSAUayTexZBV5VLAIffHty4k1IrfeF9S9G5
/UM6i22HqUbccM8X9pKiZyS5kpqT0XKg7Y7Z1LOt6HbGD/YL3gzHmuZySzVVtW69
yEGR4OMdcP1iewLz3tUhv3BJJH3DTcoi6c2FF6b6QjB/v1nYHygvfDSOrAGtkym4
zx7ODEruhO52MpPQvCh89uvgWYGbh+/3/bocUmsLAZwEqIsKq+kqsY84nvqWkbpP
u8xBgVJg7pLEnfXcLqfUsahlWNGpYLEG2HrMeFuWBdhQUdg2/jwwCl3xbUw4Ymxo
FexS9Mb9iVAF9pkrL0nOVv4aexSamEVWrW1HaWWPmfr9CIy2RdodFaJSJ/OMU9D2
SC53lWWLv3wFkQhRHQo4OgkajHW5fttg8OxNdgcVkAT9v9B9NN6Q/tv+IwtGU3Ef
Z4ebAaC186Rp67R6JbevrDJlU/RfnfWlufRWWCH4jogxEeXMYqmLcP0NNX+5ypsS
NHY4tmxn3k79M9drVvaK2WYKPc7vRCZCRU1QIiTC7/uu41XUcFf3Hgc0EkWJrAIr
43HTwRubPwJWIhiR6uXYmNAy9+T1pnrIgiqm8a5RVwI/Hy8aZ6veiOLcPH996Bb3
w36UTrMp2XpTitB0okNOGcCmtgq3eFRIgNu99JKcbXOp0LpspqdvnKn9Yp1eCql8
WXVGBQk634TTLTaJfQosognxPtVko4PcEldacDkXAB4ov28opniVSrG6bkBMBxg6
gteMpEZMNikcc0h5M2luJB1RgQ+yExywNNJNgoz5IP5dCtrhd8C0FGyduzyDyeMr
MfnDppS7hV4tCJJXN9Rv7zAFiHH5w27SBmy8+htSOX5dxaZfGuswNrxEvavKrTld
XQ8Gg/XzMT3GdtE32YyT3S46vHpI3Ga/d5hWfQLebnql7tbStrn0I1ups49/3UQV
HBV5SlOnpgmax3Q2CjD+Fi8CxpppQ01aReuJW4psY88ptc7vSLZxywO4VPb/XtsV
YASod74tU0h1GI0gsTy5M3dc9iWgRH3DlpJihVU++1wkZuR3FG95o27Zb2xnWD/7
/BMJGd0cwrEaAnawTH/j8V4i/P3ji0UXJQFl20aeoOpswLY/1PKHQXAw47CtLhWE
DdBEgwxWZOV3ySvV852axT1EYqoI5klkvZu51iAYzcYuK4uL+lhi7hTptojYdtIg
PFhn/8PhjKibD1A0ll3qLLtmEH6Ulb7euz+NxUrDtp+EPosg3Tgpml9XNEBaMdSg
Uv3krIb1EUQ6aCu6XUbNKeBmmK2/khhsDz4PRnH/fmCtLtT3pxJdHjFn/Kp001Ba
6WO6vnXxm6bwnv3IvaDy2go3YXlcv0IOPoyX3bBDsBb0zMH5Aj+0qjmlBMDaigAt
7xj+ZTy3wBXITPot29D0Htz+iUjQ9FLXmufrvA/6vweWLE/8JShSlO5R9T1iBZCo
lQLB19dqVa8dgvV532lWp6zhSA8GVMF0sHRQhHGnC+h+dwgqiss366WmmaErR83G
nhP58uRur8h1iQA8wUBseC+Lr7tK0MA+zBa7i+Rk7x3S3TBHmMfoWAUXwdEa8E5u
fggGLRqTiTilPBMmoLgvwI0QvfKfJOQgYWkx+jvjMYw4gO809hMzDDN99W4M4jm+
3QrlEFkrvDnVAb40+dKCA5YiPkF5CZJQ7+gC6bJVmgMRkrRR5WLskFr6arLKAOCc
YPQJwVBbwja4rdUWU7BrAePeux9XOrP2xytmqpXBK8EyYkMh3BjL/c13f1r9XeEq
Qr/ESUpKnhjqtt4HtDaYVZu3DUrVQ64JQ+4aj+iztme9J5qTZKXA3J4k6cPeX7kR
2ps1Qy7//IiZvvMwFt2/8IXcODU9ej9Cb9ds4wP4mAPsBhpsw/zoZ9kYZR+5zLeT
kMYtJFCT8ODfj6k8OiHioAt4wY7QtuH1b/nizG5UfAVxjnLKGWWLYQymr8aFKvn9
IvppRQNwQST6evxIZMNVvo6cHydhfSBxuf4sOtK5BRxSG0CZ9zFjmvZ8Ed6R2FQe
fTykDykQwTfNJT624jUnp7Ltd08+n7MXgPVgBkh5Z4tFXHbAckvECqOwgYZ5DQxP
Pm8lclXnD2YRQ2kfNhvrtFNgZuVjFJJ+iG9o7SdSIuCNka5CyLy1HJfVkjAyPIum
3aDHu0/A8B6FohAz3gQ9tdDUJYxKLQ6ngfEorxkoOMQ/agwwAO+Hqb1qnoqqLuRe
6kcrSAkJjPEXShCGkjJ7HpMixZMJq4CvNUR8QipZEW+8W3wAIMBfp9js7KiW4iWP
g6Zd53Is2ECZhrbOsQudojmh3QkBbGlJooxBvZ+cOCHX7D4Nf8uBkw3t1gIMiMYg
Fb22Mfugel30K+kORSxgOyp2F6HyLYOQy8mgk7pg9uFu+KzgTKmgL1MInRPkRGBX
1nF8sNYO4r0aEIiysDq6Efmi21sNOQm4Zjf4xustHGAJbfvGX5ePI2XH4QCpDf9k
e8TuR1jiZZEP7iq2WErMmRVXF7KtT6prQK3zovTOEvJH9wctuwOuh1qnEukE2GAJ
8r3blquzWbw7MYBarkn6oS8Rci9kWW8YwEReEm68Fz2CVkGbwqy9Oq+D2adiVF8Y
g+2Bc7yitT1i4QKOU2i404++xvtwpScE6rbn0lH947fDz1dNC22mJ/pHEIynp70j
aYEuEEHIdtKN/riNZStwABPjrodEdMSywTgXEa/y+4rNo9hs0Uqe9/92beB2BhDp
miIl3VHvcPWJ8oUgrC96HdeOUJOA2ZTGVbJ5EAZ8Ukk+uopvUblhMmSDjxJG2trL
K+hqogxCJaks+WDMi7g/9Dh2GVyhFEFZFTTqNXAj/brDgnkAKqM3vrXqZGpMNiGx
IhDBS1U1kKI/1ixxH2POFGF7leo4u3vtDRzwaTVkIHYnP6h7pWxlzpHlQNrk8E8x
nsvsP2GOlNpOL9E7u0fVfqwrtvFI5ORVB6x3gxek0WHYWdq/h4L8EOzGIZlKPZeD
lNCrgbCGlt8XQe1S3HrsqikiS7dmt96VYdN6WPA/OgNf7a3PLxuVt2Tpy3O6vH6K
lnONLNlozCTHkZnupnblTH4df0IRq9NQU4lqhKu7FYOqrP0QvSTh+MeY80u2koDT
sI8iQLBeuEvucCG8vOubx94kLZ/Z8x2H9/WltevQmvQs+c9t4RreMdSgDkmFscen
rCtymaA8ToftsAqVW47dKMWJy6v2tCISZYYlxeXr63JpeSDGJp5FZoU5aW6mY/s5
cpJkkDsQjMPkJQYQUsDAa3My0ddKyIUX3KXr6s2hKik8B6SBPxjeu8PCKPTOhP60
ityn1mXBQK7v1NspfXhCZMzqxkQ9gT3fUzUOrBxzfvVxZlD5Jb1+AjmfZwUjt6LZ
Y/eFOSSlGH+ON2pdnDMF4L+LqFM6hmIVXZaY14TCRohnzv/K1ZAxrf2qRaNZBNB6
GAmNW0+iOPbNSjOk+NJQQgf+Fcs1DfJevHMTgblOg4ngYw4YiXX7h01d+CZQk2hX
VR4lRDf5JVJkCJ/CBPiWmgVFncXTpAHWlZcLe0+eqCf/1/xpKoCYtnqKB7ci/aVH
mcDLfpJSYfwTLs3J+IozrfcVhbtiRyIWiF4cwbkD3DK//0OWqUjTcIWk06VdOiQq
/M5ZlOV8EwIoGoruNgBwES+BhM+LWNHFLxA3HqSNBotO5SJ3mwp+ZOEgcmcIdDP7
1YLRL+0fXDd4Nj9Frppv5WgAhJt0xR6pr1H3VYkYwfiwz1lFiVi8vsMJM/+wKSxr
1EKigi+4047sVQA99MnkowMMzKIgH8BM196uWcUPgw/gZ31W/+E6+x4xwaN/I4mh
y6213OdiupuD8LQv280yYQgAwMSo1Gmj6tWDLxVFX4nPRsHyBl8RH5UOAigwCAhw
j4FmTiCkbwBAcFAcqLFl2TbogFVIewn6JmRnWIyOy2De2+wkl66YHzYmnXG+LTML
uMV5xlpW+Zy2rNmxkFCMZNK7286uH7i7zgmfLl58wr7YjiqJR6BEQiQwwTVy5Dvq
9AjZF58lxWnfj6GNJ2IsqfxChGijLxUGQ37DxvUhgEbge0BeC74s3WcbhixybOqJ
s+NY8ix4oJHAsnWd5pSzUMrNrWXiDN4eLp6kTVlRZ2sX1sNOB0KI+Rfm1LoCHuWE
SsKA+YZZZpAn+hgdpJz9HKmxME4L8mJLRMleQi3eMFtaZmkwCKuy9PfSMu87Ts8l
UjUwenlOcB7eJrfCZI22cK1t3iEp6hYk50ovYJDgBvpl+QuUuyl74A0lo60yp8uG
4toCzHc7zaQ/J+zJDB9cnC24EZZxDcvaHnJU+iOrCER/xfzjgLcovGcdMfLm9Ypm
HhJ4/tJAmUvfs5g7lZqz1ylQXJmruNnbHWnuSiJjYcAvHdNZuuXtflVkNtDgrIAs
eNEc6NRXLR0hQDPX+9jMBX/3XBxBtcUWl6eHTX/j3xuvhfcFmcWZEkh+WlqIUmgT
qvWS68+hW27H4FbgUWoJYx0VvLKw6z4zDR5bbOGsAR21TijvMNLxAILfYga1cCkm
KdYlYnWzy26Q7u1b7yjmeTVsayuEOIFqechZzSd2rpNwJS25n6r3r06LjfBWNvq0
sq4Dx8ut97MlUmq5RUuCoYhx5SE8qNXgcLUDGxxQB+9o1eXlj+xe+sI6Y2gWh69K
nlNq/T11rI26snZ9fnN59GaYzE9xdmh4e/T8WQ2qSFRzWgE06TOIwWVnQiqe/xa2
On1D3hSat7O2vrAxjhpB52YmCRd/QBwLgrejgp3tH5nuX6XniN8rQ5jjdN7ZuUHa
HCUVGy2qEQBLem8rFRzoeACBSzSeifoKmXlFVHMyRo0i2gqrKZXZFxpkRatf/6Sc
cEaQVDY5jRPI4FHUQ2LTobBMCpLVeofoBRfKQ60/6n+ki7yxuRKSr2/rLd76eQxP
R1NOerki8zeSfzOqrLA+Jktb2aVc2xhlk2/n+j6HoN+FSX801Yr02J2iQ/pJjR14
RZbVPClQXrSuHTV+oxkwkxf9+jdyPljMkshc6LMXDdAylcreezpz+9ZrhNiLzC0o
Wt+JA6Xl/VayOBUZ40SH92gqSfBpu4lDpWrATkrYrzS9JtWQFanhAJB8Ozx+IUlQ
9nooaRwrYtz55AZGq0YG8zxC7YpHP4NvNVkL8QpT1ImLxVAFAei3mJ3mrEbW+NQJ
f+t5ukLfHfV9OrRFC091RpUMvyNaion0N9A4+HK/BeKrewDAxK9NCvOd2Vb8krpR
TMpFxCaGaD6PTc7iCjWX2kSvO988nHdPzmeIokpGZU9t0NdLCn4/WEYwWlKyY3F6
GpIotWIqPHmCwUkofPNF2K3Pkqu3wKw/OZ8Sb2Cc8jQqsQAw3QT6i4X5sBwgH5sg
tUws9p2ALfdwxV4JVaKQ7gUCWs64DWkGVTdsVbsmi9HH44I7lHEOMhNd6ZZFbTR2
aayGdn1uiCJUD7Gy+zQyTrXuedHBJKvl4P21rHySHmnZUMLk3z549auuZBu4WZ+z
8AVviSq0xTspzfG4REwTT3w8mgb/XVhCJc80rDEbnb4frMvMOLBI/oyDRg9VLkXm
XohTwjUxKshkpol0X4UY7elcQvsmnUAsxnt5bHa++KOz1UVYUzrvgh/Nkipempxg
ywvddxC3uyKC58ESjJ7eaDOlqW0RiQQfcoYHzAgX9I2zTOgA2gp11z/bN7zXu1W+
UPu6YT5TQRQ7jl1VVlTfxPzy2y6HoJcyNqM1I4m15+uR6sP5IgKwNPgivotKzYQ/
TYJ8ImtiMhpdy04MYS+fuaQ1kn3osDeA+IUzWxVmGJo0DxoMSYCXRMKBajqBz9+q
FgGXG9yBFyM+jVlWOaTQXnxjWmfnXzXJDG9RJam1Suy9hBY2MiCOzBkpgDhgRb84
p1IrK6yYD/X8KSWRvoWKthd5hAKLpkMgaTW8B2rBhHFMeRtkFo+Nw2IdeD2py/yK
rteN/sXYuGV8iPY/Dnj/3gEY86WwNJy50KLVYcnIPhqUtmrBFe+jeSYfUAI6zilP
Rsc0MkfJ8M+qfGBTmCV/96gLgPIBM/V7Mf8WyVNCsrVwRFcrzsEtTnRvYQMXXzXf
lq/U/RGYrg1K47Cd4rlKZNhuSZjzYwDd6k8Zw/v9C9OycERdomZ99dbm2sM0bUbk
38sQx1IqFZUsJlUnIMCvadlziJ62/FuDz95wHu48R6rKGfiXHIeNJwUI7PX9JRAR
7F2x3HViQO3xQq6QazdiK7uU6LQfW1JzDQYs8MPYmMRRO7uVWrmVtimq5UESZFtA
1IDGzkqI1H5BBA4bJ94dIkKCGGwikLJnfzHry7wHYZEO0oIBczu13X2FgDEfXRc0
wgenP1Opwyhp1zwKS5R+xFSRIFSCGhhtEF6weJz1EOlfy4TOYtE+JZALN6SEQgQO
DwDS7e16g3COFXJR/dT6wYHX1ssLuEnLF9hdf+RWcYcEm2wqtyniMiSzHMHpAdRf
2eqL8Rbcw9bOA5dvdOgupsgsagZKlblg7OpYO/MMVauBrT6grfxD3EcZLPkH15ak
SrVXmmatZQVaC73u6o3GUvdmD595+HihtvEyhdEgZDZMaV290OUtljJWFU0VTyii
NadcyepOODoCqzdzQcns65aEhPkw8na3QDeifIC+dgR8o9wPlatZ8cAUQPNPagsH
nfuEtMNHgoQ79hwc5/0ATKIFj6kSUtIg6V/9NgJksUeT65Cp5ULaaZpb5jffrFZ5
J3tDznWCJbYvmYmYwPOI4Z1op1ELsweYKfwIzr6BJjoZenfk71/FgAcWlaSdoBsL
UBiI/WV5OsW+DpiKcOedM5pcYOKA/WUDsoBLKmvGBXm/jPzDEt3kM94vvNnDLcLm
cx1nt50fPBJt8DPgDvaB6OA93+JqKxaEmhEpsJFXsB74HTwtpTNUKcBQhMQMhs96
7y416VL/yxyKQIgAyEwqlm/7ShVAeg4D6mqfzNxf6HT9/b0fjqcJg/5PYNyVsoMK
Ni7GIPU/42YOvYzfJwfzf0Xqb1MUhWiZKAirhBViw958GQpExsrsur+my5LZI37H
xcT+bGZeQ/fTlmdSvBTHHJgq1lQnFKxqYThu3nSoVOz+9PQxV1B+esabOetasulP
wJZZXnOvEawfwswo3fle2xC8XvXNS74sEq4KUD8MjubLRcKrpX/tUBRMiD2FpdIj
fT6aIbhUzxBQa221zAf9U+EDRSE6/6/GDM/V2+ypg+89yofsfrHmqQC/cxz4d1Pn
Znt2tvyGA8nREaCGlexGaQ2WsB6L+AK1F5nQint+liMs9zUDeN5VbeGHXqsnfbWh
SXs2fpjEuQXBlFgf3ZTTUUkwm5ZoRDO2iHGOgWY2NhaPb/c5oGsr32FGqVCiQT6v
mKMSMBQ1V257JhYr7ZMocG8Vuia8ANXT9iUm/zGjYF3knXdxfCRUh5zVGlNbJxic
5BwJvhqtg6q9lbsWcuiK7rUpYdN/XiUzsQ7fdQswsyeJWJF3QjTASwnaHKNcxU1q
MlzpaL7o5om7W+4em7AdxcgElGR4suD2pkxibaYef75x0FeH0/wBP6wKBZQ9iwz+
2AtGzCMMgVuDju0jsWQrDrZpTx6xJnwSl17OTXg6sPo7EwdnTQ18jooL3MelZ8Oy
J+7AV5ToCx2d0ZZft3Rq4+Z87aroUhuFhCT7RjIexg0X9Op4vrmaTANTcjoLEbY4
QhKsUorgZbQXEe10etMnDENxwckv91nn9DsEq4kSBbPFBAKe3mvFlZK6aAoLuCjR
7AdJL4QumEy5c9qgKZJEQ6RWiD4w8IhTWvNlmR2/0WMI9jFfStXe1XR6gVhdbopL
u+95KVa4qKk+WNzk17XDzQ3P5uUx5wWts1iTf4o5YD80oTIHbh6C4aekYse1P/Ew
92yxIbt1Hc2pV6xfYNcJDOmkiMZkSdSC5Zcf/NBexQX67x4okNsv3k0ZR+eIazY0
eCCt+r5yrpTmGkZsEZbGmuQ0uq/Ujg/CSjiSvM3UByhf8fVuqR9iP2kfFsDBOAYQ
DaEzjhnjvv+udgNhLC4NZ8aFdS4LkUoC0ELCWFBZXK78cvGFgZ5iX1f0drincLDe
/pQWPjRxa63RXMUVjvq9K61zLNEfDygVbjLQzPlu5ZdBIetvkTHpyOEOkIVRhtLm
hE1OHsdmBUfHxF/q13J1CZ9KMKofBoIgywWlzHBgKXKs4V+GfYwL4BapLKc3lYst
4soY0/PhQrZHpAtcztlQuo0p/Ks9XpGTmZfXDjkrMcUzqIwcVv2KfBys0lpGGZHf
deqdtY3L8UP5yLRHCzUKVwzFSSpONdQXochpw6Ksw4K9YYrQWJ/h0m6g7v0p50VQ
WrS2KlVtsov8gQP7i6BFrxzXeVvjbLN9GY1Wk4Tg+Tb1JFWfn0fe9etwR+04fSBQ
7s2I/3qhXmvueV39yc1K3huqoSTge/WiiPTdjEOUSTY29BvLSdhmIq3f/3CKQHdW
INSx87+47q9tQSNDWdNCEoY6r4NGKp2zmUzcFzUOHt+LlEoov27XWhGPCYarJL5S
mQmRLacD8I/5Pz2/ShdFxxwbkWs2OyJZ5818e9BM6HHJxLlvYhcsOuiMHxFgnjuE
5IRcVNcSEhML4LCJ9rCcL5D5nMeytV8A8/EggKZg0z2ceULnMlhP1iRa30cROnK8
AVSpOTlH0uT3XnM29ccIP8ih0sUUHbBc77hITWRUzsZf5ViXulziaRyA/RsxJAMz
Ht1js9rSKOq6HJrIC0VxEMnQ3DImRICQgDEgZjaA//7fJzlpWQSSYDZABllsT2OA
FcFKB16SBYfjXmZAdki/nLhDrUf0UUB8bCQPiiJ8Rq7KIxfRp568siEYipmYkKIf
xSa0eJT32euEWoyt9Nge1MEJrQJ5QJlFRza40WQa1QTugiZTW2IsdXIk+uTHCT7B
eESHLgWllQZaCGLRstbu0rRiouQnCuUN815NSTAkh+MWe/nUc0NTHov8IA6kjIyA
QU4n8MRlQR1HQKrAfwSOHHtSi2Y1Gl/rAaOa5rckT7puZhFN7k38jyNvnWLjLwfg
yuUKrquIw5AH5QEo8YRE+BxzXsPcm4z9IIY+345tXtg4FGPWV2qHkAk2F0WZdXLB
4WQALpl+ZuHj3s10x+sd8+1BLVLkoQvL2TMC6xa9cZxnnoKbN1x+GtvlXFpQrHBo
rHWY7N9aXxFc6Y4/oo6iEyaKybpzOsEoKREmzV1eZerrBs7O5pO3QSXinhntQjhS
lP1pIyn1uBvw1zr2hyNIeTw8bhiXioZ0qd30YrMMGbifVEzPaDctOwmBjHGOEfh1
eGOjHnRKgjfbZwqQ2LHM2zEqrFJSn0rNJXeiE8u8iAXx1KbxjA2U/kAULvGULwDa
m3ghyG59QGal5oJAlBAnAxoBijHLeLkOetleiXBeLyCIgAa7dVKRreeqg0ptroFA
aSjKfZh0Fh/hkiILRknzH3Oju7Vsbk5opBjDaMF/ujtaWOytHpouXgwAj0zoUa7M
gfV+a6Z5C84rFzki4MeKVnlWT1zD7L1FCRar2wKdn5almcS6hsCTe0+QNS65ov/N
zvprelV9NeiumZ9M8zoIYHljUfzUy6ac3oDdlqnPpnLUgpgWEbCTDc4UBLMNnmhj
PxXZ/Lkl/YhUOtmYLJIqXyyTT+gw280tWZ5BuCbl0w915y5ClbRZj2Q98nrooR0z
X45pdrFSfinjIzP+eRwprXyc/s8WDW3qdCph97UjZ8nXhgJfk05dGMJ4tgIDkxxk
4w4dtTraT7HA3ScB4e3UiBXed1et0eYIn+xEDwL0xm1VEgXyWnmtg9SizEVloI+4
GHzVYQM+UujbQucAvAuw6oCHqwYc7a7wl3u9bTpmXKSfd0moEVsqW+UnP2vq4H/k
qTbuIxJGOXyK4BU9r7mCbF3kyazqxUTaR/7iJMPECUs4u46wG9i8vkuetDfOper4
qCXf0Ahz9CqlDmqmDtTfBT8J+LM5oCgzgwoRvBwbuWLEqmCpNd6QLdgrv5z/spHG
gZNl8S+nNwgF2HqlPwWKH2rzDlqeyJB8wtXN9/eAHYFesA7zzqLZ2Q5sZk3PTM4n
c3SF4Z13ut7qjkQwGgDzvqWJ/eETQcnWqjwamIpkGGIdnaDqRzomqAFVyH5Xd1Tb
EvUXS1UUE4YHYq0IleA5R91OUJkWC4xpiTkI3ZObn7kdFNphu1Zs289UenWkoFC2
+u5SsBjjMZuqEZJnLzKYguxO5dBN4gttSckNGgiYoSo7z2B5e0ug6e7Q9uqOvsjW
vv2kZ8Wa10wbp5mRh7p2zMCNeT2bHAsvqseGH734sN2XnxCqN+YNt9PvPmwY0VvX
ZWZ8gA/7c9VYDmZj+dMjLoeapfGNYoZDzI4fY5BjuWcdEbab3pi2mpywbmc3kss3
YtJ6c+xwaRlXQsRiJyEl15FSnc6G4qhuwj+Y2wWzmoRu9Lz2KTGHi023oBTEqPy/
RNLTW1sDx5OItEGOnIjRyD9aYj+MIyPz8gwgqM6VNltxJTrtpobiT/6HdvEbho0N
15EoT65ckPxO+2vL6dZWTjDsHWYa+e77t+zh5jzoXG9+a8PAozI4FB5kJM4kAZ6S
qawW3KAqYEKpRqpnfxFDxzMMR5IBwuK/Pg1EVofjYz0CJ2XEcBPUrsSjNpxjRjw+
N5Rf/2+gwoTRL7Kp4wHXydABHLTsLUN8UJ/43ILIU16zlqCsg5773UGNkNyXIuXi
8j+jYhUNUJgYPzaG7Tu1dT6pbEUivNqtE58Rxu4Fse8td3NCENNGJ9C76yeDqpzM
eXS1ngrnzrNkIi1wgb11qHkBlO++zixOqznIlYggyLOjQuh7PmlaZN8QNRN3sB0j
NK+bhV4pv2LyYgbEznIfn2rphKnCjByHxHv4NETMglNUCVdoAMQxbusXO9NWS3wD
6UWKzhefYnLBMqLAdDwDPhkjTIUOA9Jnb0jbGBzmwGRYdBnyc6w9eE9KmJjDZ8f9
6lr5t+X2y2aTc3x06hoKFsvQ4jL+OEN9hWbP9Od7IVL+Ee458BqX3aZrkhTyKp6m
5gww9w/MKLjmWrH+Qyqp0t6kcW1D+sG1wTf62NcvGXj3B1UaEzX0YjGvBRY2Cj5F
dXYPCZ8Tf6I+p0/M6yVIgkCNUUmKxliZCTTLik61PsnAgAwUeXhFoPFrEzHes5hI
Qay+dIDbfRXUF8YbBBGEKE8xCJn7qjknzsAdnFpeJQjHILOEl5E6QSweGB82Jvd8
rgo+E24ORcQWdVrgt/2ziJ30aUEdhX3shjdn6LYppAsIUp9pgZL4ZJZh0ik0cvEu
Q8fYa8PB0I+gtvQmghRIIFNdUKQTc8pa6w0ojVI8ACqZFjXajnK1h/KW8Exwy1kF
aOF3F3p/8m4dKG1ocY3ql5FvlVfsGAihfZogdA/ZUWhj2X2rBFg9DPDFeY7axqsJ
WWdgQXHpKdg3RjyZx9cmzob9XtjwgqdExlnxseSjP6hrCZNnmtZinfxh+0NqGhBz
cKFkMIRfFT0aheYKb2sTulumaLmES2bRMeehb5G2NAjkjZmhWWiEVx8xaRW7YrB0
i09RR7kVVPDy6RT37ycCyAMbeNp5NfGvvdGzBiRtfqMmOlXpTkOFZG+guEhLiVpZ
+VJ2UMIAcZAVx8klRTfMR0g/flbUE5cH8wGs1vOslH9t+rrlq0Su06hg+AZ22WRG
kIUZNgX/uwMUSwjN1lX+pWxq3AcOzr9+G12TTMvkHwY52uXub+R1H5JE2du/rW6c
cj3lSQwzsvu6RAVB8vioSoY7MZDNcCLgbPicH3PGeWaUomWVUQpBV8gg9LSSMCds
8xOCV/iVrQJ+VnffOdUsiUKDR04CZsk1+2NT5uI964cYee2WtnLtaIlVCKby2S3L
AOPrCzaVAnpNPTNCINckl+pr85FNrbg4gDknLF5QUF+Erh/Ed3NvoC4I6iNK4IsE
XtGSzYBbPxKqI2/iWTwu26IBTYFK8dctOsCKnpe4sc26+795etGaYiL/bTW5zsgT
UM0xpOZI+DRDLOzS32HSYesB+z31oQtRztBDccBfqq1PF6/JzwfnkyuFiQzuBhMH
AVG16STSHC1obkbR5OjL7nQ4VQ9j4sMS8lE4rcvCyIz3NgzKZY+QF9e4b4fdtAjd
Up3/wklOgfAoy+rQh2p6i7ATJUza5aT1cqhrJQH4K9Fa+nWcG5/ycSWQs5X6hQMP
4FRozPAqwzCQsjWf0JnqwqUtQEfThke56S052hM0f5Nc6UcLcgUppazw04zY4sm5
WXKOEe397lbyhW1HDeNut/FJn1NIWURibAiNftW06zuuclF++kqls5mzeC3UChnp
rsQ2vS0ayFTqP1+SV+paG4FWmyEnrnrShkqMez9WsOGf7IpD375mYyVyjLs281oJ
UB1uxJgRfoXyMQGFuOoTYh6ebkE3nOAFSWLkucsqG75vscsjCvXEAHNEDFlBITtN
NSHZrSm3Q0g+0c0E9farV6G7hF+f+7St62YLq4h5skNWuUBVQIiOOS9i/k531zpD
MwcCbSoDJP25CFsDiwGd+3SpjSTrl4I7lwiBsyi4y+gwCRmdWwbkAWd1+il9+5m9
eHX5MtP4HQg1pdtDIPCSBl65N0AwsHcvPD1eg/hb2MronJZ7uoNxi/7pLu1293bd
x8ta5Oa7zErfTylue+miOJLcmI5MWEy2aVLlNeAr3oCasFXvRXgeQ43Ng6XFHffx
s77ji4ls5fFFWIHBORnEe/sQIQsG/UuEDxrf8wpibFJHEgWmG1eY7dH7ONjcgFMW
IQlvuke2iOzJ34UmeyV0Xn9fZge/yUz/V1TgzZmpNprLnqtMMn6ynCxAJouSFh7n
W3TyUMozg/2zafmiAILaejncoxRiINQglkVjbv8xfFpQSwKqSTjha+Eje0EzZb79
f2Co5qhb04DzbchFA5kVrtwimqOPG1HtE5hhUK7uxeyKXHpxHcyNi39MP8o9m2C/
CigKvuwkq6MQac5f6TzYjsGWm1j1eLI+tzafDfKA47jjHB+z8v2w3Fv/5+dlmKE8
dmv1d+eOlu8+3gLg/YuSGWYHM8VxLzHFOA+3UQIk0YdznCDiNrIISLXWC2qKh2Y7
fQ2KTUBnSBVVrYdOWM/l1GDh/JH/PU+scDJjMZh8TxyM8zsGFiAjbBr/etdPMt+u
auGyzoAjSrzH0v9Fi5Vatf8AfHu++h4zAfaVQBVPyBFAkOMf4PhVVs6JbgnxhEJZ
0UlQvG58kCstKFNDcinG5xYZzciNvWq/9kwK2DQvnm8Bs45W1qOh4zCpkxO8OJbr
JP2cpOWmnXGmUwj75LRLiR4Qg/B1Y6wUJopKo+FvvKNIL5+7b57QmwfSQHRy3QBX
EG/bd9RgwbLXBCpFAFSJllRi9RUoNM1DdHJQ/XMplV39Mun2SxaLLyl1qpYlffuV
DMiHzqeadRch1PQoTeoL81gGsNaDDLmrRWEJBJN7qA9vrZ1XlRvv/XV2rNDjbqhj
BvI/oCV/rPvaKVHocoQ5OO+QrLyWi78cgbInSUKQYZvVhO/Ee1M+DNV/xlHK7B7K
r3kp8DcK5Y88PN9CmqCSryh3Kr1z0PWoaPj6NiDaclbaD637oP7G212h+8xsUqBY
0zJ2neYj/jWVHYD+ceTZ7GPtx8DfIeO1C5us3ViZ/ifEcR57aP9DT0l2aWGFvWOc
ZCTluUoNyT/f6QrZ4dH8U1Oq8hYNcv99+w+voUBFV7BLvgpIinLH5axBonW7u296
2RG3/i4l8gwHdmU4XtkpATty/UHVkOhqaBCjcUF31zPurPQPOU5v+K5T/kUvb9Gm
B7qhMsthNigjDTMSsG+uuCTUJCeyqpYHQ3XRAH2jfQIK1nz7HZKqUq4aIyLJkdKr
99NTQeznoxQwS6oO2uuIazO1F4pKbI2IhK3dqB9s6pQ9CdabWPAOE3cSIaeA6GTr
Gi4PxG467+zw6W+/UwlSPIQusmtqDsQCXSlclmo1++5ZCO49BS8WSAWSdtIvub24
ZY2ia51MFw8s1jjAx2ve89r4dRxYiSUEVgRQXMEusIHV1zfoM2IgJkIBxquB7GMl
YVoAxEVU5taVh1nge5gZqKr7Dx7W9F6Lfc7ytLCUuqvpdmib14kAJ9Jm84cvS3Kn
/MmzEjphs8fvNompi52glRnBw8cU/GQTx/6M2mjauoda+v2Q3NVukUYUijFzsOWh
zuj/6q7cYVyljFFbGR/HL49PCorWmF7hW9QIXkAXvrpn8MNqozaxvT1GVFHvpaVu
YfFKsaq/koqrAZyn9B++c5IRCdyl4TF5W5eOUvavGat0NPjstmqqNJNtIYo9b1eh
6tOuWhEPeStOjQ71wf/p2HfnlJtMAnaEyJwc6Q6Y38yA5E86a0CMQwjbm58/4zvL
5DXGC8RZ4wvfL0WN/iQb/Y0Klg8PHpfIAZEFWvGAyhMF87bRXYi9hAVRViqaA8NT
pERGrwaV1DpSN3ldpa8oRrnuO/fSxFqViskyvchGxookuxdUVTDvyTzA40xnSEln
LpYD1KY+fH+bsAXiNIn00x6zBYvv0Jm+/Q5f+FIZUlAOWtOvdSNPrQNAPwXrbg+g
dGXpA5Ij5MtK/XeBYVg5FrXEA7JZ7eJjcPYPIiF1Y4GOZxwnYLuPvOGAXuMFAQ5m
BvwX3SmvzwlAU6+3BbcUL7EQV6oNaWcDEe5m+KCCbpKDPDwpP51rSYv2QlXuwUZ9
usR81UTv+vqF/7DNzSwZ9+tZd6bZqueJMgvfS76OWGY2rPnix0tcYIpQkNJ+uwt6
n6T4w0fiOrjvH5EfPaiKPgs+0jjuJTegi4jX4/HOBL/c/zXc08NdrUSxbdm2tCHj
DfnNoUAWOE9a4X0z7oS35i28vbptVuXjh7FYMzV0W/xzXkt22MwD6QmhfFIy8ko6
1/A/1T5uh8PhmQspkE6Sz9j/OVLNzdf7ENOYX8AvIDu96h4SqxkuhSPTk0pJyYCv
VsmcbDi6MjkWkEJA0vBeuWu5AaZdqRxipoISpC6xrePVjQouIg8AlF5Nk7ld4/fD
VjhUDExrFbIRoD01Pbmo7anTQBiCfUIe1rWZV3Zh8OT/GVbAIL5c90tRakwDUh47
vmcWwFJ/42TUobdBJZFnHkIV55Ys1h2t/HkteP+YOo/AffVGhXerUeZ/36VC29wF
zKc/0FILgq+2xzsPL79woxGiKlqA6yLBGPHsW+0dRxKfaskNWnYzffL1e89DG57m
lJij4MWsyZjo+PbDISA43DfdK+4jZ0rjgqgVeHAv+o/nziHDA5rx+bXkRx3/55A7
0cbk7TWaAEk+R9lMPgZ16jl5c+U50K1Pbb9lSSnIjYQsKhYhkXdcd+kgirkXWNMI
mAjbGanP35MPQ6E/p8/20+nL9Idwkgj2Fxl8XI1tAzQ+Svk6soHHa3BSURt60AwK
tC1SViXNw15ihfzry87bBTBojhfMEkdTz1DmDQc1QWUftN/1WZVpjRvJHVk35wsn
8BReBWuxWfSyFzCp/kLY0AoI+qNDtGeb4w4m63DxjqnzZzNJPNmQqNaelNgAD88P
CYqJgSHHGIMlSyvkJkYTkcI0uJ1WpPnj6v8IrsQovPn11beXaFnN71IPBBnzTSvy
bI9YVSQlKI98KJ1C1enMTBj80GSZvkIWLMOPl7vdsXaIgZabs2X8LFzsU07DB1eh
tMiWk+x+epod2RpTr0ZfjZ0/F6/OFAxvWv2AhdPZJdMEWkyvPf8dxFX+dKnD0NPW
kujW7+qvSjfWeVYomXtvaryEGpHF+cvXHPwQkWe3WuJDRrUCqNTOxOh8/LLPLKjl
B+uikRmbFv02S87iDZmpGnlKsVe21SR2omsn7bpast16D1htGiOV51VCYnJveKOX
VnpODgRD27gyk6cHdyYmDbg5b3oCiAwTQ5vMM7nHdlqnHd7ZF1flOs96zJcBU6t8
p3wNs1FcJOtVYIcF9DzcKsC/XNaOl812lSMqtGb/2OEiGqOYH0Kfgz2a09ROfYVx
V91wqOgiIPNR3ZfuKY6n8pffVLzv1PPnLSMDPvg0LuiycQr7+RfgRZ5QEIFGU6Cn
JyMtspgW3SrsOGNL/i8zXI5l/c8qLQLy+4L3GxF6K0mhcohLqvSYbcwXpGAGGoGL
OMqeH+BUnNy3vMZOEcTu0ll14ycwJIMvBPsv063Cpn+6DZVHmLNDvC2tnIbQM/+F
DjxmJsLd2AJEV1yIoFBbtq19NYahKcXOw/MgkaX+OUgGJJaY7WjKewo4Ckv0hD+t
5V3EWEOwVRTaF3Uo4cUB6d/HDwnT4x/N9VbjmIAvpncR5QXlT98UwpsYWnPpoerg
4ux7F8YiP63a2QZNbTunM4ePvZxq0AZc7baDA/Uxrhg2GKWXfJ7cJ6cv99r4bhFh
fyKd0ejTpsYgacIxIf3WlMOqOvPBqW3H+gqNuGzT61y75lVCZmORHI/wbdmLBI5g
LSmz5W0eWBp3tPEuemQ9b41sndErf3cEG/ZknvMHFdT20NYpDrDcWe5qhkr0n9hU
hsduqW2DNbFru1oCB0m4oLHi9wx3J/AwxaKzFvTIZh9tRIWH9NUPTUOTV4HRpuNB
+kVHYzr7VEwkLgSTssh5eCtajD/u/1oMqvbPb3QPrSuJkSVz1mFrkFNO+H6eWM9L
oq8ZajcOgUadsdYSEESeLOTAVy/AOXN8Vaf1DUxj26Iyrk/9+Wgagd3ZA8lsCt0A
oZXijgCj185CIGQx4p9QWj19iygZxKrD9Ws1jp05LLh+KlFR+g1bnWJinSunNiFs
A4wnBoX7I1SPV42U5ZHX8GE+8b2vbIatlDkKndJDbu6NYGzdCGNvDB5QznPVuCBY
+QCXObI3bhj3BVvM2g3K6IXlDw2ZR0oL69MUufDyqWZFmLwtUcg3Fk6jMfDtyKxh
Zin9y3UpiRWmU0CYQ1ed3wGTvmr5EkTmz8JXSedGQDBqajWDfk8/6UnTJxoTrqs/
1XUbzZcVysU7wSbcLdXx6HrL3aX0NxXXRESpIG95mnBO1dOrP3jkOhxMIVfGx3hW
qw5h+EuFhl+hszBWHU3O00Cs0gEVDQLOnUnjd98GuKvVAaYxRD3E8TmNy7OsroDI
YBV4VKznpwgGjU3BHduO1efQ9m2wNjy3swAcCzvol1SLpuOb5MVICLj4o98rxI/a
NBz/XdFUo724dhbE6oPNJd6+8qX5rv0RXuOjLUfLKSP2TPCYP8Ll34hhYHKc5xRQ
fmo7yR9TxJArMFzB4itVwuU7MhKJvgNRG+eNuj7PPvuMOS3BlQmL2ZHMoJzs/N53
1Em8xatayl4+fRnobMM/Pbu6BLybMeo8Na2raGutv41Zh/W1sl5+CzJYF5mAlDgQ
hHxfkTOXzZp0JRTgudrqL7iJWGz4C/yCHk0IhE+YQscM6jDl0gTuR6yz7Ap3NwW5
mxvXtfD6j43l5mdDmQAp7PGGYWWqMU5ZYECvtA3fr27oWTqMqB56JYMRzluv8uZs
zSnJR8E4KboFK8TRkn5ZS+4aXJvBL+Sd8DaxvdMh51VrxPKfVPtvTfyfWkM9n5zs
7MzoIDo883Lz/9RWcZZCr29Q4r9UD7Mp+lAhiflhgUtiA9vVpH1FXMEA9rNCzOHN
BP2TyIqAM039FI5KDqZsyRL33pqNm/3eiapoiusSmO84Z9HumbhQx6+AmXHK0Z4Y
4lZDoh5U01guMUv/HFWY2royX6geJ+VMaeot9/uTwu0545R1LWVGHKk4I9HI/Sky
FdEWfAQ8kjapj/eFFmZuaacNC4Oyf7qiUELgydVNLkhb8iF4jNh2n/95dr1r5jnv
onzZiS17KS2L19L+3CKpqFNHAvyBPqwbRVTGbe1b4iQsbOzGWyMkOFD1aLnvQ5kr
tlD/R8C/A3DeNojSUywcFhi9SF5rCFZyQ+g5EIg3X/ZboLlGUtoCZKbYJMuvhHCL
hdorgwoSnf7jTxdIxJFeYP6OY18i/y37VqsFUHM3mMQhjytbeg9Y8vir4gc73R6m
4qWmHkofvqWQwOarVZ74b7w0Akf7mOR8/CYXj4ksGF35zAgMP9tvMe29qG/JwdQz
ldmpNXHtN7AyzP6ILRFCuEPG8+N273JDuXwICQuHzoOBiUJPdpgenVd1tFTp887x
rSenuxjuLzh8JpdtCKhMcM65ipdbIE5rWyL8zOg6VOON9FWWYWGx3DeU5JtFh2ll
YPQgn9S9pIRyvAjXeKofpEzLqBKHbLFMG2KF9i10+l5LPB0iTYhX4jxUXTsI6Ul7
DZZQYo31CEiEUH5q0rMwbzEkyQ7pZf9ZtSnS1e/ZKAfj5ZZNS7TRkRoa9fgECFd3
GyGqKuEbHgaFVvgpUw15LAm2JgWYmQBIRCHht8QDmb0BIWhwq9WFcOzqn1f8waqH
DczZdfFz2TGp0HsnC59I7MemsFmOfmyIixgC0Vurl90SHtHFwtQbL+t/W1LCIoHA
hO7PQflHluQy+cXPe6IgNsslk5tXPAFameLaYWEFFth4w3jmQwgkolLFiWTb63Pg
f6D2LUqDGcG6NBHzBUEs5H//Vxs6oc/WydoVxs91h9sbhqYEnmkFwfd80D7qsFQl
DcAtBrFCokPmX9F/0dLu9SiEdBDJiGjYKSFTg1pZmt1LuaFCzevFjlSt3bZrUZTJ
46jxUFMEcSS7qHCJuXk7aw7OJUoKSP+wSg4W/M9WPJpnEezlWOv6t9gTrobjIArW
JoOMGtUq6zaw+sIbMQDxUe3t29tILT+TFD4X3wpZt312+0hI+4ijSgaN6OJX/WXG
4PdElKAQAsXhKSnuL6RxmE7R530y0JLAie4IGzZv1O9ttmEk/zOdUc0q/wGVH2xw
8myxFREbXaJAsZbL/z+H3bfAzPejnj93mus992j5QBSuGcOwIp1chl5eNgyH8gRl
fMrSeYl19kWNFtyWGrpxEUY1+pc5FuV4Qc/keNQbNcPzReT/w+Gr+894zYdp+NZK
mrp2H87TPKP0KyoKAG/CUlV5TfY8LUxyKmveGpDFZor38RZsA8qX+7euG3qodSxn
dTHO3gytvABg46M8oSC8diPQBy1BqCn8+w56csrrR8AtKZQ/U+4lC28VaVsVqPon
G4bczMCtIpbCi/6h2KtiuoH8udXD3M8JCws8NYKKoHkw86Hxebqod5m0JiZUXweC
T5NUHKIuwAKwKxTUybA9fr7g7AwHBtDhmSsHDbMzQuYPNJC4Vio76Yb1ySjEQhC9
FzQcDeZkK2AmPg/VapShQtv0gTwPJFe5GI11LE4YxKFW61tgEj+0iQVa/0tnc2dm
QMuIjQ5Wjz3BGhiUdjPBvMR92wlP/qfeqU+6x6VkjduuPX8sqwotoYMmd/+jAXv3
fBpyJJX/vyyXTXmFGnoKFYTmWgJYsEqKMGE/gZ5w/60y+1p274/ryG9cIFatPYgq
zHsb0KqZce4d3fQOUb/z3XvgidEW8mvaLMfKYgu1/86mFzvXLl4GDBxkaGWog5n/
3kM1p9mdX5FBkMY3go5C/a2J5s3hckycLYrllp+0/18gHAAWp6s8NAzey9J2e/G/
RqlwtlsrVyl42j7mPPKzGQ+ieD/+KaCMf9rZ/odDQx/ueP2QueimEOSEqzhdh6vx
M1d/XoSmsKzLod8uBmVjWUcjNaKVZKhhk8umZXdnrwpKqpqXCNnWZXh2V7Q2+GT2
EfuOnJg534u5u10GeGgK8DAC2JuqUx7H6EdOsCdypB/FIFpXA+486ZrjJ0ocAJuT
y/+0NW7BpdMaiNgpHb5/6sR9Wid4MA5VPT4lSAoppwWx5fTCKgGpVTLElQuTP7d1
JH4mqg47Qo3Or8br5MIGjNvKqBHkyRVVxffO0CV6f7pLwHvMQSzwN7/YxA3NU5/q
mX9lgAzBIxcpF+3yjAyewiithEIz3zkjdx211C/sICyfPvfGr9Rl1pmQ+WeTdJGI
gNY7Auh59oIAHGGYPOERD9Qr7P+wwdC1kW4Ugsy1Oi0BGOSmGCE8uKBPRkGT2DEE
JQQfilSLjIwLo7QciyukzS9/M3pincJiW5zRUvHHzh4YIYK6kGfJ2nPl3/Uj2BpL
eKHgaWxvtsd+4IwXn2kK6dRpoRhxBImKAukqvTw46lJHOFm8tWfJz9skddb7mn2q
XFMbhwKQ6L8nbwNlfyIpJd53IB2rteNN+Gm71Af0CF6XddG2SVmaxhTEUPxg/R0l
IC4lgzkwpliE7s+ETUxa4Ci4zUdsl3WDTEt97BIRrfSVP1l38SQv5zipmj24tpBS
IGANZiybvoFsvcI5hmDC+YwIxnZiHPtKtizkN2HbVtI23936FtrTntb9Yd4mgU/0
KebKanm7wUDS+f8jsqYP4yunV2fZw0fEzhMIbSQ+MRyhxUJyQj5dlmy7DIe2qm7i
fFUd51/RCmx/y5Jip33gAJQiD4rrvQntTTWsJdw3b7405H7Zx7Uj3NaSed2d7Nhx
yWktXUOJm8nZy7Bfbf9jnNiVcumlu/RRPtOqQf8R5hJoGImbQyiXaSbJh3cTLsLb
801kSUOscFY5XzGQISKdu0XivGTJcoVuO6NWie4ToMyqfs7ZyaaN2eiye5GKIWPx
7tiizIbqc8A0WXwzUrGSzoK7y5g+9cE+j/+aDSqw5kqNOsaODL6aEG92pLLlbQmI
mm0nYk+5HP94DZwnBGDaSGnZEiqJ0QzcW28dknyJyr5hfCTwh1t0yJUFYJUD53by
G7YQ/s5BeUmDZQyJ1sPwwLPJ/JHlSMcPWHxWqp9gEIedSzS+vtc7bbtKjaIyWnwu
3of/UVnS2MTBj8w2SOsUWyHpQUUeYEN0uhhs9nhmddnGoOkzeR/W5vbN8v6QBm4j
wNo11UIccdX0+Kh0pf4BIS61vMm70DAOOqfHTMfJPidlYu6Uz17QzKmcBbhFvWEX
obApTucEfiFZUchyrrCJK3x30GZItrhq2RPSXLSrf48Hca9561yE8C482atc7JkB
p8zTmpW7Dm1NbNG6OzlHdP9uq0EXRGcb0ugs65SzZUqdDs1MeVWtzKBAf5t2/Mup
2QbhRPpACKOsS71d+QYn52oL075/1X/gQhZBWvDHqiNdNABL7qDFCG5Y8z2/8yOj
nCyjNxG2vGrwLkFaFuN8FPbMZ1qZIlArBukT1amScNo9dD07KbCzIj3LEojnFa6W
VaWPIjCd8BykaHxEt0TFh3HTcReGZAg0E52g2KqZxiB2I1KdN468QW0UY/WAfuOv
SgbplBIMX7mlKxBlhZpelXV062nVw9g9mdEGA8L1EaWUw7ISDZAZcUuvwLXnuvDz
AegjPjwmfYRyFACmthtLIR+qhIvtsqUoujrZZeqKaX2U4VsnJizRaMvhJrJfGYUq
zm20gv703L2hwI2RTBy8BTRdUZsePgIfh4Cwa1l8wp1XSqKqAvOPNffc2yOB9g9p
udzQuTgTufY9SDEUGHncCv7v2EQOo8Md8upufZxNgqDB+O0FTPSuEM4oFLyBgcau
6/Tyvtj75g3YC+DN/uRGFf7F4/tIG/6D8eCpYzZitXMbTUIcrgkm4zO1hVWq6r3N
5PBehU2yq2jfbR4Es+Zno7lg1s8fmALmVt+IfgwSvtSnGh0NrLz06eI6kydCudDp
MGxRxDjXEsSLkXF7BfyreZzG6dpr2o2O9ml2eY2iLazPcpZ5Hvwn1AcSjknBu73Y
sE2VrKNkYOT4UuhpV8lZeUVPoocw0SoceGl0cRPa7W3DSHsSA98uqsNwmab8lWeq
BqovhJIdLYgdfC77/6YD/btOoigLl4MNrbO0vNbjVQjCkwba6YvCWx9I1oe0ojnj
xwqJNjQFMRid27pisvdRE89f5Pa3Atgc26SXhFjwCKGYosZl91BMwe++q3sgdkJ1
0bTAiRaaObWX4s6k22RijRJNyl3RHZ5rN9wYbsoc+v4v1drpLUTF4I1RNLiWVzi6
rn9tyZ5IdQAaC6RJyTwK3R0DVRy0RD02Cal9+pmIlablQwIPbX/8by5G0KuxZSoG
4KJH2M0UEQWSImggaq7MOIC9oYlor3/6R16qPhl7ajqxm+Hvt+0yUMbUynoz1+ex
XpXrA1Bj+tsJO4eAW+G0IoB6yRFu7jsZq5Njh+C5RuktxI7EL1SX1MxRsjF0UOfX
IAioLFtgJbSOOfDBCRUnYmEF39E5HUlRFV3miXYuFGNilDqMD38hJV87lQxWgt2k
HxWNtF60do8BW7Cunp42mIN14aZY9GPSTH9bakMdgRBmG6ozTVKKOTq4xtFihago
hzPpJPmUZDNSbqcbQtWL+tDPwElDZ4nBNaw0BV6Ka7GFbrpFFNhTaOIdRr74HzLn
w+kNGd3jzdb5J1RMrHXlxxJcIYFT0O0CFvfSxgOMMumQvFfqTD4ood7vN1puhufS
7fldTJ7bdCEHTb8Y3tcMUe5ZqegnhgxooxPvAcBVE5lwkFYriT2Hid/M1wws6Ayp
zpgoby61vGqKRxhpynToF3ECLBHCf2QJLTcDxysuL1+lGVPfSyQkAgf/lNnwKqKf
B5dHcx4d54mSKOYQWvznrKQh49sKs2ZrF1l7P+Ai0KqGUfKvI9fmbAiTDnVfqqmG
G3UqsHqSbp56vIVBBEIxjIbIBxvOpAyl7avrTpol1K9hEJyknMAKKP8lWslRH+Qr
enw9jRuNUNPkk7gW2nDuXSperLlCMhylas6wjQliM97+JjSRS+l47AF+c8h2bvKb
Dzu1Kd2VrF98GAGBwrKjGkDy88GDXoKwmqum7uC9ISNFlwTjFORlhW/emfClGTdW
7ynNIc0uXTrMVd16tOWDThkDKczKuxF0uEZGETTJIYgckVbSNgFLiG0nPJ3OyaIj
bc2PMhNQ070wssYSWC83iYGGGIkiKOHrtcAZEYmt5StqDq+76yyUpZ2erZClOjr/
OO+3ck6GXCjAYR7IpNIQOH0EIBsgiro7l8Jnni+LJMR/LQELricK1p4p/S7XPWPB
5wUcLqieFqqNmCql+U2M/ncxssSSg2IpGD9Loe7j26dinkSl5TfV8xxRmSM+K2I9
z+efgqDmWMuLt9ibvQ4HeTxaNyOiDTuNXgt/3+T558d1yYQccYgqbJw1qePFHgKI
qAYspDZxHiyYIARnFNm9pF+tyAR/ObF6/ywT9V5X8kRyFWr6PSv7Kva1sYzAPrsr
kf+Pr/oJxi0NGrXaSlF+HumBzWDtD4i2kA2rzLX08D34ps6aolM7gkx/0nUDpGcb
j8Ha+i8VbFPmB1N6Ot3kzJjE1dN9zGdnZtnIwsSoWDJFxVHCQKri2HEbaoXskn85
Wn5Q4hw1y2UesoI59gfdoyDQcCebp6gMkc5ggZTW/KsaBTQiwn+J7eORrHXLhV6e
CtrN+t9f3yyugvOpcv4+usl/s6DBwSwxtaSfwi9cuND/HPfZ3gIpqbylEhHUEFbc
BI3pVyLL5UW98KG1P2YMo+3OgZfh8UfJ8LSlHxinCd6pgc7PHhxch7JbqpmmsB2Y
YK8Cgs7RHVPMaukRn6F7KikL3lZKGRo9wqtktsefmmEdOfTeF46ViJpO0KR+PbXb
vlrylYnESCwTpmXLr3QlEerk+rqY4j9gdQ6Km6OpPYS+snRByEUIcM/yR77PPkry
EPcZWKTnzX6wvIHcq06VaqIBSF9uaWzFMmdlGfvrlNYGRsFiVBVIDAOka+/lAyHe
JoEjTWBVFrrNGQjU81XljFDEaIDOYaQgTSLWMJp4bz3EyhTQlI3a2ivw6LsVZczT
DiVeObeir0P/wxfBVDbwljFntZle4h9MdhiLeZVJqtXzIlMp7fzfybBTPrbKnmCY
j9qYJ1RKcGuWqguy+Xln76rCRwXt6EeIV8PizMmgvqhfVRXvBEQngquq8sZX38sY
5VVtt+OwkVLU0pvrpba9xMfycWhUHuytU5PpW6XUv2shk9cX0bWYHI4pvEsLCi5D
Bfjfg2qn7KuoTSQOmENMe5mvXk78EAdECX/4DUwdv4V1kbGr9tFoDmK6WBttKeyU
xcI8z9YN4wVJRMZ8D8Tv3zSDt8qjXemG0Lkd9so/nnWnh5DLMj/EcUaSYQkpVs3I
i/9jBrdhK/Y9okYzJns/lxoHZauF6v84brNEq7lVmQkHjNaJGa6nKhac0xyXnzlC
/4qnEbwCl8ylk0ya1tdy/yb7rAkMRRN7VmCwXbm1C8cRaDMhXY9/AsHacAxB/onM
P9xo96VDEOTHA68d9/zdHzf+gc5WCwiE+rOGSZRB9s/yHUsDKHLzCL3JKggiGQmG
wEaPWf12RW9YhxghhoVf+kkREmQ+rXLIwvHUV5xwFnWaCl8gAPrh9atvNXCvYbI/
zc0Ex0nys1qsQWO03W8byXUPNgLCPZSG2Qo2F3fqz3PbnhjYN0Ns11VtRfSS4hi5
zg4eQF5TV/Kp+4KJzYSLuGiMAW7v+YmwUZQCr/VamGuZJrDdlgceeycjG/J/wjLw
SVYa4YEq0KeKhQenCGe889A5Wci6WC25M3OE3Opz3M3Ml7Q0A8a9FBbje2dWW9Ny
lwZbSU9nM4jDoSjF30XMnqbeRddlQEsFXYcI1JlSJuQcZTQr19vtCjlPMU32gD54
Yn7bNU1HWU+7OD12YEUq6gnCm+Sr2tHGlgVSwydRvR2VcT0mEv5KwRYUGHndS2S2
ZTelQqGyP68VyTOR7D/wuVpvLlNqut9cvLEsLjy2X8Y2GeCDb+MgeJFZWg952F8M
UPVjg7DU7L79SO8++1giwpsYjPFQ/0V22X/X0ssakGUNz1ISJjBG3Ah9fDMRYG+E
+SxRnMOA313Pfj54diwIpJyl6hFRacyd65aYLGdUlqbofIPl+bBmAj65Nyfvl8rY
saMS87IyvPA8QLJsg+0jbGAwF26OXLLxM5329rKw4qThxWiRzVl8G/PQ1QB89ohH
g97MdWSqgpo/4KMXQnFpj9jsPbjUiXHLdptEUHfgwxAIpC8IyT5J09bdLbameXsc
u0Dqcyt5/9om2shfNvvC+tCXRmQWxPsNgfT8TfCKcddL4JtxPn7NYzOzdXn9HOS7
S/FljISiW7OBMZ6XnDUSAbx3YwRRnt2GJY41Z4cD7o+Xz5Blyyy5cwZk295Ekw2l
yzIn2x98ewQUrMXHNyDXeD02EHmrbZxXpV6tE++otYu2o7wVVdL4YrNg0c+747lA
0UXh34xqG80inipmQoEY1aUWXkYaS1iZP2rpKORh4jDkicA2e+Ph0E/QPQcPgyWT
zMjqiT54XoAT6Pnd7xAykXHD7Uyzvq6x2KD/BdPlU/0py5xj7MgWBaWkLVZnSxf+
EKhJcJhrijEWJKF2Ks3TShK8xAzYDw3ukYeBeQT6wD9rLsWUQwJeil5f8Bun9doH
7TUOsbMDm9mItwBtSTNDwJSWED10eFxWNOTsrn6GdmfOUpE5JpmpsDFK55/v7Lcf
uu1vx9hAcWmNLgzFZ0LDfo1uHlOA43Nz3RythTy3RBXKYLJxfrOJhrC4go6YCs9P
szPx3VjsH1V54VbTt4D7mnorZR8P0+9iS2lQsPlT0sYdAD3Gj3QxmLl8ao54ZtMA
dH+X/hUmnVV1JqUcrCd1kG/GWWoonyHYIwIFm1rGAVIkpnWgkYNRjsNfIWzthah3
rJ/6hFQI4uNyaK51XC2jADT0C79lbRr/KIevweJpNnlNlsqeScTnCVZou6XTyt38
xExXeRK/CbK4lhbs2jd82eM49mB4HBhFEQRcfbZ7SBSvLDctMvfvOtE9o7bMzORX
Pov6fuvYZcYbVPfDN32lg9oFZaD1DhmMalmyKbHvLvapPwbDMXaGONpJCzOtx9kF
UcTPwztM1omKgfZuyIbfhfkXtBy2sPCI25M/JBJT/BZWRtdyVd369JdcYndrvYBT
S6sRbjrJuIvoTPfX8Aqf/REuMyodz4xx/MsuKKO+aLcaCC1oyG8XwIwG9pYxdFUG
OgVAXvYPyCiN8adWLsL69A/7aHosHopXgIWpyMOnd1HhC59C1DLrGM1KK+M9QU8s
D9ugrepEHmFd7Qf8A4IeHKX/u6EtIm4u3pOIGzaN8CzNRsXAukYWfZEAYyhZuuAQ
Vj4jAvlsUB+HimjFKVUN5yO8baQUL2FIcffax+BMVKdLE4DZHtE4HnGT7meLRHe5
kzoOq58ZIqOXpzMvPiz0s5y/YnZHazen5iNisxMHL/mC+qLFv9glmaigfGrJcpyA
hJuI+bzXDlC4EcOgBtvM3ooF1yXUkthl2NNDvtI9wy0kWepedNs4bHm4fVzjK84Z
JZQ1nMtgpNIGY90mXXBf03uUAgVL3hE+BQ83s3T6UovLav8BBWwD6rP1fOhqV2gb
mtrqXIth+cfGQ0v5TPd3IH0NZTjJLvFEWXdeCHKL2pVmwm0yVvKget4CUPeK1Xn9
WgvykdyOFQYTAuDqfjrOqL0f7IKYPUHwWhY9D9tpTjqRSaU6P6zxNd2U7V4jtlp0
fRXcPgSOuX9lndTGoZIUyORsh+MBjze0aG8hJGLTjc3kBYqSTBy9tCmEw7sEbrCj
PCStVO3nHIVmAbPD66Hg3P95tN1RX0gtROq6zHcnfjR7B4vY/gyF0LFxXbv+KdsJ
PTtZ9wTdFs2vi+Y9A18ZkSoYgaHLdXQG0nvkOe6uokbb2NjtrxzQyF1ExuGqtjE0
jYUv793D+G+6ycjT3TLCtxAyEawfGRY3z8S4vSekB0k8VinaId26OFF0Q5cX+TEh
eArId+giLBsVDuWBadbwuT8Q6JRoxcuESoRMLXFU0uvVPV32UlLXDhkvxnL/Kz51
Hv5Foq4FH8oUF5ojh2FJhEXXJ3J+ghQfJBidtJi2p5UUK3vYhWfdRPvHbqZ9VeM9
YNEJG7FvSY0TulqNLXYwb5/6VuVvm6N+1DBFX8FcRprcqG/DnlicSsxR4Lqo9hY5
D5zxm4zSo5p1jA0CEqV5ir5Fv4THuMs79hWK0fKybfazyrEhKj/3Fcdn+CPWO34y
KhqJYahHcuw70JweYgK3+okWDlWnM483pmWZJOd/d7mV0aPY1051/f3VvTzw0v27
79HJ073fAEB6YFmfYdHKKhNAqFHu63bjD0vsuacCADowHh4K/Tv049pfB+RACmWh
/jVQig9o8+IJ7Hm8ss2I7tMrHVSCD6Dr5dPlhAyOKskB6aWmLqDt/MBB935LmJ0D
Eke8GvMqiCqH7DwKvuYMOynEY/CmPd8tTPSGG+YoIpBUDBCEF8hIpnp5mgjumsVJ
xKQygIfAmx5/bWUqc6WZh2UhZtxQ0SYfN8Kb9o/X7UIahRUFAbwRfMSWu3aybBTi
r6f06Gf6cVh6WdQIaRIOuMw2yaMbGiBtazZCVRdwY6/SzU33kkFyLmM0kp2oJ6Aj
Ymi+FG0LgdX445fDwubRck+PKx/UBGG7hOIsl/93OUn1bP5jdhfZEJXyFIygyJ1P
kvicKzosU1Lm2bgfhqrt3NExuKja/JWeSTuOyxg17D4BcJ5GrIBXFy+6XbqdVblf
FxsYqO3xs+YH32EMOR3b2XzNeWqbhQTMYYmurS9w8kMUBl5H26nSBPCADt54uv8Y
8RqOYawYeOjcpDPKQPMvee5qQtz4PxdKLiAz7b1eSnUG9v5I0uqMZyP7q2jFde21
phGdM8Q1R1O2r3VtIHYtHjt8kEkc8sVuXCCNGj7IXhLVh36aV9HRLXdbIINrfbHw
WXuM32L7UID266VwUdeWG4plW8PXaWkDiKNJnjPEUB2DslP7HXj0lTzNB9hLRE0t
Z9bj5/z3dwmi0GHd0JA+hEz38UpCv5u9Uu8t4+79M037JWC6NgTwlXArSCnSFwIX
lwdRb4q2uT2a5q5o6N6JvCmJehr6kXAzIztciQHE58ShtVF/NE8IHPYns2a/lLJD
MPG0XOV70FX102jzXLtIVqRgH8tUaFYs0rUJkwR+2w2IJLYKQzSU6njELngg3/uB
zFVy8eFDSD+BYvZQdu8h41CEJUntefzoQG/O7CRSAtkv2BWHmBUXWBW57wzdOxZN
I0YO014rgnYlNK4cyysDw1P8mCWJMH3Zzd/f/lsme2WYl0HJ5oKXt7NsTuX8ZS4h
0Kwc6cK6Y2O2PMzRFZ4q8YsPtyAJZJLgc8EwWuCspZDcZHj141kE9K+4qPYICTZe
lTdLFb8JiPIKdM14KPBiKJ8kCza7rwYuPTS4OVVhErwlG8yS84e4G0Zb9KUeVyzd
/zWul379y0ZIIc8UEaquVuIjoYlV7S7R2ujQ+Io3c5uOU1r9xqcjjg2WSUdMqCN1
05I9m26OLS+1a2Apf8r1avkrn2z0AFwImYptONkbPsU2uGzd79RRP9hS2RLS+XOy
CDX9BapuXLPtT42zf4PNTZ6e+c4sOcQEH/IJbGejE5ssrxOfFUjQTCG1bgZ4CWSn
aAuAZXlpJUcQiFoOLgW9d+uIOOyc645HPCQ5fpq2EO49ud22iLAy3odKczqIc5cP
U1A2g4aJ3UA8Wz7P06IzQ1SRlyiNYMXNEfHglvLJ52mYMyn5w89ZP2IQgmPVcjkW
ChlCsiY82VlcG7CocxPJlwUwzphpK7sjQAIVO+4yHroeeZPsJokHywBIabHNpsZz
7YvZmtZexMUOMjhoqAnz/cWuFxlHYEZxp7F5vJ+7kEId9bnqv4nzJZpEhU5SRAzx
OHHQCUArHQnDZ1dA4QCJR/ffKD2bYlPwb0k9OSONLb6KAq+pRZ9M30wVvKvf7wE0
jUknsA9mZZmUZjy1UBjToYiYUhWyCVm2moB3TghVn6EAyhJdSY18sTB8Y3eelGpc
yoGqnz06plHBKdxbxWRGM8cWjz+Bm3Tp+0Gb8ouEYZ7aPzPoEEjnzBwfrU/uDCIM
D3H21775FPxjyVoppNIJw5W2ps7v5Qg/5fkcFVVxZRi9uLvGnsVhL1G23FD7dyWd
H1MIJFdLDN/4Rn04C5zGKpY+/l2TUegshHBFv9L7LoTi2V6lTcVh0n6OgG2H/XLa
K31dH/XhMHZGL5pnsfakyge8HOU7T6VTvcz7+IgbYirqvpim4ccz18NcYW7tK7D4
TuHHNJAwCIjaFOsvby0yK9XsouTNVtbpJLxXSTJl97OHamDjZenCY6nranPEWbxe
nFtCzQvYNaQsSRQJUa2MGF+l9JYNr6M8KM8/3KDHW/UgwdxEsyzUxzS15EH4PpJ0
HYPUm//R140pP6Tmb8LHXXT/H/1htpoAEAEUkPAjBOQuqs39hJz3IkpgsWK3z3jF
Y4QKCG1L8vknJDAr9T605tARyysIxfKtIPPo7yllhmZHM7ncxFlTUjePsvhsZXtR
DRhGPI6XvTYcujXSJ13/dmYp7W3WsFXExE2U/rEZdGXU6VO3rl63W8rwKSlS4Gd4
0KUDXJFCG7Ui9vI2PPkboLzdnLwz4mvUdb+CaPjvboG25AvBk323geHyzoCz6pbA
bhJ0CVnzsyaBbCRTchwuIRPGoYkLtC87a6kV1zRNG8pBxeaiqd1ciaCHCvXmxURH
zn6RSW2FPFPxwm3UZu1nxnd4dDZQb/+QPc5b7VSt/LmAjDkLfVBirjZBFIzBfsLS
p8T8caWWD7QAOZywuqlIWP82bUGKLdpvjkeAbSm0d0QbcXqMUIGf0cz9+pSPFWRr
XQJOj2o0LYbpmBmj8cbnT6zD+T14eMn04mL80NTCF4F/KIu52kqed8h6e9pTxZQ7
QI/y70vs0z0TOShYphLrzWDCH/2mMaQ/4QiUKNTL7w1Ve7SOdqMbH57D7hOVqUch
TQecBlMkIZMVqb5J0RP1gFXnMj+RJ3Qo+XeLkxYAM+3pH1Obqyihfa7Q5NNUPyD2
BUTs371/igB/2oIsBbMBHo32u7MHBNuVDvDSG93FrIIsG9hFc2+2EJ/Ct7NzthFx
VqcpsVwQwNCPSKutGwpKheQkckM4AI47C+eXoenLjWkdOspREOtRn0DInQEXMKbt
9AKTQg7wwob4ycGDHpFwqK/FGM63jFwtJTcicWaq50Y6XrXGNx19sJB30XKz7EXw
KUNkTN7eqvK/mcmad23YtTuV/hMHQrRlvCNjEz60TbsyFs0veq74Gpq6uLC1SZLZ
hIAZVFdvsUdy/zK6dOU2l6etNfklV/fRT6wZN4o/dhthUYwEF60/bQOoSKNjVbN9
gE6KGhYM5baYLtoSKimY32vRGiKEubhuqu+xueQU129SuROFKCkuBzgEEFOiJ0KR
nZalYRdvj6SfwwariOE6AtLvxU6D1WxdCnll39s/4fJ5p0pxprYlt4mnr8W7Gt9l
oyMBuKOnRScCZNqpUHiiRXp7/NCbcb3gd7T+rrWggsrJY8IxrgN2WeAxk3ZhUvGT
SqRHUQbacl2MoWJf+bGVlRbaftjioRDwfYSt3VLG5wIbYN37IDTNA3pyDcYuem7P
QW0qF/mmvDk2JOF2/2qOwc6rr4xk7fKi97FeL+qLFfdkl/JfE+LX4uYjc2hQPF9r
YJliPTrFsCxEZB6TQpXOvW6pCLpZTFqajj4jVgT2z1ieIT9ww4ZHE8WdJ0rCFLCQ
CPf/1KcztOli0Fw00XO89CTIhopYCez2O3RVT93+NfLiQJPZaBVlNYswR7qxdTGJ
nBfxFAU3gnJ03NeUF4vsyOWcqymDPDEJb4qb86lT7sI7AXNpP64/5gb9hfweHXSN
4pEZLMK8NTjwynh8H23qbzxmnOen30yYswrasaKmV6IZfOMiIobU5/F+uqFYKh0R
MmL0LOx6VA5cT9F7GieFuiPKlAV3FrglWWm5XvBsCugWF5xoPQTtDuy/sj4CylN1
sTgepjoFEIMdwE2LlFDM7EgWD3DeIRAtzDJmzrc46rTYGM7CXRpwckISIHQNZGL7
ORbyLMivjZgXPnlOuZQrdCtWUYer4MzlDVm84buaZ7VnhaF0aMWQxGUWHyN3wsJ7
3/z+LCAjVY5klz9MvuW35WjJ6FiAPhfm2bbiZtxxAsZLfL1BVnCESJw/HmUNUxQ5
VjHXUlLW+SVfcTvSQ/vJ7dsAn397yqwrhyBUTPixW20TZcYTFBAJdnfzm22/XCT3
VeK82YZMpvWB6L6o/G9rXOXDZH8//Wte5+Auimnqt9Ysb1kBcnyffbsHLxQGcNMw
YySQFvM3uP+dQLp9T+8WPfAiWSlOvsR98qhQtLHXmgWSXyu6w6EtscaLrOo/dJ2x
4hzeGqgZWZtF+nRtaM7TKy1HJd+m1EimkuwUS2IK77nVyY5Cyp2hgLrsDeOP9Mz1
u6h/3L3veKVVEtQiRsvlK0Cs477fHcWH/1LF0wjCa2CUB61xrwujjvh0XiTcU/Kq
BLcFsl9Qkl03Isfk7h3wPLToQ5igh3pgSY0xS91TcY2th8CSnqWqZZeHaDSV60SI
+3MJQC1CBlhyTtdmrW8W9zVVgYeEKOzn7EauYZ3olNfOdUrFcdqrzrs52yAQxQ/k
r7u9MkIf1jyQyqZw24BQh9z3aX9Bf2YlticaX1Rw0NZHh81afXIJcbfsmtNHgmif
KlUwqRkY2OMqTwCE5PVXCrlaizv1ObPwG7JSJAyxaAauSZFgezWcMtPIIEJbOVLA
R0SuQxuOhhGo6mvk/g8tGr1JE7dnr+mocc3SV6NuAafy+StPzftv1ptqm3ldoHxd
99mzeRYi52HpI1Icu5vF4yom/maapgFwB2WNYahV6qr79+5JvcZS59sYk6AeZpFZ
ojIdQLRPDYa17N8M8i+7HOzlKuvrY9Esy2ry8TjEhFz98+0F16Uvs9nHz0jBgXZj
U3/OsspkiaznndrwzGxCRxZC+bDd1WWVQTq4XAyOI48tCqDBdZfjn59VJ0Z9CTyM
cPsUJEA1YMvIrRczyAUI7GJuMU4I2a319DfE7AUWmJk3iqlfkb65T4/ggm4wM5vT
FHNuSsbs8J6viRjHJGgfDZyZp5Tbyc8fdvXHtQjX6YVkivybKrZU+isU67+zcz1I
PXzYkv1CY6CvorJ/o49abMlLlbEfOGjH3T0Mw2YKahpq2sjWQQQWtDlw6Xv0GEg9
kscq95Cj5iWWY592HVIqQMZD/4kPxmRV/I1o/txSI93eSL4bk4fHsd+07rCgsn69
jpxbDSwl6cjmFhAZ3EMnp84HKorfxdyZ/kxT5RKa7mD58etmJM9q6t0J1AAIoB5z
jkfySW4aBSASCXVvlsH0/a/rrCLlhZdgRUEMYo8iyo/JAYlAxvRHv+0CybNgcEmN
cD53Gfy/MohmiC3z22Wse8lO9pV6SBt5zSigwmwJ8tzN8JV4E+ORv7mOfH63RkDx
NoEq1rMabC3WmF1xAAbNsCYS/bOeqZcfcSgj0TyInxK9zr+xobZZKrWYBXeot/C8
E9vl7WK12uEIE3JQrikElEbAKWSpqcx2nc11yCLGGNBbXVI2CIKSnLwqsk59DINg
9cJMvWNRG928TxrSkz1Duwmk6t6eKj6tLOYptLg8pzKdQiZ3kAoJAkeVJaPe9MTQ
PIF8ruXt7HC6KQoqz/qkPCsmN0PM2oww3g4aWGMlAbsqKXg5GOHU8DQ+Bv0AwfnY
tXYw5fcTrDMEBXrtaEmkhhz4NMJjpGZ0S0pQzZsJfp1eb/3LvQqwnTUVCbwpTreI
dDf1PoJPqvX4crTlJekqNcivLuRY60vvvBRdTCNf4n3K68Zidzu+yZHG5yeDn7Cx
b+j1EOPzpm1lN30wMtj3+1xemJ1/EECIvhDPvHhsfav0uAzFw+F1l9rqvTSKd5aX
+RV9lBO5pSfL9QfZUoB/jejaqQQ7jCE5m3Ww3+XswIwiLIxNDMQbMN7AFpyykum+
S/4jQPaPB4x/AhxD2wZ91GjZsgcumld//9WvUv9kZ2YTynNdFgpuCN3Rl8Pp5qlR
I4Bp62h8DNoZoDCwkyApRKXJIGIqurg150C4qXCMJpa7yxYNLvIxKibH3DYjC/Vf
9sVnsF6OuCPiq2T4Icrw0OPJiIHqoIFA0s9hYpVHobTirxg3OTMP7B0U6uoHdXs2
avp81zHakzbrYXM2dieK5N59u+GAntycit72Rss79s2Xekjogv94cNdFYO4ToLqV
F9pvHqEDU210XZ1/9nidMtTybYpUVREz6WogkQzddU4IwetVprk+aQajX4WfMFIX
XbnrEDkIQKg8F6i3zgd91vLkVAOvqG/Mr2GQzxwT0UN1XU+YJhyW1CvAhx1Ga/t1
n8IPrDzzK7lPjUekA4JPZ9a6cXBdA5fT7tS2fNXmoz0vB9eZna6lBgXRGcBLdVFc
2442Svbc+du9bj8wIbY38bxLH0s+i8JGEfFNIKPQWEFP/rIBA9tM4OC0P/pTxYBA
eHoVq4OnH3WsP2ty2CgnjWNiJ3HRzwusrAd3jd0MB+5Trhp8YbHWCAFBGW5zY3Cs
BBHBGsImjAfzTTPerBG98GMOIjExuIMa+MifS/WC2J8GRrPduWisdS7G6DYtZGdA
y9HhJvVpf2vdMjobHY+Vr2+jEc/1xFiVFxi+7FnXeKbCeMF/ooUmdzg1Qis1Z2b1
BjdlueS7Kau76pPktLMZ/C8thxL14hYGoqe2ZIWxsyPURRekRpNoxD2s6TFUZvbM
AMX8SwVwyI5Chj5SN4x0urnxcUfWxFdvaHpNu+TXNrKs6NFeO4m72b+j3inl5Kgo
C570je/Ooa6KYhEoalBQmysZMbmNu1tlQKxo/HUCEifXlyiXT3HzEvfz2E0gK2xw
XYQJhafk0A0I68p/ZdVd+L+B0XQ/EQcaCht0B9mfIaZbDXVI/wRGwVFcxkR1mHW5
1CwBUw2dSkSmMA96F7Yp8ERhIe4QhL3vIdR/MhMRyYaf8H7evQVnlx2Mcm2e20cW
OPIfx2EBRHk3BaPsnnXvlHPZnmxYGF7uQ9944pT885M4mrFyWDLwUO1wo2k+nW68
fV3bbRedKyJ0LUEbbnNPnk7dow4gGclKlRY8l5aHYIYB2AG/61NPtNRmgSNW2Gsi
6+w226YxHUjvozfQRN2+QxEwA0XeemZlS6VJxQU3zvtPSHEO1wjhFgT7lTRiZYim
V/XGhdTqlHYw/7zBEYtC3eWL8SulD0UhTP0QD90peaolvYNg75MAW25P42jKv3oT
hgGtCr/NtUSOxXREdjKXzF/0fh7VS0VC+vPtclLoZxKl1d36StP1Eb+ahNiJ+6Kk
JEmBMo1T4ZieUjo1RJBraNwsywXkRkOvO/WVhV7kjM13CPNoq00SPJACNcqKb59Z
4xm88IQ3xJjA5Gop0TJrQaJAgm0aCYHTCBRN/GDl3TBbz0jdP9U8K1D9NmxKN9ai
tOtmfvhIQRX5MGOzmqQmPfKJZyf704sWZ3xX9Mdw6XT7r7vQJNflsiy9P/ZiVa/O
ndUQetxg5Z5ZOucFMWM0yEemowrQc5P3XntYQsWUgUzTXTBet/wEmNEQwIvth4rj
h6CUM8eldvsbwljXMKj+1ehQ2GXQpq8A601ijAfD5JqXcJ9peYu6QOlIPaXtosHf
fs605IBY1uwccN7sY+gQ6t4ltjYb22XnvpcXGA9mKXi5rr7DibGgQsWAvK4R2FJG
DXjWLfN/htjq/16G/s65+2N+QHHc4VzQtROeSdXwZO/AfCWPLJGSNNJ3S+HEhug1
aSUTo+lKCwT9Zqc48ikAvcJBDH2N1xuZzlUW+rlTYdBysZIF90lrnXi9T+QmSasC
QK3OrxjQGIEc4mWJdyyhnQL02I0sv9r+VZMYj1Mr2a1x6AoWWCZPMcfwkETcf9Et
VFt0bTIMDIEBG4M+ppSN8DjPEXDfxN2pJFALm7L14WVgEHcoNcZGpY24l5zVtqJq
n7RH10ImM812A8qWAJGro0mqQWLTKk0wdd1q2HbxWOY48dgnc3DVCs6+q2T5cSh/
Oh7R0n7+4yK3oupACO3g8VMyzS8OnUbxU586q6jbQ+3JRwb/hk2CLWUyJMSJm1C8
cdlmnXxSHP5mmMNXT7E07cTVCIf1vUy4k2pj9EL69rXcO9yYYrrz21Ze34TLWb4W
aXSGdDpmkVGwjaH3NMlinKzCEze7p3LHnt5fBlHqiBgO6KzXYHx902BFfGtu7m47
3qybsUcv+b8KhNs4i97HNpuYciy5ppBFbdA0PPmCdYTIIxPWZLwuOfdkODSWQxk0
MO6XJyPYqbh6cq9vR/P61kUiJ7N9/1i9APvzGmp7ICEAfxLsvqcQcwPZEBFrVWL4
4ELqZzjDkiTO5JbwpO71u5jWlts+jDikGD1IZKw8qhOmhoTTM9VfV+HgycHS14bC
/At0bIB9Aeg5mgsj+1D0Xr1utkzSyVfV5w715Dkfi2oEnofbS31new4tzkDBqdBO
ZUwmC7NFZD3WA9pkZlsPUGfucU7ZzGogZJIGXGFU6GuXQH1a+vRqmjNpPZpFxfV7
01U9FRAB94zmEix7xZpB5mUOXKOD7BtLX71xtA7+0jHalElhKfiBHo6tddeQaYVD
INbJmd6BoKvokGtWLmFI4JbyqOxGDVBUrV22qPxRTJc2ez3ljGf+TGucwQPFKxxh
4rVuNcBAImoN1lNEl7ZNFvqEI82tq9fQR6PIEum/L8hmyg87pQoz68/13oGj7qak
EZgMx6uyfkIRAHUn0joMNEve8GISSwdfAzDmSmZpkiJiXd4/zdUcrjHKgpY39za4
cleuV9UH5lQLDU0KCTvx/+jtHdMUmXfBv855pBPCEsRBAC0R7D3nTWNoH6U8vjPt
A2KzNYhbtuhWcdxJNiHDoAZVf6JrE4/l5tHup+TgeJWGP08+dxx4dcvNAaBMLyda
sP+XZMcAtw6CiJoOHCtfrB++MRu6Ur+UmLQ3C5oPEKco+pp4n4D5GF6GYp+P96Oo
QhCHwOgit/zHnIpzjifBV/1zBzvS/oeGr46H7gGrCTSZTL/XjsxCYacsqmuOIp50
d53M+WHGXVWNAyFeTBX0F4Gp7J6yrwNa7uuLLR6uA5rV3K/ICbxvQHLqqt1623hq
WDzXT/aaFh3fKJ/wKObxiuSzqSq2A1+c/6+bvFBdhXOq6bbF7SNvmNSDk0EWGylI
nx9AzYyejtanipVK+oSyHKq72eH21CBu6eH3RsV9Ku+1xbKXBT3teiRVWatPj1Eh
/Qskm0ga5UohJ9YmAJrGSb5+IsrFeKF5dlImbH0Vv8MwCvkVJokUf6TSX2PRxyOA
GDDFqRLhr1eq4A/aGqFmyVNl1HRbQ8Qx44QCJQm7PnSbI70jKs3OVN2MD9MYkJwS
ZGPIHnrSQoB3Ojv+ZVpJ04ssB9qjei+93AI+ahVk16Lpadk43fdsv19/TtTSj4sl
/arCCn6td4P8Kj9r9DEezaJARg+iqkDGmnwVA0Cq9GziE5lbAcn/1/fk1F4ep7Ia
cj1Yd9OwRieGp5rgzNP/nc4SfcGGM3wmJ+WnWedNOCFcsmwLHEWYj+GQB0YUcuIu
CbVIakpvznWlxk2dKfZe4+znXb2ZOe6GN18gQw3Ioj5VX9GoFTWJQSJBNTnmeKog
gyguJ7s02WzKhhwThifXVXVq9w+reLdu33E3ufdEvFXlp5PY1CLONa2kwmoBWARg
wUIN/ZFgjs3x/rTxc/8X6EttWbslRd4LzwRS0GdDqGBD3t7qZMEUonW120o05vCW
tizGzk0MEJwyd3oCAHMjHR5xfnBS460Dyc8kkjU/rnuvv7fl5IXhG3hMMvGNtrc2
cl0QA8Mb+wqymNFgzFFv6as/xdNUEFeqj+zs/JQYbAWhyVVe23C7kySnswYrIQJq
M/RAxN+tIAAruKekOffnYdVAKNb09iOuxUEyqp+Mrj8boA5//2Byoca4WQrASoHO
p0+X8Ri+qKu+f4KP221e2dIKOnNkWBAVEQ/l/mAwOtdKdDsINoKqw78SJI7ojZip
9LIKbTjhOS6GogD378OWsENWi0MJgNIQUhgfJbde6BtyeImUpEDZf4Dl1VL3uuxH
cfjCGyxWApvWk3UHiHGPCeEVo97ijderkLEyQsOmhmalNKlhTmYD4ewMTBdIe3Mm
X9Cs/lTQ1zpbwnbPdWIr/OM1Y9dvMweag8dm0/eB7YlwIeaeYyhuz2msxjoaV2A+
YQjMS1pqF46kxM7+hgexTxzTRSfVcN/GSW2qezT+sS7bfp4jFEmmqSJsHLltLILq
+2xL7Eytu3scOy/0SAH+KGKlrLshmRbv1hyVuJiqI3hIlO75D1+widGf6T1+sheN
/CNjDSfPHrVlX05D5bMmus5+uVLHk5cs8EZEu9cQmAtoBc9PobNR1m3T0imMjYFt
18imQU0dXPjKa7XFCLCB7GxrRTW3D9JL8Oip89x4IedTKECrx3c2rqBaSQ25V/HW
VlpIhCCyIhIP3rppMURVXY9YrGqFlmOBoXgU6yd+JosoZy1P4j1MrHxdp+tJhgOh
QuE6iRj7eS2xqx7pGc8ZN/HiKqX0Ofn/6pitOOARwYzKawvRjfO7Bpg2zvtrMFiB
JbSfFQMOVaU//jH/qy94kFFCBsDIN3Z4KJO8WyYq91dsX6wn2CnCRxNRkRbNmJgg
EUBJMEwFYD+GJj3yEq/2xKLxkxgrLVVZG2e/eu1oMB+UUkKhvFXdmj533nQfG6ls
I8Q6sZXHycU6ZiMJVgmZiifvTt47MAn6hmV+NCRBB5He3fTaBSG/DcgZddsvb3MW
xT8hONw16OByYEUwQMdTjnSG3j/h8PhmPFqBFevIJDjzuU/DnC0K1qObtCeLlnB8
sqZtWGWvcJS6j7iWMXWT/OPJjwGU454ZwhrG0G9THUL3DZngBmGGlF5eeR8xYS5R
UAG0z7REe1PtIAAZbBSe7MDyJwFeiXAdqBNhnbapJzOqyDME2UgAy6K9Ie43LDPS
9orO0GbuAcuTvDbpupAGr3Rki7z+RRl5p8ZQD5pqmwifVAyDXY+hz8fJMcFgC0+D
9siLv7/kLkTZbSll+zyxbEt0UHyh3o7xfe4MOYX+FhTneSF3Tonaz65NBp8bawL+
QptdA6UKthnJKh/jVtM9Ugec+7JHM0L+uv9wsk/XKlDwketP2INd1o+fwOzmoMbI
c8VOqKJMeYM56GufhMYErYo1/CgYcUC8oXwQ9gxf4UP5tBIbO0UJFIG6dohRfVxE
TCUewoWODBnB7xzCT4oUsobeqlNcZvzmH4fr4psIEUdVD3+9JQ4lWiyImnQYQ+PF
2m1E9bn8DTEf6Xyv0nbbMjEp9dcHoAQ3ad5aSH2qmU5bepI0F29ufLB4zjX8vQpc
czw1vZVTUMsJO7tQl7MQFvFKur8EgaTtmIg9nOMB2BhbI5u5cMN+V7SGhLKgI4Q+
v/wOmK1PYzsgsGPZ4PVFUV0CgFvLA2TVSQRPrjGl5ARDvhS0Xivk9a64iz9am4Uv
LtHAtpu1dgZIndBACcLgDHYK/+XPkpmgdLBTo+hJVuGEQZbYEqJ/3ZTd8F9l/zAx
LQOkb1v+6H0rzCU7NUaQTkxZho7PpB5aPh5n4cbuojI+otXdwAVAv3R1W7xyxtGc
1gzrk2MJhTuX2bge5U5tJmvENRT6OD392lAcCxLUzH7mGD5OmwumyG0yyC1uVso8
XH6lYUvkrEr7ZWMGlTpBcE+YCUHktJb4zAM7EqXxcq/lC3742zZp/yI2qsEVtMW9
sGKjv4ebWnnsPETbW96mNwpsG8KJ9CSmD9BhnAbBrzSJ7XN3Q4gf9wo0wbWWLmL3
7fZi/SWTrh6UPWkjclLxJejCpDznitxMqyQdiLtlnOADP2kO57QkcO/++fjMIRUu
ndu9qE+iSY06+JvGlMDnOvjNyVuRhCkXCwcj9XtPzeNhi+HXRRsvBRWBZEKJ99CB
fLdwKrIdzHNrbmqDBv9AP9Ps0rCMyIInwzBXK93og+zcpzDolY6Vq3teJeOuFGlj
Js2T7EvyXSma0FQ8WVT1SUl68fyumOk3E+6W42rthLGj2UC0ma0cn43ytsK/bmG6
S+gERe94uAoafwX15pEroib+u1ZABCYy/xgEPl0Qr4av2ANiD/U8goa9OERzfvcv
7tKohLbxd5xOjJu+Vy4NwMYPxjC4Ox1+PDd5qe93YKCPFSZ2HbJMLDZX6Adx8WQD
R+pkt7qTWm6apM5riVWhKSY2DNvYHWGLjCntNarAXhSx7dypN7BM1HCWottW0X6k
QELwmc/DAnngqNtt6Tx8EFFhqMwKBD7yzC4LZviaOykU/crR3mIqZQW6/bK1cCe2
gvhYPTpmtUfgGlP/2eu17pHXqHsIjXXRF9F0anrfpcvg8lQjEO9as9o9UogovRVC
AtfI72YpKiZYGatd2l+KlxyymkMoRGNeXthj9XJk9mBZAx0H4zTLhAX/mdAByLBv
8x0hmQ4imZX3KlagttWJK64yAQ1eytNB6MYnKQh3xUIlj+o/nfXfKeGaLuOnfHDz
9FqcLZUg5GoznCIZFS8L00VnF0xd3sY2lp3gyn3wIRO3/NXv3x7hWscTNUEjZ3Pw
Cyd1U6A3P5DoBwEYW9FoG13ARM9/5S6/02eaU4X7bB86qKgqtUsvAi7tjC8ZKzAr
/CTm2laWSPbhKmewmifoBdwnOO83yu5RkbXo/ig3dZkDa0oPhKSb9HSH4KoffAqR
op2WyK4b6BwsIyfNIM8FUJKGGogCDfTa9OoOPHBvPEDAPiE5NdRFNimG3WPllFT9
FWofy5vzNyK897JI5Rgr/iIK6I/+jJNaZ6mNQcucuzgxfcSRSki3NaSrsQjwhvAt
vr1DYUEKMzKxEho1nYu8AQv/97exXEq4i1k/n9QorP0OmIILwZ9Hta0D2WXdXGd2
EOp059muUq5ujZrdK7jrtdlsm4d6s2dP+G/E8G0raKjTBGxG76HLwbp33O6godHW
hV3A8MVKIgASLfmETMe30QcehrL6YgLiSKt4X/iwPcUqUW+cR0LTacVs2HEROGiA
CZN5labreDKiZpEUs7/ucXyY661hI58pwW+2XH1YV4ve28jA8YhEf7RDlUHQRhZw
Bijj0bFg6wthEAB+rUMGsSL17wBKkDbGhxoCRihdsknggIpcFAgZKwZi0A6tD1Mi
yLBjdw7N2msXwB/uuYj+5pVkh0FYgwlV4EwX7x5CMY/vKkuHYCU11W2wmW2CTOBl
pxJ/2Uhf8vmQ9MHlSueYngLdDKXXDOuDR5Xueg9CWazO4CIq18ZX9SmoFsPXbm/W
VKs6TtbR3JNbCEVR6tFQoarLOirx9Ipb/JP3Ig42UJb3rEpidutgxIJMX/LBUv+q
HldAT2KQmcu3GHgnnIEpmXDre6fG/G5Z6ylLG11riWcLXGr710rI5tEaTfWEa06Q
R8MbH1uFl5pM6P5QAYsBd1VUrA8umL01/bEpmSIaPK7VK4mbb5ovCEzsF69z5qHD
hvjtmNxTqkLSd6JvVapQ1+2H6mLbZvEjQvtzBGK42YPz4lCXkw4QwgbPWIcjddWo
FH9GwDrIcTfgDCXQxoYP52jhZG5jQ7aQ0apmcBFYmxAHao2IAss6ruLkyxjtdnc2
9JIuKyeZZrAh3zvHnu7fToGo/Cs4YzFOORzSCJmUk2NKUf1Fhato6tPkucElzGgI
jByOS7kapc8JId9+GiTy6B2BJEk4iTONBu9YjMAh3YnVzF+rKI7C6zEIz6+227dh
34NwcztVEjZ9fehd8BLgpI944Zui3lM7CRnDfEpe+VM0CPsF+t6Lb81Zx994a4sj
5UWpvC1LuDsN2lj0Yb+ZRC1l6E68buaGodVlEBrKN2Z/GeFLDfEJGxruE5repRU0
6PggT5/ztNwOainpLhGYmUuSe1zZN20ysde7zEuB5iWcs2mDdVCTimvTig58n4Am
c3NpOXAr5kGzR4pEpY9I7GeZloORhV1JmbwUxCQHOeQ5EveNI6dqdx3PjFt8dLC8
J9H2Fl0sd2iRgQ3IpjKOVYXU/z7zmR/9fDnPzgsOL6VUfh8eZD5ux+o1pYwLfa6a
iCwBqdWT+HGj49H7NtCkUIvCnpNC+q+1FNrCRspxIutjwz6mGS0RkgRSMb3DcnzL
52vv/t1ue6s20t1e9hotP/GoqsUSD0NP1lSFXyESYlL4lMQY5VyamqSn+9ZskApg
OlQoo1JMT3WcnF4YE6ZdEMEUSJgEix6b8fBHVEvdWYrEa3GmGg3QrBRsKtRkD6/O
ipWgZQf1d6D4dADcvScSyT8N0ekRzjTAAG3AtqJq7qy0Jj6gdWpzR+RUdzJboki8
ZALuwvuxnqYbtDrBhzKp0HmwTDxSZI76Efx7H+3b27JN6deYK5XXy+Ps5e+IO0pW
wwxjy3khgtGYUDOj9A98kDkMc7QpJiSuRPhN0A48z4ksYjLT+qsl8VKeFUFLZRge
bvAPhWAcYGQXhnAUn57aUwP2Eg5M7Uda1l1VguWkdltuY5JiTiRz41dDRvQRnJ5z
iuDZ8I6AgcPhHSKpJEc37LevHGXV2cqqlewxBi8sIIH9oyIc/9EiQ1X7zqjSDcqj
m5CVP9SgJtBxewWv731Zbi5MvE90Fjt1uI6eCPFPldXElDfTlmYXiryiR0upTJCp
yzb0Asyu6h7ovtiGZUx0W3S6IllJ0U4PjRIbSXhdEm1Zwpm77lRHwgNLpZ7hXFU6
3OzspTrvFcLwD2QFcW8FuLWftjWycGO/G8NIAsTD29GpszSb81KtWR3pl1JOHd0p
id91WM0JWD+0cn0dW+aO96GhPtCocLZ4cURCCQTax4uCY93K2grXok8jK46KfoQx
DvcXeNyB13pn9pqGbb7hdIIlECaqCdQBNTdCwin1mEm21AndO+sOmanZBhRjsvJl
8gqV/DJkNYveTrWpUNZg9gnOUSBXRGanWH+Cbff24Tw7/5qJMfKlP54EQTxF0Hu3
IEuo0TyBRyE1K0rSqo6eZswbyYnGIIzhTrgBovkxqHplSZj+6yPTxDs2TEnl75rw
Av/i9R1FesOsDY7CBt6QNTrsLrBAHnwgXCRHUyyLFyiQLMTTbATzS0CAyC3UF9uQ
oizGlV1OntMb+UFQifntPwctEK5fIApe+vYnuJE9adIOPpMILk/bDi/LHcyEFqhg
R6ZcRvKJ/Y/LLxe96wdfYI9HVsxzDLfw66vbLoIH/MTTIovoFaIXGHI21tI+dsXr
YWVRo1CFl54BdjQ8mEu1n9DhB0IyZdNhyxxlpqWhsKOBw73w861FeHN6tAkTXlgn
zTnlt6oP5AxR3CzmsCfck3qKDMsW+4gE+Kk2HpbvmKXcu/DTlk6mlGvVK/KZT1tg
kRwNHhIPnuEyhTF2H+sO6asOQmhQ5j07yByF02zZBnDa8HMXKp7/c+CZ9vFOsn9D
ci6RFmXb3z4UnepY8Akt0zyOV+a1jao7y0j7tVv3EphmoDNflfIYgTFkWPwn+B32
3/Jm763eoP+35YZjEP65nXQQ0AjTzutx8JsKMyrCCbWfFFD3hLzdylnNegnxUCIy
/UZds7yiA1ss2fNJxQhgLvMtbsXBMqYhZAhW5QgbOsX/gKlhJD9u1wwNGnAI1MHf
h2C0fPSHlN0Td3FJcrua2q2p9OIIRb6+eU0bH6LmJ+r5Xf2OJUbjdl8xdnt4eRKL
Gckmm0JpOh8bxsrhAzozY3nBOyiwJ3pOtnN8ifiTa3hkoFlKq6s1USZsPxOBwLjw
ZHXhV7xGqgGAjHDsDMaijoZVeS5nlRwbIXEvx00hK0pRj5TFE7twPP5gRZfgyVva
A0INDfThGC0GuTMurvxYT5EgPPOFlrPoN4E9isdPMXjrBS4U9g2K59wg3tW0C6X+
v4fvlo5TrWTufFot2QC2ZtVXSb9LEYDfPmks03SsVXGfBTdFhk3xdQeLaQCDb5iY
hogp4MtbPYYjSgPA/bfQSf3rOEICWDRU7kPBYtFN4t43+GH0Ow0RbHYNZkMRSiT4
1crI7gE+BJqxIb6l+OQFTkdE7j5JLrBOWF10WpzjRXMjqQzWSiB+BSgsFJGD6FLs
8hcfFtSBdZSlAF6nU4KPG5YnrAymIt3hWFPlCFcXfA0pSJHKOwLJI+2kdPp6P12h
f/XptGR81E2RMra1yaQZHwBxBrhIF4x5GGK1IPkv0J0gaBexV00VYX7NZTPY6QKe
3NfevIBNp6HhuMmctRb6okN+H7rB96Se2SvjwNTbah+zd1qjfKU+DY+DCY73kptv
Ghm6We0R4F7ftDlwiYFyJy0HMY/eTO/gu3OxGbL+HW/Odl5klccVWvYu5xBlXuoE
m3Xbm1cWfXN/CcGCVvF049rIk9v5I68XQcjo+oN4L0ogG0tMTz/xAhzdeMYVrMab
QEY+LHcyVxEIxLbtDa0AhDKEYk8WPzfoIfU6ZR6K2RYgBWofVKsSn1EyvQgZEJ0f
L7BK2YuVtqi9vcJ21n/OAMzOi3rZ89qz+VnclPkbRC/Lfzy4vO4FdVqU+GMvcXoI
gCJXRjUwL4fNr6Cb9sQmqPVLvjJVB8h6rMpTBsPK+kBgNRH8esFgQqR0+z7T8JA2
YTIkIAfffoTj4jc5UxvJlxycvJsTVsyzdsBJsTM1sIEP+tIQa5l5tW8jrBROWrPO
65vLkdxqvjob+IsE5HgOyafePATJ9W++DryGf8YEMI2jS8aGTPBu9eoCW62QAal1
5iiHZm4o4w5yCvtEbJoDhOu1ZqaitC5gPyt2q5+1SrLQXHh1JK6eAdZLGO+hGNf2
91VQQNqr04HxeK5YQR/f++R26+4QSIOaQrqPnJgoRLBo+uYPtwzoFIm+qEE8H+27
6NNRqiejjPsjjT/mxpSQTpsojygudDOQWS+CwVG3FKYWLulNjgFtP7E7bhZLWyRt
78ztuQlgOvYh/0D9BGdCEPT4Z14jA2UaSzGtqmwMyD5OIFWiIyIf08Zb1Ys+GehA
Kvdy95omYELyBR6GIC7D5unjgLsjzH6PKEsBD2Lp1ekBVBceKJMrj7P/FyRfS2Lk
lfUdhDx06+zBlcLVJBQdhfajayAs9WsJVc0RZ8EAaea8MANymxiCEqUIpgLvnkFo
d1SbEOlPWxXFMYpog45KPMl2QVjpuLukLkpV66c54hZBXX3KaumwSX4JqT96NCQ5
CAGSU7frRUVohng5OpK87gyGtlqHojow/ye5XAzQ62zu2j9ESRXGgoEkR+TpYiYR
rWjSq1TVtT9LtPQc+n+XtGwueXLEqB3oYVyt8GLLnygTrHe3fdgdcr2ma8cxWYQg
4ko+MRymEiRxzft7zboNFks+2KnEwp9xMmsLWytNYACAmhetT2vnFtpevkWdJU9z
JPJWJIzQbd4yuu2Iv3BgWUbpP+Hd08d8tEaO938K23eMltOj02ZcRZTNQKA0vwjx
MX+kBxX7oBzjkZazSTYa5wc2uz8MwjD+dBElsB0VTW5nvnE/DsWTbMtSPBvr6q0i
sGJhr9hGvzi9jr80QqFH2X1HMD8Rt9UXBCHLBnM5TmzqBR90TZ0n2WstqQ/1PUpG
oaXPYWrOnNeof58fMu6d3BPxgk1ZARf4aKpFjCDagmyPVZp/BKIH4+P1OFKaiAYR
DgyLY1ieyEg93xnM2qsE4ClZbvShDIGFqvjWOdSLvwL00htktvdFAIiA3zC6D36n
JTIWveiE8OiAEzVGLHLariyCMgggG9ud4Fm/ig408CJhDGG8FAtNWUL2QmwIeE0t
YyzVuHkE+XcPaEFiQLTW5JKc0OaZWb0Zp8S5BkxYBTNe5JMfmVxiriAxuL6m8y/h
L/vuFYKhVK8qh+WpD/B1TyIL2S7xrnNmnxhu4oz/tQA5pwc8hUAzeK6+RZh3dYxH
mxKkTx00CRfPOPd+peIMWlqagLQR8SPR4ebE0p8eWZ184tF+t0SUZYVHVjo+npgJ
KeoWhzEiddGgHwDikrLpNlELRb/vu3sfcD7AL0N3se8Q8dpH9wTHgPP7XDLhi3J5
0kibrMoj6if5W8GOiR8KxPixNVFozHqHsNmQDq1TZ5PQ7361gvsHihXg+vniFqZr
ciUyVpnQrycD/lbJbmqmCESzQBvH0TO/GOC2EBQBaxq42NahNNFPPv81KwR7u0Ww
X4Ny1bTmJNNJpqoceOK3g6PpJCW4IbjmcBYeqPEauxJCun1tDE9Xe85xQQOfOLKP
ac3bYUnpsmnDvzvjFto9eFfufNbaNw3biWc+Os6NgehozDBgrM4r4pJcTjDL7df8
jB5OOjZ99iRxMzhr48s/mHgj8mOXMbR+5LpSzV7re+o5NWrZRlSgEBtkk6mM9d7g
42+hSjXxssLh6+Opjdb3mbJ5Xt8ccjUi5wPBXcazyuABgANubaM9S1TRo45KRC+B
z1RE8+wMDXTnWZmptFYzEhDzYHsUsIGQ2MSTmU+bjzvRGe+6tyD7ImZH1v5ys/W6
b+iiTm6zFGP3nsVBbm4kFY3/OU2Tpha91cUdxYb9Ndf9nYd6xK34LJ3vUQ/aGtJe
YRmT+dRISB5ogaXBF1rshNqLJCXfu6h6xaGjJAJ+3yBSl+AatLuHpb0gTGnYsZiu
RKELWX2BJj0f1o2X4h8Cw00cGan8JvMYRtaf5AvMdf9OHz+B/AmOx5Z7+Oz1eIr5
BdZ2N09Uon4oNTF8Ov0HxFINgO4zd2rnuzqq9zu2AiAHGkdniN23E5M9MUIxgNds
gIqT3tWSXWwDSmf7iB4B02L7TVuU8UHMgqmWIJita7Zqh1Z3XsRJjXi88Tx70OIZ
U0PvR4Gpw4ERlYd05odlWVdPf/YppOxXmJTVkvZvaIp1/dJBX6Gcsvt6P39KqXS9
E5SRwXFqTZePnGDmHSGMlhzkDOD8OzrbicNmKHqRLmiNYqA35U+EFG4Yo3E4gBqZ
zW8BHxLV9ecV6pk/o6iUV2ZQ2cMi7aIIEMf7IiB0+Dmf98Kw0J2R9LRdd+x1nzwD
SHr0kZ87d6f0IQrxUfnWq9eQg5S7011DVWyyxeN9sYbx+9gLTbBaMF4EbHSSia2P
icDayKRbRSKtgz37znFLQzHSt6l8SjN/nDCib1vO2oAZyVrO4YO0KRdrH/uVOpS2
+IyIa71cXgx2dJ+0k9orLbAKYOXIiR8bpoFEefiwMoXZ2NJ28cZRe88ff3sF4HGq
veuW757b/6375Uk3iYeq7/y7XYR3OcOsx993pizhitcHjojWT1plD1+5CIUUSAEU
T02gfZ0xWSYtwj+Yw8huIKToOaK4gRJTABTd+Ovz1YgwbkmW66vqJ6mlOXFmcTAT
VV2SkJED9iVo82LEGXnYMk/s7+4H/Ti8kMwGXpLFuVGOgXkXxr+jknPm0aUWp6UU
61bigo64BSnhQ9RuEKmsrwsHCux6l6iH/mjKxKvtzwKJd3Ktghx2Rzyz81NmnmoC
sJGADT7Z4XzuiKwGv2AO+PiZPwnF4/zwZsw3xGOFMkEA5ItKcVHyJV5REnPXEwcn
iHnihYIB/o7ssA6KVJWOxTZwZ82gEDm5DFvnu7aRbZK5ZLXtZqrtru9v6ZuSno3g
E12JGLObcuZl8ww0LFgZsz0sPF71ISrFU9ZF1jLRk96GAxobGTF70VAc0fOxPo9l
Itl81UJX6a/9j2dvjJbjYHuS4vOFuoBCfUFISVdzNGFfJPXnhYmkLK9j06Y1CzWa
C3OsR07HBgNbbNViH8SfF3vgKcA/2KJTbP5e/lkAAuKFqI/SzZqBlp5BeePnHMXY
RQWyyDQgBbMwHhWgAEqB+tg6tzyLNe8lq11H/1DpOEBS9wlkUl5Y4/AoTAQybtOG
BET1CgTjSTduAODw4s4qCuV6kXV3stvNod7IO9yfjMavHyoOaphOo/e3ZK/8Jpa5
c89MZp9PamG01IM/JWYpCpYONf+2tSmmRMJSDUcTZFyXWz0ukY8G81knTD8SSnBn
dDnSYAk1JwzWU+s8nvXA0420/BUb2u4zhEhIu18KoUPOa/fTmkV6Jl6vtR9iDEiU
ROXB2IObDCcisy4+K5ji/mqlMVlm2u2CrNJR2iTPJCKBtEblfjEVOzaIizmXli8z
5GsinL5BHgp12yiC06fmGO2QLUzewtO564+uysJAHwpQfzrT9xPGvzgE09yNXTyd
hB8OL+KgAuc06894bYLiUQ9Cc7k3EdGkqSWobMP8dolvo/Q9/IQoYTtW4ZQZUwtD
DuRmbmnFInGr5cOznzy5b0sR2g6fs8wWYXi/KQgOFeIQeXuj3BXqV2HtsXHWCAKG
y3fDLghQ/LL1xiYOtX+o6FlRWjtrxAeu5fD+GGIfYYfj2IyIs6d4xmxh/nRQzABx
CwRdfES1AYJ6PkpZ5vfDg+W2UWl8/rjGAQT38Ic1qe2bZ91cO3sPKX7wJd3itPZJ
Bn3Wa9RXuwHpWZzlRbO4aMep1Zb+nP44WsMpObv+IaJhSftdw6iI6az4m/uP/56j
YuRiAKtk4yKjIMVH8mElctH1PNwZgNKkJy5q2cy3UJPHqnX7KhynDIc+t1KSrbDQ
SGIEExf6vyva2qBTcMpyLnasaux68FdZB1aT4y0kfY/S3KT3SV4zQZR1wit2h0l2
Eb465+xVpU+zpPDgbSPkVPXNuG6I5cUkktFLM2/WMIf//xKBQP1grJgwEDJY/ajn
6Ir0aEhOR7FZlCj6je9l2XG7HE/u5QK/OTUdfQm/QC3A8BUkByWMWrdqhUsqZyPf
8Quh0eZNVX7n6vDaAb2M2LooU+DwiwoSLq+71Ber5S3lGcwJ3vUuiNKA4II8HVF4
rj/1v8dJx9x2xbZpne0j+GBWVSW0JEqzPWhLdZHyJ95D/iufm7JEL37w699Y1lw2
Y+epgZYAvfPmmUKAy0KdbJ19uDj8d/CbVng5uwLZK/XdfRxl/omnoy4tBkZyRxtw
wUaCjtUhqRgc45Tr+GvSDZ+I8GdyJeGoWxeD5IBwRG5QnkZN71JfFD74LCDxaLn4
QdaRgcm2V+ScCnBmBmSnjGw35BazBPREjub5eRDWjXHN5JkLvo3NR10wGs5EGLcF
+qrlDZ47FtHaNmM0AoZkyUgKkiSPExhGmstQwkFw7F98Q572Czg2b6OHkaCZDwbj
CfiK7He1YQVyEvZRRhKcqO+Y/n4mdzDQn6BJ7m61mnz7ejvPosNX2gA0VPHSrvDR
DnNnGMZgL9fTjKvXNoZeQPn0RVB5KK2Eird94jYKb4Lj5co//R4Cm/Pnro49ruBX
m7NblbQsxUCdKJfts6uo44OSIu4Bm8UykXxEQFYRDrx6iiEN9RGH0zfz1r1SYLwy
5oCNYlvmcza1U/RaZnQhYCGqssnV3jhNKlZpd+6p/DcS1XH74nZ2ifT0kW7kJZS7
qI4SRRaFgIA11tDLHOx5q5KDk3yKZPI3ah8T2QBwz5Td2UL3pvxa3HMDZTUGgciD
id5VZu02Z4/WBR3i0gTluFxJoBdH0yR2fSaXV2cJzRAIkDJVCcyKMWrLU/ze6hiD
mCRHGP8OwxFbGzx3oqPXfFZ3geKgvr2jZjDr5Wqep7pwVPDnVtNrzNW+y4/AwGZD
TJQGfqjFDD02v2UU7N2Lxyt2ozFDIwTmbFBg17o/Z8I0gYDNGlse2oeGBpZ4u+dS
lluqbrivsbN7vc1J1xsqjpwXc4USkBfaz1rcxqpQ5/xUSG/KPDMueCIGoqp82xoc
DScLG8vNEyUZ+kUGKHoolnevin2xEpBCv8EC6dCfaNhtwyciL2+rOCYRqdefEf6D
j32sWVK9lE0VCNn1BzMM3/olGAz0WgimyN58XKJCdGXBnas+zHZDMZ0tYtqWqtg9
j0qUZ2McYBElKfD6C8kCOIvLG8w3aZBz/UT5x0AOcTpy3iAQS7POGFfRFbjahA0c
G80bNQzIRUeXnXHFv9k6NX1YQlHfTIrK5ppvtA2VCnZMXMeUY82SrWDijfahBSDl
8QKydxP0hHjJILEMtho2CL8FOH5nlYLRk5A4O62ahv1Ed9k3kD5iwJo9zNlYu3O6
IKOvGtVIQ9UgGhOj/V67A8Ej9DUYMw9h//TM0WGJKEWhhcRG5/aQi3KpISe4gysX
J1rJjRochvq1+HpZWn7crHM6pgNstp9QL+H8mrqST/0PWj47+RO6kgmT1icUBSty
YNwunyg56TYdaDbNAL22QnPkDECVc5lW1u6bMiKqKw/mlAh5BTTwZG1uHzGhCYW6
tVvj5emhUE4+iFbrlmk3Tvuty28FyGYGsY7AUZPZ+JuOJIrF59XAUZPgd9mckcAv
ttc0rgiVMVmwuIpLaUXcgtbX63qQBXbD/Puyj27i54gof6zPY/7aJH/3IqsoL7zu
rdPwLyFq1wj1i5cEw0YwNlzZGNPbwjO2+9+zVj/WgnMi+/SKd/hrLDRN2c4+fa7D
GzrJGmi/FfrAkcDIcZei+zNVEg3NA2wQkLA//3S0jPEgv2aRgU06oXebA5MiGN/j
6/c0DAP5eV0wL1Dquz0nf+22qRBWLvc1rH21GHRPjG23F0+7Xz6xXDltxcz/r7Dl
LwO3ANj025I3oH+PFH9tAdEDIQ4FQL+MKIw42MOasKLBocMbSqVRbeqBjy4le8rr
IqSoBSkwP0HUyOTsxAZ9CZsoWnuuKSEsQgl8KoN7dhhW9SuQKK6RypCER82w2MQ5
WO5SODiHQ2PeEh6WdVDzsbnljVP9WF5b6lFBD48leIQpDpyV+UjNKDhomuGV0ucI
iYpKbq4GzHq/oygRLf1Kks7NlFSfF8H+e6tLhUIaoPyX9UZ4Wh3CmsJJHpRRizSL
vvtasD1zYnhXTWs4Z72oec2POkDL9n4z4SRnquwSjCbYowooCk/stxM1b0m18zhW
tNb+lv2nyJ5KgVlaVtBIrWHFod3CVbKtJ0fJ/Mqwy+8I98H9HcrNyze63tDGi9gi
1tXJXFFufAlBsWyx9MYEVAQ7+IsejJEF9xDr9wzR5WLl9L8NaM6qWtnyYh3WrsDW
c9zhMZz1Twdi9zgGEEuEuLyv8iqUMBNE1UGKcfJT/EZQ0eIM8nc4OqAAFsthsUMm
FMFaUCmNLmjX+I+jrlI+pK1hEJGYzFxHfiO50mzqawtGZ/uRv/Ur0Km+dqPWEwG1
gxtKV1LGKoedAtkrL0z2C5KOqhH3DBg68l/UnUMBohrDhS1k9QYgR2dZ01BhFKMq
ocQ1eCxUH4gT00DrffQR7FIPYQAfLDpy0BZaFxr0+bYx1JEzPFRxZ5Y89/+0mqjP
dp/0ngOeexaujbn9h1qNBE0nPGy6EuTgTh6OX21xivdEAkRJ67Egs2VKTDHgGdIp
acYLLRrARGz60GjLBkoSqkTJ1N7pHOCGZDYnaz4XX+yV7SeqA5yRAAU6Knn1ixSZ
cQaXVMIeovFeIU9xswYcx49deD7PEOz89jDt+PLwDixpkmbn4z2Ha2A/nI1sJcGf
BNBxQJAIj+fqkEdmegMLmW/ocVJjS3StY7hYWuBQePWqVMtPoQKrtVeZG8X9qGzS
6Ru7FdR77E+xMPbN0GB1OukQAEbGhHLrQmoiQLfSQ/RlDRMFuOIt1ahx+w4yDkpp
Kp+TKUvdVNg1ipr4jCplhRFd+mlj6wK/cygJFrWREXMFde/U/r5ISMdfsau4gxPW
TC5fx1ZhkId6k5tr0CS8qsKol0ASSCyIp20Fl5YoNqLdHBUCo3kSTZ+dSokvYfJJ
P2k6+TcvR8i3VkiZX/PvIUjgVxyjJrgXgNAUYqg6dBWrJr087ibpGRnrWD7na8nh
sSImKlCv7Cb0hm+ai0MfDjAzP/grFXzpxKR/wfIj7zhCd0j1T6MH6yyMTNSxKHbo
EzowRdUIJ0Ry8SYG9FfnoNQpc8XzToDpw7PWV3i2kFxvI1XP0AyrNmbEU4TZPLKa
IG+/wUvXoneIb2/TxqoPawkEQWIRCTprD9yfjg05uaauRP1JFe0PvaqQySIN5xv6
Q+a1Ydp5h/NeaC2bUG9waB9Z67gSIdVIHhXTx8ClA9OiHvcykhzuFT3onVq3esAT
tu29SZohNzKdCBQX7MMfNollhTLay4LngA7GLG2ploRaS0sklnz9IedEHbwznf3C
cBlUfhYcPT87CNuhnxz0UhM+RkZWHZyqxJnvzIUJj02ynF/ydeXoUTOl5f6/QQ8N
m/5q8b5s/O0Qf5m+yUTmxkWd4zdpg5hjV3GB3I4l8D1Bzyb0BlxkCvk4+Q9m2Y9r
wONv8D5msBInC+jMgMLMFsdgyU6la0vHdViamFmvXn+nWjVPWXQJ0IlYqKzHlsWn
dWoIMtinI2s6h1xbUceXAEerB2NLKcr+lmISOmHhqsm3qsNEKO+dwnpbiFR8wGMQ
t7QSrL/ZXBn2uNkQxZo2hlR+DLdt2QbY48S34iogKwMYcEz8b5GE2ZVNJq0uQXcZ
TfQwA+5JGvpM40kQwV0UYhwIQrZOwjUYQG7JaNRQ/eBI6z0omYIRyK4jPbPF+JKj
QJvuYAWG5H/Q6U59JYTBJwFk1cyKu73R3kcOoKyZ6llWIFmKsFJif4ZJnFNZsJt3
AqPyvXHfWtm03yvFaDtNswUw0jAFfVjKyIaDS3ZVX91oRbCdAWePbWxhK3OkLsjE
AL3BzJPiUBcfLZbyRdJpnKzQNR3rF8gZgwXK2iAeIpn/BWzwdkqykobiEsKbDX3Q
rcP9CeQ/Mn/X/3RlioKeGRFVlkY3enkXEXGRbqueZruTS7cio6AiLHSdtz0T5Wru
ZNXoiydHCN+J9eiuWSpBaPxsSr1dkTyj6VXaqHp7qnOaNDS4KY+uF0PL1S3Xcjec
g6LQ66hTbxO7nCiEOws0krZVTyvrw5z3jM0PxCF0pb4OvFTlJu88SmKpLKZGz0d9
W+s2W/QmqTIp3M1DnWrdCLNaqdM4iXXkuIK9RtSpSTJzvB4wx045W3hwV0YXRwtO
xco6vLB4aXMGOPjvYEKyvpSeB0Z5qWTQK8dSxztMmvrU0kLiiVSuQRT/Tbjuo17L
ATjgUWnWdEEti7ifcLpTzwM1wJ3ry9Y5PErmOP6LPWavdSsmf1qkh84Skjh8rvp8
9KM/ifSKa4RIRy2L4pWAksAFpDrUVqxIh+FIBKD1+97vTrDoIE2V8ADWxdvu7UBc
rVd7qHU2WT8AfigDUGMd27HgDuBxv4rOsBM3oV6NnSfL91X8hY208QZYOFs2tp65
hf7u5buAbAQFi+dzExtFJbslV6e1MpVmEFhBEUeIsxusxJKHIsnr5KUy/tU83IdO
awoqSRnkMJm5OF8s/kqRUlt8bUPLlRkFSdrPko2ISm/EAjm3DvG+LY/cfeb6ARKN
ZzZGreh/o3O9RPfLqPy6XDSI/gcGFpK9mVBeqXO9CC4XQNmQ9D3GbDZwRrWUcDm9
ew4WujjfPlRxi1eOLlYxG0YZmR4ERDTcSodOHQptlletergZVk7s0fG2JQMCop+m
6N5qa99ts+V2ZWu6yrDdv69GjiIUthQuYeIcwZIb4/c3hMmocy6BD7HyOcKfH97c
8ONF9tepCQZAYBoaF1Crhcf8lUVsOwNyaR1bWoxPnVRjCMZR3UhqjlW9RGRnrr9x
0XgW9QVCfAXXzmKVNj70G2erEMXggcu6RgsE21gfMS9XsmQwhKJ/R/xxmSHPMtZx
zOpuP7fGEhRd0T4ta7q3hT4V7dRTL+u9RMZMxOvb9SERQL5t8y7TyK78dR4vfAm3
Ku6oFkFT2WW7dzJ7nuck0JuVHTVaorIwZCWfx57cJpMgBAHOmj1jAiZ9ZtSn6VF2
EgmYXHE/kcJvnIyNcZKKjKJzMenyZBE0sysSxry4WQKM3Uzv1JSzTikbpEZo/Pak
lg8TD9AhENKYMvZmV8ds3fhTaGgXiOcbp8bzGVBXmjPYa9e0QN6nTOgSz0LVO0xO
ehfxkN3RisEOqSLZ0eVWQno25X4IDVPZXwIiWOkIjnqjdAQAxOHHG20aUS7uupN2
dAbGbiu1FfL/lLaijCAqTw6BbE/qUyxF/A0ol84VdQx+PMObwdplLVLMPbZ9mQ1p
ZPjGbKvzvOx2F3FyFkkYMvyivy3P9PiisTZBtcv5xw3i4HAsNfMVzz1NjRYckwDr
J2GUXNsCVyg6lJSJZkrPF00N0kqfegHssSl0MmlC2+zQNYn0QHusNVCXnrHzZLHn
W5d/3TKV9ux18uRSjq+OnYt7wjyMyyWFczmhifbudpke+zsc4AsCDzsltkf/ZLcq
/2f9yOit1qz+320ZBZzYyKI6lCSAMlvM9b7+2e9sRVnL+Y1qp1hDKUvMoQvh9MFp
sJtMXQ3y5JoBuX5FSc6qo290mz6AdpC5O2Tc2tQxNyt8oYBijvKpwa9/XrCrydNc
+6d3OTkEdKU2s750NhtqPOOMnaK93TR2ekSNeGbv6lpjyGFagmCPeWSCZL2ARZzU
tKdDBJoa6ZDKYzfXFIa1NBaA0LNCihh1N4qHruPi/QGLe5LorODF9z1uQxYYES7g
sOWKKeMUyxgpuvcwSMSea5+VnM0X1QoHonUjMRfNwY5Cu5SvllDj/EIkXm4JocHP
1notI5Q9Eu0NdQIA21cv8YKaU6aY1at6kRH7VCF2W08INLH4+ZmBNB2f+gjFQ8IA
edZC0sn4T/sivKYajQ25hhUykMrHyzhxzDzrbWzBjyHIfGib38OQy+lrRMttFTrG
vbx3edsCvzoXyX9Eyz5iLwPvwwUHECE6kBnncdi0YZJV4bFj0jgrw48SOy42zE4P
cAsv7vv573va0njPjqLRETr9oBQV/HM0h0jasBeBFQINaSN3aorCxvAfxqz3Hs7q
5rbVPeKv4EpbI2vweYdwx4mIjHHXRyEnNRmzPdLOh+E/JuWWe1ludkPsJWSqfG1n
8U2BQz9VnrQWB7Gym1OZiDKtVHXRVYqhavW1fZBLpKTJdSqpZHjAFeXbAZrj1oJa
MnXqv2HawbxbyXXMNzA9IDF46URfqWS/lx43TRV0UxsGjNKWcykjwdTRtU+V5wog
LtakrtvuA82OAW2B/0xZFU9czfPQ16qk66/i1ZzRI3Nf+3mKFsh0T01Gd7WlUZn9
fZEBNq8HqApQjZ3SoYHg2LVXaMZcOy3jhXfAsioI+b/4Kbssic3tYGMDT9f5yZ29
06dpbn7baRPxV9HVqkZLY/LLPHoEA8KcvGZ4YnYDnYXlZvkarqsNs1A2n2iH2VlZ
WkGyWQNBiua+y9moPWDyMEDJJvKh9LkvNjyoGJ2Nf/RHQJ/KcTZMwKi+6s2kzU/R
em9nCjJkx+BuqFO3QW86UhE+r9fbp8f39TPHj/8/10ngsAMVLLSuISSgZT87ZQAl
5X33Obg30pYqNcp1a51/wssGx3xKWOloeOvK6EHxTSLDyUSA3tb/XRXaXcXlOqQl
gj7Kj1f1ninzLRkC+ve7S8YZaR4BxrReQNQvCriNx4mr67oYthm2TLU1aSAZH4GK
Qd6mm+aUyKm5903YAcjF5CvtMc3Wicea9R+wXmH60G3tO+nMcV6qabHcqBGxAwR2
jceDt4+XX63CASMu2px3Rc6o7xqWMmu56QxJFpTpIatUMdRWbeVE69ypG7phVV79
sEbgp9+WAf+FcbqZ2XRZzyTrPPvNJLqihuCRzhUmIox1IJPB7Q+Lu9zoZVQkTXov
2FlINqoTlar7e9a89mD2aPTsI352Q5sfJI2ZOzKEfZRo3U19DqMmiNr7bH59+Jrq
RLPqcwo437VrhgBi+CDepbOhhuwTdvkdPrQ9BCCtj81KyMFTdSLZ7105tCdb7QyP
aC1ETOYFOvoW+6Jdr7gziDuwVDNJN6y92DweffUrl4uPMdTw3R2yeWrSzaNjJxiF
rGuKLepUpLQfODt+azWEzBP1iiRzz+HcGiBIMtwLN9/qM7niMQiUZEQ3nmupiPTe
ix8HLz2ktjYN3FfixHE7XtGfG7OIm+jalTggWL5HJdJmcRePLf3lRf3fpqle+ATV
HdL7MDpxdEtppNNheQhtJOZYh1STqT0zPLw17AuecGfC8Fc7yayO2ei3FZ+kDrT0
IlRXFhT2GAgyS3m5TsEFb6Wvgf2b2+qN5Lp4s5TZkb53VPrqQ8WLAymrawik+HGF
XAC+eqDLlv23BiUw6pgv2twrnExBqRJzahn7T5iLUuUd7Hw7ZOsdFfifPLjeC5OP
EXx+T7rQ5iMNhXdi59VWHtszfvoFYd54VQfYB1xJym4RX3hOk20jliC2bZTF3ZBq
N3536p2LISb6LcV3ZyqQNNp9pj+xMUl7VukSzqF76PTH9Ob1x+RKOslzAKv3osEZ
XVtopY+RgHShNsdqqmIyow02Uf/9ZoL6GDSQM+ekMadnMBLFH/DIY66W1TIQW1U5
EwhyiU0HELrZy2by/4UoTBR8tUSbwbaerYCQu5MEPtHC4C60/gjOt2dVHah/joYw
xP+TjmZ1oPQTPzdIjS8z5L4ql8b3Ro+ysRqNUbZtQd9BK7KhfXr2aicwZKP+Tgue
QbMbSe3RoKvuH8BQVnBXMRtMqAl1oh3e2R9dzj3Rg9uplSnbBCaKzIMSGnlF1twe
2DsQ0avdJgCggEIwFFcHr1MtoFY7f8BiqvSV8N7S4qiA9GxC4v81hbX/uSc0AQ06
pAScJXp09yYatQ2lPkXg7JZXvnTdSUUfaxYaQi089u6UecKjxmrafpNUVubNxPoT
ENO+lcLx1bqx7mYl+JHBopHpf745ylsnjc7Wef+eHnlWgtQa601O1TYnkQJP6mvL
W9Vt8R0PfAgueseTx5I539nfKalYZlKPEVfSGthrkF+CCdEwtC0urfvNZUOvLA/u
8glBp2I+pGmIzdCz31r4wBS1s2EdLcmBkAOFzMpgIuwy5IpfOvrJ0LfHGq4NID1g
j61Bha8BU+Uh+E2kKOPkMRd9u8WTytEP062P3kmHbDFOUc2CFepF/Q8V9Lrw6bBK
lTWJAWIeHON8uqSR9pJRmaQdxHA1A3CKuO5i9tISu5DLrdpTjU7SBdBCNHe9z19W
ddqnDG/J1fa0rt36K9ECXjHk6q/zNfHeJWUF+ns3iRyltrtcp+uh96tMtjcPclrY
PdZfp46jZVc7y/UM5QNznOiK+vmjVERGJ8V/4bukxXrZ87ZwicnDk3ZHCDGYNR7+
q/7a2Kukf+d1StxUgm9RPIRx12Ck821PWap0PcOb9viDrCXTJo2xjeFyUay+HLdJ
PJy8EE6P6Mkk6KjZ1ONfUuAtO7CU8vIRGSUW0yJX1qW79XcXNOISNbU+q4B0/uvF
795dDSohHpXwBPxvFtREAUFhHiD3ivK+KJ6bzh+quPOW6o6W6j/vRzZFge8VkxCa
jTNUKFavBkPBR52sEDkmVNWbmubcN9DBN37Uwa90XzajB33ti6jE8K4KwBG5pHbk
V2pDXhygiYbilnu6CvOQvd8jvu51plZCuA2PYcX3OgkIOw9bkiEB4CdHQE1Jh8kb
e/R+zA4NK3Rwf5ZEXA9DDT8o+InSGsv4BA9G04CXWuse4vQtZyTeFDwq8jVTaZS3
RLVvTorh9m9cktbt/+lmZ+zisfe9qOpr2b0BJIzbkhowiWzntiijdjRekgCBsGEc
VEnYOSle6HZoivCkSYEFRyqZdHQ152IPOfDnImGy7bNAA992dzjWByOx0KY0uIgJ
AbwO2hzgkAzHJEXzreng5urmbMbW7GN2Fvctivx+R5OKjSGkN4lfxULwc+HMGZ+M
biMGB53fQ927C7BsK6fshlCmL9KJeV1ud9+T6P3hK9rFjRA4QYKWtW66Q4BzwPBR
rV856P+juFFhdrjSFWsSP5md2Ud2UTEDvkmfLrnniMCmtKw6Ny4fNcZat0jGNCwd
iGAHCibDY9+zTDcDDojfX1bkfoH4NN/wbYIxW5WubE4kqNKR0J0MD3dvVB9r6/DO
xpqr4m/tXAr3TWv6bBuJw6j7pBY38dJFPj6B+N0uEPC+ma4iROcAf6Uh9hWc5XAJ
1HdbdOURxP4U3YbOZDqztHQgtebGel1c0wZNQF9QSb8ZOw0wJmDbz3IP0kd83QuY
JMyOjGY4WoYbJRp9aGBgLnKqAYTPhIjtDR9XJR30Dek9R/BzMWcN0H6MssofSdBL
SC7FAY8qsGVgcEO/1IMXyh70UWstm3CgGr7ozNssaecoVQHYPbyP3GLqSWj6IYZq
sNkNO/9a68tK9nc4ePWCwz20m7HNOZTha6miGifzZvTgAPDsPOZFYqnQ2RehyGSl
urPejCzsVP08nOjvygiouYQiXI7/9O3Luf0lsG6si1PJkbKe0aD13lelf7X95tWd
9rH60KdgjM5PY1hCHWnEu8+P0FiQii3uoUPyv9XcvPgm+qL+l5k8DjInXhPjBdCp
jtEHKmDr8/4xfoiEAJPIXd3URgE/wmoV345kTLIC5dOEpVW3TmxcWvZelYBZrriC
vyB+eRYhf7X+13lJQ2VZFWuKbVqL+Wjto3dZo6HmhdG/ICq3w8fjeTOBCcM4jq+F
jhi5/0IxtpKfgtDpkpH0rQPfYKY06X9t49HeWzpboRjHNXfNqggKzCj1S2tUUTxU
Zj3mZ9jONdyPx0O2WQJR2smEOoUGmr8ePYh7PcojamVzPt9mZcN8sDIEsOZHU2EM
7bYloj5YbNk1iQRs9eL3gUR+9Yw+TG+UbEKiCTlxMAho6L04IOBh7LKI9aEsC6Ds
E4JnqsLUDhRz88Ixrn6jJeIfrT4RQKQQdQCv5DmkvyKBFuEKeaUFsQLQ9xNq6MZY
yAocsOFzhDaqpdyLXgz4qpaMEV+wbNHNg9W5y+nz1gDRg2QA97q/hSgJcn3ocThZ
M9hepBGZO/jobWdmGRLuiQlN8EIh99HEh3dAUg2U22gB1A97Nxnha1RAtNQ6nenD
7zxE2TN2NyHGQJo+BaS66f9+2ZTfLwTIJM1EH9lskZAaxLMb8nxTtquBhD3TIPFS
Rn8lGpJhcINOTTXemlxowMkt7LzM/iK7SZYqPznUND53NP56mwgrgfBGdAOxZHRf
hmTxKNh/6vApQHmuomkQAUgPlRHp5buds8AfPWGhk0k5rQUILNIFd7DcqKy9FST/
WgRSVerSdqHvUYYjDsMU/6LIXgdohRgooKLcU08zNU1akXewAewL6ZyZF6JfwWSf
ccY6+jA2ZmofcDkQDsp5POgT+dXJ43mkKIIANhAvGrRX4abZ/QyQP10yCxtb3q1z
91blronRSvcDRx7uluEQOhXSTH1F8rlAiVrJpBO6BSn+B3qrc+KdEiPajh1ueZAT
oMSsN3tjiP27WNMof10xYfTLtZbK/rPfTpj2S9/R8c5BzwT3/HPc87/huG4JvVqD
63wR6ehc0skFZbf0Ysv0/nG8aRR+xqxB/6sIsCUgfa8m486dmrFY55oFoqy9+xP2
Kt3Uup6YPja7JgZt879Sqbkdi4XVIBXwT9jgvIYiUPNXHDGKy58b9Nhn/ZyubQJG
tWZxuMhq9YiwSOhMssBaTyYuGIq4g9AgxG1cUaLtJOb770RyIKzxebl4yPFp0DG5
x5lakwuLsr0fHSvJoS3/286gZL9q8xm1bk8oMZxdrzJc5BjaOLOBMSk5MHxMMcIh
LizjFO7eqsjYaQLOOdBJkOTj5U60qC633HJyePzpVR3sdZGaMK2b+v7VXSJfANT0
CG1Cmjfs5/X9ddv/Flp/QLD/6YJcuOG4X0f7sAHY0yKo1sBd6DPDjoWBGIi1qxnC
dTNVvpaoiTVgspu8EctXM96xgGRKEsg8xtyyIAbsbaSkqyhhAXTOVzsIijeCuXu+
fp2b2rYjXPWmD3LLmz+4rD3LqZhwjYQ3jEsZnYC193UF6BInaVjbQklltpT2yXzA
5ouNOX0lh0u9nFvA05wNQsEDcmZ/WYkM8kYPkYAskMh2rs3ZNwFEELWbQz1Jie1J
1A86OhUNEhRG57m7NbRhMiH0FIpHRYHBAwBA+9YCc97EDsI1jdBHq40WeM2uTtfC
AOfYfrJnsg7AfanVQ+fTZFg/ty1Ce43RNBEYoh5Y3+X016Lid7/a4B4QoXHzJdvv
e8jW+XxwkRiYKXU00M+f+oRqjc+p8U+I/YfGVJv592K1F6U9/vwjO8vdHgiGfe4+
4SpcqBeQdT2lP8KS0OcuJVK5ePcwYR63BEBQA6IeTh/JwGtHvHQ4pjE1ceEFi/m+
lJKZVJL5iWtyGc2o/3Gg66vujfMAJHStyriB8ESD1aHvB2+vA0MA4tkjGFzodKs+
06Ya8Nr5EGx+gswT7n1lWCJmBuUzkYK5JWhfSybG0TFvWl5TldkQ1hMjX7jHsJav
O1phGU8NtAu6ryFIKrCgidHv9RVBeaDgDa1Tf3OX1TLTTbzbpUHGtzKIUVH2mzAH
blqhgdgaNnDuN0xnmVlNAw+FBX9P9AmA4kI3kISji60xqD6nu2LwD8yAgvc3Pf4K
fBaG2OffUWtSQgF4Md1CLJP2QcqNtK4Oqz7lk9XznABC7CTa4WZ6Y/Gd8DTOYwJH
7ZNN78mlxcwmhoHEfE7i4LxauzRu/dFDTUTAeTwD9trz2Ypf6kkCkW8foJkHs0M/
oIfwCPBTvUxZY8COyllhdFWZ70nA4yftTEg7Qw5xauSZ9P/15gkx8Xmvhmlq6F/Z
oCmi9pTNaPkLfe8zCcPVViSlDRdSJgqhA+RhHgp35VlInTap47y49ryfrpk5zBsy
k1IZpOtGCSj82pangHsmoYqv4K878Zhw0JeD+ggrVXbFigmalcUB0U/jys8jtOFD
7S65VLHYMQtufeCKIX12Nco6KQm2FO/UO8SXfuVct3OcYy62GqC4zdWIZ9KGGytR
NXU6D2Y/23UPow1Vo5Tesp3pmPV/tB3EWAo/P0IwfcuMTiFQBAIm2HMx7H1VPyCj
2OD8EDouT93mHcGPTW/UGknolvzzg1XHIn6Cv69y9ZGBprurhXTHtwK65tPgJlHr
dqsjW4yrMurgd1GuO42Si3ABxyCckHH+JhxPEJEFOY/QdbN4vE2iVKx8hX9LpJvZ
4kOyxf8bymoUAjgm0R4B8/KY7LwCJlxdEflVIAkDPYdxfRtiKjo6SCzOs1bDOg+H
29TphaZowFwuiir8QSh2BNt4eR9KkdiQPziYw8zilm80flk+mOeggA2FZuiKgSbg
i/6aZ+DcXwwgaoPl+sWU+dRZ6n249PYWWoplk3SQs/QP0LnmfESjIyzmgjXQrJaV
7KRMUu7iXoSLOvg24GPifUBEk/f26VRjsJH2gprX549iym1xMKG0vGip8QP6uuc6
nq4YvCei6vE7r7dgoZ6LJJiEsH0cHt1U8etO8vDWQ5tdsTmiUFltOzxpg0zHI7ab
jzPqCSAUJWNLT36nIK1CHaraFAniUdNGm/0jnvrptyKUDtw1lD55ZCGy1H0LpHWx
Jv4WpRtHCo+7UAbLEOdk7DL26A/oiIeXBLjc8m97KRHlmGAF65OFIDkxHPedyUu5
9GN5EZPef8q+kzrO3VlURrGcDFFv3+EDOCFrnd6IMIRyk+xfPB/PBnHvLMgDD2+6
tSjcdDqAMa5PfFHaEpxbfvCDFns1nLgwAz/zPQ8cK7qX9rIFBioQT0BMvzXdHBZN
muAWi2eU3NcSuRM5Gj5XxwGZFTilscolf6YOzFFH7HKsVpOb33g5mrkfZfXaM4j0
66sbNsY+m+s4qXD8dpX8tuxCRrG5XgsbFzC5ySWGt/ApEdUaWnDB9W5Fczdd4nDL
IxcAt4gLYQY3p84EwlUcoS3izFmNuUGbCz4JEDWHHQDcrRAod/mivdOX2OUZndD6
qw/VKuVluf4JCQkH7+IAuIOpFrjIiX13mGwSk4KgtsaLaScVnaGqA4iUjslz8vwT
pwsh4xbcS2HAvu/iJlYPZY9Cs3vGJzsYxOBs0QBriY0oFhFhz8Ws5XL+HTCEr8qL
MmlhZ0IaDY9VnPhqx6zJSw4b7AJq9adCjn2VzZQVcqDdC3p6fem/lyg+0mrxy/KN
vV0YG8DJPxAhNUQNcebss4schUDyLAJOOze7vWtzOGglbFEqo2+w5lvp5WgZYX3v
iaB1NWBYwV5qn5bknpBO6NTFMa3gcMLh5FWxlqMFvwcK0jqwfAB1PH3rjlQgbSf1
KxROn75dYpypWfFKk1gtNUBOq0IyCG7C2gUf8EBshd6xZR3vI++EluLKHW8QHSQ/
shKEiwoZxAXLhGw3BU5PptDQY4clZz18I9yKcYvvaSlS6GgZySd8cQjLtd6bO6FY
nHY2aiPEYohfuK0m6Lyk9cvi7eo+ptlHjQGoHNkaGIFL9jpwYqyJmSHMxlIcWQ06
TpeR+30UltH9f8pTqlKKDAArB3c5uahYFb04TRjudP5xKXxiggDlzJG0c/XbUuza
IiDtbqazbxqaJcKNxqe66I1DAcIA2RW0GX/vUNEG4Mcbonqr4iFoUMH6XMFdg04c
4cb0NFHzbnj+cr0AVhFKEkjhcYvT/WkOq4KFvtneHKwJvV4+sd/o464AntFs3x6C
miRKlHakeKCmaCjgNpfyMw2IHvAYZyewCxQNdm1iFwx72c5/Zd+sPs6Kxy5OXBkD
4seJojOIMGVs/gfCldDHLhR8EaZhnO5WO2ZLgIDJqI4f2zEprrlABknCGXqwg7BC
5WWUes+cXikPt2GZbEJYr2ItJGJ4dvwOyeggKRvmtXIWka2wpnhUubv6RmwKXdKU
LHNb9evoePRUyxQKuRXkh0oYToZaxpVLWAUh5ddZCScmSWw6l+0bOfiBQJ3G9XeO
3+ui3Hb++P8AaeGtrZoVpE1kRrkIRvGzASM/fUdUPNdDpJC7Pv6wXwB1hFnFZsrT
BKKxtke4bQT8yJTkzNmgu9Dqbyb07Kmb8LV0MsJ3UYOJc10DOA3CmAtfuqxZSUDo
lXiTmPbNZVHs2WHzn5CDM4+c5Nz4p2B5M63U+2UrsTde3YRi4g3ibYMvQSRlVpp/
rsqDcztvC5aO4/6gU9lqyZB+Qj1qzxJlND+K0XIvuy3heETwttcI0lTauwKM9zRq
iZ8AURa951sIJTgFiE6bfFhsanZePcHsKvIB2Fra+LnDw8Eb8Fx0biMS460OG5vX
8eT1RPzQNaWWwObcLZYIONOVoY9cDRf4BHxQuVe3eRh9ds0Y4x6TALzbbw64hicG
WfK+PtHnRo2V32KkN6b+j6qlCNin7Yr9c2vbWKPJjkwf+HCZacRRyoUJK3TyVb4X
FkKX3qcT1oxkInSrcpEucwnxQD4o8g0IweYNkuP663aQEs3ZVLYgouDkMpgmqDn0
p893rtntX/LRC23J+H/ePpqStWxGevgzAdX25oKPPbKWviGXS+Pg7mAF/owAqZQ3
RP5+gT8e0YN6Qr+N7Ms81/x2xLQRI7dAsKjy7wsFrOOEEZ+C5wpn4uv8PPxEOn9k
HJhedd0ZTUbzAZAisZjm2AOCORcLn7zjtBV0Zin0n5dO+Wch2uugU3VEizNlNNqO
d9hhZq4TiCGNaehrtE+wdbqoaG39yK/a7ZRr5lle7lFhDZ+RJFnE4uIOo+uEIuWZ
b7fMfZA8DbsqkVnkSE/2Xf7a9R9S0D3r/IbqtIlB9a0JPMmOKnOgkn3yaCslQaVb
XN6LC5jZUUuWX3Qk3lVUY2qHMvswFU5BWWmbsmMPX/wuosx4irxlhePZKWTJ/R/H
aZaEHrdonpG7icz8a8QOXdb9eRYBmp/BTg/N8tmaFeaqXE85fpYlGElhTFSQtfKl
/rU0o0Um//zpVNmMDnusTijn4t4EMWCWt3gE9pmCHB2JopXn4Binmd8+g2nhWuTQ
G2jLgDDn/gVcti+ypTcANIk9J4hCCNZR4ThHTX6VnyNqDosChmmLztBLD+pvy9vZ
gO0O2KeYQDAGx8PxQ0raMT/bCMuTPcemZEF6RIzYrRXsV9+gu36DzbzzS9anRo0x
VxQdGN7i3eCLc21mzhcjJ+ze9zZpL4nPWOac8FToPa52+/IpAua42Y+u76nGzMsf
EPJb99Yy9bPce/Gt27Ppp5KaDCwI6+xdAfN/aBA5KsF5mRudFuSdtMfHfIpHstyK
wbG/KmRuLhMlO4uo+qP7+hf4h6SqfEcwDZZs860qrxSr/Y6HLU4WxLLQhYuDf/py
jeIdXWzUeezxniDTE2QNF6tMXd0qXuk4yQZoF5+R1SAiCLExo8wrPMkY/PA7LZkA
VTgfO3Zh5Jf0/u73E9VD2zfxAe9LRn8OQNc+5/RCfb7auYyh9fV6XvT5fZkAddL+
GIXM6gycxuPuKABWPpOYfeUv2T32kMG/0iLEHA7JRpaJ55q734weUb41TRANZOzt
n+FDECYV25MiM0Og6p9ALNUKndXweNJU5agn7dV0ThLKA4Yiagl/COUI+V4VpjVO
WXt7hM+AaU8TDAgHu3Dl2gsun+02GvnaioKZW8bsNrBrnWF+yIhRD+9qqW22/K/2
HUoNn09qCmmmVXb6X8WVqllo+G2gJHWytdJ5fti8hz6j+tRQhKZI26PjtnR6GdsL
0vXABHBnVakAyi/HREVtXl/tWrPqezYmIPy48Jmh52//4Tjcojyu1R49Q2x43SJ5
NoBNedTXr2v/9rs+h7H1uDU9xS05uz7nJ4bae/Atoyll8YEt/KbGPF0Ptm3vzAJb
5HCOxWtOCanckQ0VReT9J1AyCKT3F9kf5rIMSvd84EBPZBiQITdnCxNl9bC913rq
doMIVvQqPW2lgiY7qngavjKwRxq7XOhmNWl2T8ME+S1wHK+nuMBsx+TAeQ+bSRka
LIIGHH4UKSWplni/AKwexlLcMZegXGbU9IdtB2mKUR3JpHUBvNHAPskSZUvS7EQt
OhwZcI+/nUGocuXK+gtUkYCCGFQYdLCZXraIR9OUaNX2j5irOc83dsngqTzCFhbA
vEHEYT8CV0p7SkW3HbO8IruVEh0KKqFRE0/k1eNXbr8wz6BXieJmNuqrZ57xd0+N
0lIKc3RLP9GtPApIOIgGiTL9GVvnEtMYSVnkF+DeUGIydTWL85qjroQIDRpqZ5ex
efE/kGs3aJ1lHp81SgZdK67bmBZcutsrEwL4y48FIuXdKOW+sRa/e1rfcJMbnq81
NBuzJl1t9tnIWWOagy6CagGVCw+uygl45sHUu4GklCW3JHXqxNaf5L5y+Ev9QfPU
N9ocn//ycXKdNqNSU/c41fU1TEq5F0iWptWO9Zon4UnGGmQ4LcodBfutuIf40OSY
dzIIR0+KRi/nPwaUzM0kZsNO+YOncR+PDvTS0/TVNATa5AmI/BUfpNaVRm1xezGx
eJwaKE1x0ir5WuR8derUYZYTbblTiU8HRVJjVQISzhW3lZLWg9rDuf3Y3VzXxkzR
Bpjmc+RK92+vfa8QVdCiXQT3Gg72KFXh1tj8+poM1Dr573yG38ick3Z6zpgOSdt3
7zS+xgBwCdqFMYAizPsKpgAZ425HvMBwwjBV9jMlH4yqoESRCwOWd9C+SWbP0fM2
4tAo4oTeuRgkw/m7AkHfwatb+JqQODfC+Ie/YZzHP2K11b+S4twq5+41DsfuMJ7/
c7nDtcUDQVtPMJPjDKca186WXznkC5OpYDZLlVpfOaOxs/okW3KaxXfPSwWnEfIi
dhKkNxbVsNdmKAVf/iUYWDzbxylu6QZbKwgIaC7XMsWgKWTuTmGuzVEadc2ZSJ+4
bn2C9+t6+5uDvcvMcdF8/PzJu0QiZ+mgoTxw6Yp2yWsVXp0okm9OOq72Rb2wdPZN
6oLqjtTwRnHQaXtB9vhqpNlzznq0p/W0g5kyBOeeP3j7dNYg8s+5ng0b110V86RA
qlUhLYeRrYeHLkMliaDL/QadaKG2HYz3oBqhY33++NUqML4TZR6+tY6V8RbRZwjR
08A7q/S1b0UM28gz+dor7LBtCiq/l6Lzu8NgV/sT1UiBSg20pUyTdCRHXN8nOmct
ZTzCXzfPwuGwl7G0Ge25RearVnybHBq03iCF3dDbovTNbhfhNODU+rgzE2UNNqDo
QibP9d+e96qhvfIYF+F9LmWBzqXJAyUNoLOgQpz4Kp3u9rg8cOvVBnRTKr30qLHF
nQd5e+y4RMZg9MEjEWRms6LUkJJl18OxYEEMz9km87Atnc1dVlpjppr9tsyv9QNK
SFCgRFoR2OhAKZf31xEAL0CWMi/hMCUolcgNHs0hpYUCSBTE+j4s/Sgn2qccH+aT
GkXPOsGM5WtVmT4QAtc5XiW5RQ7QjOujfoBPMtuBpg/o0sVxrq5U+CiX0j+XQz6V
hH3NkxYdpujJSIdY4R/qY9Q/82jhFBp6fphk8xwSZK7cPF8Z6Rn5vYEi4YGfAn2B
oxtht7UkSbKNu2tUPZLhPpYInaVR68qJb/TtabWzFT4wAy7LJYP6KPguGkiDqqw3
S2APsAmQyNinQumtB+K4KmJka8zjDeaDHP8vkjZjNJ/iqUZn7XeIOQX+HGeIYbZf
afRO/5FgMpcd0WEQY+X3NX41jleMqpsDOowJhQFEvOY8eGeKPZ+KMj7NJvyIcCvL
iG2MUSiPfMtOcf7lxd+H2f8ADjPXOMbSCbo5CIhG33HbAEj/w1It0AuTWdw5d6/T
ew9+BUEtEkqbd0QqkBDeEuK3VlzGtv8ei+Qc3OFHK1sxFw9WjlDqpnFTLOhzyiXe
7LtI0MmyX1NlUoxqRrLUtRITbPMDba09tagYYenZ3v1OGMMylTKwddPsChm5lgPF
ktuSkaQ4jhFMClWkedHvkIUOWOXEuKoXwu4vs7eKvbSVecAjGsA1oiEAjggbGY1a
s4wn68OSQkgqenJ6wEtEPNCnmNl3X/GDszccjLqA+EH6MGVuXMIbjhhO/FEJMGwv
4kWseSotU3OxiYV37vjABWfhASLnx9Lge5w8ymMehR6u3lcJTuHS6tlySFmc8SwS
E4sv3b4CBUunaqmiPXMKC224FEHN6bDCwGuma1RSkW3BonZWxtOWSd0nXpBLsm9P
tC1uPOQUrskPAaZ2SgL31EWzYGGBi8BvPRqNT1Zqh4SRH9R7O6kD+xZMbwjBlrAp
CHi5ora2jtMn5LdbAVNPb3VloabWa5+3oiebYvnVwWlCHhc0CBjFytzZyyo9DlBR
jhk/QFCLHmR3513D5TEuJBz1D+6EEr7n6R8neCipfMeZVq0tWoveWDEBSYCghpqX
DNIrWU8FzVVFylw9nMYK7TJ/k5LznLlC1bD+96pCIQR8msR7cwshWBq2+t67Wfpz
i49y3HyZ88TPIqwVgtm7HYXSw2m/NBBSVOydM0igvBGj/edTOuBLpDcafYchOdkW
RuqUdHK8uLcsQgQtGf8lh+qJ7ftnhrq7O3XQggxZOGODcmtxBzBTPOy5x7goHcsa
oufTYSiFslS7d9rHn8cH8F7QDsgp7Fofdve5WVIoESgbU5SoY3akXi+sY9+9wht7
KyrjFdia0MYrR41Cp9YreasOuSJubFhl9sNT9uPY4ZTD6xXmCisxhvhZMpOYGkHr
QPI3Z15Xfgyno1+WLXWLJ4L4pwxc9iGArj6SexFESSeFeKfjPPU43ghXfTRMNw/q
2Io/ddYzdq0aVm+EryGXLWoq3UuYOimlUX8sQuJxIU4UikTYLJMu6sa6VsGnwZuP
9Cs5qjWi2MApfzSODLTSntwnZuFCtvxvxsr4uRLDKJQ3GEf8DwbIJ2xD7tYu1pvO
Mw+NCAbSQQRP1fAHxIR1aNpMzFlflpCBWrLfjFgTqT7I1FV5yMo/QCKtR/5KLbpf
nKxJeJRE6N7FNn87Oiiix0t9sBMjXI8q9oTd/6U+OWmzDKcuwWJsNRxK+dz9ioLq
FRiv0wkAFjFoFzjSsiqcPq3wEsqh8uXnjFk7gu6gCLyWbgqIKTxR2xrg688PHCw7
XQqpbiv8xWGCrTffbbj1xy1l/PWCHGiiGe8RbFK17DqcoftdEBZyLxiLQ1XlbSx5
8+IdQhkrpIFT6ZcoHh7n3enKSipP7pxq6sQOQtauypemGZ238Wl9o6WYpk10JEiD
DhVCeh1/Beg0yq55hY8Ug4ysAv6lU7mENBOVcEmXdi3PYs+ONP2/SbNVHQZr1i3I
QfkPmjRMI8wYHrqGlpzCRuR+emsuwXMMOF0qJbNslA4avYJfKV+5EHyLmq2pWcrk
/uzoqfHegnpgXGQ6rMOtfUqFtYoWFBRZCE88R8S4FogaS/w+9QuUE/hy2AsktPvU
Dca8GJdK2A9OOgpu/892np3b19wbPs+r+A3JUFOwtqJDWRckLivHc13RuMesTNTy
7WNwYBuhuNAtwOht2OVtEySWifdj//qEv2GMar8F+lLIplsfUqQm6+dRpO4JBxWZ
rV0mxmBrc+hH34mR6Rxz6dNxf6oYMvLA0ZJXTjKZKBcU9g+lV4mMMB2VVK8XlEJ2
ulxDWjsrzfiWFUIQPFX/5C8X2+JZ37FrMXnx/FdeuIjvzDzjfmzp7Cq6wZ4rv6oE
djlaK3Nw/TbaZ22FPGH5PP9qx4KMnn9oyu8EyyRJj+fmkXKKfWq0WUJAqpPYVe4t
06dWgykliWvsLODM5geFXgGRKaNN+nAeGDmARxwX+11Rv+rMEpchhg5nwXyVYV/I
mcbY0473fUSxYcYHvS0tEGuuWo0lReUSNCKEOFRjgX46iAo0IhWIJs4e11FNJ7j9
alTa0hKQodhKOz8LOi/EuzE7O1A+2hKnd+Xv21iKgZgZBN4b9rPZ83leCDIGWG6i
8gvWtkAJKh03O4vAST99IyfGkeEYmN9nxg2CowbGXli/ZDPYOlJSiFYSEwwYkR5e
K5yVgXlBUYsJOoGNq89r5fTR7MwGSZaGWamGM7VARLa3quhuNm2MDp6ElosMjqB+
Y8/TxG9qa2hk0KMDKXOB2QACcwFM7IYOCypHNHWkqhNryeaAqCNCk7Vo/kQptfj9
xPSsvUq40mYv9OwiVRpQyGZPeJAtUW2vCfmSZ0KDkxPDb4ET0Ba283Wow/3iOg4c
cDy8OYDe2xKPIn/ZR8CveP1BP++h+VLB6bUTla9R2qBePu6cy2ghY1/uZIeQ0ySM
gJDc8H0bbbfRaKLczaEztJKexfajex1KyNt+TIgEf6gTK54G+XE2T3iTHCuffp+y
6u59EhRUiADd7lb0U8FJ9wqmmBm0E3LCSuC/ASqLQslfF5Ds1Ubcl0yzfqHcdCGe
4qfpXCWxjNCYPPpZn7fUYLxw1kmNxU2N8Tux+YO3CGVFLKn0A2zlrtieNFxgeGAo
Jhe9awxnCPbOHYFDzMHoCG9yetOh/WCFB6vVPFSB6wHfOtdQg3oiBKb5DC5PmQWb
rCHqq8g/jQzvRbgGfLcm7OkCxV8XNR7RTJMgEj67iQXGPFNx8/1ZqvfCsMZ6sPkU
LrD76NaG5hyAPHRlar1v2vmObcWkfP2uHrXW++sKDipeOUqO02wPQcAAh9KuxOtu
Z40Oam/jqTqpwgHqZp3i5UTueTyWJHcpfVx6GhN7Mpi/W2NNGYTSWKN9rufOQfjY
WUd2QytF+rcSQhnLNaDoSbegEaQQgjHkDJ9ThdX85LDDtRbw3iY1vsMSE4sOYYRK
7Dz+ZWt7+cqjBLKmoB7dn9Xm6sadbdiL+7joPkGW83uhhPjbw3KR+WRmIwmDf5g3
X8BLpiQASBv6cvoaZDGpOj3mjRulLql3HPuoVltXLbzN8HpXMR3C/X10mVBZkzwv
k/ZDxiRvaIQ+Fa0LrMOHTmQaBVFSJj526iIgAVllMsc9Fr6QkrFN9FTVx4ZJQ3Ld
8/Jxm+koQpSAPq4iGps56FmtQay1UFkq4lgjlSY+s2MCQNLYrFmFG0DSQYuTljRG
s+3vufnhWvnf48S3/hiEV1rQPDh16QZpaPOinEnZQibsZos8ATWhiCsW4goMRzBF
2L3JqZmmVnsaebhLjtnbijOcyf275UN3bUwzAzljcDrypFs7diwdJDPRv7R07h7L
kX0L2bqwGNn5zihIGhTkgMAXYCaciP1/4KVtxyo2vtB2gvEVZ5mKO3Y7mfHJVbBS
guIFlb0OONrJ4KTCA57P2TNr9yj2ZIeGXTgvCrs5wIwxgeBkatf06xnuSL8fwAzy
3Q/fZgwiuNGj/tenTYjXxgOoLE4b9sjApuGnxOmoilo+YkRfxciYLirPoUO56bkT
FQhuKiK2aNcoyAKVlJANJmFLAoZ78+E4fX9fNxmiYpJxy1o3JSZ3DS78jyu4ewIj
GLQPgsL7f5Gx9aMTsrWbGkH6wxAI1ZSHECzhgRVCAi5Vn6VoiY7Yl5qW4NAJLO4C
6HGSAFlzft+Y0KPkiRg4+0s5bcouScANMXI8reUh+2ctc+3GV1+U7n8oRFM6YdxZ
2y7vgbue49P+YJWEi5PcWDHl8EklQ8+0j+rIl0r9UeyzspFW8AoIeW2AKriQvGGa
cJ9YfgPFqcByGiDTl8a17a7SDJVyyzQUQHF8UZbwkeDfpq+phGXanmkMrRrTStW8
zSkBvIIoAl0Nh4+IDpgKXxEcSqLQpKIAZoq4ElG+1tdBXT4k1IvCHKD/DQR7eelR
IBOoRuEMubiqZatCWlcEFToa27RDNTRAMCfF8lD4oV/SI4DV4f0/bmS4MikZgOJ/
SVkTRkZ4L95VYrD74PkD/grRH1DiUXGXiQ7QQJVHwlKIyM82/slou1E2AVcvipCL
7yrxDbGVmIHZzNdTNaIBPmxk3yfiyK9WsWdELcipVgJ1GvP3XSyA/RXALyWXvb5a
p4+bnzwush1q9EZ8cnkE7/bVyYthPZVlZhHCQAYTu+Q+UMVXSiICeZRb24/FwbPF
lwX6NpozE5HHBjCa3LsEz5u31TA8vU4KLhfy7Ri2GEiDpG4cZMvai2WfQ4lJSfj/
8uBf8+1egJnQyzBG/NhKWEOrKj0CydU/DhS9AKVKXavYgffpCJORZhBfHENl4E9X
sGlc9UJKSpI/xsfHfj6PSQGce+8NOPhgsiTDJi7OuCb1aer8Pnghe2oW0M1RfZ9S
FhnddsP9jv0qF5YivHMpGmI/O6BwzwP4UnwLHfPJwSi+eVj3lIYpEwt+DX+U6LO0
jyyqRgwvGnqXas2eU7r5zItiiD0u/qMsTVNG1mxiD2lucQm4jiSsIVhJ+jwtHqZK
9UpUYMVAAn91m0s9Q4IfuWQCGV13YRvQcP1zKwU8wBFohFh6uANMHZvovpTSjRcv
fqMps5cy0yuEiyKiHasc8c61zHWH7Y/dXQA5aMGBCRrMVSzk00XNXjKdznTI/atq
g6UstRsvO56mfN4eXEZDKMn/noh/LPZOdWf5O+DB1XEp/gwPxRGDf0aesVPEuwk1
lH4CHjn6fwtK1ykVzM44BzuV+CIldbUQsOaRXrEkEepgHHivx7CSKHPooLZUlSep
OaN69SaA6AMGA54lg7O+Jn9clC62pCtSA6GgFwPq65neoVyZrIJ/mvEKetfpTm/S
ZbKWT0CJAA1jm+MMaqT5d4C3F1OYyB2BZH0E2pkGEUoHBec2X3h1oGw/GtfxciyN
ExkuW++d1oGnlU3sav/1NxdymZVjsr+D7gX68BcCCQ8feLp89LR3n3nMy+p6IiqI
Bvep91TjgnTh3eVNbbRWbr/a6rM6pH8RfC5F4PTxuaHyJ422wTuHVueJXH38JR5c
i+a8XXTxc+FcNCRyl37CDJQi7pHKRaO3QcO6L0rS8+zVR8ksXubSHn4x1ikCF5/0
wYR+v+MfdnKONyR2ofvJmqxvLYCTxN9FDLKJMlXREK2osfXlF32ixHuvxNAceBQW
k76lPOclORtllnRQkc8IQnI4PR0QfLK4cv/dUZRG9Li3fgQZOTqdOxhV0IGSxR55
8hY+107sE3CF6xJIc8ldj1IjWtqBNN7LIPP07gyQhOIyWjiVD6MNHQh5TrCULHMV
el5nuQzYi2mE5pyuQk1zPkVwOME3o+o6VXNFkoPp+ZnT6Efa1qW/w/VRkkY4DLzC
xFuTliqOch9l/fK7F8losOMm4gwu9qUXjMjoXvsyk7VjxN+HI3m7BvOef45Jfnhc
ZXc4h1W4m/aVZhQBsCQ9/lAwHmde1FfQpGosuG6/7kBiSlG2DWP5J7iQU0Qck9Du
fuutRRriVnLPG6mOfYe4N7/63EvoExy0Gt5C+hHhX7r5mcwwqqztavBM3VFjo+y4
1VweLOB5BT30aEqFHgzrZ/f+doTEOQZ/PeNx0bjrAUhOUmEyI+H2RRBo6VgASESf
1zy3a3J6eHCDiEM6RtZCHcSkczHyFXmkFLrc+cJJrlF7YY+Kgp+jIdGE/ZRvOcV7
xjbBye9I0pPE4AegL9dAVqSkA0u3qVX19Un8nj9L90MFB1qpmmuqHo0jV+LUCQw9
esTy3lIPQTv0BxG+YXLBFp8uCF46Lz/6obXfmKwyFgvPjy1JX+r6CjKgUiA0QzRk
q9t6RGNrI13EF0hqziN3JeGrEEKDiIBZ6eurhNWve4piMF/4vB8ehH1g7qGSHnAz
+q4rjMI2l+kCelQHLiXSypG3keOonSN5uh256mkBvOpz7i7W8yBPDNJSATW8akma
NyVZK1h/BhAaaFT6KYRnxOsl8QFu6HXRQzEJpN3Ja0LlcjWXqXZdJj3/AXQkduQX
JC/AXv/TxevM7Bx41SPBHZrsjorS6ya3Hu+TofoMaYFA0D4LA9jayPyXLu263YV7
iB97+uQeaUDuyyJzeZM1iMwVD5dm+urHV3N0ZaWpqBpmuMxblIUaOB1byOKz0R5j
eA8OOKGtNkfggQPf2wBW4KYVeDiswNivVhg4W82sBxDQeQId58CclQZLJNQnzOv3
2iZrkdQ9rMWm23m2NILl42mDgDtRV2SJe0SvQiwn29DnspmzZ753F86qJVJn/jWY
1dNwGWRoAEawHEFB6ObgBAD9hf0L3BSPEdP5+KwM9NVWLQwVFasWAdRhFDitwFrJ
AAuGz4GoV6akcn2JwVhwnZz1RH5oogeris7NCLUpc4aJDL34Cbk2tyFluFY0d/yb
Gz2rJl83D4T0hTRKS3Bp5Sjf0BlePAwXXAtrOL8L397f3AQ2JRix5grGjqe9g8xI
fKXd8G4ghGv5VeErpIvK5L15a4LcQ/ebcrrxg19DZF5W8Q+8nNBHtumnT+E1UV5b
kUjYV6TdcGXV//sgPXXD1XYN1lweMrv+hBZVdMrK+nqLRTFP5qW54gDa7kvrvgVW
aeF6JhdDyz+op8H2Z0brmP+L+ddWgdOsoF1pIZ01xfZ8B4vHezNhyO4pcI9mq/v7
ZHfTMaLs1O//ar/RujaxKln2wNslqBeOfVYbf0zaoGxqPCh9qrI7jdYITs2gA31X
wrvgg9sBeWYDTppB/RiEFGyc45tRP81/KOYGGHEYJ2UpNjpPc/SundIKEBO0t7S0
NGPVMmDSj2owrRWf6QRDxBj1hn97z49G220q1DFC5jwNUmdscdSyDShG5xasSWWP
jWAn6rMnqseNhYYbKtr7A1hEGewUD2UKmtKUNwtD1g/77224sK6b1bDp534kS26z
ECh+3YnqphGTZA0TAKaCjVgp++RQ1jOjW93doWj2tP3HFzkW2UfcaDjGSUBCqSaS
8F8Ia/lkEckKvmhAvyp7stppFAdvIpYxz9O/Gs8gn5gy8hKnBDsOzpZ0nWy6wBBC
K3S1cOUwsZ7uu7LxGGN1RwhqCAQWOfIH1sCLa+7TBPXtJq3aNoZmFCNGtwWHy46Y
30+w7iGfDFXQak9qnFx3v7nwiJlXFr5A2uFmiEJyvTzCtNbsX1txwxmwA96luc8i
3rG8P2Y5KkFP2tp9A4EDPOQaYBEO9r58ovPLbCYb1gLLm/gx7MLjuD3OGbzu4ilm
9h3bN5Z+KozbIUJV+GA220zCaU4WNjIUdATfmuldQa7XIFBuALi+GZdRLiSUUDNl
nFTap8sc2EgosMnN7EwbDmk1cYvg+lqazEw7mqlQsXEhVSRxDk6bg6lzi5+awxwb
dJzKDdauqaFNcNY7ZJPBJH3oTfCLF7mFwi2rMsxTsHd1j4gpE8GmesRAhElctG7y
284O+LXY3HSUlw59hoLPbv674X7qL+iflSZFzI96i3nZMjQ9kWPMwpnH1my/oX/o
SNwvJm2REnbp8VO2JSj05rA48zh/r7cfhoHrJC+slsBCAhn7f8SN3M4xM39YENTD
OFRuwWaLs7NougzF1mbxy9JJLvBX49bwWLORbwZ+4RC7ErW0Ktbm3aggC2SXdacy
IaJHlLbY3aIQjMSQfsPvZBrasYZTnnYSXYoSlKz4fVaMjYgnMrqVMKkgN+SUGzeN
0s9p5ejwA6f5fo1WiqNIiej5jWdsV/I9q25gqKyeTLVRmv84/ia05OeIEXz2mHOS
SLq8iBn/xMsMu6yePwd3cekgvCXigatt66drG8q+xhsENLTrjjjAZwm1php3KwSb
yob0CilLKCH9kNGkv1xRzy8FH6B14T/0Vw4WwKd9AN9eyyWJiM503BOosZl0Sn68
c9uBsO4RF7feEobYAg7IIa7aaSmUvIjXMb8rGk8nWASwHDq9lSkXBSxNenSUUY3V
XYYZIN4oc3c4HFQtKmeu4xaJZlhiJ4a20mDYBmR1LilTmdgqXl1h7BHuedBKw1kn
PxfFAHpyQ6OiwPh08JU+Ov9w4CquPmsilDZ4zask9Ec285d490T5AUwKCWqGUUF5
bknnKPVYMV37FHSjQUS/1D6KIrxQZhYqIU8Hib8avVxvjAYSoN09pDT0PsE6Cecp
eJWE1tJbY4KfUSZHWm88bPBMeP8F5xUmurV05o1vEMUvpIpM89tDEcKOTzpXXaRM
zKxLzY37rVPwNkM6A4jr/AvbjKtc4sEUHdltxaK4YE4nU3dXMX0EuRBRE2JXt4DM
2DIkEbMBjzEEdLMBwOHKsgZMArLobkTQbGBW9lplSnmf2h5arY5qC1PjmkbrWTq+
wBtSixyYpdeb+Nt4eTxZ5gC+wjgTbnNaJwMyAfC6TQxGpnLM7VdP5oKpr8sSpK2j
xOLMy0dGVSLgY2XAYElunTO50XckKhVmng/d9uAMuQ2a/RMc3h3Kum9Q6KzEcJ3P
IpqGisOz/HpDPmwJW1dDBqAV6aDRjHlBZ2+fHuOwmczIr2U6ilmXRP5XSRQdmTkO
mAUuC+iZrVcCOQjWjPRRZfCHBtJTUOIV7eEop2cZh3XXdV2GVERh+4BXrTUPYIWU
LymQRKy8VscOrnEu6ev78UR21N3C8b9XzflStFDvmK6pOxcYwsh1HVc7wl1GcuR7
Fc34ZXGGywuFIBZo6/KMncVvW8nIrIEAFfVkp2DGEKmkslCjrHz9p1Twnkr0svPu
leFCJ2FzCUbcr1iqfgeKut2Njqloy0a/H4RX4DYmAC0XwqJb5SHuRqKjP46zaKl6
Fm5dBNeVgnGlBWhIFHyEB41OMXUeQ4jkErrbmvp3djocwOl9U+L9QNSeFvnNZzHz
26AGd3aJoHGWlk4EV8F1+rKQfUfq72zLfZDY1rf6Bc/+Kojmj0ZRaLt33rze8pwX
YpJ0KdzhacI1sAf7qQXBqJUThFrl2WGshxUqVCNaF3f3mB9IGQkhVcmW4WXcpGPW
vBdpMpjKnnHhtSG4Es8sEHjFaHGDTpVeMWqcSf19fHVrkHXFXi9jYdYdHO0ZM+pB
DtGG7UbYReOAuXD8RRjxqmDwF+JZ7v/7Pny4zmwVAqLfXIvYhs9KHrk/gnmK04Qi
Bu4aC/JvqjspkyLxMS07+TxvGANcXnjk+QbCgtQF7pY/ESFZB0j122FtTcLk9n5v
OSrHiZkzdtlMxS3aIiZMS1l641UoL0XZ38V5uEWudP7I3eWJ4uzaK7Xy0rwPfYoD
uwzRsAszU5yEnX2No4/a0vUpLqE0XAXwQ6gzfLGBAyNi97uCYLGL1VdnwIkf7Laz
SkCgjtzUGLljc4G880byx4CJfgfazDZCnalFhBxVX6dlOnuIt6bNhB7Q5amV66iC
WBBGC72HtcUMaRw9B19LfcfxqHYXfSJLrUCiQGccb3NyQt2rvnrJ57q/Y+PME5Il
MSxQG2yy00YwOMjbpDs4N97T6PCa+z4w6qDRJ6FiTCLc/5qi4y5VWTpq217NvPNk
DqJJaGN9sQGY0JvBfUMJvumr1CDWUlxRIQQNxPwCJBk6fSJQQtWUBqpht+G7S8s8
qBTVddV5HkdQtW5hQwwO5gKKBVBY3bdMTaiDwgoynAehQjraWx2pKj4d59C6RfPd
CLsD7/5pRK1dQhs4nZ+Fc0Xr8kCjB9m7eyhQ7NP2qjG1x7HMNookF6zz+mmn0Z4c
44ydMsxil2Ec8BQNLFfBg3yu+VAZn/+9HIbcgUgFDOYBvxf9RGJSknaQQ0ROUlxC
nAjs+fK/ueNsSbYf+07RQ3VZJ6xBQDnf7sWc8SJF8AuacYNFBbjAds/nMcbR4aOw
IJ6+79Bg1eCT0sQMdT6aqCuwweF7nrXPezvQBr/F6FgCd78NoJ6ttw/+D0GzfpYh
gZHpgTtngdHePccHx7K4ECBQcPz9YUSHIJJ0KG8nYd8PNfapEmwx1bNs4I1CuqMw
VI12BTjm1Vk1sLEzTYtZ2ytNo9Zqacyqr5fqGDjJ3fJbl3MLPNVe/SFHw/xHGkNa
+TXv04ewjpYXh7jJ2kBbuqCvBBwyfk75FpGnj9tKauKq3DmyEl7su0Y/pWK1Sz2S
iMaiT5od0HrQ9cHq5BCUuoDPi1ZjSGlp8M18qvczTQgqyccj2jX25Rg7uDM3GOmC
gTswhKSORWPZm2P3LaD2N/chjC1GlZv5GxbcQhQRjs+cnQ4AYxhQ2XnJJ4hb603W
eL9uBCnsf7W4YdMAm+avmfBKg1XT2vWQG785mJPhFAfiRUWSIz43BzJNY+DjCA8i
QF8T9wJAbEUppdb05a6marMtnGPpWPhjiYgTMd4VEbBUCkVI62Eyw6CfWoydNFXC
QRyrQBHywQ3IkK6n/O9dFb5K865ybGeFNt/fljjntBiqsYhifHHA/RxawLCQpXHw
s5pUgpo9WH3SOcZ5JaWmGMew77IIB8mbtN7vx0rvXeLHFt7qK93iobqKpdbexoyq
7wwBsZyuYvJL7D8xK6nFesY4SEzzle5j8lehUjlnpNsMj8I0DJoyuOV54gHc5PXi
XQgA4N27FG7Ieqa4+aGRq+Kysk0hPORUjJXYuJctMqp6Bte3JzaTHEqy1oR2BNRx
9XfaTR5M/v6LOQL929kBzKM867Lgbp5o0CUXocjxKGm5V2bC4t4aWeDx7qmxA6iW
WgR20Vl+bLD4dVHww+7DsxCdsj3r/dkR4plpDXzKlppoX4Axq6Bbt+sf+rrCpXDQ
mSdOuSCN1qLPKkyhLVAdMaCAchDRcNlR5PILxtV4p0dzmU9WC1ihgT7dJ6NkUY4R
Ij8ZMKgpGJKwCNffwcz+OABklNhowZ2QE9mmwf3Jv1dL7ETgo/ZPE9ffY8L7dfER
wLJyw7wmOsI4wLgvRhtqgHoqzb+qwwBEk0xjCjgwpVn7Ztt32HvWkQraHFRb466q
vXrHBAiPc5fqp5c6l3GsqBkPo2oEK1KnYs4wHcSeM5e1ESkf6V+q07/Wa+oN7VE5
nng0lFFYLwDBz24D7ZtQOyovTVLcE5yjNzHFnKBYV+ziDB3YmICvQyR9YOt+ta6+
W0yTu5WUc5oQjTqy3JIa8uKriLc5JiOjnjtNK7PQwiiXbtKPtTrs7l+ZW5FQabov
HNrlJQ7krFqSJIJ78/FL9KyPBW3MVsqb0285ApM18XDWNa91OIUwH4tMS1sMQlZc
PZoyy5h4aQ+gDMl+FZyMV897elCMvoFPZem9HQWSM6lwAU8YcvInylNihOD9e6Hv
PfhffKaL+uW+lfJRPu9MjAhzxqlNFaqDzksfGOxDwF2uMMgi/7wjvgjcd0p2PZ4O
F2JLsyareEyyYZaqk6MMiNalfmX3ZgRMHmel3+2yMw5c/zWUXmHINaTXMf236+HT
pZVSaZGTKTMo9eVeKHep99qSMd6WM2XP/l3JEFTMA3y7sUZrMnadeH4XgeceoaGg
jVjuD35VnNgcDpvzSLUvKSNo5e++2DqZQhQd/Jsaq58UM7L9sKYGYMrUGHxWJCYJ
uhmChEu8Wc+XBhM7eeyJ4JvHDVp3ClWh7SIp2zyc2MN+foa6vxLkhWcPtFz27SAw
4LLgLCcMIvmoyvOXlxNdH2h81dhftK42nFi1rlD+DV48yd0DJRO/iXcF7t5FiXQO
M3+dirK6sWRomWpM3I5MlCbmFvpspVNz7rKr+dmcglKNvpWcSzapxC/DME3ejhDO
YfYYrjC7O/LkoJrZ/erIloqJS3GvWl3XjEwFJhjiHpHM46eAioZFogEOlk6ql9gd
hqQnH14rs4u9ZB2sgMDGVswl2eSQ45PnqSDYVedVzwUhKut17yQ5wazJ8+hjZll7
R2EeQm3FZo3RiVqSbHY7hOtfeuMpMI9AitwagLGgs78KxyT2Md+Ql54sbNq+UJx9
XPMORwTLk69GnBS/mIbmhXbrZmK2H7DJTnba2v0+hhXcU2dNuHfwZMCWzsOtfGnN
6kU5r1jUPkPj4BfXQtRPCdI6sHmhQPJFT0iBde8gAc5isrPfskMS4GqEXBFQ7Fb+
A3FYLvLkME6eWt0koDaALL8qoS0Ec5+MxWR74/TT8Zhj3hJb2+3Tp9iBWowHr/+F
+E0RyHVHbas6OUBcGBj/uMnmlyd+ZUvzAzbOxfDGTODyEtNzi+OcUXVg2wpahacx
dbb0t0TbwyN9M1LGkcW1qFXtenT7ZijACi6/JDWkdGSjSCJhhUmkTnxPc3xM/giE
yJaUegTj/sP1BQXfkM6bJEEsNDktCGfHpkP7l9HgxQgoBSxMjDG++89wpXgfVFnO
C02xih9cgTtX1GcCe1JuAht+s1L9+gH6bqZf2IvruRaRpWeLtyaSpuFkXKXls3p3
9XgMEmwxKskNQXh4S32KOS+2Dz+MvXLKSwwFa0co+Z/92lYScSvAdhMjgfDLgcZr
CysbI9wZcAJivnIdyhGkLdT67fZknCCt65hL+JQFBnhLNq48biSe6A7kHLxQryUs
DeWOxSO3SllEeuFMnxbI629Pi73S/jcfRfZXeRBi0ywg4pYx4vq6d+Nyxb2GY81c
Y0Psi4zV4Gc2r7i10y2DIk130ns6OlCa20qnHe+fs0jNQFPVQa273WkL6/RUDIXe
XH1p59/3SHKWl5F4Tyeg9k/WYHVMvs6pOcXTmv4m3jXNU898/LbleblaHAIyMZqO
QaQnzRoia/OEbgT4zX+OR5iZGlOfLcAO5MQ630vXbtB4eYPGXtkZ5nXnqC45zsQO
NEnZNSdVZSJYj/y53ebBsC8Vzzgvgby7rZWNmlunBMTLVSCqkgX7a3C0gDxAYeqE
H5JsTLum41AZCdZrVY6D+epWcj6oI/LH9m80V4LFWVtz/FdZjujnJ0euZ+FTeXQF
BTd76NpJTJCltXYcpn72DgrVo5io60WY0YJmw5J7a3CiCI92voa0DA3R0EEqE9vJ
DE3Z8cF9djemQnUKJPo8YSgkJkjxNlKsWoFfFa9Rp6cBnub6khKtLPNg4xq5zsNj
wrGzEMTS4hKXE5v9+CiaMQSGapz8xiU2NaNsL2igxH/1PScvlPQzd67d2ybmC6pX
XKdrMI/karWAKdhWO96qrqaWacm+Ce58sKq4ea9jeUZ2eiHpRmlxoFFks6y7c/S3
dfVX99KD25GgqFfdDhFuBC4gslfyyAGQ/CsTej/SkTXhK+LIrFvZUyDnR18/vew8
gsiE/oohM7SBSje8LPR7+TUeykfDC1intrWI9c64sHXp6JfXTIPIjBrKnjaKtJRd
Idd38aFLB6WfvLZy7fnMNiSI/5zppYBNQlB8LAKMlqOItmcSqRp96UHgKNJy4886
y6VVZ1iCrfmhtDt2FNT3AN4YlsG8GulEGfusje1cl28te1Gtslgq7GCQpsOiEBc2
QIQfPF2CaIFcXTXLdFoxWsatzK5dmaeIHb8jGb2W1fQx0LfCdfkPVNN4tjX4CGFV
FA6JlZEJEJAMST6qwY7Rgync7Dr+5OLj2amjnCXK6w2H/eqAFWUtJePTaxTA41HJ
rlPS32PsUGmimfonUnyipoaemJtWeEcEaZ6i2hAB1DSf7YyLV0hxGF+xCK8+kuXM
VUBpt+f3fORGSi9NKYOFzoaXsaaV+ueeT6MO/wy3URomiECMR+FYvvf5E47NDgRe
f91hU8KGGu1USIv7coEYcEw8ou3nd2XirnGgbrU3TEPExhdqAPy2fTztJBQ4iQsn
vn0TJdhhm+M3qGII/vwN2gqK36CA7yrzmo7rArbnKIPor+5Sn6FT5yKFadDqTHng
B3i48SjvI/hOm6nefVyXigFlMDssW1+cHpRSrpqCcmc8AOsLmtGGYQ2R6ZWj4nWu
+DqO1Ni9JlqBDH3lAFbNg4ujdliIQi9uEiBuZicVElqltnkJ38WtUVYO78k0JUfk
gb3ipWpmzdf6K4+2YYtf3vBtxBv4I9QvnmUesLOFPJQZqCbPNpismwjPe12kc9e8
v6AEVcaQeDMNNhg1pyi9y//ow4Ygka4gCZZYZ8ZaCNjxIo+tgO8R4+bzFQI/U/+d
O7w7303cI7dPC1277Y3Ra0hyvygZZp8ap/LswAqilDMUqsKsfxn5Xf6CI+YoBTP6
zscLqrPK4O1MdOFdZA5S+ixgIkltVioPLVkQhuJPx5fH3L6S79Tqk3Kt6elRuDQi
yGl2xwjHT6SjXbrO1iEPUHKYwl3v4pdJ6osPLBEXKqXCAkiDe1MAiC2/ibLnSXCr
936icJXzWvd2udP599ldun63JyN7JwvMuWax3ptWhcj1GaRlMd27Ad2AKKhLOGgI
1RzS6CwkEtynkCbxhlbFDc3sksINJzZHjtoIYrq6lOBDOvupYJtx6KIMuokbkpif
/EbwS3fFKR3/pFZa3ziMqAhH9vwfeaa55jYg8rpwFwlXS+Fobt/Ta285doegdFYT
rQJgLx5u/oYcFNLQDPqZVPuF1Q8RwnEc7/GsiPJNvgMnDDg0pR3kHgSo6DUbV+kt
Ud/DxS0e7ohqRBJMOSM6GoXRjePObgEvh8tX101WoeO+D9UZbSWP5rHiIMxo5Fjg
lkKHIX2qgcH0iioMEgOe5mjiPrz4VtZ1Bh8c6LyVP5hYBjx8lU2VkWZdBLl4R8FD
1llkSW1aWjvCWL+O9Ob8y33Gmb8eTXRgudHEI17ulii5nCbEM9hDkB1OFcNPS4/I
UO+cIlkPombKx4UKBeh3WDs/105D2e5Z1uc08Kfk59W3Q6tSjwkZA2C7kvkhjZtr
KMXWmlgRSv5l7gWJn//U04+n1WKnvJYBzZ7AWRBI3ibn+pwv/vqgXI4b9gnGdqsI
fer5KOTVNU2nxDxIn8l6iP59+j+Gsko94r9/NRZu6csclGLY4NXfqGLialqx89JZ
Hq5VrJwyWvRXv6y3XGn8aEwoLKDs34qyupIv0/vsgSTGY9oJDZ9onuNXzg0cK1Ou
dG9n70C2/FGZWKgIs/xi7hosN11GahmKbt3DibbgsCaAh5pjvbhVV0hXer1BiAKo
8zmT25x7gG9JoIB404ekMBWCbBhtD4sW+eDcTQzRNZZ/S9yt1cy/kbzBou6PXmo3
87YdtxOLX5KAJCVVO8P1Y3JNu4BvRNGU3+59d3mQDipvNhgVZIJpwVDy1jJ0k684
STCKagCLEOni6AUS/lL18ohry0wWLIyvudEb9cAMPhNfwgdLTsnHyhap+b2+nt52
wgs/0tGuz7SF3zeCUvxi/4dmhTe5p8xiSJpK7InRX6i+Nhg0dPce5wLUAcXCrnmG
iLKJ3ME+os14gbo6Drhf0fv+qGMEjyeLWup8jpX0Es9mHQwYG7g4S/tZMKPMkJvv
kMPpMPmYdvF1ppG/74rQqo5vQJeVJJNk9nb1oBVSnTNcLu/j9AzWKum3y1Zj2y0c
Bhg1EkF+Vro/5PWz7O0WLGyNU+UPu/q13nOKduAuD12xmlYLfkIAqYWFiooyk5kD
+S0v9ZdYSmfpIOPMQeYnyNHxB+jrFOhW3xi1o5tWNoe0C8nDSUWUVUAmyjnNm1Vv
JaFrGNgOEZdSv1KD70CTmEd7O6RDY8KVFhvYxL3eEznHqXNLvtPfG7SCNieM5DZa
gwHiKV4x+vP0bXdr9ZwPdqqef0vKtBANftAQg7LskPLBGDfAj3kXAjCRo7W4S+9z
Uog6KHJ1bepXUCmK3ZYKD9+jNJhvgPlmwwEOFpMuB7qRBFYV0pjMWMFKdigt1/Rr
vM98yiossjjHg+ZT6M4VrnzlJuiGyUWUNqk0b9nObcpUUq876/8XvS00f6KNyno0
+IqXDT/WzZjlVS8ze2/NmPUsMzBxRNPjXQXXJ6aafOBx3Z3aGANdEqo7vXZAWBkx
VyTK7dxza/3fG2k7GbKpHPtaBVK7psue1ABV1eCiJIra09itJ8OBVpLdtUvw9PYQ
1KQ0zjFVnijOJfyA8BS5YzreJ50FwwD3nrMjHdOs4LGiBCqtvA6I2QlwxPsX0q0w
xMNV9+lqFHqR8Sx82rzDnzssAiR2Soyse91+U2eTaBEfspP3hmevUmJmJJAaKnvB
LSXKLelyYLMoGW24Ftf3s8lKxoXPwWVRPy2Zhd3hWgxYbbFVZDQoS0lcD0Xs3yOG
3grQ0LO8aiYwCYczyGIFzUOLXIP92fO39LacqJg1KMfRHhv1/AMQXoZT6mBAb5q5
G5WV9akqYAMhPfE49+javlUaeGKmjbNEckMRY1Azf34v9vXOzv1Bohs9/11NL7jh
cGo3PlpVgqnM80iKUAQVa9GUbI2YhUpihV+qEqiUDJ2LbsIydQiQqD8GPrzk9Ork
oxe+iElCSiusrqix06qyxyeRvgcnsXNKhXR7yXQcirX2153jMP8/u4PPbmTAuWG3
aiwC+Q4HYVW7hFtPhHGv8GQU2SYuvovSHpvsuIsd9lrXg80VzOw2lm4P9XjqoSIZ
UPBeayo+EhfOB5OcJRUWABqNJsaP3FLIl/1anYa87nCbUX46HOuY+dqw92Q+L1mA
TiM0f6p6LMG+vxEwQoJqzbtPSJoqG4RiFBUCliOJyFM9c4adV0Hgsm3XTo2FGCcz
zL2e7ag3p0KbU0sy6V62aRGqlFTtdniJI41BxFfmSxrDVmImlQOF7C9tnifF4Zqu
N5sdlQ84xsAIBmsI72N4Y2gz7DGfHnm0oUOfS3drgEC0JeaJesCmyD06d9eUSbfL
zuGGFGbQ7lZ9lugmtqmzAzkWN56C/RiOf+V424xyn9Q39r8Qci7M4HtLjRMUr1if
IoD8ypEj+Ys8LXO5SLAxDfsuNCxCMdK45fPbxmT8OPK+HctMwTZUQ+VUigmFlXDt
jLjTyVCSlB0H2VWnPQnzrOyfL/KTdEk2+nWNwGkQ+qIxJg50p6LSe5VenGY6MA+l
wVebBDRa/qSuRnsoshytKiD7p/BzlvVYxePs5dkKQ2ck0hIDwNIvSChEd0aZzWBN
CfxDOX9bJpLiydpLSnurbGd5ajsrwAksP5ZJrClaa/EJnhLoxHbvF24bj3updb4M
llakSv7z9fijekZEg9C5SU4O5CGPZre0O6yocJe0aEUYRJVv0089S8kTJzSBl+TP
FASzFTqTqMNTWiLTlS5R5xriI8s0msfomIn/TJjPiUvSkQKXdo4ywkWIsjx1NoGI
4+cMcN1EGUkN0ZxXsN003LSxAj/HTo9mBvewv/zX9IyyS7+BWGgqUXmmULqeiGlX
I/M0mwKV3BkcP2nUXyiTl82FXwScvVW1SKeyyP2IpFd0jdNeNqOcxIYtc67XlWOW
dgioBIHvY6noOPXDhdyLF/Wovev+Vr+qc++GkXKNaGEXsKni43cF3dM0KoUbM4OG
cBO49oMMWjWaiBD6OVnT7icJF6Bs+8aEc5wYTcHQpx2ZAXqxfdJq5uQI0D7TTBqd
qNLfxQCnxYmF76dIoTviy+otOIlQ92lSEgqUQOAYmP6ZKUiDeB0JQDD321KPbOij
yjhWzd4NsXA1xr0amG7cHuR2c4flqIJjfcmIG3WNuH/N8u9Ubye1WcJM6YjnsEU8
QpvilqWmpkCXnBRq6bwV70GeTqQrvs/8YXe2FCekZBA2HlCtLdXXSeRFklIwmmt5
KDDzTf7kVfX0xztgzPneD4l2WjaCaGAF4IlNTvkJJkhigFx0vM/0rct1k6bM0ObB
gd5tWWFA3ffqjshNnRgTwL8WdAY+V3SFuFOPX5G0RaMJwIjbzBCOi63gpU7n6+Su
GfT4dPJVQNmN3pjxaxwu9FL/okkM4yiqayYq+sHBFC7fYtxveeQ+WoEiI4klKBAt
5CMjvr9dG9DraLtR2cl2cqLv0wSeKOJlr3vm72iECUedinwns/5dXHRaMbuyqj41
0jAniRXE/ejrzCJEsJUkdVF8sSGYWiQWJ6SIqnjwmwmorrdY9bnG5YWLeKs0RGgN
rEvbMCATui656ldKzFr88Zb/nq7y0uYcZP3B11ZJG4KONqyc2/xM6QwjSIuQ8m0t
lq+FC+ZupeD4th14aqDQ2E2iZFZqEjIIJQ5XFm394UFvI8uaaj7Q6Yrwq1QJ5Fil
pRvHs4+spV9+ejOFgqvM6he8gigRbAkEUCFiLRwoDeUfYtMgpvB3gsipp3frWGhm
V4QuZm7vxIRcDRM1vqr31mwVXuO3VpxGyiSM3EbVNQiT5ggiMtSYlHt2LTiJE2AX
RyZDR5w6UV2vt8sb9H7ftG4YYeJWayLVwVdbqS2VDGwph/motbS1STVN0Ngho/OT
LSxUxTblmxikqu1bQE7v1dPU7R9YlHf85DGwosnLj1d+8Y9OR71nEoQKS7WqO/ti
F6mU3oenXT+Q6y7nAS0O+6Hcy60o57HOlVjC+w/bQRQSGDcUSJ4NokIv6xK4a++L
1zTFOh9jRYNiUcD8QwyKphFTsdSCgy2W9KYTBCFKd0xJxGVE3hgsvWHZl+3K8/9u
71AaxX/OBwqKSzAHPqNOTiMbGZGM3eT4wrDxtfNpA080oU/ovaAo8NH42XXagyAH
cmYskcUsFY4/cICW/wh4l+GpnFgynWdooF8r+W4XVD2VRWMZpmcP4PrNGMFXBr2+
Y5UV6z+fguImMBKIoL71sSc+zi8+dx77ZJ1eIeUDe+tQ4AUPxjgF9c2ednNzaKv+
DAYIcqUV5IPfmb9Li9oVVAJU53xoVSZcsPUUHLz5QpiqHMUcVJaq3OzsuCYE6zyc
ZXWaF9oUPmhvCdu0NONnQWSkvRwQOuNSNkueL+EDa0Bfhag2m4lX6eCYhrBALyHT
8o9rmT53XflHLBNHEvwyn9xYKmGxzYWjk2Sw9mj6kaDRstgPq3JNMn7bi+Ifyr7e
AFZZ5/9jFI4cMrzbFsgjz0KCMI5IOt3ttothNSpj7dQCAV1ujzGVQHzDsirCsRS1
hdSnNMDZqSfITNoYcPJkktf6Fy5fgAbTQokbd7+0YVJQmy1XtZ19YAKIGr/i0vQF
/woGXJjV6fNTHqXvZaEA6K2P7wmY0q88Iar1edIdaBv8jfb5Shh0MdRawLD0eUoq
R67GixEDwDOFQGpP3ezJHmjZfehBo6uPMaqg9SpEvIUcaNKcFWF02sNLUX8WsA8G
cgQsJCjLBp2Hj6YyWn1E/SSB5KLpowBH9IfYOuUcBO5CHODWEkavCb0VStY2xGtO
G+httuuJsape2UE4Jvzqb1Z5qVBmwDGJOUN8KS4mqkvxkT2vpXikVPsswCXkawEK
s4UYb/tQn/XQyaYppYO38OhV3z+fiWhl442xKxOGWkeYFiqaAXGR405APdBiM+2X
PyjONFwhtWXAG7B7PrQp0aPcGpRC2Nca7G7n4XNG2y6P5TDXQLPHIMOIXpJGn9gl
OKEiSxC59pI17qabvnfZMC8ZIDnnR+nHAt2inZi+VDCtL66UxeigJUtD8dunePsW
nXufFN74u7REmFe6O2ARnC9F4nEN4nPOvJq2XQlpb79Nshs0wpsKppa12eia5SRW
kaQudoI0IsdaxpCurQf6InpdNTDRLB/s6U1XwVyikNIAW/ZS6wA84p/wUFBpJxTL
prZKbDBKdGQ1d3hTM0qlLtjQi/VPQhujyypQGcbza2mXCrB1kMOl/E//dpILVzd4
cUMp7ltk2ZPZNnPhCg7TCdl7LfhKdJoFz/pwHx15cIijHb5IA7FYtyobz4Jx0v3i
nONr0Psu7pppR6qfh83ARzSrCNYSiecuK7QHrbOCwVIvuLUmaaIz/y25gb9vgd5R
xx71KnXX5ZOqOaVoc04GqhdImsGDXKNzEtWfmtRtvqHMa4fZMQdLemtW4g7qlOio
15lPQ9k6/DOwb8YFjIpejuyh8qKVu3QXpXmWy6yOO9MJOj9k7QYEp1i3AdXx7KQ8
hX4918PBN6+KgED1ZSkDF9KPo9jUE13AMie1/V89SushykoVzUSTXn57KagLOS+3
a2cd88fR9eE/CPoMXtd2Imn1na6Xf9DeRpgPpejOAw+WpsMN1P0N3Oz3X5CgaYG2
8wtrUPNT9vkGlDnVQ61KT2fzhKA0HDnZWvumt6kL1fMlU1Dkj6qk9VdoOXsj45DA
uAhskOTJRYutbwvNvqkdsiunCgPhPMFiYEKtRn7/z0fw+NbRXA5tkbZXg5WEYDxr
Ve9GpMxIivCzIKeHrfVT6Gto5Bv38LLh1awy3zOuuMzfdYuCmEZRHigb7M/CxOdM
4rpVCc3GtE3fkJagG/kbjS2TewrXYgqlZjM2IIYsuZK6G0gK/dx2nSw9CQ98pai4
8AICxp+7YGG9yr6xAzMeTHxfuasyHiGYEhrO6YDNhlYdVqFNJy9dgUsyz+f4H3ZT
Xxt76OlS9d1TGT4UTJF4CtWUitvIPjTUW1RVM7kbFCRYSSaTCrYWy9X/KYfaj4o7
T/B8/VZaH6gJgH9RmRbXbEiROMXfRimKwAPYuWVsosORGMbMNj+kr6IB7l69sebc
QVPfO62J4RlloEt/3J+F/2c05yvp7B2YFGE7W6VHtwursqZMHTKW2kXvGiRw/2BR
ijM02fTEJxxjFkuoi0H196TEYAZM86X9d5FTzcxuRLUihwTtNIpRHMn7ktmFnNLE
ju172cc+kiH3GBnh7P2uCRyCyMNjI2q2FQQuD3y8+AhwDsXIZAyYACv32aL6mQIm
hGzAgNY2TszDVTE4Dy1qeyUxZgXa4AJ69fZP1RXLcUOJY9Zq0ZwQKimN5KplHDvg
HPVp7gI6nSks5I5bFl8dPOhLNyPvwnHLlMv97DoT4PNN1hL7L1w2Z4sJM0RBzAsu
2vs3rV741drvjvy5FejbVVqcPeQ80Bqb3WqP/fwtPm+Q994v6xzXjrP2KnsnQc6z
gae6/IE/mkHAGQw4kcC0F6E9VgRDYj6Oejp1zHJ+M09pZnAtCMziTUqOSmVuDIxO
Wdmc/ggAxQM4K5fJPYl4h6fUWrJTxCzANNysxq+zIHlWaAjBfpDejYQ0XszLBRSN
StAD6M8NOXcLSwiXM9rn/CslwxWsXcX0pHPEug2SYvEtl9P/j/atnDKHGPfPB3Qr
eeToZtZj73x2AtVUrRzRFglh3cAGbY2flRWs55Si/vBtXOvIibYR4DQ3veG2A0xI
fPvfAEDf/Om9AVcm8NVW78NbnVXEwdnW1pRHai2RnQhUNAp9sdI3ywqe1Xf7ghLu
nxnXPr7a/uR4r4+UtcdK8gWd8zLpVW9MqAzEhs4dYMmEFnmM9SvesRy0wznA/3/W
QRkH2sy4c7BmLRl8Dss4Z0GeYijHs6DHSFYz7+r7K3ttGKpRPWIIL4fERwa9E6di
ArXOAHvumhkpoG402LVDGViNUGLxMJxB2y5AIMAx9o3kVBmtqJoS4QSDagSStJeP
U/OOAGV6lj1J1a2SbF6FYAOiOlyv+zvuQ5lWT4kN+OsILgTt4tYGzT0B1M/HBLX8
VE+C0bUePqXbi9gGS9I584cJd/dCW9iOnh1t1RGKjX340a5lWMDsLXUdALhI/2XI
DfTQD+PCrKEAXC9gIRbYaeGht5vli30X7xzL9AG/OC0KpB0+BtqiQmWD+DIFt8Dt
wHKrY4C5IjIgM1CtRpm8jJPEG8pjF0ZGHTf/bi1/s7B2CpAf8WKfqcU515RrzhFb
uAmHcKk+83rBXozvooSc3jcbZSUy51NA1kqF1Y9UeTiyCELKo6HlM892MwTpFOv3
7Xhx1EQF6k6FjeNPn12ZaNkXDnMpf93lUXViVhAPXjYPaFVuXmEiFU1yPlN8e5Mg
fzE3acejV++jwiRyLR04MP0UQCHV6pyLoZY02xowQLBWtc/fGOwdA90G1EPFkCU1
I1EYEktaJ/xPMrqXlqoF3Hly8yYOk0va3nR6uzA7Xm+mjGxuyB2IZJF+QhTMLAK+
UW3yqTYUVTbrsEwG7tgZMaBgNOHqgV8sif8WaLBs437dz3BLqGMIVIleDVFHNRaR
BJZWTZ+gnCANqfkejO53tcPh+XDf1acx/KkJK+6/TECK4H3cWWnC50JVyyez3uVQ
z8lWIq7KGCBZuq63Xrxvnbh/m5txZWDVFd0SxIM4BWcUzN/tEi1VwdRHoMwirAU5
vGkK0sJ+34Z1Z82nQH1V8CFTykvSVlsi6vp/QiP9T4S1Kloe8IQIDKY0d02iz9T/
Cr2mrWaFeem+zuF9VKrI+mJRrHY0u9ksOy0QDVzY7+TCMi03tZuLo4UDEt4DOIhu
SdYpGoIjVPCteKL/oeh7NeKhoAe4xNwD2n0LCRrb3vh/UjcFR3Q/d/HlgzRYkE8+
63MeoCMjPg+3EvqL9YXGLubLJztY/mguLolfWqLP9eJQ26/uv7ISBanyDWuhrAg8
rapqZ9n/yVGCI3AIOaa8NNp0apPMdVxHlGLV8kmkF8HEg7+lhdLWJfcOwU32FoWH
Ukgc9LpeEHFV8RVHQYU3KaU2wERYKBDzhdOfBw6Y6rvIx51PsiOn03Q5aFDFgiDN
jDcevyvzex/CNyS6dmagNwiQ8g9nRIh4ddVjKFbvGmKwBuQ1HrEz/uE6+WWpCvFm
2/5B2i2y5b53n0Ra+DB2/rGyQ7RpeQf23fXNGkByD1+Tm6ouuOV/Z/SxMXQhVUYW
0SlJXDOqVG1Cv3K/Ta7Zhxs3CCCQsYWhzdXNipLg+TIxCn9KIj6ebPDpiI68b4CS
0xhWkmRPyxTcn172uNEeyqS+qXZzmuR5STEuFGt+KSQEom0Z7RyfDmDJWJXAP+IU
eo8kOlCF3qAgkkEIoYOb72qRnljtOBQ+eACg21Grm0IUqbA7098sIpMESasq8E1t
l395R1LBC4DbDVv5sWEXeIwTp+Ji2FRvmBh+BZB4d+FjKIGggFYBzNq8s7mQLKo4
Q1miR0mGKcW893o4hCST38D29cRcSB4oZA94m/1PKX412dMkpCMVjpz31kXlx4MY
8tsZxmhix+4sM+NeeqJ45S7DsUu6V39gErKg2jknIT0IItvWtGllZPLBx06GRW7x
RGOQbdvIvhVABo8UkjOM93/fOvv5dG9w1tg01UrzBV/yMcE/ApT371mI9M9Whje6
GcjaW69+2VqeOpqfwp+4CuWqNbvaFPQA2PCaV75tFGOJFCKM0qy+xZR9Yt1j9zVH
uLBL3e/EREDaUXuqNhvI465cML9fL9SndvtGYxxkWvmHPnJ2BQ2DyaoI+0t5Da8Y
VahWnp7tnyHD6N3G7DdWyUvFuLCetmvyMZ4ho7NZmopYjyeZI6X3QI4Vp+gOCBgY
QZOvlquopJ4ZFL9kUcVLldJNe+ggGXyXN9rEsdJv0DsulMTQfl5DSw5i0aobfSgL
M4dbTryVDikXujZalYCIUf4qsUeTMsobb4jFJjlDK+/Xvpq7KrFt3jRXEWIDL3ZA
Ef99jx6aEmNfcaoucfYsFos8rRxfnTKSFmlgJ0q39Y7m9KNjYQay5yLoEDsUwBa1
mI4cGkrQgdZKiHcYs9arhIfVGGN+HxfsqlG4VpYOz5NzIti9gnI+nzw0P5e07FLR
DscLCV1/WFMqAiCp0EVim6IszLPDuCANxWYcjbg6Bi/cr3LTfOGqL7LT/b/htpQ7
zyA1Y27w7P+9jCyOfrYSzhrIsw0Qn4XHzvDhJHEJ0ANU4SWr+OH87Jool91dIh6T
BktkqHj1F1Qwf/iIgiG9nEv2jZ8r/+TxOPFz5nVjtQ2HSQgamjaXKAzl4cBJDB1D
f400E8NucVeo9ovJSLbR+b8mrK8Ouhjcp6qXwuPIPNq95wHsOfYMfhxCbcmFLC/S
U87GmNT4Hszs4vutPZS+kqVjp/8bG8xxAI9vaVJT2j1wcKSVbPjFIzAK+IOBQQO5
A8G2e9S+IXYPGYRH1Fv5vyT2uKhETY5ouMZFb9RXxyqVnobOakRGoRXYPRZLb8Ed
30+mZNjlCmGqZV8GjYjHFJBvovDIN+p/bymDW74ESskjmnI2Mq8Jl//jIocUekVL
KS7b5Ud4/sLib8gVTuWPW2COTIyjgH52D0Fzqsbj1qr1CkE734eDbv04F+0sbQC+
dMQSFGx77hs3vEOuztAOAkLHFxf3q+Kdcsrx4eYs3OJ6VJ0Y2d8YSyK06KT5qnhD
239r8Xz+F5u8KaCQvLKvDuDjP+g2ICJv9RFgZfEbSIn35G0e3MXUhjB4g2KFx3ij
qUspM7iwhWasSNK28uoVCCi0DX2T5sWK2RoyaJPyg4a5zUFBABp7gNUoWHgUmBPd
EdHh0JjyMw/eb/uRj3JjlFqr/bDDZGWpDm5HedZi+mHISiX1uUubPzZaTQSdrTYG
9XRbGncCfrkq8Fyf/VTp2IYuM1DplX1AIZOkIfj5aRCHQFsmOvj2csbAPIr94BFc
wBtB7KM//Y5QKb52yKDbESGTbwJptXyCyk9fr4Blwvay5OFepsdL6SXZNEMEFlrs
sujZ762L9U8I0XcY013B0mSMRFg9+MsA1PtnyWU9ElSmbXFSt5Htq/ou73Xcwn/D
IjODo9FmZL/E5d59sbCx7prpGz/Yj9lcO317vRsI/8679Z/TaMZHa0zH9lRildWi
Sn8yvhj4LjlFR1OwGbLRQmwBoSattacB89TzGtXZ1LdyqZkobfFCAlYUzaxK5gl3
9vNkV5k08rikiM77J+MjyK7lEWud+8zxlkNFLijWzqLuqd9ndlwBS/1ryrPC395W
hU2R2Z6zmj2bFeXioxBRi4pWR0n6LuDnIZfNUacuKPogF+F972163N9cqqhpvn2X
GUTaUKH9DWUoBzSz0cIqPa2xFNEoG9DnZSea/Sd0UNIMFys2T4uuCL9wArPJu6HQ
7QhRPNPYH6Ok2U8UNzCRiuLM/KGi5sBIGK5UblHJXhlwwvPOhCqQTpZL9pdqcmd+
hDRlO363e2H5sSAcvf4OWMFAsuE8nQwBxExtIrLbbcp0uRMTmThEKo6ZwhaxF0Qn
O+2r6vxvpYDWdAOBzMZJ3cjfu0a9MFDz9MhsdfHt+aMQfaPELV9KK3gurJ84+5XJ
Q3CIRRBf+3P5M2OQhn7M7xShIlNN70VqGewlZNf6czqPzLPGeQb8pJREtr964kKY
Tgdoh7U/O447Za0zQqwhSpw+A2VcuWZIUtX91RO9Dd1l05FXh8IYpS50oEqBd2jH
LuY1dZICZNZ445MiLXOq3BmrofZrZp5GiY56maiV4Jr2pucT0nyTWtnRhd0hfjdg
Q6FpTe2A/t5T1+cu/CABJGUqMBIp111+SMj0HAHj3w6WfuDDlaAoSnVCCjnazteF
ih08NFgP3AfuKfaIjX9GIVOPu+h1+2r2JCoif4joTkM+oOYwMFbBCZH7quQFfR/8
3TnCvJ11dWTIzoPh6RBoTxv4xlR+9ppCetTJJB7jJkRt1mptcxl5cSUOqKQJHpKu
FBTgJKkhYrnf9nGf07lleZbJg00A4+LmJ3Kl0hkbId9gJYT2IaESK3dXc6eR/EA9
5/S9pdjBAB5o/zVs8yWQe2x24NovbFE/Xuw8s3FbhYRfS2blcAmjpMS0h6UPOOF/
lnwPqj8eyBQTUHq0i/bmJ6SkuAF5+nK0kmWOMryiiKQY1mwFdzeGylUDxmMqT97V
v2xQ+8RvbnnjPu+JUl0QAK37mlJZEukeyL6Ag+lNukGsyZtBSvwhyW7mrJHjiVsN
ji9iw3uF/A2FN+kLANOZFvzMK79ad+6fW6wW4sra2kZV7190jUWcYg2iauqff48Q
hIQ8SnveVI7m0QJE/gjAhUSHWPDYYx63UTA++A67DePDmA/W+cjHY6JM2qdWokbi
i64K1SWtKwVeH7niBnE7rGSQtUz/oCphwBJGqE6Rb2I/2blm7BEI668e1aVrxPwm
5GMs51j0mE4/BdJ2zmMz2xBotk50ZnpLtvVw7+XwsXux0uCeu5DxNhXPzZXey9cV
NmBJ+lH8G7khX9FUEM/iGrFiU/AXNuagxiRcQyCiVdtHT7vpqBXvfyR3GjmDevbY
n+8b6ZdDEPdxeG10BQOyLZMILw24bFDHdcmLm4u9oz70kltZSt1hnGuMoHqgsuyn
83x+NetsHWO4/l3C9t0BcMgSZBJu2gxtqIvbIVgSlW6HDpBz8qOPN3ASPuMEVt6Z
GJqcTceQYFBrRB5IkoxSOHxPIwLFuUJghBKq1qOiWBFQgDw69XuBsGGDjLsRaAz3
pAL11sU+/JP3YEpTtkOD0eukrGTNACs5tT6QD+tHP/6gjAHOMfzQJ2+q/8RIKt/3
h7Wf519PcBtx52ch7KHDM0keR4gbDhC1UAloJ4YL8Wemtlt1aSP/p1SGmG06LVpo
mMwc7fM9TcwaW4x4+Yla9hkqw29kzXaChnbBYXt9FQDaChA5+Zz/LBXC/UeAJSdX
7BNqULNcL1nOj7DTJ2EtJ6Dvb1IjFpFlCe6pi6m6Y8MN0YP1l81sdREO/jgW23LO
Y8nexhsrF0mLpibW2x6PZSzozvaempi4ikbDbr6OkgIOWOjPbeDS1aEk7/EZDjih
2PDXO4fDiqJzDHgZw9Kb0h88B860PoSCw5dJuIZ6D9MywenN1sv9ToALHW3W/JLO
vOp5XuXFt4nv92+fuixexyvjdOgBG9gF5f39ghifMc4UDnOa2+4l/SGHVU2f4kcC
CpqvsjYELgP7pN4F9xwwjQFMWOIbKEe/ERBKRpyuA8OpKGkKauY/R4WkR4FsOImT
+qnveNJDPxeAGlxHsBpfwcr2okcDHK4hSCa7Z2V+s/0zcksQKglvlfJxInMcevdQ
QvVYDA0vNB4SkTuiJo8SqLo/PoSvxLqmXyEnDzVP21ffFqweDTp1NwFAbWE46aDb
7MH3MsqcrqQWfeXWt1GynrFBiBOlw3yLhiYtlPBQCvSoAa0eQs4j85tQL1TU1qmu
nb3BAp3x5BwLOJqWh4Svr80ZQ1AKYBfSN3V0B91+ldvKBCxqbPy2/shnfXpw442o
OhTkhSSWBrQ4M0AqRUWXkgd/ZbV3IsvqjgjRqEwpWood9Wf2fg3MagEZVL86vmC4
K1y65hzWpS9AXhHZZ3EFbj1FeSV0WORixeAUdKuqQ9nT2GfCEUCXvP9rZ2HL8eLZ
MvBH+qBC+qf2QzGvvUo4qPNGxz55+RlgTMhjS0y/JnHIFpbCA9zqRnLfsC+vlpa1
KVqJ3xIqtf8jQ4Y7UqhXI2V/n2Oxun38AUVWIwKjoMMfa+JWX3xIo7id/4XbfTYn
EwDhFLRPzdoEn/A9cZmwB7kdrWA4QU3jU81EfSvq7oT3fZRz2n77lGyQXml9gs6e
UIcADzjHSrikeWJoNHiXKojcLUIMTuAkyU3aPWj8c1/J+5GlNcpXMPG02nMH7XBc
dbv4sC0shWtxwnJSG+LEFmnliYFR5ZBubmYanSsH8EBgbkCp8lPF4eg6g5TnACIT
52DJy2wIFxOR4JcOybTjunk415hRHSqzT6P9zjZYUbd6FgF6paaH5pF78ZtH6NtU
XJBrBWBktdLeG62ucz8Xrl84by4wLmCAutgfqUlBcKqkVBE0WLLUHtmXoC2S6/nx
xX0RH3u49AWpFKksxebo3t5z6uP5LkQ6+3Pg5VNy5XRKbb5J7+zf5PPoxsbxpJyR
hdtNpZcLz5Wacp6ZSwkfsF0Jy8laMwqBKKTczdiZccS8wAg5dPlsnjuP/sYnEHpQ
ubyQZewJr2ymu2VYySZnvf5Eiu0stTc+OQcqwxZ50da8QkFoZNyp4T4R7BtLomlA
cYaAu9MuY78qDcml4Z68gIfLNvDHRFJ/xigjggkorsXAr+RHV7K3EAsW3AiUut5r
AcrbfxPLoelV5IIOH8aIkJeAC8drJAlabFP5V8/ES7tFvEeuJpWW1ta135tHHNLk
jd6VELRonMyZI4t2tb1jJ970Mn9J8eiQO+BPJ1aAsX7odiqj3Pm49+rjuBpb+AkJ
LEOcntIUS+CGGzeq4aD/ogibqLQfTZxz/+BFLpbZmoqU68yYEACLgSVkpy/X5Dp3
5OkajDZSHgCAGv3Tlr30iy6Lj7nPVErrObjDj5ALWljNzWETaY8+HFtFYznApPJQ
Fso184eAgSmJTfTDS77XVZzPP76W5lNRh2jcVl8JanuKG3ReiEUkFJbU/Ovr3AEO
f+fhlYKmeGxhdCDAZ9BKpuxC0QO2iBGv1y5LS/GCuFAJSslQeqlrOvkP7J0aYJsW
7qJvZl9uZtiAmwF0MA3Eh68KA+/lrMP4M8jDATYCsxuDq2tYHZSYyH9QXXsMv9tq
7po3AextCQiwg7ZORZY/OKbWDnryriNjjJOHKpBaDaC5oOJIPlhVc27UzLrq4s4g
QbGMHeVFZ9wKqW2L4alTr7t4FyD4srG5CU8V6NydC+KW/sZgWYih4YaVYeMg88n6
OMXSyDrxgmzX9ksW44NOPu4+OZijyCcifOKyjMWcs0PpiItw3DvwI1yqGU9h3gmr
op2xRwBVFAC7e0OVEW2wyQtaLqCOYwJKKF9Nm1OQaOdHDIKkqqG2eCP/5bqzKkXu
8/gpI9co95cBrE2yu6gqzwZJPKAVm/9fk1jSzadIjAlkieEcmd8xoyh1vRGhoUZi
nOv36aMzWtdlSfqvuR9yNgnuL1PqM3DGrIkOZLu+2CkIzcyIKlf5ljv3JkUFT+2d
8bEDC1qJ24h8wRDY+MD8kowrQK2lanRhnEJapHoF5XJ/n+w4UT4YdTz0rpkCjMi6
LGSGt1lIJj/gsvLm2WUnA529/iKXiUt6/rxfx2bkytLTTmSJfVwk8n472wtSnWUC
9l1q6F66iNnRdTMMb5FM7hV1HB37G5SaMWN+qQuvbx62px9FXKTsxRxu15AQXnCg
GFgaDUgeRq2p6dV6J/dfaoOy/jFBasQpk+LcML16VnmGxIuNzUNHM454AA0A7DnE
sLImQ5skxPfseUCEaOu+k6ieWByW0HUk/uzRloXdNPsoQO8BU4VxpAYJWUWCx7OM
Yw6bbI77QWueyTUjqz7VwcPYEUfFgN82IG0d53AZo1Tu+/EKQlqa8ItpcC7AatJz
2pZjmB+SbgG/ND09BrIkzh92Nuttkm2tCCuT53luETB3o+MEMXY+zzQOHHrA+d5H
xFAvE1h+pBG7Xpbmlp+aCrwS1LOchJ72CzoDSAFHncF/DZFTn9ncmlaeoWAoGYMb
LPFi4EYxwiqCsog47D7XSlWLpOQjneF7jG2QFiK6CEAzKKAy97oNO/XwWmHXgj7Y
dfVOOWoeClEvAYQP4bddKNob6bQIaPG+DL8xoKS+1W65oAjg/0UgxQGCCIxrH2tw
j2xogkEZvCpA4cqQfgLoegepcd3RKGjkLDfrSbNLsJcrlyteRPpEWT2bXCAHgakX
pPAzTRwKtJGSqM/1H1zKlz/OL2R87rYuPLVLh3XlfAada7MG6jhqAcTClHsLigF+
k/B5ggd9RHi/UJGURzXsZ9wtA2UUrteUWuhPLh+7vZYfxhWytW/jnQx25ur/5pwy
b40sI5roFvSctpPHA5FdB3SElQB7i77js6rA1Cx4TaDAf+pERhhcjUu0QSe5Yjy8
xm4nKoED+AGccugLVd3YktIFLfcRPOzwyGcsSaGqFA9KL/R3KS1MMqvb9OcQoP8C
a1YK6qO/tbaelUnTYot1HC/IfXJ6CtNtBp/b2Ammv3wj90bPAD3kjKkelQnBKI/v
yB07pyX9jWEGBd/KCmVtGebfLLlRC9eikkGpcxyN5VbpHq8qH4p4YWeVp5z3BMQg
BxCOENNB6NThhkn38XAN3hGgOJAkYEGvi7k4ceTwaiFvxfXBb0MgalH/RqN2hYB2
G/x8Z36Qod1VY0jdKBnk8/42dyW75EnUtmM808Ta5BpeoERJhLqzVyhMjteZu+BM
vziECzIDzhGYOzEe89nvfToBUo7lfHPGHGdkc5zWtdh5Sryd3Oy1ujjln6h712uW
T7Jv2IrndjtcSo+b3hgndUvMc5B2hT4hafSY9C9WTxhLYbYfD4oLDUB7Fl9e9GqR
e0BFVHxXTpeN4FPZC2sUV24U3a6ymbiaWdOltwIWKvi9RoJYlPZBAu83O85LZSPZ
+YkhqMgr6eDJPAFuJWu9Q7Y5/qyCbKqI55WrMEL5zYbNawXwlr3XsqrPtEjKlzl9
6OtN9XPLPnEr5FkB3ppUdaIzDesE+qCIDo8WmpEBMlXHCicWH0CpMOXkPTwwJFPz
nWgUPIk69vmIuCi8Wzxi9KTIEtmcrK3LGW9l7P3ah5APckm53mNtj934Lteiz5Ac
0v6jQMxYKw3/vUcJ75bChN8dHu1DA7ImBjp8gT1r5yGnc/wBOzpw4nusTGOGL/+4
vP0EP25CnbtrVK2wptLL3Zfkj5Cy93JVoKCcRbzl7dH6DTtvbVDj7aOWmhGU1+OX
SvWbIsMQZa/OWKy9HZRHP2ZmE/f88x8Uo4ZmII8cAil/a4a6OeX8VBikvRzhtAlo
mlwPcdikM7j8akS3VO03icej8tJf8818Ng9x4DUuP/9uiCOYLKKrQVQVoDArjff2
2586OqMbQUmraZyc39emZA6bdUHRfx1qwjjejyJofK9LaY9lVu7brqubg12/hy6h
qGs9Sci4kTl8sbGQjlCv8riw1xsK2Tp+8mA4AkOEuYidiKeQuFvaJF91NotcUwAB
Mjf50YIBzDJgZ+ZfxTofSxCvWtsYWoiiJOWWYRFyQjrFa0vkBtdqFycJuL+s9yIz
arHYRj4bpPAVZ3RKQFS72iC2XuNGQ2yJDeJZo4AqQTvA0bsCnJ3s3phl6bVbYIA1
QCZH9xJspDJT8UGk+s20vbh5RGk2ePqXgmb8XAm7anqdcZLq07ZoN3oUsFafGV5/
/E02uo663QLuO80Y0rZwVhj4REcqJYjwfbzfRgMpVKCI9GqvY6gtMbxifb+TbKeE
pRQWSF2TssFu+ukNhBZ5cK3BsbQIVqcH2/9nIwj5Ves+Wju+1lJw3v6WF1Zbp1x7
MS+M9O8vomhZ6TMzan8KDlAq6xaPBh5LUptmDwAg7sg8ImLvJGv0FxybRBwON8vL
Q2fNj8vr8w7kxcTe2VmgK17OeMx1A1FvADekyO7RyaQ4m9DqHR2LcadQPQOdWqsW
z7mGE+QcIj43fCWxvYPYqJbefhtGkOo1dU1suwhhcOMGXL4ejvRr9I3zRVWznoYs
Cr6kWS9dXo96KU7nUVxwfxRT1tWO0P+uY/vpqNBXUJUrS8dLVFNq2l3WosXYomuH
3s4QQ1Mj9tPpbuosaSP9dSpnb45JX9TdBKYipjboUbFwtQ0xEi1GJvaYdgwhYB4R
VupczInUy0+NatsaKrmESc1e1QtfPBT8XzG82FBpQNVHthyg8N20IZ/FDSug2CSc
5uTLpC0pfU/XMcKDzRbcZNIDBLFb65xAkk4QNluT2SnlsE6DsLf3DxTVB92+zhBG
eWWVaE8kK3i0Cp+cApphy9TO5ekTt8YUL5sbLkgFPqlteN1hMNN6v8xQ+7VHYvit
YkHt4mW4R8ieCSWPkmeBKMaywp2vLSdngn2ZIQPWa8r9XnisuIaHA93UPur+bL8D
VNzWmvclUMpdCYSBX+pXWZjK41r+TsKoA0DAwFGmNqFHJt38MSRrh+ZEeKUqiCHr
UjsupjP5kwLzuWa3qepIT3xywZPodSPx0UlJA3ykedhVpHoMdF7CStMrq3SlutOD
raSVA1UFqN1cE2ZOusUyteEF+jpK6884AGKWHbyO2gxWrzVwmhrJLBVUcUkGtmWg
vJ5xm2ueYNOsw5JgWTvFbVVrf7GXo+8ktqocSvTsDpX5CaYe8DvIq6oxqECp5TzY
7IY8C5jRIOkgazkI/3oyxonvzMIfc1hAGkvf4X8GoDCxWXlWaA4NcnyeyRuVfIUm
fnGYQBlaSEvWqMcUyvac8YzpfYV4pSeo2MgNk5b45Pv2vQfopETHPiQSaA5OMHh/
X4DYTV5ZTO6gM18MJEMMHZkmg2nV7aPajcjL8R46gT/TYi2cZbzIruDUH4sdCGjc
M9WVfrIIPWvKVzO4UmZQK5xMnHlCjqtiPAD7b2YkDWuzWOCPpYpFsewpb5KqoxyV
/HBDOUu1Y7psbKFoX2BAg6cBTkuLRJ5GUaVqsbxSKT+XRzxoPSdqBkS6WkZaN9p7
xpIXPwyFm1XT98K9hnKCk3gW/6vL5MJiCTXBpeYujMUZ5+oLijgln7zz4KncQwDJ
QiH7Hb/x6DzksVmC4E5rOwdAuVXN12VJIqBclZSST2ZabQvbjoinpVWztUsl18ba
bX8l/r8W2W+tvnsVLHEQOFT7+TjT4FnKqo0rHxEwZTP1piM1a7WqZje4ACMfPFRs
Zj9jc1SORTZgGHDIKZFRsJQ4lmQj4zOM0+jBns4h6D+AKNo0+GJe3ld+f7eahBjM
I+dmNStO+V7BwPjGA6ih7lOdvsmCEybubtQn5ZUBDBBHhinMZo1BmhsQL7eH9HOS
F+IfiSWUBndMUJTxidTYbFfKEBb+/L41VD5zrUnrwYcLV4OhajoAQhVn6SIQDPtb
dMC7sHhfl7UoXPVLJyYgkLLdGkWLjXqxU6fnLfoC1OQ3MmLvrK1X9jZF4sbMLDwp
g7CiPZTa6lAv0FOYP75iNym0+5UcNlCLgictBOXgw9DrawLEcfOurnJU7coS9hv2
lYi7ir55PrULHLEixontg3FXtDXTYSeq0nwAATkB7gaoIVVKKK0m8kPhRecZJe/b
kHD4WqUwTaOLb2Z7J8vOwPlOFCFi2Bb1zxDtv/qPFqfmrBiIs+olswR6ZdGHEqht
/aK91zfHdnSsHhmuRseWEUsY0inqrl6IE5swwpwQGivOEVu2dnNTpvWgpeHhZd8K
yiyDAcxbQHybNboDSo9uGf0DWyv/3z6kgXTLnaMb0eJ75uZV3WMpIz8bByghBT2G
igHauN74akkBBNq9bHtxEpaeu+Ho9mt/LVfoWmHWzfUNJ3eJm91bP7B/zTg8C9MF
1VPLpCjfQW3Jm7DVeSNRRQ9nCEUKJx1K9UidWwWLEIV1vu3IWCjxqtb0QJzEcqhM
lKjQlo+wRohBwv/tH97R/ziEqw0lJ3zmQnYIXbraJj8RMV1uXa8gRFgPCR7jfIWw
rlbCjEsDPvrm7Adm04WJK0nojnwOJVzRFJ7YnAl5mMZtuQvkxEpeWm7li7qDytAE
rRvS2/6PE9YpXfvIPbFS094NXeno5I/es0pqp87lodKBOAYqL867wazhZiAqgHzD
Yln5jl7mDEEbAnpgu51fjaUKTsYP85QbJCuXSMZOpIXsNgDPiQ2wRVcLO6aJm/8M
7jvXqAzR3tS3Tw4jXS4s+OREDL+Xs6WQoZiBIezHv28RevNONM1Up4wBIjO2Rhc5
kvJ1/Yq7F+aDlECoqnO1JDR/ANEQvAbZvgkUceZ58TIk3mb3xKu8PqCNYxHKfIRd
2Xr/ge4uAyyLegnMsR/RBIKfZ/6L0pfVA3RI6O6MSMG5/DazCiJw9PjyDRD1UwVK
6bKvGixS3zKzf4/k07ED0wrYg78n+ZpRBMmYP0hbRLBp1FOEqfg8mpt88yEAnxK0
lCgS2hCJxc00yaj5okpINvNDO/V4OQZhzvODohu+qs7XTA0waN6Yn8Fg22iDhDJp
mbx6BSNeY6w/Lvp8lBUNOCPxdjwll1XRYQz3AnaDb8n+ca37F09Kml8M1S1gauCf
i5+xSFvvJe+2z6rnoqnQowooQZVBn+JgTxzsmdnd4EZrWWcpYQFjkcqZS4UJnOHk
0ePH4A3Ja3zfPzvf2wHzQUJjGQF2UZqfa54hAko5W1v0e9MqkSoGqycUjC8vBrAN
Og99AuhAuYq4eFpOtMAyAOjnyOLEgOIY4y9A6ymw0bneIr9fgGVm/5kEVzwV0WN9
5j1CPL3JLKS3lclhoNpuAfR+grZ3wknSns7EJtk9tAZE0JZXVNwnKHxIT3lAxish
nlzWJm0UpeVd7fz+VTC+K4D8C7dro/vZn3d67qB4RrL4FpvXxUreaBV2J5E4iRgI
2rS/jTnSepPa1ngA/JsxkeXpFLEC/C2JMTN0sk7MALbq5WAdf34s25q4BO9t6/IY
E5ejyPGPM2w0BHhz4hBuQjdOYPughnT7pnRy7RVbXd1a13U9qRSVrPNja3BzHw8d
mUMFyXQgTA8FZxNawDwE5fxrCEf+NDPOitbUlt35xVeVPnogDxTT6Km4P47nTJCQ
ei5gttUzktNzDYXIBouxWd4BC+L3T2mK6HbJsgSGXg6m5VjmNDS67/zvYj8L6I7K
G5jmeOdoC5186ixM+L9O3BbUeZGcs7PJxmwST9xnW04ikgQVaSQKKRUgyzV1IcM6
mn8x6QaeAnpDx9WoNQQyKI/hqUJ7pkxAJ794UJOsfss9wTQ7KCY4qzW2Nw/ood2q
yKHQs8OHURvPfYKL6eGuq1eOKXK8QfC35H9jGWG+OFAP0IBY+YMePAWM3So0ZcSq
Yxf2L9dm7M3w4DM+BNy/hUG2hKjNyEvZg3A8e6gwok773XWrUG42D0OIUoG9kXC8
W4bI1kgfkPmS4z9/f0hede48UqYKBX/4xrB+vHAxO+hclouU0YBNEzvSy3qUnBCI
+zZZSUkfbep1/ee297mU7d45xiq29gEvK4VDkf9Iljem5gnZb0SdpCzkhJX+lR0u
TG54JwqsBhsHua9ddrtEukXiBygFLheccGlbj1FydOeXj0jYFv730AXYYzlRNMDc
YTPBqW7zzpZCYPY6Khp4BIj7hGpK3kScBom/oisVnN0ctxFZGhsbZkrjMZ70FnoK
fC/FrjAPNxOxIA6RBIBQDuzosouYwyI2bcQ3vPiG5UITkbi2olgPovN29p7ljtoD
OoELADLKJq1Qub3VWvB/rz3R4x5U1GPLAwGRzol752p2K8LCzXvndNCfMYlQc37m
AVVCpJWIijFUZw30i9/EuU8+TsL/opuJkLronXuRxEzOfY0xcagtybmTGix4T7VI
0HwK6bxXJSh/bN9ES25NuVNgSTo7fN0Qp2vzdw74KRWJp51JfIwETNcHmbVxgy3R
u7hyGdxEjIHQTA3vOMYcT0YznFLxyOxYachtgfNRrSYme42e2zugCGEFzFbYT9Xb
+gSFn7soqGY8evL3OGHosa/sgmv3QH8sEC47gvnkfbOAblwLZ677/ZXw2T/Z1L/3
0Y2cpR6XbZCTzorJgwIyKaollYryDas3em2L7EUrqzt6BLU8DPFrl9ca/MKPiOEF
dAIQ5uTGkRN9EtMl6+JYjC6p+LyzbYhkcWYFjqO00Bv6sglsBOJvYaoAnMp4k88E
8gKv/YeL5+ISYUE7vMG1Cb9bxUIKjQL9wtxneJ/XO3TlCkNpxi9BcsESPnPozPrg
MYMAV9ec9D/Twwv+7n8Y8vSCDj2SukfxwfPpX6TYKvNMB9KEA2YEoNMLHZSL/7cQ
AEvzQ0wmSyL94rID1lC2FniJMnpQxWo4v3Rv6iAuPfunx2DNecqgC809xs2RSMWB
twwpKBclugWEWL+LMRjP+vO3V51UgO6H8qi/O4t0mnf3TX3kiCnj3hd40gDj8PIX
LEuYcH902vYnAQ5ogus8yDfnxRQK8s0Vg/19/L3cgWrTUyl312B9tOpvlLre/N5y
nExY0JV+9xcd3VHugwzIxXpkCe4/bEbbe+9VneDH43dTQqiY3txxy5PfswvfS7EZ
5CHuDSifAHb7ClZEvDhUgVlJTcIuhhtEHtYgxow03Dko6DQP9Tl3F3Y/WLBwhBfe
s75/KVL7GzYWdmtUhhM3y0X9VpvWM2v5LYGpxb6sctaHArjMwX0ckCn0H3lUp+z8
ezagRcIsKZzL+nrp5n1fJDQ0+hjnR/WVUTk4Xi3tBd7+6T+WvfVbGPVRZNF/6daU
ynFIe50NwRHnM4Ie9yv1dJDzassNyqXifuR7yOofkvwIJ9EvuDxAHtImHXIOSxfz
EAPHS5Cok9DgwBuLnJ7r6Qz254+W/a3widaZJMBAsKmWqrkXNXymIsa0dfDF1W7R
iCEQqRb4oeKxOvdJn5fVt90zSrzrHRoFFARNDo1eZfQYS+HevDYtd5G74fSUWtvv
Ddf+Ch7zOW8edTDbTGB1n2gC/7VaNr6+H0/rVUsAFjOl4miF6ChTSnozR/aOu86h
8BF3lfvVYCKexvHIIqOH4BSbo4mNe7CsnhR4+N/S+zHQeP4oyX9hFEJbgsN5O7Pv
6J7ugE1Kf9vB82KCRYSH/XGo9LkUSHhbgDeOiwcW79yJOIlcgmszELS0ImgdgbpI
RswL/ymAKowpzflyKwXGj1RW2bYMLl8UboQpQG2SyYM7pNKHn25P1v+g1HATtktJ
/ZyJ/maaHD44HWPFU3bgJfZazYTr6SuCz3CmVG2V1xL8lWCULU67U8zcIK3BhvSe
5xlJiTmRadnsWAvDZhbcW1GkDAPTWf35wt8lcbQfN2Hm8F1pelxrAjDO6zGRBUbk
RDF7bminhuFq2BTPtxvl+krAykwK6pgpSv1KGr8Dvdt6i0tUXMjoUT5JTtADKYlB
wYDXEkitAzeTFYYOvQJBR9LF5bd2TwZcKyuhFfKvhLpW7nWEzqRRDScgwWC2daWI
EIiRCdVzX7peUP3lHkrZ62DXug2j59Hp0EcXdsPE3A5b+vHgH2t+bG9WlC30ient
COFNlajMtnleAq7g+Yb2puPObfLiggX9PkKVrhfZwJ9z5s1FPinbMsCfY+lnKPOt
+4u6uO65q35Rx3iaXN0mnECseKS2dhQUz8EWCYoyxorgWsbmb1K0wKrzAEcLgU08
sFG+aytfIMal0/PHE9Pxm+v0cIorSViP2prH41yasyP2UslfCEA9CoXkEDjCVEhF
WqEynDtbH057EsD0ysCTA3/PbllONGmoTVU6Okv+Y1jCW9MduE00VEiBbcnRVLbt
0TUuutKepOsSAf7PFib8GPu7R/1b7BrlVB6EkRgo+/NKyNY42URhVtdttdooYrZV
vVqeVXHXS6pnLxhUjRMlqm3lE+EibDvboDmIAEq97yDQ0+vAx1XkifXQAwbQ2u7n
9Mg7nKYug3aqF6Mr9jcRHIuiIhpTyEgJSgZA+1/+dLj7hcHw/6jazwl2hNkdms3m
OHL1xZX4GcBZ7w/vYL0M118/CY8icr4VAyD0UheMnPk9vuzgrP9VVVw2WlNlswIW
PGnN9zjR2T/d7PRwIIDL/+IZnSfZg3Dw3IY3ljN6trA1tbYt49PUQSB3TwKJXE5o
ZzcoQLyT/zhWObs0g1e3QJB9VnNG0h1qJrj72YNkkhQXbq2NJ5+PfxnuNVrBYvQE
RVL8cLEgC9LRjCfNmACRWXfCVznXCgulpyQ2mti85Vu//wiEx3jZNhfLy2iXh7kt
3I/20BYRINMWDYVqnA7EPuhfsHJr1voj0Sc3K47to0BVQ8ELy+XDvX8J2Vp4QtoX
FziCs3QFy0pJObgCvjuSELn7n9TuHurAeZInvx9/1l/zPsf3DxUT7HUS7z7jeefm
5eSrM49MKoiHMNRM9iQ5DU+xEu4OIDBtMzIItkHp2yd/lLBlM2G6yafut9gtVEAU
QWwTP7IAlLir/nt7VGp5P0L0fqyws/uyV26MFvHD8YuxCccesXgqqktg3TEqf3Kh
3jNca1G6RxNFFRdKkWRoY24xCuKhR2rzJs38Hs9GPUMMkNf16jaoPwYH44zYz038
yEbcMmdNvFNqON24uWo4AQkx3jpZvG9nIjRstJ/Zo+beF7bGLD0EHN5h+fv+0gsM
NUQsKtCO4CuN5CpqGjxWO12997XdThvtmZSRCi4AcZGtRyxsMzyNGnc1fLSMEDr1
9dStkeKUk2EZFL0B0HqO1U5GXYzlWufJITZ/S2Kryckc6eyNyoZooKxvkT7JZp65
AXVodSgcuWEVtG1R/JcWrXLFIjbbDz/5fAQnA9HKK3XAaCh7HGYWPloJoO0JG6By
Pf10ZElbGLBMngv4WiYIHwFyPVV5zeyoEo9gdEMaxpdaKCrvbFGQsc1CiP0gfWAh
lRXIiMQrzydO6MQUtal3UhBVyHL+6LsMdh8k4Gsps7ro1+syrRq1kZkHQ02R90vZ
Rpr0EDi1JARV9c17vwbi46vuPrzruVg7uN+PDJG1anST291BH8SBC/+hdn77jWfk
OIp4RocGl6iH5kmNrDosB5twR5Z+vz6MPo9RD73Hpp3j0niRtvx2BXSAEJifP8ZD
M1Zc1t62oFisiQaKK+JtZ1QvZA9YUnXFUwtBl03SFM1XtANDdsPcZy/r+GKYpWnw
rXDIiCKSpU1HUMRVNECKkh0evnVkNd2hwTsxcKmCKrldnL06rHifofdQgQg65IRM
vZtRPKdvPlyQ1Yt8NYhGacMAWMbYTkveNxLkmip4WBW5n6Rr/RJHMdNj7M5L80fJ
kySFP6RbjkeKU2d0gnpWrMjQxf9kBLMnAQjJtk/e3X5Ny8RMwf/CVTYrkl2GYIkL
/g1l86MpldCgD712D6/pU8RVhyb7crStIDUEoGiCoB+yt9OsbD1uETxSc41uk/Cd
7iBs1Hm0AhIq8Jrlu7o8Zh1qFCUnJcVRgxS2HY297Mzhn2mpHv8zrWASEv3rhOnt
1rxVb0ui8194yBMYnWQY7F7z0FGkG8K/8OJU9/NQY8RQPzjT8T/Xykw+5yprDc10
HfEmXZ7EGuEQsNPds3TwSfNfAykpDtWRltPGE4PNR7O50kRiGE8itIajpO/+1+BW
dp68/c6ex51P3mMyYEtePwFlnOCZSJriMNe662nuo8hg7YLBoQqLnbg02zQ2gII9
AuDM4T/GRsxvASGDEc7RWcRhkMfil0LJkV3fW7iF6v5hff69iWvC7jusdTxpqNkp
alTZ9RD/fWcdxqJT1k+AF2mvlT048FxoSgkz+oYmx08AAuyXb/DwGAXTMuae1kdg
f5jqC+HperxGeTjm3yK3YEXey6+ZVO3xGEJQgDVrBk3oFgXTSIlah52HVuVHuDha
3A0qGivFbuMoRXyCRCadob+IZji3uvHY1zx9A4phdtYGw/zOW24J5nEU+RwLFVZr
CrF+PjVJIqV3zwVtU/bSleame6KltugFUebnHtIHQIOjzWl/FvdfvqZiToezveRV
cL5YJVMQ20ZCNYRk+RvCmoPPHHqeJKJ/HQAAbynAom9QFJY9uVPQaulFOlcIXuD0
xv5U2EyfNi/e3uz2gWDL/LZ9lYhtCMeYLC0bCJ35ry0L7q0Ch6B6H4I6GHljlCdE
ogb2ln9+aRtrQ8wPvWLSAzE4nokRe4CmgJfGz2eXOA22TRUUj6vAJ4Rn9tNF5bMW
O5wlypKic07SREXyZLJef3/bXT5g22SbT1A0aILWWMIi9S22JRk+6pIfCaysE7HL
KdkCNyo2d9hGokJHpkaQeTN2U1UGU2REFJgQGHvsibU5KeOQYFbn1GuUlqISPyfE
rSjYKlxxOQnAKxwVAn1T7+dwEWS6tXMuRwcQtfHLrzGMexrCoxpkccx/jHtZ+4Z3
pQWM9DXiqHSgYSsELWAIb+eLK0dGJXLO6vaDlm5CKaYlaSTtqirqEzxKuyGjhrXp
0dY3ev8QAJ/c0/TnOqLQQukWdJou+UuaPlRpx+5lBwEN5A6RWzZhFarShWs/5sIE
H7mGvlvMIw8jDBIF3V4AsNKa1XQGbkeUsNlOz9O6fVa3ABGtt8BZJ06uLjonITBO
CDkp+crXkzwNnERrq1eZ4K8NmD0ipgy/p86Jqro7GKeASzHQCvNNo6W36TYPU117
uUT/LcJTLn0qJwMJAqc7iv7BpYXit+f1VWTBVraEoPfkK5K6eifkY8tEty0kc5h0
JldbZrdOhBMttZxc2uojfTO86AYTzmaXjrvLQjme/RZ/aUrKmoveWNdFjvgx61zW
cCGkMisw45ON60gznnzCR64QByQpr0wOPY8RsNd6TUhRXy8PidYTOhQjH8c9xDEf
0qjTq5nHY02P1+AGHnhJrJjlZIU5wiq68W+K3mfC/HpAdhjYgAXWRZ5VkYMlFWQj
ZAxNlh7Vy37vTKSiNWfEzVsH4meuQn01jt1Md/a8toLmhiheVxXgfOl3BwefU+P1
aI7DW/AfD4E4M7/+cmKVmWHDK6wIi/+TurMA245smMFk7JOX36NZJGLCC7pCaa3K
0sbeU+cZ35W6aNqFXRRKgZlwgPOJx6JkUwiggJ0/oEVHdXzZWcVROMv9YcxP9oVI
ORvnrISt8iPZhSZTrR547IdKeIVtbRE7YQTSx9jtlg3xUFb1kWKVA/QLhu8HY6hY
QggqoVx4bcPEwp9YaD6vpW1whwNS1yVyB+OxoXxUYko+I5WFVgD3W4/gnEWZC+oT
IDynZM2L88U+H5P4ZFDrhR7wE4aCi6ppJqdpsobVyD0eLKm7TF0htjMwFr8Z1krI
jWlCEWmDxSAupLtouaROlDZhDKqc90MMu7dUItAJ9slE1d6JZZEvqHlGSbB5grO1
qTq9KAC6UIaD92YbReMRrj+UIX6IHyJx/Ce5pdLdv0+evwMbhU4M5l0653w5DJ10
qHhjrQ2cEg5t0Or0q8KvzEftheF2SV+Bbl5V3GMf/6s2uS7wtzlsSdXcHzCAP04c
kdmlxup1AFtBR6mrlL9yJISv7QklQU1ADkzvncsVERV8+PXNvhfMI2nzT71HEzBZ
dH+84D0pfKwgZhVpAWg5BBmm16hfyTETZyUoUX1gcGlo/uzzumHfYFXdVUQwzv2l
j/L+YG6i95U2US7CIA18KQWMZkcLRnSzFRzUEq5RyPYOvPKogBEBSblBxibkScCd
ekQP6h6amhM1YPUpNA58kXaPgg+nYvsHmxT+t9gnPuCBQvJ11pWxUehmme02FFBo
jwOgpwPxKbkvjOenoaFVjZKgH9qr6QuJoDA2fUYmhS9cKg+k12hZ6OlkrKYuaZPY
Y6NlJYcd9AF09SPztdW9UugGr+leI+xkLondUyx2T3hgq8w2kv/13GFkz7wpCC0U
eXZJPraH1KNXsRyBS8s5cQxMDDa43+ElcmfMgYXaovlLRZM3Lb1Ca529gYK0OhDm
j6nZFf1GzabhMaLb1N0bECJBeG44xZTwlAM7SkSMwc4QfKI5hFTD6Qs97lotvlbI
i9xFT3v7DRWSylBBpysk9XtirHhhG6r4rzRJVEM/z7AoVfvNKt6NQVGfHUWOmImr
tQH3twvntOlZiK46B70TqDPA2YZG/Cxh0g0dORSDTbVHQELeKfB4fbiZFHJe9vnY
fy4DNb9KaxIJgFiOTXt1q436jYdoKraEFaKUQy6i79/4uT4p4b0XzFeYb8cMOPax
PhVVK9IlgZJ0bsr3fELIwiCDH5qUZk1R1gvS34CqaEFP1MsrbGtbfJhgxm7MoUWI
4G8GWRsBo3AkchZADGkcnprNAOjRmJq2tLOJZnk2ydsQV9A1k46fKYJYE7Rx38JG
pMvOwWUkvOBgjvIYjRzk/NYtLGf3Io+KIu65Pmssp9IqUJ4X26IAeQrIEBBRmOS5
o0VNHJtbZvAHcT8DHdBY2XWBuD/XnYMbLTDJDoYV2kjs5cZ8HPFEOcwEGO5BbfBQ
BRIV7O7Gl3GJyx10Cg5Wg31zsWXmrIN7NVMjQ0CF0slb8NMrRtX9xBXUlAkv3seg
u/QPtyGb2M2U7ff3QzXEArCen6HrZrtzirPAYgPaTcG9Fbe0WNPS1nc8kh3aE5Gt
Mh6FPkcf0/Ba6OIPcOG26JPEdWYsyuZSX7FhODTXv/dLc3/oZXUh3X74X/VvkmeU
cYPtTq9nO7Mq4gubQiPhakzKLJyoO6jc5rlVf4/5CbPgCNCdJDAMUwJUPF4FaFU/
XXrrLUZ7TGYN9nA+mlpaasgAXQVE1soZzEz6QZeH3ri7lFIcUu1ynSd4dD/QQo6s
wzVGght0LSCzZnMC+J8fGHkYUj1M67XXN8tXtAK4fsoDIONS9hyneSxM2RaydChQ
EmXQ78gCQ3R/XvLn2kfHXQVy9j9aENBUHIq6DwwvCVYbOgObgHLJQSkFmjzLyka2
PNjy+lzrdBFrRudV4L9vGt19ovoCfBv+EbjzsOtKNumo4+oH43KTKgYkq0LPBE07
/XRJKkR6HhbzUdy8y0RQdi4My89JhUvz3WLUHtMiUAg/lsKM8p0sMONjYl0AtFbQ
pV+ueN7VOVyT4BZFd1e8GCC8pEuJDdBDTBg1qAZ2lg2GACvBURte9YehleP0GIka
St8A2m3yI6N9g6WKa14u1tfrmiJYc5V5ZVg4c+ZbwtGtQknK/RoIONvJAYto0bJ6
eM4uWkpiaOu9HKzTAs3Ck26VAtR8Jiw2LjBXilXZRqnyGKyxY1lT1ovOANGrN+Zu
M4T6+tuXUdnOzJABTYehsYCdSRlBb8eUFZiUesfBd5+TBjkSVY6G6o+ulpEhg8fk
H5ylCYS5vsf06UbFQitAdM2hfYIGmLJ4aRSM+3Um+TennejWJntovlawS4Z1nqJp
Ue0coS2o4HaBr7vGWJ73n/UqRT6P7EL/UhZVomwCA+Y5nn9yY9KKyG4LdJ9rBB5J
PRUpNCwPY3X6paI7SY5zFELyz5Pa7CYjl0lPfOVXpar2vR6ZaK5X8O4enpvPo7Do
EzIK7yjMCt/qZASPZ2vvd2W0EQDa3eA5cS2khtLM4/1z3CWoqCqsGTPW0dB+auHL
HVpwPrxr85MT0jidNqn9GZWce18pgCVV5DcQ1JMLpQRL9TaVXnHOs+jPagshgmQ+
YgoQ9NULeFfjZJEJbOYGqWpROw9JqD/xxq4aL7crXb6d2biKQsb25eQpSsStbKUN
9a6oigR4p7YY6H4sBGtIE3MUxXCbkMgaH4dxW+0kS+ut1hpLfKyVroFrhCbSQZQF
HgfdO2Jd8xjHlCQ9V0ba2C4YeS1mxlNMOqNl85LqYBQF08UMbvj/wUyuSNmf3geW
BRWQfcXhQsIEK3cVGJOSV5M6B3RDzn/HuSMbqWNPKpJTk01CiplKChyzD/HZYmMX
k1EmxkTpETJWf8Qk5/0TS3f6vZi9MSdJLEtrSfiWRYS3a448u04ZYKGv1TxobHBb
attDxx1N/XZIQcbyCRYDcDl2zSDLhLY/3TShI8DePaS5SoMpO/3Rf1+hhls83Pwz
5s3O5prIH3vqm5SZOI1ec42KztVcVxzLhN0HkzjkL/uu45SCiDGJgtVhZptnhv4b
dNcvIr3t0a47M+SEXgEHBL6uEbA/tREX1OwIaNuUD44BY9aI3HV8JXJBptFOvuHB
l5EY2ylsNjxVB7SfZj0qaql+3JLJTuQDwxC7UsuYAC7o3eyiiVOO6X7g6StjU1G8
AVCCRhTGhhvPJFDvzOogtg/hzTp+uOk7+uxDwSsMIf9fMcQ+8NvZZNWPmJuqNkMg
m7B5O1HJ5HIsnVAPb9IjAeJfLccSjERfY3eS0IGiutEhDSRKAFiQtCW0v/2v5ey9
8Fb1rPisiC8ZICmgKfQjRV8NvbKb4RRiDtuR4F/WkffQ68oCiXp31syvi979FyxU
r40WjPpDES+ulV5LP8ZzhbNO1Kj5ayFdwX+epIMg5DmLSeFu2XPr1tF+SIiPhslZ
9S9fbJJXl9aZDy64soQjKvY0nmLgwmdYygNhq7jDnYpSocHpkpxLYSJUHnWi9BIw
CsNTkQruIMInPX7p1lldTSxnfQe7cXX2ezXT36luWEUwhRFUuuelQ3EPvtqVvL5F
pSY7rBTfZeu5eKshQI8WK4SYT8Z2VPejK4XHf+RmKas057h/AkTgq9ukcXm9unSh
7mkCx0pGQgw/FUPJNKnPPEiGYN7qo8QJ/9KXVj/M6VIr0Iz0JXSJm6ZeK7udMAYm
MfHk0st9CL/3//yI+QNIaZqgVpZ1QOYj4f2JWlG8jUdOhokXyPt31EVboNFDcEwD
GNCKu87EPlkRP5i5FzMDUeEiPIQKuA2ONXsr7b5lClZj2x0aw2SX+mLbCqMJkGL7
rS2WIxDkgvyHrTIvavViX8PozcEKvpCrHk8Exp2FZqOx0Hg6rtTGijDROy5LVXtU
qwlIpdQ9yLv9ob3XQl9cpHVP7MGgHXuDXk+FK2zKijvATxM/tAe8nvrNsrB42Dpm
di8P8SOMnhGahIMDlkJWDrBxaurTBU7tBF0WTtQNP7pJhcTuzBTRsbGWjAeG2dxJ
PSE64VoREzeYCmOTIZEc+CpoOarM7HeTg4rpKPPausioIFBh3KJnv37rNo+/sYT1
o5ZZgu5Q27VQBkjFU4g4X5S30WElKg0/Xk1WgzqhDQDUVsC56llafPoa/Qj3Zmf/
kOScHbgzIVeKx3Ecf9OciUN5lfC5b1vUKCIOpbHLsxxYKzdHaV5H+5vtgkpKgYSo
H5SsL792tDjXTAP3AGj6qqLPaNw8adDC3RyKouQ/ug7irhIWVop02AquLy+lBNuW
hjekO1+MycWT5ewVChoKJgR7ysSBAXQWXfGOsf7FmztN2+HzZXVlv00iJRLDAXbt
rHIEqbkqfmWXEPR9zrw4JoQu0H9V3u8SNYZwCvCol/CsKXl/1uvqTRx6+gc6+jAG
vOjOy5r/HrXZkLvqdv3qdYrVw/7zsZURgH+wnhC+CryhMeyvZRIwf9rpQvoPu6kf
9nUy+le1fv6xWNYIEcEvvH/dVDlI2Hs/i+lAM24G8UU0RuZibt5RaDq0g9kE8tAk
Girz8J9sEvGRFLHrAx6+5A3e2t7IAojrjl3qYYnxnX3lqxJQVvb7h32tJD5dmLjJ
9XmUgaby41bwzAYglL5o+H20yW13cchNYhZQB5LTQgYoTHU3iDG71gwOU15ld68I
sJNpsAQ6FAHsvFciImV+ky0W0GI6r5Ilaab6zMP2hWj0hCrp9MmTDA9Vt2Srd0xI
h72b+e/StCNp6wf6woGzb0Q+tWtEXl0Z25Ftjve1eGK6u97eMfGU/jTiqO5lZBQA
FGgECrb/hYIGqI926duEQH8hynAoxTRH+SUsW6sQlRxNX++45x4LsKGrV4HGwUfF
gBsluke/C4gOZ0IaWJXq2bcW6iu3f/mEgtFhyzqBkA3soHcJFxl72nJxHXLSz1Hh
84Vg9GGQu+PVbPsh3GchTEQx0DmKRLyX1D+/Aj+awASp4ZSxAY4vjJHUeKHYd2d3
Nz85ATgXj5dJTCiRlw3Xbc2ODYBpejfI7OXOe+fLj7Xv3Sp4vWq/p3ZDhnW8VWkX
THzz+vXRR3Ky3Q+P0j057RRuSNJo5phaEXjof38tOdnNCil3ajwVktiF9wJbjRj5
Hbcch/nYlk53+jERM5GFlrO07ynWdy4Kw8dB5ep/CuXH/5G0YElPKG0YQ9/afmW5
pnbe+fQxLaMeo59Jytu0k0xqV6H+/BU1zKLGoqUK7x4u1FB0gAYdMcOSFbawTtH7
dlVYZtvcBlZ/OQyKJi37Ct/0/I43I0Bvk/rgHzKA3Raw1hFsnkxk5mgjj/2M53L7
2/Nzeet6EXDNm0r+R4Vx2KGP1GwUbpUgtGsk8K/5ne2GYmhRBB8QDt4aqOSTtOvS
Jec5IErvarWZo8AdOiqONyBxXNGhpjo44CuwV0joUZpJIwK4yXaxkInrjITYRzaP
RULsfKWlCAKCPxjupgV/WSPk5WnyAyigKRHM3UfjXjbhD5uOrW3EvIczCqY/Ol6S
svwrYyTCfgAV48CXz5v4CIFpOiTzCiwPoM8JNTqgLJMhLb6p3dwYHevtHJJbEb2Q
7GtGOAlNOqUkaoUXgkCqhOZg/D4Dx6TllpTLv9avYiUEmZcPtCDb/VMJW3Cp1msj
P7va8pPNS/ZmrUoQF2d3k9LMWf4W3gdvoeRjJBkwhghZXO4F7jgCEVr7kSXW46Qf
ZF5Vwqfk/3BKFzGO4zjhyQCAgPA2EukNca4T5UkOKnGFgeivLtuFURgZOHORrYzT
c2GD+L4m6/zlgXDw3ut29LWwQLMEb07KSJvUCqxCIsXDTco599s95pm7jjeC4CfX
qXK75tF50rU+a3MRo/3oE4IeWR/WcEkLkL2T6Tp4ZyLBVFgFZPU34xTyVgUBniG9
R6YJWx4H4d8Q4W5wYdWMZfYPZPUJKBMlkPhGq8te3X6R2RJ/YfCrQdPOl4YeDguM
449S23u2RzKxK+c5QI3PS7/l+BfUb1GBWJOj0SicJZylbofambx8+y4NgQQDBZ/G
+ttvJTmHuQOhUUpvMeD5sQDHGMuMwEjwCsvCFiw1LSv5T5rbmr7Ot3N6AN19+9Um
AVEFBmI4wx8VZ+mjg2Rs1Za0MSGZefpgYtsHFxHPCwe2/9zQjbTBinB76906jRs4
Aq5jc/jROWlco+lFLf2ynhUw54tOHPHVud+xwmKE1AU0t0QBJGbiXBLdN/8jgpQG
jF1LpY6oVhnpMlHUP/mXZjneyd55OXSJ5GSAqlyY8iOr6HT1QMhbavQ6SyI8AvmG
GmsvXS4Jgsc886ecXWDKAPIy43Nyr06RCsBwg7KiGP6HFbTyrnqQJPOsRPHtTp9L
9SgX5AyLDT4Vbmff/Sx0oyA/QZwnvs8hNp2CvAtMAFJ7+zBOJvlN2Vz/xJYUevcx
n9fUEKE2Lt/yY57ryeMpw1xElewIXohqJLpyIrCcp6u6Z0LvGnPoWIHSichRQc3V
eiQfWCJtniUgzN5hBwluU7r5T+SyBQKLt48Asw4856uE26eFezUysJSQC5kHLrVW
qy7git+keZx8AzZVLO6SLRKfHro43ZcqWvdXQHJEQbaSK72c2D2gC1nEL6idiWAQ
LqjCNKtGL92tPTuXmuSN+cdouIYh2yDriPX9/ymD58fhJiNgT8v0V8/MIfBMCT3b
Z+zy8bgNqurR4HHtJXscGzBYPjH1A76gTce91HN5UBRfWNDXBgBnwCOH+usERaLw
ALyd7LFCDEScbIqLl1ZNs7nFd9Izmc5qRZ32XoNp4WRt+eh/hw12syXuakjXdNJ+
CSm4w7ReeWIlLYei3ilcN905dds8S6BYypRgVhAMsFTdOzLtOBkzNZwhpzmbE08N
8/85GBbKaxUJTw1etvFNwEZ+ap2/0eQoBExlBa9//GmNpb0z3S3wFZkM+uFNHB3V
jBed6Xvb81uUj7ftywzVeR1u8bIo5whqflyFZ/r+92ntAZUfcgzfIL6FgqTwiYLk
7McgPuJhpWs7wqfw3MHj3ekqW20Wf3vqFgJVXM83fo65vyQqYiVU/w+K9I5jd4hC
QAsNiXOzau1+DIYvf3q0mN+dYeDrHUZUZOUhLlXL+e0AZ6phrIgpBT2zbC3ocW/0
gbg3Ob63QWG0IrGVC2r79+Djfp4NoWohNvkde1QKvG1KgHZ2Hl4647ltCtZAOHiW
neQYNutVjlcS0oOLu0vv6b6OzmmJjm312eqLs05n7w4aIwb8ZDDwDcT79i5NoMtS
A+VeDFU/4mAgFHhlUBJwqL4Ul4KQGdulunpYNoXhz0gpIMkSuItsnVYi9CgNAPM/
1E10+YRnGc/hSt2n1lneq40by6d7nEvMK8Iz7U+2LSUZ+uDKLkHLncFXprHZDkDB
d+rvK4xC5Hiu3KiGuoDPbjAb0xduJKmu1wByIRW6LSKf1nLvAb5wdfKuEuSsG6QZ
8+UpMBTa0Tv2yCatSi+gR+hCeSmguGqOiuRXvN0AsvqsTs2ZwrLmHHkP/AHWUR45
WEk5WVd9yhl++AcSGdhX6AYGLu3bNQhHVuOv4M+g3Krwx1OVS4WgVlcNILiQRS8+
5ot1H69z0yankka9KyeV2Cd1AxeiqC+5gEtEbMAb+Gd2lRuO97ZYjljCLFOxQDjz
dG4wPDJHDnBeASkHUje9aZs9eM6sQU7jgdtpgszqRFXKCrBG9eOgT+Grpky1jBtq
jy81170AyvD7rZPaLxDrotgd5RgKWSkDnd/j7YoUTAhiw3DwfZSyBbLohJWZMZPV
AynBzASXzHzNv0GF5Ou3jakbqmKyJX6tijuWydUD/9tYu87Zr4wITfC29X82s1hN
Bi5+a2V9CgvSEuyrqQSuyrWIQy1DXc+nqO8WhYQ1oJkPOZUYJb5r6Ev27r2hYoTc
RRefx7SnxIL7a2BXfCyojSXszqPd/Iy+zWghH01wZFcGBIFtQT3fnueuCwa9MUpc
3VraLnHomfGvoDsSJ8yCSgqutGnSJQ7jqEnMn48Nruv4jSSm9n96O2pH3LyJBjZT
PqzCKrvNF5tfGDkGtduMclC+dVxmxoEfECBpmxQjzzTjpz4ZpPBeNPV5ypAkDxIV
nV0z95ilpk4EgWy4nKZnitxnjWpPzZLbwcNctlJXHGAIV6VWC//6jW4t72+zyeK7
S3f58mpOqn9HKZidIyEDUiUNSnv/Dn4YZM5gu5AkqIQ3LRgof7YogCjO54oSbwOC
1Ibln/aqHur9sGw3WvZ+Me1fI1w7w8RLxKENFYjVwIyJI/ieMjVK8ycoFm0q5XNJ
O+sD3BoerbXZN2Df2NN0akbvfjCxA3vC4dfnEtagsv3IxLCH8WjCzgjHqUozJAwO
8GkgnvMxMRvpPSStxFZrfCWwznywJTdykvn5czUSP8Kz+TOOD6M1t0EMa9VaqaTR
lS4VoqxPK6E1K91aeFTVey+SiDNGRg3PXm9lbv3BTewJXfc3BJGAkdEHEZ9hXVN+
djeh4a0oru5DDYrqx0AfiQYaozfHVbGLcnMvAwqGqyGz3KOjtgpmc/LV5QaJOgSj
zUCxYlDTlklDQfgcNBsq/q34UC//isPWEJMM9/6bplPBhp1rAqbPuK4cpju4UXpr
LUmtUchc45Ma0+jNwDK6cQ+LGw/VSu7NDQOvVgOA6M5Msg4HLEFCrgmiZ0dSg29D
j8hAT1hTH/phwZIRde5hNZSFZwu2K1/osWV1MVHQtExv9nfe0/SAeHeaPf/suGgB
p3Izwe7r3tKpjZL3mdhcjmlZk/8lMTMQIZhd7SjIfqCFXv96hQn+ZvO67AvLnJ0b
WhFG+KTnw75XZbtGO5/s8I8pZL9fZsjFdHGXImcRvAJ//ebgl2b6sTuX9JynlJf0
o7EvtToEOlnyvr4vqEAbtYRUkWk+sIoCUMFXzi8cjpncMl4/es6z5MkhCeXP2Ojz
FU2APVL+VdeJxc4IrzV3YMNNmyBmAk9dz1I90Zm4sce3odCgF4o/6gGYp6yOfQ6q
rbuW/M115jozjkAzh5ZW+tTLdzeYO2vlRYpjAfNT2gOIvagGNaB9VmcR8h7umrO3
mKdUeDsRKyFbEa7kzntBrMEiKG5eY4dBnHem/VjS39Q2s4JZNg8pJh37I4V9xEbu
ftsAn6LiyfQX0DJT9sscAE6mpow6h8cPuFXiUwqrjrzrkvFmavOFzlIPp4XmEPsC
flmkV/TOO9u+1CSHNinU5CDxUeskMa0iL+dnkvOwFh0tUP9GdN4JNJNyOqCmASWT
MdHMBvfe7Jdv6mRHge2cK85cDMy89sGd6UkclBWVTZHszwEZYaUFQplj8LDk9W9C
MB84ONqlrYPxsF8JnZ7/hsFSJRCEPEvr/kQ1Myxa/qPHVtPrdXXNSERTClMXX4mv
ZnMCwNr3MdF1JH+DOc3ImTZRAF5590gOJRK7RMSzRWhDnsi4clqSFl/ltLxatCpY
62TaZjroQBDgBNczReaBAlk246u8m69m84DkgjY8HWVLafYIcumPekk9kOrjEZnn
zVjtSMDVNzCnNpyEZXVeFcvUD6dyk+IQIvcxdxmEsON04J0JaYXJ0T/EB4JYpKpu
UiXmm+LI6Qlf8kpz5u1Syja6fxpysLha9z3WBUxvmneh/HI/z6YUV7T1wUkWcRbl
OpWQofHTxsjrHJuG0qVwcymiL8CsFZ0pyMsB/lYflf6eVTVvTOn41cTJvCCg5+ad
qqMP8+a0OTaAhJaVnKp2Ho7X7ZvQSoVV7mFLzsgQu5sOy9WTmY+8nhid+tYzPMcl
ieO7dMUftN59Z22N5qk+ATkGvCWYZ6a0ErgwM6wrTYap0x4fRuJMKOjTA32E7q1R
jaczxlHQTH2vHjLtSjRrGtNOpdzRpPs/+vSVjO/eyGkE95mRn/2sz6K4WBfHByU4
dUxwmXGxPXfifHxPVnHv9W3SYF75u8GxAJ9YG3q6dury8ldqk2z3dIQH8WMIAYw/
iXJU+cGmKTefve4F0BwjpdeoXeNs5hId8q1VdY94ceY6ni7GI4AOyowzldLUPAav
ADKLv2jPXSxVW8Z6PyD7ON78/IHhmVFsLDAhP/1s+a0ztxJfbq2F/J87WSZv38a9
FuJkzuhhlbnSrmk3YSw7lif4xDBOmwmFvjicxbnqj5PQAxAOMNvXzA9q886pvk2j
c2I9xV8Og2LaYUfKv54tO9voUOdV3tPiB5L4OM7MPtM262aREk6Im6k5LKHefAMY
2OvRmdATt5T5/Kqs0CBGE7DMd5oLloL5FdFIlcofEC/834ZGwcJ9rTV0KaylYbf3
V5z+fM68nSqrklDiinbGDuOr84zeNHriojQW0kp1TPQjC2mcoejZfFyabr/J1u5u
h3brIkjGGM+w2zOduQYeV293rKLnf0CuNmiin19hxVO6W6fB5H2a6IpJP8UgWjEp
WFJxc2W9RhSH7bPKZwH0iuheA75S3zsuxcvC30kxOsNiCMHnznTr/K9ctRYtS1dC
iNTczA0rAN1ELT76uBzPTFjKuSCsyUCJ/LHTZbx/iBLuefWIh+vR6/UBTyfmkPCA
nnZRBSkX8zmiYYDYt4ZHJEfOGBgdQi1VVWYVirb0NCy37RMzHk2uPCH0Tep5mB8b
Nk3YLl97mOR+cbQpEGwIjpsB+FooWIkZW2/Tyble/p2GDEbbhSgCdR7zazF7PXfY
hI6fx1VA6Ip4spfTchiGhWoFNsxqfp+mZs1YpMDGzDjOAWU/V0XtvpFyiJEG1f8A
bbT6GxYHHmjTm2UTshwwNwdFArMPCo/UI8SxlZce/j0yW18tk2+uXk7lk133FMOX
NVFGeEvlQVUfBcPgxEJOGqIYRQ/IpurbjDsUcuB8KfNg8ZaXJ+MVEcloruy2OT0l
04Jflq3esLuA8QyBqQZXWzeEokKInDNIq46aHV5tQ0d/j2hixRBEwpSE5yFKF9SK
v7dQ1hQY21Xm8A25UAo465xrJYF52zK48/IKxO4wQ+XRPwbaq4ozA3FUV1lZu+7g
ZIQMqF6Zl9CBWy7Kzr+MclOgeV5ASp/SAxwNOKjQDQw6Hqsu87iWUITI9sMTWs2c
sjarZzl00uFvDGyESCSHnm93BhuUPg3H9LBGF26w8+io2GBbMH9/e/cNbshT2Y1X
lHz1C7HPsrWkQZJbsrXhmMx9KzbpBhNO0TKbWFA2iOiY5jM5acIx594BpHgg8nS3
Zk1UvKSBg7hQMP4UFGwQNJGkm5tnFXdNecF7A/j96Bmi6yKSKjk8c5coFzr7cEU0
wy9szvqqBdoqwGHN1e50qomy0BsP55/RBkXwHQAet362x0iV7bJVAJXTNULsUFnQ
Pn3glPkqKXi5afeJEAVLN2tliNnwcV9GitewhRFHxkZYFnjmmqqENATcDfV3LZQB
gyHlfpJGRTsewO4KFBoOl1Fcte5N2L/89U1SzJOFxEBwd+NbRQhVkqjwgnQVrHPR
Xui/4B0rrzVMckTIPRXfTErdXBEhyQXUH/o5P5sMmQFz0VqyU31xTD+5pyAlOKEP
HX4pp+eEJP8mB2A+/VzaW7eXTGFSvWb5AVCkZXhU7ciEfrUwUF4omONSnngkFsd8
HzbieLDpenecp+QD8vXlk279K9QZHeiIh9fYu/KSYj8p3o9REnvKkTZVQwqnbEuT
gzYNWQjcEOR34m79zH3O0/8rytMbkyooZbkPJIHoh0jyJjNuxi8/XD2aqN/N12ba
Tl2DuU1KTyKAOcnf9OPjzeRJ95ynRLfWG+kx7dhvHyhL1wZvSuUExxlmFXWRJ8Pf
ls8XQ8Qh9lANs6ZcSGTowWxIVD9JUUNe0Bky5lr73tie6ZUl/5NIWpWkfIjgmPtp
GW8ATyY2o5rLAjbdahxg1ZzIa6+8r0TkefpRr2zQ8h+slz2MClIZgg1HNKXyI6uj
QFGCo1ey5u62Ibrur66lzlyrtu9N2Cz6wCKcQDmm//kaamvbyH8LIXxSb+TRG3KB
pRIzlddcAJLPsS8BOUxHEboCOG7ibKzqpAqWuLYX2sGUw+f1v84nbIdM3MtGt/YH
D+meySd4lh8YI7rvYrwZkbSCmhNgveHfi/ZbA7szCfCLjWmiYexOwl5086s6tgka
sSER4vlqiqvBpdZ0zEN7HJ2YKdxaByREbXPCAGxJnTOHjmzPIsoNGEKLfuaXY7cf
cH28+IkBoTaxU6BPeS178z04par8PShp1A+r6Tq46pI50z7rLakRdkHGDDP0Yc8f
oNXdm6UXFu5LAIA8WAVqQXq9rQ0bqNJB+H7DcQmVuNKRX/ws7D0b1yxGv9nF2+0l
C1PtRoky407UslyJR92/jaWIMyCXaXMNyyay7nh7bInpMGAHMgFJr8frVmJmBUs/
0uLWQWDe3Uf1uGjoOjrbC2UNRxEdrxiuqbIe2NlKXt1t1b6HlXM6CAFhPN4aZrmX
BFGavlyChFW6UIHuixzxK9jf9DQhN7v2CvrZ6ZVGoTiwbG6hqBuhAkGpWLrUjmPV
DnRsiee+G0b/gKPGvP+D4Vu+UnQuWsGt0UAagSnrUT9oYMmdNeELSAwQrT+Zc1oh
oTB5VtOgDqNIcxvxoHi+DKUrlwQ8ri7hawwHV+8BIwDIl1CzgEiTP+5WCdzdZRUY
P+SwZ1cZ9Ch+NLUVORSN2N2aTUMMkIdUxxQXLwGfZZU6EL0LDPf6SJHcwkivVaa6
0/nUAprUHd3Ltz6AG5MPWkKCKED8YeKKwNt3lnFHKMXgw4jUh3+zPDy9NNaI/55r
dw9OTapLYF8PfwGk4qEkxXMifvFhLgTU/vS9QJ5fQcuIFhc5XZSOlA3uVm+hg1GQ
PM/nOcWYTtVadyZ1f40+cW2OqGPo2aqIu0AGajMr4XrUtH8KZ1YuqsoIJkYQEnp4
5WpNO1LyZPnsrfDlq4b7AK4XQUc1o2QjnHpiXXA/BeQgFgPrq1CQ4v0WUBq47xbS
+GQgCpS72n2DZRjaFB8tDWj1CmXME26+nATYqJpxXDHiaW6LOUprc3hBH63ken2d
sWTkv30T7UByRxx30bFd4x5xFMLShd9gWETYa9ejKEMun9FNUdBIp1JTg5DzOuQ4
yDf0xqCTCDG1ZDFPw+MbREU03CAMrSGLbjZEi/dFQ1gyQzqhcZup1bEHnrKDFDAA
mT9ErOSRjyiCx8IMfS5EvYVMbTj8pnaS0EsrWKA5totKM0ckPiYEpxwH0W6eS6qE
KvMBtHsZqY0YDIDwnVK3ValXC1gNzMJ0TWibbgrGuVpA2EG72enlhdN7e22AAILl
iHFLstPu6jV7zWg57AxfJTB3bG/yZ68hDidLF4S5cxXmhNsb5MHKOq/fqjDhW2LB
CJP4SQXXSbyCbUqp/UDqWSKQ0tKeZRYEtXojiFGT2/KtFpIg9tX6rcLzq66n9l/E
YNLIecVtrFdGDFLsAs4/c/3THQXzm39s8QlJPOqgZ3mIAKH6a9wvOPpJOqSqbhof
38padCAUU6QgDDVraphyuJm8gHZUQKM5zZIiqnC7iZbQmFbnguWQSfuMYoAmexRJ
mM7KEoTzzNlZ4q5esuXj6ikejkc4bSi/vT+M90TIMRGBMPBJHyEBPXIb+iO4+E/D
Y7OwZ4KHSXuXP36IAQaBAsdnoYGhNfcCBssEA546Oy586VytKTQDnefgpwblaavN
42FzswK5Ofooe7HkHffmjLYhi46MMoGBKo1IVcxxAfEpL2+ZW5/gpzNpvYibQ9rH
3l3vWuAFaQq8tmAZ9eJnyNy+K+WCCrm2Z7N3ziMTOAGo1NtKbqW0dpXJ0Noau/2Y
ZUuHNLxzVT3XVm4bfv4EUanhSbDEOgylr5xKVD3TK13kj3bdWNFB920kN3mKQ0lg
6CQJ95RgWIGiuU2QORgJvWNong7mJl/zpz7cLbjsRmPQtOOp6z6IL3FBrmT0Lote
LbX1aYSS9fvEv0UBb10saMcxU48SeQVliGkhbDS3QpvLULshJiiRpkOOfB4M6JaR
XBuFuZm/RPdMSTWkN4N+Tr/FSUB0oRyloGqUoXxwYfdIQFBQjAChMiGQwh8/jvSw
AmAyBtF1cxGkR0dtgS0HRopaATr56F0p8n73vK5clGUhn5gEec/WrR1HH5+o+C+q
ciRSHWuQcO4JokK9Y4OVoASyCX4TnFj6v+ipF26Te4EE3VyJRh92oBC/Ua0FPgw6
eFfr849LUnjx9EyYX0Hfw7LHaZvfv50C8jpOCrOb60g3uexpw6cQywuD6XnXf8sC
0N/7SmPhcZ1NHqaaVV3s0Oqu7olPLRl7JHobPw95xwGfeGMdsasG+iOUshZI7CnS
1q5Xywv8vCG/6D7K9hSi2P5PiMcfGpywk7fi8+94nXzF5/ZCd9l0xOYC01zuUDMX
OyL40/1cv2YZy1UJs8XYZ1eAcnfS864yk+2u1NnQdvYlKdLnP35bcQqZRhI5xjNA
wojw3zwOTWEaA6EDQljEEN2HkKoYU/GMI6IiyoUaIMsSfVYlFdhWdKtxlH/AxUJV
41kUDM2yQCxRnsZjeccuxrunQ3mLjZ7yGhsx25jfuPOaI1HLBAQprlHsYaA74jqi
E+zDya8+JyKouVnIhSeL8m64dUAItmXnmh13wvoWDUdOzTwMFQyqTZ0quNHcOMKJ
kgLbhd8MbrrCVVTgRvtFKelbHY+iV97r5NCoayztoPXDWss7bmw0cOgY9DLu4Gap
vKp8D5LcOkd9pEdV6YpdHLHKjM8kOJ8ktYIzSovRsfz3LNUMOl8u4l0UO/s68cvV
vDCPHY9aJPU/w30AoEq51VKHjsZx0HBr6dSmByGKwpD1zeNQkoU0eba0dFuyzQJp
whE1wJmIiK5gk70K+agcHej+oRvbAIDuF9GiLsE+JLk8OiwSt/L+1WF6MaaxbFuQ
ihpuUWq9dLNJqu4qXv/mwv2RYxPI9kBAbaxpaCeFTrqozmZhrecmpRuipc2gw8PE
/VV55waUxz09KM7L1iHY+neN7ZCig5hQYLpPudxalFEdBIldeud4w0iXRR3ySC6d
noMc2VRn7kkXgLMHl7Tdeh2TRA8oUEVh0CPD6lbnQnEnrzN1QFQnC5idylkrEplm
HzOcxjCJwBvwaOYCgMSti04TUQdboYjgAAdJxTGASyHqbTz3DhFi3osnGd7uCiam
7fKzmh+BU7NjbykEGFjTQ+1MiLVIdGmQ7jlMdzRNX28ZWVptZbpzvEKAsvR/aw05
Mlt0+JY/6aYH8YIwMbYLPDGgN25JUjPjZzrnxaoitp2pgEnSK1xqDZD6+ZyvB4R/
EkKwvQvTsthGZLGmCZ2aDVgZ5gmT9tCWLni102lCXBE2IbL4mT6aN5H6z7fNOP29
OxaUAEr6PKDUGpsIL1EWTpif7lHKifcCKAV9ruy63rscPNDGOR73uBze0Mab6Aqj
wnMTazdVvPWt8ImIK6KQ+of5HbmKLiS5rtWYFl8WfDgYtCzFTu/8a32wO3f+I7OW
ITOhQsHd1uYZBwFJliFmgKK1vqmmP6cY8RUFZ9jlfr3kJvckJJxd3aRwLHJ3SWNd
Uw8MXEPb1exxE6J0kUvz1V8UAkRESs+wScSC6tV9pmwPf3ZYigpvSi4TvMuzZZT+
ekgUMgjPasK1wNy6vHZRcv3wkqqBeW7gQaaZPJRYbdEQ8kBAXW9xZtsaWJSoR3Ch
JdDjMvqI2+A8BW65a9odkFFZC8naU9krMCKjEj6PHAF7BdN9GWuUZz6YOF5vMEB0
xFtdQnVOl02f6I/YpzebmEuMgKGcVgs4atUhFNCiTAK6jIauE+6tYzzcSS++sZbt
zUXL+KCqtjyKgGaQdpOhTPIW55ZgCsg5yMBm0+aV+HzfWEPTUR+527Z/jmXo2imc
klGIL54+P/v1vx4EKKxuOdzfeJS4IoggpIAla0MPIkT6/6qzqDFrNfImd26E/L87
VL/V07DnBTkwVvVBS6Eb/wV5bZ9K8Mr7lMhH6aJuzi9Lh1gxuQnX6beb5IqVw8gn
sGjF/8/9JKTzv+xkOqpIS/UlTOV9RRQIdoRdj/c7PL38ivGCVikyAXYqS7Wc9rLU
mYOQ4bG6VHe3dDFfQSMN0JfYuu4RzKxHeNBr/dBFqDOxG3XJle8ma2AK1aP6e1GX
Iw8OqqJg0D75QYOAbt933xQZLHw9sCaQ82FmlXYwY4QUjXddZAQv9ILgyjHl5b24
uB7i3cSpE3yhj4O6y7fj2f2iYnx/dQm96V100TX6qccsjiA0KEOM4BdNWn0aSEeR
T7EhhzLmWgggw0mJZh/ZvInoApZdUEMD+r7uGDelKGyQ0j46q5EXGk+c8MdV6DXj
mQS8wf/5vruc8rzC9L5Q5KkjmuHTXvHjF+1RMDpOQy3KBeleQ08i1KoTdcG/qvtC
h9vqdd/4NG/lpjQSrl0N/GYsAz7BZD3UV58UZu4ta4V7NvdS16s321CjTNZSNyYU
qoXFIabkozRqdLC2LjQbn+tFXWg0q4KOvc3n9VVrHvG0bQYuVc17JmJQal+5taVH
8sP4hVp59JU/aaTPGq7O3wZngv6rjX6bLacKdkgkjIVo930cKcn+OE05VkYPPli9
GlL7jqKBXVxt8PtSbtnpa2tH/kdvKDYa81KibWgFMR0N+WM0uQ+fsVwbfaYMjFgj
JQ+PO4Lda+7g3DMWjgkMh4VhivPXe0V1vpqaahNO1jdr0HGQPuvZ+D7HOhtTB70e
Q0uu/cMsHALwu06W/M/8WtuKs++I50HzQfhOjr3/GT92nvsrqFbuZ4HVPijRCaN0
sS+QSU6uLH3zIuT/foUc84l3jYp7FMh29AZHnSluJ6Ty0bxKvNG8MU89WL41nyMw
eOrhGFQjB6n4R1/Mi93AiGj3NshtO4wzEpB9rv2PhZiaEyhprC5YSSJoQBfZvwDD
784q/JvLQ48hGHMrHaat+dXDnyswvXQFBfgxteleQy8/Mm7uR2jUabkgd4WlB55s
a3vTcp65lv62a9wKf59R9S6+emSPFu5In6ww0wfpOKOHbkX98uVHSY2RKtCfr4rD
yf4Uuok2m0aqTqUVdpQxUDW8yQGRda1ZMhrSxb5sVYZw14H54NQ6AbQ73PfYQZ8y
mFn9O05z2xxXe100DTQ1rn08p/LUfY9fjzlwZotjF3omwpRCgOOJGah7vyOObzua
6uMXE9/1GabnB5IW9Hz1qdteV4fZnj6xJ+13rjtZIs4KIqRX2V89Dy+G6jE6s5kH
NtaBf9fdCdvkscpspOcjN9Gd9xxXi2qwRQQNfMm9jgbVgeADmMsUN8DB5Wtl9GT3
h/coRxyKPyBywB7KWlXZKM4jnRxNTv72qLBDNnTBEGxefs3vAB5NuhZmw7Y8aS1I
3IkUHbXJSG8eqHPVJmzC8GFdDt//WXa0mkw3E7yspaxJ4VbuY4KotKe/BnyoV03n
1MpYTczjEIugdsrxyxJ343YBXSod9yxTemqmX7YKAt3rh0NUhhI9v9PnJUNE4gIU
OIOnqZbElsUV03Jz10V+mIaBAvofa6wuX4wEakjPbUhKsnjG9ZDXnn0zi3bvEPHP
H32A9U+n7zV3jT6dvlThCvaNHos2QDhhCF5NUP6PU5xPk/V0GY/dNZ7hv4AU1j0R
3g4JZab2ilVeyExAO5KJVAWoo3djOqaTg7hpIyQWGfsAuHuEBdfFPLxJBO+XZwdR
txE/YjTqkk/OjbWWGjefyv3pHaqc5MKNihkqR3TimLT3KSbJ5UloUw2vLi3NT3Nt
RkQuu3qs30hjyelRPc3psf+aYyNchHyD8m1jU1qmGLo7hdWe73CkP0r+cdoUEeO6
6HJ1B3kky+MXb1XjWOG9yEQAEgNcJIMU+RawM3CcllvfMFxUcCDU9qiaM5QFQrm+
Dofk1eGsAxRUuEvl3GBenW1fIQvjBf5I23Eo8zy/E6WkmSfhGth/cEQArgrvMxUy
uzPlNLfLbYw3BsMdc72pT0aoCV1gGal4g4/Clj2wauy2eButGNCDytdZX0D++jKV
YZYwjsYYTrYf9PmykfdmPra9BtCqe56e8CwplK+0j0iXvtrpVce1YzAbvjtChv/s
0lvzJonrB62lnrOPGU269pec+Q5yD9+lbDUnNveJDQjYoZ/xbEpET9uwLRObaM28
t1lPSaFiwcSzD0fKNabOJ+vRIWjX7Kq9e9U3UMFvUSSeZXEu2D49RwnDTo5YBh4i
XJG+HairlpcEKgv/Uuuh0E3KYWd5/byM51densIL+Ak/Y+8sQ5ybiLB4khbCHtm4
rz7ldqqGnwYnTdfXRioh9XnEV3rxQdqPAfKXWMg2MxB5ioIqKaZxRQoIJgdkJjHY
KxGsDtXLXnQH1tf1RcW5R21ny+Hbk0oUTENoQIEzjGmaYaj9QKpnF7MgUb61vWBo
JiKa+5dpSvqM7wkEn4YNaMBPZ3MX/dMFMYsaS5crJId3ypmV5HzaOwmBHhb5zwG9
DMmOkBcSzzCg7p8EHC4O6WyRJ01mdsQOFpjzAMC9aOhgttUrKXy5TvkP+wRY1/nS
Hi9T/DZVAAsKoZa101SuYLleUWJB0wgmj8tJaJfGgEZ6u1IEHmWkEI5Cw0wgc0nI
5QeUxrmoJqc8/uTMokFuGYyduufjhgtLa869/biNsCOv4aT+BG1blQoZgj4WwkEr
Fi8C7wNFNRR3UsU/P6KnEK/2i1PGnA9shIDFFKT4KbQt1SNmIy3ir0Ty6nFjIdiw
II7pdFxMPYvkLDK3MrMw+K+EERK4IIdGx2VGXV2NlZgzIyYData04X3xGPwyrCNM
Oh3kHjF/YKxuDSIIneDvD1C627mp6UNL88bpfA+M704Ncy1EqkGPzo6I1+Wx7E85
zNh+jCz/JJweNNvLiS4gadiYWQ7TjVLavrd77Ih7v3kdcU+e5fD3UfZCl1pKQbvn
W3rX4qNQJgsU6Nt40FOTBVBxaSR4GDUCR8okIdKJs//xjyIbdTro7VSb7Xz0Hq+G
uKfAQsv2B70S3rEAwuPETEApRCkAOS3ORzB6ewQ85SkrQBXiEjuI5N9h10cu1lhM
C6DTYzUwylX5rtLjKrV9vpksl7XR3I2EGunsAIoBoi14UmSnuVCVlgSqRKBvPNBA
h8PoV6HPmB/WxllSP7BhF2Dher/LeYAlBl7LsimdXK/eCQHX4tgNj+BBTyCmqjwl
NKIyI9kZ1KhWEeEIr1QXC98Unjh8GJq2PojfMqssHJHmrRaprp/7H5cGji1QkUBe
rZdbZl38yEfd+cwyCZKXe2wJV5wJ9DX0YB8A2xWWXyqXB0xTXTu7lL+oOwHpy+o1
/U6jwPPS4LTdZjkp5M25OV4AfGmA30vThKLk9WL6Ifb9pNQzor3qy3v+d8xRiDKi
yutyfe98wT+AghTi+PnaB03ZIO0OFVpu7GZQq+xP8FmUphxoAj+JUHlxbcNp3Eip
Ms9M4UHmE6AjHqsinMYpOAzrq0k6avMMVkvnXvhYljK2enmWfZrQVmAFSNyKUySO
X00B8ICPY2a1Ih7CUKYZgmunjYykdBDMUtkxQxTwi/QJ5c2PttGQG2QUZNYnn1Bm
c80x4E5eVcgtPGTiivTsMQYMxnfKCspdrVre4IAlCAsjWZ0RFg9b5AZ0GfNOFFBx
SAXTNaGXjD1FC5KivKgPuxN0vhCo1dlLj1oC1WlRsPuBmZgCIlIHgvBABSWnjCtj
ET3i505Rsb0+YgT1cvniQ6LrPBV0xeDeh6BmzQsp83o/vlxb58PsJJMj0aOAsruI
R1XSajFChYYCPDyNbNEWRcZhIrP/CYDQZp+ML7dlm6PcVZhtK6bUnR/sbdqxGvQR
koQkIgNzQd+Gryl5atLFL3CVTW+eeUJr7j2GK79xION1cfqdSkfht0cQi33Vs2Vm
SGoys5R64mTmeZdSNMwQm0RJOlTEOA0P5/Bt5SfJvXCFOElYGsKDJHugOEtldG6x
eTTpEtzBB3j8ngkrKnpjNOL8TC+BkkIlJJrqhAfgAECr5sB3T9Z5o1M2vH3+eVNO
UXTlwb/XCmVX4Sv067Lr4Lqo5ovgpG7A2D7cdpWpB5dsPWvuTUMiCJw6MQGaOSS/
24GBw2H/sY3JySQr5x0nFRr/OXVWsYnY2wqQ1W2M3N/waTYhwNYqzQDHn9UBO716
LaP52kEL5tpmmik7sf3GbIyjTWceY4bkGGK+w7/tBkRH34yCW/9CQuNMy+LQyyrO
ND4wHcwnKFLcPw63GezsK4HGfIJbQGfve7vcEVEQoW78w9mAQa8UTFiWt07JcG5k
429XZ0vsrdmccYxC1fmR+fw/C4pO2s5VcN6cMIXjgRfNbxnaeBoTcTkbsVxtcLCI
vtkfc9XasBci1uXI5seTIqZDmK9G0DwT1JdRIIRz2GZ6/QU1sDYjQT5XPCv7vNDT
Vf/b8JtFesVlu1abtPUXflahn7c2+uV1k0ikyMgfHVVM/2lGoZ8emob4pkaJHBUM
O115vj5WJwu5T3bGgOy5uMZBC6cAcbo+vIH0+/V/O77kxq7m2O2De3WXQ7a0AXa2
5ayQFLeOwuZZisnS6jJkotKAGlaRKpl0WrNr3nSqE02lNezdZuh6X40xrx5ZOS6V
6q48fLpcryAUSTg3CUGtFKj110e1xXseWx3SFlMrvS6Yo7Y3kqKAo9YbqWXH0Fkp
nT1klepX22+1nekmdEtz+tSY+Y6ipW4l08sKnt6yqwzFxOBQFZUJRt/bPn1vEOnN
/gncRFns6qrlzbM0+l7Knfu3jxejVv4nZQoLZdviwOVgGrL+E60xUUEzyavLWRqo
jUDLnbOnNDoPcukq2Bae9HmKNfLdn/i3AiM6vP8ok8Dv2KQkeB0SwjlvYR2kG55C
hkZqWm0GeV2usrkWI99amxayNODfjFWWn3CqVj7sRULuDLOP2jHm5hRxRv5ie5/V
rCKOWZSDp7ciIv+rqZmU/SBGt8QRFd7Q06ofQUDWww+kn8ICDNGzg9jrRfJ5tI1R
OBgTzwIpRdXmeGy4ghWjknwN9FiNaCE4kb6Cczic5VP6HWrIRFfXgck8s7WKZasg
6XACD1zKuRnx3G9xqNGcgkt1kjNw0NZzNuz1r5SfG70NrkBMGNZwzGOJ21iDCpVF
qQSJF5UrwfwEn7VxT70M08227mL3FlhxoiansNsd0RzZwNy11FBAQ4Id4+OZuUVT
tHeLbJlHkAxkJQ0jxDberuVDjDBTkFoVAvGVJaKVpR0aHLq+EPPhSzOaza0A27vs
Fr2abRirfK9nM3GHjYmATOR6Y9rPA/tB35uSRmVZC84rYaNFkI6mf0b2wVJsRJ47
naXj5Htc+QZCxOFHyaULd0i05wOahLskXWVpREI7MblVXj7Qnqwr1DtAjWtCYqWm
qc6VWmXnFPGkfHZatQzB+1vpwP3arYZYoedtmK1CnG/dd1rnVmQfedVLapOv5OLB
B9FzzA69BmETULMyMPLkBLd2ZRCQtSj5BdtOswEKU7Ky3CG2K1pPhJuAq+NTcTtd
s9Jmc88nZh/vKHYYU5AXZMJOPDLgzva88cDLQfrUBrrRZczpr5m5e62sG/Fx+ZhO
UZqiKwAVlyGCN6syuIIakfPjLe8OBTnv1V8RY+V2hRnb60ak+qX80tWgI8RGexOs
ayIFFnQi71sJH2095G8XtVzirZaUaXyKLzl57NPpJgBLPghqbkAeRhsPdd5OWQEl
mVGCE/eCrpHXk9PWPx6yuX+entPE97WRp97GshkDNnJ+NKgvZnymi9bnvWC48XE0
4/fQvBNcD7NQD7XO6c1sxJ8pt1QrHFb6KYO54kjT5ZCL6u8+N9HWbbCQYG3Y3fNQ
FwJL61RkIqP/0ddjd3OTXrnNoSd5wuwdQGH55ORzWpi4wbNsd61e/EljQw7P+7Ze
vd/raDOmwoaBRSsjZP6Itd59RnnlO20sEmmKtt2A0XLkIbmp5L6jMQJp95aLyymW
6u77Agt2pyza4qgpeelQ9TycKVhzptHYDBezjEsde3iCOiQ8uHQy761IuUxO5LIB
S2iEcW21imahAd2faS4pWO3yTsIzbf9aDdtgFrBlO2GfXOG3548IzO+bACBtp7O3
lL4Z77RN6mAe7TXP/pnMIAgCQUR6C3P0jJjoBN+gXwgV+LL2y65fnbC5+zxcvse4
9nUJq+WlqlsgGr36GjeXq61w1K/jOgTD+66zw83PxjXuSml6y4SqYVgs7ibMO+du
0rvoOKe6dxRTfOsBz0oNp83J01LerrkKk9sMhZOh9mfuANJ+Ssc0tfTMHhYGrS2g
aXqRqASruLDdgGyGu95kCP8blHjStiBb8cHsMfLxrAf9Qp6xVfhkY7LaYhjIsFOa
LwCdh5i2rFHlmOc6zxZEQ+pmZ62+YlO1WewhlpKIvWVQFjFWh5YqsqfEgJOPZDq2
DJpRvbjYaEcnimyg6TTuNcaFW/XLSwS6Zxg0Z3HLYuRWXMhsCS2NcQqxlvqinE8r
mutPtiDHGQIVFKPxupdsO9a502xTwm5Gn0InYYMGNzHITpoK5qanuKP5I3w0jqoC
/2fzgTY6I+VR6KkJAKWU+LeRzgB0T/PZGnWAlOQQc7ARWbqQX/HJSF3cXUbac9HB
U/vwyO4GArhVmPqPAozf4JYhwTpBSLHRbGUx2BNe29/ed3gDTsW3SoCa2yMK8rx6
b40XrpROFK4/+8tum2scJ9gQvePwF9u+ZIGPm4/USiZNTuJORTQ+LoWpZSe6Cr0M
0ezXXLpKkZYrRGHjvkqsCdn/T9IThmZUQ4vZEBmg45nl7wM5DKNm58TGWtLuSmCq
57xlocUlUWjdRHQQ08BlgsmlOqviJqFVr45o3s5O2xdLZ1E2Y4vza6vKphbuWA7B
/rI4wQ9t0QLogkDzC0eITVTTeM/uewHw9LNbbyjNgRWFVg1iA8ntralRWVVbYr7s
NE1DW0VQfAfXoCjFbksza9eBuC4kn3fduVusf6CJ1Lut6sDUu/MUGvFy9VWCE3Q3
B46gjqYNdGmYf54bgeH90x0c+TQUkd74j9uO9QylWRpYWMBiI/xBOGqPyIP0r1mf
CyE/VT9/Xd6tD1JXHeN8yCmev+1m9YHrUUIQwpQuIcPekQQ0lyPQ7+hVC7iL3cgk
+4Urcc/YUnf/aRGyD7x/rfrm5htqwVxQcqFJkBUutybpIzq9kbmMEYkZD8AbkBTM
YNle9/BhHFV0qTyWZXnhUCxUnoIHZv8AoqbErYkvH7p7ODMe1GtHHijn4pJjNEi8
4mTU7WiFQOSY4ZpOZWn3zai5hoPNci6mv9rxZrazZMl7khtpR5MkG3L8tf5btPnm
G6MFC3QxWr4l1a5bWRixOATzEJlW0K6y9017clLBKcB1woKgRCHL8PP/djcmxpwl
9hD2pw/gXJrkwuWXNUkgZMoSiGv1cor0bGvW6HL4llFZjRVnKlStPo+AlNk1Z0+U
LI5Bx+VHcQFs0l/UiswnO9hOSmM9qmRDTpnlbiGjB5gcvlM89PsbuH2y4LPVwk7/
vSTA2YD4H7GZqYEjTMw9knE6Xx5PHgfcq+6X6RkS1Jg17fDVwGyuZ3KcYBum3TPH
gACwytSnCIc7Z9wyQh9LpIspkQ8yVaYK0YFD3mssB9dzwrnV+tCM55DgXyPpLVG0
BpWRAVDIaKW2A1kr0/5pQ9Bj/YyzX5PByXlT/S+WeFOoi2XIyQ0ypwzLdB6YgWHG
xUku4b5PJk4TI9KOG2SfaBJRaKqgDjB5BlXZWTMZjCKkgOSCMk2BFss/sstNPkeW
cD8x3cpyWCbSm86+p1USDAXC/O0X/dL5fqScHpGUfeDyx5/zU5v4NyGKXlPskV4V
he+fSgQcPbY+w1svoRy3sV6fAo3nB78M4LKiReIpovUTGCQX/NhrxFfdxEzSqq9a
BMCaQJ6buqNaHAuz37sx3mAVOk4Sc/ADjNpxMlvwBvIon1lGSl1B9otRfaWIa1tJ
GALwiM7o4cOv970lDq8IfmrU+pq88BZx/4M5iBrltocH0NdT59l1YjaP3xR50oK4
skmTFimZ+f92ctNa2h/PTDHClFDr8Uryg2CmIdnIrohK9lLgqZvSl77N/tLCkxZA
/9/apjoxdFIiPQn+Ajhoae909uhocGMsM4XgzoDcRP0YkZ8x2C/GQk0e7tk5Rxt6
7iDrKjlcqJkkEKasjeWJvQ3ftybdP1W8Qzx3XzIQGwhVmPcpijyyPLyrJQ7p1wee
aA1J298x5/1d8iwibtfAyhMxt/iWPAed7GOuosO9ICT+bPzkM1npgJ82n+avmzGL
9C71d2faZTuvaUbmyi1yEvPQW3NTAta59zy9bvk/ZGrg3wqCwUy98NXJkmbzsC69
ZCZN6LXrQooJScgKJzs9x3/CCEr0q03hZi7aZj2u5dn9FV8M1SHiQVubk202dumi
dMEXdSu9oKZ7kpx71AOczMHqvaZL7c6q/ndT30OfI6es2FAC88DnQ92OR756OFjg
VV2V7NM2RVBAcqmj3KIkfOv7apdzKO3I8T4wVYfxY4abhYQ4NUIYahKlhvjn5kpg
6Dn7iy/gs/A4V8CGUrh3gBili64WrXBTzdcr4BWgkBd54gWfOgBjBUSHBS8AxuJB
UCOtyUz5FCQrcxYQWQgMpkhzVoQ2XgyjYZgmT8njWkBlC8WW/MzBJYfMsB7R2HCa
J49e0CEf4cKJtCZGG8plsL8g01r6W2JQJsc3sr57UUz6VzSaEvpjzPK7GZr92oiJ
f+m9eAj0NyFDHrDgWJOcOh/AeErJHrzEMSv6kucGsHGoTVH+dB8bVQ+/CnS8ntVy
E4a2QpSvzT0L1lRLrx/Ew3SnxootcgJ/QuQZUi+4GwxTLnP+k/2m0V9LDUMWpHcG
e8N52q8d/ARIJlqJ9rkn2Bz2C7WviL90RlQwJtnlUTe+ruWMow5hBzaEIceSpFKW
6dcS1B0GzJ0dstBeA1iM2H/dxLSNfB0DkZgHUwyi3Ij2yNq/fyH+LdX7It/sdVfH
eWtqff5WjTY8S55ybiZlpKm/o8sT2AuFKzJXEX0x//fo5ZH9/iv/aVHYYqo5oqko
CpcBxbLWb4p7ENGMyzlECB+3L9UUJAsNkQjW09LYRWTypl7Jum5ftXICp1lfNpra
UC3U1e5TOEY8E8VDCLMgwYW8HKdJawYtjgUs/4iP6KHxWSrnAY84ZjCvG3vUKL/m
vbqlP5thYjZSWhCXW4N5WidGEKPV42yoToW48qHEX3+yofVgjRqUa7tegz19macc
9JfNbctvl25ntbzd4JIzTGW+KXcQYspqhPktVvHq+bfSmOkfxUJHyM/JQl0TYUmG
26EDJSAmjRkkPgdSntKL5XJqpDW5r1/oV28rhz9wdRflMzfdJGM9+m5xrG8jyF40
L4o0rHurXxHHMVlQM4b4KKa4VBJi1z/My56uqlWcs+3vTqX9kocerBHC3Gq7nzMf
ASbQoyu7o38lSXsjWaN7bPQnh+gBy3JhKE9oT42CYvhagJSQmScq5HKsewdN7sH0
kCVWzjCg2nF2N5STvX0iYePlBLTqxWk0U4jlA8SRYgCtJSG0Bh9i/4QkviyesI+4
QUYAH+uhbJ69OvMmy0Iq7Xz7rVvmeHADS3ip0wSbgmCwYott2HSb6e34++0vP7pY
i7CvnYmM/pA/x/LMwAWkjhoZK3NMlMIHCGQ4YbKhARg4rHT3soL3n25J9IrsLf7j
m8SSiaDIZSoZTe+NfL4911X+cRvTxcYujfea1odc48F7bRv3n+Y9Ozagj2tz3dQh
+1Nu3Jlje1DO2RuooCO6qgw1Ci+dNUcKD4zC4NqjDx0ROhW2N4gtVMssckctXJcG
7hyEkyB9MNd12rAyIRUzbL+HCvuOybEUgMhSIk/OmqZhgSpB9UmaFIccEZXAylqq
Mmii82Z/2L7Fdxo3bfidZjvCmv7myRtIE08rhLrGZmMnij5ZBDF/09EfHJ/uH4eT
btOFgsaOyuXta/T6RbNzPfB8n9lamv0c+3wedzFpRWsNRpHVxYt+h1uV0jipWbBq
bR5ayGVTwzu7ksJyXjWwpeU4f3q5RZ2Iz54xPdahr9VQ0CL5Ctg3qgvXHpPYJ9XN
YD/bHKIv3gbKaK/PliZ0liC097mL79+76hVg2a229g0D/r0+2ZdSs7wPmUsSkX+H
DKVs+l8Jm5x4Rrd+lzATBDtCNnjqD4HxVLlCPIzj+oD7IKhTjGp6hKxFim8jOW1W
XMAkLaQDJZBEsac5TjlOs0jF9mhZTldH2PpQiayvJXfoaLAZw+q7I5kDFVLSBSFS
Rlu+B8GoL8p5OwV0s9GF+7lfpcuqVDEMcEMWjSREFj8m88XJUy0+Sfye0cgzZoUl
scTYeV2PlCTxBAWz7SbMjhu5RQz7j5Ej9TBWv2hKKd0YR9+Nwou2XOmjc/7FW7u5
1EMOgb1Po+Xh5g9dRhLOtEyG1XtbHjRet10P9IQ7pH50ikOFFQH4tVwlQuHhL33/
xOlH/+HtnKcgEpRVUAJcdd3aBlnUj1IaOjwB7OBxHO+DYoq8PXY2K1h+uA0wQFEa
v+zs3D8dAp2mpZWjhDRHEHwr6+wtomZ4cDrDkbbhbqZl31NaKDRXa9YeE50sLeRX
tJDDI9szgxEn7s176vuusDqD6DTkmLDXNmGJ5NxuxYIygsg1yxJzHG7+EoNQ9Hck
HCprjHHX5HAK9Dl3uwYEDY0KRh4ExFnjxAMWGSVKZngBsbX94476KFG9TB9SX7Hi
vFMsjKQh9GqiNC80N+sEQgCqWgcGxiF0WcHcJ6eP+EfFD0yVHyF6hX0XpHwybXqm
pSMNZfMGuR7CDs7w6jior0Oh4KcehV7sxRsyxVY/+JVbKBGmzrmFUfGMWqgtw99s
IG6aUXi7hUhL83IEaYIupFwFfd+bJSrA3uemIodqWI4QVfdXlJuVUIcxKG09lLz5
qXiIIpkpKNsYWWwA07/XuVmZxCgIg0qvrMtKecdK17jwxItvjLJMkD5qnO3ljpPG
H1q9agwDpPwVcjLf3QE2qpYRQE1j2sJVxONoZZKFwFvTr1+OS0bZkS+mKsbdMMkX
I4vltzb9R1jAfTx4+vTSUebdWS0mBPhblG6s233576xEQrBgKGcjdQvyE+E2mTk6
NRNnTC6i2D+5LpXCewpe+nvIfXnxs4FRCLK59r60HSuinOGTIoMczaSh7YBlJFLt
K1NNAO7XgLa4eia/yOyZSbZCTMfBOB/3QYHj7YSS97iytpXqGKXtjmMSD3AUJj4S
sFxPRgCGIwLa6BLca27ziSaXApgW6ttqHLFEC54XIh1ow1toB1dpaxWnKVBbKht9
b85Hn+0+hYSOct5zMiCGamPFYrfrXCLwCniHUyjPS1kpJ+UnSs30h73OowYY/F2N
rqUofyiq1qkkutimdnIA5s9ai2RP7zS5kVFeB9aIBbRVECb1wmHmd+L7qMk76C0D
W/BBTZxnY1ww9vr4jJb23iHrTm3XFEin4cRUJYhjt1WdFE7kxsy8PrXk3Y5MkzpO
7/uQhlQyt8Yxr7kic6tJaVN4QjKj6K2DjSZlKM9FoG8km1QlUBGwai24z8eryYJe
kjhfpXn/egVmgCPCIWVs+1ULhUJFT2r0OYt2tQRlpGHqnRi4qlhtdVEd9dEQ/awe
NwgTTmTFpNKrjyuS9GwFOkD6khV6y1nLMuEczl7kWd6Z/fHGZTAjO1eFKPLW+CaJ
1J/lLxy20fels/BW+qG3neKTrBWvx1uMRQJ5G2FnhTQOgmZHSAZP1qBaW1/oY4mJ
aurq9gIenUvdHBDs8S2jk//sDH5smjJSuiZJODAPJS2zpj7cFtlE0Fz7ZRlhLZ1t
rHvMpqtoDZmQtKZsDNrWwFZWD/bAZfksZjeKWoCcLM2Uf8/swQIlIvAMgnvbo5lS
DY0/95apTmKfNidNtW24gcMUaMqFyLOITEa1bLFsxkUZnEUcdvDETLY+l6k8D+3L
o08liBG9u2oEEW+nvFXioQJyIAxIRqyhUWh8iPpAPhj4dUUtk9nyX6UEdfjvKGZE
E+/qjkiHfJXNKYjnXGV0Pd2DVzyOd5TcI94vu+/yiPv70sC7UVKZVcEDYvIh4yJQ
YzhQkXRaiCp84PsftPn+NdENXGVmZxyPUItYK5cBGvBcJJDR6tYlZ88db/+Wpk//
9AsugPDMgbaC8KEWONkczkatJB3h4aWHubNhSa1kihmsSzjwDz1yYV9wHs6T19Wa
twXYrGrQ9Rlp/fjorjvln7CFpX72KXx2/ve6d07+RIBojj66POlxue1IpWdYt9T7
G0sWuwpt441yqCpdht6+mewEZV18OlM2NX9TuXgdcBM3WKKmrybuyHtBfC9FUxZA
7xpkNcsJYgEAJmBIG2bE1x+1OAxU+HuasrzZrWXHcIWTpQF6lsxgM/E6tbdFloDf
VI9KU6tmyzDP6P70l8e0P3zo51RVvBnjIg+EeyQN11f0m8A3B85+c3kmelKDVdaO
Hp+wLAzd1i6XD+ppJCsxXU8Bo4TqCANz/br8EVsz58Zvoz1RnEyfcTQQH9ZgNkEm
uv64E3HSqa+DyKyO/eECOMOjv2qwNXdh0VYPz8/EOtZ8W+RQ1eRrYwd+5LF1eGsM
0C09ZNHD5Hb/nP7K6wDROn0iqA+LHBXzRXCElKLKD2ca4HEDRzQiNuCyahsJ5gaX
1ElC9PCzdsOoMkgyHtJmhio+IruLb4u59DQHf0xDq9Hgx9eKJyDIfAyOOBcpyApN
dAW0go4Qelk/7pNzvjUtHoTjo07nmKlZVUCbmYPUJIS3jHMFBww469buKUqGdRlg
qROZHCz1BS0yCaWuQb8a4tCp97KDIF/dUMI7dpUQ/dcmsCAXrHdkvSqPH2R6jqKp
//zgWZxm8ne1jdHk5OMK4gFQaIFyVPET2Zi9+DP7lDJKtQbtjA0u4ni/5e/whMEu
QvVRRSRgrbHENHUoE73lix9de5K3rhRePG9WDUHiBFT0UwcR2VwosSSBniL6S9Yy
OEoDKtfDdJ0x8ZDeAWatETBUuT01Oi4dK6cTYEJ2lf5pAFQGz2ibP6JrPkQ43aEH
IsaKYnaNk0Gg2nQ4t5YciTXq52kuPGgnmMNM3hxj5E/3ns6Zj9iFWqUTBcjYyV1s
6oRVuo9D7+dlf6etO8V43JgzaQfwmio7V3D/QufGUhEjlUZ22pQxHP2Qm/3sC0eb
R8/jeKvQebi+XzjYGE0dQXptGk+7H4S8YMMoynM5ocs2AsxAmuXHTI4HxXcdynCe
w1rIhv0V3Use1Ozt87B6NeHbYG6U87lOIGK9Mn8hsXuHXqqI7k3VPS07hrnijyXe
wjIceYx6gDN9v1X3H5tYZ87ywfugOJWhyf2NuKT4Ub7+CknEfxhwqJLpxi3XE5/k
+Unw6uGGObTIi5iWiWcm9Il+6YF1GJ8NMieRwmh4/iEheZ3OKKiJNIvBEMuP1SHx
LPg4s3JJLUVbdh/CAHpr8LXbqEm5NK3HBHZ4X9s5Ya5Q0ffVF7DpGjbn/NCudCaA
bFgx8e+dRpNHfkFH0tt8ozGD9Rj40BHzYKoqZnckGlWBgAmDrMTLHxIEpSWaZLyO
HElr/TOLH4MHt2nroLwYqj10FmLvlUItocOTck+DBNr6yPx23AxZlQyTvi+GgTTb
J2yIGInt0TQxx3ItNfCO/TXpIMxNZTadpkGfEJOeeOE+6gj721yR/IV9yxjsH0Z+
7D2VJRAgsmUdoioWljj+A0uc3aintwTOCUQQblOw0JHGNy8J9p7VbrUu8iNXqMak
hAOgxcxbiNIrBZtjAX6UU1VV5mb/GdAHZeVfIrr0D3rN6mVjobw8N3ppNYzc0QPr
mxqFTI0tpxOQcVvGfb101r310tVUijswVj9wjPWT1vcQeTo5GyjtWsknn0red+vC
Mpq3XTfvDSbBGb/1TZs/yzz6JM55Ibe1lPvQ7XQ7QM191ruAcYeKV8dDlatzhee0
pguGduaPYqCEyABUU0fQrMo7iJjDKlDoobXDyMVgnOBBJ3yTWY/KhC/PJXL/ghpu
wsmDbd2aR2BTJcrS4uSjVkpSg6c6jW2yU/Tk5gCodba5bdpOfYdVbNDm/ayhoxW8
mOydjRmgReDwUvVIORxafY7DmMmVQN33HXovSqIcikY0LwwR4UT7n2Ygl0p6DZji
OpHRJDSqzxV4uxPLoFeQI7W9RfMQEDv+eD+5mIYgsAkp0nUJfAEWkwkKP8mKiTBU
7mXAcor5AwC9mv/77CptcWS5cf9vZiwbzLFN+5qjC2SJEE+zxJsaIzxAC6UTvW8u
6jd7rPtllMUulvgeGkzPdx0YHtlVvEJdyp6IGEJkaGqSq83nbIKvU4MUIFc7Mhlp
cQS9gtNswe942coEMGMuaCJ/wli84kSD5Qw/ghruZsnsW74syPnjuxuT63Bk+hq1
1ghPqarNcJqwQP3rDGAOF3vtaif0kSWFMcATxbiJNpR8KFTYe52K12IKKPR9AA/2
KNtmkXM1ANgA97b07kHk6fu8OtLWau8MDoKvxg5v2SmEx2Y3l1O+p1qd9hVR8jJD
9xEcJx3C3LbQruAV1zK1Va7HoJESOuNcThNoEoO6MbSD6Xp8k/aJh71f2EcY2x2c
8taRrv2TLhHlKGD7JE/QJ706dOtG55qsPhpIQwzf18dYouea//PMqtT0m6LnmXtW
1oyQgZ+59xIJiZrkwF5ljzUeYAyRE8RoleDhfQrITUVsAsJFbWf2TWLOss09nW2E
uZqLhQjv5IJCiFH6kfdnVBVUKRxexDFGCMV6xgbUBMdXr+F2x7sYzTgx8VbXPhWp
QmZIC3qRfy2iCcDogFthXBrYW2jyFt63jLd/L7llwcfIKBOtqJZutENMlGMgP2zC
yXNACh7gvwixKrW0R7DeJayIlzdKJCCiPztEqFEtULXZdyu0hei9g+35HPYqG9ha
VVISzcdnfblqP5zW8spAhmAAyJbjwb4tMacIW3D/3AESLTwvzGpsCTM2D9MWUQc6
2HgGLb3wCAZfeGcyH3E5UTE7KhYzHrCGuLD2AdI3Yy8tvtnunBygTzNmwmgciY/I
VCakUD09VdnOHPLfRoOkx1zjCsElI+PfvzIkU4CuOPD4rf2tYsHPCqhEP4WS0uKh
nzZLdmR4gyICBF9m/y3qzkjhLfZre26MVqW3c/ST7eHWPRDdrLt3+zrJMoQcKVH2
8f8xQs4I+WJg8a9wMoF/2emwrOyW7a90gqUryoyWGSW8aEJd8TW5UqEVwhtkoyKC
LX0MehpyWwZI4tcXqNNQ50k77Qqm4aBZzOvVEB6ORtQK9xsdMpc2pWunJ7ZIVKqR
XZGyCQJf/M6zqp0b6QevR7ln/bFLXyrbVEt7P0dKZYH2oDz/g09v4fcf33NddwOP
NqGxkBCzZ3OhNhJqoVC0mY53B4zGlyVLcgEM3Qf6k/whHxbLwFkRy9ATkL1C9AEg
DIlgaPiITr5pXW7mYyu8P1R0pO3z/cIFUP61ZQDck+UyZ4J4AP2YH/66sAZI8oBE
DL1ajEEtkvfPfMSTggdYe0UleGTA6qu4oEl3Y2xRprsvOzOAuTBVlYoumfWXpdyP
775YiAPdAXe4BvdjBEwswRJ1p9Oo7kqGCx8yVJhnpvXm249nFpR7N1KPE3Y9Iq8X
X5UKmZNMyXoYU+hp1JVa3qmIsQ9FdqbYNu30N1OMMAQvrpf/BxjwQ6AI/h/NF6ok
8eE8CVJtamhKDNHAPSoMUglVE26JqaNgOuiSHjAeKABO0zlOs8IG3Hh4PK9yKGY7
EQjwP4fzhHJIfKee59Fl/6My1ay0th6xh9lV7ubzabdwpalPkxdfI2CyQYyKoQPZ
9upPvroFIRVzEepjIRzKNemVFqgr1k+IyYwpkn0sI9juOeDrX/qBKxr0FNqxFTiO
hIKUAiGPGHoLFS6aGUvEljhxr3nf2eSlc4qEARoYHrxU2B9JFSUvg2YNesXfh7gq
xpQGhKCswy43b0FDxi2gdxzKzxeAiT65FgQMjukRahq3rU41rtplsaZqZPgyDnoI
2H4/Y3I8omSAqFvc/uWKIM6QN4m1qEAj+fNiDRUnzNCtq83fUE/40b+5DQXBYFeW
4ZeNReuuVvxZ6kO+7KmRDRlXZVC9DAX+6f4Z7S7chB+o0vX3pqQzvyG68QTvEV7q
d2KE315wVmNvV25HHN+l6htOq8J9bFxtJPTr04+ztywVfMBaXxtVtA2qGyxUlv0p
L8N3EhcGKSgYOHI0PLVSrKI2EBWyGDxSf5qMPUGO8EXsBR59IS+8A6/KvG0X3tSi
B04KC8elVGPxqiSUpLBrmbw3osc4CYkPCRuv2CMnQQQO2/WE1r7F0p0boyExtMMo
Lm0HRuEufwi8CJKjtDcwPvHcLMWuoWTRcHQ0blrPITuTCq7rbgG+gPKAfFdBaBPK
ex+6k1r2hivZL0poGWWy5QEZHpObdXIssIXyjGwWDBw7l6efDpSiWJini8SDzAtj
VpBj4pz3rYQjGi5FJ09m52HoHJEHFo7IArddUp4YrajcfvJxFynwISLz+0zgsBwI
SFivT7XUwrgU3Pe8HQg9ZPgXmjd9iVaM3/+Py9QB2OdrMsX2eYfZMHoIwnFrzk1B
Oi4gu98h4Ui4BXSIQOJiBDbtEGl9d3BWvf0xnckpvKdA1AKSOFJ9ZJLD46jgWKoa
xkwpfAeFSjiIz/oFhVzVaVEXSk8HD3VP0/9vS8LW9OWhlHNtKkGqSr24pXQzWJ3c
rJqs/rVfC8rahtil9TPynbPBuOxmYnu9iMnFWFDn8w1Z9irB+pOXpwqMzV2EVfsZ
w7q2nM98UQMl2LofK2ISnOXxuLZVd57hAgFoknDISGAfFissf5BhBGCzbYWbyMgR
fxv0xE4pxyXSgLS/AITDzSeLVJgWcQExS1XVWEBrJpGxJ9M3efUaLxJ+/aasr9Qy
6jQujs823xWe4GZHNrpvsI8dE2GK+Ez99qKQb4mO3yzpAEXu9pXZUBSucG/Qkd+0
x25LJRzbl/SnCBYxZEsHIyy7TSPd6YJjXFJOb7AcLIbcCh4t5TifSCaH/ui53e1B
WgAKbGHHv98AWFauo4ZV6Y9tRhaWqWA57nCxh3as6owWJJcJvp61sZgHAnndabVO
0jqpD0kXb1Zq4wgwUki5r3k3cqyZg+0/7gAb0BC9NYXeXobMkFcvnbAVM8STnLc2
fBiP6tWo/YpKFcP8gu+PmL1KL6t3Mcj/B8hq3TKYKP5wMWjFsMd17vicZpGHa4eh
j2t2Hw+xd1ODCfovqwzcJlct1e31sPfXwsA4bCBUCbn/s8vWf4JUkKkR2FPrjZXM
gpcUZMvdYr96go4K8nA2r4e7cSMw4eaoGUg1hangxCZevknT3lPasMQ3WSqRf6c6
fkiggi2gFG+mTAaceh3aqIzMruBz7TFreII9xCs4wBqbcDlLE8r6Fer53wqL2/be
IMvfIlNZbJKrYZk7nh3YBtOTwKRRX94E3TGs8hBmGudG5L43C456U9FKhHTT2qPA
1UohGnNA5boc+8LLdU3lgHQTBWR4odlGMW8kDNV5fTUeSpgIAdohKn9j797O6F72
9MWASDMUi3xKZJrMi/kHgK03f6w5aR+7uR/rI3BipZwRxdbpDpcWtIpNRgdvsbnu
4CqErxeGgRD8mkpFIl9Afs8Xx5z7QNrMEoN3QY1phyggPJWXjlRDnNuav8vyi9D9
nkoZlay6Fhg31PRgMYovJmRz5iyBKM4HVbOG6B8DAN3G44zRgFqlIXBWK626mxcg
BqCOvwO20DYBpdErouY9kumclFaMkpSYoUgoB4AD1lZ/BoIf5TKlwRo9LG5iElHF
5kmdytqC3ZuqnE0R8gVd63zoisaWj+j5LzWXrfiSMFOzExKa6pRAahhzpZO4PzuM
r/L5H1C8bcNCfQQn4EY8ekAVPkuLsSuxXQkujoy5FCwVe2ofcN7mU5+ZVIgOzXRe
dDD3LtHCJPkvXXQLGBCG+fc/PnHeDZUfrQEzNA0n6dRd450z6aH/661uhOSdDZX1
B/CDyAFku2HDjzgINAwFZL2k024bxJ2taj2yM1NIbAKBVTL4CSyFHgsRH3ljvwJO
7CUMkKy+zFB5Fcv5kqO+DYS5WKqJL4MwNkUKw75fsK2DYVKH4grAifMSJW8aYN+L
0gAedbwDpJWd4RWE3/iveIwN3HwsIwyeoiQNPazTC/x10dlAqwFyYGFdprpDc+5h
2RF46Wqpr2d7SEA/qoL1/+fLOYu+7+sd84QbrCGLUFzhn6Sq+Q6tI8imHbwaRe/9
muZxVboAob/DCoIpSJawpsIBX+08PKSizdN8AwhtKvtghF3rfzhh18rL0eXpYtik
utOGmsjw1l2lsL6+CYitPjlJN0Q/xQt5vRdcsVQKH9+ou6iwIARlquWIrU4tv6MC
F0sxM2ktIiTTbSoeoFeKALjebIsWjP56u1umB9ur+DcS7OFq5JodAIqbJysa1N6L
Omc6RMIDio+U6N8acFliivDIIhbgYVoaNu3M86UblMWp2YiKEvGiVCRzLDwC3tDJ
ayDcehdErmfX7F7/hieWQB3sGDAGUz/BmRkmm2RDZNRM5xWM7VSBAEK3vZS6h70w
p6Ea4b0/tOoNg1xrZlQjAwNPERsOYt43W6DNbAYJMY1JSIz4s76w83JF3yTKFOUt
iJDosmqn5c9KpH+lf0FosD66Rt0HNFbauGagH2VbQlm9/IEP8IVHa8ruOPJXZ5ad
LsG8hXiI7kwrZlDsE8AcIvqfYtoEfx2mwpa3oZUdZA2tRxQenK19s0dFxqp8tZ1E
DVFu6krytSQbAt+OvnbIfd+1hTN17wT5iVPVVDKTWRT73owfLstf/A11BRLPxGcD
v8jpojnbr21bVexoNXMULihRqaBaTqhk1q+BgJQRWSLe52aQ6v0XJR3+lmlCOYV5
7K2+t2BAEPKfLQ+S+hEYOyoVfHbX5KUiuDAhCXPX78eJi9APmRKvtMFEepaTmyZj
GTfcUoEr4KLS79qTfxOUJTWGkEht83h1ScWsdv+xLPVzL2Z2K/dUkxsTRnRbzDn8
GDwThQAPvwu73Y2h8DzmLRXh3EwYKCVMMPpQ6n4gCjY4PopKC97vLaLsDx10k4p6
k/KanOPFYYdA/EjfR18971hm0Y9q3+q7ys41yfAZVBI3sM3TNFEIOoFJJ9JqWc1C
50qHJZYPnQIKzZ9dwk1GApKd737uhGXDTZvtGGxkIb049+RBLEX7cFDrvn2uciVE
/EKCNerId/1dPU7pmrY17+WrnWBUUHk9k+nQc8WTU2/lT7hqk+xYQealMQv7SNqH
RF0NkT+K/tMKpXt8hKqxs7FlhSVpRUZGfUKfeLyC5g3uEZV0Xzp8OHjMAS8ywyHf
XzZ7IbnnGgIUvrEv2HPNZ8rQ7EVgFh6/ofUOQINX3whs5VOIChOdA3lPKSg5lSFM
P2KLD4i3BOql6CTNvjUaw9Lv44Ofx2UWl7o8D5P6DQ9bWIhZY7emomygUOLAuq6B
GVQPM+VBrLqs8xBlXxU12J7Z0ngu3SgAoK/tieOM4DAyuXO4J+ijEIvfwXAPqOXb
vzg83nkmt1x5ls7EwtcvH5DOaTP6JdaXm0+XtDx/6rEUMgG3GqIzLU5JWXcjrM33
cZ5Af2ipxHoQOm25jCvjonFb0BLNe/nLHecKndywd5vl/FN6ojL0DgI+P3XUNfab
GlJ+4bjiq2MZ3gZOSHNzKsr6YqG78lZYuyWGvLcN1hUNwDB5AWQJnUuHOkz6aN4y
PQFQBAie7SXjLxJvhbIKdiBxKKTPtNqnDxzK8S3hiUXMBedcwTQT+mXnmEHt5/FQ
JXzppbM36sgD/kpcDdTivohSGD+Pab6oIzZflMXli+MKmeBNP5eN0LUBryJz/kgB
v5rA3Qm6cizXSZuwHy5/M5L4GBBzBFU0rDPzKXpgprgdcrLlOWJvUzLxM2zQZtW9
Nn3YoF9xxL8zUxD6fLCs/nkLRgyMuvHG59TA/9UaRrWh2kaJjmK7lS91YjxqKSnp
RO1iu6fVNq8ziUEDN/rVS2LiqM+3VtsruJemUcsi70pK4SpLaNrZ2M+LmBvwiIbC
PCKqH4qmSeZRxNZgLJNTVKeQSectrB+arujuOi7fAM711odg97PnEO+F5UhT52Oc
+xBIV9IYWt8hXU+4H4z+qGTdOfsHRh2RMwAcWBMza/I3xgKr3lXicNtYB0WdSBt+
FlbqYizMGyCgNM7gI+rlnwrI1T4X0ptC5gyv8DkfETtEJgxuGDvvaBp0QrYvT4+Z
zbmRW4Yvc8twmrISIX24OU9MunclJrTSgH3WPjFn1hhHnxlfG4QIPACaUOU2WQHR
HQSdfUjZe2hoJthsTGkjP2zV8RDjpk2uoKNqTS9NAr7AcJkXX02xJ56GvrOODqFC
cSyBxXX0Uzmcy73QD+gok8H8Do5aWg2X3In1sCEDc98w/dVe81iqbl4Hb9Lh1cGo
+yZXWfUH2tkrFfjEU3nKMB0TGLamw+Lw6TqSBcccUZcxZwBhLsG+TBXETPaT/Qas
PXZ1AviNqBOMgBvWC3o4mOeB6kg9kfdu8cY4yL9oiuFupzWXLM6ZXpQ30Q95jqky
wwjKxjz79pUsabsQhKq4RX+4xKmL47qf+eH5AUzYhLaqI1LEa0Dz4hGdS7K7nXy6
pcfoI0O2BZ4WSly3oYbyppz8UFv7V3i1I9lfSsA22UGWI0GabWWGdzGeq9Yvd3/T
bh0C/A3TVUlLJbDWK219I9UPkLvaY22rPniO9C03D2FKipEizLiW4RpUIHvP/BZa
Ie5mQlD8stJ7XxsPGRlOiWUyU/vEwskm5znogFjcHK0uXBy/JjGLAV/cHqVK0jUD
Do55tdgyI3r70NzwPEWI//AUmbE29GtXjkLSskUxfkVEGfcFWW532Piqs4H0A/QL
33yGw+AGvDeX41DhwblluUpKQVQCLTkFKmBbo6F/1cf8sMzzGwT3Dub/Euq8nQn6
Wfih0rCh7cpR5nSztUfJrkxfEJIIa9I6CuL7he3BklGgDVjKiCA2Bv0/tKsKIoke
IabLt3/8hob8jIFwDWRn2+DLWw3Qx+kwu6PenXWs74BhH1srOg90vriuPcKfSKiO
sT0HekVay5gS27RGbOZnqgMym2SbMZIaH3h5dy5/J0Vz29k1VXT0LXRhiA9FRo6E
eubz4GepIcL+Cg3XO/BtcCnbk0VjMtos59QEv0Smf+9uxa44S2tGL45BrQYHL7rM
Bgz1rR+4PTlvH6jverhueWbWbWW613+XiyfJyEKglmBi3Kw56IrFnqPi2gXg5aaI
tisu8xMPOHlw9GhiqGWKVjipJDGviVpSSJhWkJLmwVLQq4XVPS/LfwDNC6kfThJk
C9O1qbZ1yiRMJUmfm1iSQg2bh2LRZ3h5tO5roTRP3e0fGijJLdte3pV7ttSlxYoC
5e0nZOrKcGbIG9zEfzh3hS0HW4ByauQzCwJWWfh6+wzkd5YYSB/l4oBi8BT6lnZu
QHBZTnhvA0oZ95QylcKacJLExPTAdx0qLa4wa/LBSVG3gqim7D9OqCHZyUnMMD5o
NynugBHLK18JbmLCnsIwENJt8+uofB0zK/lRDvVQ9fm6atK2ZagRLFVu3TRpUr8V
ah3hFA6ZLmkrcyOlZSkVCBfm7fVx3kJWxdsx3MqOFebP31qWPyF+MnqI37WspDv+
rFalTUE6CiASJYBbQh3mBmyDqKYKSRUU58MattnpnWLJspz+n8V7GM4ABiAEW2XM
L1ZRs/1B5TLef6P7sYpz54cpRW6YvRP3hAReMsEg+kjEGDLcir8hXgTu53EYWx0x
ol5/XTeAyrsAf2DxbSqiK4kwbkqxDOFEoIHDbmg1wXxVZJhAg46CbYQVYEhNzkPA
DisDV5fn5wmqzmnDSWq523KTH9GPQsczi7YTMDeNl7l4c+yfu5tXTJxGDI9ukPxx
6zV71jbJ2gNsU/oaS5kuDLp0v/pm1FB/hNhnbDbTxBBeQeiVR/XfDALSBmgmmO8l
MTn2/HLp22UzaizIWrYfOqgxkZSdbZMIytaQmogb788xfmdE8IjI1WuP6V36iLWe
ATV1OErAmX/D1mnh66uGETGGJhSNKusWvi+gYmcqJ5mTtwEbDg6IuLs8ry+UUW7x
8RcESR3t22ROS/mjYVTHDu63yUnMj65y13EpVlFCNJKETbaz25EpPCbMFFXIDmYI
h0Bp+ek0FbOIxIL2cP6YU2aQI4Co8E8HbrJ3zJD9sWuZF9Y/DmEgGvb79suln/Wm
ShqMYHD/0JFSEsUfAS+pmUOqiuyhtD0w+165HlVmVauX3pYqaFyTX38qwcRiHvo4
0LbV3S4Qr6zZLg3rCyT9+9GDkGDAKo5AkMJCFEDU6TPDKmfIjN8nudaf1dlVUmfY
9LCnwXfYZ+f1TTxzmWYVFWCGA5MEpKWDKxUscwRoFmfdZZ2DY8jtws52ahdtiFbJ
BCgMnBpLOKBxxS6KtQZLHmAanPcUp85QvPhVXQ4a1ehyZ93GKLQtHzkLBLqpFW2J
f5NAtypkIg5lVZVWzLfot4MOlweE1BVKx2aXCaS6jQwyE8V1vEnSjrs8pix9Wmhz
P5T/UFTz3xnrXOCUpQR6OHyIETBN6FUdQRAANH/QEwzhPAoR2Ly/xBLRMGkVqOqK
JUKMXlLbHk11pcUz759+pKr3DryJV1OHKlMTllCRIUK+quKyKPC1C9QeexLfr7SA
zAJUwEuGYmaSQB5dv2G9fcFNgTADN0lm7Q6dDM5ti1nvJEuaFHCcCHOXYsdikeOH
/JvVVQsuq9t1MiKUp2FKVB2zx+2RD9jJypiIlpuI4sQwFzGEvP7pqAmgU5F8NTn7
ktuecSrx6mD19ueqFST9t08xifaKiiSjUIDTs8wxRr8TFePNwQ23XRCAMqG5P2OQ
eYeVmCmVSrjyueGkszSF2rWc7QV0XI7tyozlYnOUD1zEK4MnCjQZsxqBM7f6Rvy9
bE652kusqnX6c2iQhwMdDDCqSvlMc9y7kSMDSNKtAEW4CP/AvL48tJpTAbuoAbbL
18At6TDvtzrblvJ7K1hzCl8pmUp839eeVg8wnTzzcAFZoMBGy+Get5pISeuM99LK
K82pIjaIFgcsVo2FlPPAe6zd10zgI4W8f6zCd/ONc3fFjBEk6cxX+qpoLxzc0XBL
+QKpcPzVx1O5K4sRs6StF6ykTzQHHIetUXPk+8L963pNNSIsQDA8h1hHxQ6K2Ev2
vWySkEggwfPjZALdHO8zkj+Oe5l/de1SJGwjk4I2mPEacD08mTsReycedgDTsCqv
2jAcV+D/q/CAbCSNqY6eAHkt2WAzG0ioYuFzD5SQ1FW270HrjaivCeYri0G+0iwJ
Z/V/xPAONqOCTHGbG9+BEH89IB0yz5yfZ01243gm1sV+b7GCctwDPi23njhrB3hV
wePcP1zi9053ZtRJPptKVY4zySg6425TLBMFwu/NXc8LLgTkWiZo5iwH7kBbRUlx
FJSIM10H0xtqbcapZXJZzCJxgzSmfsCMU8jQzAqWJxzIrKh9fZzJJyvLrSzlbhoq
DCsE7yciGil0o65BRH2B/9WuutjcFmkZ5xqM/eT1QhjBBRwFzjTUHuIGOeKmP435
Y9jFsiVj15DXEui/iOrq3MUJOlEBUahISaIu8vASTUj6lNF4UBzaf3B9fs9IRjOo
fpUpodjOPpeVki8OWt9+BZkX7MnzkStZXVk1CH2HokjMdAftkRxce3v+CG3WlC6m
HripeBp4gQlPlM2lGVwpn/kJForiGU5/oFHs5B+M66dU9CvBSOfaC0kJ/2okPs4V
yXzUozvS2sKH87R++JOjVPlXk7/3ZSw++5W8egSr44mmvZycU8XZucLfBJIRDRng
z2OOnecmLjDPsmTTwmn+sV7DMV8Cslhei78x24tea1LRgntZbAHI/ev+br+1+Js0
L0AyXoFUdIZOV464JSX1yeC/mUw2ApeG/2ojBCsk3t+WtOA81INq0Vf5ie7YZDVZ
jeJzDGSRJY1HlFLEH47S8aJAY9GPA4aB5j+js94kB+iRsjsWMl6pbRai1gHWERe5
VKlxyVgwqUWyJ+PHGlGQ9nJ2SeKxx2w8tp4/xK4JrSoBHB5lNwux/ZScrdjGoBzN
/siNG+517n/tLb7Gz2GMX1F5wjbWNUSOvgIRXFNn3qvHGdqdcO8LZMOFc8eRT2A2
+0tudQU0hmCjqMtcxzYnMZw1YpHjmUWcvmhrUt6CfAFXJaxmLjF1i3LGvWJIIhIH
GeowHMBJVSBCHUgeyih57gqaMVCMTyuvuJ/tIX3LLwEop6E1tfJ+vhvmFUH5z5ZN
ul1JDxZoDiDifsP4oajuKpSTrJCobu56faSR1BbrTk5kBjiXlUI/0MYl5XHodZEn
1mM9YS7HVOr+mFHSNMQCRPV/Rkt0G/1JG65Xdb8iNaswLgIroyEkeiyXxxaezEEu
ZTmC3+uQrBHgMTIqT3eSn0s108eyRqSP3o4znYw1kRJOWhRkQYLzs8mvY5rAMqYf
9ql5SvNoQMui3vXltHjufNYg8tL2Pj0f1pfsxub4NyqwAw523rYXCHTn4qxpJ7iw
tqumByv7SSXC6lgkOvZeYH85mkARxqMhivH+zwJHcvpps9AOzJJ2avF/8gRyrYlM
DM05HSL4haFquLTZnwZZ8XT9Ux24MF4Ne8le1FRoD0qZO4hNBMScfiD5w15aM3Hf
ouvs2D5Ew5SBuFtCDFUz3h9+AkajtmLViAo4HnSdt/Io6SFJKZtwhoPtod2ngqaB
LvIbXi1BE2W6WKtKMiX/UIIO4PwhHq7lVZQJBeS3LlXTXD2ldfePh8zqKvQWATaO
JSgv5Fm/+9opvNLg/+2wqhg3FkUeOZ4ymQvr/bkWA3KXuS3Yu+NJycRdvejDPhwQ
Xb73VUC6AcW2W7swoLrxHccrRhjOZWi0cQGUOe8ZKPrZ+tHUuxCbH6cFxG0Y5AE+
Xfby1Cbisd3plsMuAbCZdM+ko0GcAlrbckboa7JpOG/Cq1oDQ37OtjAMj4Uw0wDh
XSzk2Vd0UTpiB1vFdJY5aiMT41nbR7+zNfBbfMkOLB1dfdlGc8jiq7h0+jEjoZN9
pLSkDjo12jAuU0A5b0QQEm3II+krJdHnJqDuMGRmdseg0iSfxhDVck2gxuqbrukJ
Z5mHrhDldwerkuzoA28a6yHxONJaE9ejU13YWeH0wLgAVrTukDXHxFuWNG+je8QS
q83Tw9HeyKQQzRz39Gis63Di/r+wfDOqRCV6nPYsXlGl95EcMP1JT+aurCQ2/ZcX
b1VrdRNOtSLsIAmYESB4VLIITvgUkC3dgFafAcpoLDwIZ+LT3DzhOyLpokO3C7N/
G8ERi5YPszwQ6QpFMHfAUY2SjaHCwf5XxzvNaPZGU1ZxZf3/Y3qSX0VtGBaOs4V5
lkDEVxtoV0l11qtimPoczWgI8Zp56E2nQ8mYjya8ouZG2DKXktVpvhQ6xF7Hu/2I
MLkz8QOBFhBKeGL7JLqOwEHPTiK3LEK4IrefLWzHG1zmgbDyC1dzvmCwuqQw8Aaz
d6Hk1gcL4/wqpt6SstyPeml7ZPk2X0ka4yBL0el2m80leAjkZaLheikFwdQJ0KMf
zqJiZoI9CEI132mbOXmdpqu30QjlrAYnWBmL5rip4FIBn4VaZ7T6xzFUEuRpdfWI
JQlb7sEfKZCwFbWti2KqV3MoWb3p37mDT4eBS3q4irdDTmNpfhh5BDsjOAezKeq1
Up4O9guJY6kQ4pP5305ZLpM/a13cxxS9whUrI00t6J5X5jftB/VHqYn+Lg3BqOWC
N+xE6WF0HA+66vNaDm9OjCWEwfMOAsdIG0xHKk8MaIQrTvEOoUCICaLHhm8r0FVG
Gxa1YztNJvHmdjjQO4Yy9M8iiSQklvbyBRqlr7VeA/WFaOmF/tQip96htf4DtT5W
dGIi6dQaJmYg5dUE+nRYVVO94Ij0ofxeV9Gm9TdjfrL7ypTZgkNQZjZSxiHpaosD
hFS7V7XN/uodHsfe+lVsnSNkmWu9Vn0ui5dsDB7xlZsFp3kOoeTf/qG0+qKMvW+g
FB9hErzOspjv+Y0HgmL/U/8fTnblMU//n6a2Tqs+UkIXRrFjB8wFI12bzlGYLFYk
dSBNkaKwcP4e4d+qwxuqV5rEfBODjc8PLesBTiyP5+TvPRFc6rdq2vIqt69UUF/f
gpr+JdUHFaAedh00D03ffW3fh33gy0/YXB3UBUH6YFOjv9XR2SMIHRpweuDXSyjG
4hsgE5EMuzZPngkQVKCMr5TWgNtLH8kPbT4OxFe7EMtmrTAkjj5xiXNlI6JO9B8S
vMrwu4UgQjT7UzxxS+myImYolJVJCpYoeXeCsxRhPY6VZAnftM4lONRRHzzMJVw2
iIUMa3ETvYeIbGuNGMS0Gv4PsE2IZB1MINU+pEl3uVxf3reg1aBA+D5pi3H/Q15+
bVsxhWfA55/A+3cdM9DPcVWe+anQ1izidXLpaqMpNUiJJY153YKagoFld2/GHCT6
agjvcDz/t/Ko0HhobeRC+HvIP/2SNlmqHX7Y4ken7kXso5jh/BwIG3JKOECfioYX
kJzi5e+4Jfa3TwHIdIBNsMIgN5hQCeKD1jtoB37ZARehEEMzkvaXy4hkfm71WCq4
ABoACZPPUKHqqcH89CSorMCcABfuEQWYVCCa15zez1tqPucvatekjN09O3HHSojO
0O1xoupTvGdCIa+AGWeBtcQRpHfg/ABeZ5e8w5B/LiYL0hhv32XL4Gb7tHBp0OdI
cKZISunLwlTzx+CL2RkkIvRvDHmvIbj5uvjNJ+1DFafVkymSVbkQEaYlOaW9KxTE
oKXKnKqyA2FWTkGjeyKvJWYpYTh9vVXDPOSEM4MXwpuCiwt+QvYdEXSjLtAV3r8V
ACKyfgDQGsRl87tC7I6aiv/PkDdmgmc/jYAB5EbCVxBJ0AC6+rF2i8EoDu5vutse
6t1d7u4HZ2YqA4+TxyxBdlFyrRkjvc+Kw2OZQYweA7iqRu5vFpp9NU3y8a5sH7/M
3Dbq8lrFc/o5q4XNb3XECW69pZQG9w0usVkBQIVTf5iJEMP+mQFFCvEt88rVP0oY
Wc6AqAmFHnPjuTGjSK8LSUI1fSdYVWlmEw+JKkLJeyAG4n8HCq4rq+MDqXE2SIlV
LeUZ2DNW5exfHuXZ1DQPDdhmVgSaKJVw7zqTTrZCPdtttLm+C3zV1qYmmglMjm0k
9StJQ66YuYcOvgL5DKkYWMK1quZ9iAq4JJNyrwzDtyw2CCeRjnG1aXgZlVcJT8aC
bQMASCX7h1q+XFof/n8xvbfGTef0a9/jKFV7FDG/NfRRsf852H80EtdNiK+nkqQP
egegCZwf5wAFmkYPoJ9DcsbSpKVcssjxAQphNtxpFqyUla9mXt9WDWSnizaGct2k
FjCRJ7FP4I0XbAdf5tGjpAC3Vk9h9LvxO5cgdoab7nBL1hTBNo14L2qIm1N4fvpx
u6ctFTGav5MFatb4nCJ6M1klFO5Ky9R1u5uHWT6fy/MaM4xmy6136BmxL7yZIMIx
1Rt7fonkSYltailG/GOn4rCqEmINsys/J1jo5UOcAoQa6KEO7n6WvfCC8DT58/f0
Ic8cCPv+TgW3Y1mjkyw1JM1PQk0bf84UD/Pv7k+8CCz8CEfGMouAEWAPeQIXkc7x
QTd/4ZXHZdZ1+B5fLfhvLkodBGU5eDoWO2+Nngc7mOJBI7eU+iJX3CbxK8hP69R8
MecddN29/3r6kZifiPg98c2eTDxqtiyhlnXCo6ozjTIpd68nM6HoBYaSq8lSkQf0
X6swcKfmwB5CVNlM+KVOg/QyazTK9rWfk/L3IsUwLYyL/OSN8zVZS4Bjypnc3bOK
N58PCouVLJfbxi13idIUUuth7c67qEfPXoueRXNAAb1i4zhForaSPyFf5XQBZt/O
qUbS1ybLu8plluZdzGKWhUC7s0MNQqCwLi457tqXPXa35vu1vJBtLGlcgC4AyZ8X
fycN/F0x9w+UC7C+DA2C4gF4ukCtX/xnRMM8N7mvQt7/bwl8dovna20Fh5cLR1nd
HSzKWKcd6JdACkD2tvDger1ChyPGsjaPaNdsdrQjovbFM/FpWGBsbuIXN6dEyfQ9
SwtsW0X8UA0S27/vrhkKP2a948AZWq7GY3Q/ZR23si0jGmikCtnqMh3B2iOPgB5Y
KHYH/l3NCDf21/8iqv5KH5sYGgkZPrlQ+Nv/1Rp1dE1DMbfxuuRVIcjal1PVkh+0
ayObO3LYUpDE519k7d5pInaPd8d+hstGxaPo3svGUq+IFIqkhQVYRbjG8k0Am/gm
oAKzfW3VTaKgnqNFSv/pEfHRYNJ10C0SAhVM/yckHhvWTxPrpX4ptEnkUlVEQNHl
wd+iP3Ljbt5MSg610o4EYPwjR6bde7QjD/ssTZkavNy5qhpaJD1/7vlvNT8BgDMk
kbsekK6l3sKY7BqJ2dtIcqxTwoTeOkjTJOTaxRQIfLOfjUmuTJuholBRaNOZadm+
kbALXuKN0QMN/GcodN7UpAeWW/LzL/k7NwMmcK4PemT9wkySnkLWUFFKecQ0VT+B
RYFXpvNckMZvgmrZLXN2PWGWQLMVKPYJWMbR0mDV4ZJeqk08ago5AlugBZPS1w6F
4pWn8xAaIc/Mt/vqK2kWfNmvVPT3ubzgjMsxPMGbL5pb5vr+si8+0CPyK3a8hnrm
bYEMmLSBlhUoMQaZY1NNBCm7E6xLNJC4CTrd2xHKFw24QcztVM8mNU+zccahJMjJ
bnZCCeJhKwZhAgTD4xmPigvqSlFKH1I4RZfUUa9fJ0pUo7cyKh8IDASFxpqIDn3S
nS0m46OUy8D8+afP2x2sa3FL48G24eqjXsmmU8RNa7XREZW3N5nfF+CAbX4F5U/0
yj/rDaV4NsqM9unXnfr33YOG4oVxrWtvGHA4TShFvqkTbc8mdLIzz9Xf3sgnJa7E
+FCx13VCuT+5etevzxlRgQRK9xTeNcGBHmsbqsbwO4gk88ZklgkxjLPyyBYLrnmb
V6EjrN/7Ly0UEG4hQU8yCQQ7Yhs3gK6QnfJeLyT99BNgoGGYAXXf7vbZSoRA7Ujh
U9rUlNSMcGQK/Iy5GGiNZ5qnz/ngckb1zuC8pKfWa37ezbOfw2UejBGJ+gyy5tJu
zbSfuEC3a8KJmvm8D9zFFphnUF6Pbxl4wWoGGKbfznQ9APF0K9B+FvNBKs+5eKp8
JYAXvwe0uqO92zZ9IXi1QOPayt8qU0spcHU7IgJ53K9jMWXj5GFi9OTlRDhiB40y
HQXdD4xVu54RSg8z5lLFPXjjTN0S0UeX24nHuZFmM3UBNDrBuy9IPlNxUR9i0+Dt
XT5z9a8MjAlOg7Q1XFGBGTgfEMEuQexdLjalyv+VTf/BXAl/2TISDVxnqBvMUFjS
9N7T/gf4aS9c+xoXybmYUn4LhyRX7DqLV4kUPf53dPxpOmN9/Ex6OJCZoGnGooOr
aHRqVRuprxbkzBB6ca8WLKcD/ppwEq46MBtyTQWJ2MaVBiqm37o7IkAsRBr1K2hq
sU35GJbXIrdM+sQg9l5v7O2PeIThVgoXmZxBjIoqPjs3Z92/S+19K2M73nDpaGpI
Vlw/l3KqsjM56/Pq4lu2pNA5d8giiPy2lZmwUt6PNQdBQwangrOzeJSwhTRkEOR4
FrgAnqngbZrd1nxdpjxvNlJMhmPBxwcIQGMErKFbn97SMj+k9Vk0RtF9qgKKxWqc
b5MUl1qJTEYVFDgx5SuK9qLqtHWxMPPBLGwPpKC9xbeKzeybTAJFyoIKXrsApeI2
/raJ0nKWN34e/FNUsPJV/uKgFYv2ZZd0aj3A/QhNb47BRFmy0eK305NtmkBjLHdN
nhXCwZFoSeCVAB2+r+LbVZG/t/t2TXxTnedyl3v2JdsnCzzbBDru/125wIJaE1qP
MgwqHs+cjA9eiPB2kSV6Az+xaas49Qbwm4hGFN10aLTkSmum0EoD6E8a6MsRaXB9
E2QOwXuaSfjQgFLAP8WoOM/2ScEV7pT9qwSPMirC+qAP09/1exTDSP8Qhs5+QIAP
0Je2kbOJf07RxLEzDFfJ9l23zNT82DS6kVPoqKE4aBWidtTkkjhU6iWthEumqcM8
2HFsfivRIYC7xEgXRrcvneCA3A1LrzsSiDqU3/rw3wZSIJmhatEitMERRItYKpfr
2tugLW1FTx0oJWXhNF2ecYP8smZ86YxNjFCctCDENyv7WKcw9EHgmzNzJ4K4z3XA
4SGTg89loasUnV862xScg1SPB308XA+pPNc47LYWSh5FS0+9DfADk3grEUIdsRV3
WWKGfkt559foZINa2fEzNH6hQ0d5xuZCS+cr8Y59krlgN9EiTCgvYpqJ+lAz0E9s
dFYDGnjldLzgnRsqZnr+kUHJSXnyFE3rtIe9VfgqReivTEfQCruxzyIcUJOdqVO7
vYOr2d+QUp4zBMZX5e0rpHmyx+p+ybwU/PShgTBsigI5zBGtecu+6H9kz9jhyw0p
tvoLWqOzNzjCTa2PgJRAfO29R3qX9r3+l1T6KJSzV1L9uF0UJ5J1FgzsNzeUzcVJ
rWOhCSVHg5KDFAE/k0kcpsJe6X9Mb9zxmSUeN8UEfFA2k3H35LyQnKrrwo/dwE+j
SrX4A20cUsGGzlWGnx/Za335DyHvcvgSvrtIDJXaimMpCrt5cTGTONNWVRU2Qa+q
jmc0dJx3JDSrlWy3Qo943DaDFhye1+YOLhDRCXFWq4kD032pU2682hDleh0AB+5/
Ws9br4cAYV0QWOSjhfmoH8EPdU/ZCb6YD2l2M+cXMEJz9izjZ1MXZmcb3sPaxVMC
DrZbhRnf5rugA/vzw9HZ/yCc3sJRqfdXoGUYAk5W+zoZ4IJP9Hxws4j/P1ThjoAC
wPp7Hg4kl9UmYPaZkV3NZxdpU1npEPyrBsWdwLLhh+7eY4brZwD494HoeNOXVt9a
eij4wtbmrY3FGCDyEb2qmOnPtPcf4Z87qMXFzPvbdumDRLtqw41Uzw+mu/cvgIox
aHdUMjsA/UznQt/HTYRQ71r5UilY7KnXF69Mt0WVDVH7KCfNS2T+lGQKuuktEXFk
ESS8waer/XROVdBq7OOK0DREQF+ZV/42GWxAwOJVBc6pnufnz2OLLpIGX4rKa4Je
BKw2rC4y6vPHhPmylHIp+VIpJpJNwbdU+35OD3vfwRdXsm5VeGT7RWXSLMsY13tW
y7Mp7hgpJ/2ICX777lA+lFAbwet75nBHvi4YUecZfLYaa/rD79Sp2jR0L9gHy2kx
vePad+st9SAgV8L9ILqoQr5DvFFlNEKVbEPSZiuo4GUQRej89JaXv0O81dXXaT6j
38UFgbmZZpsrm+X+SuVYwlL3H/PNjLHuB+ylFo2X6v9TTMG9MAJaGUU5eBvBeAse
u/KKAiKQsR78l9Gfj8zBgetPzLX2QB1PUFL9GrV6CAl0jbt/gREM1/HLoiIJH8MV
DcbiLX/cEABj0KiXH3d9RyxMt/yET2qiKeIVObdBf4Zx6iGJyJH1+ehhK8LmPNO8
mfjYMM0nCGcBUPR4xUo8agYYV27qhkvvtkaDGYrsD3SPPYngK4dopbxN3q2U0txo
M4gm26YNgpfoIIDBylw7cLpRJhPxq2Y2jTjOHk9MZIqAMatPNwX+FxNM1sRb4Sqh
UGvHNyDJkp1r+kZ6Ls+L7Wkbo1IBxR64vc/EpmqO7aiD/sBlWmvQscGac2hr/xwr
GvVkIB+mW6waXQ1+6n/3wzZCOBlmVXQdtEuLgfRLyOre9iV+u9yrIuLfgsK8Uz3o
QI1/iDkvtl6F6RQV1wsXXwQt8hCeE2yUdfFo8zPh/9l1IKRBwBXorzLDaQ+Wp3R0
tMjKzu5ou1SoEu8ctNVoJFbPDtaCDADAc7uv9cXOmVtVmb2LrMsi0qOhP/yHMOX6
BGJOgMN9aehed9x0TEqZZUqKz6er8Y/6H/AqHuZRRvgavhU/V2SKPXeTn5jFxsIa
F0bnYuw90uFLY0QeRtev1aIAFj4mWecZNFV28tsJ+3M9sPqbcI6ija7xbacvVS/1
zI5oq0SCIP8v/81ZnPAVyrPDVq7qY6jPQo9yX6vDYC8orQU4voVzDokWfSv8LzTu
lRPBXcgU9kxxU+6bv/iVUjxYxp79lV8U9kAjMs8ebO9tatLqO8dojqTAKthcU0HU
gbpA5yIx8TJVnaHdFLbwB2N95iROeYzA6uLSA4lUYZyi+kAXqXUj0gdbBOPxV7tP
IMyA5Wky1ZAAlPauChFtjIfu+gWq1VCRJjcsu/VB1VvNNWGMf0pHlXV91+z5zkyP
8rlZiRw4CicdEgKEl6o1bi+ZZfSjQ74q+/9Lk92uf/10pZ1ZsjndGBWV8ZtXsIFe
PTnMAzQ9xL36KnhOy2cpVobKLB+i2JkuVp1rLIw3t5Sjwvw6V87FGInv0c6VbCJr
32tRVHUevtfVl+xGNHIymHGPIHMLbP78kWYb+DHMhU0vKT8QMAf+Y2dnZdHmsBB2
hhpz3Mh2YKpT1sE4tjNYXP5oAEhrwY6k5h0JiFO5H0qgyKxJl2Kr8/RyQeWESuNa
W9ZfRgINItrNe9rodQuCqn3a7hVZZlKzN1v6oH9OI4qp2aJzLFcAzLhFWRlJ4nkg
f4z/wadjZgspi71a//bd2TbB+yiiGr/nk6aXLdNMMk9LaOmQH12NpbRXUnvbZhUM
eVdSWXmTSsGpUzuPi9dhWenhoLxdCucrmhs/bHU/4HvkJN5TEMh/p2hxyZe0vZqT
RBia0zHBMCSp8fqrDYq3GDunxoTZxUoQoiXDXZ4RES5wgmnZnK1xqLNKsadM7V9z
ogtT2zjKZ7wuejzAxEURjbB/gIygIUe44zvS4kG7oyHBy5hG4QwLmMDECG2u3zMS
ts0X+PPit5XLwW4aQxECs/MwMaidLBIqh4SSQfq+OFvEpOTBwlf2SEKPO+IvgXRz
GAc3gB6CAySqPxuoZv+sUuXPjjgGdMmj41Lep/0naLv/ddvC5f04KgHNenk35UTV
ACk/B0Qdy5ydCj42OMlEIRP3m5Kf4hRv1M6UDsSwSm94Z/IihSlj8FIzR1FWf8zW
re1XGVzkrIkB0ZHwIJeLrkzMsj+PLGc3akeB6rawSMtT/YhB/2ziEuX1CNi63SFx
Ii/RmwKBKg3rBC1ScnPYgjtp5pzN0doKKpWvp7yvBaxjvWbaYuKahFyBvS5XhE7P
tpwHTpYkbI+kQ/l0piw1M6sE9vHUNN2v2q6ioenJF+yGUDUMsQX4fj+Abqmc8V0O
HN+7k/K8F1nF1JyHo7mShazgrpr2NK+Oy09HCmsFSsuLZtB6b2iyjXdPb1yZhHA/
nlU/nXrimQY40O7Zr3L2XQGvgitek+RUGn1wjwtMPxr50StiJilBh9OW1WXOiIjY
ea5XwUnAKXfmqyrYy67V7FIcDkExMggsYY3k2LG0zCUVJrHamiY4uhZDIiD0mp6g
9aerFmlq75mv2lN6IQZFuBVCarS02f09OxE/yo21NVBvY9bJ4iJu/xrMop3g5HCd
rhnFJWimOeKOF2pbVVgVW1kJQsVg0Iyu085ILV+LTsQn92BFqWAL9Cay7lj2Fhy3
m9G2DHg4xzKs+wfGd3w5GbRnSgelntMZQaogB0UX859QEHciHrX7PKACdt7Ce0E3
4BuHWv4lOeDjRDHj6HLwasoRALdH/R5nETU7qusn642zMGg8eYMceXAiKcj2SpDa
T0MUU/LgU3ks8xSVd3H2rV5mS/tISmUZXkfEyyLbaZF7lv+b4i4FqT3dbALXWRwY
454crrEnq7TUPngoQ28mteJeUqomNtsUX+s6NOlULJKEXWw1Qnn5zp3jfWkaR3TZ
TlAedv5+rxLbYWYogMx6iwaHgUltgFYp3ul/4wQ4bOQreu3ukg0zl00vXoCSEcwb
3GagU7hG4gH09KbMl8WZCnICCfOT09p/AQ6vhokz4noddXk4/uYHDbU5UVRgdqLX
KPi/oc/tfuaxbFRKMFfshunsoKJhxwfHNQM7ngD+KcKyvFnofnV4x9HUxDiKuoBn
0lzPzQIf46kQycri9Sq0dTfveklroPpyJPs3iyJ82pKY4V3kwHUzDY1De3XaarfP
m618j7oLtVS7BwVja/cGllDnnF/FfCb/I0o3KdiixsjkIezyfaADXjy4kdnu2rH3
tz9El48rKBwuP6e9eimaSinglAEon88mdUQEMkiqeteLLsTcX1lHMiJklDjOkRTe
7CzbfJIv+jUQJg+/G6RsH2Ut/BVxRX5g0XzCYHzmzuabCpkhOp1b01qV3Iys31nr
zFHzArlCGmVKbMzbkUau9Z1tEP4FLKB5SbFX7NkGySpJm+Y6lHsoAILSVxuno6nK
eNqkTsrQqxfOlB6rb434KoANRjWgNr8psOD+Actu3yKqq/fN22H6GDKnWz7STH0y
4t4E8NPZeZzF+jZLu4z+EwAd4vu5gL71ce/KkTF17vbobzkn2XpROvLKK/AN2Au0
UI+8PAqnYY7h5RXWOcZLqIfjviVbJccaGg6G9b7el8tElZXJ6ZahTQ4hS1X9ly3W
JgfxTHPoMyBOUQTuRkPFUqDwnwbMaqg9qYdoKeGDtWe3t3ME2Bc5MEZ4tJa2g8BC
uwM7UqDYs0r1v30PP8zFBAdMhAQDaBXavcWy6ti82S8b/YDQ02we6IhErz2C/f7i
ZPMTJbkljDPYNRiRG8dqA923wDlQg/liGdXbM0Eyz2vUvleRgRzDsBsCW4tknUbg
eEWYp0C8iFJc/SIVE7sdh8cvUhWwSA+VPw8E/5wMRkgbSHQA/3r55GuG3JV1NfCK
6/1E8FCu10oy7BthXMs4ke0F9hsdwvFp5x5i+ziuALqqLyWvtH/lszBzmnUDCm9x
XEBpi2nWyzS8z7WUh8WpJDom/K/hqmxmyR2Zm47WKyHXw/L/c7ajSBZIQmwIiQua
7rM1bOzY1k8Z4S3TsTqSG7BlsrsWLmUtUDUmngWE2No75jg9EjWVeTyNDo6dPCwD
pYnT7scP2U+dDabxbLjk25oayAVn17JU0uQ4yw9RG4LW9hpKLYxsJTDvXbxoHNsj
ogmx4r4aBaMfBBH59342wFmqzjk9z6Ljv41TqVWAzv1vEcB1FIw4098VEvEbgbqr
5d6rlB+pSUgH+KgNvVq0KWhQRVB1pO5nIbi6t4o4k0/DGnRwYX2dvfY+Xj57M3im
h5GvgaJt2+XoGZjTw4mFhMf8FFebpFwJmlgFoEateW90BGjTsKvQhGbVEkeVgQHq
H5LqklgzmevkQScO8FKykGKq187xOynEDBUB2w3sS1oRC1rRFZANYhZRuZoVH/2A
v53uAzwZ5uJHDc07LhplZRLcDqZaInp9p5fGwf0ByQa2methrTC+nVwfQjaWlA7w
CgwWJs2WDVNlIFZhEwbF2BxI4Mi6SwLWMuqKvNCWmcugEe0gIRCuE2jNZOR5hAv9
LUgAwio5IB/j55g2Po0QGVY9oVCcoswb/g19DKo/XvicwluAyjpkLP1jLv8kWs/T
QiCB64YxY/5u5zo/AiiI5JMlfuPwvv3CfRxWJiIVYYl4KduVeikli2tSdaOVgqjK
Jiirlh6Rfte9PynhJBkk3u6pcZkeTeofHHhTTznTOMLR/2crpEDT3slF9F6XQQl/
f2f9adQMPl9rFrM9oeu2RBl/V9nG1vGLiPF+2Ox6Sstx/GhROMzcR6GJNWF1CBHP
mGnzcQ/QxmNmhfWAP8b3+2XG0hFjuySobzVOO5gbr6wSCsHIw8Voz3gy05YvwTk9
L1zFmATeiXCpPkzpDQMj+w9Tv/u9ekJjZ0xNlJ3sVoeYslNffeRwQdkdaloJEJvi
579J+4X8F3Tf18vfpzRJEhGKXaR0swPePnPQ5whYHA7QKBsfV7CedDEXotshme/W
E50gnx3zyd3du7sOxerEbFe0WhFpNwl3iOcG9RCgpisAwDhQXj0tuvxqVJ9lWkp8
WfsMk2g4ZBNEZ/5tk/qEzsHqz/IBIO3RXBUmuRTDsA8YzI9sspROpdPkd4vYf4fj
VIQzW1MpNW11FpR/g0cmVOdS80n2uRuujbbz/1XUjEiCmkC5GW5zQ/Kix1Fi4bnE
jSDV7TeEDO7DwrlFCnmUf1CpGi4DVTLOBRPO+AsYUClogFdLr0ubIienCNTtQO7F
AdGEbdO2xtZUkZcwvLgH/YsdAkRkyqsO3jl6eWwdgM8/6Yst38gn16C3MgFDvt0y
ic33pVsov+rShhytsM46d3rJ554GQNV8J3YeLmn7ZG+srJnFELRMstf8P7r9zm63
I5fIfFWucxp5f74IuIsvDSycG48I6qjHdq82h5REPSpHc6dmOFSBDv3paaPVgDGc
gb9smsxb1W+4rk7EK7gEj8CJHtkeq8kiYfB8s+iXRtYwshHRzQW77YuZ3On40qNZ
AuUShs2dm84ZcAqU01T4TidGMody8NbGrExIO7JL2gazlh6/IZns01h/+MN6PrX6
QGt5jIIDbl5/8G8B/kevUIJ/OugrR+YyxXvdsWyVFUwdhlvtya+4VxDmhP/7s16Y
PEP/rZJ+OS9C1f6Dtg/utAMbiJ28S4op64xYY/jpV5SWFIkLQIj0BZ6SPcCYKTvq
d8p8J/gJZKAYBA5jeZ4Y+HtfVFtRjCKua+cXEpXle/IVTPQgCTf/WX/c9wNxLSh2
O5UB52stMh40SZJei649THffXdqonjjwih8IHOHSx72jhgLgeCCKd46I8EyNXyQW
u10bd+4gNm1IA/jklCIIl82Qu3Cx1UcxNFE4d61Tdv+dIlELacEj4TAEGiooNwA9
m4wyKopswUosVgI9LNlLZPDRGljrK4b60Qc+EhZvkpr1YN2kHc9XPsT7pkeXL3tb
Hc0goOgMVRkuHdLI4BkNiSr93lD3+OZfD0oOSynMecjUU/eR3Ngfvhx7U3/ptWX9
dAawtrDhDJGmZuF4cADuTnkL5vovcx/NTrAWucJbCoVuf5D0w54PFijOGn/LnApS
ld0b643zYeNboguKeym/6ucnpOGsFLSz929NsaOmYJhO21qpzkAxyJ7i6iK7LdVF
9OsksjMUv0oeyPZ25gVtuJUwcmuspIpK6Od+s1S9bYQkf6vWswcOTOxvsJks8TU8
oQ8zJIhsae99TnGN122ztWj+ikhH4MUjqMOZAvicQNJ+BB5ViiZu3+7hcRIjCYHR
b9L6IHvjM4Ap/4+crOioUJvucW/Ew5UnilFAldgj8TuOBIVkaWoar2YIsDLZ7V69
UWklEBAll5Uw6Io03CiG8iTtyElOU0bznAtg2Usofe7A+twiAC8my8KIuHXKb0IG
zxRLRrRf2K0VM8XJ0PB92pY8Jjp+qBYvj46uUKdidEwosc3dvu9yR0jrulZuw8IH
y1EkGy9C7Y/HzY8sqfkRSIFuNI9DDxoL5BbxuWq2ifW8730LDdVKehpZmHnQz51Z
fUqBn6lBOieUay1I6NZ/XC5bFu6y7GPAhHAvtHzSrldlgrgp1LiJbZRkFvdQr+zX
MvZ/NbN9ExYJJXrlFmhSjbYoPFRGBVQXog8BV5sIq2FoXDVwu37gHuC6bH4yk0Ld
QhbXa1gzXsM+2h6DJVXBf+2JGWz8PWq5igdyjEVx9aRovHsTRd2/BUoA/Mpqw5Ch
e6Sj1w0JXn5jfkMjTrAzqueZ1vU/WKoveDWJCNSfa4NB1U3ni6XMScL0yfavzMiB
Zw3sPXLOKedYW9TdNTPEB+U+N+iaKau+Oa+m2dQPcBxsBS0Y9P/J7RpgsEoEAVFl
yxLpIPFzby9Df+YK54CLGiU7NPmzN65FUn/qBVI4CHKQdl5Gj7iTRart2dyaTHC+
Yz0Io4eO0I2UeWKvbv+GezvgogPl3FLOUQCPwIShWJioexnDn7HLH6CCuSnLsfv4
bBBVc4OSXO30CH8Qum0tDm0RSrKUEgzmLOztWb/n5MBF9Qe0C8aH1amNVnEd9lTL
yGz7PaOopnRQXOT2A7zWI/IoMhmFsURSRJdPhUJc7sbA+O09VnXl5hrsP6VFnKjN
ZAtuWmVR81AMyu5xW5IlIzoicnK1sm4TGiK5BB6ptlZ4sLV8mLlmfLhJ4siJkClg
c5s8Tdpx07614lpkHXqXVnqQisR8lm55tNqyd+xruZESANzxP51mQ+Ws2+iGEl/b
dejMYVpm7S8J2+IASOLSAxNQHzVD667qSRaabeEr5Xq0xEhAS63xdnedABfN9TTf
HOo7GARWvmEz4dbptwsogyRLH/z15wu7cTlTbIEFQPZdmK6hqyHuOoG4JgE18Bd7
OTMNgiDhWlGkb10B5NRSgD7ZjWF30RFuQTZ5mc2I8gB48aV4/bOZa67jU1gh5+ye
YxKfPeslFI1nYhqai76GD0TBEZOXbcwsPYTQ6Y/G2NRJLQLa8+hMvWVcpi6cAXZ/
iVxrTA39hIEFMMYj8CDKIKqDWs3GIdg2BCgyrfh04JlVb8FU0bObwcEG4l1TwBkc
z2/Q4mVt3ITOC3IXglsFSwmg8up7ripZYuETHaajooltDlw08e/W3ejXewbXCYvn
6zfVoyN2vteyNdfkLqRt4PHCXuEolsTxhaXJJd67Xo9tWt3oKcmvKYdwz4thMVPN
mwVrp3vDKEYDOa17tWiHDU6/WLMIx3IpvUU0ZaE6p3cyhPQ6HUcIAnHxGO72jXeH
j4UTVZt8zaqh0PkdrLFagFVatGpH5J8/vryOwb96o228/3KpU7iAj0PRy/zUqmD5
3VyP2dm1mrXpeZP6NONxSKQ8KjwKLcX92s3znazS2EEQe8B6oIMOKlAJx4iTORif
HtMdeWZz7jZIJqC8JqYsYOfkAMBv+60LScYNxgl+KvZjYz5ZdqSnjZkTQFFCJ0T6
HHL7lCxAnpmp62YjLbUMZUTGBVGevXFx4uO3cUtfcPRJydF3yGey9xmlutckUNxU
mfZpz/cab1EwfTQ6w/un8doMnCTZsSGoTOEucGsW5JQ1MKJ7/DyzyWb5h6wI9B/e
aep9sWU3t3OnHD8vVGZLB3Jxd7tmlmBoQAG39oVyGZErRF+MgrRkozU1wLwOHr+6
IocXzpK5fRfd3kdXyWNBmjRzP9Xdn/35PalJebNbNfKxPex/eX6jOXE5O/C8eqY0
d8i03OlOsP1OS72tDgwU7lbXH62inrzoTDELnJ5Wr9Spd+lGojR4DtN3TAXyO1Qo
d7PFECPFRJKFuCY/hE4IZija2kjT/9s7FSlSJMo1bLkKh+2CKiLJ1uq5pL+cPLD0
BoviQnoPMSfT1I/awT5de/T5dpUxw61Tv4men+XNuEVI/Mo7+DtjrSZmzI9w3Lf1
cqCyl0MK9zCUEnbD1uExY2OVvyxJH+zqkyN2N8mqbiCZyDW+KHPAU5pAPiQoFzy+
ah1Tx8GToRNPctKg9w/H/syntPGqevKGzc6cwMgQ+CPWq/8oWI6wiCBoUY/YEpkZ
29gjC1P8WGB+zfEU96UX5kGv20EVRoHlSrSP5nIhB9hfH7HTGuUUgqm6MjUlVY02
HM3C0rXEkk70jfcHtLe61xTeuuhjE87uHhh90096pUxXq8YYs9tcwAH3h4Z4f6lZ
fTvzGf3LtHs7/HZK/3jdTwY5YpI/t2VOkgJMGM4gp0cXO/hRDsGpzGw+s9OIXP5p
eIRFp61l9Dn0yh/PJZGY5i5N3+53zMsvYHP07zxYghwCzDq/QgGb4khy9e/3cEOn
pBgL/KrbNIOTU0bPGkEHI4xTJ1rY8SldWncm6p+yfS3YrBfb6+NfCHnmLxb1lhLJ
yoWJ7Wl+L3nKilM0iLl7t2ZZW6ko1kbuZyLf3SqFbqhUlA33uDG8IMiqAGy9abl5
WTGdE98sRK0qQK4JQ7M0RET29m/1JW8stGlp+s3Rg24jsXhtxOJahOGXZXNjDF2o
3v+rRv4AcrMQeVEAlI7P7F1gSqCPfOjHfO+u4z5uSojj7MLYSvXRfuYsqehPpWgW
ppOmKdHxpxnRdRwCeQh6UBky0ElqdzmI/K1GL5hHU2BMQYo5D4T2oEli1tJDyBhZ
BNsHiUq5yDR+0QBbdhSkNVVbSsHeXLD75zfkHFNQXbF+waceWwqVaarNepBRVURU
zukEeWxzOggSUQ/+eFURoUs14M9sS5nMMeoiDRFpM2ByoOUm1TGzHY/zs1QKjh+K
wIDkcbS11/TOp8EasE8HfsQJh2OU319NbLcz/yvae+SO5kZQYaw2W2kRlimfMcf0
qspGQVXRF7hpRtSskwDDd+iKU4hhVM2ZpNB+PtwyZMvW5JwCxfy/BvGAUcBzDLQ0
w09MH4ekK0X3X7lWjiet3v2HG5GDCVVFDU0Pm5beNDEfH5PitUiCUxBbYwxrv4Q6
EbZz2vSHhCHwg8pGGpohpLrX3u6vv5Q8aTgj+WTsO2DXe8JX+5DccnONtIpyROgg
KaqFzoXSqMHXiD8aWExrKTx3ee4IBwqTWFQ8UJotPvtPcBuWWRi63kpzDgLCuqpi
YcJtV3fBsPY/X6tlNxFjhw6bzGxaiVwsMPDpBnkz7IGrsT913UIS2a0Bwh7c/LB3
dI55BrzNE5LVRxhqVlOw+etLcSOW50lpZAeWTEr+m0Dx5HEMaswMjpq/+WrVqSEL
obYAkC/WTWHEVefOjO/kBLRGWDTqXF/CABl64u55991+P/kvNPIEETqQxavlFGMi
SNd66KWX6WogADMF2eO96F5NoyIbL7QeGp3ftFJxQDqiGgMeUnrOvzB0CeNnDZ1s
udjjWFqChNpiLgJaY8iP7tZZdxlGtcQ3TAhbk09VxTKvmQVekYE5ma5IqIvI+dQU
WhUJCFnJoEOWfwcWPpcBBOj8SDjRp/UFiRDZ5M++m1d5I03Bd0xnVEh8jSG2RBhW
gZWvrqHezQamGDYTf8lRLmA91gv3DTUavTjWS1os53NTHdPIfPo0lU4xDd8Tn1Gk
Sq8lIqO3TQ4H675OVpqsV2DABPZHJXDyXCarnxEk9ZAmfIbl6lDdFRu3WI3nt0JW
Y+8LANF/ljC+lq5aNniUxO/bqR9d3q5n69rV9b+3tKww7f0WntnfYkHlIl0YyG+H
1Hlb9pC+R9jFnSe1KrX0RmQ2OWNcLKH8z9p0PO/9bvTIuwD5zn0TrCDAA3JeqsqU
5sceP3TqbWC2Gxf4kqaM7Ng/wuxGWfKLpuuF6WWfXHxEBzfJDyD+fD3D8ZFz0O1f
3NBhBXVZHUQ2fZ6n2fvAL/AmbSM+dHLjFDP8WHGi7KLr6ORybWMlKMokHdXJlCU7
d/61c4AD22xlcqXUzkdiKfTj73QsjPhYbY1K+HqvuUUe2cXLpScJa9FbLFRsEvwl
6RDZYJHXFNK/bPCm5qFgCa1PTjJNHa/69k5ZXQ1Utjubu1kRbuWzn9SnQAYvyNoN
LG3GOaceacBr0+40dquGCsyoVRGyaGkpqmZjOy1x0GYvDpEVi42YGXxjaV6u1wRI
3q7cSiA1JknznRM69ZLBf5ofeeu+9HmVkkcMb++MOU2eNzrn3b25nqC7UFvW2Qwk
qtKhKZ2KPws7GRsupN+Ep0lxtv563v+XUDyTKbX271pwP2FkPus1njyL8ZiAjTxG
OpKoz9f27kt13bP87KrKZ9yX2QezUhZq0RdUO3giLBAx9QXXoZe8wQO0NhHGUi+T
NbX92H/eMJWVndPIMYtClRqJDxDujqLZANZRM12RmgZwKC/cLUwFG02KBvSP3CGk
sQ2mUTVgMMy/IVX/+wZYhmo3kb08Vv6ckRE8VMJbLshgjQ3QM5rQ/C1dBuWoqeAH
jE6+FLS5LsBc5xqWnpIcOJ7MOV4aA/UBmg5aU23GOI8l+38Xws6nTRmN5bCUT+Ff
hSkA9ZYbO86yszXzdWoppXtuXL5tNWUcj2hk9+9MtS+D8Fvz73DdwEWN5qU7swkh
7g25X9CyqAsV+hcZAO+hfJ27qg+9cL/Zh/26IdR8aVk+KfuhuHTk+70AqbMbPF/P
rTucJTDZ5XJK+CHSlf0epwO0WhCxajHnwxDt/YZpnAAkmE9AQ89r6h8r+e9l63D9
80sKAspQhnZC8x5cxQZ1k0QNwCxEreuCqNDcKyt3c9FDuwbbvwwd02gpAwpmLlHk
fioGkSkVXD4q9IXXkH10I7Bt/VxxO3QF2CSYqS2JaMHXMKJWfJ+XTcpsxsUZBwcI
2xIroQbzqBb5nS2X1Fh1NITjVOytDN0BB4ISvydOe11BL7E2aDFw0JsGprZgmst7
aBFIg0WUWrzAdLKXhvzFXT9F4i1OAnPwkI7CUTp+WqlVt6Ut3mCB0pkdyZeERGWx
iZQ9AgnjD2zj/BhMxYSF8xtujmeGz2fxpuva5BtgZZe1fQoh9GDHnVLZA3t/SAiF
2cQQCYjfwAE/pC3XUrZg1A82b7UOB+lRXAaW6bxboZAU6vfhcNw0ubAfEkLOVA1w
pkcR2i4zGinIem4T2s9/tPbpNTuFgb0nf/DIHAt+7IozqdP4FmclWjuN9jg3Nma+
7zrwhdHWYM1nMTjFc0czUN4csK8JmBI9/zd9DK3A1hPTP31MGaNCbepk4wBD1+8I
IRvMQ3mKwCPCMqSuq5c3stHJ7H93UudzLzJvrw7LwBLdkgOwCKqDigvRa6ba5iXG
7h6KJaaoiUA5l8lBR6/gQcaXPEtdikf/8K+hAWAzUSjGNd2GSiFCxuKenee1Bmmn
j4GUkmfwwl/Id1O7J5sirh5Nc3MewmlXoMoKfU4Pj80LBqPACCixU9tCct/w8cO5
pOsxLkYZm8Crvqjdxm3Qt2Mi64dbR8f4B51RZT2phnL0QUGg64iUeEkAzsIaJfWU
mXQh1f6ET1EVV//rQRp4jn55zKIRhK/jFm8k4K+t5hTVgdUlwoNoqy5fHDJMEfFJ
CK2gltk9LNSHnvHScisoQIDZiS35SAJTNZXhDGouUOWCzXfPoCGEF5vLWt1nKR5M
/qqBV8udCgGod2PSSjT3PfMdRsX0WPh/J8hpK5vrXCi1/cqDIairbrdrzmXLaT7K
aW+1TJuD6nptCKWWmZKKDnNp410rNNphw5j8zXc/gSSK6QjkTCyKEfpaDHTimxyL
qLhZA/bMn5hLJBklDUoaodahSFdwqYS0OU/DTQCfDc1xZ0ZxOyCVnHAud/uCja9t
obWeMwNpQyoq3RJ8kzk+ImcY2V8t8wpeqDby0sxsKgcmTayq7cWq9eGS5zvAmGRX
QTVGyb1eQpcHDUtCxjRng8M/FToOHBigyXdmoqivw3oY3aI0lNU5KTMlu7YdF1gk
Q9P0+gEqxUlbL4RJcSHcLRRT6TT/oZvK3PjRt82wc4qos+dFjzGPU7DZGYRg9Voy
5qhEBSmdYUkJM9Drk5sTaDHvyNcP5scB5RTO8/LfaIhXS1Dif/71Idi277gNxbkX
KY12vvI/HdyaD6Jn9crREapzTZ2vTmTPk81RCz/BCaULNpZeAn3LiCoMZjuMWzaW
NhqBNF/eXRgiTqnTEphftCfiwD2wGqOOjylCO8OmTT3DQwvH2TG7LddezS6tPkcL
dcxVsumg54X/GxEVgw/kjpPYFf+Abd1PrqD8gYHfO6nPAga5X2WbB/FErDdseIiA
VUpSvStH8PLe+G+pAev67CDo5cZDJu8konMAPxM7T/0ZufK8y/B9IyOWH1Ac7pgx
T1swZtdaoxnfnFT4eH9pwet6SAJ4ZIhD+zrMsWsS3lnEz0kyVYitCd8sD30naUVA
VzmsSvemQeo46vPYAW15eaGRhJSmkJPdv8SCsjCiNK4f1aNhiSzo+hwjFi2eFclj
awdvhMIH5jiK469dZa19OiGElCO92gn+v+Jhs26PtMFzCBrXnUz9OSvaUd0vCMPu
vZeLJkD7k9VXCZrFuzjG+5frLy1CqmT2OpkqNoDeC4m/txZvjF4gEve7CHaIzGaD
EPFDwxg9fGoM73V/8keRyhbSU99FnhiG7gSqSdirUb4pkZCISl5Tw42ZPWZeynRK
tIQ1kkcLIVxmiYfqdxNoR0IpuMW7cvFDgUVjasAhAnArp9WlEyp2l2t9WD/wIpNi
NI6onr6KMjYJEfIZpDK56BMY8i56lKRH8m/gS1pDTIzK0Y7cs70tSB6rhdoW5c4f
BQryrqDmws1kooYP9YVZpQJM4Hha8+TRdfyiu4H22IEo6lK+N21JYFJch4uyBgOJ
2Lwh5W5/jkhNM+jW2cly7t2ctDihtzlF6gtou/oUpjAeA0HhEzGdOntSmNYJbirU
N0UH3Z7110J+VDCgJfIIXZa+WBooSLyK/utGTXu0Y+w1AsSe6lsELVB9qyYw5yU5
LEXad4/b/n38qY6KDFVpq00IXWoXsjpvyC1/JwdLD0jdYx1V+QaCRUoS6cdy17j5
GRH39F3/tuJuOUuHeVkZOiWiYeaqAgQaSA1fK6K9kHcqlzLvn2LMVeHTMZ0uBNa9
YqX84EOGFwUEZR2550cb4kMNzaj74QbSnwsmPT8jsxLOKuCKuLSe+h+53d5oBpZq
vIFtAV/WnR8uvi1MXB2k1Eoiv0eAvT18kP5K2vkc2hGKVhL2mOHOuZk3MzbdrvV8
pJCev7KV28U78NU/Yt3OYAyLSyy8XLCywrqZRK09kPKtyCW4YiweadV237JgbFzp
+QwtjDNz5DYXawHL9tKEansrN4IUyw04xGV9xSvOgnv4bie7rtigcTmQlM+3cAGq
lVt/P8Z1MMXmQX63At3LQCrwCBtrDoTLN84YLXBUiWz/PI9KVgPRo+rAL1H/8FMK
icc9tJN5WjwIiIKkTLPjEGfrqaobEv6ENO6N7BqoVgP7zMv1TuhMrQDc08+u/c0R
BTSYKWkwGRnQmXoB730Ta6vcIpNiD/gIyfCvnko3DE8WFHyvmlJ+QbgVQg6mY9eM
O64LWtZbSzwmi3Q+gOupTo20yoFKe4W7TA53ydAbO0xiiU3kbAbRtiyOkU494P5C
S4mGFq1LiDMbXCs79wcJFv7TPeuzRk7gaZOcPYZWS2LwcxF/1UOFuMVk86VrIsRc
gZtgd6qfNSZmQnmba3FCaR41YMXJ+fpOFn4Hq5xzWe9+NwpdfARsrcXAHMr5C0TT
H/AAA3ZRbcidvIMpMRno9J/XnJLXNMP3CxtHoZbk6FgDBnM6Onb7iKYH3ImQ6DQ3
qiQSLSscUvmqog1b1k67wVkq7KtxBF8fUIOdegMYK4aj3U/5bWzgYB+BQ7nSV+0v
1I9nifJ2o+H9vkw0Wn532taQFrEoPXxdaHaKrLZ2Ka6jQUNcT7A8TTxF0kX1AVOq
RRbJ97bVPDaLBilu06qCwL/MTxRU50tmxpN7N2lV+OcJlzMzJKEcc5AJ4+BCJN36
V7dUFFKzilX6NrFbFv+kwrpdctG0xJvdcqEZ17O44NNjdXGBbBoT/z34eCgWNqK9
F8eBlIw8waxYhB1wdmHuWGO0ILJELyz6OfGcNVOC1QYcvmvvLNL4/sIwzcNJoGxX
32/+C+mKk+czo5E8cOPB5Ksf9Wx4A5RLsFC/12+zApfMZrAl101wHJ3GGufi0zAB
S3lKlEp3Eu5kO0gY3BZlBu94dPWy9QdtZiHZyIjNh/+IDhtxYWQipD6MiTrLPoLT
eFUAY/smx9/5NRm5qPMl94aJisCgRHBaZtvCjghjvkkhMWgGjW/CCUGjLNoIPnKN
H5XtDmmWnykIDUheIHvacJwqIuGKsNxIfH7K4TLWMsPkw9k+H9EZFZQtugn9W7Ri
5IkQ4FKLxZ6/8VALZTEn6TBWTnoPQ6Rt9YVNECSXBfkZpWaD8M5m+JFGQlVrAW+h
IQygi9GcxmEiL253Sge3BJa6079CwVkNj/mEhypQC/l5GKnntuHiYx0gPPREY1ah
+AEXGifMxeaer6vV6xp//B/y/qfGc4YWrWcYMa8RiuSOKiETm/rzoNWUwDjH2PZh
417y7fR7mM/HtyzYyGqAKKOU3wNmNs4hT2P1iwLRg0OhDbIw53h5ScsFGVy+ckgr
aAo3zYk8bXeHfrBn920W2OiOodPNEJMVvUx647fGpvObIb9AUR9hkPP4FXztg0nR
PE6n2fabqStAt/XddVusBfjvUkhz3GHYrVkmBD5x9JC11xXISq6rziBT7elMCU7J
MAUdnYWs785TX3G30mPUBH7BFBSy+mSV4yD7h0190dd6zvWTCufD79C60IYnOGLh
q8ktjpwx1Ro/uZGVdGs0bgm+7WFlnDRq2IQjC99x/evkVXADUp7UKnrdoyD8dROm
UGslOOEVj98dGHPsBigpNgKUABHHop3QrsI4F15IGLMVu0KPCHZUMTOUs5S2QUY1
yFmMlRPi4+ixN2cPXNem/WbBfSduJPi3jzcGO35WaKpXsS0ASI8l1IN2jCxlH569
Lsdk95pfWHlC2xO0U4Hhz+igW/bux2ueWV7tr5WbmKY7mWjKUN35nLtLFWYDG11J
/RD3dL4UVIQFTn+yAhfbFcBlmjx+cd9NeVqc/iCKBVEjxsvwwC7DeL2VJSeigSE7
2TjhCPkCPOdv2YXwgQuAbKGS1MxCph8wDXMfR2Y7IPxAOZC9qmDO8wtho/RETJi4
FBRYfY9izbaoo+eB2rUYq4bFNFJHfXlFIOnk4wgngouz1s65dPNQJ425U7efXCp+
dRYx4SI1pdqeSVXtGJ2S7ZqXUvpKtQYSZJ6uBDNykZC5cckQoKRiU2FCwfiXsEIP
8em2YDEMqO8DFTWs2XZLlJOsVCdXd0WmtGdaXsLOzKNNdI7FeLnEpe5aRAF9tUZv
EOUWmFPJPD7bm+WWKNGO9hxcHxvN+duLEFNpz3uU1l/MSoIgqXrdGPAWBNGaTo2L
dBpluGoSj18GyC6/v7eBGcx9VMYos7ufvhmePZ6PaXj7zOCc4a/lgTlTE1ko7FB0
0nU7SluwIu5H28F3aWahtJVC4E0XAhfCNveXtEOarpDH9vyPmt3a+h0YZHf02B9O
FbpegD2J4ZwWnQwCsN1vIZVran/93mSpMsCh7o2YZk9OG7uEaxjNmgXWaoHs/s1l
rOIChG+wr1FtRB/0NTowTadSUh5+AO7mbC1sp24ybpcxGg15APo+/GU8AlbYSPPV
vSgoGe3u8lVXsJqt8WAXQoF8lsgSnrTRJxR4iKSK838+6P/4NceMq+v+12dc98eU
A/rku8TQx22Ep0v08EWF/FtbM44x7sBNC6N1oAJDUIOQIDOJ+fDxmLEAXAM50fD5
zOJI+K1JEVn233XBQTNaQE0VAlt0CiSiBj/5ARGGazvv5oLv0gh+rLQ24X+LZqGO
ysd548ePPXZqCTrUjXnHz8RyRdQQnTX6NX2hyemCierRZ3J+kQmhZwPjn/u2ONrt
TT2GN1W4SvuMwVeQGpTEYa3dwU75plwOCTICX+QXn9tQDnj665LKqBjR9DjkRbjV
t4lKcLiE73Jr4juh5mJr621TrzTozRSA/PNw1uf4ymUhK+ANJaAWyUghjRstSCDY
Ap//UPlm2mB9DdzdhzcSLMthXzxwc9cRLnZMXoviQSgY0bfTRdT9hRLUoNtCCRsi
47+vrX3PsfKGpmD1+xWR3l106Ss5Hmj0OL/p5stDPn0GzYN9MlZGu39KHuTob2eo
H+KmrMPSTu9XNLmKcNXS9ZDgh2cv9/uL1ibUrPZw3AmpDaypdGqjbsY2m6Rd5FN0
MvVP9kC0LuUQWZI4OX8tNYy4V1rWeCPFgcNn4o3BTJ0ZNoVmyEznDfhrdYt2kxay
Z/JpeMZYOOGhSmSDjPlrc5iqekfbj/kFh1t7PKIFdAOizZl2yrBfQHiq3t/jZjdc
/fDey+HdQoCjv4YtNEOEoYgNJXkXDsD8yWRrv3FKGjLnraeRPG5Ew6rVRU7vWlag
LYdQ5zwKQ8VvdBb2XFgwoM+gwvrVHBl1qd7ZY6fqElhcJGWqfn8Z1GC63k5p0WoZ
AyBS+qXyvFV4vLT33HOtLJgCcEH+goC+Z2stcnA+oTGsd1OprWsInRJlBwPT474j
AY9xpuRSQqCSU7S6GPWdklctDZ90r62SFldcjO3kp5nqaX6jKWsQTPtmfQKprk07
iOHgu84CBzQBIE3/4n20FZC+mgrWyxo9kYImODXK1SFcGPkI4nw0GjQU+pjoLTD9
5qPDTZEEX/YX4NmIXfDpmEMBhXq9ChKtJ6OkWJSaEU4HXPWmV2h9ePZtigx7aXAj
8t5fztBEZ1HJLcds/0ctNA/u2CyjCeo828gIrT7JE+FBQk86n2IC3QnUS4SPCB0m
P6V4YBsi2JTAh7mkFKoMQclZFfyaT2vh/7lhyiR7dunnp/jzKFbKX0pzkXdyquop
aeRrljbWute/lQdBlbalMrPINmnU33XKN8alFeawGsYNrkXdCNKdh9Nb1zhp91Za
zfSzNr3QCeoDJHwr9v01Qkaz02ui7+/Hp3WXmGjS5LmZRJDf4bCqw3sbPc+9BF1i
1BaS3V/Vihm7G8n37go79qt1Re412On2O0pH0MWRxrFLxwTwEn3OnM91FaenU0Cb
pwKZlywmTLW1ABKrooA1FEdZOOf/i16WBkBeutCqMd6Ps4qP0msf9ct/IozpLdxq
dmilnvyh54bDxh95/Q5ZbjRdbemmA0F9tCQHMpWXgZKbE0p1w0PP6CZ5EPxEEu7f
Lqcx7pQIGD9Izt4TCLj+qHob5NMi16tv5ibz4/ZicH3cXJ4Oflbxuup3bcrx51rk
IaQNEN84ThqTFDydYO+9t1w7n20OzwBpK6XKoje2Ze5lOBZCJMTsKC/89KUGP1N5
DtjxGCVKz7D/XPUEeSL2UFHiIYLUAuPwBuEpOHHmHkxqoh7VOLFRmFisFmI8tJw5
uNzesNvHpHjFMungMc9gfrgA0W5YmEHtQshLinUlJLCJuRIu86XVBlIozKruhLa4
sXc03LuX5RDp1lnZXuFP5H4Ab7jlaZZhhmDmoip2RTtggB2jwkM43YHwNQoVthK1
7MdUPnWSjCCHPaumyuaBtLSTWpcCofLjvGszLAi9pHL5E1XsprGoOxE+txvMoahc
gY6Ba4E7lhWfTjj7N5COGQkjk5DGNjbWcV506ZoB3nJCs2539bvYEUweM47tbaQe
hfU7N9Jalhy9reGA/t+kYNu/gp/imKOkkcl0T+FiycLQUvHXNxlUEjMjBTUvLYi1
OOAwmUbstD0XgSGy5hZXtD+oqFnAK4NmOx5P7l7EPhi19mzbboNtraDUo6tiIUrL
gLoz6pYFWcaFcwqZXwt+yNu0ItoleCCkBrqJhMAA6g8mBzLkMjfrhhLC241YfhE/
X1u+cZtHRuOgEOdUpEKjOvBfGvhIu2pnYCbv5Q6NI2bkUWflBEo2h61JzlCUbGdq
9cfPenm6krql9tm68jPQ3yitJwx7BTqWbZJR41gE34cjG+Chaqu+NCNA9VQxXMXg
8q8qpmid4Dt2vQfuDfzryxmHkghVPmCf0FPdeXxTW5frsr/TPVd6XdFsciyD0Pdj
45M2FXqkyEr2c5T5qTePIR77vX9NGdu3r+YdJo0HYwlKQBUvRAsSFhAUZHqRsMHe
dMGynEMqhHSLdmrhqn0VU6rhYSYtPISvsUfHpCoKcmtnaphsN/CKyMfEn5YeAEsz
7mGBD9SCk1GDajNXIpqrtc0+jJWGluQT0bCp0zU1bnjKbbRbm8u7HJQYl6dK7Lol
9Az8xzTv6aDRLKMIWsxVC7+DyQ4JffF+Hp6V5QvCTiq5pVDb/mZXazKhNn7ymdKZ
QMQlmhlmENeD2/0K/xrw/iwpnxK5mdjpXiYCq0kaURg5GVbWWec/yelRk/LH0ID0
cqP+ehqNyjEkSGV0rg8Ent4bkLmhFFUIexVz4oyhHiL+esBsacVzdpNZNVO7E4wU
JMvb+AUCMFSp4ZIRIATlHCO2UiNlt0gztocKc94jARa4/wwYzuDqdIsKXnv1pYKq
uOt1gQgxDon9gqjma43iH7msRCc1tJ4Xw9RLvPNIWcZiPYmu7oo69YvvcQ57pieZ
5TI7c5Wy/mRHby4MLss7ct04ydBuyDvNpVO3v7uOPI4i+4sS2QRxnsJr/NzZp2sB
Qz51URvYB5DV5iuLhbQgKB581ZmeVXWc46DaAalLm5QfLonb7D3W5MphyQCiJ1yc
0IHaLEfteZmIHLgVL/bhPc3zVv8YW5cQ3045ZQBAwdBgfRw23LPzrLXuu5wzuirQ
GvOnd8FPSxwyCrRNAMQDe/Ep7k0Hz+Y5+vYXQWSq+ahqa2ZV/R0h7Syv3z3oy8Ws
7pnst6Crp+qLV6zXhSNadO5ayVORRTD17+0XSiHQ+YDeDPvXob0B5AKnyL18rkDu
BjF0qMI62HTRSLjPSt+xyG0imwnrxL3OeyTnflTAXLk4nczOpubhLHfwNagf03L7
2pfKJft7HvBf+Jz80tt7rSzvcVprjFx/Bf0HV5W5HlQ6LiC/q4wpC66I6y4Te/TK
zMwSrvBtLqnCUrrwE17Df/0n/9cZ5DAIfQIRaJEBy3sSaSnzQOFwI1gUZiTwhsxQ
2KJzQyKcXOXQRUFzhd0bOR01bvA0k3yW5Jlk+gwJRHyUhB0Q6arEMavoRtxlWonb
7is73xaosknFheTsomg6uyfA3gxW3Q3Y1TqVUN6aXKDddJ5+rwrPNp7xoCDs6d2w
zb+5Q1Zryfxj+/Bcay7jeuzoD0qWeMk/dNqOvWujbrhzPlYLNNkw9zeec6NEiQBP
qkCQ/lNHygZNICfJXDFnMJ4FjT1BCpnh145QVvqfSGLk5BcipVHJ1Rkl6AnE/zTp
woDB4jS1a+7g+jR/rCQdq1rIGss29EQEqBtRGoS6bX2HafYH+oybJHSQbIMge61+
U3nAxN+UbSR8UAVhyyCzaFZY70buE2TQ8YxVooLfd+brTbjw4zcHsAeOq/LE2zMQ
m9z8zxUX74yHRvdhpMtwu1QNEyvKqaFf2a21B1yqSk23LdvfC63cu5TFyfWGZI1V
5EXqx67ylgxsQ5WmdX3GucmVRvzumAgG/3EudB+FM+A8UI93PhbFNRM1Ta8QAVri
Se8LN7Lxi+ZqR19X4ZEKdh6FushiIvL9u+KVgNdV/GAdtG/z/b/oyF1SHzMJ9f0M
cVEeCxEok06r7Yj2K7LJOuMUMPR2BtWGqJrd1Sor3dVXMv0JgEdzu6Rk1fkgKRqE
o2QcNhnqCO8l/guJ56xAVQFzLPXdwQDdRTa44pM80KjbelPP6/qzoIE2kbEoS8iM
IqV934Dl2ZgT85nolxV63uQE97DesZ9o/SuTrC/N+4o7jEonl6OE249ARqa68DF0
AxWcinU6sR5TM5djiPdoQaqFqIczRR2GtaxDJqCGmIZcFUiLNki3v7iMHFLDmoKQ
vx3AEVfl0DouuaeaLdNyFHdJJPN7JXb4TkOmtoGW3lJecLvTjFU8xDGkJtKRMJoN
ahjLK9NT6R+LE155yyYMETpoV/kBf8kjvhMFq01fVSsn4UmkEZFvgCIm9ejukG9A
KBwG08UwP+j5sIJiA5UilWBmp4+6Ri1V1vsu6k0+w0H3wF9i39eTCC2C+jOXo0Cd
c6f7+273Guu228ictmd6tHpSA+TsgH3sOowRzyoHi8lsWmHnMd4lWZQQRueB4rC6
3u9uyx1Xa6XtYPzE/UUEm9goKZ2lYVNgTtkbxWauTHces8zMjd0IAh+zXpPJyr5X
tf3i5eW+ctebrBpL1rk/w8J0Mz4IFvmh6aNo95ZF0pva7z9dnbgnIYEsOCYvUdft
bLNjbxAjQ+smd9V2owt1TBWSacezzNno03B2EjfjEwrq16RG/6k1Mot/smlcF3My
L7gnQ8lsboZnabwJZDxmRI48bRyAbIp6R9T7QlXSsgFXTb07gd4X7QIrUb5R8OY3
AmVUgjhRpBxVhvrc+DLWfGhq/ePT5544dshqWiC9Kn4JThPW7PyB9hs7R1NLkQxE
nO/xP6w2aGKa16NIIeGxRvTgMFayi/9Mf9K07y3BT8Yqkk3jq5ozjEdwDFWqTFMe
wozAvpBenKw7c82r2s33rCnwsRej37cIXIwVYyVN7cHR+eAFaO91XRCeiS2udupv
xa/j5035I2rLZfH1G25msTVTbtQX76wgm4I6z5QBpdlL5kPPWKGC0cc+NE6s7QFG
dTiftQiWqijRTfc1kuDkyWg8lagSOKDPoVrqyM7P+Zic2l8EhvvvLv0a9vbc485q
Pr3f1JdBqObXgWFDZTwNFTa4Qdw1/akpQbT8URf1ChM8/4gbd3YTu8OcZm0ustyV
EolhR3wXPFo1JwLiFzq7jsJEawQ8eTVN5c+XRdU9nSx1cqRm68HNdMaZk2TRhfCb
PwpQgfHHTlS3LYgIxPLGZD19AXA3eSt62lZFSRhICvXeWCVqRJoz4FFpyM6c6DRh
c2Xed0npo2CTooZZBksRwbd/0r5FNKrKsvUQlFPV5hoHzWpFWhlPhMzJToetKwLO
UBJGMRf4TkXrdwxJRKvAN189BdfGPmVDIUtmSIuG4v+7UoU4jzn722ZtIVjB5gDI
SLfkdNLIXgzajwg7iHr6agdT99WD3OqsTU1Ddk3ULQZRPdmP/UpdKaz7RG0Kmjap
A5g+p3pC/8kmfOe6VY5BDJzVytM81t/CmvTx0LZaCOHbgMq/yyEvQo+DEAhmMC+N
HqP6I0I3VgP/dBh2x0OuFXC9AuSVJakjUNRYDR/ZsO5Lvp3n7hqHYXag8kKMWkJM
VGWMdyKQlwYMtyV2o7gyeVcfARKFDBjhIVQWHvCIBp2kUem1ajqrbU3QK7wEigbE
uudHKoAnS6kUgKo9NYbdhdVgThEzwjV91WqSGcT7QCQJPXnfAS3f0w3ef14Nv2Us
nQw9LCKUKAO4LZS/EMbkAG4nkNhTnz8x4ztqNhkR5iI9oDVxKtl+2Eg4ucecila/
n+okuJ97zGiLiErEykipUWxjdNpO3xFUBVJCGwG/xCjQIUwPSODtW9eIE2gSP/oU
BZ9rgtiU7zzTccTuyZ4vPlD3JIPg/Wb9uK/KDQR6IXeoxpnkvCg1y/vSnML139Fp
n16q9RHgagkIMHksOb8NUVWngaowMXAdz/CQM662E+gX1SeVwsCxe3IKZOT5NhVY
3y0kyBVObPHf+uMmYre0k68lCEv2kvtToGlBMN5rxBQPdm+72aWpM6dUT0QBIwYC
LMUc27cYYeXJUj2EBa2ieLS/jVvoyqpoojWbTcRB9+RpcMBwug6E3cDYrS0BsYGP
Q0eg3yem0uOF0xf8nUzFEg2lQJWi2tMCzODUDLEjGlNSHZhfyzbSSjTsykovupg6
HjjD2ev9gxbhw2v9xfn1emfE3G9khuGvtKpncYIzKtZ8q32PdAiMETFUrupxwU1D
LsUVQmfP4mPcj70t543Rdt7ivHU3606yN7AXOP9CFl+rnTt/b7tbdVB3XShjwKOP
3zEmfRYMPiu0Vq5pt+8LV0glyl3p7Aejsob99iWlwdQT53ofZwRXYgoLxqKlQ8O+
U5tKu67SbPeRrBHygXy30aUWMa1VN2RK6GmDx4pLRPVtjhnKFjboM5PU2YVbb/KC
JvyVj6Z04VmFuNO90RVNCJt12K9hMH1NSL1yPUXNGxaeyapINdityXfIliOgROW9
edhDwd+Q7PNkj54EcazqRhc5OfFQAA8mABAa0Sqyh8BioxYzUXyBkC7/xeFvIHyW
yx6Lxi8CJ2I5KxzxySMOF2uRfyCGjwYPcd6Qc/Nh6H77SiPgWDYX0KWYHXy0kUmU
CIV8AiTfsu+GrqvDssDpwPqW25+C8dVQibLU6mCdNAaJZFcwTFY6hyERR7QBA6gv
QVHYO0NqMlRsQ1ItD9c/wJeshoYID1x8+0eqtelEa/tCz4Mxg0jl/qvWWmMl0Nw0
59Ueo0aNSAoBSro1W++3mimJ0BszUHPnAbXNrz9dvX2QhwwaJ5jS0pmUCgrnNY9q
pFGuMqtkeOAMnLGx0nwCBGt9VdFWGpHVcmZ3JZ3AjQP3s7Ta6o2ps4DPZ0IHgac4
fCIExWO1D9ZXjClgQu0Glzd1BNen0/50SYw3sPXDn8gEsCwh+hPYxP+df7iNU2lw
NTCRwdw6WCObbyH/BBIUor7Nn8Lzx3Ka8fxVP2svamOMsIu5+GFd6/4ZNAsOKksy
Q8AUePeL4ZkHWGFBYZ38CuMLbF/tX1CCoXRDnOg76EEaU6A8y+Im+cfV/veXObRI
JEn1VbtkaZty4j3O12EPDFCvneuxuTESIrJ7Y0hbxo2M3wxlDwn8Aqrszwiun1Xu
P3A+MIJYvKVT3Ab6yq9AYtIwhDFwUtiXWuS0RotqNgzOVaEvI+HkEapDz8s/aMsV
3fDedjlYl2ywIyWmNIst3evf4e7j4vAyeilUC3IJngPn/mww2iqRb5e8zdt45WiZ
UzmjtZlBxZN6phhursarF9sSZFZtEZp+1CEc6JxNxM+7lRcMlorMUHa300p5yBsM
w/T26eRiTy0wUd8zh0KTRgimKP3B3MBImaqLGwEYraPgw1cmnrPdiqy+AE5sYgFb
gAMYEc+iPMPsIVGgfTuRuo9VHYO2LMc71PbLIlelUqYX+GrLpSDtm39hC5H5CneA
7AGF4+YEMlQNflNigIyZmO0FyWN/Rj1HqgHEhV1wngz3I8MsA+9e6r+cP1xtABcR
UDWwf3cTFNmEXG5QBnfmnyRV8Uu+pqaWsE1wCgg6X9uROSYSTjLeebrPf+bNWEG8
/ujziMUvnROQaHjCHvjgZfEq2eWjGFy+6sDlrIUYpe/W3GQRtWSCzAvYG9dfJyH6
JXwX1/V4PgDiA28OdShsas0+M8+hVt2Ylr4r+P2nP6IXGFJxQQZgdH6EuVWvbqCv
MAy9mTWVHXsJ5E7VVyNP+JeJ39Zd9qpLcA66ehKEfok2f+dKZXfXgWgblEIkAlhq
D5adDACaMHIDovrgJFWUYBzymdqM0xzpD8p2ITbeuW4y/C9qeNzK0/VkszLqqbUk
nSyjDAHlFd6BDFcG06h7BJzjjQEO+GytVxhYnLu9K8hxjEOIAoHLVGKrXiyEg+6E
XGwyZ4dET7acBdqSJTXjOuUcJUC5f3dSlF7xzsz42aU0A5mAeOp9r49w1XlWnLC1
APtO0/QM/wa7/4RNgIZEBXkBe87ilbEMAGDCjihRugy4xeR7Pn4jtw0/lX/u1uYh
VktexFJePaYvx+DU+FhVCe8zW+AE+pt6+YcWrvrdqYbcOtDfQnDUvl0eBEiv+oZz
hF0eOAEYHoaQ0ny3lasFNqCSc2Ar4UHtYa1J1YK3etgBThx5INYLnaCqsul9FZ7B
be2BwFMYDWJezrOdeautrZnIw5ctTKWgXgtNiwQ6jtJtx9heHW6outIdKy+51ttc
wZ6W7SvWAv+ZxPmpB97AdtSQKjvzFvXgwSBL6LgDx86IeAU3FNu+MZg3lSrjR0OH
wO8Ydnjlt2MmqO/T679JdbnZokMUnF2Bv73jhVj74GyeBjZD7rb4duFDzmUMvq3P
g68v8eH4xPLWWHH51oOnqoh+NHNPmbLPusRxOgCpGMjILzt5kNYD3bzoWzdtiQOP
rodk6ERnchUbpXTA//4P4rbscG0DL+0GgipJWNRbWDwlrccPrK16vN3FfmOJvxaT
AL+NUjniiliED0kOTfnvZxsd7szosC+lqhWfCSJynU4UyCjYxYyP08ovVpd58mQW
f7kgKVy8/nJnjy0xM5Jr5joO5SxE0IuQJ4ve55QYWV+pXrU3IylfltvyFruWNDT5
ump2qBqrbSDIIYDrWi8IaJaWKTU1S/huE9ajvYu3hwytpZj92RO2/E0lFm9OB45p
jOc/3hf+SABAhcNeEum5Tokl8VA5YNpqRF+CSQI1piRDOA2OT7dR/xbQq6P6ne2g
AHSk6beOhukgOL+wVyF+vLGQdzJprpZOlKw1YlcXVrJS6v2XhUR1qABIRHYGCIdL
p+meXTXi/ht0KVorBk8bHcVH2g6qhkulYqky8SWfS8iU3Vi9tQgizSdvYae+JbQS
sgT8g0QLhjMpoG0nwbCM3nksK9nDwKLuKKaEEnb7mJ7PHybdSEDmvKsKopI/n61+
JNrfQ747qIMbGsJonBI965MbVRPxXJolj8DDxgjZBbARVnqYU30gM5+0xzocKzg8
eesV5fTgnbH/BP77W3Bvao9HFaPUE50A+QdHgNTF96/q17cR9jW9cp0LnTQf4Rav
njjhOrI+s2RCgfQGDGq0J9iyDNS4iXOziyrELHTzwFqubU5hEK509EYM84RHDLwp
7S7Ar+W4soumJwn4b00FPrho1gYGCFEj6RsbSFU+BArLZF37o1eOKF8h0++W/4kR
AEBSB6568ZfBYpivz7uj50JiGgs3X8u7U4N2CAjSh8PHA4oMA0wv2LAweJpTS46W
fNihF5voiG7Uzi+P/BXO1fAyXOwUWbhR0yPh+fJQ5D4uIP/FZVvcITBMkkdthEw7
BoNs8HqkcSqNB8bgIrObjKAqLwSDjkqqOCyVmgRicHtRTf/zZyf5hNBRDk38UZNL
mh9e9+gpzkaBhMJBd+3tFCB1DAWKFvR9MyqsnVpbYjMJCM4WbUcTEZijNUvV/sk/
rR4AvbuNtEmIo5bF6QIq6lHglnYIaaVdVR9/LfubX357hYmw19YzaYYHI0F9Rr+8
NHl8SD6bWXOW4lXVSf1iKhoOix9ZnZqIqnESOKreBuESTyhH6rbqVnJwtw873xGV
9ieOQQOeS3QWGElw6YrmFX0ecQwsiRUHi0HoqhTsTyCpAXObcn1egt6623NxxYzO
1do6bMbHfYvkthH9L7sqLfPLEFWE2elZmdMHBWeUfdzskwHnbEav+FBCaWr9MnIO
bPow441ky8O/B48cMNx9nFvCpu0HzQG4Frkovt0BK18laYc+5p/mOSikPde7v73C
0yZfknp4fuUqaLgxFbRBVoY8ZSec+KwuVoq8622OuCG3Hoz++3HrQNV+RjmXFEtY
fpsS9ZQpLeIQD52wetkREYrwJfhLDcF8Y7FIC6kBfsy8iyFbn/+qMvF1yxcv63hi
9EBhHusyqcuv2ZRuNPyb4RSVf6mx0RuoXKVQhXNb3kyWripOZRT4pHwOB35GvuWB
OoDJBzhf0mAX+xCkkzbMXoGnEZcVCZGrVpW4fOfyY688jwg2qMxdq6beO8HVNoCu
FkuruyuH4QXs1B1Z3BktSQ+AY/CNV5k1b+Y0YBLMgdUUdl3otQFJwQjdN+bC+btW
Lpl0p+krtGBVY0eAyu+d2oQsT9DFcNzVE1C76IHjOC8g5l/II2HGFfA7RhFG28uL
7Eue8UYJOyxq9L9teq8LiV4xY4CYohtw+8IgPOOaDU9Mrmn5pURkbUJsW+LaKdSb
QZeLZB8kmly3EVpJBBJtw3ac5gzcfVNvtU5RU9/3RXPbljAcsHQZ74U8l/7qvyOc
s8OXXLYLJCOCKsOULeiQER1nQXOHOeWfTYPBpiTlZsWiHzwxP/z3d7c75YQE2Toz
sUQ8Lxn5K1vrQdUHngQkqvvAcV2DKvD5TYVrF6D18qPUj13OtJ0DE00gb3F32hzA
F7crInWXj/rEcZP2XcfeKnfBWjaA3Q8qs8IAwy20mzmpBFr9Yo+jvIGDEwu+aR8Z
97BckhX3d6SOJWEEhjOAiHnT5out+itkLyeKrVcKi+H9LUojnxltxqo9fwbLfdo7
yl8yZ1c2XxMGKDo/sdlNNbGQdJnblVEZ3Ys+TfmelHHwi47TIhU8zwW94Gsm6Hv1
i9C3y/DclpqqYraTt26Bo4y5V4xSF8OV1WmJXOipOYuHUWWL0pja8ut56uOJf/6Y
oP7p55ON64ExtDXigRvFIRa2v7AZ+1lr/ZOmYjwKfrySOBWYooYxyKmMO477J0oO
rWD10HuOQKE7TLD6T/2YuT/46ToBfI5fSTmgx8CeNCFcZ7FKtn8aRbgXMRgakPTJ
JDGTVkbPUN0MLwBhsqS0RrG4/pyw75QZDszn6T/YtYdbv3a7PbsyT/XMtezCAGPH
VsjxCbA/i6xUwFK0dddkVqwNsgYuQbw8WEyCs4oHgJnuzoG9CmJ3g3YxvwjnNfRz
z9+SdpxTu9cE4s6oXdSh47HZFVXZ9LCr1GI7+nV4BMAS2Ais8rJkKtR8f3n62Z1W
9ffBOHmaQ9V/NEVYZZUmzM4wASy+Pw/oxJ8n2X+gFjbAhQSMLc0ZiYA+6eL1X0XV
rrfqFvfwVuzLGw37nu1u9aSgzMtxhbPA+yk2bGjoodCGmH1a/hrYBTGR/kSybByL
n30j6akt5XzQyvCaPpL8PT+4CgiD1h/tisWU/8it2mMYhlz3T1cyw5vEj5c1Cdic
s1HbrA/09Tq9hTpCNKsNq+c6GjIBW2O99IE+8OIWYoWwhfeRQW14M4hi2zxpVsPx
BHWmuc7fusb2cJbyAl9fpQhXT88p8AeSIIHT/FEgZs9MaDO6j1ni2Hg9JlWeX3tU
F84jjIcaAJwlt0fHtkeoi+lfQKBqdqPbCRMsSQvorexiPwKtRPaLEBalzP2r4XeJ
Zfro6YhMwlmSje8pLSJ0nftW1IwYTOGbxbPHpKfTH/X2QIFI1MiTZEQLMcs+jRH0
MaZMffLurrAdsakJT4zKm4JLojNDAw58GWtFyEHUk/PPiUvr4NOur+7myu/FalvH
d3DhfQ/C2TdqrcnM8G0oBCD+2pnqQki/h6+V9QlcIUASI6OaTLK+a1BrQCx4gnZ1
r9xPXhQXD5+XHsBxGLzDLHMwNAxOl3d1VbVjRHqjkzwISxGKSR9M/qj3eZVv+hH8
L/MIphXehL47lVTqXFbD9HcLmjtWKxfsyd6yzaemEWnYGGMXVvBbibonmmt10Qgr
YfKHbIvuWAnr9meQcHKYmrXd7QWLA9ZQb42o2MC+goWvmLL85ljAaODTTYtZfNAd
uypYh+Tsn0pym8yJ6woiaZuGz8Ass3uQFb9xS328lc1s6UlV747m9qsuueKZXXPf
qjodZVMXExTCG+QeexrIyHvDHsBOaYakjgWSzS25O4r43qSXXD09+iptqnz8MJAY
MoP660e8ZtRPjL/0yvDEIiQikIZzrFPulUVoQq7wBnWRraJWkLxDyfOod5IV/kWN
CQ9d3Pa7xTdKH1zF6ZCd8qaKlqNVdZGt+UXt7jGM9JE6XDpP+P+PGPpA3bzUCAW3
5rIfHYfRkXLUK0cqoOSl9zc+K9iv3gIdIWuzJoBM22zAUj9Ik1K1/cGTHLua5RCp
w9aawG7kjQ0YNhcEk+snENts+FSwnOpQvJrjfhc+RXL1Z4JvWABiXVIBKz+9gpAy
q0eWQQxhyd9TSTaN5SB1Ap02rQCZWmZHzkK2iAVCPRHt+vRItOvd9+Q8MUE0lycV
VTkgXf/npOi3jyNYr5vsq2H2DL9hhj2VQalnLUbNHnZR3JPE0gTzGED+h71IeJ6s
rDm2blEruPTDVdnP+YIqRhZuUxEUjLxVvZo40jfZCCuVErG8FSBz4h8R1bk0+5qY
5+F6DKzdoFMrIj5MLAgXrFE7PcDy8Om6oiXHq6n7XsrX+nGunrz0vyRJ7SmUQi9K
Xb6L8AykzNrV4pOwnh2DoKQlXEZIIpajuPZfwLP3BxOgz4zClTHgos90O4sG/cFH
3z2xTcQMaPs/vXFH7/7TSL+j9aNACLJFijFBQDsU1lNFpnGK/XHqXBjpbkUrvNnH
1hd2m1HWGQU9xiNjnQj5BjMiO7oSDflP90c0V1jI/RC7NQCRS5DhGGVPlmgiYg6o
lqIM8kfIYXIuxF9eS/3mjKcVTrIM0uoAJHKCyRGQGi5rTO11VvZ/yHDk4h+xpPcv
YiM96amqErz4vdy/Ok3F8G/HjeyFCz+4UndNBk9AQEZE+cuWwo39EaQeFle9e49r
6VEohqGmG2PaAD63Q0rnDZCRcQ28v8pxVyLQC/hsUmxg4nP1FgItvqIxlFzOAVqw
d14RITi3RG7S9f3vbFFQdRYrdMNdTEwCAxBlNooSfDeikPhFrwm8WeJW8QZmLv7m
F4GpIWMIbXCQq4ZLbVw2spCSOfZxCHYfdrV7VAh8o3yqm88nlM0dGR5Eq6AbbZ2w
BDDdSVyLh8pjjWYLiPmQ1nNE9jYWM8JFWgCzuN+vMvC+JEI8ls1Ypu9DWM3+w2D1
5knJ5kqB6iDFRdGn9uWkuHsXgxkmcuf0m/mbhLxRMlXcIVfADrpDMx8ifwaoyfee
7e+NMA6JTaq6IBmFV5/CQhw2JiKXt029hMjpgURxIs16tu4ujHPtnZszpz9T5E/3
ZNgwR+KcGZpsuwKyuPTECb3pw9Gyo92HcYMlCMeuZp4DUDRosAOxQ9itg2cHmEL8
HjJtHUexGJcQ9atcSFwyXvBWMHRc0J3Q8QsdaKJrTsS90XQCb7EeDnE6oNeItL8p
TU5RaZEmL8eDlySkABeN/fkWJ5z2VHCmagq3GVuc/ZN+CKzj25KO3mEV8WkQO1yW
FWMcgQgkCHkPm4vgjGIdl3Mv18TW1Ckbo4949cKAiCpPXcItpCZvZme1qnSy2nBw
KPexvY/eV8946ZTt55cTOppQte7pRnKB4+XmnaMRM+hLxwXqsb1ZR4aEYbkJ7q0V
J3bdgMQ6EABfKE1NB2Ewfh2FaGf5ueYT1zLeUd7+NlwkabP6fpn6R9/UuVqb6jE9
rgfzTIck6qP0y6VGB1moeleYmJdIAYayczDujekZAk+2qu15sGTrjhTrKj+/w4Ah
8+dd1E7/dAkrIyGZJ89oIXTqqjnwtnDjFVeqRcZyV7bx/mI4p/adCntb8kIl8SGX
gXNxcUVLbQFiern5rE2c7MWpM2pOyTsC96VoV90NLrjraKfMizrzDXq8AHNN5vTG
M4QFbeiECShwLcYIdfKZgWCanT3wqvO0NOz8da7lI5qMdMauOE8f9hUUeeNMuKrJ
e+C+wq2SfIYbAvKMII7itHwqHjL4mYfjHVWjDRGrXbr23bohS+Oe8VrcHUMX9YMD
1JhBIJVQgdrD/alN8jUXppzVEPVoUBW3raCpQVa7Z92VWsf0jllST0yz0k3LymRf
1uZQg7RWakNQhrhIqDOJbpKwIDGLUmsd4Mn7QlfoWs3iF+Ruu8yV+UYu4S5/WyKp
+4Gh7CAfozctxuruoMhvrzQhoUtAznMHXqT+htLRiJllMKMSYPiO/LKWISeIfIWR
Zth9upuRStNFfi5EbHEMD9eIohdDkge4qBxR2gEwe2UVquiUBvZusOO283tHy6OL
j3Sv7sVt7RhP0yeei0OLiaeP/gc1Rapm3lFuW+dvQQ1LFpw0fj/1jQwsvkYciJ5y
sRwSP+82430D34WyCbmKy1UdA6FQTh0ex7k9PVpYO3Mxp/j+gVDjmgaM2v5xUz8C
qBtYQwbIVSy+lBvCLHOSWIF9zJ9sM1G3mFWwR7OhNBJs8zgJIZUI9lk1gvX2Dgdc
B8piQ1r1jSx/r4DxYbwRGQkBRr3Copx6tkYZH/66JPi2SoBlyDi+dgW6DClivK+z
n8Wr035/becLobaxCD2qadQ4gjJOgneyxUPRrd+cfeYxAZh79XVCxkCb4kE44/ht
+GQmL2DE5EB7z1DpQf4cRWZbnMtEJIspdR4i5XSPNsedfCFYCKgI7YaycoXxjKQD
qt+bJ4nlC8/4CY0u7N3EGCEh0pQUDFoN21xcE9JjwsIwjeofAuWpjkHo2mnjuUvu
P6n0oOqf2PE8h6XnVnN+E2wTx8cuIyE+lieiFNDSPvC5Z3djm6HZMPHsjMIK91zS
C7NUYJPTzFzzZnjL1P9aDvtHbqYoh/SEXF0PEIZBdgdMywcejQ1uZaRxmiIk1QPP
SH8e2vbKgT/G5QVDT12e156IfZ0pt3bIltrrPnFFRw1L10qRXKFkqEAdaJqA5P50
aTN/NaUfhKYEFRuleNt/maF07hSJCG/dFZOfBAD3P+ZT2tfClcSgVidG1/BAB3Nt
sclxqrVSNhAQSW9UwGqd3kDvhdzRLmcvnXBJKT/5vaPab79oqvGn8+dSvKTXUzdz
wC6zDB2tb3AO16RqZ7QA/RS0k+Ulyh0TI2ZCpF6r1bpdQdanLtQwxB+/ifpKF3Lr
gOx6j1oal56JGkA9yp15bxzbqu2MjeJpcAwsavxZqjgh6XZ3NyZFKbdx0WtVmfgE
dNHcnvUM+r53T2JJurak1iKca7dx5yRnG3XtBV7WOfWLRPadXvCxTSD6qS4/uKKf
pxfU+nd5R63AP7dh3+/wgroStxob7hXsV66oqiG5/vT9sz8ozC4cCtHDsdyuEM/4
9f0fHcK94GMok64aIL13ASMtTt3XnVHJdLXe8ARSnH1t6OeX1M95aGaL/6UgeKWw
xM/W516ALj231h0OmyDL9YIHPE/eVd3lulrb9etpRF3cMv/HUr+PNIauXjgwS36u
JpImNaRIOrAzMk5GcVVdX8ouFZh9IS6iJzT7KeYRjs+C9ateMxAtiTsg7JVSdmca
PRBD3sSWGIZbe1hIHCpAapy+mgftwBwBvhT8U9Vs7SEWNu92aWgfQvO/vJ4NkK07
nOK2WMcF0sCuYqzPXNi1cIg/prxZOxyNxYXKqbcZal/8JROJup0NVihGKXxnINha
ZumWd65k2HcaJOgjrkrYI6fQeQQ8G5J/6y/7D3kT0AbF06Vi+5Pt2PT/0xWJRgfo
+2jF6c1oig8wEGsy5YWWysle6yJYGlZK7Kw5bidD3fhhRnKVN7alXh48BMVOPsUr
uBYyU6MS4M3jbS4r2oo3O9HbD28m6qG+zVKCE9HYS0bISrsC8zeywv1YltjzvWi/
Hh2o9zJ2+j2fjtSE1wjrOAAhiQaSgdBjwlAwbqDN/MlU+/OmbRi2dADp2X1gel/k
y2mNbk/vv99Rgtzk64IAASRMNJoGCA9o7nRTCylcFiLEJJ/fKqkGUhVU4+cUH30b
+zj42cukJ8LM/xXH3gS6s3lGSoeNv/hESy9N+MxxIZKkBhmTQXLJInXQjD4TQ0i5
cO1XdVdlAc+yt9ur+x3neRX1N7vr1DxFxMNfDI19PS0aPrQW5wx36rdTvkb/ZvVY
WpdsXTmSng82WcA/FX30w1SzE9mDhYBUorjItxtSdUfziONHH6CGUPrVp1I0WZ6y
jHEQMS161v+CvyUtxsqA98CMPJ2gZWtj+Hs/bf7uhb05S7iB3h3ZmhbKC853l0jJ
Ph+7NHNt5Hvlik/t+Rs/eoHPYX9bjMlvOeD6O9xWMFPSSH15u8zy8xHL2+cEsjP2
k1W2MVY4eVxlPtvZyw9Co0oHBJYCYEeb2tsUcrK5oZh5FJe8hjOXJ8QffjQsxysU
veW/uQSIfT3jNpVDyEDOafLMZKVevUK0aqf4/xNzcm7Q56BSR1rYqysNi+M8DQBA
vqAlpvqfoGQtohCRb4tO2tXIEZ/Z/qV9RKuh26bTMcjHZTiN43vgPNGLYXlN23k8
P6n1cwNGxUePpLyR3cBj8XEer7K4Xml/rBo66wyxuSZyWmP+Z9ZnOyzxF9I9xBvh
tTCHtmhB7kVR7SUand1mWK2r3zKDdN40JuJA3EMJKShCpls7a+YP+xhDCD9LR/h8
NhaU/1741xCYimzs1zRt4C1Z6RDcDAL7rlFRBwftJhgQd+mOSuCNtkrrzW+LEwuf
x/OkwjfXojPFP5TSDV+EhjZWepb7tKcleX2yHc3/gVtTR2l0DAmVuCbOQiMcBI1K
Tcgf0m6nuBz8HerMhVmdr7js353OmhOxaoRUAK156YCDrwfwpD0EUPOKMbWJPIkJ
XLynfEVanGRGM7Dg5HX0au+4au2daR1ShRzbSZbNst7pEUItbgDbUg3z5XioTsDe
0bl7bXxBjggk4pRltX53hq+gW+3zH2VJmd0ofsQ25Dlo+T0AHJknggLmCgBJ2Bei
jljcLqzDldsISX9FNCPjwoSi+R+xFXKwnWrQ3Of5Z0lPC2p3U4bWM/GPXEca9iav
ko9nyLhr7JwQOmApLaEirXTdPjuxHYtOcsbImCCIeBh+ukP7Od43dMxCJAfE48DE
zOyNdhGJOEmrz45nK6c/oeJrsfnZI7Le0WNrn1ku5JCKcs0lwZmvrAdyVRApTZGx
TGObWP3ED/Ra3LWH/lIqubBsaReJ6gXkWIoDvv35/7poT1cQSBicXPcPk8s4cDFX
q5otFGFqAlDt6yj1TqnBYYFoT7q5IwKjkvjH/0/rzlfw43Is4lvBJpzHQx0+fCQO
qiTGuFoW20HS3DwaV2ih6YBYLnUuM41WEFFSBXrmjMgB6DUANcCRVttV7qogDJ9f
wMLGRgLiYP4xiFIcFNSiEsk+3j8QnzrAfipOboeoKgcO1MlXroJeLBUrjIxcf/hX
2Bn67j1l/Kym8yxPMY3X8BC9Xl2qkAZUbYj5LZrzyyY7Ab+/QU45G8GXEXtr47VR
GNdwCGxeXBKcyYbzEOVBFHvRJaStUq6EnVoJxDqocTFtz6aUZY3QFJoxyAGth9rk
bzQ7AaEPmJsYzgQdT4+WVliVl2MKPYSqOsmhs7HAm6EYmf65zCOVvV0kj10D3ygv
uVx1B2LkbILgTP5+qPphsMsFTi4bSqDm+O17bMQwd8EQXGT80/2vtxkfj3jvCze0
h3X0eT7J5ROEA9BOuBgsBjSSZs/QmqJI4lWhKiI6fYkRy19XwGrUMZLj+lDCza33
o6/7Ds8VXf9972Ta1QFTKB4cKUxtqsk273pCbWrg1WYyRTq5cpPauYJSRXUK5Coo
Jxn0fxphoTqnHP/mukctyNZM4O8La1LvXMJdux8KGhL7YRg3GgsrHKAZ1ipEzOce
s7wvdaVw85lA7wDKp/DKaUeu8u9+nBauXC8+vRkX/q2a7acVCkr0JlzSqPDvnPZo
kBKLnKd1b6izjQ5GrBeJ5c5shv24yydBrOLnHK2vS4wSZKbZbh3QFC0NlvmK1vBT
QQ4wV5ZSSGzdGELbtQIoCV4KKEvK2MuEwmbF+aBcFWVAVckfy6ksZzoCl1bG1uMg
0cVF5SrHUipcq110ktr1W9Jq9IMWXihOR9p4AmNSKYXmFRl11p3tBUDO1MD4rj9s
nr19sZ3m7DL9VFGmU3sH9ErmuX4wJz1hKIfKwS7JcNxY/d2cT1pcS8fBltdWzqa7
3H0LcC2o6IlSKXnkLfiv8FmjsawXlM7uYfdU9PJnzJBUeoz4srOmX98oVmIiVa07
ZXoMK2hZ/QUGjx2GXKEwBH+Ve+8bZLuPkhSfA6x1wzeXhpOkOu/65ECPxqj+jWdc
L33g6yJTtDrWDpvWdbTiiDNKmtwx+2E8Iyb976dBMkhoIpqiQfyk4ys/NwaIOcD9
H19P1KxAWg0i6xm/8nHHqqrtVzE11gONQZLuUE0ZdFWDSbeyuwTB7g+UQTHnn4ee
x8JpBnkyK/PeI+4ug8ZHdLUDglWID70kRVG1VIWQ4Z4yDaRRIrtO/Ja4BJQKQgUf
T/ZRMj7VYVeXkyS0O9ldxVsunUM40153HvR1Z2/Om2MYlfzJB/GJsUPlZDWQ5UAl
cailxgQNvxFtPEvPmlJphXlzN9IkUwS8XKVOS1LnULjWvfbTAfepB6k5IeKWC1EA
8rSwJJj9/T/bnN2oR/lyN0v4I+Tjf6M8LWI+RTUdXX/vsi1t+Lb3xJ5h6IRCFLje
HnsZLpWCqXMhrcTk34IMvPwXdtfVivsQI8D2D8xdYsZpEF266/HT3/SMZ2kB9gWM
9HIth0bojm/7iA2P87Ffd2bbRe5uR6rDEFEcYkUPpqjyFdTmGNZa5jTd0nG6AuYH
4DxV5OhoUOLMkWHBj5zOC+dYud30NBZ/WCqdc7knVX1GYcl/PWO19KEIVE3EHVb6
ODid9ORncjq1ABGKr/nuFl7wzjEopYTduMthq+LoXWJh12daGe/GESyoWfj1JOLP
Ahi84EsdvHVeBqMgqfJEXsNdSkY15fmH4aLe9nkucmeki5hdiNh4fRPWaorr8JNj
+zGSdLl30lvz15p5Ar0MjGCVQo6gGJVVOB88goqlsR1r57i5PG6iWzJRGGJ6xNLs
HKQgnh/hhGK1maL+w0QAaJH8WTmiIHQLfs6qYrCw+oIWEDu8XYTzMGEMkXMMml6q
CAr3mInKLxDxF6xUmb1TDotJy67py/UivwnIiF8ajd1by20WRFaTg1x3EYX7/FUw
8YM8EzipU3TvuSl00jjsS8eYt61g8UXsgto/ocDcCa9JdEGdN+m7QpuGI400P9Cn
2t2iabrXNoSrEyrggmuZ56JNeEo6OOfjN0OyJIB5KKapnzH7i1NMponb53x+FZXt
PDwZWbTx9CZkfqQ64bF9/gRK+M3EJ1m5XZMyokUFpIJmPMPkz6Zbzr6ptmJ7yKqd
0VMEnJbkh0dAmbW8Hyz/tIr/9whWRuvZiNpCnJ2TwQPugsV4+e4J+GSpOwYMFZ44
pzAg8apki2tADVhNYCqT2rPD8hkVCSVuRXsksAQXTeD45bfm+hbKdIoMJTuP9kva
E/VwVN3zbw8cfanG8UDI8e9ZVYFshHYvoBfTfvTk/CGqwts8VUjh/sjPmCHw5J8X
1gJ8vgBbkDF4hoUzouDgNw/KY2R64NLzZ4IPErpiSnWIXCSnQ4tc6KpTvBfML9+D
N8wt7vgZdMN5xK/lXgYJVBUEpWoWe21wPXNa4fao0d4ldW0gTutV6+USXb3+owqT
Xe0g19gJpD4OosZnoC+beQ7TfJnWZcsNQvFc0XxAzoyUFRSxWq//cr0utLRf4Jly
kmZAqqab63tQLwj2b5K7minSXpe8UbNILXkgAbt3l6CXVcy8L37Cr59zUXTKxtU1
l5ZOXPC9Evxi1B3UCFGUS4gwu5xvTExZgcicbBcwzjlTRu2SgHhq3F4TLyKYVl3x
Y+Gi+l8xFRHKEBmacOOgMWfQeVlLxbmQRH5xlVbTKNcD+8K69GEqrUbkZSLzKOAJ
Pg4egv+Qi9/ejdTPLOPv8uHnz7gidZ1ETfa8OrbrjYMbtNMQrQziNHwJ+uTmKa63
Yh1wYi0w9xY+8xii6js3s4Af599JIpVb7Kb9FYT9N9twLbcYdzKj0JNjKB+ctLRz
cPMHMp4HlfOX3fURQFtvJWv2V3RDPqLmKKzxuGhCWWEtfXnBbuwznuafoi4gIrW0
gA7ArT2KyCFTurmUKorhDpvnV9DAOoiAMDtYjHezG00gnrNv7D81WBLx4Jf2M0Iz
m3yHV2z6YD84a1hydFJt2Tzlzclr6vJ6SzUx0g1+UQCydglWyshjZ3OTdLvDuD5q
B0k0ds+Yr+TZELkKIdn87EUMAvWvfVRPzMkyza3XjK+OJJtSSkFEaawcWcQ9tl4j
F50Nq5fpxvCYyiucWY3J337SCQ/dRoVXjrvwO9iFq5O5FNf114BfCoyPHPV2vvrY
9AIGSeuM/auZE/Hg//SKXsRXZx3yc+b+/dVFCDXNv3nQ9wPtT+2Thh8kAV2TieId
UwqsCoMQ10inLfydXGjxliKezP89Tqm03KR+UZ2r6jDxP9lg/PrYUKRMZV5Qs6u4
qO8fPd2KZobdsGKQh8bkLr0qE+tzH5Cl6JCuMB6gLPKu3BnZ3PVyVuXABoLUG2iM
fjFv9gHB71SR/nGnzRIHZ/6X9O1HI7gLstpdnpAkVFkHEk2jwX1+uDArgG6FHxjp
G0agsQeai0dUeMRKDK/jEu6kUQncefujTFGRN4Ca/XzRQ7nO8lrs2ge+JUSax/Y0
kxG8U6K22oC2RPLjM4/s/GK9BBZQ31fxhgr6Qz3YmVsfeqbNdaadFfs2fFEFkcyZ
F4KiQZLbWPLdtSvrKakGAIaK4oYIRICcsUmD2WoRsh7K0xRxkQI0mdLzHJkphRxv
0oFcAtCPvtfc1lITDNzF1lY6gtzuW7VYjAfB2XXufEoxkaPCEwzrX5TY+BgTUs9c
A+cnEdv0BkPL8CzMtNVifMcMGJ4ujfiLS4rOSJBOwD6tlS4dqwRLkw2Q2+fRPsts
0mHTkjFXKvZYwAgL24aSMK+MNocmIaZVnNKCDsNv32VfDQgbvpgQDKZxKatFJRh/
PJpSz3sDdB/S+bee/W+/vC77yRciVNYmM2d8mgNwuFY0uC0oGobgE8MWDKp/tc27
ABlwYh8dTFxRlsZwKhfCFJXGjgg/C+Q1vZ95bOnjudURjxqqtq0+RZOgSIKfCMx8
aX1nMZ4oid0tQfjODZutJTVb15vVrJfPZP2vic01Pnyc5FS9jWDh6T6FvnMxX8BV
IB3tNFQXX8MtoE1ITC5J9AF4K8WBFezL4WuzePzLPMR1BcXqUAIzon/dkiy9MA6a
qEGM9q/qdl3soK1pxeKcdr42k3WPVhfs9xaV5yCeTkIW/zXvr1F6d7GUZ19a9+/r
tAAixb0TBcXODDkAG/45A4vJceZKj0gXO4G7RtFfgh11pzT3FM4stownmFmUob7L
vhBjp1J94SqwbHua/r0ZaWfAdgfjlO0XkespXL9+Ku8AaqMxET8VR3fQOFJWjgDj
U1o9e9I/1srCAUg2/JoFOT6Joyp90HSCg+IXtQpF/5o1VLV64UcvsrOS1oSC505P
fegVM5m8FoLrZcYKSFDQf/IayqNQqBueCOtGiD6NrGn7/oYHcvvtp94NY83kaJFn
j815uWlY36VeuoFNuZFTpRCsBnYgznXPvPHohzse+BBfllX4/jtIt7BhvnlYxAqx
8irEexlvqR03hOr/YCQkJdUTaXwk13Dba4u702QEh8TXNAg4rg8InWIu1XotOp/u
gHXK6QV7uT9cIuBJlhSBxyMTdbZ5N/i0KlLXNHQowt0bWxQn7MD8bsdq0xoGCH2K
yzF0CeEsdIV4zg+mqnf6v7J2YuqgLMTauwWFcuNZQDGV1wlh3HG/0G/ppGFfYAfu
8NBEOfovsSDO6kCEFqipL8rZL/j6guit7kGH4eNXFA1EMW3Lujrl8dEvWugAnzg1
A2DAWpWAb5nNHRlmHXQduFiINbfFCI6cGIOZvFqzL5pY/PgOZzE81eqtMcQ5W6zS
5ISPjuefYX8L9geyVn/DhF4BABZKRjqBwYKcTtD0X6sK2gYFRdp+MTehCi/Ebqlw
t4qu9tlHrr/vOy5QfczW2ZM4WO7X0MyxFJ0pVNlxgb8bChPxiSkaShJHB9E2N1ES
IE7cZEk8/J2f6Ppt6Wa8Lh5LjI3lVjoVJ1zY/rNcFmYu91hx/x1WUs/k8AwGQC2p
KvJ4gvaIyCvo6lAh0mg2pzuD6UIUur40IsRyI4L7wSMmDmwKm+h2oMkiuZ0xhEMh
eGOEpIJ4gh66JCsz2OAJh6gTl+g8Eobh8OnDqDGm0Dt7NZC6OG3ApAUuHkE2DnCC
7e4lqVGHz4FIOHyTgY32Ux5o3yAfEOa7M8MElG5ob+Me3SXKDtjW3/dH6veSJJzH
+rglNjDuDftG4O9iXIgKB/PC/g/gS1A8YS2ip5lMGllmZ7DgJoSz4G+SdCc2MefN
y1bQbUt6j2bXb5sdfyxg8wBs7+sRYghfLSvVR5G/PcRwB8vppgIqsb5cYMS3RMx5
QOcqcHQigyPYLgoD/J+QfECFamHjZXHsSmYVsxw33kXJLXC/Adoozc16JKoQPm7v
GSDwRJcMRp2NsAML8t4Ilt2TwJSvWvKHQbA8DN5c4Lnp/KEAlIf8Bpr5aHc4SOEw
P98GxhPpgUNjmEStGg6/mthhJDDdN+MlLQcn3+GvVF/v/GdOd96vHMCB1mL9eMl/
DIhjQXi54KcjQGX5WZnUBOi1NokG7NyTDNWtDAjYdaqbLfB5Cp8Gf5jHCyyTh6IY
is6WIBJvoQcnMK/pkbizbAWfVqTtr7zL+EGTxHgmB8KXT3EAhbbTZWj5BmJxQkch
i6KMIOJVMQgfH/SuZzITvT1mlq4e1h7G+LoYE7/R9ZbHWtcerkhaSjgH+HUlgQm2
mOSI00VmPl72z4NNDxT0koCqqM/q/LaXIK+vSKm+wxbycx7DsvnQu/PU6vNHRTWZ
K3+P12cKSZDAPpZlxed8Tyvl5b9x8zDBzulJbWKma/a1rnAxZ0jxneSb5NJ8AXpi
IbHEZ+mG754xw2w/Rf6xs3qwYy7pG95nPZ320KNPsVqud7g1YKLlQVmE+8f2X45Z
9rMTF9QpiZ2GigVJUo5L8Qozzi/5P4KBLsq3xyCCHXA8nYCpB7gmF0HwmsveCQ9/
Fy04NcBvmpKtkzDwrRcihik+wM/xOTpLyCruGlXibnL/YD08Gua5f/V3dw1M28jJ
hAOxHnnbmf8eE8q8BJZCXFmXGC/2SK5mb1ym+HAsqNAAQ3l5SbTqRCLBmydADzmM
4ANcJOhxTCmstNgM1Syv+IzT5y53tod8WJSNACAC9bluG4mt9KEsGMBHkPReOKRJ
NFBIxYNWNM+Bq35BRmsUwm0+WmBCDfyndVqpOQnQVzakDj/+Z9ggfHiwUuYhf1Rf
t5fv1OSbfrz7m9Ty+q73fF8/pvDCTYEHCNxazQ/tFznDOAi8Qw87DUUJjcG52dG3
E91hHJxykphFQxLBf8ooevU5HBPrm0Mzz4o4LPQ9+TWPHu3zIWaATM3PFTZSoXt3
DkWAqWK/sFOARs7vy5oe4Pkep4m1/vYvpyS8OeGjMG74m5evdZkIpHivNhEXVeP0
axURI/rk/XO62C6985rxD6QqbYH50PWeqSx2FZ9KRog5cogTC4d+Q74ZPGeLGqDe
qZA0zA1zAjGat+o3cWHBejqMXybPtYogn6XQnVFyWvPu6Rq8utOirZHCVNfD2IQV
elNYCSY/aWIUm5jpqeqv9S1W93efbDWQ5KWFMv17ht9sLKf8QSBn1k2JyXp0EYLO
X+SNARKftJL163hYkTckKnJDokm0rp9w+p118BM0xWxcNJSrNdDSBoco+W1Ry/bf
lNZ1gTy4f8NRmYbmQVVfHDqRx9Kp6gC6RLBCsHT3nG13tYLtEqp9ISIiXq0qqCXd
G2BGyr7CzhTK++FQMtBQ9lMRzz6mb4mxMsL45vPtbvKPFTvBUn6CiIU6w125ZZE+
RIneD+Yu3O3E6IOu/NOriDTESspyNPqfcpS/eFHya/dXyX/6PQ1QSgU0HlNZQvaO
lyNMHwdikYgCRYlZUDWOJxkAGNmyOqKcqNUm1tWzypmAgLSMehuLQg+QwaNdKYKX
+1b4kqAqsckcvko0Qcza7yt9PO519ZUsQpU0P8mcdnL6QplBNC1If4xh+CBrR5nx
mwJAo9H9rErh4QRlV8JlW5LdDArMb51nDHrJ18q5WeoK2FbuA/ZaXZX0GusguSLC
u09R4WaVdPgAuqNQHa32isaoLFaY9KIkM1JGqAts4aPXzWlRPBzIOOJukjgpcCNz
ZkWtQOokU/Njg/hk9qfziZhDlir6tEN7TN8wGC44qfzy/ozOjV1DQAIMYry7Xzga
RKJ89qOA/oiLYiuSEZuk+bWpDN8fEX3Wc7cINLDNVE/zxjLGwCx0DOI9uoU8Vy0r
iD54wYUi8dMfo2rFvjrJ6N+LUGcU12bP/dtH+sCwFrbe926QcWzIbAMKcdt/sHKk
grmPyLS7gqmxhXouDqQsJnzDM8XB3rrCNt3JkTVvJZFvHoi/qqbFAi/Yv+YXwGJW
g40LCT7f8e4tkQmgegBJLLOz96UJZvIjcPy5Gkh3Ckxwws0wczpr6U8hbsQLskL8
zCnQiJ0Euu3fULnsoojiRLyCViQjzQHjcRj8V2fLbNP0hcZvikeXMXdc8KX0ngZ9
NMHIgxOLGJXOThT17u91S4Zzg7M+s6mPKAeVNp34+8sOJynx5NaP90VxazkPw7D7
terDsVMcKbU3rV0KlvNhVEe6bMlbrH9KTWHkQee+4i1bVcOFePu5dfIS6LLglT8R
tpMrYlAacJkWE6Li4AXHY9+tVH+6GB2mFvKQQilTYPcY3b00nmQBKI5yFJGBlvk4
3sraD8jo/zDkGExlDFDiJx11szc505W1EwNIIxkpRf01atvWjV6hvLyqJ1B1Ro32
2qangM3gDHCkNsgjI7JcWySpfrwCW34UTlAiZS2iCOufTH7Zch8NV0GO6YSRTBRB
rmnoIzQPqXGieCT+H01A2n7IUAwnX9/r6q6XXJehJM3w826QrGdTzj2KaKI/WLHf
E3YZrYDjXkMrvAXMCmyC7l+NMRlBATIFE9DBt+PiAOZzrWXrsaFealDjF6Q3aSMC
T0730tusGrVkYL5UCEny0dD/+MrGnXWh2eO3VpxTOT8KugANUS5pvPkgTU7V2hSY
IEjJqppsQqF4vb5Y32PSdm3YmWzLD2F1qjwZkWcX8wS9z8VN/jEA1Pdg1O8yzTEX
ySg7B+qQ5J6AjbSK9Vzbzitr20I/Ta8CDNRnuOteR4k2EGxUeToOQtHtFl/kzkuT
jOwDahJMHusOogLSIhnZai+ykThdv8UFNM/gW5r3AL+kJ2NbrKMThaEbal44cbcQ
9VIABRU2i30r7pbsL5W4LUgzeO6oBvMr4mJkHUcLKEVuLDFb7s8tAfesbXt+bI7R
iqIUeWaTIZ4K6X1hQ/r64fEBGufauZR3qGyD4Y+49fjByb/iXzz9OqYALU8z8H+q
VZLI2znw0cEVOh5O9y5Oc00FXxWfdxY4xcTfClmBsDRCHPpGhu1TM4i2h6RdIXHZ
zzTLEdIWqne0Ljphs07kuE5odFl/2RopDZpwvazO+alnbUkiGN3LsTGDL/kN10yJ
+eJAb+hoPNNH1wdvBsWfcLKsXuWpNAxvp20SaYzUa9YtY7baWhWl1cCD0fhIGgQe
UolYNhDEUP8eIDWq5xiQO0Ps8UHF6luHvwp9lde1l069CTdL+SCPMJjnqvKY3Sys
ZQbFx91EywC5sV8urtv1UZRQN2NkVgCM5ybi8K8hQ92bl6w6OEUJGzvUuTywWznd
rKOfEVC+GyCMD5EY0NFBy+r61u/AzL0ERLv2HErez53qmV0GPGgtMU0VNipEx5O9
fnxsm8vHZ8viS9eI0siva288WdKWDJUqha6bcgf2n6v1wSvjZZXJGLYHvZ+dbh6w
uFGQniHW1c0WWcwqHMw2XE1t7HZH3HlBdsddS6lJAr9Hqiv9Xtk0/c8zRcTmph4W
XhTZydK1VbgLjacvxirFnkOl8yTNtAJGOugvNWIWbZfKY29lHX+p6Qh1n6g0e8LA
b3KHmoE5WxjO3AVW29gWE786mJ9N8d+HsLUuClH2gkylGkk8HxgaHNPFdN0ACTEb
OBOj8UPPoA24KaLmBWpl3q7oThdwsTpfVEI9iISFn+CbqDdxBYh5/VC6nDYmfccZ
eQHgFpGQp/4pl/5wd9DdNZ6mD3KTot2Udw4di9ep/+amEUnK3T7OGIFi4xpllqLs
Zdw4TpNnAp/gF8XMEcDrsW5WjBBxRktFm3LqUNJYKpdhK13sRfu4cmXaoqdgRzOL
/pvTJyITfWJ63BcO+nnQ06nHvQ4dyt0s33096T9XzHVgFr7TqWYUL5/hi6MSBzuM
7dCMNGIN73FOOIYxfyC06dUJRZHVpQf9/IywFLWswo1aRWTDj8Lgw1EZ5VAEwtx3
2ajB6giC15jnOJbAbiuqzeyAFJvu0/lAC4Y50jAAjnidSrZAO12qKZe3i3fq3lyi
J/aRwbs1fyNWu8yosSV2vQS6fZONwwFRg0QDzw9tH23+IWIQqdvV6KvwlmIw12rr
QlNydi/zJZnwRP0RDXKlK7f5vsPXZuvT8jBLD883/cE+CbJmC7OnzH604ajiRwg9
UVE1cK7j2Yv/d5BPYneyCdPD1iJHdb8OA7is2LpvAHlefTyVYND3+DpX+VJUgj+M
I7rhX54ylto0MnDsM1tmIsrMOUaBN4ofGP1Idqj0qokr21zsmHVU+G3I1cWf01bI
g9QkiHeWUA4/AZt9g/PjQGwogO0pTxquZTEMWtjhtu8DuAKT56e53es7C3JZcwO0
WNoeYVzonI33nYk+GbmyU+wxy+OnePbdam/+a+Gr5NXNOLVYTOqT3+uRxC9ztrWq
wkPdfo3bkdgh0FchhCkDWc+ZCpRWrEJqcD8/5E8/oCikg5Vx0iHMVQiNdBSkAbgD
AchrFiV4pldMioRzuoRrba91LpQdlGQwdFFIdPVZShKD1/KuEWcRKMoKEcloZWk3
2n8tDQAWopw7M/zhWHNAdgbLvTGEkFN9wcwWyjMVmVXSFB13w02yRtE8OaVft09O
7vzNR+3y2iuVGMsYu+BAOiTSPgV+3kVIu/3LdlN+hsugGXlkE9c3qfH21yNRDhZ6
vyLKJcirqbN2Yg0GxHOSRZ8JAnmhVse4NT55kvOa1XuE7QUcnCvL+82At7UbOxLt
8BlRnhRaF5yIGTbxO8yHqvtBfB+GHECVsn5XDnbTz0Za/gKIuRQRVPo/OI4jhtI+
rjlJ0CdZxvVbtAl7fHCeBd3kcVfMCUkC9WWvvcaDzWUK4hMmOzw3BLFtdGOn14a/
BmgjqUxUvjqKMVqlBdDTb3YI6fUq3uzbVVa78DMNen9nD2sOJD6ohopUoZncPWu7
Jr7CEMPg6Ko0DewtjqWUwQLxXRYRz0x18ff8kC8Nulrm6wEgHzEESRrjygjYiyBA
EDPRn068y5+iqAT6Gm/CSVpYs6Hm4HrQR92vePMWZc5ZcKR14OXVSAQnslPqK3/9
bD7ytPjBucDPdaGl6k97fgQzYIZuH31qmXv2cWLdvn3KdmgHEvWuR67oVpS8KV2w
AbJERR4HMKmubUEFGQ/UAYhGhj6MuQpp/zBQo8A5m0R6WRf/NG/33gcP3Lts+FS2
adYCUuH4PlAPb8yCVqoARIgUpYseYmt3DWjMDeSoczUBgf6vXv0xlyJFRLp6lUIs
RU70DPYVgD9+k91cMvy+z/v75Ayyu5Vi9kQVfijnboR0oHbsuTudxDvmEi1yVJ/A
XkpX9sk/Fx7bPOjY8BgjiK1pW9yJdRHNypj5uOxrFLkNThdFWKhsg4teb5a4JGN6
EFCgii93gpocq75nfLPK7CdHmHoTt6ruZ9JjYkmstLaoDYzgGyF0N4fIBMPe/BXT
8xRajPYBIlJqKY8k/TdlppFHathO3JpY5/adjgIgWgoskrT/WeomC7l4dd86WH1J
IjOa7mtLYwwIeeB6vBP1h+wjoo+4HhMTMGhUFtXcCx9ylJa+cu7oJ/x0GjrdnArw
pr1Ijk9Cr5jo8CcYS0IAPdrDvEYdCqF2ldBFqb+m7pVJEJIqHcUyli1hHUhqSaik
Gzy6GA9SEbVTA1cMP2xZAz++5p3CUFf9dOS1HqrN7FBmfMRJAXWKd+BXHUE2ClKH
IoOdjChBxS6t0BA4XUc7YecHR2z6NLHV8cz0QKzrsmSZp13SkTYsIhGUr2u6Djsa
iyEYKsQNGZYmu6IsbHmMYqClwfRY7UHb7zatp0sncM03fhiK+KhHMtcoCtCZOZlj
xPuCjuej2obPl6IeQtpBSWPi3Y7N/qh/QdJPLFlt8bLe5uKxos6VDbM1x990oVLO
ubUKLbXsjJM9/4yzjwQufzizNSsKs16XSvQK2ZAG0Ku9OFwcDBDsSHug3B/5/U1D
mBLe1b/6P38q2twN0dbEJ01dfQw05o43rtVzvO6aNMl1J/pAlcCBV9Y7Xk5x4VAK
T6KEGyyCzb8AU8IZcwoNLFldqhCdStiO7cINkaYBzWr5SF16tHjnEmsH4RgEiK1b
4yXA8eVrr/55FL/qLd8++SP9mXHnz7LVLf67olVPr7uyuzRzKEyuwVZdjWDGfMn8
toFoawAipDB0WZ9Hu5/L+Qx6AFtn1Ulj7M5hYE7uHrP6Wjw50aWK4XShp9kKk39U
Oq+cHNpgB7KyMzTc2h80sE7VXEhvsSxtYR6l2jH2FjFnxGzvPEnooEi0UkZEWchn
OP2zTAjw5EXa9lP/zTU/3iIXg493cnWZFh8E7vpSQIp7T805MYlLf5SIX/yW6VGG
Jnp8xlcAJkJFeIp3VK6IX6SNVqD8gtoe5BZx6/JOoQq8oEsIBsAfheVA5wp4G+Nx
JvEXoHRP+ZhU61knV2BCA4QmAmc2tx4CmrBcwm4u0sm9bsJ8H5amjqx6j6dwfa7P
VJ7vpXpORLjEUFgzXDjdVw7HRSoMJLP8/oJtuacLZDIudCzcMDYiPfOyVupuH/5p
HNbTGWrZAD5QzEvS+CIx/+Tb4Fy2Xg3e62mTtr04gTzq0GXu4dpfe5mGtvDUEdtJ
hdejtqkry3RJeLwJucE1GdTM6j0w004lWw7aZxNZgj4bJDleeUvSVUwRO4h/qiMD
UNDfVwyU/8lILyttqxPHgOiNtCxXmLLDOoq4Blgw/GyeaMW1bxA/rrviSIm3vykZ
h4Quu81Qp6pLTT+kZbzP4XOGFMRh1LiIKpFUFKlo6Czsy56o+iqCVMkAfFc5H0zz
Lp3+kqkOQaUTxDW/fVMK39QvPmTEvNSVgrdZ020aSDELYV7gxC4wr+WJuL7LiCcm
VTFtYmNPc4mfwP1JCOmRZGmAQ2VzprI9834NkhNOsCLWHv3HUIiL5UkJvb+qUUu8
Xs3yrK/U+Bm62r/QdQE+ajytrbG2lopNsI4Bgh/eV5pMB7DfK8DA6J+ZAZXEabdF
Rrezc7EZI7JTcHI5w9r9mRWpCGcKBg6e6Ig6JJGa2odEPEzCweDkZSRl67nOpyQ/
AXJKzyiQqxHIBa+Sln0jkUXmyk60Hkawd4mXxxwCuZt3/Qu9nNyd7EYoFc4sJYeB
Rdpaj/juwGtZqMOMKy09v/O87nc0FkfAWDKSRE0kimMjkzyp4MJwrZIL00SF915j
NKbWrBbxQan5wmVOC1IZlZLWkTlHiHZA3TSrVaFADr2Pe1izAuHwDYvmkKbOg3iw
ZynvR3wJpkWYLWQuEBQVKQVJszzLUDcgRLvEXy8vwiaiJRIwXvRwNwRv9bfmGc06
CquDLDbPFaahatuOoh7+NUY26S1Nb/4WxXeHbKMp9FxuAi52+qvfhOc+QqESD1Qd
CzcPbE//EBRLHEYxwbAzk5Gyw+zBD9zwpySEO5tsKipzumtKnAwio2pjkfojnmbu
ZJvlT2RPGCc2k8m4xuoVYfdtTJR52mLGk50tXUE9Zr3UEvKtKj1fQCrC53Chg1LA
iPcez9M291TVTRnk1xmxWNtuR9WKKczGgZUax7iQqYj/9Ga1cwvERZCc4LbraM94
IHukyAgW0eKrS77NqGVQNeXFagilNudRpG+FA+mtMSSQ77Fivg6NXEKwXYDWC/jc
StYYvjIK51avBoV0UT3MuJZq8ZJw0Rf/wxACr/A+79dyv/EXy4JVR4kHmqokUlaJ
xgaXaika8dG6dYkOJEkxxPMuCkNxul0oDr5L/TSJwFeE+cNS3Oduqky8O4Lgym+N
UArt2ugtknd4U0A7VEetuwSnuYxSvbfJhuNQU2GMzHL7kDBZkyiVJoirwYoR6Xkl
LB9C1U8gNRK8GxGwuYRxj1OnrdDWqVu440FabImfEW/WEv7G9xUPQ8DpIydOlyZ8
N17woWOvAEwrM36BSKbp7SOADh0k/IJg7BOI9RemgZpk/p9SZOE7n9imqQILuDtX
Go86Kvt/gnMT01QqdrUpgGWD9eOgEUuQ1OBMwbKKuevIhdetR6oiuY8CCNShHy2W
xx5UrYIIQGrWMTWAwoiYoquCQJD4WYtM14MtOFRk8kVnXsJhuJKz5EahKUCo2yCl
lXLHEsevu6RWn8oLueqFgotpGRA4VGoK86n7uXVnjaqgXGDR46aRc5zHlYNgdCWI
XmrjzazSdq1pGtaM5PqJE2hhk3jONkfVhzieBiDe7xoew5P/HNv4/c3AUJYOgYFu
YYbAmic7A/si5ZBxpPZr7pYdx6qx/HVWiRYSCRmgV0gCYAgNSM7/OxbSM0+/jxv9
lllqDo6iCXR4nrcZnqXP9ndg2vq1nNGX2mV5ffQArnq/WvaismQyTpyYynKFR0Pz
UAjJJsPyQjj1T6XGBHuUgUUQbfUTBB/TUjDstfgbMQtw4klF5lDX1eIg/nHdyrnu
ie54Pukpu1PMtb6bFnOlvfytQy5RL5fYkNPGCyQT9kAqTc8NoZ+IqvdUHp93Tou6
npBqzYY4Xjvid+Z7JWjqSAD/A2/ev8VYZkPCNkxFqkELqykANwZiiFo+CzxeL0aK
vHCd7ow2u7BsWPHTfIxuDWSP358oT8BQeNceySjWzY7adDrSrohYhzCx7AJUNST0
PbLJ93rnqZhGN5N2IK7cnEWecLAhxxpBbQ0Lh8+5lZb+N1Wl5QOagxFpkMe2f+HH
rdMdrXfLS/bP6TTmNuCKJ1pCPPlDOqbFFL2JWpvlzXUF8D0OTBQHLvJUk1E2XAq4
AQAPaFXrrcGlVa6ePC8M3xrDZdtKMAD+FCKEICeY+TOiaS/YgGrNNysm95nzQFRN
qMuM6iTGtScQcCpCszbNcTBDn9ZwI+tvwYc5t0k32wfkGSbzOqBVqd6Xi6PyfAcQ
mr81X1NYK656PYEyzzm9obaWCbtrfuiNlFbwjKtt+FuG77EIxlCGD+tIk4qT9mFb
HzJv7fzZDO6+6OTqVX7db8M1q2XZTOTV03e3MVkGe8dIlsg7pDerZM8fk86oKy5L
ca0Q6+zePLusTLtwDJN5jvIKCDeyprn+RvByiMjX8oNmPXT29CJJW7+j+AeD25Fu
tcbRe/Zl6UF2ggrEJtQieVSXJc2TZlM/w6xQtw63CW01/AbnykE5NH8Fqye57X5f
Jffw4C80kVfFtfbUhchSxcBCw/2eVi8I2k/7iqPhAbcDeeOdJ6riPDDjqtJkkpCB
niGpqdWLlNTjyB3jsRKE5HOnFv3QV9yI2Q6Kb2lRRS/hYJgURQe+n9+zh82GFCt0
8d7hN2PIjhtAMGkE+9EvXFcpY0mmJ0+5sQDWonCueYlDkxnRtikWMyUHvTNxI2PP
ly8sd5vxEvObm0A57EdXRs8k9bRYGQPBWQlcGf4bE5Z5CYO1VrfLaXRSc55BRi+2
1Ldg6/FXf8Mk/a5Mi/fZb6shNaVWeAfkZ6fk1oYAaezk0hLWjXxJAb0GYwVrsAEJ
cGbB4KRG73sEuZcERyBVRa3JKluGpvv27QE54XJE4FBOneNoVzI+/ONzf9+P8vTj
ITOiMLzQBrg56WIpx+zU/rJbNkRrTA35zD40QJMfQb4VvIXZIPYeyRw1YKZiXIbV
TKQYtq5GAGj6l+XLn1XRjA9RKyaIrh/N5QtuPaEN79sVQmTfd5IeDpWqT+d04ZGJ
71IHMyARIBx9XL6lAS8alQN6iKZSjAUBgOPwfkHUz2LhOwUreeHxGiUieEIA8vM7
DKhSmaj/JcjoV54Gth6YS+WuC10tlVwiv+A9cE+Cbqtp5NS2SYgLnjuVAYjz7fVb
Euu3gJZR+/ac/SR9R/NK0kSsxMw+GgTEaUJ2HQOEu5j8VQGqZc8KJ2YPec3sqYFT
qdJgwhv5h4tkFjuYPez+3K/GR+P2uNdZiOcTFwMx6UTIelUgokgTw5x8XAkJkNMa
7ROiP475Zj7c0hyEbv+k7vkpg4o2wpAe/3Quirwpc/Duj4KklnjyJQhztuKOshv5
OEs4My12CY1ECzKVL0qrU3wGijxUNsZT08TqHAAEtEp00agffsBQwPptDW//e5xC
M6ze8oUesyO0N5UL3BlZ5Zzzgsx8+XKPsykgS7LdEeLkPgYNrTGihQ3dQhps67b1
P7bor8vRXJ7UsnMYqxsJXezgMhFcy5wLEQgAzjitD0UfYaeImAI062AjaoW9DtVr
2F43jifTkexacm/3ldAeJPyU92L1olRbvQHBrbPY/BWFaqepahXwycwmw6AGWFvX
14EVQag1NavSCpLKOK4SxWYEG/zxx1GwkYtuxD1haqiuLFs8EUXEOHMhTd6DLJUK
+thMpx9zVFPXM+3FNZ2Uov8HErDoy7rLEKj5KHFEomhZu5jKlT07jNFRWArPa2/K
NMKzyyE8f2kMrUVsng+VwlUwaEESgDhMJgAYFCn7TKOrJmaeK0puMhPeCTUR2AA2
U0xicZAkcQclyWJqltKQ09Rn63KI2HaCvh+N+PJr4LtMBvJTOZXvjZ+jK+uXDR0o
QsypDVVOL7Xss682GqDxdC1KLPXQDLYB/vXjUSo31c3VRTuP66qBAHvNkLimspKs
+FqrVJhenW5NRhiVhCzVuumsD83xar/b69je3u6onj6yRLT0q7xRlFCPNGfnOr0N
2P6rivY0/hNxki1i470pfglw15ddPoKE9/110V1jz0xFFsjryMs6u2Fs6c2//m3W
1uSkovSVuvvtbJE6LLib1nEL0EEBaaS1JAI6tq+dnEOttAubvi7NvblY9VESOKBf
hQfO93p27k2LP46kyegZnzHGkIp8lYDCD8eeiBT46pt/T5ZKcjQEYmVgOTPRJWph
5X4vCdBD0AFO0aNS7j6V5a9462WQo8akR1EuVRQrjwUvJdlnDIYAuT19TF5HZZgV
frtBF6j3mSUEdVDNejZUqrzgrDz/wUZeiccAqLmviUU2U3VilIzrytJ3DQkDf+lX
xbD1TuRxyNtwCpUZsxYh8KfDDxO7RXV4vN2Ks0yzQmXTMz3C3EqqBgZwk9L9BlwI
HhkpCK9tsKYonqWZFoFuAFcius1LlfdhodbiXTLBXH4D6/hF/N2hzZSsDtUBZh4J
Ei4BFjpeTYAjxA0EM84ocApgo70bJCmnHErO3n0tGS1q/kJSecYArS1c8LCCkYCU
3umF7V0Pxc1Ui/DQoiWR02QJRr6HiMaTRcn4qX5yEv/ECDSyG6txauSF0jnZSxDJ
1rPN0Q4Tl3MVyRWKas1WaZ/eU3+W+aGtDb5Mfcty1ACsyqP8EPvumkd5jD2BRZLy
c4TnOka1dzo71SmV7yJwuaHygpbxpYcol4yyVvfI7Bh2uFE3f7ooKw/V8p3ZNzWB
y5ebuN2GBOn+lRDFZjNq/MmYldniXFJaMpvmBiEBmiXI0yJHOar711/yUBn3Qpax
hDHazzKspR6t5u7mkfLad9nTw7TbUAt/GkTD5pePNlMxQn8u+8XNzX0ysmMlUKeQ
5pQVAQ3KHeswvhz1S3oLPq1sPix4bp7nGEE83vXG/8Oh3PWM2TRKInTgFpa+gHq+
j06jVtOfSZwmb4w+JDc2EmdQSnDvsX3xjqQnjPDA5OZzT82KeecfbSLITC8rB7jI
DI+tV6pPOZ0EiO9ys7s31wN4FW9k/hvT/Ug/ryTzxNeiCB6CruzdTqXFZ2+VNtMq
10iJ2Zse3Ix2cVgnaa52e3ZRKNR0iq6ndYEFRi39g5KmLdVsJHUYbd/yJfahecIF
SWMeWlNPgm6qO1uxR4TUJHwc+WiX46oHysDC6D3Wt3wgYOLPa22nEt1PpQZXio23
9GMH7A4+n/oeciljR1Cy8v1dWMz0Py7JYt9pSMpIJmiRZRQvDTAYlNb0Z7QqNi+r
4qwvhyansOo7l54F3jyR9sIUnLIlebOKlWEk2ZtlNHGt+/xStA5S1+7dDUD46clK
Uk50fLTckcrEc9kpUkEwHyssp/U326NDUewd6o2DYUShDPAtmRVXzoGU1DToX25c
0RT475BO1QLpJL9XXWMGvW0tcIPtpFztpS2LjJ1IsbFD5S6p8uzCGKbPlsGwdNB+
d/c43GF2usTBvmtIBnPxsyah67EGZqoLi/kXb53KFmD+Ybyspx4GCn6lZyfVCnP0
pNPxY8Vi/7ha0f1oRMH9UNBdF0EICG6LSSW56lUH9K8Qv5YzMIMmSxGQ3hdT6DaE
DSWcSi90RVf7iQW+eV8yEcobTHym7U5BPyVWnHDrAUBrBIJctkFJYsHTox6YbNfk
5VL8H6kSTGLSN5t9UxfWBuvRCtVb4bBm8rW2Sj+1D1kFvso7z3iyveIod78lrMm/
Nd01koGoHvuYzzYRrTD1HFCNWyZkt0/NOYv9ergQ4F3xL+ixSVc7d45MfRsysydN
eWBgTofVXV4pmsi7uEbESJBNiTASCzpOoZ8FCE580ZlWELixxIZJop8LyoWl0xqU
pS29UfNQTB3vnwd0GcltYWfPzMy4ZEdR50g+jQhEU86KlsOMq9NXiASpcb5lI4Sf
qBy30quYqUeiXOCepNf9UOQqITEmEsSiSvpzBOm/7mvDpgtf0tKdj07pgP8Azacw
zjOFSH7MHT2zu7lJ9ql1NKSVDb9aZrMLAWV/2rLTdZ0v6DXYuW05DN3yzXNdjOFH
szDIHlhnaoQRCLicNmWEJfl2lWm/IKW/RdP1tqttis1RKb1SpY+a5MbBO4dR9s+c
wHhCYrSWFv21/SHRGhI28osm5FmR7libw5YX/Y6iosjOHHOSrizdEY8SihLKoQDJ
Kz5ptvra2sNzx+tovjfkiLnV2h740/ylr14OX6Jz+qH9u9tQgNznNeZPogx1GMhJ
QrSH0efLgtlEij6L7sdHw1IaJ30uOGzoGY2MV/ac+sQXsbXQbd/1x/scC+1D6E/b
ovGyS48c0c8rJHHZlJaHJ+kkgS4oOCVGQBSLhgxfWWIRLEDNoOVAStjQwnlQseg4
yfFkmnY0XWhlb0htkzYvWUmAXK4pW6gnq9dQOvDK0pXeINLUXagc9taQ+rtoVlzy
HTTxjx/pdvr5/em5uOFQlpTqDNecDgfNYNr0cJzcBDlrRj+oV9INC2p1jx3xCdfO
6/cwmsqs44eXGkIzkwxmK7bIw3Ije0nQyRdYM5ElP8AhmaK9QfQm6wFeDXX3QoAn
FvJF9VBUCBZ6JQpOS7VgZZhIcjeNGzgKRdd9FYJoZ2KAfcyr+249PNDjNLsyIijy
ZFxxT2ZNpypESsk3p1JyNFrs+k2QkIX2fKX6yYPapTi4BP0782KEhBuWCqS6KiIX
CJxpJO1rl684pOX+UzG/94KnmPdqT30s6FeMTTW3T6qCEzazxzZJUMMt0rHg3nDH
bLZiui5/irnPR4xfAaFGia0La4n63v0zUCLGcJmnB1YgiJl7blxzfrLVkaTIiJwT
XKXvsjaOvA5ih2PtVeC8YrJg6hjXQ7Ed/6fH5t5ktNvBveogi923AkO4FxoNuJnM
MKTMVcBxkgxXlodSUXFqowYkKmHbajGcVhf8poO4m0R6pAl6TN74CDGjhxJF4Po0
ohL1w389freLzwvQxoJQBxR0ttx/0mIdLcg9yQwaYATF1nTBUYG+0/kXvE3uxCDP
0wFcMs3yeV4nHG1mEOVesSYA8hqwKRopnq6gLIMjfow8/IIppskXFESUpz4RqF8t
ywdHZLQ6Mjj/5RzYPRgNKhMohrgz9dTWiHXmtTCLJMGz6PZGG3gAaEuFzISsRcS3
V2Ah3OgDylCjiSzo/hFHYobggCi3DR3aMmhlhVF8kpr/GsBbGzy4rWQ3TQrjPVEe
yfrGGvGFKcg3+mx1rAK7wA8/nLlyt5OkEB5JD2SeDR6VQj8u9AIF0WrF3FKQv6Id
b/Uz+NJMotZgXhd3eAiLF4kRnt9XEuEFLrfZFFaxVir9d7UfUnY2aOcTRVP072Qw
yHOH1hXjUuICVaRIHWCeUx+M7rw2GrqDw5a9LX2X6xpK71PDCXb9oc1DgHmWOYu+
mI2VuCMNEeGuYi5mU/bZAMhSPpLy8BHx5Blx8fR5C+5wnuTr2vmPsRC2EQshDDKe
j3kZu//jW01+j2jUSM58EzDhyoaSVDv0Dc1ea++u85yEkiDjU5i4u2eFAEzpDUbz
obcXW5m8o8SLdn1NsQpagZQGImuKdhvbm8cFJ5qSEwRe65xqT1w1Jgb2MYXTY8a1
g6cuDx9wkFIgAAYwrYC5uQK14uBdlwYZ0Zdzt96lsPTR0+8slJjYCyHeMXj99TTY
srbPTLoTzk9BHCR1/APKJMstQ8r5NDJWJN2fvnkmRxzbhLYBcNyrG3N+gCa4jquF
LiTvBL/MztisfpEgH4SQXjoY9xraeeu4qpjsdkwlBSETBpOpF5uSxCtaej8Al7dZ
5WOzIa839yPTybQ9szvA1MboOjZMvbLGFUiYfY1EC88MIL7Eziw1vZPEOmMguN1u
CyRrvc/e9xHd2Tm4bw91oryPB51xk4VyP7ymt9e3lusoj/mHAHAblHRrbk0k8fuq
5DBgXeDM8vpiNvjVamzGzFQhtB9mYI5txIF5YFQdZf8DihzZUL4wQ36iTnUtmlRW
WB3DRX6URoLE45DTK6xsXLwcCoAHEXss8OcxND8O+NKPlACQD5Mqf0fGNUmcwl2v
TwKECXh4/FQ2IYmXiMLHZHyEU2l0VqO84mvgREFg24crysLoMOk1Xy4NF3xPe2ca
4fX3fd9v199NMWAoHKRdm2iyOKlrZPRwJfKEXGFvnRvuQWMViuUR//5eFGHBQ/SD
Z9bY/MU9MibtI3Z2HDCRp/Wll9NZi4itMqpznRNDzfVfyfz0k3CZKLej5mfDt/Fg
LOEJQr5rse7UAqMikzmM/wUjrkZVPqRS2MoEDiQowYSAeG7WJ5eZHnB0FtxceWjG
rxm3YJttrceNriR4rFo/iU4tcJe0kS79iEgbLBXEYOiJbtEhP2IGwej1L5mslTbO
RP5UOYcIJrHtWJFuyFMA5iRXz1rQiWm3t35jzIh+16/Cb0HjpOUcyXdMNF4Rsthv
0zy4WlXwgP+MF/NT3PiHE9t1cp+ibsJGDkC5fO9E3UYe7cIhKLl+0dF0Uugh6w7j
uQmJ783msmKo9yVCCwtCOdOWVgy640jj3dmN5zZ3OhgNE4H7mF6M3gjuijrgoXUt
O/OPONXzKo/ElSwuIMNJBXZz28HwkapVqTarlLW0XF0D+N4lhS2pvkJVc98afrmc
pTxkiDbO7t/RQj54MFfmYqcDCww9lqy9Fa+19+pzAVIRJIMC4jJefFICs8n4fgNZ
d173zUINAg18FmDJIeknkaXvdoPU93mS4nLVa4O7Qt8EGb06jDXD1A9nhW3v//7Z
0aWae9oezN5W4C7frCYUnBwG20RobwOWZAWMigP4W6pUYsk9OnneMihKBRQruEUU
5/5dnuWfUQOMxQQ6VZfq0yg3CyaC9HAyjJvDp/wpVYOAxWNeZi/tmn1PWxQkfJmJ
i9cCJeo6v6etjcEVbTo2OiH+0DQPzSPdiGnKCookJDtp2NbRfg2v6XZi1ph+p2hl
tpr2DYKfz7n0ZSMs86KR5yWv7OFA/fwf4WtwpiiyIll4uBbLMchpY3FVbA+Ctx1p
nrodhoZnvRkmjc90JLWwpi90QrDk/QwYRXaTDUC2cYIOYXk/TeV7cDaJvzJRbQfu
s4w9SQ1KbrGG9B3ZvUgAJd6/5fDDVE9x7uiEQAxHKhkQZu1fPyhA+bgF+tF4Ftow
4GRAmGYDYQjm9+10NpZ9eIVRRKQt1qqv//24t3cmmcjZyNk4WWHLqhSpFk7H/5P/
igySXBduqxSlvSwEg4Tku0wqilweUM4B0a4C8FnveJCfamnEEVJPci8IGvYu15KH
kG3bI7VdExtQIfm//vhoFDNA8bv5adudBVdtH/3E+A3Mjnpoy1RO+C9f2CfeC6Mg
CGPmc4ENtGhMHU79orlf/bOrsGc1QYeKWk32Kf8y3wRvfbllNMHtonHfnndv57bU
lW8Qd+vaQjw13u2ZGdqvG+bdwNAUAxOupH3my9O3zB3X/6fNmlEeU9A2tI67I1s+
GBhWGSJuYgo1psHJjWyja7Yx+vAoG3lRWa1zip7JSIYjUfChEnH9R11P5vJT18om
bTSNpaSzcFo/ZWh5JH5Dz/mMaymU38NHB/hAzQJw5xyEK9fiYbyzkXVoi4Prb0yO
CiSWxEATU2TxvfLXCFL7KhitTWBA9jiQXWN7aKW57ByO60HcSXA92vW4I0m9I2Fs
W1Oq7b3S92qMO0nVIHSd6dTvP9fDlWsqITF4PhhmTNA5Y3Mq+hLxaYk5KUIAYDzQ
tdJ/wUi13WyS8z35KqZHofSERmtjL9Yamwo5zzmsPjfVoX+2Il1tPOGgeFnk1Dz8
p2RP3Vkjf7lOBE5vL3gL9MmTA4RnjAtO46o1t0UD7JRyPdIaI/CeaTH0lRdQJWaZ
XSRIko3mDiVQBZNlcrsfHnj/1YFPcL4v166st4it6OmpFM1lnKvZuwBM5MR8I6Hl
LO8YesgH/y0C4qLJcvGkM//vQ+Pb1vt7m5Z6ytREZo86l84ay4sNYCEEHU/h8Usm
BELsUdfkSYaltILYxYrCOR91o2zBQZgmPpwPbho87NAJaJO24HOzOFb/myIf4EB4
JS5/E2RYB6gwk6Xeu6dDv4+HZcR0KL47pUB1t+dkN//ddxQR1g1DGLoepWqQz4+n
tYQCD0S651gfrrsVCbRG2p9AXORQCVQIHM86z2f1kbSIMVvOQeN9SaaHEB8zbohj
wnAEXeSyrbH1UlRumXK0X3uxSY0G+yCAmkNnNkdl0wVca0c12N6iI4o4raLv9/Ai
wRlqAoqv5t1dIU+89IwW4eM6tr4g+l7rzDiCqeJXbB8XV2BBQ32rCo83cKD8XRTu
iUxc/g9snX0hLhQlBm0IKui+t9xvO3QrbbYPricNH/tJO0E6bQGM0AZheEnqHC4q
fHO15OPrAz7PC5eLlSU+eAxRzt3tHjzozstERv8wsciARSvZM8TMhkz5+3ljKF0Z
DGU86lxQDhtT+rFgMj+MbCPhFdilu9Uc5/80V2JhEygikWVVN5+C8aeaPf8rYRfC
sVQZfQhIDPzeGiYibVP0xsgPTMtoCP6n5BUOL9MJ5MrhI4GNYmq20HH4QtFljd/U
H7TD6DOf7X6CzvyoqtMlLgl9d7Xni9xjJ2BvqDb9vtOw5PE7dnKH/rB6jlK4q0f6
IVSkZ3SIEpURK6FxdfuixU3iprn968N+9egJISF8xA8RjhFeo6cuxg7BZRCuK/3Z
kSxa5K/Q3mdF5oziDrgVcKdvyTHanlNInYz0YnW1Bk3p6Md4yf7/uU1qS4S7vRVA
ikEBADghTJkN7R0dgTh7vBq5BL8ojSYvXFQHmfWwwzL4KagiGLR3rjm9gQpcFGPL
9FragqRA2+R6qntZOhwxzWPNIRpIh/28UPj77GBMmR2KC9uomFstU9CJia8tpl5x
NCUy31UvkGG4ILwO6Meg2Ws7ohrzobzuFMuI89Oe1BqOjlxpPr+DKOyltOnSIt1j
vwlPPSuZIB55GNKEZhK3CtqYZ/yVHtDhV/0g2r38aJ8iyxPmzUceNNBaT+n26nxN
Zvm3CKCHhqw0twRmoP7/mL+G7E5QHZpvrnIW+OKzUxMPYgzxkywmqhguy8w3wCnp
5THj/p3cQl6J7QFqiIYZkLqvLimczG+VZRWbUoPQ2j2eSur2Adt7JmBzmgmpHZB+
E1HI67I76raQdjAy3TUgs43tBrZIyBJcXKvzSJKzoy5QKFYgz2eFSV0rBqVuylss
C3jNAvAB1TLWnv5qWZ6UlRKj5c8Ugq4QA//cAQKCuHPqj5yniZXXq76LoSyMejT/
EqujdMZ9ftPWIE4xAs8W58COKHn4Rx/Oo5l8T9zrf80qRN39o1jEA5tFOzj34F7G
oNScHF/czOYLvUa7nWz/VjWQ4JKl9ld0UQjUVPnATgyupcVBttFvDKW9pP3dHSES
PgT8pdGps2LQsDtEI9BDejFhhPduzz7En9VBZP/HoVM/Qxzn2sebGABVfE+9ZQeV
bxMWEZY84oKVc21A5n6cmmoK1RVySeCOLZPWNN9sizyHIGdUTmd+Sz/MjR7VOKeq
v0ZujTu+CqOnShEjU121umU1N9x1itYVVYP+4vVUdpvzyxvVFe3RidzB/QAQMG+L
P1r3vrhTCPH6xiz8h7XpgKRzpLFkf5sYO8rhrtBf3NVXOpdf3q/vBo7YcwrIbVbp
UlxrwpXTHUh52lh7Z9tFIH79g2r3WOKhH/hxsZwtGrNGMwv2Hkx4xJZPFc4hCOEg
QbzSgb5IpR203ZgtquqDshmaVUOPdVf9hWM8lRnSt+/hut/Xr5L0N2J5SBrjGXXw
hmyf+LqJ1w1J3akMc0ZQZrD1DSpenPJQatLwFkwMS+PrMNkT7f4P6DtcbmH1Afb3
CLblfmlepwZ7Nh2KfIBYTYgFE11h0BLYsJNelTYpyra4dbsexxRTVNpZ6jSC0Osj
IRruw4pL0/iEcTxqBiflSVzLKPDjey4LquP0WotldHFd29uu4UFuGveVsJ8qh4By
eT12jQYRuGPWwM1GVNIzI3WVjcZh0J6gXri5LPwddmMny+yXmOhj/Nr6RLcoqcyR
2UhgAotEkmIZviUZR5aQiJeXUzxSnCQDqR5JQ8KtU3ibTOM5ic0H9fdZQht08ZzG
/RbQqBLsxwfLfE7+celZLFksH8SgHzqZkjOGIP+u0iN6vUHWuxeBWJSnjtTRC7o2
2cEY8lyUcEAErAYNX9kd8tHUocC/sxIneclPJXINEfqMWxBmXMcavEK2VfFidPaW
WGiIFE8JTt6w1niMwYX4LQHH2A9utQwxCykmtPf/FyDxWGCFjcj8SjGk6jKsXpZz
aaaOJVWrZhGrjQXdtUhY3U/qIQnlHrvUFfKbskywgm7wvaeF/Lq5nTZJZYvPuWpG
rttXxdndpaqlI7+uS5ErZ85xGscGNm/Ks4mUzwb+fgoUwfpnphHnU0vXyZiLRDj+
+B+nXG/tJbu4dRUek6zRAv9Bjk00fgRosE6ryHIExsS3dEUnhkvpSywUh+nb7vb5
ZY3jy9CM6FBZViHIFrfFmCg+w8jEfbVayqbcLHK/oLLa5NX1v6bJsqIrqW3RlOi6
emaUrKrz6rWnTfRQYPfUqwbtwzbOi/lgN3h7GEX8oXtismE0VJdZRxZHw627YYN9
uRFHWCUpthYJ1G79joz2RJ37c4qW/SfKY1YddvmmevWyfPTkEQv8n/MOFRqYghJs
kJ+kPbRx5FE5d6bBQBkmsB6ArqFvIyvB4GHKXDnDm3uspVmhawbFVVC4t0mzi+xs
3G/2aAesdEedIRq0dUesHN1v24jV7GijfcXDHvM+rnJ1smmkye0Kwv8N1S4HQvob
xg6E94IoAk4MmBnSEjs7ySGAZARMFP04qZVHjrkiPbhP1lIdc6TFfh7j9b0Ak7rB
13sNf0hhcDUna430wZmqGXuR1oCCn3lqABmLxeBWglpoCqd9Qmti3Oxi8iEpQkHk
HstfdLPhLiystQ2ZYKDtr6/nfPIU3wU5S5r+rVZiyytDqAa14IIpvgys0ZmWibZW
2rWpRfJ2LNMCi8vrsP0uaJG9rswWyI0o82Rtu60wWpr9lKByXvECl6oFiZtyxAWb
5DWO0d8oYJ5Dhh4F+KsAuI6lwKqjmklJahXNelLwzS+UsAlcDI5PX8sdrZBAgf11
9IV1TZx7XDenaWuxfktVKJY9hhjy+FUjW0T7qWlQMeC/hYX+nBWcYHTt555VxOSz
uvUV63huT9/df8sW4Lk7zAcA7f0HNPdxmtd6o2jjlcjO5iqqF6eskIs5QGTo/Pb3
1sjR7Xp7WxE9o+JXGs3VIEm1FtfUjTc1MSowuTetUuKevveh/PKfxqDwyTvcsAnc
2kN4lolWC1iDiUtn4Oh1nFhUGW+HrzEt9f7YU76W+vGatzJcSDrcxTHTyrcNcK/p
VxMiHPbx8ezQG+3TJBO0BJT7sbcyuaTvuqZdEqxfpCuwsWOfMubDe/w4/+T5z1Yx
KEgUy1qvciYhxyZgcbHXOsmjPWQpwdsjaEiTkhtbnZ/fJm/o07bivUCghzT6rKL+
hAAmvNlIuqKEatI9o7Wxy3SYwXGKKosuVRps1i1FwRW9Zj7vXqueggm3c9z6US15
cZOSWRbEHy/QpzQBSHlqLQ1mUrD7b9XQSI1/Rk6vKLB1z1n0/96pqfTasoG8yKJD
Qm8+UnDvL1D0hTRbImP/v5y1DnSY41kneLluyC3n2jWmNFSdTnXOZGeyK7UkNd8Y
wY8DO8bEeHvQMFBY/RDUyUEgQckBXcLHTiMpD0CTQVphfKhgsKnXAtDGfsslRFWY
f4nXduKSvjcZcINictqIZ1oaW+9/pWoMJz5sPqGA4CumCCOZfFAOS7rUJrVImoES
zYtg+DRVZzPU1e82blesl1FvZAadl6hMNadFAkHJZY+h4vbibOM+ojD3pnECfrE9
Yr4EoFF2YZETaA1WR3nTBlh+NAqfdIP68jW5T4Ij2a10LrjUpreZINvhnKJGyrPW
ZUMhz39BT51pKCuf+5TZt5bp1WluAkLQPaOsO2qhLZsG1IL145hnzZJT2ReqIi81
WrgWi8cCKa8pNLBLEGOXBnUCKTdm7nnH9GU10xQIiLkOTKzlLMryRw3Q/9EaDSrq
xTZUwpTdm9Vhsou86xeR/4PvWzaEY2mDx6iSaajZ1CYbn8+DIRptt9CmU7Av52nl
fZpRiL5DLatgphWsvJEdplf4XeTX8vUHqQVNn1HZuLGA7MnEQCMafAhzFGCEeTAI
dc2mHikP8La9gdK3iJtjuGiP3OtzChcekaqO2tdTXjp6gbKp9D0jFLsFrP+Susxr
1fVi/w1xEKtKVxSqzvfhAgcFGQTVpwoYU7qDavdXCiFNSAJ0O8PlkJQWg4pA7myk
SzZl8X3qrmtxInPiw+tgEvwiRP7k33uyH4wK4v87ELCyh5IM6+LyXTqJ95TJzMNj
qnmDP4cBHbaIgPpF2yH6kVv8OT2nrRwVyKaMyS/tSpdVFvNKvtxWToT8iyPeoItI
lHJnHp6Uf/JZrvedODxM9S1Ob04WWD+k1947UUmWTydqMqh+f6ynUOGd+lNyAgcr
AE+Dx7c5hVPG+u6dj1TSeINEx43B2Hahq61BtpjVmAhrkirp+dMSuG6uWb9uQVLy
RIQGk/zirTD2JuTCvVtkEcb3gu6H9k7F4zQ9wBNa8Gk5ffB8OjkAUrVhEmEGaTqC
NgckJ0cfFZrV6p3D3B3mSpjzBXk5l95k53LlC82PsGs3BEHLSnSJX7BdTFrJUZJ0
NMSI/Kds7VsN4xXfbt/OIPHnzpCfJZ5PlapEJtb6decVWCCwWhkNLWtg+DEz3lC1
TuQmETuaMFH62+oMqfNw0CQFA61UkWtNpoXjK4ej6Sfrm6RxgkG4DG6jmx6JiK1R
aLsCOODYM1pUqcAANKe9Y/NbeFRoDT2DNG+VQYkm2Oay77tYTcYSOCtME7IoCgQF
4wO6j0Tzh1NNF8swPNjSkt3lULbdGMu2f3EDLuIeKoEo3O5Xoan6XwBlV8Wf3X2Z
2m0P4Tk44KphpunCND675Dj31GicFy0OlAvLtMWAOf6QBy6CC8UVbQBZe/+pam13
l8+1xs7YEvIzDjq+t0Bf4amPXz7zB1ytKPO6T8UEefIbbS29t4L/LvSTG42QsOWC
rEUbbhwn1lK9bJcTyPVYXDcphQB2LNTFK3O+v5/zEKaW6WEca6xSzXvAZ6rQW8ux
+iCPIFeclZxYxwyPJLFXWOqzPgm0RToIgESaUmyqhgUkzM1QG78DbkIdSBA8jO0W
N1gBTDI32h40VcWXUHjcNRcYq1OTLs/ZE1yFCkGcA4NFBZizlqOrWDf7xgej54TR
r51fWA08J2Fi9HUYi1sxTublreKE5xzGUI611f7ra6ONG4g4XTVlIOcwWF3dTxQt
pn6UeEka/Di3svNoM7H/ppRMG7wqOC/vnv1gsq4Y+nRtV8xppqSV6W8D5AtrDogL
Kfs1bSVMmtc+glLICYQFPOVssMKSM8tBx11STqwQBc2Fi2CPTFcUw24Ds3e76+Xf
LFjAVf4NA7Rwerg6dI/x/EIF6XnxjLKG9CUSduJrAeexCT9awpgtiwJyc7VwTVta
xLheSzqKOaiGiGsFVynco2XlS/XVTFcOqpYNyoXGuakkVTJb/Ycr3ayZL4IN32oM
W9lSey04XuwGz/bdnltw2buvYL6AbVVt496K862hUP3yhOT8yJgem8QwS6Jgn+bx
iyv//GPs2PpaC1+u4xp/KA8VlAJj8Y24huBTwfL9BOy2j98dTEIEQ0AdDeEWMyrX
P4Zg/h3qqEv2KEaGlWMRppK+Yn2SA7sin0M1IqkDojEPSqSDnx4n/0389No4y70C
PSnmr7RUFZcVwJI//j05XEocDvM5LwihCV2Pfe1WnoC/OK1t/lLksiFPB8AkG+bk
6dUXkbMnDL8bnHzhK0KvnYfimNl/jtT13xzKpc44LxwWmQ0KaThQR1QhoQCGdZtf
+PcNgJp8Pu3Nk8cvbH+0fBg2nu6ykKvaozONsDXuvuRSoaVWQ2IoHQoWahOSwdEZ
HosZ/CRlCqweFfmraUWc3rZQFG7ftw7EEpRDES6DeQ/qizq28Sr19hE82NPS2owO
fi+/mRBiOk6+CvMPSVq1k4lMsGHaw89vofYvt2FQKr4iJs3pyNvmHVS/nRNx2Fir
DIxhTFx5axThzuNJByvRKjJ50ANtqu5pNsBQsABafjX/Tjj54qrdD7mYrhqduotZ
H51CuJXnUomAzTQlPTo5nURyeQr3xbQebvNm7BTpf++luishO4mfFoN4CQf7nP0x
trWqjxZuTRScvqahT3RtDU33xSLMQqjqC6MnxrL57X9sas6DoGPLKiFoXf7O2Yno
gUmsvRwz8A8LMRCey7P0mImX0fQ4fkT3mvo4LyPeGjjaNXi1JmEeK5cLfXVCi1QD
Ky1NOho1zoanvRBpUhL1fV3IKU0hFEzPODLtGztf7KEXE4bS8FKQcueQxAoBHgl1
wn9X8QangAtv/pcwJa3wTfE3ROwfE+MVulSMyFhs5ra8KAa9klfnLi/9pFYDizrF
uaqO1+Ggv20ZLxCOu4EyfUAJiZD5YSHi0Ji2VoA+zeHLVUvjL5bipxEloMNOV4k4
mpwpQn/uk1QgVpIZfMkWcSF0qezzUaZM5SAMOlWTAh+bZUKkNK4jPyUoRbt1sy6C
2txxuieE50lAz5cIQCeEfwreCzDbWR2CjOfkCMI+Q4zncU3xsnXmGq+QLL7tXgIe
R9Q1bB2ZwfFfKLEFDlQd20EWhwOYWL2KkS3ZXSTbVCbjLSYHoMgFZ8NgTgeAjG7X
KBKLMy+eHDW525SFwhzQchWr27in1dIhPBm8sdqKdglkEjPh0HSHuSA8+i1ff/Cb
NrtI7pHgiY9yLGBRvWKgZTvUlgzGy4+A749KEr9FtwqZVwKc/oSTKwJqi7qfZpj5
OPeuggmjIDvcEiwxR9PeZ1PMH02WoafEIPAnfabRFqHPoz7ZOJzRlnpzJHRbE7o1
iYwvLKFFrZm384J8v51pKwKHIzmBLRNj19CfGUY+Y0l5IW1Y80m5bq/Yxcg3g57k
oTphTL71gUPFSUT5uo+b/kjf5rX04783BQIT728S6wPceAjAYbbzkQrYFgzj6TC/
CKWiTdccd/23BMOOxwKMvJqej69/eAWv4R3fQC60/hmC3ZyTVlDQR7DiOm3leXfL
1cmtFqa7lOQQtchouU6x3ZCCuYo/lmi3GTMxVaYfg5CoujE0X+2LuMkGuX0vwGXu
Rglu10iI6Ss0A2+o4rer4IOmh/+pKkhy/nhKDxg92/mymVkEXSfCYI+Erwultmb5
r+QsOEyffyDbAICVaLtovyfZbuXK5+DSFUgh0Ns4PYh9e3VzHBDTTM8LCgT12imB
kwKxzGj4A6Xv1MVmQVEkCZt+rIurjB6Q8yr9H99MVzGj61cOYPxeCRe73hOzmyKi
XGmj2VCL0j0QOsZQVbSQ44lY6a5XZKFKs3v1iQiF6FvYHJgDifFtxtKLo60uBPXq
gLqsMcM2fLwYyzFXXrp8dalsV+1nwN0V17yR/iRmKG0IG3G3YSZTS2TcCfCGi+8s
GsEFqPSXFe0LTeYZqkz81nDgGJl0aW6Zs2UDtjEUQ1/Y79meNf9CGOly9sRoyo9H
FH0+KsfeLeWyHFGDpSUfiFFf8jqunxXAltv0NFPEpn2GeywmC4kJQO1lKw+M0hOg
iLGQKlhUjmTeFKTAKPCf+lXIHBpbgV4UFMFWyiURkdL+55uzEWVFzNE0EWhxhPPR
/ALhJuXNOZ/OMotVC7t4oxpuueH8ikUFMB9Y51a9kXeEQbam/02ncpcJNP4GXmqS
11krV43IdYcz1ZvIz0HmCe/XQ7Ko7vnAsVPwYtBJ6X/edUBAfroWmXKycTbSobVt
NbLdu1BlY8aUeV68ajCRb5Kw7PyJy5+tEDcaDezXo+nX7/MeG4xk0YFP/P7GowYF
QEFx2DLpAaDG2+HG8FL9sD60zU3Q5hRidJv6lk1NOdpdJUFltvqeufZYyXf+u2ZT
XMZiZcw0YodS7WgBz05UOUj6yjqXUBNgBqeowcl2qunyre+yR9XXP18BXC6pc9tI
iZHhzDnOVioFI7UFR4M9uMF1HJzt/bBPeXV2ziWRP4rO6kNHaG5wyii7fQYj9xLD
KJ/5Oq9wt6DpgjPU9RwDaMGp08gYPpfvwTHrK3uBvCHLRE/cKB4RJXSMLDhjIClX
arGlDcdXcfR3UYiWyXY4NtFt/Wm0Abo+HkBIvoyvtYont/E4bBx/85RgDpKNx3I3
eJGorwhVP5pevsqjP3/OzaTHD9pM+nqtHbDpClOZ4pzhxVwSsIIgMhRc5Zxs7uMu
NsXEc1KSdiBjJOCBZSLYJTlJxX0xDlOwpnRgeJWVrTStYe2c1LXuVPcgg0H3tMIY
sKBG5RnC+yvQzBJB/z1OblqN6sjEKHxHgMgFvf6SDCcnyrn14vgwirI84Zp1+cnt
74pEO5Y8y3czUWdO026P4pk9VA/Js/lm7E3RBECDXHJbFy31zlvW9EhTK1wMqavC
hT9sIbiwsly5HyHc6CIRIlOpa7cEPnQ7KRwCaijYCeQxYe0aCbQ5UqNwAm4fsFZ4
9DI8neAqfabAPfTLgUAX/o9eME40IxRw4zg3hjPHD3c/EcZNFDV12ia0JiIFZ0P0
bNg6Oxf4m2DHMr06VXo8ZRx4VQpRC60Kff8F5eHnPExN+5YGEwEJIRnXuwR240bl
mRCSC6cyaNNQoAwAwc899kYSgkDBwd9IigZSfzCx7nCUPj9sCgFIdsdG613S1Ob+
65fecOcDvItTlR2/fELXvFP5GG3SFEwCVaF7hvUjK4TEpclWQmHuE4xstzDQDu8t
6Upd2Qu+/aG2nrlr1WfJsAZHQFEPsO/u3Vbi3MRVNe6L9JnCTZxECAuE4BOANxS+
VG1sdlFDjutJ+emK9qKPnHxqfJgoqQDgbrCbGYyEL6M=
`pragma protect end_protected
