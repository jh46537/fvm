��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���a�%�sK��h���/a�y���v��=��w�����:�y$f�*,�RA\��S����ћW;�U���T�Ǔ�q�0`�eѓ^����8YU?to�Pb�I�����9���������:����l	�~�Y���)���L8�|m[P��Z�ј�79Ӄ���e<���_�����^�2�����
v��;�{a�<Vx3�-�����ٍ��/�[�mg������o2����@�m�e�?ኂ��l:g(Ozl8S
�-�CW�gF�5�դ����>��'K�:���ϵA��8�l��X�0S����b&�7�%)����!�h/Sq�㾴.��"��w[�Xe2�.ƿm�?�g0ۉ.�*9D��>[ˬ�?]#��m�g+��;��Lb�W%��"�����n�F�`��VW��th��Y*�1 ��a�|�!D�+�iN����zط��S�6�:>�%���~c�(t��}��B�n�7��bq��FW"�}L����X 
�~w���PΩ^�k0G`�����ƃ���n���,^;5 ���6�P���P��sP�G{��E�[��.uކ0uB C8,�]܂6�N6?�tx[�m�IZ����X�K�@�5'� *y	�/ô���r��k�7���t��`X��e����2��e�
�3�fJ�����x8~��PK� �JU���|�)s}�$������9���:OdvgX��U��M+�j����72�

!�ML��*P^���=�Md�n��������>��O~W�cL5`a��ZH�ɚ/�"4����_�G	�(����@V=�~C�4<M���p͆�v1��4�&o\����+�?��a
�.��]|�ѳͽ#jԆu/r�LQqͦ�A=̭�<�-+� GAc�#�wWM�\O��	[]�����ա���K:�~��f���X�����jMV�K^Q-�=���zr��Jvv�ID�e�T�q#|N�+X��~X	x1
䡉|g�MN�$�jvn�I�]��{M��X�����_]��@v��A��M��T��y�r#��6r�<�W�8J+R��i�E<ꊱE�_AP���R6��gD���"��u�]ʖ�nF�CiVİAs�n�mi�ۚ� �Lp'@E��O����	!L(���|w�#��M�P��\@:��GM���u
�_�\+�;6ۡ�%4�-D *��ǿ��t������+�Θ����zQ�׫�{��T�s:F���ǁ��Mi�qj®`:�{�^�`��C��v���*������嚌 ����{S|f�@�Z��j�Tl^��u�X��h�\���}�*����۩���x��0�6��v3O�r��-��T�Ԟ!b~��U���qQ���E0��5쫰�#�M(^��I�*J�M����n��ְs��<��_+�|Q�ц��=�4s��Z~�j}K�U}߃�:WK�4��!�m��H���/�Q{��� ��4④�t��6v)p<4�6'����Ԓh����T��̺Ka�D=*�2{�B�?�˥h��,��[��g��Gg1�Z̡$
Ha��������/4�L�x�a.�4X����&�7/�EzS_L<��� ��o�ǏD�a����O�eD��������G�$��a�*K͙F���i�`�O������yy4 �HX��� g �!�w�
���+@�����c_5���c�XZ zo1��	�!��㶵��V~CƍiX8����9�
w�`��I�!sU�c�z�i7XKY���R�$�R~+�c���c]����&v�[x��b��M?^�t��s��G_ˌX1~�L����������z��� %�<4>��=\�6��-l�1��Ab�I���W��$j:T���ə��������W[e��C��h��о7)��4&cX��{��e�vP��
v��n;/�g�6���|��Vl<���J��"�{�2�c5�PhZ� �&f�g�R*��M^�*W�+(ޤ3@rd})��	n�"�
Pw��g��i/4�>��]��{�Е�
���e%�}aN��cE"�(3)Vk��^�T>��~�m�Y�$ �Y�;)�'����)���g��T�j����8�δ���߈��7��]h���QD��(<���r0D��U��p�xB;B��S���
Ʋ鈠��NL�Fܪ����Jj�S�[��m`2��&%nx�S�qB���V�!���.p��4��~4E�2;�BG�n�D���K&���]η��z��+{��6�Ԩ�"&��Kl��!+zl�=��->zW5#���Ь?��-��N���p�����_iq�~�c@F��>N���Fp/��nu����9܈�C��ǾHA�'��0�e�47�wbƎW�l�d�-���	iNJ�/��~j�ΔD���h����ȥ%�	zV!�R^BO�|��+�^�#��F�����l�u�s�8�U~��r��>�?#��ȊaP?q6.��Q�R&}��*s�X�民F�0����&�Cꗰ�����@��0ܥ�j�5��O!ܳ�dKV�k�#6B"\��b0�0?(�Y$�� 
	�D^�w��`	�c���G�΄?�������ܒ����nS�9|��&� �gz�B}K(�v�7Ĵy���r���2����e]�>�û��3��\9ك�t���b�CQ��ƪ(��~ϭ�v�?*Nm��2��Gr�,<�JEl�~ ����O�x�Bs����[�Ö��1Hn()O��g�o��0�E!��7F�pf����Ⱥ�C�^oon����[�4��,S+�OǱ|��i��?�����ցhm)�Hʧ~�1').O�k�.��Z�`��h$���I�od��d�x�6���
��K�Z��G�~+q�q�ʹ��Zp}E��G�./d	*:�Ą*��m���:"ș��ѴF��k/~�6�. �#��^̦�b.S
�Hj��0�BO����G��������0�q�Nɧ�-o-��H�R��N�ڿ\JKI�!�a�A�݋{�y�zp�n!��!Ҭ���!��R9�EsK�SK�i((^��%.M|`Y��З����eG�s����S��b__���v�r����Tٗ�/j���	~�Y���孏1��e?41��9�75��[<Y5���6��@D�Ѣ�+��oy��?5������
Un@�m���V��8;?��sW#�`�(J~�����Φ���↷U����'oD�`�	��2:'��i^��P���Dǽ,��YEyP E@)��RK?�U��3��\�\�D�k>��x�q�����Z˰��%E|h�d���_����	�D�xU_bv�����yoV=���u�r��E������I-��
�E[��nk�=Oe��},�b� �:��+�%\�Lq���VX����(�S��VQ�Nx��:�Ix��opD�U�cٝ������m^^����-+@�����"�?�'h�3�.���}i�҅Q94Qýш^������8������eG��'q��*�w"����D[�z>]��:����qv�V�i8�VΉ�w�$�ߐ�ߍų�3�7�!�<�����9�U��tJ.sA.��k�U���=��7�鬷�>3�!��&�A�=�@qr�.��6�z�aR���6t痕'��f੼�C1+aƜ��7B����*I0�<���:w�Dۍ����W���*s�����z�sy҃�*&)~�d��3~�j*�FW��4
 ���{.vko�4��nAH%�t�r?�iPÁw�J~�DqO����#g=B*��ǓwKb�xt㭲/]p�V]^���K��$If���	����:�"X��