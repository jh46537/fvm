��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,����t(��3�<���W_l]R��j��VqY��f�w6�KK�U��	�2�g�=^�x��2渺Lj����t|�g@�s*��DI�& vԚe�e�x�c^�h���H)��;�;z[<���h��U<���*�n&)\��L�e�m��\&��0�U睌��L�t�<�*K_-
�y��P|�Őh�οo�/7`�>�VFT��5����1��ɘ0�Y��Du�d�6 K�>gLzt�~�u�߸rrn�{0KQn�,.Uׇ��X��4���ai���x��l�)�L'7��
L4�U}�ʺh@�}1s��i;�5��t�:xk#?�D��,)�y�?<
��̮]�h%%i��Tx^1��s!�L������N�Qf���f�%_3?I�������zH+��ּ"Pp�j�pa�FU�Ұ�_';'9����d�@�;-�*;m!��'���{'�rQ�J�����N��<��uߠ���׃���e��u#6��1�r1�?��{�zC���z����FP�A��Z��W� "2��- 0@��v�n�I��� �Ode�����Ƹ�8����I���D��n�)I$�O���(ʥ����!��&�r�}[���.��/~�F5&9�y��4��yr낋f�c$�'nr5B~�7��930���w~6/9r@�#r]#�S�sA���������@S��3�����>�&=�^`Zb�Z��u��#V=ft� �`��Z`A44�2�R�{��|0�!����������x	S��A�k��(�9��ZnG��˵S�x��-mV���8^������a�ք�^VO�bQE.���УZ��+�TG(�efS
��i���q���)�LG�K���kJ�i��k���s[=�S��VC���!T)2���"�wN�Ů��MM�%����1�5R`�T	��؎�l�\��b[��1:��Ю)����Uǡ*��Sҿ�@���)� oY����(�{�?����N�����}�2h����r���� L��u��Q����QyJج�`����?b�P�����p2*�G^�&��7qJ�^����Pgxl0M����y����t.9�^�P�4�I��t��RuY�Z�iM�3��d�!k�Yz��&�����Ux�w�¬"1q�8��nE�Ԕa��^�/�7l��S���rgw=�E�y�<1Sy����a���PR�= ��QYl}�+R��f<�-=Ԫ�O_���qatD�,<yζ�^P�\�V�Q�u;����,Ij:l��w�,-�'��6r^�ɵ5Zl� S�	t�9�XV�=M����z��;ڷm9ɿ���UÝ�8R[�o���ɓ�7	��z���&Ͱ��/��L�W!gl�S�1��g���w���_�p��Y��(�/�dѳ�=�hM��3ٺ��j>�qC%P��ـQ�v4�`<=���4}�VC;����9�C����L�h5�ի��ٓ�v"����A	h�(�T^���[h'��%X&��_x��! ��,����%��g�W*�t-��nq�{깅h��e'J\�!ib��I���?
O �C��=��.��a�w"�8��p�&gg��Y$qt���fͦ��:ɼ�:�����n�]q�A��~��(�bO�4�;}�|z��"Du����H
�������'�Ƃl�%�PYԣR��n(#iƇ�P\ �j��
��Gv��ԸL%o�����ӥ��^��;k���w!ĝ�I�][4�����j�7ފZ�ֻ�{Px����A0��!�ʴ#�~P���kw�Wޘ=��G�y>*L��dIA'�T&u��B�Ue�8#;�@����p��>�t'�wXXd�ʻ�˳G$��"" �\))����-a@��!��`jG�.���sg�AP&fr��P�_2�Pv-���ĭ2���Ƙ�6�ځ�efN�!O
'�p��2�u��7��z�22��"0�jp��J����G>�O�,$�6�L4�G�sP�BY�5��'_66"�օ���AA�wNbTh="���vt��(�I�H8���뷹	(Tѝ���N�7H��V.�5wG/�%����m����竦�(�M7C��]ӷ�mZL�`8�B�9�X�-�D�m�8;Bq�0t����3���
<:_$=����9���J_�ؚ5�i��H�,[���@f/9��T�i�֙���d����2�J"�ur-A���	6����07oV|����D��,	���� ꫘P$ק{���m%���"w����	vN�$B�E�Q��K�v�Z���L��H}Q�.*hܤϢ`m�D�k\1��"��h~�4�M�f[t �o���s4��F]�_��)}�1��o��	���y��r��.Hp��xV�Y,L5`^9s��_���)v�9X�W�ْb��?�W-�8��89�vY��HZ�P�X���Z��R�!.!����9�����s��$,,��6��Y�W�":t u˚�D�c�̳���@h�(���@f�C���S_:W*��4̄4�<�8�W&�������]�Մ�a����Y��fFm��+u�I�5�9E��'�on�o��6��C����p���X���V����v�kǫ��-	BS`�����C���J�d������7���s�@6'�-{�|Z��B#�iL���"�����c�� x6I%�A�ˏ�O-����p�;N��r�*l�~�������A���? ;kx��w�������E�&�