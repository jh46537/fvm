// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SWUqQg4m5x+T2i3c26W/RQxLdSg1Kx6Sa5E5b7F4BAjbMR3N9La67zEVeH2/auL7
ArZUV1Bl5PqrZcXCxzbv3+lVNTb6gTIqrfleLbderzRxvR5ZUGWd+vx4eNLlqHa2
aStNJ8FwWGOGb8tE/qsqaAhXeu7VCqz9G2SOR3fU/hU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3584)
foS+PAoAFsxiFa0E7XOKc/u7xAA0MWA8VLSlMiB3OQUE/w42Xh+dDnAlfrGhS6ap
sAaorUru6WeKgRyWpUSZze7WpI4Yh4Eb0u6H3HYLVIbUThOuxUKWuW1+ke4AXHML
23UHt7+VpcBDFSJ/0ED6ikU5OAElDWQ43xtGIPzUJrhOxLWbrsq81ltKk8U1mVJy
/7J04X5EJjZcQyDsKjNiEHiYWI776kaAcGYxtERkEqhGUWe8oJylzEAqaRAZdBgx
y1SqyemAglmVYpdDdELDicmMxKAUYlI0ZvOdZcR0UyTMyagnjhxUHzgHl8EFEqoP
BhUrp/lBRQ0o8N/VBFdwGkL2hKZKV5NWGITIU04dudhZmfywTGLmsRSNlG1sp0MW
ldMIJdKcIaz5UVz8bS4zszSwYI0PGdFWD2AWunv2VoSXf6GT5HtNjz7rpHCGa30Z
lWeZ+nOdouZ5ktp7hQwklv9Y8jA+1GqBpIRkN3F+KfaLVkD9vzFH1p8HpdYAAkta
VAGOwBkqm/4t5uiDClaoqB4rWn9q/00AN+El36+WqYQdfAJkiJNe4w/teAg3Bbp2
1g3PpEtawdkwqPVkujKSi7kPD1kCwU8ptsQWw+ryWTEIL9A3p9erqON0AtXb5U78
u8Av93NNhZ7fmjzC5f6leYluWQv8e4KRb+j2zEYFOUGeFMo0c7toprPU/AfLMBj+
cNEYgK3g/loFPQcZzcMUdqBaM0fVupzUcYxD08EHB8WQn8q6s6VJaFUvcN4mR7Ti
Y8/XMzng/NI1By9ERYG2P1t3Kz3SdBDu2GvyYFagMHt3vzAfu7WuwXQfhO+TY0Nz
3vjN/wed2WjVWYuaR4hzAa4CXbG1bSfYfaqKbNMnuzjACv94+qcpPmGQ1js7HZti
jrCkRaTWV95ZUPms4vm1o0UyAX8FJd/zprFxAo/4m7pcQE0uAzG5XVPoph/Jh7qT
rTV96P8ga1Dj9xCas10X6czjbqlaSUFCO3RT15321ur/47j5rXIWgRAWI3EPVK/9
XV3HbpM0fygiff9JFMRNYOspNVIs+TSmfN5xHjL/qMlgQEJ5hHNVH+gQ1qIG8Nsf
Y7rzhaLFiEit7hQRBJU4pBljdQgRVkBdcZZUMi9EnY8AAF4RW7s2VKEiYUw/4LSn
ewGhXgB7pWuZwXJsqP6DUw0HeUd3L47lWdlnz9m0hdwbqIncPD9wVOe4LYy/J32P
Py7ZeBe6OuMHMWxC5D+O05va7X/x4+mTHO5mAF3jWgYU9qvOSusA+0VH5S06iqek
qIbxhSoKYVDNGpNk0zO1ZzLIXSbg81gAUwk4LTm6Y4j/p2wxVvU7ANcVMT08Isvc
jR7zVTN4VCm7BvhJWrghzNAPnnRq2kiVCIEGL32YhbzZ9AM3WGvRb0G2Yd5jfbyP
3YcGL0/BI7BmMGVIulJDt4vQf+rW+nzIUCqy+WMF3w7tVok1T/5wBubha3OyQJR3
VlWerLGK3U2zcz1VC9EYCUl6gXCIkBNJGS9t/At3rsqfjzBp62gw+7UDuZzXVnlv
m9D347wZh0hJu6ehkB/xstUMYLKvxgI0pe+ttwZjc2u9fOIYMxqacdXzKLIDkMsL
BfXDvrh6jKQ7khdn9MWbt4BK8syIHUpXyB4hEP94ioDCvQ/sU2pYYptvFGIkwvbC
ejKqDDSjWx4xoZdo3omBZzSyC2ZpOKqyzN2mTSfHK155qsaOUbGDQub/3vOQ7UaB
+NL/dnRJHd2ZfX/WoiMNUXuWZkF9N2WFbKekvkGtGOoGWgr0a+ZcrWvjIIRW+ntN
c+4kQGmgIc5tBdmzOeIl3SMJPxr/KYRhuIKG2xHyWMpdres4ZplUulF9xSPhKfR5
TsUFEFkVo3dzwgtDvWGE8dmnbSktWnwQC9krR1I8g7gLwnugOfMgOV6DNRy4nWZM
M0BCRIwr/3bUN+Ego49iGuQXwx5l6/OzTQuTPRZKNoXZV/bQ8Xu1h0fbl8vFefdZ
EDXQmmpCxc5Z1zqMYV1+AoE7jE1rdXh0Oc702Aj938WStNbyuFqDdOJpGCN4Zw44
FNJY1PLRQva4rPgFWTotqv9CKQz3x8ISAiSpeHXClsgBwIwAeNagswQZKq8JNLGR
0HfD10vomOH1jjzGPHlnLvz+P8wb3wuqH3Ocd7NwKWKTLEI+3ydJaRa4tdE+cf9/
C0BMpu2/vVgSoqHZKAZVjWCZYMYN8MV0WmhOT24ZYkzs9NpRUkeZ/NFm7bq229jx
iQpJuYA8o2cgnfzY6Oi4C77JSuzbJGNwCAiRk0IxKCyIhpsJbQ7xutA79HL5Hz/Q
xys+FbDnFBjQLxtSNlFYSvN3agg+erN9XcDD+DMVLewCVY9f+aG2lB6zYDMPSIMP
LzkQQYhgGSV2MwX/ecl+1I41gJOyUc0rP7XWbBy+uU1eRQoCGh8tc5zHL95lcBeB
eycKv/79SFvqN51eY2wPq2CO8VMLpRnQGeAB984+f2fUDYUNm9heBD/Jl+/TtY8Q
4khps84uXs7mWM2u7XXV0j3AtwvXBHrDSBj4Y6yvbWRsNHRGWY2sGIsZoyC+TJgn
sxBQvRVsaddV2KjtOGpXbJ/JpzmNVCwKNgJ0kM4dsC0lbJP7KYVzVGwGjpTvROQH
3V5eBZl+bnNQjXcEZYSdS3FqPmc97iGFfb2vzJls9jiwz1X/J2hFGwq6KwS03NsP
f3bQpqLh5PO09BVU3Z9TAYfuxHxqzQ9THHTWrf4fnXRSZfjaj990uU8Vh49spTOl
mdKQY/ntpRTbqdou3+VoBDlxecl0WOn45MjXFevWmho/8Xfm0FmNFTYCm26LUbd8
FdXSFNkpKRuLOJGeZ/vMh1FFkvXly6w86UekNPTvhig34f7OK0zwSbh47zcwYMix
eQlICTdlTcIDxeQjIDEbEfLTWZ/HXfzHtm+OXXVYKnyvFLgksGOB0TgwJdvSHeaz
AZxCMrtyZk3U3TY8saNDgRi0F5UirDJnuzhtEIFhn90d+EFAh3EHFjWzZX94oxRN
Mbee8FLkEnqeEvIHH2z6V+aoJxlwqzePHLK4J3V96hxs93hsyUvWD5usUN2RewXP
aJIImWeic309lbLO814TIsZVl8PEDcUXEoGJ0epAJNKsjzFmDtuiK84dw5YUfJnx
MY7vsn+DkgLGLBrAuDSVrk38UsQwtZK1+innMqF48yuytvOmUDzdNb5vXYonM1Ng
EuI9240vmoqv/KC4MhUES4eIlBnaAGVDWqd3chdDE6UkXVfWbuN+LQ3BBz9p6E78
3cXP/6VVimeoDoStSE+6T4Il38qtTd26lHL14YITrinBth4JO5DFO6kTtcYQWndp
4DLjtVF1rftQFcj8BfTerZ4/wmXSbK7CvtDAjUqkJ76LlYOpkgB77ia0F+HN4o06
caj9Jv271EfQAuTEACmsdHoZ+jrON/IifyU/QUkW96Jtq0K/OmdgvXlahIGp3mYN
5XG/wXR56aPmKJiGRNHuYWuJXTAE3+U+LVBPoVQSO+FlMSWedSLBpUg+kHdBHedV
85BPMM1Fd5BLof6gWLY/b4BxpYr0xAF6tisJR2qsrK6zkwLirAg4tA89b8jc86zw
7Q1+NpKereaa57WrK9OeNg9Y6bdZDgJrQBUaCAhnimv1KUrcIcdvC65iG6yH8tuG
KO4Qg+BDU287QYaTGXF7MHwu5Kq9J2rAravJ/GtUBL/4mtww9wCodYHCDZttYq/Z
Bk/b+4AkLJah/dlMAwP6m953Yic2kALakhvDskzYsJYGDLOQmw/8W0qpxbs+cDGV
y6sJ/Y3I4jom7Xg5sTj7F4uS+nhzzRiCTSejOMiztr+is1mDUFhQMhEO5E/VgBWu
aptvkj1Z0qjXS2uWc6T4X8UWx1ub3xZS3ysDNsAPwIk+ELiJIfpyV4+PD/WKwZSE
4p+OCc1lFBhjfkmJXSHKYZZv5U7PXtXxpNmF8o5osmsox+6mAF+MQUZadllj0uDQ
+KkfMEClN2kYcyqPUL4vyhX053aUQ1W1BBrbqr7G2c0u8LnWrpRkhYVhkpjaLGLc
BCWwjO8UKGMatF+XHTVNh4xzyfunRXOTQI7UqiskjxNKHAnyfJGWz+43j/XTjSet
MOk7UK+JSxZ8QeNpyGPe1ZR0l7Y9t4THpfehutnjrFAKIy0CFhvatvbG/qnyGedS
k6ilOXbeJ+PNIQETRLL15CsxPyJLEXUsVH5e7czPGclwchxIQvGJzd3ndpHvmHy3
EiUC9l7qzFvBKXdeTtmiPqpi1yISGbicV/2SJI6C0bLa5iVJk9o4amsd3ib1u2Nr
/TsoYgzsvgFQXuMDjyuTGDcmCi5jBndGKIwIbIBVDrLP2o9025UdA2/OBUoCR0oh
GZASgLSYQi9y4+EzHdOzoC96m4Ru4HpEg2rF5e2rjux7EKvoU6S1gVRXPfLf62Qw
yV2TEdix7IwmNx3g0lpGGHik+D5AvCk2D0t3U7PWnTo+uWwKiB2o6tvl4oCfC/da
yl5azFheB8knjOVdehSBfuVYayIb7FZEBb83r2BCt0+JcdktmjZazUQp/pP2gWqM
eROyowdwy4FNx5EBnKJBipDJ+PKhpl255XbK6VZpWPlmCb8bo7LZrMKdXdVC2ej3
m62O6gNhW9adBjW3YwQDrDZ1Kjzn4+Ex7YlLmYAWmu4VnS3/Q8OOSS/BOPzV2Zv7
cHvBwAjghiNRF9d9O7RBJzIO0e6C8KAqperTJnjcogcuPv11su83usc10dzR+2qp
UPwUkgPeimdiR9ojjTPzo/07vu2dE+YL0BP2XPzLZhA=
`pragma protect end_protected
