// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ma7QtjNX4ML4aTXPBdpgXjwizhpk1RZhKa+0qx0PU477kP/33dOOF34Gth6ywhr6
XucONr5wrgvNSN/z74o0XbMypV5QE2Nda7oZXH+FIFIq6ZGk0wb6KoHMpEDx7DPw
oYkrKUYN6RKO0hgO1D0MsDfdGXTG6HA5u9MS4BUKrD0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46928)
f2KEfkKlXuGTg+qpqBGaJQqwE11RTgd3bxznJPGmpPaYe4Yq8cQ05ITWKLgc7kSL
uhLWe+EBsKeskhq1aB/cz/G5wm2o4F4pIw+L4JZuchzUdnF3tB7e7xIDSSpcz7Jm
kmwzQxNYjglcw+lNvkLkMtForJRQ1uB3AvTueNMwecovDnf1yfSTIvX/CgHs7naL
rPULTrDLwDaMfY4i0cxKFgt/jdw0uNW9VRYNK2q7Wg8pQFC01U2GGsQrwN44EBa4
v4aaorUWZRGatS6wnJA5yfJojXlZesikCL5d7YPMsDqX8CcROon7JN5Ijxa5GDUx
iBXwamX4rUKtMK7GmSI2VQeP0OQy64cMkj1IQPi1EBlHsZ9wSkz4hstJNX/JX7R/
AFSibUxRpO0vNWuTpzPhGOXHjtW9jZiJPtzds00nSnL8I7XrjCg4pZSQmoAyWkMf
KsgHJx3Q+gkdoWPw5FvJjkcx44BFw/0I59ToYkhehFbHZ9HvvdKmEzdDhGjrEGZl
29bs3P095kWb1mr35JA9/v5mPTTRf/KbEcAluehCC/zQGF9CcmtdP5y07X+V1rZb
Ykb5YVF2Iv0gHMU1j5DB5sxa/sOJBCX08Cb6pzpAEhSMbzBgi9X2DQlEWvx+dTD6
PxvbcsRfL5dX7W2GJr7OedGGO5l1bUNKhvRMy8XnUB2pP7XewxSVNvvlyVnech4w
+fJZc0UJgLRGzAE7kULeRs836RscS+KV9o5s5xOyMNe/2xH29UlqGkjM9Nx+rQbe
MiPk1nWygQxcOZQZn+D/UoFufLy+iEINezPjRG/KluWCWHnnnfe0YN96OyoSE0gK
vRjP4lYA5LIl8M+sfPJTaNPeOXbBPNRRalE/Pb7mgR8GEHy/CaW0y9o/H1bxpOZR
aMI9fNddhOK3zkBtC8bv78KTlYnxMQnuOLYd/m3CVs2sNf3Bi8pcBT2O3E5IBokK
7Grhu66vzfP1bQiflADr+wbhylDMUluXgqi/3QOMWNBys2LJya39Ilbha4ZP6JA3
+K02AIAGtrtsOUgx37AMzuIO6QVtB27958GwpyTalHI0KCGe9s6AnffVNOMgak2L
6pbdmUUaIxlfyvft29PwtxxcO6F6kRMIu4S7kn0Wu1953XmrFe0mb46xHoDCwLRB
SrLnmWubXIFRMLHgy5FbRC6hzqMr/j2OiEf8eVCR4Jjpry6ILe10Gjd5GogJ2IJq
mgYPJPzdj3G5oE3SkHkednso9+zy21I4lFhJtLOyC9N73zra+g33mvcApiVok2l6
Zy6Dnzil1zapZmQBvkCrRPiITKw2JB8/g7UmmvTeYd5EO4vARKssbEnOtZgwD5xa
Y/Kczlv8/0HpS8TYVXYR4eITN54w79TXWX4nK2qYRCWnlA9Q09RZJ1mXUPVkD1I7
5YmUI+noPEPqTjrtoN2owueHUkarictMmEHzTWnw+g5QXbyycdC3HbjA9wtBDtLV
nx2oNen0uxBbLloOrZ8bMj+lplSODPgrCzXeqLlq/zEYNk7gtshihYmcimCRqfmf
SdcZXO486XCTOWgSj5tU2UC6XJfrDoejnpZAfgaLPOrRgy9sagxrA7e3sCJ7rzMn
wefW9KvqGu8GhaCYwd6jwBUBozeM5sdEeA31r1FxX1AHoQVJyOhz5bBEO/mt4I1S
jj73DYBkbvw9lxrse+4wsogO+oJciU6TcEgPIxQ4Z0wYqw1PPp8/7nkxFyFK6bhw
nX2d/wPbJaCfri4ASIdOL5PIghqaThXNS5ha9r30RgT9+4ZVRYaRuVWx+ty0rvdx
8/0n/nFVS8pzYw7PFrBJvaUQYo+i6N84LgIiemi14LzZkn3FUridLQbcMjKNoVaq
H4wzsXMswytromDoJD1GhEJKTTkdQIswHx9zjxf9zmQQPf5dQ5p4y3l4UORWX/6L
ptsvVzs/MX3Y3+c2Syt+Q+gZ8q/E5oetb09aBKQqjtZ/DjWlK+43FwSdW9ia2iZ7
MHnGa22P/eb2it//PDfMjBM8y8822aYxkzKVLJ9mvv26uFj9qSmLx6dYgXSyZGWS
O/Qkqia0a+rgj82uknOvm17eJpv+ql67+FKPKZCOlHjbXJAtU8l8Ge1TpJvil6fz
vr2NmWGFmZa9YvWiiyoaGGiBjjNFp7HCm/+XPcGMOXKkeonqs9ZM9UFE9NDhrjPi
rP1dx8zic2U1sJJ7qsIOCswUE4J29lvq+VEc+iEsWdWJDmA9ZYO4fpAT1eI0NPYJ
WMTKXTLXgnq8IstDVjp5f4cchxbyUcOz5NoE8Ceo89YaBdEN2ZPc6bXEn9u5cZ6p
+V0MzsfXhK7Ejdd+HkpQvFuu2WBq4uUpvrWpcLEOkZhPrML5EV4/yPI8HXQqIVuK
EAAX/HcYo34q0aE+gFujq9TnYeWjK0KnZkTbAHKuUcoUQYw2Z7zq0W8VnMgbuQqn
inK3Kz8tzW/bvosfgvc818qf3DpBgtj5lV3N4rmOFYu+0lCOMRcQVcA6nyarV7qO
zawX4BeV9M5YUaqojSLEIXCnKbi9eStnC/OziXnU5wLVA9OXCkVwsEStXzvG93Wk
cxmxVIK+5nIT72SNkbzBum/1pv6OmewDHrs99TQWqoaEmbBQ3rH8hSGK9CHUexp2
uSfQSNQGDsSWPUvxDNvnGSn0cGCDDtMOJHb9DbefeaZPjMBbrj6gcvB8v4rxV7Cf
YyTtif31TYvcWPY7NyVFfLOj1D32faB+OuWcNAAC+ySOkawMC/DPNfwddBfsjlyB
YNJBPfyMIZXrIL5M2C57Z5/ElUtWu0DTnzcPf93Z6M1iIn/2wydpPvCUnsUFs8XB
WTgNn27fPL+kxwP7S2RuTWnCA8qVEhhexAy5yL4w3dYdq6nsmzIB6O5vUQT65LHq
8SIYhYmVAZLXBk3AkhP2qBB3CAPxhbAVBGyiLxqecPxbVYPSI8LnFW7FNLHxiHMQ
QeCOd4+bW5JwrXyHJooO55YbMQnNjXRpeB8sjUhtIM8M4BuL5ckV7/G+IOSnSQQK
ck0dONCUI1lFSo38sbswaJUGIyZKpn3J/4moRYDvx1wUY++kMkuve8fN5TyktAfb
yGR0BK1O2VtFrm3nmSz30taqs8wJF52HbrGlbxmbhudEBdwdj27vxcfSETTecGjO
+egDYWFn8H2s7T8sAWbU8gysJvIH2oUnf69MYKY/xzmdGma5EJlSC7OyLSGzs34O
6GfG8DYuA0DoKqIr65XexcSIHtfXjBoVK2FFO/l/H3qx7JN1HyWdjPihPgYiFaEK
5CbIrJBiNB9eKD5GhEeHmQTBXu0RBvIN93vi763MbieAt9owOF0IipYEaqCsaMVE
tEHs5RkTY/uaT4hKBEgZNm4g5N4sQStlAJpYrQFPtQhY+aELhXOEB3CtSb6hXucp
C9vIU/7RU4s6/B0IRd/B9yUrGi4vERy/bv4EpixGLczqpemznXyH7FXBmwzXD0Ni
mmQlUEZn9qyAZlkpa2gGSvBYgTpnsbaKyufxJZ58gQoymu5rgO8sWhMPNJErJz5c
PPkhXRYF6ecfUg8cQ1rNomN2N45wF2riFqBW5jWiZbfy2VX1fKQmY90Kc9YDXxoi
ZlBSkUTYTW793VxXyQB1jiIh3HBYXuN63RZ32zcxUUHn3k+2HqwQ1kv5sdSIiwFC
voR1nsVqlabPQzRZ3vBVMCZoVidQEVvrlkKIc88ni64+eMPFt/uc9RotTN/AF0Ln
EYba38cBNTSXXystfhVKyX9MVa+nXWWR83sVdw/053cnj98JcYAtffHKWwDys+02
S6cZCN5jjSnXkDKjbOYzZynYI4NPf9L+IPsTnjxLqs7eU6Dr+Lr1jkCAdhmo15PO
w6xtEGC6K2XKVn/Vw5J6EYlxhlj/LrvDgH4j0V5iqxDUlibTXvOoMBLhV9Sb0YmX
8KV8N/WpNVVpl0NlC5Wd7Rl2KlhD46rpj3LDmItUeSQvaTiJRIyd9mAn1tISrrpJ
ECfMjec4QUGjWsdO/LcjQqcf5eta4hYXrG/Q9k7poacfRYgncg5dBQTd79/krNR3
auULjclDGAjTTab0lNgNoNjEZL0NigvPAAGYC1Cx+IOO7upQuCQIuzgOxvldeLx8
Nz/Z6sbhiaDofO95xGbV4pA5jKPHIaFOD8YkjNOf7WXxBMvyzmVedKiW21vth6IJ
xDC0Ag+sntpgvspLyujOsdh5TSD0149xQ0/1S0jUOUOe26081BNeBRiweSDqkk7g
w7KZRxtyzBp1DwXgPcrrxfsuQDEnntKX9kPVa1F6VX9Ps5fIRgLwCdOrcw3AlPw3
79c8gnutVT5u+c0B/kGbCE8/11KjJeyGBkrZDLA54OTD1KVL9CAF0oschHtjIs7E
sl8fLOH3B+nV6XJeqsSvlt4SAaHbq0H+MFWUyjy/4lg50bJEQ+5xw1akBeh0zSUN
GfqjEpBu1idW8/ZvaBCt+TSAgFJg6rHNb0v3KTPVNv/B0gA1ebuj3VZAtHNWuiaF
/YRu+iWzhUoBIWa8f8oODBnS6mRPx3F3QYM1C/iyz110JZjEjBPSVqKKdo6POPDn
5UQzvfBPOtRL8q9O/6rWeqkyrk4h6DHiPa6DWHUUlsiMPXPrR80kPZba3ddW4mAU
VWwt/MUh0uRK+wO4SzXLesORFYG63PWsGUYVCNhgvituLhO3aR4yL9VGuYPCNFPB
YNhnvj+TUzkeWF2Cgl7ATyMIypZupyf7vGWzOMvarjOcN/7uEcL0wVAzojvuoDDq
AGjqLGahN3AZ0kVoQnb7uf4s+Ga9rIECPX9QdHnesD8kWNonDuY9nk38ZUvPdGV2
0aIG/gwu2m51opwI/8Bb93x4/XF9hsiBtNd55E/sLCLPASfnGSf+5BrSBSElBDnx
RdzQEKGvaK5UaNS3i829/RD0EWVfcT/UmOOo6YN9xC4ljgWocp+xUOtJUwJYDANN
9I6kRx+SnWB6b6VnzZfMzoXtPMSqBxv3w/obLOGNf/Z4jI4CONJW/rj0TJVfkG1Y
JLOMmAGJOv5uKur7a77CPlZuuQWYneYPwQJ2/ng+uslT+jfznkARBSWA0aVj97zr
YurVw5dn1oDcg8y8jpot1M2LMeQonAp/fTFvCQl/Nru4Q5tVHPO3kFsGLQ/XceWp
Uur3/cYBqTyFvibI6jQ2D7k25pgAqesA4G7me6X9LCp8zVkCQ4A33JkjKJfjI6RG
sAFhEQ1mRw2CfVvdCKYy/Vfe4heoakgbTzKHx648m+IhuCCFcjjfvCLjktDuiwZW
ZT9T6YefeGVfBvy5Ef7QmP9kG1FVCywZnH/XsltlYGipgZDnQQpJOAFlIx5yFRAt
ox1tHCmj1SlX6tLUBSxmO8dkUbSPecI3JUyw9v4xQRkbzKe7LGPU/BnsSRYrrWlG
9LRgTgkET/uhRFq4LsJvc1rQJJQBujFI7X0iq9HsyG1iRIlQ6B4HgFXbDWRlkvUn
MC65dU8aPVFFrGeKc00dCdNikY+HamvE2a5tNKK1dUmeonQmGkoPPe+hb0tC7voS
DucC5yGnM22C+pGfYnYZP6UNEiJSgh5LqrDen3RIpoFtgVSdPAvOuQBC1ugdWXLs
gIMVjbskzr8PPhmp7UoG0y58yNmBC4dc0bgL5tc0FIkbm1ZQl11/uTiTduezW5mp
gJhxPSzxVDHvcwp0+MbmMiICGAwxRcbOZ52uc6a6C/X1U1iNwja48JabVx3h3quz
th+fDhWKpmKmi8kDDqJXsjU0IdKAbL/b8Rp3CKN2ajFnq1pspVEdmLusl1JI+WYh
E0qn1SqYDDk4mGOS02j7xw6FoKLr5w+lGvRHpLc0P8LgC5gNc2pp3kSTDAFFCWHK
+a9okcbrjDEMAQFe2lwJ7BebBjtJz005D8gsENTE2m3a+6/hVygABk4AvQHxjt3L
oxePTFbrzbxlw2U81SirYEyCKtEhlCCCqjjoPAfQTGNVHcgnzEBQqbhb0eLTDUoy
zZTF9OoJaw8RYZ5gLnh801wc5m4EM8xTRx1l/uQoTu/u2ilOywfK5bJeNHHPfBjQ
1RjqizivD/bJMDHhWkb0Uyh3WwM2iQ0sKf4NrR+7Q7oKxJ5GqMSV1HazuOqJBc3G
DkQtBX7qi4lvlFfETb60UqOo22pEwicJpxxA56MkHA/GK0NERSiU6wX/KBumF8te
XZviqbSYzEDuQzH4N/m7n7Su44kSzHX8n0qZotuA8TXjg6iZ988OfauZvh2HnyYd
YqWQZUTWNKmp3PF6uiKEFCNIn4YeJCVSSDZj6yLJN6p40im0dpxEvTf/o1+Jmf7l
tjj+WKAt824W35hz37hIfFb+YeYO5OERFqiCnNFrk90alExk97+C2764/hPynYyZ
Mamnz19W7MntCYU14NTDGMKB7AfYROPuYc/tirBvaLQH3yToMawwdLsRb2wbtrxD
/3jiaG+kpfqwEJ3zP4YZnJoY46Xa+pJljjkUE/GtTU73KgzNbnh861LGweLi/wGz
iCm2RYVPiN2ZCZGzibzpbgY2288jLjzQiQ4xlr2nPMBOFTiarXkHAONi4OG+/cTQ
p2/hOVYwaF7OO/w6jG9aEHyB0wppShh65ovvMztyZlH3dwyNsHOZJBd4wq7D8Nrk
6KuRQbHvpRY+bVDEqzmIxWhvPUtUhNrjaJfW/uhn1Z9R7XXOu25qJ067+et9AFfZ
ZXttnM4TTUZo43fUleD2KUFpRmPx1d9oQ0D4E+/dLY7YxWcGey8NI7hk71srUleU
h9RIJAyPrG7mkM1ak0V1MqgmpTBngEwXbyBj0x/IHDXcSavMYwhr3ZNmHlKMHiDf
M43MrOvt1xBj97WFOBG3jIZ4VVPAMQcOYf5qs966FxB3v/QpRmwc/gYNhw9ZIquc
nu1SwpxjocqFtmCd/ZU78dnTAzuwteS3B0aJp/UXEY/pAWDHpYC85+YxGuqh0Mmy
l3BhZ201UrCEK/x/V6Enzk7TSkze2KpfsGU3Bwez1CtXHrPo7bFMBmbrjyLPZgZ2
H79ro5BpndAzxBcwFk5jrrA/+06JiM/tr1XKxTeELnk7wVQkqhI8csqO0Am8K3Kc
yP17iMgIRt/dmDxHur9IdDXXtku18eoDDD/+MwPlDzaBg96cwZDBIleWnrOexMBk
T/z6tVCNg1Tnd8jiKVnPwhA2zrPZL0QqpDEac7O1WrtQ7hnIMdvaIx+Z0IF+ix2k
pF17yU8Go4CVIGd3Y2IEuKj010UnYb/k8mGOxHGyElwnS+4ZloxX6hnJx6J6PnWw
EIATzd6MTRUbqOy2HXohYkuzwUqIySGbsCk27iKDCZdnpd42Aqzj5YIAEm8iU+/H
OUCGj1Agzwz0kR+HF6sxFvMCP267x+HCPKcVfOzB6Nnw+aj4+wz/2UfE5Vu2Eqv6
bDnPmfaJnLSo5jo04uKmtUM6sjUvs/tbhwOiJFkaKJOxtlBAe+VrxlGAXMTwbFiS
qW2TeEOwGsR9LcKO5fFHyILbCz+DlzuYwSEwJs7sEkUjH23z8SxEbz5n5Uiv1xpm
nMfHI2zb/ECbNkJvsIpUCZlw1U6XIf24YoCZBSmHLX5d/lEKRIRD46SwRWXzVqXU
5InfFYfTTrZupv6oeBxAyNcGRbjclOoOyz1QMAFag54WtpISYeCJaYXTWbfsCbvN
bKj9U5X5UEZz+oYxEtu2cQk4MyJ+Fhwjz6rYxpJD9nfBw4N2s4zVfzBWG9i4nGDA
+SL6BTyyDrXTaZNmmlHjpSfCjnqLbOnxvtN9jox3JGZF1CzMClQKhnGWPco8wVuF
6wks+m/bDiGFta4GWOvKS203CrIUxO9p/6vMGw/RZJwL38ig8l1iQOioANcCZ8Kv
yJoE2ObNcN3YUeTssdCo6yKKeMh0nq5ZNVP8SVrZl7mxll1kgut/AwOEuexCdZrK
kt+hkpCAT8reUPL12GtGaWaEIDaxYobn6tUEvoYa02Sa5TyCjU72fVvBKC1YE4ra
6hI8ZE+ZTZE6e6jQkK0jucvyWNjCWyVvRpGmFLZ/vV8++t6Ygydl1dEP0DKlh8yU
d0gdLdKzu3iPqBn5WL+UA8AvRCDH6NVJ9kdV9zd0JygkEofrcDYh2LAja55e3wok
eNLRoSQIF45spt/zmjW8d4MnJ7efCZwUH52+sDC1kdN1b1Q+OeorqCWSXFc/YcIK
o+0iNYAiiUjGW/1GKNRIcGojdn4laQrvfnS6HIu+DLavPZPwO/B4KttTaFaCMVK0
jBUw+ks8rGfVqoEd2fE+zrOKIvd79QklI6DFiK0g/c5RHxagA7RNJtHPMWa6wkJz
IxRNFxfizgjtgic5FpnMOHoH4mq3iCEyg7H/woQz4J8A9jpvQ/M+pc6Ez9/Q/dUA
ORr9RIMvv1+TP8QSon2p+QIWJvO6zWUUPV2RhfC5qxkNhQEPJFQWfp462XgTN4QG
7jjpk1rSW6JoWiltY4JX7MNqUcdGd2jSM6hAeP3lr5hY+rvoAF9xahXgUTDn/GK5
/22hFVfHm6MGvXKtpXoAGBwh37RqbM0lORgfJB9JqiRZdKQgv4Tdd8W9FvCaERiJ
AbPSqtt0h7aQMw3AGy95ZQAj8t+ElnmBg1RA6tG1of+wwA6neXoY6M0bQMfNy4AZ
MOXAJktxRhvC0bSwN6iG0RgHQ/n4rqxQAlGFavXxTa13BvU/mzEg6s/N8ksZ7Yk7
E5Elv/nMO0qBb0E1r7PaBEDxmPOsy1tEO1h5P3CpUwQxjHW4eaFYmMiqQG3ZRDC/
jv2IhO4zbvMJyRoDg9Yfi4W8cLOq7h04gZRDHCFuWdFMwlfEjJolZajW7011KzRO
tzFFRHmOsgwiG2cHmVPBG9AfZr7DjB5xDdHYkXH36I3qD+ifISCP2/U+4p5ir8vo
lahl8drIkZjxzTFz9LpuuKnsMzXDlHj3CYQvDGDADaEioWd46GbDoI9M9ZIFf3+A
z7PmgiSZ9+UhVPYbL21UaX+LiGP1ZvR6hhzuCq1YJUTixL50AvyldAIejaBGxW42
iCRwqRjqch94OP348MKqYb/stfSuLlRGG80TyeFozDqvTdKC6e5+YoRNS+6KpeBE
lOsO+JQYJSEcN83KLdACJgQM+gsi3mJz13QSU5BNRokv89GW5957BbQ+Nq+PLObA
CoMOdw7ZhTJOEv24f2aNk2pq8TKRZECphYXklYpRWocsmlAs26k/G2DoAjw8NKmT
EczhSDRrxI4jgq9Di20IiLeCWu32cQ8Ipu9g3qsmSl35Zb2cC69fnmXCgQfGwNjA
S4pmRUtjSipNsfWSzPSv5GRbJfVW5N9oa0hhPqfDNEFG/aW82itcVPw/4jSrmlA0
2j7TrsLUQjuM+T7cVty4XOqcYzjhMhpRVqMmbfxt6Uj230UFjgmMB5ITJZKssyf7
q4/wpcbJdAlYwtJUMpWKyce71ujkrhk3491yIg+YypsEjysgT/FAZWoZFr0IwTfl
Y1N1PzVGFuy7ImZFlsW3QfuFfUNHGXRnIqF1r3ZFkboigFlY46WqHeyry/bTFW31
ieuiyp5w/dUjJFBgYgA/mwhv/wfk2QVlflUuB+j36xxybsJkUjf66cQztJLJPViQ
7UmoWRsDbmdUz1YNxMeuFt9l4i88s30fpuH+2hI0PG1IzP3diTJmZVEsPBRW5gPV
tvI8KZC2ezbDyIMHz/kuHKvrS1LZJPOZO0yvJu2SL3LqEP66mBHhEx3FOC4EYBZM
oxx2dwjsQtKSr/Hb3xrHv42lilN0IZ5M1wG9IBMLfba7e/MoCI2doO/MBzA1Zmpj
ZhR0YbpG2QRZvDltnsNvHE8ZYLmea89z/IsYmsnMqxOdIBpPWi3ItHSXRCl65pLj
BwbUJAlX9xrzHtZX6S1kBQ9NC70f2fy6Qn1jlETcw2EeU9oizmzD4W/M9H3EG82L
48grmIjjSfdI/ymoaoUTA6pPEoSxQ3xlfh0arZvOqWLGvqPkkk6RItgA9hLE2daB
aEaMntTBq8E3zNMfcLN9b/5mM8BLfPbQIcyAlw3WUSUIfx7o2cykFHPvcJUJLyGe
RJ1ERpcQDTnN5q5Hig/g1aq1c6+TVLIEikt1zt81me2henfvuoro+qj0YH/r+53q
nIlP89XEQoNvP9FjOxRrqnFX9Wr9Im6NW6od52+XpuVEcEtzfa/iG+61GJNPXrn6
HziulMsjHQEXQ4n8+TM3y6h6tNDcPuODHjHp6rBAk6FZbSrMtmXD4At3ekG3xOiv
6z3xac4ItmZTyOmFvrKfs+O+Dw/QVVdqLZBxb6X4Pj25yVKZ/Q8SLL1jUUsbuQZE
vG3Z15BKkdwaPkaq77QiACfqYOT2rnJBnLKmehcv6DTelWvW2AkGgpHy2IJLwfHU
ypgbNRF4P7zaEJEKCtVSWLmHM8BapTdzeLRQk++aP9kC2/z1dSBobsoQI9uPKWDi
RCydMrLqdKpOmhUqzkviszCmy57RFUplrAah3fo6o29kzJLFlGMOLhKLPNQpSzf7
nno9+zhmb9Cx+1z+lhCKs0sO9aIK2B7/qFX2fZKS1ds2bbnvz/vVVjga00uVYqcp
C/8APlfGIAALHE494/uwqcOq6KEAI1mN/0pI2huDjiRPVFX07rmY1o4+u16fdzoG
k9fKSvNz2F1u7wglpC4Amv8/+a3CrF1rpZAHiRQz4dWDwUp7jPU/YExCj63ZoS3I
s0olHXwQukm5L1qyuA5SBgEbDxDQWcSwt9gqEQDTLbas6vgRlk+ZM6JO/CpfD2aa
uJfTX5SYCIghdxrkIxVclAf6/hf69FekctXMW3D6CfId+1h6ncvQE/fsbwBMvZPo
Gzi0XW2WhCZbtWyE2unfZnSX8yMacR90biYz0gkIbDZIex15y1oFgBN9Lil1u/Fu
53o93Kv07pnCwBP8S2ygajfej9I2fiJfST6pb79/WlQlMjj4Pb87741/biJelSgJ
w68PCVqo3ktknRBo/bO/OvXm4+6zaY3WQZTS+cSTk7cmv6P79qWPbZw3L90NKfkv
qYgj8YeocWEJ3jZ2B7HBDGNGPfOgbJZhZPbnojUOLM8Gw7fLKXaQMs4lxlpdnXeN
ThKBZ/CIMy1Fb39DcXuEXKIPxnjtR+w795TK9GvXdq/hDwJCCOQiqGa+Nwrb1m4h
JoPFxo1+Nh+DOP55Pgrlh3cSMqI5ZvrJOnUZDd5CjAxZRTa4Ui/oHmAPJ7dd+rsg
AdozS+QGNi0y1Qj6rRYP4FbUCb/f00lEcNcQQx+FLNqJXwhUfiKrwEtJa7xU8ACZ
EbJWpX/BSiv+UAzWUUN9Vtpy306CWf7aGkgL55QxEvO4w1Gkx7DdNdw08cw+PwDP
UZ9rGGlqGumwfYjq1xxijO7cQh5XVe/tr4xMcDBoIS8/PDnZL9ppSZSw5MjGf25g
h+M6kFgSUBrSzuTkF39KXdHWgYz2gwRbwx/g3J8putnOQPR0+sF+3OBMpiyQXtXs
pAVy3jo7kxIZWcy1aAo3Y0dCMKOkizRXr7KOvRhXv1wppbOOID2vAyNf+F23ury3
zNki8IAL4yM29eTWqSiNifsSdA+1rKzjEtp/yzysqHyjAPbKaxlgbdJKCtpBf1zI
FRLXYaHMbSoED3SNVJ4MTTep+N5QS2hQYQov4fyfy90O+9364AtNUFZTmcLTSUKo
3jAvJBYu7QJi8WlFYP2kMmtbonTCtDbtabjMM5NRqqW/gqqK9cT8a1U82UUVqfSG
LK+elh5bC8jEGaBqY8bPTPtPSVxV7QmjD7RDl/gdhNiDEVVzkiVXstCsCgrDOi2A
DVYZMPItaWF95gq7GpzKsIi2JXSweJGLRYXlZ7jKBxUQWXODj9GtsSve2Wxon0Bn
N59xwuUNAcHzuY2Weq68Oi0xrivsooUALAzdwOxl/YSUCK1004DM65cOiNdU3fuM
PbhWpruJzpsdfrIRnAUXdmu51IasDM2El+syCyAXV8eAvCP26JB7Ny6Bca2OXeGy
6iZduj2ddoVNt+pnF15JLvsaVGLEDkrTHYlMw1rEFPviNSmRg2akGKKThBUtPC6h
yqyNv1mSmaNSPTb/2asCUI6q4SomzhfT73gXsy2xWqSc8Iol9bgPQOt49mZ8SMgw
xAqVxcsJSiMWBCA5YarM0VSssA3Qb9P1Y4CXK9PzsRIw/EOPMKHFYc1AtvAk1Q9g
TsMoIpBeppwlHF31H5SmfP6DWYKe/085PDUHert/mCTyqhIp4fOLA6FOxVJHZEDm
CcJm9iTld3m3jKuDqaAlgcxcvEelYITk4UaerqoJCswCAuJDl8wkBrWdHb1duqhD
IO7c2TB0RhOpAVXi/bBE6XMY/7AMgYsMaAj4zbWFHSW/z+crZI8x+yKhXkcWS47m
VKo3hSEXWcW5Yn3GnER8pqB5hniHAz8T77372m2HC/YAH6noBCW8nkLTrfw8WJ6g
KxFpLZEklihfdTA7Tvv3Uu2QS8+7XsY+b+VVvx+WReHWWGWtpcAhAgJ5Y9bk+AuE
FpgmwDSI2RpeBltMfP1e2HQfhqf29QkF7RWJBoIYbHcokzhBIWF398H6BhOGpVMx
8e+O/dkeaglR7livcMv4qhv62xRu37a8zvOh2uK2uWgNH8pkWGg+qpTs88jatc8W
byGptEonexj2AmfuXf6ZVcMDoDwNVXIpOhokf/SJ/RsdFURLWg7OkttNnKzK9Fqv
8WL8Z9MYx/HzrRDtlszjOQQOCYmKf7NeAm5s/Zi3JJpBe9ugeF1qBpV64PwHidyR
q4S38/pjCrStgjoZBwquF52BryZetJGYZPm8UFKitbV8bT+suHKUClifeo74aWe0
GYHURbBxLF6kCJkfK7ot39azAcLwqPaVF34i722S4cM14NiSwU4gMYUp0dWf5mLM
sX8tTopbXitmP4q4pVLvNYtLduupnIaKP//eEZa89R6gawwfhn31cj8Yftek12BA
ze8V+DmcHL8UF4ByJDEYK+T43bOjIhhtneE/BrN4F4sptjKZCnoGwupxr+c32ZYT
SJUwpvpKmLX+gHaNc6MjDb5Bj4CCy8x4mTrCtV1LRj4OgWwrdy8h7gjnO2IQ1twF
vvq979bItN39O3EuPJYA4yY5f7rqc+q8PLnN7saxYfpBuIfMTHiP85BXNjIIUinT
Ebmj8HFw+r9EED9gwmF0ADoUxQSSOhnxR0DOMUujPYLlLEg86E+YDwf7R65b/XzG
kJptZ4sracSIC3ZsCaPrMxIcnwDcMc6K0bHJcakIpLSnzM3u/bI/IGNwFSYKYLfQ
HcqophJaCfcK4bPu21G2YyuaT7/d/ktkTWlcTVz7nng8XbbmXrNp/yPAECTQbQTh
yYXQSpNWPhlTiY61FaZoxsFNChai4PYIU1vVEbDJN9SLahKDX19h7rzIzFNrvQ/C
KrE9Y5lJ+IrUYE5TMTrs8Zux5qYUx47eLW8d9Ukp4DC9HdENtxwepjq/l9FpaC2p
dEImHwED66QvKzumMCjZTl7S7Rcxmq3s3XnrNgBxfH3JLElRRLhIxwFy6beeJWAD
ByZBKphSBJptlhSI3BLy1+Ntf2GwCyi+LO1gcTp70yHl72NaElEdhQ1WnENhAc4d
fYAoYe7nYVwaryaWk0a1/VsBJmRqx7IQ5MBfxxNnddu2jxfiPqaHyQwcDLO5ymet
alvtLr/B4r7lSzQ4+HO7vFBDHHJckSNfW4fCj33xv7rFAQrfbvDvekDJH46K8NvM
d/HPnCYu7pNSd5Emiz130kN2hQRPDf8Mu982tX6NzWbg81QVWn5BJohM2u42xNIA
lugW4uHxHVWGgL2dYIbgpm5TBCSxWgktcuyHkL75imimRA6d23dF0ShTXChmRMHr
meP3Vqfb7rJTb42dJGtbgT9chTR/BnuHNcCwXLs34A7kpD2BfIh4j9kU2N0fd7+3
Xs2QiKl8bIFZlqKtqfpUcGSfZZ+uuE1jNBM+J/9Tg9EltLWhTmdFOdYBIhGFKEGt
nHW1mxlRQ+dUFLLjrkQc2mdGHbzZsatpgyZ/0C6G0HAjGQ8MCNaxq+fzjj3kuMGS
D5lE8cobWxcgHKKakgiK/3Fqrm3PykGYpMZUHjEXIZfu7AFx04XO+YLNk+JmwkGt
nm5efi9w3KFEdBGs4SJMjPX3YkP6w9sgjS5EOfjXRfcjD+sULjkoC8Y+SM71O9pn
ngzliLJNKiqmSJE5HQ4S1cs38ok8mvsXtY2Hn/0RzWJivFNI7DnE988o0wfXRmQ5
EFgGlYOJ+xSr4bPoE1JsL9UUFTCE8rBbNK3FpXbUwWs3A90kApEXYknSwBzGtXIT
NComy/Z+rdaCYmdR/CcdzNE9d23e1QSQxmjOH8rCyzeXhiF413924iT5kudXEN7Y
Mgro9b6SSk9gWLklWhtO7PwxWtj+g2kJGBRIJ+YEFb9yVmsv+fxbi7/2XZcYHLU9
WHlx5qz3GQCcRbnj9yqKdxdh9zQ1A/OmHFZqC+uquuihkEuLEnxefhCan51Dqj+e
rQxBgmuLs/PoUBMrsZqk9cOIIsKyUdKABht734CJL/OSBfpZhrTSytYDMp4nA4VV
ZTQku0zs0MMSN2UFxmMynfpKd4Y6ypWGXAWkYcKPjmGl/my2HimdoZpi3ekP0GJ+
8oXgJCdK2EoiWEzCXYF2q25utHZz+ktm+wt1VB7+SmzpMulVmdLexT0FLc5yjPyr
+eEUSb4Gb6pPWv3njGocYxddLDJBZx03xwVersPeckLLmahlO7tIaFBj+4yWxao2
CmGllP6iS4mhLeDwuSj4vfUSYuHSeHYuxHb+lugnqZux2nB0AXG3v3oVGJXztQNN
A4hRBbZ1u7w6+9w5TmQNo5Ir8lQy83frPKCr37yyDxqAdbT4/eGBM5VXsmiUKAoU
aSf5PzCwjw7pOloaxTArGTWn/kuo+36+AKyQTi6joshHCaC7I+z7LWue4u4IgFkz
RFgM9koCulsTIUIpAqBu8CyMtaWc4ZA/21BEG39m1H/4gBA6PBczjW/yDj1YsHjI
Is0vciWmTkmNqWPF48EISDatVmPx7pb3dv+WLqiON8Z9WCiCwMHaIx4I8jgYDLdW
amdrKp4qL2krviTT13mBL82k2O+K3+i9d370UDfa8/Wq+oVqt253MUZfVwGR/wca
a34KlYkRmqZzOFLuGtB26iED8rChzBYjcqnxGN/ac88Uhwl+UwmMcLtbU8XEw24d
KsL3Q5Cr0fVwRX19/+pD+MDgy0XI3ibEyFrQKDcjIGUehndjEkVVKjdeAMPRls62
hfMc7vlearHE8QUGbicSkja0Wl3X4wefQlKwgyb1k3BbpJZ2ybsZ7mL9dxN98CDo
r6dsKUlUS9ZU0VNdJcIFHyV2+dEGyfY8HPr4ypHZZ9ObXfFPip766O93d48pGlNW
/GVRYLKpGw+RQZCaDln6mhgLl/YbdsGLkaKxRf3ossxrLQIML32F/ub29ssUOg45
9BZMgtr+MkklN/Cp0J4isBfgqpwC4bA/+J3n45G+GJRTV3y71IRKkcMgrgyN+Xdj
jWMR78KYxtywci2fn9336t0rg5H0D88k7HW0AftBifcYSBspgJJF63zj39GvWTDv
9AJ22FEMsbwj7ngnk7YytIUe1wmbWy686/gnmodAoLKkXv6InDJ129N+HocPG4GI
EM0+RFl5iOD8JDv+iZkGV+27X7sjNeLk5FpaRZ+cQC2BuyXTsdvMxszGZdCGNxLl
yP5y7OHPxJ6KR+YDgQ7ikkpGUm+lpLpjwnDDORLxPnSsnoN4pB0bJxT/RxEtwHxr
6pSZfJBg3TkJ7v26l564GWesMgYflk2nykLbXTzrZiixgzLQkPU9ToF7FYdRYyeX
eGyQxWY4rCJY4d89YLeq1Qft3vdAm8BThA23FBpOPC/WLl7btRDa1wZdRjhUmm2C
SRI+KCeaLvgxkdtIQIX/VGz7kksu3vKTent+R+E/qhOtUCgqlICCKc7wlf3Lsw8E
JKJ4u9H/NJm4RV5WOuHkRIe1KmERG4SEChVQaluosnkw/6AVX2GAs2dgb00NqVie
BCIFtskrwaR/cbwVJ8t+m77Vi76AmX0NLwAwwMcooM4yOdT+Kb/5sxmOXwo9bV8+
zc/cQZts1DJGcGPqNTHP7WYXWMX+kV2pIUwW9AYncVrKXZ4kYq5a6MjovwvWh40F
8uziVoeuaJkOQ3cTRsKF2Yek/mpVaFgycfvmUOwJF0nifqRA7s5xNqnPRIvszI/2
7HapzuCQr1/TMy0tnw41/w7XzWZnB5yVvWdI3uKqQhyceq/j9qvqS/ninw7jOg48
6I0EhpTt0u2JgA8iNcaIl7iM/fPT5Yk5waIdHLpkplfhnK45qVTOhd2Ma/M32n/d
Rzdoo8X2jilwpIoYhNx6pWhv6V3bZzF3OXKREY7M2P2LCb0uSLs6/qxPsRxnP9Ln
r2dDyMn8BESanp2/pizl0CW/Olmww/PmMb53y1GpseFdpV61nna4vMsThd66++DV
FvQ2kD57g1Pp4b2EhPCoqfwnt9dzRDmmpC6e8aB/1efx5znUyDl8oAs3D0GLikF5
hgApGV1eKCgG0wDQW8rPiAqagor0ITYK+KP+vu2QAJRafehd5tFjCA+vd9tmvp1e
50D5CwhQ45xhp15qxPi8FnJ5W5fZZIwjIlJQRtbBmI/OVO/LbTE9VjsWRz594aJ/
Eb0DQHU4hBhMQylvSeT5teEo2e42Z24FXCKRgXt5iQwmoCRk/nkDJeqgl/iIKhVC
icjF/TaXx/uxAGlzhlc7Eb67VchiOVE7QcE27kxGtnzAOskWIGpWVJut0Fhu/GFg
uUwgijNAqSLKc+O+YPFj9+sF6dq825DB0qZcetXDZp6NhcxL5ZaUy3HBmjmLLoJe
HNg3KbZglBdoZW4MZ47wz2L6ntRatSjVP4Rw44niZk17l3zHXsfJJqSVRsF5HVkx
8THTMC0Zw+zUaZ4ih6Kie1nJH0kXsTtyoj3POQd9tIOBdGd/FrBEKVgrFtfyvCLf
KI2LlCiKhlsLA6J9jULTWygufEmtx+K9VvBd3ZU7Or2Xxat60wXjxHqaECL3k/bm
h6WvGatJQ+Dvzd6I8/gzPy72rLd+XrxN+aHpEP6DlzSHvzF6RHnjwJn2LyMqrcus
AK3BmsUrogw4xzTjk+HUTFaZx8K9uvJatdJXOZGoHOzgGrmwBSs+MyXEYE1nlV9A
6VorP4C2d/gCu4h79HOFq5ROBgny9ewAZQWUfNTt/bI+SNhhlGbFuD5gnK/wqJFD
oDO2UpeiPf/mVBaspdI0lAscJ1KAmGp2lSCzi8EAyD2RtD2ZSESCa38Gsg8LEci+
4qDBfbt1YlyypFTerf4/FAS1u8McmcBc8k4VhSDo0BWF6JCzzMmk9cQeSg1/ofyK
PxyF9nsikxW2kMQisy2tmqYOatrSjsfiMwWiXfKNWDH+aEirys4DPz4ZxiYDmi+Y
j2W0zY5cl+27VJWX7Ci+OkI7PYKEA5UKgA8K4re2XNReVFThor6mQnfJvaodwfQc
q9TdWkbPJSVrrbt9Gtjdl1Y6Ulfmn2GyhBghG/YRFr2UX6iztPAOM1suISVFEexs
jNFKFznua6d8S9PqKATlKW64mD+lop1NbClhRRf5wVQqjjGpdl3KTFccwNEnNdUY
iSBtpmR6k2W1qfvo80JiEY6Ju6ex1QCkfvPnTsLgJlNRQZ0PhkwmjjYhRpTrb06k
Dl53cgWYUVsqAXSKn7kx6oaLC4TJGWwfIRKEkaE2zreoia99mdtyTLZYomPv2zgU
AUByEZ9L1bKXBcCfvR4Zd7ktQIQQNQAUT7HpBIusArx3oekIyw+KmMqfyXMKLOuH
QvMFq8xX5eoSAqo1BYCA01mxonFCezL8fvbBhTRWcXapB56WcCNSc6tR5drUjoe4
l5LBGBZBp2zzQT5YktQHAgxJX9L+NJkxmz8hfUqzazdQu9K1ObGz8Uf4jTXSAX/k
KNO9MvKeBmEKKiDICb6LfEkgQXKARtcKHeI1Lsb7n1TLcl0H69ZMVqYkU/T6dozE
5225/whHrGsocaUaAyLOCjiPtedpYdg2M9g+Nac39Oex7nBQey67IupPEOZHyTnu
eMqghJ8vAICWpfb9giamgfAEAa77a5tsLK6DqciIuqomHlZ24yDN6+sJuZDiiRf8
7U/BEDAQmbYdgU59CujYya8cY8V+aP4sTh7LuQ248YWzISmducXlurkGtSlqlHf7
ufJkMT5QYjO9+6lGTm09LhpvGItfYHnZgiF33b8+yAuAROd0x0EI6bR9Tu3OqWi1
Qxi/qsaFFdXsltFE/+65vJHlPJm0zRiSabkN78La8uS/TQnGZXZzk+kqsAuJCLnd
2IpmMcDG4ZD+s9WJi9QkBdhIG11cuWrnulSKWPOXQLb5AUDjHuXBcMLZpa8S3nEd
X/T/Q7m9Om+yYK2o+b/FxDooYV72grVl2gjTTvJO1erabAs6GwwPvaL9FCtXxpcR
2GuJXDxkWvcmZdsFxizyR2x546XL5/aAIyhgBB/JKTjOCUVAJdirryrUH53UsdsK
yPtubeKPKXJ206CZswP1W3jaR8UGrXFNUklyu+CtKhsQz/K/odWymLfr6BTeHzVh
KLzcv6GS0HBs5/MMVdVwqbqgjrhi6Z9E2s/8kxLG3zrWAVuOJOfZUtLUVihzns/+
tUfmbdcrrGFcQXxGUBs3rH63ksxl87HaPfW3e4GYkB4ZgrO64REaq5k8usJh1xGA
gcSIxFpifCyfg70WDHG2ZLoB3xdJYmBDsRLCDlWAftfDY8XE9vecA0ypdlT/+Df0
aN2uQEtbjUUawdrFTuSma0wlozvtxTiGbS7zSarSYuGH/IEFTaRLygG5ju6Tv0A0
vNlSbBy3fO/2lj/MHl4MqhVU3hpqodCq5YTLLlM4wDAUXX6CtCRDykqfbiP8tDD0
fi8d5pKfUwVu4vKKoV0XQcLZcdRrU6RF9JuH96nwOvS1WswZ5pDctJ8Podg/xbH1
p/B15eL/sNKZZgt5/nbvAAo5tEqek9LVi7d7keyOkTKyb1ZVTHGeIn5qw9QLJe2u
uHlHhxejj6GnSMtDrvsGjhQFVOnsCISPk0sL2Uh9ngDVGTVPHzXeuJ/8jNaztgF/
DQE9XKlt40tDf/G4+n3m2eU9RvVCuL/PVUM1P7N/Tk5VBFxhhf3KPtyWqeLwh+ft
3aonqoo3l9+74h4tePmGg1IRy4TR3MfWB8D6eqxyseM/SvAw6almm/dgPSuQTQfk
ALKfyfFJFQxfD58O0Xmr41qv3EcxzY5w/czI25FI0oemmBcyFbeHr1StKI9kRR6z
UgaIHy5kQdG7r/Hv0JyKTg/P+pIOYEiLD4oK77/bEP5qwhFXOmL8NZNfnJ1cF9fA
fLNLjj449LPqnPWEyfu5pYSxITBCj1ujvZxv8mxXJHluKeOibPYYRoIHT+F3SWk8
MM+rgOaohyXqRMGlYdgNMALGUG5RI/0GbPShU/S9awaXCYIN2n9y0aHhk07JJjAX
eWqF8Ieso/VFkqrOSSGaWopomQFdD22I0b7MNNNRC+AUWFoMTzHyidwkPQDVEMK9
KO3bumhtwpfskpwadEHURA+GV1dMc4THwPWDLzhtdrrLvZeGCzcqI22cM8fNndd0
DfvLLw1YSLHLgC5SSe5ebsGlfDO8MFM/9bCUki7twqXvGe58yXF5lfSUktCA+6nt
FCzvNc7bMu0xK82Nkqw90sqk8oHPgxikVE6uttWAkGkaZfAkYYU8+YuAX/Y8TCVm
u6G6DVWxSFPAIGBWXXat66aU+RrrAeuBvZ5jnrDMTTPm9/4+gBmGwVblvIOUNaqW
+C96ZvI/tv+0MjVtbFrQMtue/EmKQF/38fXD3PMA1vGgx2Xly4QdVacf3993SPGw
jEo95c71f4t4869DtjAy7m6KNnBBDYYO/kx75AYYs++yEwAcYvr7lxq3MRYlB6vG
pM6s/cL4Ij+YPVtpwrakPrpPt2MIt3fLHEleDfO/VV7OnGr5itECdjtMiNpo9gZO
6QBCE1MDYb7rZToapSqDYPu4IR//m6tsUvM7cPuZJ6JRWOblDa+oyrRnkCvmsoVX
N99WRSTWlSx6M7MBPe8BqnkyKReQG9c53AOn+iv4hBRNT2b/oPBNUjjcBcZREAJC
rTRfCduFNoq5BT45gu6eatjw7p8ABHSiRdvyX4V9BZcUD/v5uGKA52ZFYV5k4cbb
rUTHy/62q0vn7HUhK+yS9wHMXt5xe/X7ldJTnrTse/c03ouS4jCkQUQhRKWSf/Bu
rUata+7aMVtMtn4xt4TDVuBJopHCFXj/l8mY29V63A6D9tpjBkqPCExYiBa2vyOe
SrRYTSx6MQcun0QUnbGh553Z1ACfCTyfhffYFsFJamHEOK9600R7kf/0JP/yYaaB
s8Q7thQcqXIhItclQyncutgzVA+2WVtN4Rxr9t/AN5hJCkSCZr9Ufw4mvHj3ptsn
WCzjfrvhitRzu2CTVUe6eR5ZaDwlkDLoOE0McAvo3dWJAGKs22etdjq1PHV/jLBX
AYjuISDCqd/6tqsZEkHFCqxQyz14cZv0uy2VKcX87ez6X3fyixZYigdO8CViS1Cc
IjgSBaR0beFJVOTedOuYsyRyYGWnBTS6vjv2ZlzwRRcX9HqlNy5DidTQyR943CO7
+fJqZqgZJz42elmBbgKjn4wW5y9tInNGb89zR1UD60WKATlMmaSOLQAm+xZXvh/7
tazdcvQPCG0DyRjDWkQaJgCAxrkM/ouUOXWdjnUxwOkpKlSt4gmgTUjdHH5kyDLM
dp+YvCKEDLBaQ6REsxn+Phul36DNlccEeHgc8ZUepQO+t3MCdxorAp0ZqMv4Defm
R+paqRLe+Be6XmvwrcbMpinFpfSFRtqske74p1Y0XgOyhjnQOyKec1PdGR64LvIJ
ndyNeNE7GjlxkkmLO0zmv5k9stGUmD/EFw84sMWgu69PKApDSczL0u+yM4Xu6BFQ
m1f4qEhsLYTuW6EfMWUydtDS7XHl2lactvXKhkHAjcGlgLWmyTwW0qBDcCsQWI6X
bJ/KhL2q2YW5ktrXLVbCW8Na+Qt3rGkEC+CvNFWcLDZck7qy0cLVU26VhYDNIbfA
cJjsKhabJ+5g/S1zcw2sEUWJemeqkaCe7E3mD9OhUEkWGAK0ZrBLRofhVegTah3R
SEGDPF26LNh/b3T/cQZw2+Y795IUPvPlaUiLP0K0TBt6LQMQoZy6824em108wsjT
vwBQoaXb3AGdfYPutJTvveXzYyccRNOKAEmT11Bp2DDP7nFW0Q6aFEgG/zo4EPKx
zHbFE+H72dEgwKW0NJmjXl0hh3dblImO3xge1tG6i2AjaOnyCphmbmriZWSTZWok
aHeW8A+ecqwxXO6/eJmEbs8lliIClzUyaZ3V/JhxtL3iQb92G+WxCiDzXqhXsCkF
M3c3rIFv5bdGmBiQkzf5zdkJNtCjP0GPofzXbuy6dLnPczU6RsMoeNeSprqhfoqX
Vwe7TOkvaD1hJjph5wEOyLWlB/Tdj74ix2MU45X7gTRIfPtRyq60nA2g4ROsrW/S
U/JQxyJd5nAKDeEnEfOfL2CcMPbq5EVEL1fQen8a33vqXHCtJLMDMCKu7yTcVhgy
JJFowP5D/wAXGcL7eeZd+Dqn96EcCUTJp912u5YEIu1pVZ1mtEQB5v0CXK2MZqZs
i1GhlPIUxQdXItyxPMEWKK2QCezNJgL3el8oCd6m9qAr9Fc7YoitmE8sLZUdMrVi
ilAe9e5s2/nqiF4yP9Sq+ubO6ZfUP7JGCmVh+5szef1tqfAKHS70nOoYICvgu8ad
q7ynR0Zf3o8C+6hG9U+9vl2PWqj7Skaz1WOMD3JUoCrTZlD1MO3PZAk2878LbfcZ
AQ14FQNviSrw1TCM06ykHFnIO6q7w6jCdoJf8oLTPh3tsmQLcfQZ1kHjUPZqko3t
NapDXnLuRliv6yjIC1yWA3iTIKPhXtSdFrpKVNT2pkmys3DKS5HWa/fCtuJNvL3f
Vkonou2S3l7K31Y8/zwQk646zr9RU/TR6+1rpwcKuw0p5143nDmfVC0VcrkhQdhm
BFfcvSuCTC7XhIy76HxaK1rnnfNagtMz1AXPu95MGhuVzQjWWuK58GoM9Qc9qDCw
iHh02nKeAz9vFhg6inrKQhJFZe7gT2IzZmARqgXVKBy8b734DN9xJvatrDRAAjcw
L6K8aosWHJp2YVAKx6n/68QFxe4rGDjCOUZcddy2urDF9qLVzI5DPf1G1cfQ6MDs
4ZctIi+sVzYBy+nK0I77MKe3UcAG95EWEp4W4thF1Mc7GA9EApph2jNKrNeVZtw9
g/Gd0rJMKkF1XNHMSHKLtP7o2Hy2dy2nAYIW3/Ry0CdJbeQ/AVDVTDnEuJ7yWjkP
2I5z178Aogbe92wYSiMj8tAs1zsUbsvp+U4vVQCHMtnMdxaBUE36DlUPhiOfAmTV
RoNrULwH7Cb1O+D6tGGh/I8HKmNB7JeMnbpee3SyTCOtH7qaykQ26SREAvaxWHIU
+fXYpyCzyJ8u4LZaADuFTr+LIHwi/q9gPD/N7AykycT+m1QmA1lQrWaDY6sH9Dqe
VjWUK9tJtkiftA+f4pyOJF4k5gLI8STYIb/xgWdrJ9PJhAr5KmhUbH3AYY2ne2Tr
e3ElDBhKi7Cpf16Y1/SLywCNGsTVgBtPiXmc++eZhKQqeQZzLybBG28IUi0mOHmK
vQ+sKcunIg6i8tQwpiazjy+yHY8jx4yWkjnj6U7d498fvSv+AmIF/bCRG2ECKeSq
cGuSaqpjgQwsv4uizBo4SXzJIjnJAukfL4YM6NFYgtPuw9IaxjEfJcL2ma/1GK4f
hf3bYyF9T9G/mdhnxTyBGiEkb4fJzW8MF+3+Ihu5xEHTNbGK/9ck1Fv9v4+n14ZQ
wUsIo4/tbT+tW55Tbt2yP8d/uinfpKBer21WohbEG2BQgAVcq91Zt5Drgasn5Mws
znrVt7nSQXPn9WMLcTX1C3bG7y+oGkgCijcqS6uOfQBOIj5eAO7YT7q8KFed50Pz
Rd402Knl/Hd9BHcY9jr/IOxbjddMLJHeQDIhRYYS2BYvT2OzF9OBJW5RCRQp9z6m
dKqaxjnJiH39OmV19jc5eyv+/ibTKSuAMYZwT+QrkG76SDIioTTM9OxVp/b6WLHs
4PSlBoV8L0GrHX8dPBcpG/xEEJ8bGlbF2lfGJgW/qWau/QfMONn9bMuHhsphMOsi
bgOeWCQiFTqPYOd426DLl5nNpsuP9qUNElZQkd5nq5NgP7K0O1PvZKuSh3sw/kK+
ErwGxu80F69OVj1azeVXgMVTf3G+Y1mUFs0UioeHGTHwvimO0b6O8pRfNb5Yvn9c
hy+OK9jDOHeh/6NGAmAC2MDHd4MzwfEugsHz99keaICRnPXBNAWsg5WqGk5JSKdZ
mWfCmdkUEPO5ei2wLnWjxnqc4I7rcHli/vhm1GpHAR8KeJko2dxDXTZl9k6yHR8I
Pc/BJOkj2cKdvciTtVl8sNr91Qoqv74Niq3nboLryNeRN7aeFIuryZwVjJRjgMXo
JzNVqU9ojpLKjnPT0bUveoExVXNhUwids3GrLdVA3VlcipprSZndMsvUqYDcJcQH
UISoma6RMiSlhmp9hHCDc9ObtSkLyjFDaEVOfF5wAj1ULS3VV6iiQNyUTfBrovo/
rYN7H2XHz9H0rp/V2LAXOZpXkhdzyYlwXsUiMgMLU4kFXx7fRASqh9ZTA7q0YKJy
6Cx3PEIcvreEeLqE0HHAeeIpQrSF0zpfMbOfxSme+Jq7SDXNoxVkMSoQGVG0mlM7
T8ZZpNe8V/VLNjh5oduUMDulcXX2ZGO10QcsgEitXLjKhvwaPQ9wnwt570dKCbcy
gjw2Q8VpG++mK2jmNE3Cel7ulxy7rli4UHr4LYRep35tSuGvYgQyuspXN2TBtzg2
wYntMpWkj8RbS8/Gui7ddlniIVKU1zLqKctQ0YIoY5XJVfLzAzyj3Xg3agq6ISbg
AHVq3xNA8n5uERnyXgl52gK+0K6If3YWwMem+9nU7H815M9YJlKIaM3JfmCzbEe2
OQhgS7pBY7giWWFdJ1bVpkJcZC/YcRTFthW1WndPvU3GOOa8bslmAy+usZtpkAJx
sYmwtzt/ocBjLEk3nZQf4ljw7GlSLPc6bWBb2/D1exbZdMOC4KARhz+yfROvaKup
ZdQ8vQ28TvvlH7/eVAqKERXoNbWjGaR8P9Hw6W+31pPGzjf4ei6OENFtzVkOf4L2
yesxa33sFN2pCIXvLzpQoIc2UxKljr36r+CVF3829v0no2eCBFOtybu45nxbf2BM
ga9suLSrb3zTovGPqPpQ3yNPEMk24obmDGcLeaoYgxI5b74UGTY+VvVI1sByJ+TT
BHKiKIiNr+jBo7K8//2jqial9mpp4gP3Wic49qGYTle5VH8moxAcRW0RAz74qz5W
oLcVrKygelWm2BAuTo6CRrhTrMHSNi0e7dEKisO3gvg0lLtyB5b0jNvoo44xyhTb
QqufzR67VE+hFocnSRY255vGYakCRQ6If55s+YIUQ1mEvgoe1CSkmI+eO7GUPRVw
mhJoTIclSsfcR1mB6dzPUw3iR8hLNcb+F/zG7WyIRHz7Nl4Eqh6ZhcNzrLEgEjL5
82cjdY+suwYAlC6iHaMgplp3qbsuvQ9PU7AhzGov/YyN1ogJlM6FFd6c4wDzKDIn
4TNwcHksuDmE0gbupY692E73BUgGpD7NO5DoNbZDVZPaqIPLF/WvzNwRN7VDfdpM
yG18kadbmKA3NTTR5DjERj5XYA3zsbLVurf3ByD78EdxNHm445SffyWet75QWtWR
fWA7PgQ6XN/K6uyfCrjdcsypcPQd7PKfVzHwLyuGD+0IVo/kHqF/HvAZW/PZMPbt
9ve7PCWISEBJOdSm+u0Lf76G2ykzC2eLSyo58r1SjPDmnaOOM7gsMs+G3T7KY7MC
LEL+hjMHbnosQ1fjnO+Mu8+RLIJs1DCS+iMfQ2pms+oVFGznAT8/cLU6OGymgKQL
rYJFB/Q/UB4qbpQr1wGIg0hRb6PTKjpwi5cW5spncqKMXy60pYpvbPrzDomSbSop
6pQGiDwXI2dmsYLLJ4/wUjrSE0nTBtEHAoLQ2Y8Yl4YsthZrQswrvzGS4fOJKEya
8MQm4JPLXVl6m+enCO/mlApvapgl2IRtZVO6AOStngWMPIZ1+IFijdDZ7nOcGJer
2/TeBtIEKFo/KaVrCa0jcLRJMxWYZJGoNlFu3kp+CxQ5z79cYmOCUIBupElbVH6J
tNrQ033B2CLkzZu2hTH8dsdFDuJhL+k1Z64pvaYSz9+/+YqKQcI0e3+RMC0+jsT2
DAmyBsBFOz33SyyZnvDqruItovgE1a3jsGDNoF9SDQFflhQviqvQDf3wR26fX/24
S2kIL4ztzLnLwesolz+VfBgdw7sWNNUwVaozDku93Wql2SqEQ6Xqb4gRfglWUjNM
2dJmCd5nLa1aN/jnMTiSaZpaea/VAcjjDFehKzRn3AI8swxrRsTTHKW90dnlmFqA
z8iIfwbbDfFxulms35rzdpMkjw/6v06s/0fehb9VAMO0MtiUbvqf9nlKfl4YlGig
oPi3PJu/GGLQfmaVx550QeZNK9JKB9KviHA3I+COJpuucqedFSETtnMOuruTgmyC
xWZVYhkU+YU23f5snjbQYcpFjkFVI3rvnWTtTSoTpMPfTv03OVYTYYWAugO2gety
EcgjDhb9I2v8W9bffXerLnQSyXG68QRqtQVRV0ocdp8lhHgsHF+vWJ6xRKDA34to
T82Gc7hHGTPxnXWOoaYRLKxARJ2qO755Fa5eL7H6oxI7JJAxUinOHzQPOVYB+Hyt
EuFzboTSoDVNeQ/klXOTM/T69hCypxj2Hod3G3vbFmF3mTBZ/NnJKZD+HEioeV+/
XSGuoo8ro3t9eVl8RyYpPd7cpb9szJiXyKJjCXiChr7mwVcklkgwRWiC6bGGZtwZ
2sqnrLEbtTiziofsLtYyyp4B97PYQRpcEXhT3uc6uaf+O9DBfQAKsL0c6PCoiTkf
a0TdhW/QoapMQgX9f+5pABSO5N4QUkJWlqlVsSnTlx0d5P+uq5qQ28ok5XQHrtgj
X1SflbTuvrkkFPejHcbFVdeMW2HYADgN8zwSICVb+mtpTC7yKNZL5vreV5NvpMje
++FXamlaTaazSR4oCARdqwwL3i6Y6fsM+ORmsEaC1lGy9gt8vzU43udksjbhYM7I
T5X6NrE0gUWdsYJ8tKl+Bv7U1gq7JeOSBM4wrXM9lg2rGHk7rgEhjm6HCWpEqqIN
baM0LBDxNE2LfjTx/Fh2tPDVBIV/S1fMBxxI636cGj8T3F0RvPoni+U4uNQG+f7q
tIazL1a5feECJ1HpA6TyPAlwFc9OqOwH0XZKAO1GfdlUHiUFIKw2e1UwJMkzf3Pw
26zFPeT9cMiE5wq1JMn0LkZ4VTjhhscmU45sk+mPqB0Jtc8AFG7UJyR7EFhcOEmf
RuZsaAJsIDQrvfRWxIL+rRxmwOf+NQCAUgA3+S1vaU6/EM8wt6ozpf9py2K8ySO8
qBtvEOv87zICjLMQGN42PixyYOaDcTlgiIElPdSe+ftqfeBsH8BOryw7Y/V+NulK
4QlBsYIo/smyfDPaSzTASm9tOk5akkfSy+E+ApoN8vadlQUoWhLrzlnJGAISTBia
KIL+dv8RfmxLtfo+dam8cTikGHxlLufDbIKJwn0QrdziQ+qQ3cM46GM9fxzUG5Ot
sCt3IrLXBuki4LyMhQ0GJgmG8ChD4A9JRqq94NwxGvAm9fuhCxQXcLAWlQKNkOf1
lMb/Sh/9d8J+r+o9kfnD1lDTSqa3tKWaM5EVOnAUbEJM4ZoHZs+mF+DUgKPGKRX0
iRitFg1Pebio41RWVLrEXNO4saWfTatsUr3ZRz2fgnFYfSV+/gRi/nrUHiQftTmL
x43gIJ11sRPBNBbOWQESlklhz9TiWXYZmoV0ts1xj1kZ9mWSAVkktGn5hs5fQy1I
QQCCprpcR3CGworPEPWNj1jauiNoIxGeBZxzOsb0hKR5BevxW/3QnnI4fZ3e3y3d
2Py50hEfCxTs7k0ovxjEaXNEju/gK0ItpBxveGMnnAy0ipjMwd1dkqvWJCbF0L0F
tGQ14t1wvK48pgR9FIH9s9MqeTLBVpRyxOiOQSMxuRBKqEEKR2FLigSuGeHqV/cy
jCOHOd1blcOVkLOfQMt12ELSLd/3YoqQ+aCPb9Ti8cTcjAvTfbT2QL0l/VF8z02Y
7HkvjktcSQHimkjetlxS5ggY1rg4abQMyXgATzP6nIRN5R/3IfNXp8n3lVN5+n3A
9WrzrK3mXw0QYL5GXHCcUWTZpGZSqUfTtySXm9wOwATZxn9inxHHOJD2TScrHUAA
gURGc85iAN08hRJfACr8gnLQPwoacRtKnHeg5CzVFzCXz0+HOBxhfvzGxDwCo8gX
+uTkl2gKrY3HXIETLnGmv5+hXxVhwQAUNqq0n1k8qIIOpwBqtu2QcyWHs3Te70BO
C4jWVJrjU84Ke18xoiybjVy+zkrwbFUkwQRJdOD1/93nd/URlV1jNkN7roEgj7xV
gOq0G+Twg7Dx0E45iu1wlBhpol9w/xlEN6CjYjMzcYzXa9jmpv+H1Vb4xiX/ZfEy
y04pu4YCR+h/00jKoGg/fNI8sohkMRPAYLY8NiYX3R34ivu/yXPc7LS7nQT9eTSD
a/c4BlgRDFNnb1METBTfhZ/3Zp4KG2M2+++0U2OxgOFIfvnUCr5krk4CBilRvTdz
QpT4LkGma9r3rLll4DMjhl/0oj1kNaZD9uDzF8cjN9lVMVcRUpPun6uQEbEN4b0w
1yCnhLx7BmfAYkGBpH7dcVtVIOnhXdXiuXWjOkM9EucB4YotRBElPYc/MiNCBrJG
WwTl5RquiFQCY+e27QPUJgExvqNKEdWpbIyMtZRUQG9EkIFc+hccD4uCrNWPDSI1
OK7VySSPW8SAZXmb9sUSeODVp3rqJAzImQUWQjwDBxl9eBtBP5T/SwpmfxnrmhOQ
eITAlzHWvl0/LiJHqKV55tdPmLxJ6etIxmKmHgPAdAH8zV+Feq3sXe08vY6fZjhH
ad2EOvZ+WFyzkUy+qSCMBqa408QH6SgZIGoDj5ysSLOTu+EFnbY5dT0L5FlIncxA
juHbsRPHa+Zd1SYBDXduAJXjRq0y0Lwzm9rJDuToVWUtyHO2N2bJN3k1rtN1yzdP
B1f1CxJUSGTa7YUBOuhbD7Z33jIKogAaoOUwb7t9KrW55Q2+bXj3mjxbAghRy7Wq
fpChd2ry7IMG9HRjSpwteC8IbRFxUfhufNs4Q8H4Kz8lhJ020D31lbPFD6f7GeNL
NqDy3kZVt4ob+SVPLcvYxJJ6Jx3rVsFOJHPW+j0MlzYmt4v6bLaewN78nNH1KZAL
LNOJZBOFW2Vi2c3uNjxFqoYDOFucpNrO+wx1kg/SNJQ7WIrYqm5kEc9vuh9logw7
jgMzNLCMeBF7nzy758LZfkUi7IoQ0ww4NE7fV24Eqqgz3H8Mc9BZjuws+SnwN9zX
s6SndrPPqYGUNWe+La5YOkLE+bpCZqsSoEkIB/gGFhKlyYXbx9aiWHDuDGXrhcEM
JJYTaEkMmFm5VvWgUEDKgoXooPBlVuQ0JgqS0yREDhl7/7/LpWKoJuaU/9Oo7siJ
Nkw0ymzXWDJGaCxTbIg2Y4EgM4QS+qoVyjzmN/pVJ7OkxF+j2P2F9RQRoaQk8VpK
L9/6DG4kmoifDGxBTmQ7VVqEZBeC1XbwE7Uhxu3uvbcM1JiB9TBINXKKIZedofwk
XtYWUVrUcnABejga8PT4Ia2J2VNRuWyLoHKovQ15cCgfeEtQt0s5DtkZoH36jJTb
eBSzqdNT3S3YGAx2z4X5I0ZpP+sCJjDrBplLgX00Hgj+x+nvEOfCshZZ4G4/cgWR
WBy8IimlgW/kTMb51Rl3bM2YIeWDSmkx0dhqtSXPfp/vYkb7gGIYNNkiQXVX7Vu7
nVCdU2xAohgmNhiRnT2zEJrkjsdMuVR3y5WT2Xfem5uH4KzDigDTql+mT1mkPxab
beHzThPp/qk15wJK2ulGta3BRdqTLVI97XirFVQg2cpmY9/TyBCoBPREkvDcWO2k
F68gOMBp2rInmERU682nd307vVXy9eD+H0pUeIWX2DALcQ65911hXU+w2fZOIGxN
NaUSTjfkIFOly5azwMfCy+QFeRQUciFbGr6tobn3pwE5xFgMTNrlgKulHXrEZQmb
MyFqAScLCL2X8nhvtChDmxsUEGgsYV1gx4l+BO81Mxurb6AYMygHpEtbhFfQ2fIC
gmXCbKVu6m7XAO23BdVJR0hLxF9TEEN5SLPQ1+dSJiaq3iOpYPo1Z66K7irQ808L
dyG+dzaE41AMzHtM88d74GxiUFIdWJidqON8EYpuJnYHnELK1ZS9VVt7HEidyKZT
1qenD9vCEFqGqZdfo4rvbADyjRtO4DMLgLXG5K+vLECqdy8PixYM7B3L8Bl9oClL
MrY/VCIQwAo+A5E65tdoq0Jq3E69XefwGY8UKKM+gTlEx6loCgc6zYYgEMQhpw/A
INdmoy11fvWL7oLPZA4C4s/o3k+FN0n0PX0cSn3OtCLvIHu0koQ4jHWSVxPUPeO7
dfWU9zq8rx3WjuPXYaRVy8tdwkkFK9Hu+iGtbtoo5e+PuAarKLzjZP4sNqBUkZ+T
2g7UZk11vjTcTmu/jYjNhOx36cKqJVsrPT6h5ftDoK+AhGtSktdsildJOP6l11wH
5RsOhW4oCUtmYBRtZvKZeQAm1zUP2DOGbS2XsBfPulj9NSh9rCEkN8ubadEmhVXC
3UCvViCvG9bQfmHjZB/V22zObrG1ZvT0ZxPu8lamKuRpsyeCVtr8rC4+PvuQ5LoS
RifHYhpGxnCBzEeeXZN01In2AhmSNZURYE7fq6LokqKj3/RBUVB5Y6dr5CsrKAil
kKfJDinNh92FWWeZbCwvCHMb7StH6ad+rdYge9JyiPoFoJ9WITTxPktfxMz/AwZK
j5IYRi6lHvyp87tUvlUTfdo1NTH79xlB60nqBzdXuHPql5BPpiHxIJMHIG+p3Vs1
9fiy3NSjJaz2eE9dUiIa9VWj/l8r/Ejjem4/QIoP9lnPg4fJJDbTgzf5i8oJXMxW
78BzeExBqwc92tvw6viwhZmSpA1YHejG4ksZvWfF9FL+vwD1vrYYDhjN7l4kEpi5
QHjWvPUaz0WzAt2Mt2V10uDOXJl8XSI3NprD2UfYuv2RLp0vg8ondYRLKN8YMkaI
Mb+KzMWeto+Yjtig6j2Jka6mGS/m5JJpldx+OW3kEUGlZKWyxoL+0Q/osluZG3Jz
eSZXGe9kQjiMjQHIaCY679kuIK7yw/BLEwXuxXC5eHbwAOyy8RcmMX5FVW/X8kH+
PAhy8MlDUteiIvw5x+q0bQqXFWtJGh1vLT6pBt2m6vFaeQPjxRECedZWFSAaP/6g
Sqb0tOFIYqdRs4kaJ0HuFBT/aHW0d4wytK1vF7f/3foK0Q+QvPJhLHDmwAyoRtfS
FDC9oI+b5XZ5UsOb7J2PePbpMpHAWIfBy+hYEY8R5ti28fEaBBMxtNk8CA8RE4jc
Ycy9ECptjsvB+TT0iPKSVOofRnKeZRcyxibKA7TYAo90lNE3G6JvJR8Jx3EeyNAW
W25+w3dYePhudbHSnr9luUWwLQO8PUfr+eaZyZWTX4Q5rgx/+qWRjukBWcVnbf89
aePFfvjY1hI7lWspqIxjpmtqNpvwHt93YfLzMBRW9Hcneqjpv+SeThUyLQTIQRoG
Hb/SACFMGnaUIapQi+3QlhPSEZ2n07SGRasT+tr2NkFn+lxi4vrcU/7ZFQudCRmC
l+RnHrI1vAGpf1+/xxPKCQSp+2ZsnOdEgQ1JlzjTmCADZmyjdM+Hqd2NgGmDd01o
iYWkyNtuCs2EXIJGQlFNo64LSGjHOGShVnBhqNVXfbp8Jqx9VeVVjf1dCytmSuOg
wbxeVUPl/1CAqkfeIj3ghTSjmOvjavNi4TdFIKwX5JWEGaF9ppZwJbdRTfTb7AwL
a6wlBXB9NlhZIjckpM6dZl//UcamZ4mCBamThQpLOVEv6wIVIie0kHKg2ZtxBe9+
XUuB2OdRZGrka7J2/83bNxy4M8Zot66rTgzeaV0NJEw69dnLyoEFTItNzYitHcQf
QVCYcUxQt3dY9Z/g9YgqclEtGUtL+9rcas3SxHJuJLx8wUozlLjLOfU4kvLt1dX9
AyPZ107pvBd420TovtlPOK+dDVkvylGM0VLcseb20axjyOGOkn4zRThvYJ4w6z/T
Q7qT+fvfNdtX2rZiNWLCvKQatJSX2JTkM9LGw7MXXgFTZi6KUvNEAqkMgctU7jff
s7ehsbf0wVLTEg8/aOKZ+Ow7M/X0UFqDd6y99rxFhr1vwxp3/JK+WNn6unZfgSl/
TAF6VJLfJtB+Tk2K7pK6QWjD28vtHDwaJELvQl0ym8X2eTcvXaZxrQLXzlFBZHn8
0akvo8sJkhLLdg1eiEddc/Slt2mOXuC1uIqLmzr8jlyrkniTfsN7+GoDKOfh8CWK
r0wkV7ULaOiwaQRXT1zbHJX6X3E5xrel/SFuGxmvJwE+NxnJ/CZ0gc4vBk70po2N
97yIKV24PF1VDxMOkcJIpf0VlfziCOi5rLfddPgTD8j3LJjSjiKY8V0jD7rNVkvB
ufYGBA4/5+SWnbMARjXJhyLGfGxMlJdvjP4BSb2eTlxZwcR0zsCuNw1mvj1fNcb4
9aOEIDfoqyMfnirAuQj+GifOtCKYSxZ5r87zyLIvsl/o4AFF4nk+PT+gGgoG7xVo
B6mrLlEqVK//n+VGOAMceNJeFDU7woZkjDxKle6CY6Rp/qzgTE6LfZtIb1W66ltF
vpXDwPc7C2Rz0fL5ViSZBoPP0j8cJ8gQfo7ka5obqu/ZKVmUGZIvPLrM9kdw3aLU
NuTUOh1bibO1EOUqVhMTNAVG8eC6OqEPVI7J77UDdmvitKa7d6hqffB+SuSRZWOJ
fIR7IjXBCfcC3YO6FgB2lFG+2fLQ066AzpwAtL+YB9V2g17eyTbsUJureWItTE7i
hQ++rM4KKVpDtvm2jGdKtJrop5TYTiN6GCb6JHXTQ6JFVSWS1OJkWcs2D++818c3
HDA41DlK3fq7Q996GcxXxXZDAdSadgxMZFfNKcSpzpFpw6U6G7sLHSywmbMbsO21
uxhCJoOmIPl1tiUTqzusdPL8DDtinJ8zkEpPY0vuqmzmReuYb4wYe2jpbSlnGu7B
zVjTjqh+M4AXI3m9lhcbwStZmMpHWia8awofw20n4qT1MgBHnDN5hWTDetl5xYPL
UQ0aWJ3/JEKQ0HzYq/lFwfuDEonjU9rQjFt4jnGZmyprU+ddOryh2PKPlCBgFZ6+
usAGgI6dOgaIan2UwM7Fbs3++IDFabcLy9O39eVPisZEnfZGyTaUJoLYuoAodEKm
Jfa36o5eJcibLMYqHP6uwEYj2hR5luD1N0wmsDnp8N7NmlNHnb010pCPGu6lbJDn
wTQqN9bpTivBkDZV3g+qhIvvLSPr+3IoSDBxvLJgNAFrMaV1TvTDQP3KaoteACVo
Z21VeE222agaRy/lrIj1gVtSK9o5O6r+uXgRNcss6/p4TUAu3lTGHjoVf3M5OfmX
w4wFOFQE7feIMG3bG2g0SHTdqD2H+/etZ85FXhmi88brOftdjkO78dTyvaVpy3cq
YrFhzmRi33kI6ee5Rx74Y8XmQL7ha7Vq5XmA1Fvtz+Xqj3KjEEKw72griWnUhtQ6
boG3gPEvDFLiVb2v4RpO3p3q2AQkuwOA0iVga4BGyHhRqGdOaEWetib50VR/kQoA
+IbjUBRKentGb/3VtKoyE8Z2kkPbsBSheKXjS0ytGu1wCdKKJLZ3aNdXeJ0QQLxK
cJcf5l6jd0d/rsyBpn6eqOPXMJOc9aeyIaHOdJ/pnhU+QoGpn30/Oa6CJWkQBdxk
3ci3y/a9x5F7rlr4cJTLC0hcvj60L1wAEBUMwtsvm/4D4sMNFyQZvKgMn2afbEl5
aT5L30tQXBfDc6zbxularWnDzeZJwo7lET6qkRA6Rf3AgzKW7EFTUGVkSUm04WxZ
x8dHFAgxM54dG0KXbb3RrHn+0orU1uq0qRLhRuViPY5fwOhJEaNTawbsSyaIU1Eo
kD4GGst14yf06umExk2M7kn4M92F0vaV+3lxJB26Ake5y36c6ZxJexu5/6NJIf2C
8z2KuCoff7rQ3/mV2k1CXYyiAD4qPzP1CCzMmiFdVJ7IFKRXieBWSHJPyslr5rwc
Lk4Tb8xOH4hWgAg9R95FCIaeP0AcWhM1dZJtOwjcPLT3tphpZHexA6RBs3WijjL4
Aessyre8OmCwgui9nYVhXUDDKHhxTpqzzfkfvkBQY271DgKHCiLbCupYp7+HcfWL
CRovSuQmf77eeJId7kV0oC6SvNPKg5Y3uVhLz4OHgii7PgA7RRCdr0hIMniqxBza
ULgNx+JOdq94e4O82Y9xyNm802uHL/AprNmxR2XW5CSOfCZamRPBKuXQuTDT4rnK
KydNlNDkJs6cPx77EqzleXsneev/Ee07v7lrDJrkieuVPP0nAmgGDdepBY2Kk1aw
R7C6lMmYOqAv9+iiQEqSXzsNWNXzzfrIyPcaLzzsj6dtRLLBQsoQaz55ddRptHnl
UCq4CGRORrfj7N4gm7b+904+bRn4soiwQSnMM783ndAiT8O6tiOogjZ0Toh2/E40
EzS6wrT8YZwSUGREM7hd8Uvxqi+kh2yS8lj/0ZTIngBcPAlN3xQLJMXHzEVE/Z0t
ktR4BIWlZu5MAgr4LI1pzy/Xb23UjHDnh1Jym4Z222bvgcTq0G7jnIMXsLqASrKg
Etd1E1VIt9Tmb5+XxrmyTbv5eypukzYnUC0KixutuMC55j1Os/B39TnKtUDSw5BX
AKgmhvXpeKNGVIooRhQdpaLcOvyQN4QiSWC74YMotFAW6oYg7CSs2Z54uKQ5ZVOj
uNx+uBLE6gJtsXuhHbXEgjghbTRiPqFQxXhkX0TIyFFVSHhWzl3+wVygGQ1fV5qv
A+HdCgEBb3qdYVYeQPU4V/Q8Yg+dyVGSdyFkPs+fG7HYEdmFF399mxlXUFYaB9n8
ptXOMCGqSdkfo1GcabvFv+k/E5BwEOvpxfrxEjwRhwc8lMsnO8dUIpH0AcEZfjN8
13Ft5oE56eFOhcZvVCPW871QVpwBpBsMq4N/isyA71Ztkd3aRng+nM3mJTK98TEx
3g+/ZknMEkeZ3WtRYFG14hD9Gh4VweiGsqTNAPs6n/S8rT/tve5lSpNC0tvlYX6Y
ZDW1/Rk+Z/k2JqiGz9kzKWO5U8H3Mb0fCZzCyhcAZj0PG6bYtJVQxZsSk6MFgez6
cMdfyT0yl1EVxaz9TUoF3QjXT8MjVFbrkke8++UF7LIUYLgL/ow/gKh2lq0WSNIm
Qd7EoWDPFn6G6aCzE9epqumaUB2qb5ZOB3P0Be+NpJeG9pe7MJp9AdXIe+7EAETQ
bZlWCub2u+eO30dNKx6s3FW1n6exKBZYSRXTg2lonjXP15rgNjhvvJwdpN/WLa/p
wZ6INaj/ig3ACk1AhOqSxkUwsTrh9Vr9XnQVPVeu96IbaEWvYMC41FBmNN9KSf+j
TgTWi3no8r7zaNvisPf8Eb7rEW6pGNUzl+8cQpOOC8BwUoqFyNDeR9+oljBjZ+F+
LNKoeN9PPV7KPIjHy+m4DWOOekjqe0oJqrZFc5vtWK1cG2yzXWSZXqTCqYIHA2oe
5Pu1VNWa9i9CPFKgiEwFIAfX4TCIbJIdyYV8ZnUddXDp+THzQCzvLKuKRHZA1qIc
wjpnVgOLtHE+2D2DgYlhV4MQf83gaDlGVEDJKf88y1xHAWNMmQ293G8EjvswPeLh
jTj+g/qNpFGOvmp/SWZ3p0psL5YKoqBmB1Z3X5FOhgrYoYqU2vgfxiNL+y65yhJL
Qqo6sbDnnLprKu29+1hsRC/UAzUuHqFyMCZKwg9EHOCNZ7VxIjz8mx4cNQ8glIlU
xfWLGI5Lm/TPxi5bTzRYbYn3lkSiysqMZKWLYAjgut3nyGf5+AkMV+3DJ4vjp6OF
3vLWB/jkqE+Vd64QfjD1JgoGr3Eit36uAmseCQeXPI7A/DfkWMa8O1n8gug5cAEi
blRa/+IcuPiJZdat802aQAWXcvHNjhe3zI4+dtcIeBVCQpORSnYrl+vJRr5ISKfw
XuJchyqc//Aq7xPj+bOrZydc6TNnKh1oMaFwuHd4BXo3XNv6xL+OHB2I3TWjS2zf
zrRbnlG70e1wtwsia1J6k14SEWTK2GI6B8vIhUgreAcqww3TP5Bk/kROdeJe/yt/
0Dk31h5M4uwovxSt8cFt9vqzbCJpon6+JfVZ+Ysu1y1IQUl96NHfeKmCnOYOWgAV
uL6otJc/RGs3skwIywbUTK7yVXLA0KrRaa+fu84PaFn0Gv7cIOYgDS9zF/Gr76FY
SN5ce7DED6Yh+dFVREIOZb8p47VM5qxT/7lYp+jpmgk7rJWq+FGeN6YddM1IoUnt
rPODxqskk/z0RJ3qKil2ux8OnvqQxN+CJlaJNaWCMsFylOJlfRoH37xC+3379ks6
S4pwMoyGdA8H3Kig8+AfQwipxMQAvp1gE+KTajqi1lYD6zryjbXV5mxAwyO/HE7X
Mkpv97ktTOpaCLwSjTONJqvCQnNJoNXldAlsxyh+itH1+Zc4bCWDw6lnBx5sXwKS
wCtFU1+r6ZkVsm3uy83mKTo2XzGZTWhLCmfOHFS2WtAcc32EVaPuj1Cjt567PZV2
lJi3qwl++FjWwkmqHRkuCrfZH+WKd+6kRFjglOrXwwFmDlmPoEHhCAM5kyKMUAJx
HXpFQYLFGNg42t7p/o6wtTOuOzVBBkG/pgHKp7SrIRYvM79x+0+uL2zj6dUJO00S
33wukhHj5FMTVObLhloYp8yXKzOWFsmh+sRMutO/g6yWdcBWKe3UYIo20BJ1F8oz
Uyqj6xgLhPf9VRbjPUCeRvDetI86ez1Ze0W+noW9q0FsvSiLg0cjlTVxKPELt4Va
NU3AShusmnFkhkd0iQsYsMDPJWwANqLRCdIs1dQdPk0axLZf2Swx+fg67yym6J7/
1JvcPspxYs6IyhALRzYa6KviEMg8Zmmx7AtiTDugDFEXgQdNsHr1ugeLHp1e1qBD
ylqjSbPBf8Z+bp6q2auUzf6onMI4qBzHWlWvh2C04X4hb88memxef7keiIVmenv1
rhFQj55QtcFI69l689+V5xeL5ytokwU9D5bv6kdOOzNOstRN8kJWrz3bb5b0Blyo
WlQcCup/2jbjZ9883Gx0kihESK3SNYkh8Ar+VFKyn0J/n89eNyYiScjpFsMQf74p
tzGjv2Lv0aac737tBO8jTzYn8CG147SsFvLTxfhQfGM2AiKQ2xprOn3tLtBZAIVH
x2dLZG9erhKbgSyx77ANGWY20giBokZa9lrODykFGQif1NS1yhl73p0rcst1vAWQ
mD8emjqYmwjmiNO15xjFS1RBtrwVuvicjjb0sTqI3W6A464KXZDjH0WRWpt2sAbF
aqxghNKLmyGJZ+j6SWFXv1p1vvPDmmaoOwhxOI/Nk71cmz7S38UWMU7KnT/wCUa2
WSsE7vGxtqUHAKHun4SAOqTcOk4LXQphdjXIMcc6Qw9kCRbmZzVF66Rh0MvEyUpi
t0xDXNIfK4f40tBi3hGY68YDwiw8kacoAmC53goWNCHtVuqE7C4giMw5L/LRA9vh
7vVseMeL3qXDWSx1hQHgEU90PABD2Oz0Vh0EcdyQGOSHBHcMQZAmaJqh1+HRx5JP
omSlATwKglNx0XfUW5fxSRePZ7qwGwM3DagNg6bCqgBiz5jlbBK2LJPDTz6rq4yf
tCP8MCFUgQDYgtCXipi9hAzneIq+tl7OGE4DYS74J5sLVoXIaQODCqNHfeCJWTc4
Cn8dqBxTjhZhawyQa3olWh184ckS2N4qoEj8EKtFHpXMjLARwMCYoW0jIzghPcWt
a1VO9UHaaQcMWVyG5zuhKvdOjtW1LDKdtNNfHSgdrx1wJDVBGXlWs/skZ/6d6owI
LvfMgH2J/Lm0WjkY4MWq5NYBn8K6Mz3pZokCtKiEdwhLKFgUe2lB0HMoiKrh0G96
X3vnv9g6s7MW2UXiyIzidB4577YnQje+OfdQyHq2hM3XbLTZ/xQgmKCST50ECxiu
O9NHSiVHfttibWUL1Gk8yq0SJrE3ZhPeidNK4E8vddcg5ywDwMcJgkP65+aAoTcr
UTCWyvY1g0xp/2XMkgiJGFeUuY4vJOXcWWjjcdtJ6wAXMOGj56644ckxYX2/fLIy
4379LnpTehqHdmCGVV5IT8racsn67bSJzMrQGiYeRYUR518LKY9ttC44opQ8KRKX
D4HykDFBS6OflqlOmEENyapjXK0NsmQ/MZfK7yEdg+fiH32zqx69JqoSpaoVSaws
kYH/DINSV3K1WkPPfHj6C4s0RCnqh8sS6YdE+tyoZTlUmgV/iR1HUrDzWl1KLW/1
DZXv3Z/wZZtvHHpQmuLp6SaCrmXhdEVvvfpGH6iir81tdZHdlrvW4H3G7b6kVCrz
G6aPPQ1qrMGMcYPsVaV9Q6/iKKU7jdF39fI8i7xwJe6DiqgwErklLUwjEm182H8D
ebURdK8iCLJ3BfvoC+EPwncopypW9LrG08Q78PI9IvspFISB1znqA5pgTfMBxDG9
mpy/FZlsx34hWAHOUDeQhKSX9CO8qNuCFbywRQtiAvOitW8jsqDmLVdnp0eWHRaX
WqVAbUDXr8WYJO2x5ndp+hoEOYuhnyUMC+pXCYMuJHGstgGSRK4NNReBK08MApVu
LcabtRs3P9gqHH8wmbafXSMr3IWIfsiCG5pc9ufbY2oIvsQ/Yql5MRZxlu4WjXF4
hwZb5MnXSrC5eAWXsCQPPROveaUCIRMJfCJo1fWrMtM/6nYZad+39+Jq2pRhRBge
BpXykTkKgqwc8YB0fTUT7eX6KJk/+k+dtBmzpkKWMSWNtVgmMFdM/0CEfz6JDwTq
BbI0E0gW/yWtlk/Hba05XbtUj4zmeWQYlyz8T8VRBMc7c0PgjYhhoStYixRDgtLx
TvG6Gql4P7oR54D8D++0E70saC/2QN3n7u3SifjPWKtvpSHVL7b0+zA3SPlSTugD
pTdEVwdeXOsdUmAta0DrRMwWwI0RE4hYnGkfCww8ixuBF+Bs4jFY5ydOHbxOueil
T5meDNTK73crUWwW28CS6Cg+Wcs5WbTbyQz/0tYXZBpuui0wxU4gUe3AOlNNOqE/
yfFHbxewm7XBe8GbKLUxvy6+PeaBg2w3d+qeo8Wf03rQw/eTnJBjtSuLzNaiWf79
tI/Jp/GcHmBNoKiGxFyY1G139WxU3lGo/yWpfa1Kzfpl78iLohiA+qKwjkUisp46
OiTJXyzQMEsLlshHu3pBkWOmra3dpjgL2srBqhD7UD2qlpTvokan91FrP7HwTLZy
l8CDMLRl6nZk6caELzSBU95dG/2hT+szXW/oxp28dzitxZNnJEprSRWOPA0WWyEv
MHo/gSkFfGbJhdnR7Gsy3VJMMlvY0E6++OSmCqFv++FursOK/SDJtx2EBnukhqwF
mOsBjlrd9ZK1RrLerwabyHwJcQ56g0xt+P/kUKkTFRIJ8TTu0ZujrQnQrlMaMLBR
TfqIocTMTt4lS8J0yMEasH0SecKGw3IYhDevCF3OtKCIqv8vjyZfgQDH2C/NzPJw
8KcKcfrQvfCFGYrRGxAHo0ntbwNUTdiWP8Idu9rWHUGDsVb4MnANPEFnHJUPJJAr
zjJ24btzzKTZspXfmNidOXw7f8VaVfeYrjclwW2jkk8lr2SixYVJD6yCjK8k23es
igfsjwbJHeLP1He25GjteCmJy8Oh7Ia1dMzZ2mw5sgHIXSqWqAJ4Ezv/G9VCHdEx
IpkXAXM863GTLFyxGl8P5gDJ1pV8ZCnLROz9MqzxB4ANI+ga1uVJCCRvNOxGqwTI
xa2WHfIhOMIzmGTQi2dXYA1QcraIrlB90jTpY4ZPAJWHBfbRVIqRlUBavu1F96db
PdfJESaD/OZoJ9UkyHrBD6oYWGqAUf7GdgNwVx0kkPrFVkRFRBzF2jXm7cRa7s9Z
SXveS/df5tWeJOeSo7BrRtQ62Q0hjIiyKV9PkdvwifW9stVWXd+DoPTFAk7J8ktS
EIeZOGcW39e8J/e1L144BQghHsn1xO7uhLgMPpv4FHIKvQ/g46x8rzpQ4GxOenxo
dS5sByZtGzjdq1pEXpnsbiVtaJu6x9/GUcKPeaq9eVzgIa00IVlM448loz6yF9j1
FqW3PvelztpLvpcuRF52TlsUVc01ORWTmjhsO7YjldSbAHbY/U4zsb5oZUdwt1+R
cugzji0iPc8Rbq2Z1nSXXt9G/z3FljjfwadZlkA1NmoyKBbogp+8ZcE72SokLcHV
mQiut5gExHkG0fGmb3rui377FUjQEL2D+mSK7WSsGTce7IKD9XKaN3IeKOMcjpt4
ZqfUzGaSt4WHzlatggAaFvTEsgy4J5jEOkJWQq1zuU0qj1oMkrDPGIV/OObs9c9n
RFjsH0aRgUjLmTotscsJxsa0O3Z2KM1mqhkuB9GYD77hNlGz4laMW1x8T727GEUQ
pHs7KiTji6bqPAW4AV5oJa3c9ynORokxRnnG6BJAAFUY3+tK8PrqTTEqdHK2Zfh4
lIRut7YoT6/Ww1UiHIiUPQJJUcH4N+6eU+PMXPQW2nw3ws5MxPIQVvg/tygrOpcv
oLEuzdBn+/fu3oLJ0FNZ7PD9Ca99KCT3OS1cPsMwkYvI6oZpCEa/N7Ib5eWGlfAD
w6yhDM99wmOzE3o7kx7ktd1hqNfpCBO+lrgNBQ6UHvO8QNjDxlQ/KNbOG3zne2p2
hz/hl2v/nBpCgaRGCX31LddQVXrpjT0IyZ4tfp6Cc/7QDqSplvu2G7f48TBJVbvA
qVildw8Z4GyA0y+qjsumFqEeYYRxxUpnHq9LQ6IBcqmoj3J9xLbA2+ujtYyIllZg
MA43gH9u7pqcV2n2nEW8WeaBbGKUYSa90MNSvVwVneEQYtGRnX9hynmTNmF+MiQV
ujb+azrsUio7xrmRTg5tDCGW2QmfZs8hNrJodmICO7t4tHB+ZYzFIHfHeFOA/OX2
RQWyhqPYpmX7E5qb3gX/F27Jf0cDp6LCJkdrHz7+Q7fkt8cHXWmx5YfE3jWiTvmh
QPaOUW6ToUyUeReKx4ebSYYM1aWkfw52YIALrYLXHEl72d8/7onV87VR12q0jLNg
T9g2snforHnAxiy0i02jR/oeOG6V18dCZZpm+Wuf9/nG8m+KPMN2szuviNTlm1m6
Z8iqt1Md9nuLizeawztvqzkxFvdaT/aRUZchsRd4kj0835+1QO9eBlYCdrbOqANQ
bC3cXBjwZZNdrDq/LmaUWlPpK+VWGPM+oQX8lrLCc8KZSkMKMOU6Jmccv1mPw2Fy
Y6M4pDSAnxwyzhWDmpJFXGgC1dwgGxiwBnjMwLSnW0EaS82hdkg1PG+CfORKcu3s
Gm2ivY6IaHCRoEdsY9Krf1gPTksdN6ExSCpQuTcbiHSlzaCmjuCfinmOZqdqPYJG
OrolS+3wg7v9HCDm9pgopIWFsOY/vz0657QmDtlkNBHH+mlpa7hXKstQywkzk76E
of1e1u5UgG2cTp4FJWF5g3AdgkDvZhu8851ikDm7Dr01a2dRyrsV16GlEMMt0Lrp
yaUa308KwFouBLlv5NdSkhzqnn4k+rP+2poE8QCxz9mKm2ccJR+A/H1uN96oN5CO
cjbV1YLjze50trYmZe2KU9GtEnWBnT6kiWUV1oTemT5fRqbj3qEsuB3uWgZWRM1q
QRVacIkU83CEJ0MxwEd3UJ8As3B1uHsHEB3dwoy1LjKnVZR5xoxEio9JmAkCaHzW
s8m+K5oNxnFSAyHrPi+OCdJrAneyAJB+KCx+6B7yaphaSXJ5w5TSWY26d4slIYng
RJrQ0OZVv/jpTv1BCNSxIBN2MwCm9RYi2Q+hAczy2FIpRZ7MbYxpqn2uQV9+dfjy
6jB8W2wFIjWVYTBeM9scxzlRoMWPite9T8a653jHwqIQgE5+WtwJwIpszr04wf1X
lJ52cfMY0i94euHB/1H7cVXIbxxoQXYYkjr9fN6M8GiXSTwF4ZPrKkVMGeRK++Ql
u65Wga9YQGvkNYXyFSM+swCIqqAeJweCJCE3sFF+/ZZzOCdfTgl7y6GX8T/YaOB2
pAnZo56LNxPZ/qSO1KiK2xgaHhvZ/gCStAHeajUzqXZvUwNObvlsGtuwDwDXFadC
n4s0W950R3rXF9borHTItENCIxrjibcP7kKYLLrm9aqLGm/D0XukBXs2stntyv7L
Drp9WG1P1c1avK/tQCj0HzLT052UjxhJ/BX1Ko6cJruhqphkpWoDXXSgOBh6+ygN
AgYDuKb80UL/dxd0eokmBKUPdfc3DLGXcy78bg2no9gvicnTJkKFsXNcpLirhAGP
BMc/8ReJk3CDgtN31TTTqQWx1+ggZSIJgRkxTerr8rLiIgcqZKaZ7jkXcpz4QAMM
x7xxO1FQsFGrY+Bk0b8FM2iLdhJYWpvmw7RvD43UEKKGAyjpCNhWzR90XKa0sRda
BV6IWdt2wRe3ZttQAVBUIMkK6mjDTf1m3P1O0+J3pZ+h+qR/uOSejeRgC5AqjCHl
IIhgNA+5EDjwEBwQJWIS9UI7esHCyUESor0gCr1RIR7j+Ewvdu4ssz7oDpo2pHfl
hfPey7M4dgMAN+mC5/6L2euxQ2iSb+AQE7x3H8h1E2vCT79KNWOK6+tGit82Hn3C
Thsje1oMbLFymBRIbdq4hmkYgANKsfwMV8GNWRkmxBl/zZnV9kB+dO6NtsELZFLv
elvbYd4l7xAjwNOny44vbDvpng4q6m2nRZgaQ/ysgXzev6vejAhYT9AgiIpEzOWr
JWpUOYYDhtWeErAGm1Z2R3HWE4AHWGX5Ps4RMFoi+XZJ0K5NrJJb5B6Z58LqEHAO
D8Uh/4uMGLt0qg4BsoWlfs0ITZFX4O23AZmkkXybWPvtt2yRZ7ncbjrK+jTsPqPe
pxd7CCamLnBwRLcSn+CgUiLUwLIV1pPVSmGaco4TMNa1XCYCI351jG5SO1cQFSci
hN0AlAcZ9sV91PILPLH3cupwE+VN9KWQA4jQgMAPwD+lDOejlHn0a1Ru19Z2yMD6
6TANxiQ/4wfseunOCxO1kVtu3vhoIeRcNFotzj8bSBMJE/Q2Eyyeynt818jUbaLZ
0balxB4Kg68IBUPMzPev2cfiApE3Rqnk5JjKozawjhsWMTgvjzBDZ7gfc8baL+i6
xnmeX2ZEjLr2XYG/akAZ9UufD5iGYxeRi8haFO46lb9y/wJG9Lvh2CAvMlRsuIS8
g/CPozSQws3bQ6Et2Uz6cPmRJjimGG3Po1F2dSCeT9G5RNk5C1OoQXqQUjmPh8M2
nGXcbSb9WrMsJRDCLQ8XCO/s5NPeht/2c5cYTN4dt8+gxAaAPlOVOnMBYeXofA7G
klQGiK8MQMzN8JgUQE0j2Os5UKM4uTpG5cnrqYqn0emjtMArTSfrWRNQ3KGYY7f2
OeWCgl8Q2WmqmuNczCiX/ifnq/faxC4KZzam9qZWkwKD37aq1IhDJZnLN3TQXNM/
uzsdjGjByVtvA3xyTc+6UnrTWpx+y+4WDCaQ9DdbeReGWjpCio10lEjfHVdciLRf
E45OVW8F0UKpDYsRtCv1U2sA5nZ06/Egj6AE8/x3BX3oSA0cH4aLuGP9EbOZqcNf
PbZSabW328Hr5+/jQfySTx/Vk7Or0BcjIPgd8N6WAtyxdpw/JoLN/EkX6GgmTY62
pzcwJYoikHGdvdbvupNsk9nGCl8f1te7fmd2YPhbHXp+ehBNJzSjtmODOXnqC96E
+ALg9FvMNITUwpXMpsyNPlGP6IENIRSnK0N6+4pfe9XANcnsDUV0USwyl6MxpJY8
tiC0kGI2XsXw27C6+jb/cVN3FPj6p11ZuZSvx/M63C9dJZTNpvGw9VWVzuH7H8aO
SpuQZlmsHT5lzcfSdJKB52TVh79vsEXPV1qDbOeXJXaHyB+XMzapvcCzYRGnKXV9
zVxrdzqo5Y6o6onxLp9ggqm2sx1HsTDbqIUgAy5QTKL780setIL2aN61mpJ1s0YB
4M/XbepLD40RSI3AmsJu0tRAs4KaUIYo9UCBu3tteNHtRXea1+PzMlfCVHzCr4Az
kUZRi3Ylws6cMMx7IzR8JYhPD3ZAAqmJ/PKt5G63v8u9cyRb1XegMbYGpeMpyvRd
HA7P/Xmd8p8NbxPOcwZiMbTc4Xep58xK3duvIGDXffbTwY/XbfrCzhmN1Yinvqya
MhaAWUb6HYY6wwCKDzIUojj5ijDrcOBq61DmRHXgO5ywj5XVpSP64i1oSzybckMv
WA1LiNuC3FGUKzp8ZWswUFhMzmzEv7JZfpwG+B6UkfSSpmqHqZPxZf6pJazXVBTM
mUVdAX2KqKOVPmBcTCUrK8xc5gOf/S6TbO0tWnoX8J+43wWCqWwFJX7nnmsu7q7E
mNA5IiGqg5PpmvOL+InFFKdMBR7VnkyB/xGgqfetvLCg9jX/mD0rNZzCqTA/BlAt
e+X2gaQgz6xHy70TmR7n1RVBEM13IsbYreJP494O/cGD5N6CcM4nIRTQJyRtS1r1
ikRH1S49GsdZ28I/1oKFa7GFLVqt7uUhzi6EvDv+MDBYcrOQJrFdkDhbH46WFDQw
qV4Bqv18AtrZj0Rt2p94iE0GwI5MXE+Mk28MgOHL/Mk5TQ0lIhJryUOmfbClqtsL
fgGjiPZ3Ktl9lEXS+ymrl3q9L2Aw6BrodRsPJVMxcAcZtgslYNuXVWh3CuPu9Khd
hdCnDJ7nJCBO9KX0EvAON6dTCGRLd2+laxhIHpNSNUZ1+mUm6XI2/9o9Tf+u7HsN
0GJs79+fG39G7fD8AIedq4e7CX7WB6gm5B1AKvBvVpdYAzcQoKFHByvnWEqPJYGY
QhkEkwixk4yxPmwO9cbapznEGtCvRwR4sZY0JOiyTZ3ZdmEvRadh2yPMfJUWrjCl
Emvjs6pMYsFA2PO3mhBJTiWc9n5oMU8C248d0ZYxT5XBsVYr1DXKF8JeBGmg4Phr
UQ6S7dvTOLnStzpMtE1gcjJbS+RPHjLaPeHETnxx+vnqYxtUMqOHecjsHKAKVmdA
kEZNpec2WLu7rvzghkAK+xD90HxiBYxMobnWHORwRzTRF+1vQa4NACUlkBCBdh0J
K/6Ihc1DPCUbX2VcMX3TvxKBga8QsbFk6mbMM2BfSjw7Wy/BdmQ+D7Dq7f8qBZdg
6ZgsUz69Iev4bYhrZfXOOVHjwVWCpEt5j1iBouW/SCpyem3cXgJ5l0TJ/ACsyqZC
dUslQtsmf+n+4HIY3EeMH/C8fv6zCVBT5D3/61bHx/qKIdL1+BSQbAXbOMdShWk0
kPEN53FeAFlV71J+f8+fMFb6RGiU4q0BqmXa7P+obpx2X6rV1OSFGPBXs4Ea2CUC
H0st6EkfqADJOTVb4wJ+Zj2DCaDhrfN6KewFNScyFRWhIA4KB/9nAAWY+it7kEys
/2XVz6xQTfZ8H/zYglAKMnFr5EEPVlyDgx4NSXnqRnIrV5pQDvqv2ufW9WUH4ou3
ZooSmeucI6K47vV/vGuWYf+AtG70PjK8B+Pj1Ou8yfe0O8aI534eih5mQfODuOFo
Tr2oHiIWL0v0b00s/4cvJAWfEImH1e6QQL/GM1t3GnxZ1hJrnx0qXqNYvbOqtLbN
h3JDyyRdzdRPHBcoXtkdbbLNCf41n3qG4nLCefKwTaBdjLD4DI82QFbNghbwOgjc
UNUi2sj71gFueWz4zSnFVpWjvQdVj+9PKWKj6LlYtk5jgwcb6byke6xQWeQpCjAC
EwiSbZ3e1mHB9YvVHYHKGgch8xDW5aBM69M6J9zG6FFkgETHloQDSrDYosmZM0f8
fSqzOw9tsy8wJEc725jyKlHd+q8kcXDGzKuR1JlT0K8p5sgEXljNSLGP97ZruNtr
0V+VDzzJ/gggGFNQKnm/T5E+H2Uk6QtLQxvpFc3z7vxO/Kbb73EXgJtYLA54uYjm
/0VubSf3ft6FYX6JwJ7+IIhshTfEtw7vgkuiQdbhhgvPRwd+LTnEMjLxZfHJlgQa
CgBEgtxi/kmNqXer+bovXj1GeO7pOLWGmkGgK4+PW70mCF+pLdabvfHNdiWKhghc
fH1Aos9E83m/JtYE/DZDk6MDSHn4exCiir/xeM1m0TJoD35W9B6A6VYO126xDLhI
UrAG1ermYcRsmsR6vwrmYCdxlckDLGau5/0qC+EW70fFLlE1rml2kwlxpp8F+Wnm
dLNmanssX9gxnN3i9nTXCnqfuTbr+vxfMLL6yZ3tXWFQUR/IHHYAK7O7eAu/cXEj
YFFAV+Sj45gkXZLGBvwiCo85K6gwur6i0hXcGFuZVo+NXXMWcdueMmaaxsNZoHpp
1L3bIIRw4RjAHDc92VlBQgT/qGvj7S6MDjoWIE4kUSQScQjPTQZZY1KjwEvHTQlU
LT+WUbcvgy2zhq7cNl9PTm4UEtAWoasiNv+MiOLq9yra5m3nedVlTBLmU6f5kt21
6Fbzztx8Y+2VomM4EyeNlTvC3yhMpBgKrvYxzR+VujofQFvnBhQKR7/gkzVPOZS4
j14bXa1M1KU5kD20TKABWtFo4gloaNl8uK+0ACss2JNB8MCdMjaNkz1uLs6AE0Uj
jF1yQr+4iJ11J5pHrisEubl58POL7XCYhIk7F9hWNuyGHEtddQ+ZpP0z8/0ms+CZ
/lj6C7LVXejNTIwkHyxAlXgvjzkq6u0CVTbgZJPa39/pW2SgF2v8kedrpNQ3q1d4
ejU/xR0GHzAkf8yxneAagsLKRCKmj89wLsbKcvj3MJIlYwUWJZYlKEWX8HGcU51K
2UUd6fk6ZM12EALhPz/mH84UMy+cYGZABfZymPlAcWa6/c9kWXixShmYQReKttDd
oohKnCsvLBABQ2iSoz7UPrHqakevBSBlYL8FRG+4DhC2/DhAhsGfgd16p3UY2Utw
vUELNOoeJ9+Qu/4/pJ1OTt58s3FrPaFNnRvXHwxMJGHO9g/fkgD33iaHL3E31Ofw
p/7VKVxjVqpi0cn+yMtN51xIyxA4uovx/c+Cx6fOHjTrwyeS1Qsey1Ajl+Eif8RI
J3OhvMWqPfnU/v0DMFWtapxfYpm43pq8wbsNZUeQSTWiUhL3LVmRWhnfkkci9w49
NgqSolH4xNrOazlEIk8JH9jTfUYhJD99t3V0RRPJDtKvx5sZllZ5pD6LrAlC9cB1
i9FbV55XkDSqLa+xK/4R1EKMpELaU2WwWFD4tUHRZfg7vOBagWSUivxPPRZRhujW
/hMGKzNL/sTz0YoGdp2yVUC/faEYjwvqD2/OwDywPVyZ/OE5GZsG/kxwvHMxCRgT
ecetcCAeJJIe6ra71PtkGmz/QfclIo82jDagSWvIlsjA6/T+NbGkNe/Eb+e0nM+w
hKQGYGq8CZWdRtXimMjF5SOR/ZGuqcFe8VcvplMEk0QXmB4ElFnkumh2CFsiGbp5
ntm90T7noi3Z/HinNtNkS7oAOlCdAPFYH89IY0/GudczR691RkejfbIUUUu8Njq0
NOcLwdFhlckDsizlxyNXXr6MNSmJTnIJKqtEB22fhc/LBledT26GPud7cjChClN6
BlGRRhTV9N+6EKtoezXOPRsYUadHq9MEmoPIBXCOa7GpNpFFw/ZaQ+H251z9400g
JI3RFHI7XCnNZEfVzogCO+489rbDb65UfD4HT0pWl2vmjyj8W00u56ES4ARdAQb6
z8j05kkSyoTg8pYxk2FN6VhG2zfv16QeHp0GyYWEG/dCIV8FxPOtK9/GXnHYfw0O
AhC8YyNAGEVJyYff5VLNWk7Rgro4uU+EkO6Xf91Q2sGRr4tr+zWNM+YvNjJXxyJy
j8r6Pd4CwIEs/tysDhQyHmIz0IVn35MAjbVf5YPyO4JD8Qtz4MGMEQ+IdQACmyAq
O5qdukuJlgyFDKrVDgy9Q9w7/dvQjVRIOpCAHFzlYy8IP2mGXfxHkvtOLNjnVgKj
v0wIioT6Bn8E+ZFGvDit+Z4vAUDWieYB+Z/6JTky8/dbWMtw+bZxLcHPYPTCbcHu
pdojKuc4cg2HfAEqGd3RsGzdz723UTouJqxKLeqrDpObU0GI2gq2sn73BdWbVXmL
vzSV66cXJsmPEpJT2oC/Y6YqHQh3SgJKQyxTtILdD9lfrvMHEjYRXAbeHeaVv3MB
roHlHII+2/8BypN5RmBSrsJ9Bf+VlyY/r0oUZbShBTFmIPNJ4oCl8ZTpBq3XeUen
vCDTS2hlm5sRmwzugLYeXYk4lZTVF5i08IL8j2j2QJW97hNdTEl2i84y6LP7RyWx
U5AbGTFSodz23Hc6kI7bhB2NZk2opyzWGNUryHfU5lc3duOkAtKKsor/6XvPUJ9l
PwyF+JeIw/oOJ2jpH5EdZZuCjlweYBbKx1/vopUXhF9NpID2vaOOnpOeIdzHS7Nb
wFKXkjEejrRovnCzrnt5FvRPtxG/AXB2U9POALVcBC6cis2qjCJrQZjIYuGHPGov
DH6E7+MwplFVknVjGeT/DcJKiYA5nId/UFOzev4R1Z066I0+eR7GwVHdVaUXAeqR
/kRgPU/hVdNGPuhnBQbQRUe+UvVsbGVqqqlm1Do4J8ybdRRcSW1vibAFNLw2UExg
w1slmzbyMyb3rJvrx9RQZSjBPx8KFzEg1GDWzckbiICVMBhdFy6npdVFRr/VMlbu
kjGX2SbP2cqz3/t7iNcr3YwFw+GDrF45iAI/DIQuv9/mmRdeqWzq4GhWT3N5vS+q
ZhAKhd5nzAfRFXBHvhgmNFI3K8eP8p90s/F0JU7oy8N5UW3Vym/07POqa3KYbA8/
nt4SvIWVy25z6GdWaeSQZoINsohWV0EjiIocHLN2e3UbksjeuDlvGn7+v7zRdnNz
LXNN3xGUHC6lRRZAtai9rLLz45+/xyfqs8Te6sDcFeYbaL5XKtoBFWlkPMgXC3ul
835hc8YYFVg1U+wXPyOYL653B+sCYAdk3QEHQ0u8Z3fuoaOyCvEzaoJF06BW1B2L
o7/kGGEiFUglf91XRZBNwS/BPiMhXIJKLNHT9B55epA5YlJk5TK5VnEnSmBIFDE3
vJJYsmOUcqoL2NS5+619JuvnpnxQNCWWoJQtECDxwjJkqGedFKHkjkU+DSnB5O09
gHM4EPtbMos2jLkenFGL2+Z3gN5UB0eZHIVZoaxon3FyAA8ogL9iqy0BPI+bkBo0
2tsK2TwOprazedH4FIN5zZJ0EvRoEOLJbeFiQFpa0OuGybKSJreQ1GrrOWoU/EWQ
j5Uh3bqpdC0DCsQ9LfN4ljDJI5vkqJzjc5jExn9YqALxL4JeHnZdbPgU67dbOLX5
Evxm5EKn51/JjUiXcRQzEfava0pgNPgruNlYxnvDh1cMQrpB0d8tmvHo6eY2dpSw
6v6qsNhOW+POxx4gNzbnD2T1V5HxEY33j0nKxyTwflawVdxJgro3W63BNfva6CPa
Iolh/An3M65VZgAZz7aSbN7Vt6klwkWwgYAAnXZMPyrE3842O+HExP7gCCEpYCqE
1dVWl8QCNuR14hbQcD0oKXeHbAFnC8bmPs8IfIlXI2chd9HM8fsTF2jcedbFEETD
Ew3dFLMnNQlY4W6xIZEr/2KNTJtBO9UeYJSwCw5UtoWL524iRsUs+UrSXfOPt2z7
Q4Bd9YhoqlhoQGfbRAKR693WmDuJp4ZZzZ+20/XfCH1yKe2IQXG+vwaww53CsYhk
q8VmNlV/OheHp6ckis5S3qbVdwmBKmcchn1sECftNkf8mdnLglJtJXaEzx4aOC4Y
kRVAXKtyPYW8knsDnokGKh6hEAZUbNQ88VSZiP98ztE5NNn7qUCSVVyMt/yEiPIo
wqmIm0UiI3eTIYBlsJUmpwUEUkz8oxoVLiwyNu1CsmZaLO2rCp851yLlQyEHriy+
MjEfzo0APUSEIe9lf9s9vAcIgWuWYqtg+jesoBUOXVIp16ukAPRe4yIYRQM87qFh
OyV2TKiWlhW+J0yVYGosyQ8j/irvXguGKijp6hEg6nAwUndN37OT0dto445nV93R
ILNw1YqH0Z8BQxcL+Ic3h7xrLVc9vLCXaJg4FiRa+de8Py/LlF3jRdMmB9MQ9Aso
u+QFD9rIpjC9WAeaBAkzOL8Sr0HggLo7hVLmhVdIki3oZOQmdgo+uHDTcYHGl+pc
Fk1LCj8UTuA9cpRSjtHRMJbHbWfM3ZOAkHtBE9hBNl8ifNLoeyjnIH6XNIGeWVjJ
QO+BoxTpY3OzGDA0YrIo2IQvUxxGSM5Plz9ilPcVFjdZpRNA9WLXqN5Qz70FFe5f
U0TyeCQ8aOdoqO8WhS1j7Lpv+YwL3sEARM/UrlihFvq/sovvJgpfMQGwDhr8JimP
6PFS1D9S+qBI7OoreJN0cuvwN2BPA5AG8PLS3KIqHJObx3/A3pi+3AmDwcx9e/iS
8XKJuL1uD0PQZYtk3IIyZIE1lMehdMYZhHEPGRlTSAK8Upr9XfVNteKQeMwUKJYI
evHOLIuvAVync5jAEDEuB7ZAYFcye/LhhKol5fBOJau/ht7A67bFid1Pzi4gs5QC
OqBw8CtusokNa+BsdDiIw5/kq4833qm6AeO0MdFVe77la3S1oqw84EW5l4o/CSoE
vbJON10C6smK1/Jx6tDi3dQzkCDxsDoaC1mAD4PpgBTRN53Nh31bJH7w5P2wTG4f
U6TFyU5UGLmvmo2PqdKOR/rCuK2NQ4/h9CmTzlRwEUhl0CNGJP8FlIDNeMw9x7DW
khYFoaJnc+mA99AeaZ57XK2mSzW98/SH+OAsEe5cQyIHyV6Ql7ytCqQE/vpfm+Uf
l4InulaDglnrLIMOUe0avRlmP8UFDpTjrktlCLXVTHhmZgLfhzy7qc/PZaezG+ej
cfhWkeEOsghWaNLhKwY9fGQ2RzqZ4EODv0v3Hk1nqxGtC+GA/40MPlKoyOAEMgO5
pi36ibn1oFZ7xdLg2PHda+ecdbqjyS8SEabuj9d4eSmONuH/qdmdIiCrzQfuvyCt
bLd9vhHVA+Uhf2QwzkyJxikN1QqwApLTAcz3ZFwDghGDyNOdFrIun8yOMJc7U3zg
pUbWavhYzTcQ7xZbJvIQbB1tUFShL6f+8OdBMyUO0Pg+kIqu+rg6VhOPfkMdehgJ
o2Nt1Z7ThVPdgj4LrxVRtmcts0cb+T3iIJCdUL6CDsMv+GNEyexACU1Zmt4o2GRB
ml5riP27IOt5x74BccjGAXWyRIy8YSru72rmTeOHjEOn48MWLUTN+WTcH95sp22T
2RAI8xMRAjZV2xxzabqAhGihXic7AVLHq5MjD4kqYQJIu5FIpxGW+NLM71zikcLi
CQ5CzunfiOUoqeLyawYDVgq3mAPfWZX/L/mDQ8cRhmjIk76XczEfA1E9KGmSC4q/
qJn/hLOA8zXjBfXiR90AC8wFRSFV2wKBsuPY90aoqrZqucY94zxPWps8IEZBzuC1
6dEtBXiSovs5774gftNzca6zVMrQYvMFPfitV56hX7pK5tIqSgMRnJWh9WTEY7jQ
pH7tU0xAksU58Aa1yMozGy32rQRBWrBpqlq1RCIeiod7WetqbIl/uuSFe4Wgt1ak
+KIZzyAk0B1/WJxRqGDPRxbVlmhWUq+7vmq3NX2ncvchZAIP4oStZgrf8nbwt6hf
eo8Z3P3abCRoIfeXBbjq9aouV5cIrsbpd39H087q0LTEtm6VXpRQsXQV7fO5KGNk
wlHJM2C5laAFR2r45FZ+RWttQXGva0V3tAcDdnufWwmcvDpRu4PdxdlrpoLBm+Z7
/17ffvu6oL08Lu6sLfuAVciP7IamYttw8do3cwNrEW1sPrU14IJyiC8w8YPn6QQa
f0v/bYReeXMmQsYM4CzbRZ5Liyg7Ds0PIdno/qOGaezcVvi6RclzOyKd05IK1TGa
g6lTsFoJwHDXGDYm2gnkTI9989YmCIKpI/8pYp3j59QGkHv69ZSpAwRSz9zfJcHV
Ip7V7x9S1jeDifQXiFpPzZf99+QHa8nLkRB+XqVp/y8H3bOBngdgjtSTvAVz0lTP
1ojgPibDPaVyqi+S0rW2tn3PbOn7aw6B03M9W17LkHYXmWjwJv9KxlnvZoCv9Bbo
9nbz90LhMkOyRFcuyTo9YhrLsKNO7tMdC7vehDAuSM7aWmD4eNxfN8sMxMpDs3dk
PpwyFe3jVkDSuGQrzx3I5RfQr6uHStL+dPv5XNzqORzVylndkuBF+oHv/FbIIYFW
1W3qzHmoVl3A/ULnbX5LTJwjcTLLZojFVPvAsAR/Tq50DxHpmZ3hAboyjUdhQEr/
GXpCkRjTOHNTsXHOlhyl8UV4G1m+5VMwcwaO2JeqreqDwgR9jEqz4iQecswuLsHe
tyNgTfV0wQ0q4KnWlsaryzixo3k3iYRIEefiUdSeW9yRRHy2dKu1YZs2UOHbCy2w
k1/cEVNBFP7tUNjoTQBfcX2W45q07qSkG2RUa1zN3MBQ6W34GjnNMEcuOp9T7NuD
NGgI4x7GwTTnnwUfvJO/oPgFi8ud3bLZYxJ/4fy43wemiYFOEla64xRjVyMWZk/a
aJ2bQ6vpc0K9fCUbb2/XCuU0Yn+ay6MgYZ34PeWelBZrB/fDJ05cj8OHuSwZBQJY
wiI4alU2Ra2/3yopPMXcKCG/BSvHxl9N58xRSBppBjGgraVfq1/zxNUDp4+Hg5Eq
Ty/9D08HD5Aj3oF2wrKoncplWR8lCA74d/QMWzsf0XdQRRz5kaiFe6tXA+naslyP
iSAEm+QM/h8/rxrOywyxKCPoWu4u3gD2hkeAgXhZEojrhTL+vU/Ns9KD8AOqypP8
2bFemcoFuAq/q0NTywdQoREFDoOvpHRzlYLtfjAxm6I/oZ3qbJZTPHCnDhXJePBz
oBV0xQdXKeKlceAR/smfqe06/ZHqqHQXNRT2P2yEVGVgxsZxvb+wlK7N5+M07/+U
/9XQy8mLUIjS8I+rnikTcHx9nQUMdfzb7uj1AEoJBNKa0FcEVcXh0DgiXMFrqfIH
h3rLaIZoKYchPHd6rG4PnMPjm2Yb7chLl0bLzYukppPZLmwM59n3k3CgMXHqOakp
tYkj12fKVIFo+n2relR12C47CbgkOAlbFNHeiaxZbCd1xT6dSH9C5fzd9ByH41J1
uV9Hw63JoBeQ+gbIwA893VCqRbAzJp2ghqmsCA6AKqsvkx0yvAjnOdU2KqVKUWue
gMLD2TP1ED5yYKinSQI4m47Chsn8i5j7Nz9mlhKDPl+knXBnYQe/xhGQOfxBtUJH
Fl+/rfPThlFMz/lB7IE4X9NmX7SvySvOiSCfgpuNhx/e5FAG7v204oVhu4sctvB6
sEmex4Y47jVU3KOZZ40Qxm8Fz6O6udq4rWno7Eg9+OYwWey2WGTOiMyEwpDHQaCl
7IaHiwZtDd7fBVcvFM+q0oZ1hWPmQcxzZMCpxcQ7ZXmGj8JPyAIn4q5crWyIWShl
PjFi+OKWnySAW2LOTqNIkCiVXQhgM++fX50mi2uQ4+2wsvFQU/Et7CO075aMyMbS
BVDS+Jj15/OLdRDiezQcZv3QBbXOwKpYcVCugsU9EronjUNYzNP1ymkujDSBw4Kn
1Fnpor4+tKj0U8E1/yKihm2xtk/RSOvLokCawFx7rJvxJKLBbCYspcutunTxC+He
0GOWqHj5EiL3Nh7Bhj2r4zq+W8++M8HA92rXHzJmVDiYXNMWhe/D9hsy2UulEAcM
EMv1y89q3Q9MkkRqsOtSrCfDtGu6Evu8pk/45aaDdwvpLyQPKnB3ynRQPu3I739K
JEHlXvFkWRvm6o205xtnQO4y11xyiyzkDZganUiyZDde3W9xeSOZIxiODf4h47Ua
CFlx7/7Izhqs0+9twy0QFwmEpP4i9CfznAHACESThs1gKo8Z2jJuu1kaiya08FVS
+2m8JTfFzOm+lC+8uqYYm/SPPjBftE6qH05vzhsF7ZVf1Z7N0RmVgw7ubTBwpLG3
Hc5GqrqZxJYwfKUiEE/OPL9aM+zAlJabBBXLNcCC/zm2iOOOwXnBjkk8BX+k7uC7
b2hpbk9OsOEQT23iP0Gnx7Q8EUauyoq9dNOz7HSXjtfwKWl6zuCQQa+a9O7SMmGY
8/yUjQBqM230d+1hfmo5mKLE0DxWsilfbkVt9ndRk+cT/SvErVPtrnZ78EmvKsNR
AXQll97AQtOPnrRiWE2TUve8x9e/4jpj/dnktntMX5FJY9feni9BdmIxqBuMsc9/
5gUWNXIyaeauM6VJRBB0mokHDEZy8/uwe7PvyYa2txfE/B38npCu1rMo70b5EFvH
APHR7ufXUXz1PX26Qh6MFAXdk/yLKEasWq8PWKhIIinRiR0xzg4yQHvnMBFdgKgT
NeVxdGj7cCtp2cF9Kj7Jf0+SIK8ZM0mf/P6tdi9ho8tKTbBM7pFL5Z9P74SWS+zl
LSigzGoR90WftHyc2VkKr9+9HNolCY5wsoEOLYZO0djSnqpSCwSxt5hOd9Duv5iT
97buTFTMQHo2Q9MMylgdj6vpmPv1adhIpScVzNxrqcEtOcAZipTUxx+w+ZL8Jnrk
+C4yiicpnQyaci9FIVjp1Oggx5zNRyTPM/jXNiz4GZtWVRVGNw/i5qOimvX5IhJC
lDz9c56njWa+qyiEE+X3kEpJVvS+IHQIo+oKhz8+uhduSY4AlX7OqeqR4bZzsX+Y
rDxgoFx6wnf1yA5bZJJLV9Y9d7G5Evnm2ECMfO+OaUZl+sshA3DnhVGSJ1GnMEbW
UfcoexqQDmSAD0olYw891NMVIjbran9fxggIs0NTc9wtnF6siFeJyVlBYfVf3Vof
akGv52eaRdOwZsEFfqeyWI30s3wIhhAZD1lAVRrgYv0pEP5SkWjsUUHfBFK2lHxT
TcZ4skizrPt+12Hrc4sLEx8zAGbMVxd8i2/P6lp9baR7KjQl8F/B2RtIwEZwvXlJ
X8IpH6RsBj+e3VKz/kViB2Fr3UsoUVga/BuBDPXhYjbPPvXCk5kUgN29F4/v5yTL
aCOUSA0jl2MGvS1+TGxWBMf+CXwiPGm7pyDhxcHc4sbr6x3K3XHRzd1Uv/oT6vr5
suTRZ9kYyeo2bGlJQZ0oUqP6tVUoKR/AkLYsMD5P2/BpbA16Z8Qjn3dcQqz9ywIO
FbxeUmsPbPR1NOcgK2dACC7MdDwpQpb5SQJwgyIv0j1gF0QQ/fekUhVItnR8dAQB
5fkLi5/VdO2lK/74ISJyUt0ckgCcnvrzZOfuZiSjq/VW/Nj0L3GMD8a1ItMdRvxe
7NYwPfuJ/iam+8khj8JDYKp/lOBNJufx0MrTZQpse7hNHq3dk0OC5PYHWIDna5g1
6rUk/0kuhv4FOfqK9zcqE+ovy+tEgHGbz9cJdPAa1CD2pOiMqSyT7r6OgicL8Td6
XsaU8Y5uy0FRyaDgdpSuQExcAif0kKDppiRJik2fY0q/ShBO1T5AjD/aPH0ayNca
NECLw3cGHyTv9i/X+/jQbGlb6/9OKzW3TfsM8HChj/CrVVITa9f3MD6bGvea6qWs
xWPM2A4ecVmPQ63Ro3N9PnlX/l17SeeKAe05Rluv6YjicvXXrIm4nqJGNW/e//pg
m0jGxovcExCg4dxhTO6Q2ZDoCc2NKdff3qvy5EeOPHsXsUK9EKsDgpn5beyllexw
DJmLjfBdDd6FKqL4kvxnugSCjXhCNQ+MMAN4N4h+u8vWoXkcFrMgT+7cPbj48RDh
Kt1+aM78LtnzVF434WRUwoVc2U8KI6vuY98NjlRJH8hGY/Vov5KVdd3bIexxqgOx
u8Rgnd9+5bZSStoEgtNKgdp+FbpuhcGiYRs5UPpdkWDDKtrc9ticdQY6jVH1Lku1
5fsbDeOMZqTXVgwiAUhLz4XrdvFhccrZWEpKr7eZ0rbb8M7FjC8S7AMBWxNiumFR
lBoUYxVRoC28PycOLXPyAFNTeCypbvA8T6oFzQpYk5fp0OVdSnrtUdZqgJLCBUWJ
45nWUJqZDUel2EAzeJqmK7Zt1moKnQxikcOFEanCl8JLdCCBnZfh5/BxchfX6pAO
740YJq84l7nO7EJnjCs/pWrZ7aj5e8MvTffGNbu+1cTOGNjRMxd1GpSlqGc2HZea
ktWP1PJ1bPerlXiM4KSyyloZPtS5FaOMKb/P9E226CVCaLyw0C7VFcyP23XIVyWv
JL2NQ46MF0dGylEDe24lI0ggQ7N4t0UDHW70QAbIwA8SyxHDPXkOdiaufeyI50O2
Zz+2hF0MEtM1rjhjoQOQ874XG3p054LXH929la07dNsI7dauSrzTW5u5wGandPy1
BPgCgqIO4Z/oblNZJOrrxpnP3I8d917O5eXiXENNMnBSFu6mrNFHZZMWjT9GCCJd
AtGe9BbO8icHlsfpoXNRsmqCRqreZu7yAHUc6ZnaCKMcESexJzzzvGbCbr04Wfts
PoaSt2sE+EsIwZOEfiecK1seaCmhgn05XEM+sWywz6YrO0tppRzROofl0An7cD4o
biwPLMaHTij+MOqgso3Poh7WIHvaoJhFywkryhKcDKJIRB+0sKbMduPbtvZ530wP
orfFdntI2y4eua9I3SXF5POhcOqUdn93FSGq2teWpRTSqgXBKPG1EPs8m2I+75WQ
svsdeHQzS0AOYFrh0LYGBv1PTYWzAbD9H6SuE4Rmlj1zP5rNKAAfgONJnYwQZk5V
cVwzJMZWupWBCmQEVWkdyasnLBleuT7Jn8JfbkknIX2mXITqhiDJvWN2yUEOFL1+
nl13V4ksjO43E5aMvhF1eg8GD3obT8em80W6A+N/fyizMF0RWKGCLJMSZAaQu+TQ
ki9ssch3R/tlBZIJInj87T67gqPYXXtDHxKv3NV4qO6C2S7u5+NwdIB+H7EBNDlM
o+qBU5R7PVYRTIfI9CZcIUcEnflLoWxGqf/HmF5qKxPMffSFqjxp8tPHrJGMDhJg
v3GCLczCUzL1RWIdUp/OiuWC13TgPz+mdRgn/w9NhxHoIL6OIZLOicXEzsU60rtE
9aDoN9yJiywVobtu9tZb4wgaZVMPGYxDwDLCf1HZoUmZ9futAUCfvzwgPIZ7rPE3
QAnaOWhHKNGyWzT/SRq4e2zs/Csqq2EHmU6iq5JDenqQTkynyAemD/AnGC+c1BlG
AC4zw1dF5Z1VuO52Js6o+SSMbYkjDBwu2rtGYVgnijcv1HtLI08NNE82ZP55+7Uy
OdaXxjFDn2SjaDxQSFhIhb/P30/ntkL5FCB4YKrQjvVssNsVkwI+Y2ahNb04isiZ
eyjYj0g4s3AzYmFjw/rb3Hex5sWEyC8LOjORwZvEy1NAc/wiE+/c0A0gf/TvBAEg
zzITh8J9jXhSb69pzziYdL8zg5+/WZjSvDrGmxtwB9J1IDA8y+Z+kd/VHEIc7Z2r
ilDiygMC1DyivncBFuKgWsVUM/y9O8OYaClf6EioRwhm6/uv+4sjWYhY+0DrBs9E
RxcLcptwzdfYGBSrpgsNbCCkY9FLuNIypQKv8onfiP8eLfobMqeVYKpejirNH1xe
4vGTKUH4jc4COLjsDSqCw9L6OkTqXRgM9J255ZKAM51YXoCsScfCIu7I40r8JGzI
+hp9734Xsli7IoYcoEqtd4MQx9ZJ2UJGRKpFJ8n7mR2fDPAlmF4V2KA8FSjgwIg5
ZV7izvsnGudUy8/Drh3pEBYmSHs3x+uxA2cTvbMorzXUirFSsnw2pwZAk1W79QE1
osGFeFA7jU+xT2eW2EncOvxe0fSbXdT0WVJ8Kcoipc15H5ArVxOis4enM5f4/lIw
fzpL9itP2xteoXSaUHZ1YfNPno2jsPPrH420Y254eZPWjzPMGZK5z+isk949O1Ki
1uX2DTrCahi4Iyjpm6Cg88oryY7wVgSoNa25xZvsggKZbW1Mk4QWZpxmS/y80KfY
F1fYBCeM/vGvkfCIbel+0UZP6PJCplMJ8v9VvXEhMbfnZOyN/GnpmbXzidKGg4bC
x29CECiDQQKUAGKkCoo35d600Y5uyEvJS4JP/ywj0CyEVnZadxSk4RAyLUfO3Z05
d2T/RMEggnx3Hj2rRVcmyQPIosIl8Vc3/BZBoFVQUQ7xGfKMYeM5h431DVjr99z7
ecCM1YbsJMWkRkKr3HcKRXVFALOzO8dZofarN2VJvUvsm7Wd+ypb7FwYFSOkbulV
wsYkKxDxPoql0PL9rVDuAkBdkFZEmnsGlsoXOlGQD0E1a311Yk29sBtGD74wn8Iu
8k5AfJ2gRWfyG5ApD/B7oC97UCMB3c9DfM7XRBocqQtLQ7gp+pld9fJ9JXfxUh5p
PK4v7ul9QqTFKzJ+66239X3bCTcdZxNp96OxCvLOvWgZOHtfoZbojhK3G3E4toDM
Mk0TOGoMeTYNG+rQ9Y7beR5mcJC92CnxpU0sKA6l+ek+nEx6bIj6rkCxGIDF4VFz
My/2bs87eybA/qLc78E8K1OwVnm7jRaHkdfVP8wKklC1/FOsFUnRh8OZAsE1TXoV
CumNY25o8wXedOIoS+QcIwWc9B0eh0o6yDdk+M0UWJMVeov0lWloJAfLPt857D3Y
ffwuau/hRi6OV9CUZp7hbT5HgmHfJaE5kr86PcuL7Tp6ktwTEi5x/STA6fDbSg8i
Rwjsax8IJeDHu4bL1ukkxmK2HqcIK4DR6tK0GQumeVrFgKXYQkJtGI0M9ferakwK
cZ4SNOujnG5Ejy2ad5eMPo4/lu1DVqS7donXSiAuxQfBl8UR+aeBJhXytzgONF6T
M8NTn0h9dowjwp26X35pXHsZ07xTzNx9zvBlBF4qZx9pvfh2gleeGC03Fa7ETeRb
x1NOWfMVtpOLBnWLrscCKMr4sU3NO9tPsGv5Gpgmw6jafEAHRioYafIIo+umpYOi
NRpd/WNo1doVmqR5iLeoQXmsQXRHho4Zr7YhUr6lgqwd5WPRiPseRBRHZryFGFnc
px+zNG/TgoXb36Qrguk2Oqj44ImA7vqKNJqZhhr67eWglLOuYqPlOSc15fCFH7Ik
ZGhhVgYFeTsY7lBf5f6iOYIMgEGwRCkh1GJDqywZ9zlhUPKc2UGjjQMZkeMxBIvL
HFPFoTVVucFlyLANLySl56FCd1hzLKI049G3aHqNWCIdKllCrhGoRBaCNOFvrjql
7SkEjZpanUeERNT2V6Zo5FP4IrAEh4UcfKYyenkQcz26bowQG9taTyLf9dfYv7NI
ObBKDVD1mLd92k9XKy/WzNIsaKPpW9G7CmSZW6eAIXFHDmDxtDo8XLPN1SwP5G25
qHsNrP7mbiUvjykfEne1EZzoif25FApcJH0au6U5e/5ygBPBILV9gtKSxZbcBPnN
l61mD7dQgXrFZm0XxBfiTiXchGChBHs8qUhT82GH+FUMWJFsG9JFvZIr2YsMAQOz
snNohRw6nEhz7G9Kr9p0OlXoslMg2J1SIkxOgc+L/o0Qj9qFai83uSTZjXX/gDIk
o+KbuKiCjBOSra9Hzqa7EmSAYBdOVNQOo3QnATqWRNteGSW9VFEJsYCbg29Q8SxY
jBhDz1q8D8oSJ2ptiUd7DPiXJhhba993sgANf3mxEldKy6JQsfYrLGKlh6f4QhP6
EgPJtR+O2/iP4O96SOvNr/48v1MYAXHHltCrgfixTHV67i954s3brZz49+IzlRC7
Np3wmVCFP3eFEYDxi9RSpqfvHqbstHgTcmS1IynXsFEdg21Mx2U2qz/3wb/Xv+Uv
rdy29lCqmf7wr90J/ZQ33LObdtRl9AlFfrL93v07cYFJ5ED78lNty2TuIH8r/3rd
9E3jXg9fKHTB456TvDY5/N1mE6YvJ8+Dw10hMvOb0LuVQLl8x3Q44vWFNSDVAtHi
tokockO0TJq2OLP/U4H8LKZO241/XbS5K8YIJLZZtXCmLvflK/zpeMZcV6rEEi7+
s5aYr0y3lMstfKAv8NwU/9tFX2VStfhMgvJNbS/hgYhQLn2Fd+g7vloxWX6BFLVr
Y5lo72tXG+/AdJM+SX3VpdIJA2HwNvoGrhoN/YCARxsVedHayhWMCs5Pud6ThQZA
ydrMVSr+V6kKtgdr1xn+dr3KJemEr4IS28wK/c4PqCiiRmSMbDRCfrG/Xgpe6wiR
ygZrh8Bit+Aqdkdt6jG5Y2hWk+3fp0c4DeBMN48JI3Xz8fUmq2ZhAfneBL7Oyora
uqxEAWeH5GL55N5BCsXVuDfVnpRVFJ+71yELilyLHHM5PkQKXc4vms1Au7gJw5KZ
nxsJdyBe9pwKTeHbBHbLFz4dxmF6emP2mb286GC8lZHqtJWVMYeVFs6PkSDnVYXt
fSRzIBKxxOVS8jFIDQPNtQt5v/61nmaHaVuTbkiqrEERHV2Eg13vETS5O10XBJu6
trfqBjK5hlcH/yoytoEp/X+xU5xi/sVzDF49yhxaesegXv2BEb85Lc/BnSVRcH/y
zcfUpuUeIEAfb88Tvr0w3+BDFCFaEvZzoFxxVXRM+ccIkbPxE1bSiuEprao8SaiW
LN+vILpY346qSy0f6aZcrCx1+/I26XMQQX/taOxvi6VY+9RHPD15F4xQcU4baXc8
t2Sc8I/5RvBghn91j+0smV7FCJxeNCOou13dKajy14YBw396HcxO4Shtaej9iAzA
mRpWsr28YEHDcqurBfduWblraxv5fiWaNpylsTlcR/yBctRFb+5QJWacliB4FaY+
Wqgx3cRHh7BEOteknzMTUzxzKZQZ8QIqYmVwxP0F2AaqLsjU6cEh29XsLC9kVdi5
MOCzleF35UTZ+il4K0Y2HhqF0TUJb2I+COHZEkNSat4MnJY/2vjYsd/O1h1UDbay
DmPYJfrtSK43JoDIiiftz4J05FF0zHNBrSDisgu2Zeg9DpD4gwW7VcK9apOWNLrM
5EwPJzWZ6HzYzR1YHzfWC9QS+4qcKL0tTNUWvp7OnyeHwuFbNS/2v/g+Uko/Fa02
n1ZNJ82d6GFowXY75NLb/QprtaEDSmKlEYAcJDmckUiHu3RTkBiygDosPmpj5nMe
PS/BpdEX2lat1PBYe2pjjipfoaivH7qjZIzNR9PPMrBgpJoLIxUrBl8Q6CqRECqD
NjEryoWkptEqbCQIo/kya6oKyw34Uc9jMsjWKPtKuq4fV955hmy5hAz1cpQROMax
/btP/nwpBGVwkudOcoKyGPRAEa8IcahD9NPoXddmGD90RACQRz8+4nOUILXXRVaJ
rzYtlJIuU1GqByuki69INL1BJzaDKlPjXRg4VKCw2w4tsGeI4Is8LKGYnXjsJarV
ITv7FueYIaarlktOI+bsjpQUNsJQas9vtKtb7jBUhyMwk/sIg4rxW7fXCne2dlej
eep62yof7pCfhLIylHzs/yzS4eP9ZhyqQAbA5TbDAfmCNd/rmjlnprRaF8weoolJ
j4ogz7XW+uq/7gZB9+ELoBxSdyTGV7i2gd+AhxSxM97ZbhpPaAtSlNelcWhdwrGp
XET51SobHSa5VxgCIeq2L2JqAraqewQrW3+qU94cN700jkV+Pr3F9LFq2DKmP+3J
9jHP8yDJq1HxzKrRdrCuzRWjT9rWT+YBUyrcIm+GOEBpQhXkq2/WVJ7eHy+J90qz
TbCHQBDzWgH4jBNdY7VUotN1dmIvMS3HFY2c32/g3vUskqgTe5qEeLUuYnvXynEL
EanKHGUTe+oiEHFL8AaEMhmkAMEZxgtsYu3YBBWxJo3zLJKbN+r5Bxrk2Oulr0J1
Nxif9R09OedOavQJBg6bQtDDOMa95Yecwh0UJ6q9HUMK2NKGTBa1wM8d4pL9VjGz
VxnxGukdBGB74wIu6/NjZXdfYXlvr9CriFjxocZkfNDfAl23dQikbX2T7zKfjOCK
voyZw2a8VQiH9mwhY1ST80i7DTrLEuXW/JhBjwxdF0ljYnqUWfrRHuXjv8eZw2Fi
pGGyXKz17m8bkTAcng5r2L7p6L8YEDGwo6iWv+XQdQjljIHPUKuAuftIkbBzxex5
NkBBkgo9q2JAnou7bUWCzDwkeaO71OMYvLyBCeCph1r2ZUUBclEYldK+V7KT67iD
84H+rbSzvDY2PwMWPvSJYWRFdgX72oKBZVBGx+SF38eI+XdFohBqCWtrbfzP4c2r
ho/mFUS51TIYTzI2RWGeem313GkljYGn1eboTz+vsqQS/cjghOKR1OTFuEOEfGNT
Kn8j7ZeHGKy0VgCjCB2OadUh8WZlQQPNPwXEtjY/AqhjOjUFNn1xNem8wDJAooMs
16ksYXwlOh5cK95FuafRxN5EGraeaPcpw3BWO311K/CK4PthomM9i3kNLNeJLGwW
sVpUH+J1ggj5cW6PKqGIZ5i5BSkYlDLpst/5G3rQRTdKr//oybS9tk4xqUFVyX+P
7TsFdBiakDBHrM2rfsttBAc+UZ6OSZWCNSBR6rgOkea30LlVB8DbAV2U39//XGY7
ouAJRmigVun8YERHq/wbL1RP342R+unuz9gQ75eVAGiH8gw/FIMdsD6twN3LLtKX
lrLakhn9wVZNXFydu8840R2xy2ThPS6UjFt4QoSiE4Lnf8K6iuS5s2RsyukrrRgY
BPN3Zyen4rqlfN45ROH+qO2F20U958R2SWeLQu0V+w6Yr3cX/WY1x8hGHv/jNWiS
bBCvB7GEtfDTUxdS0wvfawGGM1im+wVMhtoRZn2yVu93IYQlEpqixZFSarWyq5hI
vhHlQHSJVjwgonE/ZHUQ2QtBPq5Bq9AY4TysFbv9ysGrm5w4jduHuWLg1lv+Ja3y
60BYj5SH77UG3ywmZ74uiNyi+8uAPpwXs4bdRLPJKzc5TJod4YYqsBSOtRehYc5+
jJMLudTCrE+P/zdwJmYOPq2ia+OeMwx2fTvIe2AEVGtjMGhhjsk+bgwBIgsGUI1d
wFDw5Ve8kFttqjEMzN9JL5W6Mb+6RMSmvMyPYFK6KJdbN9QCavq7dH6xDag1G+b3
LvXHipM2t8P0CYuL9qMPQJOWETX1DVBnVD7NSX6U/lYkL/L/RcPX40SmuLzBJQxT
dRx12G2BRoc9TVGXQxPO4i+RNj2HuOd8eUJqSR5mDbII9KhZxmrgvrdUS7RZ5D4P
8+s1SCRs4rxbSygYGLGs0g4buHvSt6ppBYcqzfs/LZImrzGCU8czBXf+t4tQSZgW
5jkJgKs0BhAJXymxMlOdwXsHMF8Nw2rVnV37aLtpba/qIdvQil1HxdSJCQChZ5GK
SGabwT1/ydfSPrT7qJzh9w2HNXAeCLJW95DR0c7Y5iEA9cYS3hWXdyfOQtuL2fP/
UNa0ovyE2oCQLbs5CfJcgj9LkZxipgIX7GE/GDneUVCru1ZXwWmr6mx/b0xkiYtR
q6zK+KH50icCQn6Qn9ugtp7UjOja1y3kFYbzd2c5ToHbFlbTXnFZ9ojF/2iSj3DQ
FxrVU1HTiZDDpzCaLV6/7CzSr3e9tj6QOtNh/EviFuCPwSnYMpqrxCRX+PrQ6pQW
SuyPEVT+/o6s2+W0f4ug9XiCE9HDfSPh1S4BTTfmnb0qmnX4lnxnC6Sd8g1OVJW3
9oqzmjBzpInZTHIPvlVObNL1kTGe366DEY/EPa2bcD3WJxz7nRODHk5mldP8hQDT
W3Qae0pMOgxHisAhquk4NtqVpU7tiuyW+/qufIRWMpFaC6hw3CjsHgpndwcYaYzd
hzMJFoKSNlj7KV9iwmtHcGyzlrOT1v9W4SvE9iQOzdc3yxXHJC/sMpKfeVqyBY3m
Fl+QBaGkctUolJQ+CoazAX4bDVK3G9I/15n64YdDY9w=
`pragma protect end_protected
