��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���9�{RԱ[ж�8�����������/a��:��#Շrb�,��Y�)n��M��Ӡ�5H�������w�� �Gx� �Vg~�r�5�t���5�Ш>@�t���57�s�f}U�������2'�k�l�E�g�ܒL�������(B`#�%��ǩ��b�y�ّ��o�ka�0��4�~u���͸c"�x���3_�XlB���J\f��E�W����	�]��8� HI{�s�zq ���s,=�G�:F�V����Y�e>�V4e�i��_�F`�mg�_}j��&���\���B�꼗5�%_����^��Q��q�o
|�zyFB	�9{i������ag�rʲ5Fe��Eó?T6��}��K����JN>Cgc��Ӛ�cH�`��(B�� �l��j�*���gjdų���\fٙG�%���$�����tXS)�N�����f�td���kt��*ؽ3��t�����-w��^XY���L��K@�Y<&��F���F7=��g���=�p41�z�Y~��%dh~��5���$/_,���\d���b�J�Jc�i)vs�L��]�U�Z4~,��7E,�~�<�bЄ��
c�B�(/��kЇ�6+���?'��X-%��,*Cd\�H�QJw��Y��)�>d*5Jy/�����֌��%�G(�^`��R0hL�U����v�A�k�3uNh��V�3SIK9�X2D+�����ٟ�`3ѝ�6&�
*��G�ӗBLc ��0n���m�:Ҵ|�Srv��?�Ь��P�[-�?��MW>!Oq�#�p�V�������Q��^�b�1M����+qlu�*�v�F�9� �h#�Z2�VMȜ�ܸ��>��������E1*�z�Z�J�����FǏ��*�w�[H>L͉@�܂��>Y�Ҫi�5!���3��]�HR=�BP��U��y�^	L�w@�J��t�>��%�̥���#[r��C�ɣ�[5:�4�Ojp���_�W�M�eF��!B�l@*�j�?ηS��s��X���	��������b�c��?)��K��v8�N�Ȑ̊�[=���{�}���9������}^bN�Sq0�ѕU���𦃧�P�"��&�`[��՗����38�s��h��t	C�����l�	{i��ߚ	�c�Exr�����*��E��.� ����ü'O�W4�ʄ�{���� p�~��!"��;��k�_ĭc�L� E�g�3�[U�Z��{�q�a�J$z�4~>`e禩 �\D\Ѭ	��^am|�5�͢����K
��0���Y�̙<�P���>�r3��e��}ߐ1�G�J���t�N�!���B �ǈda=�Ot*EWn⇌������W�7��wO�ܿM�w�ړ�K�2qd!���5���.��a�}[�C�k���5ߌ���Y��aQM�W�g����ך�F��^�Ǎ�OX�8�  �[
�c}x�[9�Ş囏�CƦa����o�M�Ly�3[ua�$���jq�3IP�?r]���t��i�kڥb�aGz���Ji\��,��r�tM �'��~���:3Mq{ ����$�k$�τ�z�yWY@��m�te�6B���������⮊�eW+e3����=���5�C��i�ad�I�X����Y�2&4�>]㞿��U���:��m�M4�+=�C�xN���_�!Ď}L|�l�Yx����	%�mI� �P�D s�ʬ�b�2��o�,�}��v��kfFE%�<�S�y��m�����ьc�Eq8��V�M	T>O6���K��p ��]T
Z'��������+��μ˺�"(GQj��k�G�+T]Q���*g�1��"R#\w
�KЦ�dR=.��h!�Jw���-�;�|��V��V
ʆb�"۟ȫ$��pkL�����
p����_a�L�TJ��ꉮ�y�@ް�l�3hq�1 d��g���F��O�b�'ڸђ(^�g�,|ҰJf��R�B�������� 9��Mq��ȭ�X� �[�/!��>�e�'a�i�-xi�N��rI΍NZt��G�ِ����o��Ro��&��}��U��?�˩�;�Ɂ�o.���XJJ���@��a?vW��z'g?�C*���|k�ym�<p���<H �jIf��A�:���"�E�G��[���o�GLS6r�1��%��]��ek�"��k����m�+�6;����79m�C=1��
�tK�s��o��h?o�󫋞��t�+r#�YFQ���(4��R�D������G3�O��gSq��|��6(�9u!�X-�jy-��;�
���y��ޥv���L�)S���I��=��rqI�9X<�I�A�-ެ�����e�"��#g���&�1r�by+
����o����,X��H���%���Xu�|E)���ǡU�]��5��M�S5�J=N�k[n�q{j,o�h�ha�<�F02Ҧ
:��4e:�k��3�z�c���qBR3��$�@=G���4!%�GCަ$����]h���96��� Y��{��Ql����koM&���C��3����q�RZ�3E3TtrDiP+,��F��E<y���j3H2�=��T��G��o�A�0NcxX\[*r((K��ʹ�g�1�]Έnh��X��|vˈ��R�ۭe�"�����[�Ɛ��d[A��~�v\�j��	�_���/�N� n�2f��M2�cR��,��3��|z1g�,���+��p��/�i�H�G�`�b'�殌@:�����:��,, W#Pv�?�œ.���C��h?$T	���S���k��S-�����lf���yH��E�ClA�u�b��G|z�� �	�I��P�=�ޢ���b���-�SW�%a�ʶ	͔O1%��be���� q�}�!��I�Y�Y���ps-}�j�DI�*}��f.���nd괋qà����F��D��D�TK��'d�}�m�'��P*�������&/�u�Μq���?r�͡s���Û_�+�Ӑ�]��{��*�h�M'fn�{�N���#�T߇ ���7⳱~�L�wq�瑀Z�<���N�;��2ڌ���*�����:nw���x�e��Uy/�uⴀ�z{��L���'N�$o`�1 �����q��N8���%��L�·^Wo5�c�pV$^ȓ�Ω8��Mu����-*�F��
u��4���X���l�nc���Q�^�R)�$JP�����t��b��ۼp
v��9aD��܇���h�Ǭ��y��2�����.)��AM|��J<w�>�9+�*���2�gl�����N��5���5�iҬ�;VH��O��$S�,�=�(>l[�� �S�~�Fp7>LxC���>	C#Q�g�e�T�F�ػ�vFTi,�M��w�Ѹ?��$.3]0�C<�����_Y���~��R\`�2�h`t����'�D�8�7�}"p�2\��O��tW�u����'��rZ�/,Nӳ[�=�䟕���]n׋���v�\�����S�,���97H@�k�"�4�R��(����^��"s[���O[��Ľ�" J��~�,��!�
Ύ�ܿ���vB?TT���מ��&Wq���޽)u�O�<�붬��(E�2�ݶH��r�C<6-�f��6��c�+��n��- �	�t$$C�  ѢW03�ۂ����߃�5yAN	����{�^+<���Z�ğ!��տ�� ����M�dU��]�>�l$^"l<��;ɟ-�9MBQϮ�'��?�-8B�Xd���)ci?���E��VI��el����/v#���������T� �	q�3Џ��`8"<�*V?��K��΋*�0�{��<]5i����D2��B����y����eC�����Z'B�*)� �J��8����{���~�(����og�y�+�1�"�����_.�n�����h>�} ̓�X��~�d�%\�R�S�����N��t1'�,���i���`v�!�Y���R��]	8:�A#kHeA�c�H�%��P0&'Ç�~�O�Ƌ��=9[��+3?O\�����y�����l	�������,�E��6F۷D�i`�Ti��'Z8|��~�,�~�M'K��Ӽ"�m��D�]܎h���;n��nH4�R�숞�;��XG���-�/�-;�>�0���\W@��<�#���;�2ѳ�ũQ�Zi��G�u֏wh��S�O��Տ	��h"��)DU��6��H~���B��C�mu�C]�}k��� 
��1����-N1�ŵZ�7{��<˦���*.�j�d�ީ��_��vP��-�5n��2���t~��{�=H>�դn_��X\������$��x<�;*�T�����/�>���B�aHN��p���3Z"%��E�Y�3�k"�%)�G��uwaѥ�em�wAYg!8�Z_˷/H��Y�x���/�5[ �ZO���G��Y���A��`�~R��0�*���Z������;��w0J聈�^^<L�Kn�[�!	�#h��Bd�K�6kC#+9�^'R���b�%���Yם���E�Dmn�������m��:��$�txt��ZP�QfM&�c=� 4	_�P�`�`Rf�&�=KA�[3�9�A�$��yBf{$]�e
!�l$��X��i���M8�5�Ypl0�%�Ao��	���]�M����}�����!-xU&O�$��(������b��3kiw`��{�����%52h���p�v��LfO��c��E�F�kVc6��]U�K������@`�?i1�����Y�cc��H��