��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���c\�esR&{������o�T�e�Z�/��`%�����1�2��g\D"[ޏ�F�^�h�*�n�7��<�A(*Z�����_��'Я"���I�v�ǋ�q�s�^��\|��v��k,if�[��25�{`�����xSY@P֯�����3�^T�D��׿N�j����Q>��f�ZC$u��f��bZb��m?)��Q0���U[�S0��a/�9���g�y�\��fT;6��8���<�]����ꊈ�s�3�c�@������'�p� 7��^��axw��~~ߋ����
���3H��M�ב�株o�"kzTv�2�"�w��ާ}tJh"�1�(����4X^�C�N%�`^�S�շ^w�'�C���q� �=�t/�=b� �&Z���� �G�u�I	�s[�/�N��������$"���6���@#�v���ܔ�#`2����D�o��nJ��&Vw��U�$������u/ZL��)5�ɫ`���C����^����k�l��T�
Z��uH�R�cCZ5l��.�L�%��1E�+V�}�~�yi��hrM��B��w�y��Yp��xG:]�GD�z��g.��y3\��F� 0b	hEa��x�N��4�|UL�o��-���E��.�@�~F]͢l��F�ipk��i��L�8���A�,����]�Ǩ�@2�e<�Go������\��<�x�1 ~.�[Y�*'_�-�{	E�i�lj�z���.chTY*��t���R�l{(�Xo/�<��x! ��xZ���-�G�DqnB�YN�����Տʵ���8�N2YE6&l6�����r&������\�����[�K�/��A����m�נ��G�~2m�����.�����ʧl���Ɓ��B��4z�%�0���h����$e�YU	�����rW�P��_����N�&�ds:
`�����pY�l��`
Q����9��,�<�ժd��:#ļ+�.� �Q#,~�x������v��d���&q#�c��O��D-W^	��x&����̂��xpb��X����ºȆx�BS���y���C�*� �+w$��4,g`(H��m)h<kV���Y ��.��)�����c�Y=+��
�l|>%D�����?l/s'�gp���[��F�do�S�G�0��� d����4�nSH����(�"���:�Ke��� ]��VI������2�����_�]����t?�IC�BA�W-���4J� U��!�ɝ�EY̊̃?�-S��8��x�e��BQ�,�~ڧZ|#��[~�wD����-Ϭ�����`�	9#��lطS�?h:���(k+����\B�"uC�P��o�5(���N@�Q�gl���w 0��\q{ܾUOˑQZ�m�� ���K�k�۔���r~z���%\�"=���o��i���O�u0	?��"�gИ�/�<��+���Y��W����L��q��TMd:�]�uZ� �,?�"^�t�V��>�t�{2�0^l��7�f�H�G��2+�����b[���z����,�H�C6w4F:��A��C���
)��8�f%��8��&�=[�MQuM��G�ڠe�4�j�d�E��|�����w�{1\�o8��A	�UC�H��
D	z�k�qN3�,��S�ق4�pMQ�� c�E���d��#�fX�D�ԭ!�~�/g�	�B)�?�,WY�q��d�2PI�G�I�Xs�f�p�v;����T�ԸJ�Dފ
;[6���0M�����>�R�a]v6*�&�_i�wFL��Q����3��!c	�~��BX�Ǝ�Q�w�G�}�^��
|¨�.k��Sn��m ͯaEl��s3��Vr�q��� ���Ӣ��������8�HK��!f{Qc�S}��w{Ai���=X�/NSa�r�0q��;J%U�x���[XT���uCd��H�5+p����m��h�.����W�S��u:J:ur��.�J��P1�(z/UFۇ:�偎��N�oP8��Vj�>v���ɶ܌u66�<�~K�����A����&�/��k��N��#A��0�7��H��D����]�Ē5�t�6����|u�a]��Nr�~��(�F�<4��[I���~bp�,�]έ���������a8���nD����9�=�Kl
}�t�cv�ZU}����`�Ƣ�4�P�)�۰�ZBy���8�f"'}���b�'o�@U���}��Fj��= d����;O�))0��WXI&�����(vL��w2j�S��p��O�;L)�o"Bϻ>ٶq�������U�J%�7?U��<��]����2۵4�}Ȉ�g��GQ5�e��]�i��7��'��d0���REc_+Ę2Y�zh}�G�<&�܇}}�i��:�ތ�47�J�K�_#��7�fq�t߮��y�w"��� 1=���_�w�E9�0�)�#�h�]P�p�a
T3��Sl,Z5Z�,�\Qٖ��U���GG6�$ϕa�gu�Ӈ�í�4��9� �Y�7p�n'
�Y0�,r�t��M��}��'�˯܍��޶�X7�B0��<8]�<(�"AYd��̶-�W�q�&6y��g���G�'����s/&�����F_����4rH���T9;�v3�B��I���6Ӣ�sj�HֲwPM�Դu{�������U}���(�XI��WD�?-�A���f��;Yf���p�q^��\�v ��}�"����3(�50ZO�8l�8q}H�)Uiw�ұ	��8R�u	A9*����m��!�����A"g��y��\��:��E�Ĳ��Ǝ���W��I����)����`�!�e|~Y?y�_�����|�ڂ\���yl��'i�e��.�|��㢯y��y���%��.w���3�w�^!��?����p'0'������#�6�iI��8���e��v\����ٜ�T!�h/O	̽{ʱ��ݾ��,����z%R8�E��ϩ8��t��K�E�F�7W�;���J�g\OR��%�d�a�(W%+N�������(\�/�R�oe���!��s��˅ �4�ɼ�G���;�h �����U()rE4cg7@���}�d��\������L ��tr��=�$e��_��I�,����^�v�c!v�l�1�?D�:� �m�&1��	����*,TR��qj�������5l봧���ƛK9�QЦ�rWV���>Z�./[i�O�+�O�鿾����w_l�]��2{^R���)�J�p7,a�d�Pk�x���o���u�N>,���h�f���1`⩛T��8�X��` ��ܺ�g��Y���Gڀ2��W�U����sI?�=<���<�Z8[d��|��+ީ���	�E�+k���D��;���53����!�>gc���X�P�Z�%�Ъ l�0u�_�d��$�|՞)���k��R{SZ9�
��ʒK>��Z����Շ	���R�{v���I{&�`�������OF����P;R���#�	Bɯk����
�(/��cB�SU�#إ�VG��G�h�0<�zl-md��<F��T���*#��턭-g:���,��q��ǘ�O�1�iQ��V<�:+�,ϕ��� �����?ٻ�ފ��NM$����`L�ot�B}&Ba�p|~��R���K�1�~]����{}�'��_&aݖz���9!L�.L�'���Ai����M���'єˍ򍗱��.$Jsy��ݭ�&�+�7�ri*�����0q�bl7�.f�ʎn>P�ݓ���ή�Nӷ�_�n;���^������<AVP).f�.�m�$'�ZI�m��A��R�/���Gl=�����G�@�f{���-�v��a!�!�>\�kAO��DuHV��	�煘Tn��z0������p���L�Ή�x��*�i+�5��hVR	]��xIJ������F�p�=�t��T��k/��#���:�`�̆ͩ�Nm	���ϡ��1E�J���v�x31�{����	��,'f\^��b��Ə�k�4h�z0}!�˪�Y*A�saq]7�Ѿ��ū�Q���㣕�},�-ZE��[�	��cO�����릑/�kjS"�e�B���yR�;B�LѢ~D�;s����ހ�E�[�exb�P���l4ϋ��_�E�������������s��)~��@���8m���3^�@%�YV4�s��Q�ޏIJ�a�Vw��p���LP�~!�Iit��}#��,��5hZ�`�g��a�i�gt"�T�%q_���[LMj�F�/�vƊ����k�a�������4��b�[ 2t�[s]�� x⿁�����F����ܓ��'����UJ�p��׿�,m���߄
8�C�6�,޾�(k��"��<�s��@���ֳ����~ ,2%�DQW�O� ��r�C�I��ա(��=\˄p�r�O�𯎝@<¤)}�Z��_VCn�VP�z�ͬ�bO<�̌�7_r]���9 *�	;�O�7:p�)�����# �WqT�|���D],v�MP5FC��s/��m�3VȽ;|B�F�#;~8LA���	Q������w$:����\���AO�s����r�-|���-P���������<c�퇹�%�.�i)d������,NDwhӯ��z`��R[s&��t�.��k�@dEr�=���̕U�V��G��c�b�U�A�[�7�:�-f|��Q���H��/T�Vw�C��cM�x����`9��B�ws1|I��N �;�K��zn��ܬ�A�0�ݼA�e�"V�F�9%��.��jí$��.i�0�KO�����	���4��@�����	���%���`y�&�v�i3���g�1(Y笚%�ҝ�cu��X
�D��Z�bt������*x���"N^�FV���L� >���S|)M��B@_/31���X�q��${��Q'�lg�9��|x�X��+���&��I:�� �7��3ci�ٴb�K���)� ��҄!B�C�2�	�Km�2/B R14ϩ�C����!r4٤+ �^���f�Z@L3�Bӫ�Y���''x�j�H*�`�L.h��o�F�cO��6����0��~!��D@���T��]�O�f��ĸw��od��7�%���7�O0���7��!�}�1Um� �4f��B�ɼmf۴�|��zn#Ox�FfN�w|��%��#��Nxz�|1�,����C�
_*tn�J��X&�3Z�,� �>��"aw%�@��<s��*t�����)�����\�a})#�o��=ͪ���B�~U+B%����ޛ��_�����o A������2��;�n��R�R:�@�O}�`U��ӡ��/c9�l�@�)G��$x���
g�٣I�p	�x�q�k����'�A�_������[_�O��<F���؆�lW͈EӦt��~�W#�d-����=�PcS��:�V�ɶ.�ܭ������i�qco�}�5�;�Q��g�ŋ��vǒu�,J(<�U�s��V�b���������VD�����%�&d��������E�ca���L3�0�()mm�6�7"t�˟̍O�+W���V�P�KMN�P*��+9��9k+��V���n����es	A��1�,���E����,Gv[s�l���SK2��{�|���q�n����rK*:��N6���@?:%.��v�������.�6B����;b�	|�@�+P�d��
P3"�!�(�yV~F*���"(�l�g�iǀk|e#;�p�mq�Z/Ѐ�aB�6b5�J���W�"�C�:`�j�5��O�B���"A>��9�(�2r�
�8�ad���CA�G��;v����:Tτ���0@�?�'��舗�M����(c�/c ~i*^}���p�`�1��Q�Щ�I����U�a[t�>��"o�CU��B��6�q�h�e�D@�[�P�� ����*|e�\���/g���+��H��DVm��;��v꼢�r\���/���";sN}%wt3����pX������)O����@�������}�  �g1y�|H&|=�2C�F=`}4BUy3�.��y∂-?�:wD�ˎ�
n���v��	Į��U��bXO)<8���,Z�6 �|`	î�I{�s�5:�~�d#�tY�,�/�`=On�jq�4�ٺ^jHfj��F6�0�U #:$�=��ȇ�NU `��H��S3q'��As?�P4t��щք����t�դ����۬�F:����d����q{�0�>�g���� -�8�u�c}�?2�X=`���k���&r������ヿ����8�Oң]:�E~�F<z��bJNs�Ξ $� Jb[�$a6�8��h̰���Xc��c ��7���{�W�4&������|�PX�<�֜4!�7����?GYvE����;515��~
q���~���[�o�	"������L��9�m����q/
����픬X߰X��dB�A�y��ϫ�~rԈ-)\`���{�陞sT�Եs{�>riZiz�?���t0~����y���P!��A��Nb�ٟ�ً��?�R�{u�.;U�n�ԅ��Ff���-�ǓHW�°U�P�6�	J|���	]��d$���2�c����hGa�����z��4����A�W�y�%v�	����bH��Z���%���Վ�'z�	 Hj3z�(_E�+�v�M��)�f�׶=y���� �د�>�9��[`ܜGa�@��˦34|Y��!�ڟ��Ӂ(_�%Lg�_����!�b��܄� �/������O۟��X3O���PT�!p�;��^ԩ ee��� ��K(�� ���X�nz
��s�B�[Ck=��ʁ�D7g��S~5*!h(�Fp����cm���g���[J�z"颖=�Pt�}�6~%�8]���3/���I�G���qb�8�>e��HC���$~�2�Z,����\�=�e-'��ǫҨ?:d�k�ꬄJ�8� y�'Nw]'SXt�����#^:�x��e[�4��pPp�����}��~��=��W�J��Q��\��%@u�F72Awp\To~W�K�J�������,�Rf?c��[Ͽ�N��l m�Mb�'��+�IX�>�q��Ԋ����Զ�}�Y�M}��6��4����]܃KG��Q�J��GQ5}�m���"���»�u�ƀ"A�G��_x{��(�g	��"��Vd��\r���N^^B�����z�����̔[�
~�����əU�28> ����2�͋���phF*^�Z(�vKl3�H?�y*���1���Z�X8�N�އ��t$RILY�eO��y���S�*�`zj��58�nM�\R����(�{$��@}����}e��4|2�j�ͱ+꭯���� 5+�.kM���%>�L1<�{���EP�[��F��i���3S�%Š��A}�<~�nC���п{8Av��y�|#��0��
-�j��	ĵ+�4���`TL ���6���S�,��%� �-�'� d�p:�gM���CfF2})�zo�;٭����4��z����5��Ed��!�i�y�:�w�����5P(�������M[뽑JA�7(�|5�mGYO���h�3�%>��9'4�k�c�t1Ԍ�N,Yo�8VU�Jj�����C��7�PI���t4�+$D:)Tq��@|$�E�b��q�S�ЫX�~Q?<�UE��p��'�|��l/�)V����?3��{.�C��'Jm@�X�*�3�8�Wc
��l�{�H�1�)�n7�S]ZÚ4*�J�}�{8x��2td�%t>�QEUl�B�֍�V�L�6c-��