��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9�c���]�uJ]�u����`����#��� �]�� ���2*\m)ۣ�����/���>߱2Ҙ>��&+\����O�6�O��a=y��� x��o��n��0���� =��Pu��(��2�����?��/���PS!�*�����|�C�L��q֎Iл�1c�{X4�V�xs3VZF��#ӋSS<Sa���`m5h��G�*��2�8VʕZg�aT8G�^㷏����|���|�D�N�^�u�9�n?i��N��������!�Ǫ�i���#��D�@����{��15DM��+L+Z��.%o=,��f,��n�sM�vp�QZ���9��(��;u��M<3o`���d	���@����!�y��Dt���6'��C8(��đa����6�n��N7 /���5b� �y�'��BkC���H���
(z� �W�.Q= ��~����}�Lö"�(�~�($$r�=��%;���{��+�w�ŵ��%w*h�����i(�Q�s���}��1s�]tQ ��d�����	��{�?�5X�U��m�U�^V�����l�����rY�����~aSIc �����n	w�.J.����ɝ�^s�Kne�%�v�rӹ�ף^/g��o�!��`Y)
�k�����̄�4���ʫ�T��nk=e��a���$_x���q��T\&0z.K���/j>�e���:�o�&|��8���h%{��y֊9�dS�ׇL��-^A,��A�\MPp.G��&!�q��,���)��(���x6��B��[�V��ٸ�yq�j�1e����E�\��xZ^�V&�B�Z� }����~sKh�<�' "q���[�����[Q�� �飐�`
M��7�\��?�b�����R�L�N!�Y�N趎���d�C��r�Fe ���|����ӕ��]��$-�r�;�p�O�ʍ��v,�e]Q�� �E�СMv���<@e��(�II��T��%!��$N�s����8�W��"�q}���~5-����_/�l�bM��B�T����9,][�ƫ/<|�����q�������ش���� D�������Ծ,���ۉz��0�T렎���L����V����ZS�c��@���O�r��!A���&���E#quYu%���P�"*�OB����S�gH���L~�sC�4p،����J
I�o :$��7h~��`�\#�~�JD^��w���I��&]^-Kt��k�8�6�yg�x=�a��i\Ϣgq�A���n� �qUaz�ŷP�`� ]��4�CxAY�$MR鲴M�
.�:֓{�6:����E�l�;���TMdV��Yq=�/�� ����7�w�vO濇�<~9ʋ��ʚ��]i8�۔�୒����j��5���鳤�~X��C	߼<����W�!�2g��ޮ=OtQ�D˃�&��s�J���j)s��Fw��H�����h(V��P3��OFW��3��V%���(��uIE�H��Ť�Mo+ $98,���~���e3�Oe�_J�{����e良uPӯTb�����؁�ӛ��d���(�d���q���0ع�\��K?�/w����_Z����a�&|H:�1f��pՅ���A�K����a�y W�U�LI�B;�����/%����a�.��*W4u��Q"�"I[�`��Q�8ZnRN�N�&�J�O���ٽ�Z/�y�>�oC�/�%�}Z!��� �����aھ���gFl��Qr�(�c�ye���vugLޥ!���?��;��Y?��4��j���X�G�p5��$;��j��L6�:��f^��Z��^R׀C'��TD�˫FC��#��EocҤ���1��'���A�l�!�6��/u�X�|�&�a{�Z������E�Ys	�?�.���90&ц�l�c���t[��kU_h
�b����WV���
� �o.C��-�o0l�\��Qe�l���L[��y/��?a�A��b�5�W�U�w����f�D�&h���C���U�����>:*,� ��N"P��z�Pju쯘�m�R��-�)�R?����"�5�_t�#�ł]z��,�]3������"L��8��9k�_))�$.+�I�AoT#��潡3�S�o���ey�X&VKKy��1U�Y�^��L�[ZC�*uPX�\��F�Z�R~��ܣ�y�9��H�UR(������Y��J�K�!q�}�R��|S4���\p5�^��Ly`W�6~�Y�bK�,��1ڼ�S�I�Z�E�Z'6I>���B�[?�))�R�|rj��aU&����KDoO[��e��� �,IcZ+y�tB����遆(ps{�kI.#T���A��ѡrpA��&H�����Y�c�P���:?p�P��F4��+��@c�fG�+�u͖z�l�g�}�;����7LG�'M�a�g\��3G<�\�Acy�dK��J��U#Zp�����ޢ�n�5���F|�A�d���#Г��MXE��	��k_s[��9����s���O�"�c B��� ���Mo�J1�q�e���}J�5|�E���(�C��G�������mВ�}A�Cr]�_�����]��0��#�u�.6W��p� �;��O$'��W�l�JI8�U��I�a�1���	�����Jqn�\&��J�`�[/h`�(\B�r�^T�4{^���(M^!�c��T��'�k�8+2�u�ӆ�R|��[DF֬��"}���L1�N�� �}��/��ݟzi1x��� ��Z
G���FUڝ�QK!(�n_:�M5.�XG�Ƶ�W^T�]a\r�>o⋱���&ϻM��-ٸ\�&���RZ��ᥱ^x�[v�K֤��tdsEu�����u�R�\V����-o�����3�]�1�s�����	�Kz�ǹĨn}M�)�T��g��{v�j��EE�+^������{�[V0����:!��f&QL'�8�����uv��|-P{�b#|b2)���Q�p�u�I�C��YQ���q6���n�ځ5�D��1F���E�t(qVM���M�,/\�zɥ��䷿�c$�lL��T�~_W-�)9���_@g��$�	 �9˚6j5�9頶�ek����ʓ�^���t��M�Jс�\(8E#ь�UZ�vTنǾU-s�2��E	����֦�6_�}�\2�+�ˠ���M�A�6^�>�,����u���E��Kk�-�z7/Ǩx.��8�X/�^8�e��W����������I����
����@�=�c&_���\�͏+Z4�X�s6; ���#�AS�{�٫�GL�3h���S�<9M������Q/vp�����7�*��sM@R�:���H�����:��}��(�:��{����f|v��3i�1^���1u�F�f4�N̼z:ZN����1�{5�w�z=t�����V���m���8���iV�6~YV>z��nJ�9*^�ÖV2��v���4��|�	�֖����I?�Sh��w���*�X��g-��⧶�g*����������.��#r�+��e��I�ߍW�ޅ�ǐ&AY�F�,Q9���;�j���/B-����u�DCp�#5��mԣ����wH�􅡫��� �-�B�;�P5��ӛ����-7�P��]�fy�s�/0~>�+�d�������㌄/���xni�{�������V�9�]����L��(5+��Sk�v7��`��eUOCz/���h��յ�T��k�|��,��B���m˻f-��	B0�DZ��B0TIl"ZP�����}�D��:��bq�ظ�[N�<�$_`^Qt`��~�~��7B��?��Z�ۺVM�h�=�1"_�S�\��\jW`�vZz�������+c,�x����[[�䷖�@Z��^����_����#�C�i�f��ס�`@�piH����6�c8�����>����aO|b��
Z%�5��Px�\���y��#���Om#��k�ZB��2�4:�p�(G��S���W�HLr��q+-��59�����A�����Ն���U�#8h�#�TϬPY?�=�O�tRcN)�c+F� ����ǽ�G����:����O�T~���&�����gB�F�\門P��R �*po7E%����5:�H�������L�R�[��E�N��r�B�p
��� W�B<t2d��E$��b��ǥ�cW���Wud��Q�s��2�i	L�G�#�~0���fpE��f��@[Z�ǀ���IR�301�!��3>x-���������������)l#��9_f����ʇ�i݁dˢW+��e��a:i1�	�.�}+s"�^X��":+|KX�N34�P�>P��p�?.N52��8X���:����+���P �i�,1Bz�6��Q�d����u'zF����C�7��2'?IF�d�)�>����������%���8�(9,����ۑ�[�Ԋ������4���X�����ɓ�D��BR����� F��H�ikB���3V�8g��h�-j���܍����e�y�!j����^>[�l����-������^�lh~�@BH�ԏ�N�7K#%�K,�q����i��(�8�joWQ�ָ��g#=��C<�וQ����<+�vJ0�|D%_h��J�:o��jz�%�V8k�JĜM�_�����p�r��#�M�>;F�o}��qSdE�����ڊ�=���ŸD�8�@��`�:J[�1v���['����8nE�rf��P� ��p��\��v�1~���i��oy�mh2�+����l����>�w���0?������|�F�,���Yq���R���C<e�+D&o��9\q1K��*���Č[]��'5���/�,�ºؼ��.i��C��V<$�T`�P�Rߝ�i�Y��7���]�R�=�����
xT =c%�n4��j��9öPZu;�x�0��?]�\P�O�ʚ"�DL��H�,�[xQ�E�Ǥ���i�Š�Mf�⟿Փ94�Vuo�
1m-���[E8� ���# ����� \1f?CY�8�ҨK�[S�p�ƶ;_��U��#����Az��xŶ��L塸]-):�\�f]�$E�j�B`�[�
����g�