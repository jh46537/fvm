��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����G��l��"�Fe]=�/>�"�3Nع}EJ0���U4�q��q��i��[�3W9^�LU�3k<�ҋ�͙.$w{�d#?ŧ�.�&���\�FaAG��Ƚ6�o�� ~[Z���~s��c!��ء���]N;k����h ���ZAcd�q�4S3�*S���k�!�[�>�Gf����tZf�ث���Ta�z;TcP�.�Dz�Wt�'�KC���h�����D�����5G�j~7���w�q]M�����u��ɲ�9�#���ƈBt�L�Q1.q4���v{��і��гX��"K��8Z!żD T/�P��x^�அ�#�U8Kr�%��;���?�3k��̓��}G�|��3~L+�/�/��j��@��b�`ɘ@�}o(�bn%Ze�$>B#�|ϔ�}K9�	#����&i�='��03+�B#L3�"��$I�<0�i_-g�{(�K�)e�p��נ�p�I��K��E@|����9�,3�/���m������1������q��p(}��*������w�,ʾA_>���6����W���GHDp<A��F�P����e4Q�g��}�LpNz�52�#��"�C���V4©��U���
9�lY�Y�Kvi#�@�Pps���*�c��c��f��]k�zhͭ�}����z�2���i� �{���4M4����5��I&���P�7��b���isB a
��ט�&���=#�K6LD�l��a��\j�&��A��.�M1?C��N�;��]���DNB��;��f%���Ғ�:����斠Q=4�6��h���/��W@+�t V(����~ r���������[k���g�c����^eX�}���"J�%n'��wVd�pC@��;q���!�%�F�.�d�ʐ�Ɋ���`_���S�/�F~���[o����g'+��7�U���Q��E}��<'�5�x��m����|Z�F��E)����y�W�5^L䔨�J^1�B|�X7 ҴDv�������v�vn[Y˾�2��j5Ir�|�ؓ���U�&��U��u��<�>;.B�cmR.+