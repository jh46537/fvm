��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�u㎺��`�R؋l�)D95F0d"�s�>sP�T*?䮢�B���M��&_>�l�L�,_o�`�j:�]	�'0Y�ӂ~y1�+�Di�����	+��-��Dq�f��X0@ �1J���JtFΙ���+e�4���t�����gp&$Ҳ)xy��~H��F���r]ֆ`v��v�;������s|���#��i�g�ϭ���F�(q,�A�������;�wA���V��S4�}~TH{��
�&o�jK*�G���a�Ue���x���'�uAK�)���JN��y�-��:�q"� �<(��q��L|3��H�8oM)W?���\q����;�Ҧ2\^��r+�0���^�I'S��0J��35��ݛ������e�β�q�L8:�1x5-gS9��K�xX��+�K�Z��~�=��x�+�[#E r��#(l����#����I���<	c$tT�ɬ˂п[�q��7���V5��d�ɟ��L��8�f��i�i_��ro@,εڮ�z���s��v�Q4|�m��e#��ԸS�|Z�C͹,V1@���ՊA�\�IS)Y;����<�t0�x.8��N#V>Rn���^	����	��-I�ƣ(H<k�d�L��n{�5�J��n9�YO�>Y��^�.�\M��}0L�Q,p�Zw���)����'��ݭx��Þ���Nd�\�>�ܨ������U�)��7�䄒?rU3$;i�LX#B*v�o!����S͎���:��~�u��c���A����BB����M�z�^C�z#��˳� '�=�j�(ST	"�DT�q �*��8��(ce��f�!��·�ܝ�ة��0"�fI��V�-��������:9�7Ξ�l�V;��2|��{#�W���S�yk&�x��_�K��d��!g9� o�9N����jJz��^d�o�]6�:a���
a�O�q�=�w����5e�±���I�YS��{/���;��cmG��=������7�aPP�;����Ӊ``��$yI�I2�u�(�U��J����'����Tq�zwi#4ׇ�
���/I:2�������g���@�^�1�բ��Z4�=����=����fa�(Lh٩�+٩z%c<�2�>� 3je��[�B�<{x����N�"���i#�Y�ͨCGF��r$�ot��`G
N�>�L�.���~~�r��&F�ׯ%�μ���	���aGc!x+��)�EǇ�Yf��y��5{+������Ii��da�	��Ydi�ӹ��������ϱ/�Hn�;e�JfkڴU�ů�X�h�� �Z���&Q��������(�<��}3�GQ��`�'�O+��V��S&lJ��K���?���c��7�h�N�@�����N� N"��|��h�?V��.7�GpPm BK���V��8ct�r�����?�\��}B\�4��[��ڗ3 ��EW x>69G��4��ch]��A#�0/�,N�5�痨�aA(&{�wR�sm&j�͘c���de�'�F��E~a�p�:-k�;�����H�V�Ρ���D{8�0{�0���V����5��$,lOA\7�N#���0�
����g�cHj�}�!BR����z��$20�v��k�)�R�q������؉&��aĠX��	R����!>�Ԝ�5=��w���-���"S��8I��9�BK��35�%:�7x�1�g����j�e��Ҏc�!�\��t�C�:[j7��!���"W�	 ������td�S���ݪU���~wÎ.��8�����F�/�ڤ"L���B�ý�I��?OS���b��ؠ&�?���W�(x����(vme l��M��7��V5���U�:��ᕑϪ�_vs�h��v���8���φ͇c�|�rIMxI:����E��������h�a�OM���"!��]��?ꈃ�ȬW�`����r������1��3��rp��fpC3��iVs(7ՙ��H/�$�5q+�����@ŏj����;~�bX�qa��� Û��.V��&'��q��-nF��uJ���Y%ݠ���W��N�-ä=�gJE��L��_(�W�~*˓�����3QT��mO���.�٠�7�hEY�q�s����"$*� ��̾��.�}9�X��9�N^gD�J>���b)����enA(S��6X����+�%�
�Ծ_�G��c�@��}��b�`8?k��(���zم�.��,�:�n���[�g�H�ϥ��(�չ�۵^_��(�>V�Z �t[���qnF:���Ņ;���7�{ʎ��� ����u�� ��v|l���h>�
7Z>\p���њ��<ڤ�I����ٍ4��4�|���c����ӭ�t�����v�WH���o����	��)�y�c �'�X4�[�	1��m#�mǻY�L����9�&�fz�)�|�ݩ��f}�u�n̘-wx�-�Ôr���lc�����F16��h��xS�]%��C�|A}�9 ��}��lM&T�@�l8,����/�T�P�3���8�%����x�L*�LJZ:S�8Յ�� ���p"-�i=��=|ēH����Z�M��E��T�P�bjD@ g�Cђ8h52k�^����B��n��p)�ÒNu��A�H�B��e����Z2�����5��CB²%�8^��D�sPi�ԟ�C�9�#/�hU��(]*!����|���7G���?M	ͻ�[��Ԁg�Qڍ�?�Z��������{�*�4�o�B��ӌ������i@6�����:��̧�骷���b �}!T,G�A�~C=:�]xn�G�����{3�d2��<Hk��gj�Hv��U�Kdog#yn0R瞮�Jx-C����;��8����N�a>M���d�+LmB
>�+Ё��P���^W��}N��pP��x�7o6}�*��H-���Ա77�ڌY /��SQE�~��� �ʥBf�-8"���x<�)� �Z�Pv�戲dk#����/�����h�~C3@<�$3,]�>�6<gǠ��ur���ǳT=l1�Poܿ@�8E�:�ʙS]9�j	��騹N=Y��Ϯ�8�G��1>�WQ�֯�Ԍ����F����]�G��PV뤎�V���0�.�x���%3��F�n]�����:��>�iDP0Ð���'*���=O�z����ͷ�]^Hs�ֺ��O������&1!;�=KY���P~	�G�x	�J�:Y�JRI�
\H��)������%-#�F��J5�wtpb��`-��͝3�W�֡�
"&��F������PB0	��,�Mو��ᛸ0DZ��e��s��J��c-M�o�aM	:>����0�$��&ř�oy�7�T`y:D�
L�����dW�@���p�6�F���|�?3�YU��P���K�8w�J)̎�$C�~ ���"v��;����~Ff�n#���a4<�BI����[X�
�,a�&0L���PD��<���n�y���)Ŀ���%:0��Q}�13���I�q_� NuI,q���b��"��5?�DЁ�N%�&�0[K��r��b"� ��#�x.���!\�e�d�nG�U��\��4�Ŵ42����K��:ʉ��]�׸�Ju�9O�q�ç�G�_N���C�s ��p�Г��y���
��^7���3|����w���JJ�n�����FK�����Px��������PRu`���X{��o���[R�S��#�e@B�bf�����p��/�"�~�/�|����\'��C����e��3�d��6?n�2���㋿/W�l�Ĝ���	c��5��%�ԏ��tƚ�܍7�[ �pV$���S(�~�� �#n�F0ʌ�Ni}Ѱǆ_��P��SmIZ�.L�PU]��GD�o�M��`�������{��� �aP��R5�~Wt�4/���2�B��'{�+��^��*�ا�C�l���H�R�z�	�� ��5>�����׋҉����e���+�$�J'^�f�x��E�`/�6�s��)��}u���>�'o@��9�ՎT������ac<e��k����.�:���6e��}�s �A�eE8e	��%tB�6=I�����7�j��B��Ҕ]6����:Q.�\M�WO{���/��q���o��ٷ�*y�%;T+b'���1�?2�#�5����u�������ҝ��OaZV:�����e����1�=Jp �o�Rvu�N�$�V�yDC�]򘎩I��,E��v���BO1$��ʷ[�ޣJ��R;��ʊ˯��_]�L�F��������-�-���]4l��m��li�.wE����'⢀IM���(я��9^_�S3�M���59��E>Zo�>���W�sK=0~�%8�1"��J��[Z6ׁ�`��߳{�T�/��v�[!����������f��a��JA����"XY\��"�##"抆i���o�9_�njGa��H���0���6d�hj��M��
�DW���|���?1���IGP l(�h�%*.#*)����q�r�u��R�(/�I!����Y�(Oϥ�c���������:�j���)��8�)Ҏa�'�)�Sc*�qH��N��BV;���[�R�P�b�ΰ�?��'S��+ף.�V��6,�U}��P/�cc۷�+k4N�ѻ�m�
���+:�T?u�)�<>+:���`��6�	�f�Rp�mm�AL�Cs�l\���m`�X9i��(��"��|��Oo)�z	�)��.��oA��w/�W���u���N��x���(���z$nNjYAT�s5�Ql^1Qԍ�P � q_�$��yg�q�F;`�w��1�i� 
\�ה��H�~�~�'�fC�?�>(F�Ѝ��-��(�)~s�Z%�D��8$S�~:#�o�W�̺N�<<���9�,'O~��*$1��2=�%Q���X�ʼl�}?�xɵ�
�^�Ȭ�jg,.I�[�dSH���/��U�t��?�66>�׏b�Yk�xC�16�puȧ�����Ir��M�J�Ј�F��Y��;t���;�YV��m���Fr�/ʆH��x�D�N�Fp�܏�˕ 6�����~���o�-�g��F	8��}�$���ɂ��� ��Ev;ȴ��(����,0�$�^��Ǒ�����>�J�-'����U�T���Ӟļ�.��C�G�/�܇����\.�l��5��#f���s��{��O��.B|Jǁ��*��(���4r���*�%
o��G[P�o`�|��?��rM�y��1&vz�ɔ��.��ݸN_�]���r��[�U��Y�)f&�M;�G�=(`9פt-xU
��A�g���L>���o�AX��DX�~�S�)+�B�N�6�8��qD�!��KR����ϳ$wķō��&�)��A�Y�+�}ґ���.{:t�"��U�LN�����x��7y�HeW�����v(��l�G�i5$V71�U�7����{�o<t��R���h�0�8���^�Jm�A���Y5 ���,�	���?���kaa���*3����`e�awVA��?���7r�똫2,�o�IO��g�C�S9,Щx�,${�{��Ӻ�����7g�7�i�SݹX����& �.�q]�/ʰ�\��!�a۠WDG�^�e�k�SR�>�
�/uT�*��+m���k;�)�� ��׺
��$�9}Ch�������V�d�񜨹�(F�4"mnZ{��20]�94��P�et��1{<�X���ᗠp	�3(x�P�^�=ź�-�9�l64������$SR`��P:HH�D&�^_&���þ�NR#�	�<�~;R�� /�/��̏��̞j��EF�CX�����]9����Og��Q�B�Xt��M���Y�O���2ng~W��һhh(mױZHg��jʅ[������rM���&nC�r4\9�����vޭJ��}u�ܚff��r1_����G���C=�0{0��c��Xd�i7�$T��P&z$��_�(h9�0c�L��W+�@��]���|�>q��Ӊ;�ҾH~Oă&���,�z�3�E��o�0�Jh��I�Ѩ�r'��;m!_Y;{�n������A�[?�)����!�<��k�nX^�!V�Sᤲ�L�z�A�k^�������q�2������S_K�T=�~W0��(�bjI)�̎�9��Wg6�P�y�B���
�'��Ƴu�Ha0�u��6���QG�e�V�C�'4ItPn��(�q���~�gf�sK�����R��M�.?BA��1"��w�@��S�
&L���ċ��e���D�)���<sb�"�ί�ռ�T�ڠV�4,0פ`3�+�;
\�/�� �$v�$h�DH�zx�����g�ّ��=xA¥O���R3�>�UƵ���@�eS;�,!�r�S%�� yv}��Dix���66�qv�'���Jr<st��8t�/��KDNX�C�]2l�������ebU�9J�Ƞ`9_�v�&�*�K��k�!�bտi�?������Y�X�
7�1Z�Q�xqc@�Px�F���t��.S�n\	m��\�Ƿ��Y���u�����ݲ��G�X���@�Pd:6�HD�t�vWc��]�J|.KD��.��� #��Mg[P='��j&���>D_fJ�V�(g�׹�%E����ABy1��b�2�� $����p|� ��"�Yx:�D�6�\v�i�� ?���*~%b��|-G�P�%r�ު��;�RBMkl<�s˩�<�/i�%�3�>����6��j�=��2
ŒJ$eB���Do�rse���P���9�����(�y����2%`\0�,��MU �M-�#�]�ho�~�NL/1�O:E�9֥)+�dn�M�a�{��[�S/�	�gV�F�8T�F�D�pᒍ�����#Q�\��8�I�\�J�&EG\	N�Nxb�ȟZ\�MōI;�i�-���Ay�>Up�>���z��jJ;�WAd�T�78���;*�o����&8.S���CXTI)����*Y+ϮPP��H���g�@��C�j:S��T��3Dm՟��їW,��iŮ'+��1�R9�_�e�{�L���iԈBXR�UM�.���ܩ�Ԓ�U��Q:���:��6��W�Ĵ��a�Y��τ�7g��/�$���!�<�B���%�3��MN<8P-Pn����w�a`�0ÚzT��p�C ������ݱ;g�+��W��5�ͫ1��U��(i	�c���<�=�)�AʨN0K����~��e�63�V�W>�C7��)��9�+���6�.*������GS����?�d�bv�q��"ޓ�·$ߓ�%�o�M�Vގ,~�7��|���0�9�R��ctrA�oz�h��`���@��d
B�2v�٣�3�>���z�z�c�1+���)<�>�/r���t�</�̦�ٓ/O�j�	��*0�Zc:KTC\���c����
�[��V@���-l*62��UځR�p�h>��4��|�����2�@Rg��Q�7��S����8��l��t�)>VП��	�m�:/Q�����0*Ѐ��P���T0�ڧe�>�H�GDMEXV
���t=q� ���^v�I���v�_K�������x���2�V�䝭ɰ.p���M\��T���qub����+���ň�2�{�ŧ�a��z`�7�<r:�Lm��?E{@Z���u��J��ux�U��U�ܬ�à�_Wdz[���Ǯ{)�ܞ�n,���Q�&E�.Gww*�5����9�ݟA�r8���i�\ ��K��ƽ`�	� �G�7����|�v�l��
g�ڔ�N�� �-;1.Y�*#n}2��\�.p�\�����pt۵�s�5�S���p,gľ�J�B� >g�<"�|�'4>[A���)��v�iv�c���H�v�m*���>��}��.�wg��I�aT$mt�)��5?C#��%�Y�+�9Ę��)gb��!�Jl������8@y���y!���H�oA֧o&�OD��O�Β�_�Yr���&[)8����R	��%�֢�O_N=pL�_a>���M!j����K^U��/�wgG�ύ�3�D��m��'��w�鵅���u[���Ǳ���8����S8�T��p��/��;3���jރh�B8	2�|C��=�bj	��ӥL���
�Sz���c}�2�x��ͧ	�=bC����aŪ�V�m�Nq�V��q�H�5b��� �-�%}����rc;�d���@�.��'���cD �K0N�ޕ�Nl����x��Lg�^���Ҫh�I6ORM�00�����{����[����s�#��7���5ߑ����>����mE����a�C��R8�VD�`8�������U�a��� ���`V �Bkw�ދl0��/B�zw��1����9E*4r�j�&�0����Z!���[u��UG6'�I�t$�{��J\ʶҿd��6F_0o݄ i��\�Ἆ|�z���g��t��/)<�,���paW�lW*��ܕG^#g���0z|^��r"�j�R�w��q �,�8�)�\o��MW��0ѧw����A4Z��!��PoCJ���"���M�����/Q�_;���74�~h1k�0Z�,oV��u��W�~cwŐ��n���pI�|B�Zd@�����L����_K��jX�q�����x�������MT&�Jߧ�f��7���K��y&U�-��th�r��ՅAr�'�t���Y{I��6����]�fU�"� S�򽅇:��WZj�Mb+����67�fو�c��P>%��w�/:���U����@��i����w�����d�I��
([�ZWa����1&�.]xi�w{�3#�%��-Zz<e8иw���\��Tq�"'���S]˙���=�hQh�:˷�M�p˲�� �c��N��:�7Dm��A`�mT�FY21�a��g��Y�̽@�~thoK���S�T�jz\�ɖ���O������y"�{�IEd#��W�E���f���Q��.�Q8����X��g��'qd���%��þ�~��Q���6��w��.!��2�ݭ��+�1�c�Ɲ��6I�a����Cϲ��`U���,A9����ti$2Y�ۚ��:�2�Pq�]����tE_���Ra�9�nJ4��Z�)`L��T���@FBy���k�%����N+H|��5�Hh;�nf��𒮑x��ɨ\u���q�k<����&6�I<�Q��V���?�ŉ����-T����$mȀ�=��Q���
l����s �b�%�	�]8�^7]��70� ZF�-�K��������b|*���܈K�B��x��5�f>�@����EƔ�?�
����ؕ��M�hJ��
<q��N�Nd�>j��R#0��L�eHI髌�!��(4.<���A���S�'j��  ��rx�mg�2�Τ.���:��=��	Wj;�����6�Oo���sW*̼�=�o�0 �yy�T���S����J�W{�0JV��c�LW
ȯ�յ�!�L6I��CW�μ���
L�ߟ7+�5$*�d��C�����d��%Z�����H杻eָn��O�n�8yR� �O�t��I��)_�/E
��f.�����_5 -jO���;�Co��}#Z^v������vH>���-+�}g�qXb H���]�;������^o�MG�� {S�F����s7i�n�����4(�n���m�Л�>s|�ъ����Z����FpH�B͏�+>�|y�U��o���E{�
R�|ϴ����҂S�3O���}�w��ͻ����1�Ή�Նu%�<9�J�pA[���&7��=�[�_a8�	��r�+���G3P�pbv�����<+W�?<ۄ	��aQ*�,aO�VFsP�U�Z}�
�H,T�@rG*��+�|�r��U�Y���@:�SFtb����C��p~���[*�	O�b�tx�;0��>�$O�B�I��<�$�P�K+�i���>m�M�M5H�)��*%�0klD� (�gY�"lA}�9��P����UKM�9e��H�����.�6��;�N�5'�u�+9����4���?�[�Y�Ǩ���Ɣq5Qd9�
��S�ZR�,
3�^��c}^���w������o���	'f8���J���}_@Gޢ�&�ţ�d����>������2!5�a����ʔN���(�Cs��:K�r�绚��Ͻu��x��:���|=8Y/�>� ����}���x��qY�K_�/FX|,�NYU�_զ/�	�<�������iUa�K��'��r���k���,��e*��iJ6pf�>W�Y�� ��:'��Q��D)���/>