��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{ς��$�+���>�1�%���6������k� �����Ti�����(��iE�Η - �'��ɺ�i���E�-���q[8N2�كbM���у#�٘|G�2M���f*�EGb�@m��/$
��������'%�b�:�x��3��u�寂pB99$ў2N��k��~��ɜ�(��\J0����`���$�,�f���� �4����.���8Q�\��=�8��z`�th���R
�@P�m��|H�0K�MO[�h���@����&�ޔC#�����aCz
��Y�PO�<�Y�$`�ƚ�"���i�Ǜ塶M�Y��"PA�c�W�δ���z�J�*�5~k�
q.)&#k]�|��i��y,?T�f�s�/,�
��XY�P�2r48���Y1m wf%3֩�+N^��l(�S�O�E���+�+������!0�
Z�.v�)X�!h:�uG�6��
,�U�W̩,|?)1\���CE���cx�q����oy���܁�2-�F���H�m�?�R���[�(���H^�[˄Pq��, �dNf#D��f�	��ϴ�$�b���[��"�{Q,�����.i�k.��מV���;{��ˇ�'o��:���W,���.|�4��`$�J�W(5w�J���9�_�؊^↋��[�!��,��L�� �(P5��m�vT��'Od�ݣO<,�=UGj��x^C��t��[�+e�'u���W�}��Q��豟��6���Nk[���r��$�@��r��N�@�ō�����T���	/�9)�{FV�FI�=mhT3C�\�Z�RZ�~CX�v����� �Nu6�'歎�
�{K<%�a�#�,��K�.Z(w����3�"�~~O}���R����5]�x{�P�D�U����DS)|������S��G�NA)���w��d�����~���s�BiCԟ%C�Ye���Q��\8��6h���z<D�^��cj�;ֽ���F�襐p��1�^?/H�3F��-]�5�N^���*�tx��*q#�{��/��rY�Qn���
tܨ.�PI��^c�P�+�
@E6�j�"��E$%����V��xW.j�v(��WAv��κ"�����`f����R�B��WK���br�u���^�$<��w�Z�c��+u*�f{�����a���<>��exW[@mr=mі%#�1��������?}ܴ����Um�M�3iF���#F�\��9sG5
�K��Ѭ����Fi~��S����֎ez7N���bW�Ge�)Wp�+�m���Am C�S#v| �~h���m; �k�x��]�G��B�R9	���`:��{9�J���з�п���
�GT(���c� �׶t�6�Y���c�,5��E��4h,z�9����*u�ܓ�����1jc�G8���ۡGA=¬S��U7����G�Ʉߐ,����G�>7o>}$>��#U !�C[���H��$#��5b�\��o_�Ԅ�$���'	�f�|K%Q���qf�ߒ� +|i���zU-�nx�/�ڲ���1����!��$]<�6\��x�O�:>0�����?h5AßX���R]���j��Ie"kM!�5A����J�@S�l�B�SDAeSx�C�H�~��TjW�G�R/�m<��&>8�3��a�)����m����=�,I�����ڼ�0I��.�����: ":���^�gZ(���qg�v*0re��Q:��X`�U̼QA�I�Ch�:��q���[���T��r}��dXP����9�ba�<�D7�x|�W�m�z~��B��V�veS=ludH~Hz�~"���gu�i���އ~��T�%DN;�2)�����3���SYK+zZ���B[��� �[cH�,2"��e�3�Oo����T�u"zRD���x�����n|��)v�Tá���#�e,jĈ��W�.��b�ɔ��uG	��<P�*�Y
��DR���5�X���#��;�^BNT�>{���zK3���v�K�п]��صD����;�~U�X��F�k��(��*�V[�����>!R�"2����_uY�9tu�)�ϖ�_��g��4M��nݬn���Uݬ.�D$�QD�T��r�w�"�P�,�w6ܦ��g��Hm,GY���+q�Z6��Ti���U��o��>��B|�d�����[y�q��[~,i�YM��$,�<�%,i���fm4�ph�H53ۡr��u�ةٰ�x�~gH���^\���F�"�l͑>[�9J��Uy����hc�1�X�s�k+�^r߰X���'[I�k��ɴk�q=�]|��C@�uu1i�;1;W: �w[��k�^+��^���q��)u�`~pE���Z�����������./�m����c�M0�P�UO��4A�����p����kz���`��DC�����\��#*j�y�;o�R湼x�����t3�Y���e	&����2Q��l�!�E�ت����H��'���r���ذaJ�>-��f�5q��SLҾ���-�(߹_8�=�;�oT���&c��J�@m���J�R�?Y�$�K�P-c��~��ֹ־��4��˟)\A_F�YZ'�mc!UN�ᚘ/�<?��q �vӹ�OuM��S��D�B�z��X0�?���x��c�^�V0t��}w<��ڠ��ehۊ��w:�ʢʅ��S E�聘��c���Ǣ3���8Y�����v�ș@����m�We�>�;�I���+�t<�aJ�;�۰�d8t��t��M�pG�!����2��<��4M�����i��tj���j�DG��Wb?Q|+;g!j�w�:�@�o�3y2<�o5�ׄ�$�Ry�ĥ܉�9Ƕ�rV����2�Lwtz�q|_+��3�ȑ�p�����Oc��t��5�aLj��԰)Z\E��"��F�M�P���ߓLyPZ���-'��b.K)��Ys���8��XK�8p��g��LVY�s
��I��Q�M<�`���fKc��5о�"�����%����d�ڡYдz���ֆ���1Y:��X'�(-��æg��o�l^�ubJ�"#*���wIp`��°�&Q��L������`���|��L����7o���ܓ�۔�gsP�xf�l�v-������\/�I֐M��V�U��)J"�m�<��ʑ�d���G��g	�Q7W���[\�3�eO�|�YO�ޱ�w�2���o��0����"�Ϸ�SEI�q��B�R5��|�p�	q��Z+�x���E1H�ϫ.��$�'+��Ӳ�ͫ��2��Żl���Iq���K$�:w��L���N����͆��LU�����)�I��'؊����]�X\5�����I(�P��Rq4-;��'��2�j�"DD|E���e;sY�qy��#̀��][���/־|�cGK[q�t���Q��9:^���V
�a�YUd�0�h����UF���L} hLҝ���b���T�����������"W�I�yt5�ŵH/3�T�-��PCՙ�$�D��6�Dy�`�����~�[����}�msj�oHW�gqZ)�(���A���T���1'wL���BK��I|��$B�Zdě=�T����f�;�&�`>�}�oL~��s�9�I\K6�2����>�����MUQ0\ឨGp�uw��R���Na��m�J�q섍������Q�=}��@�o�k��0.�H��:>a6�:ݹvs /
f��.5_U�~W�
n����M��"p͞��uⴰp.&�m�n���ʔv�%�̡!E�D9���C�w�_0�s��'x��&Q����K�;����t��R�5����-�Vo�a�t+��>`�Qzo6�n�(!�/�uV�(g��mIUt��.JPoKM �%3��5�
����}��eM �~���mZ�o�����I����A`j]/��=c���9(Q�lWZN�{$�3�Ӊ.:�Ii ���o�XF����#I�8�oT>�"Z?��#M
/����� ���s������b=:�C����5�b)���idd�KJ[�POR�g?��	�<+�����^U�5�M�s4�<�J'�YvZ'g��~�6�z�ǚ��B��ݤ��w�,��ЭHd�_jn=��,���I��U��w�9U	C��yG4� U�\���^q�t%4�d\���i�/�c�����Q&.��y�T	�}���\P{�i��Mm%