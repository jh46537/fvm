��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���Ⓞ,B�$t�{����c�,�-��� k�4�	��[%��B�?���4��\�@e-��� ���u����'᣸߬Hӣmy� q�`L�S�L��-|�,���Ξ�<j�����̨O��f��U�,ﭵ�h���voҭOu���[�)n�g*k�<l��p�l�O
����1�e"��MT����t���*��<�i�Awd�;����ECF�ZC8��&屹_|��vlj�k�G3�*�萜�(:L
�>3���v�L&��p4pt9y�%o:b��A�f�����
@hQ6yP$�Q�f���{��R�e�5!�d᭟��7+UZ,���!��I�= ȑ���C˥rό�I�iy���3�V~/�N�6!�74@-q�^6�& �shn�'J|�#"����,�[����	�ε�Q]�ł�[���	8�m�}0��Gi�=mc�W�N�#��%���"���z��0��2C�Q�L���f�.���,`	�߻�ke�P����zhD���P� ��v��Gͪ��t!e�ι�`�w�Gܐ�bPƓl� HU5Β|��A���׋vdgyeˏ@����s7=���3�#�~5�[ߗGI�H�c}���of���l ,���f�sDfI��x�}�sӕ��j��0a�FјZ|��ִj�L觘�Oއ�q��̈́�N�y��)e%i�s2�qNSȷH
pu�!C@��R�8�7�7@n�1����������#Z�9���8@V��nF?�>s;`�3�&�3�T���춦w��h�Sł�mØk� ��T�s�W��~�.�X��L/'l���h�+@�G�W{ŏ�a_I��đ=f�;��&[��֞@��(er��Źɮ��ʰ!~}�	�41�2��g_R���&ki~+g_��$qxQ�>� �7__Ɍ�B׋�+1��-�=�����L]�E�$�r臨�(��.����=�`"+���m�pi�{H�$��0z3�+$ܔh�\��@Ȍ'S޿2krѻ'+�`��M���>l/��������/H�v'�o�����8�~>%ⳍrp5~��̯�;HQ�Z�@����)c�7�j>���h�G%`%�7���щ�+��1̢�����P <�"mOCW+�UJ�ʓ�K��&��m�6����2	�����D��]���hr/Z�B���FBgy�p�%��z��S��S�]�.�A�V҆�2��1��ވ���1�����1 &�g�2�T�~��n$�������96Od.��\)�(-FX���2V�U��7�_m8)�%=�]�{G���N�p���@И���{�l���M�a#!&}���ޔ}S,=��oN��4��\2h>"������;�>Z��w�B�S�;:g@��E�5��2���⃏�����e��̞rTS�l�A}aB�� �mO�o�G�_�Se�{�Mu��|��4�Ά􏰘�����R�>�3apf��/�ݦw+���"ȣ+� ���?+8Iũl'<`L�Ql+�T�F��A��^=��J��������$���Ԏ|�U��xF���Se� �_�5J��㸚a�4�}&�zߔ�b��i'Cz< �_\����t�C6�'���щ�9̇L8F�{>�$[�j������Ȳ��:z��&��{�= �.4/��t%�̙�2*��*�߅./��nD*�U' ����p
�H��މD7�,�~�}�8���ũ� ��nV�to;'��� �����~4
ϐ�,&!E�������^s�U���}�N�aD�@���D��oR��0�N����-6����=~����n��?��(~>z�9�[����0ڃ;7�^�[�|�]}ҁR�,���J��� �r4�wL�l�]Wn�cM������n����]-����u�d�m��䏎��$[U����a,b�Ẁ7_Jw�%v�X�d�!wB�+8��#|�0�-!������̀V#/'A�����W+2��%pß��� �!�&*c��v�Nls����сz&i���޸ ���:[&��M��Gn���Ӛ1�&�*S��ڦ�M�|{�Ԣ��� v�p.=��̖����Z|���r�@N��7� G���<��/��%�B5�L���~��m��o�#%:��g7W,@�!d�t��)>��p�	Dz��b����s���Fl�މ����4�nO�笄�=����Q ?��BI��|3�άp�dc���g)�t����%�>�'�gHO���g 40ɧ�� ��M^�D������@��O�{�#���.e�����G>��t2p97�D�+�0[������u�!��E�i3��)E�:i೉k]�$"�h�x���}�uu�/�����mB���K6��=���ᝩ")��+ M��v�h�ů�I�N]+y�q�?�9D��2[��Xpt�����Ќ��D��m��%g.?��ؗ���:�`e�6�N@m��b����4Ѭ>Ole�CvTG$.4�Îg�/,@Te_��Kctd��
��%��t�y!��B�^��a.)n�� ]�C� �:xZ��1Y&|T@J�O�dU1���Ixv�@G�,��7�dX�cǓW��h�]�ZONAұC,ۇ҆����k_n#����=p�Z���x�����y��r�I�6T:ޫ������c�n��_*ĎdHD�u	��0��`��WF� Q��C�H����9X)��s{���\z�T����"���Y�4BCv^�O��pu�dx���U�b��Nv��{L8���Qgh������5֌�5\�I!��ݢ\#�3��������>���vl��5V�Kǉ�{�v���{�A`C%(���qm�][�"���3U �6�@dڿ5��Z��h�LT"��R�Q��(�~xK��#֬��]ܺ6P�� �[<�,����=ǚ���vo^)4ԮzC0\��<GRI�p��BVl���,�F#��k~ƞ'��X����k�V�N��x���i!��ҩ�-򇲓� ��%f�v
r�j?�L�8�,F��#���t�T0�s���@T߸�r>Kj���1,��H�dK߬՗7�VL��:����r)��!C���ѓ\�|���@lۖ
M$Y�%D&I�r���DL⛜w��ׄ�u���Y�YC-<�I��#,r�q�h�d�]9��"�{iW�8�xb��4}�)��Fm�S��~��	䃲n�d_��d���}���b�m��i[�t�8������-ǣﶺ�E㍎\���ʾ��>����e͙�ӊ��D�
��*_�X2 _���w5B��ն(#"F@X���u9�h����e���B�Q�����s$�~5�N�&؇PQC�aҺ_�5����;Cu�����v�_TK$=����y�U���K��Y^�QN&M}��P�ƪL�1�<<���'TZ��RR������;���f^YQ�cꌔ����?s�D� gf�4��n��*����*Ngmܿ�&U��%�NE���^
�{Ir���9���;.p���pK߰e\=N,��ǒ4�Hp�XMc�����_�N�i�����=���8��G�{�;��=(��jK���b|+��ە��tt�"��	cE�"��{d*�_��4f�t�L��oK����!�k$�K��t�]�s�E�rsX(�����3r�B2eZ�3�oc2�rVe(s��f�H~�E�5�W\���MG$�F��VjIb�\^�������4ɝ��8D��w>zk� &��]~c�2@�qv7���jhy��S�0�<7zɂd��Mlq��v�#q�z}�.C`m�~y\���$S��l�����W��M�����u޷w~fx�߽3]�ԗ��y��k����~ӡ���}|����Z�å&����`,:TD{����0K���ҭ�i��Ѡ�S:
�u���:�V�k�g<o�˪��Fru9��J%�<>�,��	c��-�Nd���|��813�^Y�//˨��H ���r��6�.�m���-E�9!�~)�ߍ@y�/��VB|H��UN���0\�SY4G������]:P�,��e�C�Y����ڼ�))�9]��,±�[h�U
�8��m)�$�Dҹ��;.�l���As�Jϭ�3٦q0,�ɒ8�;ݐ�M�F7��B�c�V����i,%r�*^k9�Al��x�̮ڞ9jj�������:���˴p�>���A�h��'�Ze^2��"��ʐ#�:[��@�S0�K�������<y
ܑ�5����-�M�3�0��g�N��%� z�J��w�bs�T<��zá��Q��?S�7�/ؚ�ߨָ����X�[��	nq�x�@R���Ŧh29@�u;�����2`��|}�IH��ہ.N���h��o�����9��h�Z�(�㩷��Lq-�_nS��|7���)���W�T��·�4���.�-��\��Y��+��Ր��r��mh+rT�}���h�l��{�&�Y��n9�({�cC?��`�7�"ڕY��DF18���[J��N/�,�/,`�a� NKSY�����8�i�5�a���)�v���/��:�)�ZQ�wx|�����zP�6!`��۟�O�i�t��"�`��i~R�a�r�:�8�R�uZ�JB�;���b���Vb�8=�ѽ ̥�����0������D3Ʊ2����^�Ӻ��Y+3 �E=�3r[��o�-�j�|Gx��E�LP�P���ٛM� ��p(ز)��F� �����������O���&V��g��,�J#-���$��ب�ὢ�VUm8�����wg�!��q�hx��jA/�
�a�,@��0{n���cj·����v:�@..VX@GK�Dcà<�f��Ox���SL"1c�i61@����AH5(���� ��s$�g�	�?��2�������!u	�wk���>�K����t���[�8���X�M]�.%B��]�4$�\�֏�T�
��irб��ℂ��~�	�2��Y,��:�i��H�/�_��3������*�No�d�B#P�Q�Q����e
h�>!��iƟa�W�Nv��糸�`]��?ъ���8>U��?|�7[�l(�<�'{�Ν���ʨY_/8c�y��YQ^4��4���s�9��F�V�����8��;(�tBF���U�1K@�شki	DV�_B�'<�_�ff��k����t�_1��[j��D	���I�%(�>�mX�҃�azM��9c� =���)�y_C<b�G���V��H��L�~���?��o�>\
G.���;�Q�E T��#8��/B6EQ�9b�AK8���]j'%��(L��CF�abcb��xL�f�mIG�R�;����ն��������a�s}�nL�	F�����R������ �Ŏ�;��Q��Ĥ�q�°V��v��u�}gП�?�]��X���;� -jn�Q�'�"e�R��ۀ�/�I��tC�]N�0��l���K<�%��#sT��������2r���1��1d�》��Zg��]Z\?Ȅ��sP�uyӟ�q�m��r֙ꢚ���bO|W���Ї��3G��vI�5ʜ(w�	�h����fs2�q�t}S>�����]@��dH�,��,��Ub��+ޡ���g&t4���*�\�&�����Za�aH����?-ɫLI!�E��_C�y�5�����QͣzrÂ�<�s:�nU�����{e�����_+�����~�U9`���Ո�Ty�PE1�~��'�� �����i�*�h{}��������دi43:ig�l�Ri��E��p�\�Y3�f��\����� �(���&�1	]�uo�/�k$��A�2����5���6kl��a�.m��S���:�
=R^u���-JX,�-�7�l[K�߂�aR9p�40��<���y��T����FrH��l�)xђ��[�Ǎ�d��Da�ԯ,*�y�|em?�ZQ�?䒄��_$��(�AK�C����L1���4��`,B��f�.��=�ܸ4kx���Ꮲ}r�O �y�_�b6���x�p�&�)rHi3�[G�-�T�Th���hQ�b���Y[�cp�+�I �Ð4��A���IĭuL��կ-WQ�P�	�j&D�Ū������(�a��"����ׁ{�m�L,�X����KV$�H��:�ܸ+I6���I�C|kq�s�}&!5p�e�x��,%+�G�%q����1�h�Q���u���3.��:�Zm�i9,�T�g��P����]��m^;Mğ�m�#m-Z�g�����`�����J�O�s1�E����L�
�[E������x:-#J��o���gT�>��ϗ���������I�����HH;�|z��o����[2���ݳ$�u�izJ����bs<F�ԋFU&J�d���))2��)U;Y�����,��"eAA�"2ce=��OQ�d́W˭���Z,�dR$�$�$0a�w`�y��\�͡7Pk�T%��,�h���YHJ$�%�ˣM'�W�B��t7�W@���^��/G��(��~�Ns� /�F?��פ����5u�ߒ�v�#%�7�b���-��A�y&g�Ũ�y�^M���|�|/byO��c5ï�}֫������� {	t���\Ŕ��M�WΏD��y���9�̔�.q/Ab	��<ʴڇV�������3��%�pk���I5����q m~�2����	�^0@�s�E�O���n��2&z�C*�&A4���o �E_d��h⏁q�A"��0Qa�A�S�W	1e�A��LB.���?QaɐCI�ܑir��v O$M��6
��I���J1���YS�:^�<��'���!v���ÇD�F��R��_̕1�6�Y_y�,���c��,�y�`�@����b>o����j����q��~�M�V�B�*�F>L�v�d?G`�X���ߊ'��/�RX�UᣇL���,d����Ȉ����@wΰ|-�J'���'�y���������B�X�MTx�M����^m��10�5�;u���� �3�pA�����dh-��	_�M�2���;츋_1b��[�=/c�b��
(F�s5�'^J�Ya��B���l7��T��1�mǶ�)���Y�eٚ��䁘,Fs}Q�i)\��l�r�u!'�wB�	�Z�b��/��m��70F��:��l�<�"�v/"���ƺ,��@�� ���(����?E�.�0�N�Y+�8�g"�`�
;o�@��Nc�:��J�K�=��K��<�!�H�w�Ȼ��c�'Ϋ!n$�����m�c]#�����<�g�U{�W�+�ĺl1î`]�!q9>�20�by7�@�հ�c�h�DR|���b��u}�n���K+�ͪ/o����tBI�ĩ��?(l�rۼ:�@�&a�O�ۛ�Q��m�SÄ�+�򜌳+^�[��3O8}9A��&�|]=\m��7�����|@/AxN1ꬷ�7�0�o�J_,���"�͟�1���grA��g����Ib~>�����t,ХϯY!i����wyAɓ�8�#cЪ��h�.�
���)��+B����	ۓ8lt�s��̼�
Ps�	�?�}��"������ ��������R�pn�w|b�|.~gi���P.{1T7L�渋���Zj�j���'�9�5�g��?�ꪃD�Hs�/Zd�ai��~�A1s���]�� t����;��nޡ"�A�a�#;=�@����
�G��jC�M-��b,m^�����3j�st:�l<C
�J�d���l�4u9��3~C--�y��U�RacV���	}cz_/q�O�����}��̥�$�nx�c����ȣ��f�u:���U>r�į~Lf�M����,	e��{D��.��/<I������u������ۥ��&�j���8:��Lh ���A7�\�՘^�|��.O�뉲݅mpMB���5�t������ �B��-OD8��\�?��țn!�堓����u�8��>D���*`~]B��\m��/�_���$��/� ��#��n9�8m��P�g�`�y�N0�^���]��L��"�rl��)�o�yI$OT��V���9��:V��gSR�V�4�����L0bA.+(����,��d�6l�~SKe���b�����wrF#*�H�J����c��g��(�v8��c�9��s��w�̽�o���Oa�t�"1t���'z������:��4>�7C7;ϗ��G�u�L#�e��
2E�!clvE��޹��q�u��>J�k���'�{k�/�l��DRR&��� �5�"��;?cS�$s�����=�t�5����N,�D���W{�#�Q��8}��+p���!�.!��������Ȫ�U��6�+�(���N�UQ��g���v� �;�8�˴W���:\��"I�`����8����ݹ$��s0�@ʆ�%GU%'?�X��/�ȟ#�Eyb�K��^�j�7���Awhi4�*r[f�l�vu�:Q�}DS��fR@\�6n����+�	���%�*.��T^e��m�(��M6�p�f��a6{��xl~ɪw��`+���S,�����`�
�u��������D�6�T�'���b}�7T�Њ�A`�,pv�FQK��oA��v�8y��e�-������+���ru��7�0�`��H����Y�֋�4s���ҩ����� ���3
Ҫ_��q�.����qJZ�Iڔ�1�bC� pu'<i�Mʔ��d�/J~~����G*f�������+������b�G[��$�:xx�E9�Dp�Hc5�Xj>w�1��/#���(s����X-N�Vg���r�5_{��L'�tD�;9��6���|����]+�Z������-c��'ox.8�^.�&�-IUr��>�:ĉ�1(�#�R�yz5`�%�a�Ԧq���� {���F��7Wt�^7���� ?��wqva$������4$�,��A$l��:�rP�c�b�6q�U�Z��A��<<�IpeܱW_�ɻ���A��KK���)ɓt4iWw�lY����{�������IĐGm��]�M��Zv�s��O>����>�����%�&O֯�]�V6 ]A�ש�DD��AH�����O>!$�цxk�k�Sݸ��0Ǚ��^��g�����W�mYZ�z�iLQKWn�c�o1N�7�7����o�5AjdX���d��a^����%����?Y �
�q������@������& d{E �I�#;��0hSތ�������#0$4�����M�C816�W1��R��'�M�(�Yu�����,'?a��ٻD=��p�5��?J}��QǤ�BP�����T��䇔�I%B����W�3���b�e���#�:�a�n�40�~���?�����~���ߊ��{�2�Б�Y%���m$i��$ =h��-7[}�Sf�'N���0��Gb�dN��%�a�g�����G�l����Y��(���Ag�%���y���K�ǛpC�yk�:���Z���?��%Y����I�����I2��B���^4��u)oAw����EԷ*.� �s�+���C�s�WLT� 7��x@E!B�������N�f���N�HVJ���3Up�gƂ[�QP��Y�3*6�i�ӥ��d�'�@�j~f܎�}v/�����M����
w�-T�f��{/�V�ʎ���:��k���/���D�u�����

[���[�XD�x[��H�I��z�0��%�mr��#��ߦpt���Q��z��	Udg&Ay��7�}���~�v��̇p��!đ��|k_9aze�(�(sK.��;��X�A`5��2�߻qP�џ� *	+_��Q�~������}5���>�@A���dl��-M��,�+Hѥ5-0&����+z������þC�q�xΪ��^���"2R��u�J"��4�����hk)�����F�,rw�R-#'��ʸ�������o��m��'�&	6=�lyH�6F��(m*Q����a�ٳ�H�nI�|�T9{�֨b�.Jo)�͆�������y�+�D�� F�N��>hD�&��%��<�\�t��6�C B��?��0�ڗ%��8������|��SKA�����N��{�=�(\� 
��;�n������Na�!�>L��
.�����5��p+�ʁ�4��gy$�S��#�y&ش�.6݂_�~X��M���7l����$�&�	��P_�
@�gH�7��1�b�Du�S:��%��}1)�(�tf�<Yhl�B�m"�V~/�_(}s蛲���y����n����V�Q���8-�Ĝ�7����*��
撍�g�QY�r':��5P��TL"���{v�;33ZTW9�a #�]�J��z��
mF�t�������%�p�-nn/-mB*S0w�ĤAU�_��R2S7�8��[[{��C���h3�L�!��O~1l�~�t� F�Fź<
a��lۡm��6��7k(H�;{���jx1� �������Q[�����v�s��|�t�jg}?X���+��D�Y�Z��#�4�H¥��5�_��O����r��C����CU��9Eu��ѯz�.	�jz�N�[��]`_?�����6*bj�!N	�����E�g�f}�*G���8����(��΂����ו6�*ƕ���A0*�p�3���(M�,�|�y>��}�5{f�t�/��Xf��ko7$�>-��ĥ�ך�i^���|&�ro]��W�1AHf�h�0]�2QJ�!g�.���FP,�P��ǒ^%����3#G���� �:,;�h��(�o�Y���3(��0��v�ƌ����)����R$ʎ{��uʉL�Y��_�?�]]�&��ࡳkV8���@oJo`���Db�ʊ\����0��f/3���	>.�ɷ��]:�66��V�>��:����G�CNXD����O���+�N�I��I:}Y�!�OT,���p�o�r���GMυ�f�LSq=��1���R�3��z�A�N��Xu�i���g�w��BU�ۃ`�����@>����� ��y�A��2sp��s_�O�c�b N�c����\H"��2FG���ӣ1TΆ:	n!�!�4!1��W5�4nQ��g0BO���n7���c�HI]	��i��cN���p��`em�c*j=�-j ̃���H�U�ɰrNkp#*������'�SȚ{Y�͒����p���8읛g�C7�i� �����]�}WoD��+��˺3�m�^_9�>��h����-*(~�X����V�2��ml����sg��f#w)�CM[�HLK<�4%��q�rQ����0�ё����y�m�Tv�$I��b>*�}4�R��2[�"��:�~����W��>:K�U��/�LϘ��� ��x_&P�G�y�`[_�� �g|�&�ݽr���e�G�Th��8'2����|��Ӻ�V����
�I����D-)-���a,tEӕ�kS]Z=\3z�>�q���N�'rϊHAS���KP��V��z�/\-͌c "�I��gU���1�ʣ��;A�q����4c6�S�s���v'��#�c(��YI��H�܁=N�SI|��}�%�p5Ɔ��.�hU
:j�!�s5�����-[����c#y��ǩ�#��1a8d�h	�����aW�g��8ᨭ�
)��r,]"�~= �@��a��⺇�f�~\5²�	ū:����Џ���6De�G�Nm�҄x(��Z);?���6�}���ʯ��U�\:Z��p�3IW=���Ȥ��l<��� ���4�=��H�c�'L1�zw4E���ݴ�K�u���1�_^�hbkT`�wƚ{��ٜ'����[T.q�]^dQ�)��>ۆAH���iָ
 aS������W����U�a�:������N�G��ԏZ�Q�U�rP. �Mo���w��������E$3&��D)c%^�8}"&r�y��!�"�����?�퉛����6��ik}�� �׼7��K�;��fY�V��_��o��8�=���!�@�����@�ӝI��v��ۀ�����;�E���ĩ���=�E�{�N�ZX#LY����j�/�Pz�)��� Ȼ_��KV��C�uK���-�R�6����]��Hm6K���U��sK�Vͪ}�I��N������fO=��_���Q�aQn8Cx-�<���f@�a8_��:/�
����|���"�<�&t�í�i��\=>�=�5� �/�r7fg
���D���F��	No���\���i��.@��(V���R;��X �]0m�j<ZR����6�:Ȓ��+K���l���7p(�R#��'�1ԫ�ft"=�]̷���:�S
þ�fg�e��Ix�rB&�۾�*&��W~��PX^s;פ�9U[��kԦ{�J�k�>�
zeیZ�R�m>l?`!��ҁ������.f�>LyF-:�����������`��i_c܆˝�>�@�t�ó�,��I�P�J,�m�ƌ*�O8�H��a�>�YO%N\�C�f����0�d��VU�i�ؕ�r����.F�v���N�X�B?$L���-����[��n�X$@������f_�a��>�5��������(f�����0۵�� ��A���՟XqOگL=��'ƣ$>����
Hw�ʽ���µ����
,�6�r�֖p����W�u�,#���y}Υ���M�V��8�6D���L�Rv�¸Ӎ��!���0E�i睟��/T=���$�A�L<_wRߤaL��!
~Ô6	FTm��Ν�Mqg1"��q9̯Tc	3�/�����$����j��f�i�A��JA-��T��E����eH�����w�������R���a_��j2�`�]�i3���n�Bd7����6���K-@��%��X���r?�PB�t���\O�{�:7&�0=�G�څ��]o�}9�&�	w��1���?%�#�P|�Qd�1�|rQ4*Gz3�޴�g����a��M�k�;lo���(��Lİ�H��z��^���p0�a6�EZ}�����|Ҭ�x�9;��n�T�u���e�����[fs�̏���S��:��� J���'#DE��ƩOAO��g�p#�Ư���_:���	ɍrV�[P0�?{k� � �VC�d�xН�Dr������X5ΠH�͉5-2��	�#����u����'�IAoV5������C�>t�n_l�B*�k�C�pE��GH5	Ĝ4���W�_܀�A��t=L�y�WV(Fɭ�>��<9��dk'�{�8U)�����Z�Ȭͽ�
Gr���w������L��H����1�7��5F�+�K2�F�-�����\��7M�^"_��V��[�j�S-w�K�]+�e�w�����>��`��j��Ʈy *��,�<�$)�%����\PtAG�9h��֚V��ִy�}�=�S����L�]?:��;:�|��h����M;\�?�a���l$:F��8����Zsd�<bU���CLP<���Sq��( �$�#,�����X@X6ll!+E�1�jc����Qe�)�'��[ΗQ�c|� ��9����{��*?s,�m[?�GD����7-�i�\4��"�;��^��+H�K8�lu諆�P�G.Aa�j���I��H󨶺�I[#�hrh{v���$ �s�i��
���n���j��gT8:	�����<�x#ȇ41�U��y�`�= ؞�ԏ,$Y����Q���X�E�M+e����؅�AY�`Z��V�I���H;KӰ�x�%w�^̀�6"jDG��}��fI�r����i�[�l��DW��L�v��3����u+�&���-�/:�Y�/�5�fI��Ll+�w$T���d��l3��!(�NJ��6M&�"%%��KEW[����}��8@f����	���0,���|@�>���~�`tǔםH�C�끐�q��W�Yߍ�}}-�X���}sDaw�34G7�ƭ�o��.�Y�M���j�ԃ,C����������8@r�Zwuۍ�ܮ��V� A;��o^��R#�잩��Q)l�������ڳ�<����&c�-{R�K ֻݼ�����ŞźT��^G+8��w:�7���p�c�.�k�����.D0N,��k��Ln��=܎(��i����*��[ZXڳZh�]7�^C{H����ZOl9�wo`j�������ķ�kӮ��� )�@֟�n����	�y�ׁ�JX�K6�#d�<!$]��ֵ.�B����H��"�F���
��c��h���z
*��W��/(.�b]��&���3�*7W����O2�>
|r�� �4�9���g):�U0(G�����) 	�C�ɴE6������h��Η�������wJc��_8L��jE*�?�1	�w�ٸ����n�(�`.���}a\���H�u��z'ד�3��q'�ԏ���v\��!��㗀޶?���mM���Q|��V\I5�)̐2��߬\v;W�l�^���ɰ�e=�5�^�IS�M�t����c�|�A�|�t\$����\���ZT��_`痃Q��(�y� �-0AT�*Y�ᱣc\f��}��� י�[h76�]Ct�@ut�(�X[�"m�ʴ���0�n�gU�Z�q����hIdt���_���&�������T2�����LB�ϰɁ3{���!����H�>7-R�9��7{�lG�`�U��u���~�R+��r�w�@=��������7�����`oc���bt9�� rA��|�t����ȜR\�K��L�`]f�ź�h�dp�FXK��,O���q��Z��ş�s��n�;�?�Y���؇m
H�\��������Y�t���
�5�1�V�To#]P���	��xF���h��ֺAW�,Ŭ:�5����Hdn��w+F����T)J��N�?v�ia�t`b�{��4�5�r�h#|�J{��f\>���|]�CZG�I�o�@g�N8�|swE+z(qʙܷ�|1-#��iD790ҿ�����=�L�n����	q�*Ue�̖k����y��P�SdM��C`S�\`��	~A�w8�q�F��A&�t'�t��>�)�h=#�#U)��P,�4�P�5��,���-�c�.�U0�<�ߣ���� ͜�f����bb_��3p�RG��ka^8����*e�}�� W�i{7d����R�8�#}�uU��n�i�l���::	�_8!N�K�{8�������&P G��-*��hg^�4]�s.,疂b[@I��$%� ���k��t9�ީB�J�~�<��Iw0%�v�{E�ll0�����aU���s~���W��mN'&�~�Ћr�	ac\T�A$���j�Se���ƂI��ILE�%�ڜq�;2�	cg\~�BY�EF�J�=/�l��M�íW�P�2r���4�-n7�\Gc�Qrb�qY�NR�QTHbB��l�.hZFn��B�Db'�m�E8�9A\H�wa<k(9&�	�=1i�a�6,Ň��|�@�ǒ\��Y�$v��h৸0L����M�U�n����xE�ИJp���A���� �j�3�UV|��zܗ����2Ɖ�sB�.e}���k�кF�j�.Z�E٬'�r�^ ���q�������240ȝA�(4"�th�:�I�l�+�M�2抂c�.`����nW]*% �+s�@���COj`�c�0���pP����W T�B=<��Xdb�-��$��E	xX��˯���ktL��k2���L��ֈڎ�Wq��2��"�=�O�O"!����
P�a�EFM�r�������pqMGȯ�R-v�b�1� <Q �'��RH��A5Jv�g\��x�˟((D�_wR�� g�VF5�`>�mA�����f'<�P>����b��׋��j�0��wb���Ձ)�j��r,����x'0���;�&h�,[$�f��Ȑ �P����v�� +/��_ہ��z.�ԑ����C��pٰu����OI�ehk����6ӚK$��j�j�>cn�d3D�,4�w��R2�absP��R�3��j�rzI�_���Fy�������B1��S$n�)R(ȷ���]�����B"3}m¹���#p�����`��6m5J�:׺l6G�h��ި�tنq<�p`q��/�&Ƕ�ؘ1݊��h��E��ߙ�G٭H�,u��`���e=lX��AZ\t�1y|��#8&��(~�p��Q��}�2뛭���Q:7ŭ�����\�.�Jπc�ŅH�}g�N2�
�!a:"Ֆ,�)�g+eI��#:������"3���ZG�2ֶ�"c����5b��Խ�e� a�ѯ�|3��E�%���v!�g�ڗF���%�NQ�6�V/I�5���{����#2�(�dFf�O:� �9Q��������^1��%��L:��@��W��ǌ*�,q��H���x9�_$�*1��ȒB��W����?�5
̉�`2TPdo>�7>MM���>Xl/� w\&e�oVjw�!�l10����|�CثѰ���2H�E�
.�5�=�y�7�V�MUs��%�ӿ��cmI����A�������w�[ �k-tE;3R,W��}�Ni3s��gW��d��{�I"x�% ��:F!d�W�A����j�WP�n�^ �R��]2��q�js�1}���s3oi#bL��)4�4�ј�$��3�􏫶��y��L��&�6ݤ͹��t�J���Q+p�ͧ�`H��>]�8
faxٛ��S�-cQ���I�[n�9?�7��|e�Q[U���٘|�`����O�|��PՌNv%a0��%-j��=l��E���oC�b�Z�������.�P�=}�lט �vs�Tc%���vE9�=�xg�\m!��?`1�f���ݺ�p�^���i��_&1}[k,0*Wǽ�o��R��Be[.)�`�����<��q�rŷ�A��o�&R�]Jz}z�̠U�v3bw%��h���vT�(��hl}�@��
��)$�)���<K�\{��p�����VH��`k��'HC����;��뵍���Er��b@��p�����kF��
���m����?ŢW6DWM���H��Q	��-��[J�l�l����;T�{K�����@Yr��%��yF�U������+>�2��K]�F��Ҿ����\�58x0w��<�T�T�x'�C���w���м(C��V�
�!R4N�����%A����8��DxE��n�c���[B�ϽBb	�n�A͌�I��&&H��go����V����Q���2�5C.�f�e)��M'Çv�����Q���ڭ��KNs�;Y�@�Ǥ&�,&�pp�N�4�--"pe/�'}0��h�	6�6^�]ƘbƢ�%�(Ty�,���>u�4�g�p���S_�d;�E�^�%���u�T\�Ni�C6���k���X�kͶ��Z� A��.�����i����8��m�@I��Q���$�ɔ���U3���!L~�Qƅ��z'��$i������6���Hw�ڈ�O�أ�)W��d^��|y ���ۇד�),(�ʀ�>?��X�Yp�v���0>{��q���6tg=�^�	�����>6��2�f����t���&�?5ADN��`��xI��j��WD��r:ynM+d��i/1�\�Ǡ�"�?��ڪ�v�n�b��ax��l����N)��ͅ�p0щ�8�{����y�u"evő���2R�I�m/���TU�B������ik��hi_�N�d�R��Y�7�I�&s�z�@��NR�Q�e	�y��,e�}$O�z�|��Z�R�4�eʴ��p��N֧ d���޼�B�	�J��/�~�Q4uFԌ=����� �)Z�|��t���B�s7�6��^6�Џ�{�vjO���Q?w ����V�j�ߎ@"�x�w���$�L�F� !��˧�B����%�����Iy[��sT�ô�K~���4d�C�O��$ݚ:�\6�Ў��jQ��G��4���z,P&�=O3�U����Hf6+J�-��/t���51Q��rTp6���y���uF�]hӊS�X�a�H+؇��T#I�(�S+l���,����U�Qu�Mx�^���́�֨��z�zV)�smhǡCP�^'��j!5��g��v;Ȉ��]E�dV�(~=��Ƞ��"��X�#w��Gr���B̓Nt~���>�ɫz�c���II�zt�K����;7�����]��Ζw��{�5����r������%����/k�T��7�����<�2L��_��m����x�j�)����[����P�<�T���`7��0[i�q�ltK��WΓE�Ե��sy���:aǲ��y��ap^�5)iP*V��7Z�nԩ��ě�v�~�������� �����)�Ф�+�@x���M����G�*���0�O�
d�d����ƙ�0's2+�G��s],i3���fJ�į�a�m�b>7��֯4+~��m8L��o�_`�'��B^Ft���p�[�N݀�\v;xV�!�Mt"2o��*���Qխ�Y�U��a�7�յ�sE8�vGА ��e�(�/����<�G�����