// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XDGDRszr+IkEv8jzxaWE3NmJ2zrpnXM/vrTNFBdd2F8tLq0HI3gGtxnscVSn3x25
t65NrLZ5EimR4pUAE2wT9TyjvJsTZaQI7tnp2xGyYggkJWwrfhf/8PUMdg0xAcd3
EFk+D5VW3cmyc+OlGC9DmHsIclYR3dZmORi5xEpxRHA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8640)
YMoJ1YrxV1XGXACh0eikcAJ9BSCeoxqa6RcyJ2wFyb97m++knZwOLw7DXMSPZXSx
EXw7Q4G0xk/eDBPeK3Vqr6pdnvR4w1dOvStV1Fxlf66ujBpzOdq9D64lbPc3uMfK
SwHlDgqAF01/LD0DrjupZmCpzSlO2nDVZe7QLXyOOddkbIEUtDHIZdeXTCXG4yGk
800yKi4eowI59hzcR/r/qi1sQE0DCrajR1ZG01iPJLUugFT+9FDXod4gQHbqs5ef
HInlOYgqetmR+Qjun+6XHR3hwGpZefoo/+5qvzJs0kQSkAyhv4qG5DLfHlc72O/u
aA5tZm57vjiNMnRWSVU/8yuE+yQj1JwUgAede04meTJ3D0FxMzgmbQ6jQfjOdxhm
AzSogZ7ESLm/D2pBm0DGh4f6Xm5UabQE7Yy+PqPMV0MgpTIl+F1gSCYCjueyYAjV
KRAjd5R2gJ22fkeNpHqID4N04cIEh0h0Y83bhAr00vHPYar6wMELAH/zBQLCpliI
RaJnyRmCKwfYr4qP7L86xyulgVYnAOE3+Big8nAe0IiyXn6itgHV6xzfTb4tk5/g
EuK8u7nfMviHQQbcJc4vsexaX7gilEuBIfvAWuMC/9ExcKa4udK8k7j/LpE94wSx
hc+bmsSAOwMZxOJyIvIVzxGw92hFW7fn2F3DQjQQshuprF/zMpQkHrQpjW3cKt+S
VMt/mUB1cmXM4TUmQVFyfbTzrmfGuS+eW8zmHbbWnsMSPuaPGFC4tRo7KLF2Z1FE
eAV3NSgLD38MyqPL5zQoEHOJ6bfe/JtNzMZ4XO7tHxGcU0Fmi7aTxuWnYEJXHFr5
Fp9wqkNMSngKgfzwim+xadSGUPYiIhHXLMlZPGpMazR968YeS6QQ2zOgI6GNfsFN
3fHhWpUofKkevOcK3r6HIFvjdVViR6WcEhQLGKqOb/OKxOQ/rbdT4SVwrgE0NseS
NIuJtHX8ti6xubTqBLmuZwEK+/LwrWUJSqFDlmpICaDMtmFuLWxs5/baCE2jolBK
wea8UxNvlLF5VYEApa87wNh/k0OHr/06Icdw3ysLkBOguD+jrPaw/51a/ctA/afs
bm79+5mgmiy8yYQ211gbK6HcUEwvtwNH6fLvacipRvgb02/v8blUw8N6RTQXDxdk
WiT4J91ra7QilJnI+xBcNLsxqk52gpDmntAgWLsMiEkvxK5JskJ63+hYztvou1qo
rXMT7tnv2rjAi685+VaPRcF/IsaNtS2T2wzXJ4NXiW006u+205c+VZ81h5eIOtMo
ArSq566LQWjXKsJDOoMshS9q1uZvZF55mYsFDu0pzu3R6IKVe4yE8Ul9GNspQN1o
LZFYVwPXJf8H6TXnmEu+WfnPcqL1+OCQiitj2frJ3hLJdEZvrqsqpcU/WruqIHtP
mtUxnQXs1MwcNi91Tm0+hDnhaDnhJ51xVNKSZm7oZJmCXt/RfmpjtfpZLX0F5TPa
n/27lzxjUEWn0Z/G6egwAc8aO/pTxiki4iitT6yThDu6q1EA7L2J8Z5Jog5qmL4n
tENL4yJNW+qxB2R3x+wvpDXB3A6Z5p0xuO2MeH/a5bLrtMhS1F7+37oRNt0qoTUO
YwoU6yEfebNN8NAiLYR/dhL9w4wUR8J933q10iqqoG8Bguxd/fdckOZHqB5aSWF7
EDmRfhHvwDlOetNhisime/UhaExRC/wPUgogBzAuWlsQ0YbLDGvxp/kg6uOsp2+j
cZJCdYQez6XH5vTQdq7NszdlZ2xyv8qbcAAQ9ywoV8QchDnEqgsArmVspjXAkKa5
UHmLqDJZkKvFT/AyGQbwIBkrgDF5rzv3cUajxMx1+ghNC34iK1i24+FPMHwtJJHg
5b9ZBvbS22QZtTxhbAqADUDfQsCOTReVD78n88X0rYOjFT8QqIbeL0yfwfn0eUvN
pePHZ+aS7AyxgQd8CsNDTxqPIX4W+ZCI+lVvW3BSsfqiw1/QIpo4EGcae0jopmHZ
oktQvw56JTc+RA4AKIedUrF2hBz78bLldR+GlGYJyC7ytHfUnuVmnyMEdFMItp0N
1xYCp9Nl+mGOd7weVArtxVr0MoCHW+m2Bn03kmNQ3ZG7BEfY7oiq0f4SKB80vAOB
CLFMNnjKnO6k640rMDdLIv7Mawl36sRBpt9N/rI+Z1FGNM/c9wqOqEHY9E6nlL8A
XaTa/+aQxONL8OGZdNW1xxY7sMsQxEHCLpKRlTHUNdhUr1srLWg4sKsGa9j1xyfa
LxNtcpNtA/TOkJ++Eob0Da7HKs/lesnGTHS4NOV8J4xQOEPua5cE/Nh/Ty43wRDJ
jGEPsaRg1/ajYpl1qwLi7VTGoIShr5VvfgfjpyLBoNl+V7yGrFwqCbQKMtHloqoc
Fg5d/OfKBIN6OkIcctQgJmUBZcPOGTO6/6HB9vMtTRq5w1fyzJj/AxeGr6hL7flx
eTc98KAMB2bL7Xm6l4TWvvzUq92Mu9D/+SRdS6c31C5uLeu3W9dQLB+3brG9mH7x
K1yqHRHOSPyPTnvQ0MFXthqMUuE73uu6A2DCw7BKJ2v3uSJAMRqazpCi/tP9YQoB
SVSYKjqdIHKBzYWWtlva7jGYEKJLcSlnWh+12NudVXIibMX22LGUq63PYnVOTsiz
8nTsBcFWu0w5MFrp0a63R6BdNV7Hnpbzqf2yElRpZQtAGkFhenUYcPtIsT8AuqeU
lcpJ5VZufD28zz4TMQOqR91exzSI7r4IGv1yuJZ6mBcsotDWpa73KzZwJr8kPaJ9
ksfl744pz3TY2XtLiH3D/6KQhIZ44z4TARUaX3dJE4ddeoYdBmarvQo8UAsfCCrn
+73cxti08bg3V2fDPzUMATmpC3UBuyX2+E+7llyk2GUf+RaRRKe/lZQecg9AqaNO
hqCQI6E022dy9rDHxHQXJzp7ZMtj7TGC74Jhj5EmXxh23RliIePxkSrnJTMwxrJp
T3QukRsMJvcJGOd1RSvrwJXpumGKAypXOpHU8ov3CkKiHObvU2ADglZAfCClr8rE
qANAou4GcJZ3LQic4Apnl2oqb5Yz/SqDBL9SGK90FQze8i1zSLm9ArB9sNt/pJOb
alnpk1V6N5LtrUCIHFkwzD1bBIz+9JEpfugyFO/6Ra98MtFC/kXLOKQ9WJ2RaI+H
BLrML/vpWdtd3Dy5OjXUVKnNrSBOnau4MFDCEVJn7uDfrbEvn9MXJKirx7BVK0QC
A5FlyihYhXvxi966BGojTwzq/PL8Mo16kC/Vz7Ewo3hm1WZSWnt59t5R0FO0EJBX
Z0y+/5huy+6tXxFYIHIvSupAXNCo3J56UTc0/s2hnhlARg6zquTh6RkVpa1PL6nP
r99J7k4YZhshBYSgkvRkHc3oZP6movzs17xm5k3EylZ/0s6U1Hsax5f/081L7WEq
hwfxLAyrexbFFU/ChktGwpcSe+UU9zsfhLCRic6AhkPB+LD/byCrgWrkqVTja2XZ
XSfMIlz2Nm7atRByX2x/JCY1Ldh4Aq2sbtwL1hdTcK8KEmuF9KSNwFnm5ojqBCxV
EQCYon/95QFanoMd9wHKDaAeSgD1+tp7brJZ9PEdrsOPcxs5/TnQsGa/9/zJCEVd
NlO/EMxShB/zXaoF7Qq/mQYMSrp8ttJCOZ/IOv1NDf8AZRIixkdApTJMuPXz/7bD
EPuUoFavs2ZXfpfzUU+2+p9VV0wF7nz0D2ta6pdAJRNrSo0I/X9foUlB/GkQqj7L
wlUumirNYWtEJcSgZ+SDI2f61csTllpm+ZmVPXltXbkUgleLdMt2Mpzk7mmp2AVQ
CEKK20TMG0vaAKqeienHJH8NMzF+3Zr17rAm9Rf5TTULnzxrTyMKybhNk8z9ulEY
pY7Seni1H0CE0uqPBPAzoCdEp9fyqRn7wChyY18SRRvp8+DqSX5Ncj1w/9EQPVFR
0QfnNYFGu4D7dpCllcwUu+oso4J1Js0o0Ir2xe8r/2JBzJtts5ifPYMBJwIs29g8
PuwCptPIBW4kYT4L8IG+kQU95dP4Z2EDwQKuxBBan4+ilFnKl/s9VNFsDnQinm+G
aUHPEyXzcT22iqH9bet8ZuqSlSmBn9bdmoysNW4d6EhFW/SpKc7ddeo1xFxlj55s
yCSrzPkqwqLoaJc2fjeCQTPBochZxHNcVSr3ewgqg3yrka/idYatENMxSHJE5XuF
Zkz0pI6A9iYaIiJTiaTu8TtTSjD+6R0FoalOP8MvO+AQ7Pgrsas+AuS4YotlXNjL
F4Yk3Ruxy5awmzMvTSkpT5IOcYRZkyKIbsZ41oJwz0oRKs4OJFIqWVTJwp6l++1E
2knJ8uCTwRwbM0NjjC+dZzrsoZOSV26ZEGUdFPwtJQnb5YY1U559BOcsSUVsPuoF
hNshiXGyNYtr6Hns6sW1i1lQtUgG+X2j0aMRRTTIcetCBlvRs5lhvdUuExyYIQ9G
FFFlEGD9PfmNZ6cX+I5c5DHJ+rkZ4FN+rH+DSfh7dKCVLO2HX/6iRYS5mOgfou4a
Izn35FvkpIAY5qLl1U5PxGlG0xSOaeI0r0jjabaN6U2FreE3SgLiXW9va93pM5QL
GLhx9uU4bWkzjlQ4lbV01ANt+5WcaV2HjUlpeX725nG8K7mY1zCrHq+QL3yvAiNu
CBSxJvyhQsj8UJYCcFLCh9lpevnMFSDvU0SFiC1Q5YPFn5Qf/L2d46DoYhiPqJgk
K40D+y6L8CbgdO9T00JXd3whOT3UyWcjptgpyweoKdKxx3koptQtB14+ABIFlZkR
PA51Zg3Aei8+ws5+Opm7qhw3TSDGH2P3KQivpMs3z3gn3TApAPOpFBJywjH9gj8t
VIeJfLuMG146vfYqx0J4ENNj6ksB+VBtQ37hAMbWhAh/TAiGpKj15lES7JddpUMy
8CkTfd3XMnEqAd/BG0o9bJvzuWobSt1LbD8Qq/2r/EkhcCSg21ZcpDxSPLMn0lYV
3o0mn76elMdCCGhRZwlow3CGtip0fDvjKjjKaIeTcO8TVTaYktoPZ+XzQMmeyglE
/INVrvkvaNTMoVZa+elBVjvfQGL+RJx28nkEKPQjuPZdPERSGm4W8F2meezaR/p/
OlPXE6OoFYir2cfAN8s4NNJoCUAkLfk4PJV+PvREbLYtMC4VvlZChi8gIGuBvOYp
wEa59LAONljJxpdmImMC0uSF4rBv0ph/ALbudSvp+Gk6PERdGYJsnez15zMEW66w
55eP+5pvndYJ2QfsEchLbiWOOb5Rt526KRxXWlsc+HHVHoPpJkXkJt9NHRLTSt58
C90izhN5T+icFNoFDYu4h66ufSfuXXlYyLv9m+kbjpYfk+EEA7egLMdAGd5D/NX5
oCeCZYzq86C/HD1qqDRFKPTJBj+nBS49xRJQpaFWreqkTdGjVsr4f8JjxOHGxAky
BiL+XjubUTcwcj28RvTUKKM++FF16kgvMQkh8xQx+HnHQmy4hCIRcuSsW0EdVmrT
dZTvCIKZhTmqUvrTUWeugj2VpNHsjXzCP5ckbuBmPukY3euL+ghQxjiz4uwo6pem
Hk6bIkK/1N84enBXb7toug+2YfKTKMHnLWmPjHPBxQEuK4fXv8qwnYDWgH2O68ZG
K+JTiQiDd97kIj+HEvKZ8HdHHMiR1PKgG7pHzsyeUkL5AHXUac/zgfluoZm7Ffve
1XrJHHuNY2YY1EQx9zKrdy0p1Guut+3JACH7uM6AqvHd6TQYxNUGhhEMRSI3pxCM
BE9W5c7BEFBoO3cuBAhhm/VSlXlkooz0ZRX+libEtkfZVCFF9gPHWa/obwcGI7dJ
iD3NW5Gz39GHYyPJ2g2Efuph+YLPGOyvRMU3grerleASvTNd8870MPH0nWS9MbWF
9uwH4FAv7v9QWnnecRsE9KIlQFgrrG6UEqlmxPbpCZxpkwDfrq9HL/yacb2r0m4I
pEVPgKYiZDg9qiTG5qQ6Z2ROplhDK+6SD/o2UWxxpowA2kdW4PQ7YteKKmLnPfoB
AhdSQWm+9DDczVdUdjQaEX7+JGKRgfqhnqcwpkGVbjA/D7d6SGQxMQyxadZ8W2M6
at9lkp1ztNmQIRv+KYnuyJvb0+FwwF7pTJ23PIw62lSJF7aF241ekOQGIx8EL2Gn
oaO4GK16jGGjV2bF++3HuT3qity+2Jq0A9QqXAihG/b3THiFE3+F1BQnco3w+tfg
/1Cvaq5ftDE4s17yG2ssj8OyWm6mf9eUkhLB1+LrdK3epwjO8aUKMnqi7dA+nq+x
4jzGhsjZGgJFYNsoUMA6qnJDxZpXFpShWkPlL7jK3quoZkw2Aad3urx2XKz6+fvc
fMzbQ8wOrkDfyV8o/NViRkpzxAdY/ginBhURv2WJc0Ko5QGgobjs2btGV8EJBNfX
3ENLxJ8uKysjcvkNAKm2dj1rh8zivsexqeFj6z6UdHwR2MeVx3bYWfyF1jMKRogc
uxBNQM6Ovx/1+WmC+QyIEQolsYrmj5qdGUpeSODwmBvpicP2Jozzglvd0SX9HCZY
TsnfnEl7bbOZQUKw9hd+5mi9BvbUfo2dE/mEeNWXTFj2Oc66+p3/1oQpqIpdM2as
7ITiBwH+Rpy2dv8rN9puwgN7gI9g+YxPoDf8Lfh4Jy+oumcytdX8m7CcfRYSjPKg
TBKh3Qqq3KZ+C6ulpu/ydPpck4dBQxaFhg4QN0SZOdC1XyGyAJ01nrq34bnK5Nih
53DatVjUIx2s2ccBMZ7uNvJcF8ivLQT69EQPAryp+PHRnvk2KjwwBCBlp1SIZ/qv
Qtp2+ncL2XXhG/gYDq9aj7+++7+hUpE8b9cJQM/FtVcVK7Um+u0wVyiM1K9Irxjp
52Yi5iUlExyY1TmqW29FiFOfmERrzhDXWrLRJwdOy9XefiBQFydeX0KE+y59gLAI
FF/29lud7g/LxJqSUk4tpdjMswVL+7al1uQupJlI9o4eATb5p6AWJ75FOEncnXnh
oriaQ8uHTOXPts0BW+lZFVDKefVgVvP39J4YhL32Ad8iVJGcM1QVjt910HgpiVKo
nUk8XEr4vad4JzKgetpz7/iPLWXhsCSZUx2g8q/feNkQAXpkaQwv4UssSlL9RjXd
VTT618DB99Tb1/Uut2aUB7DpKGjZAcC5u4guPJiC6w8WWr41cHk5VXWiJbQdwsiF
f6e7H94DPMFC1TGQ5habVCafViTI98En6oO8oXe5djSOZb3GQzCpOU1DTYRm4r3y
UU8uJWzhjSfBpuJ9QPUOGWnwqvbZbTYCNf+2TbkV8OPc29Wwlh3Mx6pkvOyyjx6S
PiVN2BKSePzW++Rmf+EfAg2Z7dIfV6D0g5vG/hbGhhJM+JWKYCrDjw9SOXahKcZU
dQHi9WZEteP1Dbr1Hj8PagkuFpSH3Md+WPBDgO9sgk6l7ygqMUfPdKt6ipFAQ8qm
xF9mlG6O5BggwfwQJ/V5eX7QzTxrr9AMX56c4y0K78mfB9Zh5Cyjv8rN9vYMP/he
HnXMivRrBpfH9ICCFomdbALP9AQu0tFOnBEcbeSmZCgsqWoek9FKhHbA5a1pZpVE
Ujf1L2ryLE2uQbrkwbAYDD31eE7aDZgpGKtgLD//xBH5qNdKpeQgxsn0P58PGKkN
qqxzU+07F8lLtk8AC9louI/PqRAfMv4rOzgOXp23FDVVhBCo5kW/HkRXnm6qUdTv
Cz8JBX+RCBYpOBSB3kp7TG2Tk+PJOhXL8PdE0xeToiYKSuVv5soddc157xEXYZu+
sISWEMXlqNAVZ1vkWfXlpjqYaXuZuV0gt93Pscgyv2dupyYkH5kwMdzbq8Tsvs84
muDQGoIgifj+Re/AkFC7u+TUEZ9a0rcpMbyr5CVf5C5TgeTxXnVrNt5UrDPsW64f
I1dee+qOwXSu9TbK/gzRUY/Bc8+daLgp1u8bU6bnMnvHAk73BpjDHcK3O9g2e6pZ
s6CZ3ec0WTSX714yDd+vc7q0xO3aTeAsgDFlpQYNOp0J5RjUN6lc3Mwtm4Ncv+HV
0v++N47sZz2hihG8LGMyV1jlDrcEZ2H3HfNMAm0C4X5a1NeglIZvdC4Ue/YmSw8x
/cc1pfqc/NPtSsuguAML/EhIg/4qLn/beKCURePf2qreeaUm+speWaN3twX8TS8c
pznKlgAT65WUAHynXLy9bjF2rOEsqul6bagAY8qeT+NIA+StkwdojK0H8cjQSXfu
TiT3pz/HU94yYP863qSH7wAc+SrIb6MlpLUZQD9GZoJBJ+x35hiEdtnWlsQllAFw
ieLE29ZouKTJjLCf+oKrIDHNRKiHUgo/C4by99zNMEM88CEiVK36QRVV1++KBJdX
LNhGGjg/2z8ge1/ue1cN7HMrNZnm8U9ntVcmn7MWRS6djICMsBegNUv9dyOQHd8P
UsSWGd6DOA3qEQR3/E7pCCDlxI8DVco6INpS67ilZ/DLwE+RdIj9N3Lm3vW7H7wj
4sDcdx6clCmMmdesNPZCUiJZijBS6TVp2AYteI/mdKOFVmiiWZ9UATe+fQgfhpKq
oClw5fOOc+HF5VvO4pr7FP8CckzEVsspXq1aKGnzhmlE2E+Jr+ZkT2H0HfMgzleX
Houx+yEmYSAgGIAhuJr5eKXwNTTCrE49uiJdLErXCc242PtoLZZwQU28qiBrsDkU
rTPDdh3KXQUl/9lp/fUy63+CXw/0nw/3pJVQrbLdIlL/da6f+NFFxcxYKTt0oRcv
Q9tqjQVlaHPiOpiOfr7Roa+QQb+HpEm/ructipJYyHY3y2Jq/Fgdk92WFxORoO5p
NSJveYQotJnphQwYEUCb6966rvbVSeZ3gfkVwqvQ3BP48Ev3b0QKPzUtOyMjL373
jxenuaIvRpIHQkGTS3tG7hcqqaYDGf4ArVygKZjsD4LAlLVtS5RO7/CrwWAz2qlj
wF6dLQ9AnJW9Zr+3NMcd5GUc9V7xqLJ7ZOqRFx8iP18M7qdfXyQqKMwyxN/qsWHb
2+9I1iVirVYhZv86Te43MT2yUR/sfB2H6RAvSp6glaCmVAMTQjW/t2a5UtB5f61Y
EIPi1KLfZlqzhybxPII7b+0kRAGQUH1AQ1bxijNEygRieK8ZTswh+NxTucAfwczG
w83Tr/uX8jaxQo8cQS0dSUHLfD75xcI7SSX3ksuOZFqoRXGQHGePhEffnmDvm+dv
ObdWkJhHMmzd+93dscBpwe8iOBdIRI7ruzi8NfGaLff3/GuZe2gAslxRD0mDn5g/
mhWQgo0Os46IKp7fk3tvr7Nqq/XgsY9Haeph7e2Rjfzg8m3713XxSf8I0MbV2dcJ
EwdPifi29tgEZ2MP+DuSeKfvBoEtQuIfxdeabtYKJwF7TAYyalUgbD6iey4IzR8F
Vii1rQBnh9WYLxW/2R9HrwPwikLM9K4BDe4vdFd84dHFHFoV+KoHy4a+XgtgrdKs
KHIJ7KUfWTuwrJpz1YRZePlf0DpxiGV7eFoBVpEztfFUZxvsW7BUoVafxOaxq9FE
OksJNGhJ4b/c4ji6sgXi+1PJcR+PcppqfkTi0J/ntsh/rQt9BRVNNz25Ou0lvb7t
3uxKXFjrXedZIMaXumM4pT2fp5dpVu+EhKfUsyAOKT20W86YysIkLwtH/QcYUzAr
GZmAS9SCuBDYXUpxiDIF4nxsb9F+1hetGI29roC7008vy1v0oAKurBuJMTrceXr9
YqK7nvqk57t5lD5UpB82mk++ouqECkpMpuqbA9FWKtBp1zqihNukDaFHCd894Jru
X3QHmSSwnHWfFxjaX31qUxz7ZayCWqbMXRcsyYyvyqte6YwtVghfCnjvblC3UrJQ
xF/RhjV5JgByspM30R1i0jRu+MpztTj5qsurGddZvncMUnCHi3QCcgM1sL1R2SC3
UbYu+HueAdsINuiMvj3n61mvPF35lv8AOL64hZpK1ay0yZpSYEygXj+KeCVmO/PH
1KeM2oH97bu8MSFe2QDnNdxoRcteFqQXSgJphBpmZIREmEzgS30qDLCw+6ym4jkb
L4MVkeg3WB2kp3ZUezP3evdkyUUlHT5MKVu/uZpbK9WZEN0OpCJKvoFHKd6wGu5B
wOWy/M0eg+3sUyxEcnV2+ayT3kUtjn58/QuxMlfjx1EV3xWtEybLyeQ4Z9pPgs3U
q/uOvWKGtXoJcSo3KS6uxW2v2JbjZ61ldOgcZBBGkz5SeMhZxXGyu3WzzwgaetR0
13BINcHICB6RaGimbuYkAn4HOq8T06xVBfclnT7YwMjy9wIIRZbPVA/w4BZib+73
4jDDw2Wv3EJ2Li4HxQlO7ZFc7eF7Rhu1K6iOiZNr3MKd7eO+7OEOehf/xASZIknx
oorXcs5KarR4y4BVeNy/TY0LgeejsMZ4lH5txR36Ju607mXh87bQEXPAoFaqMHnJ
esZHdhJxkEbmyNttyFtpdCQfEnVpgAnrzt01+gAZ0TfXf9/hayMXDqui3SvHAWnn
dK+1UyqNbaHRw2jzzDrXnNn2IS5TDjqrGJ5Tqz3ttZS9I7EZRxASkirwstGD8kwe
IMGl8bx14X0fR2YZ0Z6rqsbTMMGbWNSSsYoocSWyjEYZCo3LXabV5gXMkWiWYto/
LkiWbqU/bcoQO1NYdAVtXdmy5dC0RiARfSwOfIrS2N5T3bnm5ZZ2ycI0D1/e19aM
kvo1Wwt/E6ZmOLfE1md7x1bpUCZ8pK5nuPTT2AGZvYmXbLgSCEHR+PslvWRBC41v
zW9x9QpaXZYUdPKqt4jC9VMKBZ51hmH7UiN58RU9G5dOI4NO1K5e1ui2CRrwPDnn
xTuSEaMQmP1zPaWgGbohGFxGjYVmYyUIET2SJlTBNEOkOsGVUzN0IS0FGVdb4qxE
GogTNasiZv/dAKKAYqP/ZURo5WWePa6DiphqEcXE4Q0URIfCBnic0x5Soe4J836S
wip3GJI3Fnn3sBXrLGbe1fLtI2Y7hvFnomx91W8tbW0S8d257zc1wAfYAfq65Yv8
gmCwtywrFrqtvcaysDzsT3ByenPPo99WqM8EO42XKjhTEs/FmhWflB3kot4sng2D
QzxOjC77AcY34NgTaGSA+AZoO1UqQT+k4Nre1KdjMSYk4Sgd/yhPYT+0b815CGO6
YhZufuHB95aaRhbq6qpFKCMzCQgcb6j6uAdlVdxe+AJg8eT1DPFMPefxwRbp3tqP
h9gj37+YMFV0AuTtxVeYmxzYALOPh7MUCJJdnC6xZlylWFcgVN2Mvc83iDEELkba
iqBxogqQI8HrDyvgoh5ywmLM3T5FkM8si0ujxVFwrRygnCnnVwEN9bd2YgUO0gJn
idQmi7fx9MLkOa0lRYO0FDvytt+gxHAtj7UxxJIUu433k7pdkpmNSw5OK808dZhd
JzBAhj41LBlSpzZ3YJoZX9TZgd7+5CxfN/a5pQcoR2eNjzgFkTOoT2yUZd8V6fa7
BZ7sw971e/MOMwkZd8cCuzEplSzvTjzXdzxTmjjVl3wNOJ2te/xKtZsVHvqbfLUG
ZeD2nyl0K5z3a47kb++ud1Rh4r37lc0JokDbNsdyFYemeYgqoKLH4TSABDCW2sod
3cKh5hC9kFop1+RDDA1Z+hW0JwTd2vlRzXmY5q49hBSoLyqHzoV7a9EO5UutHIRE
`pragma protect end_protected
