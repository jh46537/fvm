��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�c���G�J�,=N�{�P.�*�@�&��^[��Ԇ�Ă�#�a��� u!��;*ջ�2��n��:#7��l��8����k�D��"3rd+���]��*�a���7�a�W�Ce�L������ ��5u���#��)�g���=!5�g]4�y��t�/�Y��Kw"������u�J�M&
Rܾ�a=�;�D�.[9>��_2�j)���&��%O���b�R#([��%x�E��8[���i��xh Z�ulN�"m*��5ߡ��!���ʛ(k���=���&�}�n	�i��8�=�(=��>چ�����[��/��#�qĪ�7�������m�훓((IF�YZy�r�z}G,mJ��&���\�}ֲ�n��i���*u#R�c� �zP�Lr�U��]o���� J���Y�\�J��_ա叫�#�/��1��":0jO]�T�F~���?r�c$,����Ti�o^��f���eq�d��U[/���s������h~ߌ�o'�%v�j9���sY����2D� -�'%��Sn��x���}{<
��i���y�+N�i��.�w)B����&�`�ܜ�ۮdA��@���԰g�TF[ņ�Z�W�y��t�3�����jC��� �Ջ����4��S�/s�w�,��b��u�ƶ�>��ґtչ�J���F%��j���`���C�3	��@A�#��|���H�E̚n�s�ワ3.���lrӂ�|Q~�]��]�\!��F0�݁ʃ���Z5�;.Aw�� q���p� V�N#���m�R��6���~���R�t���[�0R�Z�aK&.�>����?f����!?��$:a'�/)�P�~w�@��z�G�g	9a�8�F�!Y����U6�<��#������ş�Y��Gٍ2-F0��eJ���XݓJ�a��dgT������� ��1�!z,�g�
�"��2��1�|�kOEV�TZ��e&S[��n�S��� �d@\�E�3����&w̜E����+^A�9,�)��������.T�^5N��8j��{:/����
�d^��U��N{�{��ҩ��I��Rǀ$Ɯ!�M�b!��~��
��Wy?�g�����[��)���lj]�.f�Q�������(AD"�d�*D5��v��rv��+����B���v��թ��� ��)���9�åCC�!��JfU�%�.1�`����nNf3�Ʉi�=���kH�� ���U��%`
e�R�} v�~Ǐ6��dq��wΤt���.υ���֣���gIM�B�r���I��|��ֹ����C��1�8�)�F1�JE�~�N�RӖ��A˿o۶t�uqM�z8�Z���p
w�(Y�t�Y�+�%���@h�����/���hn�`�p���C]����d'X�BQ�\�$S����qh��n��|��, _N�Q�z�9�.	��<����@���ف�6x�F)�4�fp$�T1J?s6�uA&o��f,y��*UO ؚ���ѷ#�7BVu�O�S�k-�;��9+p�����R<���؞K>��ݠx�Y69<�m���0�N��0�j��Ns���|ǃ��b%Y���(*�`Rs���'zN�鬚w��~t��]�*���y?J;!��ק���D�jX��P��JUVx~�����5�iE�G��+�ǻ������k_�3ʺH�1y���<o�����aɑ��ʾ���,B��t"�iK�ϊW�а���5ۘ�W|U��Y��tN�l��@GB�K�(���uq��}�R�w�5\45��	b���{wE�`y�q���x���W�,�Dmk�.��2z�M!��Sm$ov�bl�HK���i!],��.���jZR�*.mY2�k�琒+��F�G� ܺf�of�ɳy9͂������?HW��(�~��æ�vƨ
��\{�&���'$��RJ"33�Ak,�E�;�_r�z��Q��^w�I�<H���I���7�H��0������U
V���}�b���wa����Ւ4EĲ�[%��\>lz53kB"{�$�O�H�P�􏜸��֬wB���Ŵ~fB<V0�{\a�lD����0 ��
��z�7
�.������(�4�x�4��1!Sj��P��z�ޘBV��:�x��o�ߛ'��v�~�� Z2����N|0,����l��������+��9VݮF�wEa$�k]PK�sT�>P�o4�� K���
�����~&��hv�As���#W����0Y$I�О�_]�;[�m�ҊlT����T�A�K���t3Fl��@���dg�QK�Y�":��Q���5������XZ�2���8���E�w��%���,�ʟ��)6�?l?�#�q�\��������{:��{���
5�c@%k
��~)X�C<�l�و����8�f!k�����@q���1��IBT�h�z
��'�!�ܶ*K��_�ݗ�n��3Z��J="�/ă�wA�^A��p�v����'/��3b�<@��'QVSg�����8��Jǰ��6rE�z%˘ނL��;\A }�Fh���Z,�3~��a5�oj��G�BR���f��}�ӣq�g�p���͉e�@��1���2�E~4���������
A�s@n��;u�u[=�o�o�beQ�x�+�¹�_�)2�W��_�S����ᏻ�lg�ۦMQH�Ϩ�i��%�[�9'�D����)����,��j���{0�
�I��=����
囂μ%��
��>�V˪�l��1��Wd�pܔ�Y�#��#��]�=A:��E�������lЍBO!��=������,r�u\5h�44NL̕�3�[�`��BT"<Чs�#�I~��ÙX����y�S���ܖs�[���\W�8�n����):a!�m��V���p	� DL��G�U问0V�e�*%c<��D_��xިfu�CǷ�����Β�j�4���`?����܈��IW�����F�^[N�&)�)�ܑ*Rx�j�È�ƈ�K�}�Љb\�2���{3:,��|�uP����x��UX�k#!qh���A��u��BU��"Jk�0	���u������ƷU{žU�e��,�){�j����MOG�b�FBHd(�����@�2�|�8��$S^�W6�("�D8������b$�l�փ>�8���>�O{�]��Zn��|@�n�G�MǞ�2Zӫ"%���P�Z�ym�M�-��]��bB֮R}��|��ӶQ���S�w!�k��U0�J����27:1��!���K�*,���^B�2�	����8uRm�P�J�J�EB�4q���ōN"�Q�l�&���ZV��̠Y���L�BJ�oE�Z1�e��'"V���v��0=�ui�a����Gg|�q$~T��ql�z��1{V�ũ���0�DC���;	�͢ �Md4�������� �wHh���t�L�����+ax���ZD�~�\�R��62�����z�۫E"|01��\eW3�����BK8�7���u���|�j!]ڂ�)?�3���0�T��(LN`C����)�:pU1���Ϝ���?��L����R��BX_!���6@��Py`��lv]�EFJ��K�>���� �g��io*�P
ό9}���� �k��2aqâ [�ol����WH(1F<��s[�w�e�`���d5�|�P�2"WPb��YBe�>�m�^����9�7CQ7��ݖF:�ù�Qo[VI�_���Q\�	��).g�Ë�q����ju��a��<�8XN��{s5d�su�ŐJ���EE���ho*�)"h5 ;!�D�)���K�4P�h����|�`i�z�D�\ ���\;�]%7�tw��EQ2���[��n+����PPO���X�� z���#.��[���p������]�|��27��HlE������@�Q�۠"�� ��9�3\(�ŏ���nA�ET�mPΫ���o I�=	X��7��6��`,�/��5��'b7�k�������;.���#��̸y_�˩��w������C��s��J{��|���1�i��	�W��~ϲ�b�)/>�&^�ɮ��/���}W7� =�6�j��m�z�N���N3�:�9���*P�q����#.2�|MI�߷�G��;�N��u�n��CDs��IЌ��9eί5"�d�m�Bq勾����`�9�V|�_/(�Y�n�1ɪ(���Q�HE�@b��(r�{���D��G�#��q+Z�pI���G==J�t��.%�[�>U:P��ށ��kTq~��F�tG�K�-��h|4�m���1�0�߭�aI����������~���	W��Y�YW���շ�m.����M�f�� �a��a�N�u:��O.���r7�f�V�{��O���_��yu�zXF:�k�֖�鍤O����$e���9�&#O�ۇS�����9�c-	�I z`c�cd�gr�}��SnY��_���U���"{�Zx6�씄�`��}!��T�������Ͷ��͑ݛ�.�7E��2c댞gQK��A���X��n`T���1���{|� ����ob9t_p�̙�	���=� HrP!O )��dL#h<&hf\iV"����O�UT
Ӥ��p��K���1��j�.����Q�'	���R��l����+�_� ��D��~;��Se-�)��T��8��Wǩ��$��S�	��u� &m�a��7 D�X��3��rR����˰����G�bO�=~�98?}+�P�g�3.Q{/���	���a���L�-q�fT�W��Lz�-�\p���u��l˯��W�g���� �nq�_ �,nL8=2�Z>���/���C�gBX��EؐK��ʗ��`��d�[-�qF��q�8;�p��~fsf	4���Ih˗V���/�߳�<�\��Pg�>�罍�Ͻ2��8t�!la�b���Z�����=�p�%��td���p'��憈�⤴p9n�_��q��ܳ^ϵ��d�Ua��Tl �y�4�sd���-��H���+�HoZ���n<&k�&ۧ�&�r!���0^[���U<uP0�N/�T2cM���q�$x*B'j�;菪�W�
<n�!	)�AŪ����6��]K��Y�!`�#mOW���xTE����E�����Nmo櫨lǰ	ީl��ב`롥����~0��-A�>Ҁf[�=�����Ԋ8�P҇��G�fD�xt�����],����Q�oՆ����H��y���X#��9CL44�7�Jv>�8?q;�#��\��<���0P�T�|���H����@c.�<E$yp*A��혗��	���jh����:o-��Wqa<"�3��/o�E����~i�����||< D�%Y����E�i+nSF�v�s����Y"E^�;et�^lӉ2�$��-?�Io�6�a��'�z� {R�A����"_��y,R�&xP���na.��}0��i��1��fZ	C�g���?A&��7v1���`��{"{#�!3M<9����]�x�f�g
��"�[�����nCШ��ȴR��>Әщ���`��{��Ã_�j��,A���F s.�����Wl8P4�i����[˪�r��-D��`���4�?�'�E𤍎��$7	*��^0�G��T6Qº�+����{ڡI/�5<뇰2�"}����O�O�f�k`t3UE���Q�q��g�b�*t�ih$QˤS=���㒒wM̈́�s�Jd<��0�%[��،h�+��$ ��eY�F��U��2�x]%g�+6'Ϭ�ks,�������'��	��f�8e��t9�kc�J�J�;����r���U�(��� E~XD�4Z���v����e� oV١fp�/#e�D�O3��aW3��t(�)4|��e�h+:n��jr��h�s�Խj�����W~�K4����m-�.�G�?[O^��)6Q�ܙ�i�y��9r8��6r�7���e8�Ȭq~���k�B��'�ϱ���©ׁ�D}����ZE�~GY�pC �*�+ʉ(u��c�b���&��Z8�����jt5�{b8��/6!�P��E��:+��Il�;zQ��p�m?c��1V&F���Q����4Nm�	�2�+��ܝ���ͺ�O���3����.���C�a�L
i�0��׎UDM�_9�4��Uo�K����C��g�Gs����v�2�� V��wi�
0�K?oK��|bxRʌ�4Gi?ʵ�ֈ��tTr?��GB4�㌀4l6����";ʽ6�[�ϽjX������TL�����U�Wݕ\?��A3j ��"� f��� �Lfs5<^�������P܂=(p�ob� �\��֦���<}O俣�t�-#�/|���|�����ʿ�q�D������(ʔ�gi�����0��sp�J_���G{9zZ�T�ɤlBxvI#�M�s����[���%f��hܫϯ'L�Y9��J2��sߙbxO�j��4L��N:��
+�����R��1SP�}��H�