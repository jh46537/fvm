��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��x� �u J䇰`#����������T�jCQ�?�!b,1g�kG���K�J��@�v9w�KC���`�Mĕ����5T�7�9�Z�0�,�@,m|{�{=)ܰij�����{��l�K2��XD5�j�V�5�h��ԯ,��2���eӌŢ�\�
#�.��:F�3ˢ;���LxZ���7lU��+��8�c�yJ���*)QoJJ���m��>��%�=]6s��fk���æ���BT�7�~Xw��yk�~��<�ׄ�Nq�ER"p�K<��_��vs������`B #��W�RL��F������`��Dy�D/53Q��Y/�:&,T9eJ�񧱷�rU���������,"��[����e�D'��&��a����ڋ�k}�����G'�Q�b�!��ώR��v/዁~,ü��F̣9Ȼ��T�3֔4�����@F,��� ����e����\�HRz��V��d���l&+|W&��jn}�h�ܚci7*-���#q=%�v��R@J沛�s����
��x:d���;A!���T������;�~q>Cm#OيG@Y@c�}�ҺC��z�,\�r�'�sAv���T����&�a#ٴU�l�Fj�%^��)q�.q��G�w�0�7�~�M�p�ԇ������b���ش�R�[8��6��2�0�r�ppB��y�x�d�Y���߼�#���^bBb�%T��	��%�?�.�?F�#�/�K���u�w�{ A��Kyz��QN�J���k��:��;#����>T0��4Oç�p�3��Qa����N`��K��R��㾴��o���NUR����(3��Y�i�#Ãu�4e��� �}�Ɲ��b��#�Lɮj��^r�.��Ʀ����3;Y"9��,�↨^(:o���)���X�wϽق�j�>���IUW�G�=S�=#4q.�Z��A��Dg蹎�D}�pK�������E����c�Eo�O��ǥ�7T��#.��ê�®L����-��≻�A��Eia��E��ﶃ�f^����F+���[�6BG-��r���މK7p��Ԉ]x�780��#�W�Ϣ���D)��m����kV���؟�#�}sg���X����R�����;� ��ǻ�a�n˃�n;��i��rY}_=V�@IK��J��;'c�6\a�� ��+]������6��l���#0�e�D�1�$�>5��T�g�%���I�]��KU������iOKv(&�wF)^P^��J��Gݻ�BY#����4o���|��p�:룫�X$y� �cf)�.�y��"��f�G�_P�$�Ğ��$)��I%|������{Nw@�R��}��W1���>X`qg��C���K����j�qyZo�{(����t�O܁�-o�������
ؕ�3'���v�^EMqJ�:o��6w�s�����`/��߂�T�Z��^Dk�:h�A�v��2A��`W)�f}D�kQwxo:@?<��3נz�(�z�L��΀�\�ذHF�#�c�A{�>���4a����w-=2� �1о��i���ެ�Jๆa쓼/�>
-q��Jo���>�!{X����A�& a}vJ�:��"V���`Ҡ�J�x�h�!Y	��a�Wn �b���IZ7`*��X��-�Z'��4=�`��J�9.O/�*��*Rô� 2��ŕ�R��ۓ���.�g�@p��F8/^���=��S��fad2�J4JW#�^g���_�1t�3��'��$��O��RD��@�b��I��*���9jO�t - b��p����}��D��`"�E�֤ibV�h�-��&�P��?b>-E՟�+w�qݎ+�j�����n��'����6p\f@`����E�=Km��]Q6��Z/��o����߀e91q;Q��H�񗬊 :���X�{r�rz��M���hYQ�/��X Q?��0��4pEa�<�y�X����h詘��@~��$��B֣�8ĥg9"���?J��_����H�w�qo0o���Ӹ���u��?g*F��P�Ǹ�W��6��_�ujuqs{���k��R
�'�)��	�>)^+��d>d�%O�x��פe�����7V�0�^:�7�k���Q���&�;%��`�c�og��H����q��
����v�/-��1�k�=HR�d6��X%[�顫����
��;p����}%��=5��Z��.�:v[ꎅjGTD�G+�� k��hvt5�\��