��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<���?�)�,��}>*�;3~��2�l�*$�T����C�=��ʖ�OZ��L�(��i�*hwnՠ�M����o�T��J�&M��E@�#r�X����4"���%�J�=��ի��9}BK�-E�6���%Y�1ؚ�Ъ�@�̎��c���%�K�L���̷ݯ6��ŕ7j�e��G�|+��j�j	��ul����df�N�#^�p΃̲l��G=����f>6�ǡE���rĆ&�򸉹�Ȭs�	 J�Ѵ(Cf�d9F��59�T��O��&��dn��0�?r����r���|r�n̦��sɋ[����*��)������A�J���c��n��R����,���Ok�ԢtM����.�/-�&�_Y]^���;�Y8j�S�C���l�=���olx��j�)�H�=
ǯ�Ӊ ���AI���$�^S�e+;�ez��!z{��W'_!�5p�1�8����N���ĉ��ȝ{��#��A�����z�-<�P�Ν$)�X^0(Q�Dۈ1���K��@\c�����Xϸ��#�;QE@b�*UiB����WD��Y��L�I���b��LSY1�٥��G�]�G�`.�d��UR��ne�l�qNv��4E�3d��P�?<�nhLK���[�b���!�T���m��������ʂ�~a�2q����p5f~�Ňxy@P�'����| �"ӒBȨX0k��M��5G=�q&u\���Q�1J� ������K�@����e�k��O`���_tu�����P�^o�4�P��b���T'�G ���+�S�E<$"�+ޤٷ.��kN�ˌ���w�w��|4Ɂ�Az��oolӋ7:�O��(�vr9�.��*��A�8p�'Hw[�WVV5�9Nm�h�@�*Y�4JQ-���̆.fW���E
����ga�,Aj�r�4��M�ԁS��?h�����
u^
GU��*w�ސzG�G	s�O�F�jR"#��M��TT��o�t�\{];�RTt�U�İ��寤��5$�ܗ�5�ys�[̓�fI��}�ϪB�R�]�&<?8�4���|W��i�zG5ͪ4�^���7�u�4?)�=�a��pEŰAӔ�Z%r�@�2r�gD	�rOMj�vߧv��fVo��t�29�G�#�� �6��V5��6��Wcz������kt��\� (6�>�����Jc4,�Pv6��wM���7�p��Y<b� �>�1��CRc#;p��7���C`��F��6~����G�m��:��d��bϔk��vep��`���i1%��Qo14Ѯ�E1����Z�&Vʶ��!��"nâ1m�$��{�Qh�/�.��5O���(��e$Ԥ��}��Jp����,� �)�V|@�n��4Lb��D�j�o.�н�V��Mg���$��>�Ĩ�=�FM�"G���"�$�J��^1o1X ��a�϶u��ȷ	� ,9�������o)rܞ��ˊ�;���Rg��z�&�Fj�&Q�z*ks�0��No�z}tC<�h2ֱGj���6O����^>N{��L{�uF��_@+����s�\j�s_{;�_�X���>\�F�tYGE��fI�g�{��M4�i�@o�����X�oT�E���Y�ڒ�Μm��x��D��=3Vzϙ�b~���(�t݌:.����z �&�E�\�J+vv=�N����";�� �	_U��o��^�eO��a�3�p�s����l_��f�)����x�J�VX��5�+`��|٨-
�.I�r�[-�v�mh	1LQ�I�N�L��qpO�!Z"C�]Pt`�6�G6�����'��h�VP�4��]����e$��'��g�/������!�\���dxiV3���F�JY��8��ߊ�l�ݍt�_2����1TI4w�I���B�L�,����m9��Ɇ3)�h��A�9�����?��Q�
}W�6�lh��X�C�S���V}4�bOn���q���#{;�"�Q1����_�j=L���lT�h��WȬ+��G0I4�����q�I9��^w�l�-�YgEE��v�q�'�3t�5gᠨ$@J6��ÀK?�k� ���".�IǺ`��۬b�� ��h��ڦ5ے筂�U*���!)�4�k�$!o|{�/p�	U�v� �ҹHON�(����!E�����u1,Е?�lԞ68G�[�e��A�Vd�e���j�a���tG��ܔ���u�3f����<=WuY��EM�X6**������#�2**ް��k�ϓ�X�țKZ�X�v���Th���u�Q����X�Ju}�#�̨�7�.z���?�k���Q�8e����Ig.zn�H��G�S�%l�lw��x���_@�ْ��XEA�%�Bh\DA&�����|�t�=f�&��{3�d���F?V��Ak�K�Nx�0�Z	t"�N��5~��߼�;�����`�ί�ݤe{_vɌ����}��V���Ɓ����Gj��d�ˎ�oy�d�%�;��	��"���V~�H���b��qf�7JC!C4��I<���u�ϳng����X��9�0��'��?H�2�*(1¤�1�[d�FJ�*��J<޾g�;��q۷�n��]pJ�N�/�Hr�P}�>4�e���RX�¿j�*��9�.V8O�N�
3�5�ك�t�lV �,���" ������m�Uj"�\4<u��gP�DS�"����[2X��k����U�Hآ\c��(bQC��������ϐk�!��b�ȿѭ�F���p�	8�f#�s>n��>ڈ.'�3�����ό= �t�#���+ ~ kQĮ,RCHj��<;��j+;�3��b��$Uә:B�/�;tL�(t_Z�x� �����~���=��[�"���_<9;+
F��.�6���Ŕ��)�&�4���]�V܅>Y�b,�]���]_D�S5](/B�3�cޒ�BҐ�̥�O㞜;]���ab�]Q+j�Nl|�zp���5��y�ɉ�~�eP׷(��X�>�d�?�X�k��#��<�)�^��ƴ1�?%`ɿ8��ͅQpD��d����~!���H�͎�6m5#�Pj�&QN�=6�D�&3L��ޘ_31P���+�z7��+��2!v] ��?.a��W�����"�x�- <���H�\������W�y��C��p�\�&$�cXFfضX;�]LM;�9�d,Uڤ�1�J��%�- �U��E�d����\[�.��3��A� 's�	&E�XNx��#3��]x�9 �[��߮w�4n5���wd��s?h4	��VC}�zg!,�tE7�?�7ؔ���C��Yr��\dt��j�|0�d�h��� ��0:6��<���"�A*?q�7<�[�!���g���b�.�kjL��|�����-��!��03��|��۠R�❇^0!���1:<� *�yjzҦH�v�Ӵy���S�qm"}f�6�D��ڇf2[���U�v'�B���PeW��,� u�AߤI>nK��+��hu���t���0>�Cg�.��Sӓ�V�:d��qj�1]���Ui<���g�(n:��0�Ǡx5K�lΪ����7�j��W��.��9���w�bU���9C��Ĳ��	z��pZY�Y�{�OvVΠ('Y9GL���;�C](�d��j�S���c�gv�ݭ���E:$ޑv$�%93��7{�"�1�}������6��S�����^:��\��7bu���nd��o;:�O����&�A�^�+j��o>C-������5�7r�3'L�z�x'�z���f��HI_h�PdGz �ƽ�c��;����k��Cx� @���@㱎��8x��\���4j�M@�۲~Ps
�����?L��� ���Ar?e"c�b]�j��a�O�n,yK9{�4E�/${3z�&��=c�<t��"w`R���9-?/fgH���&��y�+o쫋�8�a���E��/n���s���YI��������������z9�@�����x�3�P=qm�ً�4���?�.} �\:�w(:�������)B,V� H���<5�^)�7��G}|t(�O��M���%�G[ZT�wCy�3?��6N\^چe�aq?Lf�D��`+bk��(�i=�mf4h�Z���^�L*�:���J��k�1���5�T�4��<Δ �P�l/ŗ�T��VqyƮ�O
 Ɇ���̶�ltZ �b ��X��������*6[�w]�U��P��=����o�h��q�.��|m�LG�w�j+���h�ݥu��Rua�D6�8�s����L�ĵ�66�3Y�"��1�[�ݵi:���DJi K<�+0*�ʉ��ܱ{$�l�-���7�L��Gw�$���E�:�pt�&�5՛�H�d,Hw�w�&�2��_�hZ6{�y�����O�4SWF<׼ٳSKu�ђ�4 H�>ن�G�R������õ�u/��S���G	�@���i�\P@��b�F����2�{��Q��t{������sMh�ߣ܃�j��g�QEh�G����|,C���}�ďO�K��Ó��'�l u#�vPҙ�r`*�q	Ԁc�Wqs�BXf�aߑ����(��θ&��10��XNrj�9�>��U���m {��G��
�Ҕ�*֨E?+��5P��S��v����22�a�z���,y�=K�Y�^U�qm�!��;)v�}�N3�P��-z���Ɯ)]�M��%Q�Z�jKm�`
��0TJ	��?��J������vs�/J����W٩�1�̊b��8�_x�_	e�v�i�}�-q���4��$��3v������:/�����$PZ)>�)X$�LGКd���L�cA�|O�x�ļcH O�"�����h�X���.��Vi=�� }�:�pM<~�CiZ��I��vmv��rz*���T�U㈏"��t�#�sg�G#^t/+%TǪ�D�48e'�Ż�Y�6�8:S��9��6�$�7�MǤ��y`�`e��_���K�8\/���O�/(	�rà�0�^��1)-
��*���F� �b
�,y������	�&�\.��K���;���8�F�Q��N���k'ӚPok��P]� ��c���&go�3��?��.T+�M.�=\�P�#�^��E�2Y�!�S�o�9�4�D�ҳv�4���3 �&���CR�hSǐ����V�ϓ�ׂ�(~�\���Cg�\X}� ���Ӻ�4�9���;4)�4�=4�CS�F�H��(�j��Ɩ�a�q�=�����HNcK�5vL=2�G˦ĲսO/ȽKR�jb��Z�3М�aIe����[g��6�oi	�[�4I��\4r�2Ο�� σ})�(	����I�P� �څ�8�2���q�#'����9����.ǂ�d�z��;�ny�)��83��S3<,*�j�Br�6L��	��k��^]+c/2�Y��UXqd~�wb5%��ف��e�}�_|��;���/����l�V�2wD�dj�M���&�>��c�� ��?d���(����S�ٲ��_�A�k�����?��v6n��>n���6��D��T�����+��|H�c6�I�J�5�ڻV���%ul��k��G�=R�!���Eu�:�s�;>���B����1�X���6�e�#�X93(׎�;}9O3u���=D�>3~mu5��ki��v#��*�/l����U��oE��ѡ
DRDJ�'T�c,��:���C�H4*�@s/��]�iz�vc~ȋQ�t���X|��,R�r^��6�]��޿[Gi 4�!V{�t���;�1�Z�/����D����Є�R���Ϡ�_�7#P.��NN�n<}^v�:R�T)���3�.)$��	�(�@O��}1��%�9��=�Fݟ��"����|���?�	m�F�����_E�F����EPh/�{�8�M�.(GH�s�ynd\���s��&��?&����3�и��T{�涧�_`D|��mo���ϣ'˩�7;>m#Vv��M"�w���V �s��A��o^���RoC���`' �	t��D0C���Y�=���7����.�V�  �a!�4��NO�8v�Oh(D#�F(�LK��P�V�J�Hh�Myd{�xW�(�<�z��-��~��T�L �mQ_��Wd���F+��;Z�ξ
9˹���h����(��V�K�k7��1����X?D�T���Un`e���P�m�.{�f�����V���|���HV/�^ApQ��y���;�=#�}�H���܎À�B���w2~�0�ɗ�Y�5�\])D6%�y���R���6���2ߌCI'�������{�����[��ހ\3��������"��ޡ�z���ߵR��?l�eVh�&����d���-�}&��e�� ��6g�-��2w��ʢE�!�3���$"yH5�6��,W�Ey�������%I��T�4+�<�M7p��ƛ�ᱣ,��\@h���֕0��!����G=�(nl�Hx���V�w��� E���tSxǼ�Vc�rv_'�<�P��#��-;kV4F*��ҵ�Ji윂����\n<�vϜ8�>�K��iv.���y����@UU)�B����9��ʇ�k5�����?���`"�!�&9����Lޒ[������jن	���w�; l����Iϼx�iBM�aA}p�8@i��Z���ٽ��%���ߞƞb2�����W��Mڎ�P?�ز���U-MDz4Δ���*�(~#i7��0��أڼ���NW��H�g߻�D)02�/����߄��~�!�����6@u���J��6�l��bfL�/�C&X|�U�7V��c@�]�SW�A=���<]6h2��u[C�b�h+"<ٴq��	f�R����+_ǘ���O��u1ޱp7q�Ty?��[2�qLX@���A���հ3'���ug�\�����0h���Zu�$wE:6���Q��	w��~*0���Ђ#�c}��8h���V;^�6D��tZ#V��c�U���d��U�հB2v�	f$�?]��͚�_��0淾�����?w"�f�3tjS��DM]n̓����_Q�'��Ə�H%�ҫf�N��8k���2`�P�q���T�R�M��Ʋk�5�g�*�:H���Dݗ�*I߸12��C�ȁ�qq�F�(�f�L#�e2`���w��d��[ŐuR�}�{��"�z؍-�),j|��2����Ǯ�I��ט��(�J��Ǜ�U���l� ռ�#5u�9���.O92O��v�>�oqA�#�lc���NДť���,�|�d���������R�0�- O�1�����Z�ű��`�$�)��d�10/Q޶7��7���\uh�~���[�!�\���~�/� ]�y��-N���7/O��1?��=�z���m�.�)���/��h��Y�|��q)�q1Î���L���9Z�?*D����֟����5��^��˹��e�ҭ�݌i����
��}�zr ��� )17�3G�⣉�A��@�<��VC�u�èܛc�/h����e)����:���GI��aʇ@g��dO�b�p�M���%	E�A��
@��/���
E��h(�]�8euU),`G�����  �E���/G%p��.Y�	ZY�~J&�n����d�l<#@��{��hχrs�(r���/�~�{�3/:o�'���0
�ܓ�|g���=��ߓL�Atd=��ʡ��/4[�X�����.n�ק��ag�.;���x�mI��`4��f��J�\>�{��p@��^��7��.���?e�7��5��%����9���³k�-�Q*7d*O��$cz89��e�"���v��&����r���}e��R�3��sW�ON�~%`YL1�A·	���K2��g�rbR�`h��|��5H�JT�t%Co���$T��m*���\&��Q�=o.���uEh���5�A����P���X�V6W���DЯB�� ��܌����c��N'^XP�w��O��b��&�^�!۲O�}z5���AI�K��V�z�~/C? }�N0g�;rِ'�8��9͜B�w ��|�#q9G�1q�T"��BZQ<�T���W{9�m�l��MxCq�욺M�p�u��(|x�	ӝꦩ�1uk+D���!�h��g��*���Ҁ�Ue),ϬT��{�� �ԍ�7����pZLA�f�긧ύ����z <�A�d�&{�%�Ń Ѐ��:�}0w7sBgU�7��)d���R�Y�>Wx7kz��$DH&��� �/]Q�H�9gO�^1�7�,���*� BХ�o��-;�DF�st��_�ד-�%g:��d	���û�,����-a���>�C,�	�xYͭ~L+��s�0;�uY�-�Y3o� ���:"���-�a������3����z�ON� �ub����&��+}�`f����I��d��*����`a���Aۅ����ҋ����V��*�]P�%N�QA�J<�C�5Zm�ԏ��[)}��g�G��A�8�,
�w(i��A�����
u��ku�m2E����!�\Ʌ�4��R�ʁ�m����ϥ{���fa�e%u�	^^�1ئ�v�h�蒮�mRpk��4'���6Y�;hx7���ڈ���U��}D�������y�nM��D�Aߓ����Ы�LA
//� �C,='C�i���mb8�2��p��h`w,ml\�&�H����:�MwT�@�C2OLX�]W�M4Ӂ)	����чTz��	�g1� �F��`[�!�Q��ѩ=���㈈<��+��_������pa_���u	]�Zr)��V}GH���ˈCf��/X�t�D�G}r˶�5Z���B�a����;�E8��Re�E��l�P��p��� j��Q�U�,����TB�}�;�/�3k3E��mee1�l���t����4��I%!�q����.����1���j�LjȜ-���=ڪ�`@�g��,���F�[�\R�q�24�@�3�OIG�~r�T6@n��
��W8y�H-j���׉��r��)`��៕cH�!قv�n�䊯õ�r�(��-.w�K��W��4�@��1?t���)Ą���`��!6��F��4���t�Hǿ��q��w���T�r?�PcC�p�9r�V��Ũ�K�=�'�W��[����T3����#`����{�V���:��)�S����v�ȽW\U'ӭ�.�>��T���K۵%).<��Ϲ�i,�G:S:���ÏN$�[�r	��i��v�F�H�]��+��7ȼ�����$��P!�����1vC#s�_pR��ُ��J��ȏ�M�$�T�`�ɫ��m y�y��3�~���^���I��2�Ra��E2�e�j�`~h_G�n�U��.W 7!���aa��9��=�H��c�D�n����[��B�s=�Y�5a0H�Ps��v�l�hP�r:�a����ӂ,��c��,G�<�z8&����R:�)3��o/\ˬ�D���g߽Q�+����?1cEI(֫n��Y��ߘ5`:U-#��H������v��]�|82�.��A������g�B�� M����z���t�H�lj4Ǥ���OI,4F(����~�5��G���?u��ͻ��n�C�.����׻�I+R��<u#�+ v��d�^���)m3���!��F�Z�����tlv����+W�x� ����)�n9R-�t��A�5��$o� �	��g J�����>]c�������6T�2|'�!�:��'�y�rx�KNE\O���g\<@���t-O�K+�h=��������ClC�����ŎWj��i�����}���i��Rc{gVDԻՓ�)��
�v���D���0��Z��
�Z���w�c։ό�y��?{:�C�;gpE��u�ގa5�(��ZmnU�F^�	��4K��^Ǹ���B��z�|���t��P���\'y\�����U��*A��Gz���m����KYlN܆�)إk�	�~�wB mz &?���eR�l	/h	���
%K��X���[�h%J��	�r#����=E჏�@�9d%��۹V������1G18�C=T�huRKK�,���E�1n�p��<_�MFG>b	��	C������_.=tS�����c�Ǻ��>�0z���S���1,A�B5}�Ouj���Iͱ��S�&��$��4������>�oH$JOS� ҳ3��w1P��T�ѭm�������'��j㻰v� �<�;s1Z0�,�DgJG%��B�6�O���~|hs��&���o��x�!���.��9�6ܣd�0�W�X�W�Y�
�)D�\K͹­���d���+F,Q&G���3��������u>��Ѝ�+4��~����?"һ�q��x�^��:�M��X8�I��e�(b�s��K���.￾�