��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{MEi$ ���ݬ��Bj,���C����a���Ag�a��PLW�J��"��zH4'�2Bu�AkX?�� 4�k!a�Ył~XQ�
�.}��N�杘����
��kv�Yy�wj��ќ{x#�p�G`rSF�vP��[�Z���`Y�GH�IB�ڜ�"zww���dʓ#')$1�E�c}�a� 洱�`u�l������Tf�.��I�� L�=�nW��-��$�K&��Q�{F�,@{�jy&�Ry��<�U@`��ֱ��>Z���;z6a������p�fI����P#��J�e늕׋�����4Y�����Y*g˟ߔ�Nz59�wT��r����$Z8��Iәt��N�X��A�[�i�oH竣��p��H�'���,�6V��rO �t�qY M�f�&F3J��Q��8�=�Z��]�i���1f�YZ;v��_zQL�z�
���#T�ȵ܂z�UC"v��;�;	�*�c#�|459�/���;�%�jC��[����,c�� b|+忽Q3�|�w�6Q��9�������Q�<��ܕ,�����|��h�(U�B�8-nb��aq��Jݷ�Ĥ���� .d��L5�}��oEw���4�s>p���m=�L6�C���C!��%}0�H�
Ӎ���7@��Y�����l��n+Ivj�T9��оVA�/o�-���@�e�nhI�[�}�,ѡR� Q��Xw�Qu�T�>Zmx4b/,�$�X�A�V��5����0?���]�Z\(7P�4�C�=���xF���0�����A�ۇtl�3���'�O~��8�7fà�ˈ�N����_�R��~N�ӿ�~Q�=�,��ES������#���{��w1+�;���|�+���Dv�1m��|C/�V��n}P��8A�8�W�q����V�hi~%n9�^�DEǣ��_�2*`6c��,�O��9�у�o�X:NF�4=�[�Vd~E����i�w>9p;ӽIM���МЪ�����eO�zSQrQ�#������X!q�;�����jdڹ)�Q�j��[���ྷ�����9����=����
M6��bi���;<Ш�\Na�y�:���jeR=�r��B#�@�V��z��'�p��"q�͙��ѐq�r�y�f���~F�
�Ԕ��aX�/uq �G�\n{A���Pl�Hz��C�^���МI�(���Ǭ�L��M6�b�Ā��CM&���B��L�iP�*�����|;^��h�y�n�'������f������y=�,h~¾�Ԧ����d�6��N[)�@,3n�V�%�<�93��񸸅�;�@��1^�݈��0���6Tu���av�9�߬e;��띄�;<���@�5�g��D�={iP�䦮M�(����|�d��F�$/ѩ�����0 ������C�Ka �Ҕ�~	���a�_2�9 1&.�3�9m-���8��.�/M��)A����@F|�(&
�Ʃƹ��T%rr8��c��ͨ4�^���Վ#���)����0�?��>�\�N%�s�3�eT�l��j����ECJ  5:�0����yO��A����
����������>��;���R�=�Y��Ԟ,QQtP�~���+DZ%+cmQ�_PV0Ǣ�6oN�� �rŴ��|���Ti��v'vN~d'Dĥ�q�����+�Q��7�^�>�3��y3����>!��c�=���1s��(7����o\�n����Z�axz���vf���Kf�3eg;�re˗�>{�9�W�%b��.���j��C/]�g^���b��gC �e
��C����	��ȿ%s�Yچ̈�U��JgJ���v$������p/In]�ё�x��UHO������6 3>��Lr!>��U��Meq(�~���mhP �u�W<���gb��{�Jc�#�N�&���9xn8��e�΍vnDI�7d=t#8�u�3$�S`�nd��'�_��R�ӛ ����i�6Z��k̇�C�2���0��P�fs_U��2�N}z�Vy{Z����в�	�\�8���ܔ"n��.����_g��6����M���! `��՘yܙ���| ��{zMs�b[�.c3շ<\x��ӆ�=��E(����*�u�]���Lo/t�2I"�7�ށx�A(GG��c����@���$@�_�RǯaE.I��独r+���C�����^R����{�)	�@<j�y�]�%.�ƖA��/w��I��[8rE-�x�����ɱ�+R���S]b�EC��:��8B��J��l�W� �*���Z|#@��˶#���qa/T1�=�>�˰d��?T�qt�)<��n�ϥ������y&Q�W���E(�t"��0_��B�T��U�R����������.�f������15u���Z@g1@��*��18���Ao�#���j'|a���*u^U@|��C�m��;.$���p��M`|W];�ҀC��E�Q�r�n�����֕��sn�ܥ��\��}�u�a)��	�N�l,��j������1؇��\�4�S�b��P�>�??�, �l�u��8"#�T���4>u�U! @�?,���{ ��%<����h˲fsJ˅�)@�H��Z@m��O�RU��fA��6�֥f<E�6�B>����T���ǚ$8�Z~q��Riu	�.�;9��`௅�y�&�y:���;E�����>��׊xk�암w�slZ�
�=��iAd
��Z�3�>��i�p�H���������kZq�)�$f(��C�����E�����&�G�s�	W��CPZ�A=)�3ȷr�ʒ�(E3^���g�p:���j�B��⠦�쐞��4,B�f�Y�(���/�d�yyxm	oQN=Dy	��r��|�1��Ψ4��y֝Qwo���B� �oqo�V�=�gcoޟ9ck��d��1K��9�~����u \��l�H����I��.�T�)������(,(��%ɖ�y��!��v�l| ��e�\4~(<��ǭ��j��LkҀ��f[9}�כ5
<���^�I�� ��W�ܷF�r�n�k��Ƿ����k��ex(�O�U��'S�겂�d{Pi�c>�����5��n ���	bj�HADj�=���c˗��|�Y`�		���!!/��Ab�-�13��7��9xS^�ݰ)ʳ��oH'>s!|��B����'�[�N� �Z�o.�Eײu��B���&���#X$�$@�|�O���'���	���O)8��[�PG�ɐ6�bm�1�⌸;��-ǖ�{��R��E���b���O�t�]�)�� �G)��S{B^�!B