��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�9zrv��^�t��|솟<���+Wz��ke�q;�"��������U9�:�	L��������27�u�Z>y۾�j �|W~��-܉�L!+�!X�%%�¹%[O��U��UA�^�n�v�)e��c���v��o6ٖFX�E��SN�M�8�SC�}� 8���8,M����{4
K���#�4�k}��#�.Qԟ��Ԧ�"�_6�>uo��2����~ �L3�b�q���g�~�G	�� N�l�<��}�|�XN7|� ��Y:%��(��6S!@~Q�UC��~�6�3�"!��v���,q�|��T���>\����-������@b���\�F jm�
z��?�����5�yBG�_t���h� ����1<��|8��v5��4*D�*͚�L�an?aYԦ��ؚhJq<ݜ|\u����r��h
�������yC����6�ْr����c�88;�2A����%"?���yD�ؕ�د֐Դ}�T�p��Q�;����
yͣ��Rk]�f��� U�z��'O<s�èp����&a�,q]5g��F������p�ڼw;��@/RiP�Ӑw����JlQ���������ŁZ�$}�C�!2�ӧճ���Yx�����bdX���'"k0�e��zi���˦+�Z��u 2�@2����zMs�,ڏ̰斻z�=y�D��P�c9�Ӏ��8�]���,�H����n@���O���Qj����P�"cŜyD�Ǉz��-�6�ͨ��c��O����:�T�!x�3�`
����ХK������͹F<
�%�=������O�^��Bm���\B�е��Lke���R��'�2��� Y�1�h�Y
���{_D��؅Z������ �@R�U�#�2w�ظ� ϥpՎ��|E |�j[l?�GJC�OF��G�*��!���wkL��z�Lr)�@�#�*+)�6@��^=�l���Җ�QHM��|:�w:U�(���
�Z�4-��Df�䚑�����6�>֦�H�/�{~�����r�;��� 5=����pʗD����Y]v����� fmp�f� rj��p�1 0�����g���������˫}�[��C֕��ìM��+�k��Fr
�� `�ż׏X�Q�Mz��
�@�T�����bLV+NѢJ���^n���*֍}��p���
@��&�-�Ii�{��e=F�&�bH���LxH��߱�,�?�ː/#kp�-z}�2���~�1t�J �*6-�%R�=�v�B�?;��F�Qi����C"��G e���l�Sh����{�}(��@q L�����j̝�Tk��e�7�؟S�7�d,��T<O��5���#M(R�JF2�ݯU�~��.QW"zRd�FzS���<s��f!yz�t�����=^���K�O��U�ȫ�=R�FlF`�.�\i]��H��`W%G��ɡi=�?x�gG�H�p�:��e��{��N�Ū��/�r����{���y�G?"b��w�W�ت'�T�����[����%�,���RMcߪi�g�h�2B�faJ�6W��jŘ�t5�,9����0�D����j@�k����P�*��숛��7G���|�C�5yL&��Z���N���ɰ�7sy��� �Dϲ[ci���b*��� ��$r�hؤ���aU�V1I�0����R�u<xD��H����.�j����es�K���"YT$�uڋ�WI��6u���L�x�Y��Ȝ�>c�<R�S)�3An�{��R)��`R��I��C�C�]�r�ʝDj��G]㲍D�%�"�x93Z�Da+�Cz�P��B�x{�S�K�"�ɛ����^��/�+1���E�=�֞�R�0b�(�)(��*ۀ�쐌V���MG������fC?�IYH���\E�)2n���O7�;����-'V5=�=��ˇ]�fTg������)�������� pt���L#�y�<�ɜ[&î�n�`̨��F���?�X�5�We�&�M[WY�,н�33����He��j���Ȧ����D{N&ÃXb G���nꆍ����E�8,3ۺ� �-��]�����_�u9������5�M�N��wYX,����%R��O�ɷ�*�����1]��?4c�/u��	��k�7�R�E���K�[Q��>K����1�oH���U�u�ree�;��� KL@	�*�ńN�eSf�0&(�+�-��$8����5-@�1�ށu���=��1*�>�-���%�Z����c �n�HHN�i[�)�y3N�H�dIj#�.:΢����Z��&��P�M`X%��`�<�|;_tX�|{�\�;�b�,�(��� 0�E���i^�B�ȏ����}�t��/=��?`�		�&!]��� �=�ӹ�8��X�6\��f��š�b�K^>Ǐ�`��jH��j�|��,i	6�B�rM�FR
̧�,����/ƬA�?���^� ���*�UQX�]��l��[���F)B��Ѣj�}��n��\h���b�cU
Po&�Q̔�Z�(.�$K?�$����4����o�����N����޾<K�K����cܸ�6����9�W!6��~����>�ˉ��������QO��K��.�ܸ��?;�0k��V& ���R�+��C����.Oq�=��L2���������ȑ�x�'3�6��.)	�LI ef���v{H�*qLɷ�lFa�:{-��7'đ�;�e��6��u��2��}�aӼ��T&�SctO��Jв.�04�D궆VW�ۣ?�Q�����nf��/:gpI[��Fc|`/0ߗ�"};v^2��H���I3,��<C�(��@ti��S�DJ��R"����ӂ���1G�r���eV���>ǩ��ş|R�j��V(I�ع17�!�f��XN��I2bL:�ʁ0 Y�w1��XI3�.Í��`4��`?2⩯�Y�����u�tK��ҕd&�)���x�`�����n��B��w�f@s[��U�@;�A`r�
!.���&4�`�=���\�l�Z)���� G��ro5G5�4M��n�O��2�����=>�������{��A�|5}�C�el��.�}%X�	u=6�̻=����v3��s�{fq��~R<���a/�?�P�j�&�INÖL��qٝ�F]?=�	��{F��T~;x`����ge�Iw���4Ve����-��Mˍ���v��Q�`���y;<)Q{��K��[l6#�ve�C>��љB��d�'b-��Fq����u^`=S���!0$nC�����^�7��\�v��+�_�����=��K�����"@
[@���I�6bđ�5󫺆���葮ӿ@��Ʀ-�R�� ���;�� Ԗ�";���ٛ��ū�%�7U���_�(�����H����KL��j�����B��椦|]�t�Q_q��r��|ƌ�I���6E�{=P4�ˢoe`4���g'������U�ۮ�1�k5?�G���Pi��^��ĦX;������I|�m�#)��,�6��4Ǉ��95A��i�}����l	��y0�p�xA�S��I"�{.j�$���9�}��~��8����joQ�'����N������^��C����"����y��:�ӋES�[: Pw
l�=��F/�h�]*��tU��?,~k�Z�*Wd,�`Y��^��cT�LRz4`�yR��%M�H���S�uPz
�����7*$�r'�]=�E����FdM��IϨ���>�F1��;�����D!&MV�!Zv��: ���#Ub+%�����#�)`�爔j�QMC_���Vj��nM�i�ψ�tL�̆�,z���2��Β!��
��L�·�S�8e�o$���b
��_�$�n����e�H������]��	B���c���<�����u�e�D]d8 z�uN���TA��$�"K�p6D3YQ�����
K�~��&Ȯ��m]��B�%ߘu��Ġ���=>�-��36LX���������έH� #zO���bu(�u|;���cn�zX��>�D�Y��8S��4�5��jX^��D���e��v�2��4H^2vk�;y����ڡ�+k�Kpb��l"�WRzp^��� ��d��CȢ���<&�a^s�%��ιװn�><R��w`��M�s߹�F4�F��X����|8fm�������k�p�j�.�`b�3q�m�	z3�'/����||��]]w�p@3���vM�a���{���������)p�"s��Q�j;��l@��/�����F��}�Gh������?������L[���ϰ�4��w�s|��z]��	� rN	��S�)�uď��*�+6�8�K̈�PCB 
������˚Z[֌o��:�)�B�?��ȱ�dBB�Zd~�6{�BJf����#����k$6��+���<
|�]���E�a�f��b��ߡ��^��+)̢Ιj�	��a������.�34x��%<&��)a��ka��Is����0��~�^0�|�H�96��L����{
ⳬ}>KG�"ة"���[��ՙ��@}3}�X��E� X�x������[�J>`���Us�V꿁4��w�w��v_Y��
����~��a5xl�+lj�_�����W�����_�˜�,��+��g.o�Z�a�n�/��ĝGC���Kk �#�l��N\ބ($]����n�v����1hĜ,-��>Hs�G`fu�Sr)";ғ8�����,�d~{J_�ףҭgJ�e�	���H{�r�T��x�c��CWMd��ax�Y����4/e霎�E�I�\��66*]l ������I�'��ku}w�V�h8S-
x�
ەZ���Q�h1�eI��k��x˯O����sYѱ-l��=�c?Y��r�W��|!�j=Ӳ�޽��Z#�.��s��T���&�,>I�ϒ;$�R���O��KXZ�"��1�c+s
$��8�-]b�m`�Й�+�m�����5�q��ڦ���O�E���Q�{�y��qo�8�T������Jb������y�$M(N�GTܟR�(MpOR�-��9�ӈYm2Om�
��2^(�����[%V0`1�&���c��.3EŚ��.�����'t}m:h�B��{"�����MZ6�|	}O����d�gѪ����5����0cN��j��U |tG�J�b��5�b��-��V�iA�pt�k�K?����Z� �iy�hb.0�H�RS������/���K�R .���p���9�[���(���ALg�$��y�){�iϬBy����}Kh�4��Z�pf�x,7s��L�钙���
'��b��F��}�VE�B�!%C� âC\��֞]�GQ}�+�gW/����5�oM�p�\��޲�Q��iI���� ��Q����Zt{e�/.���d�`��Z�̇W3Ed��b��+~��RB���� *�Ț�J���G��W���-2R�#��d�}㧔�Z���[�aѿ����ہ��i����Xqa�e�#z�f��]�\AMLݖ�M��G���j�M��Qݎ%�9������r"�5�ߠ������2�5��kwF�I���L�q6�̨Σ�M�5L{j�}(P�V�sE^_���LS�su�aZ|q��m�S���O��C�z�����E�{\z���޲��wj�n�g�k �"t���+��q�D��W jϡ.z���
�
MN���ɬ60�	�ѢS��R���[i"���g,�տl�>T&������]_��t�����nj,�3��ٚ+�1�`A
8�g_�.D����{J��:rb\���4�{:ɑ� �b�DY������E�"�.�h_���X���]6\,��Ů@[����x��8p��4�{%
�Rр�N�IŒ9���'\m�� ~�<A���3L|�w�D�@:�x�Uj�S_����פ�f�֑��K��٭e]�5y�ҸB7B�9:��������u}b�`�h��#�Ұ,�&�+vG	s�X��+;��,��W��8!��\[�{��N��	�@��?�ӭ~�r6� t ���%���0�.{5]U���i�S�3��F�|ۨ@�aI�tA��ǹw�7h����P�G�U_���Gj�>�m�Aj~�DG'�ō�5�Jj1S��Z(w�c����O�`�F�,�]F��#Ҷ��0��}h�	��T�����������?~\���օ�'AL{�F&�;��je�x��h��,T��.���4�j.��f�}�.��F���	���ro[�9U��l%��5�>��k~�����0{3#��[O��$��^%\�A��|�~��K�Q�k���G���Z�r�I��#�}dQ��g�D��3�%Y��ȳ���Y�$�嚉������|�L\�&�r$���|6�#����,V&)�`�^9��m���Ӹpg�B����߻��l,��(�]�,���G�%H��e��h`���^I,_�uY��H�}� Y�i�^��ǉ��a�!�r�r������Ϊ�
���S�G��,V �o�(W��L�A� ǅ|MBq�,:/��eբt@�mv#΁3E �y���5ܿ*���*��Iy��X*?�E�sT�����"����ٷ@���Ń��vV�Ǘ�.�-��3��+^�'v\�)4<u�&��!�F�PW�2�.�{;^��ˇ����E��SuZo���}+���vc����,��m]xCg�|M7���4��S1�7g��\a�jaAWed�+��t�iZT�1r�O
�p�mޜ����S$Z�؊�G��~o���,x���&���_-l����q�,�L7�-z����v�b��E���B3���ϫ��?�W�}�<�qs�h&���*	�ϬЬ]�č����_�A����3�����D�ۓ�vՃ1�o�*˵��vY� 2�]�h!��@��s'�h��ˀ^���1K��j�ԗ�p�s�	�+Տ��u�":x7�-��&������(���o�&A]zX���|�HXFx��'T��葹�1�g��s�����m���
�'�S[�����9�7uЄر�w�ԑ�9�����L^eia0����q�l����<���0���-��T3�vf=�3�U���ר�b�5�r��#�C�i��Q=x�~ζ\C?��"�}]~-���g[�i��"L�����"	��Lʺ�&��.73��J|�㪥g(S�ݳtb�$�=WC�(b�[6mt?}�\!�H'f��'�r:doPpA�	
!�ʬPwЇ��-d�=	�9<ˣ
v�������H�$Oc�F�		�O�,_F��=W��c��n���#����x\VŨUР��L��aS
�x��C;�g�l�`����=��� 1�_��Յ�t;$b��B�w����!-Iv���{��sW$wI�j���|R���e��0�iL�\�Sӭ-V��FK��}؃�=ν�~�	qR�w�@��6��H��C�N���e�+��������� j+��	�����N�3|����N5��g��)�E��2���E� �	NG�?'�S���?D������ƀ�C�%�ΜԞ���l7݆
5=�i����E��{�=�AZ",�L��3@��F�k���*먦�b��yw�"�\�%)�'7�ⱔ<����P&$Up�k$��G���W��,:Le���&j�+7�Zx����6����2�Uk���4��9��<�������*o	R��'>小2��jV���9��TBI�8
II&>к�L���GY�Tqy-�{�~l�j����BoGR�� ����s�{-�G��Z����)/����E;k35��{z���?<�%܏+��=
�iꮵ$p�3�͎N�^���,��k��`\��moP|Ml	��&�-��_w�1�Cj'��!7�B.�R��g�L�)W�5������_�5�J ����5��j�v�}Q��o75��8w"u�`���-�J� K��&�	�
�Z)�&מ}�ʁ[E�6[򧚆��~@�]ؿ6m;tU��/GS�[�
�Ҳ���i�w@5�X����	D=I���f̤L3ng����Nd�rKS�$jur�5ҠnZyPua�=�G�I������ROo������F�z��I1�裓��
|��f9��B!}�eom^|�eY6��S���V�'Ql*��e>A������A��n��n��zV�^�d�lN������	8�ί�ic(�Md�]Y�KܫT0n�G	�J1|a���`P�P��;U��s��X7��B��_
/[�\��U��,�%5�t͐>�I_���Y\{��������_�-�>ySl����#i\ٻLY�מc��a	��p�'�4w�׋���aL�a�	�Ǻ�g��Z/3c���37ZB�7�͆���)�lys_�������xs��|b\�mZ&�߱g�e�A�]�P��6��"���lK2������W�}���;�{�Ǝ1!��tf�#�F��MXA4(�@Z!��6�b�Q8�	g1�:��FnJ���c>���ͲV�7r
������Ga�}�s��C�?\��W�ݴK��2�y��RE��Z���$�;�����W�\���ܽ�Y^��B�KDN�Ѿ6��9�8��y�/l�>(�БǴ�Q���DM��-9�+Xs|P�֩�ρ7 �{��@��zT�yo��H��>3������Y�_1t�	T���N����A��;:�@Ua	�Z�;x4.��C=&y(�8��<6�L�1o�R�q*��p�����Tݙ1hd<�T|�n�p:��`)�mħ�%��C䂠�jr����#?����A�����z�錑���4R��QZ;��@eU�3F=N`�\�ݤ��-��v���+������~��	��"�Ȝs�%L���kL���*�ژG�r@O�|ܘ�Pg�cP*�3��5����%���0�(���ۧ�QKxp�y��[Ζ�E�Q9d���(vm������y�3�f�A�i��;E��SY=�S]ظ�Wr�ds�$� 5ӚW���ۿ&��$���αG�5��Vkўp!	��R�p��1)ڦ7N}`��cF["�﬍���=�Ø ۤ�2j%�&����4ʹ���l�8
�0�vߠn�Xz��˅1��XF�r��v;:R��T�l%�f�%���]챍�0�Ƅ�W�^��خ�x��o1�&)q��������(��v1S�Eq���鼲�C����-6�Z�*�҂�P�f]91L��$���^�`�7��n��ĢY��Э%X2�&x��H�� q>�T~,0�>�"�t�:��U��{��B��-�I� I\�$��24$�5v���!bH挨�qX۞ �V��&�[�Y�8�� �}��7�-��zSF�?a+�vh�9,2�7X�g���Q������[����ܶ{k�X����P��Q�t���L�,ʩo�H$�c�)�r����ΐ�q�4������$V<�����
O݅�r� �5�X��w���*�h���W�fy?�8͔��Y�eY�̱@������-��I%9k���X�6�M �'ƞ[��U��:�o�[|�mc����I�>����_���J\��;�)nIn(W���yiߜ9G{T��ú��N��)M��'�>�fkhF�C~�cwN+*by��!@l<H-��b�á2�-�^�W6VxqW��A)��Q0�D�
%���Dڻ��s���<�=�ճ��h���/5�r�ѢҀ�N֩��|NUE����Z��Nt�;����Mw��O�OP���;✺R���u��M��p�{�sZg��{��s�;�98~qSsN�|�B�X�_����q�^W�y�$!�#N#S���cR@Q��kl�����{ݤ3ҟ����Lp�O./���d�鏊�����M}�N/�jo	;���jv����(D�� <\ڬW�%c�K�>c흪f�<ՌBX0���D�v�y����[�	͟��P^LzZkE��B��T? �l?fj#�	���ry9`����w�{�z��J%| ��<4�;q`�&���gU�׹�9�ν��N5b�VD��ԯBΣ���Vr* ��Xq5T�����˘˻���J���C(��`����:>�i���L�܄\w"�yL�"���nľ��g�Q輽Qd�@�)���J�Ӽ�lஂC���~Y(���(��$�c����8keGe�(H�
����)�en�Z׋�l6s�B����,[���-��q�G���742����8��������}��V"��!�z:�/�9����"_A��r���D�`v��{?!إ���"��� ��mmd%�	�I����0\۷	
��2
�|8�w��T2���t�3�����8�U�[��^f�Lc�9���w�J��Qz�i��������/Do��}���k�����c�0�1���<%d͚�S �)Yk�����V0�������s��Q����M��/~0����KS1�|�c������ʚ�� L�2�Sa�<y��z���N��[��R	BP� �n,�;_^�g������K�q���H'��WU1���vj����P����)�C&���؃\PŨ2���ˏlA0�U4-8x�;3�6>�[�V��%r���2G�9^�z���X���?�߅y/l]�Ȗ,��<��p�O��t�,��EjS�-���#�^���n��������V})T��5p�2U����Rp# ��Z�趒 �r;`�Ě���%Rɉ�hU�mQc�8�t�7t()�����m>��y.�}k�J�aIG�p������f�����*l�eF	[4?�o���I&:���;���5)?H*ٻy����ȴ�v��0,��-�mn.�K6��W2R
�6U��2Rɞ�P�(�'���C�����zQ��
,n�q�g�bk��N8BB/���[����r������R+.T� �/h�K�?�z $'c�.��r�z�fH���0<O��/4�
�ػ ��h��5t��l���W�����G�,�84��7�:��͙g^-�_�b��tϭb�4�}٩�$�t��E��y�;�S��Q�z�^�1��Ǩj�cw1^�o0z��
&��U�-\�\�*>�6��JT��Β���؜�y�Dh�v�N�m�ci�LIKI�V҅ޫul`���v�Z�R��[r^�K4��3�B0\���SoA�3J$��N����??��"���O���{̻�G@�Z����/�so�0�J��]);�����%��y�.6���0��Vx"��o��L?`#���ϳ/ۈ�̷�5<��M��t�H��Zi���-t�UAm�ʨ�7B:x+[6��"����q�u7����ջH�ϖ����:�&U�H�_��Z:�F�.,o�ّ�G3X�!�p��Z��Z��;�u�;@؂��v�?�#)�H�r J�-sg~*�.%L�k���rk�����)}��]��v����	���b��~K���L���z*lQ�϶�D�b��>p.�ב����3��q`��5���}�p�g �p�plC^�Rf!�2���ۓy�T����>��WN	��O��;|{�|6o�,�ekө`��s��{�h�+}��%"�;�޹m*o#ȑ�o'U�;-��_�h/v�K�m�k���f�13�շ�H4ce�h	H	w��v#����ֻ��=�P��æ�3�}�,��YI�a�b`��Y03Ų]P�����箸d�?�#�r>j�Qx^��%O@�$˶2R�\`�tIj�4�O�#�[)��j�.rm���ʣ�X��^&�G�T��WF w�7�uu�fh��_0����?7��rP2l�:�a8�ڷ���p��LG���u����sڗ>W}DS�D}`�7 ���,X�J�	C��p[��\����V:�������.�fa�W�_��V�C{{�+��^jX__�T�̌����C���Y:����U%�V,�C���#�mL���Ѹ*V��.$++sŕ� 뷇��M�F��@��>#.�^Tyw��[�6!R�{1<��ÑIA��3l�c"����ˉE�\��I����]k��]p�w�<��:��{��L1`�鿬'����{���u|�P���B�H�N�A�;�`�ѧ�4>�:�,F�5$�@M���E�+E�? ����L�i�ّ�-��׏+2�#'2��5���z8m���Uc��qKo�Zܕ^��ã��g�+� w�ۀ���)A�m-k����;��p��O���4I����9@&&J�Bw�x#��U_r�᥋?B�/%pӧ3�F�-rY?��-���{M�g{)DL;��Y+"s|*�~'T��,}%�\1�]w����4�$�Aǡ��	��̠�ԑ ��+!ge1��"Y~��6��-+�Ơ�p�W/-w6�=v�'��0BV1�nJ��EPIp Ӑ�{��qغ6؜$�A��~��_|4��N�n���:�,��f�?Ѽ����(�2F ���fƃ@W
u�s�U�0[dab��IZL�׬M},?���JW�����E�:�Tz��2'�� �h��RcB�K<���-D�KR�:N���!v�[�׍�̿��!�S��)�����$M�`�<��O��f���#�8g�5f5	��{ںh��x��8��5\!���-u��F�l�Ph�0G��"e	L�gK�*���������E���_���@H���
S֍�$�Cq��G���YZ7���4��?�Js� �mv��a������)��i�^��l����n�:�.�˾��p�r�u<������G� ��ǖA��!v�1=zR��"�y����8��諴V;7@@�G�N�} �y����� ��Q�GSgué����;�E�hD�/�K��q� �#z#%lb��I��FHp9�)�ϻ�u���lͦz�s3�Fi^T�B)�Z"����ُ���ؤB�C�,G���c�I@��P��+�I�Z
{�
%���W���W!��*� ]�!���%~���iD<28a��E~iQU/��B�0�0ISd�R3����X�`�%"�B�qۨ~a.�^D�-�I�d�l!�
�����C����[bb5��@���V���w�E*�2������9e��h���bc��8��E���h$���)-��FS��ԫ�31$t���z�{�HH��l��I��\��lW�x�h���&�)�p!�iR��c�s�]���t��,|����~�M?��3���9��g�V=,C�e�7����,@s�xL��������ȟ<��