��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0����>�P@�:���VARiI�sDyK&��+E�,��RR8&(�-�`B���#����0��>�杞��9�OCg�	�@�p�����(,U$��X���࿯�j~��Ұ��y����-��B��\��Dyy]`\�M����$���P<�x�%j��q~e�3�B�q�v0����3��8��
7ǩ��K��I��3��<<��ٞE���M� �I[]J������T�W��-J�e�����GvE\�:ڢ�7|Z��(�8�.�r]R]�O����Էz+��o�%N;�B�Ze�KŐ�����	-�F� �jds�E��.�f{j��|�4a�x8nL�Kj34M,�h�r�<��o�4TO'��&EA�m�z��y��V����b3wx����m%1�ڢs��A�9ƛg[����\�#�����{�gCL�k����U{�G3M(#9��FAjG �k�XدEX���ecb`��$��hU�E�c
�û��ԂX�p`�V��}�ι|d���kh�7@H*��
��d�V�����&�����@s���h��X�u$�ϙG�\+Y�./;^aF]��S;&��gϣfnC%��,�d+GK�xT�P�����[$	q������/�h�tϖ�+�Z���&D���);��J������ySU���6��&�X9s_�mDo#'Q<��X^/��
:O�tx�Q�c��7p�֧W�tJ���UlG~�mݏ��}���(��ˈ�&���y��M���������,��xF<�Or�S�w6���ԉ�T���ZƁ�'}�N,b���@@��ݰ�������;e���#B�N�eo6�sP��R���=���j����B����Ttd��lՑ��]I�¡HM�ޠ-;�ʥ#�ٙ�&�%Z5��Y�s|W��|=���d!�)ȁ�Ň����)��.d)����*�tfY���$�"Ig3w�P' <�����vx�t���tp�L%�1f�K$�qc&�4�^�����Ou��<���3``�5��6+m4b�=ZL@�����4<K~z,/��v9~�tD%S���+sO�d$`��u�� L��� �:�|x��"z��bd]m���WiwS{��y�;�����2�Ǥ��
����	
�s�BŤ�Tهud@�>3�2�Ԡ�W^_^���j\*'� pŎ�8��e$��H� ��F񔢄��|��T�+�&z��%T�'e�JMS>��,^.'<}�^�>���Y�� �cN��u��72�����1�;:ߦ!�_�Y���0i��I�J����䨤TB���k�z'4���S(D�[]���W�8
} ���bK  jh�A���:�ټ�~�$�ivh�T^]�!ՙv{5��U�f�`CQ�����V�1�Z)��C��G�P�iȀ�D?���R�#�ھ�*��=9���K��hK��%�G����X�i����!+tH�=�o8�$��J��H`ɨ=,��<e,Tn5^b���0�:I��%0�M{�:������U�n�����kgpr�,���f�%��������Ө-yC��-z��V9����f���=�[�d
n}22"�Y'�i�#ʃ�w�a���=�t9��P�#yS�����#t9��ё��k��d�O�
e������y}	gAZ<��{.�t7��H�W���/N@k~6m�ЄQ>Q�Ԇ�Ntw` ��
o�9Ы����:��Y�c/](�ʹ�6�X*pЎ���k��>$E�)4K�3���v������_��!�`��USeqe�I��
��Y�zUᢗ]�L�UǮ&̍��i���,�`M��Tp*C�8��NQW���r�Z+���D�+��C�?���k��k9��?~���g�@p/����pWյv���Ha.|��Z����<��:�j8�0a
�B�s�'�56�!y�wKsګi4�E�y��hi��%!Q���pݣX�������]�8�)�Uc-3E�Ĕn�K��z��LJ?�(�ū�>�S�m��`�r&�R�@⪾X����&*nWl�c��ncʜ7uw�w���Sե��׽��iF儛�'����L�g�C�A%��#� �J2^�g1��}�kN����̂�#������ɇZ�>*���F���<J����v���ޖ����ӃO�����TY��F���o�v��f�)7���}Jf,{��t�:�>A����ko+@�ov�Em2���@AER�̇\3�H�A�֨Pg���g�P��$�� <c3[��56��o��8-uP�{˯�B��Gz�C#4�zK���OA�
lÚ,rv�Pڸ�dm`��q�,�_�Dԧ֒���PY]�U���b�	f��.��i}���2�`�Is�#�3Wo�y0����Q���<,�A�D8�cښ�����ά�l7��Ė`���|��kG�,R��( ss&:/c�G�i����iYŒ���T�f!]������3���L�./BO!��љ�Y� �M`������ñ�-SR��c��Ú4O\����J�y.�G����j[�N���^x;�9de�d��$���il{u|�s��z�7J�p�0~�9a�܊v��.��
g7��"����u�#�j%Q�:��|��!R�v��r��mL���MHꮃE��[��$�!��s=�@���z��6B�v"J�7�v�����U�⩘[�C�J�e