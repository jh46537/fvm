��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�>��,�t�Jq�%�qr��A���/4�HRN��Ί��w:p��'�˷34��>,'2��q�B�'�ri�v��B>�k����2(Ahb�I��Z
9�-��I|:$�a�^�^RB������������i3���k�����Ԓ��B1��X�}�%Z����'z�_�x64mhOm~(�� '��U�B3��H��.�6��K]v�(��`ჸ�<D������Ö \��j.o�ShL�v5��SԲ��z�өY߫�%��?�'�����"��@�_���B��
�k�7�S�b#5�	�9��K��b�3��j�BM0� ��@��b"u*C���o�˸�V��v�$���,ް6b�?Ph��lL��5�V��am�!7��!A{؂�ߢ3�"=4�Ct��B�b՜H�+O�X s�ڼ�R�O�Ū��������2�p��>�Ns�o�X�	(�!�ߊk&���	go���Lm"Jun⵲�^3!�@"� ���:�+u��5M!0 �d�a�f�c+��ހ�Vg�#�̑Q&.[�5�i���עC�0o�Q�u��^&\=λNO��l��b�5�A�wH~����Z?&6�����3�O�����ֱD���Ff�����X2S!$���
y*�	�0�8z���r+��y�!Ԫ���\,���������({�a�K�f^&1VF��^�+�݋i�%���%v�x���>`i�gG1]�����g�3I�/���H	3�?�E]�8�Ph�@1�\A�N��r������J�b�|-�y���_l�I��r�<�i���A�z�C��,��lrWp�R7'��"{l�-
!ۉw�n��M�=��Ql^�*p6�58����-���Ow�Ӏ�/�Q��cy��bh�6����K*^��~��c�^ȿ��R��O�\	�b�<���X6͘/�u���Pzl�ۭ�-P����Y�˼�~wkE�;v�*�;�vtN�Up��s&��5MD�]^�Έߞ<�9��;�D1��Ć��y�^va1	�� |�H(L�U>���jQ���R��p�����=&m�ߑ��ه�B]���7� ѻu��V�b�:o ���yv�ȆW]��:����6��r�ԑ��3$�?�v���Rgj�:O�f��ܿ�;T#S�V�I�ˢ:�y;���']�)��,�
ZZ�����-Rw���$�R(��Uy�¿n����󾇘( ĉh���]��vX( ���$/1ˬ!�ss��{�XH������>}��(2)h�����e���K��f��9��o�Ɉ'�p��X<��U��(�}?��3>tn���b���>Nch�ܥ�\jPVᶰsW��N`��W@�s5�����%��P�-��&��X!>�u�<�{)	6i/�BN�6��޴\�-`�4����]�D��"_脁T%�� 
3q��U$� ��pҌE��5Ǚh&B@/XR�(��ڸ��2Ǒ�Y��R��������!F9�Q���1~&��g��&7.��7���X��d��+aku:�/�2��H!�@y\�u���Y`�<����M� ����F�. ڴ�&I��1�B�8�%��a�ݛ�mv�\�.t��᥎�0�Gw.%f2�1�n�^I�*
��b'�|s�Jq�9I�eL������f�=	�Y��U�K^�k����
~�:�����=`lj(���`+_��' ���3�L���o�� ��*���iw���6LK���hn}�TE}�F�U����Q�LF�&����o7lCt��/�4_cs�ܓ�V��p�ސ�������h|X3`��|XU�;�6�̭�M�^YQ!�0�Ѐ�<�[㰑�!%��E��J��Yb�m�؅��P�]�^e�z�@�ܵpo��>ty�Ex�^g�g�A�ZM'���*���A��K��:�����s\v��Ģ��f����)~�uq:�Kh=	T�H�Q�@�N�^���$�rE�x(��8�=�k�(e��LB[�J$S@Y�oID4���S��]�'�J'26�	�o�1�&��JE�d��_��%��T�8�m��*P-
�&��(M>���K���D.��׍|���^��F0[�s|��8'PÆ}��0�@e�|9��tz���~�-��Β��Y����=F�$/O[&K��99?=4c��?���|aM7K�5������\|�:WEsb��>����R�Zk�4@#�H��3�W����4��	Ĭ��p׀�f��0'�������`���.�ɋ*�] 8����<���N��6�z�qt(�dފ=E��5e�cE�[Y}EC�K�ri��K4X�y�{A�c�+yk)���^Q'�D^)���4n�YGܻP7X7�e�:fs�@�&�1n��L��IR�Da��TR"#WsͶ�8|����_�B�V �<�%wKy�MZA*��o�*p���<�[rz]Z!�H+a��<��cº�D��M�u�-M����;���8�ĩA���E���dXl��P��?m�h��t(��[�lA^�ԯn�:Є^A��} ����5���0��R��|�T3R��%_���0<��)?C�����*�-r�>/D;�0�O����F�OD>�h��z?ӽ��P�kM9~���Tit����E2�?�������OjĕCf5�4~?��-Ԉ�u9A�5`��בW^���v�7J��7���RS�{�H��U{<!��r�Fc�� �u��՜a%#���}���r$�|H۾o�0�'��jJ�B�p}�:Κ�)�hkS�93�/���{���39��~�e���eX}�r0c��@��,a���{K�>=4�d:�f)i�/�*R�EQ��;])�H��݆?�F�O�>l�Lg���{=�0|�1�C���g��:ߴ�Yp�C��#|2�`S�5\�c&���U���xא�5W:�ac�|��>�Q���>�l�#���DG��y=��ɦ4�gƅmG\�&�	{��[�cb��R+��+��?��lQ��H�N4��W�#���f?r(��B���~IaH(���N�5]Eeqh�ok5m��4vUaśӥ�2��F�a�:�1D(;Iv��u��7 ����9]�s����8 ��_ԕ[|�����WY�z�����f��]�)��U��O
x���.Y��8��W��㪝"[!�I�C|�ϊ���^���ږр�z��mŧ�Fe>�J;�T�I���Eg#F�N1�x+�a �U0�5�T��˘�ڊT5zg���'��X5��^+!Ed���9[���Mm�jxO@�s�ᣧ#�n�2��nviXLU��K�����$��7~h(���zE��S�@��ȋM�{�����O� �}���(��2�]��EJ��ݣ� ��I�0���������&os����(�{F@�f�c5L���U�Ga��u��
���"�,�7g�̼/C�
���H�C�1�u��b�ZA�����W�6����?��WZ��v&~2噒o�O��r���}�	���ׅ�|���*r�|Ծ�*�$�C�$���'�fQbu�TC%�S���B�Ot �E�^E��e��)>L�S�I7@D�q���X�ܧZ������S-���V��Y��C�܈����=�K�u�=>\!ύy��i�@��޼R(-xK9s�}�e����%���a�t������,���>`F��h�s��/E�Ft#��f.��%keɎ��$?s��	��N7��h��M!���!��^�@}g��S@Q�q;É1��j���U�r����,ܝ�œ}�^������ �)R�H����9.uܡGm�82�Ԓ������3���X�Yd$�E��X���ƕ=իI�?�����t|�0J��@f�NE�'V�7���#9�>.�f�m���[5\M8��c�K�m��]�p0p�,)-�=�j&kA�IG�'Nӕ���?n�]uf	�0<��LZ�Ɵ
�U�D�s���^��@��K��8���Q���HNj0K�7z�1���;lp��;S���tf�f�*-:)�@�Ĥ�Vm��^���0nܳ	����a�b�,�Z��<�pd�K�IHM_��#LD7�b� �%�u�vL�MX��NT�:�OY( +�@<�L� T���/{X�.�S�^*�Th��Cʭ������ᗎ]CYkRN
���s�i�kp�BM}�}-���C�r������R&R���\WSlXks��7�ɀ*�&1�Uqyk⮵N9�y�
<�"��\��5�����ݮ�"�G(x�l��R�m&w|�B�MT��ߛtaBʥ�V�i\~��2�,Z�\���Y�E���jAST�9�.�^�jR���2�s��V�\7��we��!��,�� �M�L�$!q��٤����� Q����4u  �,���d��lz$Dk ]�[����a�R�9��5��u���L��ಮ�2!�D���K~���>�ϐ�QO�^e环*o��:�z�L�\P+��[VPB�n܉9ļ�ܴ���m�]'^�1Ew�KD�l�LG��0�P�������x�]�, �уW �ǻ甀�ku��������@x_��\������xgh�e0�a��d(YD�Dm�脱V���CW����<��}��g�^�QG����Ϗ�9�Ѐ(�)�XG�{3��m��tJt׎+K����?/��6�^��2j�~s<�=n�:n~xt���qH,R<�I>�Dz�֍���i�t2�=�+���碮"m���G�AEA:��^�d�|&ɞ�}��x��$0�B�I���HZ�&�jjvc���\t�V���J��bL��Ԉ��ҽ9�ȏ�v��)IT��C����m�3IH�#n6O����ҩ@�?vO��6�9�������*����z{8GW�N��|�π��NtC�+�y��lK�#�Y��ժ�`N£'R	̢L��M"����%�xW��~kE�)e4��=�X�e��W)b��"�K�U7���R�@ޮL�j-�%G�V���1���t/G�����Z�p6m�Y�^� ?Wc?p�'��1�Ի��^��@��Yx��K�^�~ߌY�G�4A��tL�!�.��Y7�';����j��=��I����ڗ�4�l߯粪��	ŉ����(���ǦX�����ɚ�4F�5d�搉��.������'��"K�Əg�yʞ\$��e9�zP,�kT��b��K�M���隂�L{v�
k��J��%e��V�c�W.}.[�������B�� h�՘#��c@�a�u�:���C�6���^a�V�Ƅ�В�̍�(PrP�f�Z��?+x�w���R�#n��t��]"<C��U�����#~:�f����K;��:
w;dy>�q$��=��h0��%��[���o�0:Z�ɗ\h\ ��i^6�q��J�1ڡ��py�J���()Ux1ø�0V�L�����J�0nj�������v?H�����w�+p��lp���@'F���)�Ẃ����e�Ɨ��j~M�\ b,ԓ(Z=���;cZ��;Vs��͘
A�>���{�da�#ql�
X��Tή�l�S��������&&r/��9���"x}���|+ ic�)���]OԠm�W�U��UG��x��Q�a(��AN��e�f(�'���#���>�p�F@:�8���ʘn�h� ]�n!B�3Խ@�i�=��=��?�����Tb�cK�?���=�j��=&9�,ײ�	��Rz%TA�SXiN<)�_�]о?{���@	r|�M�ԭ`�k��8 ^j�Ÿ�i�2��*1Z+�[�=�ʿF�{*���oD�1�A���:4��+��}Ww1�L,O9�eEyY�l�,Ҝ{P�0A��
����z��=���S�t3�e�[DLI����5|��fb/(��ſ�T�%E����-N���wfN����&���e�̿� ���tn���wS.��f��>E�:�[�̴�Z�o:� p�IHIŨQ��>)@%��v>��]��8�G!�շ�Jmq��Z��g-ꆄ��"4C�!M�����HwC�������mpW)��V�$Z�Z�Y7�=�6��*.>B��jU_>n#�'���U/k ��݀����d}QZ������_t������Kfg��n�	P��ܸ�K=K9�r�����sY*O,aGq���P#�w��u��܈��~s����tUw*�$�̖趹`�R:p�όK�4����]~���v��Q�}��n�Ζ�]3� G���%ER�aZ�";�[�dV١\;IA�Ɔ����{1N�@_�2�;���������yN0Un�j��Tx)'j΃^�{kua�0��
<a�^��l>�@O�}׿3ȓ�%)��s+][�y�#G���'4����|`i`���nz��L�C,7ˁ�8�+�E�6��&�C���u9��s��X�E���-k��7��$@�8��87��Q��#�#j]Ƙ>$�c-�+�}&w�7��RC�B�F^I>�>xo�i�ޏ�={�HQH����4�{Q$� �CDx�5FG�������"�7n[L�h�%����f�3=��Օ��d��G�i�-���]C�.����V�;���Ո�:�自*�������˦�r���'�r���]T���	�.�OM4uÌk{��(�ߊ�'Tc߉?��S�p%�q/��ҁ��M[���@�lCL���50?��.�g�	�\K�bO�����0��>�e�|�X���M�-�M�P��C�M������PB.�v�Td(�}k[<����+�1jJ}Z!�M�}�v�YjM� N(~as�`�~A9�ah�U\!���B(���o�Jo���L~�7W�n�7���� v�SY	g��a���6l"!��%��z�D���&c���$�Sɿj��=�h�IS���N�l~W�bI��MXϥ��6���ܮu�{%ư>��;�@"�1��JL�s��p�)	�B�`�ˈF�華"j� W �h�'���3:<�~c��ZtA.5P�}<i�^��s^�o�r �i�(3=��<�G+��V�DB 3����_n�}[��@��B�g������T�$��t��f �G|,|]ä	�(����+A����K7\��s�)�}����_�%��%ji�\�������\� ���T����
�%K���]MuV2�0!"�1�q������Ru5\
�Qp�Ӣ{$�=I������0��B�P4 �q�$y��ld��G&-г�$}+��3��J�ԩB)�<��'�F6G��Z��Y_�(��o��U�� ��W�|�PT�l�[>���D��!�p��o�A-ռ��rs-z�/ ȷ����&A�5�$[���5e|,_�\�kH��d��w�I���i����c�d&mw{��G7��BK��)�E������2���Lr�l?���v���CɅ�%��Ҵä��͂@`�O}1�=�p��ni	�����6H{���$�e�B�( ��f=�[�ć��>AⰛM�r��|�`���*�̼9�������T�y������C��aQ�ͬ51���Q��/���jE�J�e�x!
�z:���/"ׄ�XqV"�E;`��a���q�F�8����#Ql�Tն���7�öV�9ѳx%o�5>��G��^ihΩJ�"��ޥ�z�3������|������SY�6�d���?Z�dM|x#��M��d��K'����r+�s�0�b\�=uah��@ёfM��Õ��ڳS���ý_��BT�G�1���S�5jsI�w(�<��f��.�H��5�k�*ѵ�t̕E�d0���ۘ^Ñ��QHt�0�}_����t�`E'�������K��s_Rn��E�7���gg�*Ks�
���f�hH��ZzԢ�[�u�7i��\\ъ���I�Ӵ�����mg"�R����Q�����*��#���7��X���I����P%�C�%�+A5VCXw�������c�;+��A���e2W���{��5!|�e�n
0\���B��(^��߁��*Е&���?��[q��MY�EhV��/:)��&�� :�Y����@0P��t��8. v0K����#�_L>9u�c�`�r���1r����s��l��1R[ �|/K�����I�!�B��4�Y�9�LCR���@֣<ϛ����H��/b��<�Qn������g�&�'�e��4.;m��=�I���jͪd�����,��"_�N¨pH�0����SIt��v�<@܂}��w�I�� x��q�U$5��X�Yl��5p�H��6d�N�v�zFz�;{�� 
�����恾Э4%�U��e�@z�\����B/�=�Ě�s��n�J��(*���W\H}����d��ai��#^F��dp���.��f�5"�Pԥ�00Kӭ��.Uc��,�áD��L��]>���T��S�o�)���kY螗�	��[(l(�}�a~w�c�Uf����^A7�U��o��o�D�cB2^Rf[!�QR��ޝ+�t�n�0������eW(|�%�G̧���1rV�˪)�ޥY
E4g('�ط�:���~mB�3n��V�1�!�3pC��NW�����E���G�S_���9E�'��MHᘁ?��j N��aF���M��=��yyJP#{ɣf��B�^�Y�!�'�����ӦNgOZ��w4�#{8=��B��p�\M��y��\
�E�k�r�	�t��^8M���>�t��K<��P��fV){�s�rN/�g����=E�>��n��P� )$��&���2��p9&̳��e_��s?�a�~ge���)fQ�E�=#H����eQ����	����s�{w
���%g��^
F�f����*2���u@0t	���m/�'�t}����� ���ʟU�<��Le3rL��h�`�|�C�x��
����g\x��ـd�i��+�S�Bͦi�ΦuU���}@;��O߮%t�D�7�uڤ>o5u8	pI�����Ū�M�V��5��us�D�a6S��=4�P.yT�V,2�>ptxIV�W��ݛ���B񤅥!y�:����q񤀥�(��H���#S�C�ve�A��8��%n�Q�V��:��w�߉���NY^�Mq/��_{�~B�y)Z���TٓW�����?���U;6�0��4L��q����ٲ����mB�vHH��F�c������B�	����\f
IY_��+i�	�����3���HG��%-9?�QX1;�{�8@��Lꮈ��?���e�h�W
��\��H�����V�����& �Vb~dY7�I��'��N���G2&O��+�!�a�����]�@�dɔ�m��i��v�@:�0B�&�^�s��"���uO���GL,������lj�"�f7I�����O��x�f#&�d�t>���,M{����JoA��� �2�.���C�R��kZ�q���	N<�ļ ���_��U:��rk�D�x�Wx|&��K�DM���1����o�p���D�7YNd�of܊�i�S(��N�WWh�gۣI�-V����w��2�nlQ�)�J�,5K�u�z��_{cp����:-��'l����q;����lո�� &>��)R"�-y����"�vѷo�}YאՍѱ��-u��O�K�WшR���pPA{j��8����9�y#9� V��A�u���z�	'���d]���Ͼ���G�0���}�#�yy� ��bK�����.��!��<�*Z0Q�^��RW����T���}�Oݙa0�28��k�3(ypK꜍�b�R�S�J Lv�u�]��҉��͂%ˋ��`����G|�nϵ/�4q��(�u����@J�A�M#�ΉXM"q����g�0�嚃��U*��y疕t�M�>��H���q�oA%w{����8�Z�C�� ������C�U�:�+�=�r�CZ��B������|V���b�_��S[�r��r�#�q� C�I���n�h��xS�)�G\�B��Y��=��:�s!*m.�� �崐Z�iOЎ����U�.{G�D���'Bd���l�NE��}�R��r|�T�v"����Qq��ު��������L�I�D؎i�@7T�,csy@��@0ޠ�[�C��p����V˫�s�x��mU�T^��6a-d��{�B��
y��m�0�*���$s�_�����
�̱Ac�V0�CL�Pu�o��k�{A��+�D0�L�>�`�}+�(�cJ�['W)]=S59��c�}��g�uP�֍i��s�ȉG#�����l����i�!(]T$��.�)#�|y��g��� k9���W��$kv�>E����c�"�F�8X���QhH����������gt����5��3�G��U�v�x_��z��n+k2D۳��#���6Hz��j���4 �(ۄA%R�S(��;n��mg�T��M�N�n*�'~�ݑ�LT�����X?�_��!>@po'���G��h��ex�v�I���0��LU�����^��0{�6��3��oW2��=d��g��O�K_pyÔL��<{�&�{��I���PY������;�$u�]�HÞK~yQ�E�z*��7�m��M�mr1���������i;¸�rΛI5ƍ�4.�Kz ���%c��`���ѤR4���ËЪ~<��Sp�uJj�O+�g��f�M���c+��������c�:sy�g,�UoFe�0"G4��[F�z#���x���l��6%��̝}�`-+0��q]�yX����+���L�sx��^1~���b��N6�=14X$�2.�ma�T)L��h,�%�&累7s�f���t�,Mh6r����}mR����g}xg�{��ߥ�|.Z����r/h�؄��f�Ƚ����Fw�'�@�?ن�k��v����z>3v��x"*:0КS����هD3vP��Ou=P���u���������}Q�7Y��3RI"��So���+X�嫯
�6
��Ѩ�	�y4aȍ�MWFE�g��ճ>Q�f>�'�z@��%\���BP)��E/M��+W�N_�FJO�bD+�l����iq>/;{5�_H�P� �ڶ��>��`�9*�+.�$>�����^?5��=�A ��LYPc+��FE8>* =�]P��m�YQ2*�7����Hyo�D��B�T9�0e:��_��:�ר��)(����b��T�K�n*����I�#��\��+/�eL|��Z_9F�S�y��{yo���P�2̛�V����|p���v-��Vq����5��k�X��4��Nv/�מӉC���Y|����s�T����v}KȤ�{�u.z�5��$��L?/iŚ��[��R[�����&|��s[�2���l���O�q05=s�t�.�}���"~�m�x+o����$���C��VVZ�59-8����x���~l�*G���%!�5�5�Q��e��}��ꇑ��B�	�A
Qyga8��B����s{aB�^��=���Y�ÕR+Oտ"���E�2Ƀ����w@	uV˩.~���\��Y�A�ѯ���	Z��9�R�fpo%����OYj^�i6�1���G:��|耦3T�2��x�Z��1k�)�H#��u
��B֯�}a�eҿ�?Gkz�����|f(�v�J�{��{lG���5V���4W�����N�b>��aϠ��U���U��p�Lc�ۯ�m��������,�N�r*�n�,��U2�/�b�쇙7�U�L�8,�fds��t�va[@ȳZ0�G��Mj߈Ꮉ���1FE������pmڲ�b�v`��2���༆`t�t���G
om�`�Tn)���