��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���q����f'����U�S-Կ���Q@	�Z��*ѵi��s���*(�Z�K}�7�6lg���T�����'m"�Hq&��m���^_���M��Ȼ�}����^b)ٞZU'�ٴ�������Wl��:H��`P�}3�RR�e�ǘ(���/܁�g!-�k���;�HL�
Sz��j��eDs�BP���	�[�����'�E�Tt�n���oꊖz,������..7q��~�r��1�0�T��g��A aBA�"N�~����DF#Ԍ�Q �2m/DuE.�Ki��fz�aм� �"�!e�Q�<V����9�VGv�jN k4���ׇ�ӕ!iG�<���O�o(�Q�8^v�vm�7���om�%���k��'�x�j���!�O�S�3#��>�c�Ց�B@]�����,����8PJ�z�Aǃ4IF�xj����h��������`Xή��a6U�0��;�YT%2Ă�X����m�m8ex%�2�ӑI��f�C��Fj��}��4�I���E��GQ��,yFgi���$��K
?�"�YT	�V�(��i���Rd��\/p[h����h�xJV�d� �h:<��4��Ԙ#�G��P/^o�	>��́D?����5���M��C֠Ri8±k�υ٦�%JTT�r�ΝYL�-��D��j�B�\��.Z@6����C9eRw��z�&/�U�T����;�VH!'��{zȴ��t��Ͳ~��M�?�U�p�l/D�N��)�B#X��t�o�ύ���7b⋨����ƾ}���-���tI����7�P�k�T3f�PK������P�Ux)V����7���HL��V�a6���=��$�#�E����g%=��J����[.�N$�h�!�5��
��[4�m׿h�Q�C<�8�$�I��y�ꆯPE�Z�J�����_&a"�ۂ������^�mљ�6~n\�۹*D�"���F�E�w�ne���ƂG�|"v\򛕛���6�����9َϾ �K%h@D����K`�é�C�T �jw��Z���������C%]�1h��֭z�y�Ր����+��"��z<��G�8�]
�/�eIN��8�d>��7����R���#W��h�'�pOLւ��?��#�N8��F=�O�ؚ�ymR&�v�7�7F��jP���3�8�ܙ�Ԯ�FHL���� �Ǐ����f��߲�`��j��7u��cV����tg���Q�y(�������8����eu�ٟ�:W'\� ���������EG��>��E��B�����D�ȿ��5@%_�G���5���#J�"K�R!;������=���?� ¼����� ��P�%�$��݋[%=I�EF$q�)+	ë;Զ�74�~��֮�1�f��/~a�I�q:g;jI:�U��)�65��j���b'�}�&A�y�ի-���r�ʬ��oGnڿEo��c��>(��!�q'-]�4��XW��VРADiD�\���k�����3l�C=��:���85�v,�@'���Q��X�2�Ƀ�d%ŋ ��f	���'�'	�h�v��樘J�>�)����:!��+�Գ�������D��fNp��%����&������f-��^F���7�*���`c��:T*�.���'�T��p~^�x�?C�8kˑ�G��xmc�1�OÙ�
)�<��,�w�G���?�wS����#7�qlv>����Z~�X=xQ��)_�8)��y���%���.{s�jN���A����O�|�<�I�ϔX'��٥)K���B�+)�$-@{�7��i�{я��J8$i�#�x��	��#jUnM�@�cs@I�Ul'Fٝ�� �T݃P	� @_�v-;�8`6�J���I�že��Й@��n�틡�K�."���/ɺ������Cy�P󬠌���%TB]v'X{Hz��(�Ʋ7�3�ݍ7���4=�=+0u�Ȝ��EޛM���8&��"�����圼I��C�3�A���������m����^ru���7��2K=b[����>!d1h�OŬ��^GQ�����k�����I�WVGǚ	f�v�N/4�k�g�����ߪ2P�2��B���p��F�\n��)��O�GK�pT�ǁ���}|���2�2�f#��K�X�U!�:C�J��SV���|?N�~	�B+�,�"��E3����m������������z�B��į{�t�^J݁B"���<�!ޟ�'�1Cav~�sF#v���f�Ө�cJJ0�nK���=����.K�0�
�B������,�ǌ��)t��.�y.����q#��s5op3�PW���z)�Kf(��>�Y��U��r�E2����)m@>����JK��q��$ �xF��P����v���s��>8�J�"�td���{��0T��򧃬�-#�֌#�h�#�[̳>�xE1�}��� ��OA��aY��l��y�|����Q��:��_WQ�-�!��h�)0��Ekה��<n�*�޼J���N�m���='D;k ��K���&�6*d� i��}��$��{WY�ݤ�Ͻ����~��.�QI�;'�cX3�X�Ny�Q��85ȯ������0ڛ���4g3/K$#�M`,|���z���̀��;�R�q�����݉�W����S�y�Ȓ�e��!�w�eI�J���{*������d)\i��Wǎid�"�!>lJ���q�e���Pc��S���8J������H]�������T��w�/q�T9�MKB�xc��RU]sZ�E��B;l烏yNP��i$���������Z;��@ <)*0�th���<�Ҙ^t���gy]v�L�#^z���:���6�G�2�lN����Vq��ɦ}~6s���#^�'i>�n �����;����ި����D�Y~��GUp�36�zhѡ��� 'd�pc�d�L4�?�)Wi�:��S�G��s�ϧ�_�8��t���ۊ�i]��Ջ�9����XHD�*j���@��H�y�݌3�P�(݃���6DY9��s�����f<i��m�j �����'@����6�R6���l�?�`!��TG�����|�f�9�Q *_�v	H�=�)����MN��1�S߫����p�#�t��1�k�q���ޏQ/I��T�Q���0���ī!Tv�(�}*�ی����\��I��]͔9��Q~��t��7bu�T�鱤���5b�=U��t&l熌�^P��~��_Xa6U� 7{���Oi�0uy��=�̸\~񢣩���f�ٹ�6���k�����
(!y��ޜ�����?�rd?����h@eA��)`Ͽ�q� W�$4�ۓ�,���"��~|�;뫕wא����-cv	Hft�l@�97❨W�I��a���QfY�Ly�\z�4�s��DiӍ��ݩ��,<�NC��Ċ��f�N��]Y���TyU�n����s)	�k^�%����n��/y��H�cl{��*U�	���ctJD�=r<��C���/b���ס�hkJ��ܳgz�>�?���U_�&�<K^�T����Ŕ���~��j���>ڤ�.כ\ߡʃi|Ֆ=��t5jm����_s�����-��d�u�7t��?7�zp����j���~6r�b�I�q�����~Aͯ�\�D�9�v}W���=��ߏ�~=q$Ů�=,)ߵ��̄2������o�Ҁǹ��l~��A��UA:-�7;�/��w$mv���8G��t3?ɐG�������л����M4��\��4\C4UU�ٿj����|��1ѸU@��"�wW (x7PZ�]�H5�q+������:lۦ�c�
�	��C��/t_ojI��&W�W�՟���th����L���]�5#�lM��Y��p��;\�u�`�#es�F�<�"��ш��h�jZ�����d��I{:��>3���5�|�nnX��Q̖y�X6���\lH�Gqz;^��b�ӳ��k�h/��՜�I,#�=֋�j��^��&���	��T��_�De����H�^��E
�ƾKܫ��і��j��@zU�sd��'�p��(J�B������kY�`����� j��:�e{����7k<�-���ͥ�e�lI���v��Xd�y�牫�u�kSD߄����Mk��^
�Q���g�����bi�IS��\&}?�hJQ$7����ٯ�sΆ�2{���nndI0�&����Wbɉ,i?AوmO.�s�ю�
5�Ò�?-H��_���4�!=�ʨ���.�-���S3��c	���D�d �����Ȥ -��r5���>��c�X;���3E�����k��_T�Hr�¤�Y����Gb�S�?�����Z+Ƽa�ɣL�f��O��s+u�L�pLT�[��[��^�:Xa���U�E�B�^��w^�U_�&*� A<��$$���s'�8�{g��ψ��xVh�x�@� ���|�$W�i��)���zd�ݍv4\�@�����(%�ʢ�~�P�3bK�����UE&��)����� َIh&N�e�::�d���L�2�m�	h#�2CH"��Ą�lb��n �2�CUK<���kLNo��Ys��u o�%�� ���R}�4;xJ�����.� ��z�E�����l5Cz����a���E�R���0c<0�L`!��z���,x�ә�N�d�Q��/�ס�'r�6��72d��z�鑄��F-Nۇ�I4��?����/�Oh�S獅j�7=
�?�q�VΆ�_m��p8�<���?�s��y�^�s���8n�Ç*������P,3u7Td�ay�"B�h<�&�Ey�.1vsҒP���±b��E�D<�xވ�#7��n��+��z:s��:��}ɖ��J?��h�L"��U�׸3G�~�k@�מäGJ��TR�[�n��M��(�ȿ;[^�d�P��MNGs?��q�i�O�k�LY1y�|���TG㞗���o���fRau�o4/�1X2L��,��m��N��m�n&Ok߇�p1$5�:�K���evK�Eʵ�шv���\B�?��/���	n� `��K������	P`�lS��I�}}