��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&Y�%�ddؐ7�V�>sxQ�TLs��*���%;^�NW`�B��Y����5rե�E���V����W��! ���(�ȷ�$�=)�	Z�5��6�P%�ج����0E����vy����,Ÿ4�,5SX<�������)-7�P����؞-��.L2g�X?�S����<��+���l$�ؐ<��T�H�X'�-Pa=�H7Vs���2)w7Q����3T��Ȳ�H�u�)�ޒ�!��ޝɍ��i\�=p<�='as����?�eƽ�� DC4Rwd7ewn��dv�wJ��ZO�jc�^�0םP�A#J�l'�F��|Krd������o�A���I�QGER�ssYT��c���Rܧ�y��LW��N�w�v���$�$��ڦl���_��yTս]\*[&V)��TG0�W�忹b;1�2������T�#	[N��k����$��"U�_��pE�03�S,t�@���v�}����P [�>O�ք�]��&�����I��;��P�]<�^4b�~)��;>�6�M�zzo���!tL���*�à^9��2�� ���<"��0�n����FT�����p�ug�4����r�WY�[%�VVR_�����_Zi�%�=/i�w�Ѵ,��Xnk��Y���8m�>���#�9mlC��35`@���RSJ*���{fk��شZ#er��̌�/+w����$9f�p�s�7-��sF #��I���p�V�p�q�N�0�jX=�i�W\�]0�H��9X3����8��h袰�l��Z����:�i���oP[aL���i�l��M��QKR�jm-,��=��͈���
6��Luҁ�E��73_���L�)���&=Δ��8"�>0y�@�0���:m�[��QT������Q�e^Z*Hmk��^����j��`�1��a�w���^��8�̢0�m+a���|�2�e����ß@�l�Z*+�jڊ�T#��D C6�vv�:�riK
J&}u=�*�q҈��|�>�8(
:���I_^}� ~Q�/�G:��f�y� nl� oC,�W�@�J9L��U���~&�*4Dӱ�K���LS�]�ˊ��� ��b�b:"��5Q���_�E���Dx���� � ���'��r��f"/�������i�B8�^�_|�]ӎ�>U�ѣ����P>̹����N���^Ex�@�Q�L&�	v}��^��J��aV�I����<��!n��?wI/�y%,g�ȊI���?��Rv�"�hJJ\�듂��ڋ��&��#��6���L"2x�$�J�9}�Z<m��-�G�z�x�Z�
��ԏD��#R����7g�l_�֠T�_i���1;_�%6Wq
�����h����N`b�T�[�n�$M�2g�_�S'/�-s�S�dy��SٹKI�Ϙ�/GYoM�U�R�1���rp��m}S�&���m�&����4� D`�+ [�u6w��6ě�y�f�eȊߚ ���lS?O�1ִ�iM_�����z�|c=/�Y�`B @(SSv9�aN�'p�-ﻫ���܇��@`���'_����`�2�DI�_��eC͝�ia��u��v(��a�����O��HP�����q�V��i܆�Y0v��Y����,��'�d�8[B+73M:J<���[M��;���ȃ�	^y�D���k�åZ��%�#=4醹�B��a����Ռ�|������IBHB|�,�+_�~�w����D��+
��|Sh�;��u�lR�qN�<����*MR0O�M0��|����5�A|�@�}���h9�������o�YO��_T�����̒U S`�4�q�@$��Ew:<����o�v韕�=;:�[U���1=bhRh�:�KC7?�;#��,^8`����.B�&+c�im��$�r��$h�C����nh�J�&��=���˾~*�Z�f�����s�S�0��Y�
�����}��
��ig�� 1���	2���w�Ɔ�X��:/�ÉJ)�/k���~�KM��VA�UU#
�8�^&?�C��m�e6`9)�t�k�U��%cnR�4u;�@n\2H)u[��9�k������.VM�u�H�ۖ3R��	�s�j	 7~��x�u���P>c��fRcz�#8h�/��0�( ���B�� �\um���<�R����H6�K��g �,7�bs^s+P\e�4���C4�0�X��m�-0TÈ]ySU��t�Ik�OX��W�\�wz;�������y{w>��[���gF���.9Rj����k�{R?���h�$_:�G ��wt��r<_B&�<��� �@[#;l�+?%s�J].c�e�\芣F��
{lX���$	I0ߠ�8v�GF+�`���4?nפ�<STSB��s����U�M	�/+�)�
CN�%$]�.H�h�Pr�����l:��Z��m�J�M�i�~C��U�4dY���r����W	ڙ]ix1�$9��3g���T9�`ŨJ\�-n��xZ��h�?��F�K��̗ʷ<x�@��;TI�#}�����������G�e<t3�_�i�	~�B�M�!�&���R;����"��yLA��ŗ�����ی�찖�l: В)�"<9o��� �O��~X���Pڴ�%��d�#��f�S��!�ig��G��Ќ&�~�2�/�#P����g%��ҙ���KR2v��c����-l#~ỊD)g��_yz
����3����ڷ����\�`GX����v�3ȣ�2;�4����KJ��Va-�_�ɬcL��6l�T�pg���/�[i�q��7Yj�`Y	� ��	z�@�sa�d��%��yk�j��+��|l̲�E��d#�{���u���u�0t�˃��"RVm�i��a��ᙢ�G6��{0K[�2V>Lg\�t��p-�ЖYځ���� �ԗ����it���ܯCnNmtBT�:�"�7�]�.t�7�Q��sr)ʲ"�B���tO�����4��n�t籱���gz�1�t���5�!LYV������E3�8��AJO�Gj�l�2sq�B�7�x��T�{c��ʨ����Y�*���Yq��H[M]�����KY�0��=Ie0&�ѐ���DA	��..É��a���!��	uQ�����D�eSWn�xZR�D�+l>k�	��2�T
n-�|��J�a�x�^&j���fd�4�?f� 2�A�s��M�&���h�w<ZC�f�L�gB�I��õ���E���p^��Fh�$=ڰ�t �zB���{|�$��~��v��6J���r��t�9�u'�A!��*����jw����	�k�~S�+�I ��g��C��-��c��9ggݞ��تW�(Q����hx"����l%P�3�<H��~����.��^-���WAFnA����Qj*89�$�9(F�Tݟ<ԡA�\��*A��ĸ�b$���l���!����'�Lk;�Б�E��}�<��b-�>����R&�^����6TvQZ��ho�$~ap�W!� '�N�y+t�f��&����Y,�8�E���U���gu
�����r�Di�2�m׳NB8U�f���C�a��l�bd'Uӛ�$��?I�M�7�n��:��|�4��.��d\�A��l�|��̀ܯ�^��&��՗�H9�G_�Rh8ߓ"leKץF�J�;=�P�@��bLa0�P�E�s�/�w��O(��QK:�[w�]
��]|���ʞ/�/uܸ/�����哸����y��R-�d�܍
��G��dի���*�0р���-Ⰴ��_z�y��SS�~Z��^�N8	��2�&��J�a�4`���ʫ!6y&H9�Z�n��[(p
�V �^y�����W�]|�5�pN܏��ҥ�=�﮼R�A9Vl�S��#���U.F���7糞[՛ y�%�0/nTY\XN��׍
ިч@��xgu+B�Ox	����"{t��Pu,�p���8퀍�`�$KJ��zLe�:��i�<Idasy�����p�9B��i>�P��Iė��e\��A?k�+y��2�n��IX���g0c�?�*�e��ԣg��d�����◔�I�v������1�2C��;Fd�n����Y��I��"��J�Rw�&�jA6yv��vv#������Ŭ��+O��n����]S�-ݦ'�z�y'��*��:�kV�V��yQ��(�*�Qʉ��h2�S��/�I�z�,W��.%��is�߭�lA��(��Œ���~�x�p���ϕP|Shک��9�bk΄�)���i���l��*_���eG��K(���-�����l���.���Z�H���U¡27�q�Y���P/T�1g�
8ݦm��^JR?�Lџ��y�_S��lVI,�i`m*��F̠��8�7�� ��u�o��`zf��t
�?3<���N�#N��:յ,�v�6���WR|I�1T�C��z���qQ��퉂�x��n�QLo�Z ��&̐62X*̭Ѡ ���n5s�g����U�P]�~�$]�>��6]L��y'"PDi�*��_�c��7S�@�P�t't���Ea'S��a���㭿�xc��u<a3���s2�0䌐��-�p� D���(I��l�@��{]�Lx�ޚ�+~�?�l�#]�hН�Zt���9�g��f0�ތW�i���4�=�i���c���W֜O�%����MQ<L�]X�̓�(��$��B�XR�ϩ��u�ً.2�hgy脸욊� �=�w���~i#h� d�ɱ��ϴd�˫�L�*( eU+�i���)�5̇�����%جq���P���3���6�='o�Z��JS���D�v��
��4Y�	:x�����65ǲA���,Ź c"�U�y�dPi1�csT���V�C���"�����5��64K�1��/u�Kڇ�-\b�����}�=�k�(L[��@�bD@��yF#���a�G����j)��>U�x��K�H��BN��-�Ml��WErp[�?لm+�u��{�&tי�mͻ�v�kU��w}u�b�ݛ�M���{�+�����*��]��i\MG���C����[FS1�N{v�p�v]�� rr�_���y��(M� Cy'z�Et��A�&3��~ӧ�\M�;�`����`�X/+�����R���A�7~�۫?ʨSj~��yL�{F�&���r��G�|
~$u;1Q���3D���$I�@�%���Wm~/��ػ[��Q����#���j��y���[,T &|G/E�qw��`�X�����0}3���=$��nȢ�����.SbƢb�w���>'H��\g��-�dV�r7��{Nyw���8�']X�oa�|˼�z���rڒ0lU3��y�*�e���q���+���oSF��S���C�ʨ���Y���'o�p��2BR�!y��w��W�*���-?>D on�v�^�~0Z�1�^�/L�2�s�VgfR�x/�t�W����s0/C�.<u��f�-�k�W2(���k&�I�
�\g%=-�:�$�P/����i�*8E>mص����R�#����PV�{�] �@����eh��Fd��C"����w�2Q/0���*QJ|�y �8��;���R8��}�����`�9�I��Z��v�»�+h�to�Ss8��F�v��Ǔ����L/X�-�!�3J��������!��S�o���������A}\T�VS^�uW�v(���o�D�����T�F�1�z�����%}!�yn�$�	�)�P5�`"��{Ǳ#�?��77�m�&{w^ۀh��5��w��7��6���U��Ò+C�b~ �P=̦�K���x�k5���Hm��Tý0�5�g`}N�D�E?mZz12�-�<��7���Ȉ-[�sxM���jH�$4��@{E8~�I��Jk����F��	c�s��y*�`����pш���0���Oǅ�]@�GZNxod\�Δ�2��ƹ3+H�ɉv�_0&p�)�^Џ����{юÉ���c��j�+ER[fl�V�kBOd5���#�ȏ}�ʬ"��9OaC�5_��͉��_�cz2�Ƣ�)|��0��#[?�^�t�
��ɺɇ��E��51�\�O��|M	{�sfg��R�7/=�>u��~�ZC�e����q<�����VA"��%�3K�f�2�\�{D�Ѧ�{9ޞ�V�}ܚ�f�����fGѲH�p>�?#������>���	Q/��H`?�&j5������#��.�v�L�>�w����"�l	���]"���A��'�[���.6�~8���9���z�((��љ����.Q:x�A�9�x��s�ZH����Th�����幢�FN�,Y@��Ʒ2��D�ݸO�Ő��G̹�k����&�nӰ�6�Nj )���瓗`H�~�b����#�J4�uF�_3a��M��;�<��ሬ�%��V"�,��U�l~>�m��x���.��J����h�$�����s�#�E�Plq�2{��z���HU���C]����R�S!M���byꭜc�:�� �����~�s����K8�p�����	���ḃ�)?dG5׹	�$�Oa">3{�^%ǍY�C't��^�ppI̡�U}�����@"H؀Ug��66F���{������D���&Q�F��Ѷ[�!MAc.)����K$��gp�^R9�:�z��4���~6�k�M7/�4��Y�e�B�ۆ�&������X�ϰ�������R��_M�g��&f��g
���T�s��;��q��;Hir,q� ���'?�I8ŅS���o0�|�/q�����6����=,�<��5�n���(��(Gh�����qX�5$z�z��F��6[���lp-(�O)Ʉ�	��:ۗo��DL���׭</,3eETl+C��Ute��y��k��\��!�l)��	�5,e�>Z�!��m״�,��3��E��iY��$쌾�P��m�à��k�����f�y�q]�2Yx&5�K�B�wC��$�1�p�έE�zb��:.D�3-RjT�H,�����G�i��K����c��K�a8�C0���N[6f�78��=����I~��zU�v��I:�j>|d_����D��j��jPC�N�-a�sH����m�H4ә8�6�n�:��B�sPy	��X���]���RR�[h�~��6[��t�yJ��c��z��]B��C���r�/R0��3ĥK���:6�B����c�$G>xgم��Ii�d�J'�͢�t��������ʪ�HCx��|�і
)�zXP؍����[���%A��cu���y��n�&�F�1s8a�G��"ۯg�\�����r�C��^&HW��lӊݖm����:FM���j�$����Iz2��@�jۗ��=�*3�H8M��w�=�6]�E�s���G�ذ$�$����M�樇���A�����W�}�xB��<�i�k}�T���X�P�F�i^m��x��Oo��7h�����^2�)�����-�72�� CG���ίǤC���Ɂ�ԂI�w�l�
�s�	, �	�Xc����g���Z���`y��Rs�������z�ݱ��hd��ݸ� ̇�ܾ�薯\��;f����Al�FT~U��^��t�s�ymV�tg� �m߸Mɐ�a%��0@�����0.X0}��0�&zWu���Ff�۶HԘ*�x3����U�9�+�}yX�v�*�7���W��ڪ����^(�s���߃��ΐ�h�)� ~����|��U��_��J�9$�������[�ɀ|�DO5_�}^���H�+�9�ү@�,�`�;1�%��Y�G80��#��I�IAĻ�Uxr���O�C�3�at�����:@c۝���tz!_rv�m>��#EX��T����9�W�бem��	�n���ܩ�8F�d���>�f��F��Y���I�V�7i�2�FU�����eL����]�������?�i%f���BB�������+v�=���%��a��c}`�>��?)��1ʹ���T��Ϋ}�����(�d��O�T�ra@�;=v�b=�TͲ�iz�L��?���p��������Q@����2Nl-�e
5��DUؓ� \v�'����T���?�>)2_g_���� ����㧇������$����ocJ�����=�nU��npv��Lm���$����:��_b�[C�Y�ٰOF�Rq^��*�m�@��f���:ai�x
!X�F��f��pOц4�`��96���(j�fs�IN������3�	�A0*�%F����m����L��X<�Xo�+�י[F%$����f ���K07�V���lZ(���Q/���ʽ[�7�S�lY���~��Ii��ӝɊ����qlιϡ�O?�'�>�Y�I�Ls҅R�q�G,*ﮡ�"�d}���^Á�'�@�F��G�QSC=�Z@���́��7�mV�,�:���zD|(I�N�:�h��Q$�1�P[�p��MET��8��C W�DT�E\v:�8>R� ���r�G�;pgE����\�Ot�O@�e�&)���L/�7W�_>
s/�պ�ی�v�e�E��ĳKpc7�!� 3�5��Z��I�0+�?Bn�5����&�u	M�<D��[�f�H�z����&�,�Q�
��a[O�y;A��Sܓ��@'/t�o)M9v�r�%����LUǪ�so�|c�;���`"�Ol��Z��=̀Q���]6p�Σ���E9'/� ���$�!�fF��L�	�TNs��l��=�����GU�s���94`R��!k��������D�U�8mz@��.�.�R�D��^0�B(�r�u��#��y�d�6F�@�m�d�������f�8P�=�������	W�1�S#��ـ�D��*	;R�C���R{VN��wD"��#�m����(\-����U;W	���ٌ��o�{N��7k���� �eD��[<�Xj8 $�x�#�B~4�,�|���M	��%vp��'���i2}ܳ��������m3y��,�����E �3i�-��caWU/4L6Qy+�X�g $?0�i�r��=�%�X�S6�b������8�=�i��Y�g�:T��� H2�2D�6n"D[�N=���ק}r'�y�'p���]��|r3<Rs�@C��	��آ|��.Q^�7��Ɩ��ov@k3a�$��AW�=޴I#Y����G��������(��'�o��;� ׂ҃�=,t>&����pS�W��;VrRc;f�[���1:Ű�lr�61��d��Xx�e�c,>r$�V�ʒ��z��? ��J`9��l�{h&�[�-t��4�x="�#�Y<���Ǥ�@�yp:�g�����|0	B���z�k�d[7>r[ș�ͨ��=r�"��͊�,-�;wU��8�Yȷ�+�a>��G���V|��0R\ey��:MO'���2R`"k(a�Y*#�~AxLj*67�2p�|v���62t&��)�H�_�X�Qm���~�jwu� ���Z_��� <;�M�����AU�j&a~�+�����#�`��u/b�6�O�XN��rv���n��0��٫�Ě '�|�ܺ����w葷�*!+���vb�ZCm1Q�B�tv�گ[!� q^e&K��Á��B���E�|���-��Xj�Hߔ]r,�e���`��δu��\@_���靮���E`�"N��^a|ye\��x�M8 �V�s�Vr�Tai����+����L()���j������:(�����v�	̫����p�����q��X�ɲ̯�h֙����D��ko�Me���cF��K��%꾀�ݿ��4��W�֌W�f����dT�t�4F���7c���~����{'��qtq.M�n7�++��X��䊊d�hė���hr�o�����n;{	��~�E�
�������z�T-.�~�_k�7���r.��~I����6���M�6�ԁ��ի�C��y�,��X̯���.�-U�����9=Q��bZ��E�5C7
6���ES/��K����~�ai�1����m`�E|<���B��a�a{_�R�
+W0�ki�!W���~����u(��S�|�W��2����r�\�Ȍ-]�y������U �j������&d*��:1��6�B%[�F�4͑)d��'�1#H1�������?۝!�e)DB^��q��<vD������^|���|��DX�d����@3�T�P�掴M�,����W]�\�A������AJ�e]K�i�dOx�Dlm�Eo>7��?�GwS(7a7���.�N.įES��
�БW2ґh^ړ�uD0�8ܡQ�Vҟ\��o$q�v+څ]ZS�ˎ�Q��іbfky��?��@F~W� �Q��ޥJRM�2=w�$'00~�����_S���H��ھ�T���X<T��:Xe��e�(E⻭�Y�E@�3��f�Wli�H�i�����k�n��$����N�2F��i����P�n�ύ�%��!�l͙t*�nm���i�	���#|��a` �����+�R�nZ4�x��#�$��k��0XG���
Z���<��5���������E����_��ɥ����^���c7V^O��Kor��.@�2��A.��L��i)둊}��X薌�` ���]<��w�g�I8uM8I�tq�Mr9O:a�b��m&��{q���a
��z\J&���*p�4bF�
!;��4{H���|������R*�_�敻b0�+��"1�v$���^|	���dк��e�&�����d����cȨ���#�uqjD'�~DFϡ�mz=0�w�l�+ap*���� �/	E�?N=k�,�=�=fj��)<�W�����Ű�sp�Qo�Y[	�>��"Y/�_�1d3h���[��7�q{��y/hp�2�p`g/J2��٬< �.�|d`"(���puH!�޺�j�̌�f܆����c=r���贈��%�.�SK� i��
�P8?�M��ao@��{�o����%
������Fa֥�5IeɈ��;�t��=�V1V��/�9��R$�E N�P��"�w��� ?��ŻiE���'�D$r��!E���ˍ��Cً|��	]����ZsQᇐx�W���g�ͶJ��P&�+��c8ȋ�N�<X�pS��26��w���P9��:*�d%�l/^����p�	L� R2m�u��[xTe@��7f�ԕZ�Gi��;�ђ9cf�c�Uc�*�\=y��
��WXB߄S���*Ȣ��niJ��l�#,�G�+���*+r¤�Ջ�iFܼ�d��n���[����:���zl*dj��؅��d��yE��n�ʓf0��� �}}��WD�Jg�<Г ��wlBk�q'����$A�g�E�+��"|Ȱ�?G�*�F]¥ʬ�k��_�-f��ۍ_�N{A*Q3���k� },e	�+p@�0Kv�%뙴s*��n�G�"m�S��	�Eꁸ��*K�ǮC/����[��I�Itk^����v-���l.GǢ����ZW�|xa�l5�{G�%��k>����mL��񥪱�mzp�B�.�D��}�(�Q{�v�<�bn(Ș�v:�g��H���v4U�������Y��$��
dh�<�}�n~V��&��/A���8�B�Y����v�f�f���d8M�������UҮ��w�p���r�>�Q�ΰ�],:島BD����hبƧ�2��5�N׬b�?|2}������	����hxX����@����������7�ag|.f��r
Zy�#K�˱zv���톇馤�A+йm0LȢ+p#�����ys�����X��j3���ڑSk��F�oϘy�,��PS�S
NP�|>{bس��9$�|�p��*���Q|s��2պ����hd��|rK_E8����{&��������]/&�[�0t��I�������6i����2^3HjȨڱ���7�G<y���ؒ�-���4�2��d~�̳��h�{�&��,yq��{Eh�X���k,��*������l���=[�AL�4��&��{�[��?X��k�J*�U�����UE��,�"iJ;�(����	��okS�S�Pk��n�PI�(x�4��ǔ!�2����!���$=0Y�dJ�;w�Hkv&Oy�	ԣ��� ��aB�����7�KQX��ږ�Ϊ�D�9g���1��~kn4��伙���A8�!͟@�T��j�f���mZ�@c��#Y��O�`1��`�<����[5�"�������h"{ڜ{�탱X1ߝUe/(Ǚ*���0[��ӃJ@�6׵B?K���C^��*��i�_�Tc:��@Z�B���#��Cm!�R˽o�HK�GQkF�3�i���5��XZ����5��R�a����]x�Yr�P��<aɼʫ$��£� £o������y�:�Ԏ	,��@\��:�m�?ֈ'��J�k���%X����\<`X���m.�U�tθr8 ����i�%Α�D��F�~�[��z��$�I$5H��_�C��N�ΐ3;���<�L,2���`%���K"���:��:eNy<2' �j���w�W�XX�~�`f�C�D���rT��;��#9M�M�	6��:�̩�Dz�|D��w)��Af~�L��L[t�u��U��C���G���+G��T�0��lʆz)������9�����ak/>'|��67L��$��c*t�9�~���D�{M��)��s�|���Ru�-J���
,�t���VPD���T��c�wA9̩�8��.T.Iy�J]7�Y���2,R]H��/��=z`Z��b��� ��������/�8��`�˧V�{п�Xt�*aG��u%"��~��}q��QK��Js������g]@�c���[���x�2�	����^֏�i��nK�K@�j���1+��֧~��F�[� c>���8Evh�����v;�#�U�M��^�l��� �u5ho5x��n{<p󟈌0q���:7S�t�J�C�.$�0&�l�^��hJVk V��+����]%<�@x����ѧ jЀT������A���iB�{���/z�#�hd��}|3ٸ^Y��\�� [ӣ8�Y<�:%� kM�e|��Ե�?�K��si/M��ъ�nT����9�b�@lqX�g>�qB�cys2����<r�Gu�e�G�W�)A��C��N7�v=9$cS�&%����ǠB���K��������C�B�/o���/c��65�;܅F�2_�@�Va�P�6�k�r��>��'�<>��o���~�u��ٕ�I5����"5�}.�5"�-��(�c|������vA�3L�t�Ł�Y�ځ�i�1{G�l��A]�*#�ګϱ�a�E��LCFW����,�����'�,S�x���<���5��>[v�����ª�^�|��7�酞8����ok��4��4��g�p?��:�q�y����D�?����s
��0��u��C)p4)��v�r���Ɛ��0�IH4	���R�cT�:q�F�U��tScG��-W�,���)m-jT�dd�����G��@�L��%^�� +����@���sN�(��W�举�M���!�p�y2v���q��ٔ'Ջ��xB��z 5�,W8?���3J䘩��7�):��@ �\�������(�ʫ�����$;��>��қrᏁ=��,W-㐂���#"᲋i �P��}�/J���C.!%m�Xx�[��R#n�Ǥ�1L�[b0H��6!��Յd�Ow��_!���Oa�
�kL������@u�Z@e��/Odq��C�$Q�&��~#��*	�$�M{ ��1���/��yP�3���{��� n&��V��?n�[<SŲJX
�ً.��X���YΜ���0����גx9?���F�ϼ�1��z��C3ob��*�_��^҉%4 �����Ft�8�)֨����a��2�RJ
���`��N�F�	"��M=���A����f�肌XQ̤W���!��%^gB��PF�c����d@2P�S���3j&��eO���/o&p`�F!�`����4���t�f���ۓ.���B�28�3�4�Q}��3�%�_?oY����UӸ*��KA�c��]P�p�p(ng�Ͳ��>�?�Q�	�E�H���N�?����VS;��mp������h�$R��+��vf���uE����Z@����~(<�vB�R�-^����Q9̮{)R�B-��U�K+�=q� nl-�눆�72n�A�(�*�BS���A/iX�`��Y �q�{�������g-�Lm��=�J-	[\��