��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]ǂ��O��˰�	JL\=����"pI�: `�r��+i���B�Cp���,��1��o��(V�M�`SqkH㵊Kp9�=�B�(�ǋ�ƈJ-Ч\~�:ч�	�5��O����RwK��zHI�2�Io8��5}�+�㛳����7�K��Db�s�}䢓"�nOܧ�����0d�3'	�`I�7Ђ����h�4��C���:�(�ۓI��&�݋[wf��.ţ�Mw졶��׾��ʻ��/�TM��Է"�Fcf ����hw�O.~&uP>�h0�SӨPFٖ{��!1�Z'Y����C�qy�UX埭����1�ryW���,�����͟��!#�Cv�TuBjg�1��WZ� ���Դ_�;_[����&V��$��~`��� �����C�e��6��c�nA�8ɗ;ɄC/D�(�g�oM�i����w^z�'��2��C��p