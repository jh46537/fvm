��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQl�E��*����XR���J̕�����-Z*�Q�o��`�����^�\�?��b�L [���2m�ei����
`S�����/k�#$����n�XT�t�����W<}P�p���� ٽT�m��|���i�<-(��U+�n���DD�B��M$(�<FUH5"7��i�H��Ӥa�O����۷Mæϟ��f �?�s������^-/���Pf�$������q��:��b�$v���z�BVL3���#�L�D�ڈ�T�Y�![�Q�М�.�8A垒Νt%���k��,��c���H�X=̴S����b�x�mE��+�w߉x돫���>k�8�E�ژ�̸��h�a���C�_�sz��p&;������>��O�l?�¥I[q��'��ŝ_��	f��j����@�e T�$U��t��YZI���`�P��z3�Ƕ�k�)(鄟(E��8���;р�w�r�UÃ��G<����V���6܀��J6k
�0�y�>��-��{����k	w���]/֋85���&8���y�۾�✗���:ːX8(�MO�����ӥ��i���	�"�ai��LQG�7�QXWM3���QG@u%+_���������`�� {~�%�d5Ҕ�u�F�z��X&?l�X&#=8Da&B�+�ܯ���o�"A��q�j ����At^���B��Н�vi�����z�[�"���CR^�V$��y;�l鷂fS�fZ!�y��1��7��Q�OzA0�ʮw�0�T���0\^=[K��$�HT�O����!���e����6�T��ʚ`�8������r��$7d(Y���K�R���B0��F�4�5���:-KSE9�ðt]�D��Y'��qB�b�����e�@��/ގ��36�m�{J��@fV�9�j�>>sm�%=Hw_���+]�T��-�7���jf�q:_C���*�b���l�% ��%��$$MP+�to8���ʟ���gJu���	�g09��ao9̴x�/��v���Lh���9,O(�
�x�M�a�a��$v�U�G�$���Ɂ�ß��s:%'D�I��ǡb&��^��]p�Ή٥͹�?H,�Wկ�h�k�}�]�{��ȀF����y������ekV�S���mϼ��&�B�o�ن\�j���D0y��X�F��r�IJ9֋�r�i���_��dK��Ԇ���@tޭ���ӄ�*�S�筚�D�XC|����"��4���Сk������������J��s�3i��ڍs�E#�^�~�&�1O=R��@��7/'�U�O�C��e�QE1��TkO���+~%:.���PD�_�Ζ�_[)Dnsh�1�����O$���A��A��`D z ګe�H����$��LO@��k�H> Z��<ED�h�ӣѥGf�y��K%�z�O9a���$0~�m�e�㶣��>�����Q]��f# ���|�U;k]m�������/p)ߛ���q�6I��Vj�i��u�\���s�.v`Lh�ji�\�y*%�G>'��r�"=�I�2|�3�h��y��w��m�^.��de�gi�Bj��o���/��uؼ�:�k�wE\7�������
���9��Z������H.~Q��^���s�wW\�V�2� �K��I��X]���yݢ��zI�����y�bfL�Wa����w��,/'
�_\.>X����������c�T�� ���]��"YƨƭG2\������	�)mm�9�����A����	t�N/w���s�8PK�>d��vE�u�fI�!d��쁸s��_|�:��k�/4�ga15���ރ��*�w�X��`���c��C*⳿RD��!Y+F�B��Y�3}k�Y��A]��Iܳ��HV���Z����j'BqcK8eB��Q	/f�+�u^��4���ȫ3o��悘�/��
��>R�9z��m�0ƣ8��@��l[��|S�X�,����_E��]�����^�~���U�:)v7��	�G���*�cS��%����c1���rQ*D��gωq������,�ڷ6��m�P>��E}����N� A|`��=Y���A5=o��|�?�	�P�=��@��ȅa�}"^���X��)O����*��F!��m���}dj\���3��9b���w?SM�ڌ?'ED��f	K��0�qk�:@nN`-@�S&1j��G�?���hޓ8F��afTrk��dI������=W�b3��6�:.`Ԙ�{��!A+js�
���&�׭�)E8��
O�"4��q���Х�3+h�j	���l��#�~�+f����\T�ʍ����_(����ˮ�y�n��L�ɗ��r��U���[���&z;��I��-���w%��C
1y�d._���<_sc ���/��`����lRes��>wa00Eu�hvzq��Ż��JO��XR���,]l);�~"Ⱥ�V���w=�q��b>�t��Lc�rj]Ј���q�k�W���I��r���e�v�2f� t`��3�4�horƥ�+�t����C��	�p1�NFܤ�R
��X����b���{��ca�UG4���g�G����n�ORW�����ȳ������Tq��*W���9Ey�O��U�X���S��z�����>�d}m�Z�m<������7�z@�6�[O�K!^��>��������%�ԻB�)�ZKC塶�<=u�!Y��z�s?K���膇bK�O�י��{V�����}�ҽ��J��f��]�p��i7�C����w��J��a�V���6׊댦��2˃��J*���I��Jq����B���K�Xm$y����{z��|n4é�<��v��i#X\W�Ǌ`sV"���49bpo)�1�zZY���@8��l��dL��N�8$��{�P����x��׺MU����K���/
s�d���,��u��
�I跦i��do�.oľ���%��)ڡ$����M/��l��z�z< J��i>uk���)L���h؝�
5��Ob��=C:�:e߻�ˀ���&���S7�}A��f	[�X����z+��J�f�.u6l\�j��&����щ�����&�OEu�� U�ti��=f�<��y��T�*l6W��1�E@cua1T w�ٴT��1M[8L�"��n�B�����*.$ya"
�
����4���9"i-�����yS�n��|ө���$ \�k��C�����k�����ea�*��$AR�ID�^��7�"�0s6;%h*��b�9�G֕��"Z��ZO�'ݍ��]l�dfK:9�xT����<s�q������ذ*�Ξ�=�u�u[_�R�k�`Ժ)���:8���t��׹��i[�"3,��v�L!���#}�����2��o)���龊�_=��|��;�'޷B+��2~��Iy�I�5�z���;�ڻP��Z������Ëi*��
9���EH�X�5X���?΃�7μ&᛹���p�P��^��k'�Q�=t�=T\��G*1�wQ3�0��rZ���Jl���?%-:�.��ƶg�"����1҂�S٦V��(T<�5�;Ғ�9�2�����S5�#L��i@�G�n<4�9�jv�����z�!c������������AwV�Y�S�͐Ù������V�c&�8�\I�;�48$>��!�T�SC��g�Ƿ���x��'����C�Y��6|@!��"�VrF���ZR(��I��Q8��o�1tL����$������zlew�HC`�ĝg"�y�l��Fm�PXg�^)�f���L�֋�<8h��19��t
K,�<�I�2q�1e����-���r�?J�Jg�ap�j�p]��Q!��^�f_N!(���;v���K{���F�|]\�vS��{�~�bُ����Qi�����T��A#���ht}�� ����ދ��]b�)��qz@�H"d_^�e�.
������4���P-:��_]2�����zz\�D�u7ќ��L�-��\�Dc�Ҫ�"��n��&���Ф9��x�n�B��\����ʘ3%l�dl9V'{����9����Pu�G�c)+}�ڀMxm]�%��U­��Մ��>=��:�i�&�.kz�F s��a���;'X�>����:�3B�,Vs(��o�.�Y��4mc�o������1�� j�sw�1|�:Bq�t���H�C�����'^�(��h�����b� ��Xgq���@%·���C�jB��St3V��<�������_o[�wcY�'Dk�.U�~;(��.*�
4:m��	{�wH��lv��?�=��	إm�^��Vm*sƁG�k4L��|�ol�n�@H�[|'E�>�J�ѣU�+O3�3�We *����#]�/�z�������=%�֥���0�!Ȳ�Ш8�,���!C���ߵ }�Phb������4=s�+�c@���+z���w/��-�iXa��>n���s�){�i���|����5g��7\O��0�69�70�n8��~��\���)=�b���Oq����Ć�u��� � a@VUPWoW[:Y��k�ߢeP<���D�h/<�e��RS��� ��C+����-LL����>6���|i��E����M��Ǣ�q ��)�-�<����bȇ�y��5zg��`���"���FX>ݫ�u�C�?���<78v3��H���v<�����#u]., ؎��KSto=��R*�J��v��x�.j9��-�b����z�.�c���+|00�x�oeڈ�֖r�Ȼ1^
 D0�6Fy@�~h��:G���u�32vm��v7k�晟�pY��=�Z���Lf����|N{��]��E�J��utR�c���C>o`���3*��$ 2�OȻ�_A������:�1���k���g��=6y@o^5B�6�r�ق�͕���q ��1��i�ው�:���XJh��� B rV���Z>�~���c�>��.�F����ק�����1����z�
â�
��z�7
΁��
�����&��L*n��l[�'Ħ�`�p��RQ�Q���傥����g<s�N������9k��[��eρ�e���}w��F�Lw�/��C3�r�n�.?�%��.�S!���=Ј���R�͠g2T[�rK�)�tT��ݛ�� �Ō�ϼ1�B����LJ�4�~�r<a?����iqHp$��V~|51A��&^����z(Mc�� �R*�:U_��.�SET��N����qt,E3䶊�y���u�!;�:5�zָ�֩��d��ۈݷX1d�53�27|��!x������w����<� ��PS\���F��g����y��8I���`��>X�c~�p���>_#���hPQ�F��7��M49���s�-���g��P�k#�*�sA