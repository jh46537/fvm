��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK�cĜ��O�������_#׫s+St<r��~_Yu��x�vڴO�ruH�(�YF�gq�v`
�l�IcG� �&�m�qqKG߭}S��nO!Ќ�㢤�?�ѿ��^rs��)��X���`B�<a�����-H��=/u�j�xxO��Z��3�[���),����5�3�Ʃ������}�r�er!�:�ә,jus���M�^�9�=Bґg�q����/Ws�Y&y �1g?��"���S���Bws�|�к+O(��H��}[�U��_ё�~[���YXC���uyI�E�@)'h]���`?%j`���D�l���_<�����v���s����� ]���ۦ�K��>�m�3#�k	 �X��£�Z��h�w�s��'�}�g�9��X&��Hp-μ��P���^���
%z #p��s�;�!�h%u'�R��-�X��iOΧU�U�\!YM����-�5��2"��B����G7����jݦ�x�b�U���y5d�;n����&D�a�T��d�f�<z߇q~t��ֻ�?ж�
�Oho
�س�E�����:����J^� ¾7�����=&���e��#QG�T�2O��)���0�s��Î�i�pz��d �[�c��G�;��
��M����3��7Vs���.���Ⱦ,��{�TM��ы���Z�c@w��D!: m�d�a{=�LA9���u~�*
ơ��te_�l0��+Km뜪����j���TabM��E6�J��9����]�9��665���n�C��o=�E��+s̀H �,�%]�4�H	��Ă�E]h-��~�\};�Dd8������8�����%aI8:��'N��]Y��ְ�����E#c������4��xe�������ݙx��]��D�b]�I��7�ȝO��B����g&��.O!B`�L��:��>VJ�X��c�щ<Ŕ4[�f��5xu���V���j�8ʤC�����hF)� >��Pe$��V8!�H���E�8KBz��o�jС�QN�)a�Qҧ�s��9�q�ԕ^ΏJ����>:�1�Q��t���a�7<W�K1{V?�~�����-�=�QB]I�K�+utâ��8$���$��$��kn�t��H/2-�A�0���ZE~��\҄�M��`H�ͳ
�<�|�JY<6{��Ct�?�#�T����p+i��~�`���G@�p���M�땼�lM��Dr���g�ճ�&��7+f�7y����B�Y�Ҽǃ�Yܗo�,���Ϟ�����8wt�O���lu���G��7�千<C���d�D�U�H�S��8���yB�7�n��qW9eܨȩH��y�6��>}hO�<��F|�gR���`��/��������|z�K:�#&�&F����Ar��QlZ9�tTnLӃD�b/�a�A�[�M��x�L==VI�5�i�Aw�_����H(�+0cMs��m����Sh��Uf�E,��$ĥ(ڍ��M���S��)j��B�PVSԅ���3�+p��M���� HxOhX���p}du�`���ˬJ�N���J���-P��M��j5����{�x�I}���	�<�vI�3ʠ{@� �����\�S��3	�	d��m��N���|��	U�a�W��Wn�]�J2FWM`�Y&hTn�Z<A$yB�?J��Ҿ�-������_m�2O>/�t��x����q�^��=����"C ͡�4�c��9l5N�{��܈��3>�xD��v<��ٲBk�Jtu>�{7�f�5��7��7��̟�t�՗�����&��e�/���z�ʆ"y��(3�tt�+���;��5�p�d��F=�����^��a�8�q=�%�$�j���z�&���hB�����sa(XO���͆Y�L���!�����"�I�.��,�@�	�zaiؓ�qx�z�ƍƖ�8K�^��6x]H��P��]F�j�	$��6P�I���n]����(�gP�њ����z�:����B5�gM�&|i��-��V�L`�#������)�R����SAP�
�� d�f���ǵ{A��:���
�&�r����Rݺ�&U2%��B�I�͘"�;�El���)���h�N?����/��8G|(�dm��<�|1�%�n�1��F��j����,0gGe�K�;2 ٘�
��S��R���Da��X�wnut�&Z�Fu
~x�<F(`����k�\G~�̚#p�|��\@��ٮ9�z�a*��N�� �v�$��%C����cVCd9����#�Z�,q�q㋿"'}?~���z�X��E����r�~SZS���KȻ�H%wy��H�ҳ�t-�����䥕�R���4��	�$�h|6���[��&�1v�+��KI��������+Dkz%�H~SN'�F(�|E���ߜ������؟
2˅wD����6�#Ѹ��˷�k�r��F0bQH�ʍL~�R a�ڐ��㢞-�E��Z��E�2��SUַ��yaA�Nշ���b[�CFHp�`b�W~�}&�C�r+��P��bB<8d	➱�t�]�KyS��^�ӏRw�VKE�̄�5@oǿ4���cI�� �/��{����u4�*���(��~=����Y��8�=K3�=���t*��uM�sy<�*)�Q���6���q�و?�Q Y�U��JBv%Ǫ���.�
�g���S�=w>Ӎ�>���K���
o h3%$;��@�"ǟ�h�d�H	gFz�T��G�1�g������@ L-`� �y��;��?�Lfb��<��a(x (C�y�cE�N����,{�'.�O��'n�	�]�/�ǈ��5��84�'�MZ����4�QI�����ZT0S|���4�v+�YA�I�b���y*9$��`^�v,2C�.�m"Q�B�Ի(���i���kf�koT����-?�jyܷ�|�r/SF�M��^���𺴗ON+�9�ũR�t��;̛>?���
���	/��ֵ�y�с�~i�K"tc��Z&N�>�ޯo+ߨ��&�Z)�Z�*{3C����p����yvYH�Bk%N,�a�?=���a���wX�אk�_b��G�JF��~fnEٴ\����.)i@��@w{�Y��jո�b�N3�إ/4��(1�J?w��HK�\���A�o�`)�ح,��3���2��L(�fb���;d�)G��P���f� ���GJ �f����1�Q� ���,��{�z��,	�$�k�u��	_N��NjY���G�SU�^��)�� ͼq�.�y�ʅ������c��C�Z���hp����\��$(��L��T�R��1�j��!�dQ퀗,����-�tb�!=ŏ�4x�uh3BQ3ul��B��ǌ�jAԴK؛i�Hv�*_z� i�g4v��8���j�gBd%�*�X�����9�RιQ�MT!��R�U-���C>Y� ��
2`��^��-H�0	��S$�b���
��M��$|{̓��e�z��<i���i�!���u8=G�����W���iԿ��������|���&��B�+�h<cs���7tO��A)�i!�oH_>��"�,�)h�1��.�U���AT�ġy6?��8�_}g�BjHt��F������b�@-(;"Ir�b٢��q���I/-�q�[��B��U�yQ��7K���`��4/�-�{��.[�HT��\r�'Ǆ�3%�p\V�jF-b^� �_E����ﻢ�P�����~(^ih�.0! ����.�%y�Q�z����2c�>j�J���in��
,cko��fh�!]/s�D�ĳ�nػ�����~ Hf���ˀ�.診�c�a������sB�9��U�zݗLF��r�Q(}��i�����{�:+��RS�d�=���yɯ
�77]�\3ٚ?��� �H�S~��d�a�jr����0"01#Y�b�r�W� ���Wp��Q|�� �oY+���Cr�>�>���fg�^�Q3�հ��9�܈��]%$(TcF~P�9t
TD����Q�|�U��ʉ��վ�!&�������[V����g�Sh�*5�w��؋����+GgR?x9d�|�{xg�z���qh���k�V`�5��3f�	���1T=�%ei�E�Υ��g���%[ �������~6�`�}�S3����L�8�x��=�'�vbA'&K����nٟ���*�T&C� �tpҩ����Q��y��v�x���{�V����ƊsT���+�����?�.��7��P���2�8�2E��"!�5�8UbH������+[�;G8�[��9C�;�!aWx�̩,�;9J�N���R!p ��1�E��`o#.�w"�����U[�\Tmn�� �8%�%�\����T�$D�Y @fS��7����NH��(�v����a:B�<���'4Ѓ[��a��ae��-�r��?~�0W>im��x���ssZ�#��r$��K���_��p-�-p���,�g�k�h��P�AKK�<��Q�ÁK0�O�/;X���u��N�����n���l�~���,�+�v���^֚{Nm(�͒������"1_���όS�0]=$@t�<�M��Ȗ��d34g�n�R��T������2po�\�&Z��fU'���hX��+}T%	�z��O�����W%n����Z0}�;�	J����#�,�Y��N[�>�"��<ϖ#~K{���c~��GF�#LJ� {v𻟘�NZw����}b�!���Į�8ح��kXdz۲�\1��X�d�W6VB���vir�b�g(M�Ś]d�<hbڋ�8��-�g�;�?z�[[<����G������KA$�Bز�9px�2��h�BU�Y ���	<��4ꓳax�J_�;~e(����!+c���	\C�ڋnG�-
J9���+T/V�O�fh�K�I0�?��7���ߝ�ma|)��y>C*Խ�'�,��-Nq��r�4А��m��ءjH���o��o5!�x�O� .5�z�X�W>b��0.�܋r��J�a2k�7���dxۊ��A-TIوd.������i�l@�)�:����g7N�^w�h<|�5�4��O4h���'�Õ`�d�B��$�2�k��b������Z��|>yRᗋՊS�M�����.H�|IL�%���i%z4r���/�G��I���n�t�~=K`}<��be��շ�4:� qS�5C� es��2p��z	x1�������9#0O��Q�{��'�1i�.h|��ف'@ ��!!yH�M��F�%C���3�k����z'�b�=��sҢb�����X��S܍�L[�&�"A���*cR3|=I�h��qR8����X5������g��� �����Y�8!T��q.��Lv�ȓ\Ko���O�ʛ@�ŝ 22�j����Ճ,5��?gjv��[������X�LT^�lv�+_41��7��өh!Q���dI`��p�`<Z�y�O1�։=�^���8��.$/�H9prd����閇�P�I��v��i���ٵ ��H�]�+�տG�2w�5�N��\�o2c�����:b�h�� =�q�Ԛt��&,5��~"�C�G8B���O>Y���n��7/�L�Fm�^3�$*a�9����x����Cb����Ⱥ���G�0���b�5염�X�t�y��o�w�_)۱�:}���'����l�z�����f���.��|�F�0���PL�4n@c�.��^�u/Ӛ���*����?�kM:���-�M�&�B��M韋VKT�u�tV����>��%0��.��NM]^��c��|57!)NSwK�w��7A/�NT] u�\eZ�|a�n?	��+�eD�����#�Y`�U��X(7���p�:��;D��P� ���[řj�}n�|�=����g���#�;R��w�Ym�P��?�,r��09}i�\P!}�r�J�'���,����g��bMع��:֚�u/�$8.d�#�0��3uG�n�������tF'R�B�Y�R���g�f޼�_��4$�M����:e��,�����7��ћ��%��9��O��Bn����|4R��c�
��|��&��iFU@��w��UsRDF1��@����s^JH�̌�^m^x�pe2P�7̾��C@e��$��F^y�L̰t�ZQ��-���V�n�[9��B�����C^�ܟ��=�t�ˉt��gfO���k�~�inq8:R"������:k���X�Zt5.�6F�`�qY���S�9��f7���w�d�r�[t(��!o����؎n�$��Ͽ�tF�u���vcY1	/�(ET,��K3p��^���1��5<BY���|�u��멨m"oP)��)��͹�Ů��^�wS.>q�AJ�G,����4��D')�t[x�\u~��*"��"mO8��U����Z�ćyE�і��8+/)�^~��t�w/�Qڗ�/t8�>�d
[��I��e��$����s��¸�?v����~)��V	S�jZ��'��L>S��n��.Zto��W���Y,�5�Qm����+����wx�P;%l�b��]���U�|�Ḧ��O�O�ᓮ)+�:J�����/I��\�2�4�G�� ����Q���PQ���?ӿ�[+.գ�0����emb����^�˓����i���`��e�g9p���-)�@����Z�e���4ן{tM�N}ئr��J����}��(�Ȕ�q�٫�Y�:4ƟA��`HR����6�!�ټ�&/�O2��n�R&��#����яT[���D�`>�UB�i��e
(6�ao���s��g�+8;�h�i������+Ѻi�U�#S9��hV��4���Sn1~9��}�è~
� ��7�X���W�7R����܆�0=)@�a>��V&,��J�
�^j�u�ؼ
��0��H�)K���OVD ����g�+�3�F��5�lf�����D���3�F�d�,(+�q�KL^QZ^NhV�Gܧ�ߐ�Ze������5�H����oG���y�9��}Զp���!��������V�^�]�Y;ǘe�ֽ�+dٲb !����qk�s^m��u��|��bX �ND$ue��چ�O��3�����Y{C�S��T2��h3a����׮T:�y(;V����Ieh�\-n5�Z?;d	���:�ᤰ��uUը" ���cL��c.k+�)�28���*��O�Ē�%���fjJ��`�X���V�aD�rV̇�qZf�$�؅���5n/�λ\���JK`Ar��N_��F�,���ZQ� º�^���w����v3E��:��(��M.��&`P��6��GTJ"�r4q�r��2M`���~@x�}�W��M`��mL�X*� �cZF�!���_�*�`$x�����Q̩:L�<O���"<)�d�E@�񙒙��^R8}�x��g+ly~�фb�	a!�o~6��4\�csy�ߗ�5*|��m����_��-��{$K�����+l�y����#��ۣ�k�{X��SB��,vS�.�S�=o�Ǥ#s�M�&i��-2�(D6dPY�!�PLq��IG�{����YH������
e!����عb��@�a%}�! �ƅ1.��o�U�����h���k3����������� ���Ҫ���>�'��A.������9}��P�up�L��V�%xn��db.�&b5�w�}[��R��!"蠪Ma��� ت��X�@�N�mdC�ιs���������4ø������!6ҟ��5{����z���7�Xy���Fa%������V��v͘s�`��	�K����.�r�.� ɛ���Bn�Ex�b�]��x���#�$[�!�?�~��Ô��8{����wSS.��]u3�q�����SeR����`�3mH�`�v�ev��Y���:P��KG���u������x���'.0��f�2�i�?rd����^2��>�.���vǰ�%��DN΁�u��,�8���k��J��4<�<Z�׋čbAFsw
�!;J��X�Ag���KK����8Ñʭ�w�EC��b����H������F���S�l���l��?�K���%���P��|��심�K���B���ܢ,`�pw*��'�,S[�@��O��S�_��Y�H��AZPUW�[��i����v���ŢQ���Wy��l5���,��jh�r���^�D���܏��L �z��� �A?��� ,�����%���y��C<��{Z?���I�*	=;�͚-�m~�ٓX�T:S���̚���d��ש��s����FnE�k�k �����K�Ba�:��'��B�f������0��2��|����u`.�Ɍ�}G�,v�X2hX1N\�뫨��3��E8f6��/�|腈�5q|O���}I��Vv~IO�#�0��q���خ'k�߸L�m�)N�a���gi\F�N�D�5x�`]���6�x[�g���%�K�Qd�;��f���?x�>��Go��<�G�X�Xm�QVF�,7�Y}�:� ���[%,1 ֎�Vj��p��YVH�Q�^ފ�~�ě9y邟������E�S�H�O-S�����Ȅ�±�Y5��`4��vi��h�N|He�W	�_!>fs�^֝Xq�l�n2��g���.d��\����x�ʈj�^Q�?Q�� �Q5&L��%WFg�༴-.e{r=����-`������Z�};��/��g.R��UD甪����m�a��0�D|kx�&���кV��Jyw�٭�e�u:����'�G�p���Xc|<�~�����XF9��Q
b�q���w�Cu�z�)��9-��q��z>C�ɣ�[d�[�ԏ�h�����(gJ@����3ƚ��������\�@�q8�����;B�!�0Y�ae�WT�E����ô��v��ϯI} ��ǩ�<a�v��,f�n�ܑ�N���"H�u��o.�9ع6W�c��c�oТs�3��22��C�Ro�}p`c(��{���k���`3�B.��/5O<�itt�c���B,�#Gt��j3�:�쬻��_/T�j���k�ا�{s[-O5!����4q����o�C e�Ǖ�pF5�����!+�v�1�l���)aDR��)P���zkY�j�����x�Z?�E�#X�"^.q*T0�m�G<Ӳ4�`�y�;,U�����"z���2��O���jU��ޕ_���{�0�g�8u'W_OMc�%I�޶~�Y?�����c�[0G��U}�۶)`��#W���w�i�&��7�AA��'!|d7�,u������܃X�Z�<~e5ٖ�k4�\�T��F�5̷C�J��2o7-NpF��a�n�W*��Ťj�b�C�s��Ja��<}�l�dYu�m4��qV�y��}-	Q��4^��]��MNJ�����C����Wg���8�d�_3�G�Q�=� ����L��Z�L�=��?{�&۸b����0W����M=���������rm|����W9v����
jS�MA�xy�+d��O_HpC��Lki����m���g�'��]8Y�0� V6�L��C��Aʊ8%�-b��H'�Gv��K�����4q-�~&@���f�M.�V+`Y�fw(b'cm�JZoN��-��W��JA�#�wK��NAun��Z�v�Nz�H�[��]������a�$0:I�5C�W��F3�/Ȯ�ҫtI�;�@�0ف	ِ�w��;^m�J� !XᘾJEk�;"I���2���q���;����Ҙ����r�\���jΛ�l����t>�p��"�2�����PmO��hHy�F��L@#Jh���%2� u�Ԫ��T���G.��)c���/�m���s6�h�?�zY�?���zgO l��q~�b������
6����g$�7[,����<
bx���t��j#N#]t�ڜ����悛�����Ѹҫ��
��t��/%�߆Z�A�\�i������v�F�Rդ���?2��`s�4��>��C.�M9�����R�A�u�U��,��������/�T�OP����r9P/}�.04��?
��۶z�p4M�%{����`_U2�6i�k$�˝�3�����^@��D��t�d��"w��@q�,t\y��.�4��(��')��A!��_Ok[Kb�c��.�b)
���x]��hm���)
�p�
	uF�79g�N2��!q�-�b?���ă�A�JG�|�f:��j�"��~	R5�;�K����˭ɏ��MrEr����O|���V`�Z�;���ʼ
��D,�ށ�`�<l�&t�[m���j~������;��BԎ��#/������[��K�Wc�����j���5K:����e�o̽���rw�{u�W.6�$���M�䫉�^�'��&����3<HgG������U�>�z�ϗCe�\ O�����a�Ž�3H��͡u�X�t����2+��|̦(G�T�"k	/9&!�G��S� ��X$�!4��D��+�iݬ&V3qH�m��ު8�i����	�C��s��j��'�|/���[?_3 ض���$u�ŗX�r��ɒ�ߙ���z�'�й�fʳ�.@���7:4�����z�L��ɲ���	�PV1�c8u�zvJ�d��ky�M�� 董.x��
�"�M�	q��a;B��-�dFۃF�z������ИC�kc�5f�6Ċ����t6����t4ⲫ�S����xºn�]�[�TZ=���wav[� �}��n��;S�	h\��L�pn�֏���cT|���[�rW��"�q�x~|��An,BO���_V�z}<�������K7��ṭ̇��/�
2�.�#�Ԓ,U����b:��i���MK�~d$����气�ɬI�6@�d�Lؑfx*�#��-т�4����G4qI""����
,�m�d�YڝzKR�ެ{�}�A t*���YTl�9fE��X$�ʺ��(㨩u⬪l|a��`yH/u�`G�����r�n���s��UF�4�
�y�2@D3ɟ@JO<"~ߤi�$�o:8e��Q6�c�UlI�H�qVYwc�q�`���3�"�*�Sh�9��	�-Zt(����!�G�G�/�8�� �Z����%00E��3z;�����3�e�~�-T�͘ٹX?�[,"�f�e2m�NC�g�'��P\�F�'�\�Љ/RVG�q=��&��4
��67g'$��� �su��l���L={�������b���o�ݒ4_e"�\�����^.���(,�Mh���2
�1����e!�a���H��d��g�29E����^�s���z]52��'ߊ���vRw��Os{4��?/��ДT�GA�����B�w�?��¸n�7�M��9g���]�9Ɠ�ꋄ��]�V�}��=��q�ڀI�9TH�͍�M�e����T�{5�Rs[�	EH�od�3�!�I�/�Z5�h# ��O��D�bp��Dc�?k_���{��H�fp���,l����z�	��~?�h/B�)�o�W�`C�e�hJ`�l�&Jkr��&lX�sr{��i=�f����f��h�/ON��w�-^�'���Eh����8��Wz��l#��#t�\�DNG�)�,�wji��+�)�4�T�e&?�Q�� ߲�e����jUHӄ�vl҄(�ء�R�N[`��cM��|=!_�� �����hҴ���c�Z����ԩL�H�jKfJ�c?�����R���P
/Mm@�8E�� ��*�r�81Tɟ}���S�6B��x�Y/�U.%R�]
hXE�]��_�ey�!gF� g}��bz���Y�7�,vK��0��ޅj] D����k�Q
n�W�	����K����`�1��v�V�ip{����xZ,*靱z�L��j�̬4S�����͚�[ى������(pj׀A�P~��Q�����*�w��k�ҋ>Z*�&Jw���~Q��H�q�>��yU�i�J�?�\M�,�Ⱥ����9q����Г����o6ED��s���}M�>�=ފ��E�E�wtx�;}K"�։�"�jXG,ʵ�L�Ki��FaYN�'Q�DI�V�a��w�����ޡ���SO&��1?�����}�I </_a�xoم�C# *dyh31�����m��a}N�֡�.蚯hP[/�11��ۻo��5��
4�z�U�Z�2�U�Z0�=gʽ\˼�s�I
E <nLu<�AY>Óβ ���l�հ��B~h��~ė���֬*˰�%��O�wCV�$g(х̖�����3�}�F�n@u(�=3wHB%C������)�e�l��B&gU����ǳ����q�S�XL�Ox�#S�
����F�gG�z�Q���f�O�dQ>Z����s�HV/.|:�D��3^�+c��5���*83�E��=7�@�9ŹD���_����f7�]�W��<�Q��&�t��� L�1В��~�V��f��P�D�T<�c���(@CKW�m�8�-���(���.�H0L�C��#���U����:Pvy<�g�^�:-;Bk`a�Rqx�e�(KY|Es|u�y�O�h%�On�lV��G�Ec��M��K3 �
)��<�>b����oS��-���� �ԅ��C�\� ��s�N2f ��o����[OD�Ƴ[`[j�d�oo�	�=[A���O�P�M`�}Z�֛��꽚¥���B[�s?%K����/XLr�6�WҴ�K�̰�)��6�R��39�aa_�I��i�	�M��Ec0~`���8�������ǋ�<`�p����ૃ(-? �CҀX�(ѽ���N*m�.?���4�)�?vI�Β"&�P��%��喍r�}n��J?�?u�jMn�Y ��_1�$�]H9���I��lH�.X��t����Q�ae��GB��'�#8�!Y����b����b-��(��A�溲��Sz+�b�u�		0�X,�yh�e��ȏ�wC]�s	h�@��@F��A5Ѱ�����E��%d}�EUiʟ%J��$фT��fԊ.��m�%���]^Y���i���%�-��vԏi�ȱ�q�.�0�vIsv,`m>'�a}t���N�P��Z{W��[��pQ��t��.�����~�?��v0���u0�[��V��}��=R�s
|��w`]�red�cg��`�Nag��h*n��s�h��ĕ���=�Fd��I��R�i��x�O���rG��(��F���E�.�J�__"0weƅa�v4��/@{|�4�c�p)�r�觢IS���+��+������V|��V�抦]��P�h��[Z#H�w�N8��FJ��k����p�y��[
�'�?H��Rz�a�<]q>?΍�r�̖#i�I�ET� �q�8�O����M�fW�4����03%0h����;-�a-=�I��,�k�`��2U�U��M�_���Ux1��<�0Fg�����$X֤g���.k�R^�J��2�f�g,&����"ȷ�  O)�^�����
!��S�R=F�������	5 ��rO�\Á�2�9pN=��.n���ch��v�K�d�4��EβM�d|
 �w��7����i�������{�С���]��z��1�{���d�ٯ�#w/>��Yxb�h���v&��_�V�;*Y��1y����WEH&ơ�E�`��kg�o}�VP5V��v ���{�<���,����g�B~^��zɹ�#��#�^8�,�}��٠Kj[��"!b�y��.Ð��g{��/d�i@_�j5��gáM���5�_��Fܞ^���	�6���"������n"nD�k{��unK����
���]�E����
�NKn�m��=�	*
p���|�JE�s>|�'V��s)Wt�|W����t�i���B��ܛn�)�XS�I��_s�LF���(�ߎ�=�8��H�'��<���~H�yS8�܋|L�`�Z�'Q�Hѿ߁�>:yR�EDBW��bA!��2L��� ���I0���3�˫��[�B�����������_c8:{],Q�	����9����s�����Ԫ1����g�$�U�*��_��;x|p9�ũh�<�S��t��ie�QUр�7�nH��SG}�b���	��0������e9�F�v�^�֋������i�����;r�v�*o=���^�ڛ�'����co���9E5;�L�/�L���2�<�Eԁ���]o���W������/���O^��=UEA�ɢR�u��ՏR:�M���!gn�^�G�ڧ��d�ˢ�q��C5�:�"�c'𣺁�a�Z;���MԴ��Eĩ,��$]�d�<��^E����`�挊!Ө۫D�����@����<ۦ]����,3@x��Y�%9�S`�y��t鉔+���ZЮ��Z�"���w�[?��,EԶ2�wУ��;$��L2xԻ��V/�2ؖ*���z��6d��&	O>����z>�-h��:�s���)}y�� �?^;�,j��M�U�kg�n�J�&�&��;[J�� ��sz��9,/WĊ��a��b�dt�xJ%�*�܋�Vr��@��`?Be��'ǖI����qa��tS��26]ջ�&H �]�`zȔ�)��F���ve�G��uȘ�Yۜ����	orK���j� ��+�Z�DpN�hA�!���Fο%�*iLK�08aC�c�\��V�Io�k�IQ�,���/.�>��೾��y��g���}��a��Be�K�+i�`�a&�\��.NO��IR�Xv�\��,�>fz��f��=�n	��o���-[��B�_���$���B�4�r/`�Q̛S  ĆTw�(C� ��P{��N����+r����·8�ҷ��#2l��!�<�_sބ������w줙d�^���q��;v 0J�K����t�C��ǔH\����N�%g
n�*�F�2���Op*7�r���n/���{JoږY=�(��Z��=�"������G"�[�
�;��PD�d�R�y$@�����/]��Z�`�È~Ј'�@�a����):]��A#'D.�h��%v�C��K�}��N��fb2[KGI�q�g������%�D����J�8��B)w�o�����ߑ[�X�ʨkc"j�*�sR��U�<|��у�)�Mc�L��^2����g�{�����h���I���di]8޽�x#������j�ow l����u�?�Y������n.��2N�^#jUPf�j�Dϵw�3%��\��}�@]��f�����e
���.c≴k�ߥZ�BO	��w[������0'�����"� �tLN|��a�_] d���dt�����C^m{~�.|ͱ<��uS,%��D�U?ڛb�>��=,��&f	�Th|-k��Г<�O7"'�ho����C]�-�rs'��W)�pA�ײ�c�l�*>�U�=d1��9����ާC���e����.t��&v�琟ҿt���_@N5��3ɌHG�%9^���m���w�M/�CZ��.��esdN��"�]��Pz�(I�K�1w�	�Ǆ����|\H�����$Ԣ�ʥ(1�ˋ��ů<��)sf5�(�]]
��~g�]��y��c�;���9������
�Q.	t�9�ڿ!s�P���}gIZjE)PtFE�zj�T�)aa�����z�L�M�~5"u�d�Bcۑ��rHfJ��P�A)��B�AT�wy���5�A*|~v󬋅��Ѝ*~���t�o_�/S�g��z��i���7�ƒ���O��������BH}J<h��� �������ӄ�W�En�	I���V(����Y��C��9_����(���v���.�x~u����	&��A���&�dӵ��e}R�0 {/J0��#	S�0Z/B���З0]�p2�b0,n��6�E&6h��a�`2�QL�o������ ̄�Gjfe �)�\��I��$�Q��/��ҧx9;�k��Է7u�W+�>8�փeG�=eO�'	�B! b�˙q����pz�{$��ڃ��5���~~��°�P:9�P�KHR�JLSi��ę:&A)/ϝȋ��Z+wFxo��~���˱�GfXCc;�� `��́i��rG��I ; �j�)��W�E8/R�:o�=��Y�i�u���x�@�v*ӭ�v�N��mA7�^��1�\�o�н�!*�`�0%���h{��7&�݉Q�J��R�)T���<�S<0�-��+����,)��{��D��	�$��q�~cH��Ƹ��
*��V�g>����ۅ�D�]=ֽZ �@�8��o�j;Þˇt�T� ����"n�ň*��'��˵K�+?1m�|�(R$�́a�#N}�1��yh���u�۵ȗ�-[Rp@�DX��n���Y� �Ö��`F|���Ft�U��D�� �#�!>���M�1�ܘŕ��۝}�	�s���Zɡ�,;f<CUѮ�	�k*�$*tyK�M�����!��Y�k����Tz�66�2�cgdN&���H�r��9� ��6��)Y�!e0�W̨!�\��)�S*ζ�yZ���͡"C�<�����+Xְ�9���������ν�HJDV�=���I��:����j��^w�l�U�i�	?�ԃP�I(�L��޹�!�l�b��͏D���;2�J��9ak@B>�<�(r��ת�v�
?�ToiP�~/h�j��IvM�i=��lC�~?�-<M�cfu�9�/�o�a��A�[9�e��[�~CE�fW�i�H�܎�.��.���}
��p���5,���V֜��x�L�Z,�G*�a�?Wg9�Bi�jo�x���;l��gOT])�UQ;�\��
E㵉z乵�{,}k8?U��i3ڈ��&@���1Z߀��"u�~4�z����>H���(�%!l7��v<N�5H&q�K�2��*=�`?�_%�����/�`�V�&^�R��~ 'Wy��7���.X]ycИ��<!Zݬ,�6��6b�K㖲�5H��X	���V'��z���-�<�r�-����hц���t�.���
2�����ِ_�YLTt���[ګ��ʦ{!�gG!����c'��޼G@Ϟ��{_��{��ʩ��|���`W���1�Ԁ�?�N,_Q�>�����יAI�@��3)���,f�̹$���c��)l2���%�q��T�P]�CMip�0�!{B�l���@�k�ԭ����_�R�uC�>��k1W�Nfŉ���kv;����:�o��|*(8\��3(6�[�Z͜DDVN��s�p+l����ڤ�.��}����*ؒN�M*2��ۀ
z�{6o��8O�T���5�5UB;Y�:�-�qy���<n��Bٿ��Kq�������A{�^V�H���~�mhL{#��/���C.2 ��CIʷ1p�H�T/q~�cO�Q�֚ �u�@��¶n�p�5�l.�� �VEP�v��$f���g�\��l*\a��%�m�%c�]��ξ���J���3�?��^���^��!ϰ0)�ָ��]=��;.������dx�;����8��$������MRDݖ�΋�3%0�44x��2[i�������KR�8y�ɺ3g��#*�H���f�"wXE!&������I��]��(���	W���܄`���푬�z�sW'E�y?�N�{��h�<�u[5�;X���9r������tp��z �O��+�0 P딧e>���M
Y��k���7o������Vhi�2ބ)�^{�#������]�MO�k�wX��V*���)"��fǑ��>�A�28`�@*~<J�z;\�P���⡤�2����J��o�rg3o�x��T3����|0�i��9�-;��O�z���9�1[�?９I�:0����F��4[n�Z�>G�~A��"���+����*@cj/m�A�~�R��9�6��1y�_r�>�d���<"j����4���ߦ�1���������CJuW��Lv���q���z z
P�w	��k�8ݎ�6�
����Z��T�o:X1�2�pTZk-J��c�;b���f$�RZ[8r/`lj��4��K�oK�!�iRk�1�v��{,�'�ex���B�ތ�٩h
vtx���և:���`�]�i���B�	G`]�3Y���ܘDH��+?h���I��bRh�X���P��[b�h>�Z���|��T����n�[7)��N���C]w��助�-�N��Rh�R�>����jd�(i�r}U	Zmr�����7`.���f���>wf�ǫ� � ��+�F�7�3m�&�u���sUw;�Tn�O@)��I���o�23Fy��E�@x�pJ<�TT�$i~~�WѮa��:鼢��!Hp!�&�t}U+�k�"~�������'m�\B/jk�^��<k$�'�C�U�#�����G������������@�S�5ޭS��@�+���-�H�4� �ڼl��� ��*QЙ����
���Iy�,��X]=�1�o���M.cd���)�
<S�����#�D�ѩ4���� ��{��Rh��ݓ�TNcSsi�9��M��_]m�9*��m�
��5gx�op�uc��� ���C���e�7+���N�m�dR#�X�*�>���`0׭d#�O+��D=L�3��R�X\A~/@�z+�橘G�n2�����M�w�����Yԛ��l�
FS����( v2`ۘ9O*L�D��}d�6vM_G���/��_c�~��6Q�����L-�NroBHG.�j��`^��4
X��'*�%%��T�͑^�]\	�;�о���_�[^uC�r����M�b�)��ș�pwe4�9r�)��(��N�g�_��!Շ�P$�c�ACSٹ%1s���k����Ro�g��K8
��ȍ+H8w�W6`7���@$�����
K�ըP�!�E3�@��pL2o�@��~7�Jx_q���Xั�z��ZS�#�@���ADcO��q9�6#���H�W�G�M�4h��,A�6Z;41OY��ZMAp�R���a�Yi�3�{H��.	�$1I��>��	v/����u�z"�w�$���GR�y�Z�8�ҳ�-�D����T���#2z�&g=���V�2��������W���Y��uKΡt�����fT�ʪS]�5��R]ކ؟6 ���-|�q^�G��~|�k ���\�oG� ��H�˚���Ά�r�N�ձ*0�0
3���a2O�@[	2	���q>;����K��������w8<F.o����e�]�\�8�]Ѭܒ�.���!�v��J��bR\�+�-�r��M9ZE��v��>�u�F*�jI�x`�3�w{�M"���Ѵ�%MA";�����;�m4�-�* s;�*ᚌ��D)?���3��s���������o���V�ђ��	FB�Y[��!P��o��D�/ТP⏽}S��'�����-�Z���4���I�~��<	�T��7C�D�;�����,���$�D���j"��q���:U ��ŵp�[Ս��ӛ��r
4˱�|�+�vyf4����Zr+�6���)�)��ʤ6M����)��D��-C	4·:�^��$��ze	��̺!�_��	L^�goh45�����8��z�"�a𒆜�n���ǟq/B�`�,�6kh0Zv�0�A7�۳�R�bF����G��i��!Ъ��Ws�P�}�O�s"^t�*&�G��ُ���.}�ܣ���t��` u�����8�*?����J|N�Q�H�����>�&tͪ�ēNƕ�� :(2!�$�4�G��)�=������tN�UQ x^b^����/>�u1�ZWÃyW������fx��|�%&�l�d�;����-e𗔟�	��-U@^c�'�__L&(���`���9t�*�ݫT�W�ǭ��F��LޑxZ�~~L��say��%�{���G|���$TJh(�r������s��_1p�SE��*���$�(��d^�\h����1���6�K��|Ge'��l�i�I��R�U��Z/)0�r�&XF�.�#ȧ�!�'U#ƀ!��KDt=���6��r���̍���?b�_���V�^�����E$/����d�B0Rjy_ߖ�<
6[i�2�Q�Hc����i���-9���0�x�6;��G��R���\�/$B˺k�{Go�[u�W����%e"�ª1ԓ�u}��#�H�ۯ�ne�n�
�bo'�Q�Q �*�+��9�Ѷ�V��8�v��n���. ��I7��[��x��������	z���~r�t�D�$���튋���;��+�+�������諤O�d����0���{�W��Y���é�� s�HsE�ˣH(�6�;�\�e�4dLf0�ڸ�O(����A�4�ok��b��0:�F�M����`A��N�bs(o���!��i��JQ�-��e�0eǱ���B�I����/y�;2Eu��B�7/r�'<J� ��˖���*��Yz��]ĕ�"���W�,c"S����s]6_3`n"��!Y�vZݛ�/d_���c��VM��+[Am{O��GoXY�Z��16� !�[��ƶ%^	�9e���YK��`��{:�~M���-(��$�E}8C�~$[vFP��`Ԁ���S���NF��ZI�ۨ��Бv�e5ps��9%����0��ؒ��,#����0C��DE�k�*����Z�l��~j�b(o��t����ת��@u)2�"���ՙ�7�#����!�~@L���~�*�ld�y+�����J;P�/#����
���I�LȐ�)�i����5l��M+}��GDQ��e�ꓺN�s� �{C�m��I����=� �[��>XL��5r��F2Z�����?2M�_;X�@8��O��������0�ɤ�2�sG�C��M�s�,�C�,��e$wN���3��yb�])�s��+*�P|�/�&�z����+^��Ȋ�������*��6b�|�$3Z���:�j��3l��,��w�`���	�آ��o$�?�o���H�i��S����m4�����W�%`'�p0|�%r�"�����=q��e�_�3��9D;A!|V�}��*�\��`��Q�:'Q�x�)��i��Vs�n��I���#�� �g�L�n�5�3 Z��ˍU�(��ɠЕ#vZ���J4h�e�tHM�$�l8�<��n�[���#$ra~��}��:U>��Ŋ�
8�WTZ4���OˎJ�N�Ü�r�	�p�X��TTŝ�M��,?ba�mc��]d̈́#yxC� 5��:~=-͉B�3@�#"�!�iN_B��r:��A�#>�	!-t�Ն�(��[a�(����3X�<��P��m���ß����k�t��'S8a7L�K����1jx�:"�p h>���gd=la	��:<��a䀝�؅��p7Wl���ES�2B�6���c�Mz����tMD��`����ŮW�S��,1j�J�`{#��]�`��y�K��i/*�PI����IA��.���<%��0&�EK�'ѐ9��k��p�j}8��_�h���P8�p	_����j����x/���W�u�@��ߴ��)�@���Df
�4X�p_��TM	�}m�y���0���G�,�7}�TTt�J��|?���a�Ii���Eƫ;N��
f��s,���S[�D�I�Ĺ�t{��g=Fg�aT��l� CZ%m�X�H	�"�Ҝn�ՠ�i�S;c�$*�@���±3L�xba�G��"��2������>U�/g!����X/�?��dt��V��E�=₷�$��l"#L����?��C��E\���_y�̓��3H09��=��g��n�W��s�T)��5\)m�L��~5@~��9�(w�-ɧ0p�{�䰅+S�DY^u9������:_v����|:���Ӧ*i�k�����tg�Vܴ`s�q���M^W�l��S��<\�?��#�I#� /$׷gy}�����P�%a�{]�+��χO:F�՜j$�I 	��B7
[��}�U'/�����
ak �zzT}�r�PJt.��L0�&���m�ٗoރ)��ͮ`K]�|�~"Ӷe}.<�ʹvgq2cj�N�T�����l�9�#��Q1��BE�ĢA��h�|�����4��{���)'ª���5:9's��P$r s��PI�]t.N��3�&���F^
�[����z�~O��/��ډh�׷F6LG����d�R����cc+B��9·��Ć=) x �%�%y1���e�t��5�@�svU̞�M&WGj?�h�mo=�\)�(�M��@֚�d�DR�i��یn����n���6 �9��o6uV� ˪����j�)<�`��m��,���uq@��Z^F�' 7/������eB��7yq���(l-נw�D��&�0ٻz[&���*�H��Н�9������:�|��f�nJzz��bZ���ş8�D�� ޙ%���B�))n��$�K�0�̊-�Z+_0 o��>4�;�1�A��K��S�q�o2���bӋ����^ۧb47�Ԋ���:�{IE;�£VK �e1�I�3��p��J��|@���\���LX��T����][��$�#ڷ���M��9I�$����'��7���-&�j�O�ƥlL?|x�t8��BD��ƶ� �j��Q<n�=^�@���׃����uQ>�w�=���LNjs�D<�Y��� [4Pr\���9`���h���	�݂��j��gɍ���"�%��x\(��@��nJ��E���V��r�Y��k5��� \���'��M8z~9�9y����*�9m��+��B\���:�ia)$�{�]�[���hKP�w�n�0̠ZπpNv���0�H|�0b�)��ܲ�(ZMH|n����@���~�:f�O0�7U(�����1WM���$�IN��K=,���x@��,�����Y/;�>1'�����W~3�������հ�#�jR��H�2/]J�J�4o�n=���=�*��#�g�z�dr�?p*�V�T�'�E���ȑ��J�	7T�zY�bZ>�}��KO�4��.dᯣ}��*T�c;� �Q���5W���+.-�=�f���\}�f,���O���[1撇&lw;>SRsљ� ��F�M3xn��!ߋ�o܂��}bwO'?���G7tvy�\?u9�u�q����:`��l��y��kr��WpV`*��18s�|�DKaPǫ��� �����^F��d��U��D�?,��&��c��N�)&)/���n� {^v!.�-�O��_��.P�Ȁ��RԶ)2˔o���'��?kL3<S��=@ڷ�H+�]x�58���]-�6h��$����Y��.-q`�a�~�k��)��I}x��.�^)$jO�t\
Io�OF�v���y�b�R�U����6��j��~��:s�5����+z�1(��هE�8���:_ͻS��p癑co�2�l.,�Թ|���"<=LDw��'����#f~VK�����KaK��t`_��\�tD9��)�aJ?�����`�憞�ĝB�����D(��������e�j*����5@ʔˈ�1��S��] K�J�3b@lf��KYq�Z�D�dtU��x'�~�?U�Q�+,b���授yn-�u�6���%�UX�7a�:��yi�s�x��g�K-�]����0�^�mW�%�b���8���?ש�*�"�#�$���Z�g�l�{_	?'RM�s~�%���֏H?��ʺXu8�O�Qq�X��E�`��_TһO�JEGm�YE���s[��y��������:^7�Z���65������7Mq6��9�SY�..�:7��##`v-���TbW�.�=ֹ�yǢ�\d�N4���uB۾A��z�%j��,Ųs�Լ��|�Y2!��r��П�Rҕ��1I����{tr��ã�E����kAod;=��}._8Z�yT���2#��ڒ<ɯ�?e�#��K����&��S��n��V� ��ŦD�)[�a|Q:-|`_ε��QZ�]����#�L;�1�pp�/i
�0�����fW���