��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>��������ّ$�*X`F~�������><06�L���\�D>�WҎ�����r�.~O�I�V�X;w�G��ts��K�5���t�7��R��пr�.r���x{��}sbeq�XG|7 ��$�ڳ&�e
�=r�$��!錋"���ۆ[�8����lr���8Yi��9���eIE�(Z�)��VJ�j��?~�	��c��R�6���/�WC*��B�����-~��R���$=��&����O6�F�~gh��\P:�w�o"Z��{��ܪ-|$�EA���ٔ:�_JFJJ��S�B	*.�a�ꇔ�@�/~�WC(���&q����?��V~��A������(}�b	ѝu�%k!gŝ>�I8�s)�u{��>kp�Syʰ+�� 2����=��D~0.i4��SJ~��U�h��ERc;��@�p&)Aǳ)��� hU�`��ߨ��a���L��L�D���ŉ�k�^�9	U��X2,���-�8x����tg����;h���K��c곚�K �M�U�+X6e7%��4�;N;��0'�2�C�ڍ�X����j'�]T]��Ec�����t�(�s��-'���I��Y�_���$.4�6@wx�w�Qt��vu<չ�Udo�Z\F�sW|��M,�dq�9��4	Q�
Oo��u�7 �^[��+̮�P�W���h����F�K�j�S�?����v8���L����a+��7�����=�/��L�����ථ.4������~�T
�PI@�N��T)���#���]�y�8łe�$;��505�l�h㹉��^�G ��*�VΒQ�ru4�/{�DNe]1h;p���-�q3{~�&�c�L��'��L-��u���бig������������&��^v��uN���ywq^�v� _�@k;YY�� ��=��Xl~/����[?K�>����;d������*� �0��a�B�Nj��D;Ұ��N~ۥIB�X��.d�je�+�MZ�^������ഽ�I�hj�2M�����L�Mt=��VtI�.����#a��������ʆ�qGb��em����ԟֺ�g1�Hu?BԱ��j,�_�Q O>8���ӇX �6�vs�9���2n�F��c�Pb�t����By�d�����ݵ�>����\9�$7�J�����hI*��@��k���]��3-x `r:L#L�0b�n�崜j�7��A{ �~ÈYq�:�	:�����3��rp���'@����c���58A�	�mrd /!��ia�rm�O��JSHL�8��1E�B���cF��a�y������M��4��ra�'�w�E5�S�.Uu8#�ed��oS�4d�ĝU�+�� 6�U���u����.��P�3�fK1耿���-3Ӛ �;'{��؋yU�yuڨ���#m<32G g(���$�F�\N!�t^3��<X�W��bq����0
�G �2#�+�!"j'�2�����k�V�h�`�AF!��Vb@����q E�ɷT�v8i��٩��9m�����O>?J`o���xEM�H*�9B�%�\ �t��]��/�у��$��z{.cN<֘�G��v���$9���	~�OI-��m7L��V��0/�ɚ9����*�u����ER��J��s�q���jyDl�c)Gy5��MM�A�����������7�j�֚�܆m�'�o
�z��:��-X*g2�U��'�K�C;�nŐ��*� /��@�1�@��o�V���.�x(⌂]�g����E̛L��� N�ɥ3�aǞ��o��[�qIͨT
����d	����f�@��oWu-Y���E�Qz�'.����x�S� �|�	1K���\V�8�̼TĹ�/�"�O��<����g�_J�\�'�(� ��X� �X���OPs7
�8$̸���vc�����KH�ei�	�=`�E�yP'���țVx����@�yS��V��\ �k�$(?AM���j
TD`��5��F"�^G`b�Y��*+4?!����58���HI%�Ń�`�rS�4����'��p�|'r�.�nO+������m�^&B���G���Ķ�z��J+�ܬo%�}WE"��7��:M�8��tp}��Z�.���LY��噆Ud��M�O��A<q�mh/rJ��@�6���8�a���ԩzW�_�z��>��w]^�<�.I���<#�'v�Um-(��n6�wz���4�ip��Kǁ 6�n�<���m����I��i@A�y��l��Ԛ(KovV�,"@��)��g��ߦTHV�by�o���B/`�^�»��[}����K&А�v��L�O���_'2��1�2@���R�tΥ�	��g�gj#�lG�6��'�:�f��Kf2X-�.Jq3�G���L�[��?��V��7�]�aAn�q+xQ�?$�G}�:��iwt�k��{S�w��S�&�^\x,��O��B�7�J�u��=�rM8�I:�V��Htm�7ыb��ו�
&?�M�Ȏ(\~�k8ݕ�8��d���?��̓DUؔ��ą�DK�JG��<c��*�q�3��fǸ�N��	�L�dZ��I��;������ZNZRe��K9���Y�Q]���p�xX�L��J�@��E5w���$IFZ���y�p�����3E}���IX��ɆeEW]�>]^G/�0/�u(Z2A\)����6��o8-��7�I�G���(�]�`z���R;9�M�Տ���u�!�.��R��1�ˁetȊ;R�K�e���Xn��p9I����&��q�
G�X9o(�7�ށM�;ܮ���*��XF���dūOtp����%�MT�<�Kr��h�"�˪����2^�o%�v���@�%��Sg�Y��j�eY�9+��� ��d�abTgj]��@,��lĭA=ytӾN�G� ?D�:�V�Ǩ�:���A�7.3�v*D.��d%#5�`���l��E��
�k���U���yV8�2A*����q J��:�T��o�����/`��� T�g�F*�4[�f��hx�yOfNIq�z��[5p�S�b�n�G�.���b�e�]��3�6����{�J����;!���O�L�&=��ҺoU_uX Z	��1��k����O-D	u��������Z���y�%�(�J�F����x�1]�g���t�4A�T��Ru������_�q��B�'q2,[�al��=Z��W�2Nz�"����ɟ�Q�~�Y�7�:9n���R�-p��;8�ð'��`L�<w�u���J[����"I�%B�B��|Iv�vV�OQ��G^��w�5/H��Pc�f)�7�*C�FCi�j��c����eY٫M�<�=9]�������|���d�j޴��u����D����*v��}8�V�������&՜���2�7���S����Kd�A��p�m?�������F�E%<� �_�)���k�KT�~��T�_��v������s��v�ы�>�W��}2K���`�$�k �����^oJ���
ϰB�*�x��~��_�7z�;toFDrWg������u��0EE����w�A)�C�SJ�M�Rn(�X��N0��'au*���`�m�3�>(� �TTd/�� �E;�D��L"��)$
�m�Wl�O���!�� vC��yI����^5��tw:[`�����0fH�$��6i:�df��Q3������.�L���<��"ݺ|���s]P���K�L��W)ۗ�r#�rԎF��8�_k����d��f�)0���^N!7�acj�T�A$�1��'d�S?������Fʟ{@-=���i�r�(1�[ i,�����ǥ+�D@#!��M��R@O���4-Z����t~E�潀8~b�	����0��]��ا�Q�TZ�����s'�	�	��^��,�_�J��b9v~�t-1BF��uRH����L.Wc�W��C��lj�k�"3L "&e�`y=DK�=I+��h� �����+�w+��z�a�"c��kU��s|����$E)��vY�۰Ȯ�h�������݁`[o�3��f�KT�tC}�$cxO����P�v_~���_��c8�R�s'h�p"so�Ҡ@y f<���x��n��lA�9:�H��h@w	��Ӭ����7���۹�oQs�UT���^A;a��wj���8�[�cL�����{�V����d�(!F��w�}��L!.؊,H��~�o�b�'x�9q�L�����X1H��F�3����ޤǮ�(U��,���+ �˨΀� n �RBc6�{aT�Ȟ�^��(ީ��D�����+s���$|����ǚ�v!p�U�u������F�`ox[���N�O�Re�o�x��jo�B;�	呰:qa&"0ݜ׌�V=�Y�o�sY��B�3���h�ѫ�G�[�fT'��r��۳"9�c0��º�K�����j�������T�q
"�t�o��±!1�c�!�hp`�����"9�e�6��3�n(4$ݪ�O
A|�Mȵ2ڨ��UZ>�U�V�ȏM,ҵQo�����<����@Wh�X��{R:���1��
���%���=�#A�b�'}�%Y|8�e]Yԑ�k�f�O-�@��7��֫���D:Tm��O=�1�ʇ*]�=x+^ΝP���:�P�r�U�Q�}A���:��N����|����@J,np�Y���0X o�p@�{��?��A�5�EA���ͅ����N� �BHĹ \V���0��[;�Q�~���(P�����=j��3f�r'H('��O��|�MO�hUϛ4� d#$�����c��4�b��V��)AD�}_���ue�چ�Ba��`<O=�3� H�[l��m�ƿx���AW�0<�]9
K�\���	P�,-�d�tXç��hJ�Jvm �Lv?8�i�KH�ܥ/7eVp���)H4��`.88\�m ����h!B�1XL����=���&r&�G%��n̾P	��J�;�N���i�7F�W"�^�[3}��|�O�tH�%��@�]R�v�^ɺ!��܄���#פ��u������ȳ�cY��=�~��0�s�x8��@�'� n�ŋr��V�3�H���wƵf���ȴ���ă��IWl�ޢ?���p�^Da^�q6o5��]������.h���jn8
�x���a z��SgqO�A~�t��u>%ҹ����h�Fk��^4�6�Jm�6���Ə�_���?S^�}�
�0�=��v�w�_��mq�J9��9�4�[g�����������&�W�5�����Ⱥ�K�X�H]F��W����?�b@�r Z���e��$~o1��F�Z�anEjᐠ��zԱR���Z'W�o7)��WNU6Q�K0W�X��(Q�:Y��t'hz���v���:����2G��vPbP��K���~&�]@2�� C���a�	%�o��L�j6�MK�m�yT��P������BN���3+�Bs�;
I�:�뙔<�n=dDL/�}��9L �[�w�r�+�x��3}Tbķ�����!��l:������x���9�	�0M�rw6�����5���!�g7+i���O�j��z�x^�N�᷾���Et���*R�1�K�<���z��{F�e�u��� %&&�.^:�U)���ώ}ɚ&������YT����T����
r	Yh.�%y�R��cߊzh9:#�������v^��������#�J��f��`.�@S-[�Nx�������}�ly%� �5ˁ������8At��VE�?D<=��S�*NZAɀZ��4$W	"!�\,d��Z@�r�Ĭ��qU�~���"���}ei�0*;<���w�a�%�]��G��|�O��:�����8�ۙo����բF<�L6ȽL+�#�D��l���~~��ӗR^�Ԟ��U+��U��{!n��hR������S�}s�*�D��˚������7	 4n�C�k��B��|xT�e�ڿ].#�V0�j 8�h��s����P���NK[�3�+R~�U�p��i��^����G�HM�u�� �My-uXPW
(��W�-��Z�f{�d�I�����&��3�wtE��۝h9������5,�H5,-7�:����85�9�Ϙ9��&ƾX��?�9�r���.f����X��dY���i������s�_��\�KY�
!8VRIҿ�k�" !O��\����3D�o�q�[�g��}�u�<��*�^��U�?�G�=��(+��\	Ō��vNB���s�a��I�Q�3�}��
�<���hl�`{W��\	ȮĨ�錫��e�c8?v��f2�2P������?�2��f�g��rD ����$�sS��.s�FF||��l����c��w��4(˺�n쒽b ���^�|��d�/��Ǖ4�u����w%X�W�l��E��s=\P�|��`���g{ҝ]��������gR����+N�ՓV�J�d;iYϟ×���Ш?�ї���;4HDy?�∡`se���pޣ�����#���Fۋ�j��\��=���S�׃�eh�򽕍��u��x�R���Y��xDI����C��|�)Y���k�%\�6����?M������h��� ��uߟ��)���y�\g8�k�~F��F��j��7�$���w���"0%X�1#�W:<5��x�&`5=f+�n�������Bz����z�Ɯow��{N��B:��"&��&_�&bH�J����������NFp�X�q��G����8Y�DA�j�u��s%�1�{ۋ��i�9Wla�޲^��~ѽn�u�
��Q�W�"S@|3��*j�����@(�#(dl
���F#�ouer�>s��X��#���� ���^a�hº���k	`�Q���ɓ,ɮ�2��[����� �C��k*�b:ȁ���Q#S�Zd�=E�I���wgkWR��m�ͱ�9����w.Hq��rIT-���,qj�3+���3��Z��s���Ȓ"�Kl�#P� �׼�H^u��Ð�\\�/�"�N(���!�_e#O���N��<ԩ�w<�[9���8�Q���>h�t]W�#�n�qo�qH--�>u-0 L�z˓=��I��j�d'��_�
���f���=��0��	����2L�������ta�r��Jۮ���fk��]&)�ԕ�K��D�!0�ҝ';�wK�������0U����W�0[�}f�Kȍ�U�W���<�t'�B�F?��j�K��q7:a��.:c� �DzPi�Kn\"�N�R�v+~d�GSk�@�a�y5�z�˿7Ԉ�l"k��o	T��LP�p������
u&��_�)
����#N4��d�}+m��=ݴ�����P�nst� ��\�)Tw�G���k���EΏN�i�Q	Y$��Q0E�4�*Y#����)W�U:N\�K���U�b���Ζ߈ť���Wj�A�)���mk��>�sL�N������'7Ҹ�[�W�z`���'�t�W�fp2	����vgV���t߁)�Z)m�yxH�d���kVc'U���um�L�H��H��Qd�<r�#�%ʐ�  G���2�3N9�T/�Ʀ��զ~��"Y�	 �}Mb� bZ� �,b�lc�'���k9dy���fӆU��U��;�$���0����EۃkV�gJ�~+"��#�f���
���
Π�>����d_y��3�����=�s2�%"s>(U����E�,�e���Ӽ�f:���;%]I��!�t!���Yj����nKR��SW8�}l�S
ʲ1����b��%�U'ƥ:�@�)��*���q
ea C���ĉ��U�2lK���K���ZPz�;�/o��X�h�f4���u 
�x�+I*m��qz8x��e��!�$b�`�k�:�![���x�OH)�����!Ɍ4���=|}9#��峲�(]�P9]�URl�w����?��LSҮ�E5�a5��x���f�zl��6�e�͘�OG��\��/5���}�o�j�"�螚�W{č��0��r]�]1��,Ye�A�˖���-�-g��a�y��=�o�D ��(]����h-S^� �u�o���x@���L�p���=Ъ8��&ql!��>/���7��SC��r;q�
;/l�V0�"���;x(W����r>ILM{Y��G Gi��z�@�����
n��Gi)��`M&3T�Ϲ�k2]��~�n�y܌�,J|ܚ��-?�b�P%��(�d��1׿E)�'���r����+<3ŏJ���z�e���O�W��`IT#�>2m,cmCOq�,R&��<�r�TW���_5-�������vxqKy�����	��u�`�H�1d/\:}W��p�Ĩ3Mۓ�&��j�'�1���t��j�]�8jS�Ά@��\�� ���ύE�&M�|i[a3�M��B�� /Lv�gͥ1u�a#h�֠WZ����{@@�2SD��,�^O?���bH7_²򋹕~H�u��q�)Z*��0�jz��*���N�1>�e��#��Ti/9��-Mܞ�K�+?�Qu���OH�����h�8�do�Wˉ�_�"w��`�%#����DNn����n��?��+����lz��B��K� ��5�)��o��e�ąݼ<���IxKq�f�{��Z#�D;��cY���=:Z��fCD�X����Y���?S���Z� X�R�;�v�7�������pɻ|����+�Bat�r�T�I����Y�Rm�|P �3��m��TkUC&�5������sq��'W�aƔ��-S^B�V]��ȧ�qX�<�O���l�u���F�$�ߏ�窖�4�����\�w��_�=4�zɱp��#��Z��爰��D��]WdL���=n����O�=Ȟ�����Wy���9�u��q��~�D�@Q�%�i[�F�� ����姷�X!)|�T�Fj�^��oh������-�&���&�u�~e��m�s�����٬��k$�"�
ʮ��Q �D�@�F8���	_�i�߿��`�!a�E��˿�;}#��B�%�����gâb�4�.ꗞM�6K��5P������"�o ��W���ܑv����s�i�9'b�:g����	5AH@�_��i�n=���6�n��P0Lx���p*�A��K������97U5[i(F�W�NMKM>A𾧤ͱQ\l��Ī�������c��������� ��1��Ti��!@��� @3<��b��4������=�iP��v��J7��v�^N�AY��qn��d(p�mb-�|��ط6��r��_���9�f���B�"�]�Ŗ� �h��/
�����M �O?��)�����l�`�#9<�@J�iw�+�eO'6��������C����FA�dH�-�{̦��z���x�cv��(�v���)e�W�=yV`�fOs ���I�r]�'r�|QFR��N��T���խ�=��\)�|�&��*���M7;1΅�YA��	߁k7!B���^��:q9�Qs�4�q�t�;,b��mÆ��q�4��P:�2���cG."G��m��;62htK����/b8�"��red��)������9���^s�9ܠ�6>'
�Q�����-�@o���p�'[�&�@��N��]���퍛��2A��L�R6�ў:���}
�˨1�A������)���%!e~P�����p���Ο�׸aI��4!h�)����xV^�o�z�kD��-���r��"y���XU	[����o~S�N�� k}�"�x5���?�%��l�s���2�,Rȕ��p(�$9H,S���v)�b{8l�Ʊ��=�cp�0D_/�u86�Ơ�?H^�J����M�<��Xfw���\Z=���.|#�E��{����sQW����!��>v䵠CaVe��\;Z\���m����"5"J0����$[����P�,���D�3�&�[P���']�h�:³�w�0��S����j��{6+��%��FطxׇN
����g�9��[An��	yԱ ��3ղ�'�oar�	7�����\�ĬE�kK`����D�,��ih�����,U�I�5�c]=�}"J����}�|��o�z`NG���Y���XW^�"X�֌�`�b0	w*�c������y��h�1��G�7�T�v����fwyn!�;��?!�\۴Vr��_G,�����4�R���V���Kw˛�ݯ]�K4��[�H�ɣ��J��c���8E�YD�AA����ԄV�G��_H@��.tcDA�˳Z�/b���U��)X������кF��u�{��$�w�y�!�S������dE��/�A�Fi�D�"���K}�ڰ�>ۼhmӵ�'����X����
ʊ�1 �.�������G���@�����Re�G��Wf��[ӊQ��kO�icf>gzۥ�[@�g/��[�5��NX�8ag��|ʑc�)�"�+����ـ�k��Oi�{v�J�?h�}�x,��b�u�u8W1K1���Q?pd�5��T�= ���e���B\�76�\eB��hErr� �,�b�gl`ao�\�������Ό|7P�/m�ek���������@�A74�*�e��_�7�h���*���Ŕ��D|'�%pA�V���>u6�"�4���@⏬�=N^>Y��V�yr�4J��j���lcVL���t{���Ml��)c��Z>��Ⱥ~��l¯�O
�䘮΁��4�V,��d�+��Cku�A��T�� ,����w	_����cZ~�bx.��{חN��bY��X�_�T��oom�լ�*�F���-�>���u����눁+�t$�s��p��=4v��.v i7]32dm�X�n��i��sZ���z��>��-I�pwE ƛ�ㇼB �^��29w ��uy�aZ��`f����OįV�2�S�-���+f���`>���ҵ����'�ï<�Am��(7$o
B��A��J�_O=�Bس����`��f�'<  �;��3]��0��g-��e}(G_1.�Ԅۮ��Qz��s�~���^���e���VH;�I���5~N^Qˇ�LC#���{���LV�ꢕ~�*��"X��fR��KW�I�Օ��sc��R��F���#>��|����+JS�
���K䟽�%AG�u�nA(7���2�Ij0�W��y~���^9�"���(�G��'���$	��)#q^�����y�)���o�X�۳����^B�0����C� �=`HR��d�3d�� ��dPn� a�
^��]��|U���Z��ap���BM�%�=ZB���wTV:��xu�Ҍn�V<�>���U��3��F/��S�m��Mp.�P#�O�J��4ArZ��Ҹ2U�)+w�y���s����J�|Ӭb���m��т.�G��I�j��87;��s0�A��&�&ڸ��nX��+gx�>}
�<{�Zє���FƊp�?\����
J �.�8B�O(d��� ��r��O�AIƴ.K\��SRB�s5�wS(SA
u8�� ��O���^gq>�d ��Y<�?��h*�¦��86�f��{�w#�˴�F�\��������H�L��*A!�F�>8mPk�\���@���ߟ.�HT="��k��R�W�7��~���\ޕ	,��+D�_ L	Ew���g�� ?4b��Um���ȧn��H���-�,�!���8I6f��:���'��I�x'	͜[jju�y"���"�W�ȵd���ɀ�6��1,�OK�����l:Í>�NA��S��`B[�.��9'�#(�.���bn�$�q���Ç�dX��&�3
�Z��D*;�����И��$Qx��d�a�!.��DN�Rd�p;ġb�cE�efs��F��V�[��4��P��a�b��R���w�L��:�ҁǱC޻�--�y*�+��º�>d�u�����}��`Uplr
n<+ރ��r8�H_��g�p��L�����"�U�া?6�4�=�G���D��!��~af)��>}2.�%P� �](���u����D�ٜ�BHօ:V��]�&t0s�)|k��j�t��s�Gl�lBv���Ԡ�Z3?���U�Z`*H>��o�,�Z`x��|�K&k��~���y��K�-��y�����`��e�"���# �\X*���44�RY����3Y�v+�㱱2���:��)�j���O���=��"�E�j"V2NE��M�R�8��s2����`B�r��7�� ��*���V�H}Ik@x�b�n���y��$����[�e`?k�U<���HO��/7������cb�8�){��G}9�'�{����iEo)WׇM��oM$�W�+����ې4V�h�u�P�+�Q%��q�O���,&W�Ϻ��Y�[#MU7���������JlY�t()���¹,��LZT+�z�*���	0���L?�B�����f�ǉb��������.�>^��н���M+KE$��C�p��%3�\"._'�$cF{�����6)�6z�w�вם*&>y$����"$/H<Z��<�{�bB�Ŀ��)�ܧO���A� xʊf�!*�XI}���mQ��f$Lc�ƒ!=J;E��d�u�^<�#��#�,�P����L�o.��C��{�M)h`*�,��:���-Ȝ��!^�%�Ykd/{7��dP�,f=C�
i��Q؂�*��vm��^Goѯ���h�LЬ�`\`,X��}E��+����U��եyz���v�U�z�T���|��NCKԋ���@gö���M�J�8��p�狽{U�����
����fXv�]���O����{���%��KU,+�(���`#q���L��<���|��z	W=�
�'�ppP����̉2�)���dy�s�5Y��ī�ԹI�[:�|e�uhN	z�a����b'��y�"�R5�t�2��Q�1m�!�׽������N|X!�v��VE6�+��I���z!�-䋭蒂=x�mj���88���/`V����%Bn��
x55;�)�ď70����
p!�؉мj��H������^�?����b-�3���5dD�f}f�L,�~ �f[�S���ʿG*x!�s]=���ߔ�2gk&vj �܈��f�r�l�h|�m�1H"�#h.�EOC�g��l-�+�4�-]�
���;0���]�'�.��I�\��Q�i���ݏ<B�+_'��U�ҝ��u�y_.�@����|����(i���O�&&�d��ȁ
ۀ�2]K����,�?�*�C6U�AFu+O�-��"�� ��9���Z��k0!�+���~�dS1��c����R�rN>2�;�5���.v�J��u4O�$��7\Jyd �d� �^|\G���zp�����`���Û5A�*�XPA<�Wg)3 4�k��o���īB��/���BV ��q�n�3�Қh6<��!n�Yj��G
��2`,V�Q��x�C ��a��M����r��B���&س� '�OvFm�����%K�����ݰ�LSh�SCzGYl���FU
x8���S���͔ #,r����;<T��E�,���#��i��s��E�p�m2r��A�?�F��n�rKz�t�@r����kTq�cRv���c-��V
B�r��lMj8|�]YGI�`��g��Ҋ����D�����[���L]x�����%�DJw�8�H�'EK���U7���z����큿$�0��o���ƙ���;�@#/�4Q�,�k$���
�.R��S3b�?�Ê��w�!�w�W9!�ѥSm�]2�<��Y����DA�0]�f�j1��s]6�)xv�|��E�}���F�U~R7$~��֨
�s�ן��� ]>���ۖ���� V쫓���o���Q�I_ubj�����k�V�
�F=-Y6�V1�����9a5ʃӑ�'s����Xd�~5�5m�ϻ���o�[�/J*���\��lf�uF}��:>{�:Lм!u���N�a�$O�$�2�!|ڣx<hV.��UҤU���_�2��Apz�w�����W�����1����<Ή,�����"����95eEIP���(ro�gi�8q`S&��⵭�1�9���?�g[W�r]n1u9�� ����{$���C](0q�7�2�W'.(�%���ܷI�f�����9�Y��a�\�IZY}�csDMC��������X������Y7WX SeQŜ���0�[w�%������n�.8;f�ȍ��q'G?�Y��f|o_����l��PO�	���K��Ix�(��>���#��<aA��(- a�H���f��������8�	��
Dz�|J4T��mI��J��զ�(|R6�E��j�+ϕ7<f��j/s
O��#*�	s˥z� |�����_�����]=�-7Ǹ��M�C�����UN�5�l�S�,�9Z��Ww��n�VMάTk8T����p�B��蠙B��U�T�{�JJ#O��0R����{��#��#J3�t���>��s�G3�w_L�G���x+�w!�?`b�B��`��>��!��Xl�C�K�Y�V�BS4q���xS�6R�	�Q7`M
��c��m���^7�-w��-�ƧP����uC�r�<}�}G�'!S�J�جs�vp�+��Z�Y�l��(R`.?��YV���=�&g�K�8,C��J��^�u�lY�1��J����y�㘜��յ�}����C��t�c�$ڛ�5V���Ѽ�R�c��I^>��|�@��1���n|Cs�ơ�m��RJ��Y�V�ï1 hY�و�V55�ZXTl�[Q��r��B�xޑ��"i2�
��X�2N��EbB�um��r�4/�_�#i����V7�ȭ83�Ld �8w��o�j�[ˑ-����v�>M�X�,��pwE��)IzL�$����2|���+Nl��A�=T�
�H4z���t�'���SF�ܘ�2�
j���X�����5�i���������8:���	��׈�_E�׼018�$7���0��$���d³]g�͟���x�l��)D�S����H�}���V�:
��/7*��7�ؼ�m�0
��_�ZJ��p�-V�� ��"#�ja@�r��W��g¦��J�,�~�7pbM|?pgV!D��WJ��v�v7����֠�m���]k�_Tm��8u�"�t|rN$#���(�2:L�|Dq�*�/#�ln1��5>cE���Z6��m"4k�i�~��/H�|d��A��h3����?D�%B�O������?I��Z'��xEҞF+�b��H����>x����u��� ���x��¥�V۞ꑉ�ը�L�K��I^]1��~#��?�4K��OP���zŝrKBS*<W��쯖L��O�^#�ĺ-��h<�b� �B��֩�nn6��#u�_ V�EoXLya*���1 �x�2^+�*����Q��|�9��vi�,ʹH�s!��2