��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xMMh0n��f���X�h�ʨ���H�P�e�Iܷ �>Z{�hT������d�׽���EV�</�i0'�"�z^&Cn���+�$G�������L��>�'C,�H���M_@��E�D5z��#���,s��W��0�-�
�,�֟��;e�z�i�Q�Luy����V!4�}q-��)B�A��_�9�B�3��O��p�a��y6ۀ~����h��0hL��ɟ�B�Mپzds-��p��v�u>�ѿ�����b-���'AC҅f��!�����M�W���s-ӽ��:k�8C<J��o -��yv�N��F$��AE���j��9�fOR8%��/����i�ݧX�c�6�P����y�B��ce���̘U���'�q`��<��<ތ�3���=W�B�'��u�$/��K�4A�O���-!�f���(�0�����1��}Z�#c.��PxW|M��7����t®@@���P���Mh܅�#���"���_$�m���N�C���TH�N{�,���!8��#I���>��O�8WO��y{���k��!U�Q;b�d��?�#�0|���x& ���۸<��q<���<S�Gm�T	��%� x}�̭����e�X�#i�!�� ��V��$1��%�"����P9��s�Z� ��Bh����<�F�~7~S�u���B��קp�s��`Xk��2J���q��U(u	V�	#�nrb����L�%y&xZ���!�6fp}lzoQ��f��?0��-�BVǅ��b�����rC`���^]_s�c�ߙh�ث�W��q�g_�M��������H����>Y(�t����1h!ƾ���W�ޜg����X>
t�<���&�Q��6�\�煭�c��i:�}�*�8�-������Q��~	U�9�R>��2���c�+G��}{��h3z��j���jb��������7�d7y0M"�[j��_�,������c׮׎l�5�:�|Y��� ��g�t��դo��7|���"5T.�J�:�AA�cP��k�4�(]��$�r?�T1h��-=�(5��QQ�	�ʇ��,26g��m0����[���ag�e�qo��A�H,O���m�c��rE�t�ʹ��$~�.�-(Ja�C�����.m���
Y:53�����)�o��%t��D�i"�T#�G�l�E%rsv���n��&���#�c{��X�~ބ:���L3Ǿo�D�l���W�.Ҿ" �B��`�[�e��%�Ac]���2�2��X�되�i��P����|Z����g�����A�T2�b�M���7p���YFA�\;Q$���/I����'�C�Ur��Ђ,P��KTbYP%���J���(��e�MJ�4�6t}]t��x�ׁQW�w�m/Ku$����@�ۂ�G����sM-��au�r$!򷒳W����0?�4-8�T��%IT��!���k���ӓ�rH��U�ƥ���/�
mP��s�����{�S�:d�Iz�$j\���u�����$��2���p�a��QMsO�v�l��cVۣ�'�yBK&�7���~[�I>~����+����|&}D�mtV��?�P���?���p=і���{���B�qd�D���-��S����f0�4��bDP������(��s�!�5�O_1%eq5E��G�@˗m\]t���..��姴l�[S/�� �5�}X��(�h����%�i)��b�'x�K8�� {��^��(��)Y8�P�;�a/�M��/��ӃE�j�q��H�����~�<�7.�ZAq~
?����z�w�cP��|�W�O�Oi`�st�����3&L��Ӹ2�w��@+�زD'oD�p
��o%�������B�\b����?cp��5�������e�5�p�� O�d'�X��R~k/-�˅���^)�2�͑�X�y>FQ3�oa�.d���da>����'������,�3��Oz)[3���:P�M�f@6q�!P|�`�aa!�>�K)�x������G�J��!��~�;f6d� �{���;��#�$܎A%Ð���]<���}��P����u2�=5p/@��`���3t��>P�K=K�����D��n.���H����)Qa�%E��h$�3�ҽlLIRmR#��km,�a:��4�P���@�)̡x��4�0l�P�� �;,s*.�$9]8��轻;fa�!�w��|�?��{��`B���脎Ւ�p!s�o��l5@�x*Q:�	�ܧ;�4ΗĜ+����j�Z��d�b�'�T/�Y���d�C^�A���S�¢U�!s|Y���	(dW�lͿ�Cm��`!�m��6�5x�;��!C�-�Hz���&�nP�eȑ�e�' �����\!��.�<��p�U�B�cFIī%]��wim\E���a����a^7Z��XQ3�-C^e� nj��'����d�|���z��d��;ED��R4>�p��m������z@Y#�=���0�������T�����h{�AHI���C�ُ�����X_u��s��f4������-�Hjt]3	�_�O�D���	��v�9��j�9C��)o�F䠼�,l�3T�~�,J�2Q�0[@��_B�PwǅY���]�up(3H
qӕ��g���ƣׇ��B!Po,�����1�2L�Va
��W�l��=(!�a�=Y(`�sJ}�r֭n/N�ʒ	�Za��B��x�?n��
�^U�M�ӯi�䪑J����͖�n��-$I�ϫƙ���էJi#��]�(�M�"��c����y��k�C�v�P���G���{�2�K?_�+��7���"�����!Y]:��٣���'�y��5����hTZ�b�F�[ʃ��˛²e�Z2���ƋB�鞱a�Y���M� -��lb)q��	�xl��	�]�*�ظ��k?��+YNr�(;~���Y n�JJ��;ր�vlY��<�`��J�n1�?�`���	�i�!�<Tq3��b��Un���f���K�]I�Ǿ4pFBfh0��Q��������6���߾�\U�U6.�pM��gh��.��2ט>c��L[L�����!O���f� y�'f��+��A>�F�G�2�P@��Bo���t��=��n�)����dc���^��s����'�sum���U*^�ͬP??�G�̘��Y�:R���>�I:#����4�����@�:�<lZ5{CG� �"�3	Gl��܋b��!�to$�� ��m�bd�p�;��$,xQIuը>{�=B���s�I0��1�|�U�<h��J�?2��a=l�Y�����a� �|���a*�]��VHy쩊�ņ!8�>������"/_j���)^cd<���oJS�uꇞ�P"��A݅�W2�� !ިA�"�t�I\S+V|5~�����=��ljuύN 5^ 6�6<�)�p�3��V^��V�,E�]E7� K����ϱ&�r_Y'T����)V�MJ�WӅ�aif�;}.�ڷ�S�{�w��6�b.-�<�0�L����1ƾ��[)���=#����Ꞌ��.}A�Y�A���M
:�
ƎOa��9���Q�E+�r�}m�w��imӦ����k�| �;�ê�I�e���|���N�nd����z�)5$iȮ!-����\ޡ��q#/�,��{'���-yy��W����&�~��u�x�_�+f)��I�D��dV:�	Hv�
�Ըn���J�v�kH&�\���8G�rnӄ۫U7�(ob���0�������B�P{�g2�t����nw�yÉ�/��2S�c�uT!u/.�����fG���O&� e��9���@��b��c-��=�C�#P�YE �	���0��Ⱦm��BIa�U�R��9D��U/�ov�μQ��V>a�νp���j?N�n��� oȖ9zY����b$k^h-�4���*��&��F
ȟ���+Y����`F�)`��H���jer�=�(�u8}7�_�Us�Lb,W"n�翺�w(���jH��WT��e����T�9׮��6 r��oX��g�߹��jiݽ/^���<���\��_�6W>[[t9�����\�F
���EW�����ur�U���D-K!���&^J{&��%g�y�M,~����*��g���BąC61��oE���I�֭Y���C��T%��%�I�.@!�ww�]P�W�$�9�* �U  ���E}
�Xes�bV�%�מ�`|md]�,�t.Db�򒫞 �_�`B������V%R2Sr�A)���MCk;2~�֐CJ��#�( qI��t�+eld�јCY�h-�x��1��W�ǜ��x�d�MV3?�����7�:�h��<lN�I���r�&���M�D�^(�-\2hT����:���iFc����\���Ks�̞���+7�[�6�)�YM!��+�z.�CJ*��X�/��sطoxR?��4�j����6���/�e$��|��o�&�އ��%B&@U�� G�t�pͅ�=3�t��%p&Rt��۳�-\O���+��°s����D�h���c���uX�c�^7�WPR��}!��B���\-H�<������2+a��4�2p�j��t���Jܿ^F�J�k� /���#g��,�i#�R�5a)�zК�$T#N�MC�(��&���f��$M���Wr(���pJ��l��N�����н'Y ��4�s�C�5W���q2|A�kU�U�Q�Т��?؎�?!����i}]�w<@)�-����tQ������&&1��y�H�^E���M��.��X��4��"�}��"ߓ�f����P�\)��M�������o�7�t0���&���N����L��Z'�T"D��m�nP��`u�8zS�h�%�@4p�����1\O��wc>����M�F.�n�A��'i�֕;~�?�ߛ�$�d4�.!��T�y$��0yh�6�}=k����k��*Pj1x�[(^�zB��$�z�h!/����&j3Fi�|L:9���校S� �=�+<W�tJX�J]���7r^x��]BNw�1��R�ZI�r
8� M�
�'���%\�����y��E�Ղ<�Ţ��A	o�Lc�It������VLy�Տ��F�?ϑ����c�4�9ȼ;nW2Z;s����	�y���*y5A},.Qz���Zqϣ���mr���B裕�.�1���r��j��ԭ�3J� ��Sǖi�m�R�'/fy�.����K��y��	��'�X��b��H�ҥ؏��T�6�?���݃�JpU�eUaD�l<�#Sj�P�W��cjF��V".���'������_�����K�:>�Z��Ok�A_|�K=#,��	�w�������D3~)�S��rpM�X翿;i�r	']�C����H�V�A��<6K�^�A�%����&p֛y�g`\��l`�d�����WO+���'���4��$�+Y�{<#�����B����������:z@�&��������;bZE��kV�Hy�\gM���k��]�'dcp1ՙ"����`F�?�8rK��VqmИDk��
��U�;��Tأ-���� "�-��,��0����=a�۝��n��A��8ӯa��>�V=�$K��1�,��Ґh�>��v�}�2�Xý��9�C�L|����b-����{g��M����2��Y|�g��QG,Ż?�lj�<}��+�٠x�h$�/�|#�j�>�������u>����C<�4�Z�R�Wb��Z����#y��B�8���j���8�%��\�A�pX���YD7[AT��V �Ԥaf�X/��D�ܰ�֚�D|�KZ���k[lB��~~�׆��-Q%�\:\�s�Zuo���5@�	�Y�pFzr��h�A��ѡ�P�mdtG�*��:p՛��P5j�du�#P5��A�(�t����,~ƞ+ә?�����F�㯢o�?� Qa45ҬW��:�i�ԣO���L�A�O|Q�5����ӄ���K�G�?�oV����{���y̍ނ<�j��T�f����__�Qz���� h�c+�bfY�l��c7"�+d��
�P]��q�C�0�n�J
1 �)`�s'�Z�!��[+�ޗ!OZ�@��m��~���L����-���s����Y����6��t.dIj5���W������xP₤^�Ě-�0m�_�(���*"X9���X&6tg���B��S�Y�d�[��^DE��s %{��D��s��1'�b1c�}� �����B�y��h�:�RO�mp�,���7�-00(W�и(�Y>q#������[7�C}%����s��85Jڋ��U����{���r lp��������]��Q�ƫ��!�<W3WNDV=�F�G�o� k��C�=��ڃWա'
e�Cr�\K��yo%���Jk�jo1(�_���rs��a����H��ό�5�u�����T��a�"�0��<���G�{X���z����0�<��(�+d���/���:��դ2�d�e`��m��������gr"�P�(9�Q���a�Mj��c����z�B�j����E�s���|-Z�DF��%�D��gO�шe։��a�� A~���3[&g`�OSp����`�c=5���M���m*�.N[��!1�X�/�֭U�.u�Z��V�L�?�:1r�ָ�C]�ŋ��
���{甃DYl�̑Us�:�5���ڴ����#��[`!
�=�<��N�!O�L1[��!�©9"�����:�8���M0�،|�K�V{YymRS���nM~N��ԿE;��������]�|!V(j�u��z���2dY�HR�e?�����y��(ߎ�uɓ�C��%��a �W[9���d��E��"�p\��N��Q��\�
�u��8�ա�s�	��c��!{}�����,BQn������z���c�襌&W�x 5��3'�(�P���ML4~����ȶ8���PP�Ǩ+@�˩bc�=�j}ءd	K��R��Ͱ��7\\�75g<*� g��߻�4�Xɕu�f?�pwu���.
��Z�L�m\��֝l^I����Ԗ�5�X)AW1t�8�7���'�S��R��ˀv̓����/��R�V���Q�>gg����/�>�DIU0#J��k�����d;�«���$V�KJ���(G�bu��W�S�>h�ۙ_��p�� �����GG�M�.�`�K��"���$��%GhE��N��w(ƁGiO���tQ��[+���i�Un�~R������}�7�̺1N�D�O�\Ջ�z�D>�\��-�P��O����)���搶���:�y�'R}���ʙSv�8�k/����IZ��by�>���K�#�u��`�y�q~�jeD�R����f�����B�!�.�ɷ�#��ɞ��x�t�(�2�(�o�#�3��hW{��<MN�5.X�)D%�e4�SA�|Za���4��Qtf�����r���\��(�W�A�ld�����u�DA�=� �^��6t��7˰�2��<��.'���d�/R�U�Eb�f�lÒt4r����0�;$��r�L)'ۤ&��R��jI$ʷ���hL<�ԡ e ٧�<�Խ ���#�{Z&�2� ��YKɁ�^b�����V�yݣ9��=G�V��������Wt�֏�l��M��O�@	���\go.V�ہ�.n ���z�����[����׹�?P����~Y���k��ݮ�V����=�>����V��@��yɟ�=Ѭ����R3,�6n�� �M/��ʷ��^����wo�uƸ=SN��u��k����O<
o��Д��%
Xj/=���T)�~Ms;��V?l?QO����Z5f�^mZ�`Jus��s��I�E��f��\�v(d)����o��#�����֥��'Ω�hfH�Q�8���@��l�ݲ2��I)m/d�4F翚5� �,��3MY����S��4m_�k\ޞ�oQ0]n�^��+~�ϼ�Jqa�p�e�;��e��J��>�M 6q�*x�iݲ	9��HThڣ��ё����g���h�If!i�*V�4!��%2��VJ~o�� ����C����g����[�/��F5�z����	�pH��q��oݾ�
.T�-�kԔ�c�:cǺ�76�pP`�rB%��E�o�:�^�Sl���V�g��6���v�`�17�.g�p}�7���-_7�Np_���U��H���6�$�;���ZAiC~���������D�ɘ3'p2�?3�يYrp��_?N�a��`��;���.��P�Br�M��zO���r�Bm��[F��h�g @�]y���0]��m�F�*�O��L?���ezёE5���^n��*��9��I��Mk�mۚ����@C"Azj�������5��6-ܡ��O&�i��T!}IM��ڂ�������ow����F-&�y-�-ۉj�!J(���Dـ�0/sx����VTg4|㞊�`U��@H�'aF��O|ڦw�l�zz���ö��q?ЉH����*�(H���_�*�����\��qz���-���ǹ&s��<Z�X�����p�W�.cQ�V�*���I�������ӽ_b���|�9���p��ʲ��95{#��I��342;�M ���%��J�ú�A������rG�4���WJ�i9��ėQi��]��%��>���7��{A��,&�x:5X`"�FVr|����4��|� }��=l�h4	�Ui�V����X�{p�:�:ۨ��~TЦ��<�љJ���0҅�$��5,�\O�Y��o�dE�*=E���u��(#�S�4�s^�eo9Jy_[w�+)d�@�\��&���\�a������L�Xر��4��1�5S͌@,�0) �y�kۙذE�=���C�^�KQ���4/��,P�	���o�2�.��D(�E"1f��	�[$,gy���C1uM�s�<��	M݆�Mܕx�1G���