��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨס�>�6a��S]/�k�q�&�S,L�Q�1�=wޫ�h��]�	��&�ZW�-|)C���v��,�R��D��-mU�$&=v4
Hk�C8�6(z���+�AĶ.���u�u���F��_k����`�~"
���h�$��͐Oz�O��dj0�%�)}q���U�ni�1C���<�4G��~u����E���F�Oz9+-y�����Ș��R4�c��W��G��&�NS���a�W��t �Y�����j
��x'����N���y����=�����|�%�.aݫ��%��S�cD�cd�<7�f-���Z��0�Ǡg�:�&��ys��C��Y)�嬼\s�aC��yt��D�������4�L�ޭXT��
�P'/��f��������·V��QG.8Ͷ��	�̬2gi<mY̟���xQ"�0�K�ĩ*��Аٍ�D�	�kDvq�����᭭}S#��B�nac�ǃ&`�+QWv�e����هP�;�rW@���8�=h.��4,��XP�N�)��#n@�\���B��^��AaD<���%'�_,��WH���5c,�α�Bv��
���4m�.T����<�=��h��X���z��A2�\�;��`�P�9`�����6?��� ୳-G�e3��B~��t�<��EZ>n��w#�ńRv&���6ޜ}�pJ)U &��ϱ_^z���yx��*>K��G����l�y���䱆�(w��5�Rͬ�c�C6��8�5 >r���*^��5���å�g�P8�)���V-3:X��W��(�m��'-Q��q������:k�4�gʃ�=_6[%��D��_��ݹ��`V1��#�eǨ����D��� �JZ(�U?�)E���	J��J)�Cl�>`R:?�M���;��x0��吣o�䅨���}�Uʴ� u&}ȩ@���4o�#{}51A���,2�@	��b8AE�\�ѕ|DR�_����� �����WpQ�(���gc]8�|������-⶯S��иU�yp3%�$$d��5!n�V-�"H��M�u4v���'�9�)s���́SN��������P��g��+�$�$���|V��j͚�{"�"�H&2"[^M��-��I��	%�LnŜ��//luFpݠ����d�����[�u��ʌ��$�S��Ť��B��5�̄j�]4��9#��|�_���l��;~'�>�8����N���K����}5  ��#�ݐW#���i����:�N���_��#A�Ůe����2�O3K�_;' �UN@�G��/{$�N��?�3���pA$U cU�L�/��ê�p��^!��c��B'mQ!�Žy�U)�p�_3YKA����Q;m֭��XG2f4�ӥC�o���Ft��?'F�}F���*��l˘>��f�%��$��^���R�lK�c|lWմ�����Ч?ә=�C�r��q,���|E_��96�ئ��&�<v�ވ�/C��"O�921�P��=��ɰ6Ś8�VY�-��h��x4����ٝ����Ѳ�0�,]��#u�!��/��~���`(��[rh��������^���7��BN��!��2V��^BҠ��_o��BFj�[����z�w� 5��1�Qx1^z$¥�����m�N�MӰ׻^�KR�!wG�VG��'D���	u��	E���i�#��C����S^C�܇̼�'�q�Z1Q�"�OX]V,Hl�A��m�������Y�E�U����/�1f%d9"s l28
����=}����a�Y���G��ik�Q`���O���4i[H�и������Ǻ'N��3�|q�i����dY�f~u�z�t��//��ew7��JiN y�F<l3 ��"�THU�jV	j�����_{���׊B����q)Hi�Y�4����<���cb�k�)�`W��o6�b��$&/�o�^���Qg��F�a..XG4�h�5�����D\�Mj�`�����8eٯT��Ke?p�V��3d����c��O5!`�d���%b��Y�YÂ ��t���h���&�Xw����>d�w�ئ�����b�;nLXd`΢� Q1.�Ȏ)6����⯅�m�bj�6�1�05ڬ�8�dmܳ�L�ӼW�3 ��NP�13]��+zAY�8�UV�n"��~�^<��k�1�*����-�����2�YN«�)j��
��E��&8�.�J@Xn�ߓ���pV�}7_&ő�-��i��R�V|�Gl�X�W���M_�|�ްc\�0Z|#at�-{���]-}�i����Y�d��\Ƅv�{r�Β���1�7�l�6�#�{4��#6��K��s������K[!�!�&�vhRڈ'��DH�RF:�ҎϏ\���㵍����M�A�+�4�8C¤8�'�1��aNe��
����o�����(D����~5 r���淝m��	rq�%�,[D�����TX���B`'��֥�5��XU��{�d�\6�W]y�%f�t]�Hb}k�"�U�߈TM�F�A�;.(
e(��k��2q쌤���Q���]���xE��ݩ #�&��%a�u$��c!����#}G"�@�x�P���`T��dl����v�x�N�˕�Z�%�O��(aj��޺�?}���th�y~�s����������e�Kp(�I�蚊���4I��8g�7�M��ЂYᡜ'��^g[�Ws$V�<%g&$>r8_[��}��O�3l�g6Xݼ��#e�2�}�P��i.��u�R��9r�ܙ���Ӱxri7iEZ�%�m'܋�߭3BD�<�(�1`!K���9�uC��1�u)(�^�V�2g�a6͌�ĥ�ZbfgO�j����v����i"Ȇ*�6�O� �g��9������N�^/5�Kv�����zG6�O��yA���j+����8�3lAm���ԧ������j�p��#Gcp:�? X���p
{��)����sԿ3��Ro�y|���m��Z�2����"tF<>o�e-[ S�:6	��k����-(�J�*֙7E8>�^���dN�O)#rU�%$�/�u�q��ĺF�gʚ�!�H1�ɍ�|��G�$ˢ�P9�����M&������^�E�ʺˢG����s$�>��Z��%О���b�ȖoZ�۩)���2Ս�����)���~S�[���� ���rC�g.U�%O�h��wx�,���� ,$�3%Y�B��Hsl���c�^Q����_�d9l�>o��~��(R	�߈�)�5ې�:��z�5-<.�$xwF8�x<����>��ڋ�HV�w���ߓȨ�U�}d_�r{"HD���S����M���9�Rw�����z$FS��x�d��^F�w(J�x:x��&a�ۀ���R|e�7�ׯ��B�;�y�˿�!������!����aj��@ç�i����k.)�e-��۪#��	�Т�Z�S|�>��cW�NA�j�Ϋ��rSj�b�9elݴ�Z�{��"���t����؍lv�M_��.o�����s�^�==�'����A[eP����8�DeŤ����t�F�7g�$d �yE-54��E��.�{SX�l��=�p�c��OZ@��}��בu�뗍=Jl�}/�KM�>�^��QIb��4`P�z�QI��P�T����2��%�M�#3&��b�L�'=�OV�3V-k+[.�X�E��,��`���.d'��|JQ�e~*_�L	��7,ʬT��[�������'E6f&�Pķ�y��r8�Ԉ)���WA�.��.��,�~ف��]��Բ��\Vhy�C�nGu�F�!U�)w٢�[:5A��w ��nڊ��.�Gg>9��]�8�ف�u5i�yI1���O*-��$��^[|).:V���(���h��Zq$@}[���\sp�܆Ϛw�J�~R���;�F^]��8�����)4M���m�S���d�4#�&���ҙ��a��	F8BԬLuĥ���PkR��ݭ}��<?��I���QBR�����n��cY��6@�!�{"�U$������,gM�T��c/���'����đn��ܳ
�{Y�����zi�et��5Q|�mfB��!��p��R�35i���&�BD�b'��qo��SZ">�_?f�e�j:�7!�FeJ�!3L��x沢�ĹX�/�-f�þJN�靌��L�����>� 09Ғ�	fU�;N�Y�!�0?����~ˊ�'�E���֩_l�i���dnD��`�ev��L����.N��n��7~�����P�X�R-T��s)��i���u��Kn�:�+�@Ȕ#�:���3W���%�i�y�.١&)���A�ȜҳNʐ�.8z�X�'f@�<�`�x��u!U��ȶ<JC�l��7����#����瓑:�˝6)^���<ŀ�Q��R�� ����%[��K)۟6�M�l�̥�^a��9�J��ª�FƎ�4-���mR�/s�����sw���{6�����J'F�p�����ٓ\ҏ�ɪ�rDp�^��,��z�HI.�7��=%��$��I�$$+|�g���	�٪�.���g(��L�'�Qx7L���A�PXyRQ��-�.m��v��
��X�S���J��^�f8s���+a�ʾ�tV�c�!`7+NϿ�=B��%dl�~:f�k]F�Z�s.P��
�������������;�S�h�����{ʵ*��(�y������,�Igх�	��*J�A�t:.��[�����z.-���&>p2�[[Ւ��\},EIr�&pN�v̟d0���1<ʇ���3�K�ҽ|B&l�*Z����)V~�Â{Ʒ�mF/�.�d�C� g��a����o���`�p����t�L��܆�/=Qv�}^EJ�6ġG�7f�h#f��]rˡ�+��Zx�Z}#��B�M����
%?�$��&�y���I��T��,���G����?�yA��]��4��-�0�)/�q,�)�U���p2�	�����gWT�=Dp���P���0
Mقxݐb�����y�f��O��:��+�������Bɳ����Op��֞X�e�0�X�{�_��`�1��yF J|��k�t h�?��ߘ�)��D:'�?��󠨘i���#�p��P1�4S��H���a���X�����Km�C2���wt���Kx\��ݠ�D�qA��"��x�:�