��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,V����i�E�?=���g~��h��Bz�D�*�䥢8'����=M8����?:?�-6i�\������oyk�Ã�`�uߢ�U�l6���<9ِ�	;���M�x֏]��Z�](�dN��G#��iWDC8 @L� ��l�4+�<Еp^Pga�>��X��ML����q_4H%�g�m�'�f3��̰�ɡ �OU�2H�M �̬l!}�gXF�N�@�t&�����i�$���3M?�i���(X膀Q��L&� (6]Қ$�{��qɎ��	#h��ފ�$��&oe�W W�p�5��gI���c�u?���B�؎��E�G9��|p���u�`��E筝�W�c�o�QIl�hAp�d��:n�Y�ڞ�������h�&ئ%�����q��ٞ9m
�F����nY�<9�5:�0B`�Glc�DC���Ҝ����g\C8��IgL�J��e�d�-Y�M���\�.�����ϸܮiV�%cLߐW��#I�O�������w���+QޱAV@>�G�^s0��I�[� �ǿ4FhA*e�ͥq��EҌ�~��,7���OMm	��n����Ьjy����D�5�<��	k7tP/�����uZ
Q+]� � Ͳ�����qHi��F��׼?@成�1X{�(t@0v���we����hN6l�%�? -��Ax�l��Ҹ��5� ��MeKXK�~��oҨ����W���㋎2TЧk��;�"n�2��L���4v�Hy#�ZD���j`?��(&����`��_^��w��y���C}�(x��,��G��'�@ �I������ݎ�(FŘ9}1����c��C�6�2���v̖	�J�a^lɆ��ǚސH �p*�n[���]���E�.��'���_�Xj̽=g����]��5s�#�ў��޽Q
������^��6t�"�w�P !V;�� Bឞd�s��Rc���߮���j�,	5&�m�6�M�u��+B���xӈ?C�W�q\gP�}?׊i��kΣ
$x��/��������8���nihje��;_�~�A�!R����e��lhrzGn�f���d0����6s�GW0�0�$?�9��b�7:���T	oI��{eoʘd�R�|St<�#3H�.��f����y�Zl� �s��a�M�H�t���٨,�0�<��m�(�z�*,�]c`;H�Cˎj�u�>7T!�\"�d���K��p�_��b�w�·�GlSKf�񥋽j5ߠ(�����f�c�o5)ݿ~%���P}Z}����i+f��y3� ����&loj����Z���� �t��zA4�q�2$�=(u1�8���fϴD����� s�����:3�����>'�n�&3���,�-�Kj�9�&�D���"��QS�]��>wZ���햪s�΃�T���{ȧm��B��&+6P�|����� b���;,������Q���2}~"	:�LX�g�)�����Hp��W�_��'R�L�� �]�RhE������%�Gh�G d0�8�k�KM����1����@^/6[OP��r�n�^��q^���{�l�/F���%�%vz���
��8��R�eE<>xh|
ۡߧ�����%5wYwS."7Mpd:�6���y>���!Er��輓�r�s���46,�XZ�K��M�ڄ�� ���s3Ot���0'f�-P���8��h���g�ݝR�`Q��8�֬CW�r�5��i��b*�K vK�Bcǥ�������9�{�G�8oo����'y��� ;7ԧ��S��X��� ����J�����v��\S��G$b.���G��d.� ԏwr�8��C�PQ"L�$��	?�SE��E�J
ڻ/1�l���L݊�_U�S�D&zخ׭����E~S8��b��'��T���I)�3y���s&����E��"�9���k�3p��_�*`"��ӧ+`dC�_ޭ�		���^�}j�'��F7�z��
�=�R��&]~�uƘ�6�^��Aީľ�liH��/�b��C�7.��@9>����KI�w~Pns���z�R��-�pm�؍k �Ye�g����lnOF����"N�f����L�R�'bdsT�t�<������&%R��=�o�gr���H�nlm�uJ0��:��ءu;"/ݟ�_�`�0��g!�.~�;�VZ1��(�{�$�є�5��Ɔ2lTx�����N��H�
�/N¥�w`17�ٜ�@�W�amޜxV�H]+''b��hf���v�m�¯�����?��Y2C�e�v�+��j�������6(�z7E�~q����7��5���G��"@�������$H���M��t�q����Y�O��ıU�0[� �����w
6	Ac�PK����5�	\�(M������1�M)���3���ҩD�\�X܃�R��8��h~h_қvG'���<[q./�^FZ�{t��}�T捭��8���N�#U�b������3P���j�ՠ�