��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\�#��t"�9h��=�4�n��͇���@�1��(�ifl���H9���N"�-IB�~����Kj��(p4� 3Y�2R����y�x��}��5��"W\�شA�v�;��P�F�_���������~H�?��B��O������Np	�э!�w��	�h�A��:]uC���S�%I�ڣ��z���=��2ƾ�*�	j-k�/0�w=M�?�<��jT+�z0�إVf�.#����\Ԝ�78�s����М�,S�ΧT9��vz��"
T&1����~s,h�(�o�d�֨i���є������G�I� ��`9�Tx�&�?�z�)��6@�w�� �e~�/��q۶����^�F5 ���i池ݳt��Z�u�rI2�;L�De*f�,)���!`�z� ���2��J�u#T��>Z��8�o��CF�5�~)��q�wX��:-NxX�0��^h@��Q�J���S�,�n99QS����;X�֨���s�4��TmCa�=v��`Z�*�7�=7F�t9�\�d�@����?i ��p�{�Oi넌��9�+������Qr��ǭ�v�� {�O���f}���H��H'S;;���)��фoG�GȄ�S_a�1!����O@%+!mcP�|��J�#���!r'����P�G�)ݬ����:|l�"��b7~▏�OѢ�7l�����������[��@�ԕ�3'��D�f��^zV]�#=�1� �N�w!	�8)��zn��,���P7���*Sŝ�}��9�%��)��������#V0hB$�Cf�*�h�m��w��V B/�*��͓O��z�U.��è<g�d��m�S��������G'M>��q�+0������5��Ջsڹj�[Iǚ1=�6��t����4.B��n��G���ф��cǵ�E�D]hv]���M�����pj� ��1�xa��|�qe�.@��������]!kl臤�GUa��<1����������������06��xi�)�	y�b����U帋�k��e�^7v�����ޣ�6a+�;	"�Z��ݥȻ/�)<y�n�e�mV���쪄�?���L��=�=O�h"$�����qhQ��
q6��V����YE|ݍd�'�а`'�JAf�V��d
er�u;R�ܗ�pz������dZK05��G�A�ڮ'I��O�/��j��郉� ���`d�y��@D1Ԛ�I�J����3}5��ۚ�_��c��,n]�;�;�t�K����jї�+���S���h��SF�)뾜�,B5/O�H���"e���@�] G( ������Ġv,��k6���9R :ï+�C��/.%�CC�EZ��7�.���&���"?�<����u'���9�g�հK���Y�,ak�JLH�1Ї�_�^&5����.�������~�)��J�0�����3W6� :d���k!7$=��WI�0S����a$(Yl�����Ll�Y�Q�����1b�$*~F�ǎ/[�C����Sm���x���ݦ �Q�6Z:�E� XR��i���!e��1;$o��*�Qp�$�y�l�<ŧ�9���NIö���`��K����}�"r�D�����R�������y2�����s� ��#�%Q +���l@�1|'���[�q�gCuYS�Rq�bߤ�$�9��*����䞃�Q\�Q�g�Ͷo��)r2�\UIc������d}����y9�y�)�'���weO#'!�Y�]~��N%���{�C���}�`s��S�k}�\cL�U�Ğ~���\�/S]z�}�:/�ī}׶��Y���{���T���m�Y{�o�YP��%�>w-��F���ّF������xN*+��]��*�_*�e�mπ~�g���i��,B\��i��FH�����c�&�E������FIk,x�2�%���{��!��Ou�*����@)h��h��AsMm�H͏M;Hi�s���c���|�����n.6�3m���H�A ����U��ԇ3a��Ӡq2x�Ó.Tg��Z-q���g�wX2��W��{�S$Y�MD�b�F�?�"���eqEZ�j���n�C$�����ppOtF���dN�,����9��x/��N ���$muo�4��)���v��s�%.�0�&�P���G@��ĥ�<��9[;&������[{��R�M���4~ә{
��z�Q��Wİo��i�o�Z�;�}��Fݓ�_���`����_l�N/�*��� �u�R[�:�m}��:�p�;�"w��M9��.�S��u�*x(Rr2�u�y�$c�zhq��`x���0U�7R���z�ËyC�m��0L3��%QT�3��[Q���?�~��`��ތ7!��ӽ�,X�x_.G�C���o��ȏ$8�l�A��q��[s�1.R�����!�G����@P~�w�s^�dDa�VS��m����g`\����}J��"��V.�ꥩ��y�|�`UW@�l1#��>S��8�Q�&���tN�e:_����=Moc/����:͐���VF
��(�. ��"�VX>���ȱZ��s鸿�@C<��-4A0.e�`�ԉވ؂���F��1�Jz(msR2ķKM�4�T;� �#�x�Z) ��^ݐ�/G%p{�#ɀ������p@�ᰯ��oa;j�KK�
��W��Q�A.
�~��,ISxX�*��b�Gq��n�Jր�mO|�Ȣ8r0<�P�H�*CU�|Q7����#��P;u�0N6�6���0�{��/�muV�xʈ�>�}�T��b��X��8��	���~�Sc ��L �����t�����-G��f
}J��#��I�7��dB@�Q!mƥ�
Q~��OX��w�{͛ԲB�V"���!�?�ِ2�gϜ[�Kxn0�>	&i��ؓs��*ډ��z_���`?���ܚ�y�.���BC �|%�B�/d���i8B ӓ��17�#J�' �elb^��9�:�Df��rϗ���BV����ZA`NDh!nW����;2�!��ͩO�8�fke&��a�m������ ��س��F�����	vlp��(���,�,�����r���Yve��6U����8Lŧ3�	�4�b,z�g�=�~�wT0��l�)#����K����3b�U�su[X��Kn��˝`U*�o�5%Jf����$E֎���%27��v��~��=ռ3����vGvK=�]�[���yK>ܲ�K�j��Y~����B[��~��� �P
4�%᭕�LgΝ=3%�V�:R]���Β�"�ɤ��}F��.$X�~����H���^�z+� �S�/:`e��\S �Nϊ���P��$���u �(�/���ǔ� ���ޥ��p�v��7ȃ5ڢ��G�K�3�A�+�ir��_���&�:k�C�o�)jJ&��}V*�����ɝ���4�L>�o��R��Uj��dٽŚ\�s��]���~�|7 *M:��}�*�O&���*s�~�!ߖaCNLr��Wۢ><�p���r���I������%�d*`�	��߸�+M�����ҥi���xd�8$��gYѽ�7ݠe�
B�+�]N�?T�������6�v�^[�9�>���d��"�_$��ʺ�?�˃EB�ZH̢�b�\�F��BW���Ә�
/I��#����S��j�&�$nE�qj����;�rkP�T������L�O��J�����
��m�櫚e�J��{�|�Bq��v��%�"�	\=Q̖��O�Ʌe�gj�5���>M���ͭ��Ўu�!g����pD���Z�b�C���vn�|����l\�W�-���^��z~�=U��fP��`Cϸ��(���8�K��ź�j�C��I���ŅrF�b�6������tU��g�Uu6�����+���{��Wp�\L���I����b����o_�ܭH��bT���70����|A�>!��}`[��3�my1ߧ���;;#!P�r�j�.�� �ƣ��4�P�"�Qx��/�|��s*z��iwF)� ]�M���������U,*�L<M6e>~�	�d��,��M���ɡ�5c�
૨ƾ������L`9��+)�2]-V�*�S�*"{G"���Kp�x�dM��AdyH���Ce@���G���L���cY�hI��8��d����DDi�8�++�<��p���L�Ѓ!�$�nK�t0U��!T�U9f�@}��y��*b��r)g��li㏁��l`�m�8�#�>&c/F^a�0�dP�Kd���pN��F;�'�@��Yy����B�_fL�Ų��H��/Gu~ƾ�L~��n=�H�&���oe�����w=��e�ĺ��v�`E���|��}a����ݑ��}����֬@!#�~�m�X��
���2A�����S�Ӥcs1��.՛S�
;w$���XLg�f�׻�)����&�F^�J��#m�[g�:]t�K�i'��}R)�-� �K����Z^ѧ�ʶ�}膊`�Zl��ק���u���jj��H�d�k�'%�>{�V��'d��A��7��<[�Nz-R��
����護J�Q�ԗ��Hc���	/6��t�Q)�%�$ǖU�x;+�F�w��%F�N��$�/���.eqe�9T>�H,2l���mkhn�rp�n"�-6g�
�9�%����������v���=����8���`����?6�$׻2�qy#~9ZvT�?6��"�\I){��A�i�v3b_��N��F`?GO-08������� �jv��jr5�㵟��6SJ'}����8�K�05gh&��>޽��dxU��R�a2�!�5�P�������w��ܶ�Z�+хDLGD��!�t���x���8�n�,�@u.�V>�A�8}-����"	�0D����v&,P�憍h�A��ń�1��T�=�}��{Ld��jdǳ����jE��t�8 ����S�\_-W�o��E����=l`�Ǫ'�G.=!��Ulq6� �E��g������Τ�� L�l�9��A����׆�HO�~�{�!��V-K���7aA��W!��q僊��p���r#s��|��`
������ѽ�z��æ��g��b���Ļ�RV��+���w���