// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:34 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V3gr7nLD9QOCKR6bvEPnhATwdRTBarT0CnfpwcwxI0AjcBbn1eQtbs0rYfg0WbXR
9vexXXX8ESdcZgxrqf36hse4EmKtJMGPnTDUFFPqYU1aZR7NS1/lM4Z1vcgcud7v
1uIuQhzouHLz6soYDjQv3sCU++kaP34Jv6x50RyefXM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1584)
Lrglr40UW56YuzIAyCDZoSkd1kSrUwYU4l5CCPqMr9rB1qr9ERvoQoHz8Q48jzGx
5pBWGbdl7OkE/AaZWqiRpg12FzUVRCcOhM7Zyn7XfYvYcmj+e4z6EK6/Wwh63O2l
+yM7F9ALMYTdTBRxRVKiOK8lvlqPi3hQStQZKs3wuYuTnzZfM5m2WXtd/ThmggCS
arqmbfmAIFQ01fANWYaCPyElzi+EwQmd5+SCGUq4JLtOqVKpUkVWHKumkVXkmbaM
GsqrmC7jde8lm3Gc4+T+pZOkg93uKg+9vPA3ISuadxa+HuHEUXlGCCxu/wq79xi8
G90Mh040df6vLRoyokx1TA5sLLmVeJpU44J4y2YoFjROpLVM0AwB7gdY2uWu5bJL
Bn8mNhzzhuRmnLojzsLD94uONdR/mpAXYCaPHb8+z26SzDLPq11RJoVr9DrEu960
mrol/Qs1cWKwM1kYZcf67jlsgkgaTTFywl2/oVt5rDWd/SD0Ps2Focp4h20ywmWc
xM7WNpAuA+KOb2AkN9Jp5G2QkyYJnAzJCe+BTTdFPVXKPSnYUAyU60z9IMv3+hK8
h5C4hoT1O9Plv7NLSUnmoCaHMXqPYs97LGu0bpCHtURompi/nTok6WjGsMO5W0bE
16NLm+K2/rQcyWFFf4gg334Fx67YSoHDzf97NImus+JLM61zelCqFD1519X6N1+S
Q6yF1b0n1TpSMCEiHK/zi3PghrrT/8byiZETYM16RwREkEuSDSnk0ZGAtQEBcr7B
yAMx3B2CYjx292zJCwI9vy4Q4TiR8COQBSO2C4ZCpmxomSUXJzToDg30REHn/wsv
dJ6twuFh8QqfF7MvVUaBaKyqeqNQk+chzUi/Fcz5BMdCNwgr0RCwrjl21TlGtzVT
l27Dc2z6t7HZE09yu5I8EY9oFDyRiBYv1pBiQYqoXE6qzRcLJ2UuZX57ksruXZCu
6E63bAFfF7WhCjATtsDburkZfmDWqMUz/IvTHfsbdFqvyzGW6mgKdU0WkXr8kaic
Uvt7gRb7TFtSxZ0xLLudWnmDx9qBUqW8tFTycraGaDaBesdrbNo6kH846+z8yViY
YD1iIbvsLvIxfea3C+7rtBBvB+e/XD0twJ0gMW7VKMv6pMqXrOOD+5dUdhX3zNL1
G/z6GKunkKb0lO+cHww4MAmSZY3RYrLZ+xJ7orB+RBreNKh2NNBd+S6TL1BEHyzY
MvzU2FLctzZK+aX1rA3VXPL67/8prNn9ObqiWNJIPJHxiZpimKGff/nO4SKeoM9t
DFF2dS9/YOAeYXm/2k/SIoeklpHmOcLjUZdclGIS3Yc9aYwiW2HkyjU4+dBusTsv
g/K0lkV8ivPr/v0NnUtuNqI/B8aCNtH9bovRy4U8YCQVsU4MiKG1rZMlmJQEPwRM
dfkXq46IDTc7Cyb2WCM2mWqOBb+LyQMMczDOHiIzJWHE6uFE2tEtAs+4owZGFWqO
LokG33TxuJPJJBvZ0aslDEXb+y4cypzPPuBpPLYoAy61uG9JjeQ3LWrZz+JWId+0
D+eSFw1k7Iv+9qaGKZyOdfwJCOZ+NTtmdkS0rAUFvGZ3axc+NfIWAzcEh3D0ypxw
E3k6IWbWfSuPhS4bEdQ+6d3HRiCoJSuheTKCO0RhtX9nFkA2s87NyF3W8/qNdhr0
6pqo77L/PPbudQTv2szxL9nuyfD7JEeaGISSu3cYFR+cJ2iiAtivnYik1LHU7eeW
WEINWACCidXnQGmKSoJDPJhhDgBYQd8aguUp6o/sD/SaEtE6RSNZpHCj4Za5vfcJ
UdeIwcQrbckqcm4c+unotRWa7yirbYvAw5PL3lzFE+ybr1x0Sn0K9HqIbXcVazEg
dTpxFuH1sW4C8WBezIQs4R61tSpYUbp+pGHw6b+T2QTm2BDqP6W4N1oACBdSvYLM
/n4ajD5eKv/OcA586yPJJjAbZADOgzGnkwIpSTaxSGz7DH2fMoyMILAJWjU4ngLb
dB46Lkc60Oa55apMHgYQhwgIpfvZYqm0Va3ZJ+b4kfCDx05uAo8JGJF/EVQnCOEk
+dRZm45pZWT8WpLr/Rh1m1XV8VLYKA3lXJL6trB2wLVpC69A9OVl5N4+efsst8Wx
`pragma protect end_protected
