��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�]d�L=3	w5��?�N��A-�5�P����B�[���훋�^b�sG(�dt�.KR��:z��X�X�8,E��c��DA��G���\�9��=�����*z?��'�]?�VUv�.���Ԩ0���L�sB�Ξ�U;�[�B����gM�1�·܅�̵�$����Q��^����W�M5�}�<`}�]مڦx�|KW��(`G=2[�'J��m����5�E�0�d�ܩT�I�f�[9���wt��f>�eo��k��F�����Z�jz1���(�+־876�����O��|"��Y݄v ��#�<�;�dWZ3wP��3�Λ�v����6ě�M6Ш]� �ಳ \��+��1��U������
����$8b� 0h�H%˂��>�cxf�T=qE�Dʱy�B���	��cS��4���f#�7|��?3��]UV�5N�/j�-�\ְu]�>��t�V;5ߚl�оL�MW(���Y��d���`�r8).��8�.�F��V�˂+$Ї]��6"��<7��i��?`r��R1h���@�*�%k_r,}�%f;⊽���2��l��i%��Y��ؔ���i���^=<%Ж���+�[˰�����K�p�٧|�H���iR��������:X�GRۅޒ�N��cb9��O�Oیbt#��O�)���h��s�Ծ"R��|�
�*����|<�#��V5�|�O<o;?���
�2��U�4I�r\f���i����j���jN�L"+<"�m�'���kz��Φ
��zP!`��^E�@ġ�f{v>[TK���u��vh����
*Î�|0O
��_G����8j�l�1�S�n\�YYA�]˻x��v�>�s�][e3~P�n�]KU+x�<DΞå,�����e��Op-� ��߶��A��eV��~;2<<=OP}(1"�.����e.,�{��9�8���I�8��j�\>����VIhs^�N̿;h@�?�������&�^:��E����v������ D�}(��)WT"���By^�q���d��)����f8	?�Q�!�QT�b��_�ۯ?�\�0�@��������z��O��f��#�Phr�@�2�ҡ�T8�iW��FsU��7�=�W)�KH����s����7�����H4o��ʓ�7��^D��[0��U�E*�j��������x$R��lX{���l"�,1�9�d�a7��[z��BF��Y�|k����s y4U��on//���k����~\���7�4G�������J��ł��1%s�ȅ�w �V��E�.�	<p:��K����z��ȟ�����\�ʀ+'Ce�G�����Q)ğ� ��29�@�ܨ̱��v��l���fɓ�o��=���7Aۗ �����O������<�pk�f�v[��y�#�=�����=��r����#4����#��JF�����"E!���M.�b�:$��D-	��Ŝ�F4����Ζ���I�ձ)r��'�L��]���_�#��[��o9Y.d���o��(���d$l'�pUА�3d?�ش|D��<��x'57]C.����#B�V��{���e�l���A�Cb8��Vw�yi�Z~]�'u2~㑃?�Iu2��|�ʚEgוҘ�AsK�DsR3N�-xH86����=]��E���e[�EP�.�����V�4FǇ&7�z\76���U�~uB`���L}q���s965�T�1�R�+nդI�4��ݓ�
;� �E!�jgo!�4K�G=����e�]а�\��\g~<��!�2�
�ǭBT�}[�o@ �ֿ��Ө��q��4�EW�y.$�i�
g�ت��.4��9�,@�X��l S+F��-r�亁�&�Ό�����M�(e��]�r�H���>�f��\mh>��x�p�GK�C|.s�bKT������k���^.�g��hn���1�hgZw����c�# ^�]�wbN�ǌpP$� �j��̎�f6eG��k���eg�m�|����#�t��"3�_���ѤYr_��0߬�}�T�d�ڭ_������4ՔKZs��I��D�AW��`��-��t�#�+y����{)��d�4���,��'�3Gt�<��:���^[�Z�)9a�K搣&2�V6쉘�V��`Í����V�vL��N/d��ܮ��P�����IX���Q�2���5�e
���%_��{;<�����s4�&*�~J���3�tr�2�_)��AZ��eid��y��91�?t?2�����Fw��Mk<U�@TA�'���A��Lq�c�<���*z�8��F��7eiO����^�N�G6�v@�͚��/ �#�	B`��l�W:��,dj+�l7^��I2��Z�˒�	������+Q���9����蔠e-������D��E��%�F�Jg�-�\�|�+�QY9���u���P�f�!�;Z�K�u��dnZ1a�o��6��I�û����O����oE/�~#�}��r��V�0 �"��>u��u����a[k�s����������f�yه��W���xׅO]��f�����A��"��w,�҄�w	�U�yrx�8!�-Q�P"�6,-�m����hh��s|��\��9�mg����CXfC������kPw�����v��G�?uB}�H���Dx(��A{�W��>¨I�m�3�"����QC��}�:�>�a'(���At��{���iqӈV���
f㍆g_^�O��Q8���jʐ&�[�Q-����E�������WJ�L�K��#����}G�������랷Z9?��̖`b���kn �s��oGR|�SԠ�$��R�z�@hVc]�$v=���,�@�]���d�H��l����A*�x�+�EJN=��H��s��j��w�Y?V�es��vpKT(�rG�9uW�Cs�P���A���yk�!H�Ylɺ�#�F�O�_?K�mJ�=�,�]�s�H�S˨3�>떍(B�fH���]}/�cLN��b� *�{a*Û���\�s��f�yG����`"�Jr��2K�!�|BMRO�����'OH�b��o���:�ݪU�l�m���h��*P�RYG"�εز8��0)u���F�V���;$ �I�o�IF�9c�q�!K�qTt�d�Dz�
���W�7c�m;@����&F���uy������l�ȶ�u�5Mk �U<���=Ul��R��U��Ʋ�֊��xN��[j":��|���]|�״�L�0�����O�*�\�y'\�[;�����b�ǝ�t�Tق2fb�p�|{���\��^󹯠*���ۿ�U��"c�Y�?�׍�i�&R�e�pY�)���'ӷgԖ�{��w� ��>`{�7|�ˣ�� ~�<Cd'�� &_�Xk��T��O�Z>�=Ï-@C��nK��\�1@Z�َE�hV�g�!�T�j�F�,w�`�qk���!V	��4�&���l�4`1&��Iǧq\���g�fv�NC���a/��r���,�m�����!����d�`�����#�RƎ�~��Z��V����Y��>�x4���1��۟�3pX�2�lk|�Fm�n@�����u��%�)2<0�s��G)���0.OA*���'7�dGS�����a����qA�Ď��s#,��Uq�!��|!���ʅ��h���g���I;TJ��F���Љ������I��C�{�\:�T�猓̰k?d��.B�؀{� �}�7�,�1���U�&M��اΤ�n���,�J�5�zgg�|�:�����S���@�c��1����)��>�"��Vu���=�J���JQ/�I1>�z�E�T�"��C@�.ez[Vm��V��_�������S�c��Z���|�@�h)i*M��z�q�N_�@��9��D�������ò8e�[Y]�Zwk��B/o� >tR~�v(zB�x��ցhv#���P��ӹ�C����]�"���|�ҢB��ve����Ґ(w���*2s��+`I�7�D�k�e*�Y��p��¯m98禦���>-"�Nۤ"BpXdݲ��uo ��9�d���oy���R0F7��"����I-����yl�Y�`AD �Pz�w�-�/X�vZ��E�B�����_#���c�	u���6��%�bEi�ц��;��f�;{��Rˊ�~��rߤ�֘�7۝)��'p���[t�W��J�р�%��{q^P�)��[)�|�� ͝�s��������l��G0q	����qZ�e��|.g8b�*_<ѯ>�<y3\�1jO�_� ܙc��P�!8!��f��XD �
��B���h�;9��'����<أ�fp�z�?���p����F��
m�w�]��������?��O���B��x�@�S9��e�dk�u���6��$Jw��R�ʳ��b����	?e �A_]���^Wq�F���eC���c�l���d��k�ƁV���Y�ApW.$�Jpb�����1*����:����7�����9/�ӷ�&��yD)�2S�����-���:�8�=rՍ���޽�h� ^I]t�m	�j��R2��%��?��-xwWo��Y(D
�Z���$��E?�e���˒><���ޏ�`%����N�$��(h�S��l�*CI���̖�6�\�W�
6v	<��ŵlu%r�*�2��u��}�Fo��ډ`k�[.Hur�(n�������QQ^hi�?������ ����ÙiUA��態F����cM��^Eo�g���EV�YTP��CS�!��MY��믅�A�P�:��}4o"��G�0syFZ߂'Va����i���p,+Xˊ2���?��U��l����د��f����_���n���5 {Y��<����z&���kL��,����Ě�R���