��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�؆���o��9_��ʵ�Fꙣ>��IG�'���-v_�=@��*�S����k`��sj�a��ī����s�ޔ[�*
�����V�C�B��:�Wb�$6����T�θ?�i\��h65�9X�s���}�@3~j Й	]
i�+�����)f7{��oe�����
�h�1��?1p�~yb)���R�Jd���f�g����h:��'ߺE�őm�Q����Ao'	�n��R
��tƟo�:��zy��}E
gz�
��Ls�m<���nɟ|�ׄ�^��Z��wA�|�����=�_�F�T���sY<�DZ^��)��ظ�DݚN�������^�P'(ۆ�қ� �K�P���{����)
�^���슸����7vN]1mdϞ p\7���xB�)l[�j�f���a��G�mѰ��f�ӐC�rβ<3Q����~�>|������ZS���5�:��8��+�����൚<�t�eތ��mϥ��|�����&�"mu���P'��	Zm�h�MU;;F�Q%� ����`+/\��<lRzk�?���W<�G��x�.�4G_)�<��2�h��FY�9�� �v���c�(C��߄�qYS	��'�N1��0
���}�̪��	�d�A�4`�m߽Cl�/RJ2\Y��'�,y�.GJR�\v���N�`�H�k�S�����F�WL~LmlJН̛��0�;�`7�n�6���ܡ��۳���9����}�Te��b5�;���bX?��9xC��������H���b`��W�v̾����g���8�.ك��q	#�K�˝�T�N9��0d>lwV��h�˒��q~b���Ԣx��ߎ�v�Y��=0 ��RD��J� ��FQ�'�3�pr$�31l*"I��ӛ�'
0|rd���nm�����/���Oڸ8�ޭ�7TsV
Q���BL�S@���תb��qJ�)*�]ʢ*�a�ӄi"�T=���#p���x�����xv�N4-v瘖81�!c�YSuyH3�4*���Q�mm��Z)���k�vӁn�ɂ���I��2_�P�Hew--a��y[���j�, =Ԣ��b�ƛB��|���`W��ʯ 3q)�È��Mk�
�ئ;��&$�ǒ���B������M���;>'��J��kXP5i�-#�y����_	����ʩ�Z��CeSU�I��/�֞¥E�E`S]����N說��\��Tm�2����D��Q���g���W�gX,�O�wY�se�&3?{U���)R��R6�g��=�(�$��`X5�^͎Sc=ֲg���|�wMkydy�Yl=%����dQc��S��@��]`���b�c:a�	�^�U_M�vz5Q�W���ZC5r�+���D
eq��~gh�&Óq}��.��o�!��D��ܱ+��J�e��Q��^t}�[��^������+2��B~�f�w���1Y�9"|!Kmi�1�.�g���.��Ć|em�P�E��	�K��r��ND���0B9swXGZ��x�I�s��e��%�ra[5�Ѕ�,Ռ�:V���"P3��O��Jc�ەx�Q�A&若@�%,�0T"����o��y>Vр�m�c�M-j�,��T�W!ޘP%���F�`ߞzk��"94����U �W[9�{�y��� �O$� !ŷE�_����'����P�hs]%�J�����0/�;��u}�#jM��=l=gQ�-�!1���69m^%�4��q��Ԕ��qB:c_�ϼ����Ϳ+�3����R����Ֆ�R����NM�N�@p)�e0��i�39YO<��N{H�P\X�(|����j��M��&�ƚ�۔���H�Q!ggg�s�q5�?��T"E�G�L�ƿ�8�*�$Zf���,N�����A��K��!�2ݒX�g�Y��^�hm%�o0-W�u�pЈؿ@
c�l��;R����N�O�4�TK5�E�>΁�h��,=x�ڮ%9saX�rAT}��R(F9�ʒ����YY,@	��sc(�d�����&�(o��.��eh���:uQN{Y�x��/M��[
�f�Ӌ��66.�~[��m��X$�	�o0w���UL�g�6=�R�0�A+,`�y?�Wޒ­oB�M1��cVLd�C����W�H-t�5�ҧF\CzA�o.8�d����QLi[��ȵ���>���_c�>�A��'�va�����4��S1a���h�e��	�r�Dp�Yc��G�*q�_��?LT�i�V���x��Lx.�l�goZ�T�KXg�t����I�
fU���[������x����c���2.�����hɺf�ʪ�{R5m:l;1�ʥ^�"�W�o)FD'��ө/$n]�0��i�ʇ$�iӛ�P-@�1�y������c��)���[�?���,cr�M�Ub���g�b�?)w+�:�wC����h�=63�jS9T{ȭ��
�/�c��0?�N�g��+O_�ޑ�'A��4���ӡa��^�=��4�܎�r�w�����X�^��>0h�N17�u�9����Av�;���\�B���N�1���|��E�&��޳�lB�̱V����8-:�5F{����ю��0��m��JTn_�P���b�4�'�r*	{(l�������v�-#���Ut�e7o��e>&K�o� ���5���)����->h�C"��e�S�����~6�����8�z��+x��qH;�6!�82�='ڨ%��]|�q��F���؄*9��0���o�=^�Hz�77����t��?�Y#���4��)[�Ix��K�C?M|�,��B�r��A>�iSd�dS��j����~}��fL�d��\��ydh�H�t!!�G�||�[��|�sHIEP��!��q\�O:��u�+D!�Ky?�m��J�H?�m�0�F�+}T���~�����~���� R�뤬��	�H>Gmn�S��U��<��;��Q�D�Qgo?��fs�ڍ��U�cr����lG>ګ�r��R�ۇ�)����ed���>h���B5jX�7����%��HH��uK�>��S�:�Ş|���IMi�=����=�������F�tx��ٺ�XB ��n����i6���ܲ����& 5�Ն�Z�}V�� ڙe8��|:\�?�+�9Jg�x�L�wnSgó�Q?����p����������1>&,�� �{��A����$��0�],@t;s�2n9�o�s:^�k�ZX?�p���ru
\?��3뾅�x�Hg�
 z��Q(�~�����z�]2S5Q4�nV0���RJ�6a���\��L�)h��VA}Y=)�:Z�MM#o"�bb����#ݐ6���1̈�g!�k�bY����w����Ɲ�a'!�XObsa	W��l�����k�'���~´�2,�����e'��r[��=�z$fa:�I�f�=��
]��"	٣�G�
ߊ�>�n�L^�D��ҽ��,v��"�ip������^)���S$�1�l�����������a�ǲ5��1S�7�� 4M�9�T��t��r�䯷l}�C ��rÃ���wHO��UT��E��W�%���7��ByH[ e8	��N�����'i8Nd�Ԓ��rn�~g7�U�Ʊ�f�(S�x�q��6�3�ᔞ���WRU��Ra��Űp\�������4`t *��#I8�)���,u�|'��` �C��<�_�m)@�n*h�:�dE��Rs8�H��!0DF���&����������A7u���`��K���,1)LX�~+P�0tif˶hR��U{*O*p�aޖʪ
꧟�7]��.�J�{x�ZI�m��`3��Q6�b]l�wMP�ṘhK1���(�Y�T@e�>�OM=� �y��в���Ę	jA�H|��sh�+�w�]��a7����7�LZy�4�m��lx��ǂz�~�#Tv��r8P$)�l�p}9P�ʟ2kIR�K�R�\�y��-�������Ż��T�el-�<>� �F���?�\��$;�a{	~�4r�u�+�(^2��5�ŀJ�*[,��ώL���ǯ��]�����=�Z߈�d��4+?�su�k��]W٣��g�?[>�1z���!�C=���h��/���_džr ���B���S�:'��7xm�$�{*/�	Q��+�z�$�p+��t`���Π���_zq�
> �����ԟ��\B��T������:�z������C�As�y�>�`�b��̈L�N״#l���n������%�.q\}�_��L�y�wxf��ɽҐ�`���?��k<�Q�8��Ǚ�L���&m����˸bB�N���U���=���jF��"5�|E��Z�c�傁1�p%ζ�����1O�@�xj����vE��ku}���[)!���z��S�󒮐��,!�w�s��ͦ��I�l/ݠ]�(/.����m�l�v+��)�%3��2�1�%�?��GҝU��uf�)�8L���z�l�R��s�W¥-;:^�8��@e����x��R�]�O�z(��T�n�==���E?�X[�۫\���s���(I��Cp��>`���~a�><�nB-uj�B�ֵ}��6�']g�f��0��TΚi���t-���
T��E���B�o(4��P���>j���=���w���D��K��/~7V����g�Hس2�P'g�g��"��U8����-1��x��r�=2~l{b�7�1%C�fp��A<�Y���=݌a/���˿����=E�r
��N�Vq��c[S���Ӄ��i�Kx(��\m {L�jZy�y��\�A�Kjdh$�nހh��eX�u�Z�,mZ�I⦘A�v��Y�P-���a�2Bm�I�3���$�a�-��0�K�E[��29��5XͱƄ�W' 5gɻ�<}�#M����9/��&(��w	�8˝8H��Q~���JД ��Q$��a�Eۙ;I�f��Ƽ�[)��#I:8~"�$�1v\�;�7N��d��Cކ�h-�z��� ��<z(���Be���[�A��&�g㏲�5�n!t���?����M-9ܿ��zX�IN�UoM�9��\�~�����#�\H��U����t%�c�NBi�'���U�x�a��k0��)o{s
�D%��u���0�Z���ce�H���0���w;����J�XFJ����l�Ak�-fά
D����^�ШG��$5�K�7����D%��<N|ah�c&?��!��T��R�W:.�?����e�ԚXc1��+#v�D�ʯ�<���R5�`��4��K�@ߗ"9�-��+hփ�YQ��e�rK*�n71+�P%�Sn����8cI����ׯ�ʞ�FO�v�Eډ���(ߕ�^�~Oh��<��n��5�#&+i��B3yG��8��:� ��Ydn�lP�����7��NAR�����t`C'�n��Fb�+��� ᅇ�w4]�7(���i�h	�&7zU�|���M���(��@�Re��i0��8��1Y^.M�]�`�;�AP��IR�r��t[�<��	�4�V�`N�#��of���@?�_�\�r;�{hM�;��t8'��ٯ】֑j�Q{$5�]8�Z�>_R,2+66Z�^�I��&x�}��Ȟu�k��0�S��y�m�+[��Z��~�ۚ�]�Ez�B��)Go�#1J*�m��+��r6>��F���57�`c�b�e �$6A|�d
R�ެ5�`�� �E3��S�M�fm��@bB�O�Q��"@��ٺ"L8�v�.O��i�-T�ϝ����w�t�7O!�<2o�\p�>E�x���� E����,m۷fE�|Lt�ܦݔ&�|hU�h�։H�B9���j���*-��{�JO���ث`�pmݳ���yfI�V^��>"Q4k�ո:��{�9�Ǝ:�մ����qPt��[�à�"�z)u�����9�Sc�Y?��;F��1��`��� VW�W�ʈv���y_�AS���61��F�+@Ǉ���9�ݐ��@>(��U��H�L��J>�/,2%�e�۟r��*�#VU�:�~�w��"u{]9,�؄K"Ҝ�-�����˟�,EcLhʛ��Ў��y�HWD^��B�@����7V��4�0�A��~GI� |i�;��y���i���������1��.�R%�y:��*?���+g�B�����Ys�+��E�������9XT�>��i2��s�[]���xO��|`��Vn9��W\f�IϘ�������tj������5S���p����AhL9��1bW9{���fCZ${*k�7OȨ�
��В*+��X[L@�;�e9�ӭ��C7	KJ�Zhr_Mp��!��[*�w�>)�@�z9����JHDDT�$��7̽�þN	9%��T�14�ߑA �̂�Y�DK�`�>
��rt�Ԥ�eh'��)��`j�G�tqc�`:Zt?��JE.�� ���gqL<
Lf��Q�3X���"���|^�KF�A��害���ɯ0�3�����oj�,��j��^fIA�BЬ]�H��Ԫ�G���:��O��;�����q�RDO� m�AV��*~�3�WCG^ϔj;���vOi3�Yoߦ�����3=��_\���xv�}�����$�����k�b�Y�