��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb&�L�S��O�|X��0��<����V��[�^�)�I�.�t�,����O�z�u=*"�8nY�p��y��P9��#L������t��{x�
Xg?���jE�,3��69�v8�@Lt{�9w�M%�CBu���.(�{*kz�~����N=q��Zq�%�OV�a\{%y�0�?b�1Ř')���$� 0F����a�B�F9���Rd�5Jϝ�
�`�
(S���ڐ=�|��-z�Z���J�8��"�@��2������Ϭ_4��l�ၦ�t�7@��v.{�������;-;DM�ωp�g�7�ltx5kcZ'j�Jb0Ƈ6�el,'�AQ�	t��D�0����@u��M�F�*�F�����Em�ePD����E	][k>��P/����(��ʒ%>�kk�_A��/�i�6� �"k�'��.������XB�`�%���El�ِip�S�%���}.�-<��^)���oe��S���Տ��YG���w�����,n?5�
�,<�ߒN /V��Q��С�W/iB���{Ӵɏ-�8�N[��a���&���Z���ߘJ��1"p�X�z�.�(��&2�p���C��^�������v��B%#J���.U��?*�/E��4�۪�NO���C>r��ߵ��67����iA!
E���y~�i\:!�5��5LƠ[ↆs,� �|?׿CО�uUW�_��6��4r�߀�D� ��߽'�c�jN�x
��J��>���L��U�]����z!����]Y����ȭ����ӫ5������O�����2���j�DPk�8o�P���dஜ�K
6�ӵ�[�<F|Y,B��F��/*�*%%e؏n"C]�`�u'�q~M������ݤ̘�R5-�m길�)������;K|-Ô|T~f8r>{�:�`)l�1A`�����rd:���k}?ς*��`��^�n6��id���G�K$�s �ӛ:-�d�d�ڇ�f:Q��2XI��d�5X�0�?����j�4��D��Y��hqu�c7򭅬~�йFf,Ҡ�p)u0�7^�;��VO,e<�06��n����xv��8��qN��y���;#-�ڱ;���Q�d1ʆn)��b��O��T�!���6���)d5=�ɴ���N+1�$|7ְ�\C�j{��flxʒ�%@�mrTQ��wp���|?�k�H?_ @�!������/du�	E���6n����0y�0����'���U� 7�d��k��,�JB���	e9Ǣ�z~
����6��!��$���P�88;�/�gX��_6�J��3�o�hד�Kg���d%wAo{=���&�!�g�j��/z��|�~6��j	���c�,P����U��0b����F�%�]G7�@h(FOҩ��̕��^��d1~b<��e��ynU%� ���?R�d��ǿ��hX��wQY��ԡ*}	9�N��t޲r��N`Z�A������6U��P��,`P�'�b95 �m��N e�́/̧v�V�:�n�tH1�|�֣�Ԋ�ח�2��!^wͨ������V��#�	/P_&�'�+Q;O���=��ģ��4�����w�]R�h�(��^�ʹ�Qё3�8�!z�qO��͐��d���P�t�W����sB����v����\.�̟s!Li3�ܰx�U�+��y��Vl��}r~�>�/���8����(�,c%�l
k��+>:�h�K��.�8���fI/"(��s��
Aƚ��À��Nb�7N08N�9���@��G��[����^�i�G���6���Ás�?됏�Y:����;�������u
*��R�C	���h��~�`�}��[��p�o�o0B-�v�����WI=���ޕ1Pi�Tҍ]W��Z�

�8cѬ�?5��WH�!�9�ֈ��<z�<���7��5^]��n�4�\'���0�[[��5Ȑ�X�Tm��?r-��#�`b\&��tL6K��W �!�o�5��2���~�LVѮ��-4�g4�u���6��= ����F�V��J�=���k�_�[giB�����ɲ`�i-�:I9!/a$z �|�}�Z����\1��zl�/��RQz0�~�MɊz���=ꋿ��H�0Z���u����y�����ߗ��\�S�y��f{-PL��!��s�5��a��TR��"1��{pV�`��:GQ��������1t�&�3���j[#T��9S�똚�L*�j|,�E��q5�ً��,b9��5��K/sW���`'R$)xǦ����߅�a�R(9����dրM�r�������;�x[a���:����N�.��ӽ�ҵ����-�9VqL��p�|�P(-Fskj.�2p��V&�W�؇����m�u�b8��xX���@�l
8�����mc�3�1D�֩.�P�)!���S����G P����ѽqCz�jx��@�.,���L�a�@���:�*���/�h�?Z��ˆ���U�a�kL�ª�'� S������T�:&R�5q�o8���z%��sX����2cB��wE\�r� <l(܇#Q`��Wrd ����y��s����q�q����)3���q0�U�eIUd�� ����t�Y1�w�@F��ps	<Pz-�\�q��:a�
(A�d*�E�����:�¤���ؑ��oYo����c��[~	��)�����O��e���:�0��X&�=���P�IC�����:V�N�W�փ��r���N�@���w�[�ڡC�m�_��iWz�u�䬸�::�穙D�Vc�<2�6ˎ�$��R3��4=mh��/�ѩ0\k�b��ii�DV#��F�����T�YN͆�nY�K��Q���:k�#��t�[K]��f>��-���F��TI��r�65�s
�
^,�_]]|�v��������/���j4xZ��G���>-�����Ce��dn�>6.��g�d#��}�kd^��[ :��o�jC{�d���^�2A��ka��`�1�	�����ǳ��VI��aۇf�Ir���9�[�V43	��+T:G:��'��U�>A�-RM[⊁���E7�T݀.G�5��o��ie���J7O���	]#
+%v~+d-���"a{8w�a��+�m���I�Ԏ�y)A���sѯ������r~&JژI��{�������B�Y3���ùp�'ț���x �%��tu[�6~cYI�ymΏ�?������N[�:p��U��.�b]�?�je\._!�'� ��������}�EY�b�BT���0��WT�"̖��O��Ue4�A��[���T9EWg#��-�W�-�9b�����<��`_i��qCd����^��!��|�ͮ#�i�~uqى]Wd�2�`�;q��#
u�9cw��Q����|k�*Y��v���b����//��ԝ�:��d���=�T_�m;�:�!��Gخ��ĥ�*��0*�+��MPU�����E�W[و�����y2y硥�єs�2p�W�j>�z.	@2�C��!\�VB+�PRp�K�d�ػQ8�,PѼ�)P�L�0�o��d]i��Y汍�O�|��r�/nhk��~6�%^�O7�w��7��MF����4�	��H؛�G]��{,N]�H��]A$ޤ��+�nx}���b<�~�})�*{�E�Y�[1�=z}w�W�L���#�ݸ|�.?��,��+{�e��%.r���ۣ)�)�|;�b��q��-�?��{#�"M�w,�.
��eun�_��}[���vH`q͆}�ps���]����<��$�)��B�:���x~�̜��D��#f꓆[�F9��_��]Q0 �@�b�B�-�_؜W�|��䗸�2�j��MB�6~ʳ���99����Ly�bn�!��LQ�}W�WQ�+DAB{���O�l�6K�Ϣ��C򸮡�b�atȴ"�+���95��Qs�ьϰw4�T��=ب$����[5^�+�. K0 ��5��!���=L�8��.f�j����1�F%�e�1q� �p����Zr��*�p#����U�>v��m���X��_�+���z���+H2SK�b�������:238������
�c�wp�f7��f��v�C�*�P�W# ��|ԣ��6?�G��h�7S&�v�s9�ST�F%��Z_4_�M��
$�v|L� D���ӶѾ���:���c���#���c,�uC5:��9�Vz��F G��5�f�(�����M��� �|.&��t)x�.e�� ڈ��`��=NOd5Ԣ菋_��:zm�'/�