��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����,��f9t���3>��Ձ�A�7M ��uj��M�0��{�ơ�Wa=Kg��!洭D�2�&�6����2�����X܋��x� ����G1���w�S��3�C�1�9��1+CH�<3�vwN��F�T�\#[�'I���ҒO*K��V�6�k%���D��Sn�&$Y�au��Q�/���OO .�XS}���9��k,[=0�hj��V���w��:g�!,;�(���1��+�\�dn�/x�o�+H~�ёn���c�~�]�]-��A����Vd�FK��J�X�� ��"���I�i��j�S�u�,�AN������������@Z�9��\�ݚ����k�>��sgl�S�;�э�2�qEEE�(8�`h��]�Qػ��"X�0�?� �S��k��H�i�G%t�8ZI��(5��� #*����ڏ0�N�ޮ�끭�J$5��+3Kt F�����Fp��fS�j�`�y����82����{�Pϒ�����gV��nx�����8%V���;
��X�V��[9� �����X,�þ.��-���~��UX��s���B*�;������ES0\��;�~x���`��#"�º�@{Bj7��;�g������qRB�R��X/k�6��Թ=6�a��3����H�Kp�D2H�&xOSx^B��?L�|[f���e�gq�����r9�ҕ������g�i�[���:vp�OD�u�;sy�o.���F�~�
 <��+ �#��
�ܩN�9����9���O$i��q��$=�ʯ�G�2=�
L��4�(NC�g#�HY�3fg��u t���#��"N ��gN�W��E"j����G��	`P��G�2�K�0X�!�kZ���L��;�O�zlbݶ�0c�l�mj�޽+�_����pe��p��Yf:_ix��Ng�~պ��:��Jǌ�a��������&w�Uh`� 0m nyf���§�t|.�h�M�*����4�?����mת��j������;�r���'��7G/,�>��{�,���(���?O�=G��fwQ��uF�(cFq�����Y��w2����X�c�a�����!�"���Y��]�f��B�E)o��8���@���T�Y�eGΊ�;���[D�17�:�L'p��%m�h�	�d����5��p�7�,�p�%[���}� ��N�XA�I��y���~�be�B4γQ-:;��_1�#}鏻 e���[Z��p��z{~�G��ӷ��(��l(�ߍUwR�˓1�@�齀�9{<�c}�_�)f
�%	<�Ԅ�T�8j���C���z�p��b��r�����a�����bx;�N�h��RcҦڷ3J�P���,è�����y����/L����kY,Ȼ3tz������sHĝ�����`�P
��(��澑�`�3����>uhW�~��{�(|C��R8p3{��������:i�|��4�8E0����7�uR�oұӚD<��
]����\�Aբ���8<��@ZS$A��@a�]f�#)�\�+�A}����J^��3m�&Y&/�2]~��@��,�b�þ�/>{z(��7�9��+�v�N�0�V��@�u��+�Bf�D�G��	�va)�q�=��Mծ�UG]?���Ї%۝fE}'*�^UX�k�<�]�@�� ���r� �����t%�ɏ������飑�L�)_ҧ;O:c���4?2�������#�KS�w���7xT�M��0Nu�6n��;ǆ����7si$L�N�&���)BOS.��@@Վ�*@�}`��
W��E�`�.yS���\&6(��1~�0^:�ѬDd}�Y~��!7_ ���<���^���l)��)�0�g8�m����pp$���΃C�i.X��=�L�8ν�Y��D�XINC*M�M�G�m�]�y@��������i�EVT��f[`�|��c�F�;R?{<����
��M�C}MPս� ��Pa�%�kH��C��0�b0�&�\!��q��1�
������H{��xk,�`ը�����p����ݹ3 �H���˶ܾF�
a]z��T�M�FE��r�+�N���N�g���l�e,o�!-��0yp�~�|�3f%	Yu����R:��祷�~��;��[-��ߴIc�'/�d�>�{mU͜�F�
g�|� �K�YϚl$�_f�M
�mu��u������8�]�+��{
Ae^k���6ٕ9'��-��_A���Św���q�N~�����Hk��-f�C{AA� 6�5%�`Ҡ�C�[��fP���z��oB!D������F�
�L*�)� ;����g��	���{w�a{vN�%�4���Q
����p��dK� Z���)�+�H�Ί!}�Q�B���}�`Y���=����x���n�j���kDǙ�&1��~՚��6!�[O��z��~>�����u<��#�Y5}�]n�������r�iRS�5��o(؍wo� �U�/.�r��yXq�DN�]�PbO��6���,x�Y��&���c��]\�E���EA�YG*�--�ߢG��{�X��zl ��>"���ྡ�~���Fo�[F��#^B�����0�~�൘��/�H��Q�����_��m�G~�7rI0�)�3W�����$��]�);'l�A-��W};�4%�7������'�+5�2u�E}��M�Y�i\�\��y /(1w�[������]��Aj$��]�?�W�(����N�B��sH���!��ն\�<Źs�&^a]����ݖ�}��.ZZ�U��T��fS�k��
Z���P�*/P�E?������][��$�����~@��%SxۢO<�I�8��u��9����C�l/����X��,"J�b��3rDvu3�v�)��"՗�<7���./G$��zw�Z�ٴ�@�`h^?M��X{%L�p��_��@��Sп!�3��-y?Zs�R��s��V���+Ё�>��F�z���mp��k�o�vpK� *y(�ҍ��;B�y���=T8ЊVC���Y�`�o3���z�
*�����";d�nV
����S<����.�$7T[�7�&:�����g��qr�1�xi�X���TKLM�{f��gT	����������҈\��I���R�1���	߭[�v}͋�t� J�2�#�?�g��k�#��%�߷X�VE#Y�2N���:�*�ӫ�Z� =@�M�ܮ�2��w*q�3��ل��9�+=]�ؖ\��*���W���z,��YRZ�5� �2|F��y|����ɖu9�RZg� �-��D�S�dVl�h�� 8����h$�>��0vHD7��E,�b���K�u��(6�z�y߶��&�-�͢���ΧN���a��{�� 8y��9�u6Og���<F�����\��e�=��3S~���Z�m*��'��w�(�:d吀|��=����?�3B�1��a�N�^fZ�bo�}a/�jO��N�Qh58�&�.�T����h3�{n��Z(%r.��K_��M
�ï4�j6ݖ����pZku�d���\�I�E�A�\�\o؆�,9�.u2h^�J��ʴ��N�y/=�$�����f��`Hh+�x�������pF��1y:%�P�����������3�y�O%Q�7���Ea�S��,�NM9�=��L��3�:�_,+��r�,��:�����3��3�PS�*'7�ks�cL.�֯a,ň��k�ҏk��L�2=�7���D|�fF�^���ӝ�����[M�:WD���"�h��{���?6D��.�~���I�嵟�o��NNlmw_Yx��/�?��%6K(���?�4�"��pyJZ�{=[�	�]T���G8D ڕ��|Mj�6؄��U@&��%�1���r2�����azD�ȉ��T�͗�8�4eGB�ۋ�+�[P����QCꦶlx����-�Q"�A��D�}U,�ܓ�6�Ј�`�p���!�7����#�y"W�N�t����?p�)��ƛ���ڕ�VH�[�rMW�Hz�>�Buv3B3=٠�F�|�*BB�6t�����@?m�;b�^jͷ ����,d��Sm���m�%�I���_�*"�����������ȿk��:{�JTS$UpG�kh�.˷�)��4C���I���.�Xmx�F���uy�9�&Qb��u��k�W�;N����B����(=I�I��+��~Z71��	�Z+�6��;� n�@~��l`-2lp�!z:�rF�`
"Vi�Β�(\\����ҡ_�qG�w�MM��MM���d�^F)�:����3���+j������AI� �~�3ߜ.�.���2��m���9W\+���c3�
n�:o	ӝk)׳_Ȑ`��O1Jz6~��ԏ�(=���G�����x�޼,n@�	x0���ɋ�4}�v�p^�օ�M��~ 8Z��j�rRm�]�fD�v-Y�����.�6������[����u���z��׸��N�
����y�X���K"��/�����o?�`�B�d񽠸ym��L�6w�wcpM�BU,V�D5+j[��.����Y!����P�ִ� u�kk�&l��F�}-hßAE�d�p��ǻ�ʞ�eG���O���z����	)�����l�ѹ�mp���GI�o��_m��	6l�p��uCG0��~Jͫ#(�d���Y�3����ϩ�5k�ůR�d��v��I)�'�(E,
\ׄ�+܊������f(T~�|�X�P�8"MM�#���#�e�5���w��[�Ij��t����F3��a$ӄ�Ǝ�=���0QA�������ǽ��)`�o1��ׁBH����lE2$�6��i Z�	���O2��˰'а���#e�j��\\r$�z8�)��$0.'��˚s���5�� [z%���M(��6w*�!M2���]Y��FԖ��;����E�������Oz�QG��	��8C-7�-?1��ۄ������V�aN�U.��_t������g��Q��;�D�R&���@9%��'oCSr[�
��\�Y�^D��W����oÔ��W}A�:�5�sX�~PcM/���>��ܴS�&��W�ʻ�o��n=�Z��U.�^α�\�S��2f8���U�}�zM��ň��ƚ�R�lŧy������.x�y�KzX����|4��z��S�G�����㏞�aۺ�B	�>ak�1!����ܼ͌C�����Z� ;iܽs��A�Lu �u�3Ie��l����L��dC�Ra�����;�� ��9�0�j@�
��t9��t��"�}̅�'�+�|���w������	��"����q��R�����5\G�`��q����u�̛i4y��|��OR2X<��.HS�=I� �#Gﶌ6�{�µ���p��Ce"ŵ�����-��聦�3B�ju�ox��<9�ݾi�(�n9nr��,X���Dg6��]�"��j?�dL���~:op����>�(�$A'��i�fy�j����$��'��>�eʶ���_"��́�O�HOK�t�M"G.zb"�����Le�6/��h����G9tS�\Q��|���ER^wSS�PLr�u�.>Ri ����L8�_���`>QفƬA�1�Z_JN�:uTS��V;,��ޒ ��ҁ���Os$s}�u��Y���\Ϸ�v�B@@�՞Mqy�e<w�	lRg��|ǘ�jR��'[ע�1��/h�ro%ܵ����f���|d�X
���!KLCb��@"y<F��N�]�H�/iv(f3���R�p���{B��F���;�Het�L�gw����R�U����Ԁk���\��?��;qĊU3uL;�R�S^d�C&R�*쌖�R���!��4l��I�r��Z�����a#�����bń����Jf��ސ@�/9+׈�GF����?{	��� wK��~���gKo��Z�NR>т��t�S�-B"�e�+���h	�E��Ti���񯬞�<��1��#��~��!b��K�eQ>.��'��UH
%y��*��j�w �+���.�ʧ��1Yf%O�Ȣ�%�ڼ�l�B��=�BE�騺���&B��H���"~O`Pŗ�Ó��]1	��7_��y�v�=tT��S��"�K�4�v�jHb@���K@�P�	k:`���L�����\�6j�i֏ax��LI,���VL���r����S/��e��?�/���2�6ڵ�W}�Ss�"p�X���/B�K�p����:��)57�?
ɤ�V=i�q�c.x�.9Xy�
@O��u��������bf�e>`5݌~ՙw�Q�+d��V�>����u��XE�ɹX��3������ۙz�xV-�������.'��Rr�m��U�ڮ�A�ʐ>�Fa%b��܍��Q9�Gb�Bˉ�5M���8m��`ӟ������o�G����N��\Q�ծ��hB8�80lON�1s��ZT����T�!�|TE���Q��H�'L.�Qf�/~K	�>@
$y���0�MB�2���J�M֐�٥\�����7��$����XA��6�.���(�S��/�Ī�_v��ų,�MZ�	����4����7������h7Vm����r�ZB��"!L���;�|�v���P>8�t��vw�N8:C�"C��+1��F4�g��n�?ɽ���D�w`��|�]�i�	�b9�q��)�g�g�.ߠ�Nh���\�aI��_�	��n��U��a�1��v�����7s�6|i����zaH]&��݇^��]0�`*�D�cPhb��-�b9�w��r*R?6���:F/�f,��^����L�0t[ T�ViF���<�z�UX�T柹Q��4M����dE4���L/}�+sHL�ț}?����#M���(J>,r0��$��G�c/�r��	{A'� za�&Ī�Z�����[�7+M�"��b���d��F <j�.�K����k�t8�QAM]����H5���]3�l�5�����1�2�X�9d��.�JL��dfR�� >��Zxw��**I���E��DO�ؔpPTBB�k��U�(��� 0�T�W�=�xN��O$n����Sy��V�e��֨��B�Ĵ;6�^_��!:k���`�~_R���2�Q�M`��Q~�v��p�m��x_'�"&��$/Ms����@���3J[�����c���z��h_����5OTB�P��u�;�s+Q|��r���m�9����Þ�$����Zy~�۔���g�Xh��7d�v��x���5T��I{�|�\�F���VW���~�
)���g>9w�@���A�J]J�uo�%D���W-��؂�]qx@E����K6d`����Q��.�����s�v�%_	՚��0�l��ǅ?��?Ę(���4{�ay���8,R����`a�M�v!b3>P�r�D���-�6I&�Ϊ6�#6�.jū������#ݝ��Ԋ8~�H� "��Y���h!�ϔ�&�!�ji�H�%u>�:��|ɔ=��=�u$p�?��� I�����f����[Q�ջC�挚��;�MR�(�#���ƒ��0'?莌ހ&o�ad��sϑ$'w�lr�&�Z�!d��t??�m�]`���Z�6�<'K}�S�A��A���������j��Yt����dr�,F�Y����d�G�TKH]I��ؒ5
���`pՍ�{�_�2����13��,�AR�EKv���fc�&]�Rz�/S�扒bN��0��To�3+�j����w�֫�H�M������b���'�sv�]C�\}	�4d[�NÜD�=���!�5��H*S��GS/�$4��2QC�=��<��q�Ը8��~����!?�NӒ��_�7��mp���Q,w��L�5�
��_�
���Bos4]����B�_BX�b�b�d�s��G5?���c�)��m}s�����py*lk9�p�&Y�I&���ؒ!g�	U�5��8kl���/���P.��W�
�p���m�E�"��9e�KM�$�W3���{^7 �qASe'��7��VY�w:���X����]8@�%�lM��P� ��q�$���it7^���y/�o�e��ԧ(�f�ڪ���d��8z[��bb�1��wK��PT���=�tN�[��٦?�<�b�Tn��j�&���O�N�u��f1/�<�>�8�R���� ��+��o�����:lKA��(lRPӺ�U�����0�᧧P��9l�r1�	WF���#��4G�QK�}q	��ߞ�b��Uj�~�UK�Ǌ'k�:i�����[�K��	�r���M$�lR$�|^��<W�6M�$�w�ynEN;�=T� ��z%vU�[u"�7nMP±C)��w�c?���"��~S�0��Kc[�h��-��`����`Oz�?��e����bE冶��_�h�k���U��(�F5��f?ĵ9s���vmo��6��N����[{R��#B
E�kƛ>�{si%x�����Ʈ�TI��M ��O=k��#C]�#�����}��:[fK���ضd�(8{{>;��^wM[��icor�]�M�0��G�V7��s�	�|~v�o��o���zÝ� 9����`�n[��j][	N�[_�sԫ!��f &�U'�{x�К+�'6ݭ�Wdm�L<���r�(1�`�wd�����!;�����aӁ-X�U ������p��!5�#B�ӛ�˘�;ݯie��3����7�Ge�x�fhӱ��g̸7�����~�9ia����B��^�6�8!C�9�I��Zs|�vf�(��,c������O������JK�HS����6���b�>��mG�?,�;������{:��r�Gl)rF����r�L�*N�f��%���h3�vt��7�/e����W(�F��0���I����皖>z��]q3ue��h����{$�3�ɧ/�Pm{l9��X4�@�^�Z�:��_��^�@'�sB�w�*�Fh[^�Y0����r3��rRfs~��I��J%M�{�kh�m%��G��M�����`q�Y�*��e% �U��;
�%�n��8�2�����	�A�sa�Z�i+��]`��������Ch	����Ηs���8��P�X�<�8���O`���^Yz��ɺ����̞��Ϫ��3�)�<�N 𢫮 ��9R�<}1[��:b��wA h��
��}�(3�I'��*(I�S3^yn�uS{�;ͱ�x�sA �̣\_/})��)�&�-���͡�;��m��xj��N�i�y� �gյ-Ңԕ� @�P���	��4t���+��м�
�x�ZW�/S� ��4ɒ�p��\؃ �g
�Y��Q�"]_��`���]<��b��f䱶�,���>�����h�qUZ2I�F}z���	��k#3wa^�X�*�[$fZ���<����<c�� s��\s[����H�_އ�}�_ r�D��F`��j��_�놫����� �gf5�[�P�2��<�,�j�)�Ͼ���
��	ڐ�t�ĵ����4o����;��46CAi�����l3TO�@i�${���X9�|th�)��\}�X�A���>�g�!S��5A�U3MP�W��߱-�
��3��r��^8�{�O�Q�����J��"���O��TJ�n�*���áף��N,�u+�^�:��8*8�ٮg�!1��� �ѹN�{=G1���{�	���ҕ �TLb�:���W��1����@��:T�	�� �A|����^yK�	7 �W��� �k�+x�r�5�����	�K����>O�x�w�c�F�7�s�샅2ƃ��G��*���t@��pi�N	��M����U�{/\�A�'��a��h3\�ݫ�R��$��g���Щ���}'�l�杌��?H(N_�"��v��O7k��O��`�	��ƣ#�C����}�5���cgBb�P;�����[S4���C�~b�ich�0���N��y6H~ Z���s�W
�����ōbNS��}��}�mqi��N�3�g:���l^e@���M*1/�5~ʹ��3a�֟���F�ȏ�>�T6U���W*�7FX��K[ٵ��e7%RTپ�BW
^�u(�������KL��r��՛kXsZ��,��gg�G�Rb�l�=��%���M��VTeIv2��/���.�h�֎��Օ!v%���M�`��v�T��=K�94�FA�x*�Z�xI��"�*�U��y��Ҷᆌ�I&���������g��L�и���S�K���=����k�L5,V�a	~�*��,�<�j��@f!%"Z�Z��|)Q�L�6/��m��XAk:,�cO�t�*����j�}��%�-����2n�%	P��fYtk7r�>�m��i���j�#U )
�9��b�2�tȄ&6�(K��7��clr�Q:��f��	3A��
q��­$L���z[�E1��oB�)��,+A��MJj*���SQ�h��e�?�(q�D|��*�c�p8\3gq�r�(�"zF�;�$u\1�<,��G*Ϸ��;�<`k��
�ό�S'M��^^0�� ���"�����<z�]�U�b .�`���2c��h���t�z�m��r-+�h���u�/��Z��;�`����L��{
$�B��n6h�M��g�D3dU�9�͸��/4�ӛ(G�oG"p9�6p���p-7|�k�ۻt�Dk���U:���@uv
*�Y����U:`�����\_]�y'Ħ���/�����XS:Y4Oβ�+�����@:>G���n�X�?s@�����>�#�';7»]��km��V��,��ܜ�F�����JZY�.�;�����;з�t�����J��������(�7�E���7���i�OC
�K�#p#w�Ϭ"?��*���&�}R�c��<]X��__YҐu��t���U�b]�ǉъ꤭��77���N�W������
wS6��Ы��1��d���]s;�-���ڮ����$P#^�iV�W�C��W����zG�W��d�ȭQc���f>JJQ�P[Dſ�\�,�.��N�<��R����AZՄT�ܓ�Q���N�-���29 ��g�:�ob�Ͱ4�Y�َ�@�C7��:��=�\�U|@2!�w��h���<ȵ�z	ƦxE�|��r��m��O��.H��2�D�e��2�pP0pȎ���?��$�BS�2�8��T�J.;~��P\A�Cv���U+�Eԫl��ϗgc�ֱ�o�-�.�@|m���� ��-����^"�a�-�:9�Gz��n�O\�g�ѻ���Tj��w���bdB�'#�7Tb9��x��)�f���U㿄��ǳp���!_k�m@�%J��a�,%�$�v�^��f�[x�]�1�ɾ��B�������ɩ1\����V���I�~T��p�}e�F7lx�GH�r���Ay@3�Lg\���Q=L�,��UD�/ֵmQWP�'��UM�cs�	�TS�I��e�]������s�W3݂��-�1j���G{���}����vr'�o�#*t��[�Q��hN$��͖�(_e+�L2���p'�~/��M��y8�8xZ����'��z��������y!�ET܇�b�:θa�D���.�9�*��{^�~�w�n�	�@��n7�Tu.�g��[���V��;������Y�4u�آ�f�o	�a�,'┖�{V��3=�u���2R�,@{D���lU@���&L����hZǓ��!���y��S�Xo�d�m0&z-��M$6�8{z�]�hx�ڶ2u],q�2^$D���z��o�f��$H�m��>���ҏ+��/T�`�.�q4��Y�[E"��R4��Yk�l�J0��������P�2�����M�V$��W���8�	�h!��	{iz5��s:ῶ{i�̄;�>�&?��0I��H��#%d�-C�hZ�Rń����>�� I%o�n���8��":�D0���6"�~�ԽR�wz^"j�E��J��z�>�͊ש�s��(u�LJu�Q�=B�q���d�P�t�YNV�.<,Hr����L�bI�L�N��ր���bE'�� ���u��Ez�{�+��b�7��p�Օ%$[��ҷ����M`F2�����l^��2+ ӯ��>4R��0[$�8}BU?)����	�U���J�Ő�ږ�0���ݢ,�4�M�p�������5%���s�-A!��e�!�}�"��W"��b�t_��[�jw��։a_w��^y�h�qEiPe�6e��ye�c)mP����N���/A�D��<��q]�IJ�E�ь+���������2��apGw�����������c��������\�oB�p`Un������
b�]�g���	!�Gv�&��ݩLH�ϐ�O�G����{��طЛ,[�,g �V���;��U��=E�#��'����0���H��/�s�Ĝ_CÓ�9p���#��8"w帿9Эi��H��J>9b����s�˃aP�U���	ٮf�I����;#f<z�8Cy��؎�K��!E3���o�\L@��[Fe�e�\[�;�tH`��$��j���Pj�su�"6d���L��nC�΀���E*�.���|��:(i�
��kw�Jp ��Om`����Ͼg[Y�jX�u�-:��:~��� RSjߥ�낶�����?G���,���-I*�Q�<b:f̶X\��&GG��~�	!7Z��˗r�����,{�*[�b�|9B��=�1��ߣe�����A��2�R�1|!�_�Yr�J������ɉ�7�������$��탽�V�ʵc R=��c3�� u���Δ5.R�Ǧ�! ����	�=kn�!aK6�{��%���R+ܿ�xyҴ{`��y���0�.�݌V����ئ��61O�2�A�w���+��՝:�1'r�i����;��#Ox�f߭P��/�A��p�zc�(&̡�{1-��Z�Z�qn�@~���J^��@�����d���+��k��3��jm�x�:1�B�(Mս�f�y�����k�m���9��K�h ���6���2N�a'�.p]wuw�n��g{Ƥ�ٷ���H�-��^�ё�I[�F����?\�
Jn�u�y\Q?er@2���2Z\S�M__�O<^�.�D
��P�����F�5{�,_B�F�M�o,J�Y�?�VB�_�j�Yj έM,H}��q���]�`�`����tltڞb�Ch"W�s4�U'���<�h�ĸ=4ɧ�"�����&�7!���)��r���������N�H�ا���+�;6�H<��}��v�9���]t�7�
����.w��&�!�Sx�,2���������PD��
���������Vډ��J,d{R� �|G�d�7�:���p�6zx��,AP{a�z&���8,(�$�[��Ԙ�;S�����3�W��E'�­���SN��(?k�xυ?I�^��jb_��x����]�0���fn�;�1���,t���S�Ճ� *TmI�5&��C=�І.�#k����}��
K��#��L��zg��И��o k�RW�s��-D���1���<k�w���=G%v�oi���R������1E#�<e�W��t$ ����v�H�ށ�5<I�g�����RX�s���q�7�khB<n7�6k�XZ���rx��p�X�Km�d�w9Z7\F�)�-�(Jl�+�wZI��C5ҙ����ߍz�V�S�+�3׳����=���w��!w�' L�4����H�U���/�gr��JK��o��Jb�B[6Ч��3�������Yz�b�t牛%�6�e�߅�y��t�B9��- �l�������ISς 1ʗ%S�Fa�>[��Ϥ�8.Q	�6��m��bg��и+̲�1a��ΛtT81_�*��;�c����M
��9|��^��\g�DQ�#`1T����>}8c5\MW4x)rx G��pC��#e�K���0��|":�K��DH���̐ߓy�d��E�~�^6=�$�S��X�	�nz._�ҡ��!}<� J�t;���X���5����� Z��Z8�/��������w�k��|Y����X��/5�(��.������5�m�<L�x�(+	���� %��Z�߲�������L�r�5���R5&1��́��G6yٜ�V����D��`����ϐ�&Y���p-��Z��" +sxR�Inyq�'=�I��Z�W�{sу���y�V���'�R�����W���@�.6���E���S�=�s/c�C7Yq��\�&�᧰u;D$�vl���-�Br�Uj����n�(�hxܠW�3�����:a
q����ױS����g��Ė�3G3L+$f*e��䋴�{�õ* KE"��X�UJ洀�
6~Լ/���rO��s�Tt�� ;7vw���)�u���q_
�
���!������ ��Մ#�/�(`���Ib�a����&v8�U��)W�gǩF5#�x�|�ᡌ&)����}�Mj@�LY��
Y���럯�l�q��t����KX��b5��Ml+s�&r5�:M<'�#�CKO5�+DxU	�_������5ۇzK���h��nr�,l���7֝15w�\\��!ma�L��P����nM�mԆ´4 Ŧ=�4�Ӵ(ݮ��z�ݣ��NrF.���a�@<�Px�E?���=4;�=�db�t�-�H)m0���+L�\;t ��%��+;�3��ʫ����Z]����O�����<�w�c�U.^i�����$��QN.��*�����x���T�������#�s�lY�� h�h1��i��M�W��ݞ��v���PZ��Py+�>��D�! �W�3ΨT��s��a���x�+�lč�x#����UZ&>��߮��b��M~��GX3�*\�i	�	�ؽRQ	t�j�Y�0
�*�v��t=kq�Pv�����W��bM�8�"\[H"���1���̫t�B] Ŝ�@��xb�7bvL�nC�V��̿W!&�vn�����#� @B������.��Zl	���a�Q�%���x��	SH�3Z�788ڮ� u�3�Dck�����g������'�=��p;�"i�X���~P/�&�y|�==��br[cc�V��V���I^c��x|UQ5�ɬ6�`��+��(W��H� �I�ͻ��[��.��7zƇ��ή_<������r]^��.7���8���؀L���L���3��^$h�Zo@$~����J���N:Nǉq�k�tzB'��UF��~vF9T���E����.�~f�|�~F?��Y�S�G����P���I@��!~_P�X3�W�
K�vGQ-��(*���,\�����U&#�FT���w���M���@�H��Rp�}e�I���9�1:�kt$\�e܁�LYC������/¨?Ҏ ��G !0`��sw.i1�m��'U8y#g!�_o�2^�j��A�,_K+p��#8m���q����;~r��v�3�˚����i�u=�a f �i�A���Fx�m���f{W^�1��UR+R��z��_�ege��rɭ���X�����E^H�R9�?�ЄZ�D>u>\�Ĥ��2W�3ࠤ�Q:Ʃ�	S�8����ES�m�9��<���F��Q��#�5ȸ#�{H�
���Z�ڳ�Kz���p_#*/����54��Rjs�ީ��1%�O��0@�׍�_jcz��.�e���D�Q���h�E\�m�z�,�swGn����\[X{� ��2 �	}������[�4 �z�{�L�}˴u�T=���Fm�A�Z�Z�8�SBL�{�vD�XU6��M�`��#��o� �2�aS19�ŀֳ����+㻍�@[o����4zZ)�2VkX���$��"a��Mp�� ��+̩Bt�����b��(�����[�d��:��,�7���qO��W�^0�3���+VL:�[XRÿ��(�����g���Shq�i͍[�O"��v�c��WM�8�-XR�k����5xЂ�)���r��R%x`�%&�p��t���3_�]��Q�"25>i�bܘ�q��C��+"?��扱�ߖ%��戚d����sv���4<�Z%J�Z�����\�?^�:�C��TX��d �~XՆ�>����u;�8<<�g�
$���oU��Jp\�;���|!�0�~�ݰ��^��QE���֌����U�DD��}=F�-�(7~��lD������N��a��1��p�^)�\��LoFz3Z��T ���9�~�o+�@�q6؊d�J*xsR�ˊ��?@ׁ����q,
�������S$S�!��`b5�ÃkNC� �C�f���(�d�!���&�����`�.�xI���#)��Ю~�������\��X�9i->nޡF$�w'j�Y���f��,ts�p3���;�?Z�2�r���s{���rji��ٰ>΄��B�)J_�H�.&=�oS^ߜ;��[1�[���߅��r�Юrɵ��[��>䍙j��[u!{X9%��^���y���L:D��
��R�@&�9|,9A�vr��z�E^U���wh�[���'��
���f	g��0�wڼ<d��H�0T�9e�����m0������ �׿��|�Ʉ��T�>���Vp"l�B�P����0޴�U����@�o��9�:�W����[�@�9�hj-b���T.��xh��et�u��T.٬��'��Nq������ˇ _^���|S[u���S�ʙx�e9�_��� �w����&�����*_ :5���9N�4��2�a3��n��E�U�H�,j�R7o���d�k�A�*��4�3ဖ�`ƿr�#uf�7�_�l��[� 憨B��RW6,\0Mz`��2�A�K�Z���w�bp
dM�{�"l5��T~!"���iL⊑��V��3�lSaũ�<�k5� fX�ĭH9���������L+~A%�鲟=2r0p��gS�2|���µ��S��&�j���v҇�t��[D��F����Bi�綑���zO�i�T�4'g���΅�E�LG!<��LQF}	�B$M0�L����D'UI��+�v�2Qqu�V��Q��"�Q�Τ{;���j�@�)2[0��W��S%����Mxs0���iVEި�&7_�qi��ԇ��ĩ��יV.��^��l��|�y����%G�P��]����@H�-��Mf6M|�o��┝�7�Xe�����i.o6��[�8.ż?썗oț@۝�!Y{
�f�N2E$���u���~#*��c̊䴳L&��N�{*"	�b�~����b=�f<qAV���,�;�8���<������B۾gʎ��g����_�S��P~� O�Q8I����m�HU+M��6���>$�� B�ƽzBh��	�\�kK�(�M9DL��.�LCҎ��ϣ����ѻy�<�2���n׳(�^oyW��^j���5�(�����K�ʴ����Y�������b���L��>mh�|�}K~PmS�TĿ䲖8�n��f(�$�c5��Z�G��?�gT�Y����;��v���vVt��u�O2PC�sէ�
SL�c*ʵ��c�	����(;C@�.nXE��݉��F��ъ�>��#so%�|YC5vNHz��P�"_.���Ho)���*5�%1/�dŔ8,��`��g3���.TS	q0֜��iǱ�U7�����a�I|���t/��
��(at��n.��[E4�����c�%H��ƾ�+��}?�aY-���4�C'�ap
��p?��G�f�(~��3y�8��a�#���7���K�	q*+�5��^/2�B��7������}�-o�9b�5��t� �!�':Z�⻽�g Y�?_�7E� ���ӦD�I{�����)�`M+s�w�� �T ���<�=�m��pj�U�u�uRV���j��7cd�SH�tq�u+u����0(7�xpv��#Y'��2W���`�Ix	j.��ԟ��(�jx0�U˺YѾh�dn�%.�Y����+�#U��/�ģ4��WX�OF�YOa����e�Pp�����+�;�4�U���j�q�qRw}����a�!�����c�O�<yV2a��q.sK�����L���T����?�d�N"��Xeh��#�7p^��
S��t���gb���Jح+��qt~����`�%AF!u��}A�q�v��˨'1I���e��-?�8�P�%�4KT��X5�Z�����os]e�<բ�0��F�H�`�0Dժ6}����Z�Lڨ�%��9�}8�!�|�h���d�7�8Y2e=bR{�ɲ&��A�(�[�Ƿ��%���jm5�Y2��5ݠ�X��浈������%� ���۟s	���x��"�#��>�Q�E�M��z�(t�z�;��S�,2|�A��}T��4	�V���A�F�|������h�\���%�Q��N>�Ŷ�9	���{�{q���#7Xe���4^uRF�͎$dny(�W�)�b����&��d���leo[�I�?|����k��-G^O�V�Ō)ߺ��|%�Д�-��c����g9�2݈��L�e~�w��(@]��e2k+�#�Y��"��1%P ���ϧ"���թ�W�{�m�i=~��-�^�<TW�~*���į�Z��x'�遭���h�G�$��;��s�Hb����a�{��Zw��'�!�4Tr3x>����m`�E��Y��-,�~������c� hК��J��s���F������\�^J3j�Q��R�����= ��mO�64W:�0W�Y��3���{��8�`��Y*�1�&;�3��Pqu�5������^_����r6�ت����D~j��֛�`�MܳVb,��Z���PT�V&�ʼc�~��D��Ѣ	���s�}�{࿣�X��xm��f�/N����7զJ������+��_R����9���LS���X`�Ol�.��j�;z� z[gy�c�S����:v���;Ѡ�f���u%����e2�(TYk�d� o�4}�a��m�v&�b�,<滃�ēRJ��ł���7�n��o���cV���Tw��N�n&K��-}[���T�No�����p�%��̲�E��ѩ�iw�yt��BA9p�����3�J��c�(H�S~�7����Ъ���(�.�	���;VGl%���t).4,k�?�Yw+�s����ˠ��cɸ�В���*paT�NiV�^�d����n%�aRw��Ow5B���������>���=K]�K@ȧာS�D�U� tm̻I|x�Ɇ�eS�ėTr�Е�|�$�BI��%���/hDNH�I;t�ojW�ϲ��o��ht�c��D��\TG����@[����V�#���F��2ʿz�?`?[����so0�W-����+�6)k�	v����<X24:���G�)N��I���)A���� 4a#P���Z�.��V?�nO	��U���X4�y�p�}��n��+6B�X8}��r��b��C=u���VV�΄<j�V*.Ec���\��*�mp��[U�a�r�I�# �~[-�|�UXf�>��TAݖ�W@�I�ې��寘<ϳ`��E�$��k��9"+�v 3n�����/[����f�k��!��(�"E_�e�P��N�����1� }8�����) �O����F��b�'��;�:� �&O�`ɡQm��|�$�zc�����ޙ�5�E�s�ө�:Dx�*�
;�g��<�h��ã�Ӳ��m�Z5��~�=�H��X')Lw��o����T �կ0FB��GXi�d^7�,�	\{���23y�W�vF�F	� �2&�;SN���<�sy��� �#b����C�$�Ny��EBym�;�ǧ����h��[ֹh{�'����K�F�<�g��㬕����ͮs,�*G�;\a����UHџa���y~
����n�E 
 �&.n���1�tI��>{�Í6�t�.Xl��:����̫H˔U��}��(��\w���Q�~'�D�,�%R����`a#����z10��zX����1�w^՞F͹����NB���e�S�8��{��~|�
��0��v�^��ǄjP������\�B�Rz�R�9C��cZ����NL�Uӟ�<S�� *(;wl}���,�Ս0��/�qMwC�
n�%O����UE@�_���@����y���{]AnY1��"ӘS�^w�;�,}p;6�׵�$K\'�`MD��5����<�b
� �zq�#��!�e�ɧ��7�4��:��(tn�� �@+=?%-�MH���XhhY ���pi�՟dc"�:s�(���
Q���݄�S����(6�5U�}�҅�|�X���d�I9Q���j�꾵�,s��n#�/������X��4#��8�	� �d��#�J�Q��Vw��L�!x7����q|�@�PvL�4ޛ3٢{̟[��T
'��J�C���2��D/Ϯ����H@�2�<~2+sw�����[��K�zG�i�J��y y\�ǝe?�>�lc%���G_�r~p�ɚ@:D =�qó�M�����v�I��ɟT}�~�/��t��̢3^NT@ʃ�5�,AL�ۥ!�k����tGr��8&8%��$��P8lY
���=�<go?{�N�ͣ����w�;�*ݗQ>�JF䎩�+1�
-4���';nҮ�z1c|�E�ƣŨ�R�Y}X4���Yhݸ��՚��X�Tp[I��s��}������!�}�Z��J�)v�,B���ԆI̘>+s
7��tl��l!_��I:%�h��բ�O C	��}��4�W\t0�7�ES�'����Q��z;;�_;R8�S��b}S�55v̳_��Ρ�=�f��qOEc���[��&e7�ʫ%�/'	7>�H��������[�@@Ql�p�^?�tO�V�_;&��褞P2���Q��E0��N*��y_�H�t�э�!�VV���.����Q�\Z���Z�*��./�xx<��jwm�p�9���Fb�0`��f�
��:���K>�.MyA̧i:���t3`�ޘ�u�7v�.�%Y�C�+���"��a����򬀲�N�{r�}���U���֚\����'���꾕m��o{.�?���%�2��Sf�v�p�7��$��h�{'N�LůX��QgL<O���O���7������-�o}=�)��K�Y���\>����E�w+/�(����Q��K�f�|��s���=Ѐ+W�it��˛!�]��5��PBb#۬���W��&�y�$�N�޵�B�C�����♗%5��sR�)����3�����-D/9��5�
�q��S(��G�Qo_�XU�i�aA(��������w!�����M.+��O:3}��W� s��ɐ�Vz�	0u/$�-�D�ɰ���Z��Y&=ߤ�*�р������2�r�[��=((��O�� ��A|X����#ϔ�}<s�Jq�jOv�S~�J��` ��F�a�����\\��~�@��q�����Q�v��Dl2���.vC�����_��R=pᇡ)S�K�pT�&t!߷��h����'hs$�/�,]Ȧk��R��/Έ2L�m�)69u�^��/6��nc�Pɘ�4������~/�.�ti�2���[�X�% ����'��K�`�gb����c�X���3N���G-��D�ZILj��dg�RO����br_�~ n��e>!�j�&�6�Ÿ�5C����93&b�2���|>D�0�l{]:@�ɯ;}��K�����:�om!�2��f�?�*߃�:���X��ݯ�,��k��x���3�~����X?�~N(�C¿RǱ�-� �%	1�����*܎� �|��l���+�#:5��|�(�c�	��n�����q��x�U
"����o'�|���G����e�}��o���fԛn7���ܯ�X�7����-_ ]?M��Wޛ�Do{Y3/�d��t�|����ҷ/˄:��h!���HoCˇ�~���|�ޯf{q����\oL$��`��6����Ӭ�� �6�_x������_g������n��o��t8��n=��Ke
��%�9Wm�y �H)E�ű�.���y��I���R�֞6���վ��L=b�<�3y�j��K=X_|�kWY�-��M���]}ۧ��Ǵ�u��N����?�S#
�`��{znTJ
]vUUj�`�*��5�|�������K���-��+�}GS?�y�I�=��- ��]�<Dh�v�3*&�tKq�i�|~�� _�.�/>��f�0�y�-{'+i�?����;*	��eW��6�K�ŉ�len�˰�*�®�U��Ġct��i�bC�90[l�S16�9�m�Ն�q�k���io)o+�&�t��L�_�"Vb�>E6��$��؀|5gA�Dݠ�鵏��,y%�-��o��ҭ��*����Y�6/D���Xв\���X���q�{ԕ����"��:�H^孰�4U�4$��ؿD��XHX.�.�p�Щ����j�֑����u�!�fj͝]<���ͼ��r}XIq*s����Y����y@�%0R����ɀ-� M�\�%�0��U���v����o�@y��Z|zh�(�)�UA��Pܗow�y¤S^�?:_2V�+v����Gm�!�A06@J��x���}�/���
���1���ԫ���"�t����6�� ��G���"�G��k䟃݊�%3���ُZw]�h�m�,-��;���ڼ�%0� ��.��e��dͻI����?�����aɐy�V��ٽ����i�
G"��.V%I�	nۼ�)4��E�F�� O�h�k��=\�.���ɜ�C�od9�y��+\�0�0rM���Y�|�P�՜�s��D���MU �O+�":}?���m0���my�������F�)����?�����&��&P��(fs*ӏ�a8��b<!�M��&�|H;j���g��!;Vl�U�G'��Ƹ���Id�I�d��8�h�;�lm4�	�5��v��X�u@#��Ro�ćTC���ЈpoCC����g��Ȳ�U�pyJ��4[����w�R�K�t!��+�,5�ȣ�Y�o��.`�+K~�u�z�8+ʰ�����h_�ԣ�������u���Ξ���q Rv���8���DC�q�d��?��RP���ѭ�����	[�o}�Q�B�)����UF��TƐn�	���iksN5�9���D(�y8��x��a'OW��k?Mj��3�����?l?��3&�o�,���_C�:�G�ޘ����[�ك?jj���
!�:A�%ݵ�W^We#�����¡{��5gVR!r�QnmmB�"�̺��8d��04���X����5{S��1�a����0k�B����~�g$��s�;�@B���<����o���[�_rQ8j�s>�����D�Ѧ�ބ�-�֊�n��C�>�_�㟢k�|e�`,��tk*$^? [p�b\�YI�h��\m�����9�^�����zV�<�jL��%���rB�I$�T�tv��ܜ���x�m�dz�ێȍt�i||��^
��1}��{�uBE�s���M��is��n|xN���=�o���lp�&�[S/�������q��]"\�J���d��"t�i��&>��S}�E����x��c
p��hz�0a��e&�!�����h7��i9�u��y���O�Ŵ�u�gr���n��*�Pd�y�S��-�!q?�C<ЍE}"%����/�ηZ�XW�V��:�B��j�u��餙�"��CZ���_�����6�M0����C���:�d?}F�:q+���J�����?�}Tݾ��)
d�4�ׯ����N�>j�3����>D�z5z�+��U3{�ׅ�����n��)����Q�U��י����s{�Ӌ��� ����=N��T����(2���5bE��R"�Ǵ+
 �/:�#M;��O��4r�J5ؑ-I��+FBdGPг �&���P�oI�P�O��o�e��ϻ�-0��φ�q�X�����R��5O��z���/����E��YyR�=@���~*.z`��{�K��7d��s���y�KG���j
��^��8Xx��ۑM&��1�MKhx
SH����8�tV�=PV!�9�Vѳ�h[e\�ՓF�N2-7��\Eа��'Z^t����s��p`A�/�O����TO�H�)��On~ň��׃�v�J�j����Ȟ�-�J�L+`���E�e��m��j���b��C��^�u�L�ďI��]#����j;���,�0�a�#Κ�Ϳ �hp=�C�nr���@堔���'���)���\��#=���
߲��?�I��,�����Z.��`�&���'e[�������R�u�Rr��4EA�5�)t�*���q�R�a;�X��K����ty3�N)ؾ��5zLF�-�Rk��������(���b$6`�o�cW=̤�(�[� a�p��#P#P�����C�J��1v\�Os��~�*�>���6�����ZB ���xn[��A�DJ�j�E.�V��.7�VI��w�kP��^9�S2<B|���B�{(�f."FgjWx9I#��Cpʪ�� �ɸ��kj�Z�@e�w5N�g�l���B݊�5^����>��,J3���@^<�0��CJ�E�g���b<��t����P{��
��j�9�ő�1�N0zG~¶�ߧ���#pV���!F��-W>�}7����{�4����P<F�YƔ��+Ϲ��VY���H�]h��2�v.��|�v���7�T}l�ʃv䇀�q��҄U�f�2�4��6� ��)~�-=w1=P�@}�Q�)���LdR�}]�0еZ.�ީ��?��%�CJ�/�4����u*���@���/*|�I1�ܼ}��<"g���p;�^t�p�-׫��[m�%(�M�iпl�j�?L��?��k��;/6��&d���.���J�_
_�wE.5R<���ؤ��X6�o�g�GT�W?:�󢍾 	�ѹ#��UA��kt���K *�a�����v� ��;f��ԁp�����y���LD����O�Y��UUŀ����J��c!��M� ��k(%h�0��,�W�%�<���)ȇ��K�nX�#��[��	d��c5������KA�ʭ��W��]M�#��F\�wbi�� ��C\����ܦ��<��Or/�ҸDb�f�R�0,E��~I� u-* 0E�tv$�1��Pe����M*�A����~�ހ=�c�7sև/"
��U��s�<�v_ҽ�n��N̜�o@!χ?�=�wMQd&�C&���l��w��6Q	�Y �-�)���w�3m�7�lT(W,D�gL$����L��0�#k �:.,8��{�>����u_����r�)��)�z��3��|k���/���4̘���}J�C��:.��VW��Q��2��毀�����a5���������-�	��Ͱ�m)��ڋ�����ݛ㐞��~8��ebf1y�bR���MT~�2�DQJ5���㌴. dt?��\nu~T�7���������ER����5-)��-m��8\�����kkP�g@dϝnyf<Z官e�Qd��p��&Z�4�,K�rϋ��k�������ϸ@��
���j҂^�W��H1��\d�yF��k�I�;��+�=}�e�9�)MAN�HRZ�Ϥ�5OEg�U�tw@�w��`����N����N>*�$˙�>aVr��(��Mt��3\{�q�����Ն��΍_���A�{ֱ�dK�d��|�)�6@��'S{��T��6�z\}B����l�|�.և�Qk��5�xu$=\hd�&/�`N*l�U6���G�っtQ��ߥ�ҵ,֍	J�6np�R/��V%/���ce��ֵ�n�m�v2�{y��m�lI#t4Ȉ6�N���(�L+%bpb������*9#�Nh:�1��d�L��~�!dL�?��@� G���%�h�V<��x��Zo��(�a✄����`��8��>��p	� `b�2Qױ�_����̤�PC1	�&�~}�/F #���I�	��c����}���>'�6����}�N��q��T���1Hd=_7�]�a��J�����6��P�?�9]��TpF�0��YR�o�u+A���hf�+v�qEuai�8<�F#�gɮ��֮fw���T����/"'���AJm�˪,�4�����XY?��`�EAe��z���R18��b�Ʌ�dȪ��}x#�b�g�� �qf��[<[IHZk*���6��V��#4���gQ߿�2^�#e�Ju�t�e�SfU�����yC�<�m	������=�ڍ���#'c�ꢑ��ݮ�S��/��o�:MlT__����Qpn�E
�)�<�BK�T�PC�w��p�EAΞ', �W����c)MW�H{5����x<�}�2�w6����XWѰO�� ]��ĺv���i���9�-R��Gy��wԃ���A��Z��YpvtV��d���g�M܆Z�_�K�zv@�d�M�(�\��D\S&���$+�� ��l���o<-�๕�Ck�;껪=�}�Qg*kᦗS+���z�!o?�I����D� OXy/�s]E�z�|��@�]�Y�8�(c{�[�W������%�w�J���^D4R]�C�1��Gl�L.�%��RL�8D��h$T���~��wL|���eu1w�36.y��ccz��?oچ�Z�'���	w潥�[��x|}��@0�$`8Nc}\��2�J2�Áڳβو���f��>sD��I��$	T^y��[V
:� �b�cs�NZk�����7
9�F3��C9��W���yO,��*�N�=�c����o�g��+5�6���9�<�0�[�@��$�*Y�W���E�q�q�2;.��AX�����^�_$ë��n�?�vYפ:3���paK6R&�4�,����Σ�\����;x�72 =�o��k�m�dF�'3x�����H�2i��|N����7�]�f6���`/�
vɚu Jٿ���LQ�4��:r@�Zb�]s b��!��k��� �EVJ�Z���Py~%R,t�&�Uĉ|Mhz+~j (�ȭ����>��0��Z�- �h��Z��:8S�r��a�Ӳ��n�K6+��i�����}�dy�~h�4$ܞ�׳�^.&ۜ�tq����f�rIǕI����֌�鯛����Ѭ��xp����u+g[�(���b�3T^AY����W�����P�V�km�7�w@{�kw��c=�{4�|������X\?|���.<��}�ߔ�q��A�q&e�Ÿb��-����#1u���2���k�@��sf�[���T��V	�
G&ʎ;4�#�+�?�X|#��$��N���Y
�_��N,ou�0�8����ytk���j�� �E,��M�CrrW�d�տ
�1�n�_�)�q�7�)�
�/R&�O�ܔ>v�vPmĳ��t}7��;�@���Qw�3OKq �6�]ҊR�'Q�[T`Gs���ч�;-^��T��W���'���8<h#�+6�����k�x ��u+{gJ��4�^2���h�w�$i�\b�
�'��3��*sZ!�w����f�5��%������3���߳"���js���J hc�@i��q�i%+�;�>��M���j��L���E�Fc}�M�>e���5Y��W�.���0��ő��[�]S�lʻgO����5���r��i6#����Q���o��?f�KJV<F�_G{����9e �>���Z�r&�+R�ք%�h��Se`�51"�i�#W�s�1��g��g~�Xx�=+��>l� Nc��C����-���x�ꓯ�A���
�ʸz�̈mS��SYx�)���*^�V*Wa#�� �*��^�@���%������\�
�6N����;�'�_U�I��k�N�9��L�A'����X���V�N��5f~�R�	i���%�x���i��ppA���ә���c�(�`g#�p`Ӳ�^.��o}F�?Н0!�i���f�Ŷ�]d���!t�� ���`�����\������֭I���I;Y��~c��]�d��[yZ�,.�/�Ɏz|ͭB�T~%O�n7a
���o�z!��g�P�ʋ�"h{|P�S+�驈%�^������t���~<�θ뵏�J65��K^wG���H����� K�xG(w��O�t����%��i�=�2bG�n�5����`�wq]�L��XX��5;�<���$��;<��0�ߜ�@�~~^�5�-�s���?nD�}�i�˯\�[�4S;�D�+7�i44��m�xX�oh���*M�����/_岔���Z�v�Jfʑ�~Fw�&�����{��9ͥv�Vdƣ3�w1����I�$	i@��t��vU��Ԫ�dV��n#���;Zb��-ef��-o����]UC���:�n��Drz�n$�G̮�~M��\��Z@�"�/7��pLR͉�l�;��|:j�(y:�p�Te9�i5Y��-WG]�!L:?��*C}�_�&r�A�G�&�QѢ��<4����rJI��bw˺E�e��231��t3�L�ԲV0�;��ed�� >��
f�`�Eh$o�@>.r���m��Ӳn�ѸL���f�b��Yk
q����H��T��- S!��A�3�=�=�@u�6@E��	1UY���^��SS}�Ekr���5�(¤O���'�g�k,M���m�%��{6/�wUW6������)c)<W��P�����1<�F=�:��3�H�O0�8]y0W�/�W���i�=;�۠��((�Ë��r녎s�roC�*ub�=�eDp��%S$TZ�?V����oO�p�i�kW!C���^�З���?�-�5�.�Pu�Y���͋Si�{�L|>K���`�sQ, ��T�a�K 7�ɼ��r�g?�"E<*�`|����q�B֕��@m�Mp�2�Ί7��k�Ι�x<Og �P�΅� ��q�����>Gm�5[Pل�N%O����"�|��?&w�|5`��Z2;�U{qο�_F/�����+}�@��ڃN�
����ZK��֔P�W�̏*|`�0���.�h��U���Z�O�4'�T��l:z���J㡼��ceq�1"~��2��g/���0�|P�}�;��*p�%�/�&0a|u&�p��<���48��ȯ�u5n�n���͉a���}��t�T����%�9.^u�J[�MA/չ5��t��~j�F�T���Mzu�8õ�'6��Z#���9�O��m13� Ǩ jxw��ѕO,W����*������r�Y��9
*���?�N�(L?�K8�9�r�G��Ǽ���gע��,.�\�`F�:����ϗ���馛�t�b�!�;by�j]��yc��%tq%�ٿDK9w�q���5>P�i�(�"�Q�ҭQi�4>&������S�:������e�u�Ķ������U�7�Q���F��myH�(���h� �>��d��Ώ�@��Ln~sU~9�p�lU���7���X�d䛍���%��Y�S�L��2s�Cޕ\�/��ʼ-�:�)P�?�_��F��7v�u�(��-�92�^�߬%��֕��;P���UyF�ꑷ�q��0[4�ʁ�<�-c�O6������̏e����i`�K��x�~�)e#�{�j^h�n=^�Nb&����x�Ia6�8R!�UF�(��f�B-�W7u]=}�ܠF�q���w។�||���}�O�FD�� ��X�Ǒ�}3�jn�!�M�a9荰TUڮ�\��F{&�ĝ]n"8�1|���1��������wK+~NB60d��6�zw~�R�V��?��/pi�r"d;���{m/F!�C+xDo1n7T�.M�:�L�(����~��3�b0�4���ŧ@f�8�$"�}C�
�9�r�� U��O��)��Ԩ����p[r�[!]L���m�X���"��7�����N+�]�:��-_�7��7�Ͱ�]a�'Lg*��}S��&�͟��w� �c]n�ʀ,��Ǌ�)D[<�z���#�JU���o~ޜ/�ɩaݗI��9�ґ���� Ç�T���?2l����d��2�BSzo�0qf�ڵ��M�+p�ٲ��ܯl�5����#�Q?Ԑ]�7����I5OG��OO��������ߜ]	(P>E�����<G��6�Z<�/9I���SQ��q²g�ZmЮӱΕGI�"��Q`K
��9�!����^ꖠiv��Vn(�>���ۺ�Ob��x�=�2�!~� =Ge+���vx?g*)�*�zbt�=$�T����V'N�@u��Å��`�NoĎ)i�5b�Y�l�tX��=�P�F�Q=mǍ,�����f�L���߯5��B��A*����g�ׁ���r0#�POSb󴟌߱AY&w�30�FI�k"��i=��O�I�@�d�v��=~op`剫�s��)���gE�xx�ƌ��ɠ~�r�����L!o���)��ٌ/p= ��_K�ܺ���d7�1*-i���
q>����h����	��R��~�Z"���S�����	V\_u3(>@�v�!�/l}�)ߌqԷ�Ylc��^S�:�M�,��A��#gVS<>��*'�C{����s�q��8�{(�w	�{�V��DVm���V��z<A������p��u;��pDS��y�rs��W9��Le9�q,��+37 v3�`����-�x3]*W�~xDF�m.}a�?�baY��2L���:�>���n2�m/���xYD��>���.*Mx���s~�:�N�*�I5���`C����#��'�	��X[���*��p�z��F8����>F�*UZH1��7��p5>���"�`�-Y����*�aQ���J��/�����H6�m4�Ov���ř�pk���浥u"���ߗ�;=�B ��/A�ș���y��KG�o0E�_&��%Њ��F���0��
� \ �NDkZ5w�x
���e�_f\������a���yOQ?��Y�+iU����L���ݐ�@!	�B7��(��d�-�cʰ/��M]Q�c�p���7��������1�Ct�>Ky�S�/������)��:���Et&�tK�7�5yǷL�cj��ΐ'�*�/�y��r�oĎ>��'�l&�&l�1��q|r�LQ`�+��U�:�%��h�x�VxMbT; 5�aNם�<Ej��#��K�?v�c�$�W���o�ڼ�츍a�4���������,_���@�q`︹*?�������h�R�����)����t��N��!Fὒ�}�m����_r�g��/�:��~�|_�tn�=����K�������]L�w����Eb���O��7�zg�n�����؀
��k����J�ĕ.�}�]�<��ȼh�������2�k$H@;9��V5��N��ŵ�H�Z���X�}�&��I)�4�Ũڦ¹Ai��ͦ�;�� ���2#��U�$��M����2�?���k'cѤ���=��=��nf#x*���Om������Z�?�M\�v�_��L��hd;��C���6����Za�lˌ����.K�AP�����D��#R���հ����v�L���9E��^(��dɚ���JQSh��7�K��n��g�Ϋ�N��f���Zf��<g�����~i�޺$0�� ���ޥ9LY��,��޷z�����Sk��e<c��yzl�`K�D��(��u�����-gq��~mcڊ�����3��Z
���$��Jy�-�X�c&�5��6O/����H���#>������?S6�$ω|�;=��?����]U�������t&ԭ�sg˴�D	���8� ���n ��������|�ӄiz�N�����|.��/��Ǚ�YN][��y{����1�a,��A2e+�tJۢ&����ZLp��_��t��C�FQL�imL�������a�����JA�h5j�4�gȎ&����7�Cl쿨�M��>�����y��f���DG%5}Pee�?`HsJ��S�b����n��-V'e��v8����ܯ��$_��r�`I���oŉ�|J��n㢨cܦ� v3�ꁜks0�^E(S�����%��p=ɺ�s����G5��0z�q_�� ;�9*9�
���;;��^R�u���3t=\zs�U�	x�"���ɜY�����y��f
0w[䏐����ym�lӯ\����*5�Q����6B4�k����}���a��w�q B�����&�R�Azp�HB7������j|����i� � � ]�J��疋�nTpɬN�1��$ǆ���Jf�?z�>>��yH�}k�bDL#�׫
�_
����-�����L�d9V���p�/l5_F����t� f�k�����G�j�"c-��ޅ|�_��
����M�C靻+N���)im�c���L����EY��~qﺱ�������N�P-���� ����Ĩ_dļl�����(� d����O/b���T ��r>XJ6~�i�
#,H�p���lQ�)��(��*�Q�� �t����>���$k�?.2��>�'K`9�=���#������խ�?�P/
�|��ݟ.�7K�,9J)@�D1a�f[p_N��UkВ���q�L��Jԅ��{��Sk+�+'l��M��҇��?�Q΅��_����w�-��]tTN_i��\ߞǾ#svw�`ڈ���̲`��]�hJ��}v�)�_U�:*�i���I9��ҰԸ>�:�,�!6gA�-�+�����5����l 5c�
΢���-:4��d��TIj-KF�Mn�coj�&�$��GLʜ[ �x�쀏2��d�Ý����#������2���7?�)z-�'��lB���]���N9H�7�Qh��+��^��]�� ��D.
k2f������	`����7��X��\����섴A~M�^{��41�|��?��(��I�_��	@������	����֌�0�����M�up��g����φLsX4	xS����kO���(�6rK�S�pڨّ�B��D�VF��M�G��=mԻ��j�mU���9���H�3-���r�*�S��I�e�	��*���ۋ�	�'םQȪ��"6�\����hz�<ԛ�~����&�bS�7~rb��Ө-����)��L�CJ!����=�L �S��-ҽ�M�)��x��5o@m���T�Z5n�6�yt@��La_(��-O��\2�?\��^#��-[�̪:P$뛃��2�\'At�`����FpJC�'�R���D��d7J��g��m#`7��!_�n��݃ܺ�A�a�k��)�L�͑�&.�%�� 4�w^�V�"��bO��i�D�
*��=�&�U����Չ��Чy�?G�	exHx�a� qN�̚����B�@!B���+h�#�n�}�	3�; W��{C���~׬�����'�!�+N���8J)3��fPj%aK�.�񍌺�Z)��8��i������`%(Z4�yŉ�s���6��CDAeJky�ؕ�~�A�������R�j��Β%���T�BYd�So[#]�R�z^�S�v�u��J[Q4��������Z�My��љ�v9n�����哧)�T��W;�f�"�Lr��W��BZ5�!�0y�6�rU!l,r����ޮC�-�,f����]엦�AA��ꊒ�.�u���ڲK��80O?L�y1:(��c���b5��Ce"���6��5��f�e����y��~r�Ѐ�=L��	�P��s kt��_�ȯ%Pиg4���\������J� S"��ro���_�o���Uʈm"�/���_�Fj۽�0?@9
�]�[�{X�fn�F��\>�X�W�����l&� eԱ&�6���CW*��w�D��9�O0f��@q|!��Ӯ}�{��|���䟹^��K帬�R�,��DX~��Bֆ��lۢ��T|=��\�6}�7���,�J�ݣ��ʌCP�}�^a�9�X�6�~���İ�\C��j�ҾnS������$�P�m����[wVJ
A���Ɖ�&)/1䋥�=�p�j-���6'\�����m �P�KZ[�����n�ޱ=��ζ�hq6�=�IM�C�������6�9���Xng����6Q��'�G>o��(E&!���q���e,�`6��b�x����O���O�!���V�T�/è�$��ԉ#���e�y��гC8Eu����ͯG!�RhU����YlT���s�wi����'߾�O6۷�2��Hq*aY����g�B�궽DCc[�/�/�Ve}�#�L���W����zFT	�\��,��Y���	ή�i&���Y��M���F��f{���G>$pN�ި�� )>K��~a@L�S3ݶ�-�Mu�P�-����F<HDˣv��8&m般��f��F]nk�n��MN����W��,��A��`�͡�� t������Ó �yR������V�tg����X�l�3�rf̍��-qb�<��$�3I��M8�H��	������U+����_z����n=I��ƅ0�U+`�y�s/�����G.':�p|���g��;��qbo5ʅm���`����Q��P�*:�F�?+�;���cp$
W,�P8��t��:<A�8Dy�OW��6�9ҜI0:�r���z�y�Շ(�4ԝj�r�m�(&R�x&�w4���}3�?���=��<�Ӑ�5�i�հ��5��F|����7��� K��U��b��w�m���_؉�f�&:�l+0�� ��l-rL(*m�<ޯ^�5m��/x�|YnU�{���Lh������^�irx`?�^u���g�MĶt�ǯ�,�yk ��������$pqw��j�D�?�	��B
�7���tv�=�6N�C��_uپB����D	Sa������� �L�{�Q���GM^'��b<ۭب������"c�9g�P��Q��gN����k�';Y�W^KH4߈3��C�����s��9�~�5uV�-O���1��7��7��xP���9�տq2�Ө�;�w#�O�k �g�.��^u�tm�u�ɖq#�B�6��EA,z������±,�`Q� mM�S��.#��W�""��1�������������Ӑ��k�xv�\��q/?���,F�㢓�#�I�gP=��)-�� -�l�J�N�7�˸�6�S,�n�=��Ɩ����YI���t\��@Oe,�)�w)z�1��o��q���|˂�y�z/���>�|���ԥ3�~r6�ߗ��[`�~)���v+��Xag��7b��t�!�5m#ZV��n�ǧ�W�Ǥf7D��]��z��j%Vm�Ra��V�����H4��#إ�����k.�&5�.@nյ���XaOD�^��\�m�Cm��+�es�h�u-ݪ���M����LexRփ��]Н�0|������j9V�Ɔ�.=���$�O�7����Y��
v���L��}/c�X=د[/p�A��~?/O�U�d�!�1�ə�,�I%s��B��: Nop��w��v�|�̷̌�#��q���w���w�֋��w���$^�9�[XO�)�t�Ơ��M�*����A���BH�A�n
��`�^:���+q���;�I�VPߕZ�]�Z�ϫ�U��f��L]�,��Bt��Al#�g��̎8����yd�����}j�������z/�y�[�yK���̍�q49�E3��S�[��6�2�Ae&j1<z�͈)EyCa*�]6��.`2�@�;���׫�xrn]3f��W��z�ŕE4�;9����S���k,?jXv���F�v�|��I��c��ϊ��X�"f�94����B�m����?�� 86���~\ �O4D���RV���n��:�g�������pY��"��,���*	����֤`4Sؖ�����W�=��bp�2��Wݭ����;b�ͩp��Ч�qrś:��ӈ~��6�{����Q��m�a$��r��˪��qW�נ�lZHmLj��\��)���=�1�����r��֠x��x�۪���8���:	���3�����D���Y����$��[�R����/������M�m �K�3�y���_.~RO�.y��)�x��j��C�nUqm�6���5B�3��)A�/�*�~Yr	g�6��^�o���BLQJ��񵿱�C�A��+d�eb��<Z��-�xF�NMn!���;�1��:��e��l�.�Y����L�r>�)�WD�	X�WO�%����X9ޣ/!��!�Q/����q��m�CK�ޤ��ҋV�<��H���sD��oF�U�K�;5��-f�'Z�0�p�C�eb>eg:�W�Y�$�q�S�Z�D���� d��v�az�{�LB���o��iw��@b?Y����ǩ�V�NPW��nf_��>��d��J�KH��.rF�(�IG�>V1�2m�a�e�r�s&,�f3B$��0��{�3s#-�;�9�@�[s'�s��Q��/1wo4@ہ��@܋�0Ó/8��T
/t�޿�oVc�U���;\q�q��O
`�x����N�QY:�ɂ�4�f�u��