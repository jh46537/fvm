��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���ymc����#��בsb]b�k������w���A8dbҪ�;c���Bh�5u��):������P�Й��w�V�y��Y��&z1-�m�W3~��;7&�]ދ�Nrh�dd������q`��^%�2����/!t��y��U����uU;�G��R�|��+L��!L�&�����t��E�TC/��	iA:���M&)ኰ�P���MOA�R#jfz�r�V�r��>�u9�����g�D<������ws~�Q�	��	���P��sq���a���+���U��.zXu�a �P�<J�|�H���ɻ�i��h��n��vS������އ_�.鲌vz��K�a@�M��H�^�sW��a�E������W�b=e����=��:����M��"r�T���6�%h2���+�>.��\�G�)^����3QF�X�3����P���Em�\���W�da�a���D�L�&(��^�#�f6>�ɱ~�w�N�����	-׆L=
5�X�+dZM��-2�J[�B�P��Ƥ'�� @㿂�1�y,�0���c��FhZ��n��x`DW?���`���E{�;� ��Ze�����=N�V���`�}��rG�//�F�
������G-�I�I�0���JNY!ܖ�]�7���ڴ��D"�ir���!�B��*wQzp�h���4|���x�:��5��E(^��L|^&����P���Y�r/&�+��	�TN�C�s2Q��sHӟ �����GG�T�Q��B��h~/���0��ж�c;I������[6�=��)� ����{�n�-��x����x-�pg-ހ�������U/���`�<n��h�K�N㊠&8�����)�p!S�0������ЈZ�t�WAQ팰��'g���%>xd�e���Ry���$
k������1��2G"E L�v1ն���\�:��%�wFB���1�P	3������|�f*֥���	�C�G,�`�lO.���ip.�gL
8��t{F�{nD�	$���CL���4�� �Sw4p��N[��dV�:a��IQ����8��^�Qˋ��}!}a_��S>q�禍�O�rѓ����%�����*��[��C��^*�n�c#(�`\��0�P;�j֋v�0o����Y���>Ӂ�yx���$�Q|�V:ӯ���e3�L!��M�p�hC�8�w
D�,h��H��YF��ǽwm�i�n���K�sij
�害�G4SF��Z֍���m��$��~�	��Y��#��t�߲Ze��u�˓w೼s;���*��OH�w�@���~���=��۪䞵k٤���B��G�iT�B� ��}�T�LDl~������[Ϯ'�;9�����daןK���X2}��� Z�\(P�急�b����9��#*���b�`��ϒ3y8�ڲ^*7����,������	7�7��<�8���%��
�ιm�(��X�k�RƱ�vB�>��;P���X8��3JPn		</d�6��Ti�J߿ 0t�N�ؤV��T���[)�@�<~{�װ&���[r���&-��]Pmgcj]�m��V�5e������&qYG�=�{	�φM�*.���?�&!m]3��l�[��C^׬������I��l"���5���?��ZC