// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KMTZcPu1W+Jk4wGJFL+G5fQUHOlgh38PaFtW3/aij0wnct27QDtBs9QXak7v5U7F
1OXBty8qDQ3dhfmJSmy4xBrcxkXalOA1O5zfnok77qYfQdvotD8pf3WRlXs/uNX6
Mebv+X/8hpleZERubKn6ei5GIa2uADSB63AULrIuST8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11424)
8P4/xIfRUEw9/NkRq9LXz1Bn3e5Sa1TXjDP1yl3CR/4F/ANXBEL6FVXreBYhy5BO
Y4XRM5h6AzXXxWS5EiHppkH0b1puRVDy4pjXRVgjai6SeS0QIL/Re6hGzNpFCn+q
ntmBYVjgS0iIOLheLdMZ8qTyXAkefuUnoY3Qsx158bdOSg0+WTBsjrykAVY2MFQG
q8kym7yir6Cx9ATf7gwU2v4HJDmlqtCcD7Z7b9Fn2iSJ6T9Zt4CtehedGu0G1m4A
a/csAq49VlvF2OP5SM0eW6Lp0pUxwxakVK5p7IFEYfL5u0A6TRZODPNhhe8/RsuE
GuFqZoX4KbIFClLrCYy831/2c3zsPsLKa8jBzdte62IXTu0j1bdAyjhil0Zg+dwT
GBW5Qe/LqNzUT/XfdQKuK3omksxcpt3ga0ugaIG+JyQUxesFfJP2DIFEbB8mMUOn
LuP8dmWHoXIGWSIR+Sfsf2XsCG+aNijzDmyT0TP2iEZnIVDLUiVk1P45JkV4PW5B
M3jCCNZSN1QfJtnCLBh6Cl23BW0kf/jux6K1k2mcLeisT9nDc0FOsESDNjdTQcvO
9iTrUYKhfYDLpfG+FQ7erYYMT76rnxduQg1RRU5jrWrHTZY8WjDuBipVQUJdVl7i
5McCPIYiinToIgIeFrz+tAkNOLZgLRAIRYcicWA/zRNMqfE8SkdIYWiS2ysjaDxm
ntcehFM8c0HRd6e1TGvEKZDBGW38Uku1pOjT5YgTwHdtoa2oN/0lgCCIVtQK2j0u
XU4u8G1nlUBZIR+2n/daa1UpoSpXLibl5iSZ8DCMKfDAI6VcEWPJYEIZy2V3Puoa
QIRFTsn3hyF9K4EuAw15X/XEKdojRRipeDQrQBDAqnk9qZnaEXUd6p/z7tGcrO5T
XIimpVKeLjoEGVAyqhSJXEFO5gfQBrwqNEzBu39MaLvWl3B6mC5ycGTA+u8y3m2E
qlMbHFBBrfB7eDUmVVQ4EbanaxRquz0oHEvztosOHCENwJ14aNObOfGfpfPkCAlp
ggGM9nnMFHYnS82GiQo7dScA/URkUveOm5zLN4zZlVn4WNpJSALRYZ8RKAv1S0Br
vTCjiW7RwlElejL4nH8rNrcRzR6qwXnXtCxtZh+yoev8Qe0eAVUgk4sUg4a5bQrD
ARQVgJoAUoZlcdkPy2Cmd1cGxHIM2hHNGiP3Z+rPY28yAH1GPWNLkC48PZqFbPlc
w85ixoSCIcL9Rsr1SREzyS+lqE0rK9VHxnTVd+jXlMHoI/g2GPayVxQST48OTTc/
Jk6kvZM1AcbscSgE+NaYozssSYspFlW4mSmN5zoK8J+zwox/ZwmQDGjXVy2iAc8A
eJ8ENA90OkklbmjJA9o7ihRyyFlpa0om+cnxQYp39Rugvcf8rcyN4WtHxhrbZhQu
07xXjH4Mfq4p4syDSj8y+0kLIUdScVkdy9DMelHLWCfsuMX7WwKViv7pJ2QGTQOK
vv0dvWDFxE1GcJw+vZqby9hHfUHeG13bU5f170tpjpIMSmrSh0UYhaLBjhURshiG
UdNr29FaML92fh/1iNRmll2sGni4WRQrCMtZZTrgoK8FSOEvevNM/rDRC+/b4tvb
XoslsZ2TSCN/WplK+2PSLzSJ1pIyrT6Wvucs75BK+8r7NfxD1q/SNSp7fv8+Yc2H
sW6z+VXq3AVGdXApCf0RfZbDWlC+pqG1+zspq5ECfrMw4+KOiwP654+OItxJYnPR
Zbok5ZtUL+rj5FZeMYFzh58zd9Rh7Ms3kYjOD3BBpnCyvkBfJympWpZqf8hsj30l
BXPKsMM7kv7i5v2zkiDC3cGo8FORO7wwQ+yMe4jk9S9uTaL/IH5lJzc0PsKS9y9x
NAGBLANlGZcrHAqg/GD9ncRZK7GkXKXbbSeVaHKK0+SiJ0SfRaKnnyR6yQ26duq2
38hHuS5jl52QN+LRRCr3OyvHFiBa7o03RC+YAx/d0QVbA6QrjgmBh99rHsnQcZ3Z
QQIe9IWK5MaaSbknuGIFTHX9VkT/KOZ50XvIUXI3qiDacEmAWyS2TZuCnRqhnl6G
gS6r6S5/T6LxFGYyUdq2o4ISOt8Jbs1thandnlA2D1UHohtIcSGSmk53f1rH92NH
e66JJWgP+9M+KZ/kkQyAVYhU92Iut1wqhH8AEedb18hJMbPmSy2/BSJNthEsJkZp
Z9iXx4TVqiC4yFfkjQvIu/shqgPq8HKLGqEw7QS/ySVqbF6lVI95ivI4oruyGOAD
6MWs/uHN3ZVLyVZeCnaajTK+yLhQTQipH7Qcv2or2GU4nLUrXu9asCjAZIYZ8Os4
GSSE+6mOo+gCtaBUPo4LPISBaFL3/eQECUcOl6ti/qYrWpZ+l0e6kGEtpyVv9bB7
fZLhqe0l+V3tsh7oD9zkZ6K3drez4SAoLcjwzMCV3ix8HaR4rcj439QlityCbgzQ
hmxXxdaAeK49CMPju/UyDyE4ONoF2nVFSIZAPhG1iHleldHg0DPgJX8SqZDBEobT
nTdkeYHtLfEuvnJtW4ZxEQWVt1dk74L/JJtYavGD5YLzlfelLl70grhc4pfQs53l
MjLu4OoAHkdUWqHqBP4KkhByp5kdcZBpw0ElsL79hR++1fp/1CFxlrWBQOJ1Kh4A
G7xSFrFWxTH9/+/H1xKNuhbyNIF5bDF488uDmJ+mXnjpVR8s1HtB5y4x5me6P2Ra
k99vXO7FaurA288ITTAv2bMglC8mNNJO1teC3XRl6oKgnMnPSC4Qjci7uVeaLxVr
H1QYrrTA/gPfSXqeVGewUPEu4YqydXWlAT5rzDqHyLMTrjXiOYucdK5FRCeqlpV/
IPFkAn/ixy9o5UBSBIliEi7WKlU0ttCZrwd36FSOqY5UfTXiaIfHuXpqrGooiOoW
3gUknD6WEzbdP2px6T4VuJebV5hAudstsukNj3madJICVZwwVZS2PAwjSie6JmP5
Gx4d6y86dIl5FEDU6w0L3vWiBcj1Hqgi9Y6gxgNdN+J5RKG29vz57dxfuyXBwtf1
MrAodLUxvbxPGmF9qSA6hus4UXaDA+GEuJl+9/cmLnmEI+Kp7KV4K52wMeKxjKva
7qK9nHXiLPLttlGMf/d+T1Tx8zJ2RGksuCmlw8Wwkzj+CK9w5Kf6bXf3Hsg1pmHC
XKa78ANwu0paSEnBXMZQsTe71+kMreQOAZv1L18Cu2FvJ+d4tm24B3LDwZtci8/4
bZLVQjkrYuExxA1hPBCMBOSHrCJQZ6aMNydTWJ3tX0qhXwYH4Mhd2hAcYNGn5YJZ
ADkhM/eKZzA+ymfJdvWlYBC6gLUVtu/6qoQdKZbf8sSEy1PvqprZOlh6E4JtwhQl
LwD23nDgzqpF8lRWNKoxZg4JMqqlrBGa+Ila9Qo55fkeoYt2WNFfvIJrGT/YFxOm
jg4bMaXULwLt8clVu/djveV25K7aEXeNaAfkFc0Yelv4aNOgGhTWR2A9X2yTk65u
ziIlfhATKUSBaY8tFhxzmqnO/XWAPNgRMfkKfZkEBv4v6dbNeKIM+yMcpZPexswo
D4omkGCS9F+5RCeo9QD5SCwee70VU+3fYwVKjVYjMbM22UrbVkEaQVo7T7xFxxPc
rumbWkuyq8aCg2JVjVv41+p5T9rmJ6L7tgAHKF5nQjhqSvcW5FvaVtIsMmPpFeHX
W6ehxXCM5aRVJ82/MLOe+M0dJtcXYZMz1vJ2kurzKc192PxlKJ1uDfLXaVBUL0kA
505eALghUF0sLufBNompCco3p2J1zqJNxdtpllKz9k1pL36LqiytSYNvNUSTFzqt
2YxGWpkYIqYwXgeUCUJC1xemz2Rxv30azd4Wl/H27zfOa6TsYbd3LgxXsW5RSZPt
3bOzBKFsd27J8EEFsUsbdSROAE4sWtC/SHNYkY3Jwon1ablkdYtoLBXtNxIjQzcM
q5YTJzLgNbl13K+Wto01FC70RPuqvSisd2CU+c8M1LM4mYLjkkehitxQsUrmRVqd
/UvFwI+Ymm9bc3VxenDXc+O2Bqe39lLOoigfQzWpFJReXOQr1pKylEgezPodjyw7
5+gn9ezF4NQJ405GhYTdLBo6K0vvf1Y3pdi0cw0R/G9XM3mKo8hQf5qmP9+2rWGq
EeFhp78ID5TgyK9Q1wrADIUl2X2LBg3JwzQBq1znDl7/JH9Yspka28CLhUFz2Xwl
WLLiXQOG6enpzNZWaBitm8h8clJiKigylMBSMk6+D84Ir1i9vCHrkWTMWq2I91bO
a/RzdwD/M47f6H95ugwODav2wobZK33CZahazsX+NzL43xuI04ORkwQHtUrPIv1n
Nerykzh5Jn+aXYJgRnsRuH+S0oF5wrf9mwNf2Thaz426aARqLd8eRvsvUBkuApio
zZR2/s+mGccvmqq4ZpteFYphGgNfH/jlElqaBJ1ZPSjjnSttotx6zKqOl3gnXyaZ
lyOlQFJREgFhxF067dfC0afyDAE858B70TSyUkGnJaMW/nGvWdaXXjDSh1t7oA1E
mbbmlj7xVJ5E6SIW6OPQtemQgIySUfrSMr7suV4XjXdwlDQRGcLCBe7WHNXJtMzv
acWuSP1ZOpbBXnZWxs4xWSPS9GqsVwbSeTrPrhjyhfZ5/cTFaDu2KHnVpZQDnnvs
a9qQUajJQajQvFq0a8y7V/CoA0YY7VCvRQgFtK1WmvbuYPVvznKg/Ikzn+CaeJBK
g2v1mfwzlTY3gSZy3LE38dDjSLiKR1/mGqqi5pUk5UIFXCxQZKWVe9V47dQ/ZqAA
ZHZwwXT8q2HmrVouafN7Jog3fQneZqbF9/wF3gweW5/VRUOsq5e0WWleQCd9ktVo
EbqlMxDALC8F9P2Qmmyy4IAOyD5LMy/51gkXUxggpAAfAIUE1ih839mE6OnaP2p3
Tdm0hjxb74Owzcf/rTCNOGR3I9aZOPJffa+GIdS+dANwPjGKPniZmn7sW3iwRq69
aLXIHZDIh4JYrCnTcQ8fA6R8NkZ6L9HP5w8Iov+yhyitg1EqvrfO/Ux0PGYifRZc
Ysmtk7aqz06T/6S8iPp66We2TpIKwfdLuKQF/1kY8Ba0Cet/TYHXA/3BkfGL/pSZ
Sgwya+3PpmFO8QMD51CVqlswSfYSkZIIE24tqx8JuifVlIx31NY9SHKlShcQHD9E
AlE4LaBp6DuWY7xCzRliVx0jdnS0X8ygZTKrPAZNQafKYiFlLC1RjeRHM20xgHLn
GbwWVUm/FN4CM9jFw16OTC3+Yxf+DK3MaFqiuNemrrEL7b+m9R5fq6Xtg/bVTla7
aLkssD7wEZi7XwTD5i3cnk3UzJ7QKeJ/1RIqfEh/NPsBCM3l5OSGy99DproI0gRV
MCL4g8bVHOG4r6bU5F5w9ccgWYmVXTq6vb+XZxXjJyCnCwBVSDHMQG8QxV2I/q48
NsTBLjR6IQafL2DZeGfe1vR4m0X/0SZARYR6+7bgKzXCstspLnCmNJCVkwr7ok7K
e5Qb4E7DF2dO5P0u6SzoVyhop7DYliFRqe2LzhqVuLUdATQwWvmmHl1GuvjUgaVz
+menP8ehefhcaxXNk2vkbAInkLC2aMWPUp1VcXLixCpqQdnfQxVOv+w88/Vma+XK
bFROa+6heqgUX+Zhs1gDlEQq11V9g4qfHdmWw8Umk7C4qhpX5ub79F59KTtKOAFn
XNFYZNvdgfFWBxi9qf3tHD9l81xudUAo7U3x8OXwD21JySNJBXSuE/Otd+wHtfFB
hlofk7yNql33/E5KThRehRSfBm+nqoiKscjy/BoIzxCQ0Nvmjhq+boq+LSuNGDQ1
q4diqOBB8tWtg6Lu6d5dFJ1f0IwkZQs/aLc5gzFrW+w5QDBLZv94r4qlgEgF5MEW
gRExMYfr1wvIxGt8Mm9qqFbXkfdXG70HEorkQxPESn8f1QGuWlIiJEuYS1384l3F
FOXlYJXWKYpSzAINX7z4JxjIunEZdHIdpyzQ1Hfm4rCgLmQ+kxnpuCZVhueaL5/6
URVHmrNK5wB1ahWKaEtWpvdpH5hQDbZPost9JkEZAdjuL7E139yst8GlVwogaisL
uIaxMGX2aEG1Gpmkm3PB0g+0fzHgVNIGju+TStnGw85BOzhsqL3TUjaw+v5ULyCR
tP/kNz1UhsfVOBeARplO9/6fM0AAsMRDQaN9I9mnQAhaikcOuA+QTMM6h5QWz5Ix
aniYZzHkJjJFZudycGQyTrKDNUmIZrb8x6h25b3eLVq02HykZbpA+2LcXG9PXUaY
8R9e7VIqEnmhbJUpXJjS71JQSUDH5qS5gi+g0gl+MCyxN+oJMxaMYG/WwE7hxeZE
6ikhUxvmgFP0CIDJWl8s6+PjHo91lwjOz+WgERbbZ5LSlLKdMcRroB2msru+988x
5md1dJXWiyXMQpadLHCZXra0eeWz5+qKB1WcEmnM5OCay/KY0jxJKg3efgvLOQBD
uDe5mZVQpbwtu0zePpQh8UFY77Evr1tBsocfItByZTlJBz+A5ytI1vzkm0JIkaIn
FOgoYrmjYuAzGSlBNYdpthTWNtT/A5WaStVvye0vzo3QnrGQS2mhF1Vc5YUhKuMb
pMvXoDW+RlRkYATcY1WvJwEdxGSq5d6pCpSGV3Fkj8ZePUWrizuTXeaZWvGFZmJb
2HDQKVYEm7mazB6/Vyxs+oDBBQqKr9Ka2l6fuck0msLAVFpJZYbk9PYsKUmmKMTT
wG7dxbQKUy50xUJx+YvHMHLFc+e/Cujrsk6ZIEbqhnRJ/KZ5CW3Ej29OLqtEXeKT
wskiMdTPGSc+lL5k130fkoKYq3zYgZ5U4BVPHQUo+jA1eaxW0vB9NIPiL1EXKaVY
7QTsLJUtZJwmmx5DBYIZCd4jkg9ZKfqa1l1NfGY7NyrpYPI4oRrP3EYNci6PZOK8
5WvCtf0ZG2tMpV3b14llglhRsuzF3qpFspT/DThR9YJiV1JYL3JN5n/FIUjiT8ZT
DJ3OhPAIlzAYSD3UjNY3LzV9kZ5xjpB0inYzT5dGNvj3sInKfpoABq2KkYhIskm8
jq/uUFJQi3A2LMOmzgCPfLuXtXBtoKDijyXrmMDk7o1axt4rZquvy6HYlCJ4tTir
ZFnzC/8UCf1pG5TRKYLi3EndHZdSeXeUbfVYcZKamTEvDKV/jrVhGyVmnaT/lzAC
JTtstiU7Mk+jmI/f5CaUAaMe379UF0kPQPdYj8vVO1PCSewMUxrJA/IvehzJ1c+S
XXWwm8V0XEJkBgu60rZfl/+t4VAp8P0moZH6ODL5BvvJzHC27BfC4iFzRoKxLr3l
1kb8PwH2aQGxcMnsYQb08Nde31yvgXCQQ9tYSTXTDEVFYGRGp4tDWbgIFlMouEsj
Sa60gg5/aj+QDIipFJR2aMzzDBmLlBvvcpDomr2cQ6zNZYWI2jEjqJe+7NVtdZQa
xAMKas1Gv3A6vG+XG7dLGvIRgeRnSLv9ngbviy8G/Tc660lhXIpjnC0ySSacOd0b
/YDeYCqZkmc3Nre8Fa89kfNS3VENr+kE9BzMIxx/1WQ9zuh/LmVwa4XbpHDn38/H
kX8biq5zj6aWPfqWkXZfXu+HivUJIqa77jQ9xPPGrnyvPNXJDXXAUBzP8jXvvrsY
eVzsM+vqhjvtvWGhDQzyiOyFqMTCud61jeQvk3yrGozj6m5r0QzP4vwJaOvywtam
gXaFkJ/Ge6krCKTn2DTsrruslnSoDPTdgNFlM+XGqzMXQnPWahApNmCjd1+z38l5
riMaObIVnxM6ck6CUOHfmNxi4e76AHDv38Az4Q0ybhoqCAyYpEWwUPWuRPDHUyeq
Nwd8QkrcB9uGjkdvjutwfO6dBIcsr5+tFQxIeqU+KEfu8wbfXpT5vCwfuEBZrkpQ
MbpL/TQeCs/4jVMSjKvkvWOuPs2m98HcV3rEHitS6kTrMYA+JVmJjj2y9cEhjY8X
t6FQqlVrxbAxyyUNwk4q2AkpKnJwiqT7Sd8IXVekxsn2qaRN1sRP8HZoLGedNosZ
7ZCRReMP/vO5T5nBblMomwrmUTgywiXzyaox6VqwrZnvtBUiVBEfcgg/lwTYWASh
lxzytHxnRKDfU5mo9+6cXoyZDazsLOpcX23hbxA2K4BWXD/GP+n3byHp0NkygJZK
2j0tGB0EqTbJHLUpdhco21pGCRq/99thYoSDrS42i8XiCn4l6elYPu2LcmxguoLM
wDzbg1OdoN1rrOATKhkR9GFMHOPwZ23H92+DWRy6ir8YYjemD/BRUKJ7uFV2Qwje
g8lstt4N2m/5IOviFnuSLomshwaBpG40oG2t1Bk+7yzZ5kUV9po6O/tl3DCkhH40
F1k3UifcZ7Rn3wRlCrLEzCIhLzmUThAVCEppSUbO+TUk0ZbWC20+nS6V8nJDfRJ1
U84MoPeqhvPUflk/WNnUw6BSOb8YfvS5mzq+0L7ct58EEMpu+oBqXJIOvHg46b54
GyheS7xRINqFrsNTaMTBzmeaswhcjtd76Z8I/bcLawEjdV1yoLEU1O8nGjasiD5F
ZBLTAV0WvyjO6UhHXHb+9JdkyMtxnxlM6rON29FgJzUKfCxHYIayz/c6YOicaX/1
2YPaSABmt5TnKexNDI34Qb1QMrrGiqRMP7Cs97NcUjgvqIe35OwCWcG6qo6k5V+u
2WAFXDAtZTcYSh+CHE9v4B3fL3krMwgvL85FFrhObTylCuPXCDwzjO/wZ5ORuO2s
REFwyWAYKwsZhvbiosUVc8pOKPcyU0wEscJwaUlQj+nSVCjrEt50sVhzwOoq6mQ7
7LlwcDAasOlDRe5pVxNJaG4adJtYOsHNnjKkW+JwnwXUaWVMF4yWO1iH5foL72wj
Vv5SmmQsLZ3c+goUOp0gVZmAliAC7J4ZeBy/nxbO+nEDoTXkK7sc8mMqsOIedY8Z
SQaamph7yF4X22AtZxjaxEYc2bFRhUOHdZy6OgENff43OrF4rfMk5OaNklnEFAOk
ELhpT/v8mn1bTuuysdUhDMgE7nCiKpDpu9Rl8IW9HwU8et3wtvMn++uspu8mZ/cR
4YHLIOjsSpntjoimt2lhiv7tf45z+eaoUrq4SH6ZV68dLJOdYWJiyKfpm7Dpkiif
p+gacoS/GiuvOt24uEiajLocbyBNcioyMbod8BwN72rKJGTmigGG3MI3m6g9LJCw
6DRmuuBNyRW1E4gdn0UIwBg7dUnfCq49TJnnGLqQHmcTnEYSlDUdSEH/iblZ2lsK
/wI6/CXN+OVZQqH5+o9ZL6cDtib3jejcZNtiGe5OM0ZLjYUjRRYPEG9X9nO1k3mR
oq60egL4vQBONHNPmpd21Rrjdmnq6RvKShjpUqjUYAIiDtlOfoG2S4s6MVplSqWO
hUNp4LrUQSzd5f/FJ22/bFyPEZM3S/dv9s3buW4Zc0cT7aD4LA8b/J8FS2z1qu0w
AInkIbKmgqu/D3Kd9rB6AFMoLjvMCQgsHgjBhk0iLLfBU3Jl1rWBMDhoha0HlJvx
eHwZPq3qSLDpPxUqLTbqCjV56unroTRUwQaInK5pLFI36DAU7YRbZ0aKuIoJKdBh
D7ZTk0MASoVhRAqUHvnYnff4tYgYaewUa9EL6uY7l1Mmc3q2szaN6/g9WDS1RALc
vroJhVb2nVl4swSvGrEUyFZeMPSlInljUzx1kWU/LnfYR0YCBmnVV7Re8ilN6Wn1
Tl7luTyhucX3a+oQz8t3soZrcmH6q1i2AZjF/CH5Aiz+0r0CW9mKhAj/Eh6fnnbx
YDC6JrUULsuCzy/qL9Db5zQJqtnWvjIKVuU5taAbyVREe+zSzzGp6ArIt3vaeYhC
RHSTsvx7RBARkKJv3GKV/5LYwT68NRlzLZps+bXJ4rjl7eVXXhCl7ILyn9bYvCmR
nkKGpDAkg0OB40s+Aly8vRHs39K4Mni+idlOTEJfjXLsT7I7lr8qLiL7yJU4lYjS
nFQfzT/VIb3MkuMJ+RbhfbzsXqUT3kBzDqt5caeGd9P7cu6pvMRNgcofftRN+VeU
gIQrsSeSe/oTsEMrLxaoKci0P/vhX+o1ChPddHAKBtgmQ64UDg+oAiky6ie6lS6V
t/Jkl0jrVbKqNXk09ttmXP/aGT01X66yEpQxwheWmv8dhiOdz2OoGPVuuBx9VGCJ
+Vvvdfxbljj6Yd/m9uVfyBM8MJ6IVxYawjep+gh1FZnmb5ND9THMU6aL3HDtBHeL
CLmDamt75wHx7lyue6OD4fql8k4zpOy7e7ZmxkLVOVl3H17aiCdxieAGS3Quhrnp
b68lfQQysbcomAkap0HOtbtWWebqQeXRuzeFswF8CDmXt1KG13HX9hPnWOqSQPct
FFHneEqUDSYWRRW3SnGFh+qOKjdfn2U/AMYr41hq4xIwO7CSAMeZwpFgXx7B2n+R
DTSovKv24aO/bGVtAtLAnyKVPqa2YmoH+KcRcqh6rDKIlKVzpF2olx0S5DVX91ym
ZXVfv8NW9b/sSsOrU7zit6Y6oXOIXYPJdj5vB4BRm2653keq0nrp/svGFlRE+xqn
sYB++xH0532U6uz2ULR7BxiEeoIIeKmyRxvMPjSHHc/+v6V4h0hWoKHOQDbJCxAX
AoirpfMKnCn/jCLB3yiOj6u5gl86Il/eYqcZNvIHFZU9alnJKWrQKq31K9gs9pD2
zYhU4P7WQ5+hJRaTLcd+SNdX7YU2d6ngX/l2lT2ZDmJhd52pmg0ZFvVey/SqU2tl
oTknH2BX7iZbFp/HBS65YBPIMpzqGK8khGwM3YVg8syJ+gJpxKMuZMSZ4wCUZzo7
AUzyKAzu+Ft/tEAT8VPXuei4df6LyKxfx+mHwgChlsGfQbXuecl/nlJe9CoVqbpd
X/1X042B84EjV0TLBqKkbj5ADFTclFtOD177rWGdsSdltqsI/oEsjg8nNxpaxybl
nFuleC1FBLzJAeAZPhCJkFyRRo6sAX6dRiLe/MZGQz6oTnRLxGQ/b2D5PwT7QMpm
d/hwNjFiKnH0KqyeysCvtYj+BC+Ovo5LLF8ZcTXlfXT/1wOo68kEjeY7SMADgjYE
IO0t7yn9bnBwUPUOzieOE63PhWkbWWBz1DoKFJt75nbI1wkqgOKJK87Cya/385w5
rRkHPYm4MtQrIio80R980alYfTm7fmt6ljtcwiJobnQz4Gi0we+UUT3tCwbl1GIa
T/NGdsmbu2g+rQIj7xBQu1Xm31eTgrhQXh0F0hOl1yEEz0jjT3hpBbYpkpmXXsqH
cl+jUT2oWKS+8gwGGAqfGkdFtze18Dz2btwwGaC//folVQP0CIo/kIJnQ60ILcMt
7ZFrXoIzQOlBpROIx8UKsntQU/8FxHX3MWz12qQg/BI+iDIh0Py9h2BReF6/skqx
pDCc2mrDlPmmi9KKLaWlsFlnV187bEcuOYkszckkqVfnYfd4u7djNTvdb9B8NB5h
rVlOAUClzTlRMjUYL9g9/q8stj3NpSIUBcAo8bA7SV+o1sgfRXGmTrQ+CSV1pH86
VEsWyWhjGwmRSWDvMvXmEp9whS0dIPrlpgO/VPKyiciXR7GpQhMoJNb7NprsCEmO
dR13/MDqnhZmUipzrBwKBpKxq8Ah8RdMTiGUfKj+5EK+O8GmSYxtfFxgi/NEjTC5
tXM1vp0a3E6c8YHPIloP/kriYobQTQ09Th9v0ltjOf2/A8FfQMpOXIqwot1sIMWn
AE+VXYqM8GqWj7xGDFGBeK+wWxupp16B+K6U4+icomQMp7bHh7Gk0QzxPvlijA1F
S92zKESsRMDx8oZQu1B/iSNKDjGpmDVFoir//AiwWxNFmer/hfkCepJDV11YyDue
DzUkavd6WcUf1bLiTu8zP1a3/7Yk5Y0wiHbkPHRRwzQ3DeWtnc/KSm2luIklGO6k
03MNmNpWpC+w3Qay+0SxtSp4hAej5nH4GB5CCoHIpJV8gB+qWnFoVf3qxQV70zMG
hZVFwY5PjeoqxWtjcLFM7DFmsFvz4S6BpiXdLmt5tgHLyPsH0GhWSxIDRBZ8vVPD
6YoE/dQ/+nol9jUxvgkNl8Ti0EjyeatreEhmM+ViZ1qEhGFgDFF2MGFWm1TOSUoj
pO2h/9UjXXl/nA3FlSH0cQKqXMYid5gnDAdFgAMc1O52rYBvnwCcc3KTcpFFQFxI
O9F6CTquVGqy8amlnhwDXnKHI8bO0lrj/hu4xdh9/iAGsfCSIJp+4JsrZyQaSrwB
FxtsFNR4AIVod403JghWZHCqOyK+owRhwZSmGrgZiwNFHiJRJ1cwPpxFTsgxH1lt
3I1pmuu9zqqoPATb/4yY+uXn1vCCqbvY3VFwTjs6veWNdjJiROsiR+CRDkHJQepi
ml0T67RpR7UI00cWrXUxcs4+zkEOPjm1AKk9MwnZWneFNys4npEO2lFicC6Z/cZ7
R9vICmcCxUEjJrUpCGT+dDaCA1MuHLuymxiaBLJlk2b3sfumd25UJllgy6rCZc9y
CCqG9NzxivZGmDwKGQVDeh9mlE215Tknv3clauWCVvgwpacR/J81Ha8xJwr8+ugj
Rr1vJ+TFTgrYugaGdHjIlnc5vBeG47PturjQBagEHcTw4HlUW1h7ltsAkUsD2URg
ZoYJ+Fifqbk0VOcIv6QegQMUeXvuHHJ+55bN4+HJalpjpdQo6vvVkIiDZRlHIVfb
xn1nWRkhLPK/z2Iyigz/LiyswsqRUmu4i4RwyckjXMkUe2OBkIIdzlNA7+EGP+Ng
UCBnZ019q1BZFXir2KcqZq9rwuCFWMz54C4ySSHquUvCtUBNZA/Xs3kcbLk/wO3p
grCL73sGH+x6quZkPSoLxkbo7MxhZp0MWL7J0OsLlKZmsbi1577calKo+xwNWcqD
9FdU9YH3+I0My7GPdwMJOCMV5hu+QQ5sErMZKGklqxOOZkfA6zqcibwvXPn51O+3
ud6YnrT2NAgVCw3C5evmgY+sS76M/WQPPxyRFSqvJLPpgcET5QEmo1g9+XIu7cJ1
lWSr/sn3X1UBjxwitzPsdDPLv9rJmkrYkpTkixLjW8/1cLrggC5UEa63TvYtxMim
l9Hu/lzIIJ7a9jc0fIN7zzvGJ3YKI7yV439NVtwy0aiHbYGPpPuP82ELIKSR+0qr
Uk0MfFozBRmK3cM/BTkt9zOvmfDNO/udZJIj6z6Q3C0g9gxLjnS7QD3POQQ1Gq6m
BTGb5Cst8mPFfQjq/8luNfGLYMlKlNMFgeq2EWEGt3B2OK4qAeBgYd07ckxIBgW6
9qTqAB6uLPUUyVsn6GY31nPHoYNO2SPPaYN6LPebfjaFbEZv2frHY4abI2Isr+Nb
SIDGMpc3lsz/5TYBlZ2L2qPG6/JbYMWhw4a/WFFMC4GaYd+otwYScHo12MX5cz5R
3ov+zxL5r/FFa/1JpfZuPO0Y6Vciu1Y8U4Qa2vHrHV4EZZVkGnbZDaLFtRFBxwKF
17d5N+n6r6ukwYySAjGyY/Xx+o5E09tf5h9TMJVVVW5bcqFZ3IOn/Bcw/nFoupyd
0mx7W7Qh7V9BRBxyUnEzULMd/wtJELWe6ZnCNK3AOeJle187HYNSJbXyroM/+47B
kJEdt3IKLu88rN80FCUmvZz2ZhOY0RUNvNFc9oaNSPgGiOeOPvu0xJwQX+BszNj/
Cl3nc1P9TFy3vNNEuWlXVPfUv/iBDYnQMBwyj4fJAsEtn/jIuyGFTiRnVzgiufYE
PI3cWxbZFOJVr5HaKzd349A9T08Gqu00X/+4s/kpE3iWSihdjHZz2gMQHtnrpo+t
9cbpLFXlN96h4zUBbBt1zAU2Xte9Bie52CcqktsJ4zsLPIIagEM1BB3AxX7KrFW5
X14VE2XzUUYC+Cx6J4Jgf4dVwhKBDQsnb/A7hLtWKf9piqdoTJRgEzXdJKVR2Xb9
UvskMBbT3mLlKeRUpH7JQgeA7qHn+yv68qnZBAQnCztP2SJ03TGS0+wHIhWbw/r7
44P+EGcqQAj8CuJSqS7o7cjx97HNYesF7mUYKrrpvD1vS2SKGt/XMEvly9B0d86U
pmerJOK1Nsk4QsvPsYkn70jhJ9Ha/gSexmGDFvELhUeNFQy5LyApKuRQpSNjHXjH
CH9gYUkLd1Id/QLhDBSi52k8cmXzYIiLKzoKH6SPSPLX4gXgTYSYmdPLsUknHHi3
CGWS+6zDpr8VyfIsj0cZLhQ/w/sae11Sa8tL329XBk2xkmk8HjPz23DEDj1yOnoB
kqlhD/PON1Xa3jjpIl0mIxWzTd+9wixQ/cYWn7t1wKJ/EFBVaMG4of3oXVU5f1/m
fBBmQR0YzscGCI/z12HFNq2iI7Yn95woTExJ+LZl23MGcgAZLaxV67KGecCsx0+E
wZ6rV2bRkb353N7GO2NCNNMNeeXzLUw6FRD8UWdlXtuHcGC2eVs1y6IJkfdHkc32
dQuXDCgr9TsqPLDqNu9UBJMmqzEtKhWZLu0RsJKoaWx8WVBdK2oMDsAoDPxfHnYS
1YEIaE24fAfsHnZ6CpFPNBtENkM4klOvxU37icyGLttDrgERc4UGO2zXuzls1JuI
NvyHfGJX12lNqKaASArUk7fvac3bdBcXbhnrhzmp9AytYQU+aUsYzBK6t8TMLtfF
MvCSLrbr+1eehWVDM/syTqGI+MIuScLBZ6a5meMd/KwunMnmgt0GwJztF2AArd9/
bP3mk0ZOikZSKZndMNrq0DD7kd+TpzGWHhIDAzQ9RuE17cqGU03nCgFM8neurOZw
I0943Un+52VtGuhlIGs24KPgQ5jzLwJbFHaW11ewx0RHN7IJi1CVd/+dcilwiQPf
1XpRd4Jeka1dXtV8F/S5bcrzo8Ar4V04Gk31EL3yiBFzxCBV+gPfAz8BzrLWnDo8
EUFSjT/OB08QDIjA6rzujY5pOpYvx+vPxC86b2jJnt7RRz86p3wZD+UkpK2NauXH
Jr42d2ZMSwMJeWBJppsjOVz0mCua25EaABlZ/J85nzFnBUAREp/jiI/g+7Lhfyd9
3jrH1rrkjNdrCCDRsz+h7gPOSZIzL9iCI89VdxaJUfNTa9t71fPhxJp8xGrSizwn
ZWcSaw3MHciQVp/5UJkenZ90KF44vnWlsj7BwJapoYR+nKkvU1QEjo4U1rWD1LiK
bksZBYFguHEzrhlTzOIxlBvM3soeQdI+VHdg9HqOAFqCTJ8JpUFsjj5jQUA6ExFj
RJbad6DpbM2gAOTvt6WU0fF3vHrgyMmfMSMaj1DlhJgv/8emWfAFo3j9uZGZNSYJ
HRjvjvF/7tVEczkjpU7Ew0ehVdq1xkIu1QEMmR/NnJfG4tLh3Dmw6GmSoFKUTuj6
6rOBvqeGYryBF5ErBGPb8tit9vkDkPr6APyAsyIA7esE21SLqkMH5lOZGRa6LMxc
`pragma protect end_protected
