��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}���3{M�G7�b��}�>�Bґ۫�3�w�f��2�O~j�W��E�Np�����5y�G��������L.�*�D�e��BP۫l �)�r��&��6�,X��d��h�}i��dG�ߡ[��Ǔ�U��a1�G�g�Q�huy^2�4�Z�]?�8� ��*>Ԋ��S�����?� ,I^o��L���
b]&
����Z�b�뭈��ҹB�R@�:l~;�".�d�C����#�>���8�����Q���%q�U���8c�o\< �O�}��˺�p�?�z\&�Hb�#����tvID�J��c��n3l=��3��Q�VO�V��V5�����N�z�����(�����w��w�ssn�.op�ڝ���;X�3�z�h�k�.O9j&"P�!�b5�-��B2��J�����r4)���v��v��fď�*�u}�[h��M��8��%js�D+���Fx=\w���X,/9�;.��n 5�-���4xO��F�oM̞~@p�/��v�;= T���L����cR�p�ܢoQ =����ff.��5����ȝ�`?��4(����e��h�DEV�q�d3N� �n�|���Ø�W��b�K�]x>�I�Sx6���c��9���`V<��IjF�]��e�A�����!)�M�	x��yז2�|ac����/��X�E!�%�nRs'XZ}�X���Vt�ZU�i���CB���G��\�c?�?�����$���p���
�����-�a��kD��+?�4�_|7_�f0�����11Г��xC�=�s��l@�O�Ǹjf�;#�90 r_aK��gp�Z����T.�S%��ZO� ��Kv%�.sT�wܹ�bT�gJ�k���Q��tD�ھ^We^`��i��m
K�kC0��|���Px;w�;F�@h�'.3��ij�'���n�޼��a��T�O!f�53��0�˵��)�Noa�G���ѷ�*�}�4y���b���{KNt���������Y������&Gf�-B m�m1��Q2���Ih6�1� �7�%2�ۡ��ٮ�mt�I߻�E�y���(K|B���Ep�Q�s�FY��r󗸐[�q��A�k���
���]��ȇ�����	j6T�o�eC|���k�:0ȩ�� rbЇ��r=cndQ�=E��F��Y�<�:��`W,�[���݈���O=�Pa��;m)J�d
��|���V�*\����
'�\J���ś�������+��0=��`�e�Z�Y	}9���n�*�_�͆x�`4ar��>b��>�~�7��ܺk�2x{E��UxȦ����1�)��>_,;%�T��_��	���`Ǻ�|b��{��	m^�J@X`����D���ȡ%S�Yh9}Hl�|�f
�Ѥ2��%Nc	sw��aRA��#���lYJHe+�r�	��h �c6�����O=	�>N��#*��	�Z5�S�]m���~�8~G���$�e=cg�DdM��B����h0�출�k�DFN��'?q�;O�:��$�;;,�p�A�G7�� |�� '+1$[ �2V0L+h�qሹ;l�ou)���ܔ��R.���e3�65�痌��QA��k���F�[�EI�,ľ�V@������Oc�ʖ\Df���G0�awD��/����ǱV�5s �������N��|� �Ş?��%a�=WE�`�!�h�n 7������/b�?l1�&�Lj^���_�hl?��$����)K�ӈ�"H�\�<��Ui����"�,5.!j��}�5~�#�7��N^��a)��F_����G+�b�{<�J�i�S|����z��)��!�1��Ƹ�SC}cz-30\ks�[�ו�7�I�Th�U��$/V,%��.�
���3���׶�1QwOj��Y	[�X�þ�Z�C/����e����F+�`�Z=oS'Vvb%���$SK3�̡��Nb���E����U��:C���Bn�屽����ue��b�	2�"!��U���ס�IN cd�#����E".��a;��UF�/���A1̗M�w����P\�l$�-��<�s@�d6�d��Յ��z� J�#���6�����p���8�v��	��E���i��:t+G��F��u��k�$�<$*w���P��� 4|�y��'������7���|9�}d������h��_-�p��\����3�X�7�Mx�	�Z�繺��Vx��T�.�`�i3<�ԃw�!I�@c=�����x�v��TI���?erE����cf�#��!D{�b����u��u��;�P����%58���HJ�Chy�z.��
P����Y����<U����^���{&���j\N��>�@\ݴ#�ma�g-,P�9\��S����ԓDU�]6�J�Q�Z$�t���Ӗ_ӑ�I�)*FD�\!¬-_Mx��e�|���W?ԣ�������Y�2�>
���2�|.ld�[|�y�# o2�\�p5N7}m��M�!d�����C�J�����[!+�,l�	a�:o���&̈,�5��	�1��KjK:��.?��������mɢ#��S0���!�_�?o��������8��`�����A�P�.U����]��HXh��wv�*�3�����a��M�}QGoq�/��ߚ׋�Yԡ�젉j�WV�ǆc6J��>�|!�CLIq-�X�g{�3��W�L:#p����(\fˉ��`=��wҸL}�|��g�S2z����;b�N:�l��%�(��D%�����CBh	-b�Js�*�;G�R#�NS�l/O+h�E�>{�s��u�n����>12�DpH��@uZ�Iٝ,C�qD���k"!����/zm���K�u
8�A����x�D�)���ur]K5������7+A�[i�F�0��W|Q�c$f�Jv���1�E�~.yi�0��9Xbf��;هx�.�����Pxz�<���z�-YB��Eq���,��I�΅��L#ǘ1ӘH�I7l�8/�*SB},���V�euO�߯E������|���W��0N�Z�6B��K:iz꒽ԡ ��U��ky��g�6��y��+S���sC�{'������j��5���)>'a]hW9U|խ)XvZ�l�^��D�0�XY��,���A��� �s�!�������8�6k|I�Z��/�
�܍�jv�ck`d���+�Z9�>���xW.�
�,�7�z���~K�
��t���(h;u"�ەK����ˋ�mF����VQ.�M}o�G�'33�S��*���>h�h��ۈ��j{��S���$����<8nqx�.��ꢅM!R\�p�������b2 �ȳd�ˍ�y=�v
�u-�j~t����Z��K�-�Z�Ӣ��
��:݁�W��(� �'�4s7pbr-Wo�O�2�.�)m� ���jbb�#KX+]-(q����R-v���{u>�~-�C��v�ـa�,�gʭ�-W���gs�X�Rv,�A�Mb�`a�;�y�]W�c`م��_�V7"���yX1��A4a��,ɰ�r�M��h�|�}x22n��^���y���e09Q�P@����� !���|g��Ϩ���To�ζ�u��ڦ��y��ni�}�
���P�HrS�W&|=2�>%፱�.E�=�sK��N��U��N-��O����Rc��ToiT�q+'����W�͖�>�$�(�D��Q�vJ�_��R��& � `������=ܫ[�=�\���R�J$ӀPA�YI�^=�$z�c�~l�zS�$e0~���qf���eB>��C)i��-y�LY� }��S�A�15>&Sbp������0ZU|�ݷ��7��Vd!$�[@ k�����o��hio��+n��� +�������c3�,��~xFǥ�7�-`���_K�d|,���\6�K��� .��Ԇ����3���H'�ǿ���"�Oyt��Q�<��~cz�.���Ƽ��I��L`�3��ᨽ�~�E��e�0��R��T� ���5yA!�F��Q�åwͱ6z(t찺��i�
$���z��~7�Xt��ƨH�	�YiQ�ԯ��A�g�-d��38�;��c�Sm뷈@�HD6t���	x�CS�Oִ���"���e:^�h�	0�.��2���鼸��4���}��7�O��Tu��Z]m��$�F���m*U_��5�d�ٰ�D�ؤ������ ��˭��$ƣV�7s4�jqi25_�.��m
�9cq�Ý�� @�6b̡��8J'd)F9�Z�p�D�t�'P����J�w�c^����#���f� `>����bv5�-����[���,�����xM�${`��Z�Ct����V[���g���a�ؒ�<}� �ӊM�OrT�nmF�-XZ&ȼi�P\�]�y���$w��L�[iaP��t�kd�=sQ�h��ȑ4��6���H�oa����p&�� Y:kз!6!��(��w�9�F����o�,Wjb��(�.�%gd[�(��|j��h��8�ʿ@
]�%������89�~��O�����{N�mž>���[�m���
=��{鮖]�6�61�0<E�S����Q]�P�ty��Z�Q�}����p(d���僧\��Æ�N� � $-s_׉�����XQ�O%����O������Ưa�Ǆ�P��2���c�7_8�X١9�,p�E��f��	Åí���,qwJ, hG��U|��n����>؏AK�цx>�'?.�,����T���*}�/�SAN�����Gr��Э
�mQ5�C�Ƥ�L`Z7#5J�4b�3@Fn�(���w�oo��k��~�$���~�k��f��AlpdS�.�/zU��f?��N��f��_��<
��{��?Q���EU*�;��E�!��`���t��1`�ne�;t�mI0���,���j���JO�d{��L`�����F}��
"�0�1�(�۫��v�Y��0��-�)w�q�Z�N����
�m�ZOj:S�,��k�9J�[��P,c3N�����Z��|	fA�j�L0[���S�i4w`��)pȳ�v�o�AO`�<f����}C���o<8�� ���~:�f�,c�Z�M�ִU�݆N����.�,�)3Rj�Gү�B�D�訮6z����`��X�]�k�@bn��j���Y>��p��J��좆�v pjg|�r:z�&4I�L�Y�m"�Z��L8)Y�ay��P6��~��t���k���������Y��ϝ]`��0C��,�U��w���&�{��$e4�MS�[����U&��N9��3���8����P��o��I��iuc*����I�_/��q����ɽ���m����h׹��3a)?L�S��|�q��ڙ\��|g��G��5zL�r�ڪ�|�y�R��_J���a�^���F��7D���.~J�����(-i���b����T[����/��xa�3���t8ߏCf8��ul�ql��nr��@����͍�UMz�u��C��22UFZ�x,�(�k���#p�b�nE��|;8`��a-���~��b�/�8���o�Q�="��O߳�ϱ�y�
��~�mqfg��nτ�MN-qEs��[�h�M�W|TЌM�q�̱D�ػ�]����]Y�8I�QPK��7�A�x�R7���zdz���jVdOg9���BlJ �x[��q���gؿJ�t&
��� ��D���>}c��O׍���^i��B1���	��S�!75 "���:XOџ�X�`�Fa�@nD�P��=aa�>X���W?,ݡf�J-�7�Hh�'��Q�-E���UGpG��xk��Т�yr�hG
����ӣ@�7���y�y5�;�O)�Sr�-�\����i���V���'��8$��vNc��R��g}�!.ț��V)PEXA�'��K7����l�F���X��򻴕�q`���hnͨ�U
b3�Ү �>��xc����p�RJ}�?�@�\4�pC��lP�V�������wU�w.��K���X,EK�]��.�'%���ӯ�$D�[�I���]�G���ﳔ�Ѫ���"��S8!���ʟ�
n���^r��+��t<ƪ�mU�Ƶ�˭n>�T:�{WLI�$h�*H�L��1�y��%�ܚd���O�t8���e�I߈�a�f\`���j��ר��y�ֆ��l��[	,�Ȥ���Gq>)#�h�P/����y'P��q)0�a7���{9�jsp=�÷��\�֜.q��~�8tQF��������]T�A����H�Y��b1�9*6e�x�1����N��t�Z�ښ�~�jeI��3�=r
��k�¡n�닖�lp�$I,�����I�5v�6��\�`����G����.��
�1�~��!�j8��<=�:XN'�l��[;TX{Wu�y�N7۟���b��K�8=�Ϟ��sDarE�C3�)����r\�
np��Si�j?��X��iZ9����`����{��)6C0=��r�X��=6��#I.��q�W�BK�	]���1�9z��m���,�/�F��T��ڌK�ۘ%t���,^j�u�#l����^ƳXׄ�τ�T�"Q���N���g�]r�P�Z�϶���]�
ѭk40r��v@6S���<��a��)� �$��[�YӘ�L���y��d˹ߵsjM�m�����TR�`I������s$�uI��D�2TQ�3u!��a��֚���T��� Q�1�8X"v�+j�%�e��#j��kc�j��rK�9f@U�29�8D�=�u��(D�:IH��DH��)������Q�=�'��,�Ab��a��`�ָ>�CE��A8�<O�^�:ϠƎ�� ;M7Q�脽�:�kz�F0$�Ҹ_S�:���bꦡڜ46��]kR�����RAܥK�L�]��,&��Ѧĥ[
��`�My��#���Hi�� �t�nx�B�Z&(Ё �=P�@��~�~�k6u9_�3�5���[c
Ow��}�\�� �:܇S�>���AD'���`D�t�o��jއ3(3R|�-��\��v
���b���	U}����-��J@a�S��Ӻ�=d0�3���U�<z��RW<Z_P��(A]��4ɬ���!���2���.�߇�^�N�O�9�P�.�B�di��B�u����&��K�zH����I�����n�[jx,y��~|���4��S�LD�g�L{�$_��NW����_��i㨠=����~[E�أ˗K�s칁F�x�0{�f<�hg?�{@)'���̅��l�h�JzG�dXKW�O~8.(�Ǡ�7%V�����\`_��(���3�w�0���L	�XV���|}���ͨ"��2�=�4�y�#�Ex�[�z|$~�٣^-jYi�axӏn��1\VIR7�k��}4N��Ru�aT�f՛��QϤ4�m����+qCؾLMy��US:�7��3a$�A�w[aКj����Y���oו���|���H�u�%�T��|mB �Gu�fX7KO�Әڼ���ߨI��sòa�����;R��x���nOy�F�V�!��ST �p�z\`X �'>P��#�~j��*���8�ꢘ-c��(�hs�T����^M�����"L����S�g��M�ʣ�ڛgk�$��,�	�$��@�K���.r�����Ŧy��� :�YC�e�䉙i/����y4�M5\ ���ˢ�Kw��ժ�)]��M���:����m����2�Ƒ`G�n�UӁ�s80�/�	�H?��q���!�#�itEa���Zn�g�Ըv�	ƾf�_7"�$�U5$0V���X����%̍-(m�x���G֮��l2,��%PbI�#}����h3�����o#=H���C���L5�MI��V������4�ޞҜ���S�KpCM蕭��A�߫['oh8$P�~A��G5U@�ߏ���b|�(��U��qHӜ��o �&QԜ�y��D� �T3��M��N *��xi\ϦK��vUB*��,*��9��w ����:Ә�4}!έ}�'����}x�n�7���>{NIn�����nR���Ћ�D�K�鶽�ɶz����(bU��H���l���Zx��i�f��':1'9�7K	i4۔���e� %�`FCYR��{Nc��s[
a:-{�#f�\A�~�X=����K3��lTQO���LJb��+y����,��gGt��4-��"�����U�i�E�`�g����禟��F�C���	dn��iG*Q�3S.߳	<�LF�_m(���g�Y��;��<����h_�j� l^� ��0R;�sT�˻s��y�G��}���}&Z N�o�����@sv"z�_��q��(��H�e�6Ժ�zp"����7
��b����{�c-�4J�H��5AF4�l�_��kM��|Q�l�:9$u��w2Zt�c%&D-^���-|�%|Ǩ��)ʞƒ�#yR���^Q!��t5~�P�������ݜ8b.�R������r�xeeY����k���8�T��n��d��e��/�]�� (�"�����`#��'�Sk�njɛź�m�C���զ�Z=�#ѐ4�	X���&��L��6}�Z�W?���~Iν�_N�O�d�H[�Z�C;ڝJ��,�ؼ���X{�(�����L�7���d��9��q��J;w�g��?�]g��
�y
�L,�=˦"�T�r�	FD��p����O��~S5e!qH'biH
I���C���K�7�rxY�K�?�f�0<$�D����-]5f��t���6m�g Xz�z�-Ui��?�SDR�ɪ �Ƃ���������G�l�N�z��؈���L�wP�.������y䑍��)����7�(���j��α�X�7��$=~���F����œ�б]�Ra�,ڕJ��xa
1����!�k��o�%��v��:+���%�)r���A$K�������d����掮4�)���+���,,��+P�l��#�R@g�{�Q��� �L�m�֣�$�����]n�8���`��i���qꏥ��Z}ټD��D1��S�iS���@�l;$V�lmJ�þ&�^�&ҩHD
,f��?��YW��y�钼���:��[c���NEOtJ7Ru����%~��2!P�5���߸ W��SR��%�6RDIS�/��BI*r��\_PGKn�8�,
K�T<h>֟On�{�B�v��,1�s������N��\Z�lV�)7���I�S�L���Ik @`_O0�*,ƈy`�q��$�}.�2�ͼP�.@	w��|�V�!S�-�q�p�e���YX�dXG�Up�;Z��#}@�?4�}��᛼_��.(���ڙ�I۞�3�L\c�_,56�����e�Ƕ����e���<�R���n�yޑ(��v��Qj�����q�6Q����>n�7��a��§6�������9Cv��Z�YcV�����j��b�<��9��e��p��@��a��kK�@�+nE��4�T��ݕ�t��p/v�{�0�b��^!�Od�-2�}!p��yf�|,�g����9�,Wi{�+���u��C\��9�0z�����YM��x�8�W���Y�1Q���6�35�Sz��x�G�9	E1����\o�+�5��Y��z3zz��A���\�2|b,t�c�nFؤ*g�p-�b���?Jd����Rs��`8�?W�o^��)P!D�E���[hgq}�W煣S�I�R	g����!p���&
\������75��w+�{9��J8�N?�����5�a)��jL0(du���E�I��c�,f��(0*���P������dן�������t���lN��.���oo���	���Fs�|�ٝ�=�wJ��Z�w���9 -T݅$��ԁZ��gN���,���	��*잝��޲���r��V^a/kK�)���C<�i"����cW��(���[.۞����6W	�XTȘ�	akl�h� Uh���]�$����g6}T���@���\����+�	f��LmX��uQ*���fa?�i��4GE�Jf;�I���Xd�a/��(�?D9��u�K͂��	�Ƿ!�����~���)D�Ag;:��I�τK�G?o�Ы�2Z]��ʰ$x���<�(�?T���U�~l	\�V�*�CI<M/H�-0-�[���ٙ�W����G�x�G�w�H���`�O�����G/�2�as�Ŋa��;<�˝���e����8+OO	 ��5�|-3=��=ː�}����K����;,��##/���;~OH���U����<��>��Ƀ�\�����V2:��P;��6��EV]���$�e��*;��̥2��Qi��b����b�!m�I}���n�yvu���ז��h�oap�b��,�!~�!�b׸7���9�og��`	�C�\b�1��[F>v�	nb���'eu�(j�^r�ݘx�Y��
��f���O&!�F�O��nu�h���TVz�A(M X?es�Ɉd��$�a�Y�>3M|g�$�nYOHdU�z�B�B�#W��y_a@��~���]V�;����r�>��b���8�3������En� �5{���D�)aL��֚� <�K�D��Z��7��(
��i�绶����C�p3Lu��[��7?���xv�M֑@s��p�mxp����
N��xLĽ9G�4o�����ot q
�p�A�ݭ!��U>kL�$}�n�'��@���	ӚS�����^Q��]vVE��j�����v�j~�2��f�l��<X�����MPbbe^�� ��϶HJ1#;U�Ǡ�~ �̈́TJ=�����l�v72��z��_��"U6[ߴ�7[	�3~����!xh|���sA����w�qKs�x +�Q�B���n�����t����^؜éD)�8�՗�N�j'� �@Sޞ��q#[bEh��]�)���*��j��
��؍M\b���ŉ�����Xo�ꆳQ���":2@ϱ�DQih�;~�y���L檥7�8����}f���K����I�nQ4���&�q�tÏ���G�a-�ܜ���h���`�@VV��*/7Q(Q����'�jb|?e-���gv�1k��	�1�}+`�*�ٚ�>�x!(��9 p	9�����Ϣ}��.�2BI.�Y�XƗ
��`{]A�/��א?�{�ٌ��Ҩ���K僔��oJ�T�J��[qZ�6$5�C|�h����x��n��/���:��)<]��b���i�Cφ�OkC�ԝ�N
�6V��I�A�ǃ�-^��8�!b���8m}4�;��U��D�[ܕ��ġ�n2���;-�5�4?�C/I>A�_��rJAվ��صs�뻪�~M�1����J$��䔭��˝խ�r��N��Q���zB�(�MRB���s�Rl��`J]�ndmqd Em7\XE��"�_��#>X�J���,u!~���q�ҶC
?r\M�/���в�Hk8�����MRl3[q��pr.3m�h&�n��\�J�]�m<�Ƿs�:��a<&!�i>D�4�/� n�=�N���g��;�tؑ�p�m���*a���4ctT���D�A.)�Q��!�#P�:n1�>�-����5`�T	���_zQ����'�Gy1��$��V�Mo �U�bS���2F.ؘ�����TmK��uq������z�E���*��c���`6,<��*�15]:��6�\��!fg@��f���ԛA�d+Eu�4޵O%�(�4��p[��;ja!{Zb���@�����T�a G֤Ԯ�RM@�u��tX (Nf�~���R�_�uk��у4
���K]e@#2�)z���\=���@ւ�0�I|z�,ɢ"4�D�3da�˅�<��l���.��˪8��H�遟���E���i�=�Ҭd�=]�똀��}��﷏�ᝬ��`�����I5�%\��i+�|�P�-ɀXf�Ѷl���}G���c�n����a�	��q%ûh�Iu{}�Q�B׊Ua0�%�v��o�z�yz� HS�t;��9�Se��쐾)��FYۍBp>�Ey��g=m�Z���.��5\β/�[;r��M�D�A�Jz�o�����X|N㒮��m�nT����k]@(���)�u\�擠r�� �o��Ҫ���6��,C�1�t�ՏI�*��|c?�љ9�x� �G��~�!�P9:l�B@����'�����lZ*]��k\Q���Yc绤���0��C0�-��{{����!���MJ�B��L�U��)'���:1�-A9C�hm!o��@aP���8
C���b���X���)���+tz���xK�/�S���ï5nE��]n�N�1���J�c:a�$�^8�yw�KD���;��q�Dy�t.b��v�!Y���xG�Yx�MZ]ϲ�R�o�v�A�TW���V� ��gCk�O]6�;�^tg-�4�Z�I��m	�Ƥ���y��4!C����b孋�I
D�n��zin�d�Y8²�o��M k�����z�+e�Lw$��TGg{�'-M�=�p Í5;�)	��4P����v�b9y�,;���E���Rۿ��L��_���%�����6M��2J����ʡ�JN�AgBʁu1{�g<Ns
�w9~-�8�24*���|��)��)�_�g���"(8}g������֛�h�%
V�{���h�)����O=�>R�rp��`d��2�x����5I��4���d �Ӷ���Y]�h%t*�{��c#����=��`��X���b������wX��� ���\zK?�<�*a���;��A�y�ZI��/�Q��D��XQ��Y�AE&p�9�v���b���$�'�L
��lV�;S��áj8�_�-v$^���҇�u%�j���Z�@�:1�X!��ɑ⯕�����/�Xh�Zy3�f ?jG�a=�F���d���f ���BL=�g��e�@��.^�AL�u�g#`ja�"E�4m~��׶�V����Fd3ߤ�ˇW�+;M]��� ��r�1<A*/���̏���i�<�I��-	�Y~�*	������r-t��Nc$돸�LT*,<��W`���rC۫G�o�k�~���v���x_�p�z��!�\a�?���܍֝C��{K]�r�{X9h�J���#���߂;���t��M�ǌ�[dn�G�V{�9��J<���$I5Y�y�����vp���kʯ*�P8�@�@���
װ��^��V+fX����/�C��|ŝ-B+)D�ŕ�\^��?:6�mDN(V��SW�J�?6�'�Bj�^e7����"�R���>E��v CF�+@�0����[����+w�OcЀg�6},.ـd�j�$V�d��K���M�P2y���2�MO�@��.��S�F(�7��.�Y%l�!5�#�L�U3�M��b�E�fq�<����8l(�5~x՟1q���tA�W3�A�d���'d^`QX��c���0-a_X�A�&?�0�1�-�$a=R	s5��l��%w����N�N�p|�C�d8v�}��:���@�������q���U)�S��}�7F�:n���]�3?���7<N�ki33v�jg�u�(��h?&� 1#��'�<9y��ٝ��_Ib���z~	z��Å뼈� /�슖����?diz��q�m�E���𪠳�esBʩY�v�KBd�eS��ݒU�����kk���^�`�ۓT9�"C3��f:-�E\5�񣮑� �q���)�c�Eذ]S��j��JM��q�>ԏ�Q���SRb�3�vK��-�`gO�&68�J�����̶�y��+��?#�y���8��{-N�F�%
b��! �L:��>�^w�H��K5>4����y�����ANV��
�PE�.��8ܲR��9��,Ltlq�����\����& �0t&�����"�|s�H��Ϟ�_l����JU���֪'%MXeV��ĉ�̓W�e|�su���غ�³����ٍSn�E �<#;��U:z����H���p3��&��aX<��{�
�����)�*В��է7N��3p����IY>�)���`e	����8;�:�H vp���jG���g	�jme]��\�R��qR���.���Axx�^֍G�D4j�w<Zc�$�(!�ScraN�w��o��}Ð���Ҧm?���v�{��������SeX�s�4��-#s�����~���z�=rF�k��4���\f�K*_*)� �L���hԁ�&\��~�_�":�-�8챝L����K�!�)J���Σp#Pr��U��|r���q'�������o�sV[�毖���r�k��)ӧ����ʤ�r0��D�Q�镝��L�k�7Mo�Ľ0�	�(&w�%��A`�gY��u}{��k��#8l��)�`[�,�$�X�#�R8p����ʩ���lu�](Ǉ)�W��s�����pd���(��n_��<35��iZ�*+�&��,��n�6u\�6-\�v��Rj��;7l#�J׏f55/*�#mhFl2bHX��� �b�s�E��"��1�s�����q�S�ٿ�.���`��/�/8��e#
��#�-+�Vu�k).Hβ(L!]���V���=��k��y�`��<~��9���Pewt:pqW��z�ޔ�g]E��xi��7��z"�m�?�b�y��W�3}���[�g�dWb���w�RJcN�sW�|���X�,�a����	�:�K�ٰ����Э�0N��?�����������P$�2��
j�����`$?d�pFGR 	e��Ek@TO��΄�&:��9/[@=�]#��,P��fJ�WI �h-ɩ ;E�Q����Ԑnh$[�r�L�~��fW� )�������0nD!�θ���1�Ei���N���Ia߈hQ�OMc%{jB2s��ܳͣL�|(\�^U:z^L̿���#�4���^����Kk�,�!L<��z��FR�UNܘ�/�"ƞ�$`|���ȶ"�M����`�s � �y���(C�ݶ�Ȋ���yf��۫��ӧN����}�<��X=���舭1&�Ҧ	;�f�G9�|������Ȃ���N�Et�DFط�4�*R�����Hҳxm� �7O����]J����i�}+7hh`�����XS%ҡy�=�

�G��
Mǯ�U8�riyW��f�CzJ�,4ʍ�(X8��BT>z�i%9� �|a�g2���@;u��?��X
�*���n�O���'�J��	�[ ��	���p��)����gO2��C�
�z~�%x.5�&⫢�!k�w�t.>�g�f,�b��#��R�`H	��Q�e߁��"�n"�^Q��<��1��V��̼.(,����53���7����T7�U*���N{5��w�H|"�-��c�x���4T|�@�ٸ �~}�de���*F��!��'�^/�i�Z8Ei��d��G�6�ɷ[/����$W g���nMZ�'�P�)���ކ�F8ܾT�m��1��{��oIKIpR��>��{�*�M�� ����I�"��0!����~w;��\<0��C��&��� "�7�V��q��Ȣ��m�0����3f�ݺ��$ׯE%�[%��E���)\���\;���l��#�p�Z*�b����[CEC�k���FG��5Ҁ�v���5�a�^�����Ł֡'C�y��f(!�`J�,>p��y��9���t|v^�>��Z���QBT��D�1ZC~M�j��}@ ��FuNN�z;����5h(��%x[.��{�:�]�}T;�v�qo$j��mK��ʁ�TX���@�8���S�[8i��)*d�{�ws�)��I&�'�L �Pk��W̧��=*t�|5��W[�`��/�h�z��zhX�R��)��HRt�FȰ��C:]=߶�����@b@[Z<�8=��b"KNi4mH8}�Nz��S(t�}b�)�12��s/3��4O��?���^}ֽ٦���?>*s���W�O�"@6Hnn�}C�a�V��$ ��l��O���涤��yE�м�=t$I5X7hYcBMtY<�!Z]��� >�a�l�����a���V�B��6��1��5R(��{���)v$L���G�@v�_��&�s%&�a#&��� 4���OJ�.d�me�s|������둊�8�rAȾ��)�l�����8	_�5+*Ɂ�QN��u`�3�B�\_ _�0���hYi�eN�ڵ4��2�W�G|���M g�NO~�X�_Y`+|��"I���`������6C�|��(���*��t������s���a�o_͊�#��<�Z?����T��)v�/�q�n��^j?=��X���Ac��6�ֳ��D�|<�|��)��;	_E��7>�����tݻ�m��ھ�7���m�����Ʌ�Y��k�ʮ_S��!�K�p�j��|���V���u�qO�B�3xڂs&�[μY���@�J�⨔!��m����$Ռ�ԹC�aT1�d̢��&(�s���������s�
�մ��/�N��逰�f8*/�o��|(��wG�+��O����<��JN��m3R��7�B�E�d`%EU6C�����Mv��Y2"�"##�B�pF?�|R�/ܦ��by�hA�P�/�Td��P����l� �ή�q�)�! ��xZ��D�&�̔�qU
=������w�T��5�~�7�)�D< �������~BC+��V�J������X�OLB��;ك:���P�?�/�=2�=��Nd�	'���"�N �	ѭ�@i��~8�wx�ȅ^B� �Y�R��y˒����f@M'˼'vʦ�~�M��s?���*� �A����iÌ��W��.�ۊ�Z�����&5�"5�u�³k[?����s�w*]!��Θ���Sś\o��j�:8�U�%~�1y������?��1����a�P�2⺽1H}�yn�TE�>�G���.eip���W����ZW����Yq��-���J�ʼh\p�H�A�_bX�,9�<eO���!�_��>��QOh;~Eӱ)�#10Ie���<���Ŷ[�xf���h�:��Ը���ߢ��
)Y�O���U��0:Ȉ� ʳ8ڍ%��A蜆�+��UTƝ�lX}�m�8z/&�(�|�h:ĺ
����m)s���꤉�{VG���g '��)۳�II��̢��"7]�Wr���qŎ.���D�6O��fU�X�X���x����k�����q�D	l(T��(�񄋢 �x�Oɽ	���`+q5>�}�Vzߘ�[�B�q!�/��<v�ǿ��z�*Q0������P_9@�s�Ⲿ�.H��71�2��À��5�}�rг@�L��f��$ H�t�HXo�2�"�yC���=.#��3�.��>�g5��C`�[D@;�4Y	�NTSmQ(L&�{5��|��F؉_�}��b���?ł�I��l��y�քK��歭i?@yḳ�wO.+��{w�w3l��e1]z	�<�f�m#ݘ���G��W�B!����I����>��i�מ,W�#x�g�{c�A6��'e'����l��T�}Ą)=c֫aF�v��8E����3����B_J��G�l����u������o�M��=|������������h!�i�Q�Jy�`_���ŧ�(^������ܓ��e��!��k�Vxn�>1%��OY��ў��������KgcWZ�S�t2�\��4�W6�B�K��V�3�2|�6c2�u��X�~��rMP������SۈXQ}pT| r(ާ��Ř�E�?=90���=Y��dn�7�,.o��f��V�( <d
�D]+:��u��`̒X`��\�;c��k�YH�h���rU��`���5!`Y*�1�>�f_����t��� �qHo�%��0�Z.��`q]���'F��{���ֻ����^����e�,gQ2�揃�;�q̷����7�7�*rd��FG5;��_u�D�-Z����BYTj��;�h�QE�/��֦=�"N;im���+{P�U	��B�3��P $�Y"�_���Yv��,ϼW��&?�8U�@�j�x���?�$'���Kb"7���
���o@���/ЮGr?Y�s���y|K�;��«�Ns�ؚ���-^.tJ��,���'$�*i��z�H�<��=Z�na&d��X"� ��d��(`R�;�`��mwY�@-O"vgVf�^a���$��+�na�7�PY���!H>�mA�� %W%ĦjҰ�ܥ9H�5@	 6��"��$b�z�m!����ː���FY�!��@=Ϙ�qm����YZ5΁=��nu�~�������c�AdyA@��l�#S3EUn���P ����ݪ�L��������;��J��?��
�P�M&埡�)N���~0d
�.�if-0�Ȗ�H|�B��O�EH��%� �{���掖�^W���:���_� x�W���;[pR\�*��E�i���\s;��0���b�p��\��/|��������(Z5�N� ��3��J��}���<q�;�I�l��Z a�G��}�����V���[�{kZǓ�9F��/ϲ��r�˶Q��̪~�8�h���	@�~l
��������|��>leC�^��W�=~�=�"m�:z�Fyv>�N<y�k�T,�*9�(9'qR'��e�4�8�Y�J�N\�-�*��S�跍��Tr��֐�=���ʝ�Dǃڪ�M��^k�������:�͓Bd��j��W>��;��lv)��Q���%�W$O����/3�(h_v��v��??�>V�b��js���B�6�5=.+�������O@� X?�y��d�h7���$����S75O%l�j��L��!D>�;��}�\�������f��^VS��X��K7�1�g����}�Z�3O������z	��N�k֙�~m��1�:�����P(!��*���P�t��OTw{[J���_vcet���y
o�Ve>�C��[�h�Bڬ��?���gl��A��z��%#*w�X�MN��qk���#��:($��SIb�z|I����/��@��D�5l�H�}�5�R!�
�$�m]���J��a����k,��hN�����>���7���W�3����C0�b�#{���g���r��d���7̖���&δc%ϳ�U���C���椠�+�"h��F6I��S��-(21e!$c�:�&=�%$E��WCU�L����e}�8�XJ	������Jg�g�Z"sY�\>�@<$>5Kl��T�1(L.�V�yO��?�z���0�,�-g�Eσ�:CI%��`G� E�v�L�z�}�y�'��\�FΌ��h��958��].����M>d��ǟ�wU�|T~�H$MW��Y�uix!��	��F��Ez&����o�`��$���,E�t�1�=;��+"4�2���(�i�g�����O�m�XM��}KB��n���õSwNb`�k�Ȧ�e������!ojxW(ZJ#`a(p��Ee2XoE�3N�~?��+��H�f�l}V���)4r}�+��	1�K��)H��'�!g���K�?t�z�w�38�o�pV�_H2K?�`�s�276ƌ.8u���{	Uk�����V�,��/k�3�V�X=0t��k�$�d�0�P����#l����1�q1r���\�-�L��@!�K��,bg|�+�5V�W|�Pv��V��+���H�Qt�f�BFX�֫�#��%���N�gH����q˲`���<��Օ��+�j�{u�@�D�DitX�&��4�_�r������a>�C��ң@̯���inSו��!!�]3/M�W���b�\a�����Ծ��
c��R[/�� `Chڴ]��M[���Yr�J����Ǚ��q{�$��f�Ӏ���JK��k���`\_,���#�$���^K�g����*����3A��əhz�\��j3d��m2��+:Fn2����>�Hl���	�BcԻ���n��_�����h�hO�[�M*��wƂ��_o$�B��v;r,��Z�҂����WK�1-�Ƥ��G3�_����v@a��~�3�m<̜Z�aϕ��}(y@��l���U~b�^s�Ge|)��JS'����,P�u����ɑ7Wc-@U}���L0J�J�Y(�3[?�PP���";���<�c�D�G1p@27H�KD���4����Ķ����;8%(?�M*�I�L(Զ�6!���C!����A���¡iY��:��������|aN��IR������h����S�}�Q Ȝ��B?@�WS�&�P�K��L�ט�GV��S���R�ɰ�|�TV�D���[�� ���Jde�F������Oy�(1#"�h�}���P�{D7�.j"�Zp�e��Y���M^�q�8���rPy�X����@(i��yҧ�S��G�2趘)��\��G�̓������{���5��n�,�w1�M2�&s%Bj���$㹬-�VUĽh!�叉&an���Y���|r�dSx�Fs� *w����w� ��ZL'�b�^��
_�Ю�̳�E���vn�i����{�[j|�N�W����=7���ʏk��I���CU/�axj��p'8�����Е]棉�&럺-]���
�oܜ�2�ˡ�CJE���2gk?�G��*4Μ�k�����ĺ�D�&k�RN�ԍ���ꭵ�>-SOZCӵ����'GW)��M���;��6�f��ĆYn�������S��긿����uho�g�����6�Qp!f|�st��T����x��P2��	PUFD���Ǚ��p�@7�>)ϥ�ĮTׅ����<k��閇�\��s�?#�q�n6▷r�t�͉բ��#�0���z�r) �S��.9w�W�����π]�Bx2Yfm�C[�-��(|�t�e�V֩�#�WK�T�� Bz	�W���� @�����ʕ�36�μī;MɨV���Ŀ�y��e�mh^�-���X��S�u�>��o�^�T־���AC!D+�bR
Ig����]���M	�}�K���wW$8�^4�Ձz�^D,�GM&���J�힨���=(�{#04%ڐ���`�"�w?�iA���e�v/�i���.�!���� ���=�����ET<�q��X?/^_��1p��>I��+��ț�] G	�&ã{	�7���}J(����c f�_��ܵ�G��~Jo79+��w�w�U�'���:c��8ӛ���XE�FM����$������'*���Z36K�L�!��M������<���`�N������h���F�[G��=��LX@���E�*$AW�TAQ��3+�� 
;n��x���	�vH��g@dӎ���W����'�c��[�-�<�E�����`���Ю���W�m1Qn�J��!��s�G��L�#ېoa<�w�^��E����1��,�O@�G�a�2m�J� '�:�I���b���r�keu�A�W��{�$'K(Ŗ� �a�LDeh����l���u�i�q�E��6��΅�V�c�#��/ڽ�ckh���~��_�!]�=!�$p�x�k������1���%���9g<zU��HѻӅ	��& ���csII3�����aE�R���
�FV�F�s�J_T����@%=.���o�!�މ�㕣Eۼ�_�P��Ti /SJ�њ�D<�`�{��-�㎔�)�C��M�ȕnW�ia�y�@:=z�bا�!��pXz��Я��v�����4�QX��M���Y�2+�w�Ǫ	�q��erh��2��uگ�*�I~p�1��/#ˎ	�<�I�o9�PI�0�b2'hM�}t�M4`�d�y@�{O|Ԧ4�n+E�*pC4f�6Y�w�.Ti���"�,l*�5 ��K�j޵��0�ݬ�t���Ԅ/E��Ё-�k�p�d�;�|;�=�K��oi�����:g�wS.���s��kֳe��ЭPHO�ll�0��RK�1�P�~[&��n�P=:��uA����ʷ�a�ނqt�8%��4إ@E�٫��Q�����BEe/5Wm�B鑗��v�gU���6��,L.l�b��S�~Y9t����
�����5^|6�x�l�;��xYS�Bo�&���]/��g����&<��&~2^t��l����K؟2
]oʇ�"u�Gv�t�0l�$�pZk���̓7�_�ͤ������H��|!Nn@�]�)�F�r42��0��,)WԨ����jvZ���P�0}�Āox���<T���
�|/7�,}�:�ˌYė9��2���-QC��XJXqScl�t�XŜ�L��,��_�er���2��6(�"�3�b&��6����t�k�{R0���R.�X�7~�[��y��lo�Y�����XK��p��܈�3�N����2�O���t�ݢ��ު���y�F��w�%���m,��؁_��x;�����s-�����-�<�l���lШ�	����,��B"�fZ����D�4��iTu͚����҇uһ!'������@�x��aNNi8�\U��<�]����:�S�b�D��I����y�T��++;�@x�������N]��'�Ր9N�����ؘH�vq�S�=;���	&3'�j�
�������ڢ���`�@֡��]�=$9̫a��uѫY�V!����N����$#�J�-��K
�L|�|ag� ��e4憳+Ѐ(�~|�EM-�F���x�FCu��0ۍT�pل_⅟_lQ�`i��"��ry}��}\
,�������9�@.�xѕ�6+k�W&֔��i��MC���bk��$�Q��dIܥ��~�]d7�������9����v��Y�:T���9�r��Ш$��{�E
d7�x��Z��r<���!���ʅ��7)4Z^���[P������ֽ?�\JE$����M<��|'�������Ó(��x^�@�|����$�C�L6����Wc�?Y���Y�`�#��DL�����'� �x�Z7�]�@R�}��B���	3���oS�c�&a\�B���;$�)(b���>��f胢�P�>w�D2�A�)�嶺~�lZ~�%�d�8��k�������g�Id�f���SS���������Y}��� +�>0�ڕ <��b2�R��v�-��2����p���D�T�8T��PiO�%|
���V���6��z��4��*��(� ������XCE��q�a��j9�ת��B���ft�.߬'�����7��,>.��;����S����r	�15�=��H�(K���f*�������Y<3�	\�P����
.2� ��
�����c$u+\=��xo1����͆IB3�8����y��33_Z�l��,�[4a/lm��7�����ʉM F�:�#w��:�ULF^D�� %�^l�TDݤ�ɵ��s���`��i��%>x�:�2�3j���X. �'���lj���%^�����7?`nb�e'�{��4�S��t����AzVK�*"n3e�P�(�_��_��;j�d�Kl2�;i��i�Wz�Xi�ҩ�ʛrΗ]�:v�
��`�XK#$��%����Q���G��9���:�԰`������D�I�9�=��L�A�y�SU�os��X��lAy�ս���,2cO73�図��ц{8��u����c�R�+`3l��W6z����_��=���aZa�X��XUo��� r��@ NPCQ�z^��N���DX�vfDew�b�ha��[X��A�n2e-��!�9�1"
�n�0��Z@�1�i�Z,���W��������s%-e|Y�$4!��eF.��p2U��5�{����kl��\�$�2y�(bxn6`��0��p�Nw�y�f5� g� RQШV�:�2�T�� h�=8b��y�ѮFcE^����a�8$u�mF�h�`�.%z	���]�fѢ���U�����V�9�#�(X'����	d_�*,�Ƞ�z.kX��^��x��ϪVFM�R~��5�p��N�j��cR��^o��cF`l��Y/T�J�.Y�&+����n�í/��,e�UF�T�*w�J[��t�k	;�%5ǖ��׮���-R�l�h�b��L�e~���m�^v3+��.�Q��=Nc(��hniӲg�%��
[$k?܎<�ЌDo�>�b��kU�7�v!�p�����%l/��k)���b|�����TK%xJ�j�p�7���Rc����D(Aϛ�(��U"v#��ao|�E�-�n��њɐ��Cf�&��JO��,�C�~��'�șv���a�E�W1R�<�~��C���u>*mS�?��k���i~���K�J��m3u.��<r�r��!�?"P����$K���~���@�V;F�R�~i�=.޳t{t���İu~��c�{�rV��U���S��NPD���P� \���|+�8���U�[��W�>nK���/��rT@�\/P_��{��d����B�A�"�)�|���!����`�ie �9��YZ�.����+M�Ҁ�K�	k�k�Ǔ�]�#5�f
y���I�͍&�Wy��B5|�G�vm�1�k��w�*�y�_���L���,�}'�I�x��Q�	�5�,�m�Z!�;z9��?(���w�^7�8ܦ:��e����b�#O��h%�1���C�ѣ�����9���U(��'��Gmv���-�oS�m

V@ �r�|�h���	H8T�3]ЅN�;�"/4P0�iV〈ǫ�tg�+�z��1	]=y����\�!}�IN�"d�(ێ��|�:�ɫ�yMh)��Tx��� ��;~,ٗ�]1�9S���4+��b *�¾#/�;�?N�x���X��R�޻1��K�_�=�i��?�ƞ�BU56�u��*�5ŀ���:{z�,��O!�7
>�sL�0W������IB�P�Q��Ԍ�]�壙H���Q�*��/��Y����'N1-�`?�P!�{Խ�y�(��2�Pd%@j㔖��jF-�,U�3͆o��׊�!#J��r��ѯ�t��[�M<}RHz{V�j�2m��ѣ�ڄ�S���y��H�Ƨ�D.�T����Xv��*�6X tu��>+:�!�4*VZ�_oރVA׈#�,��'�ߓ悆1��ȸ�����>4�\AY�]t#x23�* �#m�b"�6H��D �����	:��J���k���ꆪV��_z��-��.�����v�$���Z�++Ä=�u��i~�V4��u��"V=��������2�}|��3�5��]�'ㄌ�}y=�Xʀ�7�o�]j�rR9���B��故�8�\}�l�]r����b��F��<�B
�ڝ��ټ#��\�n
x�1m��G�d
t�,~�I�2+��9>I%���:6�&�,���ڡ��p/O��t{�X�wQ%�!=�v��#�N��J)�^.��!�IX^`0>05-�u|*:�b�=���=_�����Z�N12���.�o��fVl���1�yT\+��2��x,���EqmQ\���D���&��J�	�C�أ�.�:ji����?o�J��͕��tIQ�dԞ֔��S���w�h���[�#>�T�#�S1P�����7|��M̬x�f��i�"&��Y��t�L�Q��\i����k�8��ܬuO%7�w�^���>p���P$e�������`�"���D���x�XA>�g��U~���j?�˃^�aǃ����V�9�2u�9⓪2+m� d�RP��5�ð��#p`(޼�N���M�_���<N��QX�ι�29Ð�1�H6�9�Ϩ4;���qH�y��ib�R
q]*W�ul�Z�4Z(8� �)�B:J�@07!��HL����\��
����}$j�ܝpa%����B�f��Ϛ�V1Z
�P�"Μ^v�F��5	/,�X���_1o�(�z��C7C�Ŋ�.|w���2�q=E.���%�N�œ��t�T�^9A��W���O�M���N��%f�ͽ�s��*^i�p�j��a�:�3!K�z'�@jDq*��hn��&2A��w�ӑ�E�(�!)�1LUՒXY���R�����&�sw��R�CTcL\�C����` ��<@v�о �.媚���W�͘8,d�U~\�	�@{2]Fw2��f@9��
y""K����B�5LiH��K� �A���!w��4�E�����22�ҝ;rr��j�)-]3ji�a�����ɿ1Q�1�]���
[)��Om֐|u�[#�\tf�ض��+�M_�]%aG�����yZ��c-��N�}�9�좷0��3.Ɇz.�/���Kuu>\O�9;�"6���#Q�V�d1d`�_����%xp2�m�[1��sС�+��yf�7{H��XS����gD���7��sK`x�ij��܊��<�T�/UB` P�ړS���9-6����%��E�ҜH����n�`�-�p�KE�v^�1>8���#��.�]����:k1"	�8c��T��՝s� ��jh}�y�v��?P��6o(��5���6��G�f�F�N���z�FϢj��cq�л��غ�``�2)sSz9�$��u��(��L���b�8�Wu{�!}��^W�
�z4G}��͇��h����r�a�M�>�3�yȝVX�xM�i��y�I<������j�b�??$����T.5����>R[fvݩ���4ʵ''o�u5C2�����6 �~{}?�5Ë;a�4w���a�$�
�@�����Z�:%(���Ut�r�a��	�;�w��\�7�g����&j�����D��@�+��#�Пrf~�/%��Z����ʴ��˫f\o�ب�ڑ}*y_��*��.���ns��X,�ޑ��4J�x���ڛ���V�ow���.�m�G���Xԣ�%n��/j��W�.�`p�A�y2T��6!�h�Ƕm�&c���̣���at6_������}�V����.{`&��Mb�F��n\��4��{��N�t�?�55%[�ҋ�t���X-S���S��Q$�����V ���tesb�1B����	s��Q�	P�N2UT�􁪀�x�mdJkz{x'�^Z�ҐP��b!ɝ���_���[����+A��*�-��=���W�H�^ndw�����[t(��/*���K���e��^��	�p�ىo h�c;��g��z13���v��Q�3�N7�	ҙ�vĞ�-i�I���BQ�t�/}h6{��8Z�v�pN����^X0��Z�&��;U';+r��0�Q;m��7��F�3\O�U	B�j?&g����g%��!Cl2�ZYg����ʔ?�@�i��,�""�F���~|6|V��~UI������c�Iv����!1N؝EBZj
��0p������켺��L]��֢�:�t=�[zdʩ���$����[���\�����
��t�6,�������2�.��t�I��df&�N>��AӋ��yB�$�ǯ���@��^I����m \m�y�� ݃>2�?�Fq�b⍣��ҳ`�����!����I-;T�-���¸������kL-9|iR�j���^e�����s_�v̓Ž`pUS�Z;�����r�n3��L�ƀAp~��k�� �V��Z�iV\�7���j��8�xE���ݎb�i����
�n���
��7���4�UW�Sxdd��0wy[f#�Z�-G�"g�l2���3 �+#��RVkN\�׋�_b��E LQ 4�� �/��NM~s�2OvW�wRL8���]M��j|�D� [j�%E�v�+	�=�ZP�'�Z��m4b<rE2w-ߓٚ�XW���j�%BG�i�Z�F�����p�	&5��Е�W{!���m�f�lY�r7�=�l��l_OЛ����JSeK!������ճ�M�ڈX�X"�x�� Z��&.c*RvGD�§#�[��+/� ö�Juw��,��Y�@x�N8�M-�R(��r7Q�������� �'���h1}ۥ��P�L�w�c�𒃴٭%�r�����_��y�h[Y���YX���D�\C�|��e���C0H� �k����J����fhz,Lt�:�.�ĸ>Z1�ouw���Q�;��_�:��,)�����M�x�H��'��{Y	�Bz��Bl�,�WR�5!e�6�*�&Co��������'�_ ��xyt&��$�������}���S�P��K��&?��s� E�i�P����� <�a����a�nr�XE��Qbh7��"���≁v�,�N��S�m8�=HUs��.�dͧ^XT�u`�k��
�ׂ8��Wꕑ�O},JO)�{ ���
I��PZ�YN��������M\�Ug����<����&�m�٢��8hh>D.��t�o���m�����Gc]��0Z|��cu};�o���c��L�&�
%,t��QiCw��p��Y��̺�;��KDT���b���PAh?DP�Zz6p=J�^������pBOۗ��:����r���ȴEE�4�!%�S�oI9My��1Eb ���(�T 
���/J��5)9��Ϯ��D�Z�`�H��$���м��i����p�@������Fb>-e�&8��JB��� ��Q�������Ңyy�1敩��;fP���Ʃ�tռ�2���﷌�6��.��:���_�����R�1+Ѵ�h0U���Y�'6���\��Q��Ze�R� ���ꬭs&�ڟ)�� �%tM�ka���o(��F�r5��d�͏��t�����>��������9t����e0n7	-��W��!����һ>x��7�en�˿���`��KoN���\ϭ����ӓ�놭�\��(� �-��)�Ȅ՝ad���Լ�a�*���'Kq����8��F�]R����/$��իN->G  R� �J#C�y����w�H�j�,��sC�%��p>kTŹ�v���'�Ҟ�Iv��bX�R\��(vIs�bF�$�I�Xs#�>넶^x��$�餵�����.p�S{�Єs���l��GIYP�K�Q��|8�y��}�(��C�^EFp�j�7U���c����ib�-߀�\�i|�)�l���T�Ӭ|�I���V���r��[غ#���K��'������^'�!B��O!�k��zs	��^m≜��q�F�	Y�+�����&/�?|b��a鷨]��0����%kWjO�����B���;�u���¨
���!ó��w��+��(Ǆ����1(�E��(���Q�ײ�@�$e@/�:���=�}|x�З�c��)bhS%���f���$󧰔4�6�;;��oh�a����%{��U��,j��(�Hv�`��ۚ�ȤT�v�2�YduGv$B,O:l���v���w%�~yl<���~��X�7��g���q�<:�:���,�W��F��mb)�_�v��ZJd�m�~�g��*15����Y_��8��9���"ȃ�����5���ީŰT�v=!��BW��pe�X1�gcOr ��|${(s���~/x��D�濯	����P��i��d;����┩����C`����b��9��8H�wY%#���]��:�s�IT6��S��|���i��O����d�̑#�����-��R^�th���:��t�/[8�׹���*���i���r�����]
4���֌�܎�#H�l�y�Q�bC:�ƛ�姌B����v���F<)�s<iE� 
������k���4k�ߦ̵O4y�s6�
����-<���3W���}�x�z������&���	^��X�f�/�Q�S�4����r�-�Ib���w�S �Di_?��W��\��RAi���jh������is;��`���y%�L0b!�s����|B���S�CB�~�a�y_$�O`b��o]�w�x��%y8Ѿ�i����E]ѥナ�]IO��C�^d��,A߿Q3h�L�BPv��ƕ��L�h���2~�#�Q��!��
a'$�w?GF\Yk���A�t���v �OlF�nx���ޏF���� ���%���qS-�x ���G)�:^>���K�h"�J벱9��!��N�9�Q-�~�Lf���H��t����Ȱv(�^��r(�@Za�ve��[�
�K<���=HJې�$�����L�m��3��<�HAm��}@���gv��z-B�����F'e���F(�v0e5m�q���h�!��g�[r���>h��x�m.އ���!�9��^8�ub@��˷Bm�dZ�Z��q7��e���Ὠ{D�ˠ/P�ｂ�N�+�9n�߭���2��.(�6�2ηO7��.[�� 5C���T�F��{��xEL藳5��C��^N�� �kd�Ҭ�A����u����a9N�H�!پ�T.Nv"}���)�L![�K�0?�W�DQ�d��U��� l�|�؜2{.�YE \���(�7�P��
[ ����VLp��P��H��z3RP��%��\Ǎ�O��������:~�Kd4��D�=dO���+��o<�l��@�G��X�{�(&+K�#�E���S���M!�j�S8ȍWMw]:B*��M��е`y[�Ԕ�������?�����-`a��"Ph��Q���P~o���d�����w w܋$�&�1Z�5I��2.4�B�ʰ�9�O�����+WL��mF��$�pv����%~��b�R�C���Z6qd�[�2�+�-Pb)x�}AG��M�U��6n,�<$��Uy>��-��]Gf8M��I������,�A���~�LüIB�eb���uZ��8�C�7�݇�W���~�W[Ǟ8 ��JF�S!�T��O�H�<��� ��-��bv��C7�0̠�I,dvA$ΦmlX�,�U<ɞ���:��zn�G4�3_��?�����4`��9.�����餌����-_0��,�� ��4��7�:��M.\.�[��t:��%�E�=D��+�Z@��U0�����G��}�����D�\��k��X�ŏ̦��E��i�xм���K<��
��;lB�Ti����(������"܀�<��% �3t-��M��s�0f�h%�O0�k�ۚ��{�4kĻD��K0����D�K��q�Ì"�Xz>�7r	Cd��j���g/��F��构�ځ���b�/52��	�4T�Pn�<��Ѵ�*�u��Mvg�=�����_��{hsh!�.?���� �s��E@��f��R��?���2�c����sv��A/��I9���D�7"�q�tg�[��,�[xf��Ū��b1�Z��[fB����t�e�P��s"26_��WwA�N��{5r͢���4�죊��$m��'�� ^;A������\l\���PI\�S{8Ի��1�ْpY�2paN�W)��a��4�rM���������ˤ����8�	�XjP������%�<���z$n�T^/}�������:AG���4�̯� ��Ss�XN���ͺ�8{mbq�{�l;`��s<�䲈�K�2�����Qp���$h�
$p��5�e�Ntk�B�l=�=YS����,�W�9v�f�!5JO�{��n�aq������3��bt���NT������P5΋4��:
j����!���UQ�D�+�w��݃���ϰ� U�����~�R��l3_Tɗ�rrb��w�~B�9�o��{�3�#�Oo��o@�kPQEf�`����ni`������<o�Iz"zA?�ʥp�}�ި�D�8(�STn�B*���������SV�s���v/�kÌ�[�e,~jQ�yЕB���`f���jɅR^+���-E�������
�0@`Ԏ���6P����*A��J�Ѱ*s"����=ç��rt�J�UTq5�*}c��x}�˂p�x�|��_�^�!�t�(��X�2�YO@>�?�q�g�R�w�*kR�F�c��=���;�XU4IL/C$ܑ�o�o�s�ه�l����QmtȖ���v���tH}z IE��������<���j,�X-��M����L�CM{�WM"q!V����Q|���`�����s��-���� Y4�܋eB)���0)v��[�mJ���A�5�o-9w�S~��8�A��RlFXJ-��H��}f*��fU_�U
x�y7�f�-3PDݘ�D�X|�a�d�T�M�(�Na��_v��mI����m��|���PZC.�ko�\�������ċ�0�/�~.�K�O�\b��_7�����t%�C�[V�c���/�f�i����j'4=������`����z�Ķ[��睈�}Z�,�"zq8�pO�`d�����<f� Ҏu���8ME���z}c'�m0؟�Q�{�GE�����E��}�J�%ᐙfƓ��B��  Ą��mCY^&bc���4��8z���z&�n���<*�-�A)��G;T_,�0JV���0�׫]FE>�	�;i�`?��FM	�-�t�K�n]�IG���!���4(�Q����!�z�,�at��{g����p�Dj������ͩ����KK7���,���S=BF�$����66����z�;���[��w�]5f�҅��9nZ���-p]�|����jPl.,>��z	�2�m�B��q9´�;�_���U*SX,y�R����x��8IõX=aس��0�u�,�z�����'��[B˝V��Q�PR"i��Ե�/��?�Y�U��;��Uc�̨]n�f�e����0�.@ଢ଼���d�aR)�5���3�bOY|��|��{�������,�����j��	�pM�&�ĖJ������"Dr�G�V���H}�>���	0�u�9L�����<i�0��iG���U+��m�E;O�.? �脅Q�ҍ7�̔~�0'���ۤ�,�wf�<7�On]va�u��3�sx�4��W:���V��D�f5�u�yY�BUl5�ج�u�����-A�Ф?.��p�]g�����5m#2��:�垍�RY}�b�^M��?�o���:��(n1�⪱#�l����h�������v�X�#h���=���U��uu������� ��$��<�ĕS�bC��PQ�l:W�����6�Gh�S&�3��xx��^�]Y�Q ��!^�)|�rfFJZ2�j˝Lߊ��C�G�ɴ�O��YVh�l��;ɷ��{ڄF���^�U]d����Ѓ5/����=�CoP�C"��e|��#�F	8d+r�&�a�\H~�ӽ���g(0�1���p6�n̬j&]y����S[K�GbW�F�j#��O!���{�Y�|#,�07&��V��񽞒�����"9ڽv��+���p�"AyUDV!�s�^o�#�gS's�_Ԁ��Vg��Й�q�m�i��@�{�Ɓ7�ZݫHy;� }"�'|��
x#�%4!������I �\�II��E<\��E�Ť3bvcg42b�Ua� �W�����[��W��hmYu�Q�OK �U^�>u���P��2����	Atӵɐ�&yYL�h:J����ꠚ��"�0>���)ٟ������B�ЩGR�TK���C��➣����v�����F6�,$�#�$a���*�=�+τ ��Q�=�[��BܦM�PA�T�v�J2� ������I�O~�a�����b7_��P���Drk������x�T��;��b4��P��^���r_2	���_�Z�3���Y=�~�<�U�M)iϩd
�_BXe)��rX2�j�t�T��xԧy�"д��dk"8L5У�ON7p:ے�!�]>�2r'�5����H������4�p�;X�i��x)WӾ�v���&��|��h�L �rROu���S_݆�ęc�.:���s�u�� �]o%�]�M \b$�9Q���ղ'!{|��Un���r��=4-��&��E�M�Z�7��S��_�`��1��a�d�;�8�@�P������.�� ����_6B���r0;�,�nI|��j7D��wg�`~�Z!.]��H�����	f���s��� _t�L�
�PPX�=�fx3��	�,2���y�x�ܸkY���ZB��ES����l!C���܋]�>)xҦ�?]��ɂ,�"Q�L�Zj�P6gֳ��L���{��=�J������i#��śM�c=�w��<4��ޟ��W�.8K�bi��!(㇕1���d�	�T!_u�"��TbpʠXI�Z�Q���B�P�ɋ��R�)�ba�Y���|�.���zQI,��'�BMʔ�	�c�C�:��C���z�wqke|<��G`	'����2�f�@�ŧfc��TԊ#=mUл�U/z�#ڸ,Y�>���0~/�E�.5����������	pFu�)c�f��1������W���u��L}iH����[�KI���I� �7��Ɓ��s
��J,~iѫ�;�r	䌁ׯ�zK��|9¸�6@�-�&�#|B�K�&����^m	F}lBx�p��o�w��ۣ�MQOT�drW�o�Q7a��D�����Tky8��&��"����D�1f��\��F���U3�}���L����i��u �����Z���f�U�uS�}�Z�Dܒ<7� J�2�#w�)���W?^��x
��fE�YQK��%�Fy{���5?����L�Mۘ���F����D��ø�������� ��ɠ2itA#��h���07hyP��f�w�)1K^�c��L�jȑ����G�D,�~Yg�)��݉j��o\��M��������u"�����v?".���a��[H	��F��?�۫�}�]�S-�+��^\��Ż8��{��.�1�[����|��+l5��ł����l�ztsuİF̨������Zٰ�K�֔�N����s#��,x����XI����e[�xĸE�6�f�]�a?��Q2�6-פ��T�	�G<���"��f��"NئyŌ��nmH�Dd_��`���j�\i�ǂ�⮧�P��j����B��>�٣��=�2!�e7�F�Ьܫ�1&E����ވ?0|O�X�(�<7�;���2*���B`��,���m�@�Xŕ*G�1�gr#��ĠQv욜+����$��`�6L���{������ڻyɭu�ٸ�UE2�;$��B8�Cr�
�v��Ғ��]�>�:�_d��s��Rh�/�3򯪰ae�%��Ϙ��{�׀��l�XӼ{!˜��G��;_?xw���I��b T��o�s>��E�_Sm���Cw9�ܬ����\��졔���O�ڍ[�ZLL9��+�X �D�I4}����,#�u:bU㢵NAa�hC/�t1�&&���z4��n:�]������G}�P(�*�����Ki=H�ښi! 
B��*�kY���'�G�l+���裵f��)�ss���sRB4R2���F�L=m�|gϟ���.B��,P?<=)-�6)Z%�=ic~���m@)W�OZ�q1�ϧ��͌.#��6����wNw/F�1�yJ���
��Zv�o���[QI/�j����qK�r
�?�yS1 zN� �?�Th!�ݕ'9���%�cLH]J=�O�{�EX�T�@�8=<��F��5N���WLE�J�_)ȁ��w}R
���Ja�r��	�{� �@�m�uf�I���M+��L�뷉�c�?���ΊܤJ#t����b&�TfG��Z��V�*� B���D��s���_|r&+�X�o������>�9PQ.i�M9��pc���w�5|�
����+����/09�Q��yXb��?�J� v���)�t.���l�,'�*if�Ⱦ�u�ƞu2������y���4RX
de�-����_�=t�l��T�t���[@�dz���V��c�ĩF��TK��ua%�u��b%��&>&��6�w�:���ݦ��~ �7Ӓ��c��S^��y������<�R2#���?B����	o�	{�l}~���vz]�+腈�����^F��Vc��4��������w����E$(���M�^����p�W1\��q�s�5���&�Y��s��Ѹ�|�N��OU��ŧ�u�ӆ$L�|J��"r��Á�)�\eב~����ru���t��ie�t�}�O����C���2ۅ��K_�(�NHkJ�htc�@��d�|1r7�I5��!�4��\�ɺ1N�Y9I�?)l$��ƋD�_���WZAU��9�˾�9b��J�6��ڋ�?Y�ӔD4w�Y~I��أti�SgĎ'�A�I��m��K�����=��]�Ncō�%��I;H���8<���~!�4eK�G9!���񺂖d/��3�,l���
�ua��+Hf*Cr���DCK�!F��y�G�w���1�h/�P4mN�
�o�ȑ�z�d�g�$zk�'��7���\��Mϻ�'��ɣ��S�3��`c��Ht���N���f��ټ��EF�]��}����YَKk9m�s�՞�B��~	�s6\]�=K��wO�1�b �mЪq��O�ʦjA�@5�{���lx� ��M�#�V��w��OxU�O/;Ԣ����Zxt���D�q�dy�ysp�/���b�%Rf)/	cG9B�BD��i�͉-��E�3��g0�&?-.	��r�v@m��<ޫϽ�6�R(S\[@Vi��6�5��S�K~���#�yOw+c�铖l���ǧ���e���&����f��օ�K���x�dH�ߔ}�Iս���6qO976M��ebT��a̓�ojB`�߾M��yzBB�^;=���R¢�\
P�DN;`�>�.�ϵQH{����ˇ́�+��HHd�K��14:�Ǹ��pq�"�p��_��TS�#�A�0�0�x�-��Q8UhS��`w)���R�-!�Yen A�0��ަ�.v�pV����QX�on�����%�rqO���S�"a�LxIK�7��}$��O����,�KȫB1��2R+mgj��Mh��b�J#���a)��e(c��.P"��}��o�乮&J���vx͒��Z��V@L�����)��tRnF�3;�1R)�?�NPOڭ�6QX�T�ҷe�d���g+Y4\tI��R�n�-��S��beT1A���>�Б�\b?�<�cW?�m'�1�E���q�G�Һ�k�C����%�Ű��!�3�D��"���||��v�_�n�ߟɗ�<a���]�H���7P�{@%�{Bb�����lXvDL'SU��b	�j�}9ԞA-�}���_ㅓjF
�߈P�~�S$�ڭ	�%Hu�~���Omz����3��#*Y����/���֝�l��W��Bm{I��_�63^u��~�?a���"�ayv�"����6�(�0R���#`�a��&��+��bϛ�K��L��jŚ��8X�+�<�K8�	�����.����=:8� ����jy��e�4��?]2AGG����D����x#�/\���˅��i�'���0:�]�x�ϼ�����ˊ�v�D�5l�V���ΧqB��=R��zܖ�Zo/�ٕ�L���J[Ճ���<p����𓲩���!-�/q�^�,���/��͑L��fͣC4�^"��I�+��~�(��0�R�#�R�R��ܦ��(�Zڈ�	Fc������@��M*�eu��]�*��g!��Ȃ�{c�o�
ze�M�����ɶy�R
��*c9�����A;��9����y�H�;�L�!�ø]I�F�y8�?-���c��
f<0tL�Q{?{�@�m�3/�,�;�˝*����C�뽛_ Y��KZN��c����.�A�XY�C������al��φ��(k����/	�����Cv��Y���;	��߅���֡mg�Vܛ;��K�2Z����ڻD����<�WH�;��o�ecN.�N�VGzZ�a������nJ�n\��:�#Il����k`d�F{��0j��֖^����l�O��{2Q�s���s����w>ۋSl��<B�0׀�u2�I�%:hUp=ae|�~�	2Ch5�\�~�>N����7χ�("�������UYD�B�9�a��_��������^:I��s�g����0yQ������=��G��*j��ɕ�Y0��w���[0��%7(oӇ�^�7�ߤ�y���I��[�$s������D8����yi�� O�k�� ��"��n��O��՜?��/1i�O� �$�}�+��UU2ɢ�.�1�5�|��-7����Fْߔ�.�D��:#�\��-�����g����q�ӆ���"��Z�ή�/pݲ�AGEޥfBm���;�������6x�vf��r���B�Cu�ܫ�x���5o��W�q�}-6Ζ�d�ǟ�r$���A{��w�)3
;�����\i6])T0����Z#F?�G��V�7�Ij�WϺR�銚s���B錅LG�w�xr8��s��z���/0q�Y<��fafy�����I�9>��F��8�J�gwL�Ϫ�G��ױ3d��^cwZ��>>���Bb����$�o���
·��U+����~�O�	N���\��jzJhl�/�ZJc�MB��n���峮:� �+CU��#�O�e�8�5}����X�/��O��zP��|����rS�8dR���[�3�[C5���Ҩs+���W��>�4�+`�G��8iWRCeI�r�B%����(����}'Keh.�� D�XX�Bۙ�Q-�ي$�����2j�#�;˙P�����6�Myy���3�K�� a.�h4UY�W��dc�~g���_��� �P�?��]ڣ9���Ч�KaB�ϖ��|�����G�(?��פaH��%-��G�ȩ�o��I^�J��y�Q,����ts�ܒ{����#��-��n*P�6K��MǙc��X��5���PBɝ1��\$\�oW�]RM�yk�/�;#o-Ű�栎@-yx�1��&�����=���g�X쳣с���L]�=����1�����eN��P�^F6ʅ�sV8� Q�N;��������d.�)�O)t>���_����I� ��{�hV#.���T���f���>�|~���`pwò��x7|��� (�t���ރ[_��"��Od�1S�����k��%�A8�����,���,�}꣦(�Q=�3Mt꒭e��>"��6P|��)��w�N����Q����z�w�F��:�!d�D��i,\Ө,d�0D�t�߷���61w��������q�ԛZ_o1��v!J��^2©�e���j�5���.�a�e�)bi"������Q�me���*0�K�uŔ��*�:7�J{��EPSr(O��zJ׭��ҕY*�7�Aq��^��;������׌v������Il�a
�3�6���t�b�f^�`�`x��CT�Dg�1���(yR-K����Sv'�/vr��G�#�y�\���J���ALq��\�$��=a���Bq�d,�<�2�����J.�'���2atUq����V�f�0rhK�T��������X�w9f���#yMR�@�Rb&���|���o ��� �5Q��7/S6M��mw�qB1�� �~�h��^��HH`K׊���v�ci�n/��ě�y ����4ބ"H�l#�쳸;Fǯ8���v�TU4aR7[�	��w@Z,��ف��m������9i�٣�I�ޞq$/W
=�P���6�V��"w7*�E�`B��(�{���`���H�É��kd�إ�p=5�Q��M��o9�$C������ �(p"���m��v�4֣�O��\�s+���;�ɵ�_��-����^4&��Y�#���j>���p/!�"n�|MqTۜO��x���0{��2;��{��C眷K�j`����s[�|j���8Z�򵕅H�yy_��	��s���E��Ǧ}[ڢˑ���3�����~��=������v�#�[đ��ݟ��p�`UCA�F��:�XP�T-��� �?��W�A��Ȥ�*O�{��Q��CG$`��7N�yf���5)��V#�Kv��z�v����P�|��d���촛�9�GI�B�X+�2`3�r�yHw옖���kĳ ���,�S���/�3���D���%.x|�+j��K֟w�U��#�yHv�Ӄ �����qR�j�	X��$v�g��f\2��7�qf8d�R�Y��(%��7��,��T��?{m5���z&R��+2J��(ũn`*�`���.��M����OD�>6��d��9�#�\vK��Se7��fo8a﬛�r�\���~ſ��!��ϻz2�guևX�Pq�3d���4��7��?}�K�r2if��J��Q蹛>��1�u�=T�ŭb���_����Dy0�@�-����&/?�H�x>��7Z��O�����3kv�dD[&��9q�ޥ�������>-3`6Kd�.'�}��Vr7B늩�y�z�������2�"�Vw����VIq�ę��WYʲ9�6Z��_	��AJ�S@,!:`5��.ڼ�5 ��~2���iYS�ۋm&��%���#�����b������i/��|ҕP3�մq���LRN[��{��[/�����v�Ã��awq�&�@�(Ϣ�B�a�e�3	پ���c(rM,f�i��W�V')^7W�ut|��M��5��=��|��{"���~5���@�-�y��Uѡ���9�I�s'�j��Z���HX���"d-��r���DK�'����B�i�fn#�5]-��e�U��<�����IQ17t�ݯ�ƹ�I��̓y`����c����Hk��{S��K2z�J��G~��Rx�@o�>��	t��@�����Im���@����ԡ[���91�����4����D����ϕm����)������}i�jǇA;��b벡�lWK�0�����埻ʼ(�@s�Ջޛ6�C�]��b���$���࡙ܬ��&m����p�p!�-�W�ٸ�(�=�0�V���A!5m�_֞8d�g�$~G�'Ȫ��]����{�� �P�1�1>C���2J�[�G̹���@ƛGQ���Ͳ����s��H�P��0�f�Ih��ʼ}�r��lh���~��W}c���5x���&p{�H�������I"�HVR:c.���;`M0��n��jJQ�P�M����ߡ����S���w�&�*�����4�Zc~H�ZXj��9�t�'p����h��S�%Θ���n:�m"qe���!��x�y�E��A��=�j��ֈ?X ��o<��o��ѻ.5g���l"�@N�sv.�]�P~tpw;��=�N D^�!� Q�%[c����^��-`�%br\��}�-3	n��p��#�L#�S��.�h�-���O��F?��0��l:�� (�N�������e����-U~��mq9�`�fk�ΔH	���my�5	ۤ
FG�/R�h�5�Gǒ<ѕXڦ���kж�bb,�2�KL� �1��}q��o�\B"ZÆ�u����(��� u�m�=�7���g^�)��J*�w����*h��h�K�hQ���e(����٩:Z�si"�bw�ƍf�w%�_���(�B�	P����O�w��@�?�����A�3���'Z���=5�xҐ�����9�Uɔ�]�l��s}�}���\�U�����߀��*�<�Z\z��~X���M�M�� ��O,�Qd�DG��P���:5s�爂��w�@͙�j0}`������j0�Ɋd�5�X�a�
�X��ԇ�
t�HZ�y�"�:�-3���ձ|����E*�q���$S#tkқ�N� ��|�K�� ��X�pN���f���q���~|���֙f�+R�b�/4��>\�G��0���*�L����L� �_j���Ё�ߊS�{�!�H1�y�'�VF��f�-��-@�0�����a� ���H�Y����W�ȉu�Xp��h {��s�.���w��q���hAǫ�ӯ�|/zHN�~�����K�og;�+U�-c`�8���<n'Z�!
e�E$��P*�nu�T|�􋀸�R�8k�k<�4��xsi%�-����5z|�?#}l�
v,�����
;��	⑇���^�w��^:X�$#+��d���>��5�l�N��x�G�j_|�V��Ս�fF,�Ô'��Z����+͇��ŉI�(��A�K�l�&�v�uLsA.��ྮ�/|�����da#_��lِ�1�"��2��2��(8�6䆦E�n���#����k�z_'B�b̳x���܅ϱ��`1W"��P��ٌ�F��M{ZaM��� ؟�4ëw�m��-(��;,I��T)V`�n��
P��;�z��� �mиDϾ傴LV�0K��4�+-���#��V��Po����Z/e�f<��jB+?j�J� а�H=4U�;��e��6%u�-�x�R���2��6�0�=#e�ꯎ����p�e'I2{�S�)����_���D�`�.p������"Ie*h�q��I,�R�Q��7`6������O�rY��rw��;�.�җ)��~�#��\�3�:��S�K�on�#Qw�3'!b[እ��X��y��&����e��3��˝�t@H��70�.ad�<�e+G�!n�l�b|�Qf���?�?Z�)p���Hfjg{��Dw�I�+ �q5�A���K�o'���<b��z�XS��}}F��MV*����Ց�Y�g˴�ߋ�̘�-�x �_�;����ND�7ْ��e�%y���)�]5�{�����tN� �y�+�f\N/�����ۦL0�2T:�ru"	�p�
�=GE��ݷ�J�Pแ.�M}6DF/�')�<Q�I�ؼ��,./��^+zJ�OU�%^x=���Z��Sp��'xEq-�ŷ2����:�D�`�,�:���1yܻ��S�MTC�ؠv���l	ugFv�sl�Ne;��<��i �'i�8�T�޽TC��D�㺭�ִ����'��}�7ߨJ�{���N�!�Ȭq�� ��B�*�_}���^T:�e�Gb���	!VQ�I٬��8��7��W����x&�O����!�p�8�-��M���\0j=����#KD��3�
��Lke�D>;Q�[����c�S��|.����x����S�Oz��&�@@Ͽ���Ho!��g�mBKm�v��v ʮ�����vi��J���L����O��?�V �*X�)ͪl~ڱ2s�_��6R�(ld�d�1Mt�CO���� �����b���}�\��r�1m{鱝q��lG >g+o�fr9D
6S3\Jw(d��y:�2v*� J<*q�)���Yd�O;�iJ����c���w{jW����������5	��slr��	"�S?;.��.����+��?�8��2O�N�=��q�{��#ٗ��@�����z�v�E��7y v8���Q��6R�0�֚�SUa�m��-x�뗥�t�U��?q�0oxz�[�M@c���$���V�Ho��b�. l���eC��qn�x�o�����PJR�����i&�I+j4rR	Av�s*�Ƴ ^-��� ��l��\P+`��N!X]%�Y{�!<��8�W�k��zf�f섩�})��$�<z����쪸�&d�/ha#��^�!�,>�G���$�H*)b�ǿ���8|�[����]W@�+��𺬧¢��IW6 65S��vq����`J�7���X?�2B
t�y�X�/K/���S����G�i,:��͂$S0�RK����
C*h'/-<���6��)����S�X]��5_v��������Ճ+�LfG�|�8��0cIܶ���Q�^�
�c��C�f{�a�-!Ϸ��C��98`$��,��틩�5s%�@��j\��l���gk�/*!tc�=�*�x�yXL�[�%㬦c}&����_v�Z���$I�v�a�UaQk	3ׁS��Y�[����0۵kx���e �`.*Z��=�qڍ�B�L,�b��!\L0풐�E���۳J��%)5�)�G�^�Ixt���A�%�X�3���3�1�S,ƶYf�ZQ��dE���������;Ѯ�������eR�hIfl Fd���ٴ��|r�����Go�06m0�SL{��.�y}!��F](�m�T)�������f����bv\1(��X�E|�Hl����k�K��mv���]���Ե&�[���*Ì��vPc��J�p���w��@���?t�� �������{�c�|\|ᏦȫI���v��顿g���^�<�f\9|fUk|��Sؖ��
�^"B"A�@�wr�]��{i��2������!���/D�ph�˫"�$=Ã��IT]�ͼK��|���L��UT�vN6ᴜo�VHn	�bTR��%Զ0�@���''M@P2�7' [׺Nǃ��[��3g����4���%�B�n>�YZ��o1'0.�: E`iڨ}�&O[U}�ݲn<l�2��9��~BY�L$���P@LE�m����*tS����G;������3-��Gpqgzz�z���q`>�QNjK>:��Tx�d�b�	zro�gh�
pp>̯q�����J��':��\�M7Kp����7�1�=��fPc�����ϐW%΃�NS��w���q>�I�|^hr�DxJ�.�$��G|F�o�l�/�D͢S�$���o^ԝ�i�V6���ƞ*�kTѤyL��K<R�"b��N9 �
5@A��|u�(�����$4��9q9���I�K���b�V/a��yJ�p���T�C��^��O�f�*��<�K���ɲȌ�A"���~����Yi~q9�m˃��K�7�ϱ��C*�B�K3�T.x]���Q����PI��0�Rt)�l2o����E��"/��|�E��
7ߴ�:��3Ą����<�M_Ѹ\���	���e��p���l�92a���[mɑ�����c�O�3O�����$o�,t����d��Q�Û1�S�?O�I�����Y�jI�jn��n�G6���ڛ|��;�+`nG	` ��o�������UIϹ�ڣ:�t/��ځ�}�g\��.�W,�q�S@�4�#RΚ�u�>�����I��˷����7��
�k�]�&�-4��dI~��~���g܀��"c�pA���rt�pn�udM�E_rz9),�6!��!q�X����@k�Џ�:�P`��,Q#��B���qI������\� #�F��Y�0��aj�"R櫖�7��Q�`�� |ĠQ9d&��/M����n�I\S��3/F↖�ҥ�융\�"��/i]v ;�P{�?<E�#r��"<9Ůu�����!�G>L8b��Nt�vS��w����f� {��+��+���#���R&&�Y��d`r�륮36����@;��W�JˮI 䈱(U���'˛��k��S0�:���������U�s ��ܛ��<�v��f�/�ۖhfV�sԯ�;i��J�#Y9����������g��I�`G�����Z�;��������1�f�R̘�F9ǖVS>�9��.�&��f�Bz�
7�ܢNl3��[\�ǧ��Z�{��ogD�6�\���'b�0�+���s�-�?ڀ�|fA�F�$بZ�cF�?��!�6bn��l��ۿ5���:tx ���a��k����ɱ��ۆ�'$P,)&�"�(M?*Gn���A���ĵ��iFKI}�/�z'hO�d��k~Z`-��a��x��i��%*��*_�pO�&�5&�2̈L*cJ8�:��u���NU�Ma�DM?Fz�L�9=w���CֱK�u^�@FI
9�F��M>C^�υ�ȅH6��Vu�:�̶�#mbVq��^��~`m�7^���ь�k1��e�%Ёkg�ɺߗ8����}X��!*��:�/]E�o��RM��Þ$�=�D`���A�ҨKa����3r��_�[`���i-�V���Ц'��?��scF���s{��I���Y��g,�>�b|��v���0���t�!�S�3���#�G oh+��~+]��8�NYd1��ؖv���= 
��U�iSa����)6�;�s�V�^���6+��߷D�X�I���O��Q8-���l��0������s6�2�j�/{\�RN�(�ٰ���إ��gA�nM(�;?_�@�5��7��6� :k-���&���Je�x7D�VC�@�h>=Ry�Ѿ���-e�%��9b8�N�>'��0==z��X
�l�GA4�Fi��i�+���h)���5>���s��w�������_LN�uO�{�&b��mW
�x}[sin���`,݋�]r&Ÿ�ԑ��QKi!���̂d�E���͋K�����ܺp��1[�5����ց2�e�⏍�԰�[^Ȱ��[�(y�1�I���%�Pҕ��
��W[��W1<)Κ;`�_'�1��h�����G�`c#��	���Z��\��9�2>�R�3�S������}�2����]�6BѴ�&��@[����[���U�VP��a�.$�́��n1��
{|jҋ�#T�7("5*u����B�{�(��6-����]���4j�t@n5��jxh��Mw�2Z�,(��x�=���fؐQm��"�*��t�����>FG}R�����0J2�������'A�q'3���E����\��%�K��1v��9��.��_U~}��t�P�}�D��d��� ���D��˨�@���(��1d�.W�H��2�)������k~GZ�>�B�N;]�I��t<0�����7�y�\�ŉwJP�D�:��4ө�[Aq]��&/�.�$O��)m�6D����"��%/$��W�d���-�!H�X��"�u��0���=���|����1�[�]V�׽�"#p�;�� ��T̄���	[���r�2x�� �2�+.]�]���X��x�V�_������3�'/`hV��|v�ut筌����ԣ\��;�x�ൿ�4�;M�`ަ���HY�(|�+��,@Ӭ�T�X�lS�(b��4۷�[$��6]���ĳ�&i���a(��v���c��XX��:�Ѓ�
�Vwd8�B�'�딷�#���E�b_��3a�#�
f���_Ͽ���GK���R����e��^#H� +��&�:�Ѳ���]<�N��93�5<|&���#�b���ИE�֫d����5RsH��%q1��36������J�,���t����,��m��i�"����ˀ_��==��.d���m�������1��EbR���X�f�AH��ly��6���U�{�*d�d���2EN�q��VP#MgU������)?˿�����Yخ��]�W(��ي��Gϸ�R�C�>��!�cZ�H�S�=S���sS(�|=}�F~�����(��B3Z2�&ݣ;0'�Z��=��%iPo��f�I�)p�pP����>�uǕ�ߦ��-�V�d���UR�R>� h�H�Q̈́U:�h&T1�>���>�O�/$%�u���ժ���� y����58��/O��~-�1�G�d&�-�ߍ�C���;c�y~���)7�c+�N zbNT'��ߗ/���=?��R/�fX+�`��F���<L���SŰ���$�֛�@.�M������Z���lOѪ�y^�m����"+��d���Xo�7hY.��/ӭk.P�!��ky��Ҟ@m��ؾBk�u���x<Z��3M��]OeVگ$��%'�S�l���
m:H$� \#��ӵ��gbIx���S:��������v!푮��Xi�~���*��Hn�5Ӡ���x��&�<E-�<����E���Y�_9�x�E�P�E$EcQ9�G���E=K�Wmi����E����:��v���~{5B�y鼨B�t�����̋ ���N Va�fl	��=ڂ��Se-A�	-�y{F[I�`�t �7=扮�	��D���R�H	�Wz�S�]9�,�r�c��*95s9:$��]��� �����tg�݊�s��N]R���M���<l&�U<P�4���*D6 ��� 었%�2Zm]���%���W���&�@�͒�k�ض�$-$��<�����_��ĔA-��:���薹�k�j(U��ʢ��P5�qo�� 7gK|;�R�L�8R(|z�g�h�櫯,7�Yh�E$cm��S�� u#�
#��1^����P�<h��@[�H���i�#�V�;	�3��;��a�=������j�;� �}����s�*��#���GQocW&(�[�/�b��[���� nN#q��o�N���k�1���p�G}��X���)�!��h�%�^�}�a=]��|��SMQ��5י��>��~��[x���>��^6����v#v�����6�~��o���<���煹�/\]W��}t'е�	����D�$��aZ!m�{$u�,*{hXW�/��]�HH4vm��K�Q�h��]�#�b~�cE��GC�}d���������]��+#�3�ۇ"��k��2�ƘQ��P�b-F���f������cY�tP�;z�C��ꯆ��{F2y(�иڡ�MbO���`\'�c�{��>y������-�jFm�;dS�j�-�9*��)t⍃�b�㤹��"sL!TlM�Q�_�;gуJĄ�7�2��J�+�1�7hd���:뽊��[:k��Ht3 �GcC�gv��
�"i�1���S�,m��2�潢�Z賭~hFlbE8��>e�X2e�O?�!iH#'�.XZX�w�uN,LmK�WKJp�f퐁�؞Z���/!�F����-�1�ۈ\����&t����E�or�~\R7��0u�d������2	m���7c��s��B#4�Vrqn9K�[��p�27h�90~��Wo3Ӭ}fb�?[W�r��E�;��F�7_����d�#idD����f,,�CxȞ��Y��<c�����Л�B�٘7������
�W齬wݺ?Y��i��]5���d�N�^�M2��a�h9�����R���1W���ΣWF���b:��M���3�=�W��J*��\ju���e����nn�Z2��
���(Ϭx��p(M`n�LѶ	̟V�#����q�1wE��?4K�z�$7,�����ҫ�����Jq<�b"rx�[;���0�8d�V&�������-P�	�H*>�ͩ�U/΀Y?\�T��v{y]�
1N���Kc^] �ź���M)p/����;��/i���U��]{�-� �w_�`��Q�rc�'N�Jp��a�q{A�e���&�n'u«,��W�ί�(�B���x:˝�/2{�b=lL��IC���W1��!o�Qk�<����# ���#�:��c�q��ئ�E;�:%л�fӯ���c�VG�B�����frBH�������������*8����S��i��;Ms<��r1��ZEzwQ)9m\s'ן𒞧L��>����O�[��TH�$�܎���h�}#lH���P�SO��c<�~��r��͂�8X=���q�L%8/�A�D{��t��~��-�;Ȍ�3�t��Z�@׻�Z~ɪ	.CG^8=�;��ڀ�6w��}m���Dl�	V�X�c$;����F/���mv$��8�Y
�����pe����A35]�]�!,/���I?b�&�ú��1�z���)��&�Aڑ��L�mj3��^c�%��ivA@�6 rC������q�,�J �.�ZMlQ��'}F�ҷ�)�L"�F9D�����e�9�=r�-�V��	��r8�\S�� �����Y�*D��RwsF��L�DY㖎$��
��v�l�k�{0�Z�E.6k7��a&��Ry.w��,Xzg�7$'q�(��z)�b�#�oǅC	H֊bW�qH��.};y��+�n����5ځU)O�_��[�5���L��LM׏�GhD;k���*�*��?L��2R�.��o��'��Z0��;���Q�Z��� W�_�F�)�7��G���s]n|�4܃��6xrBD{|�E}�RF�R):m�����S�w��VqVm�)���}���Wͷ�@kT����ؚrw�h���+{���մ����%l�vaI��~��L<k}l�5������ִx�a�"�]����v#^4�g=�Q`7vc�)2YUh����-�e�C���wH��Θ�-�F�"_U-*�V�5[AO,���Z��b���p�A���Iq�b�h(�mT
ļ��^9���K��Q��5�W�x���>��?C*�s�
��:�m2uI�$�����_��;f�鷄�}x�=����Tw�f^K[f���J��k�k����~.�ch�ra�04��^�W�RS�mY�0�3a�3��#�z�������r�']�������N��1��ތ�{���țkJ魼������Κ�I�/�U�B���Qez.��
A	�kCBwG�8�C׳W �
��A�6���� ��E"��|Y&q,���Ѣ� 0�Ζ�p
&�f��Vn��%Y�Nrb!��A�bi���
��0��CO�P��o�w.�	��fc����	[�~(U��1T���ͫ\����H�����&c�HuT��l�;qjbr�7A����j�Ub��ce:ݮ"�H/���{�^�3oC%��x�CPJ����i�[b`�"a�gSI�a�������x�]L%7�6���`����Fj�j�GH_Zɞ�&�苿Grm�Gz���V�b`6�U]X��1Nýn
�F|�TZ﨨xw�����j�C~]ֲ�E� p<��v���֚�+�d4��2A���;�<c��)P�bB=d�ɺҥ�y�.�y�B@��	u�|Q��$m��8c��;��3#N ����#F��[�H5_�,(!{Y2�`v�W��y��:�?0t���Q�Z�7�|�� ^� O�0�`}R�S$"^�EA�U���̠�c�� ?L�8�c<k���*�Z	��sx����5�+^K t�2���ݽ��ί�3��~���^'g
�P*̭�F�]���)
�ѕx�YB	�^<Q|PJ��W�ڗ51d�����CZ�4y��n�F��9,y��}���K��A���h"�'�B�JpK�"���*��nH3É��r0�~�I��Q*��O>����OW$��-�nH�Ȣ�� .	/&7#1���;�4�O�4���⛫c�@9���$s5�Y�(��M�E���5�K�?b�Q>{jik[Y��ڹ�X���\l@2���=�W��m}��4�?���e�8�)�\���J�+)ǲ�~EYa9�4��Ҕ��6h� ��#Yq���
;O|(��u��=���{���ޠrX�FD�r�: �MF���^u�~��!��\�R��zTՐ�[�yt��� 'k��U���I��c��g�!��A
U>uu�ި���ف�<r��yj�οh�xn]��O����B,n8iv��U����z�*��
������
Ӈ-���T^����N*<���7� %�[i�V`U��Ѫ��E�M�ã�"A�����]���n�
�'�[�\��_Pe
@ط �EU�ɀ����}�v1*'$�+����K���#�\��Q���}8n��H[�J]�Q��YY�����eJn�ʰ��A� �1���>�gf�d�AG�B3�A�F�(�VU��H��K�Ȓ\/�N�ʭC�7hq?���/�02�l�*xIZ����b����	Z&�+1�>��`�k"�Ԏ�g���S2�������U>����243Ug���LƖ�*���G'�rV��q.�@-_ct1�>��*����pG�yY�3�%���f;���`�$��#P�4�m�cԦ�M#��d��{�<_Y�jZN"|=
��]
$̳m��8(���7$�s�@o�Nj������R�Ұ�e�Nk��'4S6-x.�ݥ�c�;9��k�Tl<@zTV�����;���Qs$󶑥�{*Nߎ�].�G�g��x3 h�Z�@�������]�{Aύ�v'���I�)0tY����.��Y�#D���3�o�r`��\G=ې��lm(���������; 3�����em\��y2v��Hb���@�%}�N+Se�%`6ٽZ�6y5,�(��C�����g�������7_�_�ws#%ٺM�8�vxU(�6	�)̓��QD ��e� \iDiu���X�O	fWC~���ʼ\1�<Yv-`��5��n�z�ϙ7�?EOVm;�VYe���0���ᮧ����FJ�_��h7���~�Y�N�(w�[P	��# [o����ǖ$���(:�)�2�9����{(�ߋ˰h�A_�}qJ���P��`t{�z�@�L)���7�wi^�:p�4>1��0[ ���d�FC.1|��2tƃU�\á)y��~-Ӿ��$�<� HJt� Il��'ݲ�)q��f|��;��~"ɜvuL��f���!%ۭ��;��E�S�b�t��]nF�1��D�Ar/^|q�rA���T+�
Z={����f;� �C|�f�P\��(̦, �bn6Y �[�����}�O��c���q�+!v��[�	О�!,�*�{�%��#q���m�TB,wg���F��-r]9�]���E͸+>T���W#C�)��z��$~LF1{����Y�Ex�yq�i��9�1����\V��������������<8��l6�m�2��P(� ��*�s8w��2V:D`2�:�m#����z9;�ҹ���*B\���7�8E�h��\�F��]V0#	,��cHz��Kj8��D���L��F&2�m!��%��H��n4˅�j��`�x��*�%}1M&S�97����N�����%G���0{�}�#3򣖀xu�3�6x�����(���s�2��*�#�;������b\�W�����;@�x<�e+��C�8�]e骑iX}�r�-�Ր��t	��g���9����A�;W��ۮ���&��ؾ��
<�f�6/�+*��T12&���>Q���m�2�ɚ�[�����u�ڀ�H�q�$��ۛ)���YS�Z�d��}�c7�$��̉.�>�&_��ԡsW&�c5)��|������4�=˱�t�>�i�4�
TT�~F���r�hX���!�x��=� mjf�O�����~|~��S�K�&�H���?�n��[DY�s�5�8��������KyNwFg�[������j@��t�j$L V��;e�Pd���5��C�
�L�\�y���d(�[KN{h�Y#)��/��%�
t�:4|ñ�:l{h���z�Gc�\F�:l.B���/����x�~���>7t���?�]qS�cPwE��v/�T�.���° �`_�^���9\D\���E�� ��g���fp�����:mGk�KY3�����AW�A����,�F�����
���t�1 ����9�/°��j܃D[v�=C��[�
��Vj�d��ٳ��ou���	�q�>f������D��4���tN:$�1A,ӱ���t/Q�Bnf��)���:*KX�X��Av���P=�(럦�,lȭm�s����(��V�(����e��WtA: z#*��;�ި�/8d�q�QF\0��[Oh*��b�������x����P��1���6p�~_;変�n\'�c�2���{̿*TP!^�m�-x"]�W��e@���/�'e����9OǙ�j0G�q>k>T�u���yAA���7lo�=u~��TVÜf�\��Qp���6�A1;��ts{U�\�1�<�����0��xN nv�N�9���$"�I�:�zDɟ���~&X}�Y��n_Hk�(���i�':�V��z�4y����p�U	M.tNV�u��,�1�p�;�U��s�y�&ξ�̲M� )ىw)����d��y�*�!�0�;��޿]#�l⬕vŖ:{��,u,A@�l�v��mf �>�Φx}L�zW�B�L���;нg%h�m�蹗n�y������͸m����P�<�Lhcf�������gE�򫗹ɰ�WR���8��L=��f�O�BTh�BW����ɔ���
�Ow<�"#
�S	�h�7}�VIࢠsm��}�4)+N���D�K�%@��R[���sD��\�/=2 @�L��3S�jZ�������o�o���4 �vi�@�x �w�0R��}-�]�� )�Qu;@z�� `����vg�N!|U���-����E��?J3v�X�5��Ñ����٨�)iU��(bb{&���*X~L,U8=?��[�X>�J�<#�� u�jt��̙�#h-"q��=ś�����T!d�9H��B����K��P�{�5:g�R����5(p�4���Ѥ�}<8��i���S,���}v�_�?ŭ��ׇ=X�C{>�nw���0���ǁ�ËO�y�J���D(f�\\�!9�#�j�����;�+�GD�ݨ�G�5ns�n<X1NA���c�kx<J��B��"���TC��wx�V�rnl�-��5��:*�	����cL�g=-G�;%fc�y(�z���-lW @+�o<E�PՊ-=���	e��%r���cSvɏ:��%lIp�o©�L�U&�z��pW�ȧ����R�יZǥ��#P�! I��R�Fz�;�i�<�n�!��f?Kz�עh���1!$����|a����S�z���~w~~}�@'B>R�܃q8U߈ȟ!1*e���x����s�@QYOd? ���c؞.hQ�C "�,:�Oe��U �f>�M�Zi�/��ki�	��!z�0��Gi" p̊I�7�BS�a�=ոY�������3@*/���&S�T�ǉ���O�ۖ�,ᣃ�o�Q솫��{T���Q��-�2�9��@F�Ie�|6��� 	�K+],��i��Yhm�`�8�\L��2�RX���xD��J��g�{Q ���!�pVu�G&�[��X��{T-���^8\5!!��|b���P�e^��/���;2��q��Gtmמ�5�(G(8�k��W�P� ���x�O�U4��s9�ұڃ�7�H����b�� i$��J���{7�6�O���;tW�����J�x�4"겧�%�{�X�����x�u�������>���bg���pKЛ�UHL�VXd3��ۈ��D�P@De2�2���Z�d!��	Ե��lb��y$����:�h�c�T���G��%~Z3��������,��7����p82�7r!���aG����j�<��ٔ���0u������<��� �����NJ��6#�>��F��S���o��P�K��Ӳ<�Pb���Qƿp<��k�xB�c s�q�����
ēSҰ�gbSF�B��ƒ�L2,��:&�Ѳ

���D!�t������۳q=X�D�^I�����"(�6`m������R�➠y4O���#�7ՖeRf),XX�M���yl'b�\��j��\��=���v�I"HO���w��-��O���ArJ�ߴ.��On�Z��=�s��[h�]<C�g�o,�S7�}~�g=Q�s���@ȇ� �­���k�H/sd��)k����j��&d�N���C�d��sj {��Cv$%J�͛ӈRO��q�Y��<D˞��9}�e�˒4ög{y�b|�#��o��D"&�"�E����p���9L{J�;�)h��U�L/s%�͏�EJ,�H�����ka.��!��x���"x���-��X�<U9�{80�&��M$�2?ѥ@��a0!��F=�^]���G�N��lD2��4a;�8�q�Tw)�>��B���"j��~^��`��r��Hч�Of���ŗ�����_�������ښ�7x��]߭T	��ɘ��E+0�9X@T�l��+ڊ���A�z9).<82=��!<��K�z�j��6�(��
�:U�Hb!�ed;�&4�����������p�G��Ŀ��d�|��7����<�˛N�~��3�@�1�{ԫ��0yA�����v��hPf��l�����"�2i���j��A[s��ډ$��z�")\���|\@��ｦF�H���W��6�1m�{Pz��TJ��$�K����!�,� ?�JD�����$��ћ7�����XK�����tT��;h�0v&�O�f+�\�k�j ($��B和�D��r('"�׻]{r���z�|��N�sC��UR��DLhC5�QFY��^���f]�{\7�f�r���]$��A$�������#D�{�MH�x��|�2q�6zyB6��KS�2��d��V}���Y���A�k�ۆ*���m*�!i�m:��(ܱ��0�6yI[��k[��L�gfd{��mE�&�t�&4��=rB�=\NM�f��3�o(#����m���Gv(���ߊ�w6ً�&90m��j�}�⠂�ؗ���L��#R���&I̦�k�v(��1bA$㙟pE�3��+�W����U��u��Q�l�'b��ý|���|�):oJ��['���q���X����섩"�{��k+��͖H�����Ώ��䵬�Pdf�^mTr��w`�T��y���(ۭ���j	K�z�"�_jB�w�Z�7���9�l���Ѷо,�?z�"����d�Tc��fQ8��9kTo�'2]���@��`U,��SEs-���d9�s�i�i�d�Sϊ>�ć�c�0(�&/ZK�꽶;�딏I���)R�a�A�h���Jm�Ͱ��mm���LY�N7�9����f�&*�Zu%^��{��k=�[G*l�=U�Hn�`W=Oćý��&�!�=��UZ�H�iڀ@�n��4��?��ճ�@��*�}�m{n�I���H�8/�ּ���a]ji,�-�(us�i��zoH�[<o2�8�p3ۭN_�����5^�k�C��X��f��e�ϓS��"Y'�����j�p�ֆ�n�����K�Q��*�K �C��%1�M�)�
?�N5���� !�dT]�LA9���ԨF3՞�*�5a�v�>$��!>�p��A��,M���^Ö�	́�~E��?�Զ��դ��"���Q��9�=��ka��NB~y��kr%x#�u��7�r�A0�g6�|��\�kl<�,�ܿ?v�}=�U��]~�����HωwwdĿ�76�Z�
f��f�T'��o�'�SK~�z��99��MŅ��ur|�K4Ux�p��》<BBn"���4�+�Z��dt��
�7�5����0�[�g�C�ItI���KԪ�Bq�E:QX��V�%�v[��i��ٵGq'DuP�	ǩЇ������z�;!���X�G�´�e��dHҧQJ�R��0\ǘ�\�L����QW�{�r���;�l˩2�wb�p^��u���O'��8�V�
j8�4o�����W�mY-�U�t5�)M���������a2�����c�Ȅ�5��1����=�sJ��0(�AȪHxH�=uj��B�3���ׯA�K�^��i�T%�5��4�f�,�*/:!Q���"8]��c�E���w�Q�)g��R�F�ZbXY
�G����1������騐_�O����R{ �k8Q��C#�v�H�����:�] �"�� u/�
I�U�/�X��� s~�v�fM�v�"�:`�[!��y'C������13d��@!���`����K�Pl�L�aQ�����|{� ���t�(]��'B'���"l� ���:��{�ت���4̸�V�)�ў
@Ű�/8'q1T�g*f����qQԼ���ed�+���0c�qf�g�fpSl`uܕV�[���m�����~n�n,y�����He���л�|��,�2��/��r��t��&��ې!�l"(Q*WiQ����8lŤ��rDn�<��}\Ƙ
���}��H�V����/�GV�N^LI�g�ݥ�
�\tz�Y����G9���Pf�s�[���{Ϧq�Mg5�`��5Xj�&p�������;�z
H�R�6�x*��>Wlv��#����D�o���<=\g�� �!�����|���7����j༟.���4oM�?�7H8�
��A�|���zZ�Ad��Qj�oH1g��i��J$������c����)���7��ҳ�vq~0`�L�‒Ѣv��^c�߿O�W�]�����;T#�z�)*��ƙ�z6e)�By!s��i*y�%,)�����T�=��ܽ�=ɕ�����)8�_!���aA.��J������:�#7H��Aս��C�归uNlC�_����J�`��Z?1w�~�ͧPw�����N�1\�]��������TW��N�w��d�v�f���&(��.��Π�鄺���(����PxݯN%	�y��Z�D����œn�c��ζ�W{v"�FW�$_�M�5��h�������T@�HV֍6�F��dn^V[�c�*Ÿ���c/6d��N���'�!�K�V��L6�HX�(v����Ĥ�,�lJ����=e�x��8�B)}�1o�$V�*��2]U�*
�/^ܖ{��B�^H8r�,1o�C�β�oA{�Έ*�ֆ��2�D���=@[[��|| �is��t�˲alhV��&[�+?�,���C�IRl�Ӗ��/�-�=|�_}�뽨��u��p��KZ�+5[��5�Uą�̏C0
��]�y�*t2@�'�<B���K�VD����{|�o�Ըm
]�����I3)to�/X.�q�G k��ɀ�!P���%�:�j��x@*UZ��F]r�bw'6��FBrBE/{JQ���=���ﻙ=ux��rSƍ�&����ĺ������L3�P�B'�#�Mwt��N���м���?Zߓ�ˠc�P��y��>y&cN�!j���+���lbu���]������lZx� �����3Yg���ܣ��D�ٗ�	I���ua0gs��O����R<0���trL�jL4�{�\��%p�Y5>��������7����b�z�P�e����t;C�0��Q>�]3�)d��=���+�ҁ��9#�_�g!p�N��CJv_P.�qB��P����'���,M�p��WS�fٺa.F�ȗDm���]�y�S�yNˀ��f�{�Ha�<�H��`��}�L3S��:���4&���GA�Q�ݼ��Ӡ�
��V�E^VM�\H��N�% OF4�Y���\�p	׿r�X��Dx ���e��<�c���$+5W�BI����c�����ZqD�2��JƈAEyr�;���np��{T�{�v�}�LY���/�Њg���sO�0�f�����?��#J�.��gw�\�T�nH��v����ZƠ���{��
H�1�T�� ��tN;дn��y�X��d�X/�Gܟ� ���ퟟ�)e��Au�����^a\���3��o�o����*��q��$��C���[�N�jZ�� �fb�Ժ C�8h�n��(�n�HOO@�#3��8n�ه���4=~D�V�hS��������S�%Eo)�[�X}l�=B�/�pJΈ;�]~	:�	��u���v�C�99<����	��,���n&h�����
%��ބ�XI^T7t�/��Ɍ|�v����&޺�����0<O��|$�O0>T��O^@�F�t ?
���/=iY����j�0��O�]Z:m�W<h	�w�]w�������_�&��=.��8m�&81�b�J6��CA3��N�<B��qp��٥n���h�a��v#�����������C�¬�n�T�~F�03fF�p�����/Qkq�QŘƻ̗��H����5F�=-�;�5U�rcZ^&��B\�j���F[�7"���n}�N
&���.s���'��ث
���(I
��z��P�>�=�����u[�TFKq��Qa#+aS���\��26�N�vą���ۮ����a�����#���wʹ� �A5ť�X� ђ5��Z_bf���h�����ۉސ�`V��@��p�	s[�j�/��ȣN��36�k6�D��'<�B��9����[ �낪��tL�Y�S`�˿Z#� ��&���|*�ilm�=��VZ?��텡gf �qK������ܬ��B!���T��Bo��+��.�n��\��ߖ�:�Ƅ���4����c��W��!�%��*F�'f7����W��x��w#�Z���G�b�xeg�/���{��aQ��/+��M�0N�����1�Jk_y]��J�N!�?πS ��m|33,��;�=�_�������N��۷`F�yv�HrO߫#�$�u�2B���Iǽ��e�d>)�q�%�z�~��?T�`�=cI�|.7��=�!�ib����.h���j�gr$��/�*�R�յ�*����-�sݗ����&��b�e�)P���	0�<r����?�	n���{C����$��F ٺ��zO���\���ڪx��7��g����r6D��}�)?���5������b����&���-H�^�wU�f��
� �X]_�|�k��^~�%XU��.������"��Е#��#�u}e@t����=�ߧ�b��K#'�U5#�m�\^��m�)y3��RIb׆{@|cϼ٢Q��i
�1���4�gl����X1����(�:�C���G&����e�_�n����{�{�������2և��� ��/n�&A]d�sGJ�o)(�q\��\�V�L?Ư��"[�lW~�"�h�����k5,�� � m���NѰ�yp
Ȓ�T��*g��!������*
��Ʃ!��:[N��1<�U�r��HX��:�GuR��a�}LJ�H[�L�
�i���i"�����єR9��/��MP�C'rE���}E��C�;^#x 엗�u-���g�q0��,�n�:ۅg��-W_����F�$�?FC���Ƿ�M.��?��� n$������"��}���4�S+OzE~d4i�����yW�p�_+�瀆4�'�P�c#�f�f4NY([��8 wbQH��V6n���=��Rw���Tu,A�J`?��#�2�H}�X�gEq3�e>˒Q4�I>}�rP#lU�x�ֲ�v0njG���������G�+)f����4}v����e�7$�z��S��Q�b��P�`�1�s$5?�/�:ˑn�B�c�#uw'�tv�Y-d�XE��B���6�d����7�C�ǺHc�y�sV�R</Ȑ(sVV��Z]���ҁQ[/��Ek�d0�2��A�F��J҇41}£AA�"��bp˭��S�e�AD*�k����$8�yϛ#��9f�ӗHꮎJ58��p��(�����簦3Z@WN���Jy�G�'TXu�����W]!���\{�Jk�c`9Ş֓���-�{���c5$$�Z?t��S�	��
�)�)�ԭ�3d������4$,�a1�p	n� ��rq�嗾ɽ�Bo�"4/�3��!�k�D�E}Q-�c����`�g ��3mcN��n6�&�9KU����}A����Z���'�����qkO*�vQ[���!� �O��ҊV���b�A���T �C�y�`ì$ǥ|�	D�RO'r�4��M��������x"ZXj[5.�XQh�0�R����8���{g�T��ń_>�d���}1��|���i��Mw((��Ј���#�9D���>Ϡ�%�ɰp�%s�4���^���x�F���PT���#�M�6�s(&�V���#C�~=��k4�NQ�c�g�Z��2塔_c�y��"s�xv�*���'���z9R���8E��J�� ���D%
]6���YL}'�1k����$�Q�A��^?iPW�#�k]s �>�N���뮈8gY�H
g%��Z�߉^L#>bzX�fL�֔����C��x
̟�����( �۔D��++, e�D��V)��DEɡ�ж9`&(�?�6"F�͒�F�쮧���U��u���vBn�l^�^�A��\�p�$�t�9kx�Q7�����6u�EB1�N�c�Sj�%�&!�w:��>q�����vD�6�ƸE����0r��,��I��N�+{���^�CO�r�=ό�m��FzVIr�n1s?�W~�(�Z%E6�t��*��PmLJ	R�,�{=\��S���U���$m���Έ})תa^�'���	�L��h���D�-��(,=�?��ŭ!ԅ0�	x�N�C�L�S�՟TXW�Hx��ו���A4SxF�9������v����$���Dh�+G�q��s�e��+/�X"JEY��Rs���n�2*\%���B"����֪7o�Ȱ��'�ֳ�,��H�`�,���p$.����e`TD�&��s��Im�Rȗ
�Pc��ir�MW�w�Bf"/�Ү���x���r���/3�Q����L�L��3�ͥ����a�8��%'_L�T�$S��[����鈛�1u�ˤ�����6Wf��A��h�D��p�&���+Q���\0D��s��s��!�����P���&���W¿��n3ؚU��� �����e\8�ծ�8i�
���6�8�9�!�\�sXH�G}=ae$OH�o��Ă���c��f?!�
�;�ށ�F�g�ʸ54�6�����#��n��or�Ø�8c��Z�M�.�Tg)�Ը������P�y��}���;<�!D�.�ϵԿ~������c`�=�]�|k�����|�������p�*=��.����D���pR�>NwH/�� L����;B�#|�hC/ܧ�A�����g�CEV����a��4�C=/�s�#�=��������'?8z�n���>*�R�A�k,<�uu�bq�k�S*A�[!X�ן�  u##��%�ȓ+���Np���(���w��cn�<�#�e�t���y�9��|���7e�O���RNz��u�
1�U��D/{��@|V�{��1Bq���;v�K�Z� ^���,(חD�H���~� 5z%p��@�t~s
H81h�e�tФ��*�-�_�j�r��	_we�\cf��M��c����^�tr�c��x�~�'s�O�l��ZK�(L̹"Jn'm�e-MgV��䁒�I*���9����4^��7ee� �<>'^ٿZ8�d������L���=���<47X�K*�������+۟D�N�C���pQ X�����z�
�� ���a-�_�K�AHDG�⼎��q�7�u8;S��W+���U�L*M����n�rl��E���
��t�b��-���>��5���7��O�����FC�؎��D��m���KY��x��c�4����(`��40r1K��ǰS5�����<���֜�Њ+9��I\?�д��MH��Bo@T2$Yh-/� V�4��[��hxv{��y$�ź5G6dN��X= �u]6�~9�����]��rpE��[�%�J���C�z��G����nWe��9�;e�Y���0[�)���c��A{YN���m�����bYO8Eޟ{J�U�U�ɛ_�V	l��?��W���O/=!\,mo/�,ؾ Rd�80�
?����jL���庆��[��7�����M�"��ͫ!�p��BhN���Gc#�	��^�Dg|��9-����뎃�?��Z���Ki��&<�Ɯ���`�J�]���1RM&��UBZ�Y�/\��g�F~� ��69�Z�#m���KU��Eʼ� ^*�T�]8�];�~C�6�U/�ܼ�.Ь�9A�t�6��ڥ.<�Zg��aD��H����@��N�2c�ܣ�����|t������ :���U7I�˼���}=��ZF(%}�7zq��t����uc�l�M�V�l,�j��kD%�<���+{�f�®#�ˍ��O�N���ƶ3p��ΞM�^��x.�� g=��ʙ E��O �J��Aދ���ɚ^d�� (��Ql3cWiҽy�T�U���d��Z��,��lM�& �P�	d�Ohҵ�
W�_�f�kDL�����2��?	I��F������H��r�㰜�K�Im�f~ nI�b:��?���t�/�p<!�5�h��KԞ�Ua��%C������6�̭0e�&g�hs�v}L��w��Oy;Fp#40����Ů�.hҹ�e��u6{0� �`��D�E	�6��{]u���^:���؝АP�#n�:�/	}s�H���
.��F�4��U�BSk�6�!�u�P��n]�D������C�H[z!aW��h��v�T��`Q�u7��5۳ m�I�x���N�G�^�0�&���b�j�a�C�.�W�ω�����)KV�1�}x�;n��*F=�Vuⅼu�:�����}���7�3 ΖG~�j��"�S�*��-�uG�����0%���0�l�\w��J��碽d�4�L�M��K���s��G�〿"gX�~�)7������.s,"�	j������N�k�� f��*22oqY��KڦO�+�����/�z�&&��0`9������aT�pK�z�c���l�t!	P�ɥ�Y4,�}��B��#g�s�H�i�Y��n<� r����0�Z�����jLJ����#����-
!z�s3�Q�V�m��s�o�)1����in�x/������L���y��>���B7"����M��ʥ�_�{uA����P_8pm(&�w]-�3��ѫŪ������R�w�N~��&@~���RFWM�N�qu�1O;m٢3f=HGt���S#}�ξF�^Q�+�X��/�D��]ח;x����0y6E�}�]�����I%���c��E{�\L�F���m����|Ma+Z��
H]X��vQ�B��F�ʜ��@����sP���m��۽h1�ݏ0�&BoV�4��d2��UYO=nV2]�'������W!CF<ld
Px�K9�ؼ���x�b��$��,BY
�ئPNL��&S�މk����B޺^/���B�sf��U5����E9�k:�-g�j�x�S%�T����#ҝq��cm�+�t��@�s��k�jۿ?��A�8�kNJ:�+�U���G����5d��b�L$���5���a��[�_n�#c_����X"\���!��)�z�.�ۜF���~1Fь��֎���R_�u%�0j�����4_�	����o���׉�Y�e�8�ǋ�G��v�;�{��e���Y<)цɇ�x-���~�R���#7�_�����F,߬!�o���#�a��;*h� ��A>{^JO�����Q�!���s?(��5v��ñ�ќP������1!�
��C	jt3 ��ڡ��q|��.�w~�RM'>c��u	�@����+�?3љ4�>4NI�Ryx~�e�(\����{`��pe:f�l�װ�ǭ�t�@�T֥eW(l tHx0��n�4������g��zE�T����y��T��8YS��<�Tx^T ����8Q��%s������5����w#9���:p�ڱ�� ���H����9l���ܮ�輪tvi�P��@P[��Ru�(-�:Q�҃�A��{��8U�;�[�GJڴĔ
�2�%4�x�S�U�3A���2��o�oD<=<���A��.A���J����eb��Խ���/�@��qw$b��;`�qB�M>�?��'i�X��)P�	��%��N9#Э�$��g�@�J��	1 <�!r���X�nC��F��$�x��U9�Ա��ڣ�;�k�wf�m����o��!2����]m����&ʜ�6$�ơr��ҳpv�i��V�]F��!s�D��˟*��g��I�l��)��첏�]P�[-8H�sa�]- ���C�|;�)�7�=���'m��`�ߩP��n�0���A�� ��H��Ͽ�3�nƊs�הo�u�S�Î�ҳ��e��Ϭ�dq�u�t݄0�m58�R��\��$8�m��Ѣ�pO>v�i�%`_1>7�2�?k���8�ޟ���
������n�$��ɨTZ�aM� ��1���1�8i�+���[Jǃ�b����xKGF��Y�������(y���Pї�n����'ԕhy���!*a���nr*G��!�s�o/˟��mp���3�#�5i�y'}*��#��ԗT�� �kFH(l�f�ˍ��td�jM+�2�/AV�?k�S�){�J]��ci�Gg�a�<<�J���,7fRu�O�߻��mj�G�;L9�:�	�sI:�iJ�xFreD�k>y1 ��X�r������|BY�2 E�j����-�E�*
�e,�r�D<pMȖ�	��Q��ݩ��O�%�H�D�Ҭ!p�eMeM��-��d���Z:����l�u�?}=�ŋ�xw�6���?R#����Nߖ�)I��ud\f���,�ʋ4�+Q2(
�mm�����H�Ά��(W�ދ��wO�#b.��l�
���[��X����������fzO�oa��E�R���,�<~wj��h�pC�,ZbR�$P����F�-�=,�YD���ztEE���*�,�'{��g/Z������n���h=z�8*��2����x�|�7)	��|�Y#�;:�]5O�k�?
h<te��6b�F�|��5�C��(��inm	*c
tP|����$ӵȦ�G�i�l���5EB����U���=᐀(�]g/���]m\
ESp�ט?� t?x�?��=6�oĵ�4S�������JԘ�~A=�޲�����Z"Zc}@6
^ ӹ��o$����V�8��6S�V�]�C�-[v<���P�#v�}UN��!�������ʊ�%�x�_�.���Q���_�tW�O��*�O��ѧ�	��g����������b:)�:��J��n�	�Q�-�gP�W��:S~��O��G��w�A��SLأ���ߓ��(�Et��`��*wK���X��1@���g���<;��
"�W�X�\�^�v'Hڐ��z�  E]N��Tm��g��#.H�QU�m��Qĩ�c15%z�b��C�W��ػ�*i�{n3c���<�x�f~�����:-��̕X�2���hF'7=�M��S�bNpp���lCXRl���{edtwP.|X#o�g����+L:����H�� 3pd���Q��!L�� G1�Qk�bM9���,nH�)��Hy;�0�
l��Xl�1"q�OYm=D��Ϥ�;v����$�)E ��m�)I�:#��;b�K���l��)X*%sQ4���ݢ��rg�9�݌<�6,�e`P�c�'�����*ʣ��u�G���«��k[�f��d�1�h�'�K긻|�*�jɱx9j
�3k��#6��"/���[t+�&�}��pw��H�'�����C�l��'�
μc؉�!��P}�SN:�v{瞜h)5�S�������z3�0��(e�����i\���Wu��[&����O�g�����*^g${�v-tOm�*0,e/����r7h�-@:�������xʐN�,Q�����%8QS� 1�C��7��D����W�N�6s�'9�~C$��`����[�m����&�e����NU)q4�֪��&WI�%y9!��Co|R��e�r+���^���{�%&�]R�|���N�1�9'��� ,P\����?�d�?/�ݲlbFi�/e�o��[�ǵ��T��'�k;BO������c��`�m�I���y��$zѻ�m�D�檹_�q��B��'��B���u��E#�����E	�tNF��'�SX3�?�g�<����_m�hXNx4?B���&O�����%��f^�ɱ!է� �+ńx�
;���|}���QQ�R��,�tV��`h�� �R,�d�\Tڮ���X������B�ˮT�	ls&!��FT�k���S�b����G2(��\�����*�N2��0��A�# j{`�Ĳw�%'��k�ϊHeT�䫿s`�%r;S,���մkt5�$Q�?�����Y@�QrK�0��z�1�%�N7D5R�mh�� �%�ڮI��bE��>������%��d����}�~6#�8����N��YX�Q|� \�N�瘨�'@A4p)V M/h/�=�"\�c��j�CO�	.��.f�3�hV�a����g>�z�"�AN���7���Օ	I��G��x�����p�|��Zȷ&ஷ�R�ns���Nl	�R�����d�iF��(rҕ��-�W�F�E���G=_�	M*!-�tw�Cי�$�@ʔ�����*�{]+��U�P�k�'ct�!����@�5_A�)D���-�ݩ3�n�P�V��4��uk�3����v��r��wظ:�Squ�g��`|���;�������A`�P��0�Di�Ƣ����c�a�͙�v>�y�6ħ�N��b%^�:'>�]�����	�5���"�9�+�Ojۼ�T�J��-o9�&��s�S#��o ������b�I�%>o�d׻K�C�rOq��X�/��-eB��s��(�u0a�;�md�K��dS??���+���S���BZr.N����u0,l�����2	Z�k�~0~�R��zw�m���v�=Z��5���|��������{��&�P\&Cb�;�x�m���Y�Q�1��u�0ڗq�"1�/�%��	-eA:ߧ��[-��w������lj�+��
_y����"�v�%ĐQ�J|s�8R0���S����0�G}�M��׿0��-����tr+�x<9:7 �:�c�Lޞ������<esbTLN�Kק��;@@y���������]k\v씷���1q>��k��@�����:-�����T���f;B�H�>��8��:$��&U��	g3�z���J5��u?���M]+�+�p�j\G���5��T�I��+<ͱQ{��9�;�8�s��EpF1x�K�&�~Q�X��׸C�8�,�jCW�ᾩ�EJ��>6�����~�d_z�J�"|� �x�=���]N�-����p�$@@)ª����q�A�o.r��W]�,�_+���o��Q4�����젏�YVs���%rN4n��l�5���.h�����i��P�����ۘm�p�m#f^3�6Pq��aT�Y��ǨQ����� ��&���UUV�����
]��׏�iHoLWk�m4���u_9$��k>��J#_ߘ��1Q)�������xx�ީ���!��*2�|/o�n����#{��W�z#g��[�B��5�	����a~Xu�_U�,7<q�U�sp{���A�L-�4�_���×Lt*i\��	J�t�ZO����p��*;���Oҥm��k���B�s�*r���qV��K�z�-��o�\�`Zi��Nc�nq�c��#f�^y�Y�%qu���
e`~Ƕ�0��rFn�@j����/����M�B���K��^���U8�c��(��"��S�d ڢ�5��!,4@>��/^j�WZk�뻙LKvu�q'S�{~�b�Td_uq��U��ܱ����&Д��>�eI��ۏZ����ڌ�Ӓ���+�&���nlyYj>�W���#}'�Xu�O?2��*01�=���!?�N�Ր�E�@1ͧ���z�,��\щ�µ�����# �.�b���4;}�I�l@�������&��{YM��*f���`���mʏ���0t5��L:��ڨ!���-�d����5�ݲl3c� �j�?���g�Rl������t�K��~=�t��`� @��z���J�+�_|z�XPm��̻��.T������y���e����"��.I��W���p�J��#&Ǫ�銚��9����Ps4�eM�g�q+jC�U�T1�nkd��9��A&8�,m�����Z��Ȩ��m�i\��y͔V�(���y�O��hR�"����iB��H����Iy�MS�'ǖ�a�ȹp.�z����w������6kS�QL�)���#y�3���m��Q�)��e_xa����A� �B����_\��U�=(�C^���Z#G#�g��ap��L@�iܫ���ÇE�Pf˻ì�ǧI�=n�����Ҍtb�9LA�
�queL�}�	)�4P(l�!?�V�.Y	�]�x�A�ꬕ����?�8�HYJX��{����9��fd����8��W��65����٪p�޽�(D��j	R"���ѧ�C��ٯ�)�Oze9�lO�\!�~�~���;��͚�A��Z�3_�6e�.a����;�R���r�!24i'�]��K��xhw�ey�:�#�HR�i��*RӮ�¢�c��ly~{]I)���g!cN��*C��#H���hiBv&��=���F�}���}�R�I�&l>$"��\��� �����r�KQ�5�{�>�@�1���MU[������L�ϼ�� 4Eg�l�����[�Lp"������rH��9�Ҵ����o�W���ICD7���%����ή���Ʌ��4~#a-�u�Su�sb�8ƙ�©���%��K�.L��h����A��'�f�t�A�7M��Nx����lR~���]C9.�ݭ4���v�� ��д�ppp�/R��RV "ŝH�zJ��T~��wY'g�He��Zl��.m�ފy������J#�ը��|�1���4ŽLƎ�p�k�w#}�VL]�o&��W�3H"e�nTm�4Ò�� ���6�xZ}^��Ͼ�?Fk1�	�}��Q$j�oϣ�F�]\b/����=-�^����sh�"a�	�q�ܡ7�S.�mlO)J�����a�nѝq�ޣF���_��������v	�xы2�r����\�E�l�Z �d�6�C���}�ĝ�љ��|���,F���2�'�:�jN�~��[�Ӛ��"��u�;kusj�Xl�� �*���u�lֱ\j�Y���<��{�ێF>��D��6)���������^D閪�Ha["v]B,�e�c�_6�����>[�\��HC�[�4��ů��.�#M8�b}���Y�寰<�A��fJ�ڋVz;eQ���=���!g9X�T`�1�,�Q�tWS,�8��׎�?N?_
;�˔�r�%*'������S���8��5�&�R������I�C��c������M4uʝA�����b��r��iU{�.�S+�Q��M�U1�pz�8����=� �e��� ����a�S�_��?��⸐��6I��S�Q�>,E��4,�rG���Ŕ��+��e�|���Jr��H@6��ǭ���zB:)�jZ��6��ե1�T'��b�v)"�R*^|�'�xV��d�&Ri��3�\�Ecʝ���e�t[�y�&�*�6T��.'x�=a�����cy|u�2Ci��-�K��*�T*��<�B�{����ݬ�n�O��ʯ���2�^��+G�V��n����3|�_��hd
�S����R4�+�Å�t蟔Q!u�[D���3\�� Ś(�p_M7�A�$3���,;?ȏe�&#���f��t���E��þ�G���;$C�zu�\x*1vkzܫ@[Q2�n��j�vQ1��_���gAzd�"���on뇵}��v�KX΂��H%X'�P�c6�w�� �E6/�ir���;��&/b�`l���'[���4�@4�B:�/Z�#3�H�g]�v��S�3�l�5�����#���6qr}��h���):�����w�9~�������r�h��5JzC���l�Lh���
�T�艹�NVŠ��"XW�k)+X��[Z!���%����k�x�oD�5����)���	���\5ܢ-��V�c�Dc+1���@qK�����D|Y�)���|��lx?t���KN����>�[*Q-6f�D��j(w�@�9c\>!l���Ip��+I��i���H�����?�\;�2u����x�dy� �!���)'[w_��J�y��|�ʻ��y����Jo�e8`9�{4ޠ��߭A.}��P�Yj��y�[xR2��\�Mv̀yYh��(�|	��M��!R�,�������\Q�����-Zo^��~����,���J�UR D�2t��7�UفP'͸�
0*4�*p�)�V%&���[��d~�P��+D�&���>r�([D��9�*� ���B�����x_��X�-}S���kj����a�g>� ⫭�yL%s0=X��xΪ|�Vpv|.֬:yI���[�b1��ë#��˦������%dpA�<��d�C
��v�t�ó�r����������N��Xr��"b�eJ�X�u8�ܿ�Vޝ*�6&���i�G�}wl���T�ʄ����#�1��1�P]���9f�ע��2�Z[�}��Z�×�Q��4C�(" �F�uİ���ѨAWa�x"� ��vZF�+{�A>�"�r��$rX����2�u��]�a{��M�T�7���F�ߢa�%?�B#��;�dst�	��,���d��"Ixj��i�r`�r[t��R�n��2�����1�g�sÑ�Ԕ�p�-m��Q�Ħ��>6:�ǫ�Ŀ;�g?U�.�@��%b�U�ro�P�s��7�������]����U͔hY���fұ3�,�`��Qy��'��OB���~�;Z�T��yv������q7k[�L-ZwB	����8<���2��n���]�������I�w���s��w����7|��Po��>cQ�;G�L`�	X+)Y������ /j�.�fb\[���M٥�\.���š��&Y#Qu}�IWq}oc��YIe�5gqJI�FQ�B$�\\�9*f�D����/����m�=��(����$d5m\�#����r�� �'��$n�̧��������IbB?Ih1��1F\���ω!W�/���J�<|*�w%:�N�Tö�������@���L����qHv�CV~�T�״T���>[�t�n�6%�K��&v�va-(�����q+}���.:dz,SE�����j�z��u+8�z�(_\��2b!%S�Ex�l4.۶i펙H�?D i�b���� Cawp��{�7�L?:��d��KY/̸NI����S����-��2?>Vn*=�]I�mF A�@F��L�o������PADG�Xh� kR]k3B��gԋL�U��[k�Q�'a��
C�w�Z��WV���S������B]��m�|$ߠCy��V���ޚӞ��CP͠�ڦ����?ؾ*ˡ̜3�Q:�^&V��Y�yp�G��L���;ڌ��U/F��gY��܅^e�8�l�����F@2\��� �5TWe�"X�ۊ���?�ѵ�j��3CU����6]Z �J�_d��(�S|�}���H):�&_#$[��;y�KQ����������Z���s�p`�^�sfbȼ��A�!���^������<�	w�լ���Z|~)R�^�D������OJ��l��X�'�M�yP��1<�
��A���;�QOXܶ5�~q�Y-]����r�4�V|�:�����$W�T����Bs貫(�
�FWT\�	�?��W�ю�^����kq�07s��|�k�k{p	��.>�ȓ��'��Tܸ�uxm�:�1(
���|<�����D5�*;�q.��.�(\��d��R�|ݟR�<qq>��x�-��"v��Z�[�E[E��U �R�J�/��R��_ß��;)��f(1;�o�I���!��SRb���9I,�~a��i3��������Z�Ojgݘ^�dnb9�:�jЂ���
MB�}k{}�/ы���������QĽ�c�W
�y�b��	�j�����/Ԏ{�EK�Q�%��2��D۔�������-Gc*��,��s�3Mk�	��=�q�"� �8��X�#C;�,�U�#��wx�b+��b�,�d}�����ʑ��n6�|E�˅�)�_���<�p�OѾ�[����h�ĆT��_�G���W*��MĶ5q)
�A?OjN�L�{	X���L���N��&a�e>��cDHŴ��Kx���X��{�Y��Y��?��eo-�]Gk�8M���ׇ>� �R���/Ձ���ճ�w���<�SJ?x0#"�F�Ʒ3�+C���u��n��� ����׊s���
�5�8� ��������="��e�&B$R'!�<���T��S�GB�H���E����H����8�=<(�-��f�\��g� ����q|�~����_�V�������t"A�;��4���[t>o��v���s�ǈ�(π>M*������7S����.�o�l�.ǖ͇2���*����j�!.�Ō�w��涺nk�O��Ԙ�Xڿ.Gx�Y��h��pRC�?9�;'H�-�,ע�w&j����-Q1����	>X2�>W"/s�]�B���M�٣Y�{}?���*��<I�Ш L��g���]a�aO3� |����x&�(A�$|��<Bl>
Ӗ5	i�Ҝ�z������W��@<W9��E \��rÇ-��D���>��SUV�[�龇xl��=��@V=�Q|c�vۛ��u����&�.V������+!*d��CGlLlO�{o� ym���m��rN�A:��x��H��^�)f7[	�J|�.a �>z�:���r����_^䴾��<m2�)2�C�0Hۅ����8�vXK��{^��F��[�! �S�k�6�j`�����U.�
T;���َ��wٱE�H{��E��G��=8�S<Ѓd�-��5�p��^+�x�S�wo`�UM��ǋ��rԑR�Z~��R�x�e�@ֈ�Y@���u�cw,���z�so8DJCrkY�e����pļP�*r� ���WT@��oˁzÍ�~�h��D���k��7�<Er��I�:� ��ĝ��f�|���&P"b�Oa��a�{����� U��� ����4a����2^>4�7;ݧ_��}W�nZEQee[QuF0[1���geCR����%Z�r�K��>�6�㑊,���j��cL���� ��U�X6� L��杀�nYq��O)��Қ�N�t�Ԑ�iB���!���.���>>���*�e޼�5[�����o�-F6f"4�sT�����n\Y��{��[��ii��`��hƝ-�oQ�YR�b3�|����PA�AO�x�+�7m^�^��+�z�4�Yi�բ��F����H�����Ne�y6ԋ6˚�_'�;S���6��;1
K/��5n�
k,�(M�������tKBqۦ���>�ڲiFT-��BcՐ�f[���Hs�uGyΈ�6�X}J��<Mq�RS7k|�4u�h�� `�����Ŗ�����k��4D��P��/q�F�`�m�� BD�Ah"B��ZXs����M5GH���2�|.�D�˅y�F�����Nz��ԱR^�\�Ux�?�:V����C�5�wr�>ǿ�S��̘=N�}�1�L	w�9�-%�Z4�(9�Z��N�N�!����������.W�Gv;G���U��t��ɽؼP�64��(*4s��p�ךs)���Dc�~B��j�A��Q�>|E��	bf�n��H
������{�)Z�<}X`j�i���In�1���N �D�~�89�_l�g8*�'�  ��A?�3���_�D3Uis��1\0������Ν�����ßV�������1��'�Fg��Ev���A'7���H:�(�o�
����-h���Wk��c��
P��}��i�,��\\S�hu"�B~����w���J��~�:Ȏ��Ih�� ����.�ۥd^N��!��+����63��JǬ�0nxL��q.Xt�~����,M���GY�ݨ���xT�-�<����'�ش��C\O*iEe�a��{K�Wx����Я4�Mէ��Q-&�1|�	j��$ډ��M�SF!AL5Z���Ahb�H�����(zg��I�I�gG�G�ƀ�S�\�}�*eh���â��,��j�C��oɌ�q ��[7�����W�n�+����N~��i�ƦӘ`j	=��*b�ϱB�>��Z��p�X.�"
J%�[�}�\��%E�ߒ9~��<l�A1�!�����I��ԅmRKݩL,�9�:��A�>�e��~���8����Y���.l�[V�MB��P��k�W�K����cn:�B��B�$�YU��urQc�	�%/p/}���h����~&C������l��e���c�]�A�~�1��D��Jb8�[6�M8���.����:�Qh80��X�f(��̖>-�B��fM��hy��o3����#j.6�O�M/B���
u���6��
�!-^��8z|���\k� �~V~ש�"����7I�t3�)�k��hJ�_�6c�5_�֨����j6׷�H��`�r[s0kd-q�ȉ�����/�Z��H
P�0�q���P/�1⑭���]X�� ��-�xWGL��昑A�^�^߻�|
Z�������Tic%r�I_���o���yZ�C��@��I�17N{WB N6폇�ƨ�M���=���ɆE=[��Q�'D��Y�nJ�N��u��4W
���=8�`��H��`�F�c�ۺ��$ �ʷ3�d#'�]]�	�?"�2��<�oT)B�:�9����\1�FdD�}'��B��#�=�˺�2O��[R������&xͶ��f �
t_�G�G���"��*���(!�kU�20�I����4�L�8�b�&�,q�H��f��e����D0+O�� R7�X��]��9qtD���]�(ݵ��$�I��}t8��>I��7�S���z6��	��5x��q��n�[To�� �Lm�\�\�l�x�J���_�^���ըpr{hc���/K�	���	���5��e�4f6�v����sgE��ș��)�I �<��2-l�OB�Gby�$X����Jv��Ϙ���3�M;�|v�J� uv��徾��e�~���=f��).���&2��\���Bq�-�0m�͑'7��dE����ӫd�&CZ։��'3H��IM��)vCl��4�G�3��N�����n"��l��A��C1��RD���-^��\�m/���xLT�*"i��c���.m�9� G4��̗��Lֲ�/q߈['W�q�Df>�l���(8$:,�@��GeV(>�W$��,��U�s��ȟ��m(#ݛB�v|�Y��g!���a(p��e��9�������"���z=Uz"�&|ak�~��T��&����֎TÂ��VB,J�FC<9�(�ƽ��bqg�9K�q�%��,�tЮr��]{���N�P��[�-� ��I9Z|jTx��8�%X.�Z�U��1�M�M��SC���|�(�?�qˢ�h�]���~�ڹ_���F2��%����Θ���Y�@�Z���Q?�E'�;v��l\ɉ" ���^M���ؐGr���F�*���H���l��+\�Ѿ,��X<��4�����4�DB�*-�����Qq��\���1�����A���7X ����e���p�h#]x�
0�A"����;�5�׀�)+�@�N�Cr�A~0_r�`���r��� RG�Q9�`��)�{d��oEK+$��R��	ƑP�1�8ՙ&�T���8�H�?�Nʿf�b��_�-���~l,�}[��	�1������!W��p�X����5uXz�0���R��:}nd��UW��[ڗ����ݗS���&���8� �t�.�`o�B��7�I7���:�څ��n6�ea�.vE ѡA�l�k´�����14�t�y�2�l��I�a`yE�)]���GY�E�;t��C�2u����ج9��A������qo�K[8�yA�g����f�ٱ�c��S����Ȑ	�'�\pIX*�f�޿�+0\>��B�I�|�����0{=�j�oIV�n`�>�XoK�L�fg`U7b��pu�!7\2	8�N|�r��N;&>���,�b�r�I �C�~�7I.�p�T�ڐ�uJ��:�Q���Z��x�>F$�"�QrI�07�*9+�-���
�Ì�)R���%������J���.�.���ȵ���� z_` R	�Cʹqՙ����P[�b9��"3�D����GT�T�@��l���3�a����<8�l׋��P�'mK��'�}�ґa_4���fIL^<V��e�P+�2����a��=Y�_��A��������6L��S���~���]a�ʎ�%=0��h�����L��|#�3,��-���koe��CʥLX�~ȝh�Y8��+z9�j�F�"O�q.5Lp�������7[)Y����6dLOsJ0��1Ht�{'�� �St/��fA&����>�"_ ��Cb��|8�D�x��� ���j�n��(>5#h�)0�XO��V����쯛����%.e���`ILdF����1M�E5<���p�+��������ӕ�F�i���f�Q�Sv�ʉ�s�9��Y�(a�b	�1�0{7Ԯ��\&�B5��!��A��5��=��MB��A�X���ܫ�w��R
Y�=�3?e�Ys�[K+�M�k�8��1�J�i�j��~�Q�1��LejV���^	n*��g���&�O��JЉg��+�#��������kt@]\���l�&��	p�b�k��!e|��(�o!�5(�t��5��)��uۻJ|�����h�%	�R8]�ۏ�q��͐�K��Ț�a�������)�^ꔐ_�����=�m�ܠή�m��.1�2$�8�Y��3f���a�u_�)v(*�-��6~��sؗ��vH�yŲ��3/�JB<��^���m]VW�CzV<�_��؃�'e�s��o4�@5Y�-	Zuz�y��Q��v�T5�0�[��Nq�2UL4]+�-�A���L��}[HK����{��J[�����/͗�Y�l$�DUjG��&�G����WI�˕xx�|گ�n�NN��4�q�(/�ake^+\~CdU�as��G>������(g�I�e��h$S?~����$�=YG [���Ln�u�rT�;��|��K0��0;������ʣ� Ō���B6��Tf�J�6T�){��\��#3� ��Uԙ��]���gA��O�~��7�yj����mk�GK�s*<P@��S?M�u�!��Ec.},�s�V���yg�N��:�G�]�fr��X�wo%�Fw���*�rˠ<��j7��������4��H��c��x尭F���j�=^A��ڬ�i�E�׊52�OT�1O���A�&P� ���#�_��`G&��h����dy���ۦ�r����Ѧ�����\�b�k�{��ۉ���������g{��z#�x�k�M��{�?��� �q/P#2"G,҉�s�(�V��4�B�%F��)�>���Q�˟��m]�t����&�lRK^�9��4�<��R�j��e���*��6�m��/���8���w��/t�˖s��lH�Χ��Pm��z�����ڎ�y)!�̦/�*=�PXX��T��ma�� d<�!�.�c/�p�>�_?��E��C����&��)�F��>Y��S�5�ҹ^����Y2�|�b���n �,���zmg�yFYyfH�6���'�V(V�s���Y��`S�R���mNF�`���ϗ||#�"Y��Х���(u��b��/��ST��85�$q�t��,t��Y؃��hf��[�!H��
=�6��ȃf�u����k ���G���O��
p4�@��;$~瘧��� ql���4�/_��X��B�I�����\�Ksk��^d4��!�>�+�>$��[�]UY�-�A����feb�r�<�O�5�Aq�@a��D�]�e#~�;�s��, ���،��_6���ݒMK��5+<��kF���m`�/��v7GDYrЙD/�0w�]3&}�2��P���Q�d�h�ȕ]�������tZ��6ze:��yMJ�n��	��
��C�3-�R[��!�D�CrʶE�r��P_U5����\3���E�n�w!Ēj; �=2_d��6��|#��V>���hYф,��o�0��SO״_�L��z�N��"V��lX��o���8C��� /���$|�YcP����#>&Pر?�+Q���t�+j�B.^Z�ɶ�z9�M쪠4xeW�`�(��0q\���W��[<KI��8pc*^Wf)n)�U�TC��7I��x��ғ����Xa��;�q�	��+lbC7���7�A�ܵ��g�	_Z������M�Cy׬�׹�]��]/����rBE�s-9t�*Y�r(6`��<���6��X�RzW����7j�:�fx�^���6��������ܼƭw�w<Y�eΐ�G�0�.��L�uDj+� i$���Y?R�X<R�*c,%1t�;>��f��i�l9�5�b�e�I�Y㫏4��j�e�VǗg 7Ө�8�BXzb�����E�@����h���+�o�RW�H� (���Z�zǺ�
B�U�e��Nʢ�����b�u︄y�7/��AE�=��
7�A�6��j)Z�X9�=:��v��2EtOl��D5�g@$�rf����w��0�qB$�}}R������pk��(�p���`�S�O(�D	�Q�2w�e»���0%Mw��5K�v*��?ޫ
�*1u�Z"C�0�ܠ����x܏�i�i��fhv�P���-Cid:����k%�xr��S�p�P����]��T�d&؂u��� ��9���O�z�@ګ���!5������J����:�>O�;����՝�₳pɟr��{���u֋,D�f����z�,b��8h�&8{ҁ�t��^d\���pL�Q��=�mEP�fӴ���,�􀾦EE��$����؞�����t�7�:�p$T:̴s�.�l���=Ot����0� _�;ag�3d/���#���9J'"X:�����������s��W�F�4,�����cƳKn��k$�j%f��x�a�\g�q�G�؉��@?x:O���%[{cnߪn)vn�c�V��
�����C�NI��/"r�9(�lu����gL�bA���l��-ldr�A�ܜ�F�O<W���?�ri�-�mˢ��73u�s�yɌ��*Q����Et��(&��+-���s �H�����\~�g���L%��a��aE���� ��o���¿毽t";�$�h�q����]ZF����C=�}R��";ܔ֍ir�?lZ�/F����s�-�����-L�՘X��R�X1Y�	o1i��>���W7�0�Ӯ�S=�L�aw ��ܚ��B��=L�$��s�I�p��XY�r��$gNTzc�V�X
S.��)����u�0q�8F����.>#���
�2�P=Ahs�EV>][���T���鐠�m��xa?ͧ*�Y��jTJ2��ʒ/��ڌm*��Ewvb��1��$'��-���$�Q�2�Bk���IF���g�Z��88������2�#q��c���[��n��L��;��"�[/�������"�leC̿V���x�4�#������q�P�@���C��L�V~bV����GAS?����_���D�)���t 	ꉯVY��s4
�[l/�ܷ@��w�����u�_w�Ѫd �~��_�Ƒ��٬U�g.8�?�V��6q��K�Q?��'W:D ����sE�+5����Ȟ����u�}���M��tY��l�s&���}����h��֣�T"�i�)�!c�u�y4�GZ].�R�v�k��>��q�c����,��}C�6uL3}�ʙ6�{^T��,�;�\��r��>b� �X�����(�]W�one�|rf��X��(j_9@o?5s^���ͤҞ14AA�|LL�|��kP4�$���ZWKy�p�����.��t�$�Go�t9ί��	��ۯqiL4f��P�V���r{)��6�԰˧{�s𰁫H�D.�z�H[�^�9XfK�MX3��!����l9�G"/ by]�\���>&�������*{񸱋m|�?�\;»/��FPҘW8�}���Q��#������˪�fD�q�7fd)�5�dxX1(��$�\x�O�/}g&��� ������-��*e��� ���/�"+���i���뫛�]Q�3��*8��OKz�H��������dH�5�,�t!d�uI���>�$Ӈ>�x��o�U1��6�u��7:�X�d���~�����K�b��.[\����I["��eG��fT�c�X�$IlΒ���҆�m�e�}�D�R�N�����i��1�y�MY�_��sF��'8s�i�n^���,V�ы��`� �3���M��ޭa/_olmu/0�h�M�)P ܎j])#!�����;�[�ik/|~����K	3���u�C��j���bj��kN-PF؆rm�g[���	�n�тO�))Sc-�׹ib���qhiE�3����`�U��''��,P֑��2�C~{�խ�"d"s���,��F�h=��dRT�x̶�S���t��	�pgE�0�A"��-�<�9��k��dW�g��@IB��!r�C��:ޢ���l�*�ѭ�-H�@�e�X�-�\��g��;�����j�㌂��G.��Mf)�:������(��gp�� x�g?i�]��'�5���1��B�����<"S���
;�C�_+���#y[��`(OQ�4s�N��N ��laLG \��ģ���u
�[E��U.~�e�ǽ:�<�mOO�՞S�7�Ϣ�sKK�a�RH�p�Ab�ǜMJ3�`���#���z�g����"0�19���<�K�^P{��#{A{�ւ$��rE<�8Q��&�Hq����L8>�ۀ��|���#DHR�����^)�%p��y�	_��Q�P�gu�����~C.��w��e��մ^���<�|�6*�> [����ۛ9�[�8�$�q�c9��.M�q�\�- F�:�Q$
�������xG�lD�H�5m�]i����T��N۠x��L����$�U4=!�p�H�{5�| ���݊m��gs�,�1�ޝ1ͼJ8����x@����n[챲�k-����f��79�*��)� LcJ[p��s�Y�C�!���G���iBV���6������ф�~��_P���B�|s�`���v��!h�	EMh�T���4a㚤h#0�u�nD���*���4K|��2�u�D�7	�,Y��h�7H���z6Czӏ�6��VZ3O~^}�,w���\�/=��J�dfϓ�оoʹ���m�W�~o���dՓ ���F~@!WC�M?
5'`p�`3�����	��[Q5OM7�?� vQ�?�H��,>Y6E|��UQLv+i���&������>o4���C�'��P � Ke��4�x�ߗ����=��7��"�	�+�Qo<H�l^�Gz�V�V�FhN%��آUt�L�W�f�^��/	�Ԥy�5�B�3���%&Yt�ME�r���F�ӫ�_ u܋=yNMe%���K�-��@ �IP���L<H��Ta�K]!��A���F��齣��Y'?,
l�Y��tu���|��kv���r;�Y���6�C����N<2TɄ�dN�_*E���s��j���Wt4���c^B�!	oe��,ŵf�է
!$�L��$�\��B���l�o;�����(
�W�A�0�7nK+I?�uU�	����RY8�<�D��VĄy�15�}��l�4_<gu���(jA/rB)5�.~"L�^Eq.d��3bX�+it�,�E��KѠfg��6.�[�_�S�K�F�h������������x/C�Ov{]����+0s�f�J���b>w<�~X� �F�g&D�ލ�Å7��#���՛U��m�
K���;VC�0�8Ⱥ�D�><�"��,�f��p��.���cL���,VF\���ʢ���_"k�5��2I�{G�����Y��,ƅ�I�b�����g�c�����H��\u���Q��ш F�Ԋ;�5�Kg��9r�xp�-X��sr���4>0^4V}OC�0�d�R������Ս<o��?8S'S?�j*�[!tQ�x��ٙ�o�B�a7�B���m���4w��j��s;IF,�S��h�Ӳ⭲@��1=�Ct����	�Mt�({N�Q���+���V��[�џ*.��H���x5T(=�A�!_�k���tH+3T�A��
���%lvŠ�%>"�!+d.b����k`G!G]Q�w�$�@�CR�+c$m����!�P��s�j(	%�!��O�0Z�yC�@^3Q�j�)p���ܮ�}5��-�F��-vz�ڇ���9�-���fB���AlSW�߂ʸ�!ά��A�,-����e��v`���]o�$|5���ǘ4T�X.!���o���
�l�c���g��M%�� ���U�Ҳ�<�z�ūԗ��H���P��0j�m�Û=���9�)��m�/Kg#w���}�>|����<b���U1s�߱�rj'�Pш�A���f�D����+Q�B.��;��)>MƧ��\����sy@��N�O!��D�f��)]�JV��!mK����v���W1��ݎﲀ���B@��|:�?�w���fhqcęL�I���ri�YZ
ᔢe����-�6���O`�B��p����3�.�ݙ����\���<��{�Y/�H.�$,<��iv�LD~Q�]11V�M@0 %� (Nd�(�:y��Uz�f"���_5r��� ��5��O83O*zhxY1�{7��zS�����6�M��&r�0F��I�>�/��6l,���M?�wA�=\&�]�Y�slY��/�䜩�~uM8�@��Siv�$Ґ��Ĩ��R���^���_8��K��Sdư�6!�=�r`�4��t?�u��#�������c�4�=E�whZc�e�<�V��'#g��SXOV�:��GHM=� ��Ұky�^1p��(���+��U�l9�)�}���
v_1��3�⠈N��䋏]��Bm�k�I��z��Rq��5�����n�6>$�}�XRz�f*�z���$��m����p��掼�n}�3O�=���{���|H@�Ɵ�̶�6��޿	�4�ԛh���� #��z\�Lslw6�r+H�]�t7�ŕ*=;��(������AS؋0�$X��O�M<�ψS�쐌�/��
���(��*�@�g��8$c�C��8���w�S陚���m<I����6`���N����^��M���jx��b_Ku��2o
:��&�-���]������Q��ٮԮ�9n{O��Y�N8di��sd���W�8��N�0+����{RؿEȁ4=�&�c�mq���dg�����a=ɿ�c�m�����/u��!{��\���%"o�]��De���V��,��)�y�{��Vq/ڪ���T�O5�Dв��+l-� �ƌ/���AM_�!��2�fH�4�n����&���7��V ��|�jJ�W4Q�'����+�h���$z�g���9X.ދ�{��/�mg<b8 �����=�&�S�7"���޺��t�$*��7��	��Uq��?�R�ғ?G���>��� m��[[�-�q��LyL��PE�o�e�ʹ���[S
��M�T?�-5��ԡl9NhP���!��DJ�-Xga���M����C@�$�Ě4*���益>�C�����Y#�ܞ�O��-��Y�x�M(����Nմ�H
!���p��Ɓ��{�&����Pũ�.�<�C�=����b�0�~кaI���Yi����;����SX#O��U��-d�$z��%��Q�*m�cb�f�,t�:'nDk�2?	ݬ�[y��*�� �#ɲ�\ƒ\�&����uXed*���F������� &��*;=n��CDtD��mr��K^���n�ۚ��a������^�O�*������i}��6xYl�f����/����Ff�I�d���q|���'ڧ=��<��I]Od�P�r�N�4�}�.q�5��_.U��U�c�"8�i�G��$|dI y�����eC���)Dt&��t��Ҷ��n���
������q^/�~i,K�e�0�c���oZ
���L\D�����^�X�����q�֖:�Y�Bw�
�H�����VS�������� 8�x�t�R��s���K�UՖZ ���i<י#7���A�����*5
]�
�*1r��[X{E��C��Mz�~h��\[�������]T����,a�&-]R�gjMA�T�^���Br�櫆vĠh0 %��5ǯ:��.s$�˪�t~����1�\[���@$�r�����qpf��'���.[B�F���Ou��'��J#��t��4(�9O��F��
�E@ ��w���n�U)G�X�uv��)�ua* �-�\��]�@�Ew��f�����	G"B"��p�����R��L֨S��uj�o���i��������C�� aQ�?͡(�=���ń���F�PO��8~�^N)�ô�pq�S��%�X�	;�5����d�����X�������	�34��M�S���W��+֐G^�Xo�������jtI�igq��gK�z�q��Nq-�>��T��&a뜪]���,z�Hg=�K�];yHzi�"_��x�-��o}���#��{�zRөr�Q�s�% � q�(�&|��o� .��ڌ_�֭���]	xkw��1�
��9V��������+C��]z5�+�� X�b�g|��(B�����<�O�(��l�ȯ�e���'��.i�' �E���;�O-PM" 7t���sq�4B}r���t�Pl22~��U?�¹����_oQ����&�2}�C@�*���u	w��47w~�wH)v-�� t�a]W�Q�8ɗ5��dY�T�_��#'�6f�`t��~��b�O*|E��ƳX��l�c��` �B�Փbpg�.�uX��*+eb�A�����]����ѕ�+��:$��<����HQ�7�yE36\������.hw�ɒ���&�k��rFn^%-�����R�����k�A�ۙ�#�~|�R��#�uJ^eTu����Le9��N3�%v���� �AZO��Fr�K�J|�}��	�Ϝ�F!��	)g��p�y��7ǐz�ғ�L*~-`���F�k�#���.H��/��'���c�(|~����F$�:g&+���ft^��"��\�U�*��m�����	�(�׾�Ym�9��RD�/R�U
����o��l��BǺ���(�\lF��,����ׁ�7HM�a�t��ES�&<ը��~%i��N�@46�|i���m���������W��Ѳ���ҿ�?���Q�R&����겤�1�
����~R�s{��Ƭ��7�F�s'��r�L�>�73]^�<�]�����S#qe���?	k2p"�d�/`̽�����;�5�����3�!�LM4�G02Xb��ˌ>&z��@����BN���˒lň�����B�Z�D>K�����[ڢ���^�e9��k��fW$ �� &9wk͊]Ni������(T��M�f�Э���a�/��7=*&I����c�V�>=(�3�M���/dMRaW��JL�������;괌��9c" ��|{�����k��@��۸���|�4� ���Cg8�xG�&v��u�������S8h�O��AXt�u	)���g:�]�L�Yn�#�����K؛��e���)f,���m�g�"C�82�ה�Zs�㪴��K�"��׏�E���P6%�Kӌn?M�7Iu�������.�.u����ǩ��)(f�W�HOS�NA��g�ӌY��;�2�&�ж���J��E��-�e���C �w0A�#��<H��, Z]�b[��S͝��-����y<����l}�e�E,QPyxr�g)֭D'u���r0�A^$�D��|h�l>;�����~��R�'����j��8`�6{�t�ݓ���us�0���jG�e,��;"f��/��kfu���4��W3��v�W�6}�|�,4<�������j��[8�Dy�p��^}|�~�nJ��q�{�vx�m�c��I�q�����5Ȏ�9y||&a�J%����|˾fS���Կ�X+�Ҹ�`�w�T�6,���p���R�T�l�I��:}@/)pz�ۡ�l��x�!M<\ґcz(�-'��aq�����y;�7��|
N�ENs�_�p��I�Te+�"�����}�^=|����f�&,�~�M(3��H��(�G����q���j��^���j�8��+�,^�s�aC���{��4W��>��@���eO��D3�����C��������>#m0������^M=;�.�W���|����%Z#��i1��]�z���G�Y[a�'�����l_o��^Mu�y�WQ�ܽa�I�9B��\T����&Py����K��X���)�Ǡ=�*��^/kp��s�G=���qk^�K��D���T���R�!����;uDO�=�F���h��<�,PH�������g�*yy���q)ݲ+�d��a�h13�?U#c)�_��a�D���_$˾��X��CE��$]3{gB8j;9�w��~�,�V@��]=�JC���|�H��$ ؍s�̭twK��5iJ+O�9ְ`�Q���7�d[��t�h������w�G�f����,̮�:r:#�8�9�̡��r7�
�fcf~{��\�{r�K�0����V��h�^$[�+�qF�[U?�"n���$��y����I7S,��W��W+C";M ���������X���GTGWz�TF�E���`��8d&H�<|H�s��8��q����M�pج�{��6��1�`R�	h8�3���)a�� =��3Ď�w��`�x��R�x����zwO�5f��+oM��c��U�ִ����ՆV9����g~�{.��X���s��G}9�1P:A�i�����+��^=�=Q�I4��v)ʔi*D[N6BF�{aE�����۝K@}(��r�y2=�wf���N薔����O��-��<����[������*���!Q�k�MQ�ۈ�f+�;�����������uu�����Ǵ�En-�ϫ
�?���k
��qc��ar~T>EVoh��ew=)��\�p��,5?5����9��u�V,L�!����o���{@j7��Y�5C�M��&�;nqs��5�'B��=M�08 ���C�O�@�2�vp�%Ѧ���t�:]���"�R�S��5��:;ƟZٲ���ۇ�y��A�T�O�����@�R���)����.��6;[�c�W��* I,.�^tq��:�!kϬ�	�0S���A��L�e�eSH*E�V���}����3>��f�/� �|p�����O��7$7(i�x@��E~�J5ZY����F�{��ƞ�����"T[�_��?�����j�q�A��8}���E��sq��&��1���8V΄ɤA5'Vk�s����p��� ����-���hڃ{f�#^�>��
\ZbҔ�t7�ۋ�&�%BУ���v�ɯ����qL��u���O��ܚ�Z�SbxҌt2��I@�Q���*p�����P��A;?E蟢�����)-�{Q.q9%�2;���!!`d"��{�3��3w�o R��:�~_�8��ߚ�޺�vZ������}/��qO%���jA�l�h@y�Û��@;��q�-I�`��#08��C�}���d�h���@ ��7����ޭ��cM��e�QcTd͗�+�D�@@�'ܻoY`�k�z�1 YQ�z:M۾�O#��bS�Q��[p�[f����ލ*e,�կ{q���{i���!`�_#>T�#�Ы;G�"k���b|�9�����Y�u�61��ڠr|u�1�Ƨ�pKMO�y5"ҵ�����"�lp�h���/��G�r�Ay� mo���ׅDC��P+�.��e=z��"<c�K:d!P�W7��=��=��Z���ˎ��J��S�rES� Y�m$5��1�B�2@�����}�9�6f�Z�$2�#���?כ"N��a��ߢ4=&�9���¶'ؘ7g ��W�T�{_�8�!E�0s}�����i� >������"�]X.u6��:�m`<(��F��E�dW��E^���~�{6�eM��(�3�O�q�D�5lO�`���: ��
����֨Ly�Tj6���uG1��v�� �>�sv�!���������Y����x��z�$IS����=�,���I�-vф2�P^n��<V���!�E���cpX�EB�b�]܊�Z�R!}j,{yUS+JB�_��_�h�6��+����Y����R.*R�t�4�Td�J���R�4E}=皶�M8�t�?�]Z:A��'�$\=�C�p�-ϲ��ɷ+Np��A�"� �Ȕi���bQ␰��{�N��I�I���s���ky*�^)�#�o׻��Nk^�P�C����:P2��DF�&��r�ƕ���M�L g��;�;���5�W��� �\u�G�X��H\7��C�Cu+�K�嘬�a[���Q���xcV�F��+�A���e1�:i��w��]��G,�ے��d 6mM��0�N�-v��������|��z6"���kU y�GF�&���.\�ذ�;IhkY���,�a�b�����d�ȣ�u�.�ڬ�?��ʘC�B}�TL��h/L�%6�6_��U���w}!q��_2��-���
�ç��н��G�!^�)V��!/�v�*w��đ��;�fU�l�XAa�~L���i��ߙG�Ūu����|��G�U=���)m�A�<�ޏ��.^�4�ПQ7F[�售��p��l�h�wRc��Y�,��M̨���B鲲G�N��8 SH���=�g�V���\�x{�J<���**!�QG2Xj�ċJP;�Hc7(��J�k/v�3���@����G�j�CK1�����)��E��o:b���͒���;���BC0�������hs�L��]�	Y�꽅9,	������3�ĉL�,�v:۰�(t���!����<���4������f	_ƕa����]�����l�B)% ��C�x�̪v����/�+��C�F��GB:�,#yL��'V�_D�pc����{�-&0~yc����_ٹPK�ɃNU.C!aj:/}�µܜ>@�c�$�݅A���#OOA��7�e���)r�d��ư� h-���X;�?u?L����^���G�w�s�b�����s?����@Ø��#���i\n}�����ё�w��EBs(�0ڀK#��H�����"����4&�jQ�iHʁMʺ�'�}+��Y�U�c��s[�V��Aoe��;	CD�X$�a�*�l|�Q�1�$55V�Ma�o
�%4pZy[���2O���`B�¾�Fi��J�Ƭ�����k��(���������Bs_�c�֫]G�a�� �>k5!Y�$ҡ�c��[	ꋤ�5�,�tŰ{�ԝ��@\NҀ��@�sON�r���vUeS��(jb;�m��`��
�!%4�[��z�V��u!�ޏQ������Men ���|�Ն����Vx
���Z�ЋrV�ӧQ�gX��M'�n�!ݸ̨��z�*���[Gk�m�R���r1��-�I��X�|�;p��碵:�����"�0��M+=�ӎ����LS6�B���]�aci�?D�t��K�ϑ�a�74�=��{�rM,�@҆·�x�R���	����P<ף��2��)�)�˄��H��]�	XHm�q�ls�M�w����}e�����褺y��b�^�������>�r���7�'l�LE ���q#eiN�9Y��
�"��a녢9;na��K����D���7�7�uN����[��U�Ѐ�U��5!U	�|����"�'a�*a��$U�'�������;����o�WmXZ��I�����GV��G�'vG����_R�Y�F� �<%M
�yƘC�*(��o	r�5��|;�=(���C����6���6�6��0���gܚ��ex�5Yqo��X������a@�������v(iE�_C�@��A�����	_-z���6��#�]HT��S��>5��-J�{깑�� ��D�h*[Yrib|K&vX��\��h
��pߍ#r+��G3!��0��al�Q���b��F���D�i�Aa��P��R��L�xF��M�8]� ���i�����	�W�Il���~�g�nO�Q�%��%�5� p?��W�@/��f��U�����]K��ysA������'S����H�Y�}z���Ѕ������fOp�/��*Q����{[�M1���Y}��0x})�=��	���7q�d��W�E:�G�J�.~��Ӵ,0�*���\
 �\*��mQ����켆�՟�Χ?/���t��^��c�h�wg�Z.Fr�n��M��<�Kh}�Wя+νt��t=1ƽz��QW��e~�L�)e!�)5W2EƔ[xa�;�lՕ��q
nn�,�Y��_�'¢_���
e\������ �p�ݜ#�-��7�����`�2����?&"���%a�KT+Ks�I�$�Ѹ�Mַ�h6~�F&�D+��ϭ9� LH`I<����[�s=���
�fY W=�C�81�}�kF�{z��������d�ٛz�b�1��c{�ၻ�����c��lT���1�7,�Y�����,�� �.��������|i,����n��M�V���y �fKxC�k(C,\{u��Ƨ1���C>���G]m�����F˶l�����Y�����{�u^�e��֪@e���e�it�z�I��T+�F��y�U��i��Z�6���y=ReV���f�O=�3�s�k%l�"���#4�:������(�8O�-Icg�@^� �!]7�p&*�=IADaiU
W&����~���UoϹ?��sv��8��ZA秔�?��:3q2E�_��R�:�x�Z�f���D]�9w�F>0�_�L����*�Y_ ��4�!ͩ���#A�%�T�Z�BHvZ�j�n~���G���yǃa��dU��F�#�bޅAq�%�Fb)���qOs���c~T�U��;�H�]!-e/�z�fHkL�w��<%r��;�6���Gl��w6�w7�I\!'�&׾3�{q��JA1�\2��%W��Jۺ���{Xwⴵ�vd>;�h�Ŷa�o\�Mf�BuB�e�40� *�LZ��	 �Ldgg�H��{.��}��v'�؆�{�.c;q����_�A��&mQ85���iD�t7���g���[�J�\ �=e��j�:78�Qnh�n�����|�Q�mr�/���u`�Nf�u�,��9�jP���Qʕ�j��IF級W��ǿ<�1��[��*�RH�� "�mq�F����F9�W#9m�T���1h
����E{T%P
�8��9#��O�:��i��D3�B���J�t(!�?7�Jq5��54g��fC�J���,z�WP=����T�(���k^ #�$����ɰ3�qm�p���Yg{�/h��倘q9݇���}�����u�R`�Vw89�uثT� ���F5�$B�䚅��4d��.0*�8f)����v�R�\40�A	]�$��mX�����ڱu��?k��S��j��DN_��I��U�(pv�Tŀ����=l���cz-�](�<��#C��=����+9!�'o
�s��8����Bf��u����u���G��т��뺠���� ggp�.?Uŀ���4��>_����;?cǌ���8W�[��.���l�@j�,I_������}���P8�t��A��g12E'l�sX�������(G��#l81�c�����'#�6�v$O
�w/�UNBXժuI�+:j����h�5n�@$�LC�9���
y�N�����'����4������I�v�Շ�a�,$����[�>N�ι�����"vM̀VR���ha�zduOcMdC4���':�ђ.�e�œ������0�im#Ί
���T&�R&(��=g���3�c�VW���o���;2<��q>����B���]��I/`�?H�3E]"�M���v2,3��GS-1���M���s�:�J��ݮxx}�=ct����L`�ˢߊ��X��{R񮗣�3!_:Ɩ(�`��w�Î5�ʷ�m�~��xE�f;V�E�e����oí*��@��1M(�GB���iĒ�g?����=a֦�w�"ep�y���ޚE�'	J�6�^����S���K�P]QO�����x��3޾g���'ZK6�.��']4x��C�f��m�P�ʃٗ�I4�>.��i�,�=0,�,SF��'w?�Vcc�;8?l6�vy�8�ɶ
ŝH#��ob����@�gG��@vBD��hi�{cȁ�A���FdmFw���+�k�qy������u��4v���~�#%���^���LYA��E�o�R�8s���MG2`0B�����ԇ���+�����M窟rUHD�^v+M�u���*���VE�ܴI}�v?W��ѝ�Х�*%E ��i1L�(����*Ģ㺬��Ej�~r�?rѳr�V�/ƀni�C
�]�0) .�PM���O��H���2���^���H/��>ޠ�z���]����ҀQj('f/Sc����E�@Y�b���Zaj-��>,���~'\�1�9��$M����!:ŋ]"4Oǁ�*q��E^ ��sEl���,�N3���QSG����G��&^�GG�'�����mu�!��!����̊�x��=���Z���#��(�\k�<����	�\4�c*4��?Nk���@E�2p[��!�MxT� S��tz��F��F�����*k�f�%w
$�2�K/L��fpyf`>ґ��ϝԫ4v+Ή���ـ���g9">��@_W�R�k����_���7����ѯ��������w�'��D�L�����ߠ�"�*Fy�=�i|��u�p!Z�X%�P�9��}u�p�E�x}�w�ַK1[�9tB�^֙y��Rl�|�B%B�mx�������A�?ۨ��{��*�W����+�\f����֭	�帴�Q�E��+���`�ܓt����9K�ߎ�Wo"��6�?����O
�*�S-2�ғY{�c1��E^>j3���:C�Ihܓ�RQ�<9ϊb� �r|��� �'5��Z$5~���ۢI���Ȑ��B���ۨ�%G�ˈ���r�<�\�s�FV Й���{��m`䃕�	!��;�1�i������9='�2�@hMe�k��)SIe�ֵQBۀ-h0�&X�s�+K���_�ҹTIpP��OYI��U���M��~��i�6fZc�1VZ -��S��!Q".CR4/�S��1�\+p�:���ʰR2�������>�ubxN��0t�G$=�:������>S�H# ��oM[[��ᆴ�p�M��s�@���,�
�}vn��}w�vjQ��W�h�%�7��͡l5�y�C�p�=o%` V�o8Ωr���/y�Ӥ�sGC�0�C��\�BU�#�3�7��֫%�(�~����,G��f��`�e���4=8�50�d�#�v�ɝ�T�7kge~i�&��{����p>�,
=��`����؜�昬�+)g���p�I��x�Du0+����_���!{��e�����`��C��!Y�
J�+��<�cuK^T�Yi�,�d� &���O#����.���_^oc�{�+�}��(��jV�,��^���r�:B:)G.�r,ܟ(�t�����-?R�lܢ0P�m�lɨ�-�u!˺Yh�}�m�ԇ�������l�m�`��T^�lz:
��)�5�����?x���/�^���E��|��@�w�Zs��i����l�Ժ�1��>�E9�����;� �b�n,�l�;JHǁ#����l�DM�dZeW짆K���-��X����U�>����&�4�T�WT��5a��6�� %�$�BM����	հ�Gs�Nic[�`ک��++~�<��8hy\����j��gEm9+\��P�C�_�I�}��:$��J�Y�D�pA�~F'+���x�����8�h}��
�\/�Х���9H�{�i��N2��lB^ɦ^�z��e�JEy������%�1>6v̄m���',�N��^;]6�,�����@��W�f�I�Ml!��I݃whσ�j5��9�n%�����*�����遒�����#�ls�P]7k�Ǣ��,�
߬b�ԥ���-v��Wg�
��nK2���N��	`���6���U�f��y�O<�L"9�$o��[;^�C�z'J@:�&�1����EpP�ȍ�>�;oa��+6� J�\���!����R�{na�����^C�}h��� �[؝���ܾ�"{~D��n-3y^S��"�XVn��Ū��ϟ*�fi��ߨ	��%������e����i����~��y��aw5�ʽ3VwH�o`�����I�T-� #(Y.��ܳY}Y^�~�o>���[{�y��!cM�ԛ��������bc���� �G:c�h3��`.F
 �V��lw�x%Ed��Y���!,`	�X�i�W-�7�2G�U�q[z��.�-���*�:�[��$N77#�ňl6[�v�#�ه��H�y�o6�a�ɻ�Q��d�=Pڏ������;S�-��fࢍ6���@�ol,f��H���Y���q�������["�V��9G�N��أS:� +<7]�+Ak�oR�XW[̒}R,�\���BV60ur���rl����/��R�O1ׯ!y������Mn���n� U���Os}��m:��JkҐK5���d]+?9k��%|�McC啝3v�i.�uS���\{��1���H~]2�`�yk'O����9�0�U2�6�Ll���m����$��x_B0����B~7������oM�=�mU��xG�-�W�a�4^�r�>k�a"�$F?��FY�9nE��
k����.N����s\��6����L����s��=�-���[|�	�߃=�$�@��@���"�',W��\uC�y��P2�]{Hs������������Ѱ��)����~�1�Jwb-m��bU��}����+���綯�����)Qd��=����0,;CL��cy�L �T�;Sد5��30�Udz�[kO.G#��92��w�t/�af�K?ѷe@���o?��W��9����\�J����]
҅H'�Y<TK,&�7*mF����������]�����0�)am�(�*U��ݕ����c��w��t]�{��gP,3�k-)�{1�K 
`îEIݘ�]�N�!L�▆0�!�_�0A���E�,�b�T-��\�({&	�Zr��1�5�<�!�WCrw�̃[�J��v<��~NU�o�=vB���=/k����23عœ�r�h/f�bW���i�sJ��ɲ��lM� [zc��yF�
�ƅt��]ް�ʴK��alQ�2v��>n�(��:AH�I,-��^�E��Mx�X`M���yK��vt$b�J��S�n+���N��'�z��-] �e"9�_IR����b�6S�)��g>DP��Lm�Q{L 
,L��j������:a�h3q�	&�*�UҞ#�a#� �����(!K+�"$�r�ȧ���Bt(��Bs����ʆ���r�{�5�f�X�Q�Ib]�EZ{�eX�c�,Ȅ9=WL�*��A�]F�EB����@�`�7_��q2�ĒK���q�55H'Sgڝ��DO�z��!	�����PY#�fKMu���'�ݾ�|�4��Qk�\�;�T{�� �%B�Z��Č@�� 9�!b��?-� 3�����gw<$����q��F�Z(jv����u���|�5b��Y`����؀�p�IB� E���:��e�3K�	N�]�ѷ5��@�k�V�V2�8�|�i#�|P|tfֽ�0AYɭ�-�n���\��<��`w�I���,ѻ���B�Z�o^S~K˝qI�p�̘����9
��a���2�����E5V�A"J��\�}V�}ӌO�M�P��ʷ�j±�'�I�̅T�o8Q5U�]Ʒ⮅�n�(Kke\��IgE�(��1�(�Ww��p���0@�edP[q8�u7I���]����0�:���X����T��V�F����}�����T���2f���Z���_��O 2��>����}",4�(ƀ�>��k0�\�K�������k���"��\:�P���ɀ4V`cЗo��μ�E S?Y$�+�b�̑�!�b�t�f�" ��ݰkZ����0Z�*=��a�z�B�;?H0��D��om�i�����@�|���y��EP�e!�� ��컽�i]f
�jH]�+����%[�'Z����| ��kj|sC�Q%��6E<�Cŷ1*g{,��������<bu޾��e�/�E���k��
�[-S�^���2�aas[��\���<�(���c�_+�ש<�M�/�ɪ	��ƫ�$�-�&G���%n�*lKA������l���}=6�y�y*&
|Ϫ����:#��LO�FU��5�w}q�&�7��o���9eŪ����Cz�Kx������ۢA�:4�����_q�]�l�u)X<SeS�[w�R�"^hCF�L��k��?�3피V�i�6��,wI��ԗ��;9$Y{)�����o�
(�kʥ�H}��
���G�n��\��N*���h>�����ToHgJgE��,�aU�n�o��@��{gɃ�7��K�͍��6�0և����i�3��E|�������oou2�0P-�'���L�w���ċִ<����֕�>5yc���
��tQ#*F:NF�Z�m�z�旈d� ��m9PNGܜ�}�q¿��1�Lp��p$;jYs�)���tIc6A��/:֕���_�lQ.��WE�ܚ�I<��E�V��vOܸ��7L��|�^�.�9�͙��,�2��>*R�$2I�D_�^��mw*� �䣲���{jÓ���r���1cj1a�M���ߴCL�a�\ܥ5��4�' ^�{֗�r9�$	�W��ϗ�S+B|� )B�����{0NI>��סI7h^۷O���ҁ)ja%	�2�vWq6�8��!x�Hd�5vՠT��M2��m`]��u��v8�ѿ��N��\p����>�HНU2�� �8�ī�6#���j��9]<oq�`f�yl�y�����W����J�n�(;|�^zc ����a�>樭$BCfi�zH$$�_���YN����D���0�K�������+�c���j� I�ԃ�4��ʳo�E��L���@���!�����kۤ�F Q�[�u�hy�U1�;K����O�cr�%��h��IJ�K��Ȝ�|�dP]��G	HR��rHPt0A1��n5�˸�1�Qƣ���cb��G�Z�m���m���#�N�������=T��������O��t��[�Z�i�W.ɎQ:y�a;ܣ����D?�bL0�|�zD�7�������O9zJO/)���N|��G9v�/��/+}��	�f�����~zs�P���"r���q�/o�0�M��Y1*5{�-�,dR�{���������,�Z�^�'���R�Xs�>�׀x�!m���b���0��6D~b15��E���DTZ�����3M���U��=�"L��Q���蚎��m���Ae�%�p�#���_{VD��(��8/�8�fx�+?(��`;)f��N@4'w����/�ɋRV�Z�L�$�i�`�a�.P�qj�L<�
δ��u����|��)���c�|\���::�����Ofh�"�R��XSR/��;V�#9����(��7=���C8�~"i6k�����R?�����
���4��^�5��3a���F�5?���:����<Evtb%��i\,�R�CKS=e�M��P^�B���Ji�3<Bx�s��b<�"���Q��*�U�X5�5�qʬz�y�M����ui(	����i9=�񐡵�ή��!��%���n�#ҭ���}�\�w�ף�\���t���еb9�z�;F�j���e���.�Ǥ��z#���o_Nt���gn>��P��Rʵ1��L�]��k!%@�ʘ/\C���g�e{�ȯ���oD���9������>TޟzE�^'3�o�]���#��r�/am�>�/��m��-�'[ϩ�\�6`��s�s�����r|:	q�P#%�S5J�p*$�zt��㺟���|{��Ж�m��O� �Z��3��`�}��>�c�7�v_��f��i�._��T��:�7�۾��K�-j-E�y��ت���~��_����X�����	,^���䮶_� t�a��'��$k�ϸ��Z��'b��tF��t�Ԛ�2�{d SU��:��b3`���3k��{#���(�F�Fui��;w/��hϓm^�펼n���ӱ>e�Ts��h�s�q��4_'�~))��v�%-���s�XCOA�X�Я}IHV�������R�*=;I��8�#�`�N�av��I,$Vrd_�e*���<�f��;�`ݱ�B��8�N�P����a��+A�t��>��0$
<بjnyE���4 �e�6�"�H�Q��\3�V �Ng�E\�pow4x�v?7��2�C"�v��e���Sl
`.��@%��fM&�gY$w��y��_֖��@���d��3���e�(e����U-3A�T���>ʭ��/l�����aڢ8p�׶
3)�<��^��_��}g`�2�!t>��D7�li�*U�EȳI[��\E�*v�W�5��5\�mmNL�5�$,�݆���������/�Q�yx�9M����k�����&�I1�j��אk�P_�
�V���`��(��1��K[�,L|��=�a[�:�%w�/�K}���#����R�VdM:� {c�薹_�8�0�$|U�&h�t҄H�kͫ����
}�]�Ԕ�F��^����4�~�K�[	Rw1�;�����'���o���٣� ���8CR��ѱ�/MF�Ĕ�Z���W��_!u'�Y�h�e �f����J��:[��mX'.��bػ��r���^,,�(�a��0a�4v��/bc�%�x��r6�)�'��t'}�sC ��KԸ_���D(�m�(c�b��{����O��F�rћ��G�aKF��S�D�$q�D��Ȟ�]�]��������@Moʁ]�tV��ǒ��]\���ܺ~'V��L'�*G�2�U���>�����4�i0���k�ə�~�I���6"�I�=�n_���#g;e1�mm^��\�+hT�y5�i㋤�o�&{a$W��1��ރ,$)��ل!_X�Ć����l�X�T)���v�� �M��ᑍ����_2��~��f\f��&�LHI���P`���.�A�2���v�����µ)���nB	��OZ^h�W�z�����8�����Q[s�q���ڬr{ >�bD���mh�̙�$��Oq�}ޠ��8OqH�5n %d[-MCBH���wX��B�-��N�.˓��xd8@�q�H��d������'��)9X�)!���aT�2��8�#<=.���z~�|T�Y���u�����G�;c;.A[ò�d��@�5[�/�&�l�]�2b���Ӣwms�bÈ(�A~�4�������Fi`�����*��Z���"�y�6U���7���%%�m��HX�>���K��6'�ږ��I7�b+�m�^�mJߪ��t�T�D�+������9:;�D1�n]�<�J��A��OMS����"F��Cqh2E�gu~�9�֥�o�FU��6�%n�{���w�̥s^�Z���df�h=ϫ4�����(pKK�)y�^�	G�A�&�����щp��R7i^��0��'���ۋ%�U]���,�{�"��Q�g��6gׁE�֯��e9yKpx�.�G�ɸkՔf�L�fD�����ՙ���P>�*��`�\�'P�%^6Aq�w�w>�ra����Q����d3�?�NUh<6^�K��X������/N���ƎbmM�Ȉ�z���i�W�Di�=�-J���6m2�u�D������3P��HG�y����ȅ�Hu�*{���dH0e��gĜ��,A[�V}��Ѫ�'[����d���	zl�fg����0Ї�UH����pI�{{jU]J<r9"����s��Yp6��
�z���ԴcJ�SR�{������e-���o�(�q��@]~��y:��a1�3�	�<�RL�0��Ε?z�y��NA�Qg-�Ʀ�O ��5����b���ty�c�;Jѥ�
���w#Y� Vs�\;SE�'Sr��	uj���52�L�,Po���T���&����G��R��+�<`W9�9��u�n&l~��	�eO� ��{�XN>�T�>tqU��B�}�%:�4���#���JN)�{;uC�m��~dn�{`�b8�����[�_�!��h�1��q���iȖ
�� �Dx�J�v��}�7�
�z�Ӏ� $FTҭ� vŮ�iT�c���>��H-u��h���8݉�q,�6'a� L?�+eWjģ�l'�/H{b���/�f��| ���<��U��i��6�f�B��"a��0 ����l�q<V,)nw��m�����[&d�w����5�ℴGW��O�]}�fo~,	�c^υ�V�<���	��1é�(��ז~~;�}<�[�];U�Qw�����!���M��4�� #W�� g�9�uX|���"�G��)����-%B��m�9z	�	��PzX��gT��wb��j�\��+j�Qd&���Γ�P~��t�Ke��*����@+Ȃq�k��۵�pT���Ig��nɬ�A��o��Ҳ9ea�A�:�a�%Z�3*G":�˸��'f�(/��&�ۡ��Ѽ6�l9͒�,�c]�2��*��X�le]�K+�k�����p���^��+��ΐG��#H�Dɻ���'۶���(Y��׷�*���"&ˎ�&�WD�ww۸�TM�b����EQ�XAV%2��c-����?��:n=Є���!�o@�'�,�}W)
#��Bq��P| ="H^ڇ=JU,SZ���޸Q��s�*%���Z%0���q�ד��_��9H處�BgK�_���S��j]�l �����;x� O"�5�v�g������!� �V�Y5����u~*堾-�\�KT ���Y~��#�Ef܈�\�Q\��Vp�3�_kG���yWXw'(c7�%��V*/��=��S,�Ϥdq��;�+�!��B��>:�S��.���xT��Kq\/$�׊F@֜�n>���d Q�}`��9�y���-34��o����
"�ȸ[F�<�t��������@�ȁ�Cn��	�N��	�=�s�W�/������f-yD/�	CRj������»lKx��!<�OQW_�YՇY�c��{0���Z1����M� *0�JC/I�m
w�ɀ�������A��G��*&���j���
|L��-;)?�}�+AGKA�pz�<�XRR�I���bW$y�S��ڵ�ՆY�)[L�tf�|Iޅ]�u~���ԜNsZ&�������d��ӰX�Szg��n�^��։�F �h�]s���g2�9Q������.��cJ���#f�ױ~>�#�����
��v�;n���F�P�Nwރ��t�:sN��u1�=�f��������ռ��oR���i�[�Wځ�!"`��	}C�&0���ޮ�u���(���
hi�z���e
�\mw�˪�	}UA#-��j���^�r%�cE�,��A6�:"�P��M��9�ls�PGġ>��7:`h���9���f��O�'o�������T�wF�-NJ�rL*}ILZC����qx��BBpW:��T٩���(�H0RY���%�3�Dc�o7�r�ǻ�ԣ�
hx3$�T}�f=佧�����ɂz[E�©�=�-r�=j�fj�H}
3�O�Y5�k��PsSyh~[�B�W@��Qe�pD����(r�Av�I��\0b끘+TwJ�%���*z݅���6H�$���1��i���Xپ(NG=m��]�Dѭ;����t$���@�0�u9�2�e��@s�������Y��=�3��࠺�.�y�O�F6���g[�prG@t�xg��Gxu�T{���t�o�Ev����:�ތ8�@>���Y�uFRI�dۼ̡���[�o��M�_����s�D��,Nb�٧ϻ`}<��6�m��_�pz�j�"�w�9ca%WϨ��N"YDF)�uE�'�lk���](�,|�V�?@t���~&y�,���<�JN�?�X�VLy[�1N�_m^�4;�	���)�b � ��-�6Z���w�����u)�}�i�?���":��Q��� W���3 J��+�0u�	w'��3�z�������Y��Rr�����b�%�����Ն�T��޿��߹{F�5l.�eBddD]K�*h�� O�xȅO�5�G�.i�^sj2�\"�Ŏz$�6H���I��J"�@"���О"��w�JDh=&��]���qJ,��XlOw��UV�	5B�+�ם�Ōځ=殓7*�r��"YX<�Z8O�� ]�n��ʹXyE� 	aU�V�(Z�=[r�x�!�n��f�?n��#�nbN������"6�����ly*�($��T!tk���p�0�&|?_�W�˰��xUJ".[i��5�S���rD�I���4V�"����z�����$���ta�rtf��-"JV,��'���ga��mS���o9C���%��Y_�r�]j�n65�Fr<���N��vݎ�H�j�X��.�d��i:�S�������.�v��ų���֙(����>[�׶���%�ð+�T�M��@�n����ߪ�!��dL�����^��pR}���.R�lL�Yl�7�&�Τ�ͤ<�nn����_F	?�
��B��e3��.�����-ě/��e-r��ݷ�g��쑆���ˤ�I殒z׵�U� �M�\ ��\�\�)��_�
���{�RJd���u�"h�oNX�ɘ�Uی��7\�o�\)�Sr�}Ĭ�\��r�<�$V����2с
������B;�i�O2~{?>;��W�3uǂ���d=<�3W⚰7�%א@=��ہ�>�my_D�7������9��U��eJ�Xnt��V�ͲkO��L���A}���0���.�` �	��EZ��2��6K�}d��=����2��(z�((AY�N_�)���� �hK]�d�*�����Ň�s�����-��.�C|�̻���Zϝo���bw�xˊ�`3����cVv�^urS�X�Q��M���q�[8@�wl��&Hn�3@�;WBYS���n�^6��Y�xY=�[\�&�U0�ų�Н=��7�[qK!F͝~Bx�p�,7�0yrv^�8k���bK,���A��e�P��H���b@,{ڏj���ܿ�{iZ��vI��i�^���˃Yk��x ��$wt �F��pG��	CY���x�<�J��]����mq���׸�\�%H0�giu6��~�LVK��H-@#�-ˁF�/}]�(M+��M�������DB�o�!�#���![z�_q�����?�����,ҁ�*��9+�ڎK��9SK����~a?i���Y|���y�9e=f&�|YW%�3���Y�&�	�=�M�@S�?�9��Rz����i�h�{�����w-�.P7bE*������j Ü�4"D���]�@=��j��E��"ŋ)a���y�%��vc�+��Tփj���c�5Q ������o��%���A�g'@m$]�.�*��qΰ'5RlI�%�@��R���!��Y�FS�T� 5#BwCM��� �Rx��dS�
2�.Ϡ/<�7\�i:�!k�E�+�IR'�FV�Xi��A��.f�"��E�#2�1�����+*c~K�`7D��{�wH�,�/�-�m� x�P
ٛ��f�pX�q�Gq�9b�����W�6����1>2���kwq\d\?`�^D��k��WV��J��=�J�̍��6��D�_�����sX]!��]Ӑ�n�����ޖ��ٴJ����O�w�K]�]�kq�DG��X�z�l��@!}�~�����g��H��fP7?u�cC���S(F�2�x!tgp}Z���FO�^Bz%}�l"��T�f����C�x�ZFsYл��6nǚLc�יI�"��o�l����N�K�!X'�Ieg���́r}���t����`f��<RSP����$e��m��'�>Xōǈ+	���-9"��z�}��;�m&��Nנ����];�N��H�C ��X"�f@�QC���"p�z��#WUB�H�Mԃ�b�[hr `�h!1�s'�?@'O|�kAH�PE����DDrƤ��"9������o#��ڨ?��E�m��$�!}�����/��h���XK��"�=�^S������i�@�D��W������#n�
t��߱U����5(L���Y�
Y��y��jr���˟D�᝼��
|� ��������S��d~����N�%��k7Q��L\1x�{ִcY_����63�!c��6����G[D�? ��;H�4{���h����3�t@a�E�"8�R�q�z٠���@s�#��|Ou���z�Y4�̄�½}LX�Q�G����t>���}&������jQo�O���u*�EF�@�6��I�m�8��A�g,�q�%ʞ������E��-�Y^-�{T�'��\� ����*�~�=�g�܎"���G�֚fA�k#�C�nD0^[6�+�-v!�Z�V�	B �%�T��ߺ��j�P�`���+���v�ͥ�%ԜE`r��������Mp��┎?)�<2�x�d�Q��aڊ��I6)g|��Z�hӯ�u����jh Qc<��]�pg�{�Z�Z��jD!uI*��a��pÁQ��I���h �M��L��ɒj_W�4+i��Xn�������A����.[��8�n����o��Z����5��!�uF�F��F�k�t��򨟅n#�W��N7��y�������	k�};�>�I��}���NNk�!h�(z��T-7o.�g��#4�ZJ��o�z�4Ã�V�V��T�Z�S�8A&];�Z1�9\++�k�����dB�2����~t�
��VI6o�W`rJ�.� ��a��,�B����xE_��B�㗾k�X�	�'Lx����G�'�F�-�Ґ����?3��+9~�� �ñ�ԏ�d�_^mϻ��W4�����Q�0�$����n����2{�p
�m�����X����1���9�8��W|hTߙԟ��&�ܜ2�$r�A��#��}|����&$�)f��Ү�m�3U��z?��@*�!YJH����A�!��!�Oȟ�kC֎�
�h�A��I�ɳ	�����d��H	�6Wl�c�w�o�ba� ps�|/�"THI�
�"a-h������b"=7	����� i_��M��`�5g0�g&y�	\�gM���{�.�*�g�6������q�+�/(����8"3!^��n����w��I��c%���8
	�HB!n_���U�~&.��ܕ�s���P���6v�ߙ�����\߯�V�FӝX���\�U�jd�TC���}�{H{��5�#����5 ���o��s5���u���hP8��'��B��{��M��A,,��0\mn���57�$��&:��0��˩^J1�Ԥ��_j�g�|.Q�_�M=}	���\ϵ���vC�J}P�_0�Z�b��q����'�GV� ��i=UCv� ��� j��sQ����ز�ٟ�|~X!c�x�F| [�ko@�y[�JS�Zr��>�����o�
z��n��T ��hŬ,f'��>jM;$OH�E���dޱ�/�c"�p�Z����֒����;n9��􌦰��o�W
w��'n�ل�ϵ��=��!��# ��u����3U�]�^�Ю�%�{r��ˏ�t��!��B�5l���o�g9Q�pH~~g����(�`�;-oV���XE�1��Z�o��g)6���N�
�,֖������Sz���S�kuF}�B��P��K����Ixk^d�����E�P��an����Z�f���
#�a�̼򈛡����x��KϓC�b�)+�xj ?($|�
l˝�m�`+�{�s	�(a2)�X�Mr"� �:M<��͗B�%
�$L9[�4��ϔ�)}[������4�"|�6d�H�J�>H	�P5�&]��<�x=�@[<1�ۡ�Yc�����µ|<%=O}�B�C�P/��/(�Lo��%5�[��N�Y4��uns��Lo������蕼���p��wO����(s7J���9���(����������6p/4s�5%Ӷ;@p4y�NU"���9hA��`��٫U�^��:���B������`�ϸ�\,�ؠ�$��%6*���r����ao�k�@�_} ��O�b�qa���x1eqQ���1�ݗ}��Ģy9�%�u��l�u�/&��n@-��<���ˍ�L����7,��=����g�������Q?�9�ڥ�v�/�Fΐf����G�v!��l�_#�=6�Ԁ�mz��׋�s�6yn#��V@��F���':��Ӹ��Z-��� ̔5�C���V�hE�l^"�w�F��Y4�Vߘ��hJt����5_����A^��a�� 9�i`j�X�] ��_el���v{4b�V����Gfz�����7��(�m�����/>B_pP�r�9�~IuU��I'_�{9��Q;����|�,ft�[we+�,����L��&���$k����[�R����C��S��J�2�/`z�:��<ʁEX��;�~�Bp��IE���Z�>[�v��3��lL!��]�����#O/i���A�7�=u5OG0��2�򨙗r�l�4Q`OP��{x�)#��y��W}.�B�E�^7d#l^H.�K�i�W��i�e4����O�#�+u#K��,#��Rb_���AM��׹Ν�P�\-2�~=^cTP�<���H�U&f]���0'D��RN��:�QM���I���.$y�2�#�����s�8$�����,c�S��o�d�Ww�����4}�8f���)CAT4&����IDL%��]+��FBN�ؖ��f���*N���4%Bv����� �C\�M�b����D�ۥ(��݋�Q����K\�����ur-�?��oLT[�KwJ#7d?�r�;��X'z�Ow���W�o�yj��d0�	�8P�@��mM*���f�y���D�!�ځ�+��xO��?���j����r� �=
�a�
�� ��F�f�%Gɑ��Eǳ2����Z�5�wޙ��܄Sl~��b-�L������6�_���0{��!@��Ew<?t��j���y�s���9�$tq�1��Mوl��4`�bQTT����ZŐ���w��ئ��bY��5¡P�����L�T�?�ڦ:�u��j��c��&������a�J��զ���V�k�~�ڧ�SZA�k�9G7[\� �~��܋ P�������J��]s>(�x\ ��)�+�Q$�4�F�1(���*�\�����q��Q��j;f����E��� 'ȒW�o+��6kA�#Y�Q�+�`v���c��+c��*���G[#-O0O��v-ћ�1��$�ӼQ�ip�+?��X��m�lѤ�V�G�f��~"H'��Q�C��A��C#N�{I"��>�Zm��+Y�dr�W=�@G�:��ǧ�<t�P�D�K�R���'�I���Ȁ@5��u�qt�����5�**���f�r�B�ax��b4����29qs?W�7��7ׅ`�{��Ԡ���6�~^paA�#܅�Z��g��a����f��s�߃\-����!	�͎,d��4��Y%A�Ii즳���h�&t�I�H�c��?�+a��M]�9-���˗K��{��@uu���à�(&,���"��́� �pS�� �qé�#�b*=�2���j��-��x�=��yQ���qh�^9V�?*$�a ���U}6�=M.��5�>��3�R5�.��Qv���N9��V�5�k�ѷ^��굸�,`�xk��E��tS�M�,��,8�o�|���RV����#�-�԰<M�h��Bz��.����;�L(��7%?�20ya�! }+��fV�ڳɭ�f=H�1���[����ky�
�V��(�_o
EJ�.���L#�8=�S�f��?5� �����=�.����rI!��oV�~x̄��(��{�8��.R-+�����p���6VO�M�uiy��6R[E�1��j�����,f���C-�u�����d��Ro˷��rv�S�<u��|i>�T���M����j!�=��k��K�Y��:v������?��,웧�1t׵�庭<+j��j���w�	}� ��K�u������is�N��Ϯ��y�XF�.��j&�@�h�ǀ�)��N@Y��5���A_���.�BH�W_��!��dIt�7��%��.�v����H.�7JJ����ϠN��l"��]��m��=IG�%�{M���9�>��+���,h��\k[6f!�"/tCa������ݜ�2U���Zk!��eY�蓤�Qo/�Jj�n攟0˞_��O>�
f����*�rs5�������;4ln�����Ԋl��և������m��l�K(���S�-C��?k��<������)��# �m��ɼ����q\�����E$���7�=$�ۚ5�������p�X�c2�ؗ�s~�M�&��$�i�9b�Z���Q4Xؖ�nk�4�d�K���1����[�>�ń�q�[�]����<���i}�LA�x��ݺr_��X%�%�-�����TWi�����FO�C���.,�}^a��RV��-����90L��o$��y�U7�mw���;��=00��!�4��k�~{��5�Kj�;?�C��ƜIǎ�'�����w��)��j�C���AD�k�Gm�h<4jSS��،M]�ƥ����]u��a�{�%<�}��ώI,�:kdxk�&wa����G��uk����h~�/H�s5��x6�|,���"��{��8�� >7��@�5A �5�>��`̤�/�d.��̋N`��b�D�K�:��RV*����I��Gي�oN���"p0��|Bε�:�}3[��-�|�ۜ�5-9�y�o&��*�b����(���e*2����h�v'����`�A���wA��`��Bĩ�$:���� �(�@=_�0Mr/O�����O�qF��a�fs��.��@Sf�>�Bf�Þ����cV���ǽ���<܌��x���g�M�E҆����hn���nlM�~XJ���4#_��^\,c�iL����&{�2p/�PlL*���P�k鯓#}E�������vX|�`Z�_4����_$�a˲5�p_��bGG��H�J#0����۱�,O]�������H�n6Rϯ�t�Ft;Ө����!ŤEgޣ��F�{v�no�2u��2
84�m��
k5f�?���9��c�6MP�^ϧ��.�A@�z p�F�؛y"���pWT�3>Sf�@d��� U��?��7ot�jmyJX���K[6��D#� R�͂���a���c�sڻ�b���thO����2}�h�7
'�����@��q5�#�n��+����Rz@G<d���3����'��u������e�9�g�zQ�f&"�Ï�mݴ�9ɟ��?2� ��E ��E�;��c������7Y�:�����}�*"���|n����	�}`g���K�t�{p�wK'B�Bp�r\�Εw����\,�� �>l�"wd�/G}�-�������2���^(�?� �4F� ww�5� �b�$I4�T��P^K��+L
���H��1���|R�`�F�D�$�v0�Ha/�f�� �o%*���T�U$�a�t�ڬ蘻��|Ұ@��~���:�P�!P���r�
���O���Z$�*1qdaP���;1��5� 1>5�m��<�?�d�v�+Ӝ�xL��I�y��ΕQ����Y��*�	Q��w���䠜�7�ҍ��JYg���>>���U��{M����0�-�VK�J=�3O��~��#-�c�!��g���S##@M�^8��t��A�J��m��;x��@���d���H&�C�:��	��p�v�ԁ�t�ė���R$b����M���u�ҋ��˭���M� �=�Zk��M\�~�>}�U#Q1z��h��8�Z7�x�8�滋�F��+xj�%O�_�����h]sj6,u�����ۤ)�>��1L����l���5w��|��#�~���n ��3�bÍD ~���N��^z_fEK�����S99Z�?ċ�}�� �� W���*1�>�:��E�(�ã@D)֞���[!��η2y��� -N�t�=�d�ή�Kuq������[;��G�?�$��{z!T�ll�}җ�Aҩ0�s�7EE��W��-�(0�R�!�+w�1�m][�S�W9���B|7������o����w���5���;�vƾ�?�Js2�ݯ�$w�n��;�$7+Ύ�о�>�a3�]?S��w���n�$S��f�U�5��1�{���0��&2K���c�Ps|c�0�&��E�G?&?X����u�%���Z��
�?l}�H7���s󚿝8�FY�[��U�Ӳg���D�d9�T	��%-c���ߔ|�mc+�偽�"-��Ф�41��l<�#������	�d�A��{f8�:<���,�S����A�B݁��(�)Fj���<�A-���a/��PX�xh[�p����:�o=�i�P"��)��`,��/O�u4#�c
j둷O���8�����N���A�0�4I��2P�0--���G]��^�K>-��q��ԔO:�����<<�=|�))�/jT�g�� �~�� O��;C*.fR��J� ���(jAp6�"���s��MZx���%���t���q]~9�k�.��J���8�6-l��A8���j���{�D*�K6�SC��,B����_B,V'EN�97��y=��ne,�6����_!|�dV��ȩ�d�o��?�����ìKH4���L�z�L�%7�����r�I4���A-���oL_��� *L�JH֏����5{4����R�;�A��O�-M^슪͘�{�j��p9�e���!(�?�)���Ĩʤ,��=���T%H�ډ��������j?'i�,i6��/ء=Ңwg�Y~�aWma.`��anC�b�<�8���"��:�j�EEC����;��bgLX�%���Z
�9��Xo�[	����B�i?"�O�ݐ�\���H��3x+��
��쫢���D�L΄LQ�F2���J�v��q��+t=+�������04}�M�T^���Lм�:��`=DE�(S��r��AQN�ԁ����Lٔ�uu������_�Ai5����Db����N�����6٫�h��*P:��{�~�vID@71`�16���	�C��.l�IEa�-'���H&��j��� ���2,�p��
�97��\	��������op��-���vAd�����,��h&���T�<�
ZM�N�Wȭ�z
b�c�ۡ��'^���~�~R�:,,0h���E�c�� ���������,Ϛ�7��3=�jo-���N���G%��4
��d<(���*۰����,ݲ{���K��u��X�U�P���ƀׅ'Q�����6�ҽ��!�%�n�ā��2�=7zλ��W`�i�)� �H���Jψ��T�O��"��H3�5��[<��m	�~%���Vb�L+lB�&G���焺�p6��7 Y�~~�//wC�޹
��y�K䚈ގMF���pg��9<�;�n��]����̓<�:(� g�s�k����X���\�����Q*�w왼ٻ(3�u7��u� <>A@�C��}���-�T$�b7�Y�W���h��T�i����s���#?SLQ��?���~�" f.��7�><x�~aҝ�uh�������m��F�7��I���f�d�t*ܫv2�/p�i̩�p<[�oxȀ�J��ƌ/����_�}N���K�����B(���8k��h��0���Ht�Q�oeqn��N: x���#P[�r�΀�3k2I���2�:�����#{;�pjb��%&VDGOmg���ӂ{%}�����7�*���&�FL$�-�s����^���!��m�����3&�[��d���Ps ��g	�m˪f��T���ƛ�%�I�����F�%��Nv���h��~��)q�~8������(�H& et�j o[G/?��P��]]��/K#/C6d����.C%���A �*;�5�"�n�T K³�i*�͗S3G<A�����vI1$ -��o{�9�;�pQ�,�-��H�-{g� �v��)�f���̋5����i9~j|���ƭ���"�r:���Є���5�6�D��[��bH�tM{q��?[�M����4y}Εt�Ǘ�f������?�?�����������H�Hl�UU[ ��Ҍ��q������T�� �f��e��I��,�.�z� b�F���~�G�mh�d�f�N�
k���Ғ�o541Ԝ�ֆ�D'�d��}Xc'%:V� k,�?q�o��u5C" ք�t�l�tB80�-�Xi؊T�|ES"�^6~�:�AErTd�9����-�_�������\ml6$ɣ�����#(�c	8��XJ�4��~,��D$��� #�]g�=�2nx	��|d����$�B"�S��r����xA��(��W�ǟ7�Ԣ۩uހ����ѹ������?۠�R�2�j��_��pr�k�^��7��RFH��β�3�-��Y�s���۶�FH��7��-�	_*�r�>��m��ވ�薛��^ �{����~���gZf�;I�~���Z�����1o�Y��ؐ���D���v�r%lpr/[vA�`}��Q̀���%�k���3�*kx�?����"t���#��r�4�p8��a
��8tB'7W lG���+�S��'#���p(�V}
�Ň6����A+��՗�N��K�f2Qz�}nA0�m����YmnXB�uu��޳�9�N _��l--�	B�)"+,�0�Z�����l6��AR�S��<Z-8�(H �d���\]ރ�(/.S���hDXu��l~àꍭ��˟���ZW���ť��(��Q+At�*�{�nd"@�[s[�t��e�/A5�L�r���)V���k���"(�D`o��T<f/8�mK}�;�1�U��2X/�6�|�]3}D�	O��Qf[��q0��y�=���������2�����4���
�s�1�,_��8̽R�*z)�T�4�����*�'���:��	S8}t�ڷP�X�X݁j���I.����c|� ]�uD�|vc���վ�Ĕ��e�f����3�ϻ��,t��_�k��b�(���eဎ����Q��7��0�p
�ɿ2<Vk�])ǮR۬zO�1�]v�*S�9;��r>%������YI`�rg�� z�]5��FJ�w#G�87-E�0����3v�T��XX�2b����@���\ٍ���Fz�t���y��!��+sC'����L� ������{9�$FІd�R�A�}��m���j.�p�D�Q��(;h��}+�[���!u��Ю{XiD��x�4�؊#�/�����[I��*i�V�`>)ߌ�K�jg��Z���2�n�-0��G�Pͪ6�g����ꝗ���I_圵nR�Kv$�O�J~K���KUEs�N��ӱ���S0�/�Щ�)��2/^���������y�
��ހ�(/��f~���q@��ȼI®���)ˣ���|�0�V�sJ�H^���0T|~gt���,�*$t�xy�����Cq^�ү+��oD����;��"u��f��p������c�֚�D�2ָ�,H��g{��z��o�ᑱǲD�"��%�d�bG��pʟ����&7���Os�|!%�̛���W�E?���++Yҽ@�!�E�_T<Pe���}[Sv��[2��%Czmy�F�O�	!z�߳������G��o���֍n�1��Y|�TuNA��v��P��y�mB��'�2>�LQ��o�(�I�pZ~.���� GN�}�A�{M��[�!��.�I�UQ ��W���[�8��b����a]�)�@��5��B�*d�4�W��B�W�%ND�grd �oִVr5���T�|JN�yF]˺����ہ����3e�y�$�;	��
۫�d1�Pz��~�K�i(Pl���v|��m�}�RK��(R�h뒣p�pr�����n�Y����'�>��B�1M E[S��nQ��Ժ���%��%S%�j-N���w��T�R��=0<ω�BƱb�.Y<@I�����l�a�m�K�M���R���;l�����7��T_ڭ^jv�o~ �?i��|��C*"�_��񷙕���.���Օs��C~3��'#X�Q�:CZ1ᣗ���3ō�}�?rV�z�������T��5�"�؊ڀ�'n����,l��ש�y�[a�`����&\"�
r�yI��e��/���x���D�O��ya"�$f��[���V����� pѾTZV���e��+%�S�)H�?�vg�o��겍� ������Ff��q��������]����bXf�\i�����!
�9Nk�LS�x��b ɐ|S���NmpD6�q�S��=�.� �R�ƽ�O����<S)sx*�����7ޙe�#�r6��"Ն�v�!��1��D::�k�E,�PU�����T�8��0F@���v# �/��s��)�.�ꯛ�^��,	f�K���K���|*8jՠ����>5�Y��2mH�B��hO��gc��+9��J�i�̈�8��HC	�w�'O4eܟ���Lr|�a�/O��%Pn�)�V��7u�*2.��i:e}5��2�%]��\ΰ~?Ɏ
b�E���p�K- �* OJ���'Yx�a�3�΢�
��<s�W��,}�Q�ʖwk���^���?����vod|�p!Zg��YH\��+������w�5��O�1)/��N�9C��/i��*NO���G���2��0�n.�jZq;5� ���K�]A�V�Bge_�kV?Lv'�� ������ 6Ŕ\sSoM>��.�]�ߒ������݂uF7(<�u^`c�I�}��O��.�+m��C13U��;�<[�v���
�QO�)����A~4�Fl���EԶbf���~�*8K�Il�E�;L=0"��elDTr�ɲX��.t�m�os0����}�A)9����T�Q�:�h�dM�����w@��S?���:Z��o�P�km�&!T�J9L�O����0߂>���eNݸd�:֨,�d�n9p��-����0��z���>�&��`w��G=D����[�9E�a�8ͪ >$��"�����Z�m��)�,,����9UgK)�E^Gs��!;��.���j�����X���\sD����1����4j>�X�K|��^]6ά^��O��b4���n��C�x�퉤2v¡[����׀o���G�#����v`�W�����VX:t��jB��s"�����T�#��|>8���]���z����g�A�1g@��բBe�#su%^��l���ω��P��9�}�����'��dhᇼ����A��eUk�
 �2�9� �	�u�ħ��Dp4�he��Z�p��������
��!0�n��sj�נ�m�_����Jv:����X�ɰ��vj�p��[n��?��(��'�WZgT�(Ɂ�u�H9ӗ�)�aq�
�Q�Y��~Zg�᧊N��lޙ-M*��:��~��=8V�w��������V�|��Ѿx=�jm%�kn��F�4�N -@�� #	g�>IX,I���zR�*�Cq��>:�2TK��r�U���E�c����iRR����(���bsY(�ɻe�SU�p�N�h�E��D8��t�tZ��bj,�<�8]B:q���3�(`��50)q,A�}�Du�J7��@�Uw+����y�e�M�@Ĳl7��f�Y�K�_�=qBI9~]X�W޹�e��6/QwI����b���>�2U���By�I���I5�|UB���pK#�q5��@)t��_f��B��RZ;�U�l~駁U�[ft��ai� t�vo��8�����۵��Z��(���y�v��
x'W���x+R̘=��,j-[�����ȼ��!�"�D���ё8�8��㍷�6�_*3�J{ԉ��֡�q$��E��MU�]���[�(�3�h[{�R2���؇�yW��Z�{�`>`��v�1k]~g�Rڮ:3U�({��d-;�L�� q�
�w�;c�r�p�"pZ�:M���sZ��|/x�y����v��?�s<����f�p��Tz!��Ik��2J��x���ŤG�$���݊K�;\�9��f�k៞0u5'UK�-Ǟ	��k\�E�)d���wenB�oC;'� ���E6�ܶ�e?G�z�w1�ㄝ��[1#N�Ì�aj7��r�A�w�gܙ ��G����R�'�P��p��T͸��˛V,���f�3L����s<�6%߂��&�4A�'�zH���!/��8*�[L�Z�`gMX������E����5��+ʐg��q��Op�]U���ZC.e7G�\��(}�
��d��ش7X�� �u��e0�2JvWt~9������9i���J�
�PrHj2G�b�=��̸��*�./���Ua�P>5����N�_β��9�Ư������rCi��(�N��`/�A���ǹ@�ͩ]�T�Hf���`��x���v���� ��[���C{�,�c+�Ds�0�<"��hU%ֳ`{ :���#�ؐ�!_��<\4��A�zv�
�8����u�ڪ�������4���H�H�U�led�d���[�H$�B`�I}oM����|	d�r�(��6�^e2C�w���23�]zr��VQ?��͈`��I�I�$���t�t�M��?��%����LY@�&�V{�%��*/dN�h��}��'�,���8p�T����xNH��Eº��Q&).�Jf�l%���Ԕ$M��=�b��� Fd���Vm��CM=x��_v	oΎ���CB�v�d�����P�����1&�tG���?EX?��x6���Q�΍�<�����):��CQ�x���Zi�B<W.��ZJ�1#Vlr�0�H8���#��oYb_9&�2cA'�JiTy14����������D6��Y=3����3�E��D���O�:�SmA�s��᚜�B�fC��`^�0s��df�¥M݋������|=/x����E�M��5�,�-��ն3gÇ������k7u�nN,�����l�z��MQ���������k��8̽tH'R��t��}^<�7�ߏ��M�U��ѰÊ3�|�
�4&D\)�v�ͤ�c��3�_T�����p\�(�Y�%�f,�5fK�]~��Q�Ǡ��m{X�����.Eߜ���"���K�e�l�[
Bv�+D���hˆ��O�C������.<	��]^J��~J�9��*��M����#0QA���'Ɋ�3�f)� �ō����i�j������}���zA��A�R���Җ��գ��:�|G����s��샜w=��א_>l������-��Y�h���3��j���x��l	���s��c|������B�I�明i�B"1.�|�����3�on�I&~� i�����Y�@#"=���Ŧ��Z�)�`�k�'�`���)��� ' 2w�"�/�^0*,�y�t��v��{�a��N��b�Y��ܒ;�6��<�|���2��KK �p)?�;N�{��C{��F3#����Xz��_/P~K�����'�̘��CM��^Z��T����P�/M�f�/�JV{U+�MB�j�{�1��'��{��YV��c��)��*F������� �p1K�F�O�-v�Te.�q��J�MK7@0�eiB��KA�}QL�M����.��[̜�"[9:h�TˎǂE��+�#V:]j�-�β�c�k��{��+�����?��X���G���_�h��]�6V�&)B��@0
zC
4�d�W�v�c�.Bw�++":�5X����_��m�Q� �����,A�Rъ|�١��Z6-���`�0�
~z��V��'ݙ������ݦR-t��|��hHN�F�7��(�{Y�RM��/q���`	\�eFP6x&���.���}_�67c-���]nJ��{p#�����_&�.�WW� ��c?�vчjmg8�����LG�|< E�Ǔ�oL����v��x5�ڟ�\?���	��YnS�Y�u��tcg�؀��L;nxW�_�e�_��X]�j0:�Ml��Ńv�N�0V#d~�{S�����̌a�|g��i�O�oR�dW�u�O�6�xu|�v)��̉�6�G����5��
�`RF�Ҿ1S~�S���l��e�w��u�ٹ����{�Du�ɜ(v�y�a��S01���Na�cb�Rd�7�>ifi-�t����(��7sC	 B��P
gY'j�������ϘY���`qd����~p�2vq
"�P&qS}'%@�>��eX�O~�'��i�"5��l�=��}���f�����r�d5Ӥ��8������/iA�s�F3aG�ϓ�A�m��Qi��e,�Lq�>������Uxg��C�U����ͨg3��(CE��$,� f����#�{ab�S�~�d ���j�%O��*vxN�H Ƭv�ܑܵi�n�U�D)��m���J����5�����AkVY�\�'n��@8�!�+c<v>��As�E~���s����פ�,v�[s���!�ww�+�7��~��`5��{���rU��5C�}���x�������b��b�h7d<ٵ�B0˂k��%�U͈r(T�Ɋ�*0�^dz�i��Ց�C��Y# ���5��f�ǷW����q/'Ll�$�mk7/��i���_�ؘ�:�߲z��o	?�(��&!볶�:�΢�q�A�F�C������a�bvA[m�DnKՌ��R��l�9��K�׵�;k~-C�������sdʊ1�_� ��\J���s��M���mID�yÊw0k��h��^_hY��=��b��Q��]Hr1�YH�d� �ݒc���~����[��P�&#Z)^�b���\�6�@�e}�O�<�@��*���@`v���
�"T��e��<�BaA������|L�j��^I� ����=��^1�K� ����4癆�j� }����1��Z%������ҳyε�U|��9���'�X՚���*<-�/ߌ��,��[��Yz���(�@72���/��f����Y�"�%��>	j���3EڬIu��ie�u	�;�m�`��ࢆ�U�����r�����j�|n������u�3��G2r�6� d@�T,V�X�՗��Ԍ�J�^��+�z��YS��SmS�Fp1����;>�T%�d����������xb88�?]�����9��	��BLxQ�5U<4�j�˂�l�R=E��tQ�<��[X_>:)�Jx����@��cQ��K��ݯa)�R������Z��7�?��
�M!�'K���8|�yK���~�nB�El�96Y�y��l��@�?�v�W����#� ?��qDi��ފ�?��^"2�n��s n�)K��F�{�IZ���)۪Ik0�>Y�9�E����~9�LΚ�Ӄ<(OV۩�����rN����G�#�QQ΂�O��ֆ�B�"��-�h~�G��n�`�U�W��	1>����W������ ����
|�;�oT�Y'�j��VX�[`ɟ��U���.z���<9���4	���a{���8�0bU?��44����/;���,���υ�+Q�(��ޤ���z��C�z�i�n�7������U(�dȐc*�}�-�!/�(p��v?�6ص'��=K�eY�d���K۲
q�r������^����s3�S�Vow���.�租�x�"e,�O'��)k���Imx�4dM��ʶ��";7�up�p<�+�l ���3ҟib��br`ha���!e�@`�
��rC�C��Q]�3���n|�UO�j,���gf�D�*�ͳ�;�	%\�~�*LNe�8^r>���q��*�#;j���:�!q���IT���!b?��N�$���GȽA\CE�Ȭ+j^�����bm���PE�WVF��\����ΆQ��0Dq?�G-�Ak��W\��=˲����^gq����SH��:�k8%�Г�Er�>KC2��9� �U<�7��Fz�����2��Fd~�	v.�s�Ycn�����D��a�>.T���0�ҵ��窓H�|�6���)��\��
�^�a��Ǒ<q!��"sT":�_/�����j��u^����|��U��~>�T��Hr�FPS`�I�Y��x5�M0@�Ax�,p�H>�ݞrV �t+敺��/��$�XXⳙ23�����$Z�kÑ�;��|���e��V^;���Csʗ|�x�p�X9�. $�Ӳ�F��y��(˥j#ђ�ޓ�ȇ�)��k��VH?Ԙ
��rj;�'nUQ�d����$�I�	�/4{Rx>Ç��QJ�p��Y��65���g
��F~x�
�j�}�Y�lH�m����s@t�k���y�Ѥ�`he#�Д̜�t��G���V����(ג�h�HC��1�<>��7G��!��ɣ�۴z�:�v���f䱴��~���3�����?+.�,[�/�~�w����^Z�J[㾨�(rIj�t��F �Uoh������Vg���G)����5Y�~����{�v��ј��Cܶ�+���a,K���v�	)����̣{C�N�n��e�9����f�tL�D�N�¦9{��C����\���nm�7\�3$��O�����d!�|�G0)�?9�M4��*�-D�i�خ
��AM!���!�����4S$���>�� ��c=U4�b Wz�Nj���%9�����~|���+�6��ɉ�,q�[��G@��8��?Ⳍ��ʾC��;�"�#(B`����lq��������a:��RaiOw�r�>ර��v+迨Փ��K�������M��]#�o��><�2�y*���|9���Ӛs`�