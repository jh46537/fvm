��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z� ����v�?uf���z"X�:RN>����x�*���͘�䁺�^�������d���R���1�D)Q|��(��v��ǭ���z�+r�x�>AVv���z��"��QG\*t�����*����J'����<ς������`|ݯ��	�03Шq��+Bb��Y}���{�2#�1d������!�Ws���!��Q�zB�$�e�4��kS����$� �&%�_��ZV�i����%�a��ld�� "��A�?��p�1��o}0m%A`s0�����q�Q{wz��%Gl��.��K/e��C��4ך���o>�xKz��]�^�_!��v�r��kCas��聙g~���z�}%Nt�h�Rm�2�L�nϏ�;7��bD˒_8Y�T��<���]�_�a�h���r�������F}��V��$�=~c��!%)�a)enq\NT8��G�����?R�i����Y�c0�+7��n�0*��%�k���H��7�g�,�K+�xm������~3�O'$4�r�=�$�)�",6�C�i���V̱l�p�zAqPk��a��
X͓-��.���=pY)*"Aާ�b>l&�bg-󙝠UEŨ-�K{H�V�/���M#"����Y7Аm@j7���qxOV��Y1k����m)��������t�mÁ9f��`c��K*Qq����#����6�ϻ���ќ���{(K�����=ր���K��S>?D��e�c����N*CbIoj��z0���۫�ʖ�rZ�=9V��'�<,L�M��ǳ����r2��'~+�YB￷]+��#F�D<&��_�N@������ ��.����~4Z�P�� �ǚ5v�/�Z~�e8��Ӟ�NN�w�� �S����x���JT��J6�B���q��<���Pl�ײꔚ�X�rG"���1<I�>��~=1?4<���U)�B�Ď�<���-S罢5�Ԁ�$�P���b�A������A��#����A�z��%���O?E{�]}g����LgϛC�o:���Q?�A8�gr�V��r	d�����L��/�x��ec��6��Y�'`��9���ϯ��Yy.	���Z��2�u��/�����&�b"2�+w�nVɽ�dB*1�q9��+=�L$0)�*h���y�y�G��W�#���Mզ�O�q<>_�Ӯ=�-Ji�����
���j���r%K=S��5m�\���I(���`�|vo�n�Y3l�<�Mqń��]y��1Ym�v�\�dO�iyǏ��x͂�rZ�!��&/�B�
��pO���B���{`�.-D�7"'�3qO<<�ۂ�I�D@<F�M�*	 Mz&*�ⷐ�zg���b�ܼ��[� �{�ۡk	��$Mtɳ:Eߔ��##�%�,��^=9�Ծ�.��l\�X+O�uFB��<�p21֚m�CK��];D�����=Q�ܕ�㔡��e��@�������3�K��p�o�b9G�n�~��+q��d�zaJ�Iɳ�wL��.�Et���-��|/��ʼ��H�s���Jk����`�5�|:�zD���9R�읟��<sf�e��ם��G�<,�QYܘ �m���ȑ�w��S�%Y�9ůҕ	��Cx����E^�ګ���ė������T*	���]��^?���]��.���1�!B<4D�`�]�Y;���*�U����t��"�6��$ob�h;
�;+j���l^Y���|�� ���f9U��]�G�G�ñb��$?/�4����b��|/�󬝸��b[��,�p�W�b��?��7��������~#gz�9� �}("����a]�����^Ul�r���Q���%Z�ݡ�;�
!���C�w���]�+��'��W���&���|�f�MKf�ø��$2u�5�Y��t�g&^���d�XD��$�8�S��֝��Y���X�b�ϧ5AA%VK~쐗;�靯��f4� ��Kq�(����!)�/e������7&\���/�N΋�gf�}�<�>��ߡ����sivƊ�=ߘ�d�g��y�n�\�s�Ax�[�k\�ěn���%əL1kI�2�N�ɝ4C�zګ�[G�C���������k�
O�2~E�G
tM���i��K�5��I���R�ua+�{��J	���a����Y�8-��v�z9oY�W�7E�2�x���#��O�'S���Q�cc���Ӟ��f�,&V%�!����FDt2Y�p$���ͅ\���܇2���վ�{d��������͹<�s��T���ZY�{��/�����NT��хY�p����+�]�!�������H����0^����iZ룃���8�K+o����W���Ԭ)�۹���	r���ÞEt1YKˋni�.u�(ĝ#��J���-z���	g5M&��Vd�Q(���G�£$����@?r!)'*�a�i�q���a�ޔ�ڄ%R�3��ً�IT��	K[z(���>h:�90��y_ʻ>Z��*��ڜ@sLΆ�"m��G���Gpm�C	�0��q~����||TB����;j�r�x��X��]����Ȩ������(��̱�:l3�ܲx�}��G(�c�iX����
�gtN0M�2���۱����uz�{R��)�g�_gF�"�.Rꣾ��d9�d@������QF�^���)b�j�"���8�
�z��i���j�����4��/̫{���*��(�3u[�k�t�\	>���cJ2Y?�H�`��'n�2�i�7ހO}��,��҅�Ҥ�]E�z�=�:k��8�����}���j�H*��x���찙�F�ZX�9��8^˘6}�,Y��ݜQ6V����5ּ�hCOt
k���u�қ.��I�2֘x1��Q��ip`kk�O�������"=rk��8����P(�..)v����s�voܐkӠ�_a?�+}w�\�acʲ� ɺ v(z�ٺ>�]Z��bZ�NLѺ�Y-��M �F���X���Q�n*����N7Xn�"o� }��f�[�q/�}�ef��|ҪA[樘rA;��JPՕ��Y;�	��f.��4=��N.�G����f����x#��:d�˩�##�<6��5"��*v��k�/�.��V⬢��� ˑm�h����!�\������-��w�dG��?Q�ao|����x�^[1�V�]Ž���ֶ�F�E�_g=<Ra�' �ŧ�W
{��*��6�*7M���է�ߑ�Q���v_1�����f%�O5���
蚘;z�k�xt~ff�=P�	]
E<n���Z�>[}u�ю��7[�\���� K!/G�*N�+�^`�*������W�~5���p�+A�}M��<�=�*&�a�1%I�Ǩ3� �py�e�<�]��(ٞ%V��<�n�#��3�n>t��W7��umY���0�0B�?�����W���v�jK�Ų}�C-/����:�[d^�r�9 Yg�v�F�%�]��b��V{�L'��̒M�wt\m�b� �:�j� q�S�����}r}�����ƛ�[�;>b�*F
w���T\��ܾ+�I=9FԐ�vD�v%��n񣉹e�k�jM5|4�rA-X�ܯ��;N���B�ە �:��@A+��ppT��ۊ�9 �&H����&)p���:���A�9LE�a,��2�oaR�\lBi�Ws@�3j����
�ԝA�_�tR@�i���6�bs9ԉ��h�>��;�议�K��� �K���GJ����6���$�g%J��*+�1W
�d��(1��}�M���-(p�k۸��#�RMהD��Q H��B(���w������d�"?���^�w�@KitH���l.�d���WW��F�ߋհI��gX��̽,�w����wJ��f�P|:s�9b���?H����n����IM�[�)���T���wO�F��+��hK-]q�Y��hH( P�ޯ[�H `�w�C���������۾���m}kM�>mDÕ\H���4���EN8&����;���(Z��h�Ufe��A v�$h���e�R)"4M^��?j<�.����3��dl��?��2����q��SDK��w�i��|����j��6���:=r�o�S{,�K����{��gŭ�2�z����?
����H!��*	���+ʑX7H�P��
�𰔺	���Z4oPb���N��k����}��u��w��`�Mx=�,�L��$�n�a���Y	/�x�[�^�N�3?5ڟ��n3j-�A���b]�*÷e/ h�%ۇ5��f�_���N�ߖ4p~��A+�L�<_�t��/�/������6�/����j{��M:�D!���V� ���X�n���1+�9b�4fm*i���j�r�2��3\�>>:Ҍ����{?D$�[�{�����y�^1�L��H��,͋���MͷoJ+���$ә3e����^�4g�)*�ǖ�ʴ�	�&,����߄�i�w�ik�E1iֹ��u�>8����ǔe�s"���JcK����>�urE�?�
];�Ib!�� �)�3�7��w���!�(Ժ��<�DbԕX��3�O��k�����zq���W<8�ڞ��\A_�<V���id�#/[�X�&(ț)�6���ir݆�^v����WWJ4�\��f;$/���cho��M E����N g��,�H%Q�A�n�!�TXܸ�mv~j��
P� ��*�LϿq( ���K������7@JÀ�3���+::R��~�%t�nO�#v׷�����J���y�\X����$��,TX�+�g
�@�Ѡm�T������Z��;	Y�Vy ����;A�x���\S_����E}�4��*�L�n�8�m�H �W�<1�x���~�Q:�����G�u8��#h_��FR=��(�D���)��dU��ȴׁ0���d�<&��f5{�O�~,�ߔL��\eM����_��֣T��X\���K�i>���^l��NH'O༘�7Gy��ﰀ7C�v� PY�9��@4 -�	q��xh�j b����rk*�	O�0��K�k`3�[.��A��#��l ��zU�MS�ȃ����Y���s�w���*hh��w�e�eR���-��ݫ����v!���A �&��Ah0��杉�f����r��N1����_�<im�Y$dk�=_MF���f!ih���k����~��΀ܠ��="rփ��.�ȵ��</�<S>w��X0�n�����
�~| ���\<��D�ָ��B̆��z"i���Ul��1oC��X��#�Lْ:���^�*���y���9�����P�O_4.�c���+���͟�>�o��̀eYd�xv�����R42x����҂W��%���%LR��t5j��
xC80ȅ��IW��Ť�E�C�B�r�~Ki2��T��+s	�df���}q^]H>�����}0{j�}�frO���� Qqci�p��z�)��I��n�#6J�E�w��p�J�����H�&�ɯ���5R��t�������&ի�'t�O/���|��u�G�} %M�"P&�P��~Yu̵�@��c�%j����2D>0�Nc�h�-X���Ɂ&:�o]�y�7D����s�[���"��/Nq�F�#��d��3�#���vpۧ����QW@�=;iRz�+��C��N���D;Q�7 /��t%2}�&M��!ۭ����� {�!�����f;69ޡY�HF�:��`�����E�����
F	c�'*~;zB�"�-�
�h���Z�\��=z�C �t����A�%FtaA��EօbAm!�\K<�I��$����(xw$L�v�4����70|�=���Y�(a��!o��Q�ݯj?G�m�yT���Nw�)6A�@~�n�yS���c@;а��H���~��i�CΆI���	�<�G;���WܩE�c��(b��L-��x�حUt��A�M@�݃���Ȳ�:��a��AXG�lC�m|�N俣9�r��gW���QK%�݀���MF0�y�����L��u�x\�8O�/�^2)�i���XE���eL�k9B�:�̽�Ě�?m�ޭQ�R���&��q:.=9��`�⟶d�M�ɢ���J���8�[}Ac������!Nq���X0�,�Rk� P&JS���*4��<U���S���,�8U�E�\��F��R���^5�r��΅��㸆)s��y\`���� �~gP\i��N���t�s���٢P��-^-�1`�'�M���V������M� �(���?b�[�߫B_;\�'�ٳv����.��Q?�6ް|�z��Q�q:�^@���+a�u��76e���k�:]��Z���	i��Ѹ2,�i� }�z��;X��c֥�9]����:�]��{A��r�5���}�G�X��Cy���#uRc.�l������\�]� n�x�r1��ޜ8l֘��suX�F�i��Վ4NP�eIж�G^��Q�hG:D�f��ʺ�'r�ωu�"����}J�bC{%Y�j�Įs�N
��lQ�L�'/��D����ê���`����i�� __M\E�ҩ��kd(AN�$UX��<$ֵ������h�. ?�2v@)�Xďry|4
1{�ֈ@����4vr?��vu����$ �"�'0��s�;DC�(�P43B��@�ܩ`+��+EH�\O�Ø`�T�c��q�n	؍��~�_4R}�����ۆ���q�VK�DD� ��Dm:]&?�z�]��e�z?���^�J�U��SF�+\b2��k9LS�6 �T�-Y	)�k�sG���^��I�R���Eߓt޿��+%�|���z[ș���K��Z�������W��׊�S ��mw��%�9~�ԑEEg4Z�b���b�3'�I�L0�|��?�&�7o��d�J�����ygu�����J�}�����ƌ6R�g{�y�6��%��x�l*l�[�X���*O5X�D0�t<��Ĕ�O㌕tM�Y�b�6(���8�2qs���Q��[�
� ��L+��]�uBE���Ϙ� <py�+Y���3�d���C�Y����eP$��x��>���_KL{W�¬���#�l��4Pm�p�������݊�i���	�E����M~��Ԩ�@�3+��˒�G��hE�{�C!oiZ��0�y�?�W��@p�֢{�B��+��M�2�����Ѕ޼vɣ���(�Vh�?=�W����꽘�((�-߼���1>�	�{#�m\�ʼc�g]��7ՇT��M7���E�U���?[� w�B��;w�wR���bO5��?�P�yD�ʡĔZ�z�Bw�������	�I@̏MNG�#�g�IͶft��� ��0�jn?����5hPږ ��1*�+�V��)t֋��q�&#ǝ�l�3�{�-
����uR��c�[�F��ś��?�7:�����{be�u˟�� �aY'�q�[ AN��q(۴`p��i�쿜'>xӧ˘I��n��r=V̩M���sag-�=�v7��X~-���DCRÍ�H�m?�޼��~6��^;��%h�rh ̮����u�%�]j~'��@uڥ�v��C̒�jX`�߼��*��.����A%�s-��vC��o!z��^*�f^��mV�`���G"��D�u��G뇻O��t���ǡ��=hQP��v�E5���DۯO��;��T���>� Nq�[i�\��&'.p}���)�,�VET�b�h,���{S�]-#�X�.���i�L�:�1��R�â��	E���<��(hM��F��۹��QH��h�Z�jQ���c�p�!ov<�`��΁�q�G��k��v��N�h������sl���v�Qk�3eH(����$��F�ꅏ���r@����K_�	��\P�,�|e������ɑL6j0����O-t����nS�gv�W��I����P�3�D?]F�ڦR�x&Ual���쭊�n�����2R�^qwO��%�lD����p�:-��0��o%�����灷ޣ�i�W�Q;����q*�g���NśJH�$'�)�i
~}��]6��ed���'���ny/��[��[p!2�κ %�`u�؁�<�m��][�0��|��W�
pm x�:n�c�O�r��Vg`��ӅN� VQ$T�_��#@�bdQ���9F>x�^*ۊ���b]�$
�̉�������\Emo |��q�!|�!�|%)Ď۾9�Nፘ"��P{�q����93uߥ��{�?��AoAu���Ӯ����<y��/� ýPoB�Abs�,K�QY���G���P2�{�������~}��N�Z��
�疍����<;'܊l�0w�j���N�ާ)n��.*)7�Hj�:#m=��������1������R�0��	Tֱ�}8�D�����i��P���1cX%-sաd���]�ͻ��_��'�68C�����$�2��1�,��-6?-l��$`�0�/�ofգl�D���/!Y��s�T�C��F�8���:j69�����ÁP�d�)"v�"D�.	��g\QA�,?%]�{֢g�^��۳�m
 �ߜ[-rO�bC%C`�%�����*�t��fg}S�5�d��Y��[-P{1DN��B�����[�ざ����aFW��2�yO�7r�w�ͯ6am��Mt���&d�7�zd)a4d���+gٱaK�*$���`���/�Nkt�T�6eD2\|���a��j&W�g��'539��"s�V3q����I����F�������גY�kG|G�0���CD������m��[��6�&��+O�2���$��5��3�Mq��R��R��<M
�X��#_�O;f�Z�u9(,��=~��TT�m�S�<�޸��T'P�u���P�^��ߠ$I�ְ��٪�����xv��$������~ 1�%�Z�dM��C^[�	�>@�A�ױV�A�V�/Ef�,���Uc!"�-i�������z{K|�A*�	�BH͉Yxۂ�c߯�"����&�c�a.�ZZ�!K%E; ��� h4�����5b��8��x�r��-�z�iX���l6G���0��z9i�)61��mN=�;���*���T=@�	{�� �z�A%����M�$�Zf�ڮ�5��H��B�����e�:���+]<�6t��P�<4B�W�����#��RG���'���SA��p��9���vQuA �����]�ZH�e8#	�Ht��jh(���=���+����|MM�CBx.�^G�1�vi<x�iH7� }Fv��K��)���.�S:��{�j3GG�cl����F�
.�s�e��NAX�z(V	H�/�dZ
�2qRX�:p�E�o*
`��p���z� r}9�蔲���MN�����$͊u�E#��I$�� 
R��ь��kMN�zT����v!�o6V��N��l}�8c��	��q��Q(�Y������f`ㅸ@�EPg�D����隣��_N-��Vޗ���������F�2��<��F?�s*�J��A@��sꚐ����щ<������j��ЭT�&�ejA�v&�4���P���;ӿ��i>thl�Gc�A��D������u�!�W�7-�GY]�|��ք�?2~�����4g�a.)�G��h:�r�QF��C��" &�u��S�Ĺ�ѩ�M΍E���?���̀�Դ��l��9�p�K�+D����d�"�9��`>�B�E����l�͹5$��A,�%�`Q:;-a�֖��Mn�7���W��'>q�C_[G��]�Q�����N��Ԕ*�������ǠqkX��]"%!�?�y�ݻ�����$|̮�B�sy��Ɵ�Xm�1}f������NK�$;W<5�6�[-�V$s6���N0۠4K���G���}�x9�z�E���z<��e��+�`��i�R���u�X�ΤΈ�1!_%�Hv�<z�Io8`���e��������Y�F�*���/ y�e�PU�L�C"���:�T�?8�*�������Ф�l���

�,���<+�	O�WC[ۮ|�FI�+Ǫ�E�;�?sqю�Uo/�>�|��zLڷ�K��[(��rY�c����yJ��fR���DA~�Y4���J��V����ن�$�����m+9�R:�1�~��)�l�9����gmM�4�)��1Բ���V1!���-����ǚ{ӄ�iό�}X+J^��0p���:W3E>z�d&,�D����ӿ|TЇoa��%���B�R7���;.�tJ���5��f�X��e�w�k����/��E�ɣ��˷[Jڊen���\�
�K��|e>HW4�����W�h��[>?�Ģ�n� G� ��>��?3�����"+½��&yJ�tx�:��~�=��2�vF�q%G����\b�B�t����%]��u��W�tx�с�a&]��ہcG��1����s'r�)C��*�#a��9aj�O��6�)���
�C�����=��E�hF.�^��(��PѿY��X\s
ۜ�ݑ��E$P�ԗ��w���۰$��֏������hYBiH A�S����þ�p����з�#�}��ҥ9�tq~ULdFZ�����f��]��p2wW9̃���&*J���BJ����.���	���GO�� .���v�$I�'�@��"�Ky�b($<'L^F]$��M�?O|',�D�̆;؃̬�ek)=VKq+�m%.��nX^ �cN��4eKԁ�N�����#�c���ƚN�Fug�}�{� �wt�.4Sui��=�U��x�o�g
�@:0Lm��9�{�m���֒�o� Cl6��j��}-L}�]@e�k�9�����n�K%�x�[�t~���S6A�r��3�`b̞�u+������b���p|��9;�����,J
���M�h�s�`����p�'����+�fg��j���"�=�		8,g�D��K24�6�צ/H�J���ŘZw0�-�%�p̠��ʋ���S���h#��%j�+z�MbQ>g"���rf��(��[0 ]���i��<1-�����y^ �h=�M�2!<�@�黀������x��B��wM\��0u�7X���2���QY�[ա�6�:��G	H����'+O�jfԨ$���Dla��v=���SLv��ƥ �*�	�rjZ1�n����U��U_`��"��x��h��g?�ϟ	ev^���``��t����`�/+ܬ%N*��Q]�� �}x�}�T��+�N�
��U���$4����{�|I����@Ὺ��5����r��l�����~QL��MP�`ud��0�䱴}wo�����>*��u}h�-���?�>��W�W{,Rk��.;J9�|	3�.M�X�.O��O�_�?��_Y7�E�#Bn�/N��q�ewJ%{��G�f�L�y�hc
kmRj���{b���%�㯢L�����
���B4R���z�����M�c��4�q#w�p�!�����嫊,��j�K�":��y���f��T�i�t��&��f�(��/m�n���FvDjW!I����s�;`��ʮ�����L+M@y Q+�d�f]�q��:�e�?�e���%�w6L�� Xu+�u&bg����K���Ʊ���|��C�
N`��(
��O�H��9K|6t��9C���;������S���u����)�Eq[�N�����-���a9j5�E���;�Q�ĕ-��ۈ�����a���U-e�52Z���p�����<�N�F��C�s�5C%�< ɵ��K*1��A,�W?�&�i0Z���ڄ.��OOu�2kiOܧ���s��ؑو�_�v!�s���q�����nWL���,$�އ�̜$>("�oxO�E���]	�I�l1SA��F����ie��9���9���1��Us��jl��x9oz��P�2Z�Iv�^X����#g���+��;��J�:zN}_>f$ ����c���ů�}�T�X��.�@4[I~F��?Nn+����H����h�.c�;UX���pEd��J�S(X�� �["Z]�V-�n(���p�P-0����\V�!ؕ��V�M�S����a0��C"4��FgY�ίs��/��N�.��2Y~�G�&SL�f�{��{�aPDE�տV��=o����I��7}�����yzOssކ���D�P?�,w�)QL���GL���k�?}�&Sj���x�k+�k�;��g�NG'��5��V�c	�J��pO��;���Y�#�>���S�k~�N��6.�7��РO������Z�bW6R��]n.G%N����%�ws����~P˫G�ʶ؆.����~���C �e����]V����ڸ�1��Ot�����ͩtI�)4��)�LΧT�hL��BY�f�`�i�ǧ^c�*[�}�3�W*0����}�9�.z+u��M�GD��:��:�KT���-�sWl�A�[Fmď��[����=����T9X��}F�<c��M��zq���m�ҴKK(а�M�P7O�#���kU�h�/\?x�F����¢̀���`5�u��#��cb����Tg�'�)#d�|B�{`�"(�~��M=�::��Nݵ����%$��R�E����/"}��Y�q[��+���iW����
���o�>��9K�ur���0�6�(�Iu1�����?Ò�Q��#� &�UL+�N��������qI���m��̵�S��<�ch�]�rl��9��M�Ю$P��U�ؾ%�(``�z�@UB]�O��E���⛭�1�Y�����-�3�L�~b�G�0��D���-��=�7�ha�.����_��5�������~��#Й��*��m]m����i�N��)$�/��⁕�@�k{e��I�[�B(j������v}���8�"�$�9�ow��Y"%�**��~�cK���\W2x��q�ik����N��ڡ�?�Ś��"`�X���H�(�:8|��Q��Ga�X�޹��YI{O����Ġ���"@����'/q�l��տ�H��2��E�.��fD}P�G�#���(C;}��e�4�!	U\;t���bz�>���L��6LV��|���'�pX=��� Ǜ��-]5������]�`6����L���)��� 6������L�έd��2 >	��CTԪ¬�ϊ��vߙ�Z
ww&=j��%����(�x��i�>�^++Ci��M+���,D~ F���k�\GD[��E47����8i�X튑�#y}[�\ŋA
B�(:�.�y����Ȭ� �K	9ϏI� ��YҨ+���o�@�b�gQ4��,`��;æ�y2�\�DY�R���c�[�����7^SD�2���e�1����;T6��Emv�r�Ff�]�)�2�D����V|\�2)�0���h�%�$?��jI�9�l�$g��o�yńY���'8�+����,�����6s�)�X���@Zy��f3�Rd�3Hp�d������r/	#2E���.�I��_�z�E'�E�9��ct����j���9��g6}�ǗXKR�t�d�}��إ��(�j��7+1n��'�Pyf*�Mk�U��)V/
ק���#�����kn�r�-;P��o��;�{�W�kx� �Ģ�!O��Y�+'�F菂$�N �!�T?���=��#��;��3$�N�Nwn��Q��푅�����#�O{�m�;*9�M,{�Id�Q�B���>l����/y
�:3L��f��kE��'��480��Q7�l�� �Ӑ~e�WH�KƷ#A0��W��a׈eQ��	c��|˄�m����xFN�ݕF�~�
�+1lrFH�h�����#�G�3R��z�7��-���v+�������+�%�/I'NC-��y]f�%��'~cB���ِ�m�@��B����/�k��-�Z��r�lg6�f�?���|��䓠K��PM�
���bt��A��tq�%Z}/�=�	�ɢ4FEhVr���:��F�PR��-M^��w������ʦ�"h�N-��a�E�rv4{N� J�~^�9N�sf�*qP*�����R�w�E��O��ѿD��k��޽�c&��l����k�qg�
���Ppm�g�9�v?��xi�1}j`����֊(���]��w�+C�qv���EV)��5M)��7)ø��?[fP��"%{���ܴ�
[�z8ؾ�T�MK�e0�i]�Y� ��oL�*�'��CF��rQ�/���ۓ�P*���i��K��;T1��A�uȕ�Y; 9`}:�ӛV���%���~P3:�G����G��"����+qԘrn��r�v��{��znF��ᰂҐ |t�|;�AmK�����&�*��dy:mD�ˤK,Z{���S��l3���!���D���-�~^�H�C1\`ݗr1�|�
<���qZѮ_r>�ie7�v�hq�y�<G��%B����m�nk�-�I��Z���$�s���R F�ͶW��A��ADA��C��������Ϫ��FN^���`����>c�����txs��V=����z!71巌~7'�]C�-}���t�bZo�rP�����T3-���HJ�I>Ejj�Ӯ���M~!a�D�Ce�}�?�?��l�ԭ�M��>���:��C���M>`TEL���rN�6#�R�P	rq�>5^mA;�x`�.�<X&f�
$�HJ3 �h�Iy�:�	�/�Y���T�7ʾ��i� ���=�WkH��G�[��lq����`o3M��֩����z��[pr�@�2hFr�^c�ZZ�ѩ��*6l�=�'4z�
�3.����f�����L��Q���W���]��):)k���`f��̀b���e&���O��*������������y���E��A �|Iaj��僆 !��w�a:��(&re����j��N�������?/F���6W���
q=����|�j^ ůt�t$���bh�P0xz����Y)��L��ߝ��hi�sq�u-8C�Ytk���1�-��	I*��T��S��1g1QR9��4��E�w���:`��Б�9�+_n |�չ���8�L��|����d��s}Ŝ��"xa�jEJ�i~���ϺΊGG$G+n��/φ
;��N��͎F8��b��C���/�Z	`
o��O�}�)F���1�k-�/Ze4�!m�O��������e�"봐BZ�1��T�lg���-,h�E/=\.A��` ��?Z���ީك~0�(��� ͜S��	@��UR��A��m�7�3s�s.M���@�]��Ͷ��u2Ҟ����Z�Df�m?
Lm���^��H
#[r�{�B����� �G�����=M�C9A�-�U�3z��gX�.YϺ�Ǜ{��h�����[Lj)�8��`�=�|z�aaX����
��E&��3���G�)<Ui�$��UiR��*��`���%��!L]o�:���A�\j�t� �Vb�cV֥z$u+������6*�G�X�8��MMjr�F���4E�V�������ZF3�$���0��rG�#r��w(�z_�yR�·j����1~����k��R�j޻� ŷR\��Y6e- �3�CZ����D5��|Ѵ�g�ˮ��##��ሠ�����w-:]��_h���- r��!G�<h��h�i3.�z;�N:�����~�ңd�d��솯Vm�c�т���!	��8!�>���&fa| za�ƔɌ��(��������;�2�	T�J6���`��*u��)�H��������RT�Ԁ}cV;�}���W2S�������<c��;��ϴV�(�&�]U�h>�� �R{1�R�v���%t�Ʌ�H¤�`�pU��4;��F��%o�T�ܮaq���nj{�&�"̸���՝h�,m0�V^����4ē��Y�;��N��WB�6n(v�U' ���n%��Ӷs�Ur�Kc�nU4�g�(�pݵ�h����ƎN2�D��?w�	������f�]Y0�G���e�����W��I�{�ѡ�c�s�Fx	��P�d� 䩈GܼV
���s����/��R�F ����d�Z�gb������K#���_�ٶ�����O����S�_x���@Vh�E�}��I�,OMr������l��0X����P\Z�&���2�.D��R���q��'�=�=W�o���љ0���R?v(�7G�}�C�/6ɧ�ؾܖva�P�m��2-aإǓ��)� �E`�^6��=����)�v1�l��cbi�Z�$�!�nIOݨ�E�դ^y'��M��6�5!�O{��dn�Y��/"Ww��ۈ���%��cփ�w�'⭖g.�D��x�2��HF��ϋ�Ⱦ��N�s�<�1ț�L/q(�L"�|��J\�Z
n�'�$�V��}�V�b���]�����$�5�m��@�So|����-�ļS�K�m�����4���b����x"ţ���*Iԕ���1*Z�D�%7H�p��a��;����Vo=���`�����>|�gYa�x��o����0'<ـ>�X�r�m�)�Ƙ��>P��Ǜη�`�φ��%?����ѡ����i��.��N���V�6{�Q�$;��ԛ[�����0+M�G��?�����b��l]�Q^ϱ�l}��"\Ά�X�ܓaE�~�5ҧ��D����?���^ec���3l�8ɒ��,@
=�'��j)I
w.�<��븅�I]���d���*��"�?���p��������C�P�$TBB,� ̨�2ܽI�I����չ������m,��jPpmS64��V�Rac�(f��'��T����
����~��/3$�`~!!�{/�1Lg-��1�9�"z���:2�n݆F]c�g5�n�XBC���au/caE@3Rԩ-�>%2_�w�:�l�[o��yaJ����� a
�0>z�޾�]tq˪V��,Yd�bav��Qѻ�t|�)�w׃���ݜ��c(�2~���y�R�.��V����s0�Ш4;��v��ৰ�y������wuN,���%_�@u����x���ze/��B�/{]�ޕg�.`)�R��;)/E���|{�y��7�"�B}IB�aD	���q0�+��D��_�,�����a��q�zz>���ЄC���๴��G�X0��^�]5b��>��LNw����7��l5pص��]��)�ɧb;`��Qѣ�5��;]M���J���ش{�ft�2��sͫ-��X<1KDͻ ����ң������]�5<G��(vu�1�a��24�y��*��S?k���D�%��Q���%{O����g�(��^�FyA{��
��,�Y'E���C5�M��"�my*d���Hx�'(�▌�0v� bt�G�Ċ�pꏔ�~&
�x��q�ބ�`�j�������/y�0^8*�e���ғ����MN��g]p� ��g�H�<sC�}CJZ[p�_>�Io� lb�7����ߖ�ҽc�'�ߥ��	�~* l��
�`�|,������G��!�ZG;,��C�3�X�/�5�i�9�qr��l9��1���ڑJ,_Z��caMTH�̈́��)�(�C� �i���Z�?b���e]�Y,e���4���y���D�m�L)
�nM��1I�:�����:İ&"6�ƒ�Q|�c(��zZ����X/?)�v�~��d�\�V��-D'_3����V.R[%<*����|h�Co�v-�`�)�A׾�crbP�\�l�.�F4XP��,N T��� <��:�wJj���F2F�MS�����G�x����l��h�dŹ�C�Hv ?�O}OU�,LR2�,!W��&�p�R����ݲ16M�f��V�؀t�V+؁	�(�;X^q�>γ�{�(nҐO�ig�"��VI�[�ϫ�&i#�I9�c�_�|Jk�J��߲z����LsHt-�����<�.���<����8��֥Sz����7<y)��ۜ����ٗޖ���w�wL��	,՛�U�F�&����H׊:�S�Qx�5ڜG9��6������H�l@�F�(԰���ʻS[��5k�8�D�͞A6�e�m���i�^`G]��V��6SX��Gu��Og2�$�>�|�zxWO���o\�Mh��yV&BQJaz~����Vߓ�O�r�-��wjCj�
�@O��bg�o��-�T�z�R�
'JGt��0�ai ;~΋X �LIĲm��\�����0ה'$(!�p�\FC��c����w�����NǴ�s�P�w�#��b���`T}$�>�-],˛,�.#%6_[�hR[���.�&����	� e7�py�R! ��KQ�{�o8�T��I�<��1�
�1�MP����皱�/���#ݸ$' @2�D�y���mv����=�9u��g�F~�YBTD=��AY{��U�zn�i���̐�vqo	;^�7|s��Q#���+����γ������,ҴYǣ���ϩ,����j�YVك�����#Y���ئiaT�&E��k��ۣפ�vg�}�`k`-,v�z̼�m��[�,�أT��� ��� �P���W��t8�.e���{����i�T4�W��ٶ�7nl�}�� �@��R��w�LK8c������GA��t��b�|����ȝN���:�]|>��-~����W�P���$_k'(bv,`�avC@�z���c��T����:E,�f�b�Zw.`>ƙ�mphe|����(E���[{�VYS�4x���Is��3|���2�_�2	X�� ����Va�u�<A���LJ����Y��Y*��W�-k��΍���hD���
���^�>�q^�b�]9V�I�^(|�
Ӆ&�m�3s�����]�lhI��CĞ.�V����ZT���rb�x���6�魹tC�s�È9��3y���)�i�7[d89[��{���xm����oӳ�B��#7��qr��S�Iy�O�Ʀq�岮��xFDC����x�j8d��{���$;�JN�h�\�Ky���v��q���)u�|��hMOY��t��9��rF�cp#�LKy��?T���؍�,�e���EKK@l�[���s��=����[M&�}��~�)� .���G��4�EXm'%�T���vh��#E�6	�B��V���^;���4�oJJ��B��V�b7:<a׾i�������nR
V��Y�P�+���us��˄�M(�ܹ�����&g��J�ma6<Q����d��d��V�~�$ �$����  �;I�}r�rP�5X����Վp�aPh��� �� ���W�`�`� �ބ��������$	%c��ݤ�<ʧ.y����wcL޽����(�9p�v�1�r'�;�Q��(]�����c�*;:d�\Xl�}�J^���q�wa��Ĝ��@�s�6Q��x�>�bxY\��j7�OUW3�Ja�5�O.�C�k�8Z��FtG��:T���'���XT���w}�@Ps��.�y��
�k�.���B̳d��e����h~Ƒ�N�ZiG�y�B�7pʙ}"�HiZ���,5s*�3��М*X �b
�k*������p��ɹohv)���o4k]��=Ń���`�ԙ���3ˍӨ�%��m�g�;�ך�?�H�2�C^�%T���o�SՑ�/�Jjl雖�zq��{�����5Qd|ز� �J�}����P��s�5��$0P��>���b�Nlm��n����Ӥ��Z�x<�l�)��Ek@�%#�����yc�x��E��rn����$���ϰ��ϐ=w�BT
�����?�;-D�|�X���Ly�4I�TQ���C^`���QG
�)���T�|/!��ZO��u�7Y�}՝��spoL�b�k�}�5+\Z��{gmas
w��ݸ)
1���@[�5az}����C��w�W�`ȅ-ke C����r���=ژ�cgz�ψ�`���p��~N��U,ܖ�R�)vس��9��T�7���B什?`��r����4p2�1E3�gt�p�?�����A�Hvx�����Q��[� �s�[��y�N��s%��^�4�G����V�h���-��f��uwz���Yg�:)�V%�$����z��
�=��ڱCʌ��~/�g=kh�k�>j0s���T��K�ZO#��'�9�\J��!J��fz� ьG_@�x�i��1��ڰ�RYz�*�!`Z��
�W]��(��\&�t��1�+T���?�,����8��,R<���ŝ]������|Y@s������gb�?�w%_����^���Ws�f�	a�r�����PaX3�Q��X[g�C�޲d��B��eGçl�Q�4垤�Ԣku(�B2e,���DC[ �2{�k��I�:AKw
~���~�|�k��i�X��״&򠴽l.mJL�#d�!d�t�X��������A���Y���;����H\2.��r���'��R}�p'<��~�|�g�X�y�H%�S����Y�g2�g�Nރ��;{�vT�!��c|x ��m��V]�` �t	}L��'>&��j>H�7}ص������M
J�5������e��^v�jTM˹��Q:�Y��dl�ޕ�ɻ)�*FD�m����,�(٢�/a����Ս�V�7�|��hW��Kto��&L��k��
�-rlv!Yr�t<v��q��c�yڛ ~�[�VW�](�H,�&|�1zGm$�f=B�����j����%c�~��S+�g�Zvɵ�0�1o#�@����,#�/ʘ�m��zW�+P�G�/n�dF���V\\,ؾ�?9z�Һ���� u<����):؃n��T�J��C��}g����P�d��!�ū��r�+� l���ԦV1<�ِ�r#�������78��X\�i?��HD��"7f@�ҩrӭ�q����ዊ4��u��n��s��3� ��I�Ζ�K�>�_ܗ@��|}�����ԋJ|���r�gz�p��(U_KwM��;*D���L;J�7��M���m)���D^M\�� h���ܥeJ�bu�r5T� �2�
c���]f�h����ǆ.5�T�"��$��W��l�7��Ma���Ӥ�ޝ�E7\�S�������[�4���:�7u����� Xې.�JNw�J dx��D7�0�Xx?��!�W�nE���N��/. ��ƲZ� ɷ�0���#����^/���v{%Kv]$�NP��ןO|q@e��c��
3Yp�޽�n�͘Tz@j
b�]u��@�]#�d�����p���ª��B�n�Ap�~�Z�O��UH��/��R����v�ښL�<6K��T���2�%��z?�l�����@ۯΌ�o���EXL�~��!��争�,�It�i���Hlo�dܤ�xZ�%@������#��L_�nYd�bWD��dO��Ҍqܕ��+(Q�5�R�%]��aП>�q�gc��o+ʯ&�_ӽa���b��쒾l��[��Ue������v)����m�Zl����`>	O�s]���r�n��|2(Al�/�y��������9dB��ۜۧ ��U�gm{&�R��ʕLȭSk�5��4��0˽�,?�v�5w�[k\�/r��	�{���-�O�!���U"O��ko��C£q*�$�O��������7�
Ğѯ|���)��T�>u\O��ݕ��� ��~�#ѯ���+f��X�-#���yQ��Kי�S�����iiR��#��f�,�=UZ�G��
�*������� P�R>_+������3�?B^���A����^\/�ٙF�N��������3&�����,�*��϶@�� j6O����F�ycS�C��ި����!���A��)R3�rn�f�Ҟ��+%]����:�x�7�0n}x!�kݽ�B�pJ��}ɴ�W����Z������6�"ANWe�}��K�7*8	?��d,�z�#~5d���OJ:�� ?�a��U�?��D�@���Z�<�,/1�rp�G���ˊ��t� k�"b^�=�4m�\E-1?�AP�u&�s��]�.�;\��/M(�O(�d�α{q[�D�<`1x��vdy�q�@C��
0|8V{	�N��5�\=1]�2?��ìN�2�h1�����p����b���A�ܡ��M� ���
a�\5w�V��6hNd*{i��+�y��KhN�A�1�[1�S��: !�7��z+=w ��?�}0�{Eh+�^����ȑ/|7w��� ^��!����+��nq�K�KeN̢[Ώ�.�|��ʖ�-�q�2����=�Ay�O`��Y�Xi�܌D�{�v�b�ᤕ2�+��$��/�����$���4���Q�4����٪�7NyW4�x�t�L㗆�D5}�qA�|=��Z�Z���k[��
�r4��i�SP�a�h�s����&S�����β��$y!7&������C(έ�Bw�,���-�aX��0^�2�?/w��x�O�WF�ET��.����~�j�R
���}iW�W�-���]|��:�Z��K����/�h��yr[u���Ys��3�U�S����N����NK��:�{۹�"|�|�R_�c^��b�_������6�7i4�F6{���U~�0�7qS����4�ٷJ�(�7���"{?���5�KYМ`Zbs�J޼�����7�3�(�g�H�Q�@���sY)؍����k��� Ѫ�,����iW�:�����k"��q��>ȝ�y���(�t�H��S�D$þ+�S��Cں�F g���Ա�#V����o����yЯ���$Ãu f�x�ak�W�7*a@��\~ϙ6��ŀ���kO	�^��C��<����d�}g�ݺ{_���a�ȳe�C�3T���ڔ�)a�zI玴bݎjDu_X���	�=sfRtдѬ�Ka���}!(u��=6�ѝ~�P��
�K�A�F�-�QC�Jf6w3r��td�h�睧�z� wu-���ָ>0>�G�+�8��m5���|���]�����$��1Jy��J�1Zx�"H���'��z��S�=d����Sihu .O�/y��I��'����/�ٜO}&.?����-�O���__�F�@��w(�1�֎V�v���z>�(��=z�S1��&��R�q�PW�9�}5-��Wl(�� �{���gjƃ��	K�Y�6jD��[����p��5�
�.���8�\�9��y)�L%Nt����U�K��c���=ٛ���dH$d��4�M��tI�������jϫmj������{^�j�Rk^O@8|�L�W�Q>�V�|�%D#z���i1R�k��E��Ng��A���&���������Z�?2��2:ձbw<����VGz�L碣���Y�n~� a!M�55��a˚&�00V�VL���rJ�܈d�̥D�ش>����k"^�����_�q%{�_Z�P��OF���wH��b����z,��Xq,MasU
�����idN�Bq�G��J��t$��nn��a�.9k+�X[f����'��h�<=�o��뒈��J��Gh��s��`4�G
��l��{6R��x8Jd����U�0�b�|�u=�V7�`�8� Ҽ���8|�.��LV��u�����y�PR[��Y1d���x\(!�C��,5�Ծ[g���B�%Z����<UI�8 oH��)��p�9�u��� Q�q���\i�x����l�����ܸ�_h�ú7XL-��~�x�Yp2�HX^[w��u���Dn}W,�21�g�����s<2A dR�N䐃�����;��L�O�dF�ω��x��(�7��X��D�H˜���R�Φ������C%+������
�]8"
�r�3N�W�(�־�D��˳��A�a/�����n�ơ~N�/�L��
��x����D�k��SX�#��/Ǒr|������dglc��k��y���zL�c��`LT#R�es�Z2��Su�@ �*�Q�Zcd�����+$�y��N%X��v���L�aRm�a`"�8>���.��P{_�#j��:ԤS7�MXV��^�!�{(�� ��o���~��J5�G:V��%@� �a.9G�8�'<.���(9�Z�X������t�!��m�H؜��WW��yE��S�}���&��K�Hᠪ���oo�,�s�a�ojo��0����m��ݭ�f������d����VX�NG�G��cP��CaTP�x�����ByT�O1^R����$X�O��x	I��H�($�k��h��=i����E�B�C����Rб���Ĵ�CІiC{����m߀+#
਺��@���7d��]��G�1oc-u^�ED�>;���	0Ш����Uٳ�	�Ǥeo��}�Ӿ��`.xu+�4��B�:�%˃�� �÷�!�o �!��Q�iE��`
l��3h0-S�!E�&���d�o��/,5Tl���*k��t�q���{{����l�w��i�[=44��(� \9W@Z� <o����]����W��?eh���6��"��]�Sg�*�~���߃�⦛�K�V�����(��8
��ۼ�N���wڂ����8YO�<S+�>j�̱�'F<<�}ڎJ�U����cMB(K���1��I����_����D-���6�ծB��d�e�<���EZ�ޓW��I�Is4����c�ԇ�hÌlf�Y�,�Q�g��ùQч��PYwtޘ:�0��U��<u8��`/,V�V1U4��imi�=s�1�@h}�"@��Fg�sj�<�� שH�]��?�q66����jT!� %�ܛ�ퟺ�o�U��Y��I���5�E��1��dH")���X�x��t�DF���:��Oq=�6 �=\/w���]E�]np�K�Mu=j�(�t[ʣD3�\w�(T�I/��{��p�r�ɉGvt�l��r͛�y������pѱ.��8�8-�m˚��� _/�71��9�L�Q��1r<��+YH�Ǆ�h��9yz0T�e0�|�6�A?�;C	�%���\{;H�:���(����ȕ���{_�������7�I��<��f�a5�;��ǰ������;,�(�?�vox�4t���/�u:$O�s�������~� 97�N��)��*z#��e��˴����G�v��M��"���}2�P�W�[��]=ěF�b�(/@��u�v9Z���违��מjE/}5Sf|��o3�>b��	�^� ��]�"���6�8����_}E���:l�0���eRb'ڪ/�ߗ�p�ʰ�#�5�h!+}��q�$��0�^� ��7{�S �E+�|
�2��g�ќ��wb���u ����40�%� ��/
�P%<C&��e�g0�-�2~럈�3����a�W�'�_i����|M�f��ulD7I��^���!um�?zj�V���g`�TGQ�z@��87�*,�~^�&�޷������<o�Or6$���s��}�w��ɀH���Ĕܿ�iCcry	_	�՚�h l���R�����'u)���B�}�U9}@��f�;xH�X�~����+�Ԡ��m�I��Xv66so��~��,@)�����af�Z��A�=���P���{lgq'���uD���Ρ��[W��
���~jS��{�u8Igly F&��\m���b�rm�Ղi3�$�05��B����'������C[�E�OK6q��Tfzq=�B��)Z�i���.~?���<��A��1y�XMZrDM�mAl��og��Fn�hK��D���U�IfT�8�*V�I�ކZ�H�?�ғ ���'aA�#Ϥ߷�ܓ��V ��Ǌe�HNb�"Г�c���+�\>?')XS٪G���m)G�}�{������+n*�e��P�DAxR�J�P���X�"M3�~~��U�6��!��s���r�6���)�F���/Wr��L�!�3�噶X�)�2bDg�h����䍊O�����,��]��{�������Qa�~;�r�63�ب3�(`�7
c��V���j��th��߇W��~
���������3Fׇ~����?��M�-f��,/���b�P�����^G��W.?�"���������&�'-�ĊP��ۨ��j�@HN:F�&}6���H�|�� 𚞥y��v��#̎A�?m7����EXl��	�l�����u8���OlU'��ʋ�� ��i/�H�tLզ��%DR���t"�;��:VP�x��|A�P�i�o/"`�SsO��4Z]Z�\Vm�A����v^�B381��`��l�#�Gi	��_P?ˣ\@�'�}�˫Z�.c۞,ZI2=�,jL�N	�#i�d��B��Ď�՜�ja��#�4��w�`�;��x�=�4eAR�}h.���G��Vw�����d���8���/�S�J�@��nPm7��u���FBA2ǽ?��P�N��p#�l�]���"Dt�imL��43~V�H�?����*񫻱?O�7����<��Sʝ��Տ���w�y��K4�C�����~a�ai��/��	�D��κ�X�|IU���z���ڑ��M6�l)�9����3��3%��,+k�f�jd�}�NhLA�6!�+eʰ���]�LD9��{�Ma1��yz������9c�Ę3ʺ#^�N�H����Ÿ��f�^~D#�&:|�+��U\�d�=@�	�Y��LM��W_��zj�l�1�0��H�Q�U�A�)P�	ƾR֓`�v�����)c!l\2���N=y�w�g�]>q�$