��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�Y֢�08)�	�SX�����~-a)�M������Fn�[O���� �B�!����Kn����PKāG����VYP2�E��,��D=xx�p�F=�Ӽ�>����@O�g;��C.΅"����w�����4-6o���6��'��	���B���;E�L�_q�0��^��P ���ܬ�n��iX��(Pc�UBK��L�m?���W
�w�/��q�3���Ub���ЕN����c�aCQ��@�4�!n�: ���DP��m����3ߍ����h�C�����H�ZdD�nӽ�\A�&I��h~g�����7w:�<ٹ�7��t<�](�	���XC($mf+? ׈SQ�@����]���h�R
�KQ����(Ȏ���7�h�(`ƪ{�˚[0����5#]�?�;-%�U���	a1���JѸ�x�u���A�����-N�ެ�ʅI@4N\�9tD�S���1a7�ˉWq`�5m���]�n���~�W���#G�R`���9�}Z��<�ϐ�s�?�ɳer��8����G��
a��v4c�P#�:��>��j��>�˶7x˾:��c�����A�z������˓�O0���KHk��u����l-�S�4$��wE�����D�3쭐�����@O>Y���A(x�D�`N3��� KĊ	sԤdp�cfT.=���Q�S"nlu��޻�A%��2i;�?iM�hKÍ�C�џ"��̫X�1�UG��>���q�Nh�[���Ҽ��7Y�X�_�5�'���ɢ[�����c�~5�ë$o�I���.�9�t���hW���.�?��^_Xu�|��x��+��h=���؃[؁�D���|�Q�\��>@�к_gی�?59��@��_{�>.V����&K��� lM8��b�=A�D!'L�uB���~��T�A:#I۵�+�g�'��\h	�m�]Ƚ��<�/�2rLZ��9w�7�\%}5�pl�� ���E>����-����k�3?���k=�S�Y����k+���t�m��07T�U�b���fڰ?�l��y_�� q���̉�P�3�`�fĳi��������,zx�ζ�j�i9CS&�Ds�����	o<�+�o+������I���4�3u���-���oZ^������� 0�jl#�%�z9'BI����H�a�I�R���o�z3�O��9Ǟ�r@(���D��@H��Sg!��.G+h��q�J��<���9v��?O�(�V�j��t�p���/�ȦH��BQ�&S-�Y8��U��SPAT�L�j#�����hnYo*UT�`RJ�RA�ƀ[]`�0��V�<[ҟ^�ק����������럠캩�"I.d��I`��>�~��?�Ʊ�2��ޥ�r��R���ޱ�~�
O�η��)�U���]9@�ӆ��FT��g�I��*+4��{�6��Dx\mB\������4w���(v�������w˖4m���`{���oᵉ�gG��j�~�[�H��^�J�,C~�Ow��jr�kQ�k-��������l�#����}L��y�$Z�(4q���v�ֲ�n�M̰3H5lжp�zx�'9zz*?�	R��fȋ�Yva1׭�t�c��DF�:{��e���v�7ij�fõr��6U��N1E���/�;R�h�ī�V�3�U�G����r��V#�O��Oz��"�9�%b���CM���mҋ�u��%4��f|D6s�����T:��8_df��p�6�yh��U>��SF8d*޲�R��!tҏ��Z�T�{Z��V��=���>��5`�|�^%�K�u�Vao�,r�4g"�z�mvlUZ�빚�Bn�1��Gҩ��w*ܱgrL~�4 Bۀ"V�%�����U��f���K��x=(��פUt��W���T$�k���͵���ј_��_l����d�i�f�Z=ܧ.YI8�Vݧұ��@�G�ȫ5l��x�M�X�d��+m�#���gP�`�� ��C� ���yC��IS]Z&嬭�3R�����5i� b��hVǴ1:.��^���Y�T�z4@+h	u&D?F_��E0���3��9��#���7�R�B�?�wݻ
䀴�m	��<X��F��%m&r���NJ�e���\Լ_���S�r��];��)��d��;�N��'���P&�N@['G_!I=E��m6�x<<� T$:�]Q~6��N$*�����ǀC>�۠�jUɧ,95H7��5��NTZ�B����)/�\��s	cǶ��/,L�m�K�0U���PW���u杩�z]૬�$���rt�d-�@��Ij���X��@�HW{��O���ߟ�3��d_A_,�]�j�OCu���W㞘CSy�n�� $�ٝ��]Ei𪹺��Q�CB��> ��A��e�d"��q�9NhR.c߻�[98�h�w�,7S��P3@ݳ����i�l.`�Dï���kN��~�q�c؝E���Ɇ��0q�eΒ�M���lﾢR��y�0���g�:䄇�A�y�0+���OKl� H����+-��ǚ+5�JȖK�h����ϓ��A�d1�	���P����ȖϾ�0��V�I销*!�Jw]9����AjmLgch����M[���^~ ؊� R�|�G����H�#�__�^g�.E�rIRTa�+�H?��5����W"���o���GZ����ٟ[�{+��vv�*I�	��(�i�-	xD����e��_�M+b�(�׿���4��T�G�#=Vۑxی�_����$c��A���R��J�9��v�p!��^l��i!*`h�Cy�����#i��+L�ុ�tѢ�
�8+�|ߝ����X<\x�b�	ܾ ��B���3��?���;�� �㎵�TÑgE^ĺ���z�%��}��0�V_����G3̆P�1����)�#�$2]6[6�K�vS]�X�����G�M����L]�GvZ�CNr\Z��[���Ǆ� �1B��?;���ĉ-����R��t�L�ȸ.��A-��~1��~a]���'��գw\������%�0���̈�j��G�6!+�'�\i.q��J֌��H�|���M��m)���Yj��*)Դ���Q��=����t�׈8!�5������9�u	R��@�Kn7�,��z�J��M����dh`�Z��X�fH��P\�y��O	��R�x ��S���	��B�#�����������a��9�%�'�4��؂�m�pl���e��g�����qt��,���0Ȼ�E�M2���0"N��.>I�M(���w��5���1Y)���w�*Y�4�K���X�I8x����%k�:���5�3(ȩ�@�RAɧ�97�����
��K�/T܎��]/��i��CQ���V��{$j��ݕ���/���7�m��F�����BU�U��HC��ڹ00�
��n�ƜQ�)��ǚu���!�������\~�]��{��U-fn��%+_��2ua�eJ1ah��r��,���N󛶜���Xi����[�Dd 		�������6r���=�E�D�7�,�~�����T�{�$�mz:)��!1j'Hk�5=���,��6���Ie(�@�ɍ[٠,����۟��2Qw���T��s]�Jq��&�
.�*�+{q���%�����J��I�Nn�nzH�Ph�+��t��^u^�\qm�>W�d��z���RMg≑���@G�t[���R>cpE������7Pi��ŝ4��Є~ 6eR�)m��滛��bF�tu����Bi��γ }i�<-E��2���ɦ}(��%KP�&k����xb�?�d���p��܉�����o�q&�Y5�x��	xЈ����o�Έ�r&�DkG���.����K�Fd]��c�vEB���0�7��$U�_�1�/OFT�/����Jh��Q2�Ը�#n7Z��/����<�@�lm�sM��s?ITD$��`��x�x1�#%�No�rHJ>oJ6�{��*�L#�o���5n}1Ƅ���Pla�rG�=1!�f��/.�~�R&��g�i���N��~����wX�^/��us���=�c��`��T�J�"K��kxɛ�����'�\B��;㊛/{��BK�߃}��~�a�#'P�������)V��~��_Мߗm���8W�]:���K7ka֑^�k����? nj�#/jn˾\����24l���[<]x�)Z�C�Uqhg67t0T��?>�]&�[TP�>FL3�~-�������P-��^t�u�aY���v��?�?������t�����ҥ���wV�kj͢�Ϋ�=p�E8�A�0�:�C{��#�y����}��3��\��;�.`jv��i��Co	p��˴=n4$gb��n��]�B,cYW���yF�8�yz��c�`0q�����ҕ~�L����]����R���}�Xef�J���.�����g[ԟ/��D�?�b��E���x�{�3�;�Bz�'�߇h���*��Ԋ��}������1����؆��e�J�yǙU�W�,���ӂ�⣡�C�E�}�H�B���^30�Ў�>�qD��x֞�74����+��`G��DJ"{c��&�~�h#��mXt�{˴����4�Uj�G�3;�.�� ���eWN짯��K����z�����9��O�#B�,������?2���}m�
e%��l��:�Ֆ�>c��RA�
bWբ?!$�S�q�h #�;Ut�/� ����+B�6]��O>���J����Ea|��]Zy�m�Ә�Ѡ�6��b
6*�G���b����u�A ɬ�Eӻbv�" �h��ö:��U�+Oj�=��;e-�9�3�O�^{1a�a�z��@���H�S(8Y��i�RL���利�_�Tp��O�1y��=�@Å�n)���*�MAo�k/��b*>��A�PM�]���#t%C0i�7�