��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�؆���o��9_��ʵ�Fꙣ>��IG�C�����TD��=��v��ޜ�YU�~EZ_�i��ݯ����yϋ�?'�Kъ�n�tOZ��kzA2���M8촕v�IA���}OK��퟇���\�>�����º�P�>o�QSO���!��3��0O�s�se*�}��ɩY@�js a.�۹�W@`#��ܜB���$���U�(�c`����T�[�]����ש�̊�xx�~W�u��?9���z!��`h<��O�X���׺R���ؼ�JE�>.��g�q���K����Šks�b��Rp�e�S�f�m��XEU�Nh����0��<d�R]L�t���ּu, �-E(L5�x�6�0Y�,�r���pl�Z�:��l\)$����>`Ig�yIbB��\l��));��9���_����o�_ܻk��-��8H ^����nF�P������[���TM��d�Z��� ��;1C�d2�g���5Q왊?���m�X� |�D.
n����#����@g.�7������XZj���^2�J�H2�q�Nĝ΋�RW��9�������1��g<����Ya���@���j���h��gh�m���<��X&�&�z�Sj�?֨;q���+��q�&?
R������f�0p�w-�)���ci7��F,�O,hA>�Q�֒�*�G������	�|Qjւ�𗈎�?�[�3��(�չ��W��3����\��<����=���eŪy�v��3���N/ԄK�#��R���K��2Yણv�}u�T@���<m��	��~���\B�Rٰy�5d��W��>�*qm۱֔�A=��k��?ZmL���z����ɰB��N<N,�ۜ5ş �-�6�g&UE�SP����a9��K��k*e���P�:��<��-f�))ˇ�R��� �A%/Y
��.�xa��n��$Xn�Q�[�U��o�4֚+j&�@Mq� ]�����c�ȣlS�g���\���3Pjv�e�y�$�U�9���iN����Ӟ�uH(�ƅ�?v4���@����wn\�88��G���P@��,����G62v�������ۼ��$���B��_]�OI�&�I��#,@`��q��~����[uoY��c��Z��S�D�&]�ȸ< p]�3A<���.*���?������2Ҩ�$��:�� lO��s^TG�@�*#~���N�-��4&S�?��L�_�λ�b���aӚ����:��*�f�_��'y*S�s����|�!�7�0%��R{��5A4.Φ�ya�=d���`;&'� ����������{�T޲ak�����^
�y�8�?������'KVr�� ��7�|��9��$�P�GAhg O�=��P��7���`M1]+uh�����K<�B�p�9Y������/1GF��x��	��s"��	.bA څ�?5�ǚ]�Q���7��2�:H�l,h���0��i�J�!��L�,؏���_�4(	�
C&ѽ��A"a0ϪPhxʜ�>�߱Gu�"̰&$����rpCް�m���K����C�E�rk�zZ���>>�����ADU�U���Bp��u�h����x d<m�>|z����ll̓h��(� ����� w��d���A �Fj�;;]��|�~�)�Y{g��*X�
oI�$V�\O��٤#�x��oZ���0��%�2�|Ti T�k��c!V޻O�S�F��B珜E<cZ�6�)5Ϋ�����a�7�3Af힛�Ϝ/Q�騶{��EGz�����+6�:�uJ��Ǭ���|���[�.f����!�>��q�G�QwJ?0G.k��˨�	�X:�ޝI�tl��D���_���j�����_T��`ø�^%",ڦAr��X��X����)�R�P����p:�V�\3Ty�O���ng�q-�JfF�U�����/jm��_�=bDS:]D"(|nbZ|[�9�5��Q>��~	E��`�f��ɣ�g����z���i�99����QZ:,]*�Y��*��Ѩ����}:g?�+�|8���g���@�ʍX)�����������	�� Zy N���b>�&���e������F��`S��nc�tq�Z
�:�*ND~>V�
W�%㛀�'Z�Q�CP�%2���2
�Ha�M���?�� �̄�Z
�QMv����!~���\��И��r��|�v��/�$8��e�]�_V"U���/���e��{x���b�����Ļd�x��W�Ħ�&�����B��p��Z2C��,L���߷��)V�W�]��y��9Fɹ_F�����5�2t}3��x,�?�Ne1����/���*itK:b}6%�Nǎ?
���~8&j D�0Q�A��ʷ�4��u��cl�P2���I��@�n�{z�0���rN=�jM�%'CĴ���Zy�p�Sw��cjhK��!��ڊK�����$���[D��� �/q�I��8�w����j��8eLM.f�S�5��Yc�]��l̃~h�K��ӕ"�w��5Z�s�4*�&�t�/����ߗ#b���0� *[�_��Ш�rso�v�-��V7�gƎ�)�	�@�Ra�}sN��tO	���в~���ך��t��|�n����D���e/H�6��)��l��]�K�O���ۮ��PӟQ�Bp�,�r`�w3��YXBrq�77 ��E�>� 1H���Ґ'���a�qRӥ��Q� n�Sr�� ���p)�NU���)%�����¼�a��S*P��jb���9���uz�=�letq����>B�� da��\z6�rN�L�J�ԝ0���w��B(���_��9.��0��@W�-��K~>�f�2%K�-���9�w�$�7��;q��g7����C�����]x �M!�B��z��6(|g�Xz>r"��Yy؊������e�CӖ�B�G����>���1\d�l]S� �wʶ�T�G���ITT������_Z�l��%|&hV%�6��p��K��M�����즰���L����E��r�m��L0������W��8�)�	���� rc$'HQ���l�T��4��Ud��NI���oY힚�]���E�g:x���[&0��$�;�c��6��pHjKC��-��u�������eԒ���T�.i��{��W�5�$��4�yv�G�C�/w��a����Z�BUH�nuv?��ݢ���$��)ww��q�;�W���)�g�
��[�����:L*�j�e̗��U	ϑ�["�g�����L囐3�Fƿ6eO�sQ	W�p �;�xR����d%+�8����L7���w���7:z�֍�tx|tp�Yq^�-�+~ZS� �w	�*#-��',��J�ѽmx.�v��4� Ҁl���1҃ ,�W�3��.�k�=w���L���Sh'��_w9>���� ���~�7�5Gr:�:[�]5�an4��S��;��v�w�Z�,��l�lЖ��Y{�ɪ��$��|�R����qȌ�D�i�=��R�'�늕�8`"KV+�e��k^�2eM�Ύ�Dek�P�82�MC�J	B��
�
5�(���G�M��ԝU%{`�1����+�`�F��.�I��)�o9in�*x˯,� Q�k#4���ͤA�A�E&/���(�9yB�XXB�&�Z����cm���Mf�b�q�1�������h{�g6�˧�}0p�\;ޫ�LWydw2]��EE
�گ��p��Q��,%�e���]~y��A]�m���ty����#��'�f�!�����i	���C���Ex�H[���lt�;�G�%7l������)d��Ma9˥��T�%~jT
�-������}1r�z�e���,�{?B��B�rd��Me�Dرߵ�N�P���"�>�&�ט+	1N�nLTIބ���SGml���<,�n��,��qF��\��obbt�ڪ��c�e��y6�Ѧ�	c��T�Q��H�T{��ۢ�0��@Ȼ����p;{ȒM�18�.
��#�Ԝ�y�ⷦ��m�������Zu�1(�z�Ѻ��Ԙiw���- �0�mѨHB^
5�,]��4���Zė$P����<�M�c'�Wtݸ`]Ŋ����qo�p�����2��
S#�{�}L"�0	��朳.�g��D�SF�k�^De q_{�4~�.*�4rXxo�Ѭy���8��1ዏ���L��E��Nv���C�~*C����kW��W��*LV���0qK狪'�Vt����F��B��O���#�I��bH&U8�����pl}�R�|�[�8b�0�cP��]C9��+SJ��q�|S�����K�#Œ�Fz.���_�h�g�Ro�<`��^.������iz��`>��(�{u��5=�F'u|�G3�H��9{��M%кu� a�
��h�?���	�N����݆�B�]ө)&n�]�B%� S8��8�j��"�Ɋ{�ń���z����__u���v
h#�����W����PG����F�~o�5���9cKL&"�	�4A�A5� :a�������O���91o����),�y�6�6����/q ���f���9��i�^�V�GL����7O��g/�!u] +{��䄊�c�R<g6\~�ST�A&;c�?�(��(W�4so���ϗb���E����d$���a���|�y����O=�!�	�!���ֶ'�ʏ_y0�:�|l��"n^_�]}���/Y�>�%���e��-����Jf���!M8Ɨ,h�Z����=/��{\�,.E��J��wj�����D�����.��P;��5l_��!�����:���E#��A���vD�F��	�r�z�Zh��2`���@-��ah��}�+$�m����K�L	a�%�A+8���,��ΝS��w���F�D�S��oA�����񰿰6Q?��s�����EF����E܌��|�U���C�(��
Q����N8 k��!�=���*��j�,�Z(�ƚS�>[��kV7Q�B�*�G������$@��kQ�wL+-js��������9RC�=�f<��^f��X����Eh�Sֵ<>ys����)f��U'[�e�#f�G%&���Bn[����Э���x��\�u����P{�uu�s�C#c�	b{)'����S^�Bk��b�i������&Q�*���'&��#�i�j@�J��]�s�܂L{��{�YN�,��\]y1Jt.R�`�u��܈B���#��5ݺ�`�n�"m�8�uX�-F ̪w�m�*2�&���e�za�˂�]�H-�^/ķ=):�+���2���鮺K�L����xfG��`����l��<�Ul⚂��8�+�)�`�L:�� {jR�.#�_ �Mn¨��m� 5�jئ;4��A-��@�Y��v��������\�9��L`\�x���~��X��d�`{M��o�y����w@R��Hұvi4��s� ~�k�a�0Fį�f:T���'k�-8Њ��Ǡ�G�D�zx��5�o��O���x���yt�Y��u��L����>����bC#���ė�]e� ���i���aDri]<dǇ�d��p�5.��A��&���y
�0���e�b�X.��}�Cb��D6���'��B