��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM�
Ɨ�j1�]�*7󨎯c<侤�ǩ�] �`r**.}�����g�9�<^�P�_�01���?3�e��g����͏gE/ߘ����>#�_f�Nq�H�b����t��Xc��Y�?|/��Jh���La�V�31;J�ݩ��,�7�C}�v,Ȭ���ߠ���'���:~�����
��(RW�Y}4o��$���!�RX��d��8 �.nE8�AI�}ܪ%9?�\��s��9�����#��8�D���;oǕn�r���U�9�8��[�%�m�,�Ui�}������p���t���c����^��Űs@&�Y�9�:!�������oцIݞ�VKnAV�j�)�&9e����O�F��]��^'��Ǔ/�����4��3
�"�u���R���%�S���n��ׄⲗ�du�5�X*�������V\���Ĉx��|-�*?h�[?M���UP�|����mAf��.G@�Y��r��z�_H����8���L���(U�^2�G�J�@����͵�z6},�8�Y�qO��_��C�4�j �� ̰ë�bC?Ԡ+g�Q*�=\&q�a��q��Ǫ�����(���#��b�k,�?�e�Wyݦ_[Q|t��tj�GX��:�@�9��r#��j�+����E�8O�E)�� ��`�[qo���͐mo<oO��2�
�A�k�7N���eD����u8iCTҩ+��a�l���!��^`.
���5���O0���K��g�%����c��p"*�*ݐ^����s�
�-A8 �A`Ȏc���`��7�~2�z]�L��s6�V�����@�o�n�i$��]��n{�"ʹ:��`Δ�ｫ����nTx�v/��J:�W�V%�K9"�%��h�tW�X����rw-�46}BS�a=�����:`'���(T�+�8��I[̓_U;-��g�++Q�j"��׏�Wu�13�B|��f9蔯B�*��1_r�k�f�G�t�1|=ϧ��kt���4�=�;��x��;vz�c�h�sK9�+�"�8G�����=�u��`�F��G=�_n�D���k�	�դ�T�d&d��2�ߏIUx�F	\n�O����YwX����l[~�R�B�cK~'�f��ڊؒ0�i�z���Ax"J����9ϗR�{ �����`
�*äC?t�j,�Qi� 8�m�#]8���3��8(��=e�N�!���I�iۼo)'z��ଋ��`�)�U�>Ci�Lt�Jon �ڡ�D+�cMć�|w��Y���܂�� G�I�2�S����9�ǜ��A!G �T��������֛�p�h�y#��w������]xZ��@�jT���<���)�����{4;��̻�D�}�c���_��e}w&��h��xg	Wײ٘���o+1;���<�c���9��.��+�S��͆���H�a���z��V�_^E�y�()9�a�}~�ܧT�g�jI�#�K}��S���+(�(�����Ii�w�fMPc�ϫ�\`=�]B���k�������]Ē]v{/f��1
�	�b��Xf���c^���ѐov*�����X��%D0�S���O	E��qm +�C��YE��z1���$�-_ܩ��0���'5�N��R�Dy�x�*G��W9e	�i.[�Vd������P(C