��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B� �⡐*��D�k�(ʸ;+.~/jը6���1�@�P.kZ��笩� �hC�צ�'� �.��%�x�WOL�^p^��L���Iv�shI ��>�{5u�����9!cDn^D�9�b�mp�r�|~f�l��j�5��od95�� б��P�a�f��>�l'�w?5!^il@^+�>L�a��*r��w�Ś�М�0�P�c�͏�B:�I$ZtE�Cd�T<�	!3JCǮ�8Գ�1��t��>o�<��������vY�s��R 諚�̪T����fo���)�a6��l�Y�A���toq8�rݢ�$:+�~�P��# ����dAe/���A��ӳf���|�K�F�!ϵC@w؊��)��ZG����Ǣ[M�iS���Er�S�����§md���k�sR��C�����u��촒�7%&�	�uD+Y�h�|T�*q�o|�Hri��6 B* ��+0��E/��{#��+֕�m�n�3�#��J���B5��:��!#u*�7$��6 K�"�ދ��eq]�z��z\*���>�k.%�Y���9��ن�Æ�Q^�v�)N�'��RJ��p�vמ rˢ�+��S�P�{�5ymz�UxuvKvE�8���n=�U����a���N�xH?�a��g�FS3�0	L�����[b���1��T�����c޶�MM'�Hg@k!��v�9�`�d�vE�1uى7q���KڬyxȈ���n��'��,��-Ia�`��U��������B���y^dr�u����ſ9���KU�h ��tjv����Y�X�{Y����}�<z��O�ȽN�(�&~�m�H��2KςW��V��2�����I��Ӥ�����I�,�q9Y�3��8o�=*C�e�l�2�w��Y��=���'їea ~�o��Jw���-8[1��f� �#m.ժP���I)aO��,�&jq���M���T��Y!�G4.Г.�n=��U���.Yy�s_3���1=>�{�d�կ�����,`�^�_�?9�b�%��������\�8l���-�KQ��a�{��� 3M���!��$׏@�}�M�-j��+�p��_G��xu�F!i�,����E��]�Mm��xe���r�G� ��7#�6}���mJ
>�Cb�e[�~�9�h��z���p����m�t����zT��T?�zKg�;�! ��~\3��6;H#���}���_���6������;oʞ���EB�lb�xR��1�x�eݷ�xGZ%R�Ȗ8���^��}+�8��>v��������]~��v'W�'�4x���5c؀A�Z	H�S|��k���LN�[����rDL���|�RTc�Yo�%�-��5q������HSu*J���(���Z��L�Q�c*�+�D��� ]0d��u.JG2��$ ��X � ��� 
��j2��s1o1S�ّ`�{���zY�ke�ǧR��Y���� T-�d��F��䛱�(RS��c���dt�v1x��r$8���JZ���#퟿fz��;�9+"|��G���l�*�,Lh�J�l��a�a�&��u�s���1��1iS���0�%�.�[uϜzpvu	������p���G�Rl���<auB�]-	M��k�WN��7�o�AO���"��iw��_U�K��Wx�d�@��ӄ���b;��c�A "ʨ<�_#b�£1�܇!��J�$��iU�bB"sq��F�wwb����U)�K�+�c5�Q�@�R�S�$�}�
��%���v ��T^]fY=�2� ��XI�Oo�7�U�	�����ic(y���Ē��xI�c$Z!�5��P$Z��Ԯ�Ň8M{�O=/�IDJ80�S	�+������`u�Ѳ��%Nx�NU��[I���&���6�9"Y��̲��k�a;ᒫ���LC���C$�����BB�Ҳo���h����������`+\ߌ(@��.�o�s����1����2B�Ⴀ�N�/^t�JS
�/}�]/ ���o�<�cj��;��U)5z���`�{~D́��5^`�7Kj�{�Q,P���)��H���h�s�u5���%���&.>(75�P�*q�wђ�<�T�� �p�v4i/8D�Q-����[���(p�xYb�]�n(v%���.�
��U`K�zبH���(����`����E�W���e�VN9�����O�%�_�����V�刽�l��¸~P������Լ������ �E]��+�T9X��s�Lke���VI�|��w�C_��.��l^]d��T\���,�AJp�X1#��h Km�2]1�m�x��9�;z��4x~��B�q�"0�A�,ZdO�����$s�C��]�l,��rL����b) N݇mS�jiF�bLv���v���6")��ּ�����Û��N���2�<��i�)�i�B,J`�4�#�d��,�W�g�,��dǵ��4H]������}��L�6�L�Ήr�T��.W`hSC�ّ�����R3�n!�N���f`O��zb���w���|������7	s/�#S~�����|i~���}\��d�'u�DpX$X��<�C�t�(G���gj�{�a/^j���`���ju������0�iG��+e4�ٜ�a��lpHs���GV���S�1� S�]�h<3�k4�$�(=�J�R7�KA���$c=)*���e����42q��7A�{3���|��H�q�Uw=8���{Ǔ�d�Çʴ��(	z�3�0(���a����[*��Fx�=����͐���E�[c���u�QM�?�O4a.���[ե6h֣��4�[��N����"�J�TmGy��۱�<�a�VD���l�!A�ɣ���K��>�����8N;��#��T��'�ى����ǝ�1V'���m�����J�j�輨�6�yՆ���A]���,�
�W�����w@ʈ��f�s{����Ĩ
~���D��\
�C19�4u��p��"k���<�*]>�����O�i�TB������͜q�mK����CV��vN:Q�/�r!��Ɖ���� ���
����C�+����E�cY�<���S��xu��I� aK���G, �k�#����Bg�50O:���	�O��F��*Z�JWՆ�Z�UP$[g%�s�6_L��A%���,����/��"����E9���਽q���v�	ӱ�5���G�H�	T$2S�
��tn6��C�����Pf�QL;j%��E�4tb�Z�@�}�:6`Y��5��}gc�ެ�0U��OX��<@�M�A��~]��
�S�=�~h-fQ-τ�s�&�x��5k�ߝ���$��j)|��+���BPBҌ����b��D���r2�D�z�a��5"	eU��73�-��$�w���`>��Ө*/�������D�A׈�<������C�������<0�Hvy����	�ދ�z�rwkP������N��=Y��J����p'#����+	�]��_���w���̒��LcΙ 0�p=��&�@��ߺN��e�9T��*I3�|�%�o
�OXC-�B�c�;��'���*�M�- S�-�:=�)�+sc�E3�qB~��@k)Cm�>"�j �r�M�#K8���̷q����>���E<*�9�47�pA_�A�p~n=EAU��LuN)v=E���>��23=.K'*_�9��9NA��m�l�Нq�/�N���W-ڽ�.�����7�O�zK�ʉ���#DU9��A�#jD��B=�A
՝0�{퍡�8��B���pk�~��YH;���o��4��"�JN8���x9��Ji�R�>��.��p5d**p�sƒ�c�`׏lْRu��L��2�P�Q{U�!>oJ5o1𿠫s��5A�Tgh��>Hw�� ���j��64�&W���%��#{o�P�9����I6a�0���G٭:g�yl�L��^&],o����O�Y{����V��ɹ��V�{6��қr7�%��1-��;!�"~��gra�:�^������o�c$#a(�N�>
CҷP]�gMc�n�3�,Λ�f�f�ؑ��\4F�$���O��3�%�_���yA��^�f�O��Fz�Ⱦ�3es��Ay�\��S�D�ث��@:�R�y�ߡw��;Ñ~#f��}	�W�~�	�,R^>+�'�Wο.�G�[�Nӏ6}�����`N�pR�&�	�ud�i6NS��d����̪_4�8�8z��Oj�Si�XC�7H"����/W��mھ �m���H�H�B0��j���X����Lzc���(��H���U���!k)�����*����t���������=]���<b���Ξ��;
�1z���[�i�q�v��dX~L�mc��)>�	(s��M(�Jg�U (�30l�X����Wo���`��f�"�c�l$�Xp�L�K��>����d5ͷ�1.���k���9�G��Kۄ�����x��6]ί8�S��/xQ�ʛ-�Qv������E�*�=S��ߟ�&����������E�z�DV���O��0��>�g׆���s�Qh���FIH������QS-��R���4��B���v�Q�8�����dg�|h\IC�&�BH>$Z��\ �Y��$�A]D�	]��1<���FP��Z�xL!�f��^�֥���1��5�!�m��;;�=F��&T�Lԯv�{�5��C.M���굦Q~��`U�N�gV��Bc��s���jr��zl�y�K��|��mV��zm;�n���(1����v��l�����-a�6N�X����:��L�~)k3\��G�43�ioÞV��a��l��&�a�7�4��p�5r I/g�w1/3�)+|�u�&�:/���� ��fiʭG�'L%G,������]�jXmSq³���8"���em	���.*`E�x��m&��Z͛[����J�s��-j}�d\��nKu3��m�Uҿ��D����j��`h�r??���`v	M��� 4�|R{O��T���Gâ�&�k�u�R��9^O��u`�1��Ӭ?Ѣ�	ǐ�E�Bs�<��m���Pa���bGk�7��+=��ԗg5S�r#�p6��U8p-+��[��xf�$}1(s%1}��ny���S��k�2�3Chs�����h@M�;���)d�N�ޏo�
r�H���·0���C/���4T�'�X�tVQ<��z��ld�'���s�*��R\���,��JJ��z~G�fY�M,M(@ |S�F�g3��<�#c�l�6��Fp(���_�3��N�*	����zD'�dm��ό��_*�{;:��8�Z#Ӊ,*Ac�3��t�E:�K�Z��~H��c���E�S��T8M�b��l�}�`�1X�Н��Փ�It�}̶ �4��;K��2��'�C9N{�͠�E�A&r�&9 ��b�@��7�� �
/ m<����>����UeE��!ͺ�Μ߂���̭�GN�>Q�=�'�^�/�a|tZieicz�d~l��8�_��B�� �hg�x�e�� Ca7���Z#���Py�C�v����	�����{d�ԭ�Ã(�b~o߾ݔ��_�&�7(�_���I�-�Kw��-1z�O~(�Wt����e>ǹ���B��rd�xl!��/�{1J#V�
xc�8�aR�������I�2EP���v�����|F� �hf�k�*����O��^���O��r�T6xrM��U���d��:Ƌ&f�EOq`�$wDUv>�����"b�{����e� �}����2,	<�T�p~�Ra���b��曞l(*^�h��C���]�m�hr$���2}"���ل��,����y��7ˍ\N2L���l��l��˗�p`��I�r�����R��(�Ӹ��X���e]�:*�Q�_�N�\Qƕr�, ��Z.6�svn��'���Ufp�g����O��x�K��L]޿�Soֽ��w�u��d�u���c�Z�������x����}Zؖ9){�>����M!����=�����_q�B�r��t�( ,$]Q����+��[�|0����=[%Jp6�EF�P(y9��]���~�#͝j#��m�X\`_ۥ�md�{�+�0?���кŴ8���DRfl��R0����i��8|YT���U�|b�!9 �6Ι]�`�^�_���c�B�3�T���բ���!�	ӠG��$��[����/<�A�8Z�d&a!k	�����K�ط��Eq�,�瑺�G�R5��7t?���B���#�r�΂-�? 㧝�ٝ`ir��8�(�~���q�<�C����;#�� �
3�2_B1�"�$,%����.`���_qC@��^3��oRH���Ò ���4�z�3�����/�:��"`���c�l'�R����&���Q:���3v��lW!�	M�q\��=ZVC
�ϓoP"\�V=�lĬ[���,_�'
1�э�ډ�j(�t`�X�1�����d�ā�	�
8�ܪ)|V�9|p�T���G�8e�v35:����,y���L�H�+��X��o�E��n" ���u乓P�74C�:տ8�ɸ�&�؊���\��Ƨ�+�|y�'���?`;l��{�H�t�.J+��b\�֗ �D�i��
����}AQ��oI%��O;��3d!�G�t���R����@���<��_Q[�t��~�0�l��T���X�4x֞Йb���
D�D^�[j�N=�z���8��D�#(��P����ү{�q;��V"��+�����%�Ю6+��<���YȂ�:�a��	64�q�y�����-�׸�g����E��V�w��ߕ`=�J#�����׊!�\�]���<�a=h-�TN)]w��GWJ��/Z"�[.�x����/�uK�ɬU�iG��eSRF.�Ψ�9�"�nW�h}V2�^D�r�k���9��(���3N���ںڀn��y�s3��m���p�1'i�ԃ�yS
���R���kk����uz�H+�n�FJ�8�KWЛ�`(���(�⩓�w���G��RةS5���!��K��`u�"��I��R*`��xG��5�3�pD��Պw����[P�D��F�rXk�ۀ��߈Oɪ��q��e�| �F����u���_�6�����΍e�ʻN4	��d���ߑ�F��:�Y5�.t��#�Nȴ9x�~Vذ��=��v�JZ.���U��0a�!
�J������_֝�kh�h��\���&����5����Y������<i�{���V��:\��p����>l ��z�6��F�Ed�ǳ�I�R:G�Ŀ�:���p�Uh}��<͡I�KN�)�$�#�c��>�}'1/�z��Ep렌3���7��/3��˒ͰU��<���߶I��A-$��%S  ��G)�a���1�k�|)�qɒ�XqӢUp$A�P�z3a�9�紳��P+Z�*�B��y��;�M�rP�5&�Є��jn)n���/��c�;{�2��(&'�����Y�'�%�\i�v��<��=/FI�B��ב�{UС,F���|���l�,Oj�ӯ�J�U;`wJXǝwsαs���%�n <3029�	� ����)mcnh#t�5�E���r��}?����B��G�c_������e�j����;��4r<[�Zstw��٭&Y�o���V�˳�8�Tb�?l��,�wUr DO`����	wѩɮY�4� �@Y���w���R4��'���|y�?��đ�2fM���yb�*��Yb~p��o�Ґ rڿz��bU����3r�8�+0sB����I�0[����v
F�O/0PL5���h��Wn�f�Hn?D���:��x.�Fbä�ˈ�Y�o��/s;n��Z�G�;t�P4?�Tbn#��/��ի�-��f��S��)�r�(-�wOǦ�|}�F���5��)�E15(���<�<�]�^�i�N�N
e�����2���v�Td�e�GMnR5�7�����D��A7���$J�&=��� ig��$�pW�I~�c:w���D&!6��0?	M�t��%�pD$%��6�T��I��u�a^ޮ=�(����a;%Ǹ���#3War��T���KN�!�L�N@����*NA�� <�`�_	���ݚM�n^�,<����/J�Z�hI��dL/^˨,U�=��ј�m��t~*�B��z�NI���Y�U��I���#�������_>� �S���P�o�����n��;�������qo� ��.���hB�����U�7��I��L��v�BxT`�w^h+����T1�S��c���K�Jy�n��dc�L�va�;H'�b�bI�ڞ;����i���q� �s�l��TǚƛU)���UB��ږ�_	1u��F���Q��\_وi&�HJ�6t7��k&W���2(՜�t|�J3��Jd��s�A�1��8α5��4s5��p4�}(e�@����䣭����j�n�,�bD׬s�@��>��^<�Bߓ�n��b�$}����r����������V,
>ln������P��#�l�+�t�~\ڽk��,��Dǟ��/^��G�RQ8�u�fjI��Chޘ}	��)h����6A'��Ǘ� z&�u�^�fbjLpߢAGܱ����K[�jW~��: 7cW�/���;�,%�$���D�,](Ǫ�lx�Nk����,��_:,�����L��ߨ�K�A��c���F�R�Bw@8�=ʣ���Ӂ��d�Q˕`cb�.��o����x����2@<qSl��#�����۪}>�z��֒�F�v9͙��D��m��Vu��c�n�Q��ꨎ��A+��JKу�`���Қ�+ƚ�5��z�J�|�V���͇�� �?3�5�a��aQˬ��b)���\_a�3Wk�X���2F��������yO�㒟�����p�٫T:������;ğ��[/���h���^��Y\~��6��I3.Vu���/�"��v{6
�Oam��5|
@�6��{fW&�r���8����ߓ���] Q�	�/.:7���Q4-=�=k˱�r���2����^ ���֛�����x-a2v��?�bo/B_ZO�vv����)Q#�Ћ Ě���?�(%ݷ���|Q_�_���avhh�0J��~) f��ˑ�J�GP�X���[�77�*�3lj�̅��Lh�͛XR�����}�N����E��CC�F�cW�Q8M-,T�� opS�u�R�����!Q��~0G�֫&ݶ�/�C@��H:�	�~��3 �*�3�($�S��)�㉺�X��Yɩn��N2#V�3螇OݜX����T��l0���X�f�aJ��Ցܰ��յ;>�q�C�'.	Y�FtG��ߓ�i�f�&o-kWJ�hΔ|X�5� n:��7&1�ɨ���Zl%���?GpA��M-5c{yo堇b	ѹ�(�ZMDj�"*M��m��@cj��Z��z�U�r%/���N��`����m�_���:�rj��u|�ш%��4�SA� ��ۜTq�$��߮-��w���J����V$�ӕ.�s߼˖ǀ^��EYNr�}�
�|��n.Q4BD�³��#��.���ϑ��'U����Zr��w���e9�_]���YZl-_�\��Q��\��0�L�E֦�yT �
�<��pzv��L��������sЪ�y� �%�_�3�����뿌u�����HԌ*�bPNq.�G�0s僀�7�3A�2�0�������v%�o���Oi]4�����,�"@��}�(�_��R�#��<%1�Ì����*_�Q0�+.L���#]�N'T/	�OQ�/n��U��D֖���\銉�cO���3�OE�k�]d�M=����w5�X��N�z�0C/�|��C+u���ٿ���$rI�_Z�h��|�.���x)�|����DoY��}	j�edD������F�Q���M���d��&�Bc�ֻ�vV �:oqj���A&��|o� �ir��L�~�S��ļm��:��:��܁��q[ݝ���^1��1*J,,w���`^Aj�$�U�zgo�;p����>���������f~$g�
c{ˤzϢ%�ML|5B��>��L����KU*��@m"׈"��aꏑ �(���C�S�����	�J�S�]�o��4[����?\�_r5 Ei��4,�R
J¢��l��`�p�Ү��}��Q����R�ϨtU��x�E�N���
��M��m�D�Q�=�c�S�7��L��Xvt������td�N�Y�< �pa�\�X���ѵ�3���K	�K��_]5�	�g�	��Rq��T�!�Kn���l�;��Bs'~Ň����,�L�!*l����q15NU�:ZY�2����v������<���y�\Ѱ�D䬀�n�('�4��Y��L!���t�A��q�2c�y���|���~��N�8B��=a�DV��*�|"u2
ql����fJdCl��n����l�0kIA*`g��v�^*�`[�U���M��l�7 ��8���c}r�V��	B�� X���uz���4>��d bK�V��e?�\ID#]��\5�x��/'^�\��Kk�Lr��Wp�l#�4�u��,��Qz������+0�km!�i���;�Qy�=XTW~�.I�IΒ`�/wd=D�C�g��$�am��tL�:#K{���]�����e�L&~��V��IL܎+ۊ��;��A���ČZ�9|���-�Ǡ��U8cS�,ƥ�t�1M���ɱ�s%���D�?���=yR�5�~{�]��wN��g�sh��F�)&>Y^��^���4<�;
/��}�Q��in����ko��o��9���R4�s����
�a��v��j�u�D��?#X��[J�'�:��C�T�ɺ�ӵ��l�?�V�>�5|��u�v���\h@���!4QBZ�ٜU�Iq��&���J��Fq�}K���������E�#b[۩sI�:��I�ؘ/���A̸�9x<1Vy#F�l�	�2`�CWO�`/�C�s����s=Z-�.�4�f�6|"(�mlg��q���30������ ,r�5ԋ��z�]�LaT��Q���]:��7L;~����zMz�ũA�M�[ś\�޿����z�)��G� L�i�ѷ���a�h̊Ad�ff���_�Un/�+8�sA���[T_�\!����ሰ���I���ս�zlU��z{��z�<QoF2J�Y_���8�.1^��t���?`a�`�D�Ξ���9A�?ۘ%S��I[��I~��U�����a�t�8�ڜ������F=|�?N�.춾�1�M tܱ� >�?�h�''� l�%-�|vE�>Bv\���9��:�J�d��V��%@��-��r�~���)��-����ov�}�R���^î�F �.��p(��D�GkdI�먬�L��D���5���y>E�6��<C��4�lLGu��e@��8�U�&?w|0Y��
$�W���WZv��"Ѝ�]ߝ�;�V��$<Gw��zi��P��5VF�/Q�Ug+��T]&����5����4=�-���#o��r�֙����
�Rs���)а�u�g���������#�c/ɠx�Rfoá~OU8��!-2�|�USx:lT�&�6�yS�o�P�Q��o����r�����E$�nk/�$����W�fD%�m�&��)�L�W��b6��:��4�W�ʏ2�g�9��U