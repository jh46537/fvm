��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"�.0�у�[�Hd��r�vJ�?����t����Ζ6ݙ�.�?X��^T�������T�WT#T��}�)���yZ<�Z��7_����_�CX��(sU��9���8� oR���/��m�GZ�U��V4�W����5J�X�-h��d��$���6i�S2��Ls&x�~�F�ϣ�
չ���vp�"�ӳ|ЇH�fs]ЯϦ1�Q$ [�@9pNH&L�� 4�t�4���WXKp��jq[
r���:h�
y���@z�����n(���ަ�̅������c;(��8�h�~����u�ϊ�����&�,"�3�6�����JU	W��qL���pn:��[�&�1���bl��Ą�C�+�&ؒ����I����HN������g&�WۻM���%K��I�=�kx��� �;^�Ǵ|1�8g?@ٚ�.���:8�|��z��;|�&��FYU=�>�.c�!C:�p����1	�9���}����M5=9��(��}푢i�8=�Z�����*�Q���@�.Z�%�$ 3����Dؗ�SA���{q��g��d�}"pB�7�9u�AQ��6�qGx{vf��O������s��Yۼ�S�N�aXZպ�@p����O�}C/s��hj��,-��(���: �\�����T��D��_���X�O�󦯞6{A5-����� ?*���ҫ����>��;��eRy�0l/��UvE��,�ݏ�ʩPѲ�a_x���Z��`_����ߦ��2-},�6��*@�YC���� Q�x�<�g�a�<+"<e����K0|+E��qLZ�f�P�RHGX�Q~aA��
2�O�����LʦK4��#��w�)��ꢚ�v��9�ȑ����)�_$]5Տs.�pr2�G�(X�Q�$�nD�B�{m�Mم�������k`\�I葖�����E��6hi9yff�ۋ;y(�#�0��7�jq+�]�D�#?�9���V�IX*�����>@��^u� f��^�8�d�f5�=�7��S]������Eh�e���<�I��O��=���K����W�o�-��Aܸ��"��4��V)��\��PxlF�<�MR�NEJ*c��gm{4��ڪ �3�Y�qI����׿y� ���?EA|l�g�W�
�?���/l)]���U��QF���U�TnD?:�����>�	6��1�@:�փx��9/��q= ���<}�PD����T2��ϥ��a�S��|O(��ቀ3/$�_�W'�
�MM�B�I��4{L�� @!�{�+�S2�o`s����i%Y:�Dř@G��O!p�B<v*;�ls�v�+T�5��Fw��%P��r|��,�t���tn<���.�̊{{���(Un�i�5B��zw*}��J}jOC���HsVM+ԋ�z�2N����V��/�ڮ�lƶP)ު���x+�}�2�/X�P[͖Z��iCa��2~eC�����`����E.�m��)�,_�ӊ�(P�w�r���H�֙�+������ެ�ݾ���1����82��90K���4�"	�/h.K��8,�/]�V';')x����u.@n�x����CX	pZ���g�cU�-hM��I���#��½q&iu¤�Ɗ���"X�Q�z����!Rk�gW�'~Zㆨ.� "N\\�P'ݑ���5�L��GKv��]�'��^��VHms�,�ӏ�$0m;\g���^�\ �vO���%@@cX
���JҸI��Y�d&l�^h�R:8�4�^s��x���e���F�m~@�~�F~jF{��)}e�:>�|�|�o���?!Mm!��/�͆�:>J���ݼ����{�z����EB���c����t�]�wK��qce�J&��P��DV�Z5���7޴����B���A�!��P����'�`L�6GU����5k���h؛��#ˣ���c��M�TB��[�	����^�L5Y��b�зG��'/O��0[�W��,��U|��u�N�9kl�N��	���/m�f9C8gPp��#ΛV��a�5�9��-���`%Kmcw��ݮ� ��SV�S-�u�*���.��O/������,��t�UA?MR#>�H�<��wƾ˕6J}�>ƥ��*�rߟT���v����u���E�W �7����n��q�����چ�5�1���2+d5�3����/�}d6�,����ַ��c5�3<U?}�XR�/�!���В�I#��v0r�C��k{��#1�]*�"]�x곺ӟv۳��7x��ns�Fwk��P�7۲hc:�����?I�H/C�1���3y}&2I^>��`l��#��Mg�S�҂\fE�"����J�]�d�lI�;j'�߰�O�m�����Bb�S�
;4o���K�����BW�ErD��r���wZ՛р0B�P�?�m~3[��\ �}q�	�����~��*�D�cTy
�LP�^Ț~=F�|�%�m����e��I�R���4|n1���@�?d�;љ���Q�ٰ���Sk�Q�I��Z�dJ1�u:$u�R+K̵�UH^^�Ԡ���$����y���*t������Ǽc��p��� �ֱ#�K����C���%�2G����o� O��6�I��o� f�-��s~�8t�Ԓ��X�p������#|�<n����K���&��A�@Ы������������@7RX<�<��O���9�Ύ��bj�����ܞ8G˝y�S�����=�а�MÍ��c����Y������5G���PTKn^�ݴ��fb��ITZ��|q�An��1O����T�|.1:Cg���X1��E�V7�T!�����o��3f.es(v�5a�%g���Q8az���$Y��SϿ�QC�K��7��<�Q���:Ck��>�$�V�6��� ��n�n|%����G`AB0DDOt��h���;:5�k��H��t
FU�rIܼ�
%�E:�ښ�D�~;QvO-�]�ҝo�l�;K�-�P�B����T��#tj��6|�>h�_`���+�:c��b����U/񣿇�.��(;��3�+ؔZ��� M�֪P�}+b7����M���>E2��w���yMu���S*�QM;��3<�����Ύ��`�"��Ƭq,~�=�g�=��^�r�1n����p�����)i~	�ew��� ҄ۼ��n�QF��ѹݳ>���6�Nقٜ<aX���瓨���{�ٳD=��P�ah� <��"m�@Z�����ƨ.Z�}�bՁq�wG��o���S�J�n���$�����ZB������&M�I�:�F�L�aY��΄���_����P�#��c�p6�`���N}h���eB�8�儁T~;�'�՚�|Cp��/����e��x�����=�5"��˂a��W��S5;=�C��D'�j��^ <Z0F6���H8f�>;��ǡYΓ��c8������9�8-~�H%����<�����z��t�v�V�5O+FۘzP��D�]�.�	�qS[��N����N�2��=c%�9 )��t�K�
C��a�ji|�Q�,���.>[y�&�&)�.w�>�( �gL��&G�Gh�D�1�|�Z%����	1q|�D2Q�(�����\����<���C�6���hz����B��g6LSu��jo�#ܐs��"�]w����80�n��,M�������e"��r�.<U\(h���,g���:Do	��&�3F��-������Bn��3�����;	o��u^v�s���__D�9K���ĵs_(Ī{���P�K{�)̡NO����kIG�U,�u���U�-�	����ケwzNL��:�0������
7e9|��RT�x�8�w�0~��UD�g{V�����J�B
e�a�w�;M����u��`.�R2|5�.��:��k0����X��W�x�����t�)�g˰�f�E�)� �eҭ�鋈���U3�r5����)4Ԗ��	��R�Pf�d�0�v�b=ù���t8�Hh"Э��2�� oi6��XI���yʄ>�O(�Z��'`���d��`�G��"�u�/WTX�1�1h�gӊΫ#�r��f��V��Gx(��;�(�R����_K����k�0�A��P۾�M탓��G3�l���Jn����yie�Ѵ�<�'�7t	n5}R�'җ��'GZ4�>KJ�h��*�����r��.Yb��t�LVު��@��D�s�v3Q�QE�O�'�:
|<t:�1���<h'�&���L��`Ĉ�#�֨byǋ�<#4�P���Rշm���>�І��wW�uj�_'Ef,�M��6ն��ˁ�t9�}4�o��b��ʋ�'mFY�Y#4��8�¬"x���������|�=��ʿ�� ̏؏�ƌ_��mL��
����y�=�T�16��	+��z��r>�u.�_z�h�
SB���*�E*�-f��_c�����7��;^�(��%YſP��ճoў��?�5͖��A��.tU��km:�e,״s�Jw˔�s��u��o��x�Q�o'��э�D�d?��������C����nR�!�E�����t}�˟I��q�ƒ���u�t&�*l����������ġ�K��S6�oh/?%uK��X���Sԭ�_Md��<�{��<5��E������"������Z� Ѵo&x�ȑ�^ �z�-~���'p�f6����y\�������Z�v���찓(S���B��Y���Z�������5��J�s|��1���E�W�>δȑr^#��ץ�w���7��M�!z�
�����2.�ݍƛ��T�\���*�a`���i]����~��	�H�=�P��c��ןn]�U3�Φ����ԉ���!����h��gC�;�w��p婆��c]<rS�X@����pT�)�=�7&���3�C��0$L��y/�9'wJ��4�����%B�t�`�����ϲ8�������c��|h�@�k�ć�0�g���7*O���<@	5��M���ᨠG�i����q���7���v��eV�uc�!�\�����A��^� �<+����ni��'�9vM�=R0���z�@�8��q7�H@
Za3�$�Gv_�D�w��ooY�9@�� �q�������r�Ԏ5���l�C��\g-���4_�h�T;��
Wim��"6�	�R��Ɓ�d7�.�\�p�x��v�|&VW�j��C��C�ピ��R��D�šк߈��?	�j���RX'�ң���򎌈!�����W��}`(g2y�?�E�T�Y���R�0lV��"SiR�N6.�������=
��H��q~�y���/B�+����u��|���˸�9m��#�J��ȋ[e^�Lu���c4Cӕ+*�x#ꪒ׳}���v��i16zm����XԛrM�ˀJb���,�\���G�ͱpйY4�&�d`{�4^oO�u6t4�� F9���$�ܟ�ܳ����z�'�;E9}����(�����+����kV
����vV�ɢ��}���?�	�ۥ��Y@k>�n,m���1�����~�bK�5�����[b��֑�+�)�~C~��e|�/���:5��J�9-�#
l������Y��U�UZ�p��;��&v^F�g4���!_Y���,�=�`,}�aH��LDJiZ�H:�_���:���)E���t������͘�q�T�\� p��:g�,�"�Nvv+�C�^�~yV��ޢ���MM��:��~���3�a76�5��1�*���[� t�s�!�����z�J��2�~���}�Ea��j��c�S��O��k`���v�66� Ha³��E�=�'���#�I�����̀�Q��Oz�tJ_v�Q8h�x�)z���5K�� +��~Ր &&*v�PZy����:���e��R�0����`���|��Ef@�b��m�,;�6��4����BNqBnٙ�{�ɶ ]�J�!�BI�g��0sܢ�)�I�Ls{q�;��WNh���K$�����Ng�vD?����SD�ܧ�"ޖ��~�D�=Y�de�!��q,�+�oR�w$�t^ �VU4 ��I�����!����O#S��D�a���e��b#��z��^���*�o�N8٠��J��ߗ�{M�ڀ$�bصQ�Dp�����X�J<r���8�4"(�
sYi9*�")#���
��j+*��뚠~^罴e;��z��hD5erx���ܘ��1Gr��7�FL�;��Y����Jt�O�Cx�(��1.|���:ӑ���2��jnf��
�R�H�]��!�{�u_��֗��t̐�0c5��jM3G]��6��cV�,W ��x�ݘ��4���'�j�=:�u�N^_�u��8�h +���)%��Ҿ�I�ϑ�Of"�3 ���Ò�n.0u���Dp�,�c`�B�,>��v���5��]��<��V����G�����1f�tpn��_u�������6�^$�Z�'�M^�n��R�FU�i�B�E���0:Љ��K(��S��^�����5���;�ElX�>N����M�(3��벬��2�d�DՃ�Rݝ�T���� 1WE��f�"�講�Vg���������QSL�&�`X���lS�&"�##���w��o�μd҉��G)|9 ���u<6 j��?-lW?��� _�Y�`!��K��qf�d΍�kH>��2%m;W���,���Čh�B����zB����0��[�J���v�yi���t_�[�B�Q�ؔͫ�w_�u���!��Z�����l0'�n����~�O;rw�*Ҕu%�U<9�'Nn��G��0��̮&�ln�5�Whh��3X�]"Pg_�4�7�h�F]�=�t �|�w�n�����~��Թ�]cu%��q|��p��_l���|�i��A����x�h���'�4S��vܻ��[�"��s�|pZ�?`Uy�jZ��"��;�:�n��]�� ��-��e2���ӏ-�[c��&����z���7�5���S�eF{���C��|��p%�����QCG���-��:���\��ǿ���eMB���y.|�tJc���6�+7���a����PﮮU���V�uW	��(��9�� ��ۺ�'�(nV/�,�]	�_���MFL�\ߧ%`����(�ޢ�aN�[M1���F�2sR�Ak��6��I?��!ʖ�����8%r�h�H#�R��);y*����}���P<L(0H��&��#@����L;�W�� ��I'/�RA��[Ʀ!7Zn�?Mz��#�tj쫻aN��&�^��B��@�SF���^��DW��<&����Dկ��ǀm�����+FE�m�g�K��9�E 1����ey����ni�b�ں�s�Ѣ]бx�=��]��I���ޤ�g�BR,��Lv)�mD�~��B5#���b:�e3w�<s`�'[o�Ԩ�����օI���g�B�ɧJ��8ap�NM�b����<�̒!>��`��٠�!|����7V0׵��
z�ǅ�'�Q< ���
1L�����ߟ����#9����^����D�X��Q�|g��G�L?�e.<
�oC����^;�3�zq�_ʇ�Ȁ�� ���ޙ��P���Æ��5۪�#B�� g����iT�z����y�"�����R��:~B��2�C�d�m�ĝ�sN�p.L*���$D�!\}f��ދ!-߼�j���qMtǅ�}���o�anuCZ!�~�xO��2��.�q��WX==d��2�k#�"�d��.��>e5�E^&� ����yv����p��r�;00�E�%���r~�7��"fՎg�P��/2KaZ�����
x�j� �6��7[���=�\�3�t����Lz�ig
�;/��eG��vj���0o[�W�O?���7M5��U��B�>Z���ަ��lk]-Xx��u�i���+�C����:�9@=R0%�ȅka`�KT	ܶ��I�A��wJvF��Ζ�~*�7]5C���E9tU�U�q$v_�kV��]�{�OV����O�R�1��gDUd6����>
�{*d�nZ���u��¯�&E����#��ȶRp��ش� ޳�Pסx0hR	�{H�[4
UC�H�݊��55#滎��/�x��+U��)�(S��{��d����H���d.mҭz�l��4��B<��逗�H��d'z�#ϗ��Q,�
��O��]4�m��!"Q�7�a��D�������r�wmlZd߾��&����&��5�8����@#�Gɤ� e�7��Y���,H����;NK	ũ����@�,8�!�dr ��� �	�je�'��L%@M@tP�#j��c�Wo�˒����g�t�E��1���C�;Z����o��in�+K��$K���|쇷�RA��yC�N��{�8�،ƞ�Rt�k��q+��o*s����)��O(},ЛKm�x;z�^
���q|���z�y��>児?��F��wS$L�[�껻щ���l�����J�T�� nކ��22�=9�'�B'lA���;�&Jr��Q��pW�������!���!ϸ��y����3$`�e�b�=���zʩX�Wqh� �&z6@cv��J�r\C�D`�q��
���Qβi?<�GYw������Ô7�1
�-1F	�a��ո۟��-O@�ܤ���R�h]��ݘ�dנ�v ���a�>Z�1��_��u�so�A�eEU{�J 暋�����+;:(_X���#�U\�X��_�(�i����<�h�����X{�U�ې0�
�~�Uy8���G����fI����h|ȓG$�V0`M�H���lq��d	�����Gi�kX��\V���l(-ſo��W��S�b���	�N��ԩ�@���o��G
;:��.�s�>HF�IG�wc �_h;����^�<ɉ�L���h�^�����{�n�uA�/��8<�n%#s��b��臡d��&��'Lz
("�s�Z��7�40��^����p�<	�v�	�R�RP�MB�\T�7�>ݏ�&�E	4���t�I��r����4@�Q�|Y�e�`�qE���55bh�~� F;X�Y!4%ǓVș���x�$4���a�{�GW�S�eH�{Λ�2C��9���)=����xV�/�uJ�T!45 X/��֣Q��Z5�׋ӺѮ~�>u_�W{�HGT(59���,�^w�����=ܔ��2��hu��]9pz|2CkĮ~�� I��AF?N�xS�(@�5�420a֓���P����Yp��A��W�ps6i7ź�4��^w����$�K�fQY7�=ݰ���G:G3���<�,�6���R)��Aj�\�DZ���UZ��EhP����#f9I�f�TE����ex�0����P���@;�Z�d�p�uY̙�Y����mp���uM�xxO��4��tç"R�oH��g�8�`��g�~���?6!8A�F8u��ī&c��&i�4�h�N|�D�k��e{����rD�%��ٟrź`��%_EXQWw]�0�^��A4��ka�����$���!T|:N������y$?q �N�X;˚m��J�1SgY=N?`��`ƈRE�&Ѹ�R-!���2\;kXci���ı��~�KVA���`=F  i�b������/�T�*���2R��mcb�q(+"���`���ȎH����Ӑ�V(�ӆ�����Z�t.��m��'�è�6�c^�mԏE�|:?��q��و���OHUc��3��N�!�����v'e,�k���G��m�(�bʹ2�贽 ����Ay`T^Q��g
o�k$ �G�������>���ͽUy��`G��[a���0�g2/�[�n�h,7[�d�?`��sJ�'4�����l=��R��6Ĵ�{û�2p��g�1�,xH3{XsI�+�O��󤶍F�А�]}z	�Sk~
>8� q���!��^�
�+3�7�g�P�ά�
�)��S <,8����d�&C��Qsl���$����y�5�5嬍��-A� ����;��T����(��x��|q�T����m.~������}�eF�e,���>�f���a�:���iv$y�ًL@=w�Eog=@���Z@�����ޘ~�
/$,H����q�l$�'=�9\y�a�������Ym�G���