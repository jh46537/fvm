��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&���ˆ:��>��+�������u�ךF~��!�`X߇�&W���ғVu�:R�F�wRƊ����`O�뢢2c���f���03��s���d.��Аc2wT;Uə�4�D�ί�D%o �-?��*�-}EV�ҩAը]�щq��8#�N�.c��K��\ڇ�΁9�1�ar~����x+D�Tad*�F��ZB���UC��5s�I㙞cU�=�A3A������C\�i�*I(�$�P�e����� ºYW;�m���������Ӟ��2]%f�f'�߁|�;���� ǻ!8F���4C�u�j߶��SC
Gy���?�$-���K�%��Z���k����D�%�[�,S����U�t�^�1ʣm�Eيz򵆐��A��e����
�`m�}q�"���&I9�U��e��Ј�~&L� ���d,����%��}]��t��3F<c��/gC��բ���J��$s��5�2{:4����|u�T-�:תC�{�j�J�n�a̪P��?�R�$�	��tB+(Ro`K�//�Z�D�
��K@�|���q�s�lxL�5o��bݖZ��A�]�8�P�Y@���Y�7D���&6&D�0�uF�MN�h�o
=�C�7*������FU�P���Dۀ�Lp�`�e#�n�Y�����݌*b��i��B�W��<P�!wW�|���,,rT�	B\���]���k��;��td�>l��6h��?��f;p�،��3Ę�v�-��9�>��t[c��V�ұ�d�XL�J1:/S��\?Z�jx�)�I��$��4��E��91�`��<{���q'�q5.��=;�ױ�|OZ��c3.��S�g8�S[Hr���q��H���F����>F��f��t�f\�i���fZ��Oj�n�	X�ly�в��~ݤ�ѿHTtjZ/��W
}d��P�'P�y��`6����!~������tnJp�d������4@��g�;�V�C�H�-q�Sh5�*�L�'��1ps�.?�
��\U��_u��O"�ۼ�!� L�M�[#s_&C;�� �g�ofo��k����o�XV��D2�Y��:ct�H.;sbܳuj��<D�x
����q�� �4��zq�j�Y�X=�Ly��V�so%���>#jc�֒f�h��,�]���U�b{J�ei =���
_ey�g9�@�VW?P� �U��׆Η�vO|x���`���>��s#1W��rkG��pS�QB辥����@/�|\^$�byP�[�"4���U�%r���xa�*�p W)��6V��aw ���m���Y��//,��$:5	�ۏ�4W�r��d���ncOq ��f�=pT���m�Qꄃ=���a�y�Ѿ�����3�ى �S��1�[F�`�\-��Ȱ(��tm�!c��`����7irb S��pm�Մ` �O��'���e���|Ɨʔ6�]=h�*�T�P({��{�~�C<�h��}�~yb
+�<�Q�`�+[ҵ��,b��L�$* ,���֞e�z��Ҳ��L�N3e�C�U}�}��J��l��p6����5^oe����-�e�>��$C[�r��[6ʚ'{��aa�k�����:�1�S̉M�t��V!-�ʠ����U���'�&�X�A�|Č�ת�@Hh7��M]��٦�Z8���NGj��g����ӿ���5��_5���$�,^.�*� b���Ii����uE!�b �V���{"/{e��U���t`]^_��#<܉��)?5N!��[^�[*#o�7����'Q��P�a�|)K/�?}e6�I��� B�hL,��S�b� ���[���;J���T��E���Yȉx=��@{C|)4A}�H���zX���xJ.$���*���H��?�s���b�	��o�JG�3ˈ�Я@�9�z��vw�ӧcs^���������͋������L<
�Ϊ����-��.��*����&SQf�0��ߺĶ)�� �Q8�� �I�`���ꨳZ4E(�f���~�0�F*)}��2dD'��p��gn����̞��r�8�w�A>v��Q	���%��{����>_����j';T�UH �F��W�f�O���3�:�	�ޏL>w�u�G5�X��Em���?�K�Z�L�����c3�v>��wC��ը�b�ȶ�..\[���� p5�@��T�-����#���d�	�: f���R,��_�m��#��bLTd����{�c�H�����,�CF��q�s�Gy��B���A�����Xf�)���7�]^P���u6�7;+�*�3VeX簷V{)�JZ��/vǢ ��+�L���K�^��q���n��Y�Q��� `�����?l'e�+�%���_����R�J(��U�������hN���SI����Z�!��k��rfv��(�HN��LX�m��$K0c=�Pئ��S����C�����R��i"�G�(��2m:�
Ո����y�Ѻ�H�=�>LI7$5�C#�����5��@>��T�D{B��{�$6V?�����
��t��k����C̏nj6T�6i$�m㡼0ٙ�.>�BR�A|�˗��6�u��Q߱4��-w���3-�������K�����*�?�W��������K�����6e�B����4��pd�wI�u�`����׶��+-����]��GV����ϕ�/��"*�!4�Z���S���۶ټL��5r�mOQu ?����cf9$?�bf�����Cw9��e��!+��ߡx���Q�W�d��x��,�+@g}D�xB�E�6ݐ����9����D6�Co-~��[VRk����G ]��Q9��Kl�6��_��g�[���?���Ai�w�^rֽ
w;�l���T�3]�rh����$>��
�z��U��Dxʓ��D��P���m���(�<���&:������N&���D�˧�k8vR������k%FW��&����#K�O��9.�?^k(m�����+!:����)�9�M���Q��l�ҡ���jA�"���`J����k{ ���VE���$�/�������KW��L��`�d�c���{��mvx�)�n����+����&�)ߕM��=��{�S9'i��`�|nN@/���Au��$0�X����`��G��1��y�