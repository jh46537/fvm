��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��_)��%%�.��D�ֹʮ��������7@��=�y���fA-krT������&)���N)������&���8Ol.4��^�t�9��Ai�����q>��*�sv�_٪����qT������\��=�"�R2
�D��Y�$�c���]�c}��Ă",=�Dm�@ B�Ňm� �o�2����c��o9 c�)B�wy��~&�N"x��#�wE�>�J��$������% �YdT^�#���Ϫ	� � cY���A���Ѐ�w:� ��fg&�7���HE�(��L������7agzI�x�ZU��qo3���z�FĽ��%fy�'g�3�Nuq����R7l�}-P��xv���+n� #D�d��b�p�c%�������C��9^-G�w%��-e9I�G�g���|�9ғ�H_�<	�Q&����C�y�z��2�����(��j���տ��oQ�S����Bm�>�m�"���5{��� �U�^�QϮ��'֟��
g����D-AR�Ə�d8�z<z�X`��a�����8�L��e����=�þ��׍��_� ���8x/�(-!d��;3;1��r���}2/Yx1��4�{v�(��&����Kl���a�� �AV\�� 4�x�4�DT��sj'h/��]��Xc�M��
�l/N��O�wr�d3��)��p��5�CCk4�˵�и�惭�m�tԋ��M���o�JWJ�~R�H�k���`�b�(�o���u&z���]���Ȫ`�Y*�r!�,�.� )��L��miUvg�r�I��hu�e�b(�q�}��Q��ө�
(���xe��彵0�rh
���cvl�����?ù�1�M���qK|x���c�P�]�h�ZUҁ���i��7՛Ջ�j��)BD_�#S%�I6�N�*���O��Y��u=�eP��F���o��+$.g���kN�E��%g�AV��@�c��}��W� jUS\�y2_EӒ:Ku��r
=��c����ݹ��=�;6n�A{��;�R����WF�\�7Ɯ� �����L
S#R=5���La��Qb���~�ܕ�йQ�!��)�Uo��IQˌb��+ f��$\�4�qv�Z���40��tt,�0#�3l�mra�^�$6�X���n���ſZ�=�ń��5}�t��"9X��#hz,����受C�]�T��p�%ZѸ����;�nW�ˉ���q��+nO���B,Z<0�P
Ay½�\?H�f�.ug�$z�(
�������&���Rx�/�{��s�t�]�8a�=�VXj��GK�ܩ@;�4���rOkB9�������j
|����:J��JԀ�5%4����(	��w�銆�0�t0j�5U����=��>V���qU�}�'�F�v�Q���w��zE��Y�@{� T���T��֓���FB��^�9�E�#�C��ѥ���1�_�5�g�x�+�9X���}��$�Aʫ��g���q �*���zu�ǰ����m=G�Z�
&ǌo��b�GFZ(�I�Ehz@LR�� +&Δ�R�P̖�<()LRWS��e�O�˫m��2�]D��9�D�:k����j$���zYADȻ��׬h�08{����BG~*�wܗ t;�oj9��Q@o׬����p�!;�����ޔ���d$A�Z���4'r�����,e��u�Eb�	��S>��`�����os�Q�+w&cK>W��sח-�j$Ȗ.����
2���*O�������q�'��6���e���S����J�YR�)h�>�]Y�z�㾅�Ħ|G=B�4zY��%ܡj]P�1��c�l|�����9�	���N��%)~�tEA����|�"��~B=?�k�HI>m�� pk�c���5e۱�>T�x�R��MĖ|���w��x`�^ϫIE���H�S�ᄂ��M,h�|��\
0%)�}v�q|4b�J�u���vC��*A�t�DN<���ā�!-m�^�#�/cˡ�^j�5������Ná���1"$�=��UT#P�>x�eL�^�E,X�� ��e%���U�Ӳd%q�oAN��u}�A�MS�@�R��N���� �F���P_pS.�16X��ޝQ�n�l��X�G����<�(z�I���^�X�@�9`��Q�a��6���oժ�D�3���I�Y0��� �ߎc�:�_���xݾ���!+N�Uf�%E�W����L�ms(:+j��֍��Mtlv�r�W{Wb���f���1�^��b�'`�������u�ٰ8���졔�ϗNJHJ����jx���~���jd@8�1$ �`��TȪ�佒�Ea!�/t'���b/��6oyg`�����d��[Nd8�P���[d��ĺj�%���$��x��{�@�l��������	,�'#�;�U���iθ.�uB�HYHWԍ���x�ׅ�Fk�ѥ��:����ܺTB��@K���M���Y�-{)��I ���0�ݩ��+�Tp�l���uzBȇ��`0�V�y�:��.�����j�ʔ�������/G��V����K4��ϴ}`N���b�m�m���/#'ā���E���Z�O	%�`n�$��g��O7&G�2d��4{�u>�a�JE���U��e��F�����?/W�;�Ǩ�0o\+�5�K���B ~-���)-�D���[���_ZX	e�xRc�����.��r
��ߘ�Т����(�)5�Y�C�R�;��4y\g��,(��H\ɴ(`e��g��9$)Lѝ�(�/^�(���b�w�B�4�qy���:��{Bw�e�(i��`����xI��`��(����M��_x����X�c��W
���tcX�j�E1z�,+�ɤ7>�dN� �t��G�F�����h��G*��A-E9HV���m�fu�}r퀄T�cWаg���]�~���x��i��M
�����s�B��}��&�{�z���\ҿ��hk:B["W���M� �����Yg2y������0�>2�$O�ޕ۬-��-z��r�����B�Dc:�=N�Ͷ
q�^��ڑн0�t�����U�[��s�^�{.5j���&�;7�l�
�U�b٤E*Hy�'��v��:�{�~5�<��9��[��R�3��X�1�	��RQN�>2�3R��=~t 
�R9�P�{I.=:AC�W�;��4 �",]��z�A�2�;�{�
���)�A�\a���6PJ+wG���}�`�.T���ZQ�V��������k��ƞ��S���=�$�Z�����P,���(tL����Jw��]��gƻ�(ܕq࢓����v=�c��~��.����T�	sAj�;}�$"���B���������II�$Ϧ�2�Ze����8���QƌE�v/�2]�� Br�M����[�&��{�U�^���9�� ׅp�'g4�d=����\x��	��/E�����g�9��u���X�s�N=g!�#biƋpC|V\)C�2֚2=9yM�	}�A/\s��8�5�Ys���~�:���{}�C>q�=�ױ���?y_��ʹ�-5��{�b���%�K��AV{6��8/�&i�2Yf�l!��u�e)t�@o�v����rQd�`=MB:���L���]i�b��h'?�i��!���j2)3	_<����)�����@s���R8hAz!H��4�l%t�!�R�̦�LbV�A}#�Ά���o��HP��9��Ի⯤���"M-���.�^�
��R<�G�����C~M�X��WX���衜�܏U��,�^�t������:S�JC�>M ��j�s��� �I�:��K]�3aFqR��}����
�(�'�*�QN��s���N��d;��sD��|�g}�"�j���OO���s%�U��3 �K�q�ׅ.X�[�IPb]���_Wq�M�����U�?_�A
��e�{�7:�������O�Y^:1L��p�bRq)[�C����oY����,g�i����Yʦ�ƙ�7��� ��g<q=o�I��"�5��3[*��F���ulm�-|D��d��噶!s�~K؂����߻�n�X�Z��i��.*(x]�Q�+�+��g�p��d<;tq�|J��e%|&���w�D�x�_O��Z��Ļ_��CyIBrP$h���IBI{~��tr�鞁�B�3�x�5���2�Sk4j�6��ݸ�t�n$�:��ܼ�N��n�8�����"��;�����B~�߯T��ӵM)^�z���߿��=�#Y�.y���lj�i|��h�hZ���`"I���H>���4�j�/���Py��G!�)v���lL�p�Ѓx���(����e*�N�`��"��	��tl���&����8&�N�7H�EZȅ�[�ma$��XI'�A�!�J&�ۏk-��=��V�����a��:�L�^t@;��W^�ar�F�����`���
cV�g���U��j��^'��9Ĝ{��i�����9zf�2H�n�^ɕ��tQ���ޣ��Ȑ��s��
�D
���tpr�5��3��u$��s��������N��&�i��<�Wj+���Q#Cg��YO�S�_����7�S�_�2�Y���E��$��� w�r����������aa�e'\��i��`)眆�E� ��@�X������8^�c�@�nj=�&N2ߍò"ֳA��*<E6�MN�V�3��%3]�[W�V�Ld�J���05hq�i�J���	����5q���kn�mF%��r�sR��dL�8�*Q�z�,�2w���fJ� {�~�y�i��K��+�]���H�y�`���>�1ƗͿRu,��LGL�~�I�0m|�����u�O48�'���8N4E��"9��ul����Llw�Q�555�^��:����h���� �>�[c�`i�TjZ?���v6�m5�P!5<f��fB�_�@Z�@*�m������s��[w�>�gJLܓLt��#�*@��G^\��.���~�ViQ.�xe?K�2��zrU����C@�u�'���}�~� ����)U�fۣ�� �-�kޫp�U�>�xn��}�� n�
4��<���J�|Z��F���T(��zF��l�qg����BWE(R�b�>]��k���bBa�+�����w��:���#/�fLQy���<M� ���J˔�5>z��<G&ؠ�=$��i��Y9��5���B��d�+�� |^/Ook&���JoX"5�Q4�L�����8�(�.$,��ZuŞ��<�8)�.��g���?
gӓ�H��t� �jC][��*0_����稀qt@vo.u��}]�lZ[�]'�+bMO�p����Ð��Wi{�b����6$�N�NmYJ�Ǣ�m�>�(�+��ӂ=�0�ƾn�Z�3�u �uy�M@>57t�t�W�$��Fi�K!�u3���լ��"�R����ooN�F�@죴ę� Nٲ�����_��{eE\��}�J/���[ԁ��:ت�s��ƛ*�	��#���)�E��M�M!v�<}#�����9�'��su�=����wi�=ߊ���}~C����<��[��~.KmdA\�y���ˇ���t�{�V��qVT�2j��˖t"�~Q�Mt�T������1�5g*��;p��ޔ{(�)I�����2u�"48X�A�3z(g�v�Hε�!@�.��`��g�b�{4 ����)oJ��?�^_r�����������;��{ǲ�,6t��O��ӕ-���o>�<��P ?i�"�J�bO�ܒ��C[Ä@\좴�oi�g6�`n ��3>�M�ܒb��a -�$Z�4���J�'�^@w�F�r�vb��!�	*	��=��4���g�����u��e:�;�;.X!��`�QL�{;�X4Xo����Z�6q�}�����A*��Ծg�:��T��[���=�/>�����;d��:���F�#���|X��
5�o���U#@�#c���w��#�Iء��팎705DD�)H�ĕ4�h[ǊzOE�p�Be�T1��j����0|�����0�X �9����t&ђm���FF�u8:t��L8�GZQ`�[��8��	�˃�acs��kS�z��X��B�J�a�^��/�O�J���ۢ�%a�E�պ ��%�������GTib�u��D��g�X2Q�Vy��ɔ,%��@^���J}M�R�qE�rI��|Y��u�|�P9�HM$��C}68�/�u�����+ B�񭮚u��B}l��>)C���+4Q�X,Ssq�(��!+,N_-Ѵ��VT��.��Z�J�-����C�Y���*���/�[�\�y咈qk4w�7I�����<�����(�	���Q��s:��N��s����2�Q+hg C��k}[.G>w�<�с�>>�����8gfJűW�HK�Qt�5��B�K���	����$#�ɝcE�i2�t^�@+�;D�,C�+�D�e��YFIG��P/����� �P����mv�Z|��{�B��ɀ�M���O.�����/����%�DFB�4M
�B�T%:�����8P�r�/ed5���C' ��m;2a� �[��	p�V�ˌ1������s��$�7�����+��Kp&��;2��z�o �P��y<*���n��G%�1h���.�#$��b�5��¬Ϛ���&2�����qͰi�H?~σh3�]��X%���6���M�n�N�;_�{�t���U�}�6ꠙ�?����۸��K4�{
�ܔ��npCt�(����eB�eQ~z7���Y'6Uv.R�~N���z�0/e�3��^R�UF��6Ϭ�y����,>���x��	�Ne�E֥��@��|,�f�$�R�
d�eq�{�O�63���E(��#=��^�_��G_�SN5� �.o����8��ʪ�F��d�ZT�)G���Ń�����qkXׂS(�@dˏ.u�D�����+.�-e�u���m�_�x��W?�4$�|�څc0/��m�|�P@��q�$�_�u�L;2��:;����<+(n�bB$�j��X��;\�� Yü]��/���tV-}n�����9s�
��I�L$i�?A��$����S�n�S���5��N��*�ʒ�P1Z9TN� 5��;aRIq�LC�|(��t�-����z諄&F�<�12���YsӇgG��i�?�怜�
�Q4,��Ʈv�}L�S�.2�!J:�=ވp�U{��*���>P����.\�18T�:����R�\ib1�)oö����\؀�����WX��G�:��p��k��,�$���2����6h������H�U��ỿ�.?��<[֕!�󞲔�����x	�
�D=��� Ԝ��+١L���y�٩j�~�ElE��[�ܑ���9ZwExs�m�|��������l[��Rt�q4s���n�5ݐ�m�FV0���'�E��^�BaA�k�$׾��/ݬ�	���=�6&�	��������fA�3 ��׋�	+8֝��J+i΀G�J�4g@D�N��k�b�憮���X�����D��.3Q��:M�S��� �g�wķ��^�~��)�6uY(S����
&�_�1�)Ţ��H'!��ӌ�Y�)�C���S� �qLU�6���!X�P�n�g�Y.{&H���V��x�]3����-��鏆@YI�)��Xlô�킚����[��`�Qrā�M�@���~b��xl}߈6�8�+����f�gJ2����S�N܆���۲��]Vw����Ƣ|K Jl�t'+�sɰu3\W�0��]ڸ�&1�ݵ?J`h�(D���H���E˄a�q�}{�~I;����� _���b�/w[<�h�f����ⰪYyf윁����h^����5�G7�҅�uP�+�=�?�ӎ���b)�Y���zב��k��q�+���S<:J�2S�����BE{�x8P������k��uM������������ �@��;H\�C�f��>lz(�(��Ӌ���or��Eob�2g�.��YD27	N�d�������G�5"����I؜��Vpr��ZU [�a�,G^�v�n��[��u��#�������BAV�,m+N^�X�pE
H��G(-��[���pX��z�z�ދ�7X��7/
��D5�]����\]>����Rd�͏j㉃�߲������"�	���@��lX<�Vrb���������qG���_�]3�;��;j��!�3ôM�?�BRJC���.�q ������Ұ�9� ��R��k^��5�I�V�H��o�TQ��?� r����}
�aԢ�G���L��7wxH��p�|>����ջ����a�P�t��+��[Y[\��0`l�R�%�"R����K٫�f��V�L9.,ה�.{�7���䓱�:=��;TU[i�'Ӌ��Nt���}[��E�٨�(�G��bX�s7*�V���O1�f��^�3�Ҙy�x@�_I�x�b�Bq	XZ�wb����:������5�(��ك��������"��f��T+��;r|*���)�6���t�.�Xލ�Ñ>�qĂҜM�I�~mnwg�Z��B��O��t�3 ��ϯ*V�M�SJ*u��U.��<�XL
�X�ͼ��H�d�Z4�y����y�M�4�`�O�
���<C1YvŕjW����/�=F\�6�if@J����qĔ<l	l�3��G�	�)w��cg�G5��Xo��/�!dq��I�?ME�����)� ��]}D\��ϴN�Q{�w��s���j��x�O���!C����d��8sdM$Tq迖[��A,Zɝ��Q�@��^�80C�>��V�=�k�,Z�k��O�C}��[��8��z�i_�Y��'k�M�n���SL.h��KROЂ?>�~2��H�?`�[�<�.����MT��h����!��>�P:�L�L�n�"0w�6�C )�%��q���6����I���>�޴���lm�����7qi�H�_ ��L��JL�Uez��b�Ó,}~	�Ά�Ϸ^5�Op��ƌ�$��=p48%7rw��V�+�t�_��-<6�����ph(V`�Iz���U�l����2Z�UƟ�zA'&;%K�[���K��"0dT#�B����=zN�1\�R�6`j.Q[K�j�n�氞�.��\�a"e'��!�C] ���2���G�u�I��P6!�.2�+�3�,6����=T�h"�����^�|�1a(��WR�.��H�U?�&�6�"@hX��R#;#$ W�E��Z<P��W���M�DךC�/,��L���~��y���;����Њ��<��S�����-�i����{׵��[_6X�)��2uBx3�KB��VD����,/]�����B�cd�OQ7���QWB>���y��тgxV�g��ka����y�Ja���V�y�#�h)Q	� ���q�n�w1�
��|d�T��Rอ�� ����"z�Д�z;+�ڪ/UE��e���#W5�),B�T�~���ƴ	���	.���`V��)T�HhG���$�6��p�o������:y�j��R��c5����t��+�M���ҵ�X�Jg^�Vd�n�c��8[�3N�	,x(��Δ4Cd��<&�x�t&���J��8�Q����%)�i�^��z�[
�$U9�|r�S�f�n���h����G�Ra-7)�{h����p���0��ߓ��W��Q���?#�������p$���t
�Q�6�.� �{�6v|��u` �k�6U[/�Yl��Wl0
f#\�����G��r�p1��8Yҩ3�N?�A���_�z��N:�>�3}��'�2���Q�Ψ��u�}���/�i�־}����h�dB=�S���)(�}��T)�$:c�[���>}R�*�1�%:����d�%����C�f�*)M���6!.w�A
&��T��Q�*Q#��wh�T+1�O��O�Š|*A�P��l�U���W�B,ܜ͵�K��z��Ni�}�GEP��[d���������&}��׀��)&XO�ofs�؏�����;�����Rdc�b2� mrWO] ��su�%�[<��������k�2�>�.^I�,�R�KF#H��E�����s�)a6��Z]8�+�0�������b��=�B��o�����|�k9���1]!��qTݽ�F��S�V��5��NY,��d[�ۇ��]�ڻJ��(�';�(���ϛ@���� ��Fh$���cP�o/xN+�(�A���g|9G���:�����tAJ�+���G*f�_�\բ�,z��>h$�������&_�n�n�k�K�f/��Sm$���1������+8;Ȝ��/T>]�> �k �^#H�=�zo�>ldeZh8�!l?k/�n����'�( >����I)��W�ݲ|?dPr��ē�ܡ�a��Z0Ԋ<��jQ~g���S�VR�b���Sn�����|'�(ԯ��N���t���>\s��@}��=đ	�=73v��2��<����2Cg@��� �I�C���(�zUKzo3��\�bFp��c;�24�z�PzEa9K諈X�H����6�?7�N�Z���|e�G���1�_��R~�^��0ԻG��%VO�*n\0�K���z����O�����ߍ�wo�<0�5���4�'��ś�8�?Z���Y¡����<x�ӓۮۖ�,��?�� E$��j���/�5�ϰ�0��Z�̧��2ʕ\'#��m$��^��.|Vb�\P g�=l�O2	{��
��2�.�a�����6���qE��l����ςHI ��n���Q�-���t�s�5�w�z�/ә#��;�P�-�
E��P-6�Nԯ�uQX?��U�H��R�i&�v-EtJ�sh˕=� ��mN�WDxh�aB=8\���2��!����ǲ�e���3�"�:��yt��3?����&�`t�/�qA�o���װIүK���%7������x<���eL^�x?�����*컯e�ѷ�6 ?/V��!7����E�',oB�hc����j��ڋ^���s8�^��Y��|V�ū��������%��&���	�4Q�.�F�[2�1�ӿ�h7lG��P�q��;H��}8��j���a�~Yw�p�`'#P����o�L�`��^�)خ\��UEcXs��R��~�j��z,\�FP�T;�*��~CѸԷ9YS;�B������F�R��@�ue6�l���D��l	[l�%1�[W��ŰkT�䒔�P��F5�>մ;��M�E�������Mx���W�K�
���V���BM6�H>L�9����S�;��;�q�~��D��VA�*@w���O�bkwg�o}��˼��}�4�x @��kAC.A�����$s��!)՞�42���o����?�><t����f�.x�A)#V�� '�s�Y�4=d(XN�7�bNP�t��2��L>��w0!�1��M:%���)�m��ȝ�
�4ɥI�^`��Z�֍�)��?��.Yos΀�w
�8����`{���wd�紌�!PC9M΀�~��?�C�K'2z��щP:�t��;�	�O�\����9};`6����d@��~ �v�럍�����*9x�2v9J'<��s4g��ֈ����eMʕE`�m
'��g.�*����!�v���e@�1���.W��R�#�1��A9�NV�jY�=�U��=����LI�~u�`!�^��$5~�]P�+'���ܳ��H�s,��K�t��Ì����q|/GR�!�&�k6��`vm1I�N���衘a?]wI�!�>��W��&X�|^��A�	�Ӗ/7n����</��NC�8=��7��Ü���v�j�5~mU�D�jB���fz��(w<�;���e��,~��K���y�M�f�	?�a�PR�i�8����2�4���[jOp�(d��j��X@���4Ѡ׺W �e�� ɛ�c� *Og'��R��=%*����`P�o���ln@q����]���8��&0���s��]�Pe��͉ht�-Kzdd2[BGHB�d���I���W�<�D$$�Ⱥ%�\a�$�M�I����*�萇v��w<Iձ4��d��ƴ[g���xw���Q����{F�@G�Z�iLr�N��h{��;��4�C	��s9�k��$�Ձ����k�n�1:�B[:�%(O1�rP�Q@(e�q�@>R�j���N�U��nL��"}�6
�ĕ�Im�M?��?��_rA�e3m�P�]?�l�\z���v;n	Y�P��ɂ��b��ߠp�&�+�5�[�ҏ6=@ �)>A���S�ӹ�ؓ�����t1ѝ�	~�ٝoS̃OD�-VG4�d�M��B.�Q{��H0���9�����9`��&��C�y�4�Ci.�bѐt��ʏ[���7u��l�%��Q`2��}����d+�����4)=�ç�.��+j+ *��Z���)�YQ��$��aR��>�
��o{�j�K���P\y�b��> ��}�|k��w4������''F5�?��_�&z���7�� 	�Vjs~�"�ckZ. 䀟���u�Ϋ�����%����M\I�!�6��7ds7�-UJ��'�M(rI��:̟b%��Y3��i�W�z�F���<鎌Ro�cV����Pb��\�Ln�p,W��`��p#���vpN5X��_�O�Ox~,k�:d���f )M,����J��Т��[Ո]^�O��L�G�˓}�~j%C���b]�Q�̼�y�!���_Xv�Ә�9-Cl��/:Pwh*��І�WDh������;��3�Gr�{ �4+'z��J�P99�k�\g���I�P	�0�,�K�]j
RL�|̭5���ˍc7W%\����ܥ�+�	zd�m���|Q�C\�N��G��,�ա���#�͚�Rկ��X�Rn�Bշ��c.�ex���+Pܚ�K�p_��0s+�������fЉ�.P���!@",Q��3+`��3�#3cM�j;Ȕi@�\{�zS��˺��ʐd�T�̎�g)fA2�,��*����,���s�+.����v�L�/��~R�� Ij�X�$|�˶��B=����>$�y���m��xz�Ђ��l�u���ԉ	!A���^9���#���{Sc*e��{}��|ɵ����R'w���CW��ob�h��o%-ï���kk���bj,[�/��[�"ơ�����H^Z _��N�3 N�����tvR�6�����I�FH9,:��ĝXQ�Fk����"�тj�)fF�6��n���h:��:5tF�̸�2�� |�qt��UQy{K�����3E'�<��)'�^���8aԳԿ��NVA�[mj�ĸ��?���[�e�ϳy�$���'8cъ�~G��,*�_n��a�$\e��%5��񟌺3���`;#x�J��*v�(b�x�Qq�^�����)�=@,ؼ�����g���T�9�۬Z�t-~!�N�.�\t��[�E�E��Ձ&�2��<9'�&T���p���C���_]��
�y����e�fa!J�'@���%� �AoQ\�@���zf����׆� W�4���el�㳷ED��5]5�st��������Y͵ߞA���eVF��B�7=��UNF�[^��<�Cb!_�vט$w��G��3+]"\"��u[Ҁ�UO����3*�T��VZb?��W�\4�'od@(;���H��$n1�����%y���a���cDYF�#��"u�_C_�[$4-�?��*9��dK�ӏR�XH�~ܟ��][c���)x�7�l<�/�Hdo4�W��*�_�kwGNsmA�i�]fhJ�h��(4o!��o$�����e%C�۴��0���9�p��5Yz7-��Yq7m�tj(�U�����~r��ƅ��{��Hô�W����D�me��
�I�k]%<l�[N.c�l��ð�ZJ��8�9�L��pʄ��dT�k@�f"���60g�/�a���$W�g���gї>aEi���|�XY�HnnA�bKd��˸�R�axA�t%kCu�*!��\�î�� ���2v<��E�-3m&B�~)�Z��->c<�!�d��!���?M�6<���jZU{������P�&�<���N|����\�|)��R>��a���À'�{?�}�g�H������S�̜|X6�}������kO�{B�M�Zn [ăo��	+���Q��(	���*I���,�B薖�IC)�|�av����et��W���I�V�s�o�).�:��8ﭝPh$Y3ڠ:�诠:�[;&G�
��0>$���0Q
��~���ʧ4�_t'Icz�bΜ�������H�6ˠt꣑����R��/�O-:*܅��ぞ#��r�Ψ�h#C��5#�+tO2�׏y�(
�5�kYl�c�8c\Q#`�#�Y�bk  ���N06(�W��rvz%ĭ�}�1B�R���n	����v�8i-tkv���ǖ�������`L�{�a�FiW0�q��ˁ↚����Twjᤶ� ̷��$v�|Ɣs�n(8bm���h�h��9ZR]OJ���v�߽�D4�uNݓ�I��/��"���s+k�AT�gD�y��VajeJ�ݣ��M��k�=#���0k�n�0�S������c$mpf"�%����w��v��D�2z(G�������7!�q\s|�[�A�6�ש�u��]��q�@��W���>���B�!v|pdrmIi��V�ԑN��j˥Ͳ5V��	��_�����z��紀�tuм*.ak�<{�F��Co�'��{�֒n"e�����,>O�I˶��$�[�D˱D�}�S8�ꆑ�T�C���6k Ĳ��FB^��IU�0
���m���"�:J2t��w�f��=�(��X���[����O��j����M�c�Id(�?�xz��Z�]d���V�Jә|)��;�Y."� ��m_�D�4ۥL[���(h�R8ٕn��X���V�ZR#��		i"+O���СM2����k OSQ��Wi�2g��zl����`�Y�6�Ƒ�1�4^�B�%0�.T~F�*�����kMX�)���ĩ��0��@�k�࠳B����0N�E,^�J�V���9;»Wm�m����5���6*�xS���!~pC&>�,���o�hK)�޽.L�m�c|�T�I��p~�q��a%��k�\r��)�1JJ���}�	����z9�1�K���"rH,�Hr�@kڐ҅V���� �e4t�N�m�Rv{ ��8	/��wݨTYOg3�K&���~���QfVu%J�t����N'�$.J{�#~��a�/1���/�E麶��Ϭ�.Z��6�;4�"��ԡ_8B���(M����}�֤>~��t�%�s}�4l�t���C�0�Q�{w�N��<��xTK�;�1^ZKzJ�i�+��x�H�E�ʽ� �V�WU�(�n�MCh�A��Y}.5�2YVn����e6mR��mحr-*E.5/���5\9^q���).�M�y
�@ ���Mhٸޡ��pަui�7pN� B��p��1 ��B��M�z��-��n�I|����L���uk����\LyR<�*2�+Äp�KZ%����jy?{�U?��L��}���jvj/a6�y��M�4ю1��{��8$q����^�HwͶ��22���#��:�-����8}X�t�����xE80-QZD�>�Q(���s��`��
[��F����Ƕ�p��C�$�4������&Q�״x�Ve4m\]1:N�L��L��89r���$���yi�=�O�����4�dX���.�䮔�L�G�Su@^�Ϝ
v�c�ZgܶP����Ķ�}�펬�<�\&0�����S+��н̦���-:����^�ױV���`�2��T8���ǙT��ǌ<bQ`gD����e:�k�cu�В�m����o��?d]�&�e��@��YTJ�mv��CA�k����f��acI=T˪0���	���-��6�&�����Ԁ����N�]�Z/��z�j[���C�;�}����q]Ϙ�4��q�IcȰ��"��l�ۈ�N����FO�u+�s�1nk�@E��eo\,΅-τ�)[�c���҃�k�U����t0�p���8�g���0D����>f�.ϒو?�(3|��'�yն�6�p��g`���
��S{�G��"�W�/#4��R�������o�l��w�j�O:�I��M��c?�~*���oV���Q
��:���y�!�m��6���.T��>I��?`�J�j�6hԟ�����3��$�=+w�g2K���=ҋ�-�a^
� N����$��cp��-?�#vp���%�F:��UI�wې�]���cg-C*Ib���BI�2��s��lQ7`3z�ư�@MB�lg�m�7v�D̶�]��\������d͸�"#Z-����C��W<i�<۷|)
�G��v|Ӏ�[|Й�a�>���y��vY+D���4�	t~��;�k��dy7�5�[��Ѭ��,O$���%v�7�CEQ��[��x��zQʌ�s	�n���f���3R��>���L�q�[d��3H6���`����J=���HN��`!֟E�Q�����mz�rz��G_��*����j����0�&t���	:G�j��)y�E�2��{f83��჋��(,��"1�&bd,���f襲����޼R�\s,��ԁ��lY7�3��'�7
�l��*D����!�z�|UŘ�Y�s6D?oI>:b���-�H�!Zl}'����hʱ'v���, ����w���س�P�v�.En�o�wŠ���'���^kp��>��8�n=�W��:^�'נ��yo���ຄ��6��c8B�p�:���g�7�` �ю7�{@�90�O����5ڬ�	�q��v��H0Hd��>���)g'^�~Y��T:J�)>�:�߉�?`��ox�T7J�5�],WOs;���Z�����=s<]W/�Sx�/�WQ�q�A�	��)5�f�{�$�`�&Z��������G�d�wS�����im��3u�PF���@��=��<Wo���t��
3e��Ij
����o��ƛV����2���y�9�?�;-0�Bۘ�k�CΜ ���ie��D5�PG���B�dE�	�호��g�b6���9k��>����c�_q�&�O�T����yC��3oӔ���
�7��uy�~�=��q����1o��TE���&�ۡEQ�_�TS��}%�g\���I�4Z��f�;�����.p�A�0̉�޸PU�jZ�u)`PXXC�P�+y���M�cl� �K�u�A��t+�YM	���������e�K�������ف���\.�#�.���'*p}��O~�M��%{�:�9@�z�j�=g9��ٚd��֤��l�2&�3�=_��FPk�D�Pt�GVߡ���j�j?k�N�GE���?@#��|P!6ſO����T��'����z^����zR��)��Yo$d^Я9I��l6X~����r)�4U��vz��,li
��Th��*�s#�鉚D�х���zk٧��<��r7؍>i��S':���<2�<�,�ZhO,t��8;�RK9n�J��k׶�����!�#�ը�������}��&��T[�����,\;�ߏ����-�*J�iXԎED�	�Og���۫�r�F|/����7���x/���`�����;�Y������NL��s��-nu�����?�S��1�R��D�� �*�t/����d������<7b�RDUD���Q�Z �����O/o��`���0�M��hBг>��oͿ�j}�K�yJƋL�����n�~���*�(D�y��0���8T��)!��!��`˼̗+��T O��#������x�D���z�,�`V jC���ô2�1��������@b^��uXJ����x݊�����#z���2�f�Nz� ԃ���m�cj�;��W9ҡ�A����la�5i����6K�EaT�������P;,n���S�L��H��c�vd�[�|�)�w+�$E|�Q:����d.�_[;�3�Oӄ�}3�ˣ�S��r�̣���O�須p��\����2��6�j�H�|4���c �ʇ��,˔2+��S�h����"�x����v�Z��{M-��"�ı
B��f-���T&�D�)�o�7c���]vT	us�o�+���_}Դ�ҍ��h���>�ě���NRgR�]�L���������_AH�XQf��5���1y��W�z�G�ߍ���S�nK`�P����x�͋�i7��CIg�/�;p�� )��<=���F�l���+�
��|�ҝ��%�;$�ʝʿX\ҝ@��p�%�?���ݍ�{*���!P�S���BA#�_��` ^����x��E�����	�\3j�qT��!?�-QJ�v����u.���T��M��uf�a�U�����a�U�n,��0�hF0~�#0��[�{R{�W̑���:�KZ�Bf��,��tO��dX@A��)��������Un���55�	�YXԲ��]k��$��e~c�s/�����.�"�L��zJ��i����pk1 �D�|9}�p��1i���ԩ>2n8(�l�[�U���+�>vݻ�����o/a��V���s�=�mEB&ʲ�@�o����^Ό$)D��� S	Z3��%~��	�1�KKW4s�d�2$�ʧ�{�,�����n�.�E�͝S$"��=z"���,�o�( �$��I#�Y����v���fJ$W�u�,��]P�8s?�j�f�I�I�+5hO�Y���4�
�+��W;+6� ��y�3�0a�����6�ü���
�G�̪L��M�eJ�v^/�(ޡ.�~Ջ���_{6���w�bb�'�U�B��Cx�CY��G�M��]��VռKo�4F=�_���G��).��(�C�:��Slr��������`��l�)�g�������ݰJ[�����&��XWY�������o�KY;�.k�_�f� k��'0�B��q�9"��o����8UP;�j�jl�����3ͦ|P�,lm��\g��3�ES�����'�]�W�Z�y�q����O����߹��L;���i�4 �D)[knKy Jſ���E�xr-�
ԧ-���]���r��^�whk[]p���>	t���TQ���=�B%GgW��(T8]J6rYA����b�g�(v+�,ִ�Z@"��qäL�QК� !��Bh���J����G��*�b
��2�⫸*�[���刖��<e��{�@R#�)�x�o*��|è��{|�f$}QE�B��h�k�n&Zga?3�W^�Lo�9]�[�f�'��H���5l�~�[�v���DZHԍSj�5s��[Ir�H�z�}�Ld�iăq≊JVZ��hz�ZJ�L��(��X�O�y��`�v�K/vs�|�5(囁(����*����eyA�R�d�B�`��y�xԤ:�����G<'��FY�]����(^���3������ �!t]�̋DY����,nŗ4���T���ύ-ɠOs��tzA��m*����o���B]��=���sE4X�Ug�!<�ԧ�JI��o��pOoǥA�P%m�jF��E�8+�y,����b����	W�i�ھړ�	��58��.�L��19Q]��l�#�5Eh���$����ʤ3�pn\َA!1zm�J�\�+u�-po{^�p�`��@� c����75�\]>���0�Bh����
�6��kٴ���g�R�Z1O+iT��+o��XĮ��i�ٸ�/�V/�@X��ތ�ƉX.P�U�����JMy�zx�6�1��b���C?�1�*����l�O�݌½tŻ��C���esZ����4}�]p�>2
xb}�*�6��j��-��a���n_�E�ih1���&#^`�@t�l%�<"iY$�wr��Z&IT���Z�wc�;]�d'r�<���S@���j������zd.��Jר�T���S'_]u5�L>�����p�gS���#�KR�(n�6��+m�]C���0>3�?x���B�X>@ZT��x��>���n�x�n�yYVh.f��j�O���׮6B� %M�;�T8�kDp�]x�3N�j'�8��B���HJy�m����yS2���&dZmL���/N8��a�uX'�	��\���E���cs�<'��Q��<
@�?~�k��ʷ ��rS�J;��۾�-b��YsPX@�}�$��C����Ɠ���	O?�zɤ�U�(`Z�0��>\�.�Y�ѝ������(�g�M�X雍-��0�\b��pJx�+�ؚ�I���l�․׉2n��^�?(��ǧ-�������0*Vdj;��r��/�U����}�
�j*EM��ZA�a�������_Y���'�`0k���b�vV�����yħ����dr��H�p���T2����>%��yVO��@�rk9EY<���LŞ�x�eK�?%b@+Tgoz9��ƭ�&�����|��f8���4_td��g�«b^�l��c�N�);+�̀Ѭs,�(\H�l��/8ˤ�X^��'�=�o%�!�X����-���T�����|M�J�m�b���3g�ҥ�8�S½�9;AH�f��q�88)3Snz�4�պq�j�e�9>JOJ����]���?rxm�5J/��$�����ۉ��+U� _g����h�'�P�0��K|�*/B���3鶎&��u�m��8D�}ծk���J]|�?�
C��u{����'��]�TY�W���_fP�����0.�u��"���+2�`�\����K�)�*���U����%�U����z.cJ�OE�}�~��Ip�M}��;0���t�˖U����H�)���źM�ɂdE�IO���5�uۅ�����i��=H���y5<$�T"�v�q�h嬷>y#H��	��.�.�p�:�K�{�-�� j���G�⿓�:���SW�!�;���9���H,�~�6�t��t��"|�F5�XM����.�x`iH��4rШ�-�M"������!z;DnS��ƙ����?n�Ty}<�����7�r��R�kĲ�ɝ������(�����`��e�+v��~7�� ���#pD�R/=�=, Dl��썊�:ԓ�d2��.3�r���̼v%W3��E/G�u��\K�7�@��?���2_q�h���æ��z��A�X[��1x'Q�Bϡ_�^�>�'ۮ�J�9	!��Z��q�_�K(Zˤ�P?,+2�@��:��D!SvN|����1�w�A�B��M?)���^�����Ii-�-1LƑ�8a	��>��s� u�Z�MN���o�S|��"e&�eyU�Si2::F2F��4�޻���]�N'	Z�p������B�nG���e�W���ofL�}JݣB/�y��<v[TC;(�)��W!���W�=�k)m!ˌ{�Ʉl�m@��S]�C�<�D�V�C�|�G04&�[�b�k���u�^gat�Ȳ:���O�=k@��{���u�=�+6���*����֘�Ӂc�o�ؽ@�[�+��61�5�mi�������X�p��w?����� �]ʓ��ɱ��"і�[R�ñg�l�.eJ���렱�|g�&��۪ܡJo�<1�6�{],n9E�N9��U҃tc;��QӨUU����e��~M�e�ޤ�8�S��+�H�8�,��f<����տ��d����L2و�9H�}�WC�ڿ�uf�bl$rl\p���͵:�-)8`�8��>|hT�Ka�ͺ�����sQ{û�%�*ń.�CE���e����{�D������x� �s���}]��Gjv?0:����-L��ə��u\�*~��BY�I����9� �>���M�Dp����#�g�8�d$����oȅ(-q=@snb��Wg^{�̓GL@#{�@muu,i���I߄I��d{��((�nI
}T�]Xf�	mY����`��|�+a��-�n@�ŭ^�Z�"���v�m��5�����D`ƩX�tВ�r��G�j=�X'9�3��cH@<rc[އ�L鼡S���s`ʍF��z?�X�`�� �
�Jn�}|J�?o��G��1��G�>zu���J�����诓=���C#TE�h���r�xѣM~۷m�
�n��m��e茧��|�|1J��]1��i����x���n����[0�U4���x��B�{m��a�{ <��ԓ������8�ݢy+h�G�T�;�S��S�PF���xS]V�Jѳ|_I��^��j� Ԅci;!k� ^�J��[v	5}C�}ռ�є\�I�B����H��]�zV�W��6�M�ƨ�9 \K�dZu��>Hӝ{���F�*Te���Y
J���ͨ�r�3¯�:oZ"�����D�L�������^G�ڰ݆�r��'�.���t4�tm|�z��+HwWbLE�)Wp;� P{9dQ�DD(U,��o�y�����,;)���2�d�nyMK+��~����^�99Oln�V�}�$�(����Ѹ6ɇ���B��FD)~ƭ�-+��<S��É�9�j�$n@��b�l�����i$a��ʇM�j4$��g-�?T�	�J��z-�Έ��Tj������_?�0p9L�&{�+B��W��՘2�����(��:�H�P0��qrz���`��w*�]<TnIP_������.\������s:�=B�W�Z�3b�;�0M0~�k+�=�����U�93�?�y�>[Z��*�5���=�85�m^~T��)�W�J�P_�|�Q$ǖ�>��(T�� �=��(�D�����΢O�\q:y�D���j��l�>-��\��D6����P��M�Qs���/�0�w���;P�&�z_ dС<D��?�Ɔ_��P~��_z���T�1�B����+E���D�8�z-*Ը�s�8�,���2�Q��!���윢W�z�]H0ݡ�1n��zlt���ƞ �E�i+2N�􉒵<j,�J/n��,���!Df2�;0���7��<H��kfu�v�{y"��6�$�3�OcI�	��	��
ऽ��`���C�������,��۪�X��u�Zvq�2����W���6���-��NvN���ćL	�0n���a�L&�>�1́{��in�M�T�:Gs'�^y� �׵n6519A:��K���D��QM�Oc;t�i�5�G���bpF8�2����:��AH���� $��hdA�[�I��_�<lgё�S���j$7q�(J�Ad��z/|�*��&�ɲ�
@I�Ǽ��I{��ֹ��6��5e���v�)ԭ�a6[�_�9�3��ߓ��*ӻ�d
�����v�á,T~�p���k��,;D�+���k�Wb�x��$1X^�z�R�M�r�zʸ�M�]�b�Fw�X�U��>2��BV^i��u�'K~b��P�?���IH�����M�DZv~�<���5����COd}q�^�uC���5�Fn^���?r{��s�?~�$��� �Yx�� �"b&��/=\aMt�9�Jz�jN��u���=�5�������JҮ���󽕻� �0�fB�@n����&�H��9�W�n;��e��i0����1ɍ>�Ӓg��,ݝcTRgQA�v��n�1DL�4E�yp&�T�����q���.=�j����ui�O�=�h���w{�e�A]���?����1��!��ZE� ��d�wi3�%�aL���R�/,Y��Ս����`7;|�S�����~�� �o����,�K���%ٽ14=�6�a�24�膡ش�;%��K�|����>��N�[��Ol+$����8�f0����khʳܩ�(��Ƨ�5�-�t��GP\�"�1
�*Aǁ�u��c0ou.�Μ�؂���b�>���}(�W�\��ֈ�(���#*Q\Ǚ�����)�mG�6E�I+�n�O�o�[x�ǰs���%���8JFn���HcP*�Z�C�.;�����<�\|�o5(G
�6��~�q���V>O3�9�}�%>#E����ܿe<-BJ4�����?��ss+_hȤcb)��7�� c'���U��5C�;$7��K�9�y�,�c����S^�e)��K��Q�a8k�H�NP3*j �;��,[M��<J���$�;�]��~��T$.є�~㨹���ַ�Bi�շ���A�-/5B^��&��Z��yt�s�I�Ӱ��ul�$�0�W襻=�D䒞����y(���"�/B��D��֐�%��㊈�W�wS�0z�z
��vM�7�Q8춪�R9�C��C�6O�S�-���kȬב�\lnzg���'�U&�~m�D�D#dyV�<���ڤǭH��!�33�۫�GP��}�DF�8�l_4֔ԍe:����k�y�뵖���.��Z?���)�)��'b�}�q��9��ǆ�!�̦;P�Q�{҄��E��#���k�w�[��1'	.h�,��W�J���a�1�Ȓ25�Zm>E�}�m�d2H��a#�D=���O�Z�ٵ�$p���3�����Z?�t��ڲ�du,�{f�i{��7�q����>�p�X�6�l9�P[�s�:���^C��byl~g0��^RsI�t�vR������G,T�Ms���|8\]����W�0,��c��`Y�..C�2���FZ����;���O0�F^���Ws��"�}kl��W!����>�!V������؜�/��\W�o"W߀B�D���k��:���ᢇ������ۆJ�!%�f�(T�1=l����{3�Ez1I���5�M�o�&�eA|:/E�e,���d��ma��)Z��ڮ�X4x��}�Z�^��")&b1�*��&'��;�"�\���9mTC݌8�����YH����D�GZ򗐇���e1v QC|�%�
�28�#
yoȽ�EI*��	]W�]��er��wW����n�;�6S]OK�TU����F����?�}省�?�EۗLr�'�>��NW�>�nX<Xhk�ٗd���%�����a#xu�	B��0BmOR�����4j�h�Շ��j7Td� ��F�0�?��t!�e�g�٢��.�cr]L�����Ұ�!H��i�cx`rg���?���;����$����~�H�%�V�U�H,��"Utn�I�:0l$����a$�k�#m�`2Б`	m{�JG8�ٓ'�*�����_<��|*�2��yWE�V@�E�������˃��?-�}�>b�1�WC>xщ�o��D����`�ϝ���tHh
�?G௧؟�E���}���m�ͪ*��-��k%zF���c�ӄD���`����l\z��z�=�e{�l�E����9�0��;�`�eZ�K��d@2�Ö%ORG��(�\ׁd��Y�`Zy�^�̍������G���]3͸��WM��o�N���?U��Vb�����F�\��)+=����
i����⁐�B@����{�#�f,/c�&�c�

��65�]��y��}"̐;Sc��Pd^�֩�F�>�Tc�c���"\�P��
�gd���h��>4�z�*坺\T*Qf˾�x�C.���z�K~{}�<ZtN�c���p�٬�Z�|	Ji�'}|�\��̵]Kpe)o_�}gג�k�UO���[ZO�.��.Nn��ʶ)L�F��C0D[�W�f�؁9�b��ѵo�]]��t�ᚖ���M��vGO�UN;2� BI4����YN�It&�"�[%�O���wB��S������ϱ�*���<�n@V�{�xr�_����a��1H2냝L|��+lODB?:��n#�T�~���*�]�c�����r����! Q�6ȓ;�#;!\���2�����.��r'<����a��5E�Ӊ�'��|�Q����u�"Wg�bX��|/1����!��;
��M����_�'��4�#�r5�aMj�bD�
2�K?b�v�>�ոm����v��"�e�ڄ?xb"�p\��~���&�Ӷ#q̍U���RU����wA�<0<�B���O�۹��
r�(��s�zb����?.Ͱ�m�a�RJ�PSť�R_����o��Tn��&�hy�G0����a$�|��.�0$�=��4܁G���Y��Et���$beQ�Kw *y��{�<�?۪��/�**��Y|8|u���蘉�c˒.w0+D���a�1'��=8�=
�Q'q����1F����(0�v��3�?hl�D��G�;�S��"����zRͼ��|�wB�"c�L
�"�YX�����P?�rA��m\�_�'�y��.ŪTs��v�1I��T�]��O�����5d��+ލ�U�#e�Тu�2>��dH�e�u�dk��fq���)y�]�.ѓ��?��vq��0��l:�2A�E66���eF4~|��Z���q��,�����1^B�p�iOD]�<�H$���������,�@O$Zg,9}�,k���A!x���Щ�s�����`:�nB�d'�6M�����FM��I���$�q���vn!�k�^g/j-����꽢<l�d�ZW��I\a�