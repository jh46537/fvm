// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g8vtqw60el7AEtPwfboJYLbuBowOb+yjAPd8S/Gr4u35zuUN1kPq3KhYdNoT7t57
eOq644RwBkUGFGyJ8xl2pl8jqxTRVDdXF6VahEcug6Lba/Kzp+vz6fMks1y2KchS
JMGS07usfNm3+fIm1Rez3eUMrhc+WAtlSv1Rd86Oatw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4592)
m1GLS39OdqaqWO4JX4qxNJP2LE96ZcG6E9nENq4L7SjVd5QPzJzMsEerHzMCd9+V
fJMTVi8CxR9Z0hd91434j/Bir2pLcMxwPgkgERm+3CnWQx0KXAzVz3pOks4+KfVw
NqkzL8nFJ0SG2ZogniyJV/FGF2g/bVD3xgdjzqiZZmP0nHQzB/GXwIqg6afVRZCF
dUduU0n0ldtp3YosawkJQIXW6PSSmDfYFZ0r/lLYHxI/+qdhGM16T44vmQumFDpB
tgtoucT6X4/6+5qBwlQQfcVL4qFfCfYpiHJzvfzd/jkrZm3ep/sroOS2PQS2tgiy
cEjB+dYBHziqxgsAJTKd/lhtDv71+b5ZNKTcc3F2KpQtY7rT8ADunsNNt4wi/Poo
x/BxGJXoHbW09SVpWR2Os85XL9NqY40XZG1IBrU6YKY5+qruz/+HSjleFictHDhq
/WXuE0Eb+Yd9DeAWBa7z58pGVbFkWwJBUKIji0V5JYQ0xxwOUaRkncVtLX9EJk1Z
NsARrOeX4cGFZEY6s7iQe29fE50zan+2XDcR/StB+VXCsa19ZZSw1s/TIJXi0Xt6
479JKJIm4XYUvf3W4bufMTxlxWNmHTyxkEUXEGpuf3X46ph3I7FgsMmMMeXxtjlh
CQ6cQTrFJnixMOlMw3Jhzl8A+drRV6CG2uwCJgnw+1Uv5Ot5QU7wd/5cY7VJbr6g
HbSrunH+NPwPeDEupuutNegGF7/VLB4B4HmxesF7NWajloVJJB+5KDiOBz9EyspF
GumCKPsL65HTfubR8phHqIhH+/RFThi554dCFl7vPvodmb7UGW6mP3SjG/pTWk+W
Alf2+FUpc0VpFOwvgR1Tg/I0xkC7ETOzDQHzdBiqtKAgX3riSqaJgmD833YbDWOk
/ol3/6Ky356Vzjd2+EYGUXePAi3HoPLxBHnhJypEhde/cAUx/mEUXwwFrx4NMxYX
BDON8/OSeZ5FDFryl56tKEE/tXbuJgPzO8zlHx9IebOWAJuhoZ+dE4gwg3nXFum7
jEwYw0roO+sTaqaAKENd9848JpobyDqHX7097sfdvLVVKs3IaCPIO2D+Hd/8oSTL
YI3FDto9lKVtlPe8iZhct/hWmwUlMF6xUvn3WGnW774aEfEidOiJsQ+siqkG2IV0
1KVwn/JoggWPSak4QkkqUB5nvGWyUjwyV0IP9lotG7U/yjHOorGappjobnBiyZbI
jGgTYb2/TaoXK1t+sqrt/Oqsunh1YBWA7wn65Pir/o+FeTjLulQ/RL3ufgiJw+hK
fxbvooztwQMqP/nhEQlfJCmrmayERY11lq9I/fzZhBTtVse1zzZql8mlPCt51Fas
cJy/aiQD4Jph4gBxO64AGsDeaQJv3r2JmUrPLmhz0oXhvVtmyVQgM6xmCuXY/Ux8
eHfTqDPXsGmaqEKrxW9Zr1Bzi24tOv7YR0Cvpy9qUwDc5Iq1xzOUSq04e8+a5spQ
uftkdt4JnIaSFeQvBCAGwpOzPZjapwoozaQKV2OtbeUIdTSBDc8Xu+eAkyg2t4jf
j1SMjtWVoFQRTx44VOZTwRN21KlqvnwKwzxFE+TbtREMMPXRGS7OK3nlYN/l4yn7
HHFFBU30tBBbNwa/z6IZoJz/d/oXfL8/0aqB5rPMkB4n+xmNDqSjFM32nHarqN+b
PZykM6HTYScEWNYrYVm0yG0l7/F4XcCO98eTVYiB7yZNMUPvZjTpLXEL1LWKRlpQ
0e6oECh4ds+O5ZorMKXSjy0cloXdQ6dWga8gQPN3K1i4sg3THHn+fKD1k8zYeQ+y
COffXh5PrioQfIL3WE3HP0Ou1nFeUj1FLRleFxYYkQdIPEmW/zXOyEz3vVE0YBmt
qr6bJulZ06exbF6r9IQxA2vQnrwnK6CmJO+WtRwb27895d3T3B8sEc31e+WcVN6w
dG8e/DVeBtfYtLDOnyJZlR5PUYQm8esmgAJJH4+inJq2BNuP7FPvLVJCm4zeJGVp
0QamhhZM/qiCbPwoRseyQCVwEAaQDGMG8uYmDohQz8FHbPGM9BFYhHoiNeWkT3Pp
je34e8XQ/+sYxoSqfy5VZYHdB/tQwq3yomQHnfHxt8017w27Aj2HpNXlxOX0fgyR
z2C+wnEQ/J7ecG6mRAvZ+5MxopnE0RuwrWR7kmBBSOpHdhF0EcquLCfXtJKUYI8c
TsKzHWCm3I8pAMCjutKMlmVkFG1s8UqOpf5EfxMApAXIDxcQLgdUrq0QQZhTtAGw
yxwhL99T8OTp2Ea7VhNGMeYTPsZo0ViuSaE6a1oLvUzg7IYKzmhiyHNQm2pzqOyb
P0m0KLaQ2A/t0PhNibfuA4UXXNFw9f2eRFdpsX2kqcRzD/NwEdIX/vvCyObQnXDV
msyKghaXvKTfOXKl/lvvdLOFD+AF31d1EfEfKnj7lgyey7MLNrTT5le+frdUUcfa
n538j9Wces4oQyUI8Fo/1NcmaSDqNUdyYSgSQNojqpxem8QLyKTaw5yH+pY5lIpo
6162cnmd6ZaLvCUGguJO7g2ZSkUBMCHGy6K/oBU34KhYalMCi1LVe/qLOpc47s2x
3ZFl3eSJM0o3Ha8ErLu7orR6l3KWysujECP2EbC7iJClRtgMolNTSC1mT50p2xwq
3RUUGgO+FpE79VQSrcDtjyqpcl3JnN1V4N459M9jyYkr3LQ7paJBffU83PgrIqvp
cg0saAnBUIU95j4W8LThV9R1QhewdCmNz5JXiZbrbhEbxlW68SOydb0A9Ouq0JNl
VuqMmFCuREKDjRx6l9jGRaq5xetp1Kwu9l+NCZ3JdxDCi4rrBmOhYisgj7yadjG1
JiuUDCYnLKEsDR8zzl441iXpcPjmiq18BxZIaaec4OxlWCNrC5z3EhY5PD559mUi
ZYOn8BGyDMiUYDGbsYn4mJ6mcCm3lvC7IcER+/gheVZQdEsOnnh+VJYUrLWSuWZk
8kffXMOmxpn6Pf5SAaFcN+aNDO9n3S3huUjQlJRXcZvtsxV13tbBS5DOXcHnF14O
jt1KBTayYiDvCJeTaoKkAs6D6JqdPpUk1SAO7xqDv031IiCyeS4Ar524u/JSvSDq
CO4Zc4/iigFueM7xsJcqZuxOSsOmtDEOKrop9DL1q3eYPydhLayTwTVzOnI3GB8d
zGmbYcAfUg6jkQ53tvYT/+xecn715pzky6ebflz2ZlQCr2NCMSo1Nth1Bnwi5z8x
KQLtdQJdb2LRRdkvQYL+y3upkic0HsoWe7wj+D3ccmKEEUoAQROhZ9u0AzMS5bEf
afIlrcqRjPmsF/avTzkm1CEaK1Q4H0aTT+GJweQ5aObXu8zqu9Wq38MRljq0otSu
N4wBGkIgOek6alKIqK385iYqZRSOega4HQY2vzclSq8lvEmg8so3UlgZoDt5O/vN
27nOllqwB1VcFdFEDHZcbUhC7JGrrMa3YZyp8bQqrhtU/15HvvO9sMqpe/fLkNiM
zGrFtXSCrqu3tf6UhAIOBBjJsti1c6WD6mH4rGfrdnf+3WMzewZ8AQaXBmvT82ur
Q6Bp1OAqZrTL4cjp+in25bgeNEUEkHViRsFY7Smr7Et6kZzABQRwPZvmsAZtAsSV
GNs1Apm0BsgoD+9jI1pcLWPKJ/kjE9VxshuadVAcfVEL5i4LoTjUBu3JrxrYRCas
+mtjiwdzYCwUySM3N5KJMZSsXV8FsiW1WIKnSpfmMtDyCPFcVXuWyZ1S36/TKOKc
Wo9zgDc/UYCS8XqQstdUqLAtmyStB9hud+MFGhtCoYox+9cwR/r2HSXwakP0k5QO
A+L7y72w9ePTKD1aDSCHC4TrgpaHYaxl2tXIw67cmyfvO/7wNEHyZigP74hdMJe0
5dJrKpXZ9WniyRErsGb8bL3jFdMcp7Xmo1C6m78X+ayplZhCU9EpXEGv+z9C+sR2
RsXbY2UUAnx/v1byYEsPQbzkZsJXX4hATH5FKz64ZijuI15zppBI+jdOEgsNuBgD
6ael59omalkmGFSChb6T6lbmrLVkoKzZUOclT5rpdHrWtpfNn/mUqP/F7DUZIWLl
JFAIrRR23OeGF/oHN15XoJ9IVQy19BBpcPdr85zxSPxo0wl9ucGSTZ0obUeIAEi/
ku+54KonAPeTEt7EKbpaSAffzcrEmavqO+7tv8TKBhB4U6nd4Z5+J+9Th65NZUHe
we5lkKzj+YqAgmgHBa91LCzaLAkvLlunRu9p+OCSxNuO1f5/4GDAmsqRHS0hlJXB
G/AvPqCyziDfGV+9S8yL6xR4fFo0ExX5cJbSqT675jfNOZ4LiN6Ekz26T7RdExSE
buznTUk4siuBlb4P9M6fwBPbHBWGTF87FKVPKGEotH+bnjXGDJ+8OmpbSxYg411b
GKaUJNAxRl/0vjIdg0eeeJp5PQrGg58B/HZ2j9RKCJZfdz/3Va0f1O/8xJkfg6HP
TOu/9C/GFVfAehEH/0YpbP8s2ZslQJxX8xff5DrbnFvlOHP7s1OwL4Y5gnrIwTGj
38NVpiyhSmFC2WxUy0fIJFiNp9chSBo4KTOwVFmNIxY0JAAn5OSM6VVyO2SCXo1c
T6t7k1xQladYMz5fwCR8Hr5HzVx60lrRRxg0M9AZuL2bKbtcun/iDTbrzSu45hVp
DbP0Rw5DM32PqLE3BzpwBkEC0lRrDbQ3zQirqoQtAJ58YZJl20SLz3nvVz04HGcu
3GupcAlyK75pj0Yl3BvB7UHRNkbQdG/c7qC54rYSn5pzS4x7DK9gQhVbMesOZaJ3
TicZSNwo0MRr874qeKEg7YCL2t+u+AUp/79L+16bz4Pa71chhMxerbYymCh5IWBE
rZT2KeQfegEANYeF/1jglNmUcZD9FNw60UCH333UtwqaHjDUrM4n7/ezgmbmi4JM
qMFWxIry+mGAFmvLHlJsJJ6W26vmZtwX5Yi4k1OwXnCZa2PhnJEscabmtwXy19Aa
YeWZKs7av6W6F1Nj+QlDcpKlZhoEPwbdjyKzNcLhL+7WCqXh+Zl7GdHcZMOYW831
MvHD2Q/8q/aeJpO1zKV7BnFMP1cInmb6cKeBZexUgJzAcPHkZkkK4xYPzmDzBVSa
kcZYm9u8Xmy7jFHcmpK5H49LS/CmKKHeqmc4R5iZ6BwI5SOen8habSxHN/R5BExD
vPcQYztDoBiVQlzyXoBtkKTdSLIIrz0gH1YvNbOq5pHKqz2Y9l/XAgQ6BXIvhrTG
ED/nlL7z1MTeLiwINBPPbgGMHIZIsHcxtZ/trxFTR6XBrf3kFTSWu5lEQj22+5M8
1yQsVAdDpqe2pU9cfieo17Ty8FCNenQFvUACrfZ00AFoeswI21gYxJNdJ+TZcKPS
yG0JiMz6hLHo9CnP3cmFA0BrL54IR3PbiJ7SmLwasAO3s/XIOvKW4ilpUs97UC+h
wUsPhFJmkFp1j2SEuc/C3GicccygjK8Qm8LrXiDRq/Evwmk7HoyG2KS3mK2f0Njm
QjVQNIilG5loU9OOhUvQlRZVi2o/a5Q2xUXrm2zrZnhOWV8CQFnybZ5NLPkFtXLL
23hlwF1WmeprMAig/vA9RD0htxSSy2QyYO/0RKmhyjB56mapO1qsNZ8K1w+7Qo8n
rrV/ZQsvqgC/rUZI526gOSHHeqTOeWR8Y5mmEi0ili5h2D+23fZDCdQsVH3VMJjV
5PhHUFSnDTjqxv/yZhrUXMSNJ8GAox/UbShn52uVmJCSAPzWtQRR51xCjLjjuhHr
28TiEt7osWyFD7OB3hoUX24qmvgeNc5VI/y9ekklcTW6HieUgci/uPAxyDfvkH64
9+vEOGfyAN2zDjBjf06LG+tvvjM9GXyO6j2++eB87s0NEgPcR2uB/RVM8HRNjTcn
VY9ky9T4zCuJR5TT1J7yrLTUPfTFtsT2miQc3SanYdJpiIiBs4KHlpnamt7NOCOy
cUiII6B8zonGTdJr0L4BWCOW2kRzN6qdEgvobh5DxnrxEDPY6e0KiEM9BL85IhAh
hKQITUfi/tMc0/i9ug3FEuVN98tdacfRFq4SwlVFYTi6YIfc5e+uK+/571FcsNv5
ssqGUYFVK7WHGvhmdhLyp4nsGz7wHGAcnMhFjWPAQgxx7nUJyKmCpyzXZ54ktxWZ
SahHkUBEa5pZrEK5iMWVAgJdv4CoouxqRfTo1RFzZRk=
`pragma protect end_protected
