��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,VI�0=�E����pbT6oplz���5���(`(h�rr�����k�ʩ�^?F��QM/�����ӥUq"#�"�5x\�$��r,��$(a!r6LM=���N�%���ڛ��4�<C	:���==���I�)[�H�����8Žհ��G&h*rғ�����Ͻ@�N�N�U�y�P�B���l`�������Bq�٨�2���F�d�G\�(�>��`���{}Lt;�2��״�eZ� �I�o�g,.�ڮtX�N7���$0���
�&/�f�ӫ	.R��=W$>"�ҿF��u��[��n��C����w�159W�s�g׭��8z�i�y��sK�9�����ԣ�"S����8&�l��@�cJ����&�*3��a����T��Fn#>&�/ɀ��_��W�j(�ʃ�6QQtH�,��!0Cьu���E�Z�g�Y��@	�{��&�Uk��׫6Y�^��ܦ�,�j��X����"�t���z�6�3x�阖/�4��NPMg�Z�:�@��a���'���m	He�KEZ���	��.���-* ��S�Ї�@J!e,��3�wi̪�k$H�]1>�7Y$Z�q;�
�S��p#�X�ȯW�����^̬���m�$'.�><!��mz"�v�����21��r�
h� �����K��ߧ���T�s(��`��OC~h�/�#������ w#����m��'75*���+�j֬�o;�#�$H�i	���Q�D�B#�f�E
�
 Q�:�+�ywE$F�N�� �������f�U"�JJ�4a�Qh�S,t�v���M��6?hF�هT�\��O�{V����6���9��Z�t�5���3�l�x>���}�7�(m5�R���{f�[�*�������h��!&��$.�ƅ���,"$��:f�I�L?����"r�I�H��?X.�dl��Xi�㸒��͊(�9[�������W 6;�*���G��i5��X�spG��_�V#�w(��0��B�&ܚ���'�d(W4-�=�bxg�Qu��m�c�5e��Y�)�r-�=ِ�Ū�,2��S�D��T�����4 �:&�s�Z��Ү�_�.���0�i��>��6% �
�~2�W��'�[�_~� ���~j]@FEm�a�!	�'���(2�Iʁ
/�&�S�U�����$����u�W*�T�+�.D�H�-liX�blar-�I���vEA=Nȷ�IJ֢N0��p_��W��ռ_R9i׶0{c�֮�R����e� �PK?����N�Tɭ������ƢS<��H��z�Z>�p�����ߤ�m����y���Cl��>(��
�+!c�{�=�Z�0�C�p�^"��$'��x��Fx��\_�@,��vL�������ʧg,�Ӱ/Α���()���w�)7��YZ�h�_�Lh����i)���ej�B�9�:Z���yp#�oOrUa
C�)�F��՗!��n�6��	[Q�T�!��$�����uԳ���k�ᙛ՞�싆������#r�5u�Ϲ��C�SC	�M33%��!9�p��^S�^`����*;�1W(��~��)^����X@����ؗw��O֖[ծ���?��K�٢�8^������}�oa�'�͏X(���o���4�حKK�ᆰ��Pҡ�7���(��J�h�'Q���$*#�FκYG')������`����	�4D�mҊs!�#^�^�Ut��9^�CN3,Չ�v�TwK�O�!�"V�ڕ�ƍ�!����|:����-U�mر�CRu[���=a�%q����V��J�w��_��9 ���G�f1�Ч�K�߯����LiNS�����h����j�aX�>e�&|����4A�<��%~sn�V��@�u+3l��
�N� �Rnm�Y�u0%;��_�}(��\�^;T#$�Ӓ��
��͙���;.�:"\s�V�&s������i�h�xZ���r���m��!���)҈tg�B�H0�Z��Q�`n�k�vR�x��^�E��c�E�����O��B��H��S�,��R�:�^BKʸ��cPM�GTf�#��RK����	SɾK�72�_iD��ܢj	����ѕċ���-Y`��B�U.T�^i����-sO���j� B0����+�Ί
���� ��p�)�xz�F��3�����$fo���x��ܞ�*�6�,�Kmbk�JR�zQf�a��/��L�t�l
J���h�(-x��Z��Q�O �@vz�#�5�%J�n���C/~�Lj�(x�C� �wU�����t�U��s\9��-ixuR������|��"T<	�K�����B� )�+.��#��E��t�e�K|��_}L�:��\��5�wː�e*��V=M8[�fCƈu0QW��א�����3~