��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B����R����l�JxM%�$$���E`�����o)lh
6[#V&L�.2�%���1��(|6����"o���F�Q�,���-eQZ��m4�`�b(�I���w2�Λn�J�~������%@��~��� `aG<l~�tG&9��!���Щ� �;գc]���6`�AO鞱����r���D_?���0�����a/��3oE�p�:>�]������+��M�Q�'̌�����{	%�92�L�,ԋvm]�"3�F��Lr򱗼ݣ�65�R�?�}5Jj�%0Š������'�P$f~Ad
ң<Be�7Z��4U`oHj��3���܅K@��6��	����u��//���Z��ŉY�3�[37jV葝��;�[�˟h�ą�x-5��aDX�:�/�)���@F��+W�Z42a����G�>�mr��ʢ	k)�	l2	�j`�b'L�sTv99V2F+��'i����x�"�+u�@旻�
�8Cs=E��ii�#�J�K|�#	�鄊�j�ç&*�YOT���^W0��N-^P�qk�Y�=�{�h��Nu��O��>D7�� rXWey�O�%��i�_���#Y�P��i��iKR��Fu�[F��� 0X��#^�վ6z���(|c4��9���Q���3��q��E$���5����/"3����!�,��Fg
�d�?�^W���р���X��fE��L��~|�'��iox���_����/Uӏ{����R��,F_N��E��L�BYC��?ij>�|�e��L��l@��»�W�$�"�=>"m��%�g.�l|z�$��S�T�y�JQ|*����kO���K�~]L:�X��hl��m
��v0����;n!���[A��ͩD�*��#��,o������o~H#?�����Ͷ��7[M�4��8_~8C��+�Y��f�H���yd��}��/���K�C��/���]�1��*����}���f��f�]U�bB�i�Q�Y����'f�L�)��9鍇�y�L��/<��l���l�8!�ET8螶����*@ǳ���>|����tn=W�hf2�8���v�/&�,Sd�U6Ϗ&��cT@��fT��*�?ˢ�m\}����(����w����F�ռ���K��<i�����p���C���˚qC�`i ��ԝ�%[+#��Ԧ_�����p_��.ƣ�w� �I��f��:��ŵ�K+�I1��Ih����تK��dd���s�U*���ˤ����V��~��Π�'�^�_�=h�ɘ<� L�$�Z:�g�7]X91���VmڞeTS�@��!��� �6��;ڀ�����!X�J��Li��24/��=�8b���D��t�1I[e�%�Q�i�A�G6Ϲ�(�:�b]y׃��V�!�/��@��q;�C��_������n��N��W�<�����ps���y�s[_���r�C�!��1�PD��
�K��1&kqݚ�e����bS���2�%���?���
�A)��h��2#v��u�x���)����.o5�1}�����z�z�O�o<{�%�cQ�ؼ��o+�\
�.2���0�~������\���8�#���[4ѕ
���e��#>G�d��3��<�w��>O�\i_v��Tl�WlF.��DD�j�����g�%+�N`��D��	>�*ڬ�!jK��������!f�θ_��d��S�����,1�G�|������e��"so�[/��Ġ#O|���=�Ɉةɂ܄B�d=h�R�z:^E�:)�<���hr���ۥ*��R�Y�*�*}�&���	�\�x=7������Ɏ"��=��O�3v ����T:ou\�${��N��^w���m��oڪ\E��2,���{��өJ����f�D}o�hK�]=P�rݡ�TvQ��گ-(��ؾ�����dكW��1����.z4u�݈���7'j͛KoSlB��>������9.�S���~����!�M�d�ϥE7���s�t���vl&�_�m"�Us�����>vJT���d,��ب���߹�fT��خ4C��@���F9
��͝4r��&HrK$�i�
� _`"�bA��������־"AAb�HU:�}ez�@5�����D���T� |��御ǃr8�'�ƅ�Ha���_�w��%s��k����;+h��(�Z�D=s<C�D����y�2�{3e�/���� )�%3B/8)c[�ީ�zl\��H�����p��/��E�oG�h�⨀d���ߓ���[P0��B�}J��o���C�}$�������%� ��河��w;�#�[�-1���;�iUR�%�T6q)�ª@@+;_���ώW��nrR�R�̶�4=1P4�̓qc\L�q�[�I�N���y���}ԥ�	_��\���_��Su�:V����B5j���eB�����Rw�!��7��9�.�ʒ]4>q�旱k�GU�L`���|4 �)���oj̕�_�Wtw��8,�A��q���[2*�����N���2
�6x�ֶNn2`J8���Yc@�<m�=���h�����j�eS�-~�Jr��զ�|Si<�.��n���z@vf3df�v���-�i$F�V7��q@��w���?c����TSNv�;�FئW�����'��U�d���s�-,��>���A��3+��z�Ƶ�y;�mg�����>V�?�sلp��z��oW,l��zD�-)�`�G&$�������.gd��]vO����r<�ڏ�K�q��2J�%\�Z���r��d�:�;/4�Ѷ���B)��<�4��(�-w�NP��j���_>�g�yG{�>ڔ�[�Y;��ŋ�P�A��n�$�ѡ�a�w����
i ��0$��Z,Gn��2����iNݛ;�!G�֊����p�ɥ����ys��
�~�q�j�!2i9�7��f/3�ۉ@��N3-'ʢe������T�Mws�y�_�.�K�h��~H$�c��M��ʅ���)����F��u�C�<툫S��i|��	Q�9�Rf�'���O�MY��nvk.������@�AKp���z�X�*�Q�"	�(٦�!S�u��b�ǂ�jx;*���U-Ȯi�#�$�` ��c
�~~�@��a�sA�W�]�uﱭ6���U��t e���;"��a��e��`��~���n׻"�Q��mMh��`���0��O~9��8�㶓/%«��n�<�;Ix�b���SJM%� !����Fdϫ�,��7��.]�u#�*V�SkR���ۙ�y����̥��f�⹔&wV؍��}蟟f1����&��K�0���U�yW]JL.M��c��"]Wr�^b�*m��M������Zn�����W���ilིpM��N����Iyy���ј�O�;q�wBcܓd�--얝)[x!��MA�v�ՊoI�|zm�3qa���;y�G�b�D�W��$��^یx�ZK�Φ���U[(�٘~%��qL�/b��(݋K]�k��X�S����1YI�*�>	��,�6����n����D����<ds �����.���U���[�8��Fc9*��o��9@����G�Y9�`ܙ��6o�?ӽ�(�����'L��ψ�΃EzNg�g[Q��h�����ѽh���U�]?mb�i�߲�pd���T���8��\H�^Q����Cq'�4�~y���?S*���7i�#��Fa:�0.�I�p�=�B7�E��n�.P����.^�F6�5?�[r�6�@_�[s��M{���-ۧ$U�������0l��/��Xj��S?�>���K`��U���>3
?ՁK/eT=��㚖'A�EG���|�XpY����E��_2� ٤M,��2��{�@gL���*�;QBf@���	n�-����i����2ܡM����8?沤��N�|�73q{>5kU��>VX�z��wq��V N��+���T����"��}|oNsD��	:�;���42(-�7䮵�3�v~�-��Ӛ��I��[�$hfOAi���:�Jsqg��<�4%��aX��e҉��)��@�_er�]�	���v���t�<e�S�s3z�m���&�vB	G��w\?�`C>;�n=�
�'���,����إ����j�4��!${_+Bτ����%���!�$�B�zU`� <Ny��p"\�NB����m�q'ԇ�"^9xi�yu����k�Bq� ��cW0���aEV��Vs@�U�m`��������P|�Y �N,��{��s2�sj���6��s�ά�Yx�K���MH��E�w�*�K��,�Ðx���#�axk�d��_�d��5��X��*4��Ѓ"#���u�=��G|V�C� �)߱�j�}�r�����?vO�C�ﯰm�����=.�H���^<���[��k�)�OI�\I���́�r�e�8k| ������3����Ef6���oUN7��}�_,��	�����bu@���P@
`څH�i��A��jLu�:�����	=��Rp'����P2GI>}�Aw71�RR3���$uiW�$�ȩ�}7��":C#]z�a���re/h����W=���k������^���X�d�r`a����5ۛM���`�aFU�Sw|2g��)B�J[H�˃���ڀb]�K_q�v��}GA	�����!e��o
�b��[�E��Ӿ�ɖ����$��ZJ���������`��*����|j�e�G��SR+"�jݰ��0a�s{���g���p���P\��b�t���dt�@b���;&D����/T	l��6<�W�4����d��	�pK��麷h4I��6�}�zY�w����� �-����w�p���VM3�x��l�+�뤣�O*W���m�>�dH� D[����X�s�4g|ˍ�&J����dfC����?Z�N�(/��
&����͞�Xod1�~rgZE��!)(n�3u՜U��(�`�Ei���ȑ��E�W�$