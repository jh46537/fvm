��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�I�X��a22}�<�����k�`1⇎G�֕������`v����"��o^�V�&u��`���E:�t�9i��E��)��x��=��X��t=���D��eK�W�7@40������5y�����T��J#E˱m�@�:5=<
���4�[�T<��Cd@������{�V��~���i�(X\_��	s��e�&�N�Al͌ߌQ����8=ݾ&���f���*�^����Tظ��7���/��Hݜ�RPZ���e0��<]Z�����
s��	��AYR\�{= Y����p�_bӚ�&'�j!�E�.��=^�䯣m�����XR�)��$1�H	���>�� @�埦SbE��pa����,�A�c�3�LԀh�Q4̨�)-̈́�
y�Py�Ύ���x�&e#2�7��7l����=`Qx/X��͸�@bn܉N]Y!4X~/��?o���{.��d Ud�j�糦�>��/����7��ښh����Y:����	��(��>�@��i�a����νF؄�y2j�y�Z��A��g�P��{�����m��" �aa�+��OW8���G$;K��ާ��hv�i��+mx���Y��%p@^v����Xm��W��¶S�j���Mm-]]ۮ
x�'�[��*'?������Ӝ��⮎�D�f��+ɡ��l�I���X �w�?rڡ�q@ڦ̱V��9�+��r�B��/���5�������1�6"5�9@��c9MB�D��?#�����H�=����A$���gk��:�s<��5��Q^X��d��$��tdoE2����/Y�ep(�b���l�Ctp�� ��*ѱjP�v&�b!��`��1���.κ��%�?v}"D��Gm?��H������?J�o߂��,2�r�;��mč�F��"R���,�1 M�t�+��`����
��W�'ψzZ
��O��vӰ:*���#�[m`𢕩uZ��K�M��a&��V��)WHi�%�a���dź���&uX�7�JR\$��S�<`����u�9R�� �V5�X��ݻ�Dj�,��&���?1�l^�*h�O80�]BKy9I\rS FP���E�"�;b���4,GZ�3��j�ˀP�j�����BWB�hi�94����̂�ڰ���n�3(^���P�H��i^�f�-�`cHPʾdhMr{:LL��]rsŗj����#�]%I��D�s�"z̏ߍ����@Xs�"�R ���}��uCս3R�jKp��[~����*1-q?V)LZ�\��G6#��02X�.(4J�#6Ū�)s�j/я�A[ ����^&����Ҹ��,�\AÞ����䥜�F���ZR�����O��T1�-RhEO����1�#Pڴ��Q�$8�[�LO8�*#�ZfR4���?��C͡��"��ɛ��vdF��KT�t�g�>F�d�ՄC��O�j�'�Y>�l�a�ְ���E03�Bw��ߏ���ۢ9ʳ��ط�r>.F�y���x�T+v�`����)n��1-�*9�C�}l�> 1�%��F`{V�Y,�ı�-����#��c~�t�՚^�F�j���ſ{w��Z�����tDUo:mB��-}�R�?�G�x�oNd"	�W��d�>6��lk��$%i�K�P ��JK;�.����1�6w�kګxn�~�Kgƣx)����v|�^c �ր\���|3)��'#�_�9_� I��q��G��N�|���C�pc�Q/�$�4��@t)#XDjY�p�3��,��4�ʂ��jk!�_�O3��Z�O�s��~����m���'��6��p����6퉾_�����t��Y����t[�jn����E֯+�� ������?e�z1*�v����p�i��F8�  ���\o����(V�r?��I�r�L��FKݠ�p*����kK�߾*�]o��k�uXL�(��5�<(lC\�li[9���\Y�i���Ӕ�p�1pT��pSl�֫"]�����������MX۹i�V8��������`NB�,�� �+��'�~S*�PO�P�؜0�)�|��4ċ��P'�ߟ�+K�)p����O�,+����%���X�;gƽ�B��><)נ+V��*t�
��,e53w��r:��8G��V��g�<�X���.0}����S�����hx(z�J@��̅`&�p�&������9��Rt�Xy��bA�����B�%��,�ǻ� �Ej���.�Y���IJ\VK)��f�
���ɋ�?���r��F���t*A3�"�@���_z�Û毛u�Ŏu���=��%�����5��-B\ȹzi�)~<������4��5<,�A�2�4�Ʌ(%�!��J�;�mQ/QbRp�$�5���w!��b�c����`̈F�f�m��|Z�i��+���,|��,6]��/��UÚ�&m��s2x�\+~���&@�)M@��Ừf�W��?�n���0�L�,*�E��{�q�v��7�8W���J=q؀�~R>m;x���V1�Ko�R�ɶ��o"	+�_�x/�@��W#wo�=�a@의�(q�!�)�
�0�w��Ψ�㷃n�� Z�7�
����mc��Mm�����R��׌�)�?^c��6�t�E�t.�>܁�Ǝ���h��4���ֹ�6$p�f�k\n9�"G�����,@Y����S�ꑶ*�ґ�+! ���$J�5���q��V؋B�$pG ��#�?Syo�i/���]y8�-�7��b��G��I��v?�]���+��M=R���%�9��d���]��Z� �ŅyE��XL����u:oZ-�RݐO�?�}������vo��4�l�̨Γa#d@JT"��9�~¾G�K���f6?P]§��֟���$�h�+ޥ�%����B�A �l��l$��E�1�Z1����;Ec�r�����S#N�$�tR�� t%���k$�eM����d��ɧ��Y
Ry�gƬ��D�Y�f\�^�� �l�Io�e,NF��\���٢�1A�P~��8iud��_��J!�>=A�۟��Hߍ�s6�YP�f��4B�^z�b�0�͆��M#@�
�m%G�[���A������~�*j���W�*[�Sq!f|��m/��Ugc�_W����So���/s,��³Ni���BN>���D��\�WX,�� G�ϫk��E�ON��|͠�`1F�9���B�_���N����Q#�k<t4q��N5��A��%� �}{���y�Rh�����dY�0���d�!��qY5�Z�c^� ��0�݅w�J̠ &�����]��EU��D�� #-��Bzj�2�u�>���	"a�m�IN�T�j~��#���LZ�P�.�v�BMV�U�@~�SBx��[��2�C�/{��.����?�r����T>})�E��݌��6�c���V�piwa)�xÊ��SV��ф�������(�u�^͘@0(�k
�Z䆫��!a;}�3=|��=�����]����Ѧ!����Y���͓4���g���Ɋ���N`��<����L��s�,>W�Q����ÄxȦ�6�դ"EQ+��ӗ�8�_��(X��B�w�O0���$�n���&Ǔ���+���[��Ѩ)�{@�2wAH��Ff0�\"2_��S����T6z�����g1o N���T�$�pr:�Wb�0e�~U����V���˽Ͽ�ڗE�Y�)�Jq�b0�E��hIf�R�oP~��#�zd�&'��D_�M3 B���S� Y��oڨL~���u�@_��f�Y*gf�2�j�b� z�N�O>w�����t�!"�[Qԥgc��[R�ņ��W��K�W���Ú��?��� �3�/�B�e6P�Z8+���Ѣ���UƱ{8Xdy�	��V�βF�ZҜ��%���s�5}���VK6&�K��bQ.�&���"u;Qu�33����;�G4|�K�kA^�Û����+`��m�<�SM�V.����h@a��`��v�Z�wI�7����9� ���a��I�l�w�E�ENj�& W`R���S}�7H7@�'Q��n��"N�gie-6��V\�����W���5��
��=��:M�W6q�ɞ�8Z�!���RO��1��`<ºo�5��R~�³|[|[r�^'!�������Fi�W��/I8�dyRb�ڿx?Zj�})sL��,dV�k\_��-��t~��m(�;���ݯ`�$�
�
2��h�y��|�>��N2��%?�ajY� 1[t,��w�l<��<���K_�f��Oƽ�ߤכ�I�3�^�o�y�d#٠���=�����~M��x	��]mD�u009��N��޼DQ�Њt���W�-]7�wɩ�`q�iIW�P�������\G�4r�7�L�T֧Fm,(�h��S��z�A%�����I(Po洍�
n9�a�����=)�ɘB��2��d��q(2�!ZY��ӝ�z$�V��13�y�,R�V��5z�_�Q��w�e���h�M�����I�`5�m�\r��%7�s�X�b�~Q���i�n#�Ӈ͔awg7��̆�N	�*}g�=3@����{Q��-��|��Eo�;e�L-q��g�Ɔ|��o�p+.	��~-"��}�IȜ��גx:ݓ�`���x����S��j�/@�bu	-����Y���5o��K#3�L�/N�֣%�8��۟��R�h���x�l:ɚ7ƈi�5Vs`��q���*���'ۤ(�S����d�JTG�G
�A��!�y&%_PWf{��NZb��ʇ$��M�����-1XP��O*�g�[4���=�w�/�1�-J��T⛑�;`��wR1�ӫ���0��G6B�m��ȡU����?�����k��w�y�/�<� �{`ԥ�[��0U�A^�uՏ<�n�D]hj�l%�.$;D��N\Q�U��Ͷѝ���"@�.�<*e2�7nRj7$��g��vq�޿7c�|/,�qp���%���e���p٘�k��I]齷;8^|�6Q�6b��0�)XI�B��~��N���y٫Ģ���v���R���VF]<�#��t��{�es� �~pz��L�OKp/����������Jb�Ih�����la�r�0��^��n��2Ꮂiae�(zN���n-/���/jL�˧~��0�|l��s�j