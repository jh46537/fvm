��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7]�s��^T��N݃a�O�BL�z�᫛��uᑵ��@���I)��G��:䕂Z�q� y�KD`��k���������I/�ˮ�oʥ��dFf�y�fR�^��濶����~{|E�[EP��h�x��.YȔ�&+��[�d�L�
�x� �ntv��B]� ��^�[_���i�H��rT��p��mD	<γ$7�*v�ҹ��V^l��)��E�$��o�`:`4y�ac��`�龕B(�o>;N+\a.5��oe���ՈG)��9�^_G�|i,��>x�Y���=�R,������bS�zs@������6��d3Q6�_�/m�"i*���aLD��
(�6�zS-��xV�O�����'�TW�+���m�6��}��P�x;!;�$[�h�3����(Nw(�H-�?v zv]��w�M��.�pS��z00X�O;�6"�S�U�$� ��9�B��h#k�i9�y���}&�B�O�(������sH���)ย����ɰ���=�ev��51/�W���Z��� t�O�Ҍ[#�Og���`{Z�Q2�:��I$�g-l��Գ�$�[k�-��=�ޛ��_����{eB������t�r��+C�wv�1"	�˼�c�`������re�F=Nc����`C�2u����s�"G����9q�MpL��6�x�*�bs/���h�FV4�9�2�!H�+c)���u(̢�A��q���.���dcR ˮ�P-���0c�yy�������,l%�P"��}� �Z�"\�4�1zY��H��.n��UUY�����.ό�W��Et`L��@[m�d���z0Ӓ��G���1+F�\��E�kҙ�߮�fK�\��N�)�(N��-Z"0Î!�-�/[���鐕���N3�����_%��rzR�=!`Q�����r(���ĝ�R�`�ж=���Oή��-!]���u�ae,��k�:���=C��<�H��Y2��JZ�-�J��Ib� �� �"����H�1�0���xfMF�$��'��
�3�c?�&� �u�,9
i�z���2,�2�	��?.�/q���~�`���Ie��`�������e}�Z�b:)7�-K�{z��ܕ�Jb�D�#����vx���F΍R%�i�D��3o��cB#=��2�W9NXt)3T��X$�W�>w��s�y��)���9�>��Ɔ�[n�$�o���1;\�0��"�%3�_���ÉR�[��&虖B��A��\p�T-ˣ�H.Nz��&�J�K�'��C�� ��p�f_r�MS�����D=�K`�c����r�!��*<Oڞ:�$&Xܤ���C�r����������<5X���'i�
�F�?]��w��=�X"���-Q�qTBZ)F�a��� ,��t����
�x�����(@םIYnp<[-]8��� ��S}裣df�c|��[T��T���s����J�ﶡ���ɼ��
$M%���ń�T�| :vm����2t�9p������9���xzi�~шs�'\J�i{�G���Z���#dO{�;��(�[b�{*�d��~��|#UM�{� tS��='>�D�th"-Flc<1��C���1��s�R���4gkW�N�(�Jk�Y	w">�!9�0���E�kMa�wAۧS�p�w4�,Éo./��{j��h/6n���w�?�:�a�M��C��3�_��Mc��OD�w��(d2Uq�9�=[��#��/��e�U>���1��H�Q>�T�6�F=Pj!�ǣ��,G=}'��������I�_9J�1��o} W h��)/t(.�Nf�L�O����^U}u�t�>H~�M�B���1Z4ߦ�NV,��)X���|Em�f�$�D;C%�zg�����柙�bݟD��^y�Ŧg��D��^B����+"�ŵp���z|~�������p�䊯)�v�,�U	;��z|r����H˗��i��{�䷿
RL���8� ���>+��kNL��2��}��˸)��W� �[�)t~��@�"lc��e��q��d���'�� ��L�K#�L�������Nj�%قi��)�~�� �g�d<�.�����a��$�2{��3>k�nw����x� ctR����a90��4�T�.G��l+	;�l<䘓���]Ql�|�����jlS��I*x�9tP�ƈ���'����cs\���q�s�Rg	9� �)S��p���a�i�y�bmk"�[
	��_N�gS'�Kb6��x�Z�F5I�i��;�� � <�k_�6��i�NuT:H���Ӥ��&�i�O���Z�,�y��F��კmE?y�i�AiKZ-�����q/'��X�g����O���W&�1�Ւ��ȁKϢ���&��o��y�H�i�`��{�C���7[wh|��%�[Y���sZ�3�:��W�"�9�z0�M#?�����R4E!��-�ah�k��V�[��I�}D�I9�0Eɳsb����L�D���)ӨUz���>/)�7߮
#�7k�;�
X��S���)�	�yMD����y_���J��~�mi�S�[�����Wݧο�D[����%���K��
T
1&����R�$Q�S��'AH_�� �T֪H||�ZMf)jR˟NDhR�vT�C�
����$G���Nw���<@#���8x�?PGK�s��F�>��Q�J��}K��M
�7��"8�!�F���A��	��|�C�����V�`�����L�DO$�����CI���G�qB��]����G�p�2��f8��Ev���� ��$�n������ݘ��T���zV�9ÊVu4	� @�4a�<U������e���@�T))RR.�̭@��>>?A���
Ƶ �aB{��N�X��3K?��hJ�ˇ�#�)@N�����ޭ|�b�gd�W.޺*��@���n�z�*.�Kԡ{W5�{௅R���2�oX��j���kGDIry� u�X#��gQ:�R�)�uI8¨�l�gv𧜟-�s��A��O{mV��2��Z�(�\��tV��&ITV�K-�>h��F~��.:��M@�њ����#U���2��V�#�T�����T�X�P_:��:��g%Hk��T��q|�ֻp��,�u�m���g�$����@�l�~D���n�+��"���&X�C-Rl~7||��C Z`
�+�Gb����#$r&��Vԣ���&LvtI��]&6r����r�@��p�(�X�/]95�j/��ꁚ�0�j`ƒ�0
�M7��I����a����'z�]苧��5$�'�����ߦ~�����"�g�qW��աԒ��
�9�W7�s��q�-�-s
���`��K�?�ٞ�hL	T�� �k�HZ�K���j���!M�;UO ��R�J$��V���!rӲ2ܕ�0z��μ\ ��.�b7`͐`�}�q���_F���y�!�N�y����a$A�{�_lE)�yq��%���-5�g'Ʃ%�F���/�֛�7t4���q8vn#I)������\���ǷG:��<��*�gFSz\�����A8�3m�N���M`t�2���9�J>�O0��W��rG��7i�Z+I�(��E^^��S��k�rt*<qnC�秣�;�K�p ���ە�H�V�,�1_'��A���:���Z{��LJP��5ȭ-R׎Cyס	M�"b�~Г�+`W3=㼾����:�@Ѓ|���P>�~/���d5����;=�1.XN�`�u�����(���t"�uՓZ�q�8s\n�WK�H��ܶ��,�+*|���=�-��ԕ3�@�5#�4yJs�6���.�&���������wc����(M����X�:�T��[���i���,EޕM�����O������:��(��߽^���\���TX4�g!��� �W`��6�Pw,��'�g��+�,@y���:�tq<�Uw��[j;@J�&��Џ�YP~R�qň�l�<5���2�����Ȋ��U9	Թcr�`��p����gɵH�FF,y��Ĕw��A�!z�4o.8�B�O��}�vc����Z�~3h�2�쑴�sx�E#֛���Ґ,���ͦ-��1��\A8ѻ��O�q�d���.�W�`�N�����/�0�8���X�\�ޜ�Ѱ~�o/o�G4����^�0��p6�o3�4�'���K�pc?��=���.@�Y�4�e��E]�ϲv�O��_�	�4q�>N�,\nix*�7�Gk��<R�96�� #~���[�o[�O��X�Gܜ�S��5թ܎,���;��]5�m��0>8}��CV&�����$�A�C)g�ʃLR����Y�ϴp~�γ΃{���%�'�i�ճ,k�R�tX�{���@zx���(�Z�ُ�Y���k����3����vÙFyϕV���;������5pLT.�LO۱�K���5-��g�?	��Mk|,��)�HA���'�S������VH�H��ʛW: ��$p2V
��	��)���>v�fB�-�!3�<�/�����|;c�K�Ϫ|{P��4WJ̄[�b�/�@�cƎ�^,���'���2���-�$dƧ
�h��y�Os;�� 04� E�X��}�R��v������wz<ɗ�	.T���V���姃|���0�Z�(i����sx9�F��*�9�2f�5��4�m:���\�>S_&t��]�k&єh���yMCܒ0��s'�U��b�Z-�֖T>j�'�U���� �� ,T�/6��(�Jd	ƚ�b��N�3�D�3G�Q��"'�A����X¼��q�c�x�b��	��1~�υ�I�,Go̹~?�J(q�E��L�`���3�'�d��ڼs$; �
<�q�?�G,7Yz�]�>ZɳT�(�DZV
�c�Tݧ�����Dg�Ii3�?5����Sd�YVt:*,�#Y� ]4����Yi�J���H���:�%"Fm��X�4'+��f:;WX%���n�k�@�𽃜K�R�xS�#=�sV�]��a���������G��^��	��5!���D��El����!��1�����M*�9ߣ����@�mN*~y��,���@�梭eu�&Dq�((�'?�@��KY^�1���M����0���)f	��NM��
<�.F�U�
b�o٧-FC�-�A%�hVUxCѧ�x�K��tEj5�=�_n$r�YsE�jL(�BX����FM;Vt�$��_�-�����e�X�z��{��B�Q��0;� a�|� *���L������lN�Irzз�8�Bt;֥�?�<�KA9�����y9XV���zߗҪ�=��Ci����Α 5X_Fl6��&��o�CD{E+���?!��õ��@�&SK�Q��)�=-�EȄ�_Ε�UaԼ��tM�[VD왾~���=����3B���z<�I'S�>q��^����u&{�@���7�����?�⑇�P�l�i
��wh�b�ȿ��sF����b>�<�;a�y�U��VU�紅/�,��kL�gf]�����?��1��\�Y� �ߤK��
}�޼5Z0CO��4,�'t1f���#��0�GJR0L=l�h-����QXYlǙ|j:���Q��ƤCA{��$Ǽ������ݵ���C��¨-�