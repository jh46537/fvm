��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���q��՛������@�oa�R��Iz1A�#`�ԀP��Iqh�3��F�`�ҥ����c�
K4#����ge��T5��G�z�4��R��\3jU�;Ѫ.Xq��d���D��nmac��V�ܕ�;�)=�(?0�י+�k�襮=�%�YO������鏷w��>�s]��6�t�u�;]��4���!����q��
1�xF!b������.����\�2�X���`���~���4�k2Y�a�w�7=�E�u��#��_f�g�:�S|.�� �֞/^���J���,\*��p�#�0k�|
]c(��7��ȩ�'�Q�	�kR-`~���Zk8�$'��x��A1����Ko�� _'-l_���\��
+*�q�k�����V�LZ\?rŮ5�xwpP�V�22m��w�j�{!��;�Fs����]U�ӂt0�����Z�,xm� ��^�I�/�)�ٞ��O�]k�Y&�2��F!��b$�J��Z�d��9�����?��Bm�6�'��~;�?Ւ�ðq%di����k
`�꧊¥�4q��3q��7�$����~�' x��wn
�Vnz�cQ�o�GS}���駰�RY�R0� ��i�h��0��(�Y���[P�w�&�@�;���m.D��P�;�t�8U����U2t���|�ɘt->���^(��a۷}�����~М����"h�n���,�
N�pJι�G��M�H������|���a�0$p"�����u��NR����hZ�爈�<e[�4��ggW�Wɼ1ʯ��t�3fP!�a:�K#�W���	��zz�?A������U�Z)�Z^ܝw��Yy<�;�<ɍW�uj65���R|���n��0s�ܔ��6��b��;�݅DU*4�ż6x�5��ۅ�$�����8�¿���ϳ���Q�|��hT�҉&H1g�����7�
T��9ؒaG:/a��E�8��S�F��f�
�
9L߱��ѫ�1��Ե)U�(`�O7��X�ajF!,LO+�ǩ��A�q�A�O������~w	"�Ǟ�X���\�8!��Dtxm+��7@��<��l��I0��,�Q)<��$���rX5�uk����߮��й����c5H���3|c��\`Z���쑕	m�|�s�pV�4�FhU7���ϬT�Va%�/�e��m�1��>n؊�AB�'�>9\dh�1v�����%N�o@IM�'a>��;q�ޡ�T���[J��k#OO��e5XW�Bm�%4\y2��
i����(;���݆�G "��X��}��{��7��.  �4�mv�x�Ŏ�e�X[ާ�.�����A�ZW�.�4C��6�o�n%�[� �A/=#�߉�#_2>��e��jnU�_��y�%/��uTj�L���"�~��]\����Z���.8�]^W�r��&O *ʹ�8�Q���l�K�U�k?��G�Z_o��F��(0��M@J�ɾ��Ǟ>9&��N�6������O�}��~�A��,�&oq�'�N ��W��=��M���`���4��8L�]cd5�h�rOA���j��@T���RA����v����V2"�^��js��]{�2#�8��[*Y_;��aU��jʴ��Bp!|tZ�x�z��~�
iB�K!�h�)'h)�9���l�=T���5)�7a�߇I�'�_�#ˤqq_�m5��D�E��0��ŝ����h4��b=��e��3�"$�7�HM� E�]����<7ѢΟ��Z� &]�+��p�B�����l�s9QB^p�+��WlT9�|�(�y���o-��/�烅�M��� �U���z6m�g��(~�\��M��%M�˻=��%�R���oZ��}�bG��1����\�]w�s1M�_�?�!��o4;������3���}Yj�$F�C�B�:��NY�'S6�O[��ʭ�dU4M�\\��]��Ԏ�˧/�%f�E�3�z��Q7vGe/?�Q F`��}~q�GBX�L������;�%YĘh-z���֢ʑ&�I�z�0f驔�X�|OM��>�ǈ|�>� ��ҧQ��+6	�-,2�N�Y��ڢ��V�"��1���$�n��
1�����"��NU7��geE�Z��/G��S�H���wq4Qe5�9\��9��Nhʄ0��T��U���C7E0��6������3�u����js�<���M�{��m6�X�p��7�Qy�&MV���Q���@�c� Lʏv�O�{j�>-m�2R�9vk?o��2��,�������mQ�V�)tEV`}�i!�a���1�<s�_`&�У J������	bj7ۇ�J��2�$���M�Մ�K(�'�-�;�:�j���=?��	�bk8Q�p���G͌-C#���K����05uJ����&^����1N��rV�g�ƢQ��[�N��%R	�:ƉL�r(>I��;����ʊ�6Ԯ�~�[�A�nI���R&T�p{Mxe/'��G���P�S�O:#�0G�P�6�X�Iy�mIj���^��MZ��f˅�M%������ 4OmZB;�ɔEU��쐇�zp��Q�C�o<����E�ji�~��oQl��c���R�?��x��Ki���(:�y݀�0��6D�"���([9<~	Kt�Dq�Wf)��J��	�:��yy#/~ƍ��[�e�@��n 'йЦ����/gְK�q��~+qD��Jc��Xz����U��a�� e1P��z!ᡆ_ǻ��N�o� ���heȰ3�&�:��$d����%�[?B)��Z	@�EG�P��<w"�U"�7�L)z���Eb"�X�T��wE@Wϒ����C�L�C�9bƽ�Z�vľ���8%�U�ή�+�I}�0:SM.����`��2�]D�3��/S�U?���H�;Jxص��=��/��k`QM�7�D���1��W)��#�o������/`pT1�F��Wz�s�>y
��KzS���Cwׁ!����yq5� ��t_�}���)�·Έt�b0�}�PH�mv�S��"�z�@`��G	6JRA�x�{�.15���G,�6!P��x1̣!�;ؽ�������w�Ӊ9擪�b�!���������N�Yo�g�I��\�[��;a�{`#GH���z�>���C_���K	�y��v9�~|�~@o���M(�Z��j��fe
�&6��C?��uM�%�~s��Č_˦v����8D�:�"���@y�1Om�p�zIgSP�
4\�8�}�Ɠ+�K)�J}a�)N�`b�v%i��i����g��G2."�/m�����R�_+N5\x�#��SxRzv|�m�G�,ص�4o/�Ê!�_bHڀ1���p�Vj������57�_����tN�?f� Zk����M/)b�;�yl�"�K3�,ubۘ��X�����*��<��h�G��\@��,�@)g�y
X$��>�:�mh�^M8�X��Q_Ρ
��_P�����ڧ�p�ͧժ��4QK?׸��"��-���î�z{�&b�*o���v�`�lㅫ�_7��D	ee�榧(�ޥ$�b�.��=
7BL������e���+�soq�KӐ�N�&�B{��_�Y���^] �,Iߍ4�l����N���C�HJ������j//&�����U�'��eL:��9�Z�N����`��ӣ\����ЋwЄ�_[�!G�s��$�F+�vC���J�Aj�}!	lu�ZW�;�j�;?���p�}��]]ܷ��j;��� 0cz@n���{�����v�8���~�nk(ӊ��!�ȯ	�_�`�@"7�?��������?��4}x쁬.�)g�l�:M��6����YCF>����<GW�ݩ�]"��B�ˮ�Zw�2�Pf�SbxG��)��h0�*�0��mĉ����{v�O����䱷�M�ՉDfo���pP�����n��a�T./Ι�)_��흼uI��F!S_�;�&#YJ�۬Az���<��a��9��i7�m�"kj�I	20.q�\���P��
�ѓ��H�'�"`��c�{n�ɝ(�!�#�8ÕZ^IF_����=y�	㋢�`O*3��h2�$[y�t��'S��R���%��@?��b&<u�4���ӏ��W�M��_0�^4ݫ�Pس��Y���� U�`��:	�%�TՏ/3;����U�#�e��d��Z��wE2
`��!����=�~s���UH��OФ�sŬ�b~�6��M�t���IN�F�&���Lc)����F�)0Ud�S�_Y�� v2ˋ.�{��ʕR=��M-`V�_��Glr�ps��`�ϔya;�;���p�;�*A��'��e77��O�`ڜ>�y��-h�x ��@��\�&�0�����5k"�,��L��H�y5�\7x#�E(r+l���, T�����O{�LF�M)&%:�mpW!	Q�ݓWpA�>�A|����DK
PI�\5��C*l}����;/ՖEՙ;&^T1����D���8[x�ѹ�L�%FD�.*i��*� O�mlpq��3��
���Li_3|%�6�ZLd?�A:�HZ�]��F��M��"|G�dl2*0�ZgRbr���=2�
�4�]���l���^��OtL��~)NCPR�o��>��ZO���CjK��m�S!E��烑������4�k�ׇ�Ά\o�`�_s 7��O�1z�0!?���Hm�kVe6�Z��Ij��òa��q��S�I$���K��z�~m�[�;g�+�e7����/�,����E�r:Mn��,@K���v�Af�N)��)�e�K�÷-:ղz��2��=i\8��¸��R�W���#���9F�n%��%���c�E~_P���Nud�9��E�."�y� �q'𠺰@fsW����lqG���C6�D��V�L#J�۸Hq�YA <�'la�H*;�h+�n���k �=rY�y)({5v��̈́4h7���BI$'��c�ذ��� "=ǵd�%�נO�R��G���?,M���W�t��s�����/w��k�4�3�;]�3k�C#�ea���~8ѡ%�S�$�<�]s�����[��޼�P^�E�U�73��#���AJ��}�� q�!�9��ؠ��"q�����gr�q�	I��~KUh�%\��q}6#�7�>}�hF#�ai�<��D��60 eeCM�:��,dt�o$NS�\d�(l^k�t2�t]m���U��,2�a�©1W�޶Z��������]Q�_�՗�{�:������˄����/�x�v���8.�����.qCkE�
{ߣb8���7ZXX�32�L��b�H��hÕ��lIȮC��?BZ�s�e;=�ſ�fHYͻF6���������9�O<uM�����@��@�����<ӠE��W����No���vmyy�U�~�}[[T�V	����/��|c3�>�g^Y}'O��Im��MQl��{:�x�4�R�a�;)�x�^�O�ߏpn�/l��{�U�&ae�7��Y�;��9�iֽ',2�Y�ϑC:"1�gXD�8 Ը^Иkk+��k)~��d��FGS��dU�!��r���e؝�\8mD����!�)��h�- ��9�е���$�w��x�7O7�JI�$`e���m��*���5����K/|M�����	Y�8���hX#�8���[n�ܸ��S=$�2ß��&����5ni�`,b�?q�jwA`�͝�7�|1OD����ƈ��]��t�� �iL��?��%���Ơ���;7����`�ݤb8���t��+�2P\�ϐ�^I?���l��R�#�D,NQ3G$�R�]6Τq�B�q���"m��T���$s���د��B�W�.����\$�;H�z�NHQBJ8.��*F��)M���ȹ�ֶ���caJ�a+�_j�����]�Vv�!�}s-��E�x$��p�I�-d���,<���X�"�RJ�������U9,�s����6�6%]����`-+�D��,�{��~�&�y�.!�'$q攕ʮ3�)P��E������m��Sd���a�M.��K���ܞ��N�[m�e�[|�Ȭ�ǏtˊJ�b���oL��:)N�+1=t�d6�����
�JUC���+�����|��UD-���]�q�J�vD��r*2VX��zI �g"�~��H�n�\N�9 ���ۛ������O��.lh��M����4�S�xф�3pz��
qs6`�(�<26;.,�:����3�	���7�dO�lP�EH�ϳ2�a����mٜi����p�6�I���HMX���>Ǵ(lsQY�>?i5L'֍��M�L�����L�|��$�״�_��P4)t6�b�}[��}�*O*�����FB\|P�sB�(������1�i t�Я	D��ΰu`
h&��5�R��&����%�hp��g���^م���Ob�>��9@'���"<Ri��R0�@�_D��Q(�w��Tq��ݒ�"��Lt��;����jLb�g��頽gm`yD�<ϐ�5ˠR.;�%�ˏ�����~���W�K3��	�`��3���A��%�흉GvQkۻ��H���qR{fϭXb1((��D�uEv��1|8!l��������9F��`�Q0����W��ϖ@Q�e9U�Ib^�L���x�
?k�Ԉi�|?��X�Ab�|�O3�FHyؿ�j���Hg�J�����%D��.��?��C�Ԯĕ����;��T �)��BP� ~6�ZG^�*)�y��'u]P̃�.a�iT���7CocPߍ�t��}$��K��5��\ӭϧq�����Ờ�=��ab�0QSqԼ>�ap�͂�p]�қ7̋�3-ϖ�2i�<G<6u�g����c���\�_�J_|��;v!q�6 ���n�/��N�[�w�\Q���~������|�抅_�^Q�3�5���ڲ��tT���!����"��>q,��&Ar]�?�0�Z�j[��Y���@�z�	�wW���-F'��5���g}C+�#b?��)�����맰��ј��`�ֻ;
F0�OV�l��QV�.�Y4q[��:�Z�h@ld�V-@s1�� _i鏠�����R�۷��:�+s���+���������Dk0�,^w�Y�v}�5q���9*]�ql�Gue�|���dט���8��:�L2k��՚]z���V��_~����0����)����0;��p	� ��ʏ�E[�?Cf�g��x��{W ?���A+�JM��A�u̿�B����rI�n�I7ws�t-��}��6@�(��JL
�J���uM\��y�q{���nD�v.BU�&łt�E������֡&m昃���,Ҕ3F���x`cF�Sb-8�����8�-:���(�D����r/TW�W�F�v����w�o.�����Yj\��Jf���7/>�u�7x�x��we?69�t�,���^�MP��/�H�P�ϱ���#��`L\�I2^��АJ�� �n��d,��c\�^�q�/����#������l7`7k���D��Áu¬m�E��k�))XwxU�+լ��H Yj�k��Ņ}��{���(��Nm��[
=��=��K�<���&���M��B�M���R��`�k�JIC�4��gא��U��@�5�t��0��ƶ��8�^�O�y��yZ�7�.��{͈.��|�U�Ǝ�u�Q���|~%P��w�I��^�T]:�]X�e,ZPWF��{��K�c�XS �9���v��ۓ��
C#E>��%SM0Ѫ�vb;���m����vn�b��FgÖ
R6��	G�fr�{7"�Մ�qw��w����d:���L:ߨ�!�.������t�^�A�e�0�αq�^8^���V|���7iRot�T�%�������J5f�ϻ��d��-*9���K���v��7Į�4k7B�=_��om�����W���Y,�*$�#�$i�K�)H���,��O$���?�lt(��p���PG��.�2�-"畲����~t�H^"U�������WA/�"6�bX*�!$�iS�a�w�_b0�JYwzj<���ƹ����|kEJ� gZQ����)�JPE����n+�����M+W�;�:�іw�sXt�]��Sml�k���v6F��i:�G��Fx�ɓ֋$a�ߡDV��,���r�1�N�R,͘�A�^�
�B�����\_u�(Z�mZE�ž���i��AUc�L�0�����qJ�=�w��o�b�J�	��_�QXE�'<�ñXS;��f�p��$W�F���5���ïc3�U����s��W�ݼ��(�:;?�IҞ�����pby�[����{Mۘ���?�$%r����p�Oj���ι[u�Bv���~}g�gȱ�:yj��4R������f��<�p��x`����1�C�����U�}v�B��3�£����(����G,���P�O,+H=�e��I����|���؜ +OUa.����:lcy꾧�C�~�)�ͪ����H�-~�+8��F��_)M�E��ڝ���B|�S�f���1L�U�듽�%�*I�K7�m�7�]�T)��7����`S��eâ��F�	�7uC�S��7,��N��C)�ϫU���_���p��F@�b��~
O��
��Ak�tBA�j ����C���MX�H0�ⷭ�F�zPKzr� �  :�Uo�.]��%��AKr����6G�Xg{���V���wZw(Te�Jը��m��)����] �P8L��N\�9hzI ?���.�
��x�g+�V�ӭsE�]�m?�*{������1��Ȗ�;���Y[����T?Z V���s�
�ɾ>IR�j���4�[4_&�E�����Ls�D�`\X�/������S�I�zw9������^������,,c��KN5��c4����*4'�/�<6w��b��?��:�*-Ύ��|��%��'!��a!��$9�����$S��{O)�X�7M�n�K�>iy��{�����̉�������5�N�L͈�=�Ȉ�Q�&mk;I�]��J�\Y��o��x��?1c>�N�od��	�ێCN���x�'���2�n١�/J��3|�[�^ WQ0������:�����*|O�8T�&1�<(������E�����v�D��b���A{ʖkz���H̍�g~�O����1�l��	"#��y!��̥��hQ�*5j�I��I���I����0K@�'��*-�X9dP�/��g�	�z���� g\�A�c�=R���,�T�_>�%�W�9Tj���C��M-�P�~�Up���R���X������'l�lI0�3Cm(�=�2von�(�3�m#TLG�{�F=����a-(1��6�����x�%M-S�h�)ǥ�(x�<_`/�T ϕ\��m���k!��;��T孴���Y}���6�޴��\���~�,��A���+�^���|�$+�݋�3}0!�:����`�SFPo�P�\Q�R�z�$������gW+��S��ZQc҈-?FLq��f�j���-���N�nWC|�d�<ā�~���_�� ���{���Ơ)e��� ��@y�Ϳk/r�Hs��l�R�fRJ��S"d-������wh~[�ZZ�� :XMg�/��7�B����*���s����}��ž��;���� ��QГ�����w�#� �2���H�a��r����K�'o��G�`��n��g>B�W��13 I�1��|��������@�ۭ���YbQ�Ss<ڞb�����3 Q��F'4X��@�*@U�Q_��oGm� D��
7O29")�U�����z�������	����g`�D�xʟ�-[O�;~�ĵ�.^~0�c`�7�wd��N�LG�U�c���(:�C�ͳ�B��n�]�~�nޓ�p�O)P5�o#��^��d���I���w>�b�2NO� bG���U��f��k���R��e�ʦ8%֏]�����uY���F��5�!g���$�w;�����5���}Z�NۂVG���m	�SA(�&zp�P��x��+My'$$�Ī5/�Brm$�� �\�
��kG&��3�|�l%�������.5���l���Wq�H�0������у![x���qK�3�X��)�=���z�JM[� =�~��F�F�����̻�M2�.�����fZ[���R���m�o���"$�����z1ͱ����<f3+����3��J��oMSP`<&mL���7[J����6�i�d��ƒ�YW
X��.��p�9�N?����M<���W�p�1@��������S����G�A+�q�w����jhe�7B)�Β�ҶМbG0��e���CZ	~�*P���'#�@��ɐ��¢�����n#{��H��F�nRq>�&~]�v0��c3��å�&��4�ofJ2�C3S�舯����'\��Eh0Ǟ��Ʊ��rp�wx�p\��G6��T͔=M|���Ш�+�f,�8�h�ѣX4o�;)'*h'&�T,�����JU��M�c�{�<j��f:���p�"J���r�މ�W+V@]�e��\��Cc�z�g*b<����i��󽄵�`���"�8�� ������sA?X��|=X�T���6���`cĿOE�}��V;k�����U���&��β�ׂ.�f�
0�a���p�E�m�`�?<�)>ui�����U�g8��r�ө�Y�X�T�zo���}����O�����J��x��F�QJ�����LK�";�tI}mW�M@�����!�Rb{U]�ž�#ܪ��Q�����Jʼ'YzF�g��Vjڬ�/�>�8�4������p�A��7G���H��*�L66#z�ѣ���ԭrg���r��z ��a���HY� P�:�D�)�����Y4�ޜǃI{��z�����?�X�W~���P��uX���G����<�M��8jr$.�"�a��A��� ΄�`�����J���Z:�!A}
�����JfM}W3��u�B����DK��G,a�z��]�?�~
 �_ʪp���7�j�>��5-�Ϧ@T�Sه6=u��(��A�{J�
˰��-��a;QƧ�xy8G�D�oKso���Tt6 k[l*5��>p�t���=^��q���v�:��Х=V_pS������z�����n��h%��>H��O=�5p �A.'�l`��I(mA������|�Ѫ���!`����	m��I�9��7n�A�ڝ��g��'�cq�.�GHCNIʑ�v�{H�
$%EK(�A9e��.S=]dcn~���u&� �4���[��,.�v��J���S��p��j�������9*��'q�N���5����R������%�cgabd�- ���M�r��)�ɕ����v�BR<��i\!�ۨ��"ͩ��׋S���"<�Z
i:����s��?��ˎw�.L�.��W;ν������I����&�g�=�&Zc[�n�
f�F���in��Nj�ok_�w�lD�ӑ'�%�v�W�n�A�����0��������B{�_NF/<�h�������a�tNt}����Q�sp��0��öŏ���R���޺fQ�O����qž����g�l�8W�����g��uF�UԠ�BοW���SE�{�窻i�~�_�-��p�'�sI=�p��YzA��ϥ���������Y1|�@�����$�������m���(%�9��(Tn|�T;�%�s$Z�k����]�����|$G��.Z��z��|�s'�ôn4u#}���PIsݔ1�
���|tX�9��>f��	q�Uw�z�D�1��>
B�����nmČRt���q�E�ΣQ�����N�����vD�P:,���\g\��Z��c̃�-R�K ��D����W���m1�B��5\o�Lw#2b��1��3<	�{���/J��!�!U6�9M���`�\V��C��?%7�h��'����'����o�&��!g��h*T+�Zg��R�ŕ!��3=���� \8�B���E��'��P��jg�"]��Q���ߧ.���E$my���I���u�Y����:��R=U?�ˇ8��4nA��jT`��[7�N*��e��*k6�2&(���O�YUERҍ]���'�r
����H%�2�����M�wD1���K-�Z���t9gd���2�� ���v5�Z,5���!nS��C�0H�0Mu(yv8�0C��d�� �I���
ٔ,��%8�'�/qM\�������~�KI8���;�P�4�FW�J\��X�f��@[�I"�����6l�ciЃ�����\�����#�Dӆ'Y��xq-�S�O)<� �W�"r�v~�@���򽗡�S���*�U�������=6Qbo�[4I)ߗ����Q�j� )`���vYY�+������o��D�6����9�c�GZ�
�|:������G0�B�E'< Z5��>{�����'\�.�W�UP~S$4���ط���m��s{�k�%��+"CH;��BtR������`	T�d�|�mZ�N_#����ç́2�(ftȷ��a��q���R�5����b���X,��C���Oq/s0&a;OK�'2�6��RJa%e��0͌r�|�K�ǳ�MA��k��p����f{�o��Cc؏f�D�otI��Lx���!=�&L��kv���/�4*����5>p@�Y�)���� �%0 ܫؐό#_oPY�E���a�j`��E�Q�8&��K4��5��H�ftΌ��ڲג;%�����L��ޢ�L����w�"df��I�$���[��z��Ee$J6E�`����� ��1�~�2e��x�ptM��r6Ud1+�?��	|\�K���Z� �EP����Dv�8����#r�|��$��
Z�X߫�^�7��)!�Lr�Ք�j�VoԠ�4[�Q��LiB���Ok6-l��������l�]bܢ�X����o��B�M7�\�*��G
�n�:T{	'�@=d%�.�
{�uC�V�g�5�"����e�o/^��|�X��jy+;Bk^�"����:�ɾ��7�`�ײ�A��e�Viw�!ı�H��;m[��wj&>��L���|������|�I��/O�c2�'�I>�p�+:<����ů5�� =1�d��سŊ��OG|v������h�c�{��ᄱVvȱ�Go�,���l�j�?p�e{�,c*p�ʸ�I�bʸN�C�K�=�	�0=d�Or��/ڗ8����;��
�]���IX�W��L*0�����Q�ms�+M&pάqܲ��W����l�X~��
��&z'.�U��x��" 0^�e�[�I�$��j�n��m��
��7���5�tڠ2w�qʕ��p����)���^�T%S����*�v)E��7z�5��g�-Em��6��|��F�T��
��'X�<�1�B����	)h