��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k{de���ӱ��.�|�2n���Hx���]|��3?���ZQ����mC̈́�8t�m��.Ԡ�IY�����b�\���}�o��׎L��w�Q�|c��i�+r�%ZGz���룅$1�h�)�4�`U�@�v�/E(\��~���� j�rZ�,d�����3,�_��Ⱦ�A��ov�Us���w	��Di5��Q�P��uqX��^	.�u�~U�^�.�k��G:[�A���}��+s��`�Ճ���h9��:R��3%qd�{_H�������L�w�(��	��e�T��b�~ӡ/X��.�/���Տ�R�,�o�����U���N�W���m�5��9�s�������S�=��p���s�*Cb=N�J*dq?f�@[}��0����.�Ժ�S̩ �C�^�s� p'����eNˍ� * �V�L[)�S��o�6����4���!�qfd�#8���]0�.���UƏ��b6�.R���"�|h��?��t��)ѐW�������3���W��2��n[�<_	�d>靄HLX=������v(���$�9�]�7�Ob�����{|����������Zp���\Y�ˠ��h��<� i��iRx�C�%n$�Or����g��hĹ�٢D}��o�@U�z�@4��Ԝ��R� ��\��d�L|��:��)M��L��t�@��CPpW�
f[�p9U<>a�Y��·�����E�cd4�����r,�GA	QJ�f�e��`���[����� �s���I���TC�)���9�*�&�L���
�,��ӿ����7���,�Ic ���PW(�����>����5�y� #��r�l�(|�K�8�<8��`�FI��D��U1�$�ì����ĮO�D�,K�+��Yw;A����0�����Y�ߏ�ws�t�fo��%g�7�Z,���m:6��-���6Y�h3�}�ܿ}�PA9%~�pF"M�Ow�2�JY�ރ��XXS�b�H�NՃ��ĢI+i�2r{*�]�=K$�f���r/�s2a�&@~[�y�ص����2ِ�� I��W#)ʢ;qe���N�(v)#�7N�Dj5@��3�
�)*I������]�VIe�p��q`q�R-�qg8A��)�*,�U߼�D�~�C��t���;�<�P/@9�OT@��O2�o�/I�DXHX�K����||��WWȫ:�� lm�YR�s ���.AW�?^Wت!"���E�@�I0�X ���n�*r9��%�M���ݧ��E2���h \�1DQRI�gO^���Suc�+g��f��$
f��[��Ŀ'?Y��ήk=�~#�c9��ƭ�APnU�j��]�B�e�Q�A?�>��44q�X�Ȇ������I�(��N�2*t�mP .X@,�ZCV�Dt��J��'�80�JK��&"M;�w� �q�hnz,w3r?�E���Ho�e�q ���4�k#Ou�Y�ȃa���{����T��<v���oKZ�:N%U�]Em� ��D��H�u�z�hzo���HJ�.DV(�)t��׾U�L�q�
��">2�9uT�'��:.���:8|@�j2���b�4��'޼�3Z���n�Uq�����)�p7`�kl���ã�'ʴ�+�/���"1���A���3?zg�7$�$0�g����1Z�&Z�+c�y8��� y4�G����a�^�����������z�(%Z���2��2��`fC��,���q�@�R#�,�:$�=�n��2�u՘�|@Aз�w(J�����J9����b}5�V��Is8���1��O���24Ӑ}c�&l�جFs�@ť�})�s���#X���b�%/#h��7�l* 'L4i�^T{�Ԇ�<ߩ9��m�z}�Qq����dX�h� X��|-v�6�(����8:� b!��D�H�F�CV����I�1���T����'���Q��#�@n��y$z�NѼ5����C����,�2���Db>&30�r_������&��π�����Jw�<��rmk�ni5W��w�-!�M�_К?�#2�J���&�GL2��Si��B>ͰZA�M�*QT����7�;~!nP�	*Q�y��߄{�> ���:I��&��Q�����sS�|L��	��C{���PZ�M�$u�q�(�K��n0��YLe`�Sp�:���h�5Lg(����@Ԯ���C;DN�2pmQZTM����T��̐^A�n5>�c�(�� ���R����ӏ�<`�S*.���t��t+ץ�K��W�yq� }�/�T�����וo�^�Zݔ\������Iv�hAc�Z�����������V��
����8j{Nm�q޷g��Ց|��oo��G���*ߚ�ԥ�ܿ<�p�N���[$��#����IӀ��Z��	z�)@��Ύ�����NjW#ɷ��r��8O��֭g�A��ԥ��4���sn6�l��nܗ-%v�Բ7��������o�l��Wj̚[o��=��#IM1��A{��ȞY���:�/*��
1����Ο4^X��i�����"^|s�L�����5�C����L���Rč�vuLs�4��IS���`_��g�K8���R��_>c�e��Y%�~Vmq���GE �i%`P&*b�C�'��a`��҄p�
A81+�h�މWQ������.Zס4�נn�|W_
\��n�d�@�:$��-+Mde�ŗ{Z3>����8I�6jRd�;���J��K�T�vK��ѭ阿�u��s�E�Mwj���9D��l����,�3h��u �,p�����/�O隉��@�'&
�&j"�#�B��	����i���A��p�XGcf�G �I�8��bQ^����hZr{��?B�s(���۾�^�A��j�U�F\3��6���7��,B!^i��]��jq�D7�c"3�]��>�	�I�*}�)x�E��-��m� �mƿ���Ǎ6�%�ND�[zFI3�!LQ@/������zg�8*�s}/�+s� �>&i����}�W���	o��۬���n����Սf����歮���	\~���_�k��֘6S�Oد�����	���}���~#N ���zsK`�H�˛g/D#��1�s��
����R���	�i��!3�Ī����*H�l:}O���?�\�ۓT�s����'�$��ez3G��N�5w0�2�����ʢP,��?�bd~A�i�g�RRvۇO�~�{Q5������]a-$7Ѝ����繑P�h�_�\��<����نAu��Z��9R�;�6�L�4��@@RmRC Ǳ�g�����x��$� I�B����P��v�N�h���2A��eh�E�iq]�A"�w�9t[�a�}\��6Q�q�<�G _ߎ<ԥ�3m�x���5��d7FS��Dh�x��i���!�Ա�7��'�6|��`��q���e/'P#We�m�7E�2$"��+RX��0�����՟/���Ro����p� ����N���]����m�>G�]��Zy������"�2z����&���N�Zuxh�Y�	t��M���r4!Aw�Ql��ǚz�d�pes����ODbht��?����7D��#=��2ʢ�pD*5M	�Ƿ�f"?H)ey��{f�R���Է��S���#����SHά�)�ZH����g Ϯ������D�ꭰ ����-~�f<5���ʢ�#H$�{g�!+���%���T�lq��*�G��T��*��k���E)ZI$V��d�V&	ݸ���Aq�&�M�<��Ҝ�����߀ѻǱY�VJ�]�td�!����l���\V�[y�(�픗DP҉�Nh�hJ;�wz���U�|7(sO��*�	�.+s���k"�EԒ���ei�~��T�*�"D��9�*�=0�P̕��5,~2,����8�iO����v��ӒĀ����5����TiJ���Ǽ�W�M�%�� R	^e�j�>�|(�I��*�^B ��YJ��v��<`ň���f_�f��X�O$C�ŝ��f�|�x��O>,���ϊ���Z��_��~�% ��,M����K�����ܞ�v^�yO���QLV+ދ���DK6;j~+�C���<{�S�q	7�a����7 ���0Jf�th��g��F[P�v�*�~���[�&��|@8?4sT�B=�g�.R��?���$�ql�R��3[�"��+&�>���(q��r���n������%�|2M�[����|}���Lw�fe<�$(�P��O�����B�����io]RJ�Jwdl�s=��Y<t����&��F��7ɼH�$��)���#��&�ϧ���j�q��i ��4}���"��c,,����չ+R�êlA�����JL�R�R�����L-��4�����m�}GL�n&|�ࡲ*����������N�e֪N� E	U`���/�DA�J;ѩj�Nn�I^3��&�����6�����0�}�Ƅ[pT��-0���R�������2�/6(�J��қ�O�}:�b��rqq�c���V�@�4^�N��Y�kk̃���fS����J���>��R�1�Z�$fV���+~���<p%�)�Z@n\��H�g�f怫�.V}���B� R��|�����S�:���k�����x�5�Qӽ���+� eѭ��	[��h���i����re�F煢��C��g�|��"���E��7{`���;�{~���?��'h�>.�i�E�/MY���eB�&��L�/��QC:D��K_6u>���u��:K�J���?��{iyN��-~�U�Ǘh�*�aCDfKa��IP����k��#j�<Lt�&}�?B�I��9Jd���.��7�HQ}n� #\}v5�I�܊��S���ν�~���#r�k�.�li�i�<��IAN'�w�X�_�|\$�[6�br0El���)��<U�����L��[�F�1P��u�tF���ɫs�q�*�_LRu��,��;%�al��3J!2�ׂ5���.$��?I��{
�#�����rl��XԌ��E:��p���e?[�a �/��{�����{�����/�Z*�˂WCʻ�N��v��l"D}÷)��S�R�J��dx�|y��O����-��}��@;`\V3<{�d��B㏮��I�RU�Q�B��h����`�2�A����+�,+��
A?�`�^ ��՚��G)R5u/�����u���J�Q�wR,Xh%��v�) �мY:��r	�~��i/�������31�)(TYD	Î@�M��5>���J�!
Ò��e�����.-�:��v�G?�����T����I�������I����g�D�-�U�r0�*���(�1�3��=��w
�T�kq�a�y�y�x8��_���jS8�r��i";TZ���@7���Q�w�1.�b�kI`�.7%���*2�-1X�5/}k�yM�e���᫳�ª<b�Ƞ\~IY�<�Nh^Pۇ�:F�Cݿ��[�DĒOdX6xiTnmM��P�G����.^�Y8��P&3*�T����a�A5���������!��&)�/�'u=�]�;���P��C�x(�H"���A�D���Y2��ZA��o������H����ZJ��6+��b q��(��!x�v�3�m:%�"��@��O�m��^7j����Y�5�i�<,-��e����L��c��֎{��vWN�S���֘V�g�N�!4�m��p�`W0x���4Aݨ>���[�Y�Kp ��n�l>�� �袭g͹��^`�_�j�V!T"Cn�F hԧ3Xn�[��s��(x����!g��`��ʯ��������az�Ǳ`������I9xjR�!��.+�5�4�)�q��V��Za�ц�GW�-6E�<��?|z��?¥h��$��Ӯ���p�ώW:Ս�r�3��׼n�o�.Y���:��#3�h��.���Cm��2u��B~�@��I�nS(���h�ϳ(>�-�1=T�2i�Q�0����X�4�Vɍ��vLJ��\uώ^ű��J��:8��'��b��hw�u���OmG#l�����5H���v�v�3�;C���3�w�����c��żq��A���w@�Ʋ�<��N�E���3#ܞ-��[<�s���w�ֲS��2N@������<HFD��5���y���e}�Ҹdٴ�ٓ���О.=����ޡP:X���{I�4	��;��_��!�*�@�O����9A�uoN6�x��o��[�� "-��as�k�`���>�f��#�~�V��-����>�]�5{�}��x'���*J:�Q��[C_�k{c�ٓC�\��X���[5�E�W�:a�rK+�6��3C�l����q���5�E7z��Y�D�yE�;�Y��{��v���%3�⤇�d����PM2hBb�ې�V��������xO�^Y��B�)�l=�E�t͂u=}2F���O0n��d�'}�#Rl��fyG}��V��Z����U`��u�1�,ʔ����m��fV�C���]���j=��JΏ��B�h5� ��<@�}V!��s�o��̡���ɭ��������0JL=� J���Ǆmz�c��¼l�$���Ǒ�~ ;%����B�o�S�ƥP���� ��ꘀE�}F*)/z���L�� �[=-5t5�B'�v��z�}�����`���p�,0\��d�MuU~]��ꏛ)�������d��w%(�]8�IY�pC�P��*� ]��e�i ��'r��v����{�~0P�dt����x�)����R���qW�\K��ŉ�[�p3�Ns�S��#F��c&Dd
j��k�bC�9�(��M�J���g,и��/5��iK��}�輓b�M�k��D:��^D!X�T��:��双v�Du��t�����?/3"<�4-��	^?f&+�)`w�2�t�GTҶ�[8^�R�:��D�CD:=y�t3�� ��(��d�#���Ld���hhT�{C�bx��i+n�E{�w��;�e�	�v�[y��޸�#Q��ɮ[��%��w��������U�E_���"rڊXL�D����HEEe�t��"�Z��P��߭x���Fڻ$ƹe��o����b�7��u*
9i�^�^G��|�o�%��y[���nᕏ�"ˀQ�<
�ԈKnF̠�	ㆨ�P�����ߎ������_;�%��[(Kp�A|�E��n
���7�_������M�)ɝ(ε՛<|��*b�h�K�)}=f���s�s���ع�ށ)���ɓ��N�5������2�
�����;��)��t�%���G���1�.g��<�Ɉc(��z��tD���~4!��|����.��T��H$���\pݴ��X��F��5F��-�;���왒S�6�l���3x,֛1&z�9��
P�P���8�)�;�6��S+�T�ΓM��,aT�O�)A�rXB�?_���V��]$r�lL�6�΅il�~,��6�������"�K��V��$�O;�[�׻�5��g�g�,��R� ��x5�/_)vG�y\���0�ɵ\�.��"�Dj���S����K�Y�S�Np�,&֮Nx��È8Ac�U7�5�w�B
w8��p<��~�ϫ�9\	̨�� $�\X0Q$ï�h0E�� Au���G���wyW�����?O���u=�P�N}7����Sd�H��gP���IB�>�x�_�� ?��k���b�xʑ0"O帘A�Ĩ�&�JK��2�)�v 	-��tSa�^Ec��C�GgE/�q&���K7�
��j��ӈ�O������,���}!�������s+��>�\�|�,�x>�{m{*f{�{V�1���V�~ʬ7��ꖎI~vH��32ubԼø-?��0b�OsP�s�}A��E��9Qj��2 Q�t�֊���>�E]�Q�0<.;�Nd
�'��6µ�r싆*��ۄ��\�ϩ"&�Ҩ�F���cj�N]�'-y��v�B��+;�Eb��:��>�?�A�Z��$��
T;��'u�yb����,��y]�5/3h�'�)�|