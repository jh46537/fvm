��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^��,�~{�q�E��	YjpA���zm����4�]� ��|-�<a���M:����x��G�^�\��w��ϩ��}ޔo�]�H�xzȴQRQ��j���5y�v^��
y����,�Kq��~vx���o^�yP�T��ۄ�<��P+<��$�t=w�V<dã���󰂝툞#�<[r뵋:jd;�$C�Hz�MH����7�����<l�P��̲���N1���DF�gt0����*)e,����x0��++�����j�?)�^�T�:�k��X>~`0Y�n̵�b��
L:A�*�}��;Vh��!|�M�t+���c����p74�^�EŎ�a^�vb��X��Kbdj��	TO�%Gƫ�{�;D��-�q��O��wJ��Ȟ��;Eâa5?���)���GY�C<]Ш۲[�:�+>�m�35,$F�`
�EK����dotT^�g�Ι0���a �zV��D
s�X;���rO�bW3�AqC!�F�b�J ��֕;M�n�?���
�g�L�Nҽ����%��v2'8�����oN�U�:���PVB��}���7=��Z�Ԗ�bmK*���Ba�d���H���5���**2T��eE3�Q�_"|@c��x,W|д��@�@��k���Гb�a��D��*}�[U�-HU�f�cE���j.�A�,��:��[�3�w}��.,WΛ��-a��������v)OY�C0�a��
&�^�6xRo@�z��b0%���/��Q�^p������z�8#���Z&���x��+��$�<T�^��h�هR'=� 3�K�2����T��Qt���!8>���52��@Xy �2yI��q�/v��sx��ƃ�vi�6�=�v	� m��������12J;���ONKb��XD