��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{T#�5~e ���J�	)��2Z�Zw|h��i�ͬK�OǦ*Er��G1p��綨	���7E���G�eU����R�t�y� ��42��PD�B�狼��i��M��`!�b8�d�`�0��b|���m	�$n�Jf���9��^��FŻ��PuPIu�����KS�q�!�~���Q��$R����?O�rz��Y����ʆ���l�˧�a hbT7�&8zWZa���;�����@!�Q
Gm�gcz��3�?3������]�G���i��P 4�����ޙ��/W�0�&��d}��^�k���_�n˘�4Ov�Y���-�L)�U��n���rX�]o�W|�(2*���9��r�͉��+S��I�|?��<�"8�b��x�z�\+�I�9.PVW��4�]�~�0t�b���$U�S�|K�vN���Hv��4�'f�b,	�2_���qӮ<�?�9���ñJ%���uG�є��������W�q襍˾u�w��l�ۚ^٤}j�����Q�Vq �}m8����b\HG�t���p�ov��T�`���L7���!d�FȌ��v��ǫݐI���ϙ��p�֪�N����H��)�:-)�����  �7a��u�ڔ�+��t�3�{E�z��ҡ��z�R0N��I�e^
?~"b�\iUYԥ=�,�r��)Nx��Y|7Y�u+p�����n�	3Q����5� �����┹X�SH������׼����0�*R��\eL���j�\g��(��!B%���u+�/k�ǵR��8��+Ӓ�mT	����܎��F���$���� o�D�Y9`=r堧����2}ފhx��jݰS�ڀ�	�"�ue���F��n�s��j�cN	�����t�9�z��3�Ni�e�2O���$�7������Ju�.o)�=D�n�?���{�����:���z�p��2]f�_�Q�E^����o�b��l�+�#�;��O(JS�_̳�X� ��:M�O6�id��Y�2˦�v����R��'Iq�t�q��O*?J;� ��~e3r;2���|�P�E��<J������*���o�Z�]�����Mx�*�@�q�V`E��2
)��`�����?Q�K�c�zG��]?}����4ѕ�CT���i�Y��MF�td)k��M���.`#>��%��E�
�.tU�W���WJ�F�"7c���g�PU%�4��9���f���Ii�\sƤP��|q]����>h�8݉�[>��_)��v�!����y&��G��<(b��x�5�P�����aP/��Dow+Ѻw���$�@3��@�祮r�cI�Z�v�lK�;ς�ӓX�f޸9��en�9Ajl�n�%ă]�P��ED���I�ӛA7���g�SC�7���r�'"�=;��D�%��D���\|.݊�NIq�pK��<�e����ю��(z~濿��Ĩ���}4f4U�>�t�"����w~�g�,�Z>�3� �&@A]LJ�Y��F\x��zi"#�5��FM	�x�� �oy7g��*�0u�)�ڈ��+�E�;ZķQd�]H�;G.�
��?.,�Qi��N2�6�>P��*}�^�kd��X���5w݈S.
&�ѫK� ��<�"'e��ȋ�勍�ʮ7'��i�s�h��)�pd{`0JU���\r��]p�6�7�;LTv�{�l~��d��Y;�N�G������zm��X�]��U�\��#�!��xXY������K�k�nK�m�[GNv�#���>PF�<+Ӑ�q7g�z�p���Hl>����T��w~V裨k�H�P�~�H�s��ym�:�u`����H��&&5�|p��|������Γ/1ĸ-��L0�^4��YRf�dP^��w��e�CR��a�-7m<���n�1e=��(�*ۤ	^�%1Z��3����Z��59q&84j����)���/ێ��,������o�.{г�"Μf��V}�p�
�q�<Y�����/��SB�f��n5��p��@c|}
|�
�h�8 �gQ��bH���݆D(�,��
q��"^N��p�M|.�����q������ϝz�4��8�ї�iW0!�gaת��.�ܔ�Ƙ䌼)eǇ-��:IA�\��b�������#��t