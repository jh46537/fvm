��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��!N;�?'ǝ�{9�1�\��,�L�B�8��V�R?��[6F+�+�4"p���n�d�#�$؍p�����.�{¯q��ěW�F^��A�S*��|��Ea)��sz�$��O�+�d(�W�n{�|��C�:� O��U荈PjZ�h�'#��}�Z7��-?D����͈#�26���1�o%3}V�9M5@�����s���F��	+�5�������S�/	��;;�~��g��JRyyҩ�M�'������Q����4�1_A�<�����E�s������?�I8��6U�3[����[we'C	�De��m�!L�����;ܜ0��V�~Ջ�r|��˛a�1X�=��
�M<3��(&�<�<���U�p�b��)��+1��+�����=�	�"Eβ�,�������pR�Ry�+f߮2j�۞o

�,>��������wX��2�:D�J ��� ��<���h�S[��h��-(��(�s0�9��5�[t��s�Lm�����S����f�fQ
���3��?�$7I��Vٚq*�T���8�!yxɕ"��f���&���4Y�v����^�re��F��������]���g��D���?��EH���2SM�>ZT�Ӷ����k��ֻ,��9p��3��XoS���,������vtD�S�Z0#���:0��8��Bk��{����7��e�ecQ�6~�|��/��8������y�dgO��4Y���S�`�_�� �8|C����6 �N�.���]�S=W�h��5_ @�WC8��#����d���.'4����'5@4�{�;�&�K_Zhe���������������_�3��/ħ�����G�~����eA����	=1����0Uj��m��3\�'�M[*�Z��Z�Ɵ�W>�Z��p� �ۅh�T�ul� nl��"�G~ ��Q&��4E:2�q��2�E������� `��T�dS��c�V>�/ϒ���6S�<*:��?$c�.�[ڟՌ9&4��K�Lp�dZ��i������}\~�@WmA<�i�2�@���6�����ۨ�׶�އP�T��{w�O�m��.i���s��|��8-�'6�.^�UzZa^��l ��UT��B΀?�4y�N�ຌ)�F'��Na��n�'?�ՎR�,��&z�CXL�j1��8�z�����k��@>�"�DY�qjz�7	6Ep��oc1��Gd��i�-�h���T�����).�)dBL�S�uh��.zqx���U��Z�C/B��8�!w��� 3G�0�_A��F�12����k��{�Н/j?�3_�l鬁g�[��)*Pal��-=��!ʜ�U�2Ud�"a��~r�ݯF�y`��%��А�+�0.4��Nۭ*)x��o���0ĭ��)�4l��'�I���N��E�������Fݵ���C���ۣ�J�����%�)��!�V�}g<�o�ҕ�y���&�xx%�ܷe�:A�}��j<���d�۽R�C��ra�{<=4Y	ͩfx��J���8=\���f�k͑쐇RD�*�)��#M�u8S��0/�M���q��{-�(ė"�|wS�� ���� u�yi��2~��O?��Dyh��u�:�\��HP�rx��8��]
ӓ_��g�.���/�i�݉~]�	}�v�����(C�i*���i���g�f�4G zG$�k�5����[U�|��z��3�"�~��@�����y�/N��c�/6�:���`��A��Z�+��eĕ�/O��&�p�d34�������3�[�O>wąB]�u4�<=���ޝ���o�2�p���l�H��@c��Z��Q�%�#Jx, r~@������A��ڀ�ւ���3�V2?b�	ug�t�*����X�����gpe	�"S��=KP���/���_2"aK�ܖ�pc�$`e�$��D0�L�e�.�{:������>3af���Ý%x���TP�P����9(}'���H�<���6�>,_�&# �p���b&�գ���E듪�K���i�l���	�*��k�i��ei1E�p���av��b�
7YvG��`VIN�F5!�>Q����8/�ep����9����|���"�/=�4��Ք�ӏ�l�F��B��t~�A�Ɨ a�"f�������H��h�ަu�t��* eW#������ ��}�Ѽ�}�o#�Ka�krkh������Fˮ�3^U�)����m(���K��aŇ�bGl#s��8��c��"J:�2��Ȱ��/нsV�	qD��~�io.T�D� O;U�-�X�!uV������Vuc�0X�}{]@1 ^J�ŏ���m|��.)#�_�D[cU*C�C���$���R#-�����2�����^��h���_���<��ݹ�d/��rn.�!D�.|����Er|6t3
��:n3i��G]k�����ȶ�2�E���ԡ�U�����ǉjϪa�����{K�*@�#��P��7`-f�X�����B�e礝�H�Zw�V�׊�'��Gvo�5�0a
��x+7��h�BNl��\�D�v���IV�N�-����{?�a���@^�@xE#�L؁
,m�?��>X��8p� ⤁��-�m�S�Qd#�̬Z��^�cc?�"�AGG��@�EͰ݆-�I{���&|���#�v3�ϼ�]'�&۬��a���u�ܫ�0�G��W��eEa�.]K>pX���((�Q�)�i�14M�]#��1?��]�����>���Vi�CO�J荞��ر��������\����v1@�M_���B��YĤ�Y�������?�5�p�*:���Y�,,���ҡ�>�6�������w	���S&�7��<Z?KI��d�FZ��6�� O�e�"}��@W�`�\@��5���"����$O��d;e_(�j�Qh���j֘�7����.w�+u���E*(c~���k�ge˅'��Y�HcJ+>�P]ߕ��Z�GSZ/�vRH�8�_ܝ���'9�=#�E<]��Uv�H$�X{Re�8����t�%H�kt�`l(mn(�	�^a�&��[�:A�$}�?�j�%�aË ��:�4�����(���PH�[���?D"jJBD\��?^B�X�e��sn��f��V��٣�j��lE;0�ف5�0|�H"���坁߲-v zb8 ?���]��	9����7�#��h