��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,V��`Sx�@�^|z�Ȋ�ݥP~����J��j�"V�bEQ	{�k8g@&�&_j�����J���*�]��U���hN����^B ��wN���kQ+�Aנ'�zXiE�f�]�y��A�f�ZC_������}��|O^�����oS�M<��EF¥R�-�Mٝ��J�4ơHy�m�!%�cn�fؽ�%��.8�t7����+E�ђ!j�-y���m9�R�^�G���M�������Ì?������m/$�X"�Ēa�X��7a��p	2k,�*9�W�Ĉ���֦�m����Ҫ���p^�/���{�=C �x��v":�4mն������q���5Nb�����D�-<��kh��pSc��YC��kr�(�ɥE.ض���*� �A����>}t19m~7G�'T�'�{�~�s�76�Y��3��ec�&G}�WG>,�\��P��Wr5��ӏ�2%����pt ��j�A�����@ .i=�췏!����b{�����@n�kP��x��2��<Z��3��	��Lt[�
Ei�4�4��?���c���)�����+���s��XD8� ZT6��Z5���8Rx��V*UoNCX}`!��]n&��	�̩��|gV��xyt}+<J�Fa�N�������U�
�}�n��ZR+��1��o�|�����,+Y� ���6�>F�_
mP�&�r�������]8�@���6U1!������XDVݯT]<aq���V)�h������m�Z2�jh����k.�����qG�s؝����#�M ��Kk[���hG�}�o��&�����<p���������g��=`�e�'�_���걳�I+��9 ���ƌh��-N`�l��k����]C`a�C�{�}S�DD�|�(?�f6i�CA9��E�P[룈{y4gm~�m���l����-t�hNWZ@#=�1����{�#(��G�Ŝ	�z\e���gFHt|�י��0���,���K�`S�%�tk�>ܬۚ�@cH�� ���=i�Hq�8�����l"��= ɩ��q�mu�UG�������p��:�����	�@p��1�ޭ���K�8Z���Zd�8����v���]l�������9ٚ�#5t'Ӂa����*6�(J��2��Xvw�t�F 0�4�P�I�����(rg>����`"=�6��� ��Iqcwm(i��"ao� XFl]�H���RC�#2s�@��z��X ��X�,@�.��,��9ha�a��F���)��j\�$aAw0$�*@=i����T�MJ:��MV���h˒�Z���e��APH��7Y���D�("�ю=jr�T�D��B�=sQ�c"���?�EÌi�	�$�xjVc�;H�9.��!��G_��p��ÁhrAx'�}Dy�����f��]2�s�L��i7J�@r�x��d�$%Ȉ3㙢Df`YA��f�����M�,��J,F�׏����}I��z0u|����6Z6J,K}Ş<�P�kL�Z��4+�݃��bؠ
٥��<xkb�|��VK�����F%%@����i}�k�Q�]��rGƝ����F*C��ɋ���Ԛ(�Q���-�{/!LK�L���jG�f[
�}�l�P�+I���8094bDE��V�����ŀBd5���WbT"Ij��Ŷ�I�`������	���4�z�*��l\D)d� �W|�|@銜�a��$�R8v�k�z�}ү3��i�i]��P�Q��.��4j���̅#�FH?x��{i�w$�2ċ���*z�m}�f	�����C���e]0�ӈ�>{��� ���@���^R��xܣ����U���ؔ�U9�棖��Eԍ���.W5�Y�\��#��C��̴�jS�$ \����gC>�4̙ۻc�³��>�Pu��ܪ�܀и��^��M�5,�|7����I�&[�����YT������l�hr�E������@�YŎF��(��_QWעC����&���(q�Z�Z�!^qW
M��A�N�4��S���I���[G}E��I}]t�"\P9����~oy{��Tv��x�G�٬G�c	���%��P�:*��Ӹ����& �W{s��T�88��v$��H�nhf5�\��-��
�X�uФ|���<Y��	���j��晠�4ذ��2U�b���S�z�idYa|'\ͩ5�����|��Y\dO�;�[;�� �D���k٫k�T��GB����Ci76(R�SLz+��\d��<B���{�3��t[o��W+�H�ֶ��x�ߑk�8nz*�!e0}EחN�z���&0���a> (�Z�y�)� 6C`����_?u8��l�o�}Ɨ�Ebo�|��e�ar���R:��xg_�v�፻q.�l��Q2H:��'Fv6�F��+�L<%��Ip��1��2��R�	#�FI߀��d��p���G�dӢ��k�[|�L}du�AcW��O��sM�P�U<�"�������:A�753�aa�g����(׆��	9�P����й��YܯY榥2�1���,8�7(���I>�e�ãS_[�5<���y���P���#�zA������MȨ��5���{$��r����6d�'����ޘ�,;�*pt���n4M�w�� ����*@Y�X��W1�fC�`J�dH��c{�q�Q�pJl���͈(���z'oCٟ���θ�h=�D���ʺ&'=�I(d+�����]x�R1��MI��Ԉq��=K{�{����s�t��J�G鼔��ُ���d����p�nama8>���-��0-��uNi�K\�~>��|!e��_�jv����m�,L���)1=U
H�m)Ѯ
�m/�� �d*w��=��oh���6���	��V�V���	QtonO� >p��Q�zg%����ֹj��8��|I]��2[�Y��i��u�#2H*=���� �lV6A�m���jE1�E���>^�[��ӽ�͜�����Jߞm�8��AXz6Tr��N8����!�֯��B����k�/�a�Y������kZ��
Y��3�Np�'���8�ߝ�u�]�1k�Swj��h�������豤:�^��O/(��O{�����*���S��p����$�����n�
B���]�t��[#�'{��_2a�/�����#�Ӂ_T��:�n��W�#�]���\��������[�tb�)���?��S���]_J���Eg�DH:2V��:}���ul��>����r]S�69D���Ml�O�M��,����)��vP̀;8�e��[�G#>��t��R�0�|(�XsN>�&|q���j�F�k�(+�UV�3{�Q6�5�h� M�����]��H�1I)�s�p�zdԣh�8�w�H����#�����բ��I�S�V? ��i}��|�k�!�F���"=?���*�iq�v��L�aVS<��Ǧ�ׇѰ��Hn }������bxP�i	��l��ot�A��x��[��1�������*b���_�c���bqg�֋�5����/�Egɥ��gP�N�;�P��CX��"^)uɶ����.����'[z{���æ�"q�)�W��t�i���
�����Ix�Os�'�aZ0��ʸ�I�AC�(��9��
:�VW� ��*�P#�+���n��Ư���>���%S�͚r����i�dC6�@)�g��d�	RH��
������X�Z���VS]}�C#JV^�\����O�i�ۛ}��p6���/gN3��#�D)�@R���+���n�d��[��_x�So��̊_�z�fv�(Z"�,8#)��[u�ۑ�H]&
8M(dg��5$b�V�=���e����䤆J��x���]O�s���S�!Bn���+Lx� V2[PA�U�9X��ȴ5R�@��I7t�M4�P>�5 w�/��Mȋ	��@i��|������ԭ�"�H��DA����T�����xG���{g�do��0
3N�>}5�k��[�5�P���g�6�P���� ��ˇWC�)?gc�SOu�'[|@�n+�c�&��8s�*����h�|�Y��j��0S7�1�+�&Q�ȥ~N�a�P,��Z���e{U\�5v�Za�]>�s\vs(>H%�jޏ�2��+����f9|[Y��I��-Mm`&[=Wn��-�*��`��<C�AE+NA�]�F-��)˵b-�#�0�?3���
�w֛�S�Y�ɥ�ڮ��%R�2�p��k����Ay��S,j)�Px��߳�$�D�$�s�t���92���k���o��\���Ͻ
U��L�`��
���.���<�P�X�q�	��0!	Rɚ�Lם��:F�X��oЃ����@+��Ir��\6
��"�?�<�����]=�0���]�C	śو�j�C��<���[�����7�vt�(�L�5������S�����N�3싥bd��+ ���̂�1s�إ��7?)��pԨ����:	wt8��?�D�=)2��J�W����ZT�;�9x���"�xk�LG/��'�n�������x��_�W���v5�]-�C!m"~R�x�x�T�{��9�L�t��j���7}">ӽt<�r�ʅ繫�?��diB��j�������/Q��c=M��mn����&�Z��a�v������E�N��[�6��3��J���К����2�v�z,���G9Z]�1��I���F�q�u�]�ԇ�(T�|��y��m�^b�؄��X���m�ո��I���	}�^��֓��{sL�Rc;�f�+]`��'��"a�'U��?���|"��w�A� ��O{aZ�bg���.kS� ��v`,����Ə�&�&��g!ڹ]XB�T��Z�"J���9��E���k�̓S�וK����u�����]T����Oo���1���4�M����_�ѯ���z�����b8+'�{k�'srF!)�m��8�cn��4���ʗ^_�Km�YN�>�v!�	X�T��e\��wbN�J�d�-{LK#/o~ă��E��cX�sXd"
�� D�e��؂����`&��4�ɧ��������*�M� ���a��  ��y��*�����n��t�-3K�n���N|����G��ī
W�A�U�F披M�P��v��Ir3�qy~'���X�ԢXn�� �R@�W���']���n��B4IG�l��ٻ�P�l��3|L��s�Gc�r?��V�3)�L����#�ݪ�{/_�@��V�"4R+1-w%]�<٠�͋e���x�6O���|��r�x�������V�m�
�2�4"��$���~e[��I[Ly���-�g�R���mu (�z�jF������49���0/�N���{0�k����7=zC�@�g�7Ѱ�䱊z%p(�19xf=Y�������CX���$� ����cZ�i��Uo�y��Xt3N�-��^��~���)�/�|&����rϠ�Y���x�>0_�5N��O�u��K	���t�T�$����!�j����Q>W�%�~���Rp�
~�B�5������<5�����k�\Y$i%��
F�骍�a�~}�TĶ�(��f�:�go����\�������T�9�ZF����S�W�I�\+jj4����[D�������̪�y�7ӭ��I�I˨�I6z-S��dK�nٖ@���܃΀W�6$0h�:������B������6�K�.����!���N:�A�Y�,OoEv����ܣ�>cw�$$J�,�?���l� �p�b�&!������^K���u� Sy|+c1��ڌO�Cʘ�����E"ݧ�O�:'�Nt���/龹b�>edm��g6J7�<ŃS�����?�|�F8�����'?귰M*wג�6K��r�m�Ceu~��|�u�P\���d0��s��(n�}>h�@"s�M7�~}:~�E���w�@�#Mmt%nCk�]$Jt��Ԥ�w���/o����+�蟔f#�����bi&�Eȱ��RS@1�s�|ȩ���u���p0����\H�uqM݅u��0(
�C|6��Y�ˤ�V����G��1#�YƝ�۵p=;���d���Ŷ�u��%�h�΂~nWǔ���+��ۙ��3�忼]lo\>�S�'r�0�ѱ�z;��z��펴�z��d�Q��̫�gT�:|̦4�|�جҧ7+�Ppf2�n��{[iy� ۩���(�/�a��t�1z��P,��:+����"��χ|OC6c�ǯ�$�B�es9�)��j����}���/�]]�0�m'F�2��3��,n��\ �:̏b��jӜ�5���3d�_��ݟ8?fRo�d6!��8����a��A| �};��ג3�ü~72��jE�n������۱��}6<�̥�Y;�ɝ0j��������X��6?�F��^W�p�((�s�6���#��Tp4�U����*_B��h��B���iU@|M���r|^��S��O�Uv�]�<]U��*���\�0��l�.�q��)n��C�>��P��7�����brh�	����4a�H�{y*����]�72a�e�ߪ��GH�����ryM�����m�M���H�G~�$G7đ���ע�����b�k�UG�f69}�ܼ#R>��
�Z`�~�C��yYC�s��[��kX{6�V�3S��N�G����G�������1�S��IJq�"�>uњAbB���>B���O�h{�N;��y��ؼ�BK��7�9JC��"D!k����j��Ia���b��g������w�M;�t�e+�G7z�Wk�K�"�G�w3�o�_��7|����tNJt��4��|P	��E�Q�S�p
۔�ҽ���l��,���g`�z���.���O��_����#G
,�G��W�g�s�;��V�Y�?H�� %]SŻ����F�����"p�bu��Vi~dE��ǚ(Q�f�%F9�Ŝ/y��%�V��B�X8��M+��/q.**ީ.˄k�開���.�7��4��Մ�(���
��Y`�9�7��s��l��co��z���?�ݘ�.A�7�'�����Jcҽh�(Y.�)�⯵"�2��Qf��I����G�\ImoR�G�V����*'0��83��R'���S�^c�J�n����!�^1I;����o���i����In�������ϟ=<^���Sa4��P�&��Ő*�R�u�����N1�L�@�?.
w��.�Zab��V.�]��(ݳ����c*�9���@�l�!����u�6��c{��(�[�����h9y���Oӹ @*�r�ɜVC��vWO��'�/p��� � |�ZaHM+�Bh~�Q��P<�Hp�x�<�
I�b���H�ˎd��@��_t4��	l!�6��o8p-�%G��kD-��4��+����4*��7�lg������p���As[�w{���O�8|��r�o&�����Rd��%�x��O:�ά��]2v�9�����0��B��l�6����P��=����<Q 7Mg�֘������
��GЧ��(���ъ��3�*`��z9��k>�0�6���h?��`�Nҿ%��EN��
���/����l9��ԣὓ�}��H�3�
�V�Vw�A��4@A������맂L�{j�g��e�l�F���+�g�|�q7�Ꮠ�BT3#�H�ǅ[0�a��>7�6I�I��
��-l(YV��R2� ��a��"��H�裉l��ԍ�3۔s�+㶲C;ᔣ��x�7���c�>|ڠ�Zog���3��c�
s�b%�_N�/X�-���,�-Յwn�;�����01����K�\����?Ŗ��~��}Y���]����F�%C/�E����fѸ�a�ϣ��:��_L��}%E�Y��0X��j$��	a��ۈ&�Q0(�W���|�@�y���m�	PJ������,G��O�\������X,��B�g}�$�|=f���U��t�ggv	�v�Y�)��b~�T)��U�I9�$,?� �� D@���S�X�����e��w"�FT�HZG�En5x��Z�ù+,��c�|p"p�Qp�)ը����/�V���?_3�?�}X�Gg���,�b2�܋7)��2Ǘ�f1�.��_m�����%p�'���4��K��x�d��p��}r>�M�m;賍pU���@�l��ԏ|�2��ۉ�b}.��akʳ�hX\)=����<���6��ʆ�R�X�1��4m�c�V �\h� lW���Kq�y�kK��2n�����p�[�d�cu[(l9C7�����1�-�T�,A� �m���M�q��}i����CX+�	�;EFE�Ip��!_��A"����ꤲH�ja^��Y����J��$�܌�u�&��K���M�y_�l_6ZW�� f7�0�f�g��g�� z�>h%>h*}�eNw:K��$t�E�:ÿ���l51��H��fHv0�V�����D�^*��;
�(E�1�?�պ�f>2О��+�IbS����e����&���C��W�A"���I�ƥ����Ċ���e%��@�w!۝� �h)����Z<錛�/�O�mʞ��[9�M_"|0�`|����%�g�|�����3��]g����d��Ч eu�]�e�S"q�ͤ��s�����nc+�J�y ��X���7)aߡ�:���-