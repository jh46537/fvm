��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8��A��t��
�]W˱�ӆo �I{�C3槏��ff7 8��6���7�Y)`6�-�7,!�=�f�&Q��"�qiK���ﳑ�ɃnT:��J����""ӜJT��Ʌj����uo��]B1��IJ�P+p���Ү�r���~$̬�͇��!��||�XG�@,U���56=�t�we[�Ax��mԧ3C�d�u!�R�9У�X�c�m<>$y��l]�
�tf�?�� ^��fdT<�n���r��s�?��Z*�����)��Y����:�v���c��0�`X���}m�z0\)	�/O��Q�J�rV�SK���&�v�!n!	�!��z|�M�%.�.�\��R���Y�q��CN�`"$�T���9�w{��˙�������m�![�Xxug�i/�~����ʠ���t�s<<��3�54s<���\0ΗT����a��	�ֿp'����su��p+��hN�#l'�I/O��fiUJ��,�����m��l�0�=A��ݐ3���25>pE��S��������nDa�"9	~4���h�K�aS��'�B:\�`���ӝ���C��a8a�,���*��;�26t[ۼOCT�PX"��%{�k۴7*��Mrb����:ghl��Aғ;'�;�"�^$��z;ާ�,OU�bK�H,�߉2.a�N�cls�	y��`�t�g�N]	�� K��Eo���%w#�A�w9�0 �';V��:�[]�ׇ�G*�/�3�~��&_�m��>����
h�Ώ}BDa���x���/㪷\B\ 쨚.�U9����"��mn�Ĥ�������8'���Jm�j�l� ܏�f7*�gH5/�	S��4�b�/��g8���������LG#iq
d>��V�o����}�#�X7�`BE��̝8��j�T�r�қcA�\5	�JG������G��;��ym�1=�P�������GO�0����fs5 �3Λ�~�N�K���`�Y�g����Ć�/��`nH�2/�U����I�Q�pC4?��Wu>��26�ps�+ŭ�P�P�js`����y�����ߊ6-����iL_뎤0V}	Ѻdy���j��7�y�]*��A�ǒB��V�d�5�ݟur�:�!/h.��M:���oK:��E�P-z��B�t��,y�%|D
�4��wX�����9^�VX-�FwK�(���e�m��7 ��2�̿*���/0iSP�՞_�Fa����L�	U0T���7KT��\��������ϑy�.�~q/;��p�6��K��K��KcTܻ�Q^ڻH����s�X�=s[�Sq��1-hQ����m%Y���%��Fd+�յR�Tmx�����N�r�M>���*1�*w&�T�~W�@맰&�i�L"kJUV�C��%]�_f DP���'A(�ڢ������[髺��������Hu{�DQQ�*g��$+X�^n߱�%S0u�����@���r6��Ə\b�ȁZHt��o
o�"�bl�/Y:�v�p�^N*.�?�����F��R֍!?��vH��~ǉG�	Ă[��3���c��l�q���6�%�wb̟�bI�/�EB�3Ms;�\��9Q-��՜���W���}�RCSΕ|����u�B�w��y��(Q���i6�/<�'�I�(�T͝"���G���h ����^� &}�kc30Xu�G�/)*��L ��n����/hr�SY���}*�	�;��ޡԆ���YÅ1���&9�+Q�p7�P�Gf*S0c�-¡nn0��H �a��k
�@�4� '� :G�b/
I�U�?!D��&��ȅŉ_���,�
���H^�=�Κ)
����\�Ƨ_�ģZ�88�v���n�s��]A|`o�&!U�l����ˑ��Sazx#V���ހI��؃R��"**���b��T�o��*G��K�qN��QMܗv��=*�C*_s���
�uw�5���z O�WR� '� ׽k���Z{�s�d��/���ғ�����y_�ܸ�-J�1ɦ�H�N���X��ѵ{���:�|/�@,XGV��l�8�%��Lnәۨ]J~�$Z(v�Ӧ��P&����hƌ����U����1��O+y��M�BO55�5z]C0��s�'�>vRNp*h6�2K��z(��$D�3!���>ݍ�m��x��ߐ���8�+��!0&�FP����eS]u�Q���{�te�O	�-����%k���j���Y�#�����۶h��0O�%�r;��/�vP��?a�{nY1S!#��lJ�V��c�\���!�SXvuJqэ+8DC�3�L:�fRt�����]n�=>�
�&^�����"����� ƠH��.)��U��	�Ibټ�t�e�A�*N���! ��˷M�Wmź�?�	���8��_�i�r9�5r�8M��sLJ��f	�G�E�K!�U��OV��Z�z���T��N�:'�;���s������ZF�xB
�,�6O}W�VLA��I���'�����yYg�}�9{�K��s�w�`�萫�?8��U�����}���w�qנ�^,wɱ)�v�7��`��������&�8�1���p�z|��M� Xs����8� �Qo�;qǝ`뒣���OUd��#d+uMͿX���H��1����}�h,~��Goa����Y�.�6����IM�:��]	!�An�iA�?i�ǑQ-�هvد�E��=�r�=A4���7Ӷ�2lš�.������$mE}m���h%�U;i�K3��I	3�,9�>�R8k�.T����a��P����K�b��r��4�t�MI5��cl�n�Z��9'De�%Z0^�E�/��;
��aO�PUj�*��~��ȩ%���	Z�_Q�l(��~�yP���~���V3'�K̮p�J���3�y��d���<h�y���~*�*�u�B��8-���T����s��U���� �o�Ӹ>v���\S�٪t�3	�2�DC�	��e����;�Tľ����*B#�U���;����?����bׄ�C�d�=Z.x���r1�n�g� �\��6�����soߴ��?��T�u��D&_8�InuS�:��h�,���pS7����Ag�9"���"w��iʊ}����-�lh�|+9��)�a:�_��[^��"���(���H_�>:Vڀ�I�$p�a�v0�Z�� ��{p+ܘ~4���/����^�����	p��r(Y���H�Ũ<�*%3M1ܾ�\�i^K�c��t\����� A��� ��[ �����JR��lW��A������X����\Um�y����s�Sr���U����e��"*
&s��e�=x��s��[�&$�ʪoC�s��-����t�;�z�=�J{"���zmq]yr�Ř�&���0�R(�$A�
��(Ыϴ�h��X��uء�*`���0�$&
z�r��ak�=·����0�۰q���x��?!֜��M0!i��7?��|���"��z��@;�;Wy�Ή������(���}eP/����7�g0-��;TK�����F
��.2}��\$�VсZ[�-g0T�P��%��/��}/�Ni��^�$�7ȥ��'��m�Y��,`F��D(7#.竘H�9
�"�{rEt��i_6�(5��'������'�"i����j	0�C�������V���t�'۸�ѨH��`\�$��*�����qj�J@�$�	M;E��l�s�2Avp`����3�j ������ "���q�3����Xd�/����|.�%C�@��!�0��XC���5O6NҤ/�#�}����ox��0$s�!�2�o�>XW�"��O�FؗRHkh؛	æ���<A��aW9�0P�*��;���a�0��\I�z}vf�s��`��/(�}��fNά���HS��_}Jy<�\��-0���*�xK�O�����wN⪎�A\EEg��7]]K�	G��Kña��4U��K9]���vDp){f��OE�)4�F�>�cs�k��3�HBC��5D�ڮ���ȵ}�KYՀƣ�PؼV2H���w����?Wg�a&�Hd�;��+p������̓�x�!fH`۱.�R��.Į~��8$��D0��jt�^�P�	I���.�v���iPJK�ge"=C��s�híg�;jܠ?
9K�CY�D:W�e��XC��N*)��,t:	���FR�P�xU�ZR<����xxg<��{��NT�9���q�G��K�9S
sCɿ�\�S��H��]D��W����;<��s��f�/9��i���$�:ـE���_�t�D:�,��8'��d}�mӪ�I�#��W8璇�^���;;f����s��V��L�i�\��J<+V�f#�e�0��؜�W�kN%y�*�Z7�Bc���?.�r	T^���J1�����ι�����)�IZ��.-�d@���6���D���W�v�g� �r���K�����ھ��&��r�0G�v@&�Ҟ;'U��]���M�4w	�a��`N�X)A�L ��cBC�A�KE��#H�f�t��Bwr����lX����W�Ӻ��ug��W䫈��}Y����/"8�!G���I����d%P�@s��4C�?�\B`����w��)��yL�1Nu��� -q��,��	��N����=[�K`��,���4���l��;�K�(��W�VPd���1�!q��1�+zW�Jؐ��w���ܪƐ�������څ]�<*Fۆ�*�Nm&�i�&F0#݈~�5����gen�w���[1)�K.�{�|Ju�w�a����bv�d�a^F��Ỷ�2� �ob$��v�[��ӇU�%��Ll��Ն��P����X��6�J(�E�L-�Ј8!HW��y^��C�_��M��VM�Eq�η�j}�)H~�u���i��u�.z6�p��(����%O󠜑��HE4J^j�.����V�#��b�q\I��k�A`!��ܪ��_U�~-_ee(������NvZ‣����9E�h�"��T��1����a��֩ݨ
4y���o#{����8��Am�a,���m�0"	�;��g�F�r_:�_PH��x��C�V��Ƀ�«��]ʣX�C���G�2��4�cFsjWɳA�ZM(C��B��'�h��#���� �f����d/���|�����e��E�R�x8�G�,Q8��GY\�nN�� ���
�r8� �`��\�nA�\.�������@�E��Y%���!��|����FE d\��8�lm���	�ҜF_�����hW�B
mWp]G�0k���	x>�،xTs��B~�q��sxv}rzF�����i=�k^���F핹\�k�b��W�p��^-d2�'<F�0����=~:������b�M� G/YtЧ	�N�so_�"�כڶJ��,�w�Z�L����H6�w�a��N�֕�#̏�,X'���1��V�H��S��b>����h�+�:���7+w?	~�E��/����K � ��i"J��R�坆��ta(R��+����~�8�ͬ� ׁ��<���n,?I, `\im:x��� A��(������_���C~�tf&đǐ(La���y/��6���I���l��{����۫/m�H��Q�b�d��AY7�G�/�4���K�ݚ�1��Ce�`{&���4_�jxOq�2��Ϗ��8@�w7�@؄!O�D
?;�}�5�K:5�ɓ��j����3���d���y��8y>sG�S�ɼ�BzH/�q�;��L&
Z��1��L�B ���%��(�à��{�������8f�%�B��o��i�U��@}J�:��$��hc�
�dC�g*R��;��=ĄZ�E��C��\�D���k�	?^������]��K��9O,&� ���.ʁ^�Q��^��f�I/����-�
���i���N@�ֲ
�\� kw�D�׏1�%��P�N��b��.��P>���#K�G���\g�z����.e�pw���]e',!�e3���__r��0�Ab�	ۊ�p �N�d�O�c�X��˱&��oW����gJ�A�s�r|�B�h.\Y�e��
k�d�����K煩gDb�	-5�s[�?�bk�9:�I'�\�������Hp̛jM���4�̽�풂@�1\���G�Ԡ6�Xy�I�K� �*O������ߥo�Tu��(��U�u�/p\��K���o[��p�=�"�R�����������I����ݽ�
jZ7�	|	����Db�9�J?�R0�DFKUy�����lf��%T{��y�N���V�H���/O�AĹ�b<��,7��]�Z	�PU��O���d��ҷ3͙1���H�&>����V��LU�����鰼K�gI�rh���y �T�x��ɥ�S��{��u���+�,Y��O���2(Y�>c�S҉�=Ǿ&��#
���:b��:�2�3;U����;�A�����4��O�я�H�;��cE��6zN�m��=���o��ud�ٴd{��z���#�}tk �>҇�n�'�`�R5��bD�؞IIP�5u�ȓ�Y��aSEI���4���c�&��兕5���P��wY˦">���*��Z�bOWn4�;��ȹۂ_��a����6�#:)=䞟P0���/�&��ͫTa�ѐ�<���igf�:@�����E-��\�];���$���u�qI~��9��������m2���V!C��J�<�D�����dk��s�O8p���KC��Y�мm3@7�v�n|ެ�[B>W���g*F��2qU*¹���2����G��/�T�%/x�a���@�NL����9�S��>�Z�$F(�qM���-&[a��`.?\5oL.��;a;v��c�*݈X����s�9I?��`s��"��J녧r���)���h��E#[�l����|׋�h`L�m���<�~�F��X篧�d���n g�!;�̻�3~&Jp��9��`�>�:?� p}��,�f�G�FP�Ev2PL�[��1�C�z�O`:(��(����͖��S~T:��bkA�x��ZƏ��7�[�;� �Ho�����Ȱ/L�u���H�y��v@]��[zw|�2�cy���Ѫ\A@-)�A�_��f���r�1|���~��3o��.��b(��t�R�[�(�����:hI���Sk=�W�o��cɎᓚT��-������P�M-2�����$�\���͆���\u���<a\K ��Ҿ����I����_����8�~ZOGi���1310�QL���&c"4�����^��	���#?�\؜��^bR4e��n��9j�"O�$�^q)�Τ�|}0U*"�Lq���t1��a[Ş�!`b���L��yysJj�a����)���a}����AB쩇Ne�xW|s�3
:���� ��6,���Y�71ګKD�[%��	e*�z���4����Y����Mg�=�Q�fR�'��l�t#r<�k�a�f<Iҳв��+u��[�j�1R0�O00>���b<Z��zz{��r�C�=b��n�<�o��4�/�U��VP:.�ޙ�e>��"�Î��������� �/`Ij�;�n�s���b�c|����K�r�PW����`ٹ�ގ�D�z�P����n|k��_ �/�������WRn/�Ii!�yB��8���}[�Y�!m,J���ͤErp1!�]��;�19۷ю��\r����;�O�1x�CV�o0�qn�x�Go�"D��	��(W,���*��;������y �8��L������R�  /X��J�>���u�����U΄���N����{�podA�Лb6�#-�<^��Y,��ŰMX*__	E��@[Bi3G�.8�l����cg�@� �y��'BIPX���%')����f��������\Jttm��+#%$��b y~��#�с�U�U�ԋ�����:r �B�3�Ť17���P�Ͳ�(�؅hMog�,����Y��+~ ��ڈ(Y_�]�@���ZU���+.����bUE�n1ܸ�J�,���O�6(�<���v*9&��MV�I!�T�3���s��j�!d�Tlw>�|$;s�� ����?��Jb�9�U3��f� ��(�!	Ϫ��5��y46������kĩo��"�����W�q�r��Q\�7�/m湺�n�hrh���*�u�h�b�W�Q�/M5�eI�j��w��\��ؑdF-Y�!�b�:�!ӁA�1$lG����恙*�n$D6(����Y\jW��.�v	�����>�`0��M�SH�$��-��Fa)�	_�63L�DI�gǾÍ�PD��д�Mo�D�ltZ�"�B@T�����ێ��5��q����0�������\���6ڃ&��΋��Vɹ�{��}���bw�3_�P�vt�5�>�-�p�]�x�j�OM'�_�^�h0:���p4S�5&��o˜ի-ph�����yI`�l�a�c(�1	N2��V\K�h���ݢ���U%.��\�Fȉ�q�ͷ�:b���/B����=��x�ZC/���oʰn�?�J��&�p��UI"��#_�^EPp{��f�Q��C?4\$�Nr>"�� B3��ň���� b�'�� �� ����7�h��f�~���7��A��fn7�»�:��[��#��<����� �t�i��Tsgclm?�Ѽ�ht����4����d�Eoz�r����5{ʂ�%�wlz���ɒɚy���$�li9A��݈ssZ��=����Nׄ*N���a+H!2�#ET���g��D�L��&�ż'b5m�����`��Q^��#C[��A��5��$�3��`�ĵߘ��N<-�3�o��"U�"��.�B��D��΅�j�W�V�Ydw�Ӧ�b����V
� ��,��k�B����kR�ϹT�E;Mʿ��Ge�t�c�A��������&N��w�+7�a�w��ģ��C����rN�7_vk�/-�؎v�����ۘ��e����n�r���$2������*en���/ ��gy�g�fAi+��sm5����:M	!&(��|��?3�L���d �m�=-A�~i�\%Si�NU�,@��!�g��ڝ�mVS�}�=�B�����܇ʻ��>{������}ک�z��I$�]0���S>gj�m,�@X��ߡ�L<����k|�I0�L�@��rk��j8M"l1�_�&�%S��J�1^���,e���5��|m S�/D�c,L�#v�x=��I��r�Y��Y�2�Ġ�~o@��Y�ٞQ�[QĒ�+���X�^��!��z�탇�8t��D��+
$R�����1{�������z�A�g�
D�]ݦU�/ �#.�!�Nq̉E��g�PB*4�^���O퉧 '��tgs�����S����bTw�s7d�v�I�4w�;��cf���������WѦ"f�j�p0h1�Gu��-�mk�1�Q�F�զ%#�6�;G&~�D�u�zO�Ь��ܲ������@���	���[1�	2�ׄ���)l�.�cHcSC�R�޺�[��x��Y(�t���K�m�8�����{�`Qүb��u+A��5�ZHpx�R����]��IC�b�fz:��6hxC�G��y
�{�Ĝs�x��j���m�oۘ翾�Aئ��8�&�T�8����ǆ{�L��^�p���~�a�7w�!�V�d}ҝ�:����}�Z-e�=w��&��mA��89봺5W�I��-,��ۚ��
�nWu~$mi�-�Q6m�%ˮW�j������10��SsX��w:!�!a`�e4{oV�>��w�=ŋ�y�X>+#*��EVi�̉��%��Q#yl�����c�1�(m���]&f�z����F�VS&c-�۝�e��D�F�S@#�>ݛ��~v�Ja�Q�I{V�^n�o��.��~E�I� EFA�:�Yӧ��3,��{��R�����W����c�����N��4��J4��,:���.D���l�)��������D�������uk���2CQ�Fϖ�����Ы��(��1�����ґ	3��'d�^v<�'I���dH:��0˹:�%�2R��#j_V�|hT��.UYc����F�Y����H"��Baw멈�����A�c6Pt-b�$��b7��J�~V�`qz���j��{&�2�އ���" $����P
!cw�{4��:g�/c�=1��@������JۅƮO%#5�p,�5�t��&%���P�l3�;�塀��zJ��pϡo:��d�¾t>�r�ǡ���i��^&!BM�<ӱ	T�1�"8`|���b��Ge�[$�MQ��0C��G��W.�+~�
�BG��$j�d����(�҂�,�1�kJ�s��j�����2鴲\T�=�_�.����hϞUn�a�}qXf��Ñ�v&b��b[����q����D(C���P�=���C��	�s;����D����	�F/�D��u�#ް�`�%$.��2,�-��ْ�6�W�IN-�Jtvh>O��Y$���(����+�*i�c_I�����Ѫ��{�q��zjG!C��^�W�c�w� �rTJ\/m\�إ~֜�C�
�h�"�J���&`��� �q��d�9B���<���+��\$�-KYK�u�~�d��w�:5�u�	�@T���?6l5���@J~15�#��*ϐ�����7S�j���iQ�_D�����e���/�@x`�C��b�=LR=/z�>�E*m_s��Vrb�6��DNl�wipUT��r��UԘ]i�7A�h��m�6f�b�\B�7�HC����/(��P8�M���(IŚ�U�ٽq-F�y����/ϯ���GAc�̍�a�!m��w6Q-RU{�B�D
��6��?���x��j��~��QRC��[��ד*a
d)p��������,6�?!s@�dj@q��S��12$B��*����E$�5���!~ �����7+ѧ�),��8u������-���Y�>2�ޡ�azW0{[�]�C9��%V�'��#��32������7�#'B��o�a;��9Ƈ�~��g���E�6�2C���s5B��y�R���)v5�m��<b�kTB1`�B�t�0�٦��X��YJ�^u�Z�n�I>���(	�hC�A�©O�a/�w{��膆�8j�a�
��ʄA��<{�n4������a�8�W�T�S���k���o��>SӀ�0�w!-�ڼ����b���ՃR�4@����k�蟄F[L�ݺs��eV�ߒ�M�	e�'l%�l�_h��E���Q-���
Y��HiB��.��!�R�A+�ʉ��l�+���y$�Q҇g�Wؓ� �"d	�*�Vb]l6���6��������.�rY���������w�p�������kL��o���)�?%�7b����u���/�r<E:R�al.ɕ��$%�@�rdY�3V�)�Zj�s�k5j۷;�"$�pg��fG;4�~`ᑡ���-ܜ��h��ּs/<gr�i&05-�9��R{̅�wn{�_;�%޽���d~��s��x���$q^1�'M�틹6���A�;|��ŋb��s5����Bu�\+��@�l����K.���STur@�i��z�@���h����-�T��Z�U���&��$L�,�Sqꘟ����Y@���tŔ�PcB�R��\o��Af�/��%.����|�Pc.s����E=��T��1��s|��~�O*h�|t���I�dg܃6��J�����݀p�^�12�;�yT�����m�,�%yE����Z�W�������x�!V��(I �e�����r�X&�y��.ɦ�����A#������_�Ʉ���q@N�ZEY�
����|S~A��=�͵\��m�N7o���.D��R���k�t�UEJ��!�Z�l�D�Χb&C�sh�2�vM�//��h|V�DW�F�����N/c@�+�Ŭ�N��Nf�Jܹ�ڤ ���>��ݼK�����2��S6,��.K���1��9x��O��[v���ib6����P�[X�_>+�r��7�2��m	��T-�H�,E�6	'�j����W�6I���g=�C߄g�O1�G��M�����%@X����=����@���z�!��fj�(�8��{+�J*uSu\8gq31���?�{�׶�J��&���l	E,j��m��w��\�����!ө8��(މI�$���yB�n%2a��XG�Re��}�j�+ba�g�͒��"���i6~�j�w���ijtB�{��4}y��Q��TqdYWv�7��R�v��	���s5�H��~�ﵻ������T4�Q,S��ܭq� �ՠ�ƪ���U�RVxAz�Ә�C��ȗ�F\_�Uk�آ��~}��^�Y� �������i�XwQA'5`АӖn;~�?9�%�:J���S2n���������+��M�n�
�����<~���d�{_�G<d�b\Z��8������,�7��s�����x�4W��nl{|]8	��̕K�ia�A�,k�$&J6a|���C�x�?��2��׶��h/���jtGX�`f���I�:؋_AZ�����{���w�ǇgM�:�Xy�>�%c��צ�����ם�gAIsy��i~������97�(az[���İ	�C҂�oO=�����
ஊ.�m��N`ou��=?=�~k�	}7�9�ٺ��Q\�c'��q-O)�>���t~�t�f͊-c��뺔6��Q�d;���ZP5�~l��+�5A�M��_��8!���kK6�L4r%�9K���l��.�,	�3l�@��o���n<�!@柂�b��g�C�^i>o�Mݮ���B@���qH%0�F�+��HYB��?�R���u'H��"[:�i���@��YU�s�H����g9g��k��'���qQ��p�"�%	7��.͉@��v����؀(�ɳ�x	�Ӯ�� a4�GTTL��ْ�=����Y�踺~⋜�=Þ���̺��I��م�1�-"s��T��� ��E�,�¥g��q����,�˕�l�ވ�Kb��V]@���o�/��uW�hp���R��Ǫ��F���6�-�ݑ=���'mB,Ҥ�ߝ�fI%Y௑��|Ƃ��ዼ�E㮔���{���A�W�6Y�����)ԟD���5H�]�����T��Kߨc��AL���$}�t�Ħ{����R+89����o
�s�Ť�&�&�5����2���T.�8q����p�q���R;�C��Ջ{�@}q:�V�VJѐ���#1����n������k>��������ǓC?�?h���X�r'F�9Zn1؂g?g� A������qޕg�MM3�ܳ���ԩA	��x_e������:L�ob)��p�#v�����\훨��CvZ(V"
Ll�K}����pLʉ�V)�O߶S@���6q(1U�`�b�#X�E7v�%�Y�q)2�������%��^כ�l��,B*��f�L:����3��ߔ�πd��ps C�¥���`Σ��X�����貝qJG�����N����ň �{b#����)���I��-�hO@�@�{D�$'���$G��t���4��N"�oH1༏�Eo�ٻqaF����3س��9�>�'�'g=���,���N�!�_(��#��g�>S���艈djn���j�Nݧq�n��=.�V��^L����~X[��/��.��z���>ft/xt"�� �h$e	��IҪ�q��%�iQ�*1�K[ծ�X}8i8�����ڟa��*J3U@A��D�@��C��Iqr��eSj�EE��CnQ���֝��mZy�@om�J{�Uԕ��Mc�)�Z�1p�m�>�۶L�Hgx{�^
8�)������=D����		\^���@'+k�{o��o�=��j�3�Cn��
c<=>�D%���X��5>��r"<����ޠXw��E�P���S[�`����Q�О��m��)��͓��;���.$|��ķ�0�~�H��tp#7)��L����O&4�����X��M$\�奨����������q�b'��z�@/-yX�t��<�k���M�����8 ؏5�/伌�7@�A�[M�