��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""��Ϭ��U���rRj'h���������;k�4�p�NJ��)F��B�7γ=������o��?oIv�qʽ����"D�%bkw���	����D�y�����Y\���:2�ϳ0#�Z�xm�:I��!�YG�m���'�/��`q����:װ�e�_��=bE��qE�r4o�} wϽ�y��'����u�z�V���.��͈�f�d`��� 2�#(ׇ���G*��:���L\(�S�����L�p\��#sBT�t�����Ȼ�O���Թ�Ϲ�Ps����nc�K�Q� |�6��Y�/1:5T�qY�&){�?a��)���A��Z���RGF;�e]Je�ޞZ��̴vu4�͛pk�'��;`����i�)j����$��X2Cx���Y�����KD>u�SI^�d�-/�A^���*|�]w3dǞ��"���L��~�Y����!ǖߦՐݚN��̅t�,L����	^��R����uz܎7D��� �B#D;�<]���/�0~�ؕQ�sv�H`�$�F�L���z�R ~V�U%�t!g-���$��%������]��_3t3�[!5g�%��ߞ6����l�e}c�<���Z�����pr<�J�/�yJ(��I�]T�Iy�sn����uG��0�zTlX��S���皎C��y�P{�&z���Sҩ��T!EBQ?&:�4�� g��,Xh���W|Xoy^�Ap`�0�zDz��3����͍DN�cCM�lrh�Q׵ָ�O��1���L�l;ԮEP�&���O8��/	c�{ȸ�l�S����J��4���Ģ6$=��ie̕�gU�Ƚ˃�
jߏ�m9g��pq����ʹ��ِ��T��n�q��8�ȋ/�E?���x��̝Pd<� L4%6.���o6?i�9wS���3�/����������o�/N�����׶s|�T	���$�m��Z�M���#/0���OX�����jki�-P��v�5ҌӲ[���:ڢN�/�F�����.�j�H��fs�v�<KT&�{O��O
�@6`+g��|�Rŉ8�ـ��r���U���.��3��޽��p�K�`)�Ԁ��
="��b��%!�Sۈ���Ł^l���]q���E65��;�vG�D�b�֪ ���A%�R�H%2�oVc9���ʅ%���7P��X)��q��/� �����VVOhyZ�`P*D
��=(t�H��;���Wn	M	��Ҡ��\"Vt��_��r_�y�ɽ�:�nn�	�� ����Y��<c&� ��L4Տ��`N��J�ԃv'[���5��7��Tg׼A+���c{my�ˌ��{{Ȏp�#8-��"w�苍�d^�v�"�����j����U�#oJ�`r�sQ��CS��+u�9�!6�� i�]�iר�'%�0����t�eP^-�E��o���z�T��a㈶��Bf�߳C��X����bɐ�e����x(����DC�~�2aKAZ���A�ԸV˕��8��;��!���G=�v�B�ODM擢��	�ʏ"��������..��#��$�yÝ'Sg�%k�r��X�Z5 ���� ��\A%0/{���ۭ�1�|"3�(b�_L		cX�F��')p��);b�����̓껈l��}�������#;���i����v��&���:~�� [Y��UO��o�~�H���R	�ɾ1���*�YT��m��]�A�'Ø������=�B�H��n!w"њ}�Y��+��!S�4؎K6&�ܳ���s9�Wya�����B�� 󂅁�[��/(9 ;sH�7�l�����)��A��m�V�@�{N�����(�e�V�ی3+�i���Fe��a��?���83=B[{d���2��j��N�0oL��H���i�YP�x+�xJ@����uO�.Cș'�lQ�����(*�g��ZBw�~<�P�����&����
8x��ZcV�� H	��3ɧ�v��n��������C816)KT�5ڻI����]�c���p�[f[���gL��8V�h{�q�ӘE�c��!tG���Ϧ�]'�qC���U-h9S�������c�:�9���J�N ���vX���.H,j2T���@�>�#L��� |��*�,Aɘ�j-�L;�G��%�ƽ���l/A��q��\���y1)Yb��!a���~a�b��׼�k7	�3�
�Û�A�����|/0^z!�x���I^��?�Z�<���ᜮ��1n�����A]u�Fj��Ń:�"��+�|H�bVDEP_g��VI�
9��J�b���2}��K�[�u&���U��r���|�G��	��(�R��'�0?3L7�����X������Q��e7`b�]������o���|��y(]<�@�S�I���%qa�H[�2�^�d/~p��%1x'��,2ں�ŝ[=0O�4�n������g�]��%+O�P +:p5������32�"��ak,�Vtps'��)��U��I��-��"s�4X_��0V⭛CS�����~�����>rtCo����_�1�
"�%_l�k3�tk̗.D��E�]��ь�`��0�/�e����Im0g���]0sp�h2�_ۙ �!*�S5�BL^�.lL-˗	!�r��~;U7���M� ���ygҤ��[:���>�`��,òMޞ��3ٗw$!f�T���$�g3vl����8�E%���1~�K�3d���Jz`����+3,�P�'�@q����0�Lx��Э�������\H�e�*�����;�������0���rzP�{���ٔ��#oloTN?�I��3ϟ��9ܙ�/��e;1j�ĵD����0?�	��>�wQ1�
�g��!V�Ĵ�9����~��F<��ˇ�ͦq.C�k����w6�����	��7���l\�?G&���v���G`��r~�¬����$L<7BC,1[I�.�����)�/P~��j������1�<�"uڽm�Q���P���|��g���O��S������%�W�#ov���k���+v�HK3���u&���ZA8�~���r�����E%Q�t���i�T�Ȃ�_z4)B�{u�����׮��ɖ�^��k�>t�`�(������J��.��Ǟ"ў8!����F+��1Ìr��W�E��C�@�Sf�E�>��!�Sغb>�<��uN_a�xcr�u�̑Y$��Q?����p^=�i(�-~c?��b���二�����]��?;8a����7R�V嵷뜂$z#>r�>�̰C<k�	�u8�D���n[�(��Z�ڏ)�Y�8�e�d���h�=�P�4�7��y8�B�Zc:{e�*�r�(b�s�RWl���ݛ��C�@��c��)���iWŊ~��S��"s�c��n�.����h����N�:,1GM0�n��KL����Yt�0�������M���d����Ǩ�����G���*���y�27I*Ğ��S�������齥�;.]�4lF_��Ps�qp���k5PR�LCAǺ�kPo(��P�hk���/��z���Z\7[`��4�T�����W�c��� ��>DUor�TwΔ�>i�}�\��'7_,,��6�� �~���*ڷ���[��8C�[�ǝ�d_X��85�Υ/�T*k�@q�dq6*A2'yb3�}��E�0��J��GjyL�8$ϝ���@`���n�e�a0QsH�2;����t�A��<G�N2��|��i��]��o����S/�]�ݞ��Z��)�<*Udl\+T���u�{�Wu���Hs��XEB��}؉J]�B(��n �w�h�Od�E�](�Y#*��6㮻�X�'��<R�^���v;�)OF��Ze�ǔ��>E�* ��t��)�F���*�(:����vt�o�Yxrِ+���$cc��"�Iih�z�a��h�'wO�t�xWD���NpQx�u��P�_���z���]��AB�$3:I{gXE���xm��2��HO�7D[�|�\8��&V]��O�Ը�}@����P	����J�����I�	L���8+���~�1܍�w��M�(~3В��2S�ŏN<�K<���_p�UzM�-9�����o���_3U_n!�+3Us�,)���,��y+����s�ڭ�kQ����4)�����*�>�(N�B$�.:nt�{�`CF�N�h���p�@����,L��M�Қ1���[��)���9�+
����so�	��"�"���V���m2�!��8���r���?�q����^ff*�x�9��
L�Ms��;m�[6�g;��;�6��C*@�P����y�q��nG���b�� e�����4Se��-}a�d̍��B ��>!�O҅�,����B�����T��UJm���M�0���ǝ�G~�g� ����Rf�c���9��la� cv=d�6�;!WF�B�|�)�������H�?Ż&�]P�i�7����	h&#�F�x��H��rm�C���ԗ�����{��'Qq��@%,oE��%�G�i��3�vv0A�u�'���� �i��*����|�~g��{՞����s}��+SYu�s9�@f�mc�!سV�_D;�y�b��Ө�����~C�m�(4�k+]!;���˴��s�Z_�%5��A*g A@:�f��������C�t$1�85N���^%"��B��ܵ�n��֡R�ܰ�n�^yq����l�A����w�p�t��%=��V����[Y�4����̤�Ʀ,9=�7V���s���������\0I�
I+���)���'��WU IF�@c��z{!��Q����BT]�G�4X�HU�*-W�\�"o������ǝ����PFL  ����J����N�oй�H[Hr������1d�v�ir�)E���lQƹ�>w�L.#޹*8�,(�	!/����:�L���F�� k�{o2"�O��!�\t&���C̮W�&;��o|��:�ju��3g99F%8�?#dV������cZ&����,L(�.s�ˤw�T�O�)�:c����/}"�4�c���(��)0�u�%V�e7(��l]R��g���4�!��E�E��[�f�RO�a �]������I�;Q���4��#�e�2-8�����:�^��q����B�O�[M�֞W���IY����&-�,�� =��{0� ?]2�"�D
d����Hj�M" ����	X/�m���τ��}����r�^F�k�F���I����J00Q��)OIZ�%��H��q]5��D_3fx��މY�LGo�k�U�E�
�>�g�x���F4d �{����x<6����7�m����D�_�r�ˉ�D���uI�) �iDON{�A]��,��twf�� {W>�%����rPX�I㵑$p1 9�?�OФi�^�a��v�!���W�����E�ϋgRp�x���)`��J�E����[�w��F�I~6�ٿ�>*[�������1��!*[�ɥ��j�9����8���B�ˍź���R���d]v��#�5u�n���YCZ�z�gti�Tn���YOk���c�`��a-i�M��ԟ���-ɮ�NlRmaqC�L+�7�#/->g9��x�����~F6CW���<�op���&x��^�x]����0D�YkmL@�"*$q��b?�
�յ2#�'������p1Jr85Õ��m�3g}Z%���)
*�iv�6d���/���xr�7���J�=��[��B/�P�!�hdҮ�k�6�oA jI�h�DFA�vHf���I�9�|f��^L&��c��bun`وg���x
��/��3-tŋ�����}�OD'�H�F����x4���j��{��a,�?�Ht��B�Ct�es�P�TR����X1+d�T�'��eV�i)��+�����C���q��ųtm-Qd�H�s4��0~d�
����g�\)�#��xc�XST�.j��Nk��Y1و	� �*�?���׆]ӖV�c56�~r4���ۉD}���kv��=��`���);�Z`�%�S���H4����!�t�����1��c�%���E� ͈<0�E��T���y�O���wA���h>�d<xT���7�Q�}��Nt 5d}_L�m�G?a�������].{b���Ģ�|��m���W����vV+�8<�����	}-7Y�����]��DWtb8�$�����4����R��+�����_�D͞N�L�PX;��~��I��@����U\�3��h'}�����Դ4��(&C<_\6'�;y��OSB-/�+Kp!�p]3{`��W�~�'@�3�ui�T/��f�Ar_MV�נ�>�=���A��F�J%�S�nh�E�b��߼O� �*R�PJt�߻)�l���K}�~���5��y�D�qi��0��X6z"��m��Ľ��Z�<W]v6`���8ľ��x�ٸ�گ����e�e�ng��y�ٶͰ�5�E&pyu�w	�0G¤��	�&렿ʛ�t�$h�Rb���C�n�йL�4�t�{?	���F������Q�2�y�_��B�L�e��ҕ��z���QA��]�?��E����o���a�w�nY����)�&���\�xW'^��ϰ��s��\Ŀ���ε��~{�2��г��J*.��[8C)	EP
��hbi��IߢL�D�ߕ�� p���4x�(Pl�}`O�zq��i�Y����9��]�
n�q��M}R�Ie7��gVB���8ID����o���cҐ|c����ZN!��S���7����x����Ub
������_iP���A��4�5���Pp�;`��TS>����0����h.e[�ua��Q8�Z�*���m5�ԥ��Nk�&�4��e ec�c3�ׁ�����8����
Q��p��!ɦL�މ�}n)h���/��������>���ܩ��}�����r`2aE&U�;�Td�^�lʔ[Ҫь��W�t�S��z��_}}�;����S^\2�7�2��;L���ɦG�`$Z{$��x�c>8��sy�)�ּ�n�bI��`L����L��7�r}H����-n�L�am:��6���%V�e���������0!�a�{��5�C�wաۿ�4�#i���E�Қ�zi���}�]�&�%͞I)�Lq��Pl\_��R��C`��&���|�&p8���(��J�p�X&G{V���{��0�bm��\����>H�2�ѓW�8��'t�j�U>�ۡnƄ]������*S�x�LBň�8��C�?r�\�Pu��4Or�?�h(��R�2i�#����t��!��^��Ŭ!��yu���8�8�[�B4��|Rn���J��AJ��vy)W$�e�KrR:��5H�2l��T@������Zʮ�'�����v�0U�3:E�NG�2Ә�Y4�!	���A�o��~��HlB�`��JȈHs�y�vsze�X���]EY9K[�E�xn�!;N�
�f�ϙ�	���o���2FrZ7Е�q��=�K%~v>�;�g|����S�9�7�G!�����2([���Y^C�p�/bl����Xiy����5�	��s�� ��P`b>ϱ�W�m�K�0 ����{ �(C�@�'��P`k �6"pP3jS��]5�(:=�n^��4�n�w|)�s�����zk�jv$Q2xB�jx���"-3��������2� :�yT󧄺8 �l�{P�`E#��~���A�($u�j����S��nKt�5+{�{����<(,��������b�3��]L �E����R�p�����?[���$�gЇ~|p:���o�����j�f�����b	�~��fn�{��4�x!�6�]��܎�>��t�{+'� ���F�SM*L�ţ
�?��B���#<�ɫM��jŠC��#K��R��~K<��W��3:��Θ!4U�E�Gi��}���N��	��U�<@�dsxI�z���g��1��'�t�?\ �	y�����=��5��:D�Ғ�<������<��r4 �s�'�%�����)���鯇%0��s�yR��r�Q��Elt��L@���x�vA�l����3%�y_9΃C2����`�(l%�9�N~UU�/_/�:/�:
��e�D������ϳ���D�?�Ȥ��qϻ�1�.J���7���f�-
�6(^f�yv�I�I}Ѐ�B�]t�%X.ގ]�c�>���Xr,��C<�ߌ2��8�03tհμ��+R�G�&�J��}�S��&�������Ĳ���g�BſZ{[Lx}�'W2��]�T$��
��i2�vw�q�����Hp��LAI�����Ļ��/���[�O'�P��k�O1���t�-�q���8� ?KÒ&y�yc�Tׄ�Jq��1�swOOl�������+�W�+k����	�i�L�j�H�هH��|g�y�$�;\���Ky�:"�F����b���h��Χ}�HJB
ၡ"3(��WJ�۳�����Y��,!���y]1���R�S �Bt��5�/�����hV�'����N�I�ۨXV�|���*�����V鐫-��G��u���� ��U˰�Y;���E폾u~t̒�H��X�l���!J��Ey
�HU��[�vZ��Q�P��#ruх։���nsoO|��"C�E��F���
"�:m�tF�g��>��y���"b=��v��tH%�8�EZ�zR§Z����_�@��N��G����^F�h�X�+۝�Q�T�f
�1����W���1�5B��~=w����� ���e> �����w@Y���v$C�v�����-�
���u�,N����>I�l�8M����s�������7҃���ì�|;b[���3��b��2w;���{�-�	��c+�j�W��Z!ȡ'��?�د�I8��`���x��;/�̸�r�yE�����},�r���\H!����q����Ȳ��9�*D��>��P�I��m߄}&�d�[�b;T7b_"F�^�Q��M^��x�!��?ف�CoF7����%�R�����{\
��"q��Wa-U̳��ۃ^o�(�eS�yN�Ւ�zI��҄����<+yļ�IG��c��F���E��#�[�#J5�0 ݙ�z��4��Jx�.x�Os���p�B���̺��M�x"O�0JP����`���r�9:+8��
?��i|�LD8O-��mI���u��>�}�%�'{��s_���T�ſ A�0d����M�B���*��������tA�p<BD�����R�)B�<�h�D�?��M3���N���K��|�0��mk �ד�B}Bau�@8�`�;���Ͷ6���m���*i��O?�D�䁑�w�?�壸����o���BZgB�� Hy?;`4U$�8�h���7��*����ldb���_ؓ���P����'�u�ou�I<���O��%=�uk�R὚�d�%L�bJ��p����L��,�F�һ�C�غ��_sU�{�S��];�-}�H��A�m吹����t45��i��'�cV��rٰ��R�b��y쟂r�}ai��O@�}��5�Ir�ו����C�k˜:��V���`6�8η�K�KN`Z1m!�	I�Q��7Li�SY�d/����x