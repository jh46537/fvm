��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{�&�U��=��Q�'6����od�F���!��>�RMy��|����K-�#����ȴ�a �4>��&kj���e~�S��´	9�D�g�	P�pPl���tp,��F�𪄁�g��9GDSɂ���xm�/��q��df�����c��M�ׅ�ݱ榾�HX{	F��K�P��Er$�P��QNƮ�݄w��gD��h���k�h�e^�P���M�+�~�6W�
oV�$K1�#�EA�8��WO��mBüҚ�Gs YG�g3δ �3��Jn���"����+�Ԅ�Xɡѧ��F�~�'絵��'����ϔ�P����cZ=�
9إ��ν��'E�~(�q3K����t�xjÿD*���H�������X	��޲�k5��(��kܫfsJQ�����3��'He-�O%�f���P�]�%	LI�W�rq(kvV1Ɵ�ѨG�}�0)wPDF�Ċl?��Q r"ɜz=g�$3T]:��"��0�d"����f��9�LbWlY�3]n��|�.]���e��0�[�Q28>-!����d>���PZǾ���n¦���b4�Η͙�����
/�6g�񛢉`p����z��|�}ќ[�� �S�|x!��i��#cVf(�j�
��d�_���`kd�AZtI���|�wzL �<�#Tʉ���<��.[�6K�:�vC�u�P�iD�s��`EaZ�y��BC^=��������!7�j���]����S�yj��7*y��<��m������� o�-�E�~�!< 4Z�j�9�VT�=���@��*^���@�V�.a��7�@$��Bׯ�cEh/���j����צ��  ��f��j8�JBJw��WA���DnAQ�E��Ò�w������7���n��G¬O�>
�}u��S�>>a�Jh��%;K����Z��rM.�
*��B	�'q�ҿ�%���[p�kʡ��0�J%���a����#	ن�4����°��`Ms�u
��>)� ��r]������֞�	���/���3��|�m�H�I5�
��=���W`$KT����W����*٥�R�n�\c���9`&�#QZ�lN<��W@=Ggc�����E���58���4�_7\��K�����'��ԅE��z)BX������o.���T�Dtt��"��gB@Vq88\���u�/� ��
\:w(����]��9�������]0���6���\��Ή�>��n��q����I/,�i��i�!���VIUX��3�j+V�Ό���d���ʵʒ5� ��E?"yp�Raw�O�r4���w�f�{X�k��Xg����D��r�3���g�-=����6S}W�\?��p�|T�׍�W0V��I��S״�
�&IBt���5G�)�g!P�k�ߤ��=:Wl��cW].Q2/��bp�F��U�V⷏Zb�&��Ac���[,�]j��t��W;_e+��j�U�m�r���m������!8�U���u_�R�l$���N0\��|{:rEP��.��3bU��U���,�ҍV�=��_�&� ����7s���� tY���G8����,��?�<����������Sn8)�-��|��Hc�d��H�k�������O�6��*��i'cW�`k5��^]<��9|�A���z��#�C�0�k|2LwV(�L�U�'Ѱ�X.-�����B�aՁ��p������E�����.蚍�R�xt-�/�4$�$DjS��8��u�\�cߕ�Ĺp�I��
��m5/��^��s�����xo4
;ك͔�۳�cx��@���t��= �p91HvH=��V�;�������8��t|@<ս7�\p{yE�Z.1�(>k��uv�#ML�3hQ���7��&TWe��՚���m����8OH]0�\x��gRpl��][������6����$���!�g���}w*���[y*7�N�ha��/�@=��)�a�-�A2���ȣc�q��!j�EkU����M&������5�4U�z	 Y���8���.u��`�i�A����@ߊR5p�1�$Vwԗ���7�U�� OGڡ��8�x�b
�%i~��h��H&l;x����P_���yřŔ�Q&f�����<��1M�M�]i5NM���B0�=��퐚���u ��kh9����Wvl(�v�@�/��9�r��D�wQe����oɥ����EO���1� ����E��z���V�f�C|t2��l���\<��:	)�I��ۅ�_��9������/*��0��R�j������Q��UWc�{w�ː�~�?f}�(-3���yM���
o�A�z�
���SvH��ES7�Tk��T���P��PG�*�(�V��q"��}�i��w�,�\OZ��P*�wqs�v�]��2t�N�oQ���#m� Հ���HѺV�b