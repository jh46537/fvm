// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JVJFXQZ4a/H7Uvk7zSv1R4H9skVs1RXIDK44jOgOdrEjUqesu0CW+/M8rpy/U21T
KxpNzSL46PWgdHpqeSwyNiOl1v/rG68S4tn5V+P+kXWL3TO0q733kSVYHNrT2jev
iAnluKGeC5KF/rfU/2Jg5+cvMtD4rJ1TCS6SCWUUOSQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1680)
lbvlqMdAh8PnV/KutZdnaVzkY5xlmVTb9WyEtIObN2ei9CT0yzQ4n7ZwqaLxgD1p
KsQ6co1I7QW/KlDGYrLsnIqu/E/8yhxGrHC2BWppRiqdxXi2lO/kcVL25515eA9f
wHLLgTVINv4LKK8HCCHzfo9DRSn/wVw8GwHeaOIxI4O4nkp0YrR/p96bGNQwVJHS
m0H8Na4HOLlMYKdz4RLsKRgWZ9YnRouHCF/muwSNwXSGXMlSoL1TC8VdE/AH9Vfb
Qef3Hj60d7di8Ln5xLtGbb+lLT2gGiQzUz9sGHALjCU0DFBEz6IPUgOVpLwGas/p
c1oKY08EPVvqXURchZE7hefBtnxvcivp+bhuVJQQC+Jzu3aq9+bNFM4kLq7Pm5N1
/RG+7aWFjX1mAx6HXPbltZyHsQHlGJY9QkU8iyeRRDFkZ324rCFBO+rDqnQotFqN
k1Mnfd5avCwMnzllGLifoyu4ahtIZhy9QYjkMQ/fqcNLs/TEgC3f9LTygKHzDT3T
9t3hLZu6FBvB3dVEYPDCWz3Je7zAOQMtX3FqyeoG4WBH8eHUhzvy6ZXlgyf86ItB
Hwol0RifinthSZbh0xGPnCpi1U6Vv37QJbBZHWvoQSOF49ufkb2PSJ6dM5AYug8t
XrE0Kpsq381v2C5wQ+onBtOKDdEoxL7mx1C93bgVkH5DDD90onpJIYHokIgJ0NAP
6DMBhidiANggFmiaPSQZQ2ZPv2efUvxoEczrZpJE7BpnacfV8VysrECKcFmp60XW
snmh7ivYhQNN0eKDeig0GpMRvGhr2YN3OJqKB1rfgkCdfYr0HDpyLOypiRdqkRND
NYK8taGEm3FOJeORKkQ4cat88fmzesaq96l1jYic4wL2CbX/NJUzQ39CsYHs0M2p
vBXrVtZE8SpBL/gU3mMwU6h4faX6GCcUKxrFxQNvpUFarwrZe7UPbmuQgw3cSbDz
Zd6QkZmU5n2y+QciOONt/mvpg54e7cjC2ZUP5UINYFEEG+d4V31xsIfbGAV4mjzR
JFUR9TCjzG/OPMQDM2CAcdpBUsZoIWmq8PEgTvYOywyDWjS0xrhm5VJcJfGlo2n0
ydvU6xn2IAyj7OJ4TV+OvxXDMXXuOdNrzE2BIpdj6G/Hor+MQA0siiHfy9pH3IPo
BpjLeLzy62hm6egmoe9jotVXdjqOPqtAhXpkJKBbDmPz8XMafeG6fsoSQx5UR0Lq
5WM0j8SlRKBm2dZNknqmsCsa38qZQAmHJm0WL1J87XX82SmhDUwDDfgcqQmLF04q
HkDAgLID2o9Ji840OxZN5haQN/uli24moimvsNBSkBYHQqoGQh1+zbDRIePxyPfV
oSV/+Tu5HN7LV6Mz6L/iQ2l+K0wUPjYkSktQPy1XCCKsWcqFpF5Y2wCrXdyRShgY
rDnPh4qcR0xFInDOPh2CHAUUZob4Ea/j1O9RDtQOpo5tAQPuZmp7ZiGAj6cJjHTT
rg+u/umISs1LK+uT02T7r5w1QePVUEnWrem78dzQUIPl4i3MC9HHlhFHem5Lcvwr
whZVB5Oy5PGHOTVgNrTSkEpi84kQslHQEVaAPgDNc0/jL8AZEoR4ZQDJuq+MAkFD
gCvnwVdW2cx4BLMvbf2xmsKRFatZUhWbBwSn58/8ZQmW9Ob0hczQmST+ZDKtNQ9g
Z0S+T3mghIdP6t5ncM79JOmwnRcObKtMacOU9+Rphlqo4zOlIuUfTWpT6Nk58KLk
MpsK0kIz6uUDxTCWCcIYe1uKoCS9sRUpjI5sInSoMEYVB+FUvsUEaagcnmw1ejLf
N5jWmJlE5b7zpJOc2b5bTelqWlTm4FWe7c36HCH225I69AaGO3Lg1Zt+sAuVMZXW
omiMXA/icwK/cOiNU7us9wepm9b7t/L5XcMgvWNc4Cg0JtnQWxQRI1z9W7JkfST3
G19WK3SI2F3tHqtLrvmeyuXrq+XV3TLukcpme27gxokAbducIPnTHb2wAbAbtMIf
3WjOEjV6j9KYIggtRdYC6XKtMvwSGBXbAsXsg6nJd+y+2LIRVXTN1HuSe8iu0Iqw
aB8HONGAKW3RLfhV1de6AIxNvjnz9+yqYi+wBn0CBW2dzAhnwGqJIIm6zvbBPUO2
qu8Li8IKPSr/LSL6/g7igt8/ybRdkCPP8YDenjkL1jH3s2YjIG6l5gzO0YVy2Sef
s+DsfO8Iaf11ygGho4ObXNgcGUL24ZSmte+f4dMxIgZkhcL3LhmXxA6XlEVMhXJ0
`pragma protect end_protected
