��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&Y�%�ddؐ����7��b����T ur&�\��m��[�A������0�jGY4��?�EG�c]e�%������+�/R�{vK���(��S��(��2�]���I�l���G��J����ŋ�[&Յ���'�9�!�)�ض�)p��N�4�SŸ�I�B�1zE�y3H�@�H�����Ӯy���T��v������n��Z֥�3{�~�f�-�B�B����)�FX�(���Ĝ$����|A=R�p���<�8�����*��K�� �<�\��j�܆�U�C�|��,�P�SJ�L�+��աf=R.����1����x�KC�N�|����ȭ�/�]��ND�w,�w^KQP��%5�������Q 
�פ�o��1{BBc+�o��H�7a�B��z$g/�}�����9�NB����͹9�$�<W�p�1In�B�ō�,ⰰ�Ĭ�fbvVC��3'_Zʮ�K8bνnv�}� +������$������cB�t��	���m��/��~�kdӀ�]�)��z��=c yb�'"��������<P�:����U��J(-.���"�S�\�a_�-�#��,=��H~���"}�1�Uwb�br�)d�joFj_��}�-#��i6䰂6lsQ���:2�X@
���n�N��X�u���zQНf��
���dȭ^����T!�H[
^z��ͼ։��$Ø�!�P���I�6�}k���,�<�;���Q�x@�ݠΦI{��r�8Ϯ.&�3�Z�yñd\{�뺨4���o��53y^�``�� �W�	!��o�T;Å�K��� �X��IE�b9�<����F�Y�D�+4]o�ANY�̣����^z���4���KJ�����a�y��@0�1��N��R�$��=x�oz�|�ܰ�1�{HY�c[�Gc���W2��g�_깾��9����<�P�%4B�]�_e}]6:b�aԘ��N����&����;�.������q�N>6�;���5$5�_r��[َDȞ�$�"rk���ЁTҚ,����D������<
Ss�F��s���.��S$�pz��{6w'h]�2v'j��{y�5�Z�K`��us6��D��`������?�D��z�T��p>�L/��0?�Q��F+��n��fU"�u�����y�I!���\P�1Q�i��O'���~1�T�^��>_�!�5�0sԎ��חQ��s�U$���Y���m`�ZG��g��I1j�L���/T��p��C+��Z*��W�u�%�~�4v��-�p��T.�P�o��eջ�T�!�
�� �kl��y�����5[�E۰��+/*[��c#�i��/�!��P�(�[ҝ��簶C�T� E�F����\OiC��i�0���I:<�}�7I�D��~�&b�����]��6=�����w���\8;4k�BSu��7m�u��v���}>={����G���O㻸KbZ���z�aS`	)o�������b��CPÐ_�g���Ȁ=e�Q����˥��h§��G2"�V��`>�[�d�0-�'=G@���(8|�A�ixRbOܤ��1���Ю�����&�6���.�/@D>G���5�:u���V��Z��\���E�r�}��H���*�*qPޅy�
F<�Øomz7*����6Md�8r��㉎��`_2δ;P��Ɂ�� Lv��\-�B�����Y~�
���� �C ���6K;R�o�ɗQ�ۨ�=D���9z� C�e�뉒��i���xp�L�e�޳$�zuk�Z!����(_�~�����E��
���y?�"��v=kV� 5\)';�y(�@��<�xyFJ8�8k���D�)I��E�0�t�"%�<���PB�+�}�T��Nɍ���UڊW�Q���/��lË��*<���,E=����&l��&��}���GX��O �s.�=�Ú�q�
T�T�ds�����C��$�	
��!� /X������N�e�rn[���TRCB8�kR��ޮ�O�B��4W?���u9K�Y+��(���� �:� J�xv���-�����VuЌ�K�~�m��8���Y�E�x�I%}2�=#�2g�������T�qv<O�S9=<�`���R���#Y�6���)� ����fd�����k)�R�>�Ӱu�m)T��z�,uR�=�F��U�+�V��5�ZБGl����(۹i���7w�\r�9ьSklڭ�}V�_[�k<�
5��6o���79���ݵ]ٺ*/�)�%�A����4���l?�5��������h��-�#��7#,����0�p*�����/|�����m3�]2�h�bQ���Y��I���0���T�-�x]�n��y����;���j�%��Y���\��>]�X�f�)�	�ܱR �l[8����p�1C2�f �jO\l	,�fg&��?8��ڳ�@�菆�h�߲�������p\���.RN���u[Y�:��Pm+��T�[O%�}��!���-��oCNS��#��1�6�g_�H�܁6~��+�aޛN4��!�c�!�f��M�c�V�S�V8 �{�6���.'���������r�n�:>�TI?�+��]S���M�b�ڴxjr>��k�oXo��^�t2�w�f��&��'@{�?,Bm�8/H,��d p�g)�;�d����7L�+��K�X�NW����m=�x\�FB��^W#Ҿ�^������ fJ[�R��ֹZC�������k���Ç�G����$�I
*�l����?C�:��Y^Q���p�z��Ԛr�yM�M2��!��Y�Wf�%?aOS�!��f��},�q�?�%��[�|qt��#xG?���[\ӷ㘰d��kو�)S������.�h����a���x��Ծ�ap��ZZ��EQ<�R�+�"�9�G��.+�4��.��'lCi�HD��{+��X潮}̔~��;ߪ�!p�
�_�w:��ߴ�	�.�^p O{�`6���`F��/���h�)d�]��H��U�pM)40����1y2���1>�"W�Å"ZG��E[�
`m��!K���}/��<�"4��E����|������4+�[���Pג���n�����@�����@���� ��x�7�/	�홱#1������8`��$�M���ßL��R�L�Fh+@�d�gH$�O&7 �VQ�H����'|h�B��%�F�ю�n(��cg� $�s���ݗM��;��:q���զ�6��弌5yn=��y�ml�f���2`伦㒲����R������2�	w9e�'�G=GG+�c'���ܚ�:����_,4P��<�s�|q��ˇRgDw���1�X5�[�D�O��������2�ꎎ�w/
bcgU��G��tzΨ���3����s�{�l6���:�8�Mqߡ}?-q��a������zj�=bǶ�5�����ҵm.:B����b����ND���-�Ps������mM�� �Փ�#�i�l��ԁ��\�\�L��b���nd���VW	���ﺎ�}��C)��X��F]�:��i	�)�ЀW!�i��L/��{��DRs})C/��1(JZ.�S�x��s�^3�9M.�ŝ��x�,}<7�������k9EHB��p���+�a�eŢx^�iQSm�R�΅2y/ݏ(w��K�f���k�~$�N��UTD鯍y�ݼҪ�23��ӷr�w�W����&�l������H�����
ٚ�b��b2�����Ǩ�~Mm�/�$��<e~8R��-q�^��=E�̠�&��Q�`�]Y,��,�� �`�M�)m|dFz"E:@��v]�.��9�a�_t�R탫��p)65��4p����V+��}��X���6-W�����i�{�䒭v�:B����T�wWϡ<��MY�S{� ����tBk!�B1��Th��?Q�ܚ�ym��ON-sfL �1�oS�;]vnD�=�g�4��<�C�r@'�D�J��@��%_�UHQc�@�g��ayl�>G*6#㍦[_�領GR� �
�v�5<#�E �;��B{�6��~��+����� R�̪��!��/��W2�Ȅ(�R���������Ɵ��~%А��	�W�!��:J�/�T��T&�9��-�d@�yI=��i!��1��f/�=ݖ��;'�ے�y/(�Tۇ���̤i�w�}����?$���R8�rd?*:Q�'����ɣ\�PT�r��? #�n\uƘ������I��< ���I�����~t�]��8gW`Nɢ�65����Ҭ ������`H���~��D=��*%��0�4l�������3	4�ˊ��E��U��[�x{�E�-@�5j��8��0\���_�䒺��� �0���k<���_��׊�ԊVe�t�O���:��ӆV&� ܀����m�!�3RX�ɘ	d�9yo^��LNJ���#;�\�L��E6[�P�c#�6��FT��S/U�KK�7��D�|�_���|d<���m�t�j�5��Q�_����Ǖ`��:oV|�7U�^��*�^R.E&΅��t��4s7�U0�\	�Mr�p�.~�w,jY�[�(�̟���8M�f����wj��kq�@A�����]�*ۯ���������