��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����,��f9t���3>��Ձ�A�7M ��uj��M�0��{�ơ�Wa=Kg��!洭D�2�&�6����2�����X܋��x� ����G1���w�S��3�C�1�9��1+CH�<3�vwN��F�T�\#[�'I���ҒO*K��V�6�k%���D��Sn�&$Y�au��Q�/���OO .�XS}���9��k,[=0�hj��V���w��:g�!,;�(���1��+�\�dn�!��S��Q��CU6���>���m;�$��z�����So���88ׯӉ��zV#����;��lbaᩇYU�k*�|��	^����p��O�(f}�NA�	�g��5cA뾐Ki��M�QY5�Q��O�H+8a��)@���Yr�J�-g���ҽl���,�"DԞ�(����#�]&t�Y~�WR��]�ģ��U�&�� �y�]��A�v-��=���b���=�>� �UI�eͻ�_��5,����?��r#��"M1<cUc88S�"�w����
q@u;�c��G!i|�x�9V7�a���{���bi�_��'N[�Q@�.U'�"��$ɾ�Knx�_���E^[2Wο�����.�#�J����)�+F����z�H3lNÅdjO�ُY��J����Ǵ�J�*�>1!�T�������R�G!d6�%a�{�x ~�ھ�9�"�1��m��e�Q�qf�O9���!ޜ�);p ��9R�Vc;Q'����8�.mg�X �b����ӏ,p����1�)�H��qH����3�g��7��'CRԸĘh���-r�t�!�h�ݍz�I��T1<)0y0�"�IwZ�f�:�v,M�0zt8҈��ȩ�b;
g���У�4$1��Qcf���č�p|z<D�(���
ٍż�LS��sUF��_U�?�0���^]OLq�����u��	Yy�����3�5�@k���s��q���Ɲ�l-R5�Beᔃ_-��A�&bf�z�������`mT�1ɥ��c6'�q�e�՞��A?��V�j�}B�{���	t�.��#���q��Quk������4��[��w�A��޳,o"�=J�;��̾�(f��>�y�8�wd�S��bo�Ii]�yQ-����V��Y�+���~���1��D�v��x����.i$%�Ka�x�؛��_�K��U�@T}w�X�����ڠ�"`�/�V_h��d���@������i��n���)%4⪡֢&��Ӝ�@���ǨК�!6}�ԍy!�J+A�/�`#Ģ�U�Mj�I�F�Ath߻�$Ϝ.O��N^\@�}���ʱr��)�s	j�o��z������ uW���C���g�e�][D2tmɲ(��}x��{W��P��oR�h�O5q���T�%�c�.��y8�N��£U��atN n/�~�ȋ99,�%��ޓ�����J� �;� �I'�����m��[��k`�K����NǗ�#9�]���M���^f�;�Eίޑ�P�I���������"�s��>-��F6���f�@100 �%�2�-��3r ��=�@:�!
��8^��k!.tc�0Y�.�B�d��Z��)��Y^���$��X͘���G�]^{mq��ޛ�R�BF��0���U���0FR~�kdu|�1��q�������y�k����/��z�t=ؾvί:P��y�CO���=ڗV���e�K	a�J+�c�|�n�+\s���F��<�cO�g��Z�8/|˽߮>�YN]y�/k��a���IXp����Z}����x��\��y���os<oK�f�BL&k�7?R.��[@j՟T�z:�;tq�p�~Nɻ$�
e)���np!����fb_�Fc+����f�"��P�s���s�~���- ��� p�7����}���g|�:����{}�I/�"%�M��R���H-M"q��=s81*�'}�U�Ů����w@V"����[�xL{�hW1�ka�c � �EF�����5x6���)�'z�).'g�+
2�y__x���P=~�"3~_q\�����C��7���I���M���A�i�R�fx*֠^���Ff�Fi��JN��"�����x��vV�k����|^�l|���$���o��s���I	Xyw8�]x���}�����5�4R�׉�w��8�%fw��t�/��m��/&�8 �ko��2j��ŗg���?�^�W��sM��f)*J�^�6�i�˘$Ѵ�8�$�x3f��>g&|�J"]��#q�G���y�]�d���۶�	���/���|��3Y�`�ܜ^�7{#�*�Qǥkj��@�p&��7�3��U��a(h��l���&�'RfXY�o����n%R�X�D��l���_u�e��3k=]�=�(!,C�`<����H�g���D�Z����E�xȨk�@��}[�d�P>����?^~��b�ZN
4�^���"b���PKF>R��&�GA��}<AkD� '-����z�JUOS�O	��H�O�x)��z�Yv[�醌��C��h�7��v۰�vը"^�v1	�V�uDb�=H\~ǘ�zc�3nĥX`����*���
F�U�X�e=O?�6�#���[�1z�2�2���N6>|����a��)�1x�p�?5U�b.j��jcG*q��e�̀�CuDtU����T�j����雍��cK���N~��bn�g9�	����$�#��}K��E%�&��&�)Y� �5�$��f�r��@6yV¨�t.O���O&��@���U�/8�����
�ת_�����o����9!Wyrv���_���ܨ�d���(@IlV�'3�{��=+:+���z�j�^H�C�a	Y�v�7Dm���zy*��q <JG���-'D<B�]⠗��"��e���e"uN�v�k[Ԙdi@]y1aǨ!�����ǈ俶3K+*4��J����|2/u D�>�F�����Đr�pS� l�g�DeG�|����%�f='�d��Kk'�{�/��2:���8�ҟ��Gr�@��z(���^��v��|�ɞ���M���T�v�zX��kظ��)>j�<�#� �4�ʔ]�9��Ϯ�� ���*~uq���^`K�`�V!��I��6/�k,��F![x&�,:�t�AйyO�zϞ�R�-��7���^K�N@l��d����Z��\�qr^�՗��%������E���X��<�0�A��]-�{(\��۹5����r���ȟ=m7�իڣ�P��b0#��B!E�2�Z�"p�%����4cv�*��_;���3���U7h�@�"�J�t�_�HM��i-L��-�q��0�~�{d�+����o�9_��m�M�5~�j�w�Qn.����F�q��PN��(�) �K�h�KʺE�zڒ������J��Oj��1�1]��V.fl<�c�òK�3��?>���jW��C��O�'o�P�~�|hJ�bc2�m�6�t@D���ɳ��s���V��Rnx���rO��� �D��2q�ɼ��˘{ȥ�/V�x�!ZDz&
�1Mt����U��t2����T�`�%@�4�h9m�>�)�����y�5�񰤲v�
5�0�y�s�I=�2T���3���W Un��Յ�dSE8�I��`��;@�eζ���ӕ"�K��J�M2�Q�C���	��p��;��87�V`�
6��i����sfy�P�b�x����8�B�@�U��W�69��쩦�3y����蔯�1�j�u&�{���ղC��9��G��e����Iw^Ddh��':����}UU3����v�P׽5'�s)���eW-^����OY�Q�`��$@�r�;��i����>@Zk�M�b<5��ur�9/֚5	��$R6*�VNg�zS7HFVa��{��`�=��WP�ӏ[O�,.��Ɇ���*���M��1�;���j�r6��Jk^��z��f�+��{��G��})��#9�[SL��#gR�]�f��Kp�W������g�D.b�"o�?p��ݹ|�˘1=���(.=~�s�;�	��0U�C>��{3-wP�ф������4���p��p�/,�=��hu�������~ow;_x�m&��j�4W�T������dzF.�o�av�1L9rQ����;��<ZC���xm��;�֨!�R�GZ��F���x7��,�8jƘs7�ϴ'e,� :��h��o|B�����t�FO��|{>Lg�����4���J�9k�x/w��\�!f��J&��:־��͆$x=+=81锩�ֻ!a�P�|^��	�遦v`e/򫨘MC�j�+6K̠�s�坊(������e��i{�����Q0���	6�J���ޞ(�V�L�5�:|�uГ�	D���+�MRpM�ېH^g_.c�ޖ��Mû:y1C�=�n�*�����1l�A��:�������_�~�����9�"ꤿ5A�Ԡ5�����%�	ɍ�z@�^����7i* �75]w�Ǚ~��R�O�e��$`��Ǆ��c�� ��;�6C���_>��/l��j�w���������됛�a��l��aF�s *�j �\�Lt����#�'t���KJ[[�@� ���ȃ��K@�i�kz�bb��R'���T�ו%�˰/r��zLÞ$��I<4�$��<gݵ_�)l���)�Rt����TO�I[E����Ncel��3*ϰG�Sm��!j��	]T�S_�Z�5G��?d�<��0=P農K�5�$����Kr�}���)�� ������jn����7����2�y�`"���G&��w���&ܬ�Z�WRe�wy��(���o�L$k��9p��ኜ�hH�֡���$�DI���%Y�r�N�rUR��Z��>�nd΋N-,���l-�ъۺ���n�=�􀻆=�������s�F��)�>��`����ZNe.�/�L�Dg ���(Rm1֣7�5C���=��W|bi%�;�&���N(�Dc�J���2�!��=���$��21C��)��. od�yt�~�Vɀ`Meb��$���3Ж�9�:X	*��#-{�8�C�x6�r��޿��|wN��=_g��>�u6�Ş�������K����??$AL�3)�ˬ�y��mM.��[�n���Nz��z��uA�D�Aw%\�GI欪`�}��_*�r�=Q�Nr�T;�ۘ���s}N�=WM����㳟����f@����l���z����۝��u&��o��S�Q��*�,�=�d�^�]~�+�V@�Qc��Rw��j`�G�1 i\�U����
�n�W��|���A�q�lw'����|�83�*Yl��}���?��Q09�(�-a"�[�kG5���w 4�S�N"sOJnZ�s�88]J:g۬����\r&�Sc���t�>l��5�m@�,I;�b�|ϛ��0!f�+ſ_C��s� ���P�t�w����@������QU���|�I�k�2��K<(\�ϗȩ����R[�m�Z[�D䌮����u? F�沏����#�W.�����肣.͔ސy�wY,�2�|���i�B�-��K�5t��)�ۢԌyj9�@�K��w#,tl =�����{�)�g�{ʭ�9���
�1�y�ycجZcjy�fr�\.+�l#}8�<����Y��l�t��n[(�{(�U�:��!w<�
p� w�vg����9� �.H��Y�����;��͏;X����+��
}-2Y�R���R}��n..��͸]��w���M�]q١]g�9 ce�:uL�㷾MNV���\�fr^X����rx�A�v��1�����"Q:J�S�����ԆԠ�h�b�YD�	6���X�1���ey�岥��ě�8ԙq&���yJ����پ����I���eL�D{�Պ�G�����e����=�r� ������/�?�q��PK9E+�p��P��	W�l�$u"!���ٕaY���֌�R@�:=REhi��N����4�����c�@y6J�IIN�p;����V<t~��|l����R0�	"�{0�����i�@��z�9a1���1�~,���Jq��(��fI���ڎ�j\!���]�a-a���<�,���_3~�غ���nTc��<�Z���;�ԣN�O��F eH�֚���ӯ"7ԴV|���N�8�kؚΆ�m���4:V0���$�pF�@Pm��+Ҡ��k����0o<$y��8�H�jt����BO'��%��UmP�����.�iZD�,�0S�e�@�l�����3��#�pZ$V�����������6
��D���;��D]��>3��`)f8e��@Es��s�R�2x}�/X|�g��?�O������6>�O��8�ڝ&�:4���sW^Q1&�DF�tYa�;.p0�+���]r ?W	r��nF/�O�6���U�qLr%r���2���{"۰�Q/��A.�%��o8
�g�]|���Yc�!���l|K��I��(�8Ϥ2�%kd/����bG�&����� �.��
��Sx����n���!�w
�#l<�6�3�֕�)
E/7�I�c�_�y&���Ն,	�
�dW����҉d+�
W��[�]�4�A^���'w�36�o��g"��cͱ��Y`�/�Բ1�ŘF�	E^��
*��z�L��x/�i[!9�W����#(��߱a
�5��^����p�
覝��]3�j
��������	�hz=ݩ�+�{a�D���1��>��6U:���0��d#WDW�.2�MlÆI?_t	b򧏗t�pV�!]'!�fO`��8n��ٙ�>=Pi�v��\=�!�0C���e;�P�Da��*�)�F�P��x;���O�l��78i��x���r#d�s���q�>Wd�����B E�Px��T�Q	.!�^��j��
o_S���I�v��%�K%d]�D|���ګO�� �|K��H)B���z�w��gwntuS+�A-��E8dCJ{ٛ+��4|��+�l�GM�@L:<��V����ֿ=ɛdEy�ݞMB����k��C�;YR��M(w�L�OŕV靪YͿ��P�QT�ԞMAk���o��ئe�z�3��UD%������� ȃS�mo���#)y4F���܉��e��U/u�Q����?6,��[̭֚���v�������ֵ���[UO�P�x�I�Oi�o����� ��������t[	\p�@:�u��a�[78���G|���fݞ�Гzn���>����d���?�&���U��B�]A�K@���E���f/U�C�b�u�հ�����?��ғ�=����am3��k�ZQӀ� �ᣊT�g>��I�c@՜��1��x��>�G��Xz1�(��ֱ�~�$��O���W��{�pCQ-F>���ch([M~�g�!������b�w��M%�!�	u�كԮ�{���IdmA)�02�_[��DwxD*��y��X�mq��ч>f�����јsL$8�o�u��� �V���o�|��6jǯ����o*��O�4^ �D�_��i�8�����2?��ʵ�s�Ox��F�.�G�I�c��������V),l���$f�~��S6�g��9�<��{�%����0 T�}�*"�QZx�|�x�����l���h~�o?Hb��.��t�f���pIv�9��>�Y
?�՜�]� ��c�Y��e>��n�9yh�ApT�`KI�57E���V�ou$�o̲���:;F��}�O�� ��3T��aI�i*7��$8q��x|"�?
���{�и%���Bލ�3L:qV�z��>����W!��m�ƚpۛ�+�>b��Sq���%:
S$�W�;m.�p��V� aOF:���KNYe����'���bz}�C�$�]�V x6�$t�\/*���8��:�iM�jY�)��|Y�M�3��AA��.��x�,��!�&ʹl?tZ���n��Z�A���	�;�;�톭��?�@��.�����4�4�xB�
��'\:��0^x�-ً<=��ǡm�PL0�s찠�#Ҭ5�-��?��?�71�?6�Hйy����}�Ͷ�q��t��Q$0���v���O���YNd��afI0����������%h�M��k0{Z�T���R�B���.�Wh��M���U�0;9�ݺ
�^�jw���3�;8��Bb��-^��ќ��~})Q���	??񾛕I�?������B�R� �9U��#i���5TM�����cGRZ� ����F{���[�M;Kr�?a�{p�N,(�[�S���n�N��n�\�VȀ�i}���AYi���c���t��%5����M�������Z��Dߩ�a��Wr�<V��ZVP�o|z��X1M����]��CuVc���ZY��鰶\���.J}�"�툤�D�Al�S��;-_�Lj�F�J2�a�p�i��5C�wE>{��[��^Yuf��9`=��&(�p#��� �h�_<�Bl��1�9�c���LNY�c�M�����S�G%s�o�}�n��3�g��0a�V,I�Ʉ�ԁ�P��ӫf���ћ��MJx�T+�"��A��Z(���'�6#N]������R����@�i��@h��*ͪ��p��`t�!eO���Q�V�����>$d?�W��v�*OI���_�(Uy+H�}�d�[ɺ�NѺq�F�~�]���ihǱnl��h:���6j����Y�� �.����~<M��&�,`�ϚJ��Ae�������~��Lh�|b/vu��~������f|�צ�m�I��Gw��fA&wTͲ��P�~7+�_'=� ����ř?O�8q��W�Y�����GS6��^{[I��gc��Pёx���YT=�	��R�,  �����c�dF�k" krB��@ש�`@��Zd�H����_��'�����s�U>�e5�ZY�8�acX�5�B�:�o~n���|�k{�%�貃_D�9Ͼ8^LjB��?*�5kv�]�!(��6а0M���K�SQ��}]*MW-�ך�g
�Oa�=�=C'�L9D9!Z��P�THBm�A��,���ɻCT�F�YUמY*936���*�*,GR9����9���:eI�O��V���m�P&�������'P�ߊ�㮾��^���\�o���C�ӵ�ll�9+'��TS&��k6��1��f@�myyqŖE�4�Mē��_`��Z��%��{�7w� d=�[aRc�����L|�����^�E`q9�$�D��R��;�v�<e���(E�c����
�N!_8��9g|P�Bˍ��Y�B+��@m��ex�H��B���g�hJ&i����s�I�#&ӓ0����~0H"�8-�����2�'�P gzm�����~�򪎪eq�px�[)�����c���?����]���F]_��s}AĔ�9�֑�S&6���0޸�]ao��0�_�+�`�y���⽏�羽<4-2y��E�|�G۲u��ʮ��������.��������mF�ə�!ó���"G�	y qt���y�^�|uusX\t?�s:nw`�Rr���2\:s`Zߟb������-�K)����;�g�D����� R��(RA��ګ�� B�cK��ϔ�~4l��L����n�N�}����	"�r���`'�tx��㝙�a�L@��W[��f���?���mu�(�3��,��t@�d�5�*�����*�]Hvx�4�wO�"4v����Ψ8.���b'>�@p�!�%�Y�:� ޲"��;�r(�V�'�f�`�"e��1"�D�F��¾U/��i������8�l�ɕ��R�ȝXV��t�b��A��̹�������Q�i��a��]�6�h8x�3���w�Cj��O�/['��_��\Nu���V��D�
k����SHM�ö8 !뼍\��cO�ơ�%u//%�rh�u-�G8*�{�+��� ����V��]�j�:'�	W�&�3UO����W��W\���D��[��?6�W����},��A�)H�x9���<�:�1;�F-
�ꍞ������z�h &q�/(����g%�`�=���=p�{�pg�� �	�%�v?ʏe�K�T��F
Gir�X�?�c{�\�I��ƴ�����q�N�~�=
��Lt2�jC�\F<,��1)A(�����n��fZ��OWI��d[�oO]���u�0��Z�^q��>�in�#���oh@�k�m�za�h�y�6ӛ�]��kf/v �<QFJ��A�p\A���X�,*�lz��Re�<l�m\āe�^�~~�%�ߘII}�ا���
��0�����,eפ�A,��lBqp _u�L��;�,�:��ވ�{R��	�錔�VQM��y�V���{.�oyVYa��'�|����=+`�%�u�&~�~Q���l �\�gf��g}�U�\��^�*�Iuŀ�պ���˧.
H��*J0qc��3|e���&�|z�\4�7¾�OV����Y�I(2aV�}yZP�����}�Ǐu�2��h9(�����jh}�?��#K�,,G`mVO\$h���E�S�!�ڕ�P����!���N������U��'�a;E@ ,�in��Ɉ�<���hJ���v�}%���r���!��Փ���*3�L�N��~�g2f��g?V����e�����͓-��19���n��Rm�B�8����TM���Z�L�_�^�e�	��f/OHz���`��1�����b^7��J%�e����7ւ��K��L �p�3IC����^4�pH�a�	�(����Á)}�E���7{����:e_R�F��{�@���Lz-l4%q}f!,3"To54
)��|�:��	�W�L,�u�%���l�
�l_�z\`uJ~�w���-��~)w��[�>T�� ���5�'!�<v?6���t'�׮�ɦ�gpw,��m�]tX��˛�v�aݯe�4�־�訪�$ �[@砟���S��n�<�)�����C������n���c$�v�w�����m��l͋����̃]�T|����~I�dQ�����'���6lOl�z�8:r��8��NG9�`F/e�;v�w�3�t8|6h/�.��1�W���=�!Xu���1.�9�_��j��ڂE�_A�kOG��aӤqL8E�+7h����a��<�U[ޥ�D����5�|{�d�ɏ[��7lc�sl�@a��2xW�1Q1����p��� ����|�9���2�ۖ!�b}�����~�[���`�O�g:!�V�J�Ã��\��M��b���7s�4�2	�y���c�����be��έ�]�j����޼rw`�a�!�vJO�'CL�>��V:�?Ԯ��1ң��ׅK�9@��+���T�o�h���|\wB�#2�6��H{t��8�3��X�������L������ܒ�0�u@�L����3"�8OO�-w�k �<�Öc{�"�o��3�oZ^�^��՝������9��-�f[�$kw�/Zf;��ς�Or�H������O.�P�����u&�2�*򃝀5�\Zg𤴯q�S�`˼��q��&a�����z�U�{6?;�����
yĞ��L%	�X��%��+�I�(g!�����\!��gpsr���6�:_�l�E��� m����!�i�DS��(��k*J�����R�?-�q	i8�r;q\�E^�0PZ� c�"�y���wų&'��UE�l�ܑ�U߅���r�2�Q;��9Ʉi���ѻ�??�`OPʍ��D}6m����~�k��D� �9�8���	��+��ƛr�w���
���H�^� m(ҙ9|G�֥�uq̂x���M�Eln�6���'Y���r�?�b`�[S�>�0���CR �v4;t��oɸm=x)�f����:,�	W	�� ���v{Mq��r���+V��l��s�=�4��Q�/ q�����1&�v�jnkHZ��� ��ғ�:lD�S�V�l�V����6�Z%ۆ��4n�
�r�PS�h�����Po<��1H�"��'eJyՏ�
��4$aoM�O�v���Ӛ<1O�i7 �J�6i�!�;3�J°P��3��Z����vv��(ķb{_l��{��kB|�	����X��Q�&��� ��-(��I������dt��¿�Q�`�'0G��g�W�׈,�����4͖��)����ڽ��n��I�{izo���@�z_ӊ�����"�����I������p���j�����W�8D����q��z��t�`����,B�Z���I�/uN~(���C��4��ە 258Z��&��F�w��Z]x�����a~J7$q�a������YP�Ź<s�9MPՋB������=�=����8��o�z�7zpGY��(��J�*0Qf5��;!�G�W�}}et��Ab��U�|�W#�����g�͌$��/k<�+�����&n���L�f��2���C�FͱH:��������w�K�A�Gk���?��`�&N��"�[���8�(�bȡO�d�K�m�kń	�$����O� H�4�U�j�+%���8�`�qC�����,��?���z�;Dϵ��m�yl���*,�*z.�H;n‡��O��O@4l�i%�yH�%�|�%�x���^���{�;'a��oK�/�o��mBա8$9ݘ�I��W:�q8Y@(�]?8&i�mf����ű0�*��!�$!ⅹ�K�� )	���gz)�s����h���� ʻ�J1�����x-CƤܩqԋw�'�C�p1��O��#�a&Tm���������Aйu��@XH���b�;�/�]$Js[����b�|���uR�_�J���zo�ԛ��D r$,R�Ԡb�x�E����D�5��4�D(m�B���L�zB9>Vc%����'Bym-��迊8�#W{�3U�4�?p�R8t2�\��˚��8G��պ"�#�XV
�r.��
.CX)i00F� ;�*W�V��B���#�y��r:!�i|�z���g��8O��(��_�1�7�K� ��|'��8 .j�(c>�̿+63�#�4�(( D��J���O<ƛg��:/@u�����t���]��v�v���2X�醴����$��ǻ�C*QpF�5��'�j2��j?�7,6x��f����*�^	��2��_�����8��V��7c;�J�>��M�+��>�;����G�'p^i����#\����`������|��|��;{��m�!��Dh|f����5:>u�,(ty�-�۸��emgG��i�哠��G+��gj��c���I�z���e<�������Ho���_�"�1]B�����\p���fqO�U;T�J���_���TLsr��LgrH��s���� FB������vau�(�SM���U� q��7��p|��[�mKeDjdI��6^�?�]2��D<�w|��r8�l��g_RFQܰx��W����	���7���.Y<�f]�۸��0�H��MHv�(�Y'�AT.%oǝ�7 c��1i'�>wcH�
���_��
b;ű��7�~���I}�4�
i�)ѽK۷nzb#	�0����ڂ�T�Ɔ�d[m�"h����N�;K*t���6�ėpŰD�{��H���S��DE_f��d�@~).�m:��f�D�{BK�<��?�u��v�
�ħ�2���󮨼Hp��E����@�%���^@����cDy!�`�K2]�P���	�������q?�|t13��B<J��>�<C3B��1�#��gn�Y���OG�t�j_����!��Y�$��ť��QK�Mt|��)�'�c?��Îؒ���v�NEcJEu����Q���},���5�׶�f�~��YDX��׼4jͣ��$_��t���z���VΝ����t�,p��5\M��]�U����z݃�:��W��W����U��Q`��3.e30qfR�BZH$j7Ѭ���d"��#���퍱�pKO���
�=Z`L�֮KV��9�mgzH��؟;������Q����������"�[�o���������	���R�4�I� a�&D������ʢ��q4ǵ2�Х�A콀��l��h�ɏ�|E��\��sg /N��ݔC�"��RrB�����4"S�F�rA��o�����aB�ք�~��0��ܓ���Jl�*�.�0���_�(��Ո��~��9����D!`�4��ڜM�9*i\R����b"�1���D��Ps�*�ؾD���<�-�_@�wIK�S��r�<�'ĩ�+Z�@�=u�Ji�wt�l�/�>g�4�pY�τ��$R�Eߵ/���BI���Jg�<s�/����$�ⱁ_��sR��e߯�	fJ��"�PM��������
�����r{l/Dݠ��#?\?�JRJ�G�<K�y9r E��C��F�sF���������}��<��Z���;<Kȥ�&�3t�^�jؒEH(\�Y���vʣ�8>����L�?xTL\QƉ1����gg_S,�:��A�^W�[B��@Ƶ�S%����_j��1P�4}�Z��qD���`�8�n�l�L�K]2��Y�����yʗ�y�s�5��kiP+>�n$a��WE�_V��f?��f�jQ�+�����+��v��p��`t!,���	�ky�<V/��}�^��x��1�ͫ�׏2���i`Yi�)D��`y��ML�u�`�_҉���ˊ靵WSG���{x2�f��΄�m�q���(Bb$��9�Wu��j��mG���؄@L�`�zj&>9�6��|'�1��� +B&��r��S]�A�R��h�ߒ�@W��*l�q��h�K]\NI��;�'lΤ8�?։`��#H�����HBj��<�11\_��H�km{]�Ȳ�������W���	F`�i�Z��|*L��t� �6��fX�g��<��Ĥ�Ff�m�t���`�1�=�-|,��!5GI��
�s�Y�!>�ViU7��ϴ�����M���	�G���px_�Z�Re�B0=��E`��_a1�j�9A�������$��|��.��Qܗ�iN�v�4C�v$.!̫�G�D%=�k��?�e�D�ܳ�M���p.A�d+~�cՎ��1�79���>��	��ïm�	wzl`��úc�4����4�z�+�pb�I�xZx�W�}�ܡ�'X���W�&�Ė1��`a��[��!RV�l�)��(!�<Oj��h��<�T���}��z�]����؈�-���i~o2��6b�<�f�yl���w�n�D�B׊	PC�i�
���\a��,���_�Z��B�:� 1�r��C�!:�k��3��=�h/y��T���� ��71I]6�������8�)���|�=��X�25%2g��	l���^W
A��lߚ��k�k�h�D=7��'��Rב"ZLݥ��||���<%R��%�/�=���͐O$3����g� �Q5���Iow�Z��x0� +�+�'|ۚ۸��"�C���<6�S�o�Γ�BTRy��-y�:�.���0���Z�N)}���GT��R:%_蘓��aͣԓx����J�n7���VVǒ7".z�����J��d(�K�]=ױ�����}��VY���1���ʝO���Ŝ=5<��)E�����(�$�Z� FK�qDL������x[�0��;ޡ�L�y��	�����:/:y�-��7Hqg|�4�G�=(�n���y4e��2Q�4�� �M������g���rΣ��1=�2�oH���Aa�5X����C;�^�����=�#����7"��|��j|���EqeB<��N��Np�������^�`��a���7 =������NmW�J��|zj��^Gtc/�]/��\@����F��IiO�$R6=��m9Iś�-sw���ET��ڈ��&���ٷ飿��m���8|ǟѥ���ןG��f�� u�;�&�J��O���������c_�K~c�g~Cհ�'5�i���2���h�O`��!/jG@�$w�J�o�6��%���T���1`�e�  �� ����?h6+��3(X�l����F!h	�?J�!)�X�Ѯ�+x���($��zp�L_��w��ҶVp:>̞�����ޕ�4+x���K~�v\9�>�}�@R}�=��H<&����#V�W�e�':Ԉ<�g�wme�W�:+k�����=�E��D�j���݄�KnE@ܜ�Ȥ�A_�{�r��!S�7~K�
7��7 ���wQy��Pd����S~�,t!�79��q��苯I�8�`&�h��k����د��(ý�@��j��V�<)�5�S�`0�pI>�am��<��Au����� ��7�ɖ�~�L�I4�ě ��(��l�= o�t
S�� ��1X((��ȯ��;�^%�u,gy7i>jb�M6ʼ�ܭ�E����p4�$b�X�L���y�b+<6QD(�q�d�/��,Q�d����#����G�0�����l�ܱ����\����
I�4���/��ȃH���҅
6$-U�	�H��J·/xx������d�{ǟ7�I��_G��� $-�5u��l�1�xP� �^���́c%�4���=>F�h�'�Al����+.������y�M�����ک����;�������$k�"�>�� Qe�!�7'<�s����q�^ן�<e�|��������T�Ϥ����|l�p'%o9�j���ωXJ���"�JڣI��I�K�r�J�md�f"R�v@�]A�8�3�H��'�[X6D�d<h�eX�����.��&����{�58~�F�4� ��͡��b:�^:~ٱ�oF᧓hn����*nl��/�_f������Z��
Q\��p�:��%�
CCFw��M��]Z�ff~/�TZ�u���M"����i�J���|@��B	��&3���C}�7�������,�����0��f�����������ݞl�u�S�B�C��9:�@��ۤ5�&xNE�;]��E���u��n���t6�D���"I�L��!1�A�o�rؼl�(kiLam@�|��f>D����,~S��i��v�t(#�CF�
� &�mS�'19�p��g@%W�EZ}�Åt*�e���oa?J���
�6G�m���X3�v?�:��zY����h��_�̽��y��i"j�FA���o�\��㚋Z=c�A��v�(!�����)��P㶐z��:���	dkk-m��E�������ۗ޷�zX�	��T6p?��g�gcQ6�Q#�*f�nr1�$$"�A|[h��.XJ�x���ģ�a�4��e-�-�ф�F��:���R���`�B�'",�o��v3 ����� q)�c�$�42�՞������
!�=J�M����Ս�)zw b�o�<��sIiP�rJ  ,8��)�-Tq����t߈�xb;�+�5'��ie�7�{A9�P��3U(�fX�����\���έ���_�s��lFК�Kj
� �J�q�!�)0�����8���
'q�t�kx1A�g7��]��ȩ�u]/Vsg5�c2�G9� �Q��Y��_0���f-D��Y{ޢ�#������i/��X�[��@-�w��[����h��m���W꽹mC�1�LMe�p���������FLo��X�9�$r��Él�o��Q2gH:]
��~/��MyV7�z��lZA�p��1o6!@��=�yD�-}�h��tSdi�����)m����I$��!Ҏ����s�4B���fǄ8�Gb�؛�FSC)DhC��8��t]n�`�+Q�7��E`O�4f��	A�iec�_>��;=��/o{4��È��TK����<�$�)j�>Io~s	��e�a`�'RS�6����Q��vB����I ��j|��vY�����vb~�g<�b�J]�L�'o����+?�^�*�o�=�8��%A��y����CZ��M0��Y?p��B=�ү��5���?4�����֯5
�{|���s�n���X��:���7��v�-����#H`*4%���o�6u<��2����W�~h�D�:���Tv�}�=8�a, 6���}!���~1�/$<.�o|� �Xw崳�;��H.g�Z0�mg���&�eB�J�OF��Vl�bE��r��4'�Gi�V�47K�*��g~�"S�d!t�y���َ�LB��92��Kz�a ��(�)���E�`Iɟր����nQ]<�]q�"x����=rcd�����S�X��^S�Áq5ڭ�H�q.�>g���}@�BY�^;��G.�1F��"y3�51sH�h���a�:K����穃����E0�<
��j�	9ʑ�M5p,�}ۊ2v	��0�K@�e���UR̆��q?��`��ׂV�4Z\���.�-�f>1#��b�<��z(M[E�q�+�ӣ�5���f��8@Ed����z��6���֚}�!n	w)�Q\�\J��]��1�"�]t��E��
�{�
�N�d̀�'��Uϸ���5��27�p�CQ�� �	�v#ԧ/��� ���iJi���C"yf�ق��<8/�K9>P�u�S0�I"�A�=o�9�R&�DF��������y�V�����e~Qa�>����"�����?��Y��_�&c*e-8+�@`~�����)i$c��T�_�+�R�p������T�`96���L	V��Xޤ���.~ɼ(L#I�	/9_�g�^�>\�k�����M:�*���U<��dd�k!p���FGل	~'i�-���9P!�E���Z3�.T��c���eFS9S���s&w�c��\
("R2�{�؆{;�i��9
U=J��(�Rf&p��p@�oY���z}�fWi{���m�	(����%�tV^?�G�uCtR�*�5�����KA�vb1Ǽ���H�%g2o���=��WM��p@cG7Z�9��Ϡ���Q��=
+m�����7i���Y`q�R>���t_�cҐIx�X�<�ˋ퀂�qq��E�$]�a��l�$�6o���Z}!�J k	���.�҂s��&͋vo�qjN�{�`?Y�w>�V��Лtv :ܸ	��+S��]KR����`�)u?}��{���E1";^�y6���m^��f�N�ͅ�����^���'�3�I� ��OaX�U���
���%��r+�A�n;� � @6yC����$|��zQ���>#Dp��[i�sh��s2
����k��BM`�= ��^H5���)���>.y�R��@sQ?��x��Q������� �ʋN��LLN�����Z&u̞�U9��1XQ-�"�
�B�l[CѮ��'Eɇ��a�H���k'$��y��a�z�ߥ\@dҪy�D���m.kł	� �q�I)c�?o��E���k���������Z�a!�O[�M�A2�8��g*�L�ԗ34@��,�@t��@��[�k�qȶBf*\o�	}���^7:��J;�I ��oPAY�+Ek%Qq��kx��"`k� �M	@�l��E��v�磘�~ae""7OU�/� �P_��6������D4@n�jp�RS���w����v���u�]���#��8�#Q׳�D|�tȴA�S�CQ����|��~e���f��f5قg~(uvx�C<��j�]���h����h��bb����䃕�4;��O.�{S�͗]�F�U;��R����[���]����L�4�CE�нOD�ѩ�A3e��"Q�H%_x�P��(���M�(<D�D��������; �i�%���k�$��/�$��K�r��̈́���O��skb��������nDIQ�{�L�j��`v<�Xs�sM�o��LUCX�g�8�l�F"�Lu���i/�V����d�nqc v��}����[����vfr����r��:�����J5�+��6��A��$����kLd�ّb���jTw�D����!��2N젇�����O�m֣�o�(�-��/B���ښ]��2�I%h~�p �����x�7vm�1��#�lq�������4=N��h���-��[�FgF%�3U�C�[�PG��w<�EZ�7\�m�x����Qr����H�O�5s�)���~9��F����!'�,�y� |_��[9�\����FYK��od-h.1"����RK?:E�ȸK�	�U�[���?=`FR-��םV~I�W�a��$Ԕ�$꾆T�T�/�4dXE�|���s9c��k`��X����G�M����q	L7;��򯸐��E%njj���:�����mXX���7Ւ���Cg�D�(��ƬzFSF3���<�x^[��P`��ؽb#��ɻ��q��������.I�c�P;|�F���D���-M��;޼�8�ŝ�u�9���*e�S��[҄��E޵^�3`��f��72�F��l�I�Y�4�$��>�'���Q�߉�OB�X��^�t�������8��k�.�uz��~�A�"�t��ꬍ������j���@�±����$�N��VӢ5�&@�LM��'�������0:s�?;�D���,���\���dpY*_҇�7��4a����Z�-O�H|��X,�Eٳ����)�<��ֻ���u�t���ɬ8�s
��Y��9�ǃ������ �Q.��4-H�I��N�C����)��nI?X�(�쐔�Gn���2,˩��⹷�Ӝ�D=6���1�x?�.�ՙ��kE��bο���ef,��(���:�ص�N&!��Z��T��^���c��.pw�4���g�|���D*���&�n�*���b�,�^Es�	r�@'Yįsl����Q���"��r"٫~�m`9����WcW���w����I��r�����Sd��$�U��E�rƲܾ�j��ɇL��'W��TX�>���ڏ�	rԶe\Xe(�:¤T�A����V�,�<F����S@O}ئ��n����i HZ�
(��fb���=5,:��t4�bEڊ|F�a�����۞\�}4
<���JR����sч+U���7Z%W��$Vcg��C*k�>��2^��
VMP&��&��d�݉]�ۇ�a����3�O��y����v�����٭K��&��
��,��=ٝv���V�Z߁�I��P@�h~�_�$_~����{Ϙ��Ś��L�9d�d�l��$��_ol���k�D���|��BOF��O�y�,�rzF��I��d�253�&z�hG4����Ț��(���4 �Â����:I�Δ?y�h�3q⸥?[�0aݲs����mj���!%��Q�R��
��O�l����VN����T��5>1�G�P����:����|l0!�P)-�,*��.d�$J������F̧�7,pw0�$�����JȪ}��������׏yW�����z�	^0o�+QV����*%�Y�̦�Z�o>��DwJ҄����L�<)ތM_f��$"Y����J<w���f)򵫭�$$�"��3_1���8i0���hBs!�F�����z���<�lR3��U�o��v�����e����>/K@��/���	�����!���9�BP���I����x=j}db�f,�g�&"��[��)"r��/(���&`W=�u������b �����*l��Gm��J�/q�=�綹����4�4���ǅ�\�S�k��r��a~Y)�I���"�9��ijP�t�'E��H ���(ѳ�g!�CW��5�}�	�����h��f�آ]�/;��H��.�M_���6�sv��j���;nU�y~L���_W��ﴈ^��^���Ge�J����mn�y1��� EN�Vq��Z'w ���r��JZB�����Q���	��l�ykZ]�E���V���7ɝ?�D�iIi�󜳘Bq5�ΨA��q��;|\�H�\��9ĭS8]�}���"^4�@�^��u$J�"�<��A&PfD��X�aI�~%FӮ�oZڞ .���B��q~sv� K5���4�O�'mk�X�:^�z�պ{G�.�����e�e��MV��&����q��\o����EA�%���g�%c� ������ �y0�N���^���v��)�]!#K3R$��J���x��*S3�+��ɪ�JifpZ8��)�,�\�O��`�1)�����s�}L^?���QE�Rs����p���t�#]��	��w{WC���xH�S8�$�ϝ_SZ%�Y��#�'��@����txeh�kج�)� �P�#�%���[m��j+ �;�(��)*���8>;���=��P�^Q6	�����S������u�|��]�(RE��5� �����g;��!�Z]��I(U^�@�䭸*�,iOU��(g�K�Ez��M�48�R��euif'+z,l}J���@U����Ύw
��XV�9<ܗ��B�����'���f=��-����¹�en%��^ɻu���:�,�2ɒ��\��"�t��CG@��զ�|_�:}Ү���@�q���F`�16)��vSQܶ�.���s�����Y�e:��X:\��H �}�J4�W\�6n����ß|��Qʟt����X!V�Ja�� wZ�������m`�#�	����
�8����Gbh��(�O�q
��w
G<���+>Of�(���m�F��j�#��[nN%�sls��x�s
�P�n�Ր��W-.T��Z ��Q,-����fd%��]-M$[��!��b�Ol��K���{@�nY?�Ė��&nojӀ��;l}�(�ݫ6dV��8Y�\p���)�_�����E��EK���S��A?l18-�C�\�e�lx�I�i������.���C�5K��Af�/�د�%�Nb��c
�9��	QWP�C��*��bk���E.�X}�Ҧ4d�jQ*��$����+����YkWi7�7h��^�%���5_$�u�T�'�}~�ޘUu��Tۧ$��S�FEHȃi�ֱ!���������
�6�9��ަ;�.쐈�~ہ����q'b�: �!)���̑�A�D�p}��~�j��@���:�mb��\÷��h�����4��L4O90m&��pn�F�C��<\�ʳ����7=kbC/����vf�(a��kë��K�-,�)��G@�r����2���ӫK�ǑM+7Z�ڠ
���q��2�)�ɵ��4��f�@��1�w1'����+�߁4��-e/-����VXb(t����BX��8&�=Y��a��k�=�ң�W��*2zjQ�~1�HI׮�6a_��Jc����H D@������G�cղ�H?ֶ�ə�%��]{����1��lO����˚���i`���z��s'�Bm�w��j3lEF� ݋�`��8��5�m�&�Z.����]Z��c�W(38��<���C�*��Q�r�V`c]`*�܈���셲Mpy��}��L�%=�STp�#2͈-qţ0�Sl(���_J�An�ow}��f���[�{P�xd�eb>?vn��&�z\ ��m�������j�"�ɘ@H�sg��&L@
����@����'սVl�����\ZW��5MO�����b4� Nĸ�/��C[S6ii�N�v]�䍿����A����o�42�*���g=�3\�k�C���{�`EF|LE�L�7�����qH����PT��ޗϻ�!�������;gl�/�����m�k�.UV�S5�H��.w#d�P�O�}��S������-
�G��`�G���>܌gV9o��@#�^sRg�M)jlNf}jr=���f�-�1��x!�N�c#��Q�6�H9�|�6�� vov��m�c��o�L��ȯH�{�z��b:S?591<#g����ٍ��^9ݵsb�����)�<|�qO�����Z8v���m��v�qZw߃5���P��v+�T��1e4��he�f dC�šWq�fD.veK��Lv�[S�/R���
�'YDw���M	�����5�uN�ݩ�V�ʮ��r�0l9���[�m7�\y)�\��=_+Oʽ��+�,�(�l |o'�:��?���B�ɯ����#f�Q`��.RЦP`P5hE72�<ƻHB�|C�G���}ߧ�b�OG�ǧ�lpv`09���~U�0Z��#J)⃭ɥ=-wHU1k��k�e�Ē\BѼe<���]N"�^p�s���*���gH\�4��QA�\�3Aj'z�>��>�.um{��������箼����2�'�N |c�ԡSl��2�6������>���{�u��3A�̡�9��������:�P�6��Y~Jɑ$KV�	���_��bDd9�C(�>�6��4�6~E&e-Yt��A[{�wb|�7���ģD
^�eHH�w��ɕ��0Qy�@C	�3I�����6g�-��_���a������8:��ϣ]������R"������it�>)��3�{#-�e|�J�w���a,�K�=oӰ9W�7��Z�=@�K?�
��+����z������]�����.����-��K�H�i���mAh�+�-wɟ)�C�xU���030��d)[����/���u���
������ʹs>��.})&�⦾eFa�lٵ]$J�֛Κ9
�s���q��[�QmdCI��`K����=/#�dW�CE��f�5A�����g��y'=oEx�CǷϒ��yG�g����N8�SD�0�J��0O�ʼ�<�z|�lfR��6`:��2Ȼ72��'��X�xC�o�<š �K+p��\;�����t�1/�	f�]���KN�"��HE�5���b�{-Wh�Tҍ[�0�z�Erx��!0��Z���SS-�HU����m�2L�LHw��59��P��5��4�ܶQq_�گ�W��b�Na�\�@sdɴ��^��e���'��\[Y͔�Ø�N���2
��@
F�l<�"(��q>DM�49z����s��}:=f�b��ŉ"�y��sf&�t9�6꿌���Z�C!`o�[�.+��-�o�ZJa�x�"�a}�n_�2�}'�P��</�V�70�]�u��*j����9֜$X���qsE$�|6A_"i.��{J*>o������6��m���/�Cp2��,���(��:̶=Ȯr��ìf;�`<��]���[O�DS���K+B��~�il��ԡ�وolB�y��5=�~?�Ӷ"������y�����'i�0d��R�5�q�Ơ5+j��" A��=�P�hY�WTS��:#��ru�Z�����>������s�'%&��+�B1��@e��:���	�B��O6��0�m#���@:�|n�R�ɳf��^N��K�d[JG ���mQ!+N4�%�;9�����b}1�I���Y�=�\���P��SU&���m�;.I0�y���Ykg��^�(�&�w@5;~�w�	�=eW���^e�v&4�o&3��rkg��:�h���"J+�6?�$'�����P���djh��'�r��<�}��z��K��<�����#��M�/�g��9��	��V/A�؅�J��M|(������o5��$����(!�|�[l�H�tN�V)E�׌�n�QPߑ�ya���#}�§�J��H�y݇>�Fe���V����m�|��BUڸc�:�TU'�2��ǉt%�>{"��ekY��,a-���)��ג�@G�µ�hH�Kt;���mo�1G�Sl �@%z�0_z|d�]�D�x6�@��Ĺ��V���󭱻a�D�x#/+�,�iǎ�� �eTl���/f�$�0���B����\�������
-�q;3�~�d:��q[&@���KK��[R52[+��&bn��&�t�����a���΁�ad�o��q�-�y����y�)�Ky2$3B��!L��7�!�odO� 8�Y��&�'�V))�6Y�����H{Ӡ��eq��df�A[u*;dߪ�h]��5(!S�c0�)6�?�ש��!<����3�2�3��@û��н?���W���`R���.���:B(��_���Gb>>�K�;���~.��J�j�`�9�dwS�U��f1�,G�!B�.����.�܅|�����Z��]���ANiU90�j>]��n��z!�������X'��w
�/����0�w��*�C)���Qv�=�j���,����ˎ*R���*��H��_D`����Die�[3P9��2:�|�o������:w$�8�2�M�z�:=�
rv�S�Z�?G\GX�W���NM����4C���rm:�n�\�t�V�Әq��8O�؞:��(͘���'A��Hi[�`�yP��0��:������3g�Db��rFq������_����ਈ��F�}������{���{XQ����J~���3��K��ū���>I�P�|Ih*:(��KL�Rg���^���i4� t�ȕa���A*����0�Ce��L�W�g~,�����1"eA3���HX<�u����-0W���Z���}+�B'߇P��(��%G`�q�;�C���i�����!��á�ˈ��=8�k�v0�����wv�Io--^�^��=)]x��^'�`�h~w�;4�M�`?5� מ@-v¨OU�[fX8`՘ݔ���ʎ~2f���K\k�*,��T��j�H�������j�Eh�J���ua�Q�db��	&;yC�dy/���{�� FV�Rzf��=I����}U�ߍ���/AJ<�+�%���]Xj�n���%���F!m:����f�H6�@��r�>Bɝ��rl'��=�s��_�|����� k����;v�^�d��fߪř&�,�>{�V���}�	�7����n����L_U���k�DS�b>6�	���n�R�t��˙��=)K�AP����m����x�K�v"��|���J'-�h�6�50�Hz�q}\wK\j�d��	2&����!�E�̅6 ,۸�6�˽��z�YI���c~� *��Jj��r�ӧ�DP#���MY�֑6޷0C-O��J{�N����إ�w� ��QX&��`7i�}�{�~}9ϒ��ż�z����� )|�q��y��9��&�2�/����en���Qn�D��$���z	P�K�c$���z}5�EQ��C�&O;{_A]�f�,�\�����$����ų�Ë�w�;)�]��`:խyPCI��O7��f�9sCJ6���4� ���i�����X��<s��P�cE�P��@]�\
��U��Y���p��fxk$7�i8����3�����B�E��JQH�.��U�t����0d/�'ﾏ������������.u� � X���rI��.��FbW��kr�o�'[��Z�̮d�مŉIy?
N�*9D,��6	T�J3'����	Bh@/|����Up���t!�C��!�{��v�߄GdkL���96�E,�z'"��B%z[�j�{-pXp�N@7�B��Y�J����p�^�qZ���D�ҕb{��d��@ S�xG�k޵�j}��eI5Aկ?�p���,Kg<%�vlRq��"VQԞs�d+�q���7�m�ꑻ{��5����9���.7J��'�#47na���6��_5� ��԰+�OA�߱��O+���ˍ��\���1�����.u=H����`A|�����;�[���ρ'z)�?����P�dFi����@������Uζ��o���|d �^�������m["�"�_��u,x�έsr3�(� ��D��8$�i�4�֛�|#10�T���U������t�<W����(��V#���c��PO�M.��)Y���
�Kz���Q�#/�6�$�S9-ȝP�R��J%fL���V��[�ڑ��� ����K�9L���:�զ0��a�Z�Ik���Qb;��q�ٞ�:}�!:Y�R>}���L	�|E�ؙ�����Pl�\����@5;V�� h~wcC����>���h�V�)�`5�=ۯɦ�p M[����|W�k�F�
�-{^���V�����;N|�a���#�/�
fQ�L�Zi���=�Co����oǎT^����%~.ePT4��${N�R<�B��!�GX�X︋
�#��ab� ��$saÃLS�9 SP��">ughm�^�>5�{�%���ԎHZ�e�ʋ�%Τ'x7RAU�i��1��D��� ���2���rCƞHh'(�QB(��x�{^O��(6������|��Wn���#�[vNj
u��W;��v��<YqAt����na�_�*�&��&���1���^��?�Ƿ�թF�Y��(������vM��$��?]�:�6uj؂���y��v۠<F8畍v����v�aJ�]�(�S�W4~')�Ex��U�R`1�����J�e�x������NOfؓ1H��O�����"��a�;�B����|z?>Z6�3����O��1~����]F�]�rڤ9b���nR�l���'���+�^0\�N����(��;�`D<��"`�p3��P=XO�P6��l
��AK��`�ag�f�O�6�\`��A��.��Ӭ�j�߾�1�.�	~�B!�n 0����g�`���]l،u������R5HF%g�7N��  )sm�{�����oO�cOw�r�R�}
#�)U愌����Ŧ'�5Zd
5t�Jw��N��&�����>.wHt�w�hE��!�~���e3W�VxiQQ
Ff*-2OȧB�2ߤ�"���yr���������<ƪk�zN	��)u��#�Ҵ���4���Jca��e�Wdi.����4'�x�H�&a�I1q����g��X䭸l���N����@�)��*�~?����n�~�ث7�(ú��[��E�:1cg����"+ۅ��JB����H��9G�i�����v�k��ݤM��~ґJWPE�o/H�oDO��!���BW�)�P�tѯ&q��4		Ǧ�MV5�� ��v���(��8�G���ɢ�����l{0�E�v4P�ܛ�\P.ְ�_=l`}b����Ms�&>���>&��o���+�1V�g,�-�	��+"����~���9Ey*����Oh��Ru��;K�RA��<Jy$�3+E�YR��v�?K�p�Di���d���G)���Vm ��Kr�8䘍��hN�R|. ��@H^���x `t	�AH��"\+�vFtdh�c����b-�-�����8���z[;��p*}��\��-~3��r��
|�';(6ek% S��X.���ig����GA�(
�������j�zX=���f�k������-��٬�ay��Lx9jvj����)U�x2Hj��H���[����!q��6������2J�`|C�S�ij��ƌT�����4h����0����hS���8�^*��.c1(<��&��w�&� n&��i8�ԒK������~-�]MnN�L`���̈́�ߙ2���ĝ�9l	�y�~����[�9�}rG�3���r�~��8/�Ď���q�'�,����Qzôj:[��qy�O�C��w00��bG�#r9/��3����u��i]7í��Ф���=��[�^���,j�uaoC�*g��{�ERn@g��QcV���\�Y���H16��o3Fу9sf�&�($�w�m[�x�Kx�I7�K�������t^��,-]�*��(6�F'4a��0b�>}����͢ū�����
?�q+wY6I�qw�Z��Ӣ<�~o�r
x> ���>����<v�i�-8;�p͙��x��(JQ+dwH�IY=�~�d� g�m�u�J�AF�P���bR����i�sGј�ݜ}�pL�Px���N�8G�����Z#!����a�h��q�ݳ��@�����$�[|�?�u�-x���F���={��'؃�*�x��Ϳ�ض�e��&x�8��x$͐�.ղ`��E���~��$� 釢W1�Bh���}��)�0^ki��r��iuH�l_L�#��s���flh�8)cr�l��`�5Ůzh���r�9�	�	��	�%^���W�a$ӯ��,̙%���V��:�'ҝn�F�#��c����?���� �W<��M�:�:~}{~�������9,�NT��A��G��p�jm��!r�״����M��aS/���u��u���� ���8��k���O<j9�H�B�������>��:F�/�Q6Y���u
�[Ox�w8]m���9d`'����� �B�S�]�2k��=�z�9ӛ��y��eLmT�gd�f� �_(�,.�M�6a��|�w�·�S�^�Õ�� tot�����5=f SJe���������X�#�4��v�ɰG����kU�u_�k�a���2ä.˧"��cd;.>�0�3Y�O�Zk���vO��"����/�p}�<�L��J���q��h8�#���b�!��CT��_]�&]�^���k}Ϳ�]�)}�d�_K"��3o	������w�������3��j]ހF��J�z� �r�3�Y���
��(�U6XrZ�o�*Y���Ĵ��"��O������Qt.�ϴ���7R�dݨpa��ó`G�a��,j��_�d�)�{�4�V���'/�/�κ��n�p�����ڵ��G"w;�#�����+�,�3�އ,��3ԘF�D�l18�d���TY�<!4�O�k�]���A���*��/��?����H6��bߚ�� pZ7U�|4,gk�$-��@�d�9��=��ۖ�}�H�W��__9���Jc�����'Tޗ�]U�Ȥ�����!� ��'�>���l��%1
��'Gq�V�� �Ю�ix�'��������,�w�,iE_/�ݜگ��'�8����!e�c˘��^������<��-<�|���ĥ)�A]�?$��C�ij�*g�Ja$�,����/�G�G��̗�-.,R��zk�=V[�h��Of�暅���V��:��'R���v�f�]B��2�,	�֐��8>�oGx��B��l��2����=�6M�^r�ͅT>�g���Izp%�e�앂���}�4���W(��ލ@8�{��M����6�F'�}1R��ol��~��߈�eC�q���_��g���?L�:���-��Q�t��J�8�f7
e�D�j�@+���0�`�U'
�9¦,f�KG�Ke@�R����+�R�j�b��T�Q�})NLcl�5W>�����*�p2����)�S��M0(�#�0X�w+%)�O�ރ�`~��h�l��9&yn�g�/��m���$�
��\A�|�5��0I����IU��wɸ<����P���@4��q"�����˰��4����.�\�m�"�v��U�18��#�хQã:�0Nd5�����(�$���'��B����_��l����΍�t~ٸ�"%�N���oUC�t-L	�c�w�y,S}��^�%�(n;c���XC #$/::�"�����,�?���¸q&I�$�Tw�ٹ����@_H�J�u�RbTS��˅&U@k���zTg��{!�@�L���$l�i�N�þIa�Cj��/����	�D'ͪt3 3�=�oz�AȖ��>�Q�Bljn�џC�x����^Hu±WI�,s�?Yu9
P���#���,���}ǟw9����5J�8��Y�V�-����.��8���.㈒��N��o;}�
�����br��<K��ߙl��0���V������������M���� ��
���h��	{ހW]{�0�%���ά��{Fӏy���	d$\���Ek��#Cs���@ؗ�R�)�L)�r��e����k|��+�=������4[?k)S�q7!�R��
� �u��~���ѣ��2�2O���n��<u�T�s�zb?S��54�	QH���Z_��O{k����À
+��@�I(nt�s�b��ŴsIuz��!BP��w�}K5�
������*�U�����rlG� 7�bõ�߾r����6��B��:$�bۉ@9��G!y:�>+�,�v?>uRi���#��r^zܜ�����[#����4�������pBg�ckƐ�o�+��uc��l�C�z�q{��(*t��j���ucV!_h��p���K<IINg�\|��L�ݬ�f����S�K.�����1�T���'�&�?Z��N������0g����*�����+8�9G9��pFn":��ڷ�(QR��+ٴ�`�E��'ǫt��Y���zx��E���jn���±R�ۗ���DI,gf�M�M�R�M�xa�UV��4�e|����|�eX��Q�+����.�څӒ��C�q@Pèp��#�x��O���t$	���;��z�BicQ�:ء�y�_���[��JKDt�s����7��\iu���n��0�u-��L<To�Ç�lH���b�
��7x�;�_��F;��&��L�E�<g��Zb�uU]!���blȊ�yùNl�%�uZR�-����߳��ܧ*H��p����CCS/�yJ*?��� ʣ��c�Eex]"��tfǎˈ��5�lJg}�}?Ӓ����s)TbC�B����ژ=��T���nCp}�пY��%:�9����u]��(�]f�x�J���Cs�$�`˨�\�`�����dF'�W�X����k���ZF.͠�J9�w�YԄ�����F�9Q\RT�jlm\�:�@[R��\���I��ԍ/�H��}曤A�|3�H�_.�y��N��W@�Yx�`�S�d�n�:/�B N�ɈO���N�N��9u"1��d����'��R	θ��#�����c�pr��8b����k)#M:J�&���`H�E�0eNT�JO�h$��8l%Cd[U�J��
e�+�Pɺ����2��?�"J �ޥ�1���l���B ��A�/�8�P�DYHf��H8��� �H�{���!WxW~��J���+D�����fL��2ɫ,B�bU(�����Z�d��g<���r�G�2�h!C��Z���f�p��=�O��vȸ�7��*��ƤT ٪%CD���
��yl��t����>d���t�+��A�*�I���a�xI���[�}�R�̂Oq[9f�}������_�ns��S~E���Q��~�h�V�9eg���"����Q���X�XЁYhrm��xk����(6��bn�@~TN%�"T�%������^�*?ӄ�'_�-����2�`! �=c�\��Y�p�6��������/�b<C�I���c2I;hYb�[d�qG4�wqt��l�'�V��^t=���OG9���k�pOPkfgQ�>0��<-(��tg�C��zPlܰt�֠����|�X1���(l��0���n�v��A�(7��В,�L��p��5��ͥ	��-<7z�Pw@�ь�ԥ���@��[��Ӕ/(iG�������8L~ժ�&w��@����?�m��w�'��뫱t�F��^�1�:���C\ry�<��R��/>wܓ	� ��:Ζ��\lk���&b�?�Q]b���J�XI�l�DK���{��ޙ�(wu]�$~��>4K�>Ѭ��r3�~<�_rꨕ�����_=T�7Q�N�I�B��F%�P/˅X�N��n{��~�,C�Y).�R]��ܿQ�� �6��>�ڜ�+���\'L�Fǃ�`�v<��X-$[y8BL��%A�c�'5`�[i��ņ�A�i'Ig�.�m"���&���p�F԰�D�����VaH4����ٯ��<��MAw�8p�?ۈx'<��k���#��d�+<�C�����BT�7৏��3T�3ěskMi�9e���!ȏ��;޼՝���ۦo���fc��xyt�Ս���L򵚏ȃ�"F�Z@���P|�	Y���b-���̸(�㼁�j�����@��.�A-JI�R����m-�ż�|�0����sJ�f,�����kq`�q퐰N}�T����7�Q|��$��\`h�T�� d�q�B7��nf�8�$������0Ld�C<�g���72��Bx�vS�W�����>CWLZ�H��7�Ԯmr�>�ׇ�Lѽ��M,#�ۘ���F�V��	�i?��ٓ�ĎK��
O>Z���W��jSk��� ؃ �"C��F��ɍ�׵�S�J�'O�8�޴��韑��̯��{�2���-q9�QLXb-�ׄ�R�U�T0���P>6�J8q>3���R;ɉ��ޗ%�c�M�,�tk��?l/����uP���=��zynߣ��N�&�</QB������!ԝB}� 8�U|0[Ommr+���B)4��)��������q��ò���S�Z8��g*&�R�ZJ������~��P����FR��2YBL�2�9��g'�@��H���h�A����zl��/��:��5؝�}C��	P��z�!��
������٪���s1R�ԃҨ�	��=e���B����k�9�b��h�6�6���9���`z��L��z�8�y���F�p�� �C�_���I��G֝�k4��d,LRL
;tDRB	Ns��^�U��h&�*�-pЯ��?���4g-��[v�ZU��)s��	�H���gN��p�Ԥ�G��x��px^��w$e���r�fr�Pa�
�d	��wwk�8)ӅƝ]9�0�>��[���x����T����튖P����H-�Ki��,}e�"�^03$o��J�����w�R��ƹ)9�`1��TO� n|`3��*cv1II��v�L�Ѣ�v�D�{���P�����!�5�3��>���j�n^,a�v�0��}�� Y������D��\E,-��Ȏ#k1hY�xy��ew$qk+��kX#-�$���E;ʪ���l"kc�A�/P��۵�������P��W�G*D��]V�h{����F"�Λ6�;̨8å/E����c7�����C@�N-eӶ��@ẏb~�&��	��?XM�ce!\ JyĲ�V��d}2�W�ML��8o�r͹�4:uY͵�H5\�s���_cx����]���'և�8�`�5���� ~��vO/�o�Jz�a�v�*�u#��q����˵{Pxܡ�j +�W君%5A�ge�)z9���@�Թ�wX��gL*c�v��΍�(�|_H��S��<U_`Iqε~�'.����m��r܂�r��(^B�{�m[���|�u��]�b�VX��Q��1S����C��K��[�ٱ�-���t�/�R��1�Xk�s_�9��#�QӰ�����4�*�4��ͻD��(8�%�b�6;y3*�ܣ������ƽk�G-����`[�� k��"M�|N���U Y����(��.Z�6=�"���;��Փ:x���T��du+��9m�t���%ʣ}n0dE<�ye��
�����'��vN����/ (=4�L"łv>���@Ã{����)bz�+�:&jS��cGk�|%M����qbU�{ά�Կ��"v�!�m���Z�����/�`]b���鴤��3ތ��)4l,�䅆mƦ��m?P���(�wX�G�|6�t?�t�{f� ����[�b�8����/�c������'X]%Q@^9w���*DUE5p�{�d�=�Q@1�o�5�Ed$"7�����L�����^P1��r#�T1OZ�a4�\s(�u=ŉy���cZ�P�m���� ��������IџH��&Uw��I���K^tefԁ�婨X��C�|S'/���I�	�޶ȹ���U�'��oy	�sc���3h)�͜�>s�X�x�WPuC~��y$�S���	�#<2��'�-TH*ɀ��6��A �јR�SU�:��V�`�ߜKj+���?����&'��s٬����l tb����X����
#<��f�e�4��V���×ܩp��z]�%�'�f�O�y�f��׷p�4X,���e��6�z�>�@+����2��#Ոɍ�f����N��!si
���u7����3���~�}w�&D\�:�3�o,��[��g#F���_Bz��Vʯ.K�#��ꯚdW�ʴ+
*�����һ��sF�3��Z2Q�	;�������-.�A�p<�W�,`<�R>�nV/E���R ��Q����$.i���G'��q���e!SoƽJ%���!є�- �џ�;Y�k��Ә60��c��n}+[���V�^�w�{�[���#+�%�.y#������O�T������ �2�/gb+e&�����>�
������*��g`+�X9�����3��l}�A�Y��:���/j,�*����]��C�t�֓p�Lcm�u��n�����X(�ڷۙ�j�U�(A"/Eb,0P��&����� �c�����>/�$�1�̪7�V�dh'��poHAj���(+]W���w-/�<)�{�B�1�n��<�f�SeC��o�YM�F�\� ���r걾 ����faو�z��emR�W�슌9H O"�Ш )3��9J�+��b��͐�✝�����3|�$��7_=����x���м1����6C�B�P�~W���K����ڜ�D���I�8Q�ɲ�S �.Ђ��me,|$��&�9�6��:���l���u�z�
j�z�"��%&�Vz��X&t_!3�,Sۙ���Mf=d%(SoT[��}Y2�t�i��f���]�ƚ�@�.��?���D��4v~]�rA2j��]�Se�vv=��&������4��_�k���.�̊4StB�
S����񎬈>Л~�[ �Kua���GM�DR3��Xe��'��6�(�׋���cW��1<Z