��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�y�Sy�;��>��&�MA�)Cʌtg���e�8~�����=H�9����.k������U��U�Xe���M�b�(	
'�m��_�S,(
>ɢ&T^5�[Kم~�WA��Mb�c#�<˃#:}��6͕��F��O�j�7���'AF�9��'�ƹrq�9�p�
o�'�w=��v��("�|��ӏ�I�\.�V�����)���cB�չ6�t3sꀚ u?�({��_x�W������!�`�e�H�H���|�-�YY�
ꆞ �Ӟ냨��e���S�kFd�v�e����y�*D���G�>����+�ᩜu�f�x�I���*��/1\1����r�2�*M_�4j�t�'{)ȳ:�A��!���ש��6�D`��Js�[�a�O[�G�O.�����}�9�����E���;I҄0"}̙�������@pi?%D;�4���SەW�L._=,k���1�ꐀ�Y++e�����`9�'� @��a%#�Ɋr��#
g�PT�����x�����O]
��}�c\��1��0�:�� �q
�j���)߫���Z�>�{c'@�n&����)j���\84Q0��������D��0�Ue�w��#�).g���ʺ�^��ܧg^ w��Y[�����x'��l8���W�P+b�I���c����ɳi/l�^�� \ի~%G�PXV�vqBT�Z �5�E�k�y�kyz�T�V�Z��8"*S!n�n:<�q�{�Q�P�[n�t��z"ތk�=N����l�Z'Ί�1賠Lo�"�8iWN�W�P�̄U�G|D�/����{F��̀\`ث�G�I% ʴ�L���Ϋ���Uz���3�	Xӕ'�j7�EŹ"�j���u*q|z���z�x���}��-��ex`P���_м���a�y%Ǩ�#}6�1Uq}�=��Ŧ��,�ԧ�r�����yl�[�T�"9�S܀�5�ڰ�3�`�����￈:������վ'��n�T	�XA�yl�Y�fu8n{�&��v�=�;�m�.ھ�P�\���O_É���w�r,��62��O
���0�I�O�?���ڼ�6ȅ��~����W�Y��S:$tgN+Dtp�.�$��.-�&�{�<�f��U�[�\'���e~Ѡ����j���H�|�z7��QZ�������ʕU�	'Ё�y�[!6�ЪӒ�� nb>h5��tn��Yj�N�l��x�^E���T�e��ڕ�x�,hH���È���T��xjN�v��0��=~�9��#ӧ�0N�X4_n}3��Qjk-��w���� ݶ�S_Ɉ�sG�a^�2 5�J��cxၲG�O�6�R�T��K����$Q�,�����z޼��m�}�Y�z�y��o(O�	��@q�`�Y��%	���/�A�?ɕ�rl�@��3�/845���@o�M������=H����L�#7{�G�?ʫ�Lg|�4��!��=)P,�nk�q��l��T'1���b�d�O�蚈�!W��*:s�lU��l��cI|8k��V�t� ,"����KaC�")��KdJH`w��iM���S@�_ �l�	r͠��Gܖ#om(��Sm����0Y��u��J�H,�}�|��{VK��;�NNl]lop��Ԏ
�QI�����gz�	ې�0��-G��o�Տ�R�W Y8�E@�f{/P
7OVwj��>�w���ˢq�=�?O�v��a|��v�����t<@%��g�k�N���aث�hߛ(<��`#�-�ڵ�"�$��}ܧa�~Owfv����t��n<�P�4R0�եI����s�$y��?�P�q�Q�;�uGy�7ٌ��T�u۳�nb�{��D�0��
����XA��ۭL��h��:"�9�)�(�R��N24fL�\?�7�3|��G(��d(��7t`[�c���h凜�Y�"`&/I�
��pq�/<��u���@� �4.��S3�'��>!y���ppؖN\���=��ÿ��J�sK��ń߹�������U��a��DT>q���#ޒ7 �x�����w�G��C�Md�%�u$̑�����n���CDv�机		R��k�,�xw��om��q�DQ�Z�c��r��P}�y`�R}�y�Z]��/�R��6~,D>���6����;fb0��1ҳ�o�? y]5I�$��M|M�^����6���Pf��^G��H?��
�����7���6M\S�"���lY�U�3?d�����+M��a����X-|Cm+�mtL�5�#�͏n����.��'��3�*� 0��%ѐ5���!�==��K��\�Sz#�?���Fgjy�a	{�(Ʌ�u��pO�VU
:���Lu��5�`)8Ǭ�z�(cвU�>�s�c�_�9X��Kl�R&A�ZP�o�4�5�ܡ��K����=��1o�i��@�� `������0c$�n��<ϔ�΃���&yne"�w���J�%y��iἾN�O襉_J=;:D�(6�`�b�^��	���ĸ^o��,,U
�M���A	�1�r��]�f��%Wn[��I᥏L��;W+�mP�%z�i�����5&�� ^j���@�OK�H]�0nXm#(v��U�F�ObU�O'�dfO��࿻��0Ǆ���G[�O-8|UtGL+���w��[�q�? ��eфQ��qR߶��l%�vMN�&F$qS��n�]�G[Z��w�>#��v�b��I��C�2"D��G�L�z�_)�f�Jƙr��`��m�;���gVGL	*���	=�� S݁��w1�N�����!�y�vo�8���w=7+��ģ�q�b�11���(n�#Ԁ*^�)ZƔ\�u���!�#�ZF2��ٴ���ax�䙚�ށ���)ya{��PP����WYS����MB�G �'���/��[L��<��
�A�ѷ���6�]lxm�I��ݹ��#
�����?	�D�#�T:7��o�q@���<W�N�eg�C_�](n#vsl����a3�6�[��2�,�.N�[��w���^1��0���|D�����0
`$p���m:���=�`�ܺ���=s]<Q�c��ВU��՜�;(�r�%����[�����}w5����q��~���ҏ��*�^����2���|"�?Z�R}�o�Ў�֦y�!RQ�^Z�Tϛ[e@�bo�#p}=���e�x�	��\M/�)z(�j�K3#K/[/�2Jl��l4`��T�O�7;��F`J U90y���`��v����o܃�[����N[g�dt)��N����L���
� �Tx_E)���;�̀���:Vd���V�d=�X�%icc.�o6MǍ1As�G�s��0@cig�?t�#x�V�&ܯ�&��:q����� 3��Zv�C79�vK�7��zy��z8�x`Z�0���)!�����"�H-՛�3�Ϡg�Q��q�����Ě	ft��yH�gy3q�Gc\�2/��cۃ����R�<V5���E�F��y����<�~�An�wz!5~~7�gVIny�/�~����T�O�8`Nh��E J.Ӱ� �|�`�\(N���7��"���q��=\�=K�� 	qP������Qq��V��p�Q2��?HBÆrl�W���M�9	&Ng�ɞ��f�vej��{��+�a�i�����֖X�P�e�� �GP��Ǵ�`wf}륚�6,��)�A���SLu��w��ލ.U���\�H����Wڄ����3�=�H.'�֬li"�׉�iތ�~2H�'��_'z�dW|�0��6���#��m�r?�����N����(q?Kd%�#u��`FIu�����0d����OΎL�.�l�ޗW����%��QV6�C� #�@��<u����,υrm¤q=f�O��&���=7�hre����&�QR�(�$!���L �n��@I��o��F!Q�����
�^թ�"�I�w�o7�y��(�+B/�{�ő�Y�N3;��V�MscVϢZ�'�/W�t��0-�,��/e�6����Ȉ�_�<$ ��,���@��v �Q�xy�W{��u�����n�+�7���ox�}�!�;�/Fy���(�_t$v���.���M��eH��xU����W��HRաy��,	[^��E4F�,�χ�z } _g �Ó�3�C<]4[o�(?�7|��+�N�Pn�(�M�G�0�}�~:Ji�!Fu��\3^�)X1�`�6@��u�W���%�|�F�E+�W<-��Qkpܦ�+c����2�i���f  ���³�qkX|��,Kp�IL�l��}_|�8:lp�/3 ���͋��nȽ���ԩlo�ë��>}䅀D�B��61�N�+���c2��P����t$s�C��FY�e[5\,D���K�W��%���n#A�)����.��̰���o��G;,B�-�����v�sod�:�r��>x�1��֞-�#7��S�K>"<'�������B���J�Ҙ3�/����""�-�S�@f�ݩ��Tu;!J�V�	��Eg�g cT��SJzq���\����ʻ��0��4�!�)	|e��E����@���� &�q4� s͑Kj���aM�wN��~Y�L[,�E��i�t%"-R�ֆ��=��B�0�B�ė�jO�:�>�\�࡟�8�l̂�?*����$���ܧyRDi�j���������tЈq�Q'\��r��$�����\��A->uFPհ�ʑ�18œ��y*�p�xXIb�gd���a��U�kM�}R�����܎�������,t'�	��r�63��E���D���
ƍ;/��:��3}c������%K�/����M&�����7|�:���r���F�H��e�Bu'�%�wU��e�����gB� �kZOS��k�����1I�^��Q���(�52��"�iEY����鞍䄵�V_�ACe��4��1������ӯ�b��a��yim���%p���Q�l���d�J�~��_[��_Ѣ���/����������=�`9��!�W�g�1��I\���F��fP�6T�t���k�.��8*�����[�n�5�'aC4����M��$�B���G�m�U�������E�x���r%������ا�/"燜n��� j����bꮆ��#�UA%���.����{�9P��W�ű��:̭/�(��$c�$��9��g��u�
d�@���_UBN��1���2���4V�����I��N!+t9F�kx��� ��r�MD[�\�h��'�h1��wB%DR->̓U�A�ap*��:�^~?�&A�hF.�T�n�!��	Z�J��P1g���z��~<e���"�; ��g	��h����M"<��sK����G����Gt�Fn�T�j���4�iZA�����;���VҤ�P/�)����cn��c:Y"���X���_�K�ꝷ +1�>.�bQ�R������W
�A��r9�\Z�\�Ԛ��p7,x Rm$t5{̿B�qCs�5������~�7Ey\F9|gh�O&YR����gs��r^OlE��ŉ6ײ�K/g_,Q���7x�����G�����8�_g�y����ٯQ�2#2m��(a�r�!�T��Q?~>Et׬��K��`�����GV-����'���:N��"��>��9��Δ�-5[�p���3���2rl��R�>c�Zɣ�����|t��:�o���`��0
������;�Ggq+�r$�&�_~5{%�6��ٸ4�-k�a�0��WP�䤈،]�*Շ��1���+-�FϗY�E��y~�,��g#�����B((�>�-5.�@�U�['$=�R\��k���v61V@��w�>ddw�e�%7���`4��˚)S(	�L��A�;�2a^�{�w|�6�~5A�i$4�"G��Qb������6�h�)����=�S��|y��|evj�}����8�tᚤ�P���S80���"}2��n�fd��ƇvNn�8i�L��~ �gxN8�e�z��OV�|~@s����ZS���9� n��S�%�,��B�>��� �_���G�}V�4g�_���"����k�� �0_���qt�cF���=$�����`(W�y���0�C/���?�:cv�g%�>k����a��OF ������[�#N����vN�mH �	>5�����^��Yq%Eבy��Z�Nc{m�ƞ�����,o��<��G����Ǚ<�)v�Z��u\�P�v��Ԩ�:{�y��&�\e�ߝ`ch�5�D�X����\��#8yV E��-�b��k�=d�Qa��6��6h��	j��N�,ɠO���4��J�3D�z�5B���t,�
}Sh+��IXI+Ե�t-���~���d��y�S���ͭ��L�
R���'��iH�0�^J:.�@����J5Q��Ix<�(z]NN?�Χ��K��Sƈ:1)��_��M}��c덫x��(5�8>fh�D1G��8�>����e�|�H�2�|	؞e@�]0 �}sB���-����U\6�\�۱>���Đ��;{#�.�^d�^��؊�^#�T��� ��+E5�@�W�?
��ͪk4�Oo�հ���˔�mq�R^��0����O���sK����ʉ�K=�-�A'��P���+%	H��4�����D��F}�=���-��G��A_�O��J��N�% >k#.������A�#k��Nߊ6���!��@�<���`�� ���!1��u��;��VC ����)���"
@O82) [d*F	����q�(8����^ A�!��"�n�_~��z��.��]eO�休���.ژ /Lt��W����_�V;�.���u�6�I�>.��'���u��ۣ/v�M�舠�L:��
�� ���4��9�U���QP�ť^>AY��GI*a��RMfS]f�����X�\Yk[�y��
[X�6�'�x�1�=g�)�׈��b�6���i�>�J����АP/V�u/=[�#��n�����E暬��Q �@%��Y9�k3�Ax�*�c'��|(�X�*ۃ��)�L����R��T���ښ'ֵv*��zڽǁ�6f7()�≪s�'����ř��� �Xj�9U��s��Ex��㈹�4��Θ����{�Â�����DF����V���$��3���~��i��&�r�Х�|Ѳ~I�P��;d���Y�A��3T��
��F��b����Id8���t^����%���e�xt,����Pcd�
pc�G+�r����%��<�Eܚ{�n<�!k�]�J�v]��t�a�ʓD�.�NW��an&���%��?�1
�\f� �uC7�`��\�n~��g�`Q)�U��K�K�	lT�҅���S7w���J��,,tπh%���P��p?a�ù�zԈ�gl1Ռu�Ck3}�v�[�H�6��a��L����F�V�l�[�A0�'P���O���6�%9�&�l�4����ui�����z��S����N��!'[�.:����R�26�����Q}yPQ��$j���t�ʄ�Zg���"�_�9R\͍�'���ѽc�uoS��e�hS��y�i*eAFO�w�~pHE$��3���\�y޲蹇��: �J=����6�j��7����A�3��}���6 Å��e�E-��*_�*���+��Lc��5L!��^�s\A�u0�8�Ȗn���q����<�6_Bx�f��Pր/���:0�M2���!���I��(�^�
��\|�J�$��r]{�y�����k��w��8n�D�}q
.�A�'�N�{|�M��E'��e�S��w�t1`�a3��'[E�GJ�8Z�35��i���*��H�R�E3@2H�=���ݮ:af�i��z��Y_���>"I��1DVz5>p�H��L�;塷![p�?3jt�Y�C���p�7"ߍ�STp���L(�]�T�GZ�Ufa~@��e�s�	�~V.��;����A�-g僡�	���0D����S/�f��B�&���h�2��0�f)p�H,�Q��C�0��Ü�6$��g��̉� bA����k��6;r������v,c4�0
jB�rIkvB�8��tVo� `�A�]��6
b������诞����Y��3uB��7�,ȮЍ^�I`W7�^�_����,٠��v�� �������莇�ƗM�ֺl�Ԅ@n�$,xL�|JX�/����dl����`�Z��q�͖��F�ܦ2�n����̂Odn
���f�^$�"��v>	r1��f詖��q��9�2�5�FQIP�E����(a���f�\��tu�:I4���2����^e���D���x�n���� �N7���h6�h~�/�<��(+OH������梧�uYNņ}:�.ο�7���7 �PR��i��f�z���^�Qa%�t3��s%�֗\J��}.��Na�ښ^�5�@�^���K\l@Ã���J�Qv��s�X9��z9��������N���Q�NQ�'�b�f�"8p�)_��'Õ#���%�^�\S�w���N�x�eݝGB����J�P`��i�&�"p��v��_��󡿢fj�elO�i/G霼p��><�Au��<�_�&�h���d��V�]퐸�"R��w�x��"��F)*Z�=�q���ϊ�:�EA5��4��W@�T��l�\�[�F�]�"I�#N*�p���x�M����'�s�`��I���4,\|��l?N8�W|�k7���Y����z@Zl�>�HK�C��ZV!)�m �4���WVeJ�ci����<���Q�O	�X���dep��ؖ*�bW��Ґ/�6�1B�S�I�yS��y�ѯUX͇�P�Q4c"�H
R�VY��ίt��������Ƞ��D:�ȴ8��2�]\>����:�L�E�l
�6�����uQx��(��������k���#��}��L°�2m!�	���7�Ft6oő��1�T[OJ��64�US$��`JV�u3]+η�k���/�\e�����=���(���6��o5�|0&^J!�5�A�`����};��>�䝙�M����&����ŝ�� ���fw�F:��ђ%l�g�X\E�k(�����A���B?n�Î"r���7F�_�L����s�m~�
J'�K䖱�T�P����.6���b N;�\�/K���b�ʏ~S3�D:���T�ch,c#a|��AXH�)��I8��S�n��Rv4 a�h�f�O�5�*�?/�X�_g�*��j�
����4��  ukl��H`�[)��Vx}��1��>_(��\�B�j�}�c�l���������['�k/��N�a�kP��\�j�J����եeF�f�L^E7N�A�^�m9�g�����Wz`�g�����������)?3�����ݰ���b�����m�6M���+_XQq?p+M��p����>��n�&:ɉ�,���,�f�,�['��n���xP�}�]/+�K��{p�ܹ������^�(9?=_x~:��*�;�N�6�/!�#C��/?B�q/�}�M����<)x��*g��h�e�B^2G�)a�����ߛR�;�Zb
Lg���r��B��
p�>�aZ.����[�f�����Ph���W1?(s�|�c6N>o߈��=|����U�� �oP�8?�\R _��漲��<�ӂ#���ը����^*1��x�U��j�x=_���{ױ�7{��FȆ��m��O�h���d����4�'*�)bw� �����L�
Pe6�^�n�������X�(D�゠Ng��Ct�J�ǋ2�f�H�Y6/����p�e�{UTS
�h��ΥZP2��z�' ����T����@v���t�xVjq��Qe�jN�9<5y�7T:��;�%�UQ��6���W����Ʒ�Q��3�H��挕'~\}���U�ia�׬��-w�rin��(�Q�$ztƙ�.��&-H���"��k&O�H>_�{�3A��8�X��Q'���I9��ǃX�L���0���/ ��5�u����.8�KG��i��b�H"*�H�T]_���j
B\i��p?����rQ�؃�w[,��404�N�����h&�4����0e�Z�*4�v.�)���<1��@#���N��� 
�iw�iL�%�ʾ��V�p�&����E��'E9�}<xM.x���fe�P%�B�eD��0�ͻM!���4�EAM7��M�YD���:d���X�p���Q�%�I���@�}nh{��+�fP߸�}����6f����:�]ȹ�39���:D�c3O���H�%�yA�Rz�ݢ��4�O��i��m���?�p�����x�ĕq3���!qZ��%�7P��ah���ؒr�#󨼪-3�2��{���?�SD�� p�'��(ɿ~��S�~�_�ݿf_�#.6��9�#]�?:s��;YҪ�X�p����w��m2e��K�ޖ��*:��+��LC��-��,�$]a��aA+v�
�>V�0��^fp1��`���E�kגVd��[$�F��-Hb���'�/\-�z@�Kh�@�����k�n?H�C�����ZФMA����\�����S�fzj�z��)�`T�qck@���J�ri��̛� ��^1?&{��o[�6�.p�kcA�����0����d�TE��{���f����\ȍ��(}�\�
�0��/�A�lF0,`���y���`�=�({������,��,���`�)��ۆ]�a\�A�i1�{�m���䓋�[�-%��d�������哝*$f�K��)_��"��p��z�ܳ0�9��Yy�n�TIN�!A͌��3�,�̈��+R��fz�AۜS��5A��P���D���q?Tj�Rl�¦"���Ÿ���r_�[N;z� ����Ǯ�*�K�H���F�Ӡ�\��a�Cg�	�>5��'���u1gӷ3���ɔJv��m�'�������[�*}>s<̄�'�fq����M��4�/�\2�*P-��^g�qݎu)D���Ǝ���9p��<S�� �A��b�m��<�t��mqm�"H�ng+*y}�"�I9 �}�?��(S�!��1����߿�<���g��G9��[	�YgF���� ��g���*Q�	�6���!��J~e۶�Cـc��Ļ,&4�i?� ��#Zl�O�4��P(*�`�޿�>�q�J!���a2��H�(�,{�Q�f�fQ�ʋX��%�"���(�
�W���0�+�Y+�{(G51td�V���� _�	��%�����v>4��nA����9B��64���A,�x+PZej�$�5�'��H3��7��Ux��xa�)ԋ�_=]��l=�c�3B�Yr�.��GC�F��N���;q��֘g�l��5�;��.Jⳃ(�2G07�����v�u�{xeM��i'�l0/Tδ�-6uw�Y�-~C	�҃�.�d`�y3q�Ŝ���/�����+���	Ʊٿ��qݞ[��U� �^�Ӛ�< ��X�u(�l<�9�b�H4{m�33S�[GlV,������6��A���>��E~�����m����\Zٻd����Q���n���3t �bƳ^C'D�,l�)������oC����Y���)��|3�{��G��r�`w� 1)ʚơ�W�m��\LA�E���F��V#���6�W���헱=���{=�G\�	ݔƐ�ndw	�^��oYO�{,�4<�������R�	W�� ?�J笰~ű�P˟�N�6��K1�L5Ǣ��E�?4�/�u|[CA/�R�z������a���%h�mU:�Ԣ�&��S�ٗ����ԁ��z��,���2��L�DT�j�V�	f �i�㫺hC]8�Bm�
f4�)�p������գ%����;��!�_�쾩� _E��mlN}O4�_~�-o���zN����l�C�L[1����2��x�͎�c����W�ALwϐ�*�E2�ۄ���� ]ix��M�TYwN��eg��w�n�	Ԝku�AENf	�2�����Wkg-�ԑ��z<�OSt�D��I`u�l�����F�&���r�S�������Ɇ�p���MbX����*4u����d�K���Vv�Hbj^�U����	s�����Æ'���]LS^$'F���n�
��a�<?}JK!%ڣ�.�R�讛�H���� 㢂�h����UY.�3�j�:��gn�W�:��,Z��7�%��?@^]�G(�.Z*��|�`0$�̩/g�����+~�g�+��T1H���R�	(���Z����7_@d��	�}XZX#ȱ�Ǖ$m�iS�$f��!nI�ެ?$ЬU�o��Ǉ�.Q*7 ����o8�N/���c�SR9fe�B���B$͎A$��l/J¨�;$U9*͆��\?y@�+w��ٔ��^!��ӫ���J����`���v�1��&�%��iC(�X�+�:<��@�/<��10��=��H��!M�~j����� �&�R8g�p��`�ɼ��]n:p�����j��V� Sߺ���N�����WS�4�`k��:N��!i ���j��0���� ���i3-�*�l}p����o��Z\=�Ֆ�^��y�7J5c�9f�{�0\�R���3&hE���Z�ͮ��v1��6_�J��\I�5\Y�7G�
Z��H��	_����>�FCmdg(��#��">ɢ��k�:ꈴa���O^��>��j��Pl�1�3�zc ��`a������6o��,��2��̷��T�z���2��9�SoR�>��d��bi���|F?kڥT�YǑ�� ��I��kf�z㛐��ZxU-���!{a����O"�]����o�l���H��b�o���Z0f�G�\��K�P��j�<�(��3Sh��\p�~�?��=&��nF�S���Ӯ�b	��&*��I^Sn�b�]y�ӣ?ic���ө�Q*D�n�ޱ
Y1�	p�t�<]��ȓ��9�;Ѫ�Zk�0�U]��aC�;�u�"O�#�<U�5�֧����s0�)�ɹ����ߧ�g�P���Zt���w�t8$�Sɩ�-���Od��;��p��;�Fc��ќ��,�#]@��(n���Ś�1�=YP��)��ګ��)&�Y���O$yR;X���P�ē��.L�,���BF�e �>a�V�3�H����v���T�)�Zs�*�UiY��qF�5?��E�<�yq������u��P�y�n5���� �{C[��?�N%S�������N����Y7X��=Zl�F������߃��T��`
�d��2���D����O4~5l�I�}%��F����p�����:�v���p)�UI�����8Y(��M`�No������DK�uǶ0r����R(��SoJz�/�'۩��e_��|�Bh�E�2�a�:=_@�X��ý�x�跇�_2z�Pb'�vI^�N[����6lb�k�1ACq��+��yj�a#����	�	���zJ���y��-�)�~jh��R��Z�(۝xj����}��*Ak}���>_��(�^{<Gf�i��T	��^�n���0*կ��?0gQ�Dq��Y���Jb(i�J��i=��di֮H�@�_%�����V�i�යD�]%����Ʌ��K�.���{A��Y�S��Q2k�Q��XpWfi�f����&���޳E��J���9a�Ry�q����էM��K�$w���YjW=��Ie���j�����̸���U�3tE��#U�����^%�&�zN&�&����)oۗ+_���ݙ[�g���܏G0u6g5ܑe���м%���/䱭]���\�p˛�9�5H����(�czW���n�-(�)�fU��E���c�4���a�$��p�ϒ*�)�1���޶BV0���u�p���"-c���i+K�������m��*<h@~�;O�����i T�K��d6I��Ԛ7���i�>i��������h���%�ױ�p>��e����1�A�3"Z���{���q��e�(�{\}4	���i��A��ͦi ^!�wg��2�C��)t�zH�qv3�_ϋ�Ǿ���*��O|�{�.���DI9�'z��	%��@*�	V��%��.R������,�޻��]<%Q8s�dYU���	���ȍ���q��L�1�n�k��������6�u��M�=W������/|��PP���C�'�93d��t�T�)�Y#���������O�n�@u��ǁc�w�R-UZ<�q��ٚ�}=�{9ǠԘ�)�0�S����b�(o��&�;SM�3����;	��ΚVۚ���8-&�������Z�1�e��� ޱ�;.�(E������	:������>� �dz,���xe���0�@Y������2�xf�Q����=��$��-�]��z3�
���~#F⧌����ۮ`23��3��J�����HA&�.��M۸nĤ��{�[�NO�<���gQ~N=aa���
�n�m�W��%�5��iA��0s����L]"��*i"���;����u��WȅK�I�%��>�����'��r���BJ� �4c��@��:Am�ALBL���s���xsU��U�ذX��x�}gxP$3E\Sɤ�� �wi2����-�N\� F�_�oҪ ^6�,`����� A�+�f`�h���k_��"R��ٽJc��g�4���SDpp�Q�9˦k �i�)�e�,�/�5������Jz}.�#
|���G[�QX�j������ad��U��ل'򟖁����n܌��z^�x	'��{�6U���;�xM���WbYs7��dyd�5��h ���o�ә��z@�?Èϗ
%�ʥ8~���yp�M����(^D}��P����:۲&�3' .���[췫�J.C��[+8=Zf��;�[$�\N�Hr�I���>�Z T����jwߎ��}
e�^?Ӷ�R���s�MAh}��`�ށ�e�nDh[�DAB�S����\jӦ�^Lz�8vYST��Ɩii��RI�������g��ы��E'�|G������G�&�)
���bl}m�S��u--�j*7�
ì?�[�V�b/��Q��J�<!����ҵ���fd�!�|t��N��{��V�kީ�# ������t��4������pq{agS��ُ�s5bk.�<\�i�0MY����T�t�r鉩:O��� NY��u�3+.�p�ԩ�^��K�,�A���F+%7��v��1��RY}SaM�L��Ბ��.`C+|�E����d���� �[��+��ˆi�����teѮ�I<��/�<�A�惤�Q���~�_����z���$�W*4�1��꘣d�w�T�'_�VJ��z�ђdo�ˬ�օ���ycHk3���������`��A��w!�Y�2?�%��!�_�W�^�O0���˜��l��u��}Qv`�rܺ�Rd�P{������#��/8��Y���(��	J���o�ĕf���h�mH��>��|�N8i� �[�:�n 6N3@��|`��(���Z��Z��pE��-�HN�$�����*6JT,���52eQ;oprJ6.ܱĥ\����Tw�g��!�W��\k�~@.�gs=dW���H	�v�]��ﻵ�:k*�9(�����m��J%�0��L�v���w��e��G�c�MD��Έvh@�N������c���܃�:�-zeP�1*�͊@(����ZMy��;�^�YɃ���?N���_���A]���.�*�n�5�4K���b��"�:�8��hٓU� ��Cb��5=�A���QT����"q�0��dݽ�m�G�����y���gX5_u$�/ѥ��-$��W�J�ș!��AaTB�G�if�jLV���y��ߢ�{ǖw�*�'z�h�<��_��T}(K�O���ki/X���5����% �*�p?B�n�1LJ8�F���`n�v�љ�t�~����6R/�,����Ђ���sy7�G�