��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQG�.�����t�������Y���{.p�i�O��dg�~�D>W�Vp|�VzL[yXJ��@wf�,D�.)�ot|O¼�*� ���>�g��?�C*^e&ԣ�'�k�����8Jՠ�Ե��|���b{�ݸD�g����y�h	�
.*9If�`��zb�*i�J�����4����c��UQ8���K���V��/�*�g�Q/%��w��\8�S�dY5�d�kM)h��T:�>�R�XJYI���6�/����q{�ҜO����~��r��6a���ߴ����,���ƽ�+�7^4��]V+���E�^/5_Ż�X*�o�	n����&�j��|òGT���$l =	����1|(n{Փ��w���x����b�ahiй�3bsV5�gc���u����� �U�$�*_<䉺\��&����U�9��'5�OR��Ӌ9X����x!�x ����Ю~��Ń��~��=�!��`�h_R�y��d<�h��z��j�"g7̶�����B>�K>z異�t-���3OC[�:���xN���v�J�Ԟ�;�n�5���fg��[�O�Z`���/\ ֦��tYI1��*�&����R{R[����V�c%:WW�~k�����U��g�Pk��!.�����wMvT�BY<ͦB��z�?j���lh�E���V���:�yk60�	�0�l�H���R����I4u�{${!D�md�諾=��#Ѭ4��HP�i��ӽ���Eδ4��WY�=� ���]ulȫ�o�FY�1+�j�#Si��ĈKʄ��>����G�z�qw��PI+���x��W�S\����"��1��(�U�e��?�f|��cW�x��B�}d��4�]�B��0Dr��)N��,�kg�X�Wnr��n������^�ǬfJКT��?Z����� @p9 !6����4��}N��6b�!�c#-G�k�`�z�.�=h��u�&4�-��Q[��n?�ko�R�`�2"[	�A���b�t��=�����^�c{�0����Z��1Ŏ%�E���u1��;��!\$��y�&n��3�k����o�Y{����������c�V�r&a�Ω��D.v�D�Vm4�yt3*��90CT�2��Oz=�,L �h�G�px�H`ک=�nC;x6�f'|��=�����%������!1ri)��܃���}>��|n�P�6JWH��|���物�qn@���rf�%���\*#Zcf0%����<�yފ��l~�Fb�V�Dp���Ub�Xr�ϬOe���7v4�Rh�4���^c��F.���q_L4/cO��N�T1H?U����W���{f~4�Y[u�~g$`�>'�/�-���l{@��ռwr�Pi�N��96)_:���0𼳥h1��t�^h�����7�*@��R�Ļ���t!w�feA=�&3r�:�5'�ꈞw�\k�ů��)�8x ��&;��VT{���[f�G�;�-ͳ��|���;|��*="��/���D�WR-�iGnߋŰ��x!�+�m2�[��fѹ������l��ح�ta����a��Yq�k����"m�������2ZG���*�w�w4�ܔǂ�(X���\�}�k?������?(e�\o������ʃ�8�<�h���Ű�|��^��֐����o��B��*���#{�	 N,�XQŷer�_������)�0����O�Q�N/b��x����#κ��z�]���v�$���}�e/蘜nRT	���NEy���?�K�HFJd�p3^�"ň7�mSm��`(�L%;��V"&o�6/��Y�CH.�� �:T|S��A��u
)�;EE�9��Is�G��w�_os��W�i�O	�W��K9��W�����?p$�
���q	ߏ�?p�����f
�f@�b|�a�Y����F�6v�%Z���^m��\&��zh!��_���t"�sO�ؠU%I�)��G�I���F��=|�h�}Σpx�,]�q�C����]������������8t� .��BUK�n�~��#3���Ҟ�m�+�F�ݸ�Aa��׵�:&F ƀ�h�\u~β����<�����hذv;kIlSS����pI6U�kuv�t�v#��F�-�_(��i��Z�H��o<���L��T��Uu���l�b��)0ߜ�t�$����0�XN/�g;���A��2=��d\O��
smF>;�fmx�o�(�K5����	e����n���Ӓ��y�W'�p��n��S�516��׳�4�� ��#���r�9&ϓ{s���1�}t��q��͑+iZ'�G��M��BA���{ڧק��#UP=f���|ϱ��n/�[9���Ir�S�
4L�b��v�6�H,�f��e�C苺�7�Sr����k�q�j�5�bޔ@�R���ҏ Z��\*Z$�-T�����[ C��DGzR��;�]�����J:�����X�9��3�z�7� ��<��P��?LO��HY�b��],*�� �	C�"�*$��G)5��g7zZ�
����y%ޭ��~�����T��-�n���W�11����FW�9o���~����=����
5�����ͨ���<kT��X���%G��{��#���r�A�v*�+[�b$�/��s-$.F@k�Y$Nx�4*l��v>xmj��b�g)���]��m^R"�\Z������d^�Ut;��q`�\�4J9��9�fj��TkN�.)�	�3IuCM��ٞ�;GswF�����	8ES j�A�V����^�l-R��`�N���l�,��j�P�IA�r3�� ��
'|�!nGچ)%x�)�NC���h`�n���p��ۣ���h��e��$g��ԧ'�dA�����D�� ƺ6L@7*n��bY�$�� ��S�(���9H2iwA�.��7s�a\״��_�r�7�������������6Go�S�x�\�yQ�����5=�(��]q���y�ׁ}�����E�����õ�,���<�ՏNJ��03�IAA$��{D����q3
��������L�	xߋEԛ��t�*�9�'���<�-}J:��8��&猏�t����D�eeC2SB�
!6ٸF@��:U�bTJ9�ݦ����'�sR���`�ٔ*:P�Z3�\��?�a�+$?)һ�v=��������ւ�M��I���h'�����d=6nLi׼O~�^���y�c�3	���B�6��Ve;˜�_��ܶ� mر��j0�킐��b�����M��vdJ��>mi��A#s(�s �pm�s�]8����R0T���c�1��h����îU�ޢ�8I�3�'}���0A��I�����g�ȭu�bur�)���ű?���M$⸲��i���آ'���
�ԇiܻ�pg`��>�������3����@G[���PAhG��,Mc�G���﹵�����ܦ��К����]U�ɩo�ߪ��R�?���O�$&�1�,h �Ԁ�����aNΆH�+�L�~�Kǀw$i�����Qq���(�����v$9PJ��v�1�~l\B����N��YY�d1X>V���m7��e��iE��={p�9�
N%�6^nZx���V<�J�I�qz�SG۩�5�7��t[��Oc���k�˙�@{��֓�k��^�p��:�����W?�2�b<0,�������b��x$E��_� t�>B��RM�����b��n�%�6Iz���k8鈉�>���)7zTm:A���,�E��O34�{����@���c�����V]�?���wqٛ�-�tGE�[��d�cP���F>҅fW����Z���.�BT��V��{<�k�a���t�DD��)��+��F$Y��������������E�DпP:�*xX>|L���^3���f�zNZF����K���&��5�R�(���E��i�O�exc��h6A�BA��\��ȁ-1��gdG;�q4~=�z���N(����"`"�.)�M�>�p�!zx(5~��Hˑ�$&_�}Y$�����&�݈����Wy���X�L�m�H��2)E�l�'��%���th�Gs����bvq��I��4���d�A�7�'#|^�ցn�k9�<�
K}M�M��R�����.������&����HE�0X����Z|�FX���x���i��ђ�k!�~!�)	�=p�s�;��H��cY?K��_@���'���ݝ 9�?��v� �h�d�7-���d>pܳ�N"�I"+�7�?�P"�I�O�ų#���}h��s�"���іo��l�9i�ˏ/3Uj$r�*���N��f8���>i�gOB��Gv4`�=�	���oI����2
�-�uţ�MO��Ns6�rƇ<a#�E�t�`g���)�u)2�`h �l�Ҡ������O��`�>DN*�8�Z���9�٥�c�#���{�j�+�,���?f����8r&vT�זI�W\`�E� �����˟o��;p�䞬��pS�xK*G�Z�~�&I�l4��ِ�c'�XŰ��6y�޼�pszv㠩Jr�?�%hq�b@��%jp�lM��BԳ\���X�~�>�ިX��!����_2?XQ��0��u� �\�*{�Zl(o"�Z���I���Fe�%Q�	&]�m������彑�����!%�	��-wƻ��z�@bk�w��=׮$q�j�(Q��%��{�sy�;��3~�Q�~|�h� �z��e�#�Mj#aܮ4��b�Kr]t;yc�ǋh��
�~�"�hE�&�L،���S�Z�w$&��W���UY����)f4����;5E:g��{��@}���.�4��j��g��e=��-8�ޱ��䮪��X|l1ᑑ*[V?��3���BKe�C�q%��	��
0E����~X��}�ö�;�Q�ө�0�c����L�Н�^�hX*dS	H
���&	�^9�D�\���	es�� ~���`��o.�~�P�*��'9�pW�oD���U5�Y����,��ۄ���gu���'נ{������� ��3.�'���jޖ������i�����̺��7_�wf�P�R'\����j�� ?���T���LMR]�����45s�F��g�e���rq��5kh����9hv��d��v�}�x�;�0Q	ǽv�6������4��L����]�+�%�gi����_�mP�jY2�B5�nS�(�q)(xz���z!)S`*��V0V�c��z`H-���u���}���ӒE8���ŏ��W�[������9�WC��+ou�nC �Ş3�a�g���H�&��x�����vC/H�	�UK���Q˰u�[�Fap�G��UG%�FEr��Ӗ���}��ޅbe^��#K��d5�.籼G�.���L<��=2�FiF(|��Xv������4��%SLN��Q���L���X�b��LD���Z0ܭ�