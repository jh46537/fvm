��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���^�T-��!#��S��v��\ixF�u�qb��tˤ0k�u%�k���?��)��R���Ǌ�Y�t�IB������O�O�R_���(}��i�F�ӄ�`厡S���IN��D1̯�'~�wR�n@p�7,�� &ܒ�q��_Ma&X��p�/��5��i�Y���N̑,t����vl���f��;Ny)�pi��gK�po�/�a
��J���*7!%2���I�c`�n�T�?�]0�ͯ�(f��B<"?]<�`���z��-5OfÏޣ
t:��M�&d�e�����Z��8H��p
�tS�a��&�	v�� �Б���~�(�ύ%�s��v*C��j]���X�)�=�8�fLb����n$�3��m�2��䥏G����16^��|.](G���"۵�u	|�A���XY�3��I`�:k6WB�-T�� R��;U' �m����<-'�X\6��\IBCh߼� L�'1}��v"�/�/P�}@͉�x?�(R�g��^K�[�4a�7��Dh�~�f�AlâZy!�6�+�N�/V�U��.�('v��q=���<�n-um_�Zk�1��_�U+�DOɷm^�^�����T�;�4��2��\�[�j7�Aʜ]��]�`��{�4�溌k,�^~|��2Wp%6Κ{�Dg�9��͚xM���?��k���5�ν�A�3pj&����r�@4����:Rq���o�WT�k��Χ�ۭ{�h���������lp����
����7����]]��IB\�*ӀM1adW�D�hb��e?�I���S�h�ysB/�H'��h��h��J�{�v�&s	�vh�� '�[Y�H������B��%B�0#���y}V�e£�I�b�T�A�R�	o��b?{[ʍ:J� ���H�Ŵh�+6��Te&��&����)H*�j�x�2�Bi�t�٦����2��^��u�1ԣn-|����e��6DnО�����Q��|jw�4s�L�7���
m<^�ҥt��d�tY�>�͘$���Ӗ�I���t���T�wo�7�;|g�y�cQj�E�NVz"�ދR�%w��[��l�3z)�%JM����*8�[Br�;�A;�5,=g	��~9��R�s�u.Lo!+�.�i���(M���Uu����凨�$�Ђ�=�\�S����N!�a�zg�ǝ�TC5�>'Ԋ^p�82������=�0ol�^��]�/[>￞+窳����aT��&�}�i�q�u��6���R=k�*��J�8ش�fd�Ζ��L՛��?^GIaۥ/����\���U�Eռ��b�z���id�����FG�B��١� �.�~�)�
�V�n��ڍr{�@���XCJ����M ?<Z�)hڌ3Y��������V@g�
�o�Z�` ՙ�G�7�2���ZX -��D�
��k�ZC�b��/�s�2��Ab���̬�G�v\�%��gP�'&gƿ4��,���,��:0;�0�sOeRȨg*G!����i>�ߪ�>���:B����W�k�g���܌S�����/S�hɳ��%k��	�5��K\f��7#Nih�og8U��ĝ}a�YX!���ә���x},77?���T�sțA��dI2�Ff���e���P�/�"H$7L�VNzH�+yK��ӽ