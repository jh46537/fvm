��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�ӿ�J�r���>�҅�N�Ŀやq��,�����r���J�?-�O��?B��<�ce�o,�`��<�OSA.��=��r*��n���X���
�*2��g��gY�HG�2���Ý�[����=�ӷ�k��ם�k8#,B�z�>>KQ0��a�3����:�s���)��A���p��j���y�<����Nد��.l$��Hz|�E�"
�7eX�(����I\sL��
���|I��
�=�X��3�a���ы�<�-5�v��gJX���=/�ٞ́Y��V�h(�
��B_O5���cɊ�-$ѯ�9;�mد�C�����[k�kEP�� �\�����!�vr��~K�v��K��[G�f��0C֍�h�/
^	�l���m�T��1��W�;!��-P���-o�m���Ć#���S.��b+�
�'���*m�vq)x��[�)�fгa0zr1��:K�G0����e�҃�X�'��Kt_0L;�h���Y�dBq���h{�ie}@78��|�#�N"r����YB��0J7;'0E]f�1()��[�=L��ݏ�UO6R3�i }���yB�H0���ę�����s�<)��w�����d�?F;�Pn'�íE�+tǁv1�-7��pu���s�7I�}��}@jm�B�7s�
0p[�:NV����Ġ�[�{��2~ET5�
k��x6�u��_�����>�o��8K���z�Í�c�;4��L�&Kv
��P^�vy�KAf��@G����G���< ��-|�Ptq�9 	�B�L&���Aª���Z%aY�H߯��/�e�pE�����m�h�]?�M̭^���<�~w�.�G}a��,I37��0V�/�=x����%�d�n{Й^Ý�<���@�:�㗒�{��=�3����Z���ϳx%���+{�Z�|��8L���(�u�>�����.O	!',�%㊚p-��~�S�c[=s�w(�� Ӳ��=b�')-�}�g<��s��K�Z�9�{��J�� ��+�����OMb���B�;��+�F?�M�P�M�.��srp��M��}$��B��{S�	��~+W�#�+�EJ����zї�2�W6�B߅��o��
#�1�1󟮭�/�ۯ��ÂC4��֕����h����7=�I,��JZ����%lE"&�Pn��3xy��W��P�9�����FM�|�j�Em@*����N�=������i�����c���
��AK����aM�ig�;.c@ƈ<��"�ㇳih"�+��cĠ�����,���
��ܲT\4�VV9k�b)i�l�c��&��в���c:'�Q3a�4@#k#D��s����@uA% 	ԑ�;��W�s�K2��|et4!��#��o��
�����V�h0Α�2�؊f����8���|Ǘr��Td�
�x��,���`��˧73�9��\Ƚ�3�ޕJ��I_�
��N?�-��\��E	��W�˅���6��g�;����8��r�̸���]=��}�;=,��m�q
�Y�,��%Y�Tk���X2
�Pk�oH=�=΅Փ%����_G��%R�<�L��	��$sM)�闊���Y�;�F���0�_]���zX�S�W쑳�QwT���� �D�s��`�ʁ�\��M�%(�r��m�f���a���[X-�b���D�+tW���U�݌�sU+�,�eo���}D���3���n�i����)�I���i��zO�dٺ�3 �Ҿp��f�-m~&�^��b�,n��y�#� W>]6R��+s����s|��F��Y�����%�.|IzP�p�KS�gTTʣ�6Q���w�V.Y@�;�DYQ�%�"U��xh��6I���W�=DO2=�wI�u�O�:l����]�i�A���8P	��&��N�]��,�渠��G��9���3�*�L��ٶ�9�]�Q.�T�	��1�g��MTDثͧizT�[�r�
�	<�{�i�9��9ggX~݁)�\6&��`,n�6:�(� �$~2��E]����n�lP��;/���,G"�,	g�M��Zu`�ZSJ�X� �5#�E���{�3�V;`,Z,mx�z�]�;D7Zw�)u<���c|�>1�h�������X��"���Qf�R	ܽ&�T,k��!��ːk�%�O�Ӡ�I��~���^��bQB��A�9�GEg�D���C����q�
��@�c�9���A����~�����Km��cO�Z�����Ph���t��Q����b�1~De=6O�om����ZZ�D,6w2��!>}_%b���8A2F��+l$��k�
�߷�D����՜��P��	k�j�2�k�2��x��b��)b�O����̞�q����jͼ3�� C��absy�*+��0)W&p�u;���d�<�{*+q��z�����ʇH:Q>7�z���y"��K9ْZ�����	KY�u�0�����pr�l����I.8Gw����7\Xi�B�1�/�'�Oj�L�SH���]�j�&���6�&^L[���O2YIP��5\�L�jN�P�\���NU��\�`��R�A9\ӄ�������d~����̊��!�g��N�n׻Cu��E��-��\~�ћnV�S��m��V�WKޒb�iM��S9T�P�!�������F��?�'N���0��hj�MJ��<{�v�=
���a��e2P������`^�����9 ���3�!��M�h�*��d��I��$r�hg�B�%O�P�e��13�����������Hk%,���D��t
��`o��2�*�Q2 2 ��U�u�Tl:������\/b)e��#�Z�F~7?��"媉�+���XW�Ol��O>��	�}^,:�t T����TQh�\���0�=a𺕄��6��6ٱR�c��5]��1²�'{W��jS�����[{_�Y�t�7O���e|�����Έ&o��3�?�b�����Ĩ��k�w��~��Ku҇�{�J(8�,Uy�v��Y�C��� c�ܽN�ʓS�IA���LF��6�e�H9�xz�7٭t �{�(�*S�|�5!)�-[�l��Q��M~�5���En'��>
]袠f����vO�;����3/�������J�8������J��P[�HG%���Yiz��� j=�NO�ϲ�D��ЕLv�����q����r�R�ASm����^�ŋɚ��r<�Qf̼d-������++J̸��`�
8�T��߲�~�ptcS�7XȁS.ӫx'��9��mQ�����ƉF��N�X*�Q�u�-|����eq��tY��x��
Z��V�*��� T��K"j�?�H���4p�Q��9�n�j#�M�l�IǸ2���4g6�]c����"��He�T4u�x0}d��<��T��@�($�e��#&��tOF�Ø+#��	a��q�;[��F:�R6K��S,q�s���4׿PMT��4/r	#�t���'�&|Z�%C�#s�/8'-� �	pz��#W��GN��u�mZ����IƟĎ���I(K>q�Z���Gg1k��u�Z
����C�02��j�>Mi�D��#��e%|��R�x	��?�S�A��5�o�E��H��hu�y L���"�K0U�sZ='�O�߄�n|8��U�u'�[QI�9W9:��c�%#�2/q��s",U7�ό����n� .�.���e�+>��V�@��)Vk�{�\��'"�lk;X�&���<%�fU5����@�^v��t�XKn:�A��n������
�g�%�_ق�d�Yq(�	�I"�R~T�<�A��V�j=��ow���!œi�#7��'dZ�����G.�~�d�!��
��A��J�_�|�$�F�d_�
v��͞��d}VL����\Q}ͼ�g�;�	 �	��
m���O���M�k<G-o��݁p�b�w��V�.&�9�*N �x��x��-t�sB�aa]s#5�UtK�9�\u���8b��kM5��.Y�c�к�J�in�%���ҽK����e!�v���턹�tn`FF���/��;��Gv'߽u�J�h� �E���@`eCCg���b0>C}@@�ߖa��,�<:T)q��� �	�AR�rP�����dՃ�C��L̏��{(�[�L�0�|�~^-��4؋�z
����jyc�U�T� �QU���oȝ���3p�� ϤJ�χ,�8JϺna!q��>D4���\��i#(Vv�3^.�J�φ�E��9��a�>3K��䊫��!�RE�(��艣
c��:T��G~4p�'nes�5�p�;YUM�$Oy���ǟ�����ŋ��>8%���K�Y�|L����0���W����	�dA�'���� W���Б�po2|co�G���Y����(���ĵ�{'�~ �Ȗ��`�o���#�m{�U�IN��}l���5���f��P��>x�j�x�p��쏢�N ���-a�b�Y�Hx� óR!���D�� ��.���.�0����}�6<h~��>���	�9Ղ�]tc�`�9�6� g쓹���33k�5���N4b�/��n)���я��NL�%�n�����U��!읓jL#��Z��ùt/�|����9����Ƴ'R��l��,ؗր�:�Ԝ7�'��8��-��{be�;�r�ֆz�V�F���C�%�`�|�9T�IZ�<��I �g��GZ�EGiUսO;�K�7�I;%esvm+����TPe�2	�6OG"�ǽ�����|�L�o�e����:� d�h�B�ÌV@6��tV\�f�A���50���4�rLat�q�i��HU���c��!�n�C��/�AS�|��1au��xIZ�s �;�$�M3����,Y1��1�oT�i���r�B�q�<��!ֽcELE���::����RP���b#w-
c�ܿ٣�|��o�T�GI%���)�}�.B�E��cJ��I��D���yW ,%���$ ��{N��]y�^ Y^��1��FgYk��`���4ڕ�,��>�wbc�楙%q=��6RSA���Sz���r@Uж���ǲ���"6꫰�a�D��Qa�O-קn���r~HN�"��w���)߰w1��� Zґ&�b-�0����%�H�ȴ� ������@#�`lZ�� X&X2A<r��"�<o�eG���]O-��~H���Q8��*6��.�B_��_v�4@�-&�M�83m����Dٺ���?���72[�[�U��&�}�7~�OW,vQ�n؃��>��;"sClu���K�-
~�a�� =g�i`$�hvؐ5�+�i���I�ӗ?�3G�'PC��˔�J�����,�M����)q��uB��� ��m!8�ջX��o������.zdX]m�_]���Y���ɚ�.^��G*�U����0`j^S��t�:N�MWBsZRmgUX�ct� �>N���������.���{9�k��P����8�.�P�Gڟ@I\5,N���뢛��^Ѷ� 3���Ҙ�SA�22P�G2�}�����_dĵ�q-�Y �x�/@9�˭���^�VC^f�� j�dh���[�Ӊ����o�}"��y0�{�O@l,�D�)>Re$�"���tT�;�g�.~�p���w���\����ş�XϡB
\}��*0�zsW{˃��3�z-@&�j�INg(V^�+ ���Y�Em��Y{Q���I�LЃ����[qZ��	3�>�ք������v����<:ek)=w1lM�Xk�;P�Q����f����=��j�~7vD+�M�c�.�QS��,N(D�d��3!���{/!f���@f�������MR��}���1neI�i�e'OUmW/��lL�����,R�+�f��r��K��J�e�;E�����p$+/��4t}F`Bf�� 3��Krç��A+:lj���w����pW�� o�5�0�v��V`!�B���_�X��[��+	И��8C��bVSO6.t�k�}7Ӧ���������GD������K��ҽ$���"�3��j��$@�I�.꺖��4i�!Y͛�,۩$MswVo�N-]Q3�y��[�8byoX@�����M�����5���x:On�pp��y��3�/�|f��З�'X�v#��=�b��Z�*��Κ����_eU��ja���饈�����_p����
y�J@�H�x8����9�s�޻���G䵣b���BT��ֹ���ޭ�ذ��Y5y��‖��B��8e���[�A�5����^�&^�.�5�( x��oZ��ܪ�*�i\��:�L��D^�?��X���A�^%��?���������阙�u�V�I��i��j���
�`T���X�Y����q1���h���D��tX�[��X�
|�v��?w\��4\��]�r���~���4�+��R��N	N�J�9�ܕ���tJ�4A���3=��??����䢒SrL�i�rF��)޼N)��Л�#��X�Nq>���냹4��h����wr2�6��t)ϕв�0!ĢtQӖ���ʾPn��Z$�>"��A���ׯ�7�Ic��;��a�}9�sq�,����Jj|@�~��H9R��z5"�ƀ�j/0�/zN~zX�c�`�B��&苖���W	�����?��5�����*s��KS� �:��d�+��*Ղ,��D��I�xCr�K�8'��)�N�t�
*)G����5��ql��MT�����f,M!N�j+)�	��0��9u�	���n=�5��H�)�L'�n��R��@+�l;�o��kG��Ϭ���U �Q&g����u��1gb��O��������]�����T��bZw3t@�}��-c�h���;����h���@����ݾ��<���]�갷�}.����ٌvp�6��)����~���m�G�a�/��0��P9X�}�.�jE=� �@��.��E~g��p�>��I7]tJ��v~�봶�iP���"9�lS%���e�ϟ��z�{� �����h�~�z��XUi�~�1�4&Xj���D��Ŏ�	ke��aL�N��|���˭ަ�)t�<���@�ƛ��E4�t �?q�K�TPp-�=�=�������_x�Ma3�ɸs&m$���b������V�
���O'��m]�t�0�oyR�F��#�W^����hROE�$Ӌ�<��և�뿖�V�IH@�I{ʇ�Y
�Uӂ�@[6�������j��|-��;O��%R���%Q0��cP���mPQD�F�ě? ɂ�ӀX��=�7�է���j�}=�(��c�6�P��b�*u�%�l�Ϊ�Y��%� 0�CQ�z�0���#�J�'�?XU��������&M��m�����~��:#i}�Q�CqWjZ_m�c29��F�"��~\�s�L`������7��E�2*,�k�ϋVyQ��Efm @}��ج��3��7�L��ٻ���$��ߡ�?KØ�N=n�(A�V,V
���:b& B� &)��P�o
��K�&�=n�Vəp��3b��k���D�9N�)	��>����
A;p�6g�N3JZ��h�U�`'zC�H�Z�.8�"!f�K���e:�r�=�fV��h�L�� ��ơ!�p_��B<��o��W v������Mk���EvNߢQ!�tܥLq���Sz#YY5ǳ���1f����A�t��j�,�����Z�G�ۺb$.��DX�m�oW���D?�;���
��UB=N���;o�������L*>����@yK�kH����0��R��6}�fu��05fĉ���cR��q�f��j.��=�o5�>��g�k��X�S��z_�t�b<d�ѳ�!?`�(�f�%2߻Y������?D�=�kt�n�%Ʂ������x8/��TT�Sj۸��g�1-5���w{|�,��<3��冮?&�o�8�uV���s��)U�V:��sK����cFԵ#]���T����Ҋ��6b��ϫuk��i�Yu��8`��-�B46;\��W��4?X����tu�����bq?���H��a����x
���L�)h\#v!��g8)3`�vI�啘Lg7�%���FC	2V�t���W�G�=�<"��>�� 3HWk��ӏKףmc�s�t�������*v_�&_'�&fo��+m` jZژ�֍)���&�TN�^�=w�^<U��V5�]�F���~|�8�X�q�Do�H}(�a�XQ�.Z=V�-�Z�ƨ�H�tD�_+'ԙC聤��'����&����
ѩh1����U],����ep\�E��S#ʒ���S�����Z�ǵ�2�t9� ��\oyW�g��ǭ�tv^�`D��aS6;>���}�V"v/�iPw1V�7È����L/�c��v%��WE�1��k��oƥ�(t�t}
(��cjc�$+�ϔa�b��zFvQ�Ί��̛�\h����!g����̐-t$��D`>�˄�����\�G�]��I��6�k�r�w�aCu����:
�������9���Ĉ��O�������L(�ӃC�НU�E�p)�|�>�!Qg)�4v����)��lk�K��==�M��埏��-|B��>6��tv��e~�Z�V]B�`u�Q� ��6�^"vNE���'ṿ�s���3�>o�K����ԫw���5�"�;q�ت$���)]��Н��,��b�G�BP �^��XR�Rz@u�Y�6ے��FG����7<�v��M�o���de�H��$t�#�>J3��%�FD�F0&XB��ޜf��.X�����h�2����m8���X`����H��!/�'{�~(\!������Q���bc�v�h
��q�xQ����1�T4��鴰��D�8Tc��6���F2���?2|���4 hX��4��#�~�xI��0����n\h*��gc�]q��'�(I����朝�Bi9� ,��{�������cpyCR��)zJlz�?��#�2�aB裳�$���e.r��W�U=D���7d�#P�=��c �"��K@Y�Sj
��V�̀���v�lZL:�b4��t�5����?�S�Rӊ0��!�Г�%3:ƞ'�.r��*̠����6:^_^V$�2��/���]M$��?�(y��[ͬ�|��':۾|��_T�E����MF�EAYJ ��P\��'����#��=Rg���������Ĭ�4_T��0)�N�cء��ѫ��Qڇ����p��g=�A�d��(|5�\��?���Φj�.��]��d�#�,ۇ���p(�WA�	�aK���ñ������t�꽐�Q�����b���1�p{�D� Q�Ns��9��*j[E
rC3����2Q�c_���"��5lM�9tW=#��v��Y?���,�+�����c�t*�M-,�hr'Zr>O��kl�-�hzq֫�b,��z,�S���t|��Ot�EZ,T������>��V_|���Ԭ6�}c��T���W�ϯ~��@�Q��6۹�+^�9
֤�8yDAV�ٙmw@��# 8 �f��H\Z�N[��I+�G��W�B�:^��Z����h��-��?�6���m�����XQ�/!H��a�Y2���^$Sل�[�#��sɊ�̣���&�"���i��ޭFEa�TsC�(e�$�c�-�����n�L�nq�BA���i��)�? �Su
]��| �]ʊ9]���О ��u�9x �Kl�*9���Gy����4v����xxV�8�:|��7+�s���W���5���}��K���&�ԖvS��Gu/ã�m�A�t#n�'k��"&d0�Y��5����Z�Pt�^�ܤ�T�*�*VN]����+�Y���d�Մ8G8��]+0��$59잽���~��DC���ٵ�+��O'��1���ۗ%���-������τ��cZ@�.Pމ��P��&�F�L��z6�u�Λ}��C�<k��k�`�2?s�5��s�,�ր�����{�x��x���{D��;�]qg""���z0���չɍ�9���7�`��mU�rԧ�8�p��)��g;���bJk�~�sS�+�K�F��v	��0�t���y�i�s	;_#}~XӨ�,5R�23Z5�q%36#>�� ��a0�\��9Fh��x�ͨ�ݭ2�(��zv��ۍ���d�����!B?ջ5,�Td�ki�P,���uV�@ �[����d�,v�.;���8��o���d[*�;�YK���I��|&�g�m9�c�a�5���B*?�dk@y�����B����!�SJ*.��:�=@F�<&5ā?�QD��}��gHwޑ��%q,��� ���Ҍ�v��#����4����]G��aN��t�(��@!��0�ln�>q��M~���W�Bq�z���q��d�~�VCX�ޠS`�%w��n��	��$�<���z�4X� ����b��gڒYr�}�ty�3&:�T�mZ\^�dXG�C(�A'����:-��3�R�R��$T�o�P�K4L�عy��AC�fkc��j�K'b&�L�N���3�RZ���4�����W��o>7���k����z�^�������M�/���Fƈ�Nv�H�b6��/:�#�����_�Q�k�࠺]�·���Z�C^�Ds���)e�eJXg�D�J*�Q3i�MmP�4	�ᦶ�������U<��fT@���a�^��N_��i�nz]l��5��?�R���ٖ�5�Sp��??8oW�^�o^g��T:k��"��YYfv���ӷ���@Vui� u��4�H>�c�p��+�"	އ�&���Yg�&��H���L��J�+�7���!β�)��U��]ɩ�Q.0�q�͊j+e�)^���zIc��z�ls�lGv!p4���}ڵ;-��jT� ��ѫ;yDKha���w�`�{��l;� 2��y5BR�eB4�r.�Z��͛�#K��m�t-�������� R�3]�ՈƳ�@��c�5{\� ���8�U�=�	�HH�~W�u���92�] �`�JYFAg�� F���.8G��Lc<.ê�N?���&^H�>�%_��(���ZS�ʳ��y�-��~m��g��n�-4����ݞ�s�����)V���8�D~~����ȝ5�nڡ�.f�����jhᰗ�C���ۊ�u���z�|�<	� ��LDk��iO5��Ώ�<*��w�����Bm6�2�ȅ�f�x�iC�	Ñ+���� ݬ��`xC0�Mw�y��KdZ�����|@�e����<�q��>L/oH�0���#B��	y����_ ��[4��U�3����S����PDe*l�_�F��Ds0�11�������l_��"x7�E�&�=�Mq���[��\چ���|�j^h-�𪐉p���h6ꅕ����Ж�x�Ұ6�=�q�꛼S�i�/���V�_\æ�m��דb�]
�X����@L�	j�`�0��nc�ʁڎG�b&:�-�-%����".K+�ri��`���c���5y`�m��}F-'�`=3;�E�@E}��P�v�0�&�K��FC^�nN�Uߵ�߮��F�&�o{z�����̲��H�)ioB���]�˹8J^����Y��\=�O9�,��}���e�0:ztz�^Th8ݩ4�m�ؿ���Xy'�2�Kq`��٥��Tx�^A)F=�؞J2hY�oC��L�/���ڌ��1��5*u�mFki{F��2=|2����0A`h2%|�BI�[�D�U6Aiz����6�Ƹ��U�X꿲@.�Fs�<s���y�t�����u&���0�8���Ӯ��sht���PC�I��z��:�����]��{,R���U�e
_SZ�W[� 
��_{}��u�x���u���mձ}:_Ԁ]~�%k��,;�Or���E
���u��ȵD����AOv&H�Q%8�m�C�̤�'.��uzY�^c��v��-�'뿙��Qy�3Vo�윰O��&KQmC�-56�=i�:��yv�W�w:��I�uc�����`� �ފC;A��x�1-L��A/�j� !i��L��Y/��������՞�]��ƽa�d��}��Y�ޙ�ˉ������@��ˑ:��e"z�W����|���f
 �1�
��)bI�����5�WP!<��3��2V��܆�0�Y/�8?D#z]tl�M����(���9�8F����G�S�X`ǽq� ᳜ܿ�;�J�W{p�cJ6b�$z#�kK։>?<�{��Hן{���(�<�'��[t��rvB�(i���(�BG�v>����1 ��aU�˿���QA֜�WO�$?ac��8�oү�����j�氤���Έ���?��_Zx)F�}c-R�6���Y,��Cm3D�R��M�J���i�z�T%�O
&z!�|jյ�"��ƣ���3m�sz�3��I�z������B�7��#�;�P|i��3����>i=�EC�f	�u��c����*j�}�n��B/?�V�ר):��!�6�j�s�j�.j����%}; ��vXW}爙�.j����@�C35���A�M���'[��c�#�_�;J��%rT�/S� g��Sۆa_���!5s����
�	:P��U읩`��.�_�D�)�[z��,^y;�� b��5�٫�^`�Q�N�?���
��Q%��6�oy�:3q����ځQ.�Ua�+U��&����Sb�0CC>Ƈ�n�P��u�yG`�� ��~����J�������2�9IJ�T�k��8Y�.r��k��|�(� x���'/J��k�ZN��8�W�)��rwW|�~g����:�79�I��@����nr���P�d󱗻�}�i[0Z�}0�T!�o���(+|�����e��?�ӒI_2Q;�Z�k5*5ٖ�|n&v=�b���d�%�8�?�.#��86vn���~%�OO!�����S�X���!O�����!'SB;����\Th��h�mm��靧�7����.��b�)���%2=̩h�5O�si����F��v9`�aɑ�gk��0���@�19�@Nt���v�9
�"ָ��}�5Mᔨ)��]o$��HfXr���#k�6Q�LO��܆�������`�U�&�A8�1�
���u�	�)�5k�"�\�OR�8Tf���q
�&"(������]��O�s�`V�W�&ɝ1�Qx�K����7��n˼ZLϤ�0	�b��
�
��8$g�G�u[9�I$���5�%9JC� �:o&t�����w�u���y�K�����^z	УTf-"��g�׹�Z�Z�񸟅��y������pBw���q����n��A�����������.k񋑮�����o8�e����c��J��?f$C�f"MUψ�ҤP���`Al��dC��E�Ԋ1Ac�?��La;��㲔)�Dz�5R4-(�/�n6"������2�;���{�?d;�8�*o�]PK�
�nt� �W�5#:ʻC�*������,��[��'���\G)��)������vS7!�`[{�,0H�)��/�o��'��?Be -	*�B
8��v(�I9�&ՠ��|(af諝��3uЫQ���*����\FB9�Q��ȴ�q�ĩ��%=��yKY��鼻�i<
<���p����;e؂�A�Q�r̝��e�0�����,hc]�*E��ಠ*��������k��}���ر�g!E�ήT,�%�퓟[5�&���d��4�QzF^P�����?��o���a(�]������z��ےG�\BT]S�/���j��yu~H�r-���>�J�x�wf�-�&���pp��v�n���P��z���d�vq�--��xjf��=�3jwkYv�b��9�ȵ���mJ�\� �x�釳�f���0w��>�� ��R�!��)2�����K�h>-JyF���jn����@�Y`SqO�	��8%}�F�Ϛ�zЩ䝞���|���k��P������tp�6�lߚ��˧�ֶ(���l���M�Bl���{T��,}���"��c�l�<��V:�,t3K/�H�R'hؗ�	p���|4�ͻ5��<����[g]"R��(6�K~�u�)Pf ��s�D����":K�����w��9>�WïoƱ�	���
?�j���.e��w�ʡ�'�ry��m�D��ݷb;h7��t ��܆��p�m5��"5$�o�4I�X���)�~� ��ztJv>a�t�?���!��ﵲ��o��5��Spx<�9Z_D�i�,"���j+o��h"b=�z���'�V_B�'�H��@�b��C�%���|vȔ�t�	�8�ҁs#}�1F�¤d�Y�m=u�̭��jZ��O��d�nk��=����P�d��{�5���� ��;��3+��߰q�?�(?����,�n	~<���\��q����g��q|��coF8pP�SX�я�+������qw�Y���"�8��k1���g�r���/Tm1�	�2lo�e�'�wPB# &�t&��Ǔ�d�5H�	t@ئ����m�O�N�^c�M��}�����gDo����v�1�[�8��^�
6�n!?��;5��zp7.j3n{R�[����=�<H�z��<#lifP�Vg?a��$�T�Ǖ��0m��i�*Ǫ�K��xh�~�;���4^�\{��v~�¶�L���0󱔪ق��p���^k��t����.p. ~tT��BDq�#����J6G���rǪ�#���@�x�:{��7!	�rE6Ph���������h��(C]���^_Z�`�K�r$��p��+�^���5��
N�[03�!s�r#�`�*={68��1���{�A�u�8�+.T�+7TE��q󺛢����^��o�*_Y� W�PSR99[e[����\�^M�߿N2���L��Q�-�&�p��g�"DZqsOgՇV ^m�|0�R:���Rװ����Sp�f����	��'\L�9:�`v9 3vwv��If�P��m��U�\6�c3S/:�Z�EF�q�|s��dwd��*Pfw�{F��Ri�|�G�&x�ֽ�Lv*��mz��C��6��j.�qC��[�� -�������(@�FFQ���xy��A)C��ƣ����-�pi`�(�p�D6�y���^H4w�\Y�([���pd�$�#4|-���C-�ӗ�g1��+u?����R����p܈=�ع#�U}�b�W��^\���Vˣ�v
�QKp�r�w���1KނD�;���nFSH�b箸Cm`�Xf��Et����]"|8���� v��s��p��8�͘�)5H�Q�g0:/�놚Q�e�7e~���6Nj��U����Y��Fh��f5h�M�gz�v�`�ƐY^��t���;��=f���3�8Ct�`J#0cc�嵤:��Ij�aVyof�����E�2U��#��ŧh	���մ�d���ڹ�?�_?i}�>}c�[�(L�G�@9ڎ}aꆋJ�[�Ȉ��-[|��0��֬Vj��Tyl�@�z�D����9�W 1n���k�7���wUh�%�!Lۨ$kA��P��`�j��������&9d��\kLˋi��4���2	W��9����N���|��+[m =���������6�qB��p��' �Nb\*"W�PC�����3v�,��ղ�ڑ�z�~��J�C��S@M��#8p��+���T<Nۈ�xz��,�q�zy��6G<#z!ת	'�=�T��`�xd2��Z0],�7� ���RI�C,�'��(�|dL
��D�LOϡV��rwq�3�v%�
�3/R��j����Wb|6"���Ѽ��P���j��b�wꩡ1&ZT�����l�`�q
tw���w��1}\�2�WE�K;��t���Rf���P3��:���@7Mt��-aG�C2�~>�y�Zڒ& ��'���y�|��&�|D�j�\���e�����Q�!9���ݹ����؝�\���)��[����V�H�?����T	�Q��*�4NڙV�(l�$����Ǡ_��A�35����eɡ���0�W�m�|�
c&����gD���.AW.Z]��Ê4������W�+'�o�����i�#/��S��oĆ'�?}��j�d��Jd��"ۅ@g������<�ex���啈�����8�7�ꥒ,l��i��b[��l��[���l�[�R���"l�܍Q]��0��&׃���q_�3(�E��@���y���[o��t�Q�5�T�M�z�n|kQ�[���P#�* N`�2-�7��l�T,�2�#�!���o�	�G|��̭������ ��3�o`���I��Z�X��	����7�@7���
H�1��p]�By�I�;D�?TH��f�]<��JX���b�l����b��DmH�[Rf":T����-ro�;2���{W/�s!`�Ơn>MU��e�to{�$�&i\���؀�5���I����BrX[=�<��9v��#�!�������M %`�/�X*�B`܌VT͕��v�cS	ƙ����$������_��� MX�&����[���}/�=y��n�OJ[͝	
���R�>��P��q�#~��h��??������>g-�$'t��&m�B���z�D|v�X�������dl��(ey!2��D�}��Oo	��g��`\Q-�H�]��~t$Br�Fgߐ륊�ytl�X"�&��t�U�PYH=6DQ��m� �g
[n_
�]%�2}f>畷��g`$�'-�n_�)��8	A�bd�u�'�D��<�:��@���oπ)j4�HŌ¶2�|. ^'���U���g
��@��O��6�t�|����k�����t>
�p�����_$|�Gx�V��^^YA�R��ѓ���p���d��=Wz��X��~,��kNf��ה�V'cvo$2r����?�Q�A��"=G�$@"���|l��x�O�Oa�nߌ��?B��J��J�T`��� >9U�E�]a͸�e�ϡ(@�><rrHYZ�A�61d5n�j����5�ts��WQ�i����tB�n	��9�ߜ�'��������aa��Kž�O�f�}���M(m��GJ��g��z�U.������niUn*C}o׹�n�Tブ��{rZ�g�*����J�l�ܮ ˔��,�`/�� �2��B�"L�>u�tf�_�@����Q#�Ø�l9%���.�O�����޵Yƾ$��&%����4PB��Z+&�7�l6w#R|�ݴ a`�%��i�NL��ãO���z���q;2�� ��������mw(~!�1�>�%A+����f�J|��I��r�8َ��'��P�mj:~�Z� D]���\ � ��U�ͧ(H��N�>���³����"r ��,�O�$۔f,!ªQ9h!Jϰ�K-�k5d'�������X�쎊Q���:�4�M���_��
��A����]��Ι�?�,(c����<e���ԏ�_���|"cs�B��(�IxH�m=bn�&���:S�S�m�<|L��aV�&({�=ۧ�ݮ?�1�`��SZ�H��C�v.�!��TF��5܀t���&�TN�\��C�k�="�� �o_�4
���3�DF�G�;k9� n�Ƕ��\�9AT�����O�K���XB�]�N�M���1D��BDF�9�*KR�D�a��!T]N�Q���M�	&arb�w0�%�����xQ�a:�y�/8٠��11n��Np����tB�t����P��z�4���LV>��l?B5N����Kx�q��v�~Ү�;(�bM^��wV�x�e��I$��r��1�%���'
�ܗyL�B�/���n�)g0�(2�$�����)2�L���a����k���L�v3�VC��.��9s��"��2��"о1�T��e,$H�<�6�>�v�G0ųTf�=�z֬�odftK�[dӒ�X��\MU�!ռ熍@~�T!�z�����~�s0�6M`�b(�Z|byΜR�l��۳x�E4$MbþhUl~r�$�f�=�����>�d��Q*�b�P�&��Q��I���6F�����d�{_9��!�
!�a.����Ֆ�Q�WI1�p���V�{�0���j�Ҙ�aXKfF�y��fJz�ؒr
�g�0�ǿ�O^���%e�`^������ғyXηLH����JD� �R)�|z�3�7���GX/���,��}f�),-`[�O:��t�}p� ��B(>� O�S��&N�v;w���y�d`����ё�h�s��ȫ�h�� ��@6Q�gϑ����}AӤQ��exO>(|�������� �:>����ɦ'Q/���z�.�㋅�D�/y�4Y�!pm��k���_�Q�5�@�U�JԢ�8G+��T��\�%�ɿS�{r�тFK�N�
��'�I᪐K^Jm�#	X�;S0M��y�~�1�2������r�[��<B0d�|l��ҋ���$!�C�b7��Z|��p�wCN���s���^h;&#�n�ce�^���;��ݮ�����~Ё���O���V֑�-�o(�q#:ز��h�g%�O��I�]__�4�_���e��r��$C���GN^R��̠F='b�O�i��}B�2�/���/Bj���1���7*�V�.�r�)p���Rq�!��6����mI�����`O\�K��m���z�M%a9�1!��&��j��a`�+$��(�yӑ���NY�����oclE����������o(�#?�����uhJ�b�L��SC��J�Nq��o�$�zT�FEx��Y��W������}��&��Bd�2��ǎ�]1a��n�9�Pz�YtS"���Y�l^X���̔-��9��(���^�ש�n��sɦ&*�N��*�^�\�X"}�"�uT���G.��6.	�7'�J�D���~���	����:�|�y5�I�C�Sp��,x8�h����u+�Iv��M ����ECܘui|�W)奚�s%��ȹܱ�lϠ5�y���6	����G���"�ڧ���8Vp��D������1��`������Ćy���)i��(�_gJ��r����޵�d�cp;�*���28ɂ�\6��I'x���Q�gEJ�)�(	Xm&X�t�,�C]1��-�0�|��$�(I�a�`�_I}���i�����" X�3r�=�g�C*��z�p�C���q����p��=��h�����VlHVhZ�D��{� x4r�����L���FQ� ���	(5�9���bxr��\��M�.�t���
n�u>���D�h����%0
[��Z��&ݠ�Q3���*)�'��T�_c�-�n
�h8l�Ȭ�6ƫ@�wej9�����qS$6�F��b�0��)����T��������H��^�:�?�-PS��5]�scf&��h�CQ��S��5+�0���vHj��p�V���/��:3�_��5���ԛ%�~$Bk��6}uȨ���V���L\;I=8�Նr�H�b(����Ck]����a3 �5q�p-f˩E�d+�T'sT����%��Mbѭ]U�8������N��۱xܿ�����m�;�'�L}�b$p�&-��4c���W?��C��?2~*� Z,�8!sa �9���m�P���*�o	�VT.D;��
_�Q�ۖ�4Ba�M�$\>F�t���*�2_�.�0�[< 2ξ#`���T͢E{c�Oa4�j��������5����j{t�8���$Ck��Y�Q� ��w��iA��O�AU�S��z�2��N2�+@��e��D``���|}�/H;��<�	�<���xd�}|�1(�����mO�Aٖ�w��O�<���&@��o�9�_R��a�"8Î?��qߤ:.z��4~���ᛁ���bah����@%�:�|�ꨡȖ���/B#`���k�ĽB,�P5BPg�4w�l����X��ܿ��1�>|P��+\a��%������2uG��ڣ�����������W��i���@^IWZ���*�kN,s� 3:Ѧ"L[�X5r�N��ǝq��TA�d�u��4�উ��)X�6f���{~��1��2H��/8A(r�q&P7lX&I-.6.�V2yo�N}��q@@����~�k옋51<��m��ԉ�8^Z<�/���:��Ai����l�5eZ)�F��ڏU�K#$�Q�S|�sNJڧ�4����5:��+��c�3yb�/�]�c���)��B�� ���h�T�Bk=ViKF&��2��}�0�ʚ�&I�J3bQ:�+��q���ɹ���@�I�R6���9Ý)ͫR'�q!��Z,��K ��7�!Og�9tB��N�������U����p�k�.L�(H�"����nW�%�<?�PKu�og,�HF�^Y�F�M�y����n�p�JP��Oc\q�:������V�5�^R���Pm���.���=���֚��������~�~3��	�Oj+d�]��d����O���2vK�J��nj��������Yԉ_�u_����c�˫~pR>�-8N���PLj��	^c�)-��[�4���y=���k|&���Z�L����g��ٓPyYh�{�rn��+q�-IT
�*:���"���%󙨮*�Z#s~���6N�O�d4;��qN9�Z�i�6���R����"�
Z�*!�7I!��Kh��-��&h�v�,,r'�@�Y��Ne42�z����5ݙ���c�e�7��5�h�G&Ö�ݶ(�mUz�I�_�A�-���!Y��d=���1?Y�[��f))���s��ɸ��ɉ�i�E��bd��K)�?F7N0vD��0��R�qO��q�w~*f�4�I+���J+w>Mr>��8�z*���^�{~b\l�׻����[�����d�n8�<r�ݹ2�q�*��b�W}V��ГE�s��a�X���NV� �O&{��#F�o�(��Ӝ�O�{������q�f$�F��]�6�F��uL��Ft^ /��{��>�?�jq~��Fas��9p�=�v��\�����g􇫇<�T�g������Y�����"a7
��2���v�'���n��W	�����A:�r�-u�}�mP�avZf(g-��_{��n���V�8΄���$���H��0C��Ee���������CSG��v��CmO�Fa��ñ~�r���k��C_�տ����E�ю���W`�HV�����I?��ٸF��ʴ�����|x��Ǔ��p3���*�]�v���ܳ�CGk�7�gN嫊�:P���`d7�� ���v�Y�W��,(��nO�'֓��M��ĝ<{�$�s8�o���Jڧ���եgf#�~�s��@ʩS��;:���_�"�`%Aj\}�,��Ӗ
����Et.�?y�AZ�)z@و�n�w>����+��̡xʮ5����&D���տ��b�d;� �&bEw�$��%�	�Xo�K=7p��-8�p�m��.����f�C%��\�VΧr��\��NZ��y�!S�w�Y�%ɪeQ!6Y��^��@`��F�pc6�~�o���Z�aKH�S��l;�	XnMP�Bc�-׸Nm]Y|���a 	/K<UB^�_ ��k�;��r�O�Küs^��Ĳ�dײ�a���$�,I�p�Iv�Y��~'a�ɾ�|�G��9u/k�  �n�. �L�RV��,��=L!���E7�+�\A��X��-����������xE)?"�iR΋�!���6��ϣ��͘�Ag��4nz�p�"O�C����

Ӯ� �$�]�UM�$*-[~�]�	�1�� ��X���CM��CTV��a�^D��/�i�e9���
���ื�!��۰Ol����U� ܋̝�o�v"hR2J9�ǿ�$��f|)B :+NIVY��)D�ݡ�٦?��C�k$2�9�z������}HЩ���9�s(U҂��;�'ٛ����_�`��R:�̀hThJ�D� �Z�2K��G�f��3���5Q��^��.T�����.�� %Q�A�t5Z�:H�V!V356H�l��b�-\j�p�2���iCJ�n�c?��c�q�xL��2�ߝLlg�3���#B�;���F��W���`����پxο֠�ڏ������OLԎ�o�*�}�CZa1���/��:�f��%�w��33>�F2o���1;�Z�|!.iI�I���@������q�bË8hä&k<Z�����{"��#v��R�մF:A�H��|?���o��I���|2�w�H)(�OIO�j�����˽u\��L"7l��zND��3��*w`lJ# �$���.��N�v愤�Qλ��Lg:��6ՅwZ��X��p��h��������h�^��|-�fs���<Mj���������Bj�"����(�h�ܿ@�V>�q� �5����A����!�-5���>~Y�s�!����ؘ����V�&YG|������T��?�l���'9�|;�ش��:Ma�7O����S�
�ؠ|P�����A�}cX����v���A�g&������a	|�/jum�k�-=k�{���b�+5u�!K6����;oܑ��G�K�q�̏��nT�'�.-���� #����K��f�Q����M	���?��k�N�Q���{LC����|2#��zJ]����\����h[��֖��q�W�SϵG �`�r�&(�-ZN/m|�ب>2�\���<��%jP)��~�=Hk�����F�4�#7��s������L{�􀼅<ד,��T��I�,4��p(W�33��_ߘ�v�b�����E���s�Yz~O���n��0k�������v�L���Mw5v!۩��#Is=��ɧ[s��A�/��.�%:֞�S�	�s+�nA���.�5%B���xϩ�F/H0��,��hL8!9&�8�Ů�=s�,�Jy�fZa�g��!LI�I���Y��DD8�����p�אa�:����6�cg�8�0�\!Rk�+vn����
 �=[�=-����5 �D��4�#�!�%������^� 'hlހ�2��<�o5��+2��cl�qa��1a@3`q���2�u2�2x����K�
�y���ѕt>"Ҳ��j)QV�)��"D��3��(�����<����&���ElY,��g<���Ōx��8�Ͽ"ԁZ���a7 'n�A��14�ߒaPCGđ�������0����yT�'�W۳�ڿ`�Ag�9����%���z}�]�"��[X����@�����R��Q8�%�[��W@��!A(�[Rم8�5%�?��� ��J�d�%0��UvDǚ�`D�F�����h��͆�~B[w�l,�r��q�tT�h�`m(���YX�H���:����ϸ���ͺ�I���X*�� �Kb^s�J�c߿���޺	�PW^j��n�<f:=�s��^��>O܍�
�GsW���NZ�u�^<�����x�bn�R��in��1V�g�];�x�:^d�S;�-�-�dJ�ݜ�p^�j��TIc��T����T��0 (���sш	/�6���Q�y� ��GS	��}��J�eI#xoҲ���P�$5Q=myG#.s��e
�EC��*�h�o�|��O��!Fn��%�A$܎�|���M�X�{�$��Cb�B�7�FC̹�_�9y��hF�?3/����-��������#�4��㰙�� ŏ_��6�%Y�U�j[��ӟ���Yu90B��D��S�l�-QfA��f��W��,�~�ng��L�� ;�`_1�R�]��g;��ԗg�1-�U���N<���j'����t��4ӛ�>�$y�ڭ֤��~�v��/����%zC[�I��M}�d�a�	�%xC���B�}�=�� �ҺfʎӬ��tt�U�ıI7ӱ�)}�E�-y�{*�;�6��Q�{-ު�~�m�k�ݣ�4��^�QUJ��iMt���	�g���3��?���D)�ܫS�}�����,�~�˃:�a���?ʁ�F�kF�඲^�A^��DV`�X�vdv+���ᢷe����e��?��Do��ȉ��@�6�FR&@RQ�D���Ҥf�T��P4 �
�3�Ȥbc�&ӭ���$
���aL
��h��UZ]�G��&�8wa'5�pi�@��Usx�s�	��A-���F���<V�$��xs!�{��(�?�����@��Ƿ?�s�O�}.T�ǆ�՞Za^�O�7��'#���~��2�O�E���2k�����9dS��a���.�0�iP��@�2�d�đ�@�������&J���2E�X9y%&��Z�2o&��"�$�s�`�O�u��ʎFGS2	n��-��z�~'w2� �M(�>��֠�م �7#��e���?�AC1-n����ٗ=?գk*���Z'�Wu�iĸ!uT���B�Zb��7�om���KT��3�.���#ș�J�/ �,٭��a�0$���n��ҵF�<ݝ��}��HQ������y(<�ఔ#�/�9~1���z=B������AJ�ή���ܽAs���urxߙy���J���0W�P�Y���Z��ڬ^��O��7@Ii��Ƥ?�$oG����!���u�^r�������t� $z?�d�I�q�c�''��-���$�{-���DP�.U'�;,*�9�ʙ�5�`�QX���+]�H4��bۘ���n�q#����vZ���s��/�[�|/pk̿r��ưC���L����-�����~��,hK���b���I#ko�C���M��C�K���j�:�|{�:a�(�G�(�)C�6^���r
��ђ�T���=�ulhӜ���N���I����Q�J��^��UV�����Z`��÷q���p�� Hߓ��ؠ~�҅��HK���v"e�0���d����yenl�bW�;|��#e&1e2��u�e�]-	'�I���d�FJ�S4�[B��2A�e�^�d�GZ��/E�T�
{���KF��7g���c�{f�RZ�Ԇ���݈rxZҘ-Y2髗
��9A�@.����[p�_a��&�?�p,)\#�����v�w��>��Kf�}�����ղ���!�I,'œ�ܱ�駼Rm�$�W��~W_��h�#�>����g��+�������;�G��.��T*�A0����s���^��ӯ0��I�T�J�
�l�n�]	��"I4��0]b�Z3��Ҡ�T��s�oq�F��{�ՄqաR��]`
꒷�=�u�6�4v?�+CNd����qj4q�d��M��S���E�)\)������4�t�ɭ�ȏ��^/�|����$���CY�g�H��|[P��ϐ�²���eYzz8�$0����A�w�� ���J��̽���6Zw:	tr�SD�}8��NG3���%�8�tF�k\�pb7��ɖ�3�m�a�2��4c�L�7X\����'����JUW���M�5��u"��u�V��O:�ˣ�5L�.�4
��07\�]b�-�����ʾѢH�h�k�FE���Lj1�7��[|������#i>�5�)��7A�� Ta�)uA��\hB���e0�I����+�f5|�p���(f߰�ħ�F���>�Cҁ����\#��r�Ӑ��������c���#��b��M>��.&|
��k0��۽�=��'y���`g�o7O9l�zT��0:#��:�!3�J5���?�>�$
%km�������X?ʠ0���i.��"��;&~w�i���=<������n8rQ�-�}
C���(I��������Q\<s͊B���sr���$)�Hd�c�K�#��D�b0n�(Qww�0H<U�Ϟ`g=t��![�5\Ia��� 5����,���С���<k��U�o�C�}W��{�����Qm(�h���Ҏo�����т��l��#�:�.��6�u*%[㩇�d�mGWHT��������q,�\n(��1`�ɂO E�1���@���b�Ka��G��F���&��C�����IY�;ӳ��@r�Kf��4$J�u�z:e��j��H]Xl��}R��ե�[�@D��S��U+���7�JA�Z��ʾ7XM�����)���`Os��b�΂�a'�w�l�=��_;˝S��=il�j��	���`��j�n%I�}��*�|�N��	W����Ŷz�-����M��>�P�R����t(��5�4��}�� �!/(w<�����5�m�i�$~7��\~���z��5�-s3����/�o]�#�荃�o�j��~���J̐��/cQٓ��5��>�XlN�cb��8T�O�xnV�-�t��怷ѵq7�v
n��%w�w��F�M��6o3�����¦�|�o���Y���h�	j@��	���j�-cF7(#�����N�SL;K�{�i���V����8̏/�گ�p�Aj��F�y3����/'�,Uh��/����}
2`��i7�Ϭ������.���7e&��5h���U�]P�F���dO;��u��B�uV���u:
�.��Q���kO�e�:������ ��H�������a�lW���L!V!��m��ڀ�Fl�K��'Z�����#�:>��K�����(��O�!WG��eZ�okQ��,�]���8�Ϡ��ŧa�7�@�!1�%����\-�5�f��a��V��W.�L������c��2��J�֌[t'��i�R3���sץ����3cZ��ش�V�D��������П��ԧN���!ۖXW4�c�m�7�����/5�S��݅ј_[�v�[������!����@�~^0��O (�L��:����om�3'����E� ��g7l���/����4��U5�T�l�i�d��9"��
�q�W);��p�X����[�m>M�U��{9Ln�V�~��^Qb���d�J�����M����Tiw��X��̰ҳ%A��']R�I�jghG���l��\�����g�M���J�� S�󇟣{B��e,nvn�Bp	�z �c?��(���Vu��Y�x���1�"��#�!�x�Z��ȶ9��_?�%a
J�p4Vo+��[������s�c�ռ��AA�Ć�@�{ۂާ�a*G �U`��5��#�����_�E�9l�Ti��%&ҵJpVk�w�i�Br��'�ٗ�6QxX�-/�`f���	�Cۻ;����q�~��X�k�F9��pX��������e?�2�scU|�;�n����� ���l�k�&o~����
�����P�]V�d��nC����e�9���ے;:�e)T=&@��I���nm���^����2`��~�Ү"��8�7���ʃ����&�H���U���!�}��Ńg���~����Ai��z��\>vXDpc���~N�Ԡ##��Ut����Xx��䰉P�����f�S���b����,/���~_~:��m�(L���:��`��L�ew�+��)�f4�P{@B+�Rp�$h��2qC~�,��,§�� Τ��7v�_u�MB�9�G�7˂�m��B͙t�9�jc��?!�a��h"���ih���@@�*py|?3��yTi�H���Z�\�i>��k���[�	��.�Jw��*wd||�YӇn!�$����_g�~�t����ԕʞ�?�0~2yS����|�'�������qa;P�VO'�Vzs�g����`ߝh�V/�����J��Xef1��EkO)�cH��z��H�M��]��i�گh��ql,��o�t��ʉ9��R��Qb�j��i��O�_�\5��Q!�P�Go���-Lk���K�
�zC"�j8��f'gg���!כ�7��i��k��9�-��1j]6��S�Q��?������B	���O��R�ӛ�o�<� 5�_*�:f��KKK��v\���?��	xz9�꥗E�����Feb�.'H_������]�N?�8\rQo����p���nwZ&:3�U�q���d��d��U���g����.q��BX�����p{�&8��o@
`vڨ*����X�6y��N�FF\B:L�ME"6�x���l|�[�5_c