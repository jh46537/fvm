��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p����A�Ȫ�o����jW�-�#"Kn��
<�;Y�p;Pk*)�y�ZxD;i%`�(�N9i3�A�ae ��������>gŎ�ò0�*a�t(�;��r���Yj]-ҕ��ո�W���]K�~��b=��	n5���EЗ�9��iF���K�sUa�D�c��'��@}S�W�a������e�(����8�|[���-���M�\��x�,���>K����v����)b<Z�HA���7�CAъ���lhl���6u�)-}�ć�xZF���!΀��Ss���8�`�)�wX��q��A���O�:4?��v�X*���'��܂[P��Tm��� g��R=��`Af}f���hPe5��k��H��o���;E��2�!��W��Π�ԝ"w��n8�rV�k��]�g$�����j���}M�pJu����k����gf�K�(Ю#���w\8����W��c�{3���,��_jO�m��>��wq4���+��u9�{M�-�EN~K+�<�K�&��ũ^��,�o�54Ma籺Wp��[n������+��ݹ�)��7�sһAV�K�S_U�B�*�g�sj�Y�FF
�X�~���KF�,����|Q�'�A�X�F��?	[y_ HYil�
��t�
��٠��:�F���t��L|7tH�F2f�Z��G'<��j:�]W�����x].[N��$��ڤ$wf��ܰ[�~�������vj�G�@�k�����H�#���%W^
mQx �G�v�ۍ!�D��78�w�6����?��>�BҜ�<���RŦ�G"^Ŋ)N|�qcgEt�o�����m��3��XSI,E��զy��QW�8G��:p�d���^�[ZX+��p}���I��їc��N�~k%�m�c��
����J���M����,Q���ig�/oc|v�=�vm��/p���|+ET�e���j���8�&s���Y;`��ܢ�����ƭjᔗ�rt���Ϡ�#D������a�@�ӟ�[}���W㜻|����:�ճ�R��w��FH"�%�Q8͈M���{u��ŕ�	��K�G૯���̏$�=��b�Q}]�=�'�n�ad�����h(k�	_���X�ZE�hέP�e�fE�ܸ7��H��Q^(Hxy�}@�L���������i�Ne'�Í5�Җ�N!S�m�/HfA�<��r�
"��3� ��,��J �N��[�r')����!��X�ڛ��NNOZ�A�Zvr[�۹6�$��\���X��,[����>�y����B{�
A��h�����d!$��L�<���X8�q��G�d��YN*޽�sY���4�G�a���I�D̯���sfK~�1ib�tL��\�[:��lz���P��qal�I�z~@����J]_cm����b��7��)�C�t1b_�PF�&(�����Sw�sn�)�Π��"���hrʵI e��i]!�X?��Ѽ���t�<ͮ������M��r�I�g!f☽��������/$Mg��>�[�C�t��>����V�OO]���d�ai?w����������R�+!L}�e!m'��)���'�#�L�֗���5���/��w�d����c|W���h9�CN�������WZ�����*�i'�G����%N�۠�z��X��Ճ�Z���F��˒�-۰���q��E;6�A��@=���!4o�R%�te�g�YBx論�Ɍ�����Z��	y�M�m����IMV��}���6f�H�<3�^�~-��>��UikA�����d�Y�������@��@���������-�K?	OaͧEi��H�}*�R�Qf0jw�Gn�H������E��O�]Js�yS�+���&��Ԑ?�ۡ�׾m���<��:m��d��e�"l��>�R���&�`���7wu�7*K���uNc�W�Ə(X{^�N�{ktw����%g�8&�8�ђ����6��=O^��~�*����e�R �+ԍ ]���SX�����x���	(!���ThhD�(PU���5_!���In������|�k�d3M�J�z�9�Pjb(���e���_vuۄ���+�П��Tpx���5���xK�
����2����G��*h��H)��q���y�U/>����"ݜx�%���UΙ��*my���K�����Z5d�A��D�o�ϗ�����*�?�J�y�|� M��Ip��.�r�gH�ĳ��9�o��p����s�3[q���-d��U���_ч���i#����VQ��M�ЅI�E�Lx�9��: �yW���;P_�2�B]Q�h�9n�ѤJ>�*�d��ǟ&�B�=_)��
<J:��W&>.8���<n�a�(w*FÌ=p�)����v=ø�TQ��^�1@s�T�pxO��LrPr6����@IJl"���4R_>�.��ȥ�h�ހZ��~ɚ��:zs�D����Z@j��w� �-jmO�u<)�J�aU���l�Ӵ࣪�1�_f���#�͆6����)�%����֍��O@���+f�[��ЭN� 7�,+q�}�x�������}m�D�ֺ4P�_��D:�A��/��t���t�$P�Y	IS;�2�TMߠ�3��(go�&H�4 ���%��U#Boɿg�P����7 tbJ�̒V �ߦ��!�k01�	WT��Y��$����Q�����"