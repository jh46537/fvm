��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�0�w׍��SΪ]�����E��>��顗���="�Ct�QJW�����j��I�����1��5\W�(���\�D[��u��=R�1����9��f�\:���e�zm��Y,J��'X�බ,|_�"��?H�L�"�]�!.�'�:l�y6q��`液�KP��W�uc"�@o�vs��K����z�{���)N6�!E������).	��YЋ�i�;�c���7??�vа
3%5�E�k��#�o�$�d�+a~�e�$=�H{�h��-v+���x�9��s��M�󊶪�B��W$2zF��Ԕ&d}rD��DD��'��&W+)K��pF=e��p��ձ}u6���<ψ�����8�_���9�U.�9�;�#h.'��@�4T�.�|'��<cRz�fڴ����Y5Ǩ�H�T!�Wrj�=q��C��w�G��5w(��GF����XG������O��s����Ǭ<��*>'��T����;0~��b}˓.�)~�~�t��F&�P�8}ѓ.rd�p7����I��$��;8*��t%f�Xӏ�5�zT` ��oHaF2�.��]xCȵ6#��H`��(r1�ޡs�0X9�u�C&O�\EOʥ-%/U:�g]w4c�F6-�z��h�����K��>�3<��wH��)j�l��5�u�)� ��rŞ�G��wLͿ.���`���9�)���(f��R���8̗�����K(mj�)�r���W���<�I��띘B��RU�o�f�I�w��w�a�ւ6?�G��(m�,^x�~o#3�)HBV�Y��&�j��#q��
�L`Zcn���}J�v��⣃���h�i�	��Q<���S��,���15L�e�(����%�KZ�����K:S{�Z��KO�\?��sg�_5�瑹"K�)+�MP�yi��q�������:�6��7`�	3M��ޥ�yw3�D�yX�P����PR�2'��w��[O���}}�_�� e�ig�2�ߛVY ���Z�ee�&�x���~U-Ջ5\�4�)3��lP���Ԋ�(sn�*O㗉�`��t��q����;���w���>WV;~^����Ka�ǃK��[�؄o�̩/<S@�t0=����'ꚸZf�>�6�-�xV	������c��g���-�.Ț//�V4��w��̻�����"C\���?�P�Rn�|z�l.����5�X�K��z4�@���lrt26+�H�������Sz�i踴I��k~���2�5�����"��ΐ��;d��^:��EХ�slŠ��BU#Bl
��Q�/XbعPa�'�A�����G[U��,�%-�-D��P1s%�)�q��G��B���%����<_�!�u�|/~�i�vv������ӣ*J.;�A�1:K;�,�Kd�oQah����>�k���=�s�V�v|[ן�$$�U,u�0��I��MR�2�����l�51�I_G6�f&��yٹ�.c�]�\_R�3#�����\m��&�$�5�q�Q	//0(�$)3Mr��i^���������4;��~��@�RZ	��MDC1|Y���+�:xprR
8�k�sߊ�ne���TCr9�K9�z��ح�Xi%?��.�@��G�Mݦsk��s)KAx]�����'<ł��=SD����P�~u�Z���~��S�dG��]_b�ӻ
D,����^�:ju��v	�2�=w����[u�_`t��F��:�?�<|����uJ[e��KB�G >��{L�X����f�\���I�'�n�8Mo櫩���Fd-C��Jo>gcj��`\�ϧ{�g4�����p�&�Q��;\ߩx���{���挟N��8Z���C(�~Ud�&�5F����(׭<#)�y�U�{����*T�.g|~^x�:))�dݶ��*ů}>�F���So�0�e��+ݕ�)�$�T�In0�z��4��g�K����̑2��k;4R#�o�r"�)O�|�M���Գ%�~�����Κ>J	{�^h�yŞ$m��)Y��<f��c#%�#1�IcΦ���A�k^f���������w3#�mVJ�eOÃ�ɬ.w��x�N�s[���A6����~��|�U�EZu�_Ï��g���D:�B��k�D�&���i���܎Á�G_O��4B�<Ae0��q���+9�q͛�Z�����<��_/ߏC��y��Φ����E`�F�6"���gHf��ݦg^�����y���S��̳���A��f/���y���<Q;n���E���S HS-��m VF�}`8U�3h���):��1�qB]¥�[�����F�,+w�gZ|\r�m��E���#~����֬�Vي���	Z�dg:{(pҾ�S"+�'�R������V"��}r��O�����M�k�#��(�5Yd�T�?Z-۹8-/�ѝo���*�-\_j�b�lu�hs��z(��a��)���u�;�As�4�s�&y	lH��ͩ}��.w}�偽wa���gu��r�]���4��
v~���b