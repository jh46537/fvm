��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""½�c��ノ�!]&P{9v#ɋ*�j���-=������$W�yGy%�DL ����b�Y4/WD(���d5빂��P_�afRw<�l�HO�.���D"�f?0*��%�Tϼ\	����Eiq�92�"�3�FW��jx��{��l���~�H��nA½��b4�x�Y�V1p���%4v��_���6"ߺ��ɨ���ſ�R�LHͺ˔H�,���w�8d��u_R[��&z�!zȈuG���\�$O�8I�1PRu%��*�UN[AL�0���yn �QS���L�T/��A�����W��z�p�����DP� ���(�����)�4�>��=�@k4�k�A�%VQE��q�}��(]��u	�/�H:cI���-���2�>;��[� b8�Ru�����j����G��R�:�h=<O��@�����Fͺѐ����E��P=���u�5w)�a��A[�b�e�>-Y��p�)F��T�u짮-�A��t~����l7�QG�q�	���t(m�Smr�At��7�zv�L6��� hd8-��P8Py��r� ��V4���\9"��Q)24F�"f,H\�u�N�C�l�C!cF	�8+}p����Kw���3��1�ԃ1oP�\\��g�_�k�|f��h����@s�ފe���)���ؑ?�a9��e��?^�-V�9��XY������-�R�b,�9v�'���H ��Mv��`i�s��׻j��nq�ߢ�Br�jcT�n��8�~�o�l �Q��Қ��u��ϧ��s�Bt7�Fas��Z�k灍ѫ�֋��cV f�|��A����)BԂ)�03s���f��]�,�g�kA�p���Ȼ�/:���!r��
�щy�(F�7v?��Q^=���x)P��\�t�i2g��ncF$���]�qz�R��T<��

e�̑��{m���$�\P���I�t�"�c���C��>���g�������DA�/���:/���ʀ+�7���߶�{ۍ�f�s�o���3�T��w��ڪ��{�8xYg\�ε⃢���2e|ذ�-���z�tqkm�����3Ȑosd;q��;_��:9��m͏/�]D�d��J�]SJ:"�ӵ�t����t��&'xZ+
��w�:اѼh���� �ҐSB���B���{�c��Q����7ps9w��"�8	խ�ٸٺ��3p$��N{0���\q�K�W�oA�a6[u7)N~�pI�4-���r.�b�R��Th=�ұD���N�"@���{(����2����^v�F�E���<?�*��h���Q��	�E9̲��:���4�/�枨%�8�E �u��v����#�Os���4�B.��+0�"d�ͣ�j�����@<#Ւ��?g�:a��1�EUo��@��oKn���g�s��V�-���0��/J�gϵrY�o�d!�d�w���n���]����Oz��y�} �Tl}$���d����	���ch�ŏ�$Q�[���ٻZ�&lv�Ώ�-��˓?[zq�� ��"`��R�8���Я@����g4M�՗��=ܝ����#�J
[]������p�v��H} a১��hK0��Mn�埄�p�3����"����I(�<\.�:p�t6L;�w�W5Bn��?��lZ�N�nn�g�@nx�����6��/�5]N4G��W:�$�9O�e�G���4��Ji�>��K�ze��
!�iOP&��&m�=CD�N���A�j��\�#ƥ������R"�74���鸸5�#�d�|���J��0����v��1�L:���������G��%T�n�7�zל��9� 
�&ʴl;7��P��z'f[��7{��������>�Y�UƗM�|��h@u�ƒ��=����LT����U�kz��8I�_�=A�(C�\����>y�����w�ğ?Ii�ͳ�l�g�q[$|J�(�zO�xx
(>)l�E��(�g4d9�nO��Y`��n����4���yv��~g	]��9J7q쉴���lT����VP�s�2#E���Q;�C�n�W�m�i��t.�]�$R�2��8iّ�}��J;��q�qH�6����,\1�u�*�{���⬶��jP��]���u���朂����d��/P�R�N�c���T�׌��I¥�T��Ҁ���pW�vͥ�P���md����E0���B�f�~��kʎg�V�AZN#��YSM6\&��zW���]r/,���AKX���/mV��]��8�~�/~����ɧ�:��!z-ر��7L�! �O7��:�ӎ�JP��[���������hi_d��6X�f��iP�w@W( �����6cx>���0:���J>���MM�Jv�	Dqo��)꒧�?���꤅Gsݘ��V"�4�C,�Ď)6O�ۢi0E�M���0=R�;4�j$�x-"���#`ifD�տ�,uv��璒}#Ϧ�J;�+볢1�TVh�TE�oߪ��l�M������	����_Y���E�n��rs�nO��1��l��(c��0�.+�� %f�ܝ� �1	Ð�g���lt���|�1�~<ʿ�U�-:{�5~�t
�g��W���N�m:[..�"��bS���V�q�r�q��hó�!��.�1��u:qy�G?[D����;D05�{��>����DB�ɜw/�n��H���@��s{�z�U%��G2ͥ���;k]K�i�L_�@�z�-���^W5�� ؜M�C��-������+�V�|\Վ���+�����.St�e��n���)�Oc?
�t��xj/U��*4o���gnwU0���zz��{E���R!�B,@��h���e���M��8A X�KVJ7�g�Z��_�2F��A�@&�T�ą������d��x�5��&����؏,���<�1���7�o>��z
c�'ڟʷ���i\����ǪͿfP|�M�L����bE�N�lѠ64��{�\�K��t���v{������آ 9�6B����#����_"q=m�ӏ�ʭ&�����B��7�T{R�� ����O:�F�}��W�(�eô��U�dU7c�ӪD��@֑� ��g�Q���Z~k��:H����7���<��Y���<����w���y��b뵥��|Z�F�y���Z�(�BA��ɰ�B)�t�(�J�/�+8`��iШ�}�m%	�x��ZH2������.G �6V���i�gʆ��<6sz鶹�����4��qj�(���&�_f~��_�!����ՠs�)��?��iy�[<[l�� )��z1���A>�ۖk"Ҝ�5i6%�%.� �#2)�KĤV����|J��aQ�~7���3l��Ř�2���I�yh%���O'�j��N�̷! �� �����ep�q�_�Z�[���ō��	����j�	͟q�L#��l��ZR��E�԰�G����DĄ��,Yj��+¨q;���x���ABLݶ��$���?�����''�q�͉n#=x?��㽞acib!$ dDGe�
���c�f��?�/ ����K.��o��:����2�� F�9�[OxH���� ҍN��*�cv��v�����2\w
�F;���U\i�1/�K��4W[��B��ڇ�n`��K�1������d�s/�@i�\0�eL�pu�������L����q��Y�-�C]�y5�ttsz21#ȱۗ�u�o��D���vwb+�Ѷ�W,��s����MKKt�yAA���;�Z�42$���^C4�fΚ�Ì��ﮮg4zV���%6������X�����5�؞ȹ����>^8Sˮ�z�c���X;��P���Ɔ��̢��G����]�`J�o�#A�N��\���X��_�H���J�
G��,�c�44N����躑�ڣ@�i�ŹI�<��s���`��)|��\�����V	�� Zyj��{0�g��C��k�=�(:6�>t�4(/�cXfG�"���(�(B�w�
NH0 3#�9��T��>�O>���	���SuUN� ����Y�T���E�<Cߚ6�JwM�/S����g}��,j�m�,���6\H�$\�Dۈr6�`�Zw ������w^=s��G�Z���Bz:T�&Y���3�W���hӶ����|�j�s�~y
�Gq�_��%����$C�B��KhI��3K}1t�k+�/�W(��s�'5A[�Y������ѦI�;j�Le�߼.،��;$d��%��P3�����З��=	͗mG�'5�_"�Pq����˛���R��XD�9����`�xA�m3��L�8=��P�Sk[�3���<��_ ̃�L�e}(�cS�B(�N�[�uU��9]���!Ɇ��ߊ?g���mr�Է���gY@��SF�fP��в>��u�J���ͫ��iL�)Uhy{8�͌uݬ�kW�L^����3RS�'�v+ ����qg�u*c�Y�W23+�o%a�,�7�1$
6�G�<�C�v��3XB��H��C�r@�1�n������y-���D��4�r��D:_����7D�!�JbE�6��9B�`�x��&C�k�IA���:y��S#{�'!�o|�!o�������?��Y��ejx�[.���pŘ�v�R��xiVm7c=��+Z[z��h��%��uD�T,>���0Fj?Ћ�[��}e�.X{J:ֽ��/= au@p&edQMx��z�-���馸�Ecxmτ�%$6�CFzy4y�E�B�KF�}ݳ��M��0�0�Ӈ ��y��2��W'�Iq����p��l�\�Ɔ�����f@R���T��S�`&����W@�Gr��Xï����5���>;E� �X�!�g�$?�+���ZT���w+��
:(MBIٷq֏�}�ğ�Rs�r�/F�z0L������ ��q��s\=����`;x�Y}O>�F�r^0:Z����}DH��ð�o�XM��m���aR`�SW��q� ��(v0 �^�Į�Gd��m��=�@�D|�l��h�t�Ñ��4*;���+�}:[���n#|�&�̰�f��/l�-~o�rs�ޡ�}ల��N9��˝��ӈ)�����R�
���Y{��xr8�'fW+-��+�ħ$ :�!S��K�L��b�V�QJ)�%F̎�j �ij�*X`��#|P�����S���a��:��J�zg��ٷ���m8����M�C�����g@`�S��K��&�%�W�������|�#���24Qv��_�_+��h��W.��A�?PUs��vO��\(��jSuu!њ��LY�t���@��b�=ֻ����=�d�C����t��ccԚ*U%����6�Fjћ��mYks���������N��,�ȌM]��Z��)m�MkRaLB��7 �T��e1t���b��K	 �<`�;D�!�A;q��84��ܥ�8e�FE!����Ʉ�*�~�׭���
@\$����"�ep8D��Y/rb�y���tY�_C)K�V ��@^R��k/�qN� g���PWa�&M�H���_�"���-R��$�{���ΰ"r��N�i�?tv���!��h�{X�3_�����~N<��S���*X��#f���5��e�����&��P�v9??>�֤k���ZrFY��=����)sI.2�<��Ҹ� 9����PjjF��%�dgeIP�,���eH9�N�M����Z\�$1V�̊��OvU,� X�U�:���H>߄�:�����P� ɗ�,�*�%O���״9�f�=JXC`.���2���/�߶tfy��C�UP��q]��hsM���!��)d��
@<n�ӑy���IyQ��~���bwju�T&�V��Bcdn%��ٕ���Z2,.CbGB�y�S}�y��mk�3�^B&�m���鈂��Ӻ�?��ϋ]�CJ��JL�L��^�q���]��,��(5V��z��\�tADG#����f?�b^\�\��Ae��������p�o�U���*�_:$�n������ƿk?#;�KY�3&��6�Ȑ��'"%��{PUΔujB�r�ա�.��I�V_���jV�o��5��k��5�c��%/�\6B��<��%�
�B$��<�ڳh�A�Ma�����!U�����w��5�ا׏Ծ�^&+wۣ=�A�#���Q�U�A��g��5#�^���^��~3
�0]�%���]}��7v��N�X�\e��Z��?�!�eTu�b��6Q���(�/8{�`�	ɨ��(�.ɜ�u��=`��ε�V��rJ�ZTM��B��jt �2�͝�vmH�"`�x��m�K<Z6��>����^8RQ�o���d*Vkޖ�U�ߥd��t�]�����jȓ�P%W�����Yт��t�4�?�ugٖ\̔���%�~'�?���<γb��Hi�fu_���mr�79��(�DP����op,Ҁ���cǜxi�)�JY'��O �$�d��r��#^lj�e�`J�Ī䲈aL&�>�W�Y<ec��&F�G���R��V��H��ȇ=~��k1\��D���˷����ѩ��&�Ӝ�U��-=�n���Ҏns@���:^9��ˈ��
W欃qG�ҙQ����}���D��8�;�Z@g)x�����3��4e�����%�c(��C��/$�6���h�"B^����X�!SA����#�G��s����.x?�/æ�>��pB\�$�[��KG�����r�h:�v3LǼ����H�)T�� �]�	���L}�<��f�m�.ֱ�X���.�a��$��{�5��UG�>���<3_)��}�P+%.Ԣk��Ӝ"�B7Q	sOyĔ!1C�k���0���}�ҏ�!2"�;���P�X����[�<��y�W�<��o5�!OYI�O`	x�Ÿ��
{����a�cA��l�����_���+A�#3�6�i#�pQ&�ܪ>�]�����"�)���ۿ�V��f�Qw���}"L��V>�(a,�}f
����b��kL�vy~y�a iV���ˎ>������#�&R�ĄD�4v'ī.�[�{��~�^�������x�x͟Z�0'����ƿ���~d.�nT��^v�{K^�a�w�������x���*o_x���� �Y^4v��.靭T�j�qN��@k��wU�U���J�8p-O_Uԥ�|X���� ɯLΊlZ�����Qv�rk�B��x(�U�4o�\?�hm�S�8�}�v�̂�?�?�a�� �s�LM�W'8����{"6�����C
X�����ۭ�Rv˔��އ�W)�&gw��I��(=脗߽��rɭ�>�M����*����zP�u44�e}�Wv�`����4�D�I1�\l�V�!~���:�cFl�@��솧�ӊ��n��C�D���9�?��b��G��K"�MLBu�<�($UN����56�?Pl�2��������e��v���X�&�&j,���j�Ʀ_)A�G(�ֳ]Z^� C`����[���|���&�]��k�)�s��� ��; K�
?���a��\�k�]I�/�I�(��%���v=�p�-�Ye�1/61r�4PX]	���H���c�w�P\�I�>�*�+�&��
�n�%�����
������/]�<�t�t���^�;*�Xȍ�{��D��SH���"�7P.�����v���������������P!�����f����ɸ~�.y��H��!J&�"0�aZB �>����ˣ
HG�R�i[<�2	|�$��j]��`�9eM�z�*^��
]u���"�6��p�L�g?��x^6�i�v7ՇKm]�]�c[�@ʔ�=�=�F�]5r�j9�i�],���j����X�s�H,	
 �\��%Jj����I,1�����4=K�wS{��������0�ͫ��p�19���M0��Kh}�;_a��P/IҺI�%�����hM���<�>������HE��䕱z*byl�tl0�?>3�n�4{��X*缪(����;����l�qrр�#f�ZKk�AK.D��|y���A���w��:$��F���\9�>E�E���:� c�7g5�TE���̸^��<�뽼V	�~�vs������*.�lFکs�����l.n�n��L;���,�/|��i�x��ZM�R�.���A<&�0	L�E uC�2mK�'��֖f��3假�j����^�&ښh:�b����k���j&�������ڶ�C-n V/-洆��&b�n���޾��ӭ_��Ӟ��Y<B�ӏ��W��R�rس}�)�����wn�̛�,�B%\���V`�g����i���}�/E�A$����<�+l�'�X�k%~�_V�<Kp��v��پq0��z���Q.!�tK�7����?�t`#)��2+����V�����-R�@#u�e��]j��5V
����b����b��$\ %�9+�C~t���c:�L`r�^.~��Y�Hk�b�l@1���OH�!��M�h�]�qA��$bP�I�O�!y�+�K		�Y:�s���_^J����NHr>J(�"k�9⥨�D�a^���:�0�ǌ �WG���YS!��Y���
I1JX����J��j˶Z_W��7B&�Z~F�дY�KrG~mk�+Z���gJK��+{t��t6���M�MZ=��>8�U�O/�c=�����>*�D�WByNv�P��Ŕ3�R`�fy��	_�
'Sh����������%֊.�B�$� پ�� w�r�&��b�C��˖���;�>����fDsET�{ag���eTD�LM�c❜����(U��62�1��b���-�v�L����'��-�y]�/T�-8���!����n�˥�v�e[a���!�� S�D���F�����B��5%��|Bݠ֕�
 �պ��BD����̽p�q����98
q3y+�=�+q^�+��K��U��^��Y6��oy�$uC/S�gH�m;h[�S#Nm�3��l��mF�5/�IA�c3�iy�0��TA�"���5n�>��k$�"�	���%��댎�*�f����܂��� �&��卼��(��t��\O�̗*Y�xO3|����r�������M(��#��Y	ޱ�赘�zZ����NK
���;�s��_�8���.�u%e�ܯz�8֨nc9������J5�24�������*O{�Ơ'�G�T�V��3����l�b$���nS�N��U��5�� �Ћ;Ce~�C���A���7�hPݲψ-�p��(9Tx`����G�ǅ�y7�iԣ�]p�g��L�3Bb��7��-�s\}�t�la.' �ᓤ��h6x���+����./�&>��7N@�ӝ�����߽Em[�k�:��~Dі3E�G6w�y3?r����K�����rBO�qJ���!�+>}��r���o��s!�z�*haя-��l��I�|��#�DPr-ŝPMk��}��+�us}�$^!�'��@	s��OB��"tż�	�å�[M5/�} ���l�<�n�)����k�&��˪��\��zU�ڗ�Vs..+�D��<���Ɩ$�jB�Z��gj,�c똒���+eBwf9qneS$Y��)�E�����t%f@m��,^O� ��i|�_z�l��}�S�З��_d��G��3�'�bs�')Z���il��