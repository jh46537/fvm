��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb,� K�3]p?�$5	���Ai�ZѬ��s�J�`=��XO;��&;�W(߁U�R�x(y�H��&��~iT�M��ƕ<���h��}6��Ӥ��E_oX�z�L/K=�qD^�`Զ^7>�L�\��UQ�������vΏ�eC�m%���uLF/�����rjY�<X�*�/�e�JZE,wmdc���a_���	�{�ڪ&~Ϳt�3�8���OL'J�X�3��Jڵĝэk�3|e��r��X[��b\��^'�)|ź�:w<{��WqiH�.�F�x�ƹ(zO�q:ػơU�����O�����Yt��-�"C ���b�u�q������T��ʩ�b���,��� Z�x7.�@�[q��3���ҡ�>��X�ksk 7%]���!�p6VR�l��C�d��j������^�R�j2��"#�_{�z�#�!<�e���Rǳ�3�}�Qj�״&���y�E�Phz�ɯt�4Qb��ʸ,�\��T�U���� ���KzM����'s���/w����Ú*5��OY!d攬i�����&S�[��S��fpp��̏l��q�D����7nAv�0=�B�a�4�t��h����tn�'�}���S���{)�S����p���/pX��|8D���<�yh�l8��"t����%�J�z�A�]|��eFp5�9ֽTU½���j�?����#�1�qa/R3������+n��i��s����^��ԯ�[�-!��V;�g;�M
�7bk0�*s��dk�,�.9
r�:��G�k}��w��<���vP��OO$R�+܌�1�DR#ϖܽ���WF�(9K���މ�6}ތ)���pp%Б��'�r�;���
|[�on1\�f1��/�zS���mQ?�e<*K������J^����n��˂CY=//B�6�.䁿:���oN��j�]kK�J����� g]���8K��ކp�������ւi��F]�3d[�Ka:x�fG'.9��p�otM�v62�$����Fr���� X�(~����ѱ0���*_|���̸���p?���/,��# ���6�V��ݘ(A��Q:'&֐N�^>y\a$: "6�6�%��)W���fwT/)���1�]�
s>B�a�]��4�l�!YK@׏�r*Ꝥ�){w�B��2����c���D�s�W�P�)q�k����k���]bV��X��RbĦѐ*�@�x�#M6T읕�f W"aA%)�/څ5x���vh�w07�*�i�/�LY�Q���0�".��)��ꄛ�T{�����W[a��'I�u���o@���T���7.�K��'@�l+H������5!�rO�t�1'I�Ѕ!�G��ڣ��Y����BnYr���|��t�Q�U&tz��Sn���Ba�Hx�9��RiR�"��|~�4��L��G��5�`xq�ǫme%Ȼ|�%�,��t�b$ �����K��b&��O�Z���+�_��p��ը/|^�A�@ڊ���G3l
�h�A���Y3����'��0(H�-�y����l����K���;_(X��R[���m/Ub�?"�T,��:!��f�����̀�
Y�T����/�L��k�5y���J�ѩ{�ܙ�<�j�	%$��xK!�8�G���ݖD�O��E2FR��%<�pywk��uH�+���b7܀o�"i?-�؁&�%�x믐UQ�X��~�-����ɱ'���.b)��Vo�������ȫ�C	ڄ�L9���P8���t��|�U���h\���ފ�D�\c�d[T| ���_���ۼZLNhe������I�|�GOՓJnai8���� �V6��Pl�t��!{�N�0�f�IV�`��&���� Х�d(QGq� �B��q��7�[+�`��m�Wx<F�e�G�T^�p��@�5D��^Y�߿�S�H�I�U륹~��w�Bŏ�8������]���(6�
��I�Eo
]	����[��{�ϼ]$�p�]���n#!��M����j�p�p��`Dx��>�T�[� ��AJ_oG��3�<k?���d�!�3���*3C�pi$��
Vg��g�$�3�����s��=O�N�f�8H����xF�f���n]W��J��>���O�S[�ax_��S9��i� ���
��ks����M�#��u��a4L5�A�i�u��:����ǯ��%�#
��'7��D���
)��x�j�,��4��	#�~�t��&Ɉ��VP��&H�%1^h��g��+Q��<4��'~ۈ��*id��8�"���C��"J*W��[��Bך2��+T�Q�TK�����������N�ʑ�:Ā���`_�6������f�"�����b�[$�Ȭ�I��j�ɸ%'+�u7�SG�8�믳�r �8X2�n<9���^�Hj�>�r(������m�V~�VT,���~��Y� j �H^u�C!�����n:$/4���K�b�n_*�@<����C]�5]���>9a�	v��`B.�b��:��>0�Po�a�ig8�١&(�B�
�3*T����Fb�5�2�©��&�X�݊�'4>6�wx�?�`�IV{����f�)aJVu:~�w��$��z특���Y�ΘZӄ�f���A%k��ת�S�}�E����XH;`?|OhK������>qڜ�-�+��H��=�(ߩ��N@�r��x-&��V���0����7 /�� �cn&Xz���ւJTN�gI]K��+G�j*~	}H�3�}]�sP��Q�h�]�����Ao�2���Q:"�)6�3��B}_��p�Ԓ���W  Z�`Hu^r�\&T'�}���{��"�	�%�4O/�ل��0�IN{o5W������"�������ʭѱ�(����Mx�L�m¬�PL���Z����ƒ|�i�MG����z�����euk�G_M"�v�<,}����Lw]���>�^����u�EPN,0�YG��J�]���UN��Nϱ*O�A%&W#|0b�]�A�x�
>}�Z�O�2)�?���&�:�~G�����ٺ��tTT��Ȼв�q����_��C�6�K>�%����������jm�Uq�G?�4F�%?85rM�pG�2y�4�D55X�C���z�ɖ�M����L�\e�}h�I�5��w�XA��I���$�R��|�E)W���4�C��h��j�:8Z���fՐ==Yj���x*T�)�K°��v+bv<;&�w�=-�m9�`_��
�H�g��0J	���q;N��t���B5�
J@�p>���X�!���8���n�)�;�G�	m`)��pffr�� P�K�ΰ��&.@sM���T2�:15��E9۾���2jC1�dA��r��K=�m�X��QK���))R��ݐywY�u��8�?�D��{�ĝh�)�e�)�ٸK+}�R�df���hN�}�h5�7�A���]��ۣo��Ù��0:���o\��[e�A}�%7�;3��:y1��3
A5R�hO��cmj5�6��x�S�)1�*�~r��E"$��j�s��&�uY�k8�,�M�ɍ�M_��S��In����q5�\k��+�5M&$��$]C]�J�q�db�5�y�鷻���c���E�l-�&HT�Zv��C妚��i
�ǀ(�� 0pT�����Y��e�����~&��'�kXu�3�L��Q�=]�>�IF�R+հ� ���)p�Q�G��V,y�6oZo�;⿅��aU4t+�w4y��{�~)?���S9�@���dC��&�N-K1g`��t���J'gV�~�{������˿M��E�ޙN���=��h Uo;(�s8�k�m���  �@t�=k�an\�סl�g+^��=����d-s7�������E��ߎ^Nf�ųۨ�Wk�(�9䁟�0޽w�W?��31i�F�11�5�q�I�誫�ߧY���\��V�S�}�,c�yw���!Q�����ʹ����w�"j#,�>�<ӓ�����,��jh�yZ:Xiȸ�H0�)bL�	�>�*
�����P�J���c�k{w8:J���5&`�0�Vm��9��<�[ï}�|�,�s�}a��Wa�:��/kR+��+�a2�F��A
�pV�����
��B�P7`��n�G�kaMA۔WA��FV�-`͠y���yU���X��5-g=X̿�"�q�Y��8������������ C����F}e�O�U<b�$��`�W*��도1;Y6^r�x�	Y��W��){q��P!�I� ޺S����[8*�Z"�lDPvP����Mb0J-��I�*E�Bk����_�a�(�������ڴ�L���j�6�0���U��'*g�[v�$����ߤ�����YG��C�o��P5�{�^���Y�j[!��Zգ)���V	Ӣ#�K�v��_H��4y������%�F vh/�6몏����i�9�`�G:�ǫ���� x3��2̹?2L�ө�]��:�ä!�L��IfY<h9���=���N�@Zh��mb�#K�,@dE0ƺ��k��ҫ;����<vs[d����9F��@����@x�Ҟ��O�0���d�V"��2�\������h��"y�9�jx�QZ���lJS�.���l;�L�	��b�|Nk|'�J���W��ñ�1� �e4�a��«ʘ|�tϪ�T`�����iL;�:Q��E�%,�Kk䰓��
��_I�����~Q �c�@�����pT���c8x`�cm�[Ab��л�����B�=)��Ek�d
t��u@�-�������y���D�8$9�k�b�ܚ�|'ا����۲����wk�!y�5�>��g�<����<����e����8c7�.^3h4�П�T�~�u�ގ�/�W�i�`�a��B,s�y펐'I����V�z��s$;I̯���ٸ�Cw�����|יT0��l���t��gx���M���L��32���eI��"�ĥs���aK����������U-u�R�zM �=��Z����!�z��a�A_�G���ɼ@Y�3�j�> 9����HK�.q��<˔��X���b`�Kyy�
B�W�A��b�NT��v�ӧ,��G��>�u3����AyA�o�
bH�ᝨZ�(�C�j��϶����O�I�o[QҶ����{%C���VܷE H}q��p�>ڮY�煷|\huMJ2
n��{U����M�z�P4�9o��A��������9���@�84ˀ�S�z�/1��&Rv���Ԝ�Ž��D�}��$��բ?XM�Dneİ��ywy���}��(7�6h���[J�,tR1�X���W�����b	,�@��� ��0�k���r>1��}�DE�`*"jr���ʇҋ��7	؄>��3#�[���'�h��t �Zw�6� Ǘ�d`e��o�U���Һ#hRt1xzO�-Ty��'K�oB���W}��x���rsW�\NfQ��rƶ"�"�{1���y#��>с�K{�E�S�R
Td������}Y�)��v���\�腵��D�/��S�y�+ֽ�O���.	7��>����e���ؗ96�+ҴSi���hdF�R�u�]�C�CU�6�Ԣ����<���%�r&�?GY��(�&��N�j=�{g���v�
�9��:ޢ)�׫�Ǧ)���֌�� ��H��R'ݖZ92ًr��L�ra�x����oo�l�
%C�X������>v+)`!��ǲz�V�lw�Br C`���Տ��/�.�`�����=,K�5��y���������C�jچ�y��r�kνd2u3�|a��'G�!N����9"�`�U�8��| ���P?q�9��[���IV�X�00���Y� �i�7�*_Ld�~1GOM�<����Å"�ѓ��b�W^��x�o/Iݚ�'J���[�>`���29����xm�v_(�nC�\�(u�Ќ{�2y�Y�ϻ�1�;�z%Ģ�6X����{���g���0Zx���qI��8���KԁQ���%"�rp���	?ݷ��s �b�<BCh�@��TK�b)��r���[��	��3�n)�A����8���(��ݑ^"��ۧWWz�7Y�)u�a=�-˚��_�2"�tC��/P�t�A�g~!