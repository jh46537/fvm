��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�_PN�2��,H_|O}��$7m�c��`�W�mZ��H���wz'�K�s<{(�*���w�%�:%�o��<+2?�=�l���L�G�n�y	�f��c]��g��77�D|��W�םfʠ�� q4���z��ص�n<S0z)��� ��]|������&(J��� #�eۑ��Nox��c6�)�瑹)Y�����sTt��p��T�j��凞s���<F��s�4����:.��� f Z*��R��?m�%�����Uf�ek�6��g���-���Ny4
�Z���l#ꄞ���-�Df�d�%��|��i�C��ٹ��o#��b�� ar���c"�Fۃ�l�9���6ތ��[�҆g����A�O4Q����hT�W1f��:
�z\n�s�Fz�#E:�9,���D������q���0h���z�E	{D�L�3�������g����z��̓�O�j��`�<�JÁC R
��ڔ��ھҙ;U�! ��T��~�ˊ�jT��T���j�}�������q0�{v#b��r-��n����R���]�CD�kǙ�$�j��q���N3���Z���eq�����2�a3U)�����k�� B:s�.� �}[�,��*��P�悡,O�N�B+��O@�6���G����1^)�˖��B�A|ҥ=�_H�� M�nI�^P�F��(%K%&~>���.���C�
�ft�N�N~Kz�@G�K����D��Br��-U�<�{z���z�0�eX��Hs�v!F�>��i�Y���V	kc�v��L�OU�d���~(�:�Ϗ�f�W��1-ޫ�ǰ������{�w�^��Fo��pV�^�S�[Y�z�T5�Hw	U��+�����X�י7<���� �cUL]�5��b�VڏE:4��T ���2�%��bq`����djqI�f����aG.��	�y;^�)�bJ�m�8�k*7wljw������pc����eo�� U�1׆afW�T9��͛�&Do�M�s;3YU{Q����a;e�sJ��ص_�o����9��L.Q7�d!}Zz��;��1<h�J�#�����D"�j���}`P��I�o�ڽ�K �6�6��9?�����9P����7��_�]���/��VU^h&��_59�ߐp�S���R	��=��d�g8P�Q�	�����Jw��A���~)��*C!���F��Тlw=�6,�5�0;60������og�f�iu��ɭd�"��-
��m ��[�R*ڼP/i3�ɘ2�3���G���6�LPb�~�%�S�wWE�'��Nx�5BvKo��Ab�<k2g+]�-����mN�]U_Ȍ���ۘ��G�gq>
���U��T�'b�ڭ���2���z�=��g�]���4����>�t��&I�*3�{�L��q{��'`����%UOn� "ֵ]/a�!�Q�z�In�\.1���?�e�r	))��M�?�CMB+&�@mz1������DJȮ&����M�zIf�xw�uE��%1��U+}�)k��8�e}��,Š��-�
mښ[Y�d9�-�x��2�R��(g��{��d�0�.��������_�;�H2�){ b�͆�?j)��'R�ݴ.���D<�a�ؙ>;��4���Om�Ȣ���� �l��x�z����@�1�C�o��9�{"B|I��ɼ�(��������L{��}�� ���*D,�<u��H	�ѩl�	��}��O����ӆ����7�i4�I�*�&�B9�y��0���gpd�\< 'O�B8U%\��9C�����܃��1��Np�����!�3��~SN�F�3��u-�	�p>TD�8����q�vt0T�}�z�JP�!u�3�b<5<�G��-���D�s઀���2d��P����WG˜ֽ�B_0taE�����q�`��ȥ�R���w��𒔯����*��;"��)�&�1�25��f2dw��'���(�8/yBg0
_�ܼ~�7S���κv"�^0���!��dQ�L�r�KEr<�9C���򚸋]CMB���5�Q���Q�����]����y����39	W]�>�����̍Z�N-p_��o��A{C԰��#YtC��B�%���5]ެDׂ�d�m��[� p��6��-X��.�al�v,�	1�FR[k�������FOJ�btfۣzQ���j$U6�Ye����f&f6�3�8�����ӵ�� x���jK������ʢ�-a�����B``�����.ls�:�)dG�ؔ��=�zcn��:�?�F��e��7����\�5���7.�@݆$/���KՇ�b��5������"�@�>�8�����؋l�Mx.�v[��PsKʹ$+���E�r#\�Q�����M��`��A�j�9TsGl' �%�����yh�Wo�e¢r��wQcQ�)%d0ҷ��4B6��zj�y�uȆ,c[n'I�����A����(aE9��1z����t/��N~FB���9!�$�:��0�P5$�R��d�#Sӭǧ��4bO�	n!Vk �]���L�θ<��oV��P�/�5y�`o��u��T�a��J�4Е�}{��:���<��FܶC�������E��z��mk�����@Bl�.*��t��ʍ�Us�@���;q�%s�r�2+�u��XDYR|/$�=�y��X������Q}�Iz��c���it�����Ѣ�-�/&@�dp'��{��f٦�� E�=� �1tw��I�*A�Ql�Pg�lKx4�TF���x����������\@�
�G�vw������:�J���r�`6���qh0i�|��� qǬ¼����X��ID�6n)0�K��ICi�s�v��p�"���k��`dܕ�-���P���T�� Z�qȴ`�/`Z!�uck�s���ƥ���K(ѫ�q��7w�3�Ua�$`�0�-
t�^�*�:�4wi��+�\N����-Θ1d�j��K:���G����s�xP���Ͳ�)}�/V2�q�vd���]�c;��#�/uR��]E8#p��4\2������F����۝:�v��A���x��߂�h�p�]�|��o��pի2��<�w-uL���{>�0���՝?L���?�d��κv��"��C����K"z�<��P�9�㲒���f�}���f��TZH��s��l�RB���������dL<����]>�B�ח߆N�]�b�L�/��.����E)�TOE���\�>��!�?�!l�Xۄ��p���������7�8Y��9*p ���LL��g�_Cy��(�8�]6�Ūg�LA\�>}��-�8�7~��Z6�.��*�k�� +̋F�k(j��G�6�/�
U�z�Q�^o6B���xd0�_#�G��[�3ĉ]1�����D�!�Ot
Y�N��?dpGXÁ�����o{R�hi�9E�~]�� ���+�Ǹ^�@�|o���V�M�r�Y_.gJb�r�F˞����ռ[��`�,�k`N�f�����o"�G�,�
��Pc���c����(�9-*
���'��*��e���g	�q9�����$Z��{[�KڢAUh��*D#��E��]�ތ���[�Mh�i�}�*�Ȓ>4l��';`��X��d�d�	�$��K^Ҷ������U�?t�7�Q��-��@�����Y�b�2�V+��b�t+O��A�ju@�車��6�f!��hs��{孳�)�w�óR!N,���3�Db0�#Ƈ3|�*�>���^Z4�e��+ooF	S���mI�4����9��M�)<N\,�3��gX�����՗{WCI7iPd����>c�������ԉ��7���I�?tX׹y"�;{~�V`�dW����j���*|)�+٬>+2�6�v��~[�,I�P��z�x79���
�D_�q�J��:�`*Vp�,�z2O��Mp�z(hB�kz_C*����͎A�*�9���q1�YҰ�g��%�1����+�c���Q�=9�m�V�� �z(�D�9�ĳ���5f��+WK����i�Q�����0�1�=�W{���
�����l��>�K93���ݖ2�`pI_e5�aQ��D`_b�Q�^����/����;N��t�o$�0�D&�Ur�H1���~��CNY�y�~�n�`?gGF��&����BK�1J�#1Q��'H%`~�LC�2� �%�\�7��:Pu�������)�c;	̽�_Q㋚�N����A��^M��h��q��s��ŵ��a��-�1+2T���&��l�G6�.� x���ao�&��r^��>{"[˂�N
�m�pE�+�й�X���Ȉ����=lQ��O2y=%��q� �zjO�!sm|��U�S�hj��$d秫�a����:���,�U��8��v�4_y"�cVR�$�;t�+���	dz��h�����I�q����ǉ��svނs��ɾRI�k��z���om։��?��l4Z�����8/�cgǋ�R�� �W��n;�Y����^'�fj�CNɰT��)T��Gs��L��K��Վ���7�}Ӊ�}���i���0帩o6ǧ8n6���>�IxoYQ~��i%�Y���N�64nF�;��޻���Ϳ*}C�:���qP�ne?��1	EнЗ����s��hw������l������5�wl�zҽǟ��Q�[�TSWtP~/G�^�����k=�DGs�P@_&�~G�W�wjDAz��O�[��HVП�*����(�k�uO=�k���qS�>$
�u���^d���(,$SQ����*4�=�@<�r���\#�T�~WBMgF���;q��;��2 9o���\�z��=J�A4�]r�@.r��#��>ƃ.Vc��H�k
�'6�9K�53��~��� ��n���h �'y�m�"���ٴ�,&?]���FN�@t	c&Ub �~�cSaX��}�i�'"[`��e�(�E˺�x�`�Y�����V:JTپl��w
Q=z��2	M�,�� g��E���K�`i��/���9'j��k�nT���?YVƀ����be�������(���j�Nd��~�vF�c�S����I�
<$��R��v��H�0�W��H��?!r�T�Yw{㒳��ДeK\�(,�(�)�K�Q�a����,��'�l���2^�!������:�TD!�e�H�ɬ񄶫���$II&�8��_�a:+U���]>���d�&t��8��i��DvMˑp0�Y;��LS�'�e��Qu=�	Q���{;;����b�'�kٓ[T���9�� h$�Q�[V_@Jx��?����ʑ��vJ���p�ϗ����qZ:"�γ+�}I��Ĩ2
Sb���I7���~=V8�q	��I�?q�92$��2�E]S��� ����w���k`�t��U�V��gu���5Ӫ�O�rj��(��*��x��'O�)�/8�g�q���E6�����4s���(�Q��O���|<=�!ba�N`_�2c�Mx&�6b���ax�
?:��~;۾aw�|
��P{�dr�C�)9����q�C,3L�I���2���py��)���3����/2M�?������:�r�;
��FF�U^@�,iui9\�Յ"y�|{Pew-#ޝV��w]_^�p�n�h[�@t՞Y��R�ߔ�M�ܢP�ìT��p�����z��@Ht��uT4Ʉ[tQt���m���Ԥ	�?c1�Y�빙2�Tנ�׫�Q�ؽ�+ֲ]��A�}�y�d�f��h"A�$�u�	Ο0OiV�~��|�8}�������d��i�&����$����*��)�0���NP������fn�Ϳ>��]�`4����N�ܓC��N"��!��.I���J��	f��-
�:
	v.VjF��Nz�?��BҮ�����-�JV��B��M�8�$�Ϲ��א����,�9��+�j�S��=�;����Vj��˞� 91k1��q�'�a64O��H�͵���D9����>�D]�\S*\�3S���94�鈠&����T�~�G�`s��fw.!�X��p��VsA.K8<��@�9:B�CR��7����'J��m�[������_+�.<�P��,��r��X��0R�=ߧ_ulE�������+ ��5jʪ��Bz��;��(K��8٥E��"e�J�$�^�9f �'�������^��ZL�|c��B�<I��z0���.�*����8��?��&D�6nz��I�|F>S��.|IQ���Q��������3����͔��Ӡ$/�n��A> �.D�����)�|撝<�Ic��H=�@>?Pw���C�n;/�G���9e�>�6���#;w�v/{�C�e��j�9�����WH�p� ��f���בc�#4v7��mk�c��b�)�q�Y_:)v���6![Zq��0�����A���H:����TF�&��f7�kqi�+'�^$����aG�_'��{�H@oW�a>�9()�V�r�~�e���C^��`��t�Ϛ3�`?c�Tk�[��-��$���H��Q;�l�jMw�y5p�sK�4���<�<9R�#�������Tο�Vm֣g31�[ ��	�o�:��@��9�p�[�v�Xu�/n�4�6���=�[�W���O	̓�/�^էO���79��j�2�$�(�S� �+�t%#_���lu�{r�Ց!�@��ҍ"�PW�yю�
e�0+��\�.�þ73���ȭ�i2�j#������)�<�+�y�GI��,��]����5T�گ$�j��\��H;E!>Z��/�'��]#����=o��
���\U؝���MVle��z�'��B��+�����������c}����nc�e�yE���Ni'6����r�#���@��ܕ��=���h�p�%.�����:�ưW�~t���2m�]к`[۠����1S6��ks���?��u�����*0G��TY���<�Ŗ=��y��u~�����*���/�F�z�D�q���a�O٣qu>u1�H0v�"w�p�c��C��z~� !��M�Ƥ;�Ӯj�u��1<z$���V��}�u���ޖz�������tܤ@v|~�s� �
�k�l<�oJ:���㋛s[��2s����D�uk�X2�#ly�?iS\�It���N�}��������\���3�b��M�n�-��
%ѿ>u�8�h�mB���1�Yp̣��*�j�h?��<+�JFC.�O
��\y��|�ϕaj
P�b�g�G�[/-�m���U�eLE�O�R~by�Fw�i����@��jN�����-]��!Vk�ڃ�G���$��1���E�v@J��fpe�j��� �y�z���`�R9H'�́M�ɗ��[]��*���^��&�y���Ț8躏��hMv�Zx���rP�I�2��.ʮ�z�>�C��v��S�*m ⏟=�%����P<�4�K����|�>���(>M�$p����a�B��7ĳb�Є��c� E�\i��M���7l�l�I:��-<�����g���zp�����CjB�.c?�$��l�`�%��ؐѾ��E��y�'p�S� �d��]��ମ��^��n�%��������ܻP�0`
3��
��g��q�XhO]R�,�$��G!0���t�uY��4u�s�l�u��������(u�L�<a{��1.�f��SDy�IHZ��~�J[���i�ǤI�ڢ�0���T;`��|ܔO���Ge�aC���� ������$�dwȠW	������Qin"�R �&bL[�K �c��7 �I:���d�@L8���e`�`:#c�<(Z����e)#�?4w�Y3;Fq@h��^���ȭK�\�>���0՛S�-w���>������b�]$��!�F��x׍'��c����WDz�"E19�ۀ��^lGd*��Vx߸�MQ&ǃt70-)׈��@K�9vޗ��r��p���9������iksn�$6����e�e�ۮ3����D۔�V�71uPt,���6ӣ���U��~k�$��Ń�h��d���S7� N*��5�뇋�����J���!�N��:�Z�ס���H0�3(����u�h%�垈��ǎ��.XKlY��9F���B�e�;������=�|j6�g
5(v ��Ĩ��je����J�sX_e4g���^��W�c8���A���5��������:s����a_Z�"�8����	'E�p/N��YΎ&X4�h/ԸN���Iˬ��o�����q.�8�8�����s�Ahmg�C�2.+.�E�y�5WkT趲`�%mvC��Ey��0������gʃ����/G*�2���9~U�S$��c�~K���c+�!V��"��jъ=�lc!F��f_|�"���|��?>�+�A�@�I�<NP7>L���n2�<��Z�k�,:X���'��׿u��u��l$�cX�(Z(h��"O�!��ڰo6��$-֮I��}���&{|��U���Wz>3<b��G�SUTc�%2"Ѻ��Y�N��}u9���x+�B(�z���M3���K|4�lk�ڤ+�y����1��`?r}����A5�Y��An9#�dxT�F�M-\����g���.��n��h��x�-��T*t��/�m.۔��g�D�^l����'�6Ȭ� 'd��6V�$��y�zj�☪�W�1�XHwSsX��-r��P�앩�h�J1|�#��u�?A�L���9�ń-k�Vz큭B���e%�:�t�r����1�VMGQ��
�&%���@1�����N�h�2�K|����cn*ϔk�S��Ԓ����Q��>֟sm��B�)? �+��GþY����TU�d�c�K6�r�?�?r���2�xsn������^�Sc���lg�Ecy�ߡ�����d UO �w��
,�m�d��J�'$�WT��ê�B_N���tI>���V�w�51;��U�*5,G>�}!q�O��$/&�[ㅢ`Z�L�u����gdM5�>�!���]�>�B�j�n=�<x��5T��]_�2�7�~n�y��;�g]a<��m]�l�z�@�.�����ã��m=i,*Z�&�2�*rN�aM�N���	���Q)p�]ٝ�n빗Xx���f\8�uA�-����9�OR=0:��;�5�z��\�4`���{>mq�.A���e���(PȔ�!�Dq�p�TD&(|=�#D<����*G��7��:�]���;8�/� �+�J�/<F|m�v�ۡ�,<��;k$�/�.t2�/�;�T_6�]'�wqp}���[$,�#݊t��^H�����f����З[����ge=�uU�5��:���Y�ALȣ@ޥ{�B��Ɋ.̓'x�$'eW�T���~�U�D;�|TML����e����nA�����~I.�!����9�P^�.��L��	