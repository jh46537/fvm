��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�z吴�)b���ΡrϷ���	�J��Ȝ��ݬ#��<g'�"]�w_�,� ��3Ե��V��<�Xmd�����&;[I�n�N�K�7���bX���f��6��u�����rq���V0<������+{�1$f�Z�Mu	�"�韣��J�#�bML���9p�k ��Ӄ�G��j�bA�i�[jLsVkN0���ɐ]xOU�p�f��1: ��h�9@�����{��Sck���0p�Ќ�{�����{�{#qݕ\�	�$�%�|�PFZ�9�s2�%;���_fp����nu 6DQ�EMc��A>��x��L��'ϩ��y�<�~�:���Ad��f���:rU�衙��*����6����oD��2������Z�&8Ӭ�G��k62G�Gt��/�=M���`��$��$ �����(�٠�>��A�vo����,!\;m3Ǫ{���^�@�d�&�H�LI��:�
��Q�X������7����=M�~��;{ip��!�J���@��%�����u�QN���]�}��H��ǫ��2H�.��}#F�@!����	*K�U�VB@�y��l�.�z��UЗ �	v�td����Ac����>4u�E�FK/7|O���&��\���9^;�E�x<^��N�2�>�hN�D�,�Q���?!L�9_�r9�f������L��5ز|p����tu�n_7�;�r_���������4�_S'�V^5��G�н��UXic~<9ѿH���c���H����G-f��)l�6�Y0�'���#���aiKV5�m{�S��<��cc�4�­8��Kct�m=�;�۫,��p�}~� �O]`>�|��Г��ʇH�<�F�w�'S�����/�[ʀ	@){+an���I:�̏���}����^��MB��l���TX8+�
����M6z����)jE~0���{�X���7�#�r�>�?���^�"��2����|�n9��-��,�}Sr��r���$�yS�c����l�#�����)H���@P3�Q�Q��4��>V��7�����������W�H��p>4M6;0u��m�$u׻w����g ��)@lg�0�[	1�V�RId86SR��޶�X�^��Q��^��Ӣi'��4U�BÇ����b#�a��9~"�/�m`�?&j�;}dwi9��0>q��1T���!���`��X�䅖S�&��Z���gI�kE��j5��_^m��Is ~�[��ɕ���ɱ�Ъ`U���ޝ�!4W����̊f�͕�O����d=��9C�NMd%�	&. `�Quh�m���㨛}4rVa�åF��b�h�d�07��D�g?? u?��âG�	.w���q�ꀦ�VN�c����//����ne/�B sy�lz�0yV��e�c����QoI?�l
�����C.�|$��z�Rj]�R<�m�E� =�?���s��������	We��R>3�[�z���lA�C�t�.Hsη)�ʦ�бS�!$����ζ�Mάn�?5�f��=��-���[BW>�jaрdt0]�Ea]a�l��w��?��(ouw�s�@�h�1<mP,gv/��ti}2k
����i�6��3a�3%酥���Zǁ�p�<�#̾�H�;�B�k�m���Կf�R��CvU#�P��G�VpHq