��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb0(����	zik�0���~�2>+��$s7k |w�p�J!66�څ_��s��8fK'O#W� \�y�>4�O�����?!�'�����{� �ׁ�a-T�z���?r����K���+[J�0�J.�����5�(��#�ϸ!���8
�:�@}��0}��N^z�7$!��;��ԱFҞ�~�O��j�/�q�h��oVt�]���C�IA�����0�e{ݬ\.=�D[l1Γt\�RI�C+�|=;oN<�~-���N��6!�B��c��4R�z��T5U�9��H/��4wb�J��[��) d�v�ٗxP<\���t��>�t�����'��������~���v�?���d��
���$�
J;������ir�Mk���f2w4�iW���h�J�HkY|�6�J?�����ޏf�|ɷ!=D��t`��Y��8g����8r�;p�w���a��̡'��{���<��":��ж~)�`ݜ�8�3	����jF|ח�5�^]��1T�;S"�|�1�Kb8]�yr��b�C?�9_�y�d	�K�	{�>��Z�X���5���Ɛ`u�u���J��
t�~M��b/���`�����`O0D?�v�K<��6��a�73��ZK�%�P)a�@^��pxa&IZ�F�ʵ��x0X@MWs뫿_;�B���N�>+�h����4j�������a��Y�z��.~�_"Y9��z�Op&=�E,F�0�ߗsk+�;HB�Zi�4g$���
��9t/��n��pxp��n���!���A����b�z�ad�}�nuD"to�=oZ��䥠/B��.vûC�4A��O��?�?���ǡn-Uy��� ]FIޙ����%�EN����Ԥ|��e��i�P]*�6 _:����2{�S�b�������q��|G6;tv�/��l�ս���ٰZ4���D��y��������ꚵ�:`���p���ԃ?G����It�٫��,��a�,k����ka1,&��<���������7(+(M�?���PĲ��C�[�.9�����|U {�I1���c��b���iU�R u&9��oѴE{��LI>BY3�0~AdS�a�>��J�����?����O�y��B�g�^�����}�Ǌ��B�8�DfU����(Ϧ�N�6S���g����Ql���tIYni����t���%�$'����pNY��Q�of(�<;E���w�"d�E���?HG��K�~b
�^�Z9i3)M@U����P��G.���r��Yx����c6	�T�1�M��ۉ�ҁ� �,���=�[#\�(s�.��6��kć����]}9?�����h�.4���HV���Hv>�5r%U��t;&���B=�WQѸ��	��pU�E?�_$�I�i�
vMK�����'�$����مԻr�w�J5�9�i�*��&MT�
��\1Bڋ���ĕ/�+Ôǜ �g(��?����;���و�af���~�9���n�"��Ny�93��]�j��t�$��aI��4�]�jK"w��?"��>�o���y�j#Mû�nѸ��K�a�^�6��K���(��/M[�D{(,��		{@��bBzԽ�0����%�$���,�a�:Ĺ�9Za�=݃
M�����H�:gz�u�=��IG��P�B�)�j��[�g�]��n���U���ת�8���I�Yv^�g�X|^i(����A���	U�G�z����\���T@y9�a&���r�s<yȊV��8��o�>��O�2�K#x����F�EI�<*V�[G��c4hLA��ilq�+ڒ��W$�榔x�����c�.�ٷrG�zH��[.Wd*Ј�y�L6����dɅV�̝Z=Mu�ѷ���ZC�_*�f8��oUF���s�0�N�&eD�b�G3���jc�w�O'L&�j�Х��1�ɤ׷K�����&S�ˡ�7��N~���	�@f�����Q�Ͼl�ј�B��%CI����b���Dӿ!Y\�v���R�47�GN��($(���U�b��(�߱1W.&
ڀ�������	���q�'9�؄w��p� ���Z��H*�x�7�U�A��P��iyafj����}�iK���%�ݤ�M�M���I��{��8��0�ߌ��)���/	A>�G/�GZ-a��h��W댆1J|�;9�<�؏E��5AnWj�
��z8�ݺ�B��U���4g,�����~��!��1�����q�~��TW?��}��`�[M�ƫ���X1HLI�v��E��MڞzD�o^�+��\����-�kw���0.�p�+��j�KU�ק���yY@�4M��9%�u�~�v6��է�^�����N�As�2^��1���!jF�ⴴ��~~�R`a����|g���i
t�z9��2�"?W��CjV/RU��*��'M��k��̺�G�ɓi�� �v��$G''���PD�<�̥�is�
����
� |��۷����F�ܖ]
(�"�wY�C׿bb�9�= �7��X��0���=L�	����SHę9͒a�dz��4�{XY��Y�qds�,��T	w�;^A�b�\]EP)/L�,�s�ENq�>t������~���r��lR��R���E��jBWX�}?G��ү��yEzl�^�ϲ�Q�htD��h��W���SN������<��[��f�� -��UNq��ђ�W.�'�X���;�v�/-�#����3��_d�cΖ
1�x,�i��`��}��(��L٧b�P�Ȧ)zL���o������X)4�XS���Ty��i�$�,�_�=mK�GF��OJTQoq��g������ޝ�������|e�X�w��&]c���*�y8��nn#K&�*��+ �����@�E�I`��l�)11�F�;��N^��`\�Ӧ)x�l����(ny�4�@�t�D��Q��}G �3a�k�f�nIQ�D���; rI#	M��g���2P� S����f����{}�;X(p��#Uv��� �(W�[�UM��#bo K�g�E�<���$E��Z3]7=U��0�"r��� v�)۷�^��O*�۹l�&���m�*bp��n��MN����A��T���n�4���8Hi6xP��,V��2�w�	p��R�7�[�e)��=`/�o#W	o��Xq�bV%�Pp]"ϲFs�S)��h�W]!�VAD�����!��S�J����Ү�|:9N�E���6	>�ާ��Vk0��F3!O�es�����r�O4�Ƨ���>��J�cL���,ư��r$C�Σ7��ǍD	���HߛU� L�aa1l�E�M���S����x���� j?P���.#�u�:c�C[�`ִǰ������4s�S����'�t�Egz̒8��!�h�W�.1^I�T�������$f�B�F�跂U�� �|�G=�r�}�N�M�F_X����J{�bU��,����ݵN�i�]|$��Z�q.'F�(��ஏ��Up�����������Q�k��ډ�9�*L�8 �խ˜�7ΞN�d���B���1,�bЛ�d�e�yx����hq��P����ñ�~Jդ�e~�9��ғ�[C�6m�9�I�U�L�.~��d�s��v$ ��kH&��:(-��bW�3�� c��/�x*;4�$��D�=��]�xL�>�T��Ƈ�{c�	�ou�/)~y�د���[Rq�A<ēv� �M4��t����a�f����
"f�	!q�ɢU��%��Q��ڷ�ۖ��(C��}���Ȥ(|Ϊx�3��A����QX��'��H��g���#'��Z��1�(��L�Py�U��2�'  �#�y�݌��<��~1�gb���,i�e6��;5 i����{�^ӹ,�+����[�I�-�O�D�0�b�=?�ut�KҰ=x�:K��~�m �i��y�(���S�%��a��d��қ	���u1�?���C1�.x��>����!�ޡ�Ԧ����il���Ƒ�o^�>k($Â�b]O�U�g�{��e�����F�!��������3{2ۘK�H93�ݲ�� �����;z�mK� ���.礲>`�fI�fЅ�u�7s�"��uˏ��Ƅ׽k4�.�Gx�)��c�E�k �3;w����h��;H�� 7#��Zl�3� �d�<�d�2S �xy�'�`U�h���j�h�'�RI�mG?<+g�Bra3ޒ/�Y�7��>���~�H�y>�F�kt�C�����C������}��[{_$�6h�����>�W�w&b���dxh��-ӷO\Ի[�ږ�����kMymA�4��< �H?����G�o����_��\�{�@�	�k6J<�g3���0Ѹ��S6Y�>��#8��C�`-��RPM��F�������C?���u�b'S+*Q&� A�Sը�]s��ø��K��2��D#ǽ�-�$�Wi
K+酹�%�Q�>���i�n��&C���*��O�9r��x�I�Y�Q�X(�L]&�(nZ=ැ�P�sH�B�~]M���(��&qP�E����b��B��S������
����Ջ3�ֲ�]���\��d&���;�����f1SNw��B��9|j�-Vv���v��4�L�[E�  A��J������S�w���l4���X�~o߱�	C�(*��0L���2�JKi� �В �(O^�a1$K���7�%r)nY�R�"�Hz�I)��Hs�	�d8.�I'�w=G���mY��/����e7���ѓ���Э-߀*�u*WB�g��C�;�N�5��4w�hf]ʿ�725b���J�XF4ɜ��аGģ��3��iI����� F(����ѕ������N�q��3����h�&���6GTraa�y��
��Y�柾F�O�)� 5p�����Zr�U`�=���T����Jl,W�vq��U+�i���n���3�ߙ�����_W�l��g��!^7�C�&��c\���;j�nt�(=��ΰ�t���!�(����9��O R�DI��������hZ(T%���hi�=j��,�^�i�{�á��c=�-Zňf�<tui�|6sy$$#9���ҭf���	lؿ�1|�fe�'�H��s�N�`E�dd�/�*Vֻ��x�K�i`����l�	�z50�G��,���\�[�����!����\�WtM�iF�D}e��ۧ�b���"�\ ���7��PI��JR\~-Ȑj[�/�lT���,��p�u��\�̣�����S󂧷�����;��0��ΐ���e�'3�`����i#��fS�$+���;ԓ5RK�]M�����P��������퇴)C��v�Ž����|h?�ςŜ��F�|�.���#��'���}�M�=���Ib&���{r�/��ty�&�)ۤ�ȱ��2�:K��JB�y��b�X!����9S��"n
���ByO�±(:�;.i���
uy3�J�A�S��ӛ��0\�w��ﾙ\�DZ��k��J��m}ɗDh�Xے�?�'�ky��-ZP[ޮ7�Js�����WP�>�Gr5�V}i�p�[ vA�+NLNU�$3��P��Qb.�7
4Z��L,3?�����
>c^TRMx���J��oT@;�O׎�v�`~��1��L�M�䆒0��h&������fA�|�yR�3�78V�P�*k��KL�x���Jq�[�G�/(�{��ɴ$�)Y_�)����N|��
l}����lr>sD�2<�'��tQ�����_����Ǽ Ltg�I�p�+F���P�"^�bat��x5�\�e��,`-�[�Q`C�Yi~'U����DZSZ����` �8,W�"��]�ޏ=��6�K2����N��L +l���<lc�9@�&P�BNϮvq�ab����8y�I�D$ģ������ $���E�}Fʦ�`��X,��2؊H�,�70�\�$>�~�ug���H�'�V9h���};�K�����7_�3v�`��	�g��w6>�����O�?s��{��~�/�JR��t�m7Ex�����G��8�M��5�L����ܳ�* �����"iG줙*�w��!�/7���_�Y>��tU:|�8I�>T��o_g��qZ�}}���vS�F�@��gܿNW��R�i�z�l��h�q�Z�\3�vc��{�����A�R����M�ݳ5�o���G�e�����1?�B�v+6��� ���B��U�!���=��B�M]�
�D�C��T���z�6,������b�{ըe8^���əX|<�����,���ǒ�9��D�V���7�F�����T|�^�rԛ�~��'���@�uH|L*Y�;��a�B+A�THXd���x7�	Ykq�f�%�r}�%��}� /G���@�q�@lQ�[��d0�c��z;7E�
< �<���sh�a��q;���(D`�Lq��F��v�w8��nY����fU�!p�>����@`��cj~��OoȴF�4u[���Д����Xǀj ��4�>!����-t�@����u[�5]���9C�7λ��~����^|�n>O��a��t",7�1k�4�(�U�9V�D*�bx��ͻ����Ν���,�l������������T�H~���F�|��11�x+���V�c�9�>hD��7���0���D}���y@u��o�$�����̬9�ɗB3e��@f�j�r�`pR��(����cAZ��)�����7XѦ����1���aj��炣%��Y��T�΢U���n�&ӎ�����s��^�������V�l�	��wr9���UUg�%�K��7�����"�?��Ik�'90,�����I�|34��b�q�2x/1����).��H���y��{U%8T��Iվӳ���̖zC��(��i�#�$���,��?)ձ|��_V���v��8�q�q�N$u�\�2ϯ8q:�g�J�1`ږ8�c�>dV"���&;��������b���K����ˮ���H6�����V��ԃm�[�a��iU�4��U@�8i���q�1����V�(˥蝢�����s�MKv����"!p��1}_�x��*���F�8�5��5���u��9�G ��B�$��wXWW�W	�!b�L3������3yy��R��=�ҚБ�)D�(���c&;��d���Z�%��Z���7?C��c�WY�W]J���h��f?�K[�=RC<�z5�kwAβ�S�	�Y�
ړ�q���;�۾r����Ԕ�{���oh(��qK���柜�8)���}�����% �V��K�n��l�y��걍�@R/e"c��A���GZx�5Ϥ�Y�v�K1��\
�v�o	�u���������Vu3�f��c������4y����ڋ%����7,ͦ����b���f�̈́�<��3��t�>5�g���f�.q%��~����3Z�q32�h�9���C0Ͻ��;�����\�{Xz"�>����Æ�.xgLBR�J�m� o!0ib��elUZ����Е%<䆵��eGG�YCs��O~����V�4o��e��0N�Rk�$�@�x̰8O��xW*F��;��sn���k�� �D|G���|�1���Ћx蒊B���<.���^A��#k�EWD;I��`����-��ɘL�,��,��m��l� ��&Ђ��<`Ǔ��Xo0�o�q���ɄN R RT�������*��?J�[�5̛��q��ma���kd8�v��M+�͑��h��j���*��7ֈ�;}8�܅x�~�i��n<����%m��x	l=���mZ��WjZ�G�C9��(RC:���0g�Nzn*^b�ZS���� &WJ�5$��:>d��
Q�"?�,j�������!iʉ5��5��7��_�W�\{�uy$�U@M��!���A1�э�p��Rd �Z3��݄M0�!IFm�鐷�m