��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z�����#0n�ҁP�+��k�cH0�M�ʓ�g���ं�,��fY�0�����U�
����bU���;�j��9!+�	���1�����R�z�������
��H�A0����!� A��2������^z��L�ʐ�j�y���'���Yl���Ϭr?󈋾�{���]J3�ڃy:c�ό�-D�U��G�^<���"iS��D�YM�������0��J­x܎({�c��ڳR���]G���(�U6G���JŮ9�f��,��p� ^ Y�c����p���K r�����@�C�$��g�/|�1�<�9���wr`8F=)5I0'����QS6jB��m)[&t3o$�\�g<�Y{t��f��i��zqN���z!��["�3'Sw��$k,,���A��`�]M�~���m�8�jPip�fR�Ii���߀= 雳�DxPdܡqɋפ��	8���׿G"7h����˗{%�u����^t�2�KWy����պ=��~��s~H.�vp�a�#�n=����$�XX⤌c޽���F̯�.�v������4��"�}�y����P�����M��ٽ���d�Ig!C����n���n�-��<���S ?w�T��+,5��1=�X�_�����Z���Y��ob��U{C 7J�����7�;��K���X���#�z�r�i���-z8�W��6�C$�}���v�` [�aj��b?VX��}
֘WW1n�����z1��)�@�P.�K��bP�;��W�
�
5啚���=�+p���CK	� A��	�D���ᆨ��I���n�� 8�c^�F ����F#l�p�ۙYʔ��P?JV��߀������{3k�*M���V�fd�!�G�̰Nz���Is�=�9�p��~K���)�a�w6��3�>�������ni�Y�]S`��9�52&c�D��K;��2a�u�G�_vE��v��!��$�~�[ �=��<ʩ;��Ns��e�{J� T3��զ\�uM������P�W�$WQ���o.$Ap,.�C�2��1e,��󡣂�A�r�\�	�O�g"���+U��ǘ��[,U���ѓ�a���=qH��q�,�%�M�xy�!��j]a2|$(ӆy�#q�����k�|��It4�1jTs����{��O�#�In��B4���YƝꌉ�'����i��S^0���!�)�������� ��@t%/^���Uw*�;�W�¯a��r�$�t�i O����o��A�x�&m�7��S.Q\i��<!5i��P�{����Iy�DG����\��eX6�A������F��w�UE�rhq[�&�/9�=��oƫCؐ!�?�B�kƏ��O��9�]������gR��f��ȠQ�"S"ih�i�<S���
�Nf!��s�g��2N�*'�Ep�8u��`p/�8WG`b��]l~�䁛1�Em��%�����㮗�7���{���|����gd���ݣ��f�g���2��$ڧ(���g��s��	)�U( es������ل�Vh�74L:H^w��R �
u���)�o>�;8�2uBتE+i!��_�&�A��ж�%E4�=��Ѓ����C�a�R� :��>�N���/3
Ub�z��x��+o��G����e��r���Ɏ{��C�)'�t	ZN�T{W��«W��<�y��V����-CBWjd��z��d`?��F�V^Ǩ�^�z�At�^�П�GSO,�O
˃t����w �B� ��U�(h��d����%|�y;ܤ#ac�n�Ei%��Ƶ�݁����o6k<��xW�����`�y�"T�6��͍t�{�#�j��()�gY�[?Q���Wy���1GEWa0�}p�%��H����/�L/3�K��9���onc,�ml����Ϣb�{����,�J�KQ:ʺZEc�SU�K�L����4+|T��u�����֡Jc��-nߊ�^8Vm���WA�ԙ���>�@d�t�D�Wtт����r��,�i�ȀZ1h�XI4�� D�����B��6z��Q"D(�Z@��Eh?���yu��"�ݲvk�r��U5���}X��̪r;�,?͓���q�4��#ޙ�6>���T�0�����������0�@�zۆ���W����=ʦ�U������\��M�k�|�h�ЏQ.�o�5L�4��f[Nbj�u#�u�jS��O��4R&���7����Y���թ[^Ol��G��ň��s6n��g'0��A>��h�������N�2��n����H�6��s�F�&���j�Mɪ��&�oa�^	�#Q�K)[���~ÉkޑP]���P�Z ���y�RӘM&�Ge- -��B��{�}:ٌKbq��A���P������;R/񚑗�w	�1\*>�SU�Q���Q�՟!�*D��,#���t+�W�ˈTxmXpu�P���J���0��'�����f�%�K}z+����͛����������o��c� mc�J���朰�,�(��C�.3>��gh�8q[��-�����};�����uT~���ްe�͖<0�V'��Է��v軆_���ӱ`��������(+v�]9�'����e��G�*X�^��_:׹-�W����8u�t!�~i]~�N?X@X]9�SQy��Xj��MQq`r=���9��˸�8�G���x��@��)I\�T�Af�mP���s|���Kј���m94�1�$J���x>c��ݓA-���A�E�	�)Cc�����T�i���i}t���^�� ����עc�9�[,!��ƻ�Z�(�r�"���LW��7���
���O.Q/"
I�������ܘ��7�,@���i'�˸���(*+���&	���g����D�w�Ä�)'�c�<�V��� ʪa�{�����l��[9���(�@�~��W:2/�,�l�y��{�(�Ƃ
u�3\�����1�n��(��u��m��SFn����*�YN��mw�b$]��u>�K���Ӻ4��tWy�RZ��;U�d�;NtO��-��T��Ϩ7ս�l�L��KO��?����8�^�$��.�����W9��8��j��=���x=�i����A�%�}�>/�Ġ�(9͍y<���L�ţ�6�����Keu�v�J"��ы�U?�M��Aґ�U�z�q�
[�R8?}�$�����bd���}��^sƾ��~Ɯ;�疃�[d�ݡ���97;�?"��Aw����@knQ�i,�'�қ������'�¼S�9�D�|��7�_>(�~nI(4������y/��S���86*?oE/Y�g_��}�'��!ؔ!C��b�0�R�6����dk�I�O�y#s�Ȟ�Ɖ��x���Z��\��pJs��5 =���Rژ�r�V4�5㾂�n	[ o�ڔm�PG�  ,Bc�6��daO�9*����G�� �M��a,	u	��P�� �n���������%|��%���%Hh��M��2yX�)�	r[�j�D��ft�8O����7�>e��,���NIY����GTJ��pGV��$nt$��k��Q��y� �A�G<��S1��1 ��3$)�wE.,T���\<�k*�Y�֬��)��.r�G��cHҏ7WZ��}�BH�p�� ��4�����J����ȡ��Y�u������Q�²B�ޓKCC|&�N\�}tqv=#$�N�ѹP-��7R��I-ƆZ�����dϻ9���p{�4�qV�X�S�;㱝���xxo�������0Ϛtb+���U��n��%h�R֔������"Se��gD���A���v�N�ڔ`�9�Y�.�"w��1iG�+��n�Ξ��S��v�R�ᶌ}T�b���}K
DRI�U񷩊8g�no*��r-'rN�Z"���a� S���T:�	��
�"�H$�@*hu���j*~Z�lK� F�d��X�o�g��o�Ξ��.iʗ�Kb�/�"��r�G��s�ICV�rfB6J�2msB_��w�D�P���n�����z�Ŝ9ҜC�e�o����Y�+=>D�{S��RYGO��w��W)n�0�,L�):F�@��\�4@a��Qѹ���4V���̎��@��gG��i����U����Yi���.�e(R{��A����Fk�*�g��� gieӤ��)1��Z���mK�,����ƈ9��.(H�+'��DS��~�N�t��W�{�E����i0f�@}��V��/���WTuA��k:5b(��V{Ԑ7�%(Y&K)��Q��� Y=V�Q#W��j��x�u�[�f�4�%�|A$�D������S.�]�#9��rx��HGz����p��� �O�øk2�o�ܼ��P�<��٥� <�E��w9�J��$�ʡ>�Wd������u�"��$[~��t�������d�^�<��� �w>-mS�&��W�w`��xF��7<��2ۉ�Fd)��M$}�=�&��ٮh+k�[�LSy{R$���9L�9	҄�2c����^l�knn�I�Z�R|f���:#��JfӛȱE�Gs��J���k��FO+���g��.]�>���Q҃Q�lr>[sb������֊[�[�Z!�b!Cb�a�O�Zu�D��E��J��-l����az�ORd�������d�Ar�ޗ����N2c�6�77\@db������&_A����5���?6�A*ɞ':��	fO?�_�������U3	RĨ��~R�-P�dq�Wd�f 4q������*�Y�A���,[H6�; �?N6&��7��	��:ڊ�X��+�i5d�w��72�w��|֖�o�4�CֹQ�(�%d�CQ��h��6ՊO ��)�*�Lj��ʯ�`��:qh7�@}e��
���͇Cy��ҽj�n�Am#D�+-3�MѵY.�xY��9��+C���k�tC��i�H��n��#�$�dk�y��B���� ���T�lͧ@l���mtէu�/)��|�z�^`Ƚ��9�N2-u�t��T|=aph*�w��.�@��Zij�+���g	V�DENW�=e����bq���.(�fF���������ԉ/a��V$pJ�y{�--'�|���Ȍ�EAJSa[�R؊�p� ���B����`��I8Ϯ��ǟ���J�	e�z˒�2��� Ye�Iw;'�a��.n���� H�	�ȼ�ꭁ�M8
��$��~t��!ᵜٗ7H�Ѥ����ø	nE�/���L��2�7��889�8�ɗA�5�����{5p�2�6��1;L ]"f}����
&�B@��V�q��d��<ԙPB���4԰)9��<.�x�~�������Hi'�9UEx1��'3^���B��=�[z\�~&{�Y:�YYHǁ�֌�"�� ���r�폚������T<��дS
O��M��Z�;�=�=+�lG��y�)�����BԨ��5�>z��/qj_�m������vޕ�W�� �R�H`x`����"���v��ȟ�s2�.��y�U#����Q�&Zs���FҤ���CH�G���]��[���l�W�U6|B��s��-�E{�R�	�lp�s�{��<\�!�#$�ݴ��*>�elTWD��c�2��_�!�=}.�^'j$��w�7 ˍ5G�%I���p�?[����Gb[7��!ǳpa9]K��I�����h�lI���eרĿƙ��O��P	wP�k~ ֬��WPM�.~=��]*[BRwh�Q ��X�v�f��M��*�\5z�X� گ���4���8c�}5�kQ}������fO*�=nƸ�<���&*ȩzQ>W'��i��:ѯK_��Afa����^i�	�±1i������C�X���kP�i}���@����F���:-�Wa��O,�Ō��l�ux'��i�O����t�NF� �&\`XzC;�u�5�H*)���]*p9N
��b�O���6��Y�B�*��e��Q�ku<�0N
�(�@X'wH�AC�i�'i(��Y_5����J��gn{qk������z_���q8��)���+���U��u5D��oU�0-��f_`1��&-��� :�T��#YY�4�ݜ	�3
?��i�l��X}y�Ѽ���j%w/%��г:٧e���-����(6x�����-=oHW�da�b��38[ە �|��"�ZY	�M_�4��n"V�Ik�~�z��dÞl�L"��qf�t�vFq��D���^�H6�2��Np���L��e�y��ϕ�-Vr2K��7�y�l���;;Y� �r@'�e$o��,�S	:��r���&�i�]��F{ 9(�}�	�5�Bݯn�(w���r+5�Q�}�M�5���t{9�N��̀�	!,pM ��P�z7x'��{��Ú"'B��D�Zg4��W�G���0X�b*�q���ݞ�X�+�o&��X'���5��2zh����0ӄ��:��%{��a�	`y��txx�t��*�*v� ��>m�o�:U=�6��X2?�76�1�D2���})�2c1 ��!E�@k�t�s2+�R�b6&')C,�Z9�{���W C4>��iV��糑�}�(Ò�������|�@ֵ�ǳL�hC�,�G��.�r�&��Һj&�}́���F�j���.V���MNHY4{S�|��ʶ����L����#1;PT�����`~b���ҢuWݎ�R��l=^� ��5ӫƟo�P�Q��f� ����i�>~sa\�0�Wq���Yn��}��PS�ll�}V�A��_�8� �e��� X�$�]}�����,F=8j�ձzGw�f{Z����1EX9�,k�y�n�sp�4c-^oEX�X覵�vK,�E�W"Dp��]@nv�L�>��)Dټi
���I��܈:�/�'urqh���&b��	�h&i\�@ґ[�#?�8c�%��v�P����ݓ��5�[%�.z`M"�����p��/�"�\�tOj�l����;�1�s�����7�;�4�W~Q���g�u9��y<�Y���Y
C�!����U�����AS�����t���0J�?k�����Q(X�>D,��_�%�KǇ/%�`��R��������i١��\߅�M!ˆK�+x��W������N�x6bV`ȴ�gxF80���a��{kO�4���������2}�t�6�ԑa6�~@	wô`��L�[+��`.�0��v@����5�6*|M54�D���/q4�_ ��7yKOv`�W[
GkCA�?��?^��5��N�rۻk@
�ͥ��*L^�g���ǣ{��$Vt���6���L���N�	�"��fN&m�8>��㚣��+n��A?H�3Y�~O���>��h���4kx� �=t���������c��p�|�HcL�|u�Z��y�jzi��Y��1:*�`1�2F*�2���z.q�/<�*|����T�N�q��5/gJ�1:�}m`w�WM�d�����]0:-_����7F9S������O�(��p�:4�JT���u�ꣿ�C$	��DKuǎ�ߐv����͡h��k�ia�i:=u��u�i�k�6k�܄B�݁�.���i��T�Rq�.`7e���sj𽇞Bzވj��ʷ�Xo`�oi��z1��;s�g?j���@�/u��d8=1HF��f����=�1eq�_[u@�am�Ħ]�7��;C#���16>�r8n��^��ߔ��"�2h:�F�U�{���As@I��:��qh|j�q}ɽG�4(	�ͱ�P�T�}�a��]A�j�m'شR�G{�)פa�M��Hx�����D��FL"��1PW4���t.pǙ�s�`���l�0/gx&ǔ3o�9z�ԧ��,��MY!0%<EQ`���\Еw���y��={�OI��39�*��H��
'��!���jgzȫ׆��~_�+����j/7$'��J-��V#L��jy�`S���APW��/�����O4�݋�J�>�z�#�\.����6��,��k/�6�y7>�LS�D���髒��̈�6���ņ��kEtX���:N���z4X�
>o�Lc&7�:A����z9�a.f��|��0���Ե������i��N����E��r"ʲ�T�%�P��b�һ乩I�
.`�HYo=JJ86��٘(�Bp����Y�aB�wh%�pF`s%����&\^����?"I��X�QG�t���7����2gt�����va�-S*64�Ǥ�h.�ܸ��ZջR]s���W���i������{��K��`\�?FZ�䑞l�m�4x��<"� h����ZY�>e%3j��;��,
����`�H�;?E��g� �=��NL�;\��b��K�q��a�~�.�<c��R�Sak���ix���؟�I/���0ղLt?1�y�O�
�� �>۰�a�1rQ�׮���Џ.əc��,�O`ɣ��H�Og2�@���!���$�X?��E�M���8	�"�/Y^c�MÖ�_�Ix�YH{W���2RrkrKx钢3#M�;�$����1�p��&s���*d��&&E�d�qs퍇�fC�N��üx��� ���Κ�^ƙB�Q�LX˵�:^0�e��`��s���>���TΞ�Fv<_�ʯ�~�(99gѨ
�;{x1�Bq��D;;�{��[�5y3%a�	z����騛�r&�0�:&�_1��H��o����RO\�-�j����Z�W	� }׺�-8��)]Gra�:U_Ӫ����Aׇ0<��0l2X9�b�иN��c�R�˒���g�A4��!	���E�؛�V�=��zL%�������M���<[
�H#K�K�8���<�umn��x*��q�Q
�,����]_��Q`+�/��ԗT�S�@��4��ߙ����)H6M+
�f���Z!�G՝i����s����R���y�]��Όc��Sc�5�K�.=�k����
��l�ݑ��J��D���8���&sxI�Pe�c�t+��!a�'cvg���Y��"�A.����RuR��e�����߄)d�zG��>�n�O]���Aǆب�|�,ew0��	8�+ۄ��9#�9izn�� �D���4;4!�M�' �W�D�ޚ8tAM�oI}tZ��W[��)k~�]�k�DW�9�K~c=2@�v���5X -���7�즨n�oDY���y`hw�	�m9��}	ڷ�M4�{
����4�$��cV�Ҷ�\ǹ���5	�J�}�����jy����/��a6��EB��a�_68z�q0��Nmwb{����#A��Si��=�Ӣ��A#H?����*�k�s�^���od����LP��r����U��kTYB�������ִ~g�h;o���i�
�<���YP3�D�w_�;PO��Rbe��8�J�"ω��`�~2��V�P4�
d����yvDOš�&�'Nܰ<����Zt�S�c _ps^���~������Q>����l�zvyȏI,���Ĺϼ�[��+,1�{�f��O7�!B2YY�z� sU��Q�r8h��{�? �t���s$��T�w.��1'�8l5Z=�2k�J�#5yR��10>��,(�#�c~� h�I�Ks
c4=R�땽��q����lX+Y.=0��3����%5c��1�4��#G*ъe�<��$��<�h�;�����ɡ��xt��V_f�m�;��
�����id+�}���E��N���~!�t�w_�QAVb]&꼞������%�X}:L\�7�q���������5ͫcbA���i��#��uT�ُ5�{jŶ� ��҂�=aK��4x)�U���"V�n�I=R�vM&���7�h��<�%�_�;Z5>��Ac ��Z#Np��%D���}ze��E-�d,�Ħ�V���೰B�y�L�J��j��14�7*P�_0u�7�LG�#��*& P��~�H��i��<���t}����@���X��xA�a.c�?��8�;!uiB���x��)YR(n�~?Q� �P�F��t�ɲ\�t���C��S��b�S�/ 8�z�O_����)7��H�s��a��xਠ���~f��++%E�8�F�B����"ؤl#�I�>3Z��5WB��Fr[	O�-��-�B�J�Qׯ�w�D;���p{���;����b�Bf��|�2�&�k!(u�C<ɰ�����c�X\��{ ��;"���AUa�P���_��QZuZ�Y�:+o�a�w����1�x3����hb�_�Tצ�,�Z��^��}���wb,�B��Bj��ui�n�B�Q�I?���^(R��z~H\[M��](l*��=n���І��	X��ڢ�l�:�8;��7�ZOT;(��"��Sͱw-�W��}��?AG����q����)��8>���'�Y��ڈ�H��k_;ɝ$�7ɹ%Y�'�k�=>����($���,U�2X=�$���p�]<��~ሪ#d��/r�Q�OOR�)�ha��^IeU���C8@�h���y� v�*	W���RN�{:��	�1|��%O���[	�eV�I��܇�k�8q��u��_�tMAH�+6��vM ��5*t�,	GJ�0�P��c��.r�������\n�x�4wC�:iP��c�]��>����_>��Hb�2����Q�����|�)���uO0������M�6�*��n̗+����DP����r�#����v<�a~I>%Ź6���3�	,6vi������l��F����ح����c�T=�B�H�u�[�
aS��|�H��y�S���D��M��x��y���0�m$j!_w��@?Ș*8JǼ����ЊP�uD�����"�/տ�h�?�����η�6�����WUZj