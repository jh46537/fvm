��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�3J1E��Qe����ε��@E�T�R��� A��� ��i]�Dѝ��^���&{���{�5M-���|#:v${?G�?�'��g�qtw����+�ν?v��㴪[rm�)z���E?��?�U�p��7������t��J4�Ԑ�=1d���`j�ʈƎ�L���S����ľyuY@�Ol��l��������&'�<��Z��
;���?���I�R�*�l���2cܳ������dJ�\5�H��H�O�a��@��2���^�.C.���g�2��s7C�`�໮4(r2R�Sְ5�v)6�3-�n<�l�X�&��Y��e���Inܿ85�fݯ8�Ȁ7�n�`Y7L��uv��^{)�$1c	�z@C
X�q��.v���na�4�cy�-�4�`.��Y<�;�Ǜ���i�osy�84A���H�Z:�#�d�ꏠX��~��1
sbM�U2�Ŕ���&�1+�2�QHi<��O%�//��_�e�7z��G@���//b�X�UT޲}\�Ybb��2�C:�GP�6XV,񎗻��8_�.Ǐ���/��/�M��5lX�tʐ��:Ɛ��GQ�Ju�u�Z
���J���HԻ��l��^a �$
\N�#-�J	���Eԇ�FeZ~`^*V�|#=��F��y�~H�vyK !/�.�)����F�/eAެm,� ����\��Ta��Y�B������\h"�����0R�=��Mw�vVyˮ��Ԑ�)���#�r���L|@�����@'I���&���+@�2N;e����6�p�sW�0Szo"��C�y"\�p�#wK�8s{��7NB^I`�)]4���[��a� ��ތ��ש����1�>y{�"i�D}���+�4���6h:��^�ˋTwo�a��.织��<_�Y9�5��qxt^ިg� ��1��a/6+����)�0�_�U�:| ��%��c!`)d����F�Y���bgJ,d��M��_��C���<�;���X��d���ǋS��LN�
Iut�mW��c_�15�r�DU�#m�r�A�Mj�Ѷ�����K�J]�b�y!t`�p�jv�Og�9�Hַ��'kSR5_�^Q�>� �X���	������#�0Q��?goFhd�NS��)�z7��}�[}	����_��'E�y�ٍ�m�M�ź[�g]%�펀�A�T�D�<���{3Ў$�Wo�1�N3��vJ�ۛMG�3����6��7Ӱ��/<\�����Sw��/�>�]�-41��^����9j<�_��p%/V0�7_��b��56h�����LGo��&��_z��l/V�w���OGd����I�$�f�˚-�"ѧ�+�=Uz��'"��? 7�V;���;jZ���P�,�K���@�_�/��g��U�;� ��sR�R�F�!
�o�z�P��w��Ȑ��E
�C����
���/n�ǅ��Y�:�������G��3�0{��ª�_l*7>6�������k�c���QU�G�:L��ju� �PƳm�b�r�����n���h�I�#d��~�ȿEƖO=r$��ګ؟6�{q�-3������u]FN6�X���e���ֲ������WldX�W��5��?�����
�,yQf�֬��4�`�A��F��VA��Q	bư��}B'�G���f�c8��J�ޥ+E`�R����9��#p�b3��BjX��mXm�:������bk�z�����y+m.(���g��@����'�����pjo��
�f��瑎'!�s�L�>,|�<��X�M�E�R1����D��n�@9!�]8����'R��$c�C���Qi����ot�m���24��z�A�ƴ��>��^�l�(`d�5�v�pm]���A�3�Խ6�%����R��+_���i�a#0֕��f�C����[�cJ��1�|��ua]�Ffge�&:�q�۱��FP�rC�7TFIJ���J��ч��r���喢��{FU[��6�*�������{�,1����¬����y�׫H4��;���a��(��p�����AE�2�Ϫٺ���T�t�.�o������j����������9Eh:������.��M����_B��d��G�����v~�<֨�N��@Y��"*�c�
��t��D���4���W�����3x���īi�=�zmX�w�,��a�X1p]�lv����2}�� >a��pV!��yb��B������ȧ�)c�5S���~{�,s�%��0mi�}C�+3׃���e\�ԫ}��>���3�ܮ�\B����?�0��Զ­�΃~}A�|�L࣓�M����F�~@9Ig	J�0H͠��4�M�d�7��R�l�
�#�ZL���	����x~��iN��&�-�Z�2}cϤrW�E��#d�����'B�C�X��+"n�{�&�^��]�ƥA��Eu�%is��w�$̙z�X�F~�s�IZ���nB�s��1.���Y�;4��D��P��"�q�G0��Z����8���q쓉�C�ǀ���*�� Uێ4A�!x[TpJ������?�a�`�'rG[$�
�W�^"~���`����1PS{�١p�N �g���
����ud��ΩU�O��#�����[����+����H�b}�*�{]
%�V�8�7�&0���?��m��E��,Mp��i~e:ͲB͉v�KQ�S�e']�+����D
�K�<b�
_�\!���8�QX�J]���1�qXTp]��ǃ��N�56�AQhd�Î�պ{�;v��s�������{�lG�QL���f�Q�=y�t
�w-�P�\޷���͙�W{p�bp�	���&=�:�us�w��?¶IR&ְJ^�bҤ܀K������χx �:]d
���m&K.8�{���z&^6� ��|
(G���ob��9!�ra��?ܚ�����f#4d�4W�w%^�	�e�i1��+d:ŹY#s���BSܦM�8%�{S]�l��GAB�0�
`����v���� 5i����T@�n�I��Z��t���j_\:��w"=C5X�ra����o��F�#�}��9ł`h۽���dk(�>k��0��hD1�O���yk76�X���������'�nX�/]#�l��أ�*�a�k�d�"`ǜb��(N5�.`&{��Ɓ���#�HF.:��
�b����*�B�
p(���O�S ,_�ќ��;�a�T�jϾE�|���0��?�N����������}� �� ����ם܍O�{�'�K����<����A���[mZ�,ڦ�&�ޙ�-�1%�
XMV�SG��_�T>SH�6����	�|6 �h���z����}4����9�~[I���J���]��g��qJ��`�� 'b���j�_��Д�#�1�~6�9��$�7���׹��*��?�n���Ԁ
�o6(v}%��h{��a�b�k���I���):���6"��c�Fk��ÑS��Vц��mi���=GiE̚9���#S.��ʴ�yV�䇩�,�!��Tư6�����Nf�&��3��5F��8�OJf�ebn�ˉ��6<
gXY��jo>ZyO1�;�6�0���Е��$����H�!�|镤/eeL��nG�����JK
̾ľTr��$�p
7�G	��7�¾m�Q�ֺ�<��
I��2KUo��P0��>���/�|v��dA*]�<@´I�/`�����_��}�11���E�<J(������YZ���Ǖ�zBA��"��;R�:C�#]�q�7�9
h�QE�)�Q:BN*�UD��sl��#���k��
�:;a\�^ �mЅ�=�]�2�hU����F��]�x�vV��}���_��g�׀��J�b�����k
v��j�.͎m�X������U�w��ڭ�Z�����Ǳ"Sь�ɚ 3��>�٪��u8O��l_4@�:��&�ܠ�u��m`�;+�.ԑPW��HK*�%�A��3B�TH��W�kM:�R�?N����=w��㓸xQmciR\��M����t+�W�����4�xSm5��s�e<(@i�-������疴�Z��=����/���"8�Z�-1���<ʩ�j���s@%؀�L��"�J*�}�K[_�Md�p��@���l�?	��D*�&�����R��=��/JSo�(�;	��N4��V����~n0��CTO������<)�?��\Қdx4����>�CH?8S����L�rͲb�o"ٓ��q+>
�o4���`L�'�gu�8@����!��H��8��ﳈ��2E��|G��=A=���u�\����m���[�<5��^�QD�#<$��h�o����u�*h��uj�+���[���(J�o����X�9�h��}q��:��>�Y�#�v;����HD����]۾�b�pU8'����j���s�8��Z��n�2d�>KF�T�X֜]Dm�3>���?Z�v@4�ĸ���XX"���t��E�����=� 
@�������۪-�.MJ^|f	�"A4��t�,��<�%�} ��ѻ2zd;�_:3���E�ƴ ��5�/�</B<��j^��j"�ަ�|Ź��1�)����K�C;N�Ps���u���]O�s~�l�����6��v���ގ�޳��G���h|&_}�ƣ�}`���=l!�jBj�-��n��KN�����a�TE�A����$k�UH�t���;;Ә]o�_)�C�L�M��Ȯut��{��=�ڄ�T��U��P�h��7�H�|#�@����~_.��7�)���.d�!(�͙3���F�(�}�P����8u�Y�T�.��s�T����t,�0�ueԺp�$�
:_Gq��p,�p��f����\y���y$�l�C�M�h#��xb~^���8�У1� �t�TE��La5�_��(%參'�|}�ٗh�Ⱙ�YY�w�t?�K�^�����g��
H�>�x���y���ȿ�L�D,���rQ��Л�����S1�O���.���4�W����9_*H�{ܴ�&CCU�G5�m��`�2uE�)␫L���)�1_M�����@�bFH)M�G>�@��'����11�6���z�BD8�7���;��v��E9n
��cj�����W�V�x��$���5�m&��G�f[ur�B���O���3�1�t�������Ӓ�1�b���y��]`�0I��uv]bg.gb�׎H?��D��h��s���N�G��,�>
���wv��MTdt���ަ�6���uDLy�jxf�y_�!�-���}�^�NM��7�"d��u[�hVg�N�^�����sC�?�۸�u
��]�e3&r��t���(ŋt̮Ƚ��75�	ͽ0f:h|��Po.I�!��bxLz��ū�+��&j�	�ɧL���d���K�����؟ԅ�� {��
<~��S���5����7�Ş������š�,��_g�:��I����D��֮�ê�@%3�8*�~1t�O��Ϣ�-)�Jw��c��·!���`a����ٽ��So�3FL�r�5m�d�:�ʱ()�=x�3!�o�%��~�����D�qq�A:A�+���ς*�ߘ�g�������!�zZP��&��콆�N����I�10�W�$/��@^�1����A��}�&��7\��>�-gS�Z0�Z1n_})�����Nϱ���^�?�E�� ��*=�;V֙�*?�ִ�Snl��&K�������-�f?pWx|���!U�)�޵�=,)�
Uv��mq�>�I�M�5���q�lZ��I��j2��f�zJ}��qH�POsz�d���	|�������3y�9��p�=����"��"���5츷�/u-Y	R�;�>-M ��!'��G�z^�hU%@ˌ����*}rR�w_R�Ї}�1�}����w /���������\	ښz�G�� ��#�T�Я7e3�i�ZZ���H��J�����'��5v��)�]x��]��[�f��L4���Y�l�?��F����?�kF^xt�a�B@�Rg����DĞ�JJF��`]펏T�h?��vz�qXm�5�Gw$�ǅ�3���C�!�����8���\�@~���]<��
��P��O��^��R?���z�,xQ��%4oQ��d��E5#�������yf2��i��Fq	it���L�V&SOu�?h��D�e�Y	����NF!�p�B`�����Vs�y��PB�l
ڟ�;�N�=����bd<ֻq���}���B:p�	�uz����'6�$}�!(�����+��
>�TJfy�A4���2�0C%2�x��,�/�¹�N�?��A7Ē�:�4�"��:n�����֘/������8��k���_���C�������#U�逝�>�6�ut��f4��=�������w3���4��b�}�CKhټ@q4x8!�2��$\�!�~���Z�����p�g�$Ύn��>�g�[\����5M3ˣ�g�bK� ��7��m�=��A�;A�㕱`D$K!A.��h���X��t�'��P�i��HM,
�p��Żo;�t�{ޤ���B���|��J�������$G����-� ����_��X�W�Ut�XF�3�0���=ۨԌ��"w.������'�e�l%f@����SF�٩f:����A��v�����c�=�c�r�3
���o.�Ci��i�}�%�f��#�?{��ϫ��&�����nS�E�K �c^�+��M`������
ns0̽�=]6l�eug�!��m�j� �=x��v��΂��eo�M)?�Y5ь.k���Q�;�̿Q�D�����\� [ڎqW�E�h�n�+��SYn&�?Z���}�q��i��}X�[n������E�p��d��S���/�)70��1t���M��g��8�!KA���د��Ϝ6�f�Ce�;��]���s��w�p�:PA ����2
�h���J�1<��<�f-h����s<�'^p�z��ř�;:U��1Rq�����b8�q�N���H8t����؃����M�X��:L��p�<g-v��ʧ@��g��@@ڍ���Æk�D�<�)�["HGh����e9� f;� �N�܃i�\(���J���W:æ_r��@.2a� �1��zv��. ��<�\�+/�/��u��>����L���'�b�%0Y2\��or�S�6�H�Ҧ������<6EX�RZ��{J˫���4!���ַ�DupT�E���$A��2����D{����Ӂ$����ݘK��<-�*�� ��Ca�^I�Ĭٚ��Ωg�q�J��Y�3����>��Mh�jQ�Z�Q�c>��0��G�w���D�>�L��u�3��ak�������N�E�:��[I}���j��hF����H
+���D�u���z����ʥM�e��_4r_�~�2S�X��v�x�l��7�"�:v����,!z|�O�*H���V�%ֵ�����`�k�ž� G���܇9�k%��6ѯ�8#�q9��c������-�S��'HEX�Za�c�s����M *Q�'Lc
L�1�� G�i}�&`�X>S�,�%-m=���h��Y�N�<�ṙ�Z��R�����)p ����L��(D��,E����h�����e ;��Αq�����	^�o�n���(wJ,lr�X�v��D�IS�DGlv>|�i��kw�>H߂��m�ǛG'�� 1� ջy8���t�*��Wϻ׷4��1\�� ]QEך�-��0e��U�-�dk�&����3{�O��}��@p��+v��CڜJ����GAd$M�=�́;;�Z��i���66�R��}�J��g�7�P�p&��m{a|8n�����v�������4*մ�5�ǌ�x+ĳ��
�i�x8N�ÏVȈL���<�4-bQx�\�+��>'?؃PD6}�I�}@�p�Qħ}I [E�m���#Ϊ갳��e������f�|3��9H��Wi����Ӄ��nыA�$���{�Ӊ�h�ގD#ܜ)�œ��'5��=ߚ?:mX���X��/�%�D
_����t<T�S,GZ�{?�(ƛq�Bwđ�y��ʢf�����wLZ���n� )z� ����pA^����Q1�a��\��9�Q�yOb����0��E��'� ��N>����3�x� SQyi��sK��Œ0ֽ5E]{����92|B���ۛq�dV�%{�N��og䳃-�e�8��0�B�N6]I��B($�TM<>l�߰FA�2���yiQ�pc���?gT�0���+�P�׿q1��H��������s�Y�,��B�W2����d;�[��gG�fZ�VZ@��z�d�$Y�&v'�ӭ)K����(Gnrq6�1 9�t���%�����)aǴ� ʳ7�s����h�@�a�v�̢o��������u}���y�E^���.(&-Bƙ����/���| A�`Zl�B�t�L,~����p퍥1�r�\�#�	`L]�W���1����>��*J���^�g����Iq��J�'~�!�v7��J*��I0�*�*�g�^��Ub���oOPt0�������($�,��I�I��g��<2���^�#�>���â|�3D�������I��qa\�hy���̨��+�3d�����E*9��P���Io�,o�ɴ�m~�ћ'K`.�"�v]X����1�g��	�Ti��ػ��8�Ǣ�h�����Ww|>��w�'/�3ݻ��(i�X��ٍp�0�4)���7ɖ�vi��j��s[,lM�NdD�n��Y����_sNƠ��3Ni��A����/���`����(�D���ss;����1��*�QiY�;T_0�+�Ǩ�Ia���=��d���9<�CV�~
���L��~}M}B�Fkw @��^��71j�!�ֈ�iv�z�#��ɵ����܇N����<H_U�Gڮ'��Ƌ��u���f�a��3_��ֻk��V^���=*��&H
?4L�P�Lo>��"��\P���q ߎ�浕vʺc��)?b�"(VK@�K.�4�� �p�hZ��!w{���2�N���W%{v��뜴´6ʻ�`���e�a���tKQ
du����H�Ǖ�ٷ�śc�����=s2b ���r�a��=�ׅj�Ey[&�f0���`��.v�|�#]{Fx@-�2���*�f��g����w7�m���ۺ%�>�{;ۯam�[������Qu:0-�=Iċ:Er�b(��LX~RH�T{n�ĳ;�0����uP	2C*γ��)�K⋗�5	��B�Q�?������v�i0��jw���c�����v���DoK>�_�jX�k��fu�l�n��/�j��ٖ�����"�a�7B1?��}=߭a��c0tP��4�C$�U��O�xYd	/����d��Y���G�o���6�Y.����3�o{b|ш�X��&wm��˼�Q��M��Ku�A{㨜�q� IIt��>R2�tSO�Y����sX�Y�k�6(}Uj�~`ÆeX��J6���6I9ĉ\�ޝ@��b�\�q]GG_M?��I�7lPOvM�(�����L��FI���dP�=����(�/\�m���:�.�\�Ș����@�JEHK�[UJ�f�tb�j2mO�y��.	���y��.�������I�i�^Q�>���ҩ�ў����%�qc�?	�. �멺�����;#��Z8��KC��<-4BK8�?�"9���<(��M��7p%�.lhٻ<�w�%<�_@�έ�$x����ѝ2�9jp�J�B<bN�j?K Xψ����+�����Ngu�lT����l�Hp����u�#�ٝSӤ��`d��Ѥ��)F����?���4'�!����7���`�0����n5�}`[�ep��>\�X	�@ȕ���Q��e��|��i�/�s�W>������(�瞮a�M����m݈j,��p����Z��<�U���ż0��6ےX����V�i�%|�eC$)��ہ���_�䬍��w:�TZ��8����0�#�K�d�5�q3jo{z��`���CZm˚0���D�q�u�gW't%* ��1��.�p=��Mp������X�cW�祀:T�:�\T�5Ճ&��	�p��2����5���j�o�7E�4�<5�F��������[��n7�z�nZ$틣FU�=L @�����
����T�,b�c�7�T���vX�Դ����|pY������!��N�/^�9��G)��f{��q[�gz�=��h�|�w�_��
fqޖԔg�n�)��xINf�P��+,}��,E�݀�7����7����� [Se�u̔tڅ��jt>�A:<�	�S��*�I��J�C;��uww���~9Jd6ӟ���И�����}}#���5;wU���R�4�3Ԟ�m��tnE&d��~�H�l�3|"��(F��E8S�?��}Jz�����n�Rʒ�7+�tq�MFpC�W��==����bb�