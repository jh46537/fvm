��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK�����i����Y[b�����߭4�lFHi2RC�#WK���"�1��"�
�\�0������>W��
�7�(�C��I����T��m@��z���p�4� Ý�O�D��i)�k`�3���D� T0��)'��H+N�^�6��%�:�z�?�{g�Y=��Rf3%����(�c(�Q��S�2~{��M�o���@A3��;n���c�fS�cӁ����	�da��D��ݱڬܞ�_��߳g�q˞�N����s�~E�6�W�l�2���B��V!)/��m�h�����*!ʧ4�+��R�Ï�A�J��w�eH��C[�|��7��t�V,���t�;[�:A4B}/}x��DmH	�U�@g�����_���� ��R�?�0�Qy��մJ���ZB�dfj��o�.	�"�N˘���������sZ�.Ҧ`�y|#�ֶ==�Y���4|H�+y��	CD���,�J[�4� Fj�Wqs"�o��9�'բ9�'r���L�#B���|{}��?U�~<��JA�O ^���M�����вq.�����rCL:�v�y���l���A��?����*�[��;$�	��������"g��3Rx��x������B�V�و$F��f��w .�h�� �琰���V�������9��|nj�U���ت�0��D�P�mY���X��4���::�JN�f]n˘����y8��Ae���ۛ x��bŞ�!�&��8D���!ڕ���!�ΐ���n����Ի����b�b0-��|	�P�+.�@H�
�~*ڸw] k�W��@M-�u!�rs��O��&9���-�`7�Nw���aMB�Ă�3���A�,'�8΃]�"��/cP����4�K1� `E�@
<�����2א/�Υ���|L��������no^�QGHAˑŏ�O��c�\���>�@gN��^���ۂ��)�zG:&�t�%�~`6y���>�ަO�ľ|�F�?,�� 	:A��ҁ��8�q&%}���n�s5S[Uϩ��] t6����}E������"�j�u��Eȟ����>�/���cr�y���J��Gvˣ(Y�UjGJ{"`�s]~�V:�)j�D=>SID�v����,H�R܉�c_9|ɶ?�P���D�(�vR��Q�&̎�T�D2~��]�%4���&�%�Bu%�3������d�J��x6Å^'Pɫ��y�A;�6�H�XN0�24^������e-n����ly�?|'2~ԡ�:��2{��z�J�����3zrFY���	����wp�&O���E���P
�2h{�kn�b!Tw"5��K��a�n�P�f9�Y�,O"AøT�D撒8?���wOl�&	N�2u 1�f����!~@U�ߠZ��H�U���)ZO�ƠAm1j�1�������t7�gZ��M�aTb%"�U?�Z�.	]��<�-+A��� ����|��6?$�n�JB �"Z��W΢I���
q��iقÚU}�M)��X��f@��*�� 1�O,4�C#�IN���&F��T�T%o�{�Lc�*W���1=+:@&���ژ ��0��W�Ŏ<V/�Ɗ�3��y�{�R�";}ZbQ�TV
�BV��	ZV�� ���m�L��������.4�OpG{����u�IeS�m���7��_��s�s����Sx��2GW!5����%�~%���u��UO����RnW�Q�h�*"Z�u�P��F��&�J��u�5�$�f�=c[6^/�����(��ygL��#���Ckjoxi7��C3r��Q���	$�×�;��2}�Yqw��$�Y�~�F��{"��V�HXp�������{�R���pm�=c���$��#2���T�@�NC9���#��n�t�(�ę�#��^7ǹ̈́����p�1k��V`�:j(,X�@yp]$��_��1�`aǍ`�~�!�p6�a��k�l_m4|�����U�{H�e:Q]�g.��i���+�3L2��أ��T^E�-Oy�+&0w��Ecl%�B����l�V���E�P�!�Yn`yw���A/��x�2,���6]�V,�&���h?���C�m�65Y�EbM�ϋkkƞ�����2�V��Ej|�)-ZՐ��)�.K�N�j�ޏ/��Z�U\��]�$nd{�)�B�a���ك���Ƥ��{�i?�9����%i��i��@̒e�v4��9q���]����Bq=�s[��en�q�~w���N��7�>����⤞<����ԳG�F������pyl���F���޼��8�Uq_���"nYǆ�Gg����L��T���8e>���:�Z3�غ�yn��2��R�h�,;k������.ã�-��X�h/��=g����PM%�FYU�A ��y؝Mw�]S�8���4�Q�K�L�#��?���5��9P�AE�����֒���5,��FQog�⠧��'��A��2��&;9�$Է��iI��>�[4�{�㖣�M��+������l0`���V=����&Y������y>�)�d��x���N�!����*���@��ݣn��eāE�N��-��H�������A���K9�Z;��\��+��J��}w��#��Z�5���LɑC��V�������y�[��lsH�	4�� �H��F��)0�|��Y����[��! � ���@����w)P�����&�÷qOR�]9=i.��4��]NK1^����=�
��K3��Zqs`��R����p<��d�&MU�>���rPn���2ֿ��@C
$	N\A������ҴJHeZ���t�
�r�}A��D���/�+�����R@�}a�7�+x�M�k���c�gÇO�F5�J(=�_銬"H2k>���Gy�V��^��A紾��;�gY�d/<�eÏ'���0�Q���~�#X@�&�'���� �4��M� a�f	��}d�&./�{��5�̝�Xb�T�u�C��SWS�V�n)��ڞ�o�T�ר����.�l�ws�?�U�����cJfy:}2�0�%F9�X�<e����Kg8r�8θ���A>$��uU�r� ��MZ,��z�����T'>����L�̴$��S��s��|���2�o׵��
5B�]a-8�.&cjǠ��̀�3���U҆o&�|��vE��A��'9 �Ӄ��čG��8q�a@)�,f$Q�v��|.\�����'�y�?6�������{��O� �:�=b�ZS֔y�
w��.�mu�S��HH�M�׹x}��%�<VwROE�����<��8n��AJ|
@�TK#�֧ɺ�7�.��z����|Fug8�ae8��n�sf��)�\I�ދُJ8�s�|7=1?LY����K{�w=�O�zn�g���Q0ǎ�Ď^r��ɐ��������ư�2\��a�;����5{���+�Sx�p�ܚS+5�����C��@`x��l�L�Y�jTX��v:9�����]٩�<:3��<�8���c�0�����]�zb�%���n�a]�G��x�b� CV���l��+49���D��!wX�G�Ö ���GzYoJ����������׻
�����)�Z�w��k�vP )glc��d��w�6[!�������uh����׌w�g�}��9#%���y�e-_a
�ܕ�����ff*y�s�z:G�'���"��s�0�I)TGN7+�	���-�X��w�\���FN�H�V��}/Up��g�\P_%����V���t�����-�c�`��K���R=� ��q��YNW�:d4��빦�a��|r��nS[~y��n򔍔I�
��);v7�H��g�^b )թ�#��I���~�t��妽^c}�u34 '���i	���cX9��p�sS�k����x֊�"�d���B�-�$v>G��oJ&>�$��'x����+��vr����(u�N�>�=-h�_�3�u�W>�%k+/�+v�}�����-�H�{�gb��@�y�|��f��9�@�'�r���e3����Ԃd����O%:t|��3�����%�D�} G��UQ��/-�i?�h�:�z&-�O�O��cl���_���]>��b�	��B��g�����mY��JIG�P�;�ȡ��O`s��Q��A��R� �w��?z����;�p�HnX�b�� �^㿇%1�PbªH�%h�)�@�[fi33�z����t��=�C�7�o���3��'=6���[
4�U�MN�Q��m�!���[��F_�(+zt.ﲷ�s'�؛�xD�@ 4jS��wo�75e���ɇd����ͭ�ss��D��Y`FXz��� �4;�]K��,�Hwo���pQ������J
v������:�C]�#�n뉱!3�6��p6o�S�%U����p�_�1�"�P�1"��uI�q��~o�S~�ЋG6�P����CIw�6]Me8��W�DƯ;�2v��6e�:�r1�/;�:ٵ
�
EH�o?M�)tz8k��ˌ��r�G�Hq��4�ά��	V�2��~���������	�Ā�r���T�%�l���_ֺr���,u�Y��`.��2lD�NbHfb#�(���"�ؙ���>���o�L{�,�G��p�6��Q�af��q�;k�9|��^MCS2�eq�3[�ՠ�B"���6�����/ I��J��V�O��*Џ*6�?/�i��
�V�Op���CoKDMFVY�J�������|�	�talh1yK%�B����� ���'���3�1Z7���qU5$�
��9��[-x�1S�B@1�r��	���t.�tƕ7�
���L�����ַ�V��%x�cʽ[t&[M���TuE�ه)��qF�6�Z�1��RDO����,��Dh��4�&N�O1\p������w��&@��{ ��f�C#�h�V������W�֘�e��_} ;Ŀ�3�e�EԹ�s��䪋����S��U�JҴ{�*���Ybҧɖ��7�1������k�l��
Kr�P�<7�T�cFK�M~��p��$Da����B�|hճ��g��N1��s&MXV��w�Q\�3�=}嵻�W-N���̸�OUڬ�$����W�ц?��&�@�M�J~������&$��Kg<|'Զ��ъ�T���o�k���}0�Xo%h�-����wp������O�󥏼\Ze>�GW����d��L�2���~��:���f�RZ2R�K%G!Li��nv�����z��������4�l������L(B^:`���VJ�睟�p�v�ۍl��7ZIP��q-� ��v^+���e��D~�2�sl?x;�CG�q�?�������
'�y�е��=�o��l�.�2Ѩ�����g�x��y$'�J{^��5�d�]{�i�@����o��0D��&�.�c׈���Ma��c��|��1)������t����q�A�Ǩ��|6�<T�>�����FD�r��圧��k�Ǹ�=�����!@���5���d���]0_�����oM��7��q������N	p%tD%3R4ۉ84#<��y�{�G�"u�{o���q�nH�P���ן�a�ƛ8o�� �>Ɨ�|%��}���_�1�`�H��B�kt��}��z��R�@j�O@��i;LB�ˊb��e��s8�ҍ��H��y{������z�c�	���7�_�G&Cx���������G��X���k��!�ʟ2��H~M|����E��#�s�il>�7�x���	c�_7��BRȡ��>r�UZ������s�*Ӧ.�D���j mN�4HO�����i9�ƛ# %{:;OI�$��w����M 4�*o�~ou��7b�h'�Q�C�$G�x�K����=�Q�3�����xꜻnը4�Z�G�}�k.�;w='�e��BFWfҩm�]Y�H8����B��&��= a@!U�!���8��@���3DQ1ݭ[(e�����q�v�Ů��Ǽ���74,׳X�xT�����ݲ�F/F���/;$y4��A�������7�Ǯ�-׫BVk��A��4��B>�)_%0��{�ʭ�O%7ӫ|�v�Y�C�E�����{-/�I���t�"������:��&�)����n��Y�
�pu����}O�gP�V�+��̋~��\}�zg@��3�ɞr7�m�w�����&��i�,ͫs�p���r�
�2T�,��v���i���~{�|��Gp`��L�{�Ae+S�bL�&���}�0)���k-R���=M-k��3io���Ѧ���Oڻ�\���;��!K�&&���bw��ʄ�����,���H~d~M�g�#�+ߚ�g�`��r
,�z���dx�g�����#	�+���%�[�p��"7"� <�KӖ����~�nwZmE�W�J@{�qF�'+�A�"~2�w�9�!j�kRo4��T�v�UG�՗W���h꼴T��ڍΑ.�4,ޱt��1[��/}����P^[~��\����^˷������.�t�h n4��-'�MK��)�hfAWι����٥I��#����s�]�z����@[ul��z���\�M�P�U��BΌ�:#O���g����}�f���h
�0E��'b,����iə�|��(B��~��e�q;-��-j�4�"��x�&�ηC &��RF�<ꤖVC���?C�QGՃ�t�X-����gg�R	��
%}�3\KR6v�d)Ԉ�� �7��=��Cq���: 1X����mZ�%�q���=�5<�:ɚ,�L.A�lƭ�[�3c$�h�`J���W�y���s�h�L����{�N Ǜi���cƵX��q��A;���9iw���Q�V�@	���� \�ք�o�jw'	�,�m����� �ހ�z��I&�?����s�Ʀ���2�����F��T1�w%�)<�4���j�l�\׺.��J9S
�u����m��|�5�[���~�7��9��
�
�R
�9<�2�O�����{��y���zI�O�燑U;/i�S���"l?�"���5GF��fA>�?�����!��ABIuu�0� �(�8���瑭�;�͑���U[�?t��?�c2���Smb.ϋSn��=�\��ث��q�q��4ɨ�Q1Nʊ0A��] ����w�@ܻN�hW�(�u�|%�u��z��Ҹ2B�;켩�ӹ��c�/ �k�?bU�à���DaD���}�r47
����Qp�s>� ˏ�id[A�njmU�9O�ȯj�hZ��[gs-�D��<�Y%��%&nQr!*�.x��<�q�Õ�h���n=��?��C�ꋟ�ί�;�����j��x����b�|�w���r�\�d�(�bo�pB]T� kd	4��Ȇ�mr��oͰ��^j�����=5���} Mp�e���̹jl��r���l�pge@f	��~�[�2�"7\���(�H��D��� ̀ٚ� ��OV~2NP	G��VU���5Q_�Lc�}���r����"%��JˎM�Ok�"�zz���3��݊A�����kMs�;cȌ�2�R�R���b�|�5�|#�
+�A�4w�z�$�}Gao�����>��b��T��ގ��9�"[�Ud�sx#���@`�gO����A2�V6B�7I&F�:>!���6#rv�5�d�6���/�i����I�.+�:ex�y����{��;`p��.����)�
d���[+�{�X!�F0yo�J_�B�Z,$q3�O����4�]�`�%����G\u�,�����ř���Zʹ �3V1�K	���¯h��2���lP�e�N�x����3z$��V�:�5P���o�\���7�@
���$^	�ϒ.�=Z(�"�Mub8�`z����#��{{��MX�����逷c�$MU�<�cFi$���ȑ����8��r� �چG��}�����F�i/���β�E��5��01�J�=���k�Of����n��ΐG�Q�֔���`rZI�����#�|�����S
h�&#drh���rK,�q���B��*!� ��3UI}�S�2.f�6�7E�0���d?�u/�V��򏟞O=�Qv`d��P�\�&��^P����������7��Є� A2S�V��H�正��j��������'QG��|wby��g�0��k�4�a}e)�;�R��������̚L�O�X��UY�ߍ.�h��j��6.�O3��_�z���3�6"�aȔM���7a8�&�+�����j�<��v�\ӿ"�먹�<��Q7X���N� ���]lF�`��ᩭX�������ף^�,��4;x�W�h��m@	q�yVou-����h����-���WS"�,a��6�9��浳�E�t�3
Ntu^^Ԟ�&��@�}v��K����k[�5]��,���i��� �7��Y�����G�%@4)/�����, O��y�c�6X���>��ͨ��C�_��+
z�k�R-�K���Z`��v[�xca���P���ܦ��	����W��r�x�*�pD]��y�y�?O{Nym ��}�?Z"؍�v�С��	�n}D���"���<�Jd}�(H,%O��@OEqҭ�~G5��i��R]��e�4|�R΂=�M�h��:�l�(������N��ɖ��v/)��AQDW�

LL��E7+H=��L�����L�R�,Q��u$���H޺f����h��K��>^�Y���-!����#�N���|�Z�9�P���0r���_+�K����
��;��|�:Џk��MsנDj�|�|�@L�Ӻ�҈w���3���|��oy��T �u��P�n ��Z��1��Vm�ź���̫�kٮ��P��'�6)�K6*-,,υc��dN4��Ñ�����Q��+���<���H��꿦j��m-��l��������Ԓ�6>~aK]���+�q��c�p��(0�
o��C��l�w-G�#�s��g��wͣ���-���z,�7�,�S��*T�Db�7��&�9���F��v����V��K��&+	���a!O�c�\�|3v/�����{��u�rq]^E)��+>�l�Y�4拙�%��TNw?�8��[  W�ͥD'`���% �)X�?��?7g�y�	e��6�A���~~��V����O!b9Mm��I��^����ǖjIHؐݿ�� ������d�},�Ą[<�BB��Ӄ��x�A�c�;�*eYRQv>a��u��z���1'���Q��|����t�|�o�xh*������r����L���v�g��wݖ���_��f�3>��K�\��|s}�6,�_�@N@�:rl;�Kfd��g.;��X�k�p �g'3a��XQ>����X��R-�~Df_H��WB�b��o��&�U��2�8V�g����f���Wj)���sjB���f���)�Ѱ��@[��2ܞ�YN��c�X��^T�-`�b�T�g�tw�}zm����q˝���Ym���T�͚զ� č��ÈT���xI� .����A�����N[[�1��gU9�x��I^��~����_^u� ���]�7�T�P�@�6 p��j�B��q�l�5c���Z�M���Cƞ�♐�
A�z��p$��QTH��0��G}	�#3D"���t<�������{���
�yRd=�t��q��7�S�;�&�o�h�U�+�͆܃0�;͎�����3��y�w����G�%u��e�N�e�����?���9��w�*	ў�#	�>�tۨ+׶�O��lL�����7��c��}�X��"�`�sM����]����C#W~S���p*o��H1��2��=u�t���=�V��e��ʲX�	��u���
�7�X�r!:�&���#&���G�ª]ʥtJA�N���Ɲp �2�~n�u��s�dl+%
�ײ��{$���
P!�Ude�G6f@.'������Z��P��X�&��ث�]��5��ٮq�wYW�^�(�t�	/�z���J�{	:MV#��j%M��!���#+(��]-��)��g̍�HD�0Jˇ��mA�O�
ɔ���c�n�;�T�۹(�s,aiLNy�{���'j+�����oQ��0�AlJ/����b�!�f��;��VpNƐ�vk�\��&��g�#���j.��W@r~fݙN�N+�,̼�˺���44���U�r�?-��-'\CT	�����Zǿ��yܥ0�]�uK� �<�	�_I|�CTp�c�7��X�	�jSv�� L1�=9��vH����!6���*P@E�H3e�uЫbSI�5��s��կ01��z�P���s^�:Q�$	ɒ��^��-O����qBQT�3h��F~U-�)-<A��x���L�$zII �z�7�?97�HF�J h�59K0�[����b��Uf� ��$f6�)ê��Z��ơ��7��\���$	ᤪDn�u�ie�zHI�m�
a���|�=kU@iǹd��X{�>���՟-�ëC�I���-�d��bX��;�U�����N�go�.i����CLs����J/����m���8�O��.�C`0�i��D4*����OŬ<�TR��D�Ir��hƥ�Ĳ��}GmĆ؏���
Ӡ�Z@�_*�m
n�8��U���������Z�d�^l.��� -���}�Q>�cK��d�,w��*dXf�B�1�#��u�^�b�����¹��L�ޟ�~���<E�O��NK�����)����h��c_T�I�VK@;��zqIv����v��� e�ݴ:Va�w�s��7�ւ �8|�� 9���~Ӝ�8��9X��.�~�G)�$Ϭ�#!�t{��8�:��6n`�贈�ϗ�D�CByz��
�;�>��y��{X�~R���8�l��O�ٶ;�����#�f
)I����R��4.�@�V������<��c8PC9%	��ɦ�5\j������h4�?���/5���d��D��z�e6����v�D&@/�-B0�S*#h;�Go�jXy��T�����Π��yw�"%	"�^�Pz�>�C���l�b?}���>q�B����{�K\��𺪜�O���nF ��������)XT��������jz �)r��cM��L���Yy��rAY֥���`KtbjMp]D��z�̠����$�.mM���i�S?8L�EV����� ��������7l(�W��\c���wB3	�0ǃ�͚�Wɨ�i�ِK�l�N��{�+i�#i�p����+��V��X/2�TGT�(���T�g�\Bi-fwiO���W�w��[\�v��i�(y�^�h���6H!S�W�g�0Am(l�b@��J`��v�;I�g�s��g&?%pzY�s��ö��W�*G��<_{AϹ� ��4����U'm�nY�$Lt⏆"�S����w ��;������`�?�C)~Bb��,Cq��VXk��>RK�\
D�t
)˄w�u��F�Л?��9�~]�P����=��n�
��!9�-�MU�u� &�p��b��X��hu\���s�T0~D�3�i�1j�asJh�8��KoU����W"ZZ��h���pBrm�4�~���`�K��%.6��g���j�+�
����J��n�4HA�!*a��n��?��i�vp�#�������h�kM}�cp儦��=�0S��S���K���|�	�-�r��%��;�fī�]�����#䚸��?�����+!�zKV�cR��#t���p��� �q�e�
����j��[pԾ
8q`u�<�S@���-��O4��W\'V_��G\� ֺH��F�ssE���5���A��j\�k�q�FR� ��AJ�4u�-A4�����@kr��@u��ݟ{��g��
�n������}MǛ�zV0'�\�M���p�&ݝǃp�����K����wO|^B9e�P+�Z��];�QFCMj5��i�ؓȘ.�Ͼ����@m>4���C3�Ԅ�bnE׼$h�Nk�>��Y��ݴ���e���</���t�a.��p�{�dJ�t^���C�P�r����:_Śr3�Dޣx
ٌ�)�[���e�u��ߧ��?6-?��r�����4FNY� �:�i#�Ҙv��*h��bŵ {��=��۝I	칕'5�C+*�ؒ`,K�у���&�t,�*y�]�pH$�Ld1�A"���=�<����Sa�S��Ax|�I�4���e�α�0�F8"�&歑��IN��~�U� ��z�勰�����o{�{vʟJ��������2��&���S9�7���wL���Й�G��d�i��%��1R�����K)���n@/�t��D 8E�J$)��W'�+�Y��a�R���앩�w�î�Y"��6R����@RJ��}��nD�g���D.+s��m��hح^���`k{L�fE�<.�N��W�;�!uu6�=�Ml�,l;�?�Qa�$�3�KA/L�.�H��Z�E#S������G�}0���0 a%F�rN��	;��z��ȼ��*�����T���Y;�?�+��4����Z�y�&:�
zV7ǹ�+:�Uì�T_������%}zdW-Y�,jIH6L��0>y9�A��A#Q�7~�.�w�<0F$�w����&$��5�-
��(����RkY����6�vu<�w	� �:\N�8e
jEhna�D1���#CǏ����hi�.p����a�M�C��:LY�-�p����o;\k��<dÊ�E�SrZ$1~c�1SK��f��f�>�9�H�e��22�,��~�x�a5���?5�J���b��hn��K����L��J7b̏��j�"7>���>"�"6��J�����2O����nZ�Zw4�c���Z�o���j1�Y#�mdX��|H_����fU~e���.ب�P�re�5�-^�k4���Z���@t�ſ1mU{�D#b��3GQ$��'�<Ow]�s�7�@AC�]�8�י�M�z�B3��0��;�PO�ȲZs��g��7��k��&�	��G/O�+k����<��䈡Z�^�\EuW��h�)��eq
�+5fT��J⅟$lV�ͦ�kB��
q8���+�����a���[6�4P�F�>r�.g>	0�*A8��ݩ�4ߙS��_�&�8�+�!�qO��=���h��
��^���8[�+PZ�װ[���ď����V�0I�p�W|���xBÈX黼f�uz�~xw%R�D�l��?a�Ml���Dr���0�,��*�9N�3_z�~;��v��]��C��(8����)�DHf:лL��C,ox����~�Gd��Β.���Αv����*Nr�҄��sι��)J���|���L�[sߒ��YB�8T-��Ꞝ{hM"v�}C��'M�}��3B1��oW��D:|Ե����Y�|`�o�@�wF���>w������@�:����~-Js�C��w���%#�����
V�}�%�@�5���C�&����$���[v9�$h�k����>���_3�g��bE�erj>����E��-���*p[�i:��X��	A��*%/�|�l"�R��;�!�QsQ���,��k^����,��]x�5�^tRDO��[�Q��B�<3I����bYwa��[A}��pյ�?�m�>��ٮYǪ(�b�,�1�	�
6�_���o��}��}H<����SDg�=#�|���b '��D'͞��i��⑄MGf�8��-�����v����k�=f`�Gѣ����LF�P�%�=6K=�$�b���y�p31�]�-��?X�E ��e��y����T��D�1�`���z�|18�乺��;?�w�.3���;p{}ۅF���.#A�V��߂Ф_�j�e@ۊ̮��R}�
y�]�X4Jm{�(7"��%y�:��zD��v81)x�-%�vڤ��M~�t�s)/�,���%�������҄���u���	`����K��<��4��ט��r�GG8:�4	�#��S�;�KeZ�>D&�RՔ�<��[��nʿ�K��ȅ��	�C-�8���	j;��n�U�K;���WXf }v(5u*�q�<���K�/���H���1/n�{�3�'��x���r�𴢂��%�o��qr������ˉ��� ��qa�3��\�����?/5�!���0�w�������l��_e��Q&�p+�O���Eˎ�A�v�����aߝO�[�&���اmA�A�Y@��0rfS�x�%���_j��E�Gm�+ik��M�?��ch�=��R�/����]��T���\"��w�m�� \G���әe�u�N,��o�0��z^�Y���K�����.��N?�~��N��3�1����%�|$jG�Ӟ�]�cq�Mf�FI�"Te!V�������#�3�ǹ�5�}G�=M��J:�y"?`𔐪T�6����ߞH�9]�� n9tY\b$_�)��>�����<�p8|�uph��Ag'�R(� �i���b\�������v�Dx��q�&N)+��=�����
BE$o_|��)F2l�w���7R��������RW��&"�����.5�J��8�v�t8��Gy�&�p>�*�&m}H�S�d�3�i,�tZyxEb��D��l��z� ���l��y'�ģ����L��l%{[5�:��m�q0�@�R�@V�J�!�u^H��!��~J�|����G4��W��_+{�2a2Vl�W���#�h_X����0z%�t]�v���Q�Q����=�Z=���̚'K�Q:���Y���d�����{�M+���C��׬E�R�^F��i�l�<=����c#"EI�s@�(�	��tY��"��JBA�ޱ_�yxˏ�&���K�`���!Co��n��O
��ٴ���ot���yD�G�2�P�E!�C�O�cu��7SĖ<��I#��޼*U\K���Cr�:[����+Y�óW���4v%J��/c���������F�	�X�+Q�^GL�ō�aW�k�>�WԷ�J6L��}�^��a�Uq�{�=�N���_�K'Y��ո˘\��w��C�d�4"�-'��q�c
kVi`L�fp����&�-��N�S�"-�C8K�LC�T��V���q8����6>=�X�����4������R�w���5��/6=����܎5?���眆���c9��Bn����9Z�֜L ���|[��7��@���ʪ	�H�wK ��'�\�����7�2�]�?����v�,�Z?���9��\w�8�P�k����f��v��&T�G�`������u�b�z`��* \�&
X02;�h�x�8(�a��[*����h����G��܏�m��̗�q�4��u�Q��Ҍ�ѽ570��ʅ�mJ�Ō�2�����eK��n<Mcl��~.G�~=�y����cx�M�^�U���j$F��x�s��o�>�]�&,U���i��@f��lG�b�e�n����PVq��P?���5qw��
l����f����XJ� }��2����)�fu��CS9��Ւ<`����a�|=D��r��dW�9����&yJV��s�����j�Ϗ���~��D�ʶ��:_9�o����%�l��b����63��N�����H��#wW9����'"� 
<,��Z6A�c0D��A<��_�cnڳ�KZ��->��Qxrl��+i]������ڷI37�C����a^���ӏ*OfG�36b�����}�J?[��W�����rI�o�ăG��L�F���ɏ�\���F�3aX��z?D�;��о#<`t�0��Ұ���g�*d�:^=��r4��a�]��f�x=T,�!*�V��k{-�rǺ[�	K�|�V��m��["���a
;��c��cl;��zߤ�Z���h�vk�3����]�ƳoA��u��].�Os�D����+)�O��ӝb�|��l+oYH��R���]<��~�gh�T����G���:�o跖�	,'�-D���1��"Pß���c��t��
�-Ev��i*�{p:�FK�``���&�/-6��m�{ܳ�'9Z�+��.(��bx��? R]1 ��oq�ͷ����N?P�SG��W��3�kp��^��c�� �i=�����Ak��^�%Ԁ�e!蠚7nZI����D+�+��j8	k���}�3�Y�d�"��O�ˉ�Ά�����z������Ci����7�߅�7Vu�J��=�ePyO+�v�zK�̓|�K�9�ū!�3�ݰ���)���ƞ����K���':���Y�QS�3G�E���U6�/k�_�Z�Qy�רߓ��̏K�E�������Fi���b���F�A�$���#\r࿱O�����bG0�
�h��g'��,a"^ B_��a=��z��0��۲�<������5R�(�vЎ�y#�TZ�,��G�����<����R�p�;w�|���]���}ُv���������d�����;{�r&sD����C^�Ժ�(���S}��P��52�%�OA����0A�PO�.�09�(;,X�!]{�ƓM��T}D�� �5@����0�ӻ��/��Xo��iT����h9��b}��{�t���O�c|"��Lq��������^�Q����(u�W�&C=�Z�`����G]Ϟ�?HȲ���{�����c�E�����:�:V�|��]��@�5�eX�-�ܥ-;8�8�RN�	6�p�3\+: T줤�\R����t�$��G������+�X7.��w���B��i���?^8�Ǝפ��G����D%�W�3_ӳpB��_�Y0���8إ�i��x�����8���\n��s����iY�����{�H£�U	�ђ��dW-�'2_�5��K���@���5k�]��@���O�����~�q�I$�=��c�|�����-�NkX�H!����S ��r�;�y��RZQ�Ș� TZ��N���ː(@%�<�u��¤��B�[6�x����#��"N]*����0TN%�\��2Q,P%�������廍��<�|�>!�,*rY�h�"h{�A��ٖ�AL�w2�1�[�٭xj��W�z"��(W�Vʢ�h��H�H�s�� ���#�mz5���G�����fD �=�q{j�̽������6��Uq8^�o/Y���I^��-bX��a���:�~�����#�,�Q����(��G���(�|�����]">��A����u@Ά�h�m�ħ��)n���៩�g�|�fp�Ɂ��~��Z/��FsV�H�i�RzY�kZ	v�HvKեn�\U�J�eZ���L��D;~γ���.	����I�4��MU��8�i#K���W�����&�?����t3�8ώ�B�=�1{�ߍϣ��+22��fD�aL`�K��o�
B~/!���9�7wN�h�w�u�{�Y�[��X�/�J���zF7�2��=ۓ2�ђ�z �ó_ϊ���_MS�`�L5��*b�V\z
� ��O�7C�+R�:�M&��J��������^�b� JA� ��rN�e�r��I(�B��[���w��{�V��^d���3;���]D�$�Jw����0#2�R��l/�4���畢�RHN��[�k'�o�V���lV�R"�c5��e'�	9��v\���V�;�:���"2�f���"��ǲ�ؒ�;ٔ~t�P�Nʃr�8�������2,�2R�JR� c�mbP^�=R-�%P�t0�;�Zه�C�AI��U!�rK��9�e�`���˄tL�C�zAC�|S.f��6���O�wy���hO�9�������:�ܹUR[����V��  ����� #��<��������-F�\�QB�7�u�!a_��d�h;}J��^�aG�뛍�i�c?�,�U~�nW5�8��!p=����$���@��-
�h0(л�D�[��Twϰ��So����.㔒\�!���~B�a�E��t��t1@7��O��}{�a�I��E	����4C�;�pe�J���|iU F)&�]j؇P�*Q�3�u�e+5HO������1���;U\���,��)���'��FC��C�U?A*�pNn��TSc����G'��̔I�`Af/O�D�l��������B%��/�`�K��݃.ٶmt�����?7��M����Y �7ݘ/��-�һ�\�ŀ=��s͌�wY��XњDҬ��Y[n$pȱ�J����P)���q	�����rj��D�/b����'s��N���P�g�l����Ăy�J;�7.�jt���/�'����#�"�������l��"ǆ��-S�3:6�Cj�a��SJ܈Sȯ�T��Du�v��Iâ��J\ia���ա�J�D�mW�9�wj�,o�	��z��1zz@�=!�u�M���͑}�k!�N�N,�`	l�n��m2v5��D{׆����U�*0wя�"���1��_��Ei��Y�z�;z=�׌��!�Js��p��%;]8�H_o��2~���l�@d$D��!��c*�R���M>F���/!��R:�m6�p}m%�e�߱��
�g�H�|���%Wf��$�TΌ��+\g�E�(o�e�z���� Y}��#ۧ-_��n�z�9�w�-�Azha�{�(cG�������L�y��lZtd��=�	�i�9Ҙ1V��2�Bg��G�+��c�{���q� mvO�^i�)#��J�)���[�¥ӝ������4�X���-�@�����*\*���#o��&�X0��|L�`M�(�)�2��J�ix���_[`���I/��B�xK�@l`��b�z���~׉��@?�<S��w�W��u	�͇MP���twz^k"�س�=�]�cW�~�B�;e��(S�B�l�]@Q�k�pL�����o�b�_������%-E0z�̈́9�6l���|J�q	�����z�+��D�
����G�l[C�$��)��66���&~��;(8W�&?/�S��7�xcӑ��46-��~y��&:U�i��Q��&b}��i�]����̴�Īn���w��]�NW�c�:ͥRں�[e�{��`��#�k�5�u��郷���K�;�����T��e=�n_J���t�zV}T�u��\j�b�β�}J���\,�*q�v�RN($ϰ��Eh�iLEnH��G�P��u�MO�H+KJ��=gㄡ[>K�a�%�6#�l~�[���}!3s)�0���/V�,Z�v��<9B��㮾�{k'^�"�ӵ�B���E���y�	l$������U�-�F�bs�\�绱R��k����yѼ�������F�@�[��d����ei��ߚ�n6�2���qk� S>�X� �.+.�Wyv��_ZIj��m��z
� �ig/.R�ց̀z&��Pa;�2�n>���et��\Nģkz&�i��&��7 *�c� �ZB�G  ���Ǣ�&I ���_m,c��J܄������i�B�4���H���$���X����I�PK9�})�.09�3r��Y���F�I��B�v���R���Ir�ߺ����/Z�t^4�&(�[l�\.&�O@kE����$l.��{���$��8��eD���(�?r�e���������h�*�N
B���LK������ͼ��j���ͦSKc��<���%��t�^.�q֚��d��]|����(�8"�@�M��Kc�{�޳K�W2�ԏ�mJ�c)F�KEy,'yP_�ܴ��~����N 5M���g?�e�`ᴌ��#������z�֨$&�K�A��L6���{�Ώ��s�(||z���L}� #� �Q�6�3C�G3�<=ݸ2��Ѩ ��6�ˢk+�Q�Q�����P�x�VIz�k��T��U�21�� ���_�8��uGj7ғirk��S�C���ڠ�?<�I;Vqu)i"��������*�Ɍ�W�0�BY �V��� MYxfueh�I���KKMl3���_���(u���E���E�}�T#
#sZT�m�\X��.e�����M271KD��
�^W#��#�BN�d���4���o��A���+��.t	�fB��$�~_�Ķ���q�YS����1��OW@z�9bw��W1%��1gp�Z&2L�} �ΠǺ��>�G�w�a���@�ڕ-�v!��YPX��N5�\��吻6=[��(��܀��i�1�*C����hVd������L�D�}�@m>4K׶N��l�	�?s�.�K6+��}� �!oG�,r�����!��������tb)X���T�H2��hۭ
p
_
�1;�=�C+2�<�t��|D�؀x�r���?Gj,5Xi��"?G@q<��ii���8�B���/3���v��i�/��l��:��:d�.���� �A�T6�
��γ�Q�&�v5�E9��Xs���.(�y(7,��kdZk��>����F�&!�Į��'s����������b�SP=�>Vw�H� \'�Eٙ�Ń�c���9��@`�jb�I���#���Y���O	���>C�b��N\��!��9�hhh�8�v�[�����\8�t�d�y{�l���-�|��}��s���
���F��q�����̯;d��'!y�-&��6G��� )����8�}��>*��*y$���,g��{�q!I֯)z��p<�A�"JS���pnIo�'�T��Yp��ꌏZ�%OLu{�	����λ��������C��Nm��70 �����!l_|���n\>��l�V���f�v�^�Ӟ��K����=WRq��G�3�_������T��_I��<t�-_ 9}��� �y�w��s{N
XV3$[=j6Kb����$VRQHy��SG��_�h�Z�*\��E��S-�DWN�
����ட�r���|��αAOi|NoLy������~�,��M^@.@��~<>\#_��%5�����mh��O쏗CԍP�<�Z������+���<_`'�|�մ����F��7OC�	A�(`{1;�T���� �44�ّ���gU����k��e�1Atߖ�
3�>ORG�?�(�H�0�q��z�([�t��Id' �Z�����8j��H�v�x_��R5� ��$�	;����s`��eWrX���ɦɳ�M"x�)�(H5:�+��8��H�s.�">���q���8L�g��� ��@�Wr�;�S���x�Y�-���8ec{"�Z�
#���'E�ԁԊ��ٖ�K�F�T�����Rh�4_֩H�� �DZo��k��Η_�ͪ��J�.+���<ZԦ��x]���0ҰND/j\d�3���S~T��C�׶)�H�S�*S9#���-�e��&D��G��<q��}ʧ�Z��(�1T�����	�� ��{\��:	�ʭ���ù~��m�:���a`�"� w3c�� �����Ü�q�E�����KbWBD��lm1�̹������@�;��붢5к4�a��-p���6�*aģ�
�6�.:z9���K��l�})I�������qq���X��w��n]^����B� � ��W�ҝx^���緗 ���a�Z)M�Fd���J�5*�u��q��Yo%�I� ��C�t�w":�(���E�o����Ũ��@_�s?��UFo�vsb�E����r�/G&��Z��c�D�!޺ uMǁ�D��+l\�Yւ9VMܝt�D���Z�����{:0Ȭ���p ��\�c��rr v�ʎ�4!c;V͐0��!	s`���׎�q6�S��tY���@uY�-�Sr�6�������k�s��X�[��2�M��2�-?t�x<&�6T��c��h�GL[.��!��F��Q��u���C��T�s>w9�?�#!�+�;�FH;�����M��$P�Iz���V�z��r_�s�HU�,�ѵ/f��	��U̹����H��f5b=��8eT��T"�x�;v]�f�	�p�/׀P�M$F4�A��SE�3�@�21������.�:JS�T:�`����d2S)�|��7��]#�G�3�|���?���d�n�S{L�djp��d�r@5Tn�$�
�C$��qybW��,՛�ό�Q���OL����l�(	ŏ�rR��}/�9�)��!��!��șO�U��R-Ѿ��RG6�a5�$���$`Y� �䂥Yu���!ޒ�j� ,�`�s��hh�"���y�P�����t�4���VٺRYh�C�x83�	���tFW�r���y ���LPK�d���9�0ߨ!sq��HƦ��^B��[�~���ʼ
�4P��k��7�8��<��?���j�{5@h��E�䷅�"�΂K٢��[UB�o��g���ek�o-�H���y/v��y��
�u�	���-4\��\Hjd���n��E�M~��v�X����Y���`hr�⧻�aN��@/E�;.�(]��;�1q1��~�������\	�ȴ�_�wӅך�A�X����N��8j�sj���^t&�u���,r��B��M��6��|ņ���yt;�Ɔu���#��f�Y,-�b�Lo 
�X���S8��=J�UCkam��`�Ѱ�Kp
�ۺ*T�PK���[rY;\����҈�(��e��X��
^��W�Ѭ��-.g��FtU~İGL/�ʖ'R�B,��03���Ԓ����X:}J2��.d��/���}�)d1���M,�F�m�`0�7%��7�����G�c<�sz��9T��܅h0C��5�Ѝ�W���};�Yw���e�0썅?�e��T��v�3YQDr9��$����� ��l�,s�&�WG��F�L��_Tz6�8y�	���΁�(�D�uݛ{Fa !�5xF�?�R:�Ҕ�$Q���C Gq#�>y$��k->���qȠ�����ʛ��R[{qp���q^���)�U��ۆ����ิ��%*b���L�y@_�I4C� !AԈ�+���7�֯���5��ۊ�'�>2e�(C_�Oc�J�7�lY UK z�E���j���c(�w�������Gud�[�U@A{o!�!��V�%���I��lM��f(���w��^E%��C\�@�E�ה+��/o���F���Ҁ��c2�-�#{E<���VT�x[��Pc����X��U�����?:���f$���?lQ��{صcH0l�ƪc(�d����(��1P�?>�@�	�jV"J�r�_�s�~��!}���b��l�tt���AAȠ�\@�8�/Y����3@��"�:<��g�#��"��Y�AKc��������Nd������a@�det�� �3��:�;��Mz������nM]DL�f�
�;Q�H�Fz	>8M�'Ɉq�9�h�l�m|��$�Q�Vo����|��cI+�
QT@����V�9�&��wk{yR���)�N���,��rg'��`��4b[������l���U6�sl4c���ڂ����Jf7Q�T~J�c֧k�k�#^�:��Mޮ�'��y\�J�3�)'�SLb.e�d�oƱ���hT����?MNB��QI�?[�)SAI�&��x���e���Xba$S�S�0|0!�~��7��?VʮG��^U�U9��Zj|��mD�/�����A��E��6��U�҅�)B>=��m��fcl��n-�2Z	����B��U��fQ=�fF��=�1��w�aЧE~ǲm��{�X6�k�Pw-V^�{�Cqq��bu�q$v@V�6�L� \�����F>Z�E88b#C�]�j�]��_�:�ba�b�J	W�� =�Dv?U��Q �D�VLUWO�Χ���;c�F]X����ܰx��'�1���r�8ؼ���"ZG_؉��^">�~]��(��*�ԡ90���f0.Ӫ%Mq�6n+��ü�K[���=0�,ǒ�'��/Ʀ��¸mcwb��7�`�=�3n1�LKe~:gr⑐�3U/��g��|q~8�wb�89�D���k̡����9Q������L8]q��.�a?���N��" V�O��)��0ӄq�B��N3ܛ�u\SE�9��N�L!�ah?w���/��S�&��������>�U$%s=��	7B���������[�E	�&ᲶO��������=G0<���v8_O��jj ��ݠ�{�����჆qe��6�f?R"I�x���O�1t��\��?&DggV�*Að_�S���ˮ�c��N f�!(j���7)�/D"���e�H�f-�4W�E��c3}�K�q3�m.O� �����wc����\�����P�H��&9�}�q�lcE�����UOV$���luq��r�����2��z�\�b����pv��a�O�ȴ�Nx��5��}`+ԋbjS-M�֯U�)����k���������L+r�#F}�����N���IP�n,
��6R�6��=,���x:���x�P���Y��@���݀&+�l?cLP9v"���B@���S[I������N��#V��n	*S�ۉ��;'��uot�,�!��3ie���DX�|�K�`crC���{h���hn�v�3���8�3դ��XogT��6��.Ύ��Ӏ���z�e���j��|�2�� w�m[~{�J�v��m!���2�n(D��z�����xq�\�L�Z�xN��Z�Q_���2���;�5�e���ecUޒ��/+M�����>O�$�2��pL�1 ��z����(L�݄GƏ���q'���oev��GJ�]��B Mh�*ꁯ%5�3@��z92�̫�O��i�,�A��w��;|Z91#�_�:y�n����:�d���%�
��X�p�P��M����qf�u�*����4���y�g-�԰/Y2�>�P���#�#?(�����^Y{,�	,~X�����򳏛@���e�"���3��<o��3�K�o-���.?RI�����S�:�1��J�H��aR�����9{���vV4<�b)چ�0�P߱�j) �s����>P�^�]y�k�� ~6�q�'ƆB��5j+k��f�)��:x㙢y�5-�kC�l�q�	Z�����ֲδo�����+G��o�%t�/�����X6kEcTݵM�;.��/��f����1�����d�9 T����%#����#���AT�G���m0$�8��6�ѣ���wX����b�"���O�!�n7��2&�P�������&]	�N�Mڗ��H���@�B_I��TzM�Px�`8�:��ݭknMK�h��(�1�����"�y��jh;aSv#i�6`c���p��6�;Ǒj���&{~R�˂�5-�+	u�8 o���F�]>5��O@E�$)2%��E�vC�lj��<8��P��:��D���;F���Dl$Pf�K2������E�4p�*s�R�ҍ�i����񩌱 ZP�3t�i����@o#Guy�1QB��Q�$���vת_bCH�)5��{b0���	��a��F�:��*������b�tz��Ǐ��N5�̭v�[@j��6fbu2TKt�eR0�B\ȥ���M�{n��[������+��v�4�S�
����:V�2/R�d�}����1�y��T��$y�m���I��D�8�v"f�P����:t��D�: ���p�}6�HWq7S��m�܄�D�����y��n��m�u�[-������~���L&�� �;pa����#��U@��Cg����L�WC����1���Qt�yuAW˳��A`r��(�������/E���f���A�6D�Om��Lp	y�
^U����ϕ���,��56�S:�K���9�� �y�T�i�`Y����h==��/�#]��KR5���U�Tń��ev�
I�\�`�GN۷����`�~r	���{��q�xGe1'> �0r���>=�g��ۯ�w�[��cz��YӢ�.���FeR���%��@j��7��Kl�E뚻��+�d�,��5�����i�2B�Y����`Tҋ�|t��4z��!�i(u����k��ȹ���m7-�\�%�C��Ũ��1��g�y/��`��w�K����=eI
k�M�֕�<o�x_�^��o��R�W�-L�C�8�_�M0��@hYa'&9�ҷ����nyߪx̧$yh�[5w�5��V�qz��xL?�Sc����A�[�u�wLR�v�%��E[��:=�AT�����G�v2wx&8;�-]�^.��Z�m�Q� 	S)���M��n|ܦn6ȱ�$!V�v	J��t{��1:A�����=��5������ ,���]/!�u��Zt�ʅ2׽�ΧW$�e8]������(}��qᘇ�ש)B������1��c�M��#/��I�q��r�[)ε<@�e�䃡���?����{z��������Uw�S��
�F�J'O�Y'G8�?z�+�s�r�b\"�d�Y�5�P�[n��,�>���xV)1x1
	�UЫsS��y���4Tuc`ȳ��E-U��0aJx���͓%��ǤFy�|P^A،��]���u�)���ND>��f������3]D_�%�=�2;]AC�s^�jh���N=AZ���8�����>�Y7�>F�Mbc�AWۏ2.R[6b: '�H˫�Ϥ�y�	ʯzP|�̐�w���?a��;�/6e�_f�x1ֵ86���ōj��&$����}`�C���ȣ>?q~9Ҥ�b��0E�o\q@X��)"k�|�I6��7�i3
VpÐ�s�Q��3o���8<�#岿��y��8b�o ������;Xsg-�U��|�l��e����2�t��?r�O"�t��'K�'$�i:�空����3�)�#~�x
�y�_�%��(i��j�Sx�f�<1����0.�\	����/��ߜ��lR?2�{$+��P���9��fӒ\��	���	� WH4���c�b'auSQ�|ke��)`��"ˇ�y;�R��:����=��y���-z���#6�p��=��(�7#p�-��L�Y��4��r��f�
��Ke�4 ��ăP�!4ݾ��k(�������t��nLޤ��Ua��T��߅d�GxZ��c=����f�`�!k��[�0�Ԫ�JH�"��	+�m�vN�;}��u�h{Pb�U:l?O��?��ҝ@H���n6!~��g���n�����/�I�p����(�4�'�Ӊ�_ \J��!]��jc���;��)d��@�+�������dً�i=cH�#�>�ܗ��^(z~5�ss�깎D�QX\��Ԝh��BRm �XP��I�;�ٲ�����W���wѹ��3���(1ޘ�Á��� %E�v^'��	�H���F����X�.�cbI��B�D�x�-���A[%�8J?��R��B]2����b��e�����쫒]L�p�iƬc���>}}V+�+R(d��O��JRG��^VJ{tM}/d�|�^��+�r߉�v�Lw���yx7.IaXw`��{�f1X�^�,:�8N�`A�?��.ʽ'�s�d�yKCT�'��Q*
ٴ����H�)Gc���-��͙J�z��JC�Zv�͠��7S�`K
�uK"�t�ﻰ��0,|���X���E��1$_��B��AԄ�=��T&��R!
��]�����9�8��$Ó�(h^��������PK@g/|V��s��B�&��/}R�8>�sy88?�i�t)�Ѹ�%n�\��?���4��V�6��vl0)��(�����}� �.Zn��1����;��ABL?!_��$և����~H�����r�^���dV���e���%A�k9wR��I�{����i���V�9��S=q��H����<J,.O��ː$J�J�E#��К`��$r���N�o���ZbګI݂v�-3Ӣ�;�u�I��X�4� ��M�a�d�������O?�H����c�}��)s���f�5����?#I�^e�P�\ar��l%#3G0(�ц6����Vx����k(��-Q4U�<]dbX�}5xS��Q�AeA�棋º&M�o��+#�ۻ'`���k����wۆrh��b����oQ�L�"��C�e���Hf�P9������`P�ƿ�Z_?�7o��N�����CkH���a�e[?&N��2}t�CKS?_��71C/��T�C,kk3?�%�~i����|� ͰXZ�����n=V�)�'�,�E��ND�'��d�B@�P*��Q�����n[NT��ƐyT�\��̉���>U}A��x,O	 ��6�U��	��j�_���� ��{u�~�+y��<z�<αR�^�Oj� 3?��ߨ���@VD������X�Z�����Ќ-����ߩ�s9s��Y�	$�F�)�~W���5U�\���׿����H���<��K���7ڙ��u�)-��(�<�m����u""��ogk�ߐ��������E�C�a���=��M���rAk���1A9����4��~(Z���?-��˚�$<�{>>����.e���>�ƣ*����q���� ԭ6V4k�syo�8O�[ل�	��Գ�:^s�s|�V*������@_9.n�ץj ��2ʹל�#���?�喉��6kǊ��C g��7��`��?5J�4��� `G�������z�c[�$���ʍ��VRo���9�J�$���8���%B�%���ڭHo�b�!pn4�����V��T�W���4'P�pL�}ۉ���'�d�+x`f9��74 &b�<��%�Z�:0��P�OYi�v��v�`C��)s�t�܀Ǆ��;��9�t3�
R|7I�3-�A�4ˍ��;��Y�8�+��R5�d����ɧ�kQb�W��ԝ�#�/��V���u�I�?�h$���>�'���b ���]��d��rR�߾<R���
��c޶=);��2-��d���'�%��t��+�oz��S�u�L�E����tY���1�V@�9� �RM-i�VKR�3��и~������?yw����D>��	��ς�x^� ?���݀0f�D���+b ���Yu�bY��
5TK���u������2r2q����W�� 8T*./�Dg�o��*��y�\�Ta�}fQI�X#��7ݢ�=�pS�8kg�����A ��W�jq����4:���w�0���,��[H1@�\�<�̃��ċ���a=�F�+F(�/D˺�K��t�Ѹgl�D�)���� �!��\�ɚ/ё �� zS+��8�R����P&�<�Yw�By#�P�5Y�-5[��뀄��1ƺ>��g�q�!��ȯ�C9JWr��L�j�W*;�gu��c�|���Z D\�����������yn�m��*.�v�+��Q�֧��1m����d����2g��.�a�zn�����fj����A��c?8���泪��JAm�3,�`yU�(�Hh��&~e��E��P'�ӱA�`gM� R��� ��i*��u��Q���d���$|�&�����R8��ڡ�f2���#���]�ƌ-����`��F'����!�V�E��s�D�IY����4�'�!���-�w��.�RZ�5L��y��CQ��l���	���K�V��,(�-~�L�Md�@�A�26+D�����}�.jN�
}��㔜QK
$���HP��U�cDm�N�����h�℘e�� u4�,�*���Pˊ��@J�N
���-�eb$$�vk&\�|�L<45� �Z8�'���b%�$��w��"��r�C*��AZ�w�Nl�s�t�P��f�*�B�ܮ��[�Oc{eEG7��x��f���&�+��'e��O��6k��;�js#�a+�y�������J�Ius�oT�rO����ᇆ���3�)]��VG�MF�>�<�� Oc��~�C�PTZ�t,c���~ڠh>�LXI���|5��J��w�| ����ީdu^'�#O�6B��A����Q������h�sK�D��.K�(�)��x�}c��t։����3j$}��d#�'����,[�i*�Ft�#
e��~꼕+d$ף��'
rd��Զ�񷡚	2����\���)�p�v���L��Wt_��+oف1y�: �bpg��߯�t�ܔ�uS[Y \H�EVR�����|�%c	ւ�x�ar��s98݃u��3��	�:i:�0e�p�?t��N�uZ)9$Փb�c���w6���f6fw"�h�6lq�T��٘4#E��������2���`'� 
���;�njg?V��I �*ʙ?���ڌHU�3�$��?#��Ӈ�o��9}��nd(��%D����8���Z��C�ƍ�U������~��N�q��#�g�)�cW
��+���04�>d�{Ԙ}��;�p9�@�`��^C�e��v1��-���DG�+e��r�1{lcsF4dܐ��G�8c(�����>	�OP��
̗��
�I5s�BjZu'�x ��V_' �S�jY$g�w��V�K�U��O(��H
t�m 9��+d�z�)y^�P�c�xGb�����(bS����\Cm�Q�b,O���+�'�G� @)h�LNE�m)��̤�6�]�u�F?�Lܸ�)����bT��H�$�_��7�����n��?9��/P@Ve;�s���
>rޥ�eZA�mn����6��*���0]'`�� O��s�)���"��;>|R���XJ�5���P�]�b<�!�ΝV�����8��Ng5����>OF��c!�V%�^���~��-�u�F9�5�q��_Ԋ����2��2�����Y���9^��'����ga�Y����Pc�n^�N�SX��K�T����
��(����@����i&N�����ȯ��9������M2ܧ���bu#X~�b��I��s�\XL��ݨ��m��S����*�g�P��f�����+!A'_�U-y_���ۿx�o��I`��h���$9����]�p�\��08�A2��Q��72R� {}����^�}.^,��������}�o��T�(�;vW�%]�`ϔ��#y��ӫ
�;�AT�ٻ_����y����
ݔ���Cc!m�t���������3dTmV������LU��W��fۅ�G��&U~`ڐ$Z�9�r`(������� ���^�{�(���Wh� x5�� 5:fzi�ְB��6a�raQ&yx�X�� f��!�-/�`�y`�z��C�`��N���j��z�v߼hQ\��Olf�C��Q��K���V���0B@�gzA�"��o�.H>Yw�A�>>��iB\?�W�Ljc��g�-mJ��!>&^���`@��Y�G
qL_J����5j'}�
V��S��	a3/ꞟj���K�i�7*�#����G!p�hH��2��Ŏ�[HK��Ԝga��Y�����]��6� ?���r� B_E~L]Tg��H�NC�։rc��nAO&%������X��
�dھj����}�Nq:T���Z�:*a-��%,�Z%oHU�H�Ls���n/Р@Y:M{����/?W�M�%e�O�W0}�|����̓��,�E%��B��U��T�)�L�HtU�����v)��":r�����ܻ ���@wPyp�y�k���$����ʒq�� �xi�����~�"/M�
X�'���|�<AL�/�]�0�0�{7{�w��ŉ�O?��.�;�#�g�r�)7	n̐�Iǿ�����$��k���-�2v��n�t+�W-5����Hc�����rg(2 ��f��r��Ľ�F4q���`{S'��[��h=�Rmh6� ������0�
��D00Gܪggh�\��� x��u�I�l/z�@�H�0 ��U�X�4	8���R�H�`o��Ij���F�t�fR,��)���.Ύ��Ʋ��-v�1G3��zA���T�)�w7M�|��X�v��^=E@�.�!H�uyY���ۢ�*�6���}�N� ~V�&�
�H�T�5N�J���{�/[��r��W�_���+uz���'�dȢ"������=��%��D�M�.��@�ON{�ȇm���Q)�<�ߑ!���=�bQ�:��)7� EQ����l�Y���@���r^g'�qd���O+E�y�M����¾8�LP(�h)��uxN�3)�/��ҡ��g_��3#���'V�횷���6�G�mvfG3C�%� Vi C�*i�edڬ6�7�Ǯm�3����KDU������3t���$z#��xO���./Z�Ë(jk��~�����͒{�bO�����^�����h�����Z'��M��L ��(E̗��*��_�_�H΄�+�=��q��[�k���)n�y�Q���<lўE�JO�U2�o
S~���ݤ~�#
w6�;������9X"�m0飻�4f_=~?�3��~3}�,�c��$v��((���'��'��yc��|*�"���]KW�D���/�S?[?kd�?�~#;�^�
-B2��FFҬ�u���Q�j1��ũR#����yV�P���P����	�����h%]J\�Sj��������(��=|�g�ƥ+:nL�S�ø ����fV�z<A�T������A�*B���"�0!���G{hʛ�6�[�|T��#��!��'#��^��u+<.[m��<�����3p.���w��l�^f�����!ɠ��M�W\�v�I����[�%��S�
�7H)� �mM!�AcT�6-���坷K�k=��Lf���˯���
�;��G�>~X���G�$Ց����p^3�*h6��X���c�w��v�pOA���fx8���n$su�ucCl�M^�-��-�J���6�B��[�Jnpg�g