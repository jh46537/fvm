��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�u���Z���N��P���1)v!��/A L���G����i�,�?o�˃����C�]��.��S/o��l	��%6��е�7�4�t�I�A�j�yʪ�bI�#͠��D���)?�Mu8ހT;�]�V�eu�����	;?@|%��'��N�Q�#Ћ��)��L��+��?��N:�|��~��U���uk���v��F8R�� ��>�ɞ��w��!�9�{����,S�:A�(`��D��	��N�Ͻs_�ز �#½���ކƫ�@�.S�܋�����ܵw��K;��C��*j�R���8S����$U�c���az�����J,)����E��������l}M>tHʕ��q��]Ñ�J����٧�%��]C.��F�<�������,���czmi���U����+�~�/sZi\���'��G���q�)|�|���W�2��g�N�*�Bݥ�s�;i2��,l��y`��j-Qs���&EI�D��]��-�-���u|'	 U�����>R��0�z66Gz��|	��{bM-E�=%�EF/=xV��	�ө˸��u��T��0���}��� ��<������� �x,ؙa�����$���.`�ߧU��ګ;�3k��l5��OXY�����I������I�&��e�����u_ߦ4f3abt�A�"۵%/���A����a�H%�]�#��'Y�l>�����OQ��"�[xӔ�7�;*��t4�>yw����S�����JM��2�s<\��E�%����Z;s����(_ӫ���-;��Sn#�9ױ�@��Q�[G`D<џٶ9�-뗙�ݴנ9�6�����O�<�k��÷�OzX��<���_	� ��`��N�z}�wB������9��e
���K��>�G����VO�a-�Hb+����L��5x$1�ʔ\8wǮvs�5�A��s�h)��2��(R�ʺ���p+*K���c������ټ�rW���������#S������)��H��(��!?� ��.I�cB8�'ϱ�8E��c����AYh>ȁ��VE���]���m��2��N�$k�"�!��\�;�+я�C�ts���u�0���d����hх�Kt�ۆ8KxS�ɒ��/��H�f�=�D��K��=���	���!6� >y�1/�y�D"Vc��-ҍ�ʀ��%��խrs
!'�Jl	��\�����4�z$Ws� .����&��F	3^p���S�O��^+$i(��uY{4���W�f�=LF��ܓ�J5����.�E��B�@�=�� �$3p���+��"'`�mBex�;b���j����U�0�F��pfA�G@���^-�/�b��/��R-�"*��W�oBRTf����G��.�㕗#@�;��4�����vM��9�)�H�I�<�V�g��cx�Q�3����c���_��YN���L�'�'��n3!o�j-�����]߇uh´�%`�"��+F3�|�d��L�k5.�""��q��!F߾��9�d��Jl�A�(39���O;&=��l�ms�ǡR�f�A�t�\7��G��܊�I$���.�	�OD��t��U.b{�^��:Y�`���Ҁ�Xm����B"
x�_�Z���gܙg�i�w���������VL�V���ؽ��%�	t� ��F���A��Gj7Naخ��؉Z!h�M��������<�����yP�⏁��v栅����+�vA�م���y�?T9j�����A`�D��dn�铋��H0�ww��']14��!��q�eJ�MD����;���b?��bǓ��R%����+�iJL_�6�A8��6�&T��ĳv ;�\���V����-iy^l؟u�K~qdB�S2j��SA�*U�����ݱ�dn�e"������U�陸���F��>k�2K����J5������^����Y�b�C~D8�^�;�'��K���q;n\�2��<�{��8}�o��.���#�7GƷH,�5�s�'S#vT5�$���!m<���2��+�pZ��E����yKE���N� ��wX%~���-2��9�^�m�R�+g[ǑH�Km�%��<�.1���U"Xuz�m6�*����U��p�G�l������S�����g[d��K��xUZVB���e���J�-�CN(�"�+�6���QLW5@.=&H �y�2�K��E��2��f�j�@$�� �z�U���A*Y {�1���C�7��F�_��� (.@����pQ�\2�����'�K��Y�J+�
�e�	S�*����O��nP����HA�HQ#]���(Vwnn�:�\%t2��v�&��O��/_�1��Ƕ������O�����-�7c;%�:$|�C�t�AC�