��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&$�*�Y��nO5���-���i?���c���q����r��� @�H���%��U�/G�؊�c�郧��D����q8���u����%%֌xK��1� �e�.�D�@��,V{[�Cʕ��e�"P㨟��:E�K�|�[��/j�x��;���X�0��	��sD<�g�C��m�h6����#x�2����Ζ�������~ٮ�	]{��PrF%���&����]X�>��A~���w���d�A�0ø��s�cu�p#��n�1�!��@�It^N��6L���KUkJN��^s�0}�h�L�Ƣ9M �+q�����ќ;5����Z��� A�i������'�[�.5�^��-�֧���6���C��P$�[ը�y��T�k+�zO�������IM'W��Q�.�����E����J�+c2�f�=��ɪR����`���+��Q�gśr�8��~��Ӌ(�O��,O6��6��AӡW����,	-Ԭ���!1�S��8r;�a��^h��9����K��i��3���5A��G�PX��^�D����k{d</���}���W�
��
q��?�u��'3H�OR��'��}i��8�k��T04��}�����ht���CD�
lY�%��:7���̒���\�{�k�q���Ě�vJd��Bc�(�ա���o�[�~��:[3�:���/a`���e�<Bڱ�#�+Q!*�m�D8��S�V���X��힡Q�y���bm��to�W�T� W��@��E�a'\m������Qc=�ېeѣC	��ěR��}�kc�1�M�	��M{�eʬyC=b�F�%��Eۡk��Xvׯ��ve���� �J��cb|A+t��h&�.��4A�`)�y@W��dO;E�;}��R��G�)V��!�VU��b-rF��D���F'��K�8������IԢr������&�>��D1�mS�-E�mW��g4q#�싳Gl��QPD����>�k�3f�3K7�A���[3
�SƋ��<�|Ӵ��?�3ߎ��O��׷s0���X��BJ�)�m�K��fD���<�f�X]\����#��v45GЈW���l�z����?���n�W�����7{�/��`{���&�;;�8�Я�#a@$��?i�Q]��;q�(i�H�&x�G�;�^�+���!cd�Z���`�9�I�&�2ky�~"����6$no�刮`���ֆ���L���^=�����]��%=��+5#4FǹY���L��bt/F�u��������z���ITo��'�Ϫ����Y�E�m�����ȼ������a*7�����ȡ�%�1�N�;�ݶt\$�΃PG5�$�Hv;