��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�@V����B?:S���/���F�U��1��;~Fϲ�9;w�=F���{��7;���UZ �i����C���5!^FZO�B�-��>���V���lrE�^!��ࢆ��Q�k��ԏ�+�I��D�F;i�̃�*��2��T�NL
�P�2��T-/���7�l�'b41��E!�l����N$dN�Э�'o��;Ft0.�(_7R�6���OV���?!��j/M���#3��q�5��]��R�N���0�ぐp$�H͙����:��AS@�
:G�<<�i��rϹ/���Æ# ��4;}��uw�2�fl�K����\�7��7 ����M�N3y�1P���&J���e�z�ƍ�84��P����?�k)���뗧�|ȓN�R��߄� �k���?��6-y���Ȫ���$b.z��fl��)8 ��;'�/jB�FQ�<�`>y�bQy���B����%|����S�F�#�;+��!"��1z�nT���V蠆�/��_1��[p�K�s՚�K��t��eE0��I_w+���G��\.��Y����\��
]+t�m]��:5�|�k�9A}�u�QҬ�� ��Q���}
qA[q��7���2�?���3Jԙ<��B�-�@2f!C�:��f�������g��ǲ��@�f�������� O��d�b�D�m~u���O�]�î
���3-E��e0#.z�C��&=)3���^�c���)eN��[%��B���[/�lJ�Y�l3��K>�����a?�Ak���n��Oو uo��b��aDx���6��_�
��>�X(�������tk�}7B�[�w�Y��+wKN���]YC�3j{\kŀAx��|B��Z�� ]cR�gX�ڕ���4����Sk�`j,�Ǧ����o�E��)�$�0P�4�S��z��s�x�Xm������o%��+h���k��̍�r%qu�O�9kk^����~�	^�Ÿ4�eX�-^�����'�1a.�c\0��#ST��ڑ�9�5��^	Fj�ݲ��lޭn�8[Z=?k�3��J�C��F ��+@4n�7N�i�dC\P��Fdyk�GL�pЃ�ܐ�w����j��G�-r��_t,!I�i@��9�a�(Y]���X��kpr����s3C �>i���b�����SF``�1��9uJ�]=�iKL-�O/+!�W�M��a�?^��%5C'Z�^nSՉ���MA�ם$3�^䷢�^�k�r`� ��BVn�D+.����-H���k6jiH��G*;3� �%q�6U���+$ԝ(�qU��LN|��WP˘��y!J�)��+r![��Bͤ�^����x�<<c�G�C�,7�sz�z�hI��D$�
�"q����<|�ZAK�*����]��ms/��f��ksyG@VӐC�~���
!X��^�Sc���\�>|���X!���D���r1��9&*�}�{@�щ����y+�Y��/z�P���\�@���v��G�E�]�.ɡ�2\�ק�lBu;?Sg�&Y����E�h�K�Ǔ�n5}Ua�9|�Oq�*�\���O+|-��ֲ6�9�}�jZ{=K�#V�Q�Y$����!.j�qQ[
DGj�a����|��x����N�5�R��/[�Kd��,������?�qϰW#l�[������kz�V�E���1�P�"��e�ӫ�L*ˢe3}�Bh�r��-��t��3���R��`���N+d��g�E��WzIJ���wm�+22N`/l����v��yh֨�[{����W�dF�7�J��G����-Whx�ŗ�G<�nh�T}'���Wāڕb ]э���AL�w�!�(K��x�F���
���s���|��+d�N��k�F�p଎��GI7���W���6�Yb;q�!�`����^S?��o�jh{*`�KPk�%�ҫ�L>�PϦ�����:U2��n\��@�@sKQ��+�����L�CҚX;��0��և-�����!��P�p�s�� �-t�񬾬���;� ���\$�`�������˲_k-�QeN�d|gJ�}�9�����
�����O�u�	J�zRK��Oƅ��q��̳�;Z�ۻ�T���Y�Gq���Hʞ��.��B� �g>�L$�z�ro\5�&��b�o��\L���v�J�Ӌ�%��_�{��ߙ}����(�}V�I��M+G�]PRA���q]�8��R��eQa����[��2G�mH��{80�0�bix1 ��sb 3L��(^��(�jDb��!�n���`�a���'��=�E�F����2	�gԫ���=n�v�k��nA2�G�
ېNp׈���9��0�)����"=�.��ﷲ9	�f�_�AR��A�z�2L�kU��/��R>�
<��[��7�D7qD.DU�hi��k��+ B^�й��~��X߼��"jt�����k���e8�m�ko�-Y��&@��\��[��!�pw����n-2H��Q���h�!`�ڦ�� �g.��He�I蜭��\0�f���{ޒ�-�	MUw>�2��ML{r
V��?�%��RTb��E�ŭ���)�?�>�g�E�;4���E���D�Ԃt|s8^�7n����O?��W��I4�j�>k�䢩g�*��[�"r5(�	؅��՛}�w��[���� WΣ�Pf �GĥQ+U�Q�>~p �:/��_&8r��=����jR�<a����lE(S+���8l�SZ5�g�-�B��`Vߗ����w�Ԋ*N����X��)O��$(��)^��48����n	@�E��OFSS�yG��,-{8�H�䘀�Ѳ�[��K�T��r`��[�[i��{����M��1Kk-�~*ԱM�� ���;�˧0�U=ޕD�~�ۢCvVE���o*��D�GjmX,��;{��t��Ժ�w5�����ϣ��W���!��*Fa�D�je�2�xX퓁�Q&�m�8���Ҙѝ@�f���(*��ɖ(ȍ����g��t��S��Qg�(����8e\���&���Tq���^�o��Y�n�lf�CsT�U;� �hltI�9!���]1�X=��$NA�Zc�a��Ѵ���S�F���/�=U���!#�Xr�n��%�ۜ��J�2,�e�����nW$S��j2a��V?&�in��#��_D���
}&Vo;Aa���e�J�Pn.��O6��Qn�9>�k�m����c�: ڽ� w��|D����:������o\8��Y���&�M�h���n�H��R�� �.�g�h�Zk`B��w	^c^u�X�d�\�W|��}X[���-ʥȍ�ev�����@��6-���j�1Q#̬��=��`�T[�/�v�������B��!~Qd�J*l$)�6�{c�9���xo�3�u;��f*_#a6~t��z�E�;z��oh�@�z⎹޽���Rm���q2� ����w}��eI��a(�*|�8rK�ź*����8�"eN�A�3ʽ#{��R��wQ����L�&?!��`�0�]EӦ�������y�p]"��@�������o{�HL���#��-S|���m��}� �(9GuD�,�3�$N-���19R�6�J�N&���D����y�3�1�\��)}�o�3���]��
���� d�V���S<4nG�u��o��oE~&^��NK0`<t�s4���	8�E3{w�ow���i<�'ɛ�f�W��%��7���̧Ÿ�fUS�C����D4�a�7���VN��=���Wc�bW�`C�'�D�kXҰK��Y��C��C�ٟ�`q���'_���o�����VJ�IR���含�3y1����p�5�l O���^���j�R	g�Rv�9��I����i�}�������Tx,A���!���>�O{1�%�#��V����U��aRJF8�^��!�l"`��Q��X��hcs9k>���EKh���xP��J�Մ!ҀDJ�6T0��٩E��ʓ�;-P�T))C��H�١���@6�#��Ȧ�'��4��t59�S+2�?�M@k+1�0b��JX�>o�0���
�`*��1詽?��(�Ֆ�c��z�\e�*�~ZjeaRy��	q��qGԧl�ċ�ǚ�4ĸ!Z)߸ju�kc��ڪ%�V��ú���} ��t��^(�S�(�O��$x�Ȓ@HՆ?�������l����w���.�Vu�#qQ�DQ-vJ�X�j�$?4=��=��}{Qm�+�4�c�E���{�o�1w/hB�����#&&��}DG�PD��)��liH�k���s0s��O��CJ3�e�R�R����Z�x�lϴ�-�*��⊙��v''b��`0��ת9m��ର5�)D�@��=���6�GGDn�����{�
�ա�Tq'��0B:F��V�O����b����=g��܍Yf��fS[2`�3L��6�'�'L7)3-`����m����Pz�R5m� 3ot%;$��� �"�I�?e5��5l� Y`Va���i�$��ٞ ���(C����)#O'�:?�n5��{�om�#	?0k���;����8d�^�{)�1���;���� ��B3���!ȳ��'�]텚�UAܫ�qmX7�Ǳ܂�|_�^<u��Ӻ_]��<"��Z��]�]�ytn3���B&Y8~	���U@XD�����>�P����1 ���Ӈ�f��� �jZ~��R@���k���I�������[Տ��X	��ɫANd�'O�@������]�Y)��3�X|�����P�$V�_h3������R����S80�%'�F`�D�>C��q=�6��g-|�]D`~x�X6u��TR|����6�r���Xku��Q�~Y�jXQ�������Uf�L�R	bw_vJ4�"-஥^��cV��6��ɫhM>��3u�+�'�HBN5g���g�Q�~\S�=��k��7O�IYg���hQ�<	:�H�D�	��۾� ��
!�_���ԍ�`�*$���qꬓo ԟ"���M?�Pb�x��U�M�sFO��(N���F�J�4������i�0��ɝ�[���"�S����UD�@	2�x�z�a!�k����y�hԍ��?��"�ɋ��E�2Q7����V��݊��o�/�-¤�"Y�~��L(�n2�J����[�Ρ��Pg�P�x�Q�0e �/�8c�uFn�S�k���������%��-BÜ3��[���o��t���G��M����V�M�Â'\h}f�Y��vi @2H8������%љcP�A�=��w�aY��]�+�=0�,)��	�"��( ��Ct(��k�&=Z��/S��䞣�"W�NZc��")ߕx-�#�_'a%&���~쑦�+g�Ǯ'.Ha�6� 0�hU�7���	#]��@n<��u�G�1�~�� |���ho�g�3}B3�4sD����Mee�+\VPq��dz��
�݈Ip%3Q��1���	�U<���ą8Taqhg�Sx5�hR����MA���Tޤ��W є�H6%�R�$���G��5>tL�`|��f�6�׶��=�j)r�.�`��*8��?��^D<�