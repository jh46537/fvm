��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,���?�a� ����$���Z�����:�1K�-ۭ:�c���p�1d� X��5{���~��|��U�L@��h�����$E�>���ǓF�0{�<D�0�r�+iqM�ޭvt������_VH@���K�&���q�MFLO`�ꔍY�Ë.���	W�B�vY`��9^����%T|�%��q��q䕕0�E=H����g�6�]m(�`�+�!�p\�I�5��`G��׃��J#�� �q�9E�W^n��#A*ɭ�f����O���_n�����8E�B�@0n	����Wb8���M��k����`W	m��`�2����B���0d�}Z�� �
�����
�u�����թ�t���k�ۗ��z�2��m<�jJ㢝^փ.Oɉv��ܾ����n��J���)B�:d�&��n�D_�ZW]��A<o6�S4�p��@}qjKz�7�<Q|��7^�>����g@�X?w�1 �ܶ3��+b�C�_�?�*Z�o:�����C����ڕ���.����ީp-�w��P�h�͙6�)��/�c?*Y�F���Hō���@�`.��@R}P�=N��F�l~���|��'�FE~􈟀_h5`��j�u(V�5�1�`��S�ar[@y �@�����ͤ�����7_�x�OŇU�0°
�U��f.m|Tlt�#�=�R���e�����-��.��4n��137�(�G��L��ȸ��3�
%�9���rr��ݖ$�1_�Y��ah��F�@Ζ+o�foV�rh�i#�EF�&��		����K��r?+ �*f��`��T��(�C@�}Qb=a���V�V��\c՗�����P��=:p5� }��A����C�0`<�%���}�.�v�1x�iL��I��}��1�Z��:��׋�
N^���V��gR��'R��!a��CQP�Q��WH^lBeV�����/��	�8��x�{�gBu���?��:��� �]�.���ʠ�Vk����~1H�������-���*��"Pv[�K �Q���8^��V�k/7��C�a��إ�>0��6�j�D��1E.&�tG��t2���rhH�嶂��mNE����өx��-�&�lt�N��?Te����r��-We����=Tg�Kh��D'���7c3}[�Q�<z~��'�2�XO�+}p�LJHxm��?�������X����Z0<4��@Lё�n+��)�c������*}�;L�GS��|W<o����gb��`��=q�����<��6zoȘɓ�(�I�~Z����n��o��V'0�L3:��8#��-�!�3M�`��)�N�iș��Vd�*�AŊ5LI�Z��I���?>�;`x*�u{�����	��-"��1ez�XH�ը�e"q����1�9�Qb�):o�u�+ kͷ�w���~�oSk"�l�p�sG�IP�������5��u��>�Z��\hv����VV���B�����;KO�)Q����xJ7>�ҍ�����*�<��9#J�CS�*�&>����s��2���-cs A�9�Z/b`���6"���
 M�5��u�fC/�ZWh3�_
%�� ��y��4ę���v�X�	�b����{=·C���Kt�4�?n糸sܴs)���Ku3t"��)�D⒃������z���i|��ᶥll�Y��;\���ժ�uy��Ü���d��?h����"#k���*s���p��"���R�Aڌ�Wt�z	�3Ix������kH�K_#s8��hB���j��<W�q���Q���L����ʢ(r���
�蛆�U�E��G�cA��N�����e���"�貶���$����4�
�`�����=�3b�s�'2Q(����TN��T����K$�!�9}�^�QH�VE���|$yBC���?����q�܄9�?B���R��<� �v�� Cд��e�g.������O{�(IN�t�Y�C�}7@��S�%�6WE��6���N�[h����:���`�б���k��ڃl K<�A?ejY�!ه�}H��y�,���mT��8.*�,ͤ���v+0
p�~BWpX=ȿ�����}���jJ�NV��M����s��t�?C�$^��f��"��T�(�E8/��F=��5e3����
�mΝڵ��r(	�Y`�k=a�Ɋ$�t���u`�Y7u��������P�>�~44��S��6j���H :�!���l�B�8����	N�r�<!x�M)�������b`G�P�0��O�x0Y�|B7��XK�X�mXq��q�,M80� �\��:�����r_C����a���Y�9�!�C��{��:ӧ����}�)��m~ԃw��F3���Ikd5��J&8=�r�iDݙ�]Ѣ�ѱ9�#���EkMGD�o��/�왥�����r�pu�{��<=Fɔ���q|dSБ��O����?+(�3��a��Ctwd��{��3�<'vk�~դ��V�CaH���*N�tD;�F�a$2�~��`�C�LlM�T }�\gU�؁s�p��x� []Ar�u�{����{���������K��W�=( "�ɟA��į�$��	�:^(WOɁϮI���pNS�ǤN|+=n|���ޯ/^���� �e��w���˂��u!3SI���4�!�檳�Ρ]M�z����