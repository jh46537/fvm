��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-�3�y�$9�踩�t�_�����d���U�!Svg^��}e�dۦka�wA�*Z����;�(�x�ή��4VZ���N��ޯC5��6�ӻ�)�c}�J�;8	��*R�cY�v�m�]k�O���ap;��I�A"cu����f�<� ��Ee����̨�Pɱ*��}�YфF�~���K��'Z|$�K��.�n�Ͷ�0�y<���<�D6��9���o|�Q}���+�U�y�b�9�y�qF����5��Z5�[	J{��Ů	�M�¦�o��&�*��VW��y8�b�w�T=�˒=9q4:�n� ���M990L����AF���0_���Ť��(�Ym9td��0�[s�����u��M<V�	�̯0���W��v7,ey����=.����s�����h�X�>&�RG�tC�T�z��e9�9=��)��wK�*6�9�nɢN��bOͱ�3`	G���k�%��	��o�1�'���J��r�ėZ� q����"e ������f����1��aU�N���+�n�_;|	���C�u��R]˄WB��SvI�].*⯔ �Px�ȫ,�Yj���0�_�e��؜�%Q$��*������������c����hNڂ6���n;	.���+W~.�����f�	�3���ۻ7���D�Z��c�H��ív/�S�<�X���h~��p��x_�"_<z�AAG>[�Id�'�bˮ;�_��+���HE�&�K7��O��q� �<]� �k���AR��`����hG�z6�I%O@����xB���^�z��B�B�vA��H W�}���+єB!�ƴ,6�]�5�MQB���Z�k�R�eU��Uo8�]ɂ�b��T��������G>�!R�A��iǶ����}f����w:{��a�kl��1,���X��E��.'�G,�S�4z%)����b��h���� ��KPJ�{L���ĺ?$T��E��C��&O��>'���sJ��U��Y�8��&����7ù���`�蝻���	'1T�����Z�%e:[xc��K80�BV���=��`+3��2%������_��7D��J�Em�Ø��
���̢���MRv��F /q.���'��q#�]�鎅ΰ��9�ּ�[��H�>��L �0�1F���)�w������$��xJ �̉l�M�;�~��_�=�⡛m��*=g)��1�i%�����?^�#����.ۖ˼.oǣ��Ɣ�5atA߀�س�B�"s_CT����8DD����C��+G�$.Q'���b��b�a�3���%�*+W[r��ʗ��ӎY�j�f�a����7a�eූ�q���sL�ۉ�m����N���C񯨑A�Tt}4���wnxA�Y�s�����XKN���U�X�4���]��[17 ��֜�о�%�}dI�F�N�$��A��B��B��|��暍��<cṋ�j�Nʹ��;0��8I\����uy�א�ɞJA���YGC���c��.g`��(
-�����nzD�ɢV�Dy,�����F����j�^����N�O�G������}����MJu�7�_�P2!�;Z�Q!_����� �� �?}��,Z����&����<)k����o[�,�܌��*�)�|���Vƒ'�O���5O�C�;%��PHO
	{I���L����_>#�(��t���<�Z��B�(�<�37��:��j�Ft�zh3ω�V�A8L,��q�5~G���Л��]�۽(T�n����Ҿ����h�?�H����8Q�g��W���ba��=0�f�ζ���A�4�~�UDcGTb^�݀�	�/Ӟ����Y���;��;�~�E>l�|�ا�jM���3�����n�A*��{���<rP�/�{��0�{�OX�M�wԵ�Y�{�?r\y� �i%�����>Yۗ"��J&ڢx��y['9r�k7�����<^��?�^����8ƄjzQ%�*��"�����ZPg~j#�m}a`i�6E��"��r蚌���O�݅��;\���Q���/���;�&GG/lH�Dd������X+Tj���{���t�fo�lKs��l0E���\==��zdy�!m�S����U�X�{ �Sg ɥٽȨ�m
Y�(hN���Q��m��V�]��u	���>�Ď�7�3L~a4M�#ko�2%6�_&��gC\rd�Z����b\��w��p������F@�� Vi�{�՝#�p\��>AC�L�_@&4I[�kݒ*��DD��N^�^�@8�B%��q�\m(� ��N�ߛ�B5�\|��ӌ��Ub�XZ�Ʊ@��`!P��M!#�(jvI"����ϓ��ե��!���42��\��V�hR���݇?FѪ��d�m(2��DǱ%Ӳ<0���h@�_t���H�X��,ii>��:Ķ�a�z���TK�^��i[Jo�sFY��X=�ԥHy���NA©�G4;^_x����'ai�9�	��uY@{�wvi��<Zo+��CG�F@%��EV��YO�xG�"�~a<�N�/�G�d�� ��g�a��r�h�>����
�Տ &�E���R�@Gx�Ԋ��;�-i���2Ke�B��ݙ �h��sV�*ڔUz��)$>��+�i�Py�׷�Ð�{��$�[�Wg%��R��d��su�W��+��x�� 	�m-�t�I86#fU2��hz.�Ǐ+kڒG���mI�~Q�8�I%�0E*H~U�;Ì10�M�>�C�)���V��v�;�u��6$���ݭ���2�Y��U�˶�K��]P��P�:�>�i�v���Uze,~|� l�k��������+"��Xl����tą�|�� {���CzNj��r$���I�;.�k�}H��ɣ�U���jc���@f����*Kl�%�&��9C��{����wF�T��ڵ�������
VWIj�i_��E��:2\_gL�F���]�&���ϋ���R42+���3�j�cظ����YGdP�"͛��C�z��t�i�)�0�Y� M ����V$��@�²
�Q� �&)���b�Ŷ�*vL>�&&�t��e��b���â=���8|c ��TO����U�����=X��0��07G=bmG�;���|3��%eW}^�h�h15I��_Ҳ� �WRt��_��];D�L>�.^�t�"tP>����j@uaqRv��j7g��^��-jzĩ�q>�������1y���L�li)t`��c����6��B}��������+p���l�����E!Y	��+�I��/���ܔ�a�7jk�q� �M�d���-˾�h�Q���S��%�.�څ���]\����gT0�Z�,����t����n1#�=��XǕ��8[�Vs�P�}�s�&�șv��qs�@��ߡJ}_���.��|�o�XK�f/��П��
HN�]4���ߎӗx��B�*�+���60����2R�
�ҕU�*�'}�`������� ȥmVab�/��Ŗ��O_���h�K^n<U� w��8CdE"
�9d���0�)���o�5!X�jaG�BZt_�v�Qf˃���,�~�VGN|h�Z�"�ހ�8��%���&^{��8��O��:��of�n�c��	�e�b�U��D���a��%S����r]Gka&{�u�\7�����>|��3}���Ɔ���4�Δ3�t�d���1o�I��� ���Nge<7���`M��XD�i�1j��bs�"G��܌DB��7x� ���j8��p0���Q�f��p2��Z�;g��a������z���bb�����ڦ�W>x �
�瘎��j�V��[�z|/Is�WK��l^LUy])�}l����u���S��NA�΁�\�%�0Se��1�dx"
��#wQ�dҠ�"��E�T� �� ����mx�*ρՠ��'�ǌ��qgu~7��:�7�z�*%�&���a^��Z ~�46�\��y�iE��3_��s�f}͢)����)�C/�����P����J-�ev�k�G�;=a��z0���B��^S�\Z���%~�4
��p���?���3�ܝ�J"Fx�9g:ܲ��d9@���w����p�Kk�!}�Bр���$��@��|ĩ3�ݮ@���`�2�va�����lE5�����L�4�H͡3�.ä�iF�(�[�'��>1��:V��G�o]��.�>~��̞<�tOv:8$t����f+��Aڥ�W5IZL���v����g�	�ІNf~����#>�vOV��g_�OMҒ��D��H��*#��7w��GWܲy��8��ᩥㆵ�|�K	w�eu�Cc���\��5���!������T�����e���v�e��#qe� ��i���[��=^*���Z�Fvu]����'�{��	��Z��}3�;rLOj՞=�EQ��Ha9���"��rny�2��:�/diXg5���������ع��0hLW�[��y�^�)t	�'�	���t����X��ޗ͕�Z�3�'���8����>��@3�s�5�G_i��۰�+���&�4��0�K`	W�J[��;Wd�{~?�:�}�7���aw0��"\�q��,�{�ƃ���b�"D���j$���P�f�3*�w�tf
rԔ�Ĥ���_��{F�M�{&��H|�v�Y���4���̐$�1~�ȱ�736�j�����՗o@w�k�~xB��"L>> �ʨq#Rbe����o�� ����a�7���ʿ�Z8oAt���I<B���U���5f�*ɍ�Ф���R�ZL�
d�"T�:���KM
�eMD�GSx8�\�o')�7��
15m�Y��bF�T�,$b�s�u#/!���NHZn�Y�@��A��7��h�숫�W�ci�尫Ȏ=Y��1J�t�o��ol�$�i[J6����Y��u���j=�{!Q*�0K���'5|��*����Y�A�5�gxN���a+ �C4i����?��̓]�N䐶L�)���:�x�o����HK�I2ڪ�֯�>���Ԩ���1�pܓ�'ko�(XX��C�:=��LW�S��[p.5��o�����T��'�T�� hJ7Ɨ�^pSo�f:�ۑj�3b-��E�*����pԆY9��@��M���M�m���^s�;?�6`A�iEl A�3��2�Xc������ڭ�ӽ�^m� �
^ (+�p׆YN���陾۲����L��L߉�7O{	�t������M C����C̆L{l@n���_ 2{S[�T�� G`�G�2��#FkP�;��͆p��&�A�G��RJɯV�BS�59��wޕ���yƊ�TQ��.���ni�n1#x&A���C��>��Y҄v���WKU��5+<P��m?�c<Լu�\���,��Fu���j�~�'��`�Z6>g��7��ۥ&~��|y�?ސ@!�m�䅉&h$&N�V�E�WSp&og�� �[{Q���iL�\D��yKC�Q�j���Y�w���N�?J�I��~䙲Ƭ�G#� y!Ps�X�,ΞJ5�t����L�h__
XՂ�O��1�0�𙹔������ ��$9��u'�Ԑ��.���n�9����Rx��Duw-W	0�F	(c�W��B�rNS��y��ea�C��"���d��돛�6�Ph~;Ǿ���
�d�H��C�F+��5�Z�WxQk��8��W:_
=�P������o[+�����*RQ���
k�Q++��?K���Q��ܵ7?�->�V����#�#�ӜY�M�5��vJ��i��#�bY�]P��X����L�S��^K�����pf��y �5kO���'Mձ�bO�8�".�^���J-Q���j��£�+sO�(=6 A�J˸O�eʦ�?�w�m\j+������ b��:��a�و\SԦ ��M~��\;��&@?�x��J��z���Xb��\���*�Vƪ:�m��"�/��6��*R{���0�Z:|*Au*&cwXB���T-u�G�h-�d��^y�j�"q��K���?�LG��Qch��Hs)�i`�����=dLl�Qv��7b�i����N	;=](��uq�lK�:G>��X�7�]�v���f��t�C߂������8+�z�����ނ�����|��@w�+���c�� ��"�DJ��������!i���3T"]=��f$�{(�n����t|�y��S0HB���7£�+�$"��|�?TH��,� λr%��W�rˍ;FY&��k�C*0[�^�o��^�$˰R�o�����q������rpa�XgT���e�\Bhˣ��nN�y���|�m�����͔t쇁	%g��)xq�m��8�=/i9T�`��!,��z�*,��H0����3��n��ˬ'Qx���t{A�c0����ɻ A�e {z�(��id�l�� ������e�V0�+�r����UI)$�eK�p��ق~�9���!��k.�,���������z8k�}�=�e] ۟�罳A�Ky����H;���rX�A���ax�Q<����8�nY���
���K�����+$X�/��x�շ8�5/]G�=�"��Z�ۣN��!��pS�#��v!�Wñz���.�t��]9-l�7HZŜ{��h5���ם
}5��I�M?$ Xo����D1�
o��vS�}�����pp*��p�8]\���Y��'��p���]��g�͇V���A!^���9��Ď �U�0{'�����V��H�r���,�3��|�lM��K�U,�k���0A����V׹~	>���C�.J��Z�1�HS�!�A���yZ|\z۩��,(�J\�0����i�O�ML �>�P�e
~����3����f��\^��6�����D�KUVq�>���i$�qg�~;���咋��J#Ex���'2q�`����h��m >�Xo��%�o��>WO}�"�4��>PT�����h��I��ʿ�X�e~��9L����)B�h��'���]��+����)��?�	7@��h�V��5/���8��W�5�Y��������s�]/''��	��b�<�D�5!���m>�lk�2 ��[5�^a���ff�s>����9��Ce��}� !_��C	�$�)����>* c���8n˾Տ��1��`�\�-_TԟP}�BL�����Q�)1l�L��*y�0gަ�5qp����ĸ�ȳ�Q�1�Yĕ�&%��Y�i���n3_ҧ{�VeE�_|<��M�h�\S���K߰���k=_�m+���g������B�2�Oz/{���-V���	K��M?�,�:�!�e��n���I&M`��4���J/٦]N�=0�mKF׉`Cb �j�e��"��T�� Ǹ9��4�̀l�pL�Иf*���w�vϞ0�J�-f��7�վ>��?8z�dq)@U�� bZ�ƭl]T�Q��K �}�����1Гw�+�[`�T��8�k/g���-��s���wAb�܈�=�E�6aض8�Փ?�yv�M��"Uoy�_D�8�k�z�^�5�2Fj�Oͥ�9�n���$��/ǎM2�V�c�d�Io�̴B���D����J;�@w�.��>!.�|���iwK7��	��s�1W  ��)�X���V̰̓}i�3�T�Ԛ�X۴�
�����GL&j���``)\�%�_Ҕ?V�P�&��x3��L%^՚�NB#`� q����I��}굙�:��P����;`Y�)+ybSJ�֌�r�BHT��L�3W#�x�S�c�s�o��ҀU�w���5WfCY�s��UR�D�կ8b\ �y���\��?�݌��s��ſ����H����3�bp�F�%��ZI}>��J#��P��-�J��[���H�E��ɪ�G�lp���h	Mn�S��f���������h�3�,�hV�g0;��:�GR0�J�54ȺkcА`���V��I�"��+k���?��n;��V*{D>ؙ�5�
�<U���b�@�	��h�e�p�;�cLѴ�;(� ��[u�\ԧA������6�ұj/g���*H|[R��i���B�_p�.��m�έ��M�T�V~�v�Gx=HSF���]�1��B��Z� �ӓ��5h�{�4��R~�/a���B�|5���5"/�0��Ȳ�:TX[#���!�^9Ο���PF�lI����YD����ı���b��٨��������{)�nM�b!�T���H:&`cr��&����T���]ܯ����tlO�+�8�"@��׶�_�n31���;}�,����Z���[�S��-�3ɹ/�(����]��RKD�b�ܙR��j��vc<���U��ļ��w��3�El��_T�2*�����^�����v�,WvG$[S/j3����s�l�����px95�ǯ)��:��L�{yf'a	�-���l��.�(�O�VK���,G4��`����_��Od4�؍�&N7Eb��u+���.Kݨ��v~�&���6�@k��o�񴙉'6�y����n�s���饵���v�M���j��m������A�P�2�_IS�l�3cs~�;[�S��$�S�bޥ K�{����$�#&8rk�:MZ������N�B	�A��@��o���;�9o�����,��0�s��_2^G`����(xڕ�t�"5�