// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:19 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JT85Nls5WYb5wQEqdbMWY33/Y81mFmFXm+dc1pSD06Ys96JJ7kkPQRx7GrRFtQI2
7u7YaRebzMDJYAWNAx4mdHJtWiAi40XY4C6tXnXfpZp896HNkTTaQTs5900dt4Xt
zqT1ZuT+vcU863GGW07r48cuab7nOvD3zzvGPDXRDsU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11104)
RCrEonas6XvO1xvc/+KxcH99b+c8ZGn+r2gxctLCK9FfbapMQnjqML+lHFfNAD+D
z6uRbWq9ZCvHXkUar7LyjIrme3zNmK0giY76USMWO64VJVas9YqDZlGZIMyEzBRd
cW3YUP8VO2vDgSRPYRQvyTaTo2cMid6q3K84NaSBqsSChBkSRJV+ZnKBv2Dz1StL
mZ1aov6pGX2WO6pWOKSGaBskbJJ46yBtISJg2dQkPFQHtbT7SuQholHTRb5abypw
FcWnMngZMW9WcJeqiMn222fdlLFkfQ+Wwy8uA+jimt6cdonkH12AGL+KbjSP0P7R
9RiuJQnupginVvS7uJMRe0wskch2zacPbELIsJHb03pYjGQHZQ5BT1pO73uhZ7L2
cBcjTYTx7cgAWY1KVyI1WQDFGXHQjnbcU4k67nswK/IUjodbMK/29yeeIAUpn3lg
nmjqP6MCYP9ynHkEKMKgfIamQGEMZpeeFpHphbseWBCHB0fL0raIwMgzaWuA3WMc
1sIsutRVGzIGhBw60hcIiuxdXHvo8OzoRnz8LaKMHk9WSTVA2FA7+Uqsbn++Zmre
jIyn6FiU+dJIvPcZgpH1p2F+l1/Uqy7M9xpt8PzoMkULpfVUpu5PoDwkLxhmeQus
/o4jAwVtBoSqh9Z2UXIkto8Y5MJ6a5VTJFHgozlsWDpIHZAmZhZgvq1DvWjvA9vz
i18a8R6ydTYFpLc1/FXhh3JWR6FjYenYX9VPcBWw70RpbG67a2q04smKe7Cq83O3
NKoJ4QiLpdLB4MXmFiofMgyMJJVuj7yu2McLEicTRmpAjHmrD5VJMjJM69J5zZ26
cTA6eNZuckkdehgh+AOuxGnH1AQWxC4l8DlLkjxlDalwk3EMGY0Jsn64jmjAqzNG
wZPCsdCNsQNEb82yqbxsAVm3y6CZMPjmp8WpOK2I15I93ByLB9wngTEBhBZ+2h4+
Jvhm/Mmf74et7J8eXOgyK7wB3keRelESi++Ky//qaee3C3b5PpCJCR07HZOvGY4U
MVtrLf9JNXzUrXV934mxfILhOagrE7Jfw4Kqr+nLOxwcuiuqVNxWKzZUzaSALDnk
0tirTqGWBhj+csH67fmV5QUKRUJRge7DbesuIXYYmYDseoJZv3iKB+HnC8ubq6UF
Qn2xEG7NGoyjDZjfw5/r4tq7c27ISrb6JOGPabAnGc078CbkdUqhB8Y8lFADA8ea
OV6o1i3+dNHYhfWj1BsLXrQGov5oIZQXo+n1RqPEEu2atJf+9qHAnS6jAVISffy+
bWxV/Q8KYoAG6Q8x0ZlbufPpcXPWVqX7/wAyL5M/7JmjD4cPjvLUykyVVDZ0pIZp
s9ZxZFQFRLgEgEROAI8IIdxqU1r9WfHS8HZZbivgsmpWj/EYnG7VPhfvOxX1ML3D
+39GzYGsMKcMJ2eUR6qFjFVH3TxVibHuHaLg8hfDBiJJIqbXSnvymppL5UGmF5NE
GG+6rvI5MjqcVfHHTrQhcb25tlcl+HHet16I0uqERxO14R8tB5HqIaO8Fq48DrtE
rMBhK/qkz/LM+r25gVOOVB3d8okurHWdtpmGW6d5hA9Rq/VC01dIvrOtl0zkIiQv
sXmw2x7TA+IWOgn9EZMhazgiM2m8m9SPgedYGJp24Vz7NaD4769LDWKD5HBck6Aj
bbcpNL2tlHYKRJUnXM9G9zAxVUd2wBK1ZNYm2BuaQYlDc+gDoWjCkpsCpu9AosNk
Ff6AolfXt0W1subVrExtiPVlaIUWGQXgCEfHS9MaPb5sMk2DILa1c2C6B6azLNiA
uwPcHapc3o0HM05zcoXvNuzK5mkrivnRdftNArFgoGrZ+UC5TODDdaeu87nq7S6q
Qi0jrmYtiaCzTiQyZzNx+grmbNGYm91srU0mF1UwGeF6vdEKlfiSWLoZvE5mNnsF
cC2zee/lOU2HSZauB6J1bB2gpQ/08oNnNU8etS9LarQ03FtFL71WRhYxZ/EO6M9E
vvxuXduIq1pUqg4RrbHEje9FLyOfEYZV8HGXhYg5S31IokgE7A4Mn7f4mEAp9fk+
CsPlRePrXj+1pbubJUx50CAABdK8lRmSFZfUnlT2ryrsfzyO8fgM3C/5XgSGdaHb
wpnsDBYMjbS49vB71oprFd7Oz4HIPv2/fkc1uDKJLBnBXqbvoHL0dhcVV7fstNxu
yKOE+/VGdTmnNcWAOIXzGUdfyIz+y3sR9jeB1ENTlh64BUX0bIaV/aM8bOEMDIzH
0rbq+VvrSys93ogIoITzsifvPW1KHDPJj+Yu59cBPYgKM7xddmugszeLgZjNvSC8
SPFknJsokrk2EI5KRnJkXjSWAgCRqie6SY/0dt5+JVP1l2fT5M20tmsynZE0ueN6
coIOZySgTf2F6HjdBsXTPnETDBfvZsRUyRrLkFbbENZx9jaXkUqG8w2dJGeNtMdE
iDjh/3hWgjKRd1G2tSoEfQEGOV/+K2xaWT2J6zB1c3V7XINLFnU0ZqDxxfjAg70q
R4XeyFKJbpQdgXdDRtE0sEuQuCo4h2kylzOyjlvjjOs7gn43KI0O0IsRaYNt7Qf6
qazK/hluCrTk5B54LRzhqp+SoqjeS/84aAEWydZ/Ppct1jS3Y3e5vR/7DqSOWNos
D5maxHJfU3rzK+iwD/Ltvzz6dl1xQIcUUbfVtXcvAECTVAQVfBr2TBdVgBI5Tmil
6Y2YNRyqKuGErxr1WPzZ5tIymvR5S1bT70axW3UwZD10feZWjCwQKaXt+gxkBO1B
6tMKfXvxcnNW4lu0SD67a6x+vZsN2CUG43lnHro7cOK0HuXfpfQ4TumH7YVknrRd
Ca8afCI00DQ+rOfYzTtP7SgISwYY+JpekX1Wa1+HEMe5Qdqgr9Wlxgdl5k045Qvz
DKyD4VjoHPHa5A0PBGV2CZzy8zfgwxiZWTt3sxpB3sGWhmPZmctUtaw0ARw5FUW4
o1o6LSavZdQzV04HLWROT9FGvqeAhyfnCMuInZwY3t4XE0VMB0GscJW9sOtXNUxv
O4Ipul6AVZT83SJXWOYdwzCsb0OR8XKi4uvHelTGz9rFOzJ0kZGPKPJrBslJQNCW
VJplA1oJFoXUDiIxeVTXe8Nz4gxJXL3s74zV5wnU35ZcMAtWKAN1ToAnviOAdqVV
8+822G1fpT1Xdbml7R5VCusyi8PJLEbOSzK4hxJu8VmFMzi+X8ULXBIbKeioZDng
NcSMElLYpLhYHcpXrRnhVGWtHW6dy/JjEfF/Dnp5moa1tldNRv+DvDE1asHMLK8f
WXAPmxGn+kC1e6YmM/sEctxedU3n9xjPtDxX/k7hxLp7WZ4ZK+b5lW+I2ytuAr64
Vn1yfSfxgdQB44M+QSma95v+jIuqy4jsfMPGwZu9BUaSoyWUoSwjdQ25B2VCZ3rw
sB+G5ATBACM8RSuTo0DNhlwy9vn1SuMzfnpPSMpT3UBNXjx5DNud1AizMxgeqrVJ
itsBXmrSduAD3zzLxxolQhGT5ohx2o8VMdXe3VB3KHsFssf1hsg9dtQbb66yRkpT
PFEwfgIRh/529CI0eOfvYhziqxCI7TOTW5iOci5qj2zk0+5MX6ippxV9f6bEJVS6
7OsVPT2YD+0Odj+i6sjfdeZrafmTQRPHJz247OiGZe3/yEzZ9joUmemGQ2iy0Grt
niEpIgKWyWbmj7wHrtUrvkS0Whal9pK2NDmIt89mLx6igU+O5ELYj4jVnQXUHPJC
JwxkiXAOR3ZJzsKJub2Kon1vhkE0HXE4iShGwbWps9oKryegclIvbCo32xHi2aJp
KrEtzXhqxCVexG901V83HkK/W0N3yAJCLZ9toK3Edcft8NrVFoxOa+4YJOUtUiKe
7ALSqOb2WN37bpYdBPRFKhjsRV0alhSewPhbFmVfVo9GKJCFK54J7GYG/lPGGFy0
UuSqUgjZTMZ3XrkPQ8ebiBEUE531vi2wiN5oqX9ItffbQRYqhQssoG+DvobEB5PW
B2WisKL1dKFMkswIfYPWlGtu8dSdn4YFq51bOdHs3G1fgDQL81UbfvCJYGwmfAQM
2CqPyEQnlSLpFyAvHV0RgWR8fl9EGiLah0lQst20JQnaUyNFI+c9EZy1FTaBO2ie
3+/BV1XtXGz7o2BNCmLWG5rxNk17svatgYehHu86m1bFpY69sk4x4Ezf/3e9OR8l
D3K/8hjSAfjJttBbRLekPSKDPHoIbNeo9aL+acbUTJVVKI77AdMUHaZ/skc1ihfv
BK2Q8eD4mstRHQqM8GNb/x8mQMkIMMmjfx3jY9SwSdAPJ6+9dTHzF+kTURicIxny
ca9YBzwyJmaaryhTPw8nDvFmVPa5A3Fh9PKcFogLE+CZAmoDLW64Cw0FvNkTTB21
VO4j/59P4gLkOsKfjl2jiaNjdVSANhXTNc+krzd3FIaQUgujkEzlelvaiQDYr3ZV
4x5ib/o1uS45+WZmJigDtnkz51xHvpyjmvsMPdVXqaHmtTi+3zcUaBfxTJ9rMutx
9jvAkKi7r1FOLTiWLKJaqoVDbHogMg0zQx4EU7FdzImu9X2NPxV3fzXMAIeDUamN
/1qO5KylLfN4cVW6zGoKlDQXkYlYDiOzFAenNRbS97tdJTtT3+FNI9FwbkGqCUxK
i+JGXcMuSssl+4Qkz390THrO2mHwyYo/OZEfHSn9segAc5aF3jIZx3JzV21SCoUf
8x369ZMt9o1WWO8oeUE/cTK+HuTufqUXyrLSINwXXYREZFfsVWkoxtjQyDTcobmU
vj3Iy/oMm2jb+qUO4sKTeYeAQQxoiaBw5eR5CPaTe0LWVvmBWxaLUBZM2Wh+yKYS
Lii10YiinT8ef/VdZZ4x1Ch00jwkyEv7jGCd8CNQFQ/DTB1pas0SvbE72jvtHRgX
ZFTzEYRZwjnGRDU1wEXQ3LQBZfYxoxbZPnw943giGg51bBJ17KWtPWFuXZbhf7Mw
i1K4WP1NdUSijxFCxaJtMFIJ7ttZHiMUsQaRK24oyOfl7nVbW2LKXA3iG/leOqhg
V15knUN7DIC7O2XJJ1ADvp90p45HioEXTNzd6cX1lT8apjm/L5whuRebh95fMBRk
owvywMGnft9jZ7aMcWfnXIoXjjnyDHAfTSLt2X47N434/MiQgdgJURssqwW/UtgV
A6V/J84mr3KZDR5Q0CXyweEFGY78N5iN0JSkBqECKjgMo8xTORUi75Y8H8cWvZcO
AhLMF3+coyvGYRFWvr3aIvCE/cPd/Rdd3zrq8GrBJGBKhYGxA+qkKcxiH/7zhJRm
8MCQHOkX25w4MxXT+2NgrHfelLdhfRvx6lYCE5d+qmSWL44xJx+2t9prq77oiID+
Izx8a+Aw9sVGZugPNYeqhrdeuQwlqT9TWSyuHUhENK57MjWbr7xk3rW9SlI1Mgvo
XlMAoPfh0tnvToFcTd2ZSzRRNI+I0CQqJJCetu+CckSX3Giv4oPz8B9utC+4IX80
qbP/ET6OwI46F2GFBPTe4GQmSRDuLyFkP8VkDVnmBL6yIBFcO8HFkQ8Hm7arCnYQ
U9vOavRjjmnnTMEvFh4L3ijCEs/U/mqy3XadOOThDpawItIufWau0n/FStqNZcwO
Fqgv9tb25ud144dxITTXGxiwau/Gq2bQwvqsMRTAv70cqDSPtWILz2pTBPsUqZAf
D0yR68SY5o56WoIqy/uoHNblJV+/oO/DR4T+LAoeWrIQJ2H594OW/UQwSRU2UrwB
psXS/HBZZ78lukfGVVH0pnVOu7T+ZG+/6ZmGUNzYzcdMSh8Gg//ODdmZJQenmGbx
s6RdFBIBoH8n/JOTfw7QkGXklWD6b5zHgrFtcPnRzRTrifqlO66Z+WvOYX0XVMoo
5Chvbqa4fm9NoRAxLsG/zfsbX7BPxZvnMfVTgCVU1ChKpOtrR+KNQOJFnAFUbokL
kifMjKYG4oZqmLbUh25xvLmzqZscdS7bi7FMlscVFLKkkXIkKRAwE4vUurf07rr2
Jk7syA8s4WLP66p8HImZuG5wLqK2mCKFJMyD9k2VvFwsrPytFkua2+xjSa1P/gac
6uj7aA0aYWLy0rPBHyYGrXC1nSlT0nm4EjRTved16V6cZqx4ZY5CRwPUajdwfEiO
jewm0OmdBSC2WLtrwitr8mL3uWq8OH41SDv9/LM3X3c5q1qUn6RaU95wHeWkQqQB
AtnQOFC33xG5Cl6C+GGQtQV3Sb4ufbYVJ3pAHMDuJ9Pe55CBxcZcE2s7tmAr1iIW
m6cFuE+tjPwcLc7l+hHk7TjDm2HvDIGFUoqaBEl9BULbgIhGTLdJO5ypGqBYn02z
Gq2n0dRo+c8wZbu4A95BZayEtf+rT9zUZOZlpaw4JOeX5vEdTtA4o0rh30Mplzq6
IYVWodmcMQUwpgpTcRI8xsmZX6q5Hgib0JHTgyMtBIDWO47nZhCyU+N+XtNB8ud2
oLz/4ow+vlWwyQ8FAR/nElU9b3D//EJrhYJCijisEON6xot0se+CIfXy86Fs9E2F
tjgBHLEJSD6OStzVT49Qsjk28fnXW+IYWN/bXa7FBJFo3DGKETtZeVuwwqVnwc4Y
2dYMx8ckfBrjm9soSNjyn2xOk+qluuEKZsbpTQACKTyYnYwCJ8/wvwQowl6UH+8z
VFxmeKxbBNs4zBAXXNoY+SWWVGHV4eE5oB1mNQNoQYnMUFaJ2sxCz+vXtN0sNEhP
0Ue5kCj8yMeAPGRfRBTuJtd8jJvSOzzWuoCCHdMeRATP0XnloV1rU8f+SaEPOsIC
spaMd3Tf/DKVTS3BJKBCjqYMe8Cyb3nBsvfS2oPnLYrGtE2Cv9i2RD4oBgmiHQZK
ZjUtjZGIrbNlyV12Nd+Xn9qRCoZ+8XhyuhU2gjqHS/DXtuB6HP/wNHDU26Oe1imw
lFOO+CA6oI9kA86Soj+w+nuQ9KYHiwSlgYuHe3FzEExYY7Ro4gT0F6QTVZadcMtv
D/BVWnYyjYKrJiH2JSYCvhgf0l+cuwnWJcAGVH4QpaTMI/1lUEex5UGzrH7o49Cp
qA2sLhmDQQZQkP7ZZToO7PzG7L4ntfibHg+pYCzgiKzQrVQJTEfs/Q3YObrQeXok
WAJQ7uHteO56H3/2MEO1ROHDQyz7wNfGrE5NxbJf56N143Hj59Jaw/8sZlrt+B0r
S2HqCnXHWyjgEOm6pftMRwW2Qe4HktCS+ZcrhfCskmz7DD4ptBtX1O03jXlypC+Y
8ydQ/pHgU9B4KaA0vLemfK2efBHT1gBWUhnEKd9YkAOXowc6FpXg29QoM/khwaeR
EWxR+bvgdfrYyvxBQE79y75TKtyKKrx3ysjCNixqqGbnV2enA4Y6eLKqavanPPeb
qISEMcyuhjB82ncysAIN4gEEop14jn49NrAs+9J3ihPfhXsVV/zt9Bj6+S2cG2wj
i1aV2KvMjZdWbY6clf143OGIOMz/myN4F7rYUJEmG9997Zp1TLn74pG11x1/D/5h
RuD3yMO8eu8IkGvvohalif6XZeWON5+xK4zIIxrxD586LSDTGSBMZZ9DnllVUj1d
VqDxsrsRcrkm9WqtIFwK/SgvsA5Rn39vriasDBH/gA1niATV1VzG3Oi2bnIouugV
sS7Y9HWPOE+VyOgZIhZfyHpsdGfykYBaONyUHi+Iu3KlytLN2JshKvudB5CBubPl
ehs3/Pvzx7NmluopvO20eS5TEVHwWVqvmETZG98ksEtCqZo2n9HDQM8wTVIVtIls
A/CkPiKd3Y/Y9I5LdQ1lTZeC4nZauT4V4FvDbeRxq7udrIHrPuhvUTifKkgh2qrI
G5W+/WwyOglzmVLJkNpfwdcdlMZRNDweziWFscNdUYWG/AGQSeFEFBgSj6xLL9Cx
lfpVp8oMlxaOZKQWSX6xRWF45tBouF/UXBcqjGRU5vm0RwssFDtbPXsOUTSgfrTB
jx3sgH0FOFcKQZcNpjoKb3nyoPi9uWjo4eHzUSn3rJeUWlRiT3aQg3V+oHB5S1xg
QhV5eNVeDfbK96ENTVQavvn8bcMZWhRZwkhxSyRa8Z4zVX6LNg4XSBURdQsfKEQ0
iUcC2OCGsP6FxyzJLc06U64oe1VXtFWBiNdPoCMms3WK4TV0fWdtRfDVjdoQ8dfb
+NKtQUygfLgt0gjDRIKVSQ2vbFfh56tkS0tTy+oTs7LuA8oV/UXHb++NbxIsFMZP
SAp7NuWBRc15pN2BkHB1XhZ9YQY2NkxPCOdjk0c7kaFg2DbdvJGLct9ZUjGRjb3U
SL/zPtLHyJUDJV4ASuyG6Y5GwioJy/vBnlzIk9LO/AK4zvgZYPyEQ9391aech6WX
52k/CYPlX4/0JbJvJ5Pv2wsrOOuwxCiZDRmpE5ZyzBwE3Ohr7Q4Bp0No/dYdGMi3
7G410tgxn8Z40j/5HJr2PJig+pJBjMJ9F4SOJhyVHfo/fs2pTYBQXq9y6ljv/8u3
iY56sblJmIFs31KRyb3IMb3X9uGThhKfzWzxNoSMJMX9SEmM9ds2vV0LWSQ0brNV
T6nIvhaNDfOlFp4hCiV6yrpjBE4JREA3X6mFgNPamdj7iuaE9QzAh+JMhS0Ctvdd
va7soFNEUtVPHZfQUnksnCtYQWMm3KU7NjP/nxq/oRyp/WFuUiJlBOljux0SnRQs
N32ZgL/rb8Q3RGSvGuN19IZfx9p+KHYdZdYMqzH5ovEe5D2lGtSbAco59ZUa3Hcn
Z8HOg5Qc+6qrMEl+hCPe7kZEOmX4R22ZkPxmW9OWpNUDSQIaqlV1+1wI9TCPRgh1
y+EWLJkicuoXIC7gsH6rCvEfJdUjrmeImzgHSiY+1hOaDmt/GbRIQgg887jcGWW4
tfaXqRJGaaXjB+CJaYMwz7wXTx80gMTcGHqpRqohljq233VkkDnu9tqq9Hul2HFD
NCm3t3LHLG2yprrt8tp6in907sQXokXMI+fJl7gN8srl8VdQHomuQSrjJxd7ZUJC
9U7tR/eoOISouQeRwqCCSkLjPHslMftSDOUOiemtXiHR8bDoAk60NE5QgTPqBCQA
v5KwgLbs60xvikX5OpgRt/I4szll/ubmaS6RJSA/aPb2EQsyAoZsTOuKI0LJ0V4s
TAy7/WNzIvR3Po8j6hdHjD/ox6XbMpRcAa+IoSOBwxImjCaoOWCWQOEe8xdh8Lzk
YY3koXd4aYhzzzXlB10ap3ShgQOuzapX4Cw6Bm3GO4eu8oHNWrWf9bTK+Cgldfir
UA+9akKud4Ua12rrAErTnt6UCp8b8Gn4bdr+qxNEpVay1U3hNFhTwCF03+rA5QDq
r93mnWqXEKxGDFZz7tlMc91mh2i6gbuoOuHrvBsK7bT2nB+gEIjMIfK1/HntuChY
oUr1QUZUD1322pGE+5FocG3KhBNyhz5dJLxCznARuVjHA8RbojBp3U2P1meLeU1u
ty3YZJK3INM26Z0heed2diKcFd8T18TmZA2CGQ62feGk7mgQwKGmeRMEhzHhTTvI
92JZOt/Hjjj7qkbNeu7fk5kZnV/OYlYvQ/Jf4deSaOPTCUjz1vP5bA/8lhoNYHOR
CuKsn/tsUG3tXWjs8j4Xj42z6wJ0cQFVu5Mj1XDcDg8i8s9i5Cz/aHkdUsjLaGyK
ncplAc4G7T6Lk/ttb8MuWr6eo30iSJmwTJLz25/D2ZwjYp3Fjj5kziqrAbZBi3sa
9mDivWOgyCRDgLpeSDFLiK/W86Dpy9VJyqxjXTVX7j+Sy9ImNZSsNdQgmptZ6zse
+Gop1iSSm4gsN8D8qO+4T/FxFnBthcxxSABawRWe9+85SzgVsDMaD5yHm+M6gFpl
9kJt3iMMCKN9HWAuDmSXFZXBsXnkXeOv2Yvky4Z/k66M7dZkSeSm6sS2xbz9TCPg
YUzTfwvM8fC3mp6zBMDsKkIYV1oSdaMyt7MFOlNdEUSBAbgH0hplDmwzaUc2BCZM
dUNCxXFxd91z2Agxt4p+7zp4rWXyMoaJxg7qm47+cVgMTctAQHYwWBaSrJ33oGCn
hGoY/vVCzE2Go5DAkQsaVkxXE6FFaqtEHlFsberkdQnWP5ziPBvYgVESsjXNfO02
3l1kLoxmAm4NyXMom7g81EIoBZ1KAWtroZQ0e6qqJhrQum78HMxJpl2yVBqY5x/D
crBS5ZVbCia9mfPGnTVjZj4zxd9JbMr0C55ujbQIPio3tzQ91v0KcM3NzJ+9ba3h
bS/OIB0g4os+YvQLhIZD0Ab8xyALUbMgCwa7Qq5tfJH/N+xD3wbPQyWZZVpo6l8t
lijrw4NFNuUkZe56+L2bHkAiJmneXPyQE73Xj9gH3f+sPT57Ib0Res9IDS27QN45
HqXkJJZbqzN9XOk9SpwkD09uoEnpbGaKbQIrljLlnYjfJ5/pP2HSzHqM+duUaesK
Wic7yIsY2YmWwi8mbvg7iWYdafQtxzm4DP5YZH9RvNjeCvA+GQbHJgjew6rEYQ5b
KnuaHVJhyMB9i+cqo1Sp50xL0iacQCkjMzz2Qdhii4lydOfkROrbRNcfSBUk7fcy
InyRMHIP7Ca8hym+3ivZVSfGiYVB+t7DN3yzy5bkciXIH8e9GfhTLStn9bByTtiV
Ljhcls5i5xdSx9MZ/li+OMUXuhkDiV6mhRvKdSz0CAOyjn1bIF5tvUBFGuv+liRT
RTuEboiGDh6r+0KAWzeW/UwlOzAhWaCE9zETBML7qnkfzzKSHKswizxgoBHE4q5k
ztplbzYw89kj6t14bYc0jjMaXAvWlHk9zzV5qTRuGksL08Qs0G0FgZZBL5sneo0Y
rzccUOmlJyaxo5ENuPPxivYyMl4K8iqlWY+rATixhVCiWdJEM9ziSS+PXq3CUohk
R76yLgLuCmHVoa3wJ3teHgDDGRacdwxAPH187lIjI1nh+X2/WsOlnXYx6qvRjdT1
zE6IkvycjORzen7pFYItQghJqoUng86j4iEbzExytl0IWtDGeLNG+fRQj/NHKdMr
0AaeQa/W+Qqi8g3GiW1/OylSCsg5f7DLpglCy/UasexM5ac1E/rQSZNneUgW7ltc
WDSlxsnWvXXxEKuZGJr2oJ2Duj1ZjfVaJeLljyOR3fSGONwp02ehDw28xEhDGERq
r2Hk4b7Cnk5afoW8rZvDmCXpYwOBokUtuQnSJPN3JJPAG4QBHL0i6/SO4xFidPru
SWhnRZQ3WuYf6X3jiHKLHZFTNJ8MM2rjA+rJfBvscUaHuUUDao9io+Dqk+LnSw6N
a2rhAplvhKQvFJVqVvj7BEQ8Y1Nh5fkoBSq14s/g1BLZ8dNHSpevEt8t88zFPFFb
HPSSMF/wmT9+RZhRWsQqIg67h5GXIi21vuJ2sLhHB8rrl1Our9Ergx6S2fbkjOzZ
BuaWC0p1zLDiXQEkcsXmkpQirfDThHduPEZDlnMuXAe7gGb81294CrunT8EWvE/f
BIbELvoTFd4tLFOewxglcNPjVBVx8KTDEw/fROykrz/MziEPQxlozJGVPOdMdjGb
eRqSu0Wk/YLGCBrs0VLpsrmADi0ZiS9bvtc1cO/NGuiVLa0VEzHwO7FP4wNdY818
YjuEJD6Ket/B5II/GWK41tHm0sPx+oHY0+3TdnQIvE0xXZkE2Qyuo00Rp7aegQVe
oIZuj6H3dUp/nz7heBEj3D1MqJeSR1Ht+/7pyGXE7sNvKoqUN2c2ibAmyZX8n6K4
RUAFrOTIXhjnC/K+eB9ZYESzm88Mu0sf3iebMtrnAnHF1pa36pZmOe5IISZBA8BW
0MUEAhur4FCtL7k447Hi7ZFsG9TDTL91OUVww2AWjaFOTVFVhZyF0E8W8lhxquGK
45j/K1ektROqSsY2t1e53nbIsLVEVdkr7bmGL1IZwywIRAZvY51FwaDWuY8coh/d
zgs5i+6ZskgHvgdo9CKeQ/vqOEbDRDt8srsNYTR20Ct99XOOKFtj/4TQgfkifgSq
rAz09qS7oEcU4zhwTH1TcEfsM9qSIZbvrAMYkjvnZ0pL9pvAmWJcwBotDrlfjKWW
+EjtevUEp7SWB6IK80MyyGhlMqJame6aIOZACZg6BVZuP3Xq78hOXHl3uJEEwr/F
//gHdt1IMAJI3HqqstdT+l/42UfZ4L9DJsBmESE0nRVOoHL7wOWHSgT9ApTQBEWG
Vrwvmh7fMKNcbm8xysnP4LlfrbSK/oYGb6JYs/QZh+0Vb9BQjEJV1ZJD/hCszIv9
zSoleNvvY6OyCSF1iHKUD6IZe9gQPanuu4zoRpptZ/UeUrm/sFZKEKkaA/t0d+0w
QyLtRUDfkjcJG4ysQTiGBlNm1F42UxsVqmKIZtvShZvvYGDkLICTKR3YetcxuOIB
9weKyIxT9qBg8XZ6aSZC3kBvsqCYf70rT4BshtmNguh/cLM79YXR4Q2Zx2G9eqgm
Q7qAJ2i8xwfl4jH8621PquWsGhmqM3gSkLhIK//JjKiuvTJFGrwNm6Fn5h4UCSRp
dXiCUpGKXIqUMPcLGWwCod7zihH/u1c9uA19Wd67mKRAzymC+MtgF1QiYM7+i2/k
44apC3KjH9X4uxWM7ODYz0dmHLNlDj4Ln8SOW3fthU3ASv7YqmLyf0mX26ktsQib
r+sU9DCvrW+dgcDgovfFhtKZcJCqqUkWZsN4j2Y0e76W3QO4HxC0j0yHxvGbfv+X
rRY0DxRGvBUXE6xpCv1wlDPaGgTy8XsfE65AQRZRpp8YLbfN1FTkcw71BMK1cq0t
dgIQoO07N5tjm94iqwiKMIo69ia8aV2sBw9Wfc4P6odm6q4yxm7aqJNmAJ3iB0SX
KoALuLBwC8dCtccj01jO4PkfIHydF5R4ixlYeKZAniF0Je/I3eF1QuOSdqirCmFR
XH8EGo+AaOOPRHOX7GMmPPknyu3v9F4p3ueUHtQHQQJjnP1z0e1zdXJfuD3nkdfe
mAYBg1EcyHxduEvX4iRe/RnVbQNG+9we44bqy4QPTq7bvqq2E/1gWa8hz+C+JZdx
V7tFJpcZweI/hyFxjnnIn7NPiK27nZHwQPCPJdvoXFNb82d431r8hD1WiZBFd81F
KKwXsTxK1cAPB59jJLg9pyj7kNmGb4VcZXHP8ECCM3EViFqBqMiVF5WFM+qWXoTK
/In3+wd0xCpB1gKbuXJfxjaz1WqmF0i0NfyH4RrvGNZjWrKRTgpLPPh/ParrLFlx
+iIijZUR+hhZkfUhOQBw/aP2HJA7WoBWMBu+dOos7tuBA8j1/DG69QnUBiu8YB6w
o73wXr4tDuyNDB0dioJAmOL10rVZ4IBqLDnK9TpKuuUuvL4rGB2CA23M6ELEeZTl
urrhpnNdtb6i9mLr6V3uCm0JFL2dOIuPOXOAZZvh+CUXWfJh70l/cZ7qDU+O3VvQ
3Z3pkMlF5s31bLHALnpAdqhR6HFG95S7qHG3+c4cEeNEb0Du10Kiv+71HSkF9G+E
t7h8Lp1joSl44rujYAKkGBZF4mAYE4FIm12Qh+mUIg3qPtIQFVrF6KFSGn5bFgz6
OOl8KrOsA0AA0m7AiFzIn6QQTZZ+qgmLyZR0neNqMwMounHq7Eq6fUChV33fqFFT
Qu3VSYA8+nhyAwrdNRYjJM9w4W62eEG8qaHD6riwbhW/Umu3UmYWNdepkd4/ZA6L
VknNbckQtFxEfhJw9w3LwPrqBjQf6n2DEzggdA158ApAA3728nsxNAwllhnTNJgU
O1jHHuLYeyTBpqkQln/aCvpOOj/g5UnyB869BBF9ZzOIV8BrEUwLesQzbzCF65RU
B4OHYXlahasjzatIuvA+4aSsAE6gq3UMd7qI/nYOnSY9j2a0rCd+2aT2GR1QUbNQ
SauvY0ffx7nCd6vKb6JNFDQJQE3DpzgrT8cn+QV9qQkCLVsoswpdjoYVC6aqca4v
s3I+UuT1OP8emmETlMQjsctLxfmL2BbG5D1bDA1KGK2V9hD18zxsNYQIqlMgF5Rj
dANkQXGmZkXJ4NEphazgNWtUnNnp7twaP6G1aHBv+5MGTfYi4HTx7WlZ5zlfzu7C
evOhlc0R5c5ymJyx/MRgpQecz5ZCgyUXew+Urm+Snkvj+dpmouu7R+GjNmikRTd3
bj7ql6vTzMVetVAeLcZ6txvP9KQqzhiVJtzuPgj8AHmAnXjCl0685fejDOvTfnVn
pTBKRMkWbLjoRjfh9N/fw3TMnWaysOTJH1GtejhNxYAKpKqT/PaHLDbvgFFIrlo1
7nV0Og4Bp9cWwkVaAxIa2PghUL9zeLI91jf769F8kQYjSfy19hwrGwSmgERJnZZf
kUUszukKf9ZYxqn3INT93hJTyzwdmyVliAc4JeJMbgyPPR0lPvlT7YjbbSv8t7ja
TlZvnwfx8ihjsOMynF5Nlzu0YUkHKBJ055BLxInDBlamN7cSEP7KPonOwB6Gif/c
aretNqFfuLsx4ZZHNgkkWkhU3Q+yPGdCAysXhUshbZD7JAwyujU1/JqpzVQCitdn
59eiP1B980a35btuYUiyc4Bde+WCbwqQZ2ZIr5bimeT0STtmnPygPO55jg/pbaHn
75tWRHuVykqrBDa4mW66b/5BLH3CbV4GLwaixEotm7eZ7tLX5GxBEa/reJf+8tLD
/UUDTbKe5iKjjDwwMmKKRxsQcKx1AGNgTIkBwnaorGJdczorrPrqA73djm6OUZpa
ZUP9yxXCPYUmQtZZpwCJ4CRTKZLncW6HgOvQ7dGr1mLm/mdCJ8I5nTBaNAqmalhn
u5O3CsDYeYGBrWAxLNF+YVSlUVaenQ757tJSs2NScy8PMIkclqvle1LCv7VScsgc
w1AUybfFxemvuQS5dLoCoFANAGkxoMWAvAQJtjrsw/Mq8gg2mntopktVmJS1wGAo
hW/jyc4stjcNaKsn3UqOp30teyTc9+LW6WzS/blFoBPErl27FHUOPKK3S/fiFOHH
wTEgLnOrIms3WUqR3muFOg==
`pragma protect end_protected
