��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���Ox���0��?T�}�D�yBl98�锛�l	`�ġ	d}�:��PƸ����~��R��o�K�jV�,R����vy���3����O���Z�����g�̼A��v�{�7
��5�¾����B�C����������r}�:ش)qqa���·����BW�4����"V�CL�zhXo�e��6kT]xl(���%lT'�W���'�N�V#�L�`�`�Xy�6$���:��9I��ì=P��uS�I�w��������F��<��s��y�i�u�����ml�G")�O�4����}�,r��𯴢}�鑪 _@�y�Tkt}��8!�JŜ�>9��C �gl���-����{���Z�*� 9�[�B���c�M�͠�+�G�Yy"TGz_'l��2/;��	^F�/	b2�ܕ�Z���./k7iǶ�>��R nS�}O�i|�y��!��I*��@�%��v��%E�D���!Ч��`�:��b��8�o��a����'�:R�&Р�˞n�����n��.	�����n�~Ge��E"�L�H�E����BG�P�"
��Ao�X@�o.�<ص�]�D	ؼ��w~@�h`��9ug2�4�GZI4�i�:v�����)�.�r-Sn��LҎ9�2�~�H��I���%c�<J�
s��6EX?���9��[:��䢽0gӛ;3�G���db �p�ǲ��4h�	���w��e �I��]oF+��Q@T�$�����i��x�Wz�J~H��fԪ!��J�a�|��Y�j\
?���fc�����J+�N���9�us�^��Y�a0Z���i�[�;iu��}��/�6$C���(�1�ͭ�^���g�]���}��K��A;clOV3 ��pc�Q�p5���:V�����-�4��3�5 hZ�h���]�Zn�ᑈ�b�y��]�	��jn�����ݛL�e��[<�2�h��P�I:.p�@�H��˓S��r-���j�H�KN���R��Ж�)��Զ�z��sy��ȇ��MnD%�t"�υ�ê�L�Ք�*�\�ʂG'L{B�׿F������et� ,]��G�[�;)}=���+�C�U��?����c�:�
����!]�'(��mquh��J8+�=�&�������� J{r�E0#���=n=��Y�9�!H���ٔ�;��O_&�$��i�Ɗ���ռ!���J��0N17�@��x��g�Z-{#�7�r�z��~�Fw�ޝ�Tа�TX(����u�*�U�ȭY�.�8�a�C��8(����!�Y�?.� s�[�z��.5��O_�3�&�zj��z �v?��( s����j�D��ܦ�Ym���-5XѳP��r�.��|m����A�K�V!$���A4W��n�o.�Рd�����C'7���������wߎ��Q�=eDhb'9�^��p��	z}.���.x�=,o�#M�R�c���i��G�F���3�(�jx���g�,pt���#����p����X�J
"�gA�4��Yr�k��ٌ�g!C��Z�C�T��?��%���``�'Jo.r�����lX���O^��2�'�ї+z]�[��
���@�[0��q����4��@��� .\{P�n�܅oȑ�j+�:/��dZ�W��J[�mKe$&7��w�D�]�s��0◡ �Ѡp|hQ�O����˦;Py��5c�q=Z;|�.P�_��4N1���d�+���Q���t{�kc����edU*�W���?��CU�,=A3��<5���ϯ�0�9�T���L�9���nl����E�XC:�I8;Ҏ��c��LT4��A�֜F?'��*C�(ʪ�M�"!#��S��r�� ��l���;��:�6�<|A�.�u�h���n�	�:���I3�e+?���t=飕��ÌP���*�D�+`�噯]�aU��N*��D�lB\{��ջE�}������5�rPե��]%�cu���uIV��[.v�e4�(bs.A��xV�)�5���4t�����\��,ȫC��w7a嫑�;��=*���j�v=NL����0���+/E/؎���-�G�@#U���G+�x�7��r��jI�b�8В��<����u7�f�W��2D�}�"�Ջ�L���N�H��L&�E�<!��6�ܓ��,f��X<�(���;5�a�P6�bq��~n!��)a>�r&uG������w֞u>8 *%��W<�H��C��i3�.�B�����m����A�?�3��/��!c�h���*;ƀ'\J��z�4�3%iƔDD�Ī�D`h��}��FM�=�������ף���(��&���ݑ�X�*��OOP��*x�v.����G����l*�7읧��'�:�#�~���«(����2p8~�W�`"Dޥ*��Gv��_&XK��Z5�.�]=wd�ט��R r���Dz;�D?)%F���͊9�@�S0UGChV
W�6�|P�����K���#eD��-3��Ӡ.�W2\
��s��$iý��N�s�?�.�Q�$�;��k�"�m<]�,C�dT�R�!� ,�"�V/������K�%�aut�$�-`� �"W���F4*q ¼z~|�7m���n��U0�s;�1<.*nj�/�o�ϐ�=����{��H�`�m~�	}E�n�,o\כ����nck�q�2y��]�,!}�DQ_�wr	�$aϚH�5̱�6шA�\/C�Y�$Q��&��ȖS����}(# ���0[�����u<��lР�6��(7t��4����E7�=I0�R��^�b]�D����}��FW��2��,aN��X���C���}����e�Aj%ԡ`l��*���I{V���|g��x�l̬�Ү����\Qe7Lo����0KB)���+��͒��6�c�w���z���V8u$�1�A�ԩy��K0��~�$2`��;y� b�1�g�)Ϝ�w�f���X0A��i�E%G�͚§]���'�Ɯr�f?u���j�N`��S��P#�� ���
�8��,psx��1ԽPz�}]�F�V@NO���/)T��~[P�"Խ}3G�^�T�H7��M�9��L�p2$B$���2�=%���޴ p�_�I���O�(���%6	BK��S ��R�M��x�����س�rG�QJP(7� }0�-���W�L���J��}��񁫢��0��N��+�+4�"��g������QAQ����]�2�#�',��a�/��� ��iHӺ0E�ܕyjti�C�>�=��遮�ɬ�U��@41�_}9%����K���z�4*���)�B^d��µPV��k@#���K�Z:<�T�%g=��h��ʘ���ۨ�ƚr:�D���G�a��yexd $}�"�m��0����p����#\%�^�t�C��<F�9�����0o`��Y�jw�D�}T~Qk]Ji8I/��wOx��8���!!����x�'��⌡]�w=K6H=j��	�Z�_f�|;P1v��ΰ8������V�#�����D�X�$�Aӑ� ���_ܯA������ĺM nݣ"��k�ۅ. N�&����R��U�6�Ag�Jy @�8��}�"&�NY]�9�o�WGE
�saw�a���HT鬳d-����v�c��&�qY�4$�iJm���.�{^�����Aԋk9�n�
5�]1�ǥ2c�#�'�$]q�4�|�:e��0�$ї\�||���D�H�{�#���q��f�3��2�Sͼ`�D�[�	Rj��c��k뵊��gh�L��B�EX�p��l��ۭ8��]h,��a�dx��-�j���ҁ/� ��
|����p�6��;�Z������STV51M���)�w4P�B?Ʌ�[���'H�;�fr�
Y���?h���v߂�1�ǿʬ�������0��s�`�t�m2��j�5�O�����ĩ������iȂ�:�J��)��hP����$�R�@�vI�Z��>8s���_������aI�^�j��2�#�6o{f�"�V��\��1�ޏ}SN�ϟج���؃��T�q�"��K�;��2�t�]��-�ʰ����V;��bE=�3y�3�o3��_Β=�=��k,��ޛN ��F��b��yZ��y�D�|��� �2Ü�Z����7Gc�*`�^@�TS0P�?��mh��&8d�Z�+3��U����^����BA��r ���3����M��sL��`C\5�+��;����d]����K�ӹ�K�T	c ?)��G�DO��3"���#��@^��Ҹ�9�1a#f�dA|��F�њJ�7�.��f �~V�Կ��N�|aP���ń����j!R��8�p�����A��0m�yq�����g�O1���/���a���u�/�T X5��xm�M�5Σ�f�͘^��?0/� >1'ߘ�
!�fY�~+�\�;GY~7��'��&����jH�x(��q7ԺF?*�F$�mP�Z��������߭0-�$�Hū�>^�z"w]0 3�.*�E(�4YZs���1Ӵm�L|�UX��,����|������~��b��.�d�{�r�V}_`6q �0�s�oc��nB���R�O ����AE}G�61�~"��a�������3F2ZR)+U�8![���D!�N���ģ�n�& �!))��=b�PW<�����ufcg���Q&���YX+٢j\�-[,`Z����Od�d��N��U��{�&�7�p|��-��ӘYG"2�p<U�o�Y�'�Sc��h	�U��)�L1ze�y4'�*��C�e�:��;]��JRGv��V�hV��z,'iHS�]��j�����N�؋.o�������b~(����$Y�Xr3�4yjY�}�����|�(`t�U�|l����
���F%uC�@<�^w�r��L�cdH9˓܅y��RuL}�$7<Y9)x��Y^�B��>1��g�v���Hl'���˰`I}G��O����︗cB���s'��r�j�#�(�/H�n�6���w71+�}8����F'�x�aH�����`1&��d,���u0�pr뢏@��� 7�y�$.�L�����:H�zz8s�$���W􉹮*�B\�,�d�+�?����Z����qL��di:��6{
���Wl�lN�a�zd��y�L�D�2w.�.@>=��V>Z�X�_[���$����e�+�K��u��L	q����?��"�i������G�/f���H�wh�Ԛ����l ��~���4��]�7j>�#�� b�D"���ն��3�|���� V��N?�
w2=��E[�a�����r�m)��~���i���z��a}�z3W<J-�qUI��P��(-�)����d]%N�6i=\���qZ�����w�WE�q�v��0�z�j&��aϗS�7���� e���]�e(=��~���c�'�U���z�孢>��F���I�������x�MU?��v�6��K�R�ˈ�����m=t�*�R�G��۫��CJ2�[�(�kq7�m[����ъ`9�S�A��Ju�e.�y�K�K�=S�h�]���x�e�e��r��k�dF:>����*9}�絍�J�C���!�)^��P+�~e-�U�{0�4x
=�^��K���ڿĿ�����Z�2�s�:���b�[٩�Ťh�ra�+��S[1]X~z6�7DoӘ[3��3����E�Q�/;�?�VA�C�Ʊ9��;3�Es��t��>8�h�e�Or�&Ά�G��_���kSs�f����nY�e,r%��wS��l1Xo�cN�����~��׆�+��#j�D�O��L?��������K�c����e� ��L�EXv���`�9���T�3�Ɂ�A���,�}���̫�8��?5J�!>������*?���P�nշ��f�X ��1nZ�I?NeD�k!в�6����qp�Y�������(1=��i���η�m{u�����_ވV@�v�|2
ZB.(~3��h��i�-�S5����r�#�|��\�����y������ȍn�D�-ꖩ¦9�F"��P�8�څ��!������@�R�>���ޞ��>��%P�6��f����U4����|���Z�:P6��%���tF�&G̲��.���0��~LG�P�r|�%o���A�گ�O����Ebn�X~/��M��|��Ԁ "�$$ݘ�<L!:~��̐�d���"%)FV�dr�7(���Xv%^�mH⦺~�{�D��h��
�r�ۤ���Xzy��/;uP�J�MVX��Ɣ��ǭr��|1��ܱt9P��:-H���@:�n0��J�Rd���+A9@��D3=w�L�!��6��z� ���W�P�5O�������}O��x߯��PE\�×����{vRf��9Dp�����,���
i�o"Z�3^O�چ��=(ܜs@������T�R!� "*I`J�74���{�좫#�n��B���G3�7���wz��W6���Q[re2%�j�z����e6�n�<s�u��$�{�JF�.׮����8�?�M��H��e��8��@��
��=��iڑ~�"#�JN7�n^ko�|ެ�q~�|�gk��fUR���SqUX�P�4
��y�Q�L��GMw����k�Vrc�d ������%<��:�HC�X܉��=7�~L"�!Cw� w�W�c���P'�L~��d	�Ag����M�Y#)\�r��_$�����h� z�bR3d�)F�vx�h�L\ˤS�L�F8�G�Ռ���~	O�]��Ce���N�7�����m��ߺ�CM���۞�E�J�2���#[ho��M��h�P�vm��zO�QY�u?�	J�DE�Cʂ��b??���eW��1g֭�
仺q����ѱ���Q��1@|oT��)J�e������� 5X�}�2�L@��9	�_o�{��=����.
l#H����=j(��@m���
��,�"Q�p{�G̀6"|�ԣ���x��`��Ӄ��Pm\�J���ʛYG���޸	[i������t�UEv���92?U�l�t�2��O�};�:#n���Sx!ޤj��#X�1��� ;ͷW���ԛNh�
=]R~����)Lfᴝ��8QA��C����a_��⋨�����[Q{.��@g���.��=-Ĵ����c���S��r�!�ZyN�� �eSǧsJSxF�s��¤�"s�����]ոL��Mw�7"G0ث���?)��L�#��]���O��)\<0�+^��H�u��L��!n Tu�-a1���>ò+�Q��~�d�`�͋��)VD'��	�,��Cy4�v���[0!n÷;���4����6�Nw��G!�����#?��,q�Bܬ��m��������5���E�_˂��S��;���WIƻv�@q��=�G�0�˕)Ƒ.�-Yb�Yj�1O���vX��xA�����!�T�.�ǂ?��1��$L�0^����.�Z��>Cxn�c"Qq��Η�/g��N&�I,%[^ݬR�R'j��iij,���]'GzZ�9������}ȿ��l=v�Lr ���3X�<��z��(���M#y6�%-�A���߳�1�M������춻<�c����5�\��q<n�� 2��D���a���-9T�El��!M�|�s���[#����j�;�76&n�э�<) �UT&Uf&�CP�Z9�&�!d1�w� dL��._Q�o�@4#A��5�W٠0+�4ɮ|��?Q2�kH[�(��U������I�{r͸w����?TAs��26Y[Fl\:��A�Ƥ�
��,/IwԜ��A���j�J���$����f��$���ȴ�vLz���J�6
9�� ��I�:K!�s:5�qk��p蝇&	��	��RNsx���l�~4E�?u��p�} �}W^E�LWMY_+�s��B���R��͐ ���hU-z��R഍@d����A�=�4i��W���e��?A�;��\JL}���Md�!����B�K��������La8�赿w�:�&^�&�v��Q��Y"&���		���X����@����f]�� ��b��*d[�w�տ��'���Ac�� ������$QsD�9�kͿM�J��֌�w��]&�����\N��epN�r��kƢ��7�F ���1�&�I,�)n;;\#��O�y]R�9����D1�K��o�=�i�d�,�(Vf�' �HZŦ��t����Bt�p��Ǯ��1���R<�fd���U����j��+\��ڤ�:��ʏ����?7�Gs�;P�78���  ��0 �kU�O�h���J��>he���	*��Rq��J/�{tr����)�0�
>fo1�*��]DV����?d��Ԍ<�_ʛ���]�;9n�s�[��P�|D��Uo�i��|1�����D��Z%O�+	�7��ء��h̚�����\�
�[r�x���/=�OE��o��FW��y9�IX'B����LkX����{�@�)�v���ˋ�?;���['`��
Ϳ�.ԓ�S7��XѼ�[s��'�X�S�Y�3�<���'�3�e�gT^�����m��9���<�7�(N�����sXm1P��%{p]蝙����yZ�'�|�g�x���-�:"�<�s�M��7���RÈ�����n�pG?m'���̬��Ò���"�� �*��F�N?Q̨���~O@�c���f��5"ZƁ	��އ��(p �ME�s��l���T��3M�DS��ۜ�1���i�j ?��(� 9F�0�u3ά�J���k�$��|�ܭw�pJ}�v���2q��]H�B|��~]�����C�c̎ה`�t���DO�����;D9��(�^�F�{#uO�2#��ׁhu*�����{���X�<������č7�3OT VBB����TjsM.�NVB�d��5�ho���8���Jb�I���[�؍�1�i����K�N7�gz��Čf;)��ON#榑�]:"&[��=��j�$@A�/ȫ��4��^v��ĢW�����E������+^�8�$��!���<F-d\M@���X!�ϫ�v
�w\�w���`���v1�~=�2�;	6�4!0���W!�l��O�q�D�=�z���'ېnVys��s�.W܌j�l�H�
�GM��$ CBd37/X�\/��L�<��Q�W*���=����5������e��v`�Mc��5����T��M~���ɩ�i�W%�2(c�x^�������	�|5�L�D� ��M\�~6%B�)7��?����a�Hwa����5�M��$%�8��q���]��Hw�L%Z��/�Kft������Hxl�1�>��0�3'���*W�u#��ỌUѪ��,J����k��r�<�f�cr�y��t�B�k�OpyEO(tQS�G Cuu�>��[��׍�����w# �Q�1���5zݡ�3Ξ�R�+)b���k����#�p��a�L�7���D��x6�}i×ȉ�7�P$I<A	�N.���U�^��Ю��vzsbl���{�6DmS~�^�t���EI����4�e%�&��%����>y�Y��~���2¹��t�FK�{s��u%� ��As:�����j�I�IG@"l�3�}޺�d�]�GI.�9�!MCoZ���4xb���jU����l�
��
�(���)D5�0�9zA� I�����e�#�<������3ϭT룼8?ƞ�K!�\]Kd���C����V&���`fq(�����g,n�7O[B4 �T��2�i�Ȑ��Ċs�ĭ���xȎ�z��H��e�,��]��خ����5�Zb=a	��и�w�<k��T{��OЄZѧ��<�?!X���|@���p�%c��C_&ʡ���8W�&���t,$@A$�a��bD�N�1���<}<��l	����"��2V���a�E�!��
_TӸX-����'m}3ޭ����e����M�k_ĵ��,�VG?C���޹����Zf�9�{�]-L�5�}=W�+��0��b�e����h�`m7�rP����N��>ou#l��w-e�&p�O���]��U���db*.�53�<����32+ٴM�`R՛6$����p!�,��U�ס�ޏ�h3�d�zOI� )���5�/��1>�g���b���f�,�w��K:����G�n��g�:@ӿy��f��=g&���!h�w'6Zn�gY��7���Y �%7V�i�d&�����	޼�;����n��h�W�5��-�k ��l�F�
\f�m$���5ڙ����Cb�QL�3�����lՍAkAǬN%q�ǁPOc�/���_�y�U�ˣ��!��#Ù%?"
;����ݦ�K�)�R`x���r�=���#`A`������	�^���V~S�D�Õ"W�FWvu�ud%I|3���*-`Ԩ�E�6�R'��Ny9��dŜ]lwle
˿���#�A���������u��H��k[��Fmښ��_G}�����5�N[���qp�`L������2�� !��,��9�9��L�͗��ĥ}��.���^U���jH�8�x툅A��g�Io8�֓I��ł����y8P�1
fxݹ��7K�(,�j�`����|�=��@XI;�}�PZ,��y�7�"�<5z6o�Md{Z�G�w����o�#I(}8��/L���Q��X<3��۾r&;?u���_}��\C�T��22'V���(��������}o�-�QY�啎4�w�#�u���H�煍	������*���pD<J��XZo�y'��'6�
������>i�5�0�1���M�������rÆ�!�Vk���D@k���-ȟ@eR���1��Q��}���0��̲���1�d��#@!�\O:IÙշ�3\��̼b�L�d�:�%���2G���>�fO��j��/3��sZ�E�[*�	"���D9-��� /�v°�k��]M�b.��3H0x���/��K?�NV��1�Fl���O����E��$lo��gD�a�|q<�8�e
�p<�?V�B_����y����_�Xf��L�̻��>��h/*I;(��"g��������t>1i�zi��7{�E��|W��Ve��ᕜ�%�����]<��M�aZ\�i�C�u?����/H���v3M3�L�ci��w���1�,��,$�!�/L���!@>Ȱ��)���� �4s��[���7#W� Nk���!�^G^+�C%v���Pƹ��c�b��6��\�P�
Un�$YIִ��w*���	Ea�|%��A��t>����_X}��@~Ӟ#��ս@���|��5���U$���1m�<|�)���5#�;�#��+`�-\�|x����f�/���P�'���
�I󓌶f���_'�ǝ�w�d���~���
��l�gu�n����P�x0�&�u6*S�F7D��ԍ�����k��8P��0��-��*�s�fo�G��G���m٩��*x�����>3T�W�?�kː7;��oxz��O��-a�f&�(v��$3�j^�zc�O�^�����;*w��ANg��^�;*�/� =6���Kˋv<P��hS��J��,��.)�M��=�Q��	E4��}��[| ��p�oUʼ�6*V�\�d_M �
�DWds�X���%�������Ji�ёi�N�c	�����IMƎ4��*��������ROT�O�\����;#���_��v~C7tݘy�V�����2�D��]@��>���~�1����S�X5_"�?��/{I@���p�[��'G�����`�4x~X�����#�k�~>���|�����fb���7X��T��\��<�Jᆤ�Q��&���Џ̊N���f����8��C�"�jr�ۍ�+��aRN������ߟ�x�L�*��W7ٯ��o�h�j��=8)�)��kB6�Ӭ��Ր��9�����n��ũ�c�PA�
N���yG���?b,
�c԰�&?��ۂ¥��rN>�P8�����Q����@t�C�%���ܱ�U���a��
݊�|�Q���kD�&�f�w��*K}1l�d��&�*�U�]'��	:�:s/x�ť��&��ŎZ ~~\�i9�?Ԟ'�S1YHW�iqK�Į�ʡ�������Je݁p�}4
��Kr!��ˇD���鴠3�P�z����*>�|{[ɧ�C:Q�C�'�vY��*�&�#f������jF�I�L{��Xطl��C�Mv�R6���v���L�LZ�Ȱ~&u2���U��i �h���n��@PÝ*�!�K�)�A��iw�OO߳JG�h!�`���!�Ъ�2��4�O2�X��s9�.YIy�SRO�#�-���~��*:��ng�h
R��8*4N��,��U|��%Cֽ��2(v(�I�S�ޣ��Ô}"]~�p㧨�s<RJ=ȻτT��Q]<h�PKT���O�҂��~�˘�:�?��sF������E%aDTG.���,������ёѡ��QJ�y���Dh*�Ğ�3@5�o���H�tY�NL�Эm���p��Ik။Rb�ݜ�T�F�,��}Џ��`�#m���K�?�7��K����t�3���:9�BwcP��R�5ax\���3����c��?�
ZD/.���3u$#��k���a�
{�c�(�Hl�M�Х�Q|���ل�0$ Gt?�=��j��uG���I��k�5"��'�z�R����)4�|�j0+�00�`�B���}�ڙJ�;�_�8��6�����\��)f�;DI�L�G���Ӌ�i)���_�dQ���� ma�NK�����酣�j)l����dC:N6cIC����B6x���/N��b��z-�Bh�-�x���\@��l�\s���&n?H�B��weGXN-K��rD�m���{�
�*�*��9�q����=c�]�\g�_��ESt^��N9[ jT��۟�M�D@qNx�Gµ�5{���jm������狂ƭ� ��7;���o�O�Z��g��qJ�{5?<�8u6��&o�s���yV�<�j��88��1���mB萢�D�3��o������n2�D�E��%��N�a4Җ��sn�AK�S��;� ���5U���c���4��v�)!&�Ц����t.5➦����GS��>V��ʏd��5-n��j�먱��/v͇��T��L�`��?a(�l%�G�ɗ�<U�x�V�*rT��H6� T�o�_�(������G7v��w�,{��;�J��%xo<i�]:�|��%��߇YoM�3�R���R���+C����(���`�f��&L���k�oUS�-��^�v��@���	t8
+��C����&p.-|�R3_4���Z��1�'�aSX�Q$g�ʲ.IC��)%3��7^��*K��h{f���W�myyա:T�i����hs)z*� S÷�iؘ�$����b�����$��= ��7�j�n蔫���^�/�<�D+�e�ŀ`�v+�r�ת	a�l�7�%l���\�7:[};�}R�a��Wzt��e7��T�Rr���Q\���|=����bi���?���8	2�b�x��j"O��!gD�z�o�}2�4:S���pe~�)�Dq']���~�~aq�&ك����������N]��pn�+�B��b��׭�(���Lڨ�[���Q�ը>8~	=����yi�l�#a�u7� G>(Z��5��>,�ް��E�\�*�h֪:�P�-]���k��H\Y5�y7h1H^�u����X�Y����5�ۻ��c����zخ�uٻ%��
�in�a,�V^���h~�q�9M���D�>��8�{���?)5@�U=E����*����Fb��3��.�`�̯�(�WF�e<Q�`승j������]i� ���T����`�$�ipuy�g����+9^OX�hG�pb�-�t)j���kX�Q��k�o�KH�Mi����#ɬ��z�17��c��LR��z*Jrƿ�Weĺ�q8�U�,����2��H$�(	��lh�W��G�D�4��f��e�v��/\j�������b_o{��D,~L�B��N�4R�,�Q�4�d<�@�[I�?ٻfH�%����w�į�����A5�����PN����Od�%��MHҎ�T��:�ZU���S�gJb�]����7�HY?xʄx�]��S)�"eA���$�]�s����J��VΕ���jg��a�6����:�f�Ks���w�C��dh��b�.]��$�U��ٴ/�]�����XM}�h�Df}�ǽ��?��&.g�l�f�j�"�#����a+/I5����YW4:qO�W�|����(�=_s�Z"7��'��c�q�],=���hv>���ګ|�ao�7��TM脄/�\����|¢N
"Y+��������Y�mr�����#�%rP�L��V��qó�D;�:M�f;�Ue�7�R�qE^:�]r�[��>�qE�Z�if[m��a��n��C$�����_�45˿��=�
�~U�xJ��_`f��I_���k���.���(�����}���+w[�wL��C�]����wa�P��akcF�:��ᅲ�Wu5Kg8�lű@�!�� ���N�>S�)��ϛ�B��鞪�f$�Rj3��W�5�JbI��:w� "��}�<Y5�B����m�_ˈ�`��-���''��4�Ԣ����