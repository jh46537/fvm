��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�Y�f�ʴ��d�m���8P&B�� ��
�˿F!����i�xL���G)35�У0�Y6ɓL7ɶ�4[�Z��K!�Rʶ�������(��骕�Bwr!.�FM�=��zL��K���� ��@�O�iL"��:�
�'������l�x��|�ߵm�~F��q �t�E(�FbS�	�i��>=�!�Կ��_s}��2p2A!�gҲ[��\2<E95�.��S�����zj
k�d����a��tP�a&o��d�Γ_��P|�kJ�g3*���3��ۭD��q���2�/L>��n�I�����sk���yd�nE�I/�=]��1ۍ��#T}Va�Ĳ}T�S���}�:��r���Q��mP�L_�mz�3m�,^kr��B�vN�@�$�z�&gOE�o!�$�@��F����n"��OS��h4�+�Z�E/Q&�(�Ok�D	��3�ǣ]���=���Y��A 7��^�?�����*=��������w_=���g�!��R��i��:q/��=~��,C+(�Ag�%=J{p���>��޼�w� �YiUm�g@���H�jn�Ix+�=���6�S.��F'	���{a.��J�k<�W�ht���V�o�wVZ��<�u�L��װV��ȁ �8�N!� ^|5�$�~M\����Z$�3��^�ˀ��Wd�vǵ���ˌa��+% ��Ҥb���G������D1��CH܇�m$�q��(�uS�_z}�`j��}Z�����C�Y����/��R�4$�1_&��W=�[찙�t�F����_F�(�`��!���>�ǈ2pR������C����#�1�bѢ�}��r�����syMՈ8���� ىnƵ��IHB�m/ju��h,3���૏���д�[z:���M6����8o�c�G #�9�z��eN�$�QwY�����m�=�I�Qh����G-�+���g5�<��Z����?�ְ?^K��>�F���*� �ڴ>�c��ɷQ�t_��H��:�Pkǉl���41�e�<fũ���J��$,ϧm�� �6) LM?L�س�qa�]q�����0+�F�F-2|�S���7�g��RG��_a��CNЁ�G�ۀՁ���	>qƪ�_��G�n���`���<l�X��~g�9bM�o凸���n�J�
�^����-�6�Q��+��RvD�d�C2�v �?$�������<�j�Y�Gr����0�E1O�$U^18S��Y,��}�������
]\p9A{��5�M��{�L�����ŏ��AQi�px�gQh�
Qk��y��q(_Rn�9�$ξʄ�c�ԾM.�4=�ᱎv�6�b�A����q���^F'F�wl	���I�]��3Ӂ�;$А.H�`�����0��Y�o��|��5��Bԗ{�Y����|�O"���\��kƍ�cA���[X�L���l٤���^j�_��D�4��-=�F�:�X��H08���u 5ڥu{��`��ف�<��ه��] Dm�u(��	X�q�-V\R���`�H$��H��C���ҳ�V���x���]
�ڹ��|x����Ot�2�K�E�@��� \"�^Q�hs�W;/��")߮<r�ӧb.��%�.l���B� J*���I�r�'�KJ���Ba�����*x�Ρ��('E��j�y���um��j[u�/�����G�ϫG��!+��¯�o
0��
�U���Di[�7�ڧԠF��|��+�!�Ho��[H%,|%4E�|����Ї�lG��RZ��M��gMCm��@+f_���Y��s�ay8{�k'*�k����c���>�	ɩ�e�ߧ0�tu�C��	Ǹ����hUnn�Ә