��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�=���,1�jӛXT�d݂��L�#��{_@cV�(���HUW��Y��gaW��l���9��6��?E���d����EŅ�����$�(|t g���O��o�m�wy^�e։����|�fk'�tC%��$P�v ��L)|e��� �T�Q�W��;U��4~��Lw5��nk��u����?��O�$�����j���d�Gd��5�l�zf��ei�aJ��"Z�63��~�b<C�r�0��-�,M�a��k���B�������d�]�Ս�B��"��hP��YW���-�{��"v�Tq8��d"n݁a���&OL8PVlL�1�h�T�v~٘?0�Oձ��� �
�.���i+���~�H�}vV/ׂ�g=���۪�l��+�؝$�Y��vX�[��ӌ�K��i�>���{+3�P��w{B��2nj��z��@���1�5(ހ4z�qߟ�LSUb�y�#L��D��F��*VE���6��N��
	�<��~���Ҋ��e|��3����_gM�H��S����!Ed�$�z���®�"iw����,�欵O�n>zZNm�z�Ӡ��XT�ɱ%4�L��m%,(%��M��'f��&�1e�9�W���*��i�3��v@�Q����3���ɲ����9q������D��Ƅ��T�AP{���˖>D�)�{�h�5�U�e�&F�F�D]�LI�E�{��_����/��h�}��t�>o��}%�N�m$h�>�q}	4S��ܤ�#��^ 3�q���Z(����O��Tej1r?��6f&<��T9�g�a���/(7�����j�JJ�<�N��l�a����]J��+Q@/�8]>�<��4�-��$&G�;볼���pӵ�Քo�w�����#y�JCod��	`�6f��+�6 ~_���� 2>ϛI8Ά��B��I#\�_u����F���]+�B�(�j[o\�!��,#�&�5�J�Tb�cjb4�wN+�tϣ2?a6h[[ۺ���C����K(�񅝟��ᆺ��t`���/�h��(]1{���W/����m\�6���N�x�j3cS�>kC+Zr���#�����1�7�y
��|�
�����R@#�2n�%��7���;� ,Y�3S.��f�9��	`�H|Yv�u�?�Rg&�����d!P�[ީƖ]�|.�+��o��7z�Fn���R�d���?j��f��8׆�Cv��Ä�U�w�×aM�Rq^�D$y�:��0���L9��{a��x,.�K/�f�ƼS�c��4@���:;gj�4�ϙM�R�|!�#����6�b��	��y�{ P���K�e�����Z�!�,BT��	��֩�ʝ
�d|�~ �"�j�U	��ҿdҰ^]��q�y��s+S��d����ц쎄y�d�2	cF�j �.=
�֠�I�ً	E�O]	��+Dן��DvO�կ)�)_�Q�#�y")�L��'�!;}.�����j�)A����K��(E����a��ߗ-}��8("�o�Ӿq.�t���J">�|��.oM��4)��-�uǿՁ�����Z@.��P�����yjq��!���=N�OŎ���c��B`1r3A���ZV']1�U�	�Y����1h�� ř�@g>�-1����wI�p�ROD��k06�yڍkr|����׺�x�0n��(Y�����1TeY�����9�&���}>�2�`��Wõ#���;LǪ���dT����dS�|i򂁄���N+���;].���7P�R�c�� ��J��2Xvu�"(]�h:���c�_vKu`���qh�DJ�Bq]?���@#��"*�gB��O�S3�/w�ٗvS*�n��I��\{$���[l���(�`�P�￝B�I�Fk p!�ȸ�x�Y���<5!5���m����ba���z���?R��1�B!]H�)���!�#��{L[B�e�<�ѣy���q$�
�M_�:pK��-��H7ШS���U�k�-	0b..\2F�Bb�A$��dMv�#+*�G$��D/�s%�3ӑչ��K�Z{�rh����>�\;&���:<l��҆m��P�C�	��=�H��q2�����Q���30��ɾ�]������Ϟg&�*�?˰�nڴ��g�G��f�����i8��"�'�Gz.GS�W��� |o�7ųh?3Վ3�m��F���:l���Տ4Q?�\�"+v������ނ�侾�������=�>�}���b*h�Ȓ��e�I��IѾ�ٿ��Y�}Q�x�ޯo^��+��
;�ҴI;pf!Y�������?����^���ی�*	m�`6���G�~QeEx ���>T�d\Lu�F)8,Hm���]>�Ay:���>���HO�p^Ix6�ukHͅˤVRbqc�&�Z�NǼ��M�-]T \U��4�� �/O㶟h86nO �,�Q�V�j��r=�@
V�r���d�CE��̆zHO	���u0\iv�!+]50��}���R�T7̞gV�_�GU��+��Qw�8�0m���4�\*��2��Z!1U����	P��nh�:::y����fE8�g�����R`
����щ�1M�yu��%�w,z��h��>c7|t��	�c�r�A;6��(��!��h�ٝj�X*��%{PitPw����X%��k������1�jћƗ�zzP!{n
gݩb$�4k���1Щv�S�N����\q�+:cB(7�MUͫ�� PW�D���`è��F,��f>���6��c|H^tH�s+ϐS��]�r|�9p{o*�R6o[��h����+民��[��k����
@C��oz1���q�0~�S�u𜖠�:����mI
���s��µ�����Pc5�cz�E0,�zGś����"�p�Ĩ5B�7�jx�g#�׆xQ>��3��h�H�`�tg~�/�@s��!QGQL����O=��/O�VWN
{p�z�P|����@�T3'�)PT0e��!���-G>�z�w���w+����(g?��0x�*���s)}�7�֛V�)W�1�P5MV%��f/8Ѷ�����ڻ.vq���G�ˇ������{GW�v�m;��h;�x��iM[��@h�S 2��*?/u���@��<>��iݟ <(��c�f��U���Snt�2��ЭU`������Q���w-�[Ɗ4l�l������J<r���Д��s�0�������&��U*U��ȷ�*����Z����N�{U;��~��@M2&}��,͒��;����Ae���ŷ� �U&CT���K}��C�?w���Q������f���r����~�J4�q:S�9x�X�QlO�����;M0b���L�G��y��;�+8�<bk��J�2=@0+BG
%�7Fj |S�=e��#��h��p'��f0�b�c���E)���R�"��(����M�Y��=6��T���\w��8�`<�NY�)�|V��,&�i�Ѧ���V��� ���$��8�Uɚ	y��nw�)��C�o��q&��P~l$6�9��\�wׅ��f�=�����.��E&��z�l�ط����0��&���&�`�4lL�*k#>�
p�4����[�2�HΧQ~��VIǾ$0A&̇3��}��8�g�%)�,��M`���y�|8�����y������r� ��"��ݘ�H��-	�������G��O\��MM=�ԅ�K+�����a���9�l��0쫯ٕԆD�jO�lרɠ��O���}iՀK�C��[��^�qY����1E%�LR����;�P�qT\��e9"	`��y���t�5d�\�d��%$� ���;�o��
	�p��'jݼs���-?	�D FkJ�x;�Q���*�������Զ�[t��^���?ּr�D�IPv�4�-��Q:��� ��$����za�%���{|*�D�x��ݡH�Z+�\�]͂W�l�W�0���8}�jAi+�\�ȢS��w�Gw�=O���K���ŏ�:5}�6��$
�v��=6,u]Ѯ���gzuW�_?HWV{�*&~�v���,_��t#|�����T����Ӕq�t<O�*�ꐸ�М�.D g��i�h���5�C'����Q��M���C��ۥJ��=��L̄@P�����ck�fQ�9�W�mf��q��M�@�2@�I���	���zZsI8�W�N暲����s�xđ�&K5�]���8[���$��pe?��rR�pi�v0�.8��� �xM��X~{����W�]��չ�f�S^r%0�Uc����NU�j�Z''�4҉'�\k
L=�r].�/j�Vo���&{E��v��.����/��=�[}���`�خ��n�j��L��^�E��Ɀ|D�[���Axi)�Xi�En����(<�"�%<(��Cy}e�}%�l2�t6���GO/�*�F�r�)zb��䄉�g{l��u��!� M)`G �f-d}V��Ƣ~��&���;2��}Us^�l�K���e{�ֆ��a|�%��@�D�������*8� ;��6g�Oaڤ���E��K�
���?��Q��r�:���Z��ü�����du���uR'>�t��4���E�G;��/�l������"�)�2f xȭm5���L�Xh����\�z����_M��m����8��pvali�Eΰ��K���K��R~;DeT+��K�D�<<?䘙��������m�S�~����h��\���ʽ@�d�^_6���'a�R��I�H��5.���L��gm]H���g�L0,"�u�[�+��h��wH��Go��!��^9y?�"����5�j�9����GB�B���yOԩH�������~���/�>b���Ȥ/�3]_� Wa��% 	�G6M�J]d�D<��f�H��(c��]��Di��ϗVVL<g�SBd�Ű��j�����VBT�<���}��ZkX�i'��*�P���HW.���W����6�ɥ���Y1V�����<Eh\���;h,��������څ�꣗Y�5�r��x� @Zp�"R�QF��=����ٖ�@��e���$Y��b=�/�a�&e�os;�