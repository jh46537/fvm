��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�Y�̞�������m�h�b����̘B�^��C�mE%�Z�
V{����è�c�;rC1Aű�_K8Qc�_��Ȓ�)?T+%��"��қ!TR�Z���|W�gD�̲M�"�:�,g.�kdΟwp���j����X3�Z�\���)���G�{�lM��������h�!�<�-�;0+��+섂'M�E/��L�����ό/N�88_T�5�\O��hg1,��me�dF�"Y�-��X���NOg�pP?�K?�ŦW���	�Ĕ���������YS���p����Å�9M�Spx1n����{�7�C#�������7YW.��?N��1"�s2�H�ƴ�H�˜�����H9 p�Z��{��T�|���n�P�&�
�1���xE�#H@��OF���O����uQ��fm.{p>�������5���n��GGKlp�j(�ͯ�Ur4-u ���ִ�&�t����T�Ƙ� ��0�o���b�eJ~>��n�~������&~� ��grPj';�&�#I�dMm%~�]�ޜ�Se�xp.)��t�#Ax5*W)� ص�bK}�Pf��RE�磬FD�ݛw�ں:�5�� {%��w�w���sINpms����2�O�b/���/U6�й����5آ����0���A�����(`8�%<b|��Uz�̡_�#ԥ�	��d1/���e�����{Ɯc�bBx�����	��?������N�Xk�ۓ��0
�U*L(eʠ�*,pVB��A���.�����!���&��{��n B�{�iT�T�0�{E�3�a��6���$CX.Z�S�!	�9�!Dy���1^7j�M����~N5��i�j��h���� āܑ�2�5r:�f��لs��R~zPR�)�~�!"_�� m�b�/���ZQ�`�Z�??M��+��.�U�L�2��*8�&�u9��+0:�ـ���;ɡѬ^��-��>w\�i���cR�Q��3���� ��	����̏d�k�U�'�1�h'�&Ȑ�̅���B-����� }[���(y��=[�$ܓY�I_�l� �r-�)3 ��)ݻ8j|������=���DR�ݖp�Dp����~��v�k���$)�o���Q�A�Ϭ�i�Sk�&"��
�wNJG��Pʟ�{���!��p��ѯ�<��dO5�a��(�N4��3h�A����2��:�ι��{�	ӷ��U�K�e��7� K��͋���-�|�l���qN�,g�?l�R�)P�<��PL��{C�p��K#�
a�M_B�7UTB(]qL|ދ��z	�V��5�������P�tV�n���N����g���c"B�fc���꽠�Wgݖ�vJ����6w0��Դ8����q���&��I��8��	�����f
q� ʏ$£�m����0�&���"`Ypw�!�u�Ǘ�*��k(��e�ZDI�������IR�n�����������!�-v��`��M�M���{����4����d.�>?H�%�^9�8iDF����؜�/������"A�-�	c��Q7]�v���2�eAƊ&�y����� 	_�}��܍Ġ����Gj�֑�](����;�����igg_��97�%�����-Z�c���%&2$����΁�V���b�W�p�����d���H�p$l��Ÿ���4}(5���r�%-ݵtT�Qv�j�'�2�?�*$4F�y��%eK+,�Y*���`Y��پ���&.=���c����OP�8CE����0�P[���{)����ź������停H���=i�h��5S$�dIy�=�l�������ۇ+��f�,9�;/���2k�u�=1C2�����V0�ƹ�ZV��K,��>`�o*@v{r��!b8����P"C��a��|��r�:/�ҥp�U���v�8=���%�UpW#���U۟�J������~ׁ���ٷ6n�=N������R�$�����S����b!v�I6 R L墻写ŋJkJ�o�R$.�m0LG!�Ú:�j�|���M��ky��`����ք�$b5�}v�
(�j=A�铞U:Z��(_AN(�ӄ�X�G!�(�m����kV��k�Tw���J�iCl:�Z�,ӧ��թ釦�
�n�c��~rA"���o_WD3�f��[��H��U�V�Jޗ&�U�D��3~�w�"�|	�X��o���2*ܽ]_���D�o@�xF�v"��#�R�6�Sp����Ay.tz���Ϙ���T��������p�a���H|�=Gst�Z̺�)<s�0�-Md�r��\`XOQ��6Md)������$��ɘ��{����j6�eHO�W��3�5���&}7,ڭh�ޙdh�2�9XĦ�F������)>���{W�H6��&Ϣ*P	�3�%����مLB]C[��#��x���~5�&W��}����f�������%3�;�x�H��Jq�Pl���4����|%Q��k6�e��m�!A�"������bJD�n��Q� /��e-�wtCF�N
F��??���2T�S����V9�}�� gr�� 5�%!���H�$f�B�"������V:P>��)ï���*~��ܻG�(������k����z/$ ��R=A��5��l@T�]���#�o�)��C�CF��X1��E�v��xj�q��?�����-Oٛ�	����9��p4�	l݌NjdهT�