��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���cDP�y�2A1y�n��#�e�qI�/��u�e��|��;�󳆷��N�Н�$2.�vy���e0�o��(Z�-�W����cq��4��>v��w �si�)`2�+]����
cx!r4Q-b�&�h����ņ��Շ�:_�frHp����@�a�p_~��p<��Q�,ww@HU�w�<|�(�����T	�'�{ˑ�e�Ε�L��������y��A�ԃ/�%�L8S5)۾��{~�[)�� 	:�#F�A���Uyv�V�]ƅ�p�(w�j�&��714n�x���N��p9a��؍�K�% ��1^ ��hM���؛���-׫�4��"v��DS��
X&�nB�K��YM������s�*�@<��vS�R�����j'�4��;�>v����J��5��;k��ٓ�&S������6.�͓5KI���\�?�V�Ɉ�Ϋ�`�,�G���$8��7��D$'%��u4���&/fBn[��ѡ|n�P�a����
Iu���1�y���>rtB+�#���2����(���+�9ymc�pw�����*�Z�8u!�;gL���5��焒l����������1mp���1v㑅�G��0�05p�r�e��LҦ�_N>�{PrꙡO�B�/@�=�Q��O�~E��ώ}W�� [�nA���O�7tu2r�ig]xH��~K�-b�����<,=Zz
-�UNr|m����Bʝ)�x��k �����	lp�7�e�P������O6�Z/��a.��������z����%�	�!0n�>�k��4�N!}R�� G�j(���ѷo�����qҒߡQ�	ho*nA���� ��7GN*�1U�����Ǖ��V6�����*8& ���y�xT��y/9�"[X^_,�i���lW9�ʏ�����:�����+q]gJI�Z���P��)Rs�eA"[{�ed��^z���h�d�6���OLr��*ǽ��w^�(����Z�a,�u�3J��MngӮ&g`�</䰎�3f:s��W A��ÇO�ǁ�^W;@�ܢ
n��6�6�R��'S��Ʉ���1���;����h�Pg�@��&��QSDʳ\L�e�J�ޚ�S��*64Ed��L��a\q���SWsZ�yb
�G;��������ٯ-m�	��{m�e�J����h�>e�¤�ǞxtPݴC��p�k	+w��s��u���SgjY7�$��.7dN:�C�qs<�T4��+׽�}E�lj{���{޻0J3�lt��>`������/�L\)]0g�����>o�ճ/Z���<T�~� �i_�>������YƁ1�7�?��Y 4�1*}�"��c�/��L텣��䃅�#����Oip��MIP?�I�%�3�JFP-�N�4���{�%�[�ia�}�	 o�\gN���3m2�����rb�� �{y�j���yϔY����kr��?�GD��`�����UI�J���]��)u��qg���X8��Gv�����]��
��7q	!x!xԚ�4�EU!G^�h����*�!��$��LvL�1�^�#���M0��lЗ�s9P��0 �\�2nV�c�zhΊ7 ꏽ���d<��F=�Q��x�ǲ#�����&1v�@��e)�߷WO-�ʮצ��%�v��C�ޏ�C���b�$��U�R+ㆋS���}�LpR��ަ���Ԇn\��=>"4Wg̍���e{��2�d�A�]N-��S�V��˩�[d(���&ldn�/�u�3����@nĆ�ĵ��}NkDg��n4�f��N��&��fwe��F�O�I}z��/��>s��R�{��)�y���0 Zb��a����)��J����|�kɰ���s��Zh�c���d-�0��/����Q��\@k	��I�g��-ԛ�>���7%-���?�C�2Lb�w�Nt�����{�xҬ6bs�����1m��%�I.���D���d�{��]�|�R�A�\f�c�f!2=��W�h��"J��33?J�� �\l��&�1TM{
�ҽ��Y��*�/%��P��n2K%U#C�h�K؝&Fj-��l�?�f!�pؑQ`�4��jq�_U��]�#�m��Q^��Q�F~"(��tF���܀��V,�X�h�)�*v�r��x4����&,��gy��52^rK�G�ʴURM"��=����{�nH�%]�:jH4m�X-W�ADL[P�v[���65zԖ�i����9�$�K�Jg�H��ϕ�i��Tʎ�XT9D�_�4GB�6;|�M6�nc�A�3���¿^M�\A1�;aQ�N��撤�E}Ul3�S�0Rսj�l�uz���!W���_ߧ�&�f�e��Tk�4a�K9�ϼ�d�ퟺ�P��+�I7�6���q�+I̟@F0ј�� ����O�sz&^P�]��B3���h~Uܣe�͆�p�^\L����}	��#�|���O��Ã���Đ��<�7(l6W�����u-���F�(в�ة�&�L�Ypx�sw=��.��pZU@}D"W�l�T���:I6W]T�8)�j;�ò����"��3"���]N�ٟ�w���X���9J�>2l�D�_?��Rv�nkT�����ɢb�s��s:���8�ǆ�tL8�*��<:�m½��GӡT�f/wdn#���q�l	����jz����tV�R I丂��~�_�]�@����#8�)�Ŧ�nJ\�'�
�u����l�AC�Q<�(�=8����x
.����;��������/j�$0�B��u��X���>��C:��A�ا7�'$���\��:����B�B���N`����)<f!���q�Q~�l��S�N_�f�|k{� SY�;��Ъ���Ђ���5Ao6�j���
��]n�K�M5���N�~f�@��:��	��wv�WUb�ߚBHfT�Awe�5�8ve!3r�W�>�/�7|���	&gDn]#V9����Vo1`C��_�D�7���#�ݷ�?��7�����T�$�=�'����}�������O�愱���T���b�]����_����(=E/}��Z�2�,�w�؛S� Qn�#C���V�RA��@�}��MBIM�L���ec_�J��:�v��S�4$�{��X6B�ѧv�&<z��9�;��L`C6�L�C��W��<GMI���c2�u�V�=�OP��'���Kr�3]
pбt�t�Q�j�Qf!<����-�;V�ɀwO��'�טX��ŞQ�5,GJ���&�v�������P�w��NN"�Z���)KvBI�p�-̭~KB1sk&�j�± ��4�V�4�$��=:�T�g�Nk�D�8�+w4�����Lq�RzJ�~au����I��n��s�jU924~cWG�ȇTݜh��TG)	����3�+1��|�צ�QYhde�R�;�iSVi�<.�Sw��u-���ku�� ��4��pf��t+uc�C0��(�C)7�TO�c�������Z1���đHL)��OD4F�'[��H��b(�����`��a�x�5 �=b�„J�����'��]��y����j
]$��B#�
ty�ո�lA�h���-@��G�tJ�x�D�V�I�.1�m�%�Ƹ6�g/� !8m߼.BA�]�wEf�ϟд��S�"�d�{Ҷ@��1��� Cr��U�񥩀��Y|�,���m��@Ų��=�,�R�=]~�+����Cid
���'C6Ĺ>u��]}v�pcZL�Ŀv�1�C��fF$c�a�
:��E菰[v8V����+�ts�C,�~9����w��V��QCUL�ݫǶ��ē��`/6�U�ʒ���K�i@�\O+�T1�z ��;2�߸�
R�rR<� �V�Y6\z��C�^½xr|� ���$(�_4�����;��W���x�离����}�n�-UK��q**����2܉�/���(Ev�W�I��0q��e�D��dX	ƛ�%n 'ǗZv���h�;c���M��t	�yr���*�Zr7��1R��\��LYB������T��F��e��D���!=�N
qp�X�:{k�<�-U(�T2� c�E��r�8����ч��@�]o�%�Gp�/;�����C}��m��F��-�\d�d�h'=���5:��5��^�6�O�Y� �vN�!�u>�](�`=�)Y��>(�����q�(%��_��ݤ�?3!)1WɅ|�[)�}���J��2T�����Z��6T��s��g�I&,�g��N��A�r;v��J��3���a�/V��<0W�&�h������������]�$�
� �RJ|��cH S��>u��E��4T������[�p�Ԙ�x(����C��8�����(���q�����%�6;�����UaO��g[�*�^�25E�j�Y7Ɵ-4K�_1�M��G���x����S���l\���Mi������(������������S���4uO9�M�-�:�y4��=����[���"}.k�Ttq��%�u[�(���į�u��h3�B�\v���[�Y�M����xB��y�m�P�9�pX�!~�Dm33�$���3#(tSVA2�J���E��m�1Ϋ�)	�L[��Ɵ+!7G19?`���9M�x�gDt��H~��詼���9�p�IH�G���ɵ�1Mq��_t��u,X 
�uV����x����s��H��2�	����yL��y|QyUh����9X����pu�^��n0�	q��;�1\+1����!l��h� ��(�C����v���勰�������%��Y��양����L_[��4��×�"���b$��G<�3�a�Asiڢ�
b�Q�<3pw���$C�c/R��A��	�$!�����lOA<`��NU^
(�7�9;x�ˍw�+�#�NL���3)E69iB%GTi��M0�ye��T�Y�z�2��������N)���g�`���%��i�t.�[]YZ��Ԟr581��B��o|J0�˚��_\	���
dn���՞������U��t����W��=X���#�nZ3o��J�w�	��.x��#��1b��+�챍�r8��U��&=v�&^GX�s�NE��6���Xzg�$r%�lI���N��E3B���{���UI�gmBY�F�����H8�a�gh�������QV�RS =y�rGŨ��c�5�?�-��D���C��/��l��N.Ň�H�wk�.����Z�TrA5ts�m1�}��?o����֞�cE�[���3sV��5A"8��!߳���랢
��=>1�<��#�W�4����'UGr2P~�-�¿�?87�]�ӟ���y��Y����3S3ߓ�1�Fuo��X�̛5������>,��6%w��O;\�2|�F=`�� "��ˬp�<*X+���"��-��xG
��Y��̺�d[[�߀��/��~^^�v|�z$f��H>����r����GQ�k�w��>w�R��`V^h� y����3�����!&mP�[�q(�֟7�S���f�?�m��(�n�]�TƱ߸'!i24������*��VO�O��B���3CW �z�(�9#��1�K���3�/�_�F�?x0u� qg�VVu�]��M��Y�����g���a�	��� D]�z��
?�k���PU�<(>a��s*�9M5��l�:"/�o�c��#fꅝE@tYɳ�a;ڨ��@�0ݔ��G�5E)i�D�!�B�x��eYe*�)��c��	uu3���X�/_f�{$wl�7�`O;�R�a����FN�Բ$m5v�Bg&��
�����Ht�%!Z"����%3�1/G3�d�QN��4�Һ����r�����T�N6���&�E%&_$����x��ݒ���=�{�<J��+������\б9���)��������%���{�x�����e����>�;"�JV��:�q�#W�+1S�)M�;�����q�*ئ�mG�д������^��D$���X^i��c��1�bE��(³]L�O!w��Գz�E�x�M�sHk�֊���{�0/O�W]����M��5qqO�����J�v��z����!����8���;�ܶ��
Q��O�VJ\��#w�20�n�Z�X��1��ǥ@����P>-z�6p��	PbV�V�߳���JX�Y�� �_�Ȑu�_���"?�%�p*�R-��L ˢ�t7��������������lM�:7�r�<��r�B�5�g���,
��T��X��W�� ���Z>���n���u��p)Got� ��$}�v�K|��%U����u$�$���ʭeԹY�[��l���!i�FB!�湮�:H�6��n}���|��u��W��{���;M��^n���w�	�+��g`H�{{ĸ�Xgo�h�l�%4r!���KP-�v������f��'�(?|���!Qh��VƂ�8������4�"�����bg���wěc�d��>&`OC�se�o�}��3���������U�>�X<>.�����f�[�_zJ��׿�����I��A9ޥ7�U�����Oc���D,���8���	�H����P����{�6`��N�¥>ϧk)<B�S���-�-�
��sYP�̧��1C��Me�Q��q�Y!�l�������QV
��8�o�) t7|����D�ʄ0{��Ũ�W�ڑ�ʳ���u���n,�9@��;(⋤o����
�ijtD@Ҙ��),ڒ�����v��sF>v$��n-��e���Q���u��i�'����1�t�p��Qu���'�C�/�?���4t���26=�d� �W�REDy���D������3�*�<��^=��#ڷ�D+|d�mn��Q���X��p	w�m�g����IZ6��	�ɜ&d<ȋ�eO%H,�l�I�Z��0:�׈��R�V0�򶶠�N����+��P���w�K�dͦ{����a4O�p�����*����+���/5U���=�
�����(�uJ�c��77�'��f<):3�X��ɻ@�ba^�P�r�X��o��� �����d�r.���}"�VC����B�5�����Y��^�bx�.a���u��ق������L׈�x�?� ȇI	W���؉UF���*
"��}&f�ϨM�x�(� *O�2�Y�@���q���BT����#Z��Q0�3ls�'S��y��0'܈E�
s�P�܃��\`�l��A��o��#u��B� �uހ�τ��|iI��6v����/۳�\"'��]��a5����OS����>@5]��NMl?:���U�]�_�/O>:>�?�7 yT�C�4�*��T���k�'N8&Tc̡2{^�	봾G�y�ߤmж*�i��0�r-��b�'�i��&ό��O��~�8�z�w�.��/����j(Rk���� ��v��n���la�P�
����#�Ha���4� ��$��f�1��P��P1J��щM|�@�\wp1��}�S&�UT��5��$u�o�/�=Ԡ�l�KY7UU��U�r���] T8jZ��r�UT6����������Yi�ݝx�L����}�]Kl��^�TX�r;��5�J�ZW==h3`H�ۢT�2s�1��:*
�Â�jw���(�3;W�Q�'M�^�<bg�T�A��u��R���p��g������99��sȃ}�"��o9��[�d�j�@�л7�5���vJF��_�h�+H�?2z�ac����i�