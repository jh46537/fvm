��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C��_�+��+��^���vZ�r�Ln�ҤpVCQ>د	Y��U����M&K�E�N�F{��Tx�H�|Ic��=ƍ<$���C�q�HD����9Nc��ǵ��7��������t��EsK�L�ɏ��������=L
w��?�A�;�m��V����]�u<�vg��I��E�^����9���A�7��{A����ssWR	��9���t�t��	)�nZ�ǮA��#�V��Z�{�g+Ӄ��>z�O�p�����aV��(��Ԩ��X� %���,<�q��DF��T@���`����S(Y�D�/e�� � EH���2s
0^�8i:��F*F@�M}*mN41sv@R����cN��[Bq��d�PF�A�ÿ!���w���=w
"䇦�p��_�i�>��������6Ո����/DK��#S>�uu����ٙ�0��
 ��;'���V��w��5#y�*vR�Ɉ����ىl�h�
����N�K;���H�B���[md�Mc��w�N�yrY/��4Y{S��k��Sb[��d.XAɟ�M�@uբC�a�P�h'g�#(7t��4�A�mԬ��-p)�g��7����I&��N�$�A �>�u(l�����C��U{�t�C���m2�A�>�Õ �_D��x3�T�����T�����ay�o� �������`�\�db������ϛ��o��ڴr򓬰I�;���\��6W�Z����y�h(ʍ0G���q�^��plI0�O�R�[>��s�L�g�g��u�T� �=7ׂee-a0�Vܺ�0ų�JN�Ƭ�~��&�A�}B?l�^X`�|ח b,�(�w��R���v��m�"��t=K��D�4v?��i�c�ӫ܆Z)j���� ���I� ǧH�RJ�@����5d�m$����������i���H���rII�
5~��
�燋�H��B�U	ѡ�{F�B�IHO:/�T{RE���8�����B(�؛Q���x��rN%���:�$��0�����mtG�x^�����t]������e0Ò��#�,���"1�1Rո��lK�d�uX��#p���e*M	4���������^�Sϝ'7K��/����fA���W�d����<��q�E�2�N����[s���w�i8.�-lw���_���
+۲7��׵��1.P�����p���&�6N���b��f��4���.�;�S�z/�+~�]��!#�������>j�J
|b��/<���"��<�/��LD4�%�O$Kb�=�f=c���8{���<Z�|8��h�w��h���"_q~�Jr!�.n�jP�T-��n��Y�u���,DWƑ��i²>UJW�L�z�2*�>��F�t����ҭ��+�=[�<�1ΐ$v��뭟����������Ԝ��<9&OmS$�	q۱�y�ex/�
q�R3I3# ��FJwE��� ����s���)志W<���o�T���.�*3��[Yv���`͏���;B'��#����h�`ݪQ%�~�Ĺ�ր�OW�`O��$�%��J�@�b��Yu���	���)ɨ���6y��3eQ�� F�����A�k�u�rWe��ga��+�v��Q���+��Z���;�k�H��|��WӇ���!�Cǹ��#�D�rD�Mxp)kT'r�4-6�3�Y�:��w��,�b���:;���,�n�a�����5v͉��>t�.��hDW�XЬF�N'������J��o���w$�]��!����>�Z�>[���MHEY���u	��w���Ql6`�0��I2b΃7>g�v�Ճ�b!��H��9.�N�?�\�W�
�����xJ���KX� ���j����qЋ"rf����ss̢o�D�&yn\�t�l�	�	ݥ?����y3���=�,���(��d����]9���#$b?5b�W����@%�Ȏ�<y��y���N�t��Nb2��a"�F�6���R��<;�eOn��+������r�MI�5څ�	"�=&����Oǥ���9Ll(��5n�噌A���W�+C��<2 ���xn]�BL �ǲv��R}�]e�<>0D$::������5
���ic�hj�����5��&6��Ɠ�|�n����p`�U2qڬ���b��}9C2�/��m��r��p`��E:�i��������k����PQ@��(�V�~k�.^��=Z�<Q�	n�{��'�,�~��p�#�fR��GeP���ߓ�q�]�5a�դ��lwb�I��vhR�X��n�.R��A}/�*�&�=ԡc�rE
*Z78�����Q�?�P^� q݌�kY&�D�:\ڠ��pP��B8�u{c�C�]Vi�Wq_cc]9����ו���0葭e�n7���S����kގ��jl��
|���Ȥ��^��k9ԅN����%:2�S_w��r�9V��;����Ln���J��=�q5�3���2C�L ��Ĕ���Q	����n���r�䞓_�p	���|���`b0�L��Ɖ�mj��Av�(o��AW����(	�����/��Ԃ�2 ��+������a�!o�ڕ��&w�L�m�ud>�k�/�6θ����u�b|��q�E��j��4�U#��}���4��%��+ ��1D�T�#���t�ֲ)O\��-i��;��X_rx��(��qD�k�s�.?.{������zk�gS�����H9BP���h��:��R��*0�KF��*^��*q&�E�Rͯ��,]��~�-@{B~�"��)��r �߆P�E�"��L��H��k�b��iZdy�6J�G�L����]��R��y�af�y-%A� Jv��9ji:��kv��N;K�h�Qu��W�r��2��"0؄�`"u
�?Ik�N�<���cv"���h�墥mnQ%9O[U�&��6�q���Ir��8=�����i�}=[(G�	�iU.j�E�x�s�w���'���м~��S%Q����
�8�Z"^��VbK~fvhc���4ZP��i��ې�f�Ia��y���~x)l�����[;`����Y����KZ����Uj:���ð亥O��/�rڬF)�2P���bK�����,�9�ĸ�Cf�擔��J��������Ǹ���ZG�2��2�S��7V�óM�c��.$�uC}A�.�W���:����~�
(�Z��̢�2&��;��f�*�-�mo!��<�h��NjE,������c�r����
��=j��_N`��\o�YP�f�*׎�~�5ݓ�rv���L�&�G�U�ѡV
�f��󥏶P��wE��M��̷o���A3%���O��3:���E�DFH��TGMf��p�J��`��C�o�}&F3��|�����nf��^�	Lǯ�	L�W�l�Ғ&��#������mr�L�RQ���Q�Fg󌘻MTP��L��q���?3�����d�rk���)���Hv���N_#Z���u�a:��t�-k�G4\5>��y���Ï�ʰ/^�T@��6'�

@�|,s�����P��������$n|5�:�6�u�bV7K�5�H2�1&}և�D�Ft�Q�ò�Z���0Ś��I�J(�m�Nڷ1�K��D�����(5ؕG:rV�c�
����K�r�9h����	�$�1xedOd����̱�ٿՎ&O�|&�%C��ju���[�e��L�	g�;�����?��ߑ�r��T�7/95�jMBBG�$*���w�@�2����=�����ic�V�c��	�����v��&Љ��n��1�A�����4�M��˕��� �����FU��}Q[�;�?�^��^s���a�jjY� �^��܎������� ~&;�Ԩh�0S}?��gr���Kwd�s@�>����+����2��s�Ъ�!+����?�Cc��ڞ&(4fl0��=e"���k�N�m������A�\�!��i�q���˓K�M�%8JI@	���7�Z]1C���HW�V��0��S��E�>9ǡ˷�)*ҒDz�W�Ȩ�C��x=5�����?���D�m�JH7e���uo��6+a�+v/��aF�3��!bi)&G	��ߍ�')��Ɏ�F��aS��.u�:�����������hEQ��ݸm�sϲij�d�]Q��n?]OeD�J60=d���SxSl��_���X|�*�.�\��d�������.S�gB����ea��郏�z���.�48�oSh{��هlP�3��:��I�U.���>����L�@]��t�JX=n]�Y�{.�\��th��P �۫����#EE��,�����?�R��5-�ɔm�
,F��ev���C;�HS���������
���K��/�%nq�mi�������y�_���vLm
�l8B_Z��	b�Ā"��w:��^F�үU���=B\	��н �'�c�CE3�kE$� �B����!+ZG��@[�M�v�HgO�S�b����La���7)6��#��īE44'J@>�Op������D@H��K�߇��D\�6B�Nr1�%�cȟ�VU��܎�XK��w��Q�jr�1����^��0��ì�o�B/c]+3�-o���������7���p�b�
�^�L���e/�X�6��Vd�33��A��(H�� �0�éw���"ڨi����}�-Z��Ze�l�-��Z��w�)�G����,B�~r�j�5{����l]��H����S��K�W�IƂ$��W��z�8��\kV�H	B�J-���_���>7�}*������?3T�	!��:������7��Q�ӝ�1:��o�-r&�΀ v�h�Wo����:i/,���'}�F��훕��ݯ�dÆ�ۣ�\4��2T���x&5 @A�=��t)ӍT�m��mr�|� q��[6G���bc�ޱc��ѣ��#{@��S1�Y����$u6am�
���G\I�>���G�b�a���	H��h����bt/��qմkb�!JC�� �1��|,�������-�=�ͤ���W�~N�b�Q~>��]tǻ8Kt����$�_��	��Y�{Zw����'�{�I�(��|+��*r�J��I��y���u#Ogdx��9R۟�bh�%����K,����}{hr�sv�(i��}�9*`���%��_eӟ�4�w���d�5=�Y�E��J#�߆�2E�t�:��yT�e#��~5mp���h�-"�w�]�i���f�]��@������YI���c���G�[�e�kȪ$|S�K�ZkV�1^r���͗o6�o�#J�2)j>&��e4k)u[Zh��g=VyL�M�����N���ȴ���	"^:�3��(�2I�YF*֩'�B}�}*�C'��ER�͡@dK}�2��p��s�z,\��i�PZ��n�}��G`�q�z#�mAĎ����3�����q"��a,�ӛ&l��?�����>z`w��O�*=�uƲr"5ۮ� �"l��gv�o^� @�+5gL�e�э�@߰I՚��$�I��r���\��Ke�̥�v���b����orXs>D~�Y%��:�L���?)#��z75�J$���DUp�R@�
h`���4�[�EC&��J���'߲b�B�~#it�5���1�A��/��ו��q9v���ep���0y��@��yD��.9U����:��)���Q�rw��d$)Z���{ �@�3�=	��Fc��p͏�� "v�!�(���-O�x*5*��X؄���!# �v�S��X��:�I��Yu-�Hb����e�z8�����g�S��'$���=պQ���� |�n���~���R�,ٱ|�7�!F��m�,�/�(?'vr�HT!��n5��S�2` V������~�������
�g��U>�)�X�u�*�DT�t������uU�G!q���Y�+�˭��q|K���z����h�����j\�y�ޣK:��v�o��	���P��.����wN.T,�4�/�M�����R�=�T���XVE��7i[IU�x?U�q� �q��!̼�$�u�Z2(&�k���%İ�Jč��y@�±
U˃�Lp+#�jZ���](.��E���=�[��HR)���!,�ώb!�~m���FֶvBc���7B���"C^�DA�
i����ժw��J34�����!NL1�s�#�Ip?q�EX�3�N��zB�Px�r���/���l���v�e���b\�h��7���e'�������b�������c��m8�r��
6�"ݵld��bxu�SCe�����yӷH��[U<��ɍm7�𰸽��UXsk�?>^�5E��;�l��TY�-cGdȸ�[w\9%�]��b�w)t�e��=�yɝ:F;>;X�V�����ctA�� ���ŤVQ��xr����&��s~"�f @m�t�?�>�ʱ�P�߫���u���̅aذj͸�C�:!���ّFG/“�>!�pzҴv��9��O
if��!o�`���Nm$��QU���Na��H����d�@>5Z�%Ѫ�گ��A�qnz�V �����r>C�P��'\�(
>�.��*d��z�5Й��4d�7l��g۸�5��N�ْ���f�u5���N�0�O�Pb?l���"�G���ک��T�K�֣�nO���@a��N�R�u�8���l6T���A���f�n^�m2�Q,1dg�00���5�ԫ$��W>�=B
/�9x�ZL��G�%j�1j���_,�Xɣj.��Z�W]/c�Gܳ�IN�xqk�Cۉ�r�<��^�T�!�6�\����W�|�ѥ�y��u���F���܆F�[�*�Pf�ɽ����O�8�5��c�h��|<�9��na}^Wgȱk~8�q����!�s�G���`H�3�л��Ԏm�-���̾rċ����K���Mv��.6- ��e���,3�l�����!�&a��p$g�{�3W��(��{#b���찠�e�pl��Fsa݂b\T�oԠ��yW+�ZrP�S��Q��!�qf[W��W��-L�3n
x���(�5�N%v�v�U�$����EH�L\}�Y/>�d����r_:Nw����h����j��'D%�{�Sl���������ME#'#M�%�{@�JЎ�U@Q�%�G����*B��<N�(�GNS:�^%�tB���e���CY����ji��k�^���� ����o�'�E/%qA2�(��"wi�ǧ��Kk	�&��Ӌ�%�eϗ z� �������E�k�y-EP���p�RQ��#LY��:u�6�`0`�b�Xn߾@}ʟ�`�7����/��p>=6��1:�� ��%}�?óG'&�FK�*�Nhˋ�d�apq��z�y��b���F�_�</�(>]��@��L� B�&�{mcy������5H�`�~�ɂF��L$�Ok���o���<�����*��MQQ��Z���V.�1�@X�^��d0������4�Ɣ�o�W'&���-{pf�8����Ɇ���������y��uCE� R |4���������@�?|����CѦ�2��j���+
��6&�2!m���'��������&,�k��c�,�
��YB3Z�5E�����p��?�`��	�(��vِ0�&���z������&�~Dc!z�y�%�
]_=��J+�;��5��;J�{�$].Y*B1ts�2
�|p��D�$7����/�o�{�|h�،�m��
�Q�b��N�w�9K�1��.g��M��$�4��ޑ�u_�f���J���d����0�QwP��n+R#w�"ב��C�l�5�(�R�<o��v���-�69��7�h/�@��0���6�&�����	<c��>)AD�bYn���V��Jlm
e����O���&�ʝd�0����5��D��۩��#� �mE�����A�Gtu��fL2�=�'��?�`�N�#(���Ikg��`���{���mzv��x������e�SH�$�6�Y��(�0K�%�k�DʟH1�S���� �/Y�cf<�(./�����! �/���ny"�$��U��?X���o��q0䨔 ))詛{��KZ�E�E��I��"�⪵�(Qھ��b �m1�I��s<؜g_�T�r����{�B|�λ��C�A��[��NFL�O��!j��x�$���kT4&�^��p}�ņ!X�"�P&��8��_��Af���f`��ͧʅE������N������J�e�	��^X�W��g�� ��+��Q~����u4fY�p���u|t�Kj�������:��FH��]A���
*41&z�ӽ���h�x�\M*�R��h�<(/@��8�O������ݗVNO�J�M:��5(:L�g�H��7��\?���;�4Eg8�Wpb)��	\��m�<Ӌ��������{�1�C���A+�y��;,��;���z�ЄU�_{)@78��A����4��
��1K:�}S)CM�A~h���:ߝ[0���g�?�zf�:鄀K���&�~� �)��`��@�e�,�;i$H�\����K��7�6@�>I�ް~M�B� ��{d��YG�'�w��~W�F3X.����i
��n�#�_�ѥ�@>�� N����j�1�f1���ʱ��򃀛
�P�阏Z���A��cu��HF�gBB�m���HГ��R�b�L(��(ƨ0O�1��E�F�(��_q���P�� %�%5����T������⢛����J���|��ګ|C$(�]�%P�^7�=�#|��2�-�� �ٲ��m�h���ꌩ��6`��B1*����ϊ�R�/�*d�*,+Т�X�Z�Ӎ9iSudr�I���P�<��kc16��3=�ɶ��}�k��5Jւk����'���0���3�y�Ť�-��/y�%����}��ҁ���d+�Jb#5�;qѯW;w3�?ܸ)m50oR�����^-(� ��o����YcQ��VT!�M�>w��<؊G�Bj#���s�%F�� rr��Vk\�N�*8�?L�E�lT�:Bu�tX�
�̟ӈ1Ni��^����5�o��K>I
[
��!�x-]?�f����TƘm��s{Q���0�tu��M[���	���;����|����
N�,e*���z��alm�ޓ74�\q�~XX'���a����)O��	����f��>n�p�_�yZ(CC���y��	��t���'E��2���T��ȑ2�����I��=��^�<���J|�?��X�|q�5��P|5{H�4�Kn��I�=���KT��s��{W.�_��:��q�
�n$Plw�A(o�0_��K��j�^%��f�ٸz�PU4�^t��`��d��:���\}W�G�-�IG���2h�A��i݊�������ߗ�����P�l��T�S�8-rH�T��9���K'���)ˆ۾xaq֬�|z��,�����FQMS�:�	n[������ؑG�Q̫{�������+$_߀d|����ர���[
�Rb�����o����	�w��C�1BZ��t��9�c���`_E������i��A;�<X�%�O5��@d�w7���$Nd�MR�	dZ�L�i~q=Kc#9������Wv�[���/�
G�F�U<��җx��E�䝳�'ϱ���',��~T���|
�R�lc���!����bo�Ѧ��*kDB��$&�q
t�f�2@