// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:22 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZWmv/OrGGgU7vDW3JPGaJl7gUBbS/xyjnd2R3EjzLAen7PMt1r8XQnzVR+89fcUr
1M+S7asyqNIxviXj1wNTaTxpY1lmKTYl0tIpf8NI5i4TUOghwnR+oDgc04tMKE3Q
oi7sE9v4W1oBJ1OenH8eR27pToe+lQEkwaoI/8n7WKw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6672)
uNQsfomD9zNgtBk/097hjbufFCDGHaxYgHyHOJLmXlc5fh+EBaRLXU1VFCGnuGgT
GsLWOwJgZOmx0sRjYODh1escFIm+4a9qA6t1QT6e7M0fUQOA2cWWwaOIbANN5qiH
fPFRUj1y1VeAhtBuwM8WgSwY2n7sCPl2fk8UFITZ9q2X6wcaH60//Pw0aLfMM/kd
S4ll4pwTg91ooKCehBZrySeJbq0N2tfQo0lk/1lwZvfRtjYoEE3LfNPPMVYVSwD3
QDAsIsGuV8bpaocicgr1GGL5vAbhZUL96Anz4byo/8vtY5/CmQi62zRoBzhuHqV8
3jJy/1EHzXJMsWP6uKqYXkO6fsTRjOY0ne96CeIN8QBLUAiLNOtrmJfQ+Khf1AyO
7SstGfW82917AvN5dyHwW7yS2z0uqdgx/NEESjq214+zkXzzphxmhO13F+gvOmWg
6QPXXKs09CPLt3fupzVtR/sJbS5DaBOvmqNWCD3uAIXV/+PolihYzhCHZt/qfF92
56xdCUf5tMj16VX85CMJyzqHHKi2ZOAyupTYI37un/NH7V97B2gRxfSnIKueikFW
A1Hjy8LZrxm48xg87iKr6jbBatAMs3iVsZLD+Em5FgxVwSwEBpyz8UXeAidEXPE4
52ghyw/FnI37Fom59uq1iB363D5Ki4yz2O8Y+lySpiYorW1dLQlNACcvDy+V0GqM
qvyRptA9zzQg3993FVzgm8aMaybGhzE4f3tyENVx4FlWJU1XqvEuuOUdv6K8006I
qElQyFCNQ88zySf2BApa+DXrpeiRGb+bM0HrQCCW9i1JnWA0yeSLHML8BuO7SjJF
0QV+gjRltDyDPlffIDXvuH3dkWtAevQ6lKIZXjRF7K2JgWDkyrkHnhSD02gcDfRX
H6AlcihmnSo8UBvH/VcHjCaTnL+ScNZyIosyk953HCAl1wV9b2naXHjU0CbZjmy2
j6w3tlo1B11hr42Ntn+YxK57YIXW2l2iRBXgZ0q6Gn8z1oPJOd7X5fkwrWm+HvHZ
x75XfFRh9sOrLffGPbN075eH2z6eTN0hYrmFInNuW3PUVZso4aqVRy1EHcE424OX
1+bCQtW5+rkD0r45rm6nBx5D1c7biAlToophp6lBvFgQjyWxoUPkmWwSzeHC6C4K
59EdMDv2wDUrR7h/2rwL8lk2GLF9w5OagzNKq6ALuyn2xNcpbpbnFNepTyPStHLR
ZpK1LbbS7cpq4IXyBu9+1fyNWozsIg0HiNoinAVx5o92YXPC/5sEA/nqh6BKJLw6
LallLnYykN8d7eP4TchN8bVGY3+7TceRV4edf9DA8ngrWvz4RTMS4+TZjKasYQ26
2lt6xbEVRHbLldUeirBzs7JVvHVc7eqHkSt9FL21s52oBQF62aYhyiLVCLvsfA3t
LJu3+l9Eg/krafQUgfiVJBIYVOse3Vp6hNftM9aCFZ2h0cynomf0RQZeCbI3oFQv
2bTzWrRUHj+h7uewwykAXBiMV5GJ8x2o1DZBP3Um2pn+50iD2MSDAeEf4pV6Vlxy
LX4MD+JNm69CUKgQnU5zXAecFxVDaf/+r/8dL0Rux0l4FYM+2Kx2agK29YWiSa2D
Tpl4AJ7HHgPfQN05V53frcFt+RZHGylgx+cAjB/BYtpQ+MnISWDbuyIeZRji0fgJ
N/u2sLcdqAngwKmejzjOF0POR9PxyTFD0uXKowRrcZE1aDzPysWoR60cS2uE1Qt+
bZp7Hn0IrCWvdhtA5qPZOqtyWtCQOCkBZNJ4+Tug3oFqhya0UhQ5QmNl36o36fK2
a5d++X7cJVMXMSBMuuyo75PWcVfg/osT7WSchaKiW7vhMXgLQ90KSzoKFmV3xfya
uZz8XwjiZbeCg1zWJPQx+5Sdbx/50nSRRl2a0/K+4rHD8AblsQdeAKMTF+TdtjsA
ajPXiC853pggBVql/3Nh/+Jy6eCIFL+M8swYl2/3zv6BgT2Mhwb32fJBnoxxicOc
qhGRapSYSmQVNuJ9AuvfOqy8R8TbnOtZwUJDmalV+0hsSmqreRNJHMRmgeJdGBPf
P/sx0nQXKNgqdwg5GChAHP+B+WmXCdmajlcij6kEjI8YL0MRYiZiJm9YwwE7Z9OW
ZH3wR6L001x2hRszAh3HMNHfFwhqsbXbBdG9gI/bJ6iIBSkQhzWWrhQMYuBg1KYi
lN8vHXWofb90IJEJ3nli9whNYsvgACeK7xK0USJL0W+7+W5xftUwjJg5aFKKHOEE
TfJTVXOk442a/C3AgvD9Ea1cF4xIqCDmxXPnrm2/j7z8spchAETXNpOKW9YpX4xi
PsSf5wQZLqXDcPCYDNtXb9fsnNx9yz10AhDjxgoZLuh1Ypmn2oo5X9stiLIKih7s
TzjJle5ypvXtBllt4OMfVUqXPb2Pif3XfAIoe//o+roIFJcP1xXVLWG9Q0noL3kj
E7wz4hfQYFpfA4mCo5eP6j+V8UbDaNuI3sWKKqnLjLfG0XGrVnR55Jg1YdBc5HW0
tDr5vCxps0ye0lWBfd3fnsALXj5oYwa48nHJrGi9ucnObtjnykr4F9xISLrpI6db
mzBswGtpKsI6Y/fV4quigmHiTj6rbFfgsV3vy73EwxlvT8Sr2Lli/10wDsk8w2a6
1IxsAE17mlMXf0BcbndgDVcKd6o1tqH6ffOQ9iyaEs3SfsoNEytEOc8nkvnM5vRz
WiM+OzloGNqvx1U8eN2mrtULudhnz3c4Lt+DxULkCCUkZZOFOY3HR1FDccGV25VY
QBjBVSW3Z2VB9nQfCGURkhz19metek9NadBgDo1eWAhL5NGMuFuFhOZrbI7getur
s77pG6cgohUbgB289/NI9nUqsvSgJZ8aZS2Vd7GUVOomAulEsTZBQNszL1wgKS11
p4BBFT9op+VX1e5mTQE4DBmPYi878UniZaLRL+nY+/yE1G6u3LYBnjjHbWBbaSgR
uLX0B8uH2YL6iJLoaajpkEWfPq9WutTkEVi0JTxfbe1ZZlBn6dNm9cH8GyiMEG/r
lHtWU7HytfmfeblC9xDpnuWXEU+UslaCKTG2JFYpsFvsds5Nr7HGYTeHD/3LEMt+
VmZ7/F947qAAqWAu1+UD+e5VhzzFvcYSbF/y3Mrte0gZ1L/mKvX+1Dlr+2YxxVOX
qCqPRRLOp+Wi3ZuallkX+jrOTEe+JvqM3shlc/n6Ch/rUhm870zNpR10LzM34HxW
mrKA4/0Tqd+5ZWYQNpGzeJ+0fXx3n1ijM+DUZXEaFcvXRnWoy4Rl+By99hfMQIfO
5i6RavMM3AmvYoZFlrGHK+sbKy7h21ugnOY+K5CLWFFxlrkDfIEc1AeNgdWYXlqQ
Wcxm8BhNXSXNtWBfu7aGOsz6wBijUSw8TUeycWk+7e1p0qr4oTFZgZK54MI3Wthl
gzcwPeuu8is1JeMKUfIx3yk+9G7SYwQVoh0rdr5JyECLMcRSJYMVzeAMUa5l05cK
Zj8DxoZQyPbJVDwL8IRkRbKlSSBfJa7TF/2TPBpdZb9ZVpuy/Qwar48HtJvBqbrm
JsWqMSVYjbQAXIVg3YcSRkDUbU/M5AlMTQ5/ZWRN863nDJ4QZnLbKJe2sFWUNl2y
9z8lFFxMM1uem42DS2Bd2TPH+KL3FUCAnJvwkx+SENHxFc3rr/cYAbdFejPw8lF4
aQt7jFOtN2sY/LEeo4845jLftbxWQbKu/AumQbwA2ADet3r1q0dqEptUx/Bbx3pZ
ni62zYXbqsB7SZjUtoiEdijhG9fujW2TjPjfX5/hO5HKQsZDk8b6FDJugpUMHDRz
Pb5TF5vKvm1wywu30QXRdLiK0VcZ8Xu/tSAbNTKrCr5tfp0CUQHpfow4LHiLhCJq
NxO3ianW0RvqzaEJ9F3w3zKD8dkUUgisbS56R8JVHrlOVVWsxhlY9g+OaLJIdNvt
y39ZSnuTYI2PA+KCXyiIVJDyOavaUt5+g7c3P8umo6xZIyjZm+NnQDk2q0Y8x6aI
2swzb84SoHQ8hlHw1wnT/5MWk8uAwXyCZknkbvkfeyrUCFvoJqmJ3v2W4hoHBekq
Ai7OE2yryuISLjoMLR7sZVMt6BxmLRNj2ZatKa+L3V8aigHVJcHg1qjh+HtbVRph
2m2h3ppuPEJf7GJCwAqvOpivHm4hPXJMCDvfWzHs5L+wBYxd5KcwR8dM/AJb2SVS
hlC1W6vUMmOS0KstEXUWHgH2ZkGPs6Hdq8gF1oR5vYwZr4DvvQSAGFH1rRGYjr2Z
IymIbvxtquPRJuS3+Wo+9h2i8bxRNeVsUgdPLdjjv3jqN2YMHY2ulFXTNEIy8925
X4F0K1Bz46WT3GrVlXLF+AXgTel6IGfh5I2dcDN03hLiR03jLmrHE53UvI+DuLbA
0OVshKdLmg16jDQMVfuLL2UZRU8gzPOBYvx8o1zeIidBt7PKsN9PSyyIqXMBQ6U6
8/nt9B964eTfwvS0kCp4xfE/ZBWmNtmcfScVP45h2VOk+EnnPweRTZvv03IQgElT
uJuvOfYLax29XthMRpog9/YWzRTWHs+PW0eSdX6wlKB0FpB6rmNl0E2rGbr9K2Ci
acZUsRBwHCS28Qp11OgfCIcVMLDCK7aw7KCFUoT5nMHREFKs/annsIvDcK7xLa5J
vypvkBeWMirykKxc1FImDRMLNbsDa40Ewe9vlN8r/FsrA+O+K5XL6LODFPlnHVyZ
/9WW+21z2ikvP5JmvIHnQ8weVwrp9x4PjcLMD/QwNbVM3Eu4SGUz9njyBG3WsVIO
J1Cox/Ell4ZEh3S9GsgUE+nDL735ob+wAeBruDZBRaqCknrW4zMPCwZOVAPJ3a6V
7jPNaefq1kgjeO6skOnX8paL2a9Cg4mONULXoFeEhRTWJ4lL/hJXLvdznRGAMv0E
+Qp8S0DIlm6k3E7xCdXVhND+m6nqTquY3xrJmVv8jgf9uyFuYne2IE9BFWfG8G5e
QnL0dITPoKNmS5deFSScCJrnjFUWh5B9AaxLNEIDKOGdocGiP9x67hi+jx9J5xS1
IMNtzgjRNBuAIV6sxJMGfHTEZ6bAMLjRD202jsuvCYSI3MuQ8L/rUfyvy7IDgsa3
hylRc3y2SfZIOqJK73kXGyoMLGZJf3b6ttJwULrhju2H/eD7OjTbTXH6AEpBWKDF
+4rQu7osc/4DiYrlUiPAPyoREp+y9+Hm2QvEekOhC1nZeKqhsMY7DOdimKI1TSub
Ah71/a4tkRC86Gl+4gsd50v8FjaE8uihz3wNP3hsMNqUnM/T8mDfD820SaTTJbaV
PDFM+/SJOO3aOawtxCrZV+asq7aMDy70S9PfMkc+TLbmTZj7BiqtfQjb3fkZacxI
dQoIOadBWu4fhvNGQZf/YUDJRSK+eNhxrHFNXWbXMHBnlnKtwErFNho7JwDCIo6T
NI4cOe/UzrS+N45SYqdGIpydXNbmLTWOckSiRqQi3fMePJvF4IqOEeqHNkz4iA+y
A5xItaIpW2qWBCBBqGyxqNU/gQx/LHhgg9AjxbLPnShGEJVGl7zueyDRt2ncFubO
rrZBzgTbwt24J9AcDEHO0NoivZPDsPzdjI3Pi2LlNsEyoW1T7AODUGY+RKGQgOzG
5Pz4nSSgs9pnRVWpeOBVRCmtCd0xsVYlpZTC+21WRrTMnDg1Sg1CF64M2GeTLDsg
+oxNaWHCiqCpRWHgeMd0qvrQkm0IV9mfdMbkgS7RQQ2NVbUzZKdJAOtP2bhDtMOd
6HXEPCNZ5ccS6bscUq+WzlXub0Y9X7YCTEr3aXPCKXPYXE5yVi9Wg7xuiXCaX+ek
Px5J2IjLHckrmVFt8hd5wMWu5kUnrHjs94M0u5hU6V5fbG+LmxDbQSK9Tc5fXK4w
73JlPk81YdYsEwY/M3oziDo1eakHk75tPiVuyy1AoWzOpHvIocJoUOtgB22cNpTR
1Rsr9u9pXCE+bOWoUD11ajDkfXNTpKNm1wwx3/UKMcN+XCRavIHVBUPqiv833kHf
+vsjqlU2QAKEnGKOY5y623GQg1YFJWry267tTlF6YOx34Tln8Y7YRiGkTkPcaUgL
nBJmnx2bNliWdwcLmnULkA82no6A2Hh+4zD28fYBrMul3mKge8rYh+2EMO+jWc+F
/+wKFEW+HRzOkBujjnquXhDACrOaaDqg7S5jfDKwGF32OCEgJUWYdBmEMPdl/VkF
YOecBQO7QrLbLl91CyZlI3fGQemMWx9mMePCPaMNAfs9+TYjyllEw8OgEzEvZcP9
K5Ot5WB2OS8CimzkdGbqw3cMp47VY4FLwyHBszeiRcunxRirZoUj+/19N8H/fd1g
ewPcLT31yKWCuH4qfVOhvKOqXyXWRK1jzjkUbwt0VMo5SrMCDPoIcamMxyD98wKa
7EEhhPo8LRwX0v227diJk0thsTJnzZxBRRz5KRJu6DWVcBxErQFQPVJhlWxc6YTY
SZ9NCfmMcZmOprJSTkC9zFcolqFgxJaD/F71P+sETN7e4qNCsGYlJGDbe4//33Hb
/TSgld8GrOwME0PF4cPmt9do8gfULgEJVRvcyiMWN23ZzRmEYz1O3+BuG5H/YYoQ
sNV4KHVOZqtPW8ckBBc3WoYyRcgSNvntKb0Kj/oo0YT81LZaFAYqAzSN09xXjvI4
a/ArL5dW2JDnRBwGQ06djrAhn6gOw269Q1XXQts3Ht7BPIdUnzJVpoj7RNVlYefv
fpjzLWObglQJTm1G7NjYB5sPwMFElKBgOJJtiFGHuDelf1hZmYCiERHP3w6s5rbW
aVl4AnBSyHm4apr9apEOWrJFVOg1ejIrDjMrtUDPbhMxnjpYjNBL+qSpnAKAbDiE
rxRSvGaLi9X1advv7O3GiayCwwP6z2TCWOEWKrRC7NJzXsACpWKu0EovQDt7eoHx
WByHkZAacM/6rqrGAKLS42E/H3SA6zUoEZoL7tnvzM0ybguvHO3N68RLsWmikfAW
G4SP7qqgJ4nJGeLGu2z2ujrMhhSJpuXWA+c9iqAbJAWSrmpWhRYHIJmcyV2iO6q4
BambK7g7ntknBx5h/8kVIyUD0nZ+FmK4tyIh9gFGVJfzOsjX/jBGxrVrfy27/gzE
0y67PJqLySrmU8X5B85JGbrWj+s5ePHeyWBra3wv991D+PQOCmCk8UGRH4ER4Ccb
R06h1j2H0PRLSLJakO/dgA1PTTBpiJbGLiIGEM6q+l5kpODkgqWRSQ8gdw31VXUe
vRpWXOjZWkMDthifdHxYiGawIP+eVltGrNYoqadvL8MpaUgYkSBN52kME7Q9o20G
poKMGwT+tTT4QBIZ3eoGPj3GF2WU60gIlggGV7wf/QUdPOO2+AQXuJB1jnj3aIse
U9W/uiFNpt4I1aG+j5Y6E8B8lOPQcfYImkDcs/zVze5fDPoAbnIeL0JeaUzMfdc/
HVMNVuhwn8m+mp41866d91RKOcz1tajqZvhl6RIomNJMVNA52REwLb7agTrMGBnJ
rYHL3dT4+iXXrwlpGhe5rT+TrJP7UhabduLjyiO0Ja1g7h8s1Oa0SL3vqnUDlsZv
VA+D3BsJpNvWKQT5tiksaDM09Hcw/gGVHRtOwDUz2oKY9wpCGVC6TNXcMEQFt2li
lKblSdd/bYWj8ksQPn98Ti3cqE+54lEZWaRi3EgRKF8LdWAPpIlIpbm0XDvrbQe5
Ex05SrUu3yBrwwBKtiggGK4J6oxCwyYlEFxnLysS5C0YmChmm/XoTaRwtjpc6BAU
3Buwlmyywk3dzEb9SOqjWaNWdUEIEZNY/xxcrdMxas5zM3DxJReSebmdYcjqt2OY
Ip/mRRR+EioIF7BfnkCQv8B7m4lMbMh6AzBiTF7DTNpCuQg9pAMPMRzgAlvVYcpx
vZwjIjzLqgRJ8KZE7VYNwM9CsYP3iWvfYuY+z5jNAIlmeQTElYQifpJ0QFuKzMXm
cpdhNZedryJOSeu4Adx1DLVNtf6pQgFfhPdc/swSOOgQa0AnA3sQHs4MRKPCHI1B
yFwBEb420yaeguuJNMv+rhQwOj1cfB59xu+P3ge8gIUTKif9Eslj+tYMwvirUQsJ
neegB5+TA+M7J+4r1BTmM357gx+m/PAxiZkWh30gIt5LzrqYsZ0EwkPeooyHCWT+
JupqP6/JamF/4tuPzjMabziS5LYuqwmsywXMhuxyqFhyt+5KkiDBemlW7z+unWSS
BENl8D15XqT4db1b6VrgE8+r5n2dPpjjbpV1DO897Nx8FKnF9fXgo9f3eL6bar5L
uEhss6CqfP4n3vkjrnUkBi/xLfX9UnpPNZQCjtLyauV9N3fcjE1Iwzkr2ivN7I/K
PI0m0us8huTlCA0eMrux8MitOdDEqO7BnPcVejbKOlQ5cW5+yk8G1tpRYJfH8s32
yKIPe6STg4bOOAx2GjZPiUK189YR2ZElIo1hXV6JmNhaGEMyNDbG3Yxz1EKp5kgS
x4Ntq3G3jI/BnfAds8zacSvhEW7k8LqrUDGiKWmUsp/CviSrWt2M8x+HVP7jOHi7
L6Sykc/305fhqZxKQg/3b3OnerQQ01IjxUQuON3J9vCiZo33WkumOip1VVN67Mwj
R9banMTzcbmI5Y+8uy+6cfYmyDPODwIIG9+4oWItzhTF2nS7n9C5At3sqEzhmGF2
3pI6xRE+PhR28xgW6F7hafX1UYDQank3hmLbMLHnL4fGfRTmeMr8P94MNm/69QaO
skm19R/Cj/WCoWSfnmcu33kraZVUVeGN+oSyhym9tB3UpZJ0QYF5el9ezmxz2NY0
lhPixlfHB2Idvq5Ty1D/T6z5k8HVjTQMbdBjM4WH+Zd1cZnDXwrGZqmLkDUoSp+b
TPdvCTIZTzYQiHeFBbdro7LVCoaz3qyMvP04QH2qh1CH+3h+PHrrZl+rvaGxoknK
iV3bv4M7ZkZNelqovpB5m8kyShuuj7XxQFHBvUaWNojB4M1XW428xwZCwh2n8yiN
`pragma protect end_protected
