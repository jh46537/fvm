��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�������s�h�qQ Ҵ�pp%�bs�!F1���|W��ٍi�\��չˇ���7Ge�+��9�*m@Mm��A��/f��XT��݌��GP�s��Ɔ4)c��f6�}jwS�����r��j����Īf�t�8J�gmdD����I��h9EWC0^����T�
�we�g 7H�����2�^/����t��PY��Ivs�b�q@>y�%K�~���*0p�w������
��w��{R�8u-C���_f(ZG��|���/zg��P�sIY+�e���<8%���⌚��8gn*rp,����_{���W���J��fM����D�~ۂx�Q|�hCުŶ�_����[�����������=�՞����6�����o��B�#A�����4��5s�32.�^�`�!c菂Q�h�;�wטvm���Jy�#�d�d��_ǫ&؁�	_�Y��O��k�r�P�]���{_)![u�����w�:�۵���u��\l�E�7�nj��V������`�1�M�k(6��5�Z�ʰ� 
�ΐX�oI���>����G����5d���c,f%T���`Z�� պθx�L3#y�("���^$?��R�L Tç��I�p�;N�0�)]pA9�6u�}�o�l4�4(���ۜ��\;�~��>��Θ:������ˁH4-'�[Խ4І�z��@���B�+���5�"��>x�2#+ؒ��)��f�5�hRB�n�))K�+�;������1O������<��MᎸA��ӓ��W��7��W]ۍr<RS�NJj}XSߖ�0��*��;�!�����0��Ԩ3.�!^dܑ�.W�����L���\�d2�?�?�(�n(����HB���Ws��٠�A���7?�Mh�]!�H!����VRF��J��`�bW��]��Z$t+�f\\|b"��`>�C�Y�%Ǵ	k�-�a}8���+'��0�To4'9�ɬ�9�,@( �+�٧���<foT�G�Hؾ��8L2� ��s=��ݖ�[�o�D�ܺ�6إߓ�ᓏE4�!+�׆���K��$74�z��]8:��XG9�R�+�㓶�w�����ώ��Jٷ�}[I}����f'��%ۺ+�"���2N
d���N@%7���D'��v�H$]/íb4�����o�f�='����4���0W?��"�y�H�J�X��[r��j�1E�����1�����M�u�,����#�YuWpO�>�,Ƙ�

Y.������Sv�\��`���[ݹ̆籇���ޢ���Vw��xE�@+
��J˓��3��jBPl������ɱɯ�"�`�Ĭ6����I����r�h����U��q�!Q�!5JҨ*�%N4�7
��I�K;n���Iƨ���.�KXv]=a(�KM���]�ѹ��~���xp�b�l�uq��&�?�`(τ������µ~U`��I���m�����e��l�n���KX�G�z�Dm���؛>���nþ�w��M�=�UU��+��p�G"G�ʑ�=��p]�¯��Of�e3���p�)�,�w3IER�����p1��pt� ��7P.s��chyI��������xX2҄yu@�仜�!`}���`��Y�o�%E�Hs�k��xJp���o�	T����d��-Sy�p%�&)i���Fc�rr$Y����fA�p�t�ql��
�H��͸�ƣt��DW�i�9��̼�\N���w���bt�7u�?OJ��U��rP��"�Qn���Y�|����7=Ξf��E餄&\|v��(�V���x;}K���*���'���WQג�k'�!W9�淓X��� g�?ȴ�F��z��U���\￙%ꝝ��t!^��-z��J-�S���;���XEˠ%�V��Ai���Ԝl�r��R{�k#�F��ę!�x�&�8ϕ�P�;�b����cg�%@��l�>���l$��]�H(�,z���C=�b��z��!�ϿK��f��/	��I��y%ſ���:�Q�O��x�b�̂-_ (��n��q�����ϋp�ؑ-��V���ZYuT�J���:��1�z(�tkl����1P�)�p�ֲ�~����)M�'��DY��%^�Lw`�c+��n\́`�N�˥��(�8;�%	�BV(���S��A6SvDN�\|8v�l�^1D��,�z��D�1��E�{�>¥�c�C.B֖��4h�k[F�/R�|��)ҏ���?�ץU
y��X��e�P}�Ǌ�Y뙧�+nF"H�X�q�l\�����áJ�\��:�wڝ]���$����sx�7��,|Țiy,H���p0w'4����D���:�I�=�-�$v�mGݎ(�{����2��֖PuȢ�E�M{$�|�:�@�U����� xۛi�2�ų$���4*-/�n�>�u.�-@���,�,�OYp
�p9K�=���`^(�h{.5��2��L�N�h^��v�0s�B7Q?�/����;����I&%si��̲q�q`�j�-��@���l�8dK2�d�lYJ�<�a�	���y|K�'8D:}��C��� K�Ϙ��+�F̢����2Q��5w�#�m���%�(�<��u���M�]�u���:�Wж�:F%j�R	E���TR��!��a
>�I���G���Q�[�BH���x=Jxd^�L�д'��,x [-�����l��]�(���w�47�vCf	��Im$l���#�`S`�O����H�i��84���5{r���v��ю�( )��Gn����p�X8�ѝi���V�?���v��y��wA�I�=�'�&��ֵ�
CK%�M�I:��3.0Ż�Z�J鐰u����7�s�/N�W��$������~|�|�=T A8�Аh��R$�I7�E�>g�m������E;,�!v�!������ch��pm-��NV�W�S�yPrAv����AW�[_l�i�"-�ץj:��L?%���f�� U2M���oM8A���+�x�3�Q�f�5��M�]�9��P6,�c�WD�A���z�hԶ��p��=��V�(7����C��Z:ʓ\k�l��H��kΓ��>.@�O�5�twx�$�SK��Tc��?]���?~�u���������^jC�@τ������o������^ ��F������/�T�'C]������W�<,D��{+$�S[x_m������S4c�A�a3�B�b�A�uZ�a_�h��UQ^7?m�ts�rz6�p�7S����cY:E��l�H��II6Y6+:aF��|
��0j���!���X"+ES�xK�HU�n/�Ɍ�v�+Pg��"��^�s|P�k�����9�{&��8^�l�U�!0%UĎS��Fdҗ�h���:�E�}�.�
;�F�x�xw Q�ˊ�$j��w��Z-��gxX�.S�����퉞�D'i�� ���7��FZ�ڵ�K�I�}ߋ�1�H�& ��J���:& �ڐ�IC�wv1WE.��"�:��Wڋ�\��Ɩk~��-&�g�.B�aIݴ�~�A6�*�����R����AJ9�R�z	m<8�L��`^	<B\L�|��A߶�W͐�����c�(��N�K�≝�z��ue���	s�C}�
vܿ���ԅ����`a�v��h۔K��r����GBp�Z1	V�pD�����x��Z�@��͚���h�v����,�l(!p��mv����'뽇�m@_mb�D�r��y=Bh;�����ГzX��?�	O���G�? ׼aQ�r���H��R�.�����
WX��s!d9֗H����R�� ����\����'\�9SJ�^���߀�X��Σ
�4�x#Ζ� }��7H�ؓ"�en�����W��_a�'��	�����)2�9ر(��h�Q;���\+dD��|�y��0݉��v��&�)*G��(D4Ι��&�-��o�=틪�jo]d�z���W�U�cR4wJ��{Y��W����������"}�_�����?��>�̨O��+�HhF�M��������n�$��h�����M�k��DrV�>��݊����+7��|���#�w���!��^N����vcA�W�1C����[͕�I�}�[��O�r>^�l�6B��tko�k�d'A�E�I�	u�	$��"���+_�R�����2��/K�񤿣����vcj!�梨fq��.��~k7f�suVu�%�Q�o1<�s�l�l�!��⩊YA���Y�w�H ʹkYW0Ë��m�� �/�EM>��`�e���E2<3<���,�h/�.&@k�l��|!\��̮t�h%&��1�\��~f�����^i�1��K�*p�
���� 1b<�n:�f�?Ԅ�]����U���`֮�6�,�v5!�u���QP�d�!�����,��|v���C�fP�9)a� �Kv����{8�{̣Q�"�v1T3b&�8e`�<b�7�w��b�����?`^K.��(j�}���`��7%����U�Z>O��h�\�yP2���j^��j(�~R�PD��L��9��I*����}9@��J�P� �x\M>F��H�Q�^���8^�-�ͼ�c����+T��}�'����"�myt�ڵ��F	�<K ��v��Ɗ�-�m��c���i�z�ZD�ػ���Sj4���������Ȭ�+w�L��&��׽�i�]U˯'>g��-��i����Z���2��m�Rة0Y�Ϻ�\Pl�x���=J�UN�U�6�r��?\��5ך(^Z?�("��ahB����e�qSu����5����Zm��Q�����P$F�0��.���J`�.c�8 ���&/��4�)�N���G}�|�v|�����l��i�Rc�	`6�x�z���#pd��zl�)�~2��^_Vy�J�k#�>�]+����n�`GV�r�J�u.�_~�+7m�Р6���B8��|h��Բ�� ��`�=;*��]�l���0��2�zX��e���ӫ�Y����8'r��TG/���%4R���T���y�A�9���Skv���u"-�P'g��R�������|���~K{�[�Ӟ-?�+T�B]*&�d� ��\�R�$ӈ4���""��\�dFĠ�K�nͬ�S�t�ݮ�v���_���qx@܎Q�h��؍Yi���(�PU2U�C�z�� ���S��'ֈIu�'�W��[��[��~�DD�`��fc������N�z$㆟o��*�g��_W���@�����Ss��F����ړ�E�q�G�Vr˸�.��h�
��� q_{�]�~_,E9� ˫1��jP}���p�LXgy�K$�"o$@�Y��LXrKv�S���K�:k��hwȏ�J =}-��+�Y�as��U{eK74��W9�g���5�t�t�������wAA���n,�~�|��+�@H����)j� n�|RWQ��O$"<*�&Ͳ{�:ev# �^��Yj���Y�z�?Q��篍�ո"����3��>�lc+�4����n���k64����Z��ղR�?B7G�L_�v�?�|#PJ]��\�I��.fm���}G/"��T�!��:�X��`�(��M�+�j�����`��	>XR�����婦ö��2e<�S�cp�7�.=�ȯ�(���<x`Ax�C�M�����p5~2F���U7�
�|�MG�IG.���؊P�.1��"$m�����y����Njyk��kF'���-�"D*4�������GDv=�^�jU������{;
+E��q���w�7�vˍy�8����걔ce�b��9���&����`�)�ع:^Ɛ)|��hK�7�>bΗL�>3G��z���@�Ԍ	'�S�-_�=���U����&sB@mUoh{�4���?�L�c��&oƕ��Nj�1�������XzpM�=[�k�U�(y�/M��N���>�{c*�K��)F�7�:s��":����0�t���A�X��tO�Zj����U�C7��$�vE�#�X�Qo}FV:� �Ͷ-���?�>_T�c-����J�Ga!�+�Ќ�'-A�����E4\e��k�?=n����֒<��P��'b���-�zz9(�D��=���� �~��3!,�D�1�IZ�_��2�����^�^��j/����[?p2ғaX���.�F�dyxr�Tښ �&8�����V���$� � F��w}Ps$����qi�H����C�E�W 1��Q�/���'p�Xvho�$;�]��)���O]➙�<����R�3f������6����9���/��e�=k�BQ��$�w[�2#K�G���o���^����mڮ�ո�/q&p���W��?CJm/��ɾ1��E:��)z�)�7�RL��橠���W��#
��� �� Hq�E�2�������HC���0�@*��"�_��`�ҽ��|��W�7&(�%��,S��:~�P_-0��2�h�QUbn��M]`��3�b����t�d��� _)X��u��!8��L?vr�:����]!1� ��3��CAuP�?�[�d��|~�;<�5Q�
w9�):a����rw��gb��ՊR���m��mUX�����}�����ѲO>���(-ʵ_ bo�K����$3m�d� b�����9��a��Pꃑ������n/ƕ� vSd�Q�)i;Us���*҉�r��CI��w&��"���m��~7s�*KJD��XBS{s���e
�8^�S�K�[�̎�'�����&�W
4�>�hu���d4y�O�G��ks��r��Rv�,"�W�X��L�y'Oe���۫VF�̉����2kF����>�s����鑠߲��S��Xl�D�#8�*�R��S����|�ej~�����V\|`�ؔ��.���7+-�s�Z����Ǹ�:06I�޼�R�8ɜ�(F7Q�q7��L���N��Oq��<$(�ե���q0���x�5Rt�ի1;ZՑ�~wO9_���5�C]_�&�P�`�����7L�(��k��g]HZB���f�?�W|�M�b��X�U��K��U�M�H�<>��TU�ƴ��Sjڲ̳-F'>Ul�o�����KK_��i'
���u�?�Qc"���'交�'�Rt�L���{}�F4G�/���:�r+�V.�]��8�N��"��&�qi�{�+p`63%}���E.ˢ֥[kaJN�f��C���׮:=��/[ć5�k�U�]�y�w>�`���P*A<��a2۶����yC%�&;��|�!ÊbA=�ds�k�F���[ӭR
 �.�o7�} 
�"6�� ��\Q���F��w��q�Z��|��Q�G=��\7�|�QH�{���3[6��$�>'�\0U�7���u�[��@�h����T0<�3s���h���t1�z�(�|�z-��,\��E��C��̵���b�w|P@�U��m<eو��DV'%�8�*�ͩm���4#��V�y���^�/),I![���:�ԃ��s�~�7Q��i*��Й�3Ag�%��ĕ��d�����T��+,�M���֖ۮ�T�0�����������>����[M�FM�/��Z�<���F=��P�p��F�g=���k�"\�Zb�+K���c$�-��K�2d}�	[��ػ0�N�qD��`���M1�>e7�����Ҙ�_n|��O��U�)x����vn�����"�}A�Q���1�k�u|�a��5Vt�}�/z5�ށ��+����v�������U2���Z�e�y?�4��h��V/���I�f�"7fe���@�DY��[��ʇ��:A��ʢ'u�ai������NG^���V9�=>INQ�9{��U�6�	8��iV�c,�l����~���c��Ng
 ���g\Ĥ]cqw|�-";9���5��şPY)��A�ݐQ�p���R�K��0`DC!J��J�FN$T��B/�RBSYu�����0��WZ�� hZ���y-F'�>��e���jJj�6"%Yp����".v|nS^K�x7Y|�X�f1�y��U�'t����XW�ơ>ЬK���P�w����5���e{�u�8�Ms'�t���Y�k1���f���N��{Ak����'/i:���k�/k\+܍�%��fnPΌ���]Lw�~���v�th���J���ǃ�ɜ�d�e��Ӏ�ڵCz��!���.B)?E������ۆ4���Ϣ=h*�J4�~��DS�Wэ���:��O��L}�}n�t�-/�,{�<-?�0�	]�(V㩄�tt�羷ss���IU�)r,����C6����s�#�-	���G���!��SZ��qW[����%cQcS���z=�c�V�.(�]�j��Z�)���aa*N��|����T9Nv;����[^L:u<0rc_�U�eB=��s��������%��*�j@ݏ!xJ���� S�"��Q�8t�ÐS%��s�g����y{�nb!S6�%1�;YQ�M	���L��P'&<'5ÐC?��cgj`����t����ӌ/�-�J	�閙ø[%�p{�H{�4r��53��~d���
�%���4���'�\�퍟^����l܈�y���w?���%�V'Z'�\��P&yMD�lr����3����g$a  )3��\��k<˄N ;�H远�²)q��Y������:���JQ
�ཀm��q�;P����.���%�QHd�I|��(C��#��f��3+F���ܹ)�-�iݣ72sB}�;;�wdM�����)������,k�ܸ�8�i�By�շ����i�̗ZjJ���VD�Ws&��٦��}��e��vw����>l�@Rbu��b��_Y�x͵��b�L1�~'��2$�K|��!t��oI�� s������F��FPA�m�~\�_��> ������Ā�ڋ+���Q�.��@`����� �`���H��MR�D�/���(A@/[l�1����\[������^�	l>�������qfs��= 1���y.Uk�3���{�jƹds���o%N��l���r�X�Cϙ��w>�]n�.A�Nn[�a��Y\��7��[���\D��`�v�NbdG���F��{Wh���������8���������iN`�����:y�ꕱ�R�.�݄i���N�諑B6�m�P��W��d�z�4�u�f�#)�y[��tҋ�ǆ��;�|���e�R��d�q�&��&���EBu��Ϋ!ߔ����A�ˣ����8t��D���x�>/˼�:�T�6桧?f��w�o7� -,/~>���
��J�:��6��Y����ڿ�@9��:ђ�P�6�Ε��a��Q��lk� �|Ÿ��ܛ��jͪ�
a@��0n3�bM�D�2�����U��p����1'��(�[�� ��c�2RFB#�̮~h���z�s��{�,���ɯ&�!"�XK>�H|ņAvp�Ρ/��~�â��hm��;������KN<�b1�X�J�Z���$�r��y(�P��*F���8 ��8�;�d1��2�T���6 cfe)�6Y���ڝN�;N�Y�_�+�pq�hO�?g���
�0�z�<�K�Y���oM�@l������N �����_�p��1ǧ��3�e	�&Ы;>5U�w!����*:�C+\jp������s2�csJIҼ�YoN9��[]�pm�ɉ�G��`l�5"�V�c\$r��Q!h2��A~���
T� ����eɖ0��{��������_��i��?M(Rx*mF1�ܪ��0z�T���FA�b���������ƻ�A���yyD�Ea<i���MQ�!��D:FPG�/Ih���|�/
r���̔,���}��|��/�n��z/�
�#h�ZZ$H�b߻�:jd!�Q�C��z�����4%1M8'�����@i�'�03��A�G���ʮ����bD�2�����L��¶N����`�81�<����,�E~��4鰿G����=ryi[��A��C�x@"�T�@,2�>)�{�(T��lf�i�IJ�0�R�m�>|fb6�dE�lH 	3!f�9�L�+L� �q?��D`���A`���x�9]��b�if�����g�&m��7�'2�P������������Hȋ�����C5l6�Ct�X��VJi�0�c6^&���D�F���_8�L�g*m�:��7=�Ȉ�E۵��K�u�O��]���`�b[ȟ�� �������+/�5,�mP3:��j+w��~�N~���{���7fPu� .��N	�|s������.���|k-$6[�as�X�s�W�,��x/5]�f���+��$��)���!LK�'�6�����]{���D��qyf8�5#?���X�~o���ϛ1�#!���I �Y[�9�+��|������Qۥ/O�kzP�:U�H�����JkC�^�й޲f��q�k�s��X#��80����g_&���%�'�6�8�� /��>�<Y�-�$� K  �.l�Ϧ����}��A�P"�%qK�g�C5�/razJ	W�B p��5S�ޜy�Y'��_�<��(� Z�,(��|�Sv��qh�޿c�½�)�=�2+�	8����:S?����;K��s?��|܄PLU��X��3%#�ջY]龴,2�/�����h�d���>j�d�nn	��?�ZWR_I�SM���a�}v��z��7PMq
��$�2��F!��X^ٵ��>���t3@40��]{ g/"qM�%�v���cJ��ۓ?Uc����ӕCk�aN��V�JD]a`����	1 +�}P�ֻzer�� ���4�:o�c�KS�"i�7M�|Q=�#L�������b��u��(��{��	`��9tM��n�rQ<�DT.�T�}�s8���z6��z����<�P�����A\i��[�&H�/W<�O�,eH�
P�"l+	��4��W\y�45'�N	�vR�v߂%s9af;�*%��F��������f6ш7��}����x�;+��}ZC�"� �� ݕ3]�݌ <�\�aQ����2���Z��-9�i�7d�^'��i0~�#E#������Uy��%qrZ�;�?�d���ҸI��j�1	;������J���֌��������8��[��0t��+B,ْ��;5�xp�Ƒ�RQC[ ��!6�Ts�_�D�I��H�W�y��+=����O�|o�1	�Ra�7�6���w�_&�5�>��LH�)�-�"�i�EG@)\��#l��i5r�e� oȀ�2���Ɛ�u��Dj���H��	�m���9�s���>�â�oP���(v-�~�򫝁�"B	d8�n����	O��ĭo��*7��wϙ�z����mk��h���~ 
�iPY53q��A;x1�rr4�����3��q�N�hn� ����fi�^֗a��-�mX��;|���jm�čC�S�3��|#�'r�y�]w]2��9�c8�H��ܹ�.�5����VQŃ�� �4������Ƨϧ�D���&n8�BƳ &�|�ea�b0������:�;O�۟�����Ase�8֏���7V{�#�w�J�9�3'�Uco.�?��3�]��> t�3\k��:\��^Y'����R�F�౼��7�*a	�Ӌ������°�j2�����1�㋗�B�a��|���G�ϊ�6kƍʹ��K,�3��hʶ��ã���݃ bsF�BE�|k��(����q��4��0��zv��[�I� �빚?c�"	�c�/��v�_%�]���M�t�
����P�2����g��ݨ��q��7a��@J�=}v�v�X[���U�V�o� ��yi�\��Ɇ��B�ḃ�tժ�-=��߰�۔.��p���޲ˋI;A�'�n��_�o�T!�mk�唢@Q���e[o��FN{����)�c��яA�u���*��s���h�Щ��� &�9.��+I�K��U�	�!2m�Lɔ��&�G0�f	����n��L�X*���{������ yVQF&z�=�rK�fݛ�Q6'X�I1��z��꒹�(�*cK���� E|s֏TG�RVg���k#�����9�{�]��kR2"Tl�;(�۴��c5��Ҫ�!��Z)����/�Dq��*�j�sN��X�W
��]
��$[�ޔ��6�u�sS�	��C��u�%��:�ʱ��r����y��BUmm�_�#a t4�b�a�w/�^+��vy{�An�x@�N|��<���Lb,e�~ЊD���Dp�<b�)1$���h��v!#�o�oƾXP�t��^���"o�ط������k1ՊT����IR&$H(�15�	ʕ+���%���67���P���jzļ��:%�P�T��M>�}ATFtYq�V�؞>�\�x(�?a�`��1g�$��<�{v��U��6fq�\��䛉
�������9
�h�tc��ɬ,YDK7s
�l�7����m(C� ��C�����3� �l��h��aE׏x�X�����PJ#�W�>�y���-4�Z��|]Ssd$G6f����h���P� PT�C(m8^�8F�qk)Z�n�Ҟ(�ϵI��J�1����K���2J]h; �Y���/�`�8�Zh��bv	��F�4
�Xr�7	yN%�5)b���0�W����$u�0��+���aW=���
E8���J�=�Ƿ����u�O���>��ax�"�����f���R�-�2��j"i*�*��)����#g	{o��]c��l@��G�d�@�Jտ��J;$�Qhu?�O�_ J���.|q�#���wJ�t��� �NW����$N�m9�='���B�>�f�@�@�A�좝$����C,�h]�i����o�����D�ݩNQ�1H+Z��ư���.��N��J�팆�-�3��3Ҷ�$��8���~�q��P�~��A:ڳvU�:��Yq�<�>���)���j���q׀��6p��Jl"[<|8(�(CJR�p�e�v�ۚ��6�ޫ9 zI�g=$�%43Aeaw��w����F�8T ~I�˿B,ə�y X����0:�Dx3t�ȁ�L�(d�i�U�3LS���%��!�8j)@��9�̸=+ )����`�ɏ�\*�w�$���HsA]W�ƽ�IXc�&�4���&�� ��\��e��	òp����5�T�����Bۼ�,�6�y@�>���&��:pI7�jXD+֊YS��s�W����飯���uL�4��g�&a%���[\�Ou��h�y�G~]R3�{_�`7���*>���g�B��ƌČ�\�x�li�;rqt�؜��f��������
��f
eF
��_��7�X �^
�3�?|��n�����j\he�#Kɺ�D�&��!wy�4����"e�k�'�I��qs��pP? �8_�ޭ���y��vO�Xk�!��@�E�?��m�/�����~�f�n�|�7,����Y2:Dj5o�����n��bK<(A�?_�aD����J�L n�\�+�-��+�hA"����Ŗ�9H��KD�鬏����  �f��ڪfw)��8����gZs�]FSت�^#�x��N�:Y5���A��\��P/z�7��ȕY))�G�N2Oڋ)2l�r|��Id�RD��o���S�|��/!YF��‵��"�����J�NM�2����zj9��L�ʫ�y�&C72չ5�̰�8�×���Z?X�M=cބ��a�bo(t*%�? ('�c��i�6Z�)�?_3S�Z���#��A�e>c�Q޽w�zr2S��ma@���O�`|�VuJy�ھ��*~�=�%V��8�N�5i
�2Sz�0<3̤	8릙Bn1�I�(^4zosB:��Sa-��Ǡ�����O*x�A/�Y� �hց��5�:�@%��ŝ]����j?��3ޢ����]��"i�#��Կ�Î���q��v$+��ë��W���gY��BNaW��1'k	$��0ܱAҕW����݆�f��j�y�=9��|��o������G\t�nR�|�Z�DiȗZ�a���K	����k(���]�9�O�l��C��WR��@ޒi-%
G�G\�LT��Z�� �� w�NrzQ���o��}�z��H*�4����@���ŤK"�zp���+�N�`��������:�棏&d}��I�r�=��Z:�qT�!1�]
/	J���N��Zs]u��h�~O[����!��|
ۭ���[rpMJ'�bL zU�5���ll�#Ӈ�K�g`�d���w�,"����yE�=B��Y�_�����"-'�}���p� �@���b��5A�Ey��"�Г�����-W��
�}�?5&x;d�H֘��G�#�Fv35D�r(>�a6��j�Y7t�J��wNϼ�$���y���r�`��?�h[�`=�d,桍���ux|�p>���>ZBcoðM�̌�;��(_��<��qEu7q#�9�Ķ���mT��	� ��,���#	س	<���.�V�.3��c�z����3
���(�49�[o^�.L��^F������t��O��C�8�(�~�� \�C�ezp�Ϯ�̓T�c���b/�z��~� n�rN��.�]�&���Ӌ���iBB0j���_�5���	����T7����A�W/�7��U���`y�����$n���Ue4���b=��|=$H�p��$�����-���D@r��Mw���`��>���%��&Zn�=�b��ރ���4Va�֍�8ڂeTϞ�bF�Yp��j��D@s'\��a�c���5>Z{f��~ [� i�ۂ�t����`�tv�@��s;�l�n@��S���p4��8>�Ys"���Ѽ=;�p^s�-��~�����J,=l�0hj��*=K��pU�=(�Il�(�g#4����@H��x�k@��#N�y�2�N����e2 ,|;{!�ғ9�ɒǁ`�����E��8ܗD���*SE%G��X���`c�Bno}�Z��d\nNĜO��\�Z4ٛ"��o�+�K��r�\����IX{Ȇ$--<U���y�'x���Sq�-��Vn�[��tIO|�2	��M�w�u������&�U<u�7��/�oQq<���Uo�W+Bܑ.r<9�{9�m�[���e�8b"hB����i��np�:e%`Ӛ�����jގS�\%K}�1 6������[~,��%K��<6	*Wn"L��c��=�H,З�B$2�aü�_�@��]���T�N�� l��p��&��Ș�0F��'���F�dZ����tO�A�n���� {}0�P�Ƕ�DK���](�!27
{D��}xv�EwTP�_�� 5";Ƿ�����7T����ſ
��j���X��o�R��v(`� VQ����Zʳ�1��3����O��Ĕ�8yD�ߌ5�ڨ'�f.K���wHE:�U��р�_��Ly�CE�ӢT�\\@�qp �?Ղ�m���נ��e$2�p� �:ԛ;*]�%��K�A�7#m���:\�I1>�50�}�:%��H^ʅ�0;�]�R�q�="�[&�h��lf�"x�_�5���N� ��,0�苃��}M|o�%Q	�L���I�ā`9�ů������������)��J��r�tě̟��\�&�8��Vdr��hA�E�SMa��g�� ���|����Y��L^�b�=�w�[W�L*:�'��e��t��<��W`\e�h�n�����,B9����6c���%���)Y�T��_5"�y� �誸(���}�تC=~�+�b�.��)���`�G��v��!O����O][�aJ~��_.�K ��e]Ti��\��g	9���>W���G�	W���<6N}x@�v�㨑��O�ƕr"'��O3R�?�E�5�`x��Np4R�O.�'�J�Ot)�X���JOǛ)�Gɔ��}�c�[˅n��!��K=(�06U�y
�h��鲟2�'ni��jd���������4�ا�����w��y��-Ɯ�g'���n����C�s
�a�@\�'�T����k�-;>�9a�E"��\�J�D��W�?�k_{��$~;Ȓ��'H��y����������Ll)��R�"� �(��U����JFϒ�g�4�}��Ն1��_� ��h� ���AN�lޙ�u�i��<̝��,|�� �@Do8��>���~2�����|��^��WdL<�3+�u�'����+����9�J/�����m�|�4���ro�#��l����
��S�I�=���҈mk�D[w�&���7@�[�fz�o4 ��ڕ�����T��E�-W=��L���)��MK��1����1�B�T
:P��9^���`'�!x)�Y e���ݐ�"�"(b� ��Q]��r�� M���D�4?d����6Ay�KS�g�B��-��Yج B�0^%�N�;��j��4��}��pU#i�(�H��a?]�N�Ƶ]`�JE ͔x5����m}s]r�q�k 1E%����sc�g|�^���жӍ�[�m�N|��(��h#8��� v{A�53��w7��+׊1J���B寜S�A��X�������u�ޞϢ�ϣ+��0��̜X���$1Y~���"�L3P*�/(4�,U��C	s-'�-G�D$�zG��B�>;�1��V�ʟfX���nn������粀A����>�(���#�]e�`��������e��:��XqE��#N���}������_fa��bR�{x{��Ҏ�ϝ�{uC��G�*Cl�Њ]���P�R������2�`��/?�h�⒔���|�?����GIp8��x�q��@�;NLK.��׵�����]3�.�WҾU7���v^��Cw��q��ʀ^i#��9Z��j����ug��|�\�<��<h��-˝������,I����"e �Y�l���1��r���%�z�	!JY1�����7sSm���e����fZ��l�p�?�]���J�2����e؍��w�{.�j`;&��}t��!��1U%��=E�}�?l�����9?-ʔߜѾB�!�lZ]r�  �Q �c?Q�"9�z��t��Y�qX��?��Ԏ4R��/�,ǿ|[Uf���y�X���Z�z'�=��ZTT[�ҏ/:!W���֕y�fQb�����T��@��#'_�]�ʟ#�g��/)�3ʬᣩ.��lovC�C�(�z�|�l<|�}+�?]n��Qg�䅯�H��xr���K�P�XJF(�T�5��vmu�%�� +e���9t�"�_��r�*:�]�K��1�Mc���aۺ"+hW����:��i=[�����:ܚK�M<�<��m�웩";�9��/�m��A| "��Hʌ[���ʫs�e9�jE
�J�d��o�����7�k%a��L���:܈��O��L��6Η��ɤ�ʛ�L�ޘ}�@~���(����h/�m$�57����pߜ�8b�?n젗�-�D�O��Ar;����,��x'\��X�`��K��(�9��f'���]�d�U���;yz�W��^q�>�	��~�/�2�o��	T�LD���W�q�7%���?U�-�?x��'S)h���u���eL#��*��M��m�=p��d8�L�X3C�,�_�B���~���,������è�@�����ŋ��S����dz;svU�_�pNA��8���7�˪k>�/�n�.�7�6q�o �9X���C����1`g����4�kj�t��(66�֮ݟE��M`'#�ˢ��$��]v���,��C�A��c�c8�l<�kg������� O��=�H�Hl�i��E޿H�Y +8ɒ)RC�p�m��b�t����8�V`�.��V��L����YQ��f��
����A7'tNT}f�`@����)�N�5�EzЧ��َ�u���j�&�e���z�ߨ1���*=D��-�d_�6�઼�_�'X�:�~�w � jD��t�P�1��p<=�me�]5�Fg:;�u��	��e�,�v|�f��7�6<ʹJ]���s#��*:f�s�������ts�����f������h��O�2X���@����Í�=R��A�j>ҝ�j�=��:{-�t���ޑ�X쫪�����4A;����TA��޴x$)K��k�b�z��N����!�?%�|0��6����{l�6o<�J�C�UZ[���:{������ K��3I�y��O��?w�HX8'Vj��(���G;�K1?��x�%f����Bl;��ge�=S �����������_�2��E��3��SQ9��M"D�?m �7?NҀ�\��)�Y5��6�_�};��H}���r�"R8�E�Z���[�����<e3\�d��ȍ�Y��1��d�o�*�w�^�I��O���*8(��-�������p��p���F���q��gq,zz̋+�҅��G��w�dm�A��mb�>Q��bfY#C�tG�-4	P��}H33�r����Ћ2�`Ǯ����;�h�	
D��f��t�|s7�ݦ����ch�m��AZ=]Q��Yn�"�&��x	+;���֦���:������#`-|`�k(�("��PA���:C�j5Y�$��`��}X��'a�c�i�{ʎM�z_t��Q|�xV=�ԕ��� ..�ch��iu��)��")���CqD�tY�Cnm����w�/'w'"9�g],&�g�/���03�"��UX�$zI�����+�n�{JK� ���ߊ䫹��N��MF>mß�(B3�t�q�8���H_�����
�����\P�)уn֎q�;zY�d�q��ߡ��p��c�jx),��[-�3ޣ�\�%>�y�0UI�s8`���v��Fj������z�y��, ��s�c�����M�pa���C;��R�A���>!({/���ZU�	G���<�3�s"�ռ����̹��jr�&�S!�E�Tp
p�ԅ=	_�,?����k�<(&����W&ǫ�8�ŋ���4�h�Y�mE�"qyY<T���f�VY�O���ug�^34����;ck,�#���!z9[	S����!<���@1�l=�C}=�*I{�嫨����|���ײ������#GD6��fP�%h�[@a�wI#�H��УC�៺�jag��X��e��J��#�m/��}&���,h"�c�J�W��T~s�l���(�c��u@� �x�[A�X�cU��%� �%'��Ɉ�C�5������H�?)��j0�\�Z�TRr-����>��l�g�$�@� Sso0��<s�Ͼ�РN?Y�}'���+9Mb!��͛Zȼ�������B��� ��G��!&Ů��4rD��/7m�5UFu��&o;K��&�����%}����Ue����8z����>.��7���i�7IV�f�=��W!�J�kq25��6����N
�9�@6v������Ij�rY*2vIf8m-Jrt�4;\��t
UB&�T/`pE��xt=j��b�p�R��
UQE�v�}�,a�U���m�A�hVNE	������)_����x�Z&Zi��e���V[�{4�8k�X�s��5��O�/��j�{�W���q�;J:��{=u�%CI�K���P:}�}��ڦ��5�P;H��ۈ�Da�R�+g�o�[��4Kb=�÷�p �q>Y	p`�$Nț�Khy�c�އV�B���5�/�}��,bGS�*.��g��v[?{>�+Ȋ��m�,��%��C�@��hU4��"�.ِ./B*�*���1mFuB�
�:3\�#�s�5ؕ�EQ}J��y4��D�
EQ'�EK��nַƥ8(�U$�����.�`�1�2�DL}(ir��iU�BT[%��R#F�)���g��!��6m��r0����ќ�FOdS��y�	�l	����Hђ�{���|��k;��F|N��q�cn�m�J�<�-.*~$�EZF&���ltkt.��1"o��}lH�iXud�ZY�����ƘsNj������t�RJ9N\�0(?:��d,f�7��q,Y��_ Zk���&xJ,7C�����K	�9oGTshe㻒�����a��_f���X,��x��~�=k!]4ޭ�rA���[4���w���>����A��(�~��&�/��Nw�_n�ئF��=�.��D�<�[�|�^��Ŕ��Pb�9����*]��y��z�J=P��o��q��Ev�Ӕl �&�D���>mI��.I �������:8���k+�p��Im������5p��.�4�yK�����U&p2,M ���m�3U�S�Pĵ�W��� *��~�5�}b�̛���{�}��g-��?�wl�u����5�Q	)���eA��G^�����Fx�<k�=/=����L�Ļ�K�	�R�m��@����7���I�~~2���޴s?w�-���^�H�����F�6��³�Y�FQ�Y�Zrg��z-N�%Z�EtzZ��S��^�X�G�E�%����<�_^��[w:� ��ģ�^9?�� �s���}��dc��