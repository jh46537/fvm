��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c����W�3��1���[�!���s[¬C���ۙf/)�'M�]����ῲ�!�hL�;�Y��jw Ήf�mU̚eL�!5��]!tsk��Y����F�y���QlJN,��ސ]������#f�f��P�'�̜9�q'�<b��M �.!�d��-kN%r�]�ٟ�as�j�1hVqjJq^����^SM�a�Nf�R�`�j�Wu��	����KD�����A��=���C��%�:ކe�)l���!M�<�j%���{����<���㏕���lv��7�3&0dp�vWU�ڣlŋ��o;�:c'���(��?71�K {*K������i��9�L"$v�����Ĥ��U����^��/�Z7�������^$	4��E�5��,-�x������&���Vm\:F��1DE$2�(d�-�oЩ8bS��c�"bBaE�Ωىc�^�ii����}��Ә�$Ǐ,l�o"�(_b�<G��E(�l/n~��D��A�Qvb�dl���u+66%��0��Ŏ¢f*�l�x���.�bKr��v.�i�S8oQ����r�Pw�R�%Xf� !��u
����"� ���5����*y(���$9��C&'�״�y�1��g1�b�:?�f�|l�_�i�₁���shE�(�qM�70�`i�%)���5��Y�^�ui��w�����!
y�pNİ�<bGe�<��Ԥc0�_�R:���z�a�JG�)�d\~-�Sў|��̽w�Ť�qUS�$v��83ϕB��F��yrNI+�is1��!�-9�`E�j�]9S��DT^�.3Exb�ч����XC�|n���H
h�n��>D!�燮�ήm���u�z�$�% �] W#ӗ�Ƨ$�(g�����U�l,2��m�W�,��/d�e��+�� f��+9,����`4��k���E|9+�z{J����%W�Z��U����,�'����L���v@�9��4�Ccc:�qO�g���eV"E�qr�ȹ�mN� o�	�޴�Z�'T��t,Ի�Hr�� �ӕ���v����h�S�3/�KQ[���k=�G�>*���۲���"�������59fÆO4�����z�y��Wl`�M8�`xT�/1��>�'%g3�ݬ�c��}�>��+^�*4]<Qjo��P�zwI�F�e�ߴ�.�H�M�V�jkԇ��%��>Xܭ�;���I�]i.�-�OC�t�-+u;J��x}& ���))Q��E��~��ĩG���s��G�3U�`�¼�?v5Zhސ��rwQ�>���4�Ra`4��rh���Ҭ��6���q�SYn�ډ`�s�Yx���"8��{1�N\�*|��`&�vw-�����`�z�]-� d0���1�IB3Ǫ������[T�D�9٪[U3�!wr��%3�����"�
�J;���9Z�h=�.1��8]�V����9^��r�G)��R{�D�JAi��ďGK��=��w���徇2�W���!ϳ������E���7>ɴ��f�4���\�,,��oB��@F�Ҳ� ��~T�t����= ���:ao��Cݏ�"��]{���qXm�E������# ,��NG�Fs���Yd�9�_���g�07�rݽ�Hɢ}s秈�x�/C)�����H��w�'E�\�Δ�0� ��E���W?�|��[�0~z����c�T0�s�3�[�s�����
�=��,.��\&��i;^�����|�ݔL��4�5���-7%�0�é�� 1і���gU��Gm��z{H{�\��b�g��(\�F��<�3�ѳ��W��(��l���G�8�T�V��Ɨ�ߢz��B����Ü1`���B���Z7`��X1{B��l��\ X�YZ�e�I���S�&�Kώ�S��%im �P1$�/[�$"a{��5z����������L����X��ΧX�r¾�$�eP���t1�cu�7��=���E�*��؄��*�3��f��:����/�������5P���+[El�XI�=��B����[t�R�*��P��lŧ�����z�9Ý����<�X)��A[�&�
)K^���GP'1�t����xy����Bu�P�ŝc�[�cW�TC
M�ߨ�2 �,���H� j|}@��z�C��i�/�LGh�E��i�Q���7D�#G4;���U)5��3�S�<a���4j���\�!��*>�2/B�t��m��ɵ4���3_��~{�z�ɜs;�4�t�]��v|� ,B��7�!Strx���c�(p����}�������YZ�H�Ʀը�+��s�#ȓ���[�1ë�5�f
'D�	\F6�C���dz�JMi�}�}N.:��_g�:��[�x��I�,��TH������}͜��'�!��{�0�ڮ��Y�2Gc�fvY3�Q3_*�"2%('wãYI�O���Lўz�������__eٓ������ƨa�MފE>
`�P��YGF�����L��e��t��(Vm�����P��p��"��.Т���L,����X�!��4�r� nv�)�]�C�!�=�Htҟ°���(�o��ܔ��Bo���^��p�I��f�T]r'��0��tjW�{e�4�ҵ����*ע%�:�'�0��E-�-�D�����x>�I:2E�G^��Gv������O���q!�V'C� ��6Y�Vx^����y�n�tx���Kz&q
߰2H�"�jJAhf�z�<�ʾ��
��{1JB�`d靅XN <BYam�<Ƿ����?��֙��yҚ�s(=�Ij?�:���s�ʡK׮)��~9� �p�0�I#D@�IH��D�"*I�
�:*:v�F��'�H����CS�����E�e-@h'�3�)�AF�v�������*��ۺ�֚�XJ̶�Š�C9���i��p��:d�����ƣ���1�C'\�������|uH#W�f�J���(%xE�nQOx����x��CRQ�AX���3R�W��n6o�D�c�e(l#�(��\.ð�D�r��-+�522,�:�<�=�����:%�I�@�� M�s@[�c���M���#�<���:'���<�������~C�4���ޘ��r�:B�J|�☗�����Y�{W�>8�4^�0�O3�1j�./��ϹIV�����z�Q����M�M��E@��@p]�n�Ȭa�>���2%A:��V��� ��B�?s��m��������(��^7@F���5������,���7���P	c�X=�W���Qe�ų�VA��YǊ���]xP���QW]�ـ�`]w�H�m«U�G�m��
��M���$�{�:΁�Sp�Ը��
F�}���	�}��1͡�����}f<�.�H
JTUR�q��ѽ)��a���{����JZ�F�贈�]���1�ح�ѡ�rx~(�9��j�/�H�!z��8����W3Z�r��s4�ꄱ�o��~-*s�t�R|�[��1�G�gӠ4���EM����	�0+�<Q
e6$?�Q6��s�B��<�96�p9ᮇK��.ʡd藾���z�`��3�]y���+�J*۾�=�|[in�K��U[n �g�OD�J��\�P���W07ؒ�������0��#�?��?f�oۭDZ߻��/dּ�(rC�T��J����$O/<\�/��>0��~LT�L��vW�0��)�%�!)�\�Q��I�����l&N�l'�ѴR�mFv.��" v���������Q�ǖY���[��ZH@��K˕M���� ��#|��ZQg5=2%ȫ���K��+�� JjC������6��g�z���{�������P�����WE�p���^������r�R1ޛ�ڮ��`:6��`� 	6�a����~ ���57�r��O�e$K�(�/F6�ff�|�����M��T�;x��M�eĦ�
������
�q?S�����A"�����l�Whq�KD�M`�&�x��ܯD��y�� ���+�������9��6��&4�g@J)��!��`u�7�c�~�VG�l���\y{��x�G�Q����Q��T���+�9QB�b��|�L�������:�Ǯ�	\2����|�7)�$��wz���+˗|GiO�+�`Zͦ+oj������9O:��MC_����˼!����Y���|:�O��j��EkEAef9^�>O���s��YpGd��r]�Yڨ��y���λ"�Lb������|��Q p���s+��x�D�V��я�"���н����g@�n�{dmE�['�#�ߡ~�ҕ�Iqf�.�g���PKY/�8���%9� �l{n��i�ĶoW�ibV�x�A �;1vņ���W����0 ���w��o˹a`i)�bDcӕNJ5��Xxi|���R�l_:"`G��b�D��+���O�Z���uh�*�E���CV��]�^u� '�{��(wi����X1\h���^�8�ìҎ�QX�$.�eWudߠ9ܷ|�=$k�w�K�X�h�&�s�*�D�8Ӂu�5,�-���"���9EbG���d���#���2nG��<��O�?����՟��5�^Q� �,��^�s�.���5����	<�W�����O���
t�dg������c�	�V}��~���ۑ(N�ps�G�)oWF���
0��nB�w}-�	H� �ԧZ�����[z��9�t\y01z�d���D��(��n��T�y�L�m���4\{CM4,��\��B�S�ܲ)HK^����?7�.M�&��G�|󣉶c��]l���
-�!�:��.�vǰ����!?,���L�&b�L]�b�2.A�*dD��	�I��/��������,¬�s�:���oB7��#��Bg�2r��vԳ�Q��@_Pg��">f�J��ʣ�����7���������l2ژ�F ��1�x�;��ɣ�m��ۜ u���� �^�X&;�3h��w$�ߞx`�e��!����s�M8�@YBIJ�PY��Ţ�s��js"E���G�02 ��RZ :ַ �w��+�	���h4%�<Wykp