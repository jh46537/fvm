��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-��߰Yr�ʋ|�^�	�Ij���1���à.}q�ꕄ����!N�s%&��v�\����� f�l�}�|�(��@�V�#�S �WKV�#2hl@��l����+����M���>��՘a��b�v,��v�Z���t<<xc�q�h�犕M�����s��`Xꑎ��8p�z��C���ǂ�N�BK�#P����F2��ջ���X��3�ɵ���}_���sG��F�e���A5/�G���^n�X����"��^�����V2��K�?4�1�LF���	b����=N\�(3�[U���|�j���O�rD�y��-�/��60R�\�!����~F�ƘS*)(Z��Qü`$i�Ja2#F��V����
I@�k�By���fq�Y�*��*��2��^
�௠8{�3��S��'1����t�$F�D>{����
��q�6�~�7G�Uc�-�S�W?%c��]�� �]"t�y:���&]B��X��r {#$~pz騻*�⤲;hT+�[�+��-�-X=$�z���<~=K�6���l��+ǧ(_�K$��"%F,ˍ/	+`�_� ���z��-��>4�E��=��4��@�M�c�^ZI���,	�Nqp�m�G�E���a� �jX_�}�嘒�c�]*��z:FK�6�06I�����% m$N�����^�x�Ơ�1D�('���ܼV6�mRF1�2�OӮ�0�v����U��w����-+t�*�׫6��T��c�ȓ�cg���g��+��0�r��H$=����i���	<O}u����Տ�Ǫ�����Ӑ�l�����s�����!�?�q��+X�$3eXj�ㄧP��;3o�I�s�$k�(Z$PF��LbZwߪ��w�],��X�O���QM��ò��O�|f9�3J|��h����`����s�L�֏�+������q���]pI�Oe񍐃�\���9�0X	�Z��_��ܩI]А��\c Eza�B1��t�攲����p��O�e����%
)Si銸e�%"H7H��X3���<�\�c�E6h���c/��8Ĺ��]?��Ǩ{Q�z��У�����t\��>X��v�G��ԈV4n�J�v������+�}j�?���Pn8��y���ܕ����e���};�[/?F�toN,ed5*�<��=� Ӈ�;,��ӻ�S��Y�|$����hP4�Ԑ�e�!��uj�ju����8��pF7�>F4����!�G`�|��A��u�����z��-[g#/�IR��(���c�Mq��V�x+H���G�zqS��6yD!VO�X�23��&'<��핽��>\a�L6�,׉����>~�f�Q]h�왢��)��.�c|�,F�T��t��H˕e%�J���*"Y�/��w� _��/��}$��S��.$A�X��ۖ/eE�e=�];�yNJ	zQ()��.I8�&�,I�v����H*�(e�!"�H���IGb�����'#:b��r&�X�Ǿ��h;M���9쟶���m/~�B�;�	L�VV�i�ikzҭQyeO*5%�zS�*u���'bZr-��Xx6����gQ�\�i�V<D�~H�7���a&�F�l^5�o_�W%{�*/a���C1�߂�H��&������ -J��C����@�mk�h�H��bI=��[[�!�%�(�r�+=��>�o�kgzgL�@�~q�{Tú,�:f���MC����������zmo^C��d�:�ڲ�0��}Z�8�8����$�UX�e���w���b�@�Bf���	��噰���?����!l�k���IX�0@�f�\���[q(���}���IY,BD�4ۯ�HQ�a$�h޳h��,&	�6Q0쌂,*䖿�Y `dKmE��p@��#�� %�Wŕ�4���#��b������m�Fʈ����*��\.�����ޥ�01K�U��Ω�*m�����Ftv	�����qJc8��r՗F ����= ��T��+����*A�ړЌ��W������
N��v��1������"���^C�j�#n���%$rDۤ(�`�y��Y]��x�>^G&��*{�̢덣>���!����6-*��/qW��}�DlSQ���m��TجNW��t�㥈���"��<�n������ ��T1#��9l�]
4�ذX�Q�l�������^��:�ȹg������w���R�Ӹ� �$�*��׉X~��7�_*7C^|0.�H� ��f���$C���W���
7�e��	�R��t�iYK�4
țoܟ#�QN0��,�.��K�.5��	����@+�#����g LpM���[@�s�S�8@���Yt�A�r"x�5���l(T�B�١k!s`.��
�=6l^I"�[�������Ku�8�Yp� ʊ�h/Y5��V������Ԇb:��,��5ї��PQ�;��
�����.?,!���h��<^6wK��)��k����y�dd��QSu��܈����������<a&Iŧ�d5Rb����FA9H��e\B.oX�$��	�AI)��v|7]7����&��O\��"}�MO��$C�xw�����J�k3��z+|s�A�5�̀�=�AӾ��5�g��Hܴ�{�j��{�����u��UC}τ������z��y�E���ɷ�,tʌ{�O%���*����pi�J*�g� ��s��i��JF��h<g�5�jLꄂz��^��s�{�p˴kQ�U�%)�?��1��w�jn(+@�zs�;ߠ�qk���?4I�v��,��z7��'�]3�ͼ�E�
u �[��u��X�.vr�tl�y�u�#`��1<��
f�[Y�$a� �i��u�P�yc�v ���ʋ6�KA�<h&p
�C,ή�#łR�"UFd'I�Tef�������--����Qa1��z4ʚ��`�U��S���Az3VXo��V��A���)t�$��	s��j���ɞ�.��/��2��&㵰
��n��#-�7Xy���㲥.�
��S�:s;[`uat�zRRe2�VW˄��_�X�mg7U��$`ZUR'�[�FO�V����Ǆ��߅��b�n� �7�o/>�P����xR�#�Ӯ=�ߙ���e-$�b���NB�&�6���p`���Ȋ��>�=�݄���w6zTs|���C��7�mj�v�� d</3��)��y$�Შ��̶-��920�d��Յ.�X�گ�]Y#���"�G>��x�/�[����PJ��g�
f�u�߫@�?W�.����K��Gq�s��tQ��	��Y{���ߖs�a�ιGgAB˔@\M����h�$lW^����������Z͛T1�r�F+��)Na]�����:�7��p뀡��xxu @A3��ȏ�؂����@Ż�m�nؔ��ߵ^;����K��
��w�`�P6e���r
kz�y��F���ر����=,-��%y,b���Ⱥ0K�PxNIu��N3j���9�,ݎ0��nz+�V��C�D=�K-�,%mү{�%��H+H\�y���g�?��aH�Φ�����vH�UE�E��j�q�2L﬏h�Utx����#:$�d�'cȰ��smQ�d�֑i�0�_����nq�W���_�"wĸ�Q�_���������@���v����|0A��sj	zp�����U׸�1�2�:��ʧU��%�n�$$k?��<�X�,rlTu?|Ynb����K���$��iI�1��,�eq!���C�H�f�j�^�����޽;*�\q�(�1MBΕ���zpК�������&6�Ô�cZ�&����"H�%��1HL�
њ|�Ze<�$D�����N�g-����@�	����bB���6�D;	uÇn��2�	��e`;���I$P*!�|J�O�w[��]��gK�R��p�^G�:񸄖�wc�Ԇ�	�L���Ԥ�b��9���s$���d��I�?��"|���O�+S��7�m�Љ
�v�q�T,Χ�)��cB@h_3~b���
�]k3��p}d*�r���EbgD�rhBt����Tep�"���R�4"�ڜ�;%�!L;��My�#�_�e�d��E=�# 8�P�ѕ�!V���=�*�`k �T<K��Ċ[��
�f׍a�."	��Rޔ��Km�T�\ӏ��guJ�w�7�P>Z���v� ;c
l��k7g^M>�w����L<�b�wrM-3��Q���3�b�7A��Ө���q� ���|��d�>��@� �D�6��_z�iB�h����R!�;!���+!w�<jB�nv0�a�dܛmv�����ч�aj̎�Ĥ���YL��H,T�8n��1��\D�2�g?�!��������ZW���V�%Op�U��4Zjg�w[��Je�6s��j�,3��P��_28�����t�Bp,6��)n���q��cd��^Ճ�_U�z�Bh�aw_�F<�&Uvk�f	�,�^�%R����P�/ԁ��n����"���4m�H�ՠ��j�s��l�^��'�h��0��"�ٚ� QE�jr���D���4ۼCA8�{��K&*o�c�[,eq,��5��5���ʣ��j�Q�M@���ܘF�M�(��(�iZ3��B&�G�D��Z�к�wB��~+S@0ڞ�w�����s�1�y�\k8y߰�D�o�z���ogn5�G��" w~Ÿ$h�\��;�W
�QL�<�7����{��Y�,n0�x;m�"�(H�I{���2<�c^a��;jD�~X�>=�Ϭ��0��r.���]gs8h���:�~n�Cw%�'��p��>7�mP��G�O��\U�r�l�j>E�䂜���Z����`�ɼ��+�%oh�p�6�����1����e�Čc���'YQ���5Q܆�o�+�*�RU��TQ��}K�/=����R>�H++O�������eۺoNΨ�h�D��=��uiS��K�Ã��j�Yy�&�j�NRYiЮ�;!�7�[�m�QU[�IC�ku���t�P���c�H��Ҏ����pR�MV�t�J����Y����1��OS��C�E�"�P7�hpE	*TQ�����	Y��k��Q���B0Q互�]mM��\N�d��y����UL0wߖ��o�3��6qa�>�mk�
C|@D|DQ6�+�-��JkB�(P^l�J�G����I�����^{��sb5�>�Ia��?T{*ZeRa-2ykPi*k<���CY���KF6$�l���b�u�������3.֓�x�o��]��
���8T�o�}^�c��� ��7w�;��ۘ��J{�B�X��+�Pc~�Iu�ä�s'��Q���������46o���Ԣ�D��������"yUՊQ~E2�b�o&�j2�̌�'2Թ����pd�y�Tu�$�[$\����h�Ƀ#���
F<���A!�uU�����1���X'E_)�{��-�����ܲ��0(q���Q\���n�L�d ��E�5�b)�~* �X�g=�D��j*H&
t �a���p]�[>��ﵬ�T�Za����@
 ϸ[��HPcwˮ���<q>�6����55j�/��{�h�c ���Z���L7��&�e-P�ޅ�B����!5㜑�p��a��ܚ�V�~�b��8d�;s���� n��*�F~�Ys>'����iO_Ţ19n��DHDZ�>T(��;g��<������>�