��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���_���W=1����o �6!�z�O�]E��"�X�	&b뼨Qt�>~fUn��b����=Q����t�̨�?ה~_�=�Q��$�͖VVZ$Ѐj���λ�y����\�Sl��cA�F���Z'���q�sn�-��'��0�.ۍ�'�,\d�Wu��K*���68�`�T�ɴ�{��T�hlQ��Eω�C�owE�}oP@����F��y����;���4}���55�TU'�� W��TݨtZ�j���%I��*3Q22�����ݬ	r3Z���\��rc��L+[Ӕ�N����
j��(x=�Fp��m���hH�+i���53��;��R�j��4�����%"��.��(`i�o�[��J:΅�*��v�2��1YPHx7�@�ǁ<Pj��ܒ�VG�w7#����0�o���kb����i��t�}�W0&�;�%Q��ҩ��s��֤M�f��Dވ������F4N7%0�-n0�=vÌQF=���g�^�2�hL� /��D��SpI�E�\��Kt`fPR���k5T�S�7�~�+�/TP��M�+��^�z8�V��O}i�Mx�ȭRm��d{�<�:��q��v � 0/�U�p����4�ScMw���\��:��C�kmT�/��7���pO��C")LDҰf�؉�(�-C�����bY6�vD�,��X~C+Q����npd��4��C'A���Y���a��Qg������T���9s=Z�>L�!}����ţZ�Y�j���x!�gHI��lB�|����R��y�9�8�Psf6J;}�xq?}����Vw����SHތ4CT-FIW��R��Ų�XZC&>fH粬5�:>���uGC��a\j����#Ӏ2� ;g��J'�:��J�l�c6��}��6o�5E�{��������f|k-�ί�����vpW>'zk��{�]/"��݊px)�Mh���@�i)�F᱋�Xr�Ɛ�A
I>�>7«�0O�u!��8E��	2�M��$q� ��y;�h�*����/��OKwL�����T�ϓ��~�d�0�q-uu���!@C+0H�AHz�=J����Y����\c�\�0�����-hD��#���C�~��+��^H:@���k�x�yU9�>zf�sr��p�x�k"���.#W9�lʾ2.�TNX��}���9��l'��z*�N�7/�}-R�1�toF�L$CfT���n�8|�nmhgN4aj��m���X�'-��a��HH¬}6Ä��Y�NfR#7;�ު@h���LqT���h���
��-����h5�K��8
%��2�&����מ�9J�'��k�,o!�v,��uU��|\h��U�<�`�"Ȉ��1�M�`:�O�9g�'���>R#8���g�ȯ�v%�d����Gh���K�a�������MDq��q��){�M��9.���M�x�G����r߯!���2&U�-W6�hHw� �����[��3���zf(ߢ��-j�/p�bU��q�>���h��Bm{��Ԉ&�@0�B�d9��khz�~�,<���Ч� ��W�"���$�C&G�Ҽ��V����ĥ�%���!����C���.=�5%�j>��<~a�r��G1��S�+�u�����}��L���rbv����B^!�N�1�[�n�@�Uxϔ�],$�e��?P[8���f,�� �1�����;oG�N�h�<�<%�RVT<*�[�����ʃ��<�c�{"���5��/ι�#h�W'�L�*(�W=�p��H-��K)��-g6"(}�ň��SL�A����?�9jC����o�l����-/:�;_��XgY���#�95��z6�T����Q�}����Plᧂ�2�����h��W���zy�ä�Q��Za�d�+2D9�NnnǩD���yTGSd�G�yh�x�����5SOC��i�
J�:r�y[>{�j)�� *��R�"�4��rʩBb@{��]΂��C����5�>1�y��Ykx���.��E<Ni��Mڰf~\�>`����@�3b�����X�W��L��!F	�!��Zq��]<��arY��g(B�ʵ؄5	�u�ۺ�L˺�N򪌀���w�s�d���-e/A���)��V����O����)���.cS����Gy��I~�:vS�Z��x��$q���U���& pS��DՅݴ�dR�l�o�U��;!]��s=tC�f���h2R�=����3��O#Ða��ᮮ�q~��
 5v�f�$��U�������m��gv�g���S���_\����;,��Gr���ȣ�D��2I�e�t�[K#��ܓ ��>�C������,q�<�̟wc�u5��S�zd�q-dw�"P�LJ7��Gùl?�e�K��#��
�|KKd]Ygw��#m�!>���h!ܗAyfF:�Kt�D���n�&���q��u��>^�4	m5R<�P#�`���V��q�v��)��+�"I#
�#'M;�������+*~����d%����=L�{.H�����0ȑ(\��/�4x����J/ه��[���m��~]?�lm��=s��6�7z3��+��#/�N��.��QgJK��]���7�$��k{v�ف�}�@j0�Ol�c�;�"��Q%~"ܛ\��Q�7�	>�E�]]��L-q�[���怠C�׉gd$��� S���>���Y�t�~4	]���!Z�����C���ÿ�88F� $�uЍn�H6!t� R8�g�+c�_��4��T(��� ���)�T��j��}2��!Z#S��4L	 S0��WW��jM������Ey0���?����{���-���-�#57'AG��H�9�Y�}��7XG�ޖ��AS�_��)h��x`�������������gמڒΰ-��Q��[�"�q�D�L�]t�-(lb{Mc���9�Jkr�u��З�6��Q8J��4���[���U#O8%D��w�$���~�Ԍ��4�%�V���}�h[��\\�{,�M��W�;�Q���'��;˽O���5�YF�r��B9�y�"AN|�[Y���e�SWj�C���ϳ�어Z��Q��#b6W��L��(�V���[�&p@�C��DO��FlHj����Ł�P�=l����v��5���`{�n���/�gCd���Oq��_"��� �a�@w;O�i��(����:�2.�L��rEB�)��7//�F�.���Gt���ƻ� 4�����	���
M	6r#�����#���V��@K��)�`���J5}��S9[�mAG��w}f�~�'�!�A�%�v64�����{��f�*|����Z�������m�y�CPك�nL}��p~��:˾<�D>b@��)���m[� -;�8O�ɺ�p�T��z�v���Mw�"��x?6*���'D�@�������cwT���h�.��zonx^���",�!���^�#�#�+����A���� ��͸��S���P�헒��q�~�V�_�}r%!���OY!�%Q�gM����G_v� ��Q| i��S�IM-x�OE��=�m��T��8>��Ř66t"�թ �H+Z�G*_�a���g��U��O�43�*f�Л��a����I��6A���R������Q����})ApO���*q�?�|�@��f��|�Y�sy��A�pQ�5�m#`�j`*d8�g~�������-.�__Ǧ�cǻX���ЕA~0p��g���!OHD�<�p�QtL�'B���n��ܳP��ڬD'��?bq��E=��G� 6>	����"F98�P\��K$�hs�^P���¸k���̊H�>7�إ_���h��%j��w� ���z.�,�ᱧ�9�MW��V�=�3AM1W`�7�z���)�rIs���:��1ګ5�?�����������*�Q���(��%sքcy�၌3r����2�)����O-�xLT��!#H���ށ��?^�=�V<�|@L��c����� e���Қ�%�e	6�9_h���|N�^�~MQ��;?	��ǌ�}|(3Ktj��������/ɟEr:t\��oE	=B����z���N7��i!�6ځ]���LB �T�6wV��O�r���&pj� /��C�?�4�'d�!��Q��l�4P �U���2|�x;׭���mf�έtM��=��-�.PP���>�ܣ)(J<������,!,�V�����ѱ�?�� l��F�t��)���fG�P���N�R��CQ4AiZl�>Ȕ2�fB������s�x�?��񴳋z
3���`�y5�Hi������r.����K��65��c�_Dhx����+��:,x�3!ߦ�ӫiK�x���0� 򤳗����9�
i/�"�� |�;+���U������ˇ���<�G4
��i&z��Ȅ�dW��,�rTj�D�ﶁ�
3 A&(��nA���խ�MF���E���7�?�9�mp�=~ulo��e8Q\fT��]m�q�iZf�i�@���ǌڕ��D�J�@�Ã�`*��WΉG��Q&��-����ㆸ�Z�;m�����ok���#�!G���5}o� ��g�ޯ3Z{!�+�����s��r���L$E
2����B��	n��ں�?]2�T ��EԡS;�7;k�YC�Z���"�4�<��.��`���(�*O�}�Y=e� ]
���i�|�6��G�j'�mS�~�Ty�0��P�f�>R?n���n����'��]��}�v4B�K����v�� �ݨvGh,B
_�!�f�����z��bAz�Q���yȬÞ}|��ls'P��K����y�S��C(~�>��"�E��Uv��t��0[m����fvU��"���+���%&L�F�?�j_�t'm��u�s2�El��j���W�O�{�7�	C��4���;,�� ÿ�����NJ� �O�����ly���`�M/�
���㞺��P�69�A�W�?�b��Y@��m_��d36ݨ;�; -�3��RG��>�)N��M�p�EH�1�1hA��O���$0���K�$����f� tO�
w�>|0\��_A�P:��h<�Y]�ـ�P�����p ��mHuaR]�E�N᥸xTz�F�~��ld���v
p5�o��#���|R�.��tF�of�F�~s�
X��W��}���Iܳ��!��_91���K�
��8'���4��^Z<��oRL���F�7f�ǉ�^|?0�3,�j�l����-�:PD���Fc4���~���0G�4_����u�u"�y��y�F����lwܤ7��&��9��i1D7p'�#�j�w�|��M�!.�[mw�A6ܿ}��}�/�p����3Ne��#s��H.*q��R�l�o�#k��\@K|��9�T��4�y�
�m_ؔ�ԉ�%uU�Rwڰ��eC_�*�����T����",4�0����i`E:B�S��L-�����?���I
$Aʓ�ٻ�1�7%������Ȥ�Q����U�B���O�m#Z�v�.�#���d��~��:p߷t��؜���G��xuaO) L��]�W��L �C Г�W��|�^��q����33X)�'������{�
$/g ��'����f$��+^��g^�&�j%��8/�bڞ��6!����,���fkEu���U9*՚X���g�7��㝺�'�ypb����
j�O�@��K������?Ʈ{!���*�*=�0��8�5��u��i'��[m�@*�h٧z����e������_~h�<�� �b:�����o��������*y�ψ�u{��~�i�w	��p_�!��oc)+$�2���<}=�S��j��E�	UJ�rH��̩��g���8֡`�'B�C���}[���C�-�Ǎ`�K�<<X�a�����,Y����^-4V4���P֦T�@� u���$����ڔ����+���d-ĂzY%��|���.G(O��#�Mvo_��t�729��f����0яGat��ǳ�
�h�^�p��#󃒹xE����?bQ��_g:R�(:y�ޒn�W�V���v��������i����6(G~�گ�3Jk��&d�0��;���/@9��itVwxj+����&T�q�UD~'0�1ն���_���q[5���DT3U ⱵM8�����k
x��͕��yn�B.�5#��a�C��Q@�%�g�6WQs +4� ��K��C��o��9��S\���?<v���id�6�8!DC���?��H��������'^�2�W��w���0��~��rJ���?W�s%k$h��u��u�r��C�{�Vd$!�E�ݤ���'3y��_hX�4w�.uۮ����U���i!�T�0n;*aϋ����������d	m�-���M?��>�����(�-��9�f��ʻ]nz�/�6��w�Xj���p`��tO<b���Sit�E�u`��O,&}Y��z��:=���!�pk�#h��+=����*2E�C��o��U�����Y�ժ
�w�_����w���_(�@9i�a�;v���f�
ˬn�튽����4�g�`�+�He~]	�!T�9n���Y�mn�ÿ�q��I�|}H�:Fχ"BPT��z!L��x��v�{��^�(�^�0���zDY�\" ���f����C!�� Ռ��+W�Ng�i駈��.x�T=Vi��)}�~i{YA��,S��AI�g�
=[�Sy��E�m<z�?�n�]B�IZ�?s+F�X�J�C'�Q����s�J��W��X0�j�g�Or�t-�c�UD�2�a!�>)3��a��jR�e��<�N��٢�i9E��0N����%Ik@P���� �D`�"=h�U>�f������_�¡��:})���?PKV��Jn��f�˰��GU�w�P^V��|]�8�Y�<J�6��.�V����i�&�L�5�q{��� ��*9S&�@�]��E�+���,���b�i�n�d^��,/vz�$�in+��Y�8Y%9�t
���ٸ�~��r���VV�ۮ�t�[$�p��gƍ��+-�$�b����\�d}L �4�7G��.;g�ehd�`
�֩�~B�
X$Y��6�^�ɜ_�����g��G|�n�rx�p�b�2qh}��O1I��1tk�l��P�_�sS�o)r�	�#l�e�x�`yYH:���a�cWV|q��(���&B"	߫]��F<٘��q����JK˩E\�D�O�����ڊ��]&��'i�:�Q;��뾥�P�u��w�8���m�_h�3�`�pyf��I�-���	\�^8&V<�:�}����Og�1��!]�y�q�+����K�ړUƩ(&�Bo�l��s�]l����InW�|�7&��c�ɏ�I�z�]���KN���o	��z���d�ޣ́�>z�ɗp���k�h'�`J�}������s"鲯Dlk�YE�!�j��M� �7�����ܖo�W�D4�5��r�{���)G)S,1��L4�����М�͋E|�ʟuv���Ȱw�r_�z�Ӳ>x�U��2���`(�xK�M�$%ߙB�0w�BE�o%��@'fU:S�t̟�=�D�$@��*|��J�鳽~tN�B�q]����"2"�G�7�CҞ� /�?�7�f������K���RŅ�>b�ή6F�M�~�k�K��?b��9�Ġ�X*�R��"2�c��4� k\ق1�l �A�<����Ď*)�ݭ�s�\\B�����<N���!4'�	����+�o���J>����VD��N� ����Õ�%�����F���f��B\nOHU���8q��[b���[�'t cU ��:�&�z�鼞^�w��'��0�Y�g����
J���"YH������c��Ɩ�z��lNt��;
6�Ɖի/:���V�}~������I��ۥ?
�c���ˎ� ��Q@����~I{�4г��r0��J�:�_M���l���7m�Y�9�hX^�I�e�.��K�m<���~|١{%�(�6�Fo��N%��ҙ¥�ZB�|d�,�C��fDT��Ә>��<!�S9�n�Ŵ`�K��N 7��+�L�;�nl������/]��hÆ����Y2���k��hZ�����^Yë!�T0�K�N���	E_��(���Ta�h�~�`%��n����}�b�5���}[�Ҧ���kG(� }��X������r��"�y�=@ ���=���vv�,k���pA��&�p�.ù��Z�$��An�E](�1���%+����@!��R�$�n�P2�a�}"�ޣ0捤MGI�!�<��6c�����o��Xz�9�3�5�As��-V6�1���r+~����0X��"�G�gsE2�LO���P�p���RL�<jD�jq@=V��'(Nb�LQ��M��z����!��,`̘�XnO���<�i�����
5�.,��=F%�L��2j{�e.�{�!5�T���.�wr��2����@� ������R�E0��e �ߌ�A%��+Ӥ�@D��j�9�{��^�`���<HR�q�|�w��UC����\ �z ,>ӒQ�4NmC�:�Q]�ө�#�s��&�p6" �b�9�X.)�H��k��R���Q_�.�K�Fݤ������9Sq��FU���Y5�U��ʹqhXv���*>~�ݮ;Zy�W��ZSv�${}E6�/�nˈ�@�䓘�=�ً7���T�7*b1n��z�o���1V�H=�V��,%������.�vr6��'i�͊�(�J޿H ��"vtBO�w�epٱ|0�\9��ř�d��v���u��e ��ݚ�YO�oZ
�'�*������/�2H4�'�j	W�bB��]	�(W����������x#�����v�
��<��Gf#בP���9�F�������|�n��8��'UC�j�([4q��.�����ԕ�����bd[���&�.	V5o�i���6��u�U	B�*"L�utiK�K�G�le@��7wG_�M��=!O�=��x���?����x���q��X�n��-,���S��/[�r��ϵ� ����]���}�O΁��	��	�>�A ����1���|�\�Hq{ ��z���)0���K0E��s�V,��`%�1)�+ ����Yd�7&@%��b���Z�ߧi@;ѥ{*�ƶ�ֆM�4����!��x/9Fم�[��exF�rsıA�}=��5z=�}�TR�B!rͯԧ)��"N.�\"��$�n]w^�j�=�#vO��qx>���&J�R�Z+o�cw������a��
I��nn3}�ܡ��9���,8���[�:^Q&H���hv'�7��v6JM�r�����1���F��š��hQM��\�Z��ϥ<�p�9�����܂\�ΦaK[=^�R�@��i�?�Bb����� %�՞�O�t�� ��p� ��-��i,|��.��$
��(�m*�O{�iU����Md��g�냦<���=xj�/����aM22xM|W]7 �	���'��[�=��V.�(z m�˫[N�"�T>����G!T5�6!��!�z�nկ�w��Z�=����w,j�3�Y�op���Y4���<o�ɺL���_��8!�{r~�yKZ}��m�Be:��6��a�g�� Q�)��ҏ��uJNh���խx��$.�S��!ot
�R9�p�O�8[����u���ԑ����}#[�7�����i��-aD��&������6(�.�Ơ��h��U�6~W۴�t��JNI�ҁ����$�S'j���ow���"$��J��<q�͔%�gƌ�I�����FX�{ԙk���i�MSH\=,��������]�eZ���=2��_�u�!SL������$���#�̈��$�5TW`!O�c_�
����D���c!{,�o&��zeP~�O���?o�WV���gc�c��P�͘�Q9z��~�|�{SvM��<^Bѩ�����n�"}c%b� ֻ��!^Z��N�H� �����]]1W�~z��,:�
��b��\����?tv{n�N�H8�qU��,8b,����YV�������%[{#<)ֆ$�(����+�Wɉ��/�?u��u��$��[)��>���c�<>3�C�q������T/�5w*�<�a�ÿ ���Vw�)���X�(�(U�V�M�΋�KU|�T�DY��V_VZ�G嬩������B�s���X�i��Аa"5� ,�Ӏ]�r���	�Z�(���t�ĦDb��u�(���p\��uo��P�A�P*�8�m�1m�قw�NY$,�o�j���V#�Q�u`�o��}D��z�yԝ���T��c�Ѓ�J�zL��Cl�ŭ����~\�������Y���?��mO$ �$�4
�ͷ8�y4�N5yh�W���V/gp3�?=�B|���5��c�a3=;!7��1V�J�d��i9BW��Y��	I�Y�b��:k���%z9���=���홋�r#��z4�{J�CT��h ��:W�$hӊPޯ�^���z=Pl"na����n�d�J��U����5�E��[���`A}T�EC'1���-Db�ٛ���	��|�4���;��l8$�O]�[L�E��)���r^��\gO
y�g��B��%�ǆh�D� dZ�^b�+���B�U$�U�:7�z����Y�(��i�ƕ8xh�>vdp�X@΂�|�/�vH�x�ɶ������jI��m���;���h��;���k���:��>,&l�jW��^�׏�����V����?'
n%����}����e�4:��.��fK+=ܢ)
�P�-����.1a3����.�3�f��qM�e��g_l�j D?�,@�܃=�<���$0}���a ����#�ԩ�n�k�BJ���04�z�y��eQt
�Z��Is==��H~��T�)�3`���;�O��DlYƗ�=���;�0
|K���[����R�G�:��׿�{�D59�UE�gέ��}����Q#��y�"-0�ٖq�V�&�,�,�.��8{VD�Q$|D�uY�����fPn`a���7͢�w�Ȕ5g�Pu����FD��y�!�f�1��eW����Xɩ��͏�O���w�)on��/T�k�R�{�/l��T���7����&0��{��8�`z�&u��,P������n$b)�k^�v¹4MM	��L�ؒK3�y�U�sU��f��svP���sp�CJ��E�x�Sy4w���'��`�tp���*��Yq� Ӓ����Ȑ~�͜wH$��$���uIq�zD�b�/���/P#��ޥ,�~�R=�ĩ�\g�� I1"eEanF�٨��^���'�����Ro`蹍��wh�Y���F�ɦJ%�f/�:�b<Ⱥ�������L�v������Ћևjx�R�jm*yP���q)��J�cH��!w8�2��K����Y�<��٧V!.F�[YY�����/G�k��lr�UD�^,ө<���V����tʔ;���*;7��.
���.��xm�g�|lH|E	�4X���4��`�	RS��"+�-�G��Zx�����a!k�ޏ怡�u���I�]��8n�t����B�+�4}�(x��#,��gҎy0�ڨ�3C���\�A}1���|��g�����M(�P�	q�;�jvu������k�Q�*�0��?Q�Sy٠�\�3 K�,O��]��M?u�Ӵ(�T�&�紓>��7U ���"%�|�^~��r��;Toi��(�*��&���W� �T����;����g�b�
�~�N��0���*�$:�P���0'o�6 i8�/�C����	�
��U�v��C�o�%�t�X��ӝ��s\a.5���x��4�#���&�TH��/�&���A�/	;a���y�ri�b���_�S�������E�j#ɧ�F���v��������7��5�f�*�������JL$9���٠Z�
7v����,�"�%��El��E��\���/���
���`nd`v�` B7-�0Y�VI��R�*�]���0�9��T0��3w�	?q�pJ(b�<�@�m�(R(���׹��K�q����c�i{�'D�Z+)`�@_���ޗ��@Q��.�N�(^�[�]��3�[ֵdٙ�`��3����u���1���r������r�sa��?��  �E���D�-�̕�ϔ��~��$b����)���:��Ƣz)s���S�OsƳ��R/^+3t�=)�qF1	�6yZ�mG���!ځ1�.=�U�m�[���=�ՙ|�Tʊ4Rm'@�{,a?��ͼ�\�>7�(YI� ��(O��vF>5��)`�̵$Z�2��Bq�6��4�	�r�(��(Jf�ӱ�zz�vBۦc6ϊ��A�����&ؗ�i���P�aK�L��U�d8낶ܠ]��Ʋ~BA�m�������ý3�T����>��_���xL�G�Dɹ�a"b���ێ���>I�v�9n:G*�Ejj��i<x>�7J�jS�K�s=��VU�D���a���^ChC�_M���a/?L���H�PW�@0J�5R1��f/��]t:�k��N��Q�qϓ��>p�����6�����$�q�9�C�z�1�~�K:�G�^w�߶]����cWTU"K��}��X�+�KT}�4�s����E��������0�b&~ ��+iz�<e�H�����m\�T@2KOY x4 ��n������"���Z�9▫%ZG����+����z�!N�Bt�=���S
toc�