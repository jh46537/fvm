��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}����=����g�'d�+[Zġ�*���?C����%�����mg��+~���zi��tyY�1��z��Hr�3��r.��!�D��xB�Aq¨8̆vP��V[��ɏ�Cv��U0��V��9�w���h�ª<<`&
�o��	�Is�#��d�����2V_�/��pE�xD��Qi[�8�J��%����K��RV�P_���#�0x��^ 3�`��S�bqr_CuC�Ә/j'ڇA������1��#
p�5eW�n���g>Y6��}j����c8�{�S���x��A�����[�Sfzl]�o�=�A�'D�h�QE���i�֧@�{\��ԦxoY­*o���!���6���|$��{��'��0w�.Bs����r(zs�U��)�ݵ�AF>s�!��Է ,�km|���Q�m��n�$��K�HX@�0�?9/s��}�UJopY�#�w�iT�?o� �pM���
H��o�+�etZ�}����wr�4��ж>a��OjR��r�˄�w3l�O�/2�1U����������خX�K���u������<ݔD��j����]i(�l�%���+[}E����E`�d������]������#p���=>�͸Ke?a�Y~�1�&]�Fa� ~m|����"I$��ǚt���4YR�(��<o{��]Ŋwq�U�P`���t�Es#��������	�)�;N���y�gё�����f��̕L�}V�M`I�3/�r�J6w�j�BO0�y� &��WBz��B	���O��vۈ�꛹���.0򯕙��Y ��q@���f��n�F�=nMY��q,?���>��Ɠ���	�x�.��{q�)0T-L�K�{�=���p�B4����`M�v�Am����3i��iT�_��!&��0g�bUVd�����(Y7P#������o��=��������>���?dd���<�~!��ַp�0ַ�����i�Nb�s�a$�H�t����!�4�&N����/���@�����L�k��Ҭ����[��B���]�9�.�ܚ�Jc㵠���*jND��(�Y���#B���F�n̫]e��D[��z߯u��)�%�t�����}_cU��5Ԑ8E�-��ngLȋ�c~tF:K�\w��9'm�4ם8}WQ�%A�K� ��8��h9`�?�/�&�'����uD��R�g�}��y�$vl�mս��g���e�CN�5�r�`�<3C��7H�	��؇�`��2�[g@�������9�V����8�81�{"G��qt)����ۊ��� B�r��C���}q)J�¼M�Ω���e�+[�i�k�C���)��"�U$Rz�������R�'c?V�B���#�1�Z����mQ{J[�� �n��^�_ +<�:x� ���ɵ_ �`+�;�s����KDj�S�ӵT�K��Π��S�i(/���u�.���+�@"��U"��[�"��'[A��;_2c�ز)y����N�7��7�·U&v�O}@�6����2^ƕ�(�4���ш�d�X
�h�}�2����S��p�;�?�Ƴ�-�嚧��uD�#��TAM.����/�.��E������d����xE��t��o/ʞN!2(��~��qHV�]y�қ޶)7ӂ��hk���QD˺¥�`�̣��ָP�`c��eȱM6��\p��]G)y�7�v(7���2@���<�������1~>59���E����B��7�b����^�.���3���IIfuh^R��M���@��Tӭ5}X�38+���Fr\uM���B�b~l� �Z�$Q��7�X����Ϗv��v�
�:G�*:;c���g��!"m�i�ؖn�X�Ɖ[�'(�ZW<�IB�y�.�J�	�����[�$��N�y��D�_m,3�6-���1���)V�ؒ�����(��	!yi?�,��EZD����a҇�{A}r_��fӠw�K���H��y�m��Aw�� ��!�v�$Gʣ'J;�8;R�@�#Pz��u��?aڂ74�-�C\�vN_���� g#��Ǝx�����Q�q��iӱyD媜3ը��!9�g-{0�ꕌ�RWo��=���6c����M��a�QNF�p���X�Ki�q!7vs#�n��Sr�Hh�#n	CS�֋��H۠����v$�A�~�$��aҩ��H-l8Oׂ|O�9�\�U�30 �M��a�NzQ+�#t6���K�b�][͘�/��V��h��:��_��&�Os����Dl(�
�@ZY!�W��Ч�h�!��!B� ���w��/���A�ݡ|��m�:�Bk׈��G�P�?���f:?p|%
�p�&�[{/L�/s�n���paS`�2���_�`{MѮ����-��^�y_E�8xc3�Hc�I��񬂾Q�7��L������R4H5d�=sT���tȐw�����ٽ��ѩ	�=��&ۻt�Ʃ_\��N! ��,u�	,9����l�טṁ����Lw���>>����?�t'֢;���p"xr0��̞Yj�G��X�L���W[�0_u9�t��+���4��m��a@ W�7�o[��&'�1WI
ȪoX��R�L`��l��h9N��~_<C��7O�@��Vk�.�����L�>����l���y�@i���A�{滥���%���.x�c�`'Z�BLi��x�}gD�֒��/ٕ�����{�I�p�@�G�.��'|�3�Ep�wiH�Z��tg�m	~X���Q!/�W�ƨ�ms5�8`��↟+��T�u��X�����d5�'Rݽ̋Ԏ�������P��8�=#�~"�;����JF�k�|9�Re�c](���I��.������+��2��jՏ
�L�on�&�� A�k�p�4��S�˶��oŏ2w�~H(=�����1��
������i|�a􎎖m'YN�*���7��!�!���z�@�W^�v
���KQ�P �r�(�b�:���E�P5<$-�}�E;_�<�;Ր�ڪ��\��`!xp��`y��o��tc��l����tv���)Gny��0c��_ Ä�j圭��/b�F%[��gר%-<g�,S���͂�:t�a3G�ȕdy|���]̳a9�L�
�<U벳?vO��)�Ů�9�����c:��y=���e�$��3�y�A�O�u���c���:T���(�~t�g�c
�Ų(/��`U���g�CAUQݱ��D�z�ر�Cs�1qtmLDzK9�^����T�ga;ي�.�#tn8�����F��A2���2'�ren����#ZS1�N%Á׆��ˋ%�`�A9:fK3V0��"S|T��w�}��h̅Dp�o�7x�AL�o���=�^E0kpe�@���_$"������E�M���XK�wM�j'���*�PV_mTPx�Ǝ�3�|�-�H���F�ɱ���{�� w0���(�!6��C��&5�"�� O�D�3>��@� Mk`�W�q�\���E��ձ�ڸN�����zWo�P�9���k���BA�����|��j���g/H���+u9���'�C���,��>���XZ�����o�5waT?7�T��i�����g�!���UZ��ES�_.:��S��pD�X�KC�FԞ�4�I~Uq(�Z7���Q��
���<�o{15U�4+�1���L� j�ecz�&j�6dK:��x��<�iV
�7��]�ҫ�e�7��H	W�s+���'Y�5�uf\!1������JB��XcW��A�e:6(>��tP���t��x�Ko�Ɵ)�[�� 2� �R��sI�γ�BU��#�!�����t�!�a�m~6<�ɓ�P�&���+\ ���Hێ���X���ҟ�E{�=�v.|A�Ԙ�mͦF�^NCub߮H�j P����켔Cqs HF�y.16�Ե#��nW-^�3��`dSo��I�ܖ�r�I7n>�C0JS��ג$��d ��@���6EH����&�LV4�5����
�$�����[>A:�{y��h�7Qt~�P��$JG��ܬ��v��T@gÊ��ۉrh��p������%�����d�̔I
���h���v輠�՚&�;��gv�8V*?������<�W(�����G�5�γsS-��C����t-We-��g"T�^���,���T1����!�5��Y��A��.,Z�/�%����� 񈀨�X����nn�sެ����M�J�k�Vg�?��xy�V�:8l��g�)j�0��P�E:��
ŏ2��[���2���՘8��{��p�}��AD��P��k�y6��i߇�]�`�v�|6�Cu�+�pHp��t�;��z9��.�pU1z/ȴ�fM'������`D��SJ���]�� )!�p���q���+��� �8������W�i�>p�9��Z�������ҹ��[8�������:�{�	՝�FB�)��%��wbOߑ�W$��t�%(�==�/9oX��i�����Ē�KF4Ϋ�f��v����nr�սc��#;�S�4�_�a���1a5z����k�����o�)[Ċ=pn;��ۨ�v0�Q,�n)��-t ��g�ڵ��ΰ�&b#��y1�uݤ@�@FmP>��oC~H��⸾N�J�5�d\�&
��K1��$7�5�[B쮍Vus��`Ύ'��n��:���n�lw���.��i|�٢���[�Z$�v�(��7J��tgk nRB�5k*~"�xMS�26`U�0��Np���c�n�F��������("S�[��w2H�i�<K�݉�J��%D2�d���1���F;�]HϬ(��Ē��c�?���P
�ջ����wPԋX�qͲ*��C��^Z�(������y�E�K�Ek�r{4Gj�m*mp��i6t����z�)�5اCNZ�K�ɛ���F�1Li)��P6�+�m�S3�?����;�4�/']�)Y;��QV�d�(6���������YV咘ok�i˱w+��������bm���E�X]; �Vo��^��ѯC�g�-G�!�"s7�oB�z�gA�&s����v�J�֠A>���s������/�X����Q�a�iP�����u��nH��5�U$�;��&'o:�$�_��Ǳ&{�������tD|�y
�C�t�>l���o1��	�gݧY���^7T�4�>��a�<��~[���y��p��q����Fծ�:Y�|/�D��SN��W���|@�~d�������l4�F�,��1VS���[���:A��7PjU~���[�E�F3(b.؇��[��[	Y�x?���ؕ.�$k��7H ҳ�q�ţJ�B��/_6���d�jIh �m���rG�v�/��ï�B)6rړ$�<��9]�q-{�E�0���R�p[G���f��C���{h (de�36,�1͔��E&QzLO$�q�� <^�ɛ���ŵ�`�J��fgX��ӭ����>9�Fۈƻw�-���C9�U0(��]Qy>}���y�4eO�j�#�9,W'�!�:�2C�ń����N2֊���$��I����s̅"1��;Uo�~��Q[��OqN�&|ɈW�(�pmB9f[E+ԗp�X�zE���v��y�\���1��*x畁&�����c�:O�G$�I��=u����4��k���{�Kp�<Z�J��7�l��:���G�%KM̿>�pbO��b�֩G�[q��	ϞL�^��Z�?*xAd��À��yM����k0n�v����	����b~��#�w����kJ�һ���1�vڟp=ʷ"�Ri����� �ߐ%���|%䗫�?�_8jx%\�:�o�g�*�@Zm�HQ�����a�e���친����g�./	V���@�t]@�w��@A9`1��1'����V;�'�طO��&Dp�1M8r4���[���t� �q��M[:LFV
�Z�(`���#C���L�C�~q���M������b�D`C[&�$Q-�P��=�/]����~�[a��ě�>�5��K E�4TH#v>DZ�����vXP�DQ&�4�U[�Ԙ!�"�-qhX��R�����s��7�6d����i��\���y݌g!�q ��2��7C��o�/
Ԝ��m�#�h��D �-�f�4]NR�B������FEM$�P�mH����j�D6����=|1kf�>���1�tI���Sv��1f�pᶟ�!i�����	�/ǤA����
T��r�R��;{���Ϣ2�uU���>s��~���R��j�L�8�G�Ɯr)�n���]~�^g�	�K������k��tH�C8�8��v��A��irA�ܤ�Ӹ�b�r�cG4���Q�⽺嵇��j��� P?doY����劫7v�����Oe �di��Fy�@1p�+��.Rb���n8�� ���2�^^~u��xD�b.�dO|B����B�gd�� MJ������	��$�)
KI�����������kPS�bN|Φ��T�/�5�UxG�1�s[��s�Jt<^9��O76�|7�|v8�r�_�>P �/w�-�����M�� \ �����@�5�Z6���� �!���.�N=3"��A7پ������=x�q�,L| ��N�U��|��q}�j���̽x��#��D��<�U{=I$��9Y�3�׿]�ۚ��G3��X�I�nRA�����E�5��0w�!2 ?��W?7�7��I��T�
���|0�O��}L]LU���>l��]�/�\0
 �|����*6뗂��.��#�AN��Vx�m��ܳ�T>�Cy�����&��Rg`}r�0����?i�g"�A���{�)֪j���ȖR��	�=���eE�59l��îiC'��A�3T��B����U8G̪�)u����'��c�;\g%d���L]��1֚uX<w|�f�ԃ�b�Z�#f����^ġ9}dTɤ?ɵ���^�[S"<���xЗ�=�	�h���<F0+I:�\����C*eS���2&č`SĖ�e�S������.��d|��S7�w��S� �As���ieɱv���q�0�-��%�nE�k�-��-�o�A��H��1��+��@*�n���o&w7�����^��{ґ�k�D$+e?Y��JX�lMu���9�Iζ�_�M5�A�pp�����ċ��M��6�7�IDbĤ60w:&.{˞[��cV�xD���f�'q��Ͽr����P�=[��m+qL�R��4�������Hj�=z��"����~{�6���"��$2�8�:��yy�#>�:U�/N��j�i�%�?�TO��x�Ǘj<#�fg�/�)[u�5����r�9�xb!��'W0Y�Ju����1�ےGg`�K�����N��7I�h��8#ko0��̠֗�w��̭����0\;�Q�l�P�U���Q�0��%c/�v��= �?�_Y�)S��� ���u��Swz범�&,�]�l�ȯ�3��
O��W�X+Y��z[db{IU��VT�Ղ�� y(г{i��)9�n��2lh�2KAYQ�:�9���Wo95�d|J8�L(�[�ݯ���ɖ�d2�uv��K
���A�X�eᾘ�Գ��go�1C�U�iakw)P��*��Q6��2g{��u��p������V
pD�3y�C?o��Kv7�A��F`�->�[p�z��:n��ε���W���2�W�~}��IYS�-)R�n���=JK�y��K��l���L��K��ˀ�����'�w�i0RR#�j��Q��.����������d1�ѳ�a�niv�U��?�dk��NR�!�H^�*V:=$ZvOO���T`�kf�NQp�qcPb4�h�=�c��P�01������'��ϴ�X�瘙˶%�~n��'�^b���t�9�Yg�.�8�v�f�	f�v��}5�N����㦥��bE��@v�$=���
&p����s�-����*���Q��)����t���i"q�m�����'.�A�q:�K�Eqj�Y"��e�\���8��mߕn�֑�_��'�J�.�
p�Xъ���ܙ^�k�c5����"���ɼ��9r_��'�-�:�����t���n�|.~FhsѰ{v];�K�P�RΟZ����5ɭ�T�"ұL�WXH�K\+�%m���R3˧��pf} �f(�O`^��7��ű�IC�z5��T�JyrZ�jF�������􅓤5�$��꠸��a� 7蘌��\�<���N2�l ���Vp���X/��
D:`���O���]���'�,���q���Q ��e�O�S��v�*�J�}:�h}a(�J�yY5|����*��"��O��_ �}޸jX���p�n΍	v�e��d7 �D��)-��G$��Z%���4�7U�aV,�9��ڡ��ۺƥ&���Tb��S>f���R�3������6�I�M��S�|%_��H/(}����ص���~��hQ���Jo M̚GI����|��G��;�6s7on���~�y�Tu	�(8�5'y|�y 0�Bs�z�\^�o,FWRL߂���[���w��|��]��¦�+��ٝDz�N�$t2����O�d�9�M�r��&E�������gC����V^{z��M��c��>W9N[	�5�}�c�n�6q�	G�$��i���t���r�.� i�'����A�R�a�p-I���%� q�]o��g��E�	�R<�l��9bI��0�����$T@�xF���L�ܤ�O���X�U�O��ɖ��Ӧ�8�W�m��0"�'/�-����}Gܯ�:�k�Lָ~�ȧ�H*�>����?	��٬t���g�4B<^�X�ִ����	؂Zѽ��=�,�0N�m�Q�BjĖ���
���u�|�U󏸢��)7��$�js�t����/ U2�1Ð�"6xy&}�� �sX�'�7 �]5�����nӘӗ���yd�T0�W4�r��̆�R0{.���rP;9tS}�����ut��+I>ҟNu�oJ|�B����l��@�$��r��,n�'�	hEL�f6�zAI�`㒭;&*�-�	��z�>��B�������c������暞1GȤ��f�Pp�T��^h�j� C����Y���e����r̸NŪ�=�9|�frx��YEe��00�O0�X�W
�Г�XH�y6���F)S���])�� kb���Co�n	9
W���QA�"�����]�߆�a����<�L�,,��#]�b�����M��V��DX30&z"ׄ�Ufxzq�-c1�.�,6x5i�V�����j�V�>�*)G�̽�ܘ�F���������g��$�T�����yN�ѫW�h9%*�4W�i�-�ÈjM�b�}��\��448G�����tB�C����J�4��4@hί�V� �ņ�[�Z���G��ʤ��R��P��e'�y����FW�;�%쟽	n��� �V���� ��O�gWt��=��~`�����?�á^����y�ĝr]�Q��N�{�(�w19�Y���,�Қ�)�;|\G8�y���4�l���M"���J�ɉ��!�5�@�^hn�ٖ�I�����LҜ�,�>�-� z���}ȳ���f*�r<e�{�-���℥��C��-�^��|�����|S��p-5�[�Y]����)kQDޝ�@�-��ζ��m�4��m0�)D�fB��gv,]3/V�ʹ:]&��>�q+�Ȑ����4J4��:?�e3*
��)��]@�����FV,<�֪���4;����!��n\��:�͑�/��\�=���wr9�d��� ��+F:��8����e���{�7E��}>[
کo������hL^q)7)g#�&ZPK:��'���I���Z���6�bcǰt�z�A�/�b0�0��V\v���7�s��o;%`����:���A�p��eC�R���`Q�����u�N��9ƴ�q����4����<��jz�a��XCE�P�/�Ҙ�Kw���a�;��%W! ��H����Ֆ7�V�. �~9w@X��ײ�Q��Y4��L�V���3lr���0�M!K_��Qnl:��G6��@Cb������_JW^r�ؼ^z�#����;����%��n$pi�J�01�an�7��l���p`殾wI_6R�RL�[�V}I�>
�7,ӈR;N7\n�,���Uh[	�jޏ)���EB4C��K�d� �iwaa����{o`��}����!���33"�gz7���н$Zנ��i��Eh#�_���9?��Ч��&����ia�P�)��z�QÇ�s�AXx�!t��D����0�zy�A�Cx�=�2�3��V��ڱ#P+*��,�H]g�`8��!*U�@�ZG�Eп{�z�{0�����
���v��*3�8l ΃�B�@-Wv�K�(���ggzH��� ~���&� T� =F�o�D���� Ny!T������g:�9�.�A]��m-ڱ�$���>��G}���2
_�bɒ�Y���H�{����:�Z%�a;��6��.�
�V�
��A���;����6Ŧ{̴I�M(#z�^�N����\��ć�)/Y
})٥'�B緮<>e�o0'c'N�%I 	,/�醣n��� ��� �멚�U2������i�N�y&C5sW+N�Ch|��K��;~�fF8�� �E	�=ӣu�sb�?�n���\؃�;�g
ҭ�ON"zM��LE�O����1��$��,��/qlI�:T��_4����3�_"�E�)?v���y�H�P4�C�j��� ']��!�����1:���E�R��"u�vX�P�b�T|�I�3#*u�W/�7ѩ0��z�m