��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\Z�;�j�A�D���£�d����2���(�C�rY��K��!�}�mU�K�6�( _��B�7�$���zY��۲�69� �Ǩ���G^:��Z�Y|CCҖp����x�#;����"�B��؇��tyɄ�=/ZIqG�W~�M�0Є�p��=�rȧvE#1�BK��S��{Y5+U�k�`�n�%1M4�]X�`M�W�z�9�/iG��b�ɾ��4��@�H���H����$1�s������9Q�D�E��zO���K�Oմ�Ic&)֞F<n\5��+u��蟫�La�^�@x[�\a� �>`��")��fG���б\���j������r=�V�:�A�gw~����#�ݚS�X��iA��#��`��%�Mj���^����&Z��7�G���N^�Y`V\cK=�c+�%U����ٔrH�}L�K�Q�}���Lu�"ޜ$�
���^K@��m	�ފ�gw�<m�u4j\^nh{BF��4��4�?���F�we��	�}�k��(0��:�ȏ4tă�]��v�;�)#��'���6��z�TK��fhS�w�z�����̘��#qY��n��>�q;�������\Sw��K9�K��p�}1�j�C�������0�U�%YP��5�PH���Lm�p�6��#5F���97��Y�]�a�ߗ}#�Un|n�h��txuݙ�fCt��n,"��\c+3�NX�oC7_�?*,E:Mx8��i�T>
]xIr�V&n�p�e�<>&?-Yi#"��°��z�CLX���� ֡Kʹ�d�������bݺ�sx��o��O~"�A_������$�RMr+�y�%j�aW��?K*3�͎�R|��O�l��2�r�c��6J�v�^�jXC�'�k��SI�؀t��(��gd���������[��3���0W;�֦~�,�ׯD��'%v�Ġ͟��z�}�a챣����΢_o~ao,���?h�wm-�����Q5C�(͊�( h��]0#�¸��c�N0H}l���iG��_�:�E���uX�ƥJ�6_y���s��rUe�;#�62p����P�,�ƅ��?��|��FDEi�(̣�l	o�v�uק���-d:�ZP��e�~m�W�2����V�a�whBD�󽁑V����{+�w��`�u��=�`�R��N7����+����]V,�1��Lw��������H�i,�ѕ�{w�s�d<�����X�ك��=�{n�h�dd*rƅH:� ��d�#��rP�+�
c>�V�/��/^N f0�W��j&譯ӎ��(�&��I�}bWdj��}2D�@��.����M��5���2�(���F+�:�s�v�u���i������<���O�pw*Ĕ�;jA�����I��?d65�S�DR˹�!P[�0h�~���$U�\2�;�W��j��(;{t��C�BTPd�7�l�Z�t)��V)��Q�n����"6����ݑDi8��B}rh��ӧ�'7�"�W�Z���I��/K���jx�*��@�E�G]]�y�m���l@l �'	��7o:g/;�EѺ����L�H��$#j :0�E�p����d�ﭺ��e�v�9�H��6�Vf �آ��ﰌ��=e�\��ͿF*Ц�ӋRP]�ň��>�<	Mw���Q�1:ĺ�L��U4J�HO9$����TY�'N�z�P2s�M��7��Z��[B������b�8���U�W��[�򞎢UcO��t�<m�]�r���(�q���-Y��x����

R��@#����v�SL��]R���Xf#��. .��m��S��'u�](+�^��2�GӍ���U�9�-hSየ�X67!,?]���Yd'f���E"�`TR�ހ��Z���
���=����D�|-��5�+V܊w�Yf�V�t{ׁ�˸ת��N}1����lmYyi��G�~��/��P�U*�Z��Q����`=	s��S�R$	s$���#�J	E�k<��r�~�셍��e�^��Aro�6hud<CD�fD ;C���_����ӎ(�?�k���h�;��'jx�am������vv#�=~�70���2_K�ٌ�ե��n��7C�V�����e��(��b�����~�Ԅ���^�v�-��u��T_HO0^ׇ�F��*��$fL��\�ۗ�ا�Q����)T��k�q��hG��t�_	sB>c�4O9j��	g+]�-3+و�3���:�$gE���#ڥ��]�ͻ�F�6��B;T��\���Ɯ��I<�(�-R>�~�����j%qGɳIjy�@h�'Qxܗ	��"�/X�"i���5���3I����r;���Ir�̈́`�V�<��N`Ͽ<�8X��M$��!����ㄨ���:e2���\};�����_��Hz\��IQg�����4���.�U=+$yR�]��Z���]}<o?:TN	rŇGK����IF�Z��␡�#�r��i2v�tVepS���� �X1����#"r��s�M�$O!]ji޺ݼGѳ
W@�����F��K�]�|���/ �_S�S.�#�6m�%�E)S�i���e<�3�3���i�r0��h�3osB4�����?!��KTZ��<�9�a�&�_�Kǉ�r����6�M�T;�΀K<�S���>�
�
���IZ� ��S!�/�ʌ�ď�
?!��Ü}�S(�P���	�5�2l�5������M�G�&����Q�{!��a��.*A@��_�ö����J����M�{��؍R!V�P`:���|�|��MH[��x�c�(��q��l�����r0�G34����3u$4��B
����!`.��6����#�5��.�|WeΫ�r3vݔ��كӡKf�aE��FHQ-/�'�P'"'�=6�:�XH�>��`ˏSJ���O�/>j�"Q-����g\9���˥X8����wn�.��������5|t+��m�PA���}߃��n'	��(����L��#5�	��@|
���7$#��Z[�#j����M�9�!#�� h�u������!. j���Q;S��s��]�z�(aW6�x���׫������x��T�3W�����b��֌ξbl�����6�@���׏�o�j'���a+�����;�R�cx*Z�A9ٔ��U�Vmu5�ڔ�8{�K�<�艧�㡍v�u�]lf�,>����:�!��Gd=vzn�8������P�X�����;�޵d.�n����q��b�ދ��<T=�c���
ߞ����f�X���g�Hm��� ����?��o�g�pZ������z�揕�����\ye�u�E=��+縉d��3b��ފ0������#h@��m��)ͅf��r��DU3Z�~����G�	Q�Qk�fB,���1�>�{.�y{^�m9\lS�I׳H����A�gR�u.<�C�fYo�>w��m\�b���U����3��	Ru�{eQ���$��$����,�/k6ܠ��gv8έ�3�%�׻ͫ�Gm�O\?+�B��:�PH��t�WV�飃���c-��g��Mp�פ9�qqU�Wک*+�W��C�8W�D.�C>3IMX�}D�[���I���P�h'�ԡ	�Kb�A;�+�8t��ڰk�<�~�[H�<������~xo�G�'�ܥӵ#Bl��W�lI�����&����xѺ��aP�	v���W�r���9��u�e��Lq�b�DGj%F����G�w{�'6��ȷ��Z�t{�	��&�\^!	_��Ϙ�(>�=�Z9ЇN)$v~}h�Pw��jn5�2�#��o7r��Qk�j~�e��:�a�#}!��j-�n�bW�U$�g�r�I+�[�T@��E�f0��-��������&r�H���2��ՠ}�%P���7��u��"�W?��'�>/�I?nC&[�Ð$/b������}�MC`r��%+P%�3�,9��"�ĕXz�J7_�rP0�!ӄ�7a��T��:t_?m^�m���սj4T��rh?�;{[�N��[�����*�$9#�:/Fz���py.�<��#�^�I) ��q Ҡ�z�CĖ*Owړ��\�c����\�x���� �[F�J;s�+��Fb�/g��x|��2��N��Uct{��.E*�Z���4>bEq#QMP�#���^�BI��͑���m��<7x��8 ^��0 >M·HI�}��1w�K��6��!h�S�I)�*Z\*��b������;yC���Kz��J��-:P,4��ǜc^YҲ�v��+����>��6X�0A̪Q��Oc:�+s6{��;*��+)�T	q��(�D��T�1�&̮7�p��� ����G��><������θ WL�x�'.H#
L�̧�8YE�����/5��`�bvD�l~��ȹ����5G)L1W
�l�ɗ�nV�����i�Qi7�N(�����.�Le�+<N�J]c�O\g��#執8-&2q�F�雝Y�9�H�3�Q�S�����h��I�9�;���P7����2l,�8$��l@A��@��'P�/9�d�h��F,�5c����O�Y+l^�B ���Pp�Tq5h/GJk�ޫ	Fx��u�P,����ȭ�R��2�E��)��5H�6����$ ��}=����m�yh��ߓ�_�o��[����9-��U�/B���(K��X:j�x00|�!V��Pǟ="�rFl� w*�����Џ! Mҭ�l`���u�7�h"���phF��*c�86���AՖ�s��z!u�Hy9�
��%������5��w�s�y'�]Z}K��\�i�kճ���(�­��.������/�nTS�9��������*
�T�#�Q�+������7Yo������L�| ���^�t~�t{��Eh�<�>��;W����}m�B�qM�t<ԃK�@�N9ػc�A����	.j���2�aeH�k�m�9�[L��,G�)Cc	�N�h e�):��;�mє�n�4*����fl%�z�ƏM���/X|����Qa�0�ջ㐨u�V��X�灼~F����(�'�Ykd=����?���z��x�����1�z��&]b�=!`�;1츦m:����c_F�ێr�g�~�ϋNO*��n�0DqM�~�j7T�*D�����܂���k�߷�h�q��I���f�}i����`�q�ϔ��{����N���X��Ǉvm����mh� a_��32�
>[ӗ\(qp��=��P�{&vɮa�A��/l�!��I߫�Y�.������N�6k3܂�ai9S��[}~�_���_ѷ�������>�4�}���,�2�C�G,a����U~�Zq6> �u�X���e8�HT��;nmҬ����*�o��(��@��K���i{t��q�(�L)����/��j[.�(����p���d�:H��<)*?"�-�֪���!���tuh1�ȉ�o�cl�5�A�M�-f)L�\:}���T&q�^�����su�s��?w	$ug3͸z,��ޥ�>�+�>s(��ʶ���4�e��ؤ͜]���G_8G�/�e�
�g��#�)<��$ wℬ=�Èm;kQ	nzv��-�W1D :�Ad�*]�{<K�\�eU���L�cj �Mʶ[	E�-|7�E��������c��@([2��Ō�{M��7v"��v�yJ�HF�}�V���ͭ�k�y}�$v_��[YI���>�Qί���0R�l���]ms�]m�L��g{p8&M��*ᵍ�H S$B<����.�F��5�F�g#�R����2d*P�8x��+�f�H]���y��4����*ee:��Y�΂	���Q�q�:��è�؍��al~B[���L�+��z�>=�|��Z*���G�j����Um%z��m�>odovT���ˮ���b���xd�\�F2x�kf�"�� x����yp�F������+%� q�a"�.�Vr��wD����_$�f*[\C��@������5�]������}D����*Gӽ��L�b���r%P;�� hv��-�b5�48^E��mZ*`���p}�U5؋[����(F���h}�W�.q�@� ض!���~e�����ރ1�3UzxL$�V�8�A���>�IV$��^����h���]��>��W~�霽�{�沘p�?j�����2�� ���A��t���Ņ�0>�&%}��@�$�"(AK���$�|$����e{�FW�AH9q�,.�G-�P��7��-�I@Oc���9
�4��VH��!����/A~�#J�U�"p��S�o��+>����;������=�*_�F|U3�����\�N��w�w8����U.��5�=�?8SJ�ޔ9�O�!u�Vg��sF\Ý9�I`��sbu�i����>�?�e�!C���[��u�e�i�"�c}�%�>gp�y߾�� ;�б�����vU*�W�ނ���|C5�Gɷ�j���1��b8j:�Z�#��