��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�9zrv��^�t��|솟<���+Wz��ke�q;�"��������U9�:�	L��������27�u�Z>y۾�j �|W~��-܉�L!+�!X�%%�¹%[O��U��UA�^�n�v�)e��c���v��o6ٖFX�E��SN�M�8�SC�}� 8���8,M����{4
K���#�4�k}��#�.Qԟ��Ԧ�"�_6�>uo��2����~ �L3�b�q���g�~�G	�� N�l�<��}�|�XN7|� ��Y:%��(��6S!@~Q�UC��~�6�3�"!��v���,q�|��T���>\����-������@b���\�F jm�
z��?�����5�yBG�_t���h� ����1<��|8��v5��4*D�*͚�L�an?aYԦ��ؚhJq<ݜ|\u����r�SK��&�/lW�hH�7��B�p����ҩDH�l	e�u��+��m2w��ݷ�Gpρ�2e��`qnNNV�6F��cQ�F���en����{j��p� r�uR(�mܙ�9�k�3�v���a��XQq65�A���ۣN�ֹ�>�b��:�t�}�>�O^%<Bݬ�t��O�Y���~�F�ay�bt!^W]'(�	dC"������᭬��Y�8a�(t��������^I��JLh�̀E�6�l�X�U:@���:��*L<}E���ɴn�*�KRe2h.q��{�u��ί����0#��R�t$�&Ս�f{]w��^)�Y;�I�U�$�==k��c��Gn�u!i�K? m�ea�3��߱�KJ2ME�8��-(=k�`��J컏��z�1�`@�����1n�����e���Ej?�/.A;X��K1��F�[(s�p\EQ/3�v�������|�S3�ny������r���a�G�����#�����]�O�-t��Ҝ�7�( hW�P-}(9�Ó�I��ֱY��Wv��U��TQT��c�7�W>f�!kp� '9�$����2���1��b��(�r ��]�!i��n�Fr�$K��K��fu	�#7U��3�^{���=�j��오�}ȿ�I|a�[���U��NN��i��.���O�U�!�U��}�~)�Ğ̚׳d�Ey�̮��aX�)�H�*fO,o�+{�5��N�ff��n<��B\.w��df1�#�~8'�����P}iD�߰����Ɲ���b˂I��	8�>W�@a-�+.l��l扶���w+tB%Y2��>��i�X���'_�tL$zf�xz�B��c6G�zF��k����&@(pX���"{ezOe������=�ŉ�-����@���!~�`[�xHF`?d!����9�`fwɴm�{�϶�?褐�A���Y���_0�5��YY�p��fX�aACq�%B��<����ì�S�I&3�ހ��3udL��Q�2:��� B��{ �� 
���ަ�y}?�sP�lgq%����������	�G1�woY���+�Q��H�W��[�'z�]NZ�KĢr�G/��KZ��_�>�_���(h�C ��L��vI�;����v;���ɮ��]��X�!����2,�^��'���9t��8����9���j��@�l�@MK��9�m:����`�/��9.�y�{=�'�)��{v�N�T
|���IANd+	���[��A6m�sD�&.�d�IbL�I��Z+�"�u��0a��)����7�y1%i157ɴ�G�J��&e�et����uy�X<�:IJ��0��u�I���ĴI�X{�[�)y���XVhưW�r�'�#�ƿ�H���潐U��DW���PAm��ָN8���3v�N)1�{;�m�ᖏA:�A�<��G����6;;�r�;�t�e8s�x�[T=�w����̸Ms����`�z����h��M^����l�0h$@�{���Y�``���5��ݒ�zG�vPu �q�qr��Ke�},>��晟Y��/��45JޫqX<�=MXL*�̈l���{n��$L�� R,�5�4�L��n?Gv�:�-�?�G��]�6}�������V��ө�-ع.ZBߘ�v.=Z�]���� f-�	�e%Z��r���%�]�8�V��������wL�ɇ@w���;U�j�cN��@:����`R�v�xH�ٜ��s�,�f�C���w~N�r�~��I����=�SF�u.���fu>���\��xZ#�Ĥ����^�cs�@JPYw�rk��(��[q��l��[$g��P�,��!���\�
�~D�����{����8�,��x��V��(Oǈ��@�ͫ��#UWH%K>����G���6���sm}+�M/�'"!@.�����t��/WkZ�|	������rHf�p���+��U���[�����{�.r�ɹ������8c+c�����YeVeO�by ���R��g/^�q����AX�m�����sA:l���T���w�,�4K������^�0�#�ʪ?
���jѻm�l5�~��'̠}���^�����#k ����Sq��	 iK���-�yP�/43og��^ʴ�F�� ܪ/J���f�	B`2^�N�ӗ���/�N�Ӧ~5ĚN�
��< �WH����,��N��9�H�wP�������*��!���I�cx�2����u����`� �P~N��y}9�?����8��YJi��57kkFH��]|+fi��ŭ������hG�j��H^����g'�������;j�ot��gu*=��r���FL�v@��Y���l�	��� ���
5m��-8^H5�12j�YE�\�c�mM7�>��,ᥙ�R����'g)�V���/�x盬ɗ
���}'߁-ڰ��7g�������8)*Q��r�����:��j�ϟk�{b�H��u��:��g܉O���V-��)����	�^�����W_}�<:���w���z.^g��������0͍C�:w0/�u����,�-��T��A����������e�}K��\��n<���f��#��J������ٝ������E�٬�@`� ��J2�%sŮא����iUӀU�Яf5f�p�5�Fd��O(��HgC� e���җ��ɀ�}��ى���@H���m��Rj�l���=�P}��}��ЖvS-����bW+�c�w�@�ph�σ
��c�8�!Y;3����|�ӑH������64��S�����F�z։)��(��̏v����̏@��O����%��HӐz^�Gf9�7C��؍���z�v@�-)6Q�Xk1�Ytd�Ϸ�>j�z��%��2�,�i���� ���j�:;��D�Xt�q,�<�E����)��M��'�Ze�<��v�>����4����b���������v�)�vb�D��Ƀ���L'$`�D����^��W�vL+�~�]^�[u���:q� ��@M��KS���w��]�o�jD�UG@�T�}\@3��J��\.�]f_'{��!�^(5�V�EMְxU]Թ�c�5L����%HiȽ�:�c�C���\��Y��L �G~�6�����V���0�O"W��.[��s]>"�	��y��%�������k��{���
��"0�����\7����
s7?��Nփo��X����I��\�[���=�V2	Hy!�Y�.h&�,�:�N���"M~���eIǌ#=����U{.2I�E����1���2���I����R2[U��8��<����ږ� vsG�Y���8r�(�K`�GC^�8	��ς�q�ԁ"�?�
 ��-��%���A���w��D��IO��T��ھ�{p8ѹ�w*ĶO�2�����ZolM��v�b��\�w�DR������_^����@��fV��M���MrP�^�+�/�X�=�
+sjo�N����J�1�0l�w�&B}ti��i#���z�,Aݲ%5��ץC�x 1�[��ОH%FJcPM�L�?Ak)G���+ގO���v!����n/|�G����'Kj�ĉ����Ε�])�ϒ��`�eS��ۃ�����,���˲�j8��d]���+��2��"^>z%�����hS����у�1w,D�-s �������KXs$�]��x��R�Z���a	�j׻]EN���G,�n��=�^:Cɒ��@*<�0	�,ڰ�&D���> b�������Qlpi��z!SǇt���d��Lq�ZB�vm�1�DB�F����}	�.��z5�{�"͏z��G� i��ζy��ʗ^-6�2g�T�P/S'�L��oB�3o��|�l䗯�`R���M:Bb�y¨~����M��w�T�WB���I�F�� ���*
f���[Z�"������N3G<%Lھ���L�8}E"��/D���bL�Y�� %)�(�d�:@ه=��-&�t�r�J��4��X�S�hK�����'�c�@��?D7AI�P��K<o��,�p�����/��1�.��+@�.O�������b��>���5��.������5J�n�܌ &�{#S�w
�7ɠ�;�ًR��!�@����� �Pd�4���囪��vO�Ba�AUE�����f?��6�)_ ���s��.Q���0F�O_8.t�WJ�gE��4HCdtMn�n܆5�x_�,86�@jBC���ny9Pi�4	C6.
�mkʭLw�w9��5����$&�.�S0���""�����R�P�)\�}���jR���x�'�C%q'<���ȲE�urWx3����֘��&=��d��K	�G-��C�lU��Y����i���{6n0��2r�l�x��[��+]̝�j3�����e<�$�o� (�UP��x�"�N�K��%��>���ϟ�*/tK=���I�ӁT�*�wA��(M����Ћ��?��K�N|����P��%P49�Wۂ��&&除c�����dX����N�-G���׹���m�K���9��av�z-�x�u�M���'�c#iB���+]����In��_�����U�VF�o���ձ�Q��io��j��?1�����F�]ZM*�Y��jn���q0&���.����4�S�u_���-�*i'AB<yŪ��FO-�bHj~�(RӦ�o�L���@-�y���#��w��ڟ������\@����K}]���[����R=̹J����o[?�.�h�(�be�7���$���]G){� ��3���c7xE}���:�#����o�'�:["Y;l߄��W�Bi��K�=_V'�	]���H�rY�3<jE,+q� {�5�f���Ϲ�J���P@o� �e�&���bϩ�m<�S.�BB@`��3t�|l	0�)�F��dt�Iކ�?�R�j�����;���g�	�{`�
���)X��J�0�#z�uN�%ѷU�����z����!e�Waaa �B0};�nc����v�p����P\��3J��l,dx��卭��p�=Ǭ����qj�8��f_���	��Ԓs���K�([J碵�W�K����_/V��$��:W-�8��Nzߋ�T�9&a��GW|H���hI�*�7��������ҽ�xp��7P�S-���̧B;kZ*�@��ڢ��j3���Z��6�7�����e��G��x��7I~Dz<�ɸ`p�6Y�	�T*Б[�3��T��λaR<�_,�6��SY���r����Ųq�N����\�,��T�$��Z]d��t6N(v/PՔ��L��$r����Bnb��D����jF!=��Ǿ<�]o���|��W��b������\^	<�;��7,���^E=�&�)�d�K�93O^��pj9�1�X�����f����]��i��s����.