��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�{���dʂ�V(��p���ha'nc��c���4�ft*=���-,���&��i���[=���p�%/�S��	�����l+&�I΁UD|Ă2]�18ɹ8�<�\��#g��X��
�۷B�n���P �HKeF��uy����@a�,�p~�m,�j\I� E�T���yNð�+b���2��,ǅ�����Za��e���k�ƭ�"DJ�h�Y�$dy�&��tdzH�ĿA=�*�ѣ"mw�غ�?���]0̧�f%6����73����XL昆 �t�;��Ni�(�&�Z����߮$�b��ØؙO�cjR�Xk6�T�K���O�� w��3���(LV>�YoM�(�Z�ܾW>x�]�V��I�b�;����^����q�	F�>U�k�����v��v6���g��i�E\��zfE�o.��[\F( g e��=�� 7f��p����̭��#x����._@
�u}��g:�l�ԱK��Z9���F΃8�}z3��w)����*B���];|z��Q�gK�F�Y�BN�v�J*s�uQ��l[�� �}DI���5 vzR��A��C�dz��DC�{��YaI���a����*<���D;��x�v���q�I7L��a�P&��7g�����w�t}Ra0G�>�l+�Xe&�YxDO� ����+�о+�m������"dA���	��?L��	A�_���������S�rS?�o�=��oΦ�CH���;<��?�O{���5"7}��|������i!�ԓ.z���_��;".�TV=�E@�P��4#�^X�,�6��ƅ[8��53�o^y ��K ���m���g�cz�2��u�� 0�N{�\�ԒSG��\�y�H��������(ɩ�@�Mp��]�*"�	��ZZ��9TF+��A<��p���S�༦%rl4�Y�����s�p���/�w�e�O�B�� �@
���Bhjuz֬��5?ٰPj�U�3*|a臼���kx�y0ߢ:������dN�`�
>|*B���G�f�Y���~�xF';>k��ECQ��E>����.n?�ux��i���x]����{��)v�e�Jc
�ʺ�Lό�M�����w2)��q��j����ߓٙ��a/sk�c�_6�6��@���@M�c�������-}�n거׃�0�1�{Z`y0��3U�M`p}�W��v�]���2�w��{MM�gCw�Q`��C$�7�cB�Ѝ��;,Y����@�P7���(f��bL5�;Kg�s�ǝ�<0U��0�"`�
~<�"������yq�0o}��F����e�De��A�i��T�<,���G����l���$m&)���ս��Wxb5t$�邚�l�_P�3�U���,݂�^u�s��&0��e��JL��E-�bv�����������nB,�b9�K�ḍ&����2���~�!��\�����:l���`�p�H��e�uO�i�V&����|��*s��Ό�h@�뾚�>YF�p�zl�nz�c2���y�+�U�=[BG�,Nt��};����� �^O�P�4a yv��;�0�Z�8� � :���@\DT'��J
�B�p�"�$C� J:����}�Py[�� u�_,p��1��a߇�y)�+�B[G��:h�s  o|]�������8̶|��1�-�Ӟ_O������d�h�L�� ���'��Q�cϟE_8{P#D�L���Ak��g��*h�ѩ���#j��pSNC�'uV��=#���b^ҟ
�I����jR�����'Þ������O���U���`J�9GqX%9��CfeyU�;>� +�i���N����mgyT].�Ppw=Z��S��݁������S�Gs8��O!\J��lfvy������4|U���O��.c�A��WG�*Y|"3�f�������r�]�̰�)�db`�nj�wQp�[��i��ˌ�#hG����;xf5V�N_��]���:��m��+u���(�����F��y�=+;r��i��c��C��2��e���6�	�d:u[G	�S��v��J���GH����Td)r�ن��*��yy�D��Q�Tu���+�8�|E�#���L���il8N$�aO��/���i����-�4�ڶ1�=ll�li�H��%�q޵1�r>�2�N�Ď�Цi���gH;S��a�4­$�+��D7S�1u5Ӡ�̵�᝞��eG� Ōx;���'���N��3<*37F�s�̴�u(���Њ���$i�R��(3�^V����Uu��ԧ��ɤG&�RB�0D��AM9���4+�g���e����!Ԡ	�aãp�4��UO��`��n� ��Y�%)܁렸�ߒ����_�op�2WX����|��)@�Ա[�����i�b�o'�/��5U#������}�ƶ�Y�d���h�5"�%��jAE�t�|>	�~����c:'�ECR�Y(�Bjݏ�/���
�; ��u���U�xfڲ�P���da`����m[��)��Q�+פz�O�r�*8R�lj��#9���^{���¬�J,�~�HTTY�����%re�����o�`Qsی���j��V+y.��LǶ���p�{��V�dL��v>x��j��>?�������=S����]�6}} *2W[K a�_����#�j�T��^[�S=�p��+�ftǮB�"����D���Ρ;�?L����T�[�eG�� 6n�ԥ�8ʩ{�־�%�����$R�+f��E�,ť$Bp��θ��o���C�I��߳�[��?/��)�9(5c���Է������ �!��KcׄH�g�,y,��U��g�~�w�}�(�Ūr��x�%�{ &#�9΂l�#p��;\E�h��]�4�s�[(;aT�	iE+��|����f���]?��e�UzBMi(��hl�#~/t���4@���U{���I���W�4$�A�>�ٴjd~�$TA�9 9�}C|m����*?{����֝�XRiO-�I�n.`R������@�k-�`4����8�x/
���+���5/�.��P�?V�;����������Nɻ�m@e�ea|�b��]	v��x�\���\kƳ�7<e�0/b�ɳ*u�,�w��!7����E�W��
���3�b-�2���w�E��B�K�y�ݟ����´�<��(��o�v#�!X�I��x�+�xǂ���I��yp^����6��[�ur \2N��w�K�=��
\ğ2pf�΂���.�Ը&�V=T'<)�=�t�FX-����3�-7���6��'��}y���(���l��D����2W��^����O��e���
tfV/�<^�ʊ��&!�٠Ƥ��ߴ��r�ܚ7y�ox���K�>�r�������~!>��@B�x�(@`�98���/�'+Oz�/��1�ِ��5a�A�_�p�O9"�=��?c�F�駍o9lw|%i���Ҭ��RR��	#��-�
�wv�f��|���4'�V����i4�:A��0�s�-)Qy���`��.�j��z�軘@�#����m�p�>��L��U����mQ��H����P���k��d��� �*!L;���9�Vц��PU�W�`�8 Q��wtgɓ"Y�},$^}2X����]�`p�6Nz	�j;)S
xMu�㞕Dm��3I�F(��Y`��5	\u�'W�1U�iY�R^c�nC֝6y'�{(#l4$<4���/]K��퀋P��#�����du�������+mK����aЁF����)#��#���5�l`#o�Yu�4X��=������]0� * �d)��/H�@�A��;�5�o���}�`�~@S��ώݜ�f�G������NB?��_^���E2�g��I��e�s�@�����Z�U?YL��}0��Y0vD"z��G��;w���W�Ɋ��[��_z#GY�-�����P].����<F?ëkd�����Z�F��ȼβ�t^u�-���W�(�	j�$":���^�*Ao��04�;^���5�fn�<��E�m.��&"4T�xi9�B���{� �[L��|���8�ἂ�T6�v�~ٙO<�}B��ft��B��R)��4��%�|3�ɴ����$h�m�FB�)1Z��g�J4Ԡ#qx$d�7�i�4 «����J蓑�?���W.!A�Y��/���ٕR
P��U�raFOz��m����A�YT��K����U�5;$
ņewڥ��\@���dM�dG�\�.���w����JG)��&��e8	�[چ6K���8�!�5�
�NE�H a9`Sn�ّ��-��#�����m�bu�z5=��*��N�#=�2HGw1����X��]��ɱ%�e�[�(!Pr�I�4P 
���O��nrY뚈��oV�WA�P�E���q+X��w�R�e�|��o�<IBoS:+��s�F��E�]��7If���B��=�I9C�v�%�w�$�Q�Jk�4Ж��p��)��F� ]�БO
[!8����l�zCO[+9�D+׌�,���x�Y7s��X�femO� � ,*�?�%b���r��PJ�FU�%�h��i�O�d�YZV{i����n�&7:A2�Dk��v"{|0�VO�y�죬hi�3�rs�_w�w���&��DOQb�Z;&4����-�̘�� �&��?�u�L�G����ۀ[����������V|P݋h���3�ѼK�S1���Q�Q��	��$�A�C�G���<���$�o;'w)����@��T�M�9��W:����U5"�v�m�iK�w&�)���r=3&/��ӣi��U�NnB�H
%1!�gj���"+\%�H,��u(���o�`k2� n{�׀�-�ą/����
;+X���>��<���Łk��V�g�<��m��8؍�sTN.����8RK��c�We��WJ����g_:�|7�ʞd	����$��|ac^s��w��/����Z>�JF�q�{<�H��5���d��޾*���Q:	��gcLЅ�ԭ�T	*�ߏ"���b�Z��c��q����l���s�ɻ����[>L�`q�N�6�t6]y���l��<i4��k�q5Ϳ�Gq��0u� ��a�R��֟�wO�ቤ�	j�;sh?Uq���