// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JKMyHWFFkPZDaciUA2OR1TUwoqqqbGw/e4ejqsDh6x5OAYUnXhU2hqGqisZEA0yJ
Iu1WKOj9HSQYGqU8RDCNYzvxnA+OuI24MiHWjm5V/05qhkDz1B3iMQvKwzVIDL1O
dHQoIry5ZVteUppg3bPjdl6z5MlVHlQNUx/7hNklovU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26448)
VB8gb0E2aeXupQj4yynQpFKHxr95Tf901UjrcG+veu7KopE59/unsWYACqTyj5u6
1e2qyDGt4NKGK+TZneIHamH/TBKWn8QJKZTlS7O2hhD6oiOv6mh6aVXVvmvU/ysH
fPQKFTpAhM9uRxrp5NxkkrfE05lmV2k+OhraVDwtsPT+7aM4hGYOvrrrUasN2f/F
TEfPu3xTsX28tylWlCjokQnbUtGMOUcMQ3yL/WxY5ugBOJLtV+MODd2Ihvg2Rl5V
ssLFX4lA1zrJuiaR1Yo4strRvlzI0sy2hvEZRk3Vuz5RDXx0L9XQm0Wm5WoDn+lu
7wtGHA9pQps2t2zlK8zJH5lPOBMXgliSpTeFv/l6dZyfCqSSmGQ6tBV8UwQNaZQl
ZO6fisBVr5lyl2+Czr5zbBnGrA2uWjUJB6hJtOb6WoRVhtzF+RIGkl3lc7bUgesT
Vc6s6XF9c26eSMG7O6KpyWyhZ3DVmkWvlisaMrenhwFc5c9994AKIfBGR3mq1wlr
ylE5vgtKKPkGovhtxhR1bTiVzo0v/MlIZIvGDv1BcGv/WhvGHKWTA3u+XgVEQNff
Jp19CGhKqJW68FuqER0T1bq1daG7WThzHRffLARSPN7bHsDf/utrfkOFdXv307WJ
RnUZHpBdR3kKbZh+NrK8ddCxx8wq4TjeGOS07iTnyRnqV5KfsO8lNH98cFR00MV+
9CKSTsu5f1SxpuIJOOs2mSU0NQ7TO34zN/ghL5jWGI2w3vg6/ej3VCQfAfKEeqgE
HBQmG4yzuFlnctCVOPOsrE6RGgZeA01CPxeVnsGNUl5VTZ7yc/d7iZ4rkGAapOqb
nJb14QEQ6s+jxRgBzLtJhpQFpgrkGGD6NhHRD9KZClj7QTNn45AzffyXtgM3X+8g
mEw66We9q/OunL2Mh5XhwB6E+JxbS9mQ2uEpAoLu6j5GHLF0ko22u8TpR2TfIj9Y
2s+EiZKLm2GpOcWk+LI1iNLhTzxuVANYMocbRKUDZaIPT+kxPOWXrSD94gtoFyjm
uBbPebMMVsRD+QUpu+K9W34+IVzXMHsJD7GCupsgJGGa9Y0iOcY/q4oGu6bbegzP
pEGkoeP6Gp8ZozuHnXPzQhp3iJPrQaYSedN4QLeBFgRxUFeDQwMpi+YrgciwFr2h
spyK8GQOC15HyqTxoNzgIeW+WhiJMFkb1CyM0Gb2pmCEbIoabo1kXXXLhYJaQN9F
2RAKJN0T/ncyIf1GCUIg5SHnloEJPbBXsZrygzlaFjd6WHNO2AkOZ7pwsR3iYP9r
w36TfIAwKImtATeb4EpZlUdYY0gteHNqcC3u3k9O3/Jy39DRU3DeapChsn3ZuzpE
1UcuIjEr5omMrP92WMZinbfEBnoYWAzqwBc11nWTFi2n9k27J0CzasFi18z9yAVM
gYk0ciqaPZsMsBtUiGY/geNv4nM5sB51vWzMgyfybilpjK1vstYv17epCqJORv1J
XgoL8/yvui2VrsK3ThxELv/2Aro4pryEmbj+h/3gIgJWhwVVtqd1pydgbmq901c4
My3KQj+V1VEqJRTyhXrAfc2OW58bQzShv6E6WfCu4/ZR4jCPPhHhIw4Unh0+RRkH
GsLvlcZWG1P82S3P6AlCFsPpNr+LVFFDiE2ObO4pHvvktk97W3+tH3oCjGeXOapn
oEDi5o9KDYjuoceBG0WWlbS+2NYVWldwmB7e0iB0xefVGoxDKTczvXtPXV9l+AOy
Ok8XnQSV1+J/5RQNKs80el+2Fsmw7ZU2CEczvChOdKWfAQndm5lcw00ur1P5brS3
JjAtopF5mwHgVg37BCWqX/TNRoFIu+UebFRo4zBvbRKsSqmQd0d+3bfHLainGjAu
if4s9CQNoRqwGELY9eG4KHJw66dG86n++BHjKHXLqNrZ3dXM0Enxg+zE/ymVV/cM
gtEf223+d1uCZwTY4WV3v5rBox/TioiwmH8K8PK0cWg2lB7xi30jNltvPJz4vPsI
fOHrYNB6ZyOk2gTbX7c3lRqwXLZ4d6/Wxc/bLfmYXmZPq2ewZR8oV+MuOSWttNWu
hCIdFCKXTMxRJA1/Ge2SoxlGAru0oqyJGqDXrc9saIYJTFknsrmE99AymjYW6k/D
l4CQOk7sCjJC3AUdl1A8YLdhXFFvhi94ENpSCs2+bwScWuynST1BZk23blOdt9x7
54x/tyNUV365/9EafvISBTbko56kuNyzRxd9Q1x5bH8IgajP/3+ArHXRnruQaNm7
O9NLuIHAoiJJ50pFL2pixSYRDY94/+Surkj+rlt+DpRVo0MoL01qHJjmo5HGBQnB
kjHR660yOtIUHIq4wVLq7B/dvG9YuBgIV//czsOwp8VtX1q6gNAZDOfPQ8D0Xl1c
peU5hQ+6kw8cQv54AJFLl69Ghw53EQZZcL2622apIoV16LuGpesNSkwwAE9tNQcN
OMjIKtXImLQF3lqT8PlsPGOmPT8OgRQxixGOJoacx4BVqGCAMJmev2TfS9xxtbkN
3Ir6wwgJRq1dFGY++DHJrEFqqwaD4zmPsMLeI2jA+vgmJiuJcl0WbrxT2mrNycn0
xqaPVjYMeGpzHSjdAlWrFMcw+A88q9cpexleStjMYwtxcAN72nU1IOQqR3VFuw2s
vHNNfIr2Ots4KC3IwJQ86/rqmApnS6DSfq+ybBd90oft6Lw5Z9uKhhK7XAat+ZSj
NuNHgHE78YjFOFqi0PSzoKtpS6JnckSJnVolhiS15OtuiaPdCtYcUprlDeaHa6hX
wdwo3Ujtqz5KgOD8963gESGY0FYbKdFHthcI7rMweltFXMKjTpjfSXFnT7uBvdRM
AxHPZsZy/RPm9RrvS68WictcF2NeKUipO1DN+lrBL7x2sMu/K4ztCVA8UaCkZqOR
zNlBTLqn6MP0T+1ZIgQb67NJpz3Jtk9IK8p8sEUywLBYlAHcV3Q94nhgCfE+TnAr
CPG+xWUXmmyuBCxxoa2o94+t0266FyXsHPjf8GB9/7n1Ug4z2ZYDz1bl8wg7vemi
cGi0tbpT7aF12j+iDALMDpXUO5EGeSE3vlwdXdfGw9Ijdk0F2DyGQSzzbGIQ8KE0
sR4CiUMd4Kdf4WDz16AbDYReUTQateWpKdeEsi4ZAPtowpWrts2epxKDdZxXwCFb
y7N7/Ru+k+8u/191URNn51crBYsLa8p0A7gbQFrx4cpo0QtxbqlH0qug5SDC2Y4K
8B7t63KlIdF/AIJOCEKROV4jUYUWJ1/eElJuWSRPp1drTlVAaQp+mRpx0SOrLaIG
7l5duf0GqAorsYfOqL2aHKzLBvaeCXGdPcqZQG7fdWDc/GsrYhnJAlpVB15IQSrn
k/2xoJ5IKixfO9UyfDjiNcNtoBqBXqLr5d5225muQKURUUhvimCGUVuzHOZ+k2u5
UVePq4vLtiAhH6vnDgjNmyF3vtHd1JHLFWqUmnMaDKIw6qd6dGftVAt3mgz5s4ZL
gmIF2s2/g2OljuAmTLf2/ll3KIlJUQRFrWSPzEcBJ949kRkT+9LV4uJEhH0R+Jw6
ztnotmjLSHGxVHciUhEYHOw+D6ct+HtkhUar7IXSjUnI3KkL2De7eNWyO0t+JWOx
dVzQpZgBomUnkEhVtkvn+B78mk1rMFlXrzwp5Au3i0mXHLWIB5r0JKvADo7Il/GL
nDQ/vcgeIWnLgJFOtzetFIJ5QCGI1yDE0UayP6XpKZxdxyngz+L9GxENJDi4s9Xw
FMiUzu4GujdkS6fEkOch0du7Szab3HZdP398CeTYmxX0lo3DP3ZsT1yh0Q+B5Do6
8xorHCEh6OMCPNg9vMzalyYHGZW0c0vjEMdTg5qwVP28FsPtYSH6TBDVPGfIeK6f
ygsmULJtwVnxCLFCEoreXPqpDM3pWsJziELZ48WriA3S2kgWmhbK0iiKydPXHBgW
0DvY9HHrJb4ZxwXxVSiQS27qsmmDr8TmHs8vgydsscbo//xb6hAKS5YnO+Qp5Jbd
ApgbGikj7wP1F+6J0DjuGYj/7RahO0n+5LiTIa2aqRDKapLrlfxXIEAxMN48/Rxg
Nj8LThqN8UiiteVmMKlAtIhZdtefiEZXWLLMi/kaDmMgOxlOTbDINErW2M8CuwSH
43xLsmlPofmaC/WzpqFYgiu1eFyxMO4tdMRpR9CM/X4LFC1uj3JmBAx/jLN6LoLR
oadok3ikRtxw2u+eqW9Z7mYTz0EJmr1EP76TDcOJ13nar5TSmOKOb/9fykYXkcO7
8WoBHo3fowEUrNJav0e2LO7ZnRSjm40IZxM57+mPJmwy92xukSGvXCmOoqRozosQ
Z+Qo4AMYcQOUEu/F0PFqsoqZyjpaXgDZ3iXXEaH4ovUzZ0ukb/xodXq3O8epAwkc
tht1HMP1e2bL22HZAkMlh5SogSaow44CnT69LYuqm4LOgJzHmh2wbGj+zUrKuYdE
XTEEqpe1rJhGKAdmtx/PLDsyIRq5GLTt2xgtyTospSKaZhbCCMijD7n8uLlMwkZx
SxP26oGGCQw+KJ1xeBgd4ab9X4Q+Qu4aNuYSfxRx0uhqeXy4tq/syGqii/alnZ+t
Iwtysl/O6aP2E8dviVi2hRDLtIlrd81Yk/HHbIg6kjcX45pbinyTBYBTDm/eQqJG
05T14whAVmfnQYO8yk0/OzfV7AsHSaMnvCeioaH1bjpPICUIf3+pbTUIPoMqibrE
aDAXvS3nHTZkmN4AMXh1S7EH2c/X/I2cNxbqMW9MWk1hOnFQRN68ZJpqTrKpNazV
NDXybvF0s2nRXEIbjSorRxrxg3bNM/g3ID+960nLN+1McI+FAmq21bUg7CyafSpF
ZHKXAgLFW29k12vXBlHWMV/NoAeV7vUBkV5hpmGZfnpzfmOfauivVVTHKS2mSypO
EnaHIfB7DY83OaEnF7PSLhKPxNaCtD4OPJgw6w5jvGL7RezwkEY6vYn2kIYLSe4y
eoVl9NZl/wDtq5GIO9fU447PJSLcxPBmAyaCH5u0GrvSZ0aSdPoW+bhqHx+Vn/O8
pooabO+gQl0G27XPT/+2nmLIpbXHqb/l2GK4CnAxSBkcgVOO4t/3ss9TlPTT7kKw
mOSaT5XF8zZwkxmEdV3j66by+a252LjnusJOjHf/RjdbYOQ2gEobcsnpfRVmUvqG
SdEDh2V6l1VjQxn9flpD4LRLg1aGygrhKMgbFE4JN8GORyuSnijSRJQmfDEATBF6
a8X0yNKN09l844kx+E7gLEZ0HsNOuOes8ozuPD9WDQCPiWbPYj1cwAo/8S3aQWkF
RvZCFSosUSapmM4RzBuwjdjWDTzEfZUGnqKojkec7hqDkgxMrAuGgFrfUNnNDJCR
6Zi39AueDpLeRc5nXI9tuHJvLvDRgH5DaxdwpX67ADUOURVwRaEKHYbVsPm6kuZu
HUPnqtJ9NCtEZ2FTwoBEzAJ2xJKrif/S+DEPQ7wOy2vh9Xxfu49JZsbwF2sHjBTy
9MitYqZdUGfsh/w6HpOwSZmfxoDNtCh3z1m0iJo/cu8pgAN7UgC6kYQy1B3G6BuH
wu/dwkqExOeE+E255DYHYu0a8c2EUkxgj41l5deppS+IiMjb02PA/cSQEMPhvr+o
474iJgUB9nZZQFvD133Pl4TrUBL7wm91uJ4f+yPNevIOZCnnv+SO/La6zkwwXs4i
rMM+V9b/UDHVOdAYLkixZ557jzUTBhFtjbYHfkWrlzfE7mrIeVqXk9WiWyKh0y7w
Ay1vBvRG6fvAukBBTfAenohK9nw+33sHM47RfQbssxuwz/CXCb1eyB+cb4M/2AX8
hNZ4GaaBwbtYfciGrYxZipIElHNd2Loj5ddvSUnDvxJtFcOmo7OUnkcb8oVzjAvM
jsuZxRuh0k4r+V8qw6ye26eRvQIWnRhObri4EPOd/P3Se0tsUSaffUHDAw3DTU9H
ISp9s63zHqdPwkGyLhluwQkv0GTQjrTiz2ultbYgo2KnrzWMa25RAXdd7raNmRL6
hqbyWLPyeZuho2oFnKFEjXLeI1TUaQw/rrcBvW3JAK1gm0FvecX6w57NmVKe7EpY
hKaeRGSQqia2XKEoqmz2nJxjddn9DMs07FLo9Np/yyLrwGbEXui51nK1Y7Q9ULQy
NbihdJo10Hs3LxakZMOLBwezkdBp+463U+sJ7RQC/aivs8Y+Ylhtf/5/VEoCrAe1
U5t9O2kWuZC6A1CnWgH0JnyVDDpPKx+gUNxC9FaYyBs2RJI7AKuQoxkluuUCv4PD
0IrPnbje1HwdQeaytAzHeKzd2vetcJ+goqn5wWHb9W2LBClVNHwJ71jfdHz8/wBi
4dlQhAUOM96/LynwAJuRdGu+AmCi9/djzL8/nF3tpe7dZVt5cdHQe25rlz/77FLh
RfCxvDlICmoomgsowRtnVIgdyuA7d31QNWz+fPKbIUbxGDSOgaqr4AgDVWD73Q2B
jOycLMmZQ2pStd+HqpcwkVg/aqTMsQmXRw25BBlvjaV6OLDpHWZfwScv10O6DYOF
oiCqzq4RIWv+wucznChXYhKiF2MtW7Fb1Mslnb68j0Zfs3D5vpCNAfpRiOh+Rz8N
tSmWml4BxW0nbG+vQQh7/0NfHRY2DEG4k4KqI0e0wo+xsIBjtb6QzGroWCO88rbg
m6iVuGNw0l+GCCRXDL7LGqGR7dpzUNV5FmIKLLQqzJxE0OWTJwESPIb9F98OIh4Z
AWGguhD/nYeLjg2QslfiNb7M6VfjtVSA8ut+t2T64/K0cWINJcPBfpM1r7W9iK7X
ehLF0CY33d92U24ME5bXFsGOLo7wQis4f3jL+wvRO3NktjV9sfcUIZW5WOVnJ05X
9faY1fGzW73YCgjHJYpolUf7rKt3ENiWFhRHiab5WhsO23TdM9yjVjT4uhDrrNtg
j2nCnqbIWwEfDOgF0Jf5hcUzKhOh8LSJKuMn5ivSmqdNj5qwTsuIGyMt+KJvFqHo
VJkdAN59TYczi2MavFjf9BopmPG8yyxhefzR3zu75CzShE1uyP4hYWLvzc3b+LMv
2viAE9JgKS4opQSgIA2XkkO3OhuzO6LXz/Bxr5G4vL3t7I7SkAgsyR2lV9ygMOJu
Q++0haVXXr/KE9PXgl3q30ZmreTpAsV1hGl9uBsbVsjtoRl3szgzHxhyj8BrwS3q
yk7KoVKN949iEdkXWz7kO4DHTGZ7OKHixOiYrFt8Mvfxu3maQicZqwIDzd7gpBlW
GbqbXmw8hdpkPSD8t+18+7KgNkLxtyd3wqCgeWpAk27NvOHSn7fO2pz+YmPflGHZ
RR4sK2cHrRASYmvXCaYIfcjy9lK4XuqVMHtfIcL4lTTj2icCuZHG+Apt4MNpAdk1
LpqQb5SAjV6IRaKJaZ2ohH0nsSDJ0T+74pQsn3dONEtVQoGG+K5frYB5q03kgF4T
bN7euzSSXLyZrt1AAW/SGsOkmxFc7537/wBJ7FvwO704wfkUgiFiv84Up7WgOx5s
t/Y1Fwowg80SZlwT401Dq5IkgD+wOt2wWBhE+w426fe1+eMMq8uynpBf8DV/bTYk
un9fW21YcjhYE99q5V8XEfdozTFSgv9Vt06x6Lk9GJ7P6qKZiIWeXxfee/8IFrRR
DrBWQ7CSERYM3WP92F6aY00NuQUmUayf4My5jVD0AYiHJzfwx6ZSpC0KkY7qw+r5
2Ep6XnFvshcRLxOPmPLOQUrw7yXsa2yovHJr5f8JhGQN5fom06aMui3NN8vH2xG6
ULhLMGhTs+/jb9/gN0BRLD3ikmYyaKUzgtciTfPP5VwvLLv6No61k2deE3JRaWff
W1sBm6jvcAIx+czAwP+Ke0cGlNwnIhXpcn5NZsd/+Eegtx2isMAgGvzP2KODG71e
LRG8mAIH76skNCQdBXCGzWRCJaynhXAu3oM+Se2lM5UL2STBooucXwbdsSGOUXOx
4iVNFh2B/F4MAGqQRu2C1BTMc9cc+bODvbOQOFKfdacmu+/kHDhFODigml584E7Y
x8rhmqaTjy2bKQ5/RCzbhFs9JTnIGz4blEMcp1kP+JsVuDwKNzkNwmIoFPt9YJSA
MyCiRwiWpy3C9RlN7hJ1YQViURb281rST9gajhwAoK32DQcVcKU/oOooqezyQpJx
d4Vh5zcWSBJEcBeUMMlq2TZShPGT8bMvD+HLvww+kc1bFf40EOjgci50iK1o6/T+
TRqB7l0tBHL1zuTQ5ZfIlTk3UW9+8IxgbnOoVuaqRuiYaVVjyDhhVMX3LljzU8aY
Qzt5jRkqIAueQ59MiOVCnfTab+qxFyGBeXE7DodLXtI1eG9iRH7IQm8OsaYB33O2
kg1KtoRhQuK7dnBdgXTP7AhsCPMh0HSxeBYA90hWN9c6X/Idlb241SrRO5r9mD0Y
F7IyxaDfmlj9Jh2ELoF/5ZN6EtVxt1B+z1h+5eJketnKZvLUNxChP19aquRgLy98
6/sYifDMG/ruBX+C/bsAPe5rVEg5z3sQ6ssRZvdGjx8UlxjmcZLX6IUbmVhCCYGM
eRmGbVLxx2DYJSF0aGJKjR4fvGayy6qTSI8aRRmM3XCDgLa1nQKoDeBYazJl++jk
QFKugkmK2v4SvHy8Vv1czjXX9+twTrpDZi8wZdcqsvT6YJnRizA/KjLBM8aPgg9L
hRKbdwbcSlGmTqu1c3cgBDDAEutl1WRJNYsTCHpR3jYsEynDGkqbDGuX/Zh/BhAS
wbaYJP6jPGhJ9FM/2PS/7go3lbXs6Vppj5RfpRshpj3RYQVIE2PELNpJbttMLN9G
Bd+jYHSRHu40vTfDVIHfUC1O/YLeYT6TCSb9K7k9vdOI+voh/MeZxgjwREqDsXLZ
uMKayNzbZKIjro/q9Bd2AXzMF/563WFMZN6jFI8X1sUfJqoNxEfs9K9uTr6BYcJP
LvKgkV462nsg6WAyTClVKQOa5kuMZRtGz/5/wn0VOZy6BkADR0mGD2/g19K8O4n6
ZKKoKXv4m+OOP4Vafgqf0N73L3NxzSYmo431ZS9TxkvvBfh5mUNMImGOXpKnn5Be
82IhCo08JNA+8smi3x9VKBblnEfhnwftvJDvzB0wCuZdb0B+C5brJLj2BaZNzSkA
sfNuQRfq1VB5a2jv1DLQrBhPWT5WjtQvEuw0NV2ZUIOf7MnkD++7R0fTJuKOQlMt
5znZRtcw/aHLQ/Zn858VhGKe7qX63oOTIHz+gAdEnPrQKbF9DISyTsFEHlOhR6xq
sNiey1R+pgx9vxCFyKXLQB9AoSWm74bxNhs9cQ/I1Rl8k82F3rDDxWLcd2DMW/A0
fEFtFuS0nK6x8JtR6jPcobzm1ekK08Y0Yi0ECVqxLLXXUemGQFDg0bqxUyq9q/0l
V7oDGkh7Azdjt6x+TD9EiA17lyrIf9JZv6nOI7EvmmroKqo8ZxlDKOp8z2SIRjmE
kOYQHCmlkAFQV4puV/qNV+IBgP1V3GYEztIGkq2H3o3WDOYV6HIiVUyKGqtM26+Y
Q2U0gayNp1o303HnGteBls2g9+mhvOdiD4sTLH8T7dVIC04fhNrtqEKWADAc2C12
ypZnNaCM/K81ek7h3UmZ1r4932WIpz8d+nQEXNaLDuCmAYf+MdMRsS7CeSouo4v/
Qr1g2BVPTuS6IWYiiDfFBBXPxgV9acS1jPitbVtz/N2jpyvJE7IIKzvKYi+qnz5h
IxWQzauosMJcKCg9/NuqOmw3rKEkUFL+K+QJeezzV0e9uHWQHBy1k0OdPib5se4f
Pno57y5LdtWjQaXiuCgl1waa4q1I5CycUhc8R5MPy3pXNqEI0TCi9An7m7Nj7ZVO
K6XvcPUvcFjE5jw1H4BMWoTHeu8VdsNz013oGFvRYrcoeAF+g2/NLRRjpRbK+QTa
PB51gFuQdCPMRwIkd8z9GfyoJucoZAtZqURL0mnuV+oVR35WOX8VfOLfpGqqNv72
PkiOK8O0HcQP7LXGk1snUxr5CGBfHaLCyww/dPlYFAdd1YF12jpOfU/w/G5YM4+r
rJv7uE3LHrAoEMcgqHIjKuvX/Y+3NAW91NnVQ5LfZaAxs8V0wvRxdJck05XpbatK
FIN2u/AG6ExNlYic8Gd09lBCrraUrASesfTmL+XCtq4dtGTxDeuvX2lPbRbSz8/2
giaJJZ9bQY1cIJF9CyzJRPIcQrTsxR118Mu81Ze2h56WizPtJd1UJz3b4DRL4KPV
KlsPBn0E7MHIfVEkEkvtKeBsWJ5cYR50bh7yTO7HQQGj9TnfmqO89CaiXnPn8zfC
mu5gvDpcVsVOVfu7CDjdKlOXKKIL/61LEuLKrwL9xN1/HucMmWGHLjjnqxoCKwRo
5RAjqnh20ItOpLJRsed4OIZh0SgteMy+6trMNqN3wIBJ7ojSK59YLDJRdZelX3JW
pCdZFVrsxlePVkD2KqeOSig98i0VG+2h3qyXI/8PfKYIdjHhvoGC7I1D+cHdVS/6
UDAlV5BjdpaT8J/L+4dV+f/GxQJV+UUUCdINu5V1C36uqtztUDIFPDV0vkaZt0Gl
dwTDzgHVkrSeFbta61gCmhcW0DMl6jw+nxwQgc1QxpJCN0j9ITAhsOXyFsFHuj9z
M8mQ25nux0T2ERe2fJMsxmfSlw4xKxTsDthtofpfDWeWs6e6NxeMMUxbJNjELlho
OGgOZiyWz2Yo5XG4SaCS1sqMkIkNT096kmWJZQ8VMss/I2jVnuRBp2l7ZOAXNYzY
x/tu/KR5U6929KgIfF1pm94armyXeiNsS7/eAwfiWW2j+qPIrERcdUIIS5vxCA92
O2AF0SpjyehCm0pnPviQqMH2Ioh74UOo97PTBrEnO/FrFFuihF8xe0YVvu6ygSqT
hqepmTqIcEVkOfjJcxjjabQltbMWylgxOOOVcOpEotJILxkOCz2v8WkscHDJY9hq
s1Wx9xXpdYbFrYL3MvjypIAhnc5VXshiHIJdx6mbQgU+JStlEHOLdHcMGiNK4pwQ
i/XIBYzE4lQ2dGS+gMq1DlZT3qmfoBhp08cq+iSw4lrYKouRH4vaDQpCywnF9P7K
S/e8EvWQsABe56kZwxtPjWeAj9SBK8m4wrAvqqpZnx8XqJavwzaEUKqo4wXI2j+X
xLG2CMu5ySTtTqVZqmXHXSmMfsyOJbCnrEKTFmUVhtyc56diHQ9Si4zsdLUfhWnI
5BJe2RV9RcVfiBmSHEDz//f+89eTQ/izdxz6KEQe7k2xsxUZYVuxintPjNQNCdV/
3NvLCbbnWvLXRQFhvPaczZCn6T6Nm1QhMZYfJec+m/ttvMWj1oCCUNi9jnAeTNtp
TRboE9/X3hS1HW5/hfWFajz8Lw9xzRkHFzio0qiZRQadtag1OWpVPItKnYB8St07
KttAfrnY7VsAfPneJLJxnTfZ/7Lou09Yb3f5WiffKRy2XjopRIiRFKHmfQnMtvf9
KHz5bvpK+j6K+NGouhDlYZr7RGkL6whhXBL4zPH8py03MGh4hUeH3dDUTZuge+Az
buslNI2otndUT0ARzUJt8j6wFRpgJ3EjrREyDS/S1bkVGdXueVpH/iA70S6fLKTA
9sqeC078hViSqXiYn7EPOEb/o0740dgGR8jLkUvWaKTM+upWqhrRrqBzj6H5QObU
4tj62ZWtyMXxYx196edsNbTPj9PFVO387Gj7sZVlIA1jjMwwwY61aTZ2ftPWCUxs
uT96fxS8ev09EwI/HsEQxcjsyz9+LNR4cDj3r+tmUecu0Xgnbzuxbe8rfHEnTqh2
hr8H+Imr38jdPMmdEpNo3YKM69zij53mECv+rarMCuZbJb4clvSEe938dn3c1hsb
UaKmazZSf4zHbhN5t+n9mRTU22jn/XuY5iA581JcAN7JeGcJbfYXRVZkY1kG2fba
+JiweUHRI6HfIDZbO4enQDiHxpxuWJ5Jv/DLTQp0kGScIcwy/upxF6F9FM31oD6P
C+6an77TwoVznq7OZc6eyq3ICrJiNLZVIrO5tHrMU8NSKGy/v30ko7QnqQrAftkE
hNg9efLTkq31TYztpNJg6e+NvM424KCAEO3+hj0u0+TlfKEoSaonquB/OiGgNI7/
ejc3NsV16Vu43I2kETD4Z6Q/cisGLh1/EVK39GNLIk8wGfgNxNZ+ec75y25ZVtev
gRJrzvWP/yOAH9SfbxRH4d7lV5DcapZ+T06Izc25Jgk6un+BOSeeI3KVkecAVBSa
TmdMfOWOn0iliAYWvYKHmUUtcIJwA3em+23nDmmqSmR//C6BKr5vOyMWzsTHnlXk
Iwkh8H826dzaGHCoqToiuvwd4vUCKznSqFoajDSxXGfsJFPZbm8hX7Y7nZ4gn+bY
dEJGD1RffFGMkE/9ug0bgwGQDGyF6fvPqPZ0jAAdtRFmmDdcUzDWfcFKM/PKy7Ux
maj+ajWmQKXNMNlbx8kDDH1JD0rmlYbQ0AfJnWyZu8tpJsl4joxvBrI2lv8K0DJo
C/s7r9x9iURIiYKebXLhCHAugMXw6AduhgV2YwGSmZkO67PAlbMscmiyOna2lHeF
JxZUL+PjgwW9eoVcH+cqCs4FydodeU2EmjUcpYjCvtTiekmeB08CZFaczLYmnS8A
YOVmENP+L6yUBR7MRXAjTjlf8Z6EGmJWz2xPnpf20RnY6nOMbwLg/7bBocZKyXEA
YwuJygRXl2jgdLn9UfQo1gTNNcSKnolhVRb/Q+KQ7VGWWVYDFI98nAtzX2u9PlTo
0pKkrRjeDHqFY27ARW+z3r9dIfPmJmq9eFAnV1D72piB8S42QsPyVS3O1XkMoIq/
lZKi0bQ07qxcWNkUFcdzV+yVze3SP76Wg3xXRHO2o3lATZMvNHrGAoDYmPE/SyWj
PEdx+tmqopDMSuJ1DPXXHUrncP7bf3fSTCBj4t9AEImG5ZhKhw649iV35iG4bqu3
v5mPVMrLqgDxTptzh9VkNRz/zmejItsMjs3a+ymHbFDeY1I1XdRlpPf5fGVPFydz
PTmQf+BzkMMn7czno/tayHEe+K4D1DQAp/JBPb7+ClUO19ghapIJHJHs378Ng0Vp
rjzo4VGgTBBtWrO5CP/KjUCPTlsFv3X2eOMV/ZEDzsih1/6Tyu6PcqT6bKRXaI9K
Wf0yCv/TUgpQl5ntTXBGVVFmpRFwC6uS3Oco44pjYF5FJ16UM0WFFol89tPjJQhs
lRwWkv/em/12gs66xR2LA+I1doeijK2BrNrvbObtBOCydf5wonnXbVqvWFSufQ34
sfpZF0/S210xJh1XL4M8IaQUXHzf9U4P+oFaYq3Iz3zvVZwz5b6NW/EfTurFsJIz
UAPkc5cHqRzDwV1Z2LUKxPqgP1DIimzKgvNt7YaOgFvXaEP1kepqDPVaEg90Pomx
Dp53anWJRIN/nHOBGT+6fj5z7PfHkG3977COvuP6I+owdojGYZXtm9MWPw68+nLq
2f6o5Vn95bnBtNoZ82T60PSnRyIQZkoa95uc2nUqPtqErjM0AFWr2Mi+ZJFMlt+n
be0CCxXaO1Ii4/wBkvh1bwSeC8q6APJ7iEXKfHmeDJMWwJ5sL6VDSsuPMLMaWayR
wp7EYmPef00ORa+vmd2daDYt5LVDYH831LQPIzEfdFE5Y3JqEEkO2RLFR+e62E7D
wS4h9LEEVYe0sQ8k3yFx3WqwQl5D8EROVoMi55nCbjXPezGgjLnwbMhm5s0p43Ou
KhA8q6uCs6RBzJfDP1CoraeQW4DmmRkS9UYBW+OrQQjhQfn7c969XgXEruDpDLJe
XDyG1A7CP7Kvg/dFc/vA0kG6pJVbAuOxPKlhiS/SthuA213ikIT/blnt6fpsYl1g
BBUhIr9RJ9x7daWy94Uf7wjljO54VfQYO2na2JDRL40Ij3nZaVBYkA/15SYS4zzg
O0CyHaoT57vuiVr50ibw5USCs8Z9SSd2IhHoqThD9RbLE1hg339geF02F155/lAy
ea/sXWKf7fO0wQ+xxrZRTffhwHvnXcxHI6+LULsOqPoc0jdqVHBW5aGf1dr80f3f
uuUmb5x38q9Bg5cgseE0BC0UcOWGDt1Xb7rKBy3iDdXt7bu2l/4l3vLr5PFXqGrS
v9pfQdR8I4r86Ry/sW8fptRF5K+lEI0bljxCcN591K7d28IwEt9x/3VGnt//eGYm
9JSre2c7uKD2AxkkblQibm3AWaDnj89lI8pRXBf/UTmHy9gV1S3IT1+J2eii2T/T
RLtObbdyoA2avhqTmMPz4poug7gCs8uoyAAMXp73kZhiqXIkyCF+Vpvq7+G851CP
+9peUXWESRsUnXuoRtLWIHoOfOQCdTkJMia6niGdc2/7ihKW0z8FdLaYO4KqwLMf
OPFwp4ok0hV5LdgTFOvAcm/jTOtCtQvVVOxFA0/cXeVLdMfukPhs1uDjQeMHZHFY
SK5rAKa2II/BCtjST786HyV824yQGnIW/MeDH04/gNY6D5LIqQIPaMuqgh2JRR9h
QDicDxlJXpGk0lHdx7jpO5rXTSXx4LMiXUGlDDH5nie/P0kZlxoD7MZ6Pbez40Lt
EZhRliHXSKzRBWZwRH2lRVP6QO8H52xi+IYFXeVQke5+LK1RIhGH+0vzn8eaU1/y
rr1qrvPUp8SlgslM61hMJvDFybxIgcySNqRPUXicIMvfVLiTNct8Uj7gpE1FJR7j
yPk5iih3GwDzPO/naDq4nms1P3cik8vUeJfiC9gocyQdBeHDchwjbPZ5bO9FcB63
QuTOPhEmjVFOf77m6+Jj5yYQiW9cEjWAa+JnqNonlgg952VRIU+lxRF7vpCpA8wu
5YwYNdyqo30oNxsn28DURjeRpWkql7jMN55IQwC5UX0c4kpd7Yj0osHORu0tlbPq
bE6EethLBAX8PmBk528OJCDkJUaocSYIezfOdhWWaoQt+n7IVFq2wgw3bV6TrJ6G
MskXDt5GOHkwdkzLRnpfa7ilKOlPhcX/CzZF2puFn7NRP0f5DXnYWJ38aHckIZon
obSzjtv4T7/88NTNwnomUeYdNKiN2dx0BzwLuprIrRYwM+FZ1ak/VpHRoezKOD/W
I+KnKhpBUywUGZK6L2lXNMIRII8ZhcuP5HFfd+vUOvwzQDIGC1MD+X+bSkrjs2yQ
p61egprOFUeB8893Ton1siGI1frPm//BKqKq2wuKJcy/I8Sz9n/FW5B0tlFfl64N
LbJ0qWzJQFoesAn8e2KXO2h3PvyGiQEHc/jF0rGXkLWEvNW/BzGV92fgEAlZtBfF
prSyAj5QeqGf+kmplmM9OVqsJS8DaMsfi1SHxkkgk4tHpA8VD1wM5JpAR8DgCess
enysrQmSEbHwSR91/b8NPwlP6yZp0xuroE2xeshOFjRGMZQWCnjcraETmqXABdIP
hrahZHx9BNmMnjSOZ1CB+phggp/HnAPOOM6SeClj8YkbM7xmJNfHx0s+E9y1n7DF
yBkG1AqGZ5iOcKzhVCw5jY2J1Pyr+AxabEAjc3E4nb05RluKFVHHrFaWq6vRKeA0
FzDiVxZqU8wlmeqgbcnGlp5OcTa0FuxxX1m0j9PTQ1dtfpBspAD0Kfz0XKcyA317
ePpkAxOKA2u9LT0T8iGlmseInyoXldOLSvN+xO9tSqNlutTHRRqHReQwTR5HZCdj
nkmcsf8oVsx3uBt1xG7ckKjMv2uPGJ9lMZqUPpz5KpWY0jPOfxp596beK6A0AeSf
F0BK/1OBN1zIZVWu0c6EVnBWMSJPsWA6L7ReRk0M2fk8j57pCP8AD053G9x6SAV9
Ne+YZD1754WVH/y61YgnxiXDS5Bzih6ALiaHtcfKT9QvgSTRlWMxXA5YI/mUFIuA
/ml0oNa8Vf4YbJly4XTOKarqHVDCkyh4f27GpEyjA0rYyXPNnybqW1szcmMJMKeg
E1HrUSnEDIxQEhgUQR/e+b3PaX8AvgQW7m15wvAUXTc98Xsj6drjkewlUUzc8mmM
HwtGRnZyZJpTJilgTrqO/AEAqBAlESi9r8FHEu3HaSSa3tEkhOf6r5feMWQVD+22
t078sF4wowc25R3DP5ahvoxVhw/RgR7g6YK5bVkwGpCxV4RO4yxXY3068YFJ67z1
SNeMaq3PRaA8368A/6lMtoVpS3VIdNC7ByylwInyNkfOkeMKrzjtwwSvI6SSAHzw
P1mUaDCLn9Mu3Ja43/43EOUvFfuK50TgOWkKZe6GWKiiZEunh7sc+RwTn4Iuqz2l
R5hjdX9WKjpAvrrOct9C5Tl29wGVRaIfV094fnKCImZKmSMQ7jgOVgopIozUcVSd
Tj/en7H5DJOBBhgD/U0Xvu+hFjHFaEqhWAAppeDwlOWbjelXPwDh9dLGFUUxIaKS
QGlnIboBRK/KmyVOgOD/vFXxYYtVwW6vg3lS79D5yN5tJ4Vr0QMSKUVQS6jV0qEJ
NCXoba7inG8mdhBlCw5Xq5IeJii9e+OHPqJ6lQDXVkhKd9CWm8rnL2BVKThdZr/W
s4+v8WUc4dvBqEje8266/Z4/PYd5kLkV+9/cA25gCEFXEiJ5E6+KKYkVSDzDyKBT
joCZT5XWVHzKarvfDDaqhIvHcSqMbMFosOYcl+xCc+yLnJguK0nQQzRbZ3gW1zCa
9zzXBitnkXlM8r6gFXawNsTSCXw3xPeUf/lyIdmxxaa0Tj1cWnxxVYqzmUGw6at/
wYVGzhmLarjnERPC1DxS1mpcLKMsE77q4hOHrFvrIVxQxHE0TE6KJji9eAMVmYTd
ONkrfIYlxGNlKPLu3DVwlxQZA9PNXf07tljR+c26Wz0Xq6vQrM1DINgwSf8/zIyt
oIxR5jpH7LIW1fk1TGo9REfj4sf58wF9WOO5vrnNsu2dn0X84dsA3DVHxw5/C9T1
ZpclU3LTjQBPmxGIMvB3iBPJxjfOBNXfYrHkmR3Iy1JANLo5fnNT+jdHXTPbguyu
fLnzzI3sujaiY1GEET2nGd3Gungi5IpoS9Naqe5f95cQLpBtkz1SPSA+bu4+jNGT
zMhgRXXfVabqDBKgY/3IjdUuRnvUPNY+HgGWjx6HpM3j9C03Xl5OwDJ1cm+d07HM
0pzZRPO+R2FpYaWO2bXS2yth09SSqew7lqTGtBQVmMbg7c40F0uL9EJwAnqR/K6F
EFPYFR92OgCohb7udNQ/cj/vCH3hXcP4qZnWwMDXzlXozCPHf2h41jN+D2TjDakt
y00CRBq8fXfzFdkKTPE4rCbPbw76rS+A5a5/DZqscOO1GCWcXe8rJQHRUxUT0i6m
JhA7gug7ut3y9G/tlbj/LwI/NiRMI9NrXvO3xMh+JsM5UXmbK6TIqlR4bwabijF0
AcmcRNBcAiUh2xMzAsqBNLzOY5Q/hhBWMiEfON+0X6c3+GSQW57LYWZLYvFwo87E
FvF+zwvFRTy2KHOllksC7VKLooS8uWnFEOAtp7UJJyUVQIVcQcJW2dddlscam43L
gusWHQrAGzIKSBcDoKKu/sIyieH7KNiGBIQRkbQk3fxsRd72CHVY3GswiNbyRG5p
tdzjqzdl9L/eFhoRH/hCEDl0kPX4Y4yMcuxgcsqgbFzZkUSW6WbSlecvGNlIQXxl
ryqwyb73+7LQBl7p+Gc7tKKD59P60TP2GjMPS46zfPg2Pvy0aqG3KCexFJn3zTCV
qMUmCtxgz0JtRKyrkmSa/QNKwbHPP8a4vnxYf+pL9MHawpVQV4vTKOVsHkpbZLzY
Xnhq0XkUTe0v7OWF9ZUDUPOXYW3s0ACJ7rmPJseCU1JCtwQGB/cIZw3/Rce5C60u
Fh7+c+0+iMiiomX4UDK4oRhSkIPPxi9wJqVFs7DjZYkcmfNeqZTfQSGdnHLBEaHe
2T5zhg5oXusP37BfayFZe8ksVj48zIrkamOV1DA5atLJM6HOQYU8T85ALfgquVXc
SuU6rPZfaao8M60jwSS7tgrX6cOixC1yeZzW0tKh9JdZtIa1FTTvxouNOJGP3Xx/
GR9zgGagRlecB1IygKEtgmbvANMhow8r8CXjQ0HSDrD9EA4BAS8+G7wzULRf5JvM
EcMfSHAwRFwATrXIIUDHt18LzAZ8EjIfdyDhX2GPSpaXI1YxZuaE1t76OJ84vE5C
BfPMdIaajP4OB8ihQbZwookE8vRLUiB6NcAywx1Ii8KD/MngKtryLeBnVDEX6Nrg
TEHl8RphQosaCnTkVV8zjMPEw2pcM88bQXTNEvoxZtbwN28mIabp+MK40nLM3Hhj
sLeK8YcL0gA4FKazfBjE39Zz4VK/y97D77pxu1/SqALlgRBYetERzxFpd7Li0kzA
9t4wzgjW3h1OCRmPclw0ypJQEn1k/BtrjNA+XxR36Hthy8q5QElx3cAVtQI908K2
ECzt84KF3PXAmJdE7ZJRJ0tkbMLmySegPuwrHTSNkwHIPgjUtLOr38qpdrx0gybR
SM+PgRegiXW+ynpXAPA9xOXKPWpzzapmc+5kuhyvKPusY97oHJd2mBwZXgTP/fOB
p5aCMsbhSSR0LrnS4niZ2VBH1t34z5hcQzrdKuJtYziUrAE1z17m12ud4zAp3o/d
IsuuPzl8QsfIp42fmyLuMpcNk9zv4D3Ur8TnULSxrzyJ0yqinvavfizshMqF25Pg
b84A1ygfiAq4h8E6dlqKXZHDYoGgs2ACXVCg1zRuAPfVNYoU/yfYJMi+k48kSl7r
cc3w7XAosfsG25Egc+hkeYaDcg0lObCcFjV6zpXTjc+csOkl+7XTCZdrI9Fqw400
dPxTFJG85lgFeuhr4Kt7H3ZwXPm6G/cJ/iPfVmV6WZQrvqDbRsBOZuhrIuVKWLDF
8IbS53xtJb3M5QMh+4o2vev9KDQiF4cyr0Tcvo905k3ikhqHupBbbppkKvWx7kZP
3PfJ7Y2yyK35sX+YMi2q22On3sqQsRMRPM1E0a/YB9e0Caff2yU7xAt0uuyiWU2M
FN5M/lI8Gz2OobBV1LNQU4FFMiu19U/0YSCF7xNMTgpQ49FjuOWjfFE0bNF4M5fV
iAJXs9376m6dp8R9MpnC/2NxgWo14iaPJYSrZEC94mzjAq2i6W0wAGcSi3M+TFgS
Rh6N7US/XoqEzhpRIhXEd+wWTmJtEyc6iJaLst7xUBaYAXmddmcjH7Y5hM9VLTXv
KNhuSXLVSZ10jMmaIyooyKNVi2SL8muViPukDh8N0l0mTPJtz2Whm9wiWmv88UBb
3drq0OTUWxc/3gBldPLEUfnAGbO3NK+7Toqdfy/BfPq9BTyYifxs2qEejLM012RP
va0WpNvt+4Bv5wHnT9IOX1QhU40uEtl3dzPA2iLnmQ/4XUkqurjIXtzIkq2KOP0z
WvCcgmSXbM9ZwwhfeoLNWemsBH3E4T76nHVlOEkqH07Tl2r2Onr8Lt9hpqXPlyUW
tfzf73tOO2sYhvvh1/YbcqwI8WZ9XwElVwlgQSZGJ1b/+aucLyugit0Cgf53Bk2T
gtvoFjqgMzHlUWE3wCCV82FJqk8sWtPwV7nnompLvTn6KLdMFoBq0vO5/Shj86zE
YhNPBQoHLyTU+ua3/L1RpxwA2Wg9FXsazsnhF/zhiA685URHY4w4qE8s+umCJEsw
+wBl4Sk5D0OM6h5DtqppBonNWaKeUdLRSjAJ19ovowcOowY3RNYt4Nsirjo33ldx
g2EIBnSRkN5+WXT4OaoB3vcbGtEgph1x3BldUmH7TMVaxdBtyqzSjG402PsQJhjj
AY386xKLmSj+3Z3X1IHUCj0HP9n6Y5B8jOzeFuLQnaRvWpHceQCJyqO1v12LPcGr
38hoEZrpjqar6XBciYqE8cOmYKY5+cnF17raZMLL3TRxq66zAzAmR0o5j/2b06Un
Wjcl7O9eVgMQP4YVmdXGSA+rQ2Ag9d/ps1t6QBOj9MceA8IJfk8AxCo+N1E5ym6n
iUZ3TTfuhPT7pCiyWE/wzz25Gs+9PUVqYka1orNH32LqOZ5ZaEC6ZZwFIvr7Btkz
fmRTasYXJ72DWf9IBBLORUw9iTVVyqOUFvlxfzdALWQGVKKr8Wf+O0vu0OOU/XK6
Nm5LTgrdfKH8608pS4ZUvotm3UjXx+6wRWa6Of1LckhIN5euRpfmrTLWsNaTmyk6
PN9HoXrdXrm4c6UNlnyVmnhQ9JHnCaRXosZauyrOx5yHAeOvYymncPbdVvDOIgBk
eV4cgk0aN9V12x7wkZOXEIzMxm4JvN53Yw1fJsruYkyLy+RpWQm3m2vV4WCbAvYX
f3LCcTyq3U/kZ0OGV85YHLNNqZnmCDBDUWUM+qeCBXfNLFeF3dFqQ1UcJ/9WAFOA
y80bf7juz/Kmulgw+gVlW5yL2wz/23R9JqaRGLvEM9DtsZRpgawWby7X4yNSF+ez
n3miyvI15gGf6Kq/kpzZ4FB9GBrGQOAXajCUcjcx1QveZhq/lSW8G3/MgZmIreig
yzD8x4bUJNYCELNdqnaSBPhdTM2Hoc8ev7mZOiyjwBMRyT8NsaVEgQTacl5PV68v
MyANOR0FIWhbk65yV+e2mssDPCysHU79+0B7pJGzu7itcpx+PmFiQt3S3TJJdGvf
hbPf/Og3VXCVrD+KtUFih/ghmQmkj8YROUI1q8bmZyNlzFNKch2yBBwHDOzDkCmj
pAtJpfitNhb8SKzxheORwwu75Td4RXT/vSucESNd7FLixEDbMu+GjOOBiu4vaUPD
2b8qzqpRzEhELv8zLWD6fTUK5j7TaGF/wD07Qh8dj+9KTV/Vr42icPKRr/Cyl+xc
oWmPDZ6kSs44gEmUmFSKBO84hRY2okLbW5aBY2H3WvVrvqYbI2ruKsqgfR8SSRUU
ySLZljfRFK/a3zKh4HKh4DG4L1JNei7wZzlqDVqDH7bQYZ/jN2pe8XB7VK+S/pMp
+ow+q7EPiS909QjxlOIjD09dqRuChqSl6mWgKpk/9zCLcgoASzrc0dffXikuiJvs
8xNJ4RJpoMAEyrc4sxt0Lujx8UnWm/BhHhdmQMxHOJm+evX3zJcMl9BzNQnhDf0M
Gxp4xvwHVqwca4UN4W5bUNLo7/2DceFcILht2xZnAsrOv6Pbow0ZZBZ7au1eIP/x
LSyFLivEfwOifRkt326by5SthOxVRl/T9VWMJs3hSSyAc15y1fSkWr3x7U7mD1m6
VPo04qmyjr9zCEa1nTjpu+W9UlsYEwAb2qY4e7q7aaH8PpjcKUuLhzeaFV0Q4WyA
08t3FGa1xIkFqkDtCzj7+RfQCI8+WJK5T6tSVKaFMX5htHesUijKp47N1QRae7xY
Oe4kP9xSzBY5b9dSWAMpZLDocWxL6TJLt+gJA8bICMsgz86WeTeKHMFU9eQyBiaQ
s65RTxFT2E0zcI0rbWFAb02Xaqxua3Y7h1evA4ymrfH7HUE/FN+VEn07BD5NeRDf
5yAI2Kyi+2tgFjb62p48HweDa9+gw5w99xMK5Ee9zcLYrqncUUPTiYnwVqygnuqA
cf5UVIo10n3L7beEjDM27LzYe8ZLSS3y6bxj7GwdugnjSN5oRpd4/nxpq2tlqY1p
wPlTRB6EnlxEwN9Xf5SvsgFzqiXvufFlsx+CgH8zFSVBiq5b6iNxGc+KVgSgx1T3
716XEe7+L0Q/hfdbAC0AG7IIToqKzGqJ9jojxzFYUjExihWiLO9lByg7AXNMUdNt
BXlCySWIznSDeje1Km+uIcqfPpb/vUmWEfGL36B7ib5T1vpTU2CI4Ddqs808VXuo
+ha/+WBl7yOw8y20nH8mWgQM5g+J/kNta6sjfKwMfHgNvXhMbcaT+vBtfKfjRdgd
rMrU8lrvOG0q9hwqRsjGE+xucGt0zI6YM09Lw3SIRuWwAy4NxHr0FiD38WxV4kCo
izFDbcIycEC+ufJ/75VZniF+SWwj4VCukIZn4zCXqG4l8+63a+h+Jzum2kBFz2/j
spLFeebEcbgIc2S5HvKeYRGXt2rIfLoQ4aWxX20DB8WQKVqZKvoFwQNNjj1lsGJY
IvDe0uaDEwsrSTwQFSk1v8Ry5ykH7je5uZ42acYYzHQ6H6+Ni9mE1KLTQUkzdw5i
MubaU9FTEoFu7zFqofE+uxAts9B4vd2Wp6qD83aoQc35IkEcZXE7Dl9jyAvuDJ9p
t5BD43OyliKQWMA4xDj8chiH6Gve529JWRKDlcRgFbJ4xu1bDny8FCaEh8RiEFnG
PZhxzgLn/3jrj5FCYh1kg+SPFLCprDAAJPC3mxGgVyKZ9BjFxh1Mj/OGOPIV2MuM
cpru/kFL+IWR85nInidXIf11dbTx35yJfACyX+9upAdDVv0YWWIGUHB+iPXaUUJ7
EIx4kpYYK6grBRsX7+bN6NWesWZ0EdxhZ75iM6ckxf0i1MVx99tOOc4M2ESEQsqD
293hEZIknIOPCFnZThctf+aQjndVXPw8LkCmAkxWCeSqvyaqTFkCf2W3u7ug0nA1
LMVbwyzmn5tGYkDoKGFEsaMbf45tOXnbhEBc6I5P+2Q+s1inubxay4uNcejkRQL2
DSNMCSSma0jPO++oVZfKSy5AFyVXaslk1/C2Tbp3HJFIYx/JayCg+cSAB55OYZ/D
+MUZ/2IhwS9cmTrMVrXhy7gliaAN3N5AGGcilYnY2pDXoFGNB65Z7Pwi5tXflXz/
If8AcHQDtw/FjFE4BjAl9NlefrY5LjJuwUU5ervzAiqX5zJZL7XD16u7z2o3zj9u
z+rmxIFg+Y9JtHcfubCS8kpGZbCsxit2bXt0qeIFSD+r00EPzhjQ10o17Ub8cvIS
YmUARuLGgrXjxoNgfJ4Tky2RRp39jOVXEPQjxqomAI4A93eLoVfxkNBtpfX0Bi8D
eTwYdvn0rHB7ihPchfRFH7kdCwECgH/OQdXRuGKEHPoFnOEn12M1M7Ik6XTfFaAY
8yp20fHst+IY/pDN52GxgPlRzC8ax/h203Z2FrqEHagU5eNMOefHezOxGj2W2Ec/
5H9m3Rk7WcR4qyrUd2CZgjuAP1Fyd4OSzTE44JfVNiXyXVl5R/zP/chQiCtXWtu5
TAgf4U82sJhqzMSNj4VYKsnKe4vPuuXLrRMtA4us/PlGVwO4AXRk28+7XdLCKeCb
joy0AqcSYzGOPue7mPEPjPBfQmB9+lZnf3WFiyqa5HRY1lNNuttcZFqA12FXsUln
Yvtd23biVIB/YKRS2yfTwcVCT7zsvlrkBYrgWPGBINBZP0sQs1DF8ePl7MaOcLBL
4vNwAQFrDb6GQUL8ng+KQEL281H9CZojBUJfijQXWrYh8TseZShktq7Qv+sTln5m
aN6DIcj51t6pnkI0vsMcQqnb1mFrg6zt2ajCo2O6EX6zLjQLocbVPf+LCkGM7WGj
dHVOjcT2KPUGV/PxepfQTZC7EQhzVVHFJYJB1HOi+xZhexFo9yiapAUEfKYmhlbd
Kd3X9kidVQPH0oNFRndPrnADXNC2JRzgIfQQthKjqbC2/s2ck2Ykbe8C8NonLHzb
QiLrCxJc5EDd/cLBs992nP223qEC/EpwxVcebUXpQQsjos12YFfds15MmvtZ6fqX
xwRw7EDTqd1B0zEUbYVqjb+6YneI1kTJBzU3f/e6G3LyB/9yAFM0ZAFsMvU0A76j
h2mX6+teuCk68Oek3cpOqvx3xnJUmLyG/tO1eMT5spxiMw3J46mBNdbLC1akwcqW
RQzTkfsro6sx9h5IvsR/Mqst5S32ghv4lIHOv4y2rp+pXwt3QtMAoIEMDWJLj+5w
071eNIHiBh+LM8WCUmJS0EX06BrT8fDtP9tW19ch4vYprswbFL8Hcq4o65VXQKuZ
JKhCbVoOuIDZfsLuKiuMJwwzCG3GAtNQY+h2p1ZpftKr6b+d3WWZjnlp2QgI1qfe
9jLavfIjdcgnmyqdKdIK6UIuIrz3NaqYEl0mOHrS/0LGh0dV1sV4KhY4+UvGti8l
xhGAzYVbTXbjD9g1YLtoxMf9xJgBDFj2a8sRFmzheYvxojQlUY1APMxcdgqxShZG
3gWGHEx72FhoyXV2SRAg3OqbkM/6WF2quN5QgcTV6UjXx5In3LU1AmvDJOJ4opOV
lIcTEItjoIMF8JWWcHu+bPlt/U6Q5Nj63Qj9A/CPRWeWrKLPRjspA+cfilcl4AnU
aM/cwBQ0rZK/TDXBOx/ir+C4W5AFKqcZmt1hNJzluPeErpyQR0FfI+F68y1LW1yO
RLvmPstVJTVQyj1hPvi3kf6efbhANMkVsXtVUEtD5LaWZT0nF33+7zH89TeatBqK
BjxOGobRWCof0oS+McekEZUvQNZYNhhBtZcW4LUMBcpzB+6410RFSICld3aKYb8x
WSsa65zGyDHlFrwEYpMe4TwVNai457XR1K69yv6altAdl/OwY7+1fNF57qqqr5RZ
60YWBfYSIGjVopnak0sKX7Skt6/fNNT1eAjRQXsg+OraHRqu86kCa6GQcVL/BzjP
Z26BZ93hRVtiEpMyFYdKqyNMIpeDFRZvqW15R8OoiaJGuIHH1JZ3CQ0km8BVpDtq
ezGSFALcWoXWXZr3r4cnh3WnaJc6eL9CHgtW7svDwYZkuzduw0EtVudXb620mXkE
I9opM5GvDQiaM7UNRlp/+tYvL3bvWbfloPtff4Tr1nblpMF/4DV21C6N4aZjKY73
lk9gu3inYsuLuOVAt7f7aTp30phv0cB50qF6LniWNTxEOVMV5Urw6AEfuGujr2T2
Kgk2DUjwBlM2ql6F9ncpXXWGEOGiXWZf7tsPruAPWBwuTFFq2sk7kvA6l/E31CJE
iaU6GRmOV9XgXKXxfp50/Auxxwm/7JwAiCUPFTKl9nghYyQBrYbQJoycRj/U66Ei
3Q8b+nh5NuE9wMsAULfdGD//VOCg9fabGHlY4+29owRdNEW6Ej38i8BrCHHo9tpk
I3KvtlTXjVQe47SrMvHNv+uCWfYwn94T+W+LNj2OY3+es28AN33waQ7Yv3D1vmc/
1d5ARu8YzBYHuCepKzISt7prxLtFd3AfqAiuzO2gLzlMN3wvCV5T5e98ZvBk4R9b
K4CbqR0eW1xz1i0BrJp/rwQ3ZhiCl2owRarHbee0aZqnTn/BnM411+/taxpAMgZF
QQ9VlBGByXIAi4+2i9KMdwVI+AS7YBHzMx6zBcFoHo4N5JdiEoEX+aFd1gii1GJr
qP0zDeGdNzR9nw6wVyGKdkn6OQGoqMh8XNE1rE2EaT6pEl+odS2hXPVyIbZeWRuL
4A5ERGFjJVZGZAQ8jwYicEmslsX31tWuO7FaHPEZHElBzf+7q4/TqXHk3pPg8qkG
YhPyEZPxJeJw0SIADaxBIowIKHHrZzOHkufjWqfEj39uFf440YHsPxyDAoi7gNDU
oxiUwzbcJl4QGum+ybYDeLlVXtEMvLxVCeveTcvGSyiPOvqtPzkmSwB9K3XwLBgN
XvrwkyTCJWKXQQJSxYIc379MLBzR95VFCWG+eyFH2VsQWmBRtO4t0el9cpk7lG9O
gdBIbLPErIJzQSJ2aypvCm3oZIftpUA7fRftFAphyIBuO2NOZIVlpmo45HjbCn5Q
c90ZkojFQ8HKjcN0uC70GfQTHrd/lo7YfO9KLjuXL/njggfSZ4eVGbR59eMDzQ6G
ppsN2h2tfitLCkcBmuf9tSf9pjM/fK6wCCDs1kr1XQBTM3+JQEBvXtCYzrc0ljna
R95NYro7p9NZPjGsjUAjMD1b+BOeisIq3KKcij2hXQ4xpgdrKJ9TodmzlAqeWlV6
uN15kvCgl/d6RU4DVVd38Jr++kl1s1CwwTwG9zQU6OfEZk18Ho8/OkJTCmlwi7c8
O3n9/KENCMlkRLraoMIwhNco7OF06cFRnajK1dgcCnSer6+RCJOnGu0a3ssVY99D
gEZKahaT9XbVirEgj5G5xRzx2rq1EQCm1AqeswzJGbC9odPkOw1Pi8kdIxVZG++W
tg8ianmx4UfVW0gQbH2JSir1Ww3tr9VHgliuZfLBKsyMFSVnZLU86Tg+YpbtHOEB
oy6PGmNY92kFWSN88x8s6lfsepCEZHDZlBQVH+hOzRW2XoK/vMMj8DaEW1N2AGws
N6rYg6nMGRCVeTB+gogL/hvMBkXYEc3Xy6viDg6WS/1Rb6EOFROScMhyYLHD1REK
/xClZwJLXKRHQnp88Xb6gD7IoLOa47lnEhL18M/O8qBxSNL30gZpWXUNgB9vTes3
0XyU5NSxWhIYxgmE9jSdJeTNVKmWz21g0sTEx6wqpnjwfcvxd0EjSe1Dc8wH4PLf
5KZA/Fow3CBM4FAYa2r+5yjRDAYVw9XsxA/Nc8jXQNbsQgzAi0EyrOGDJ1meUAhJ
Zaw1U5z3K1mW6JLdwjtQb++hVZrIJpVyVv+HDdzlpn+cNc6wn2HB7wfmK6pxEOCf
NrosV9lKVLn49Lr4y4LFe4D2yaI1VCj3H8aXwgD9EjEPWZLhc2t668+G/DsYSCXS
baFfx4COX2n9B5GKktDG08oliZpLj8C4Totvw5qBDF1am89/d+rvvMvliYpIlt+K
L+HF3hTwV05kk8yykhibCb7C0TFNoIWbvnml8BY1Jz5iDzR8lUUxVwV0cXX3iEkJ
Zn5fXzBn1mUbQGJtSxFlDm8cAPnhn9ppA4J8X54gGhBpW8F74zvrII5+B9yalP8I
LdUVk2nBGFEqolFCetBLv0QaWfUWLVW9zRAXYflM9nEobHdKIAal6IaC1STZSlag
DgXRfIKJHzSJt7ZCYc8Nosy+/Fv7Xj1zDC/jfjOSc7unz18oHxkjxLh3JqMMzE0H
+ek1aSlkE4QpFl3KBdoJOFOJmGCd7sG/3KwAYGqPIc3w67mzn7qR8nEJkI9bKBso
mEGeexHhn1lPKseLacjWccn/ITZExEaikG5qJH0dbMWE9nlZXG4qKTEuvjp+XGtk
yAY1GdjBaM40AT9t+p8r20qcFDFCQ/ZegCC8kb2prOHwJj1fNgSkr884I94koU9Q
AFbHYrXQS7Phy7XHIGZIINFo3GwZCUbKE/X3paV9kdi0ROc81GDOwn2/1/k29nw1
tmlWQxF5dExmC7+wqdL6q6r2pgwf7hQHq0JFTGd39t4so3AgUuKDOh4JottLIBur
PI+Xki2AgqrcF2iTgpE/9idpoTRX2hm/V+RaU65ZnqtuTd4LIl2rtttbGScqnGfO
FnBKdSP57cbyJqdA16Yz64yXdT4vS8ExN2EXpP80lpzX/O3/ePsI9Kknizpqww42
Gk+xXXlH3lu1XAZoLwCItyKfIyDR04IPjbwLlw+xuuOgxYheYoy4vLiWETAgCe+g
5/FXD804oFK6W4863jFv5MQIQ1ceqZC8j+Ormm/9jypoO2xovn32ir1MHyJ7k4rH
8a6iyimGB3FeHEqzZQX0K6+53sq6pBhNjLE4BdbqpjwLRRXVXAvLV3xfKj71O86x
2huJUdanKUPIQqTl0S77j9EzSsGyrz8fIpBsTOtHesyt6VzK3QJNRFzjhKU3nI5X
ai6p6cBcvlJXKHQmtSqQjgmIbn7cP83/tK5RcAlX7DLAElJgXkS9mW2NWejCAsYn
DeHwMGjiSTIWfmpeeImoam3RrFpMCwGvVdyfNX6r4AbhSOIcHRFReNZ3TVGBBGrm
gi3BZ3Bi1bfVKq/kL0vcMmIdDBOlfE9JNi25dHMkm3HoRJbB9gPuCP4CyPSi3jHT
X39y4unjl/HMGQdpJRAg9lwcgg/FHfZnKK1p9xj+zrIF+uyHnosGVXiWV2Vj6VRf
39dEfjKeqy99gPFxrFCYZdj9QYMPySjidj261YxVhgdGJVpNOukFcyV9Qm09LR3u
caazSU+bcL+pWsFz4NjtHnDrNnPieFlW4k5UihlBVqc2GrWijtwFiXMdhzyYa6Uf
I4mJuFwRVmePBhc0K+PYOs+6o7XxYKsAtavoglt3EHCflU3KJM8rSKpOrfcu8/jb
+j9Fs95t6BGGlOJA8t+gH5z6OPz9yRr5QXcGxoFo04SlxlRnCln0RXwf5f8fEwk3
6efRqJAn8xr3tWw2S1azSJXsWoP2LLdjEediJ+1uwHlCIsFYW527k+SeIPWBRecg
FryZTXf6eMITZwvmEvwaCWH1ka9QvLSQM2clzLJxU54jTXqE/zfoUX7Wy8vKHXkP
M4ZGXa4CpzO1fKs5oJkA0m5f2mWSUNVJ584NON/9YJxFP/XEBH3h/MZeEBdG4f8P
REucdSBx0kd4VtDX/4LlWZ6DrKTBBtfdt2VpgLrxDOzvkCUN/tngJnjOpVUQyikx
U3qrmSo8IFQu2cuPu8xDkBosxgUqqzmRYDjCKGjY0WMzFFsZN0ns2g1IfoY27Ng9
72VWK9ItQYX5CaZWE13QAMrOv/N/fFDt7U0bU5LvhqRNbH1JXKbDrREXXyAskXv2
U3M1bV4DT9QyRefs9YdD+5prDOEoLScRs72h+7UB/FRZeyxnjt1YqagyW6kdCTKY
wcLkSSqlvUrfviKggl3c5AQ9uJCrgeDdKV4K4gK8T3hIaVOAJgSFTeU0ZH+yJPlm
Dfo78WUrDu3Q/L6pDtHhqWSXRx7bvcXozA53mgtZ1SGbwehJVdvGtaSC5t9eGwrx
ZGiWY6IV6Gos1j/cm+u62Zy5da8JYLLS44gKlHG1lBQUvorNORVakIiaZXC9pOV4
mPPFk8xwrN60rlN3SRkhvAyZi1b7s+c+cSMN6DWTNEryLpXaO65Eu6/+abulg1hR
KygMHheyNOgvzN/F7FcLJb9hm2fyhWxNrwGeX5fJoKXq1IHHQTCk3GvL8faXVeCz
bQVU5yH/HuiF+g4EDVnV7GGc8RNGAXufWXVnxS5/pCtdQxZ16QlRQTWRkgbwjc8W
YOPFcSHWbNr06gA9DCKrrH0qrjjNhi73BVWKukyK1VCDVhfvo7DmlNKvZNifxFbL
Av8oc2M5wnVkFwQ4X8K1Hq0MKw4VLsyG9GiKmg/N4txYk9d3w+UzGD/mtRS5OQFi
mfEVhLKmy2EukKcG82zlSW3m4aHys8iWUC4UL8j7mHgK73YnuOlLok+2dAWrk4AV
6dl3amSzTpdOgk2OnR03R9/QqC3SBzDjF3MnNmpm2eYoxC+gGC6nR70org3/QdmC
xd5LndzpOLnYEGmL3sTRR3Hc9C1FP4UufBLW7Fuo34R+L2u9s5raQbKGlE90UoTg
l7FY7sSE9rsR21toqr0EdR4lYUnVjck7YGTnEmkaLwQ8887RJOZkuHMxV3S7gi5/
UCbu49YxFAwmpCCFfqxSyH/SsLM+wGs7UP+CkoGpOg4vzQVSDOUaXNXt1DWDKGpc
RCXJ5NKuLHRKhEPxUCvrRjZM9grplUgIysCR++INQ/xY+M/HturNbPRPx40Yy/EK
fxlKaCTiMvmC8Wyp2HANIxVX3UIrsz1yxBJQJIkY+FN8OyN+f15TAbc/+mrmx27V
HKF4VLubM1jlZwSbWl7lRNmI92WDZx8jrvQvGaSZG6MwDoQS5yvFzVdDEzBWKH4I
/7XJFy7LxxfIts0eeQH53+Bqg/KNEv4gmSKVXsYQRxsIo8k7b7cf/w08ujnPTPeo
sKDdGYlUDBMCFhEgA/C8rTbqHa9gI8m1riqBJhnx/AEMvWYtahSRbZjK7cgHujfv
aUOe8aO6vKcRrsXblUF0wLvqqOw7eozJuRn3tW7WrpRHyFs1qbyFr6SSnvmk0EK3
z85gN14elo5+m3Oyr9iiqd/zuqFYjkHJM4XWuydUJjcoT05SpB7469CTKiC7LZmc
FZygIs0lTcq25MoWzXV0+y2Mp3F9603sOTn274T9UWNgRtfV37ONBdjBh8igB6fr
WviV13FDpWqgYTlhULxrI3ebu098n8KvDuz76c1YadM6ZJjkF8r9PCnS/8LyKDOY
9g10YB+pdLV6whksWnNaOufMJFUCKWX05RpnXbq4dYE6wstTpN+6Kr9tHib3Y/3U
PO9KCiV+wurf8NUuEKLcWHf6c40YJnALh5RFbYlEwm9zP0A/PDHMOQu99bYMO5td
iF+p5tZALo018AAA9Da5VbnA1HOnNP3VBD0KT5B5SmUovidvWa9Ki2+UnSkRKxmH
iKBdGtGXlsbhUe7DKR/rM8nfCax+BZPKkXOBNWFcW0NRuEAQySYZzoN5YJCdcTE8
pvU7r/6NCxUqdF9g7cVVRZ8zd/J8RPj8Vcgvoe2ES2+oMPxLW49PJVmJXT6/Xgpn
jHYbFBfJf1oVFy3DkzI2AVgVDQ9lAJem72Cr09QDwKKZce/nVHHwe0vtmCt0ooQK
Tu9g+ezblzYB0Bh03zjuUOG2PB7qWq9Iu1pkw7is15FCAqvDSZuySKlYWY6Bvx+T
bI1nK1QpD9FCWksfxb99pO0FKgMjsZHw/MKBve8MzQ1muN4JgpaLwi7GnbZ60jeL
Emlk11AvxZJgS+2fd8U5f/steFFbFMgJQWQDcOtIky9YvHFzb9kRU1aJ7WcwXpnP
N1D0G3N1Hlyq/YAIF88yecLxdidlKC9KisSo6x5esVfgV5f4kyivDPxC8ahnxHBG
1IH36Bn5WwaYPeBKOZ7Z5Gs+5U7U1c7CJHdxdu/4Oo/LgvCUPyBPPCfbQ2plcGdA
fN0x3oK7U4GSX+XmEBce6yOyHKUrJ9VoPLX3S5hXOKwCJW7X/8A2ACtW4905GTFO
GHAwQHBIZhCaM44hMdsGKtcMIPVvLX1iGe5uGVW6UUyMTRxQgBGR38mk2Jm1r8PI
5llxSUpEryIavhmPDSTpu9rFBMQ6qAlC+osqIhnzxTJREypGBpBhnuSFFVACHUIc
8992xqHBQ631lA+bK2IJ/tuVRTCnhVZVLxaq1XR2hR7Lik5mpTxzHz4wL3owqtNe
KCqpxWdw0rNwn1T2Tuv384p/2kKK0fDgY1ntTAzm6OtO4BqNYvc1cere5FRf2cR+
oumCyGw6YUhguyl52TQqyjPh5OsBlRCR/htb0Yd3RTWTCKW3sz6SlCsxkfQEHGXw
DoEO1jxL50fKbtflETRkY/tYcAmqw0tf1PUwGuRMwNxH10dTSaU5UQ+XHZN4pyyg
CH3JRIGOekz6LRwxcrs7qtr3E8VA3nQEOyqgPDdKqxbEg5NhD8T3UtO4yutn6+nj
oBBxu5fEx8iRsshYRxbX7xqOmc741J224m+S1RDYsBtuPTKp70JJg5TGEjcD0Vm8
c4/o17QSOL/l8r5kdSVIjieIBbmyGnis0FomMrQUHrqhyUEfHVufSnfxihATVk8t
wUdgJOIY/a745wzSczAnON7pQvLt7CtIy5hqrZaToBENtD0oWqdpSJfSBD3KokED
O/1wgc8VsKmS8RjKa0/ly+m4Bb8oXE7ZCL0bXLlHN0u6Ozbkn1yAbjQIJupWoOl4
5SgbOafYjdMeSBIsECAYDkADIt1sN3Rs9uCOU25pM1qxBUvM70te7mOqO+U9eXab
xpOCi2gns6bUy2wIiqKDe4scUWrAXcoET9iBv/XKsODvgMXqYN0nLHLohkzE9h1Y
rsBcDXWgZoZwkjcHhhU+UXpF7NBuBiOmf+reXQil9C0ZftJzRbv+sbP84JweXEtF
km/HekxyBKuxUoiUM6fuX/noL6mdovefTz/YsKmBqNEaEMAohDmE2L3mElx8APE5
+vlRCxlN8ql/AFTnE2vRktPLGJOEGugOKhzNN5CD+RLf1f+/VxAdLQoIpwjsp8v0
wiuKia2ezhFjv2KHqp+OBHENqVGNhmKd6q08KktjAWqtHn8xYvZOV4vCy5W+J9aA
CL0lVr1m0BzWzaV4RZUnPHpfkfw3efBoTh2Ypd4jFKYoRA6jYM4ykoxYlJnTEt9m
HDroMvVMbyVGdB99Fm4wPMt9D4FdJdONWaBhSJdt/Cf/s3eLa844yDqOK7ggKT5A
DKE2wjoe8VXPVf3cNKJl0TbO/LAC7Xl1VbUCoGnC0o3ncmt5pXSgrZqPTBHxqcmc
wNz/48sAag3U1gyrQdA0LkkR+l/jjyejfS0atHirSLXERTQDISCfaSjE6Z8fuiUG
UgFC+xcopC67yM3y8JK1uhyQ2qM0D8AxIClQX1XurTJD+8o0iIizOhVkcOHuRhxB
eoWjofnwfHN46QLHikGCI/bE7UIy79kfa44/l96+/3S/m6CcMvlvzZqXcEPm3CZz
ekxha9pscDsQt7GBuitcUfthRF+2mF+osBS09RggivkK5xaGLkSA4+d0MtbkJZDY
N6/PpIfkbBDRoIF44pWOVcF/Bq5vnRGusqrrZkFGIWzap4ZyJDetBAjaBnOWHDiS
+puNNgRo02SOcSv0E2n0msJVlwuCBHUmlwRBfMZ4qUsbTFHbMU/e1ETxMJRj6+hf
jFYRAjabzOxPvh2w9tTXCjMpxR3nxQpDAGXnukXtSf9zuIRDJFNdwpBxaapiB3N/
T24/UJTRBeHOztctNsB9EMfviFwOtc5ILAFVPKryI4Dp7ZTtX9Nu9W0BF+MVfemw
E9thlgRaLJzMenoOscy+ZtKaGROGkhaOD1nT/PpisIzDokxAphoLsybrXjKGAV9I
PJva9yPQWEu2STwY00/M1l9Yq+k4ZemmTnpGyzPD3qgsKwVuDci6xI8e42KEf54+
M/DereG3HqHx7G9eSvG3zqC+/rwCGZtuf1cYKqXQzojxXSSpThIhO59no7qpdwgP
qBc3lgnBWCsIuncr7SReOeC8o7uWl/c18WRT//bj2cV6H50ZITA9Rfqp0a1aRV80
02g6fkQsqV/K1dZct6kM/aVKKNBubJDspIe9wMA2VBUfmEukKn4RPftjq7cMlXKb
glUkE5EdUfxcbU/rtxojf5h7eIi4oT4EB5G4vxsXKjkW0EjdVGwfdQBQNr+aI7GG
02d9xO9UascXV3h2uCt8Esiol/wpuL/jsnT5d2ULeR/JCMMeqDBOt2ElQMtTCLi0
J2xfvKON780aYxQmmdl29OjmzzXccFpHaAObFScR0DJQq7aRrLWKAVKoXbBmu+Zm
K4pre7lRj/Pw+cWIVxLoTU5B57rQOBTa1gtdddHyxJwge1RlqFpXuV05s+Tg2Cw7
QnsjD6r2j1pyKWXqU0Qe0H1P43y45hueuZVzZOtXgUTyOZyjMQFgd9ysGaC/wE63
JQqD0Gn95rJC6o6lV/5lx9jRrFQuYcKnwrNtVCy8tblu1KhCeNmGjzT9EHcFedR3
7oMqz5rra5hIDQoQ5uAH9We3WNVAcZCj02E+JahesjS+t8Utnf2Nh7TIP1Mr68PR
gfUZl9k0Jgzr5AA+25MYXyZBVC4brjWgm4aS/3gLlLZw8BPKygH7JdIZDOs0Xw94
O/mt31Iqqg7Xc94v3yI5Fwsq/NDl55p8GzOByZ7Zoi8X30QwJPOI/ePY8UtUbMGx
mQQAXc3qCdHi+JZTidSBzUFz8Tm8lw5doCyegSkN9pSfRM7Vdp2d3TWGo107hAPZ
rRUYUqo46CTGKmce3obdFINqQ67c/Eof31MdfJMOXIJaVcG0F+qeb3TPy1l6gUnY
hTOVmw9hViPTPsSPlY/uRNhB2Uc4Su+ibgyOGJLdDTJtbW8AHuKz1ZU+7OqQ/e6z
mW07yyxpvTekU8XL+S6utvflgUE/YxQ51TvQeWpUbTbpBQdKZMCrOVWrrCdvmyTq
5jifzVEMEb3hL7DQ1121O8QCklPLd9TZNmM8Li54FP4JGuvxwBayP9qCRm0vUMNC
0qZ2ibdm3orPaXK1f6U0IGRK0gr8N6Rg/o8WjEe9aeCiLAliHk6yYTvZU6vHelAX
Yht1KAEWo2KMrzN2touVtlbYHOriQ6k8lcuKruGXpyBcjrOrafOaes5wKLcLbrza
XyLHLQK7vtXxTtjZRj5gYAC0U3mhMkRwHcWcnc2EAL+HocbK2sO7lF6SIP+3WBSC
/i3uGPXZZRun1yh4nR7Fga+ppRJnEouMeQqxepC9B1TodzOvk8AO7vDfie8ngpIs
IJOcOAIzVleYzzePym6vPAQitBwecJAlbXgGr76WQVn4rJVA2sECQmlJmsUyXaQL
e5o+ob92ja+juy2/6Docl1nVxjS5d8TUA7fNIK+jbGfWEu1TTi2jNc/vWxofcDpj
IueeaV0QWLj30DYcS+1B86Z8vA4kiI1wMBBYokosFiHEr1Z2DXu+sTCLYr6Ferpr
RuXKCFq00TzuUU8/gHa6TK8n1mu/ZF6l5cwmTdfCk4eNozvb4V1alenql0KgUFsI
3+okWRT1XJeLB9zfHZIP55x6iWaQ/LcoCKfl6uvWqGYdht7wNaFGcRJeHUS+Zfj/
VD+FlvVMQdOpfaSeBurtjQaJ3xxqRmFkqd4pvJwZB+6p6eIgegAdqrH6/kBqaw4m
YZAnE4icbjFBmLrR5ppl0l3bepUaqqESDKs30Cp6UZlRxTT3vk5oqu4GVzEdJXgg
+zp67XoOOE2zMENuqPxsX/enHLB8wcePNKrmVKd7ycphBiWRkyZVsSGtmmtv4fkp
dOBfk0SHUflBvDAC4X2jTq07xoVx1+bf2vKrZn2FFi+X1zmQWIuSEbMv40cGioWR
VuPJitACE009EnvuaQ3DQaKg9wbh2/LNOgAupOnRGHpVVYaK3s2xVJJFfMvfAOHx
OA24eY3yt0pMxiMSTVGiYJQJZTLUTBB9pezl16biK0gXq5Ea398mBasligLZJydb
K8EyPWMtMZL3RIjeKuMzrr2YwwCM5VixRS5cJ5owRBGghe8xpoOJouP2vJFHQ/l2
L/lNizlhAFC0SiZ1INs7PE6nXhx5B1vlsrtffFFFefmwx4+RhYR/9t44q/SMKJBl
jIJ9CtolN1EAL8uxL4gKVcZXeCR+jIdIR7GVL6H+9WMqYZ6a+KUXnUldtRZFswN7
QDB5j++v6Zk4gQ4Ux1IO9OsvkPJKo/sXrswVO0UOK5ti+9wy8UDaFtPO48+begHW
G+HbNWeddb3lK/PdPsxiVVkVJCAOxw98GaFSy2Rl/gtV0xedeml0KU9MVG9D9aY2
G4k4cwlp2Z1QQy2QMI7SnSnvncda3hcIJk3TcDWMzhVwK4uONzMta4cQJ2p/ouVO
+jV5Cn/vsbNJeQ9/PJEwBHKq9wkUynWE6D471dkeWWKPrfQYroZ1NNzspfMgGkyl
owaHMuQFUoMFQsETupqsN8s9E17i3Rg4VD0dKQEvh6zhqEcDEEV9kbSLXt9M6N6+
hirLZKH0Ei0OeQO5C1U32k2B1uleiAuTYJkWDKA+W3rWZjpfwnpEyic4e7+14pEu
lMaMyWrq7zp8pfqH6auXo6EJatek7mHLHAIKRfgfvDdTy6cjvkfEkDozbU0ZyB53
GjJO6OvZRJf8V1LBkUYs4uNG6QR1UEK4U9ZcXo8PrEIe2TA5H7V9WdOwrS/j1KAY
ioswrEa1zPm1aLhkfsKeoKfhQG2dvfneLvLrMgWErj8+1dUBCOmkLvDM/pE6b5O+
8bD0+9puoCIJrzuKz/f9p2yAEQwbBoca3v9gLmhkP4p3qrScnjwVLwLYGnD6K+DT
NmznLSBIKVlEaRYdM4k0Qz4vTZ2qT+ZmUKKulVv6Z+GW4ZH3InTcx4R5zH+nfGko
50r5M0mdoBf16sTLsE/2KgeZXsCaMR0IVCpesfkkaEvg8nQFCWitX/qkIWthQN9T
`pragma protect end_protected
