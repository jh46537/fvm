��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�����jA����'J��V-�@m��Yx�W����'�4v0΀�A���^��-�1~^��R��U>�RBv	��n�-۸��Q���en<|G��n+B�m5>,��q�4h��Ӫ!�j0h]���eB��w@�!_3���:�����!ϩ9��WkUwqHt�C-��BK���&�U�����0�P��236){o�+�d=e���R\�-�4�Cv����]��˭��|�v��#���j,�˻M� � Il���(K �OkFYa��m
s��l~b�m�٤p�o4C)օ���&~!�XzttuVI;�+0~`[R���������CU1j7s�H`&2�d��s*p��s�B�+J���\�rj��O�EgKԥ����#{��,��e�x-!��;��Z�Y~�ʳ����S�|~���vZX�s3��a>����)g�kN��x�^g�*�����TJ�����%�uu�����;��<`�������}�	������]�D��g$��uK���������KW^��K�XK͡%=!�\ۢ�����Y�|�d�BQ�z�2u�����W���;��)����$���5��QL�j}1d/ޏ�w���1��m�ʕ��єܣ�ձ���c�E�8I�D��#�@����-�;�u�.c���\�4c�������pH@��6Z�L
"j�^&ܭ�-E86�cT��9O��������Ѡ�?�w�^�02r8x6h�whE���Ք���$46���܀ꛀN/��}��,�#�'
���9��;�1�T/g �^��i�<�q�2�&�K�\�@O�!Y#�z�Q\«Pi���`ryÈ��6�5�y��4��H�C���[���$]$��y'�"�^����Gw)y���뜁v���z|�Ui~�n��ڛz�}{$Ӣ�Py�Nq��my$(h� ����LN�����Gp��KO������KgY��2���τ�?��;�ر�����Ά-��g�<m�BP'�G��w*�!�|��j�s*����ѩ�p���@�h��rkm��b��}h���\y{�fGw��k�p�6��lr�"�1WHk���)�?l�0
�j.-��q-B��B���=�>TJ���Ro"= #��������d`R,��ư�6Wg�:��]^8F�����.O���1��1t�d��9/���By��� ��،��C�J�шjk�d/9�	Ym���PFm��[�
.��i��j��ų;�?�&k$����-v���1��ؚ���p�����Ցq4�p�|m�<��i�VU����@ܶM�5��uIF�F� �2t��iDx9��]��~�*v`�ѝ��R�����+!��DN�5��ӱ(���I�4���<���E��:S�A��#(��P
�����~��!�o ߔ��VJ#�wl�J�j%�R�y�W��8hɞ˹)��zMi��S�&��B��	�i������e����'�"	�D�m`"�X�Py+����sM>1��Q���C/궷�?� �š����|��n���A��qd�wP�9J���$]+��X�A]/
���yۏn���G� �|��;�pB�d x��em��ᔑ�������P���s�g��B��C7�.rQk��2����w�;���5�]���S"� V��B�1
�H�$0r�S5XC�(�z_|lO���˚ܬ��ڝ�,v� �&W�8��R(mW��0ږ�%`��!��es�	��A�3g��4��8�S8aП�����f����Q2SeL��&�o!�X\��
'��[��0�.4�i��MYJ�C��A�sݎ�fpf�/�]����E���֚M�?Z����Lq�	��HJH_��f��Þ[~�)���wP�&Zu)52�/��������˰c�]����SÙc�<���5�yо��0�����av�8A,L��Q���/�Og��lX�5�L+�S�OxԄ���\���8Į�����m�sS�g��9�������ʳg'��B��G�/]�22��YX����yY�rh˂zn.	�d5�Q>�f���̘R�Ӹr�.���l�^���2}`�P 6�a�2�w��P)���%�0U�	����:�6�K��>��8�cd��
 u��pA����
G=N� &q�T���!GD��ʫ|���1E�q`��<����.�� mM)q�F�X+ֻ�tD9�������+6_rW�/cƟW��OŚvKr]I�h���9Zo��Q��Ȉ�ǃ�R9R!4�F���H��ѮS�#�m�"�%�I�	[���u��.�}��B�P�\.�Y�]Q��p4��n��-W���'<�Ym�w%�B��VН�,��XAu��c����U�=�(ܨ]⟼BE��R�,�iB%�3��E���E��3�R@���\��l*��3F�M��ك�vU!�,KJ^�O1��?��N�e)����:(�,��X��=��"�Ə���5D,�����������)� l�6�t�R������pg���,�V3���u��?j�c �z�� ��\�9䋞>r�K��'`���=���ha���ԧ������V��mV\}�X���mF�q�B(P�4��Q�u�0��pU����O.vB�/E}�D��˝�K��*��'�b�*�����������U��%9�HS�Y+�\+V83�)��[�ǅx,-���K@V��O�n.B���m�˨�r,Ci�u$;�c�O�y��W�
x���V�x��`%�6�ʦ�9݃�P��l���U���i���m�(��XpEx�a�c�
��d�9�S��1�!�
��b�d���Y�f���-�LE�k܂��kN��*.�ZU�SI�]���:�""�2��{ ǖD��sT�6A5���l�wh�pa�_�'�(o�����.��.q��'?]��ӀҬX��S��/�����rլ�� �}}c��Y�-��f����+��Cr��ҳ �I�E��+N���LM#��g��x�k�m=y�(���}2R �=�c�.=��H����w��m玅#�3�o�-<���K��_�*��@?+��$�nsl1�G�B��fj�0���Q��H�d�n ���5���"��C�m�0��u!����Vu�!�̌�DR��X���s�l��s�_9g1�Y�]��L�u�ZfG0JH_/�Ʌ|����Ht�����Τ�"(�lm�Qx�^�/c�M_lװTsU��t:vC�L��~tĦZV���#1F�HƁ��Y0�����M������@���/g�},���坭�'n|`���n��&�>��>h861�s^Ԫzz�Y�V��$�N���r�J:*�^ƗkNj��<4�hS�-$�ȓh��V�6/K�b��\o	]�E^K�4O1p��Xz=?��ϐ�A=����X��(=D�ǽ#�7��r�o��U�5H���q��"�l��wl�osL�P����_gҾ��D��ԫv�$�y��{-E�H����j��s�x���lp�+5	��J3¡C���.�)������@���ZU��L���q6*^�(W)H�.��9J��Mf��� <knJ��3鉙S\�"��{�?�O�y�}��0@�G$�0d"������Y�n�h�� ���&�� _E[���z]�$Vt�>2��{ѡ��E=˓E�:S�Jx},>'#$/pJ/x�-�f�>�qZ���W�N"��yz�P���~M@B?f����3^E���D�|2�x���G߽�,b�~f���@-_U���P�3y(A�A�$u��u��H�_�#G�M.�shN{������#�kõ]~П"�a:6';Ǘ�]J�T�8�3���+R:0��g�!��p��4�WV~�OT�<�s�;M��۠߻�\���#��Y��2P�*v��_C�p �`�7g��FOߠ�w���aӘDUAA�+i�������*t�c6��F�zB�x��,Z�!)�5�'?r���<�|�TtJ/�c�)K>;��q�4c�����,�D�v��u��ո�%b�yr�ܾYY������P
o!�V� �1(j��j�e47ډ�y("�4�D&�j��\Ʉ���{�z�Ɖ�蜜g0[�-}������Ҏ��I�`d��J��I���Q�9ˊ��/�bA��Z����-��V�h��dk��>�t��?�Rχ�θo'Ň�Պ C��e��MjVZgȶ����]��0�4�$V;�F����+�rW�\Cw���2�{���B7���GD�w��>����1�ȟE=16�
�4i}6EF <J�']0�V[Ru����B�p�H�e�>(y2}����a5�{�o�Z,uZ_W3�^T�^?B���k�Ւ�����j[�	H�lwhvK���ޗ��ӷX�n.���o{午q5h�k��jI�����A�ן�D��:8��X�Kt ��BaW:����ý�d�SS���D�Ս��:Y�=���-�{\����j�vU�K� �'�r�>�sVAȦ�R��TE����E?��l��<�/��}�L��g�o:���2�&,ʓ@Uu P��,�S(W��K?��~��OC���]�d%=oP�17Yv�)��ii~����ғc�
��VY\��3*_#_`�|kWЦ:�$Y��.T�,��A��ϫ��:�l��u��JܢD�HD�7Aߏ��q�!���.�s�!,Yއ�&t|����:��S%>*�;���I�|DF�ݺ�D@*G@�+��JTn�FQa��qF��J�O��)�pww���|td̻`TSܻ�+�����_ӷl7R��$������0]�
$/���'*{X�`��u�2����8���7�~�v�M]�k1?�p!C�d]�#�D�͎��M���7�)�l����0����ʞ����Fh���2�~$B����&��[�J���*H�m��q} %&ec�:�#��nh�;�fá�&��5�U	����\�\H\7|f<�a\�|�c���KR��S���HY�G$E�b�S�3u��bu��<H��y<�f�ʑ�Aܙ!���	�##-���0s`���
������w��b_<��i>�Ͷ��D4��h�	�p7`߆�Ӈ�n*H&>)����\D
��p}���',�d%���T)��uY�����B8:�p3y޾d�p����C� ��=���6����f�'���ޘ�ɍ�}�v+�fu�\��A��nT��Bm$��p�̯Z�����f�/S=t�2sY����#˰��2<���o�L>2�ѡ���޵x�^܉"�I5_��߈M��K�����\[�
֓}���,76�����b��Z��̵��9����C���n�04��Dsȿ+� }KJ���A����tA)&^�V��DJWͣ�^���m��6�ѕ!��< d����>��������e0���aW�C�w�n�}b(�������܁ˈ��A��t�A�����ײ�mO�axB%n�&m{8�l�#+�u/w��!'IS�a�dKq�[�9��a�M�ZN���f�I��^�
���"�����To�Z(s��z���~�4~1f��	�%��!�)9=��}kS�У�`��xB�s~��f��蚤���ci�^�;W!,T�P�/��t��x� (V�'O�Β>����RH	cV�J~'��M��S�<� �fv��Kn�c0�oYsAp�~��D�RNC�,)N�s�/OR�A��JLL����^J#j����������0�m0b�SU��f����L�'̝�Ɨ�F����n-4�Z��ٌ��x�a�ec��B�M��w
l���FkT�����HXU�m��Z|2�`g�6�O_���?�&]�@�>#M�X�3�Ǌl_PChV�W�;�rC���������ߗ��o~S�����\�9&p�X���Z� L��IsM��_��
�X8Op
N[8Hm.��Z;���nT�X�֪Y��@��M�D����k��^�'�!���?���l��f�O�9`��;Q$(���?���|>���wE�
�cJk!H�xyL������ߏ�� ԧA�k�}�^q�Zu�����ZO�P+��d�?'����z7Øe6NPL"������Ήm�4Հzq�q�Y�f����`�v�.��;-3x�����2`R�j
��a.o�'W4�k��WV�o�t\Z�>��k��+�,�=�P)2*�ut
0E�;�_w!�(�?or��ΕPڻ�a��^h��k�>���=]��z ��qdK�֏�I��ޮ0�pN<����l�4��!-�J��!P��X�h���Hλ�j�sf^2��7����4Ll"��"��5֎����v\����N��?����d?�˹�k�ɷ{c���` MmDK ��K� �y�~v�����Yg~�E=�R�wN�4r�U���N��zԡ�~��GV�_���"��n�	0���	]_ �����Kz��;�Q�_-y�ٿ+�:�%�惻�0�����%�+�}��S�������6$�G
\xsT8��a��J�iIq�u�]��؄�RD�\S�UXq>��=�۱]B�玤��d��cIziȊ
y2�>j��p�������/�?s�9G&%c����ӵ��2�����:�. �(Sq�L�=17���g��Oa�����M��b�n���� T��\"������'p_37�˛n#{��z���උ��I�r�vDɄ�<��i��EET�r@�>Ob����GmHͰJ\�ʹ��`��܏��`����Wi�G�<�[a�0�U�#����GD�T$�n���f�,���꿗%����lG��|����y� T�s��Μ�-,Y1}��n�`�-~>�n�x\ C����E0Gn%o��#��+�&��p�.��Q����x�5o~Gv��62��+�w�Z�������	��L^��!5�K.�	����^��h� ��n���뎅���S�y��a���m?�&���,2�l�VN���ː�^�/��=��ق�2�u>���v��nf���q��G�8�h4���܆:ٯ�4��y����������&�����L0:� ������T)�O+�)M�����/���)l���oG�hw�L�_0˽VHޞ��c�Zk2`�2y�oi/\�R�d���v��
�|�7AA=L����I��!���h���$��u�iZ|l�Y��o�=O�ч��!��سA�+���8�̈́���,�`.����SJ�G�9\q����l*4d��������w�%�����KB�z��u@[�l�ՎR����P��2_�o �G�h:m��W�@�r5���v1�!&�ܰA���`RIz#�)`.+��j��o	��bw򳐂3w�ઌ1����pg[��(�̅���*�Q�hy�XO�����F��O�-ü X��<֜��2��ZƋP��q"n�i�a��u�0�Q�ho�].�w�^��F�q�J�am�V=�|�q�G�i������:Q���܍s0]�������e8!'�t���9^8�c����K��sI6쉙E���0ZJ��8+��Ms  D~�R�]&־��P������\��wWz�?�>
�*5��%	 �dW��lPif1�
 �`1l7%��$W�1U;�쿂��o�zn�c�h�Awi�=�(:� �ĤaX"d����%<K,��I��ZH���m�6�,�ȮU_�!d�ECwe��1|2�aʎ�w���'GZ��$f$RD+��~���:	�v��	�vn��3�ݑĤ8's#H��e|@�R�j�[�������R��'G^���h��n��`7,Y䀳8���y� $�=|�퓬������� 3yȤ�A
���`�j�n�@m��;�$sR��v�}���RF��|4�,x���@ �yX��u�l�H�OD�������!I�b��&���p�uMʇ�\���{�%U:{[+M��v�ω4� '^�e] ��M�����ݴv���{������"��#��ZE;H�G	��L�V	AMJS:md���&�vO�NE�䯖��@>�r�,j#�;*z1�!����yݾ��D��>�KH;�. �t�	����\�.�g����h��{� ]���V�ެ������ ���y��όl����i���+R����ѻ}��`H2�hJ��M5�2��X�hy���"8��-���>�` 4պWHX[rg��=����ʽ!�2&��IGm徸�!�ߩ%��ì;Us.\"s{�' C���Զ=�j�g-%	�T��㳉�
3���bkE�j���ʷ?�ԛ��S,���R���?9p�����0�x�V �̆��@�(c|��j�b0�0��:,�7��ij|Ik{&ikR��2F!���sB���>^��%��*L2̼�Ig`'�g!Na2v��t��!˵�]"��DG�n����^D]�\!M6�^C�����Xs�1����O���.#��lF����°�-����S<̀i�?Zqe0�"ز1�s'��fƂF� �F ��>�<E�	K3#'ՠ_�V#	'4U�}���ߔП,\�鳟�!�`n�/�ƌg:��4��5.�L�)3��6��c�ZmzDT0D{F��x
a툾��>�
�2ɫo7	���(�a[`�?��T0��I�*����2:S�Ә1ϸ�xf3,����	��uTiˊ�i$���N�G�K�m�Q�`���6(�zd�#ġ���p��_���	e:����������<��L�T�?�r�
dW?͘k�%b���i�)N�?W���`z�&�BD��b}{{A�7`h���Z;Q�7.1�����V䀼ԀN`�b6�)�m�*мaU�~�
.a@>ז�xI��V��."��4_n���xyT�]iL��I4�Ss��/NZ��ŗ$��%7>M�M��2	Jl�O��L���lG���X��#T��q��*y��x��󽵮�E�o�ڦ�K|�L3eV���R/"c��[lE ��-ĵӈ���rR╿�K�s���o5@gz��x��H�ݞ�3d�ЏzG���<I>"L�� UC��~�q�5z�Q�v�.⛱G��C�MVs}x�>Ў����~Y���w��_`WI_ i�.�z�ؑ�Y��
H=F��t�KL!�����&���E���<�+�@f�D����C�
(ϰ����<)�q��@#�R
�[�K��舁5����q*I�nYi�L��"� F#>���j��KѶ�݂z�U�J�3n ��������ER�������Mt�9�۠7��0����[2���o����
�'B\.3��c�~'V��5���Q��T�/�Z-f��aw���.�ݹ���˛+.���p�P�RA�u�>�,|�'�/��ɺMX7m��VKt �e~y��!˽�v�_�`D�.�Լl����cڳ�B4���b��Yڡ2�^���FI0 �uù�$�Icg��B�v��EOk���,){V��Q��Ae�8�|��X��s+������
��î_����@T��V��0���h��	G٭��;$PI&�X�!�֙���@NS�%�ݟm��.r/E{l�{{�&<�x'7z7l�HfN�,��x���16�dȉ]P��\��ѷ�Jq�L�6�m���e���O��Jw;�9q�*s��É���.��oVG&Q8����v�F��XV���R�a�ݪ�4g�]W��Wy$2�ʕUL�"!!'���J0��٠�h�u�1e���E��pd2��ʰ�ݓK]��J��n�ݙ����J�),�ʻD�V��J��	���Y�f�Pa7�X(L���Ԋ�u-^�r�?��#����m�ARN64�L�Et|f*���Ä�� �Dm��K7��<@�-eWh��>�T2P��H���܅�m����P>��r&�/�ғDĜӓ9�?������B�<k>�љq]���(���
���K��<r�/�T��]�t����d�Դ{j��b�'#?k;0j,n<D$�֞��	>6�WW�F*ڡ��u;PQ.�P�_�� �鯸J�Q�e�9�b �i���[�>�NY���ڳ�i>X�D����-�Й�Y��f2c:{�x�k�sp��"�}GXvH�gm�׭�Ю~��`n(�e�)Z4%#M����wzfqU�B#ޣC+ob"*��
4�G9~�!��Lr�g9��R���Z����ք�)Q���2��n-�5����$�a^�X���C����e�&sH-����>^�ԏ����X�Z4�<�k,�MdH�J��Sۨ��D��ԈJC��Y��~~��
�:�A�