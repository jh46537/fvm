��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&Y�%�ddؐ��e<L��`Ȱ���s�M׍�P�0�Fd�?����a�!��N�QЋT���X�~��%�Q�[�;��#f�o�TqkMN���I����X`��k��Y	�IQɂue:#��y�/	�{�*_]���a=Z8V�: �4��V����'�z[��
�/��>\�<V	`E�l��UI��ZR���\���H����� ѵ6kG+zY(jY;+����BD�B#T@�;~<A�}��r�xg�gw�F�aX��헆q���A%�ee���1�1X^�qŧ��v$��W61���4>��h���uj(��K�@��-Fz���M5D��bu3{z�cn5�j,/��ښ�� ��c�I��Ud��J�9A��A�ڻg����К4�](�`�ª���(�<R����'�h����{��ix+�ٰD��zk��j�pc������]^`I{s�@�j�~�-oX���a=�����#�u����� Awn�Bd���`���������iz��X���\�C���g���J��Z��sA.�0�|	�p��u[SΞTg���"EO��w�Dv2&Ε�F�f.2)2K_ӆ�%�«T$r��t�:�"�a���괟&l0)�@r :1���ɿ<��\�n����H�A�;�
��<NRrr�Q���Y���|�J�,{%X�Բ!į`F�Ev�Τ�'|T����⨡�q`�d�}T��/�g�z#otj����h��u�6�a�
�������{B�#ķ♮��P-�_k�D�}閦5���/-�*M�β�n�O-1���sF���[�.pGIP��@ג��Z���k��H�u<x�&n��Q�=F��爨�0�x�g)�'�0a��;�դ7ʬ�`7f��m���/�E*:?����cND	4l������kQ#�Nf��րL�a㧟E[֎=����6O/J��>��Ru��ԭ�[�O��NFm���y��{(^��!�˻��#a��1	y��E��ǯ�`��I�s$"|3���Q!��[�g�D�<l��t�?�.[{hȍ�|9��͠���N"hB�%�TV�����U��Z��G�m���r�CQ����=vס\�v}fL���e�_���JiF����W�����/���Wc�������;�`��i�#3�*�b��p�yºǃV�Ԅ$���lD��9���0ɽ=���8q��<��:�1���E��}s2�tgϚ��1ܛ[��Z�2�h�����A�P��%	��,��s��� �%.�����R(�� 9X�aD��j�QD0��:�p.sS�-U-��f�c�������2.EO'󣍙3�w{!����4�]g��a��N��aBU�C�c����]�J�a�lhBK�҄[#����
���?�"`?� �Ȑ9�8e���xm�A9n�?�ϋ0� �m��{4 Wl�K�1����<�G �����f�7�D�t�ү�!����Y���e��E��-��ȼAW �A��P������6���J_��8�➫\=r��Dq���@����iRq��m�q9h�]�fps��m��Xa
�L�Rު!����&����#���e�)��#:��5�!,���9,�M�c�NNĝE!�[�݁��-1�Yo�il  �u9�+O�@V8�ٌ
+�/Dp��g�?�����-�G�o�����T�4��R38��=1�2ā�{
��Z�:�����e�}Z�e0C��i��[�0��2��.���c��qM(Fwt
�QK�e�L���?��CXt�
`h�D�S�Ȅ�~����Qʭ���"�ᷩW	Uo�S�%��Y
'��J��o"��<-�W�����u��ru:KX�ȡگSSi䨧��_�Դj���S��<���W���G�=�S��\4�6'�� Ц�XG���@��&�%A�YQ�^#V)�����!F~�!s��|�d������1��v§��\9?8em!y�^�����T�iº��@~͂��S�ԏ�	�g�ύ��Ӟ���7#�K+,+��<Q���-���6��2)]p
��L��'�[��Ҫ쿖���ֽ���F�����VY�X}�PH�����8"����Y$h��G��H�w>��D�~�	ߒ�V��7����Ɇ��M�"�ߞO.�520kh�HӐ3~ٹ>X��GM��̨  ���)��7�E�}��P��p�*-$Т-�TDv +*�!�#"��N��]C��ICj��Sܧ���@I�rg��J�2b����[ɑ�8�6KH#�ؗr}��q=)x�����u����q�]D�P�o���Z�b7�o=-�箕�N|�vo[ؿ����"KM���~��]���-2��4���O�ql��S�J�����������ԓ��T��K
��&�sh�+�����["��}��ݦ�@�mO-|�h����DSx~��D���O�����-�UU-.O�6�Evk���y
��k�Z�����P���/�+c]i�9\�c��GLW�w��GF��hxん�t-K	%�@���b��e��p��Oъ<F�P�?	X`Y�(�癝����� �ٯ���ag�S��P����N�=G$G����>w&�%�O,mJ�D��
޶�Q;��W'����H������_	� ��#j���G�U�@CI5��XA��ٛ9 t�ϖ��a����ؾZ`$<�\�u��d'�c����[á� �HF0�e$(�����������x��?���piO]��mbd�%C�\pH�@Y�K�ۍ!M/�r&�@Һ^�V�l«�>|��!��2�,-�Y�J_�����p|�������D���΋�]�p�w%����dG��a5|�^���yǛr��C˶����,R���O��;�;&zs���,��#`���@8* `B�����$cA^_��0JI\�?���X0���Q�ђ�����g*�ǆ��Y���B瓱����^$%+*[9�J�Ca�!�8W����KGMݣ��@�|���!���,��>'-|�'�#��V�P2�E�R�4Z�I���`k�i����Ć�n5�ud	9��3�`'S
�3|�WݫZ��;�gߕ���]�0;�[�rЊ����qB��1�~��iS�\UN: ȿ��R�Q�,�_4�zE���s(�@N\�kB����Ò��.'ѭ�l�Wb<I��L�t��.��j_�"%!�\CL띪��˅h��>�	d�a)�B��L�%�7'����79�	���$�Ç88N�T|Hf��Zg��}�P}$s�� ��i*$�F/K][�_@;P)�)�
?�����,ӣ*���p��B-�Na�	v3R������*�2�}��V��#��p�Qe֙&%�g���`��g�RW4=t�I˯��:���E2��P�Uݛ&;�-�ʬJ&E/���`2ʛ��G��av�3+O3?�������܍��?T}�3Esn�I��QX���1n@��K�k�v��L0,���
�ʨ׃���\�X0�l��B^SĠVkQ��<c���|k��J�H:�H�I�/
��ID�g[�2���kT��x���Y�?Nn%��%��&�LT���R%�d8E���y'I�_�+�r	3��}�rű�����k�.;-G����ڏ�ƫ�7�dh�� (���P��I�ڤ�f$��[@����)���G�M�my�D|���v�N>4����4��Jp���6��񲘐����
��9��όp����y��`0/�:/�	x��u�
��B�C��G=��0�86y�R�C{�~�NTK�X�J�)��>�p#tb9�U���>��Ee�J=p�uJ�3٠Ξ�I�&�0���ۄ@꧀D����ת����]���d/�Ƚ���u\W�Cܯ�mB������_���Y���/�}|�Zt�����/�t�s9 ���pU�����f"�"7���9� K�s,j�VG�hz���H�{�&ƀ�KwsX�c�b��0��9����ȃA�Q��^��럇7N��{� ȺG%��@�<Z�e�%&� �-Oycc#H��I	�-Xge\�"̌�׌]�ɫ���\��m��4S�rL��3	�G��U�QkKdAҙ;Z�< b#bH�0=<����m�wě~�uo(\��Y�>]���]���V�<�I(cߒ�k��a6A-0��β�s�bS�^�� EDC�����m��)�D�2�{u����;�2��>���w���N�1)&P�Bl�c�lqA+~Y����2=��H.�x��+ M��'#�0�խwFJX[k�N�H:x����d	�a���N$���5gR�/���8��Q-:
�v��/.���}�os�[a�zH�o�vAm�2w�a�Q�v������d�'��MA�Ԭ)Xn(c~@���!����i#Π����.)r�tP;�,�����܅�w<�U�H�x%�r���Pѡ��_���|�$���%� f���Ƽo�Pܛ	��G��
��!��Z������!��	*.�t���y�5,�p�D\p�6�gE�du�^�����#HzO�X!��E=�n��T��'�T���� �[�e��� ���#:T�LÈ� ���2>7<��<QH��ʃ��0�
�r�\6��*-qhɒ���������e�w�ž�A�֊��c ��������m��27���r�Ŗ����:��`���*�Ɇ���ad��{D����?� 0�d�pr�ZR�3���Fɛ�"�ے�������.�5�@����Q1"��<����1�]�+
wAa&Nn���]�-7,
�bU1�����>�h�_�;B݉���Wu�%��+�W�_$;�c���@�\����p��O*�� L�RS�p%�S��[sA�- �R����p�w��Y/z�V�R�g��ۆhT읎��]~\r�3����m�T<�*6���<w� �ӍE8�9�W;':ƈ����%BحB(��J|.�Oa�����x~鎗7��#�S>,�z_Pɨ�6����2�9������Pin���BjzUB�"=�=�I�$
iȨO����{�g]f�wZ���?'�Rƺ,�a����\�D'�o9@�ɪF�JL��^EO��R2��Ysm$���=�g�S�yF�U��:%����XW={]x�s���� ��u���ft!�᥂pdmW#n��V?4$�F��9Щ���<of�n����tq����ڜOh2z��#�j+qC�, L; 2t���}LV�6�sa�UL��y�e����CMR͠��um�<k��h�*M�F�čC����@��qN����5\׻%`�x�-��AV������_��PTvy,�)#�knS���p���>9I��g\Q��"�R�aS'1%X��A�هw�@6�(�O�˗� 
�
d�re�=6�����q65]o��j�b�c퇫%c��.@��U�UM�S�Ƕ�Q�}Z@�Aݒ�^~;,������s<O��� sNH��*�h�2�G)i���2�i�4gN�)t������m!��K���������2�Q�;gd��aERi5`֞K#b���oN^�Hݥ�(���Z����}_x _lh�I���N�vz�M���;?t��ya�ȧ��t��t(8h�5y�x`�����w(~�j@�){�	l�ӂm(�($�s_jz��$�4CI�I9��Y ��{���G`�\P')~	o:��ļ�d�XJ-��ؘ5e���;b�������g#��'a��*)V�:��m-�IN�^Q:{�EmMo���L�$�]�R��S�§�����j%�c�)@[,����
�p��&O�{�$B�e��̧��xͩ��3w�˕Ym'n�@��-�������׺^�����N�p�Ks'��P��>� ���7�@<�P� �����M�<Iy�֡������WKU�l�%��%�w�H6��tA���'Y;��j�vb�]e�+����O�*X������Fdܑd/���v	^�nlz��f���Ǳ8M�������]�l�J�5��B�i���D	Hqڿ.��V��D{4��@Þzi�W�EɭW�DtC8�p� �G.�b��r�ˁ:I�\\XWid�B�0�l��۪QZLi*�Z�'�D���~���׮�I�+&�%�_.��0 �BZx���Y��\�����^O����r}X��H�)�zX7I�q��y�Uԧ���
L!�0�t�'�p�>�N���Գе.x�=wE����1�"�8����[�Ŕx�'6�:C�_�N����
*�#��u^\�U$�S�i�k��E�&<�ݨi���h�e���oR����xI�E�V�&$��5R{'�c��O��\��߀_.�C�#kd���?���3��)����+�9r�j	�_xc�2E�8?5D�ē��ι�����9� ��E��2?�3���l
�r@�O��mp��
k�!jT���*	8�t��T'������?��Pr�MoρR���^O{1�>=�?�Z����[�99�"`,d��1�c����¯��M�'s��&�An	��JM|�`�M�:&����3f�^�S�j�A��6U.�g�X���q���3�W	g����Јt� S_)����0=s�Sx��F:�@�=O���|rU�'�P��TS���Ȋ8t��Pz�G�Ր�}q�m�����"����ld�\���k�sM����]*5pԱ9'��{@`c}=c���$(�}�v�Z�H�!1=� $|�V�A���YX�A�z�NBV�g3�?�4*U�\9�4�,S�}�Tn?ٖ��rv�^�������e�`��AR�-�!a���w��X㧋����+fx�	��	�	�_C���#5�K�/��Mc�;��1%�X����G��ڟR��TQ��?���95��gv9�����-*��6�'�\g��c�p)����YѦ?�Ұy<D&M���-�s��n��$ޔ��|�W��2�.[�]��f���uG��e#��?j']����g8�^ejo��C^����
�Ro%2p�%j� ޘ%b�U�|Q�ËZ���4(m� ��D