��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<����d3��i��:��@:$���;��U��zV>���=c��Pz�z2��`�����~�צ�\p��yp��]5k��q���8AK9K�Oj��� ��n=!h�*�N�b'��Np5
� D*ْ�A�Ԟ;nz���5��R�9�kͺg�!R��)���-�{ڡo!3�;���cQR����M�c�I
�n�&�ȟ:Fp��o�%I�L��k����ZcFW��4�)�3��c8f��N����X�̮��l�PS���sKC6/��an��l����и^~��
�^luDE<�g'%p&��"b�����;|^&l�^S��U�A8�Ź�x9���HՁ\Zb1$��Q���A�Վ.�gtB�l�w�k���a2�e�����;܄�F��v�&ZJt{�8�YL ��ID�gԅ͵��j�fI����{Vc��&����ƀ�Q�s����_E�'p�j����<G*����@��"�$��:�a�ٌ�����F�Q	����"�|K?�K���LRN}�j�:�ڢ@��s\��<j�u
����(�~tB2�uCC�l&0�1�C ���4��u�ym���$:�i=d36�k�g����Q7��T��L� ��p���a�TD��5�\�j���Sz��ʣU֒Q����]���?V���y[�j)��:#���EB�t���=y��6y����i�|��G���G��"�L81p�''~.��~�0df��U/�mb!�\'�6t��\�+�"Զ�!žM[�k��;#��+����*��
�������߭�M�:�� ,�����a�����Ԙك@���t�����`��J@�-��ISA�OOY,�؛Ų�w�>�_�p������H�����ḣ�x�S�Q[�B��W7[ܞ�3j�j�Z\�m���l���oq�=��qo���aLZ��fg���D-��WGԹ$,#�l͟N7�@0e7f��������?��W"s�!�h��	�GB_��Z�x�S�;ekc��ݼ}�!UX#>M�*6�`����L�P���?|"�w�aJ��K�j��ߠ����(IE��ܮ��p�HRlS������c��>�ʼ)x`}�"�f�:�(H2k����,���J��ݱ5��K��Z��B�|�۳os��O���h�5����|ԩ&��݄�m	)���
��o6R$�qJ��Mf���H��̴��MH�[�(mñ "��U���~403"gd���]N%�'{�&I��m��x2@�