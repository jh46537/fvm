��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,���?�a� ����$���HY�P�'�~��p��+�6^�EUu��
�P��89���Xs��	��C���׷)w̼���3-��iG`]"FTIf_"���E`ѭXb�bk���j$�{Y�Q���8�:��R3KQ����6>�Ir6bQ��74ѓ#�/���f��g�_���cR��'�Xk�&Y�v��Եs��+3)�I�β^"�n���o�ޙ�Oa\@?_�@n����s�-�̹N�gx���a�'��h!�k7b�@���}|�J��zp�YU�^+A�j����3y\\ȡ��7$6��E���0���:� ��s�ܡK��c2Ch��&����L,%�i$b��_�zb�ojx�R���iI�i�F���d�)�#�i̧�vm!@	#���Jc���l��t��y�~�>�%Te�U�y��*���Y�����-��~(��J6�1����F�;�z�[�-�uDg�!��U���	�[Z�v9��V�J֍��	}�����9-��j{�:]N�h3$�c�o�t�c*�`U�.$�>ڹ��ġ���YBx�r�,(�<�Rc26��G��Q��t,�q����)O��:dj���U!�v���~y�o[p�W�?uH	��:��giN��,���! `c��"&�/+Ӌ��`<�dߘF�S��,�!�/&�>�My��j��7���^p;[�~[J���<3����mE�m(�ص�Q.����`���'P��O:��w,����DCiJ6��p����m�G�����^Q[a�ʍ�����Ǐ��(�������T�A�k�T6�i�y��/��m��;���{@8�@���V�Q<�|6�qyV _<:A�PHUw3�{[�����ט�ٿB��\V:$���_,�W�-�%�+c���l���$�Pĩ���5}�2z�
��2�Fܭ��5K�7.�;J$
(VA�e�}�ܩ��H��ⶈL�SY�1�Q�����*�� !؟6#Qc�}޴Y�׆��*ȭz��P��d����ӫl��i5���	�I���Cg�K�B���ۼE(L��������J�����ķ�1F��2�>c���H=ݸ8>H�)H@'�D�"�� ���{���������*��٩�Ԡ���#^҇b�.J�&��h+���C�B��t�j���]��V1���� ]��U�aMj4{�8m�B���p����\ff�}9-k�0X�Y���bA�\,��B(sq� Y	����>���h�6��W�gyX�0��5n}�W���n�P�OwRL��Q�4�/v"ݢp�+e�H�R�vj�?��?��KB^'Bm$J�-p����,��j�±fln?��(ha�䰧������QR�|�sI���:���%��G���8s6/��V�7��!\�Ҥ��MV�I���|��8�p�� �z�5F��	�6 �8QȘA~'�e���5�p_O|�P��B.BY���mm�B:0ХAêY䕷�A��}��;�z���X��[���	�������(j�L�!����_�`�}���ϧ�	�Z߹S�YB����y;���F�ʕ	�����.�X���7bk�3E忆��=��9��ނM����^	��w�J����#T"$p[,�& ��V�!�Y���h��,�v9J׼�S�V�����8������e�:�m#�X*[����_?l#�������k4�dK?�ے2���ؠ���7��~&њ�@#җʹ2{JJt�T����N9Jg�<����dU q� ���_"�v��J	��,j��Lɘi� ��7�G�li�dK�.ӂ���Mx`��8h3ϏV�]�k�'!5%�.n�
i�G&	[CU7pC�(���i>+�}�9'1����NWW�;����Y�B�7=G$���rؙ?���3j�t��WR���.%�h�s��G���^f���AGS��J>�0{����S�E�JWAȧ4F�7b�n���$��K�m-��n��q��S��;�=�?{�@h��B�ϑ���I�*��Zh�����c�9�૲�9ܱƂ��-�J
�gm.�S�b� ��rLX���z��w6�̇�����y�K��e�O���������^��*X�W���p���;z �4��㥇I�9+�