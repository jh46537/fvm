��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{�H|��6	x��:Rg�J`>�gPnLG-� �Ÿ������l���K\Q ���=������<�uO�����~��+V�	Q���K�	k7;�T�µ$6�r��:��7���"�Mh�����6��/qh�q<(����4G�
AqpÌ��3ŝ(����=��6�@/� &'5�="�@#Q���|�@_���*�a���������&ؿת�Ӵ�$�̟=�J���ŘgOE��\��k�>ɵM0Tp\��`�`��8�~C�4��c PW�R,����Y��ւץ6{I��o���$��jtϩ2�u-*p���?���4nz��6�$�ro�>�{���������sv���Z�`	��&���ج��*q�*��6=��s{�9��q��Ga�̦��z��F6c�g�p
�@y[#,jl��H��)T������q[E<����ά'��"�$�0J�6�����;�
>��0��0�jȨ��������ˇ>;�1W�j&tv����?P�oF�)Cy��j�'�ᕼ�IF�h�@	���e���;d���h-�������5"�%��/Qp���Q�說@��b�7,כ�O�!Ç�:��������5����Ùą����W���w����K"�85u�,�Z�T=屹�s0�n�����_)Rkӡ"����:�E������dim������2��s���;��E(Z4Y�Eb��!�)o���Բ��0�*i��v�ԕ�]s@�HQS����
�gҿz�2y�-��V8��zEb����ǔ��+B���J@�>�,D%�^�K��˛�UZ��掵3˘��i�%8�wo��:m��U��xl�A!��Xb�<�p�y*�o5��k�0��U	�p�,k�n/�؄�֌U�C��K�񇕳z�}B"I~S�- ĵ.v�,�kT�=&����F�Z���O�
�٨1�/BH���-�R]��eԝ��r8�<Ѿ� �;�ˋ����|��L���t��zc�E��t�S���{pt�΀�p�C�V,<�/㟧sPg\e)�ŋ��Vg�i���\�ػ����I�s��W����Rr���\��n�?����}g���ʍ���w����#	A�P���u�[m��x6���r��	����g��3��l��~D�EH�s����@�Ѫ�&�IBm��]u�oN��a�oQ����a����~�9�?N�z�{1>-_e��2���h:,z���Ez�=M��ɸ���WgK�G�O[9{�CǱmu�#��۲cFa`�M�PyuT�Ұ�����@d����À�[(��7�^Ɍl�_�8�̼K��p�0U��z��"�����<k��"=������o��v������
�{�u�f�_ �v��I��4�W�qeV��7TQ3�����~�p/�b�:z���(��y��؀Ǖ��׾���`�.9���n���W���]��\I6�v��_��[�����`�e����w{�.j�L j�"����������<�e8�Y\����L�^TP�������39��0	�I�����&V�dT�n�����`�����[�AQ�fE�l��v��>�ڮ��dM�R43a~��u@�WMh���F{�0����O��0r�p�u�l�2S57��*M+��-9�&wb����K�0
c��d���}�мFi��(�-����K��j���ԛj�����;����8m���w�����G�8W��F��L�ñ:�Kc��/W��/n�m=�q�Zc����m�y��n
n�:s�1� L���:y�;��0�isA*��lԾX�`S�Wg8�N�'`����x�'�`]?7�$��pk�"��5s��?ܠ�%+�cJ��T�Nx�=�^t^�t�Ke�&?\�b���eY��W࠭�U1�t�hx9 d�e��4h�	����%�V3��4au �r
�҄eY��-=.]�K��a똠�醘�a�*�!w	������n�a.�,oRF��/��hhZ-�К��,�m
���<�=�kA���������`�J�ަUnM�iȢ�-���r�:����ZFU��`�v��",zD0B��z�j�6���NL��L��Ym����ba�h�����;��=������.#i2�u���a��d`�Ƌ��W��A+��nB���fCA:�H����^|��u���F4�SY���@tk+�us&A�C�9�mR8S�ʨ���ŵ⒌c@gʁi�R�P�K�o���?�s��ȑ��A�l3�Wr&�ٶ�h���ı���᡽���Ȃ�YRvbz(�>[=E�l��<�*�iX}��:�*�|��C��H���R@�ۺ�~r����Α7��ݳ�S��l��:���[�����אԎ+���{j_��VQ6\�baڽ%�dU�8�u��N�A�ֱ��cw��:r`�;IP`���ҭhd����d���.���D~���:SA՞��?�(�`lm��7��F

p��ıW�j���p��X�ե�e~��:9��U)i�_��6Ē'�M��	���C�\K�!���m\�Ee$���j��
4/�S"1fl��5ud�qM�w�V���9Zä(���<�*Ɍ��+g�F���<�h��]��P��00S���������8Uވ@R�8�ē�'& ]���?�w�T�!+3H����[�2�̸���taZ�k2|5�!k��ucΚ��7c�'/�թѭ��N