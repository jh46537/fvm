��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�Y֢�08)��k:�ث�����$,�:YƚN�bK9�p�IV�UC��$�Gǣ8�yF��D^��a5�{S�&�`l��ve������ӄ�d�=lے��+��j�Y^z�]w�#�k����u��0�]v���ޓ��#N�ݔv�"�GZ��>�:��I��
>�c��6|�OI�����Y-d�S�={&k򶾌��禩�}c낪��3�Y+��k	e�����תа��d�K�%�0t�X`)ϕ�H�k�c�f�������bN�H;L�ɻc�DЍ�ª= 5^�	��f3:8Qq�Gړ��^ߧ�U��@cFj�ط�	�C�?R����5�`\�1Ǵ0Ie�X� ��[t������X`�.�[�]�fTۦ�B��C�W'߭)���⚚�YȰ�ǁA:��њ6����R��;���p�;#5��|���"�x�(	��p�ֿ���d����@����Z�8(ם�ي�5�12QHKi����I𕷎��	����&#�b9 ��ܬV,�P�"[6��[��tU4��:�{i��8w56��b��_׆�L�0zXܬ�1@M���mB[�ɘ&��:,~vK���߰�&�������X���b�c�<a��y���7$��U��b"�В���z��Ȧ�^��'�۹&o�L�'fz]'�,,)��h0�K����Ϋj�5(rC��9��9T����;��ƌUtg�ԥ9<�f��v��\�ե{3q�0��s��¾�"N����QI�,v�2���Y����G���jL�p�"���/Vm�1��w��Q���3�24a�����# l%U����JY^.2����ǉR`��)|��\y3|��m"@z8*E����5��#J�^�D~T���b��R%c����oL���9��g�����M �ae	�_��h �����p�]4���-���z��I�S���q�b`ei��
��a�JV��Y~��=\ȼPQ�Ϳ�c�J�� �����F�:����:h���f�M���	�����//6i���Üﻬ�[=��㉈t<��4�p�OOΖ��G�)�u`g˩�I�E�V��w��	3|��H�ҍ�����KiBEO"�|k\5�*[s8qPC���:������O�|���W�r\~�Y���i�?+���p��0N��׾o�Ci>�rj�;��/Ҥh��������܅�{�J�4褎N��ܩ��-s��xH�_1A��rӵ}0W!Y��%<y�%a[�|WsC�����X,y��\�b��_��R���oaf��a��:5`Q�����灝+4�TDD��9+]?C�����gwXt��v���BU9{O����+����z᜔�ҋ��o�Ƣ0���pJ����W��z���	ha4\Ym)N�d�˩b+9mW:����%�� ��M���	-�6ily��O9� ��F-��H�+��}'�%�C��G�Ö�S��`�b��Zh�r��%%����X����\���6���sÚ�>V������z���`j��h~��
N�N��7�Tza�&uYW:��+��I�͐x�(kH�>�L���wG_,��EXD�T��;ܻޗ�nj]8��_,�$6���&�������^�8 ,~��5+"�h�`�^���X�z��YAL���w}�Wě�2~�t�����C>S�=<LC�o@�R�		��[n���x��n/��%{�}V��ՠ�p�lZ�E��{&Ϸ�np*tf����H�4{��G�72��H\��T���Eu�X��-M�V#G�4����C�;�&%���-M�H�B}^� Y�ۥ��E���[Ͷc�Ş�� ����z_3y���0��y9"�H��Cfޫ�!��zz5u�i�W4�w���%[	�xwHA����D��Cq��ڣ��N|.ڏVU����uY��Ȑ鸍F���Ġ|�[=kpP�mrب�%t���&ڙ���1�3��jq���~�4��~�\�jݒow9di �C�i����ۢ���9˚����EA��yg�[�i��!$������5���J����P��(������USd�OI@�:�_��+����������֠��(Ag#��8�-�y:���۟�h�=q�u��l�N��`--��Z�$E��k�i���e��%,�I���@&@�a��f��L8A����� M��_VW΅���|�&k5a�؂&S��vƢ��3\>�D��ۓ ^=;{���`�kd�b�4�w�d�k%y%�(�(����U't�b>�����?��̎���|�r(r6eT���2�U�L_&���@R��<@*�ԥ(��;Kxi8�외�����5o�rNF?^l�E��`7i�ф�w����v)Rx�D��s�Α�����g1
+g!O�4��E�RtX�gҪ~�h���5�fv _�1�T��
[omOj�����nP�o�%��ѐ]ł�1B�����NX�@e�ጿ��0����r�H�xx>�}0��I��Z�b�H����#$�'�m���`��[���cQ�#��j��_]��`h�d�P�v�����Hק؛�� T�	�b�����C����=�d t��E�^��.7��
ܨ2V��Hn���^ X��۞G,8W���l�7���j�z����Ƞ�XU��P���rǿbc�n�<�g+m�l�L+cTģ{�-[��f�ue����.#��m�ͨ$aWI�����K���}U`�<"��ךB��өJ�aB�^D�c=+��?�4��p�IKf1:?����J͟F����u�2��g��V�	���J
F���E}��9U��b�FQ��nc=)P"��%�t5�`�,Y�{�.aĞ���`-�c� ����Ј�a���1$��F�+>jIR��cS����a�=.�CO>�s�q���DWF{�����;��W�l� �[������ DΉ����e�tH��3�f�m�R�aF�&��Z���X��pֆw2�w��ڂ(֌v�Ԋ�� $Y&�NԕbˌW�4�*�y�5z�ʠ�y������@�o�I�.&�yj�����@�B�C<��=���[���i���g�T�~���Xd�u��-WK��xˠ�����*�3�E�yB�M���}*�(�w�`ʢ �'i��Ф�P�S��> ��QûD��D�Hu�H����6�5.�-�<*�W&(�N	��D7��!ogߜa�$�ub�9�q����h��E�3�s�@-m� B'�z��i�Z-UX�#� ��"���X�ǝ�rR� Z2��4X`־���;����8���ŋp[�J�X�!��+�6�2b?�Rz����<��u1'�M7�x�%gx�eC>��X��$��_��DCU|h���7XE�r{-���7k���Dr8�T4��eM�	hhd0�}b���l�Īhǆby�<_��cʋyɤ��dpP�*���ՀS�����d�S�q�ڦ=��[C��¨����u�ݎ=�9ё��{
x���N���~v�Lt{e�`��Q��~>o�s��ҸT,��ο�Q�� ��%�~��o�����٪X#�ο�B�|6�����&�XA���w%� .�TmY�Y����> H?M��	�ڸ��VA�Xd�v3ɶ�k:�V�S�Ζ��	�~;���֍��S����ev���ۣȾs����8�k+Մ����}�}Q���O0�M+�gj������j�h�%ʇ�,����tOJ��S�=�%�Ӳbkl�ٰP7:�݇��X�\�m����s�*V��<}v%�c�3�K�0l�q-+_�Z�W[��Ε*qY$\�)���F��ks�Ɔ\A�S��3�+t1y��O�ǧ)Eĺ��pAj\a�6�vf�Ϫ�D�~����k=���b�<��2׵j�d����p��n�U��ΤBy�`��!ՙXC�Nf4�^P1�ȥ�/��Y$i.Pe(K�u�#w���p���+��f� �!�zub<L�S������y��C�_N�c�*�[�G߯�)�O�b��>�0�!>G�0�3z���
g<�,�{����g�5uã�������E�������8��� �b���c�ӡH�u�����8�X�[,M�0�Oe���3��aa�g�}��ˠ��D��ǂ�lۦ`'��=}����#:ݠ���V�V@�ór��\�[\S�JJ(�=�}��5[h�imH����fY&�
:81���Dz�h�509��I�~�����ė�W��\Y�pHܒ%�j����Z��v��?%�p��oԚ�#��α9��B�9����:�~,r�a�RK7�i�b$�l��(ۆA�H�@E-^�>Pk�t�b���Y������Q��5S��� n��>#;�/�]x��g3l=���|���-�+��)+Z|�W�e��_X�$��trwʁ��=�^�=�"TX=[���6u��!��#^�s�(~��B�䵗��*��5����Y�����m,���b��=��؅��11��DL�[Ya�����iy\�0S�5�@��7�B��"��d��������c��Hx��o� �:vD� �� �P�ۧ�A��Ç�%q��ə�k�
jf(͹�{� ��1�E,��m�$�N�K4�_�����`��з�9��}�V�F���HfO��[t�ặZ�8�?����hs0WL��Y*g9F�-i	OhwϚ��v��=f��gOt���	D4��E:��$��߄�\E�	sa��e*��'�X w';����`i�g��y$$F=��{ig߅g�M��l��0!Kh�]>mMv��Býd͛z��f1
zw�j5�7r��}��W�p�]�Cú R�E�������v�\y�O�/��T����	&"k&"z�o	7��
ۯ<�)3�\"#&*ў�`���VM7mgH7���eهL��8]^��-����[�QY���S�
�츣��޳V-�	�����b�3\Fӵd�4���R��?�T����&�B6��9P�jSIPW�F��m*�E�S2�e������E{����{���G�e&p���
��S�;�R�|�,��^�zӹq��޲X`Ŏ��R�+�Rd�@�j�T��/Ǘx:Z�M�L�}��J�>�z �:�K8�{&_�����1��cᐋ2d+�nq� ���n�Mu�q���
x"����#h��[8�j�$�0n����%��\��C߁7$���!�csٟ1f.�:9#ǜ��l
*�J�A�����Mp��D�݃S[.k{��c�b-��D�,�9JvNHP6҄�9*�pΟp�HU��2t�Yka눐1G-�[������Ob{��$K�Ƙ�g������6LDf�p"�\_MX��PŠ_)p���sI�wz2"P�Ӳ����-���3�[��6��/�F���.�	�`We�d՞�BݑԼ����ʝ�W�\T�����F�A��9�k]99�T�A�?7=F�_D����m/�T5����NZ�zB���M&���`�d����y*qGM��_g�6_*��Y4S�%� ����2 �nI��v��u��J�Ѹ׍x�בXB���v邍S�Yze��転�'&5�v��:����W�`5�>ΰ�4�o���#��~'S�;r�{�$QW~b#���oT}�=T�w�|���W�Dh���8K=�� &�;I�Ϸ�//��q��/Ӽ�f0��<B}�݋�J�*��S�l2��`���r���9 X}��������Y��廒��4�J��k���:�8��].�[hM��}�R�8GE����7�?G�.�}� 8!�{��������F�=�璲/\��o��3�y����~!4�A�f�1Q�d5ΊB���I�3�>)f@�Ek���r��Q���b(�	���s�,��=�/���Ncp�Rⷃ�|N+�+K� ��R�}�i�rO;<l/�4�`WHy�:����*9̼�Iu��P+�=��F�3�_C�Ҷ?3m|���^���[;���+,`.ߐc�hޡp��V~���v��[��)�?�'{���r>Cv��й�n'���[���K�� �X��׭|�Il�]�쇴���C��n�Ÿkf�t�=��{��{�'#/��৊��0.ׯs4]$����&��j�rv[1��L�5T�4��^h�t kϫ���(�����Ὃ��hJ*�4�]N��V*����p�ꎜ��:<���`��e���<��k=|'ϊ��/Q'E�v)<ӣ	�8Z&-��X+A���=��w/C�:� z�᱕��!-A��@�|;��s	�{;�,�G�]e,i�^T��dC,qãz[Q�G��+�	G��kvQq����u����~Q*�[,P��Niǆ��p%9t2�b+^�vb�ݏD���rO4i�Xz^�&�{'�=r&sNiQ�G��Dm��J6�^v�́�`���E�J*J�ң��A��Sj723s� D)Bv�(n~�D��T>E�Q,�˾	��P���f