��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQl�E��*����XR���J̕��������q�c)�lM����<��t��X�_u��4s�w�(/:��Ǡ�E�?��=0*���r�:������
�J�\k�ne*"]-X�1�ʸC��6�*����_C����I+8~�MBE����O�V��_�f��UјW��r�R�Y��?E�H��R�u��M��URl�B����*�9��C��y9iӆBԡ�tM���X�D�g�^%qA���Psٜ�D�Kd~��m��E�6.�>���N�0�2�T�!��:"�k:p�J����q�C���1X9��n�В=��ѩ���?)�=�S���^�ie��{G2.0���@{�|�����r��J�nG�i>k�Rֆꬑ��JeGA}���л�ex�mf>O?3���	�3>���mm|_�_�n�C�~p���R�����PB㔛"��H7��̩W�/��za�u����"Da��
6������БJj��r�ռuh�zL��Z��5:�U�ь���ީ�6�?D>��%�-n�o�n�h����z��EDM�O}��[:=�\��7�D:���W^3��i7Ħ��aֹ�fH��f1vr�]�?+�o��bpVǰm �{ӫ8DL06�a��ࡑk���o� �5@��
�֐_��g�
��e��S(�Z�Ú?�t���rM]�Km�H�C8�`v �-��d-��G�6.c:!~8\uY��N>�S�%h�G$�>�Ү���K�u�_=0��[X�k��496P~M�nym�H[4|"�0��,T���w�׸0L�J��/�ݕ�]�e��d7"�d�x����e��5<U�'/�	j��"B"=9�YM��-�;���&H(J�|�U3G���#��
_�ޮ{�R#6�~��X+�<�q�,tV���b��<���:D��$@M߈M:���C ��ٹ{vʅ^��-S���\ay>�M��!1��"ߗw�ºnL���]
NjW����Ҿ!S�3�w<�.$\�l�@՛2�p�U�\@c���D]�kѣf�T ��?���t��Vs=�?M'�ѳ�꺿�M𸥰 ůDG�ʖ����R��a�U�ËG�`�H�&èJO�	�B�d��:���������2}B��H_�����d���H��Ѿ¿��vz�/np��u�	A�uK�SByDbR4]�δ->�:L���{6���P�W��"�M��+�����U�X��߯�(�=DE�Y�뙆rH��E/�����̽?�w��yѠ҆��i�Z1r_b���1N�-��z��Q����9
�zt�w��g'#��ǈ� }�D�W2��^x�:��$q"���$m7�'f�'��I��]w����
��N�]�,�b$~�,�.�nr�E�*mz�,%�����\p�0��o'f����o�bYY&��lx�����/�G��I��ّ����
L�\^�́E�L)=�J����#�\.�|�?@�/ �S�w4��N�S_P�{Y�O���n
gd�#�_k��KV���쇔CK_���"c���%��[}X6I|0�f�0W������VB��#5��?=�������R��2%u�Ò����/ܮ��m*�gDXV,�$Ug��r��Z�� �bQ�L~�FV�P�+�>n��z섎�,3����	j5���Z�wta�d{�v�"ɷ��Φc[u)lQ����,�)�wR��9�4ͧ��y%˔�P*`�Z�]����QQ	R��؀� ���v����� [
�y��ٴx�`H&�m%F�_o�A����2�c~=饙ض��B�"�|�׏2	4�`��}�.^��Kғwy�L��K+�ǖ��_����mC���t�|f�ʆ�eLe;�'W�j�#Otd�8�􍾞N�f�8�>μMd���2h��
�}�<@�����*h�(�Fw��*���f��b(�Z������5#
�k2%�٦�:�Ȱ��fv�e���	֕�[A:��M8f�0�V� [���Mnۓ�N�9�B�'э>-1��3fcy*�q6�5�H�����AFUƉ�P�~��1Kn5�}��|�* �H �rF*�?R#��W�je�t��~� A�:�Ē��.֯�uZ�Y�%�.��8��ˇ��c���e]� W�u�Ц҂�~���ӗ�-�9*6A[�Ͼ��C�!Y��@����#� 1�����{5����&�z��i̼q$��.����m5"]��=�H�8���9�������S$L}�{.���dHם��_���})��L��Q�'v �|"-#.\d��19��t���f����H��A,8ә5�]Lirp��v�O��n���cU�nN�`��w�����Ӑ1>�I>���:H�/.R��k�n��\i4�΃�V���wڏ����]8�N��{��.����/�;�XhuKF�=�Т��K��Cjn2��)e���)��X����jgx��1����8��5]�O�r�J	|�*����߮���/Ʉ��J`��\���5��,��j*�G��H��buw�հC�`�P	I�%���7��}Lm����ù-rf8�o�[��E������K�$�����DH��F�1��kԭم�uj����8��%�������S�����W�V6�n���j/:�>�rg���򵹔���/|؊c�Z�Fpx�x6���H�f��K�ZXD�I>&fqu�8P�"&b�=��~�� u��	 V�U��/ˊ`
{���j�ɡ��o�b'�}s�p:��i�h�;"�\�?���`ީ�l����`lq �@H4�)��%->����5R;��B�a�����5З�P� �Lƞ_ ��ҵ_9��Ā��r[^���FD���3�sx߫��y)2
�G���t]���Ǐ�%U��용N��|���� G
�1�F@��,��t�@`����9Up��1�S��1���4�y4���V����3̂+��L�1�iT߁D�4�N�|�W��n�Fj~V����
m��~f��a�B/]��9���@^^Y����'N4��(�ó@��Y�`V9��rT�pǷ���P�؉���P��bn�v%��Ϲ�O���e��M�{�B��F�����Y��+�{���!����&�����.\�!�:� ޣk* �I}ܑ{���I�zv�#��tOݠ�9�)�@k���R[-W, 릜8�=}/tR��A���9ny�g.�UO��\ݏ���:M�Q�
�竊$����?q%�3�C�ylf�z1Κ(�ٟ(��2/�G
��t���g�k��J�S���.a~�ھS̩��̹}[�y~ �7A����e�y��^���.�������_9�;b���=]@Ж��A�U�c2]��6;>�6�I?;(Y7(�쑦�����d�wnӲ.>¥7�l/?�S�vk��G���_Ѹ�L!��bUOM
����SA�Y�/�N��xpcm]~�{Ͷi%P�����rS��9�ۚUA�`%�)�qzt[ג���m�6�Ƽ���̀W
�8%����U!�ck<��Њ�E8SgD�!k_��?�	Ҏ�R�Xg�y�?8�T��G\���#��?s%�I0���o9�H�޿�o�qW�ԞX���������+Ǽb�����A7�1m6LF�oDZm����v�	��E�>Y;�/1�N�qQ�������Y���٦�P�E,%�T�11bRqq�+wD����}���QD4�5%v��Rdf�̍�mx�����K���x�o���\����=3(�ֹ��Aea���x	/���]T�
p�M{�Ȉ� ����о%�V�Cu���C��5�j��3A�U��f���CΦ�ѻ��i/z塌P��V�T$�;	�1D�㜲�Y/�	���qvMS�$xօ[ۙ��e������cPK��<�$�ꂗ��Q��O0�D|h�)��Ӷ��bI���4.ʥ�BM���*�t�d9�6��4��5���æea`|��ı��Cޱ��?�"o��1�����|����ǡ�qݙa+�	t��	նq��p���:�`��C��k�J`�h�����@��/��T���+%��[�u+k�d�����*~��[�Ì�Y5r6#��MNͫ���sڸ��!��P����G\ ����UN�б�����(�x9�40��D��9������=�X��G�l
���M�c�57��ujCt����ھ�f���i͛w�x��S�w��`z;6��.�P��w	� �Rֵ�.��X��mm���(�����24��b	��"��.���ܬE�\��y������w��1����i���m�i���pN�������mq��x�b(�"�3�W� �?�T��p���Bf��������zX��8l�U=�e��gu�8����4��Jȧ�F�W�Z�n���Dd�>�W&�} �G�Lq)�R����q$���fQ5**WV�"�Jar\�]�@'�V�.R�:��&(ƹn�[�H����m�?w��6�{2c�h����qY�)�T��M��k1�k�������nޟ�;���*��vO�5�a�6S�1M$�Fym�.���U��E�����d�3Ey|0�t&W���e�Y�s@���$�U+��5M���`Ӂ�"-*m�5IFȺD��F�M�'��&
M�=^�-5�<�]׭ݛy]�`ѻ�҅!�\����1���x�M��@��D��7:�J�����������܄�m�+AkeO@:�.�y�D�����4m@=+DEP�톕	�m���FQ������J.����k6d�1;�L��jJ�V%��E����{v��@#V�ʞY(��a�>�����4�1�+�"_(�o �]����g�C4Yf֫�Q�)o|PQԍ�b�QtҙVDk����j�G��d��-��9�r��(��m�`O�#6p�]���w䋈��@!�	�74�G#>:� N��<���@�v9�h����N�O�^3��;ط>C��|�'}}�7 <�3�3� ������hd,���~-��vej�&��|E�.���f��^)�Bn��v`yK z�H��pBok����,Nv�XX�NSn߾fU|��w"��n&�G�h�#k���T+L��u�<����Geq��y���s~��VTY��%�3���VY���c죍j|0FXk��)U�*W/���5�Ky�6&3G��S�؀��5���������������>C(.2M�;M��8߰�������Q������"����$�I'uQ��_;!�l.����^zM!��b��:��n�Id�R� �hb�6Xty�I�澐��}��[6VV���4��i�1v���(h��9P�f����;�W�Z�=�����<��C0����%���n��$�|V����2��_�{���&�OK�߹�{@a��(ǈ�٠/B=.9s��[cO�W�O;+0v"j8�N�˘KCX6���6���HV�N"Ʋd�$L��P���:M+�0[2��|�B�Z�t7��GCT���]d��<���7����B�rn�#w^�lRŹ��|�LR�/�wA4�|qo��Z�:��kv=�;Ki��q.��C�}��Na&V	ԇꬆ3��IjӚqglk>f ������(��
_]m�`B�����������7����{��>��E�R3�ehr�,w��:��F����K�y���6+WGeϋ���:ˏM���W�!��w�0F�G��x~V�RΗ?�@���+|��y-ʧ��'\��4�7wf�0n���R�u���4�<u �����ח\˩@1��3Ea[ھ ����5d=4VŶqvd i)�Ť[��Z��;o!Fs�� ;ޕ��Q* ��lS���p\@�nlǮS��hs���xN/�|[:?z��Fe��q\���UQ��8aZ�c�֓��P)d��}8�;h�RIô���g����>�Q����I�Sw l[/�A� a�&P2x��eao�Fp�LJ�A���V ��۪�)�^�9^���=��
:Z᧪�"@���&n��-#�R���|5Y���_�s���A\���_4$$X�b�֩[v�m������ �6�A8�݆�$[a�5���wLWӝ��y�5�Ǭ�5�]���	વ����|�vf�:�� T�k8���� X=��ެ���
���r�h�4��	��b�P�i����g :a]�(��Cԍ+����I���@����z��T���<|�K�P�d�拪�}�,�م���Y9��9f�yq]v@(���<ܤ�ۿ���%�e���p-'෰Q�?P�1�^����ɏ���a�1��ƩP��}j�1�4d v���VI--��x��_?'�bX�Yu]�2��E�g���b���f�Ԗڈ�!�3�r�����o�!��*<�����&���]9��Xkg��И9ڡ`\�߱"�z~;`�oR�����J�K�P?�/�p�9&�`ii�C&��V��E�Fo��Z�C�,��ϡn�J