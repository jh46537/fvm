��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<@��݃VQ������k�w�
��T ���6Y92;�R�3�C��7$���]
�	��ݓj��t_M0�+ob�N�VT�Ϩ�m1�8qV ���$ۅ��|>� "컃���=}���$�]Q�t
H�i��D)O��Z�~�6aVg�?�<�0i"Tƃho��$�3���0:�U�,SG�v}�R���/JF��>���uV~�}���b�D�P�E�s7�?�[��Fod�����4�LLȱ�N�f,h�M92�3�Ҟ�61X���$�q�Gr��R��A�3�~hP�;�+�-�=�z���B�3�$��1�s#���4�6��t��j >w*䌯�ean��`H�[*�#�x�T������96BӦ����x@z�k�ۇ-ֳ�A吠y�?u0��)TЋIY��~�$��S�C3Ή�χ���VHgB�0W���ݪ��'�t��jk�_��r� �/
����P�b����c�!� F�,�hx�S7�����:]�
�_]ٞ�"��Dd�r`$��VvU�j1���N��<Q�KuЛi4в$���V�tjh&
	����ݡ異�����P������t=�ա�>32q""yP���c��$����M�l�2��MLO��<���v�� 6�߁�*�v�tq⿺rh�
�ߦt��Q��R[g��;<�v�"�(<��_�۹�v��&)�k.�A�ʪ��	�T�l��a���J�<Zm��;X���Չ��! KJ_o�0)����eA�:YR��5�^:g�=�Ҵf����?����c�w�}��ހ�D�,ѡ1�}�A�f��q����}�<cB�ݥC��ob�I���X���a/��_4��Δ��g
�10�cY�Q�h�����	%�
��T@%�,~qR���-�Mm���\e�<b5-ۿ�tLF)�g�-��}�0$PAl
ޒ �Cx����]d.?�$�������� �����
��������V<��pPM"sv`�M��?t	�}S���� ��I�I æ�#^����׭|ȳ�l��s��(����ũ#_�g=Q��3���F
|(�O6w��Cf���x�v�j9�l� ��v���[x�z��C����-�����,�����{�jm�s��'7�!H�҃���>�p��c�
wz���,����c}V]�3��r��;�;��v�)�뗌��U����K�N�QmW-�跻F�T���iU#��j��y�+^���&]�C�T�roy�B�Hâ[���³�%�?7������T�'62%Y!f׬����r� ��\z�����ǆ�I'��3��g�gs���t3I�M����F7��#Į�Ԅ�&lܡ*���}��^�}��c90�\�� fi��`���C�5G��6q��|�9�pֹ��p���S�Nf�a_�~�L����:���; !D^Nڏ�����t�U"�j���R�Dat����GS�� H�Y�#h�N0�ւH���=(�� /ߍ:���������~�$d�dt��ڷ|�2�.9w�
�Ȳζ����YF��#/��7YH��Ɩ�<ã;���k�H�ٛbkʟT(��獊�9�ԆSe %m�I�~ZZ�� 1�{�L� 3�5�^��! ��uh#��3�r�@}��z��Q�U� �ʇ�8w'��I����oF�Rb�Ϻ55ƚ^������nD��W�C��Z�{�hH�@�qR22��{)�|����{uB� �]_��b�'"�yDn�߽��Y['�r1؝hk@껾H0�J86I��S��o4���r{72���}�!� SO�JO��Z(�Yva<���TpXM�h� \�)��|#B�����bm�e��/c�>eC~�p8QQ�m?&�<���W�\���Sg+�����I�4�J�uK�Q_��l" �R�C��@V<;�F��6.d�v��W�^��*���nϕ?b�-�<cq=�	�E�����iֹ%��T�m6�Ⱥ�'RPw��d��WҸ���N ����Q"-����K�������E,1iy���_MG#��2.P-ǈ�6̺�����3�4-���=�i)qZ�����Ep�'��]�Dz���y)����2�G�.�n�yxB'B�U�70�����%7y�>vo��DS��1��#�1VLm��P<�SZ��z��r��`W��H�l��ݾzN��!xi�
���*��-Eލ��?i�!u9����S>������`q�(e��F��S��c�Z#���[���C�����:N���R�\_/��N&𸮜�(m~��qq���/=f�Eس�����ӎky)<Hw^c�T��'|Ơk�-[����sht\�Ժ 2��+�T谑JZ{$	�p���?���T'��t�A0zMa�Π�`��q��J��z�@.�4bJ������Z�����%(�ջ+VHz���lmL����vΗ���QC�&�5&�s*p����c[h#e-Q�37�C���V�dߏ������{���9�܌��31�(�>VI,��#�����=(�:�_2��J]/fDAgœ0�a��C��'Y'��o��z��>��\�h��v(]���p��]TR�,�PV0O���]~���'2|@@�&EID��u���VkȎ%�d=�T��d�cph�P(rU����Fʂ9�y]|0�s�)�y%	H|�$�|s3���C�"������+���G���Q�&��7d%�����2۲.���-vA�6�������]�D��X�r����� 3[\w��h�Qs����p� ��