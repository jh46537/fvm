��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�w�\պ}���'d��qx�Ba=��1�@t�lo�ܦY`f9��GU��O����5y�k�wy5� e%�iHF�K~3��Z�������# ��d|��̪�����PAZ:�;� ��Փ�?�}�F��3LY����U!a�N9+
�\�:�-��*����d��W�L�vb��+�Ԋ��r�����WtUItq���E#�N]h����޳�ᓗ�C�����9��~Ć�%���cuu�6������& �Z�
�)6L@@E���s�|[Z9ԍ�1I�!��q��|�\�-���?:�+]��h�;[����b?0�+M�1v�:Ԙh4���^�6�W.�^�(r%e�޶$~M:��S����bs�YJe��5A��k��~-];����^Q�
0�~�ɨ���3�)�|��X�kXk2�����WB�z�)ɢ����1?I�=2����=�baU�t��&�V�{�
�n�n0<M�a�%b�^�2gd{���\��y���@ǨX�F\�:��a.��%�d!��������/Rn��
���.{eı��̴��J���� ��C����D7,[�gn_�K)IF^ڽ�|c�aQ�P��6�:I��jޡ=��Rs #4=EU�N��;��^��ϖÜ�AM)x.�U�G���"dB��7�^ўR�m�Ղ�Xݿ~���9x��"���I�Pz��89+	�{���'P��'�#�Zh�j�`���	bE�[�=Q|�q�s��b⅛ӝ?�{j������i_��H�!f�=��s��VXM�����tv�O���z��?�aIH��.`�x��uVS�g�ԥ���F��A�>Z�6�$��#��7��_{��B�tQ7����?|�������2�fj���D�5]���^;3;zuP ��hZ��#$\d�_�P�R�QԻ��|}�zgw2<��XnV���i���P9�B�$<�`�b[7"��Y��9��!�z��&2.��jM�xV��܏�t�l볗�e-q��*�hx[�FQEc"(xr�.K-�|��'X���D|���q1�g����2k�JK���=�i	�I$=�Zd-�,��i��ұɗX?}�����f7���h|�9�ه������t)��Մ��a�	w��ٜ�Yے2�Z�>T�	��5�_�U��1��B�9���F�Ak�l�ԉ���DL�n���fv��rw���M1����|������i�?��w���� 6�߯E�p�m}x��mT�gv���Y�ܭ,�+�H/)f��%�=d��#S/&.t�.a5<MMz����oc�"��8���fO��6�+�b��?�ҒE����|:-�]K:������V�^[PHe�'�}�:��w�'E9�|�T6�2.�����퓅��@��F�������چ�h,��>D'{���=ȱMz9 �l�ޝ2�|@Ҟ�t9@��&�>�~�9�1}큩�'�Ў�,�� H�z�/'9�U�\9�*W�z��`P��5��u�[`��.�RV��H��B�h)�fГ � ��9�����vl��R�9�ZTN#�$/���}�s�����!�@��_F��ǝ�!$�=BGy�6� ������Y���.0����E��m6�����,#	�z�?��$O�⽇c|gR_��r�v��/bUJ�5	8���WI����:\�+��1P� ')j��/�}��t�HD�K�V��	Ө��~���/-*;Dj��{�yLp	�nMI<Ц������I��_b{��
׫���#z||o�"m? �6�x�NPTÒfd�u�=dz�V�)��,cR�e�����?��~ ,N��`���ր(p��������Hc%���r,,c4?fp/tQ��S���i�mh�~-iZ�P4��1��NTg��Sb���[��.71��,=�@I�"���=鐽�0��9�W\�K������n2�� h�E�\o	<6j|=�7�M�)Q�t�����V��fX$|>_�;�7:�;4�Mڴ���2�Aa0�fb��ލB�������/& 6��u`
Y�h�ɸ�b�:��Sq�Nt�z!�Qȏ�����)��C���|�p_V��5'��G��w���'�ّ���%MX(<�ƽ1h-�=�\�=eXȠw�Iq��l=p���˼�bGg��%yLy�򚞣H���]%�;t<1��@^dD��2�p��5�w�-W�k�\?n]{������ ΉX���Ж�Dbժh#�������M�����\����
��T��/T{�G�'��*���iD������1c�OL1Zl��<Z�$�1&c �{b��b��}¥_lQ�G�1���\%�5��i��DR9?�g80���i(�������C(�΄���K����>��
 o<�����UM"�1L_P3.X�F�d�5W����'�C2p��xG|(��^�	��I��A�Rk�{Qq��k�g�S�F+"���hRh.�:$��у���ÿ8a��G
J�ԺP�~�j�<�0�b#��`�n���ҙ�WW��":J��s��+%�P\P�#9�Za�������KV1��ݰ�Bæhy*c����]�ų,Oyr5�r��� 0�Z�?�]yI��7������-�j�\����t�MB�klֿ��f�xT�
 ��g��F�O��	螲��"{�xeA:��ڪ��C�nۣ`���`��N�=��T��i�#S۹�`9�%�=ra;���E�@㓰�il�i|���aR3��c{�>����G~�撍[˨�\���s4*�=�>LƏ	���������!#�nZ]E����Dmڴ��2���F���NTbu��� ��S
ٿAQ_�krB�>��P��e0����&���I�1}�Xoݾ�(���2
��Zacɰ��G0����X��r:'�/$o6.����'�s`ͭt�ao��O���cw,R�Lg�_Wr�!���b�
��"5���4}�O��PEՅBY��~:�
�轺[���j&l�h8a��Y��˲O-@�Y���B��m� 2
�:����:�8�l��!B�6̻mIv�G�PU�.��!���n󍈍��%C�ߍ�/7,���<������B��������ϭ�.�nFf1!@�B��yo��a���v^ؐ�Y��KИ��,��
�RB��Y��Gi�<U�P��cq
hZpm�B{��&�/À�y��;1�f� �����U������;��*Fu(l�F��ft���e��à�쭱ݲ�a8.�"�����zA��$;4n�0��*/T��ih�N-�xSd��Du����3�:���0�N�A������(0���u�ԑ�k���p`2�[r����SB*&�����u��2����ߧ�N*�����G�9Wګ,��q�0~~�~��cf�T��J�vxx��S�Q67,{1���C�_��b(Hz��/�f�p,��g��<����B�S��8��Q:�1�v��,q2��W���4ö�KmI4�=&74e3�'��V�En,���	N�6�=b�m�[By����6���{�4z6��������}�����E�������Ө�<�X��|����3=�~Z�y���WGY֙�����l|�r"K�l״���(Yd��%�Y�?@8d*8�B��4D��bW�|���ط{���9�G<[yS[ʤL���[_�[��@�9v�9LihO�	x0��-��Y;1`���{?��MO���+��E�K	u������]��TT�,�DL�*5�|�Q�9���/�^��ci��@iI�j���X�/`ĸ|ء��s�G�*I��v9���
�a�y��냳"6PTR�p�vyn����>��(X��[i����j�ˋvf
%x�C�ls��0{���Ⅺ./�u��ydϫ��ޟ���4�������W��+�A��O��*;E
r�z�7ȥӌ�(Y�v�s4�v����@U|���\���=��4q��WO��7��"���`��jYk��P"�G$c�h�l�\�7�ͳ�T��� n�J��$}|�!�T+� c:'\h1�?4ҙР��ɥoX���Y,�E��i����)����2���D0!����'������n�=��j�8�Q@��=G�k3�����I���4}7� G�:Z�E��iW���Y��n���}T���_�pQ��ͮzv��ߪ���?�ٳ�Z���N���P��tF'F�x�� H �?h���w�>RӋ�$I����6b��'��5�=L�P�#��-)��&�P�c8ƃl��p�/<�G��:���񡎫��P�*�H]����˼�*�4� ��RMo�W@�Q*_�K�9�	�ܲ��/F�`GF᤿���I2�e2b�5ƃރ�^�P����W?����4���2�;�^9:���|��Bj-��Ր�͛2���*�n$�F���<Ch���pQm����`��(!��q����ғ��ٙ@��N���(lo�,�3�Ӯwc�XEƑm��Tn<����L���?r@�sϸ�o7��6��`�3��w@p�Q*���/CTb����\`Ni�)��`-]����Hdwfο�����q��mu����,���Br�߳ƚ��mldg\�����*G���<�r%W`�#-�m�8(<�|BH�x�,%.Nv�O���E;�ӈ��/��ز�J�!����7�
������>��bֵ��͍6���2ږ�|����I$��Aj��ҹ(qt61a@>��s��nzI0������_Dۏ-6���!�9��&���qW��t��k���jS��tȿ���C96Aa�ݏ�Mա?�P�8\����$d�7J#�\���T�/��%�S8���ٯ@�ɽ%}��P�Fry��-j��pj��k�n�����b0r�h�G��D�-��:�տ�@A� EЩ㢧q�	�L^!��P+��ˁ�>��&�n����e@����ge�7P�|�Eݼp#rj�O���Ӣv�' \V�C�����zt{u0<3>�܁Ǟ� ���~��a�F�,JPy�O��Nswe� #�7J��m�/ �^�D��^�8�� ��y�KY�}ڠ���z����\"�k�R�(g�l���{���>��3"HF*�R3�Z"6)R�������oxy-#�GG�٨���zQ�A�`��"����F���[1t��=�>/&��I�����6�w�$�q��*�{@�*|�����3C�>@����Ѯk�h�NOx=��l�c���[]�Q,W��N�N�9�+��O���7f�^2�0���zڬ�^?X$оfwˢ���?��Z� cq�q��������0���j�qpp��3�yΡ����@a�����aܭ�ғ��^�V�*cr]��wz��^�a���L�B:�s����g%1�mr��1���4�&0Fq�