��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�"]P����'�*������@���m�-�2R}��k���+J�����^�X��=��H�����%��J3�������IΠ��-JF�n�:�ݵ��q7�Y�u�e�d��愋����;q������'�����g���8��B{����$X�}p�&s��^Y��y�7ܼ�z����ީ��3f/�śW4��k�����TO�i"�B{{� l���4wJ*�+��5O���&fWQ�"P�e�ꥠ�ik�$�mS[ͿO��d��0$/־�셦G=:�� nb�8��e�"�Ŋ-�����#��qR>#%R�� �nG|�Y=�mz���,t�R�F��*�n.�6�-�s8��>6>o읝S�d7�F-05�����3��?)\���ǜ�ߞ��/��RS��W0���@lB9~|'(;X~�� �$����,RD0���'܌w5m�HWe���ñ5�lC��!Q����$鯸Cf����B�%���*���Z�q�S#��.:v���Ijp�:�:ae�S��D'���x0F+7}i��ʓ��-�Ŧ���G�-w]q�)5R�'ɑ���x,����~~Yf�n��0]�������!/�?��qa���/�M�gR�U��ˁjeSՋkڲ���.ZE�a@��]]d�?/>n|9�!#����._���$����Y[�~ۈ�reM�s����I�^�y%���[J�����3wܛn5�Nd�FFܔ��޺r�]�+��F�3^xV(���&�Cbd�\4�'"���v|08(�W�r��N��u`�����A���V���EJ����E�E�7�;�Z��ɂ�GS�kd����*d�i;��5rƣqg3������Զ�*�S�������I=B������}<��q�t�vɵ�3Ͼ=VF�)q��l��L����2��7�)Z��I�J�_&p��.��4�m�\����T�nF=s�VP/gx;�U����C�Aq�i��B+^b��H��?2y���H4*�sM-�n�%�O��i#.�M���+\M�����&��s���3���1���qo@Z$aN�T��E��{@�*/��b���*"�$h�3&����#���!�
f�[8ohrl4;t̏*tʻ�߂��"�N9��>�('|!dy��-�Ν����&��z���P0����JIK,�j�8�j����G���W�/*.�� ϒsi��ZBQ�-�{V=n�5�������&MV����P����f7����M�^{�4�Z�Q,
Błc��el���]c=��Ꙛ�#>j�Ń��t4�\Y n��=��p�'�XF�X~�r����<�����a����
�K��,{Ⳳ�.\\��H��]��~-�x�>V�SC�K���D���;�(�����(�w1~�ϙ]�����G�ï�A�:m�"��p����;"�-���l�/�Ӂ5}���zf8��<ChLBr��w.~J��.h[�V����E�=ɫ'=��ٵ�8�%f��Q����!��E�����#!�L���RāH���-^\�w�	fw�Sn/P� ����a����J�_PgT���7sr2	ӳ���)�G4�%P��@��'����K�]w�V{�h�����J�j�fm���Dqq�7�`��*[�<��V��s<�~ʺ�wq�T6��]*�~{8KVLN0b��zq�G�@���Ny�q�|P�@�L��|��&�豟��I�kb��e��*�ðJ�l�V�+���[��[x�(X�0�g����$uu�%��=WXރf�Ӡ���.�)q7�īG\�����z#LX�n��X�{ i�܇��b�M���t��K�ڭ����b4��Ѡ�[ ���Sq/�������1�,����A�b�]X�CE�(���ѽ�3ַ�0�@[�ѧ4���<^�R24�ܔ��������Q��U�[�@�
����7�y��p��ŀ�˖W&��e<����S7�Lh����pv[�=����7$���1�M�RV�>���Shv:Yݧ���O��GG�%��Å��w�Ds.���I��'�Lu/U|���nL.^c�`-�g?�:�<W�6�إ��/�,�PhYz��q`"�r��u��i�'c��fb)�����w�"�