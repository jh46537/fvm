��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@���C�X��?�d{w]��T�-����0D+� j{�ą��^~gOs�P�s9��L9�<���٣C{�ag�ʖ��LQ��aB�x0�U	��@\|Y���%����0�w�ȓ����!�]R�m�Xu�1s��9@�0ąkk�<|�G�CN�JkL-!�#G�gLƇ��v^���D��I������p���Ԇ�)x��@��q����d��Y8�$]��L��c�.����d�*~\ҷ_�WK��&uI#�I��!\6���U�E�A�n�4�~� ��/^Q��	�v�<7.\8;��)�uQ�Q�,Qֶ3*��t���f�V��T�BT�8��Dh抢��f�>�ث�Z�|ږgq����/�� �+p@�����*�����Q]�G�^�K�����^����@@Yd���V�����c<�k�SB)���fY�y�}�����c�HE�Z�iڈCPr٭�(��m*yuz�Dc���[M�F�=n
�>�{9�fV5�:�{�l?�����1��ԔZ�S9ON:��d�@NR���O,�i��b�B��X3���m�hS�/m�ޱ:;�8B*�C��pű������C�+��M�()%2����ީ���M�%jR<}B��d��0�_���y&��h�mSs�sg��ԛ�?���V}�<+�ؑ�]�/�i��2:��1	k��a���b"�r@Y�2�,q���z)�v~)��@��)��Ql+�6.E3g��vgJ;/,���S��R0�*E��̀W�M�x�3�x�]
�"�(��$�@v�Q ��9�s�֋+E=�##��ٷZz���x�ͳπ���n�~,1�ʰ{$]�Y�#>GneR-#��_���)���B� �a&���}����F/�&�m]*_faΦ���S�1"'az#R�;()���Vt4�H՟-���%xS*� 	h����k�e���O-�:�T��Cw�~,�!��c�R�s|��û�mm���utG��:�֪lN9��E�buO�n\Y"�6�=y��2/A�ڌP�:�
��>��-�I��D/��`C�lZ�l�;���{ҧm��E�E6wk�����%�evO��A��cu<�fv�F(�\�%4��pם��U��3x��-~ �v�����2e��4����u$��K�M���#ӛ|2��a?o������3߱�>���}7+��T���b�R�I��	4��2�$H���?|��N�oF�I�H�f���w"p��#II�en�T�Ʒzs��?��J�����9���p�\�%2c�N�pm ,%ɬX�^�E���2{7�6���<�|?�U��۝lHT����[`<��ي��?뉪��D���)B������)�:��qIq*&!�����][�R�ǸR,�ŢdjBq`EG�6Ύm�s��@�B�;A!_�����o�2A����l������!2�>������5�[�C��V�:&�E�4������{������@lD����M����% ��z?�䠧X�ZG3��q����5��;��s1�V�/�|����D*�E������J~QD3,-�).[6{ۓ`<Szz+��z8�d�n*u����8%Ct�r�#�0i�M��(:�M�Y�ċ�B��'�����|n���u\����q���;�O�Dg���!�t[+�Y��(������d���'+$%��6�{��v�H�o��.����K:�Ֆq��|y�{�&_a�q.?�r�?n�9�c��T�D�T҈T��^-7	�J��+#�760��x���e�|��m8^�h���Y#_��m�s�%���N�ZtN��]�d6��v�;`�*Y���-�PSxʒ��	�����U��Y���YB�*����� ��v���#�tZ��;������z���y8���+]RIu?ۋ�󯸺k�Α;αޖ�v����J�h�&�R7���M)%(�sr�<�z+)l���_c�M����v�E��ď�A�>k�����D��2ZZ�D�G��kV�uM,MY,�0�����G�o���=�sP��:���x�2 -z��6z����1<�v��>� �R�(��4��X�t����Μ.j�Tj��ң~*��v����es�Z�v�1���U��]��m�
���9��h�w�3�_��� 	�a�/9ކI����%ՠ��tK�]D����L��SE�T2�աY��r��q�x�bN���]������6}�)�6�QH���Տ��6��ٺ���G���N���G.H�,�^�D	���כT�)��w�L�0�t&.*;49*k��jO��]����_�cϗl����{����dC����2`���5W,��<��_h��ݼ��:�ʷ��f ���Y�%�+�YEl-���0��)h_�>����f��
N.mr���yz~:r����~m{L��A<��ΰ���h�`��|�d�)y9]������#�5z®l���j��y�AmS�j���YB{���>�bzr�՜%�=0&�Qq��w�L���=�)�d储�ĳi(1J*2��Ī�����'nj��X�^8��n?K�Q�0[_��Z���G�r����ݛi���&��q	�QSG��}_����T��}�����@!f�"��sq��ሑ��{��m@6���#b��65��ܤG�s�@��*>o���SL��񒢽��9E�j��b�9�?@<�~fiwE��xB���[V