��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9������t�qp/�{?t�kF�VN'���'�.>T\}��hk�K�,/�_�Vf0��t����-�6�M��;wUW\Y��'�j��r4�]�i��ϧ��������t��dul�'����O��A���SHc�>�!}�����~�J�,���̥�y�����.Q�J����
�|5���J�3h`��4F�̓�V�kLՕ�����E�1z���a���?�K範���_�;�+��+�u<�����7�[<����h�S��	�F��w��O��5L7�b�}Z�yD-nsK�yϚ��}�?W�C�%
��2IkK�x>�G��(3�+c�3	 ����b&L�ڤ5�1m���A+�Qr�Y��v����t� ��];����$�! 8�j�0E�獟��� d\u{\��.��������o;�##ay��i�z�Mo,���������6{����t��/vT2�l�+A��c�lz� ПRT�Ty��p0���j�A	�5e�;Q奐�L�6��ίF�s:�7�k��F���x9%:�RKП�"�!W�%m޶�������||����Hp�A�?FS��7�S�4z
�)iC`K��x?�����W1�6e�YQ���۳�/;�O�r�lj���#�#��SB��vT�9� ��m����\p���g���w`^��)(W��w�ykde'�q�Ć��|�ow��Ы�b���D�̾���L'D>�)A��,
�J� ���ލRa�`��sq��u���[�~$�����Řy�D��?�$�"dT �P��)ձZgZ糑��B	�ܨ�0�&B�x�3�sHT��t�S�<��8���IO\3ۯ�Z��҇> �：ń�8����ɭ����XT�G �:�}��@�L�k��&J��e��x���==�Tl�Y�OՀo�l��v.e�U�:d�9$?3$Q�ۖ�:�+������-���he���E���6&������$<�ݯP�1�K�Q���g@E)c��;�ft:`-�I�͌�j5R��ɛ���b?_��z�E13�� .(�զ�����k�aCl�f-7N�t줰߰�r��&�����pXV��8�2��S?�ȥ:k�r`��'q܂�+k�0��Ԑ]����Ts������-��π}CD��?���J��(;r!����O�ӭ�C+f��_�V1���@� $��g@ճ||��F��}�I�B�FVG�:�`�TP�վ(��E�-�S6�U���.&��I������oF�����$��0O�缿�i���v�z9'�t�/�}�����kp��#s��q�A;^���6	gu��Ό��ؽ������^��#h��,�!M�y�� �	� GDYf7kj�]��K�,��o�zb.���F�Y�ύ[d�i���Գ��ҸB�����v��G���!{�EQ�����?����kfOkV���Ӟ�q�'����������F$��:E�E�O_�\z$"Ǚ�M;_Iת)@HұB�K�II�ײǎK������g��z�Q��*��H���+�
fZM`����1�Y��~�v�ѹg�u{�s)�gUu⋑�q�<�
<2��NP��_��5x*@t<��k�vD� Bw���E�k�U;��e*��<�t;�놽iG�
��o�]��������(�ݼT7��Z&y�ӆ���x&n +��F]���`|K�o�˝�ֹ�_��|,��Ug
+p�"�;�|������.i:�t�˓���C�x9�A�7����$����|��<
�F�%�+:m��/X�T���������d���ʥ$!�̎���Wc�����L�kL\�.CĵB�i�ѕ~�6wqi�"�̊��@w��7�:��}d��S�!�u�t���Gm_�jFߖ�!�,�e�8�4�87;�!�|�(5޶�¤<��zs>߷V� =�|I�Ѭ�v���n��&�M�M���-Ј��9u�_KQ9�F�I�z7~�YiNmQ�E�-����������SaI���.a\�s���(K��4 Q���%�����dc���*~�_EBtԞ���h�=M�g�Y�}2�Ц-><W�<A�������a�L} $ePo%�i	����_Ϗ##����(�L���]���V�յEw��u��/�