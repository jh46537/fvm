��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7]�s��^TC#�yM�g,�%kڅHе6��&E��1;JB*_X�o�	�{k��o�%����1��=��͠��k��(�r�F����=� �>BG�U����y�l�	���|�띐	�C��>�헐�^�6$?� ��&�-�)����:'"sVa��1e��dLw��&Q�2<�,���#�n�y4��A�S���Z_���C�8獦P����GW"͛���~�������b�Q8֯�yD��bL�4�j#�%L�wΐ��ot��������{��iM���X2R�;T�H*�j�$FX�v�MX9��˂صtP4O�иGkzgģ>���}-�����}��sh�|�S���%�y��8�� �-2/�G�q⼅��:�����)�C��E)9��g?Rc�:T�o�u�qd�m�}�«ks1@ιT��&k��8�E)A��"�ճ�'���}���!ZѬ�90.Z%7\�62�8�e5��a��{��v���z7�����6Sr�� ��`!��G����(��d�.jI�(�q��]w���ѻ �7�G�O��%��塶���Y�j�rĠq zkE�:��q�����]���<�Q�?�U��
����j�籹�C����E���� ��I�]͆�|qƐ��-�Ky���~�>B|T��Y�A�|6E��T�e���xM�i�Q�O҇\���  E+�vE 5��E�1�`��ӽ�v�)���)���n�F9�)���JF4ⶨ8>��ė?���f�`�\`%��Q�#<�E����|�\��>��3��k%T��j�y}��Ä��m�"�u���֔��T�ki�2�0����)p@��-����ĘP�5����"
����0�ϲŐE�F3��,��it�^l�I!�Ƕ�J������z��4���ec`�2�aҕ0h � ���YD(�v!q	��)��/Q\tl
��E����.#��*?N9t��X�@��k��a�ݑ������ L��d�7��#�R�2�t������P'OذS��~�sHO��Lcb��9�{`X�zk\;sm���i ��/�c;e/V���g~R�i�P�pOȻ�8���G�d��h�3��q����dX��y�56���)k:})��iE.�K�n�6L?����iu�)����D-��y౻��D<�r�8�J��R�M�)�;)���zݻ�/Ak�W�S��_(��u�RG5	 4��b�]�]Z�kB��^|g��wIz���o����5T����+�㤹�W�����;QDT�K��\w����x��Id�iz�=��t�]@����e$XJ��=��"!��{S���d�w��]y������t�4�NEZ��4�>X�|�V- I<��	�0[s �v{�Ͽ)e �qz=���+���n.��ɏtS��Ny��2Ah�����.J�J敚�F�MN;�>|�<=�p�՜� ��c��՞��Λ�C�5we� Y~\P�]�4>e[=sO*w0(�F"�h��жz8��LV|R8���w����ba$�atV3@�t�Daތ
�#q���Xl#l�Z:���w�����Bv	�y�V�5>��U��F�y�O�'݇{�|���I��^�'ى>s�>U�~���{1g1`f�\�8;��U� c%��X�7A.n"3���.3]`*���cs�h�)��.]�Ң��S�B�#8�7R~w.�M���,;TA5�N}�o��ϩE-|o!r%W4�J��ܜ�B���{a�	)���׶�>e:[[��n���r~֎h���,(�#xL��1��m�p.��"��KfWb�����!ndC;|������o�nz�{u| �;��K^>2��`V��*X����T������$��A%;7��2�P�g�ǐ�bT� |�Q�~�QP�g��fxˎ>i-KAYh8.Ty��,��$v/8\Ύ�u4H�`��'�C�����=�v�R�XT��XC,g��<,��?E<��c��H�[F$�Ͳ�<EP�Y�U��H�C��H^A�)�����Tǥ�-���Xe,7*#�ͣn`F�<�m.�����*0�4�)|�~�1(�_�S[�:�J{��{�ύT`!9dC�9#�9_��F�����=�T~��_qp���w�+���k��2r�Sْ���a �%t]U�$�N'��]O;�K�}8I��0j�|;X>v&��#3sf�9 w�����㫯��:�����&}����������ʀ(���Ԙ� �TYɄ�6�_G��,mS�5�p���:l�S�S\]�i9�ɀ1[�J|<�0c��'��(<8�K2�{Aj���l\��o.��%1�)1X,�����}f��0��\M�q�>΢'��.�����o%1���ϧ��Z�̹pYaW�f/��n�M�0)� o7y�����O5�j�>�:x�1�q��
�2rFI/�rg�Q^ԛ'&�	)]Gk�e7G�O�=����A�-�}9G�q����T{�~#�${���n0� nG9&���jZffS7�"�GB7�r�"El�f@гSV�?���,�`X�9^ٔw�L��K�����`�X�v0f�Z9q�Wp��zDN!z�#|�����;�e�N�c*�ځO #F���t�1oH��Wف 7VD�h���#�T�! 쮊M�>�ҫSP����U����g~���g6�j��pJP{J)������D��r�X����oZ�\ �4�X��.�M�m�5�Ɓ���@�l#�5d���S=$�A�>�W�R��sp�P\S��9t��&-z�J����� )݀;Ă�W�M\�c`�Ώ�Kvl�������.y\��ih�>/j� �o��&&N�4i���1��m5u�G�U�PqT�2.rb�v��J)�:Q���=��צ�o�f���RD"y��u8������v�D�P�`Q��r��-y�)h�w�f����(E��J���+�GB�_����=zF�@ܢ�,uN7��~�$��(������i���Q�bq�~���ELX��{<\I#P�	�JJ �3�K��-���v�D�o�g�r�ѭQY�(7j4�zy�� �!��N-}xֱy�As��K����,�v �PQL�%�J b*)�����s��$��7#����@ͺ�\& \|��
T�Y��/�8��(q�uǃd�ţ�eLp�m�5�p�0��jM�^���Ê�x�r�����fh9^�z*�����r!7=�n��g0l��(�}KR���vXv�J�������p9��:nm�g����X%�4�t�Q�.�+�`q�*B��N���G��N�m5ѥ;$�-`���ݹ��)����e)�:Xl;U��L:RV��}6W�����2OAuS�c��jU���� ���
����#���$�l�p�4�Li��3Lex��{���-�O�2;O��T'
��%<�G$M$9G�T��nܬZ96��;U�LC%$NA�O��'�VS�K-�e���n�QR!���r���+����3��Ҥ+|� �aǧ��z6�{�fU�ox??�a
���$�p��Yi�*׳�O>�\�r����>}V1�>ǖI�TIm����Kp�t��+�!��/�t��S�J*�����/��-�����ئ������Rh�� Ћ�G��2%���a��t��+gAL�ms4�c�zu*����EdE���";7_���Fp_[��W�s�� �2�d�}�W�Oi�}�9���9�h��Jn��i�#�!�";!L��#U�6����?�$ݒ�˻
i���W�����F:�9i������-��;ܼ�� ڬCb�0���}Ȃ+.�(e���3e�^�^��cX�7�Ǒ�z7a��>޹8���h�<8U��f���E��z��(4��-�v`���xZc�>U���S��"�k����(�["m�[�)������.�Zt���/�p����Q�	:v��K�ޖN���.O8��TB�]����d�s\�t,Od�O�D�u{f����V@������	4pQ�F�>ӛ�C����Ձ'�U2=���5�6���( S�d����$A�F��a�T5ks�����e�B�it4�f��&�4�w�N|৓;
v
߱�C�Uɮ-�Yw���o��.�c�E�J�31N4~S�t�<��$	��$K�8�(��rc�f��p4,�^S�^���YnB	H{�a����$����;����*x�009<�+�r;����Z��3�^�N���˷��ib���7-x��)E�b_D�ō�Kߕc�%66l���b����Tt��r"� �3���x��1uO�:�f�y1HbFb~8ֈw7a7�Ŗo����Hc��0ఓ@�|�{�B��,w�պgL���HǤ��~�SĵԿ�i�&W�Q��y��G��j������_������>r�"�QC��7�/`������k�� G� Ӌ�<g�����^b#�w�4F�(�(9u��$-[�n�i�ls5K
h��E��+%l�d���\.U�(�Ar@;2���`��i'^o�ak�Y�ʩ6���{{1���*��,�X��c��S ����u�4^�%]�i���,�ZOW�?�'��|IW���.��ݜ��x/�J���z�H֛�Ym�'/�UN�X���봇�Q���F�H����#�dJu����l�r{�MZ�5��O�D��>����z �#\�����h�`Km+�O��������G�����f������g) �J�;tB}�@*Y��Ǉ8ҽ#]���ˠ���jA���3Wqj��==������ߠ���1�߇�r9!�D��Մ݅$c]�	�l ��5V^� 	� :0�H�5F��-vm���/_f�
=)$%Ԣ��I��mR���t�rh-7�c�����Y�O-<�\JB5����5��c}.�Q�ɋ��_�&͕�4��z��?��W��~`�ٶ3Ԙ��t�?��E[N6�ަ�?O�4�.C�jPAT�y}>i,ʹ��	뫙斥�%v���+;�(#����O�u��$�ڌ�Rs�����Ǣ����Ϯяm1��K:[�;���Ǉ��;��6�65�$���:�sk�r��hL�`%���4H�m�_�/^"�^�}��[1�u��4g�Ka�|8�&[f��Eɖ�|�!��AX����=�F����n�iI��O�f�y