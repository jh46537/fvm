��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�F��Pۖ\��C�����ց�w�8PI�Tv������}�_�`��G���~� ���M�F)��W������sxf9��]�<��g�)�@Ԇ��G#*w'���;�V~/������e~-s��)�B~P*�`���t�M��
�-0%���l���>�s�q�HX�=�(T2�6�J;�pO�  ����(��=.[�9U<��5�fs6���X-n�����+��C�����R2J�Z7��E�0 ~�^t�9�޽�{P�GhCm|^��aw���R�*<䫬9a�5K6:@�Jl4.��p���k�B��F�9��%׼��K��~}2[/���#��U�(%�)b�]IOAeC����`gVhl�()�v���R�����n�Td�\�(�R����я1O��Z��Մ�݁�W��7<}@^\B��O��k(�N�Y�@��v8����H�Wl�w��q���MNEhbq���ې���s	S� 3�����=�5��Е'L�9�i���C���:s"k��XHr�?nd��@/u�� �����K��ټ(r*g����Y�%vw/�j� <�臆��_��dH���R����S�n���]2S{�c8�W�R�|�{^?�)�����7 ��K�b�j/j΁�)��s��ݬ
49��	��K�˰��\N�'S��;i��l�{+j���`�m��_��:�FG{�{�����X�58&��_�1d>��_��X�����h�u���̻�-]�=5���q|�����Ic=���~��zc�,�W�;�G`m��ʷQ4��: *n����^�d�������j�J2�!	��h��H4c�����Y�[�xL�AY-�f~h-��p<0Ͼ����4���VuG�AJ�ez��g&�ԍ�4���II�&����������b�(�<����P�dP_��y-_�~5@� 9ڷe���v��wqT&ϡ?�qܱ��	��i�qy
��ʸ�3��7�e�5��|�APڝ��4�'���c�O�r�����)��Z]D�:lhz����z,�Y^:_{ػbʻm%Y|B��P�
ZM+���FD���Dl߮��-�U��~e�����:8�@!_�Z�����+�?����H,J�U����y!���F6�E�QUAx<�`��c�3��@�۴m����a��y&nsc��A���7	Q��w��`c;�ʆe+xF#�!/���'���F*Wv�!uk��33i�_� �8����/BG�GdEb�#�R�nIAP:�_�w�y�%ÍŁ��em^Z��;�ޙq�΋���������>(!jYtok�����p
��i�_w�$`���B"R�qل�1L�!��/��>���J�]�1r�N�g<H�r+:ZлA<�`C(�`��ķ�OL��7e�V�_��ZK��������~���8(�/�L�<ci�B�G:O�O���� �u���O�iP�AXX�>���_O����X����\����xr#	��z�Z:ϧe�g|�d,�C6B\)�7D�&�Q���TbAt�^Uюt�mj�آz���Y�$��L���k7y���"����hm�*3�"Ej���������]xl����a�[Dt�T㢌�/�s� $��`�*�nB���Ʌ6�-� �����C9{�g`6Y<^�]���U*\� �	ˮ����NEZ6U����N	��Sm��7
;��F���7&ֺ�t��LB�� �+��!f��)[fԖ�M�F�|�������i�7��.L�F�q��n<p��\MO��W_m��\, [ܲ���e0'�����[�V�nNޖw�|�{>gq�7�L�-��d˞j����z�z�j��q^|��D����G���*W�J(V� 2:��Τ��j>Bi���0#��}�`��uS�����Y>i(��,ăG���R�I놄`�퀡o�A�AȊ��.nH���Z߰ז8gcJ��(~��������s��׸&��o�kTL�s��肬�O��o.˽�\"��%�Q�rt�� 㰊��t��/�,�!�ΐ~B2cf��	R���=c�o�a��:zB��� ��|�&�!N�Y�
�Ly�;�aD�Q�Pk����E���h�=�h$_y�<|N ���
Xj��"��gtl��b� ���Rق�dI2)����R�r�v��4y��˻c���c<֭��A��ճ�IZx|�Gn���	�雾��Tv/=�ܿ�׊n=�S��&\N���f�����{���� �i?�;3t�R.Oby��d���M@��-�U��*���0{� &���=�_�I���!��遖|:��
Ғ^E��e��]� ��yX���j��a�:ql[�����Ot@�>����9}��Lm���������D{���1�[���d~q}��n�}ǮPnMW�u��Y���Ӳ��$�����m����w��my(��x��U���LƸk�u;j�M�h5t��3����ۢ�3�<�>N�Ya	Yڰ�)7��\�p��t�}���bD�>p���B�Q��ibqHY��Cˆ�J�"ws�N`��NDn��M��#4�]��7iõ��4<;��eA�`tڭ��W^�b�(��"VTy���b TQ�#Z+��u���=��a1�6X~M����X���8����ɴ#����[|�E�B�0�W�h�1��>�{����ar��B���.�X�\~�?؋>T�Xr#�/ܔ�k׌�Ղ�B�t�<(�i��I�%���)�K��h�*��ą�_lWۄ˦ �Zz�����w@����(�;bJ�b���N:���l��X�κڈ�������L�ݩ�9D�k�V V:�)��Q�U�pr?�=�I��E��BTd�OL�(
����N�_�D��PsS[����5�ҸSծVf˕��?^9�b�yY�:r ��:'�h�6ض��o���W��N�i~B�g�i��o8X�D
F��bC��Ta��,�h��N�]�6&|:�g�%��:���dJ��b�h�C���`�M�����I��Tw�4��(Aϩ�ïK$W頱��F�O�ѩ-�6An.nZ>J�n�'OnI,�&�>�����Q%�����k^�#�W]wj����� ��aB�*އ�Tġ��{�>����i`�al�O�_�U������c��w�(�}=y�.`��l9�og�� n�N��ӷ�ܲ�~��o����rMa���i��99C���U6<ټ� �Rp�׈��k�_�\��=0i^ԭ�G�����Q���ޙw���U��u*E���J����Yֆ���&<�h|��\cB�%�B�<s�Ш,����f�՟?�&�3�U��0vʾ�����o]�)����1���5��P�}�̉*(8X�Y|�M�>;Hl����̍�Шظ��mdԆ�X2V�ʁY�fl>�W��g�ǰB������ž; )y� �ⶇAt6�����q��è1�����i�$��?��K�Vq���ᐫ@���n凬�ćzc���(���}Q����|c�C���\$�qhi� ]vب�||�DQQ�ͣ�fV�b�L����8��j�j�1�	��h0�Y�Si�.ψ-̀��W�	�|�ck�Ƃ̘�es���6������2���֛e����ͻ9�u�Q�j~
ы`�Bc^4�n���՚pn�������C �I��e繾��pG<u1zZ0����?؀&g�;`�A`GfW��ߓ���B0�C-BLxTb�S��H���wMb�)�M�ו�B����y��]~���z��)�4��I�{4�;!�5nyգ��Ji����&��u��t�F���+R��d�����v��(: �����1F�ޕ�N5)�Xs؞y��io��wIj��%g0�"O?�Ĉ7|�7�l�OB;����M'�7���ļR�57+�h��
N&q��[�-�ȶk� ��R�D�,�Xs�6x�f��G��	~#쏓��|5Uv	Om��rQ,��Mre��3,޹�f���ʙ?����-�+Hw�������wr�(�J堹l�e/(@Q�HC/���N0?��x��,D��ZX���+�����{����v��}���y޿pd	�ɸ6?����ntr�b,���n��l�boݨ4媻[�=�ߜ��g$G�!&�O�޽�u�ekh�`��:O���P2^�r�=S׮���kSᆚ�0�=�؇Foi�p�,.͢����׭���,�����n�V{B��k�@(f��`�Q�cgn&���x#�?�Q7��B�=�f��a���j�99� }�_�l��>�I�p��,A ��L������Ⱦ���n?%�k���¹Q��Ai� ��$�@WrU��2?��~�1��4�;����6K��i��S�g}���>;�����^�t�/i�-:������v��v�G����˳ �tˣ���t,������~��h�+�GT��K��FM}��(��ℰj�t߃,�������9*�6���BTt�Y��$A�l��X���_���NT�kr�.��(؆�C߳��ș��$U�-���¥SMs�Gh|8b��&��;;�_��d͞�y�W+��i��J(]�~J�&���;g�g�(t]��*�`'nw1�7���I�p��T��g�xp�ZTt@���Sȓ�kr��ycj8���VMAm����U��4A���F���ʕ�J��O��w�H��ۧ�z�[�9��=n&�/g��C0d����
29�i��6��H�_ s'`�\s��������\'O�U3�2��9�M��V��L�_�`���R(jd7Y�a�@B�����	B�[1�+i?��Wc8����+����݊��ܲ��1K{a�u��(��|�ɮrr���Jzck�^�]��Ls��p�+:���mb7w���CF��4�#˄څ�Q�^�/��/|#��E������UyH���R����Q?!S�W��9ƀ����#J�F.�s��tKf�26HM�q��.��.|��+�H8������u,$�L���X}B���Yk�Ђ� �;Y�:c�8!p��9�6J���U$e�B����_�&🿩���g�$��1�9�Wеs|8LY�����p��T�+�zsM&�?��܉1ϟ/�?=I`���C�w�Z^���'��7�Kl�@!O��i���¦�b�u�J��x���rr�kߦ�j�o�/V���$�|�$)Lׂd��]�]������+�Kn"����b5&#f��/x*=BZ��c��)�47p;�:�i��ǹ��T��Mi��
���rM���� :�)L�0��*���O�+��/�*�^>t���ɳ�A�<��ވ��G�g���Vf�{�I�u�� �
�k��4FІo2��CU�X4c�vJ]9��S��S䑛4z�p¥��6>ix�F@�"�E�m���o�'In��V���h�e�6fH��+�C�l��m�Ѱ�g�Ǻ��NA!���*��s��iKO?*@�؟�s�Z�%h�|��$E/�䘾��� �s�nT��� '�ń�.�U��Y���ݷ=0�R�޲�S:Ӎ,1e(���Ӿـ6K=p]��AO��vb�5���ƕ��cA�%`Ċ��M%m�ٕ
����g�r��(
;R��}_�W����=�G�ҏO��xx�c�S�����3�����hn�������"B\Q��Za�P&������k�M:�Aotb�;x�i�����*��!��e�X�Ѷ�l����ѕ����6#%2��\(�m8�!��j.sXZ��.��vn�!je{A�G푔�ZA��/�f�ｈ����n�� �q�N��\ YxE�B�����e����d�9#㮮�=�P�{�Ēƣ�	<,��g��˗��ş�Cchv�_c*w��Ԗ��Ԃ?��+�w}���@y���}��a�%�'l>�̀�h�o�p����^�G���1����:�`�|_���E�W�2kZG��]��sp9i�}�T���(I�1�����_�v�3�g�w*P�㩕��2}�|�w-EH�-�_q੾o̇�<��מ�&WT�!��[��Q|�G�8����쬭	H�v�zT�ɝ��@�[s�Oxҡ��]�S�]p��pk��_<��b�P�Mzv~d�<�2Ǆȋ�
��W��S���	C��N\�$�or�:1~U��Ey� �m�@����@6d�Y(����HO<�^��$�#��~l1�M��a�\����� �SX�,ᘙ�f+řQٝ��ȶ�m8��\��'�"�[U�Y�g��,k[cvD���ϱ���{�ݎhȡ��0"p1���"� RP� �~Ihk�nK�e�EB(�����a�{ct�b��U����H�R4�&p�'�	G�sW���*HaS�F1ԉ��כϋ��!��8'���z�D�գ�.}B��3f�
�]�a�S�qW�H����l�-u6�R����4D)�TR	��0�$��٬8x{Q'��3��Tv�,e����n�Be{��N�07E�Pg�<���Jd��,�;�
IŬ��0!s8�q��5ߢ�l1y�ع`��Չ�`�8�n=K�$�:L]�a�	��D��X<K��#�M����|<�s�pKf�ekS)���ch�B���{�(q�b��x%�=�ݨ�q� ,QBl��`�%|�lA�f��`���l4�n8yr�R'��#(�� ����W�O�ќ��\��Ӷ�QM�J��!lHjob*��;�u���y�[{s;�I)�Lu�h�9��-�i�!�%�s�{X�v�ـv$S�*B�y|5鑌<2��n�u�[��)�"Wj�x�+�2�)Mfª���E2H<��A�rd(�Q���y&����p� �L;<�;	t�=�?L)Ƒ�}v�4oiW�3��kp���む��=���]���u�_��DER��#�.���X+�X�>yD�������Zr�w�6�������5�c���_�.o�u�T�ֈ����w����\�c���!�8&��
�����ы���#�&%�� �$�T��تlK�O�-1!�����@kj&1Yk���}��6�4�V{~�oD��ٯK�c���;��#�Bgq��A���W�$6��NH��_$δ�v��tE��/��m�5~��r���lp޹�����"n<72MOހ���	��q�L�>jK>���q��!ځA�Siȶuۼ��l�έF.����/����̴�V��.��"T�,��6p=L�6*��"Ӫ��]�tS!#6�:�����-�{*Zn�,�[AK�WVW�a�eڇ�ȡΜ�}8�ެ�!�e�[�Yz�̍�q=Yg��}�h@���u�W��lQ��?�/%��>v�v*>zvQ��ʞ�JOXBI�(a����	��3��8MM���O��m_x�Vu@�u�,iQPX)yr٣��[�جm������u̻��{�� d�u������ƒ�mr]�Ur���.�
�]��z�!���ǛRH�k���.^�gZL����
�#�0��ff���R	!�(!M�����zc{a����4'�؈�u�M:�E��շ՗43�����+��/��}H�r��L*��3h��_(�b#�=��.?��t��-
�Դ�BK,P�N�-TU�>��&iQ���q��_�[O�VFZ��en��փ!<�.7�[�
<ˌ#�#��n����	-���f�x7�0$AVF�MK��;c�et�n4 ى�ԪY��|R_���-(�����M��Eۯ���|O��E\�����Go�C�f��}�J*�-&����:Ό��Jf ��ϸ����7�H6�~g4����
:�u߱��@D7c����E���`�(΃u�s1� qO!n��yMG� >\;�8�uM�ӎP)9+܋(��8�'������� �����<3���W5��'+Dq���Q�N��B�-�_m��9���C߹�����h��}G(�o+��S�e���]h�yآ�:��k���}�S.�|��o��;��E�V���B?z��9/�Fi�]�gQȨ��J�ɼ��:f7[f����x:ĔR/1S?�XXG�Id`~ԚDSe�
��[��m%��_�����`�78q��<�-,C�	�\[�I�?���\�Z���{�HnyA(��Bur���;��5�t��=¯�{��M��d�$GQ�n�q��ݶ���c}<���������QL��Ihq����K�Q��a�S��� �$i�ʒo�{Y��3}��<����.[���J`%8��?�m>&�p3,�;�[vL��M5hJ͓�%cr,lR�l�(�iS�&�ѐ�9L�y�
�!k���\����%�I�`^�_V0�o�`G�,��.��QU�Np'a�U �%����X4�j�z�#�>hC~ӾU$����8t�b����x~}����.��q@�z�j]�&M�&�iypd�eĦ?.���.��RTSW$���/�!k)G5��͕	�㌚=�K��f[�<H�,���"�R��=0'���D�g�u�݉��L�' �^�@N![tM�dt���J��<o��=�v�Ԙ�*�Mf(�|���'o�c[�6�`G�B>eeM�Y,x����
-&4�&���~�u��s:6rRo�N�ὭiN�n���߃'2}Գ�m:��<�����]��O�e�L���W��~�TٓW��0'G�2\�7�ʚ�o���������4?Ҋ�*z�p���X�*D۴G�Gغ��0D�m���������rC��[7��������-W��a��BD�1NKE #\1��B�1�� ɏQO��6�� �~�FwK ��t�t��م_uPx�@�R�-��v{��� ��L(>ȋ����
���-�����E0f��0���P� Tk�P���0��8R����e۽�B �~����a�������N�l�#������O��◒L�0�Y��w��h����$S�p��cu"H��==�XB~+�G��usg���a.�/m^����E������܈���~5�٤�����:J�1L��?��d̶]�U0ۙImp�!�@knY�<�l��������[�I��$����`�鰶���K�)�A=� �d?�ͷ1u��g�	��R9�K脶,��UhS�)߅�%�Ǡ�c�&�r�[��
O{�ta��Ɣ�IG;��=� �����l|�$���3�:���ǅk��,��$��h;���3�tC`�Z	6KHU�̋��ztM�9�ji�YX|��j+)�z�A6���j��M	���ԺD~�o0;���vVN�/$�����缰���=�� Ќ�D0�,���b�D�Ʋ� Bx$'�Ĕ�,#޽�g�U$�ѽ�[�y�S�43!�xv�}z�H@D7�p.}Л' �;�;\���㗙xu��]v*Ö�K8����<"�� �S�,��m��<
�0��t��~��� �?��?I��>�BMjm�7"1�d���1\CP)l�֙;&��%½[B�t���34�#1�>%�Jd�Y��US=-��n_k��U?�Û�l�
��:.��o>?������tc ��}��*Z5��[�������&�K�)_X�ț�V���c_��ıp���:C��N�:��Br�y������?lVɟ��Q���\�����	��0��a1{�-:���j��<2y���s.)��ј0�e�(�}Yr�Ga�q�í��+��]�͑�;:��Q}����zd��R	�y�ЭȖ�ϧ\k!ӷU�s�=hV��m�=�F��A2BD�.Ɵ�V4fV
̵�(�}a'@}.�������;��5$���yA��VA+��m���Mc1EYW� �p�zV �'~���~��Ts@V�����r
��A�1�Y�T3F��~���5F�#/ˍ[
�.�`�k�
�-'L���2���K[����@c�D�H�޻Ú���{&�U���.�Ʈ�.��u���H>�8��ngZպsFH���I�����x������>�:���H���#}� (�k���1_X�Rw�B�i�� �wh!O�.F`��(PWX9��J �����2�G�{Rۇ^�s���h�G��SG>�&�6 M�y�Z��r�J���MۘE��|%�=�n��)u-}\��u�<˼�މ�MZA6B��7�҈�������
hDG�6P���������4�g}���F
���v<��z ���vo� Qբ���Jf��9T�R�o���E�p��e�fmne����B+�-�BM/)�}���rS�G���RՄ�t�.�-�3�h��4�+Q~Q����31p�	/��=u6���0<�B<�����ds��Pk<�ɮ��+�_�^;c�r�0\�/�ي��*������8KYEQ;|�5�P��9���Ga}6 ͦC�����4�]�dl������:
2)T!^�0�{���,��VN�8B[T1(��̓r��d�u��#KQN�+�_�~��u��i? }�ϩ(�b2lSӖqLӿQ�n����Q0pp�E��mȴ�;� ��a��2�!̕Z����W3�ni�{��"�T�؞<�7��7C��?�!:P�k|�&�b���A����g�Erd���i�k�$�1@_��g࿍U@N�*��{�Q���uǍ���҈FʾO��y)�Q�OAC�8s�c�'����w���_&�0��ˤ�5�ԝ���X�em3At)�)����y,kW��6�M ���e��%�� ��w`?e'V���G�x#d8g�Anx�<�Y�B���6�g���/��S�G[�ۉ;���&x'�z�-����>(ؿ���c
����,�39�nBD����N�W�˃���#���Q�Gy���Q+,r,����I��R��g�P�E+>��4����g�	�ɁGI��0�;Ո��c���DQ�:|��-#�H6��l��J[Cq�F���h~Yq�u=�0څ� 䕬xd��ZY��+�	�>HUg��}� ���n�-#�:�à��u�����Pz�6)&`��鱂g3�׆��7?�����9���"�I�3���A���С��N6Ɔ$}�ݝ��U�{���l��U�W皃�I&B9{߀H��+�Û'r�$��aC＋��#��[Wa�I�~����F��_ꛑ��@G0�:X5����J-w�R�A�y��Ɲu�=ш��gY׼���frNq�Qwε*�ޏMV:|	k7�ҺUc��:���b�� }�Bm��W�5����F���� �G��Ւ�Xt�$����t����Tٳ K�ρ1��t?PI��ף)`�K_����N𧉀gD'����Ԝ3WV՗z/�J����Z�q�==�"�6����۷��ڠ�)����#An��S��5v9Y<�8h��Q�i6��'~L��T�������5�.}ㆣ�+<3�Q��iq�1��f4�?N2ROezW�я�u�Y�pj%^)��7%"D=#�&ߟ/�ue]�������Me�l��U���������c�1R$�}�hcl]��A�EE?�{��e5��=���)���=!~tW�U#�K�@��rv��P�6�<gz=�ş���ؤ�H�{�s���;���8�2a8�>-J�rAz?�*~�M�}��p�?^�j�g$���4��6�1�w�=����]͡���ڟP�!��4,��,,o��7��Q�ue.��������$�����	�5���#M��a�I��N�*���-�ꏚ�����fK�{C?vD����o��s���L��;oL�gY >3�\�*Ď݊10��kk9��kg#��q�.n;
�Ur���'$S�����U/��$����։&��)á�E�G-��z�5W8Bj�&�M�� @u�\H$	gw�M�,��U�ݧ�����
�$�LR_;R8qT|��<�pky�5c�w��� �� s}�k#,Eź��;��̺�:����z�g�K�t��SC��	5R���w��҇Y��1����);�|����[��l���A��9X�\Y�MT�PB�g��1js;;�)��f<*���4<>��� ��B�qpv���>h^�Dh�Rl$7���7x?l>�Y9at��S��r��sfI�� �����JM�.,n)4Σo�o,�Þ�V�~:��?��\aG'�WS���uS���;�[�V<=5��},�b�W�
e��u������K�$[��<�HX��a�W�~ 4���=�Z����sGu�,{���vK,zL���e�oM�T:�GS�Q�ue|�T �m��E�E_�@F2�7�j`�l�R
C=<�J���z��d��e帹W����	�{X�
� ���XS����i��Ցt�xb���.�9�$%:eJm�ڷ����FzV����M�L��mP��n��8Q@ǧ��獻
G�Pu��0o���=��fx(�^��-��f�qh֛Pe������s���E;1!8'D��jY��c�����v��������oO��BGcj��e0�L������P���C2� ^=Y���p�[=�2yV��B)**dWl���g!�q�w���ZD�y��c0��ϧ:���CTCa�� ��]=�f�%`- IF�# �.149V�M��:}:*Ί�B���G��D� ����$���R�t����ί���I�Q�z��)
~U�O�oL�V�&�2l���r2[c;�ʯ��ź4�'��n��=P���]�C��1�(��?vW
��:<���	��'d<�q�J��1x� ,���Q!8�nǝo��G�]�p_�)�n��ɽR������O#�֭T$����,3�e$:n��8
�R�s6f�?ɸJ��9�L�u_Ǵ+]�5|������Nc`3)�=n�~�Ї�!(�b�4�*�d���0� ��%���M�;�.M%��w?��w�����>�i������]��w\`�������o)���wWz>\�;Z.�׳��5�vz	ˑ%\)��5�NE�D�pnA����O���{gG�yg��=;B�|�p nu�S=�Z�B��Rͱ��x�0�O��W�a���GIT I8����	��c���GǤ����m��o���Ӽ�	�����w������V�T�Te�y�H�m�
5�ǵ��g㉝?�"��О���&�=ߑ
ŶƊ̴� o([�*h�Ei1R���AL�_�_;�[���C�����3�8������H��������dy�]ԃP�6��y��a/dt��P��/��D���A:~P �L�c���;��C����NR�H���Bܑ���#�g}�<�Ӕ���:C�ah�u�ij\�.�pn��s����s�,�^,�	gzl��̩�<O��W�pj'�Y~e���z�R��@���iꎍ�:団�(j�}]��~֕�\a�Ms�1hF^����D]k�tcѝUIc�
�f-9�
����-w�	�w����x�Z4~���
���ɶ��e���.����+F�,ftU�x[����VLy��W���_Ɖ�D
�Ӥ��B�ů�	�Y��ʈ4�었�����ĭa��44ir�ٜ�9d���W��#��i˘�:�1+���2pE�B�]ߺO�fKl�ޜ�v��gƽQ{{,�:v��|�v�ݽ��d���X��f<)��Hu�J7uѶ������JSi9�܂�G�/��d�બ��+��He.E��vf��Bl���8n�+����;��?ɥx����?#>W ��~�z�bb���ϟ���Ģ�D�B���m���Ɩ�#� g�l�ُ�u��gt�'d��"H�c�ɽ�S�β䊯��:��v`,8�ߙ�	`�]��)I�]�5��Y;+�(�[��ֈ*����&���(
��ۿc��3 _��C���ct��+#[숞���S;�L��4�<��2�Ǵ3���&�s����67�G �C�Fhj������ޅq<���Y�¸S������E���ys4��́�>M�h?yV$�.@�XUɅ�����̒'6��nU=����gLDq�X.��&$����ݰ��d5�~Y��ctvi�����1� ����&Zm��P����^��uʐ�I�,�����w�W���bu@����
l#���;i
?�%1!z�R��g�+�� ���O���cJ0�=O6�C���#�sҶȣ]�tk�b��|�+O�ί�BRr��Q�����rd�i�6OT1/�4b�̤H37�L�\��lز=�B_ޚ�E����Vg��c���hZP�5�j̪=-"�$��)P�p���>�-Z�bdr�AJ���?3��ByO����@G���a���y���㞳E��|��06C��fp�C���FIՔ0�(�E���Ky`��a0�
!�@�z��/Ї_�����\ԏJ��Fm��\΁�'#�޲d�:�r�F�p`"���xQ���J{�"���#O����6+��dp����o�����ⲡlk�����E^�ll��0�@�X���1.Sh]'|��j��ޢ�E�K�� n$�M`dk8���u�g��+�6��o����L-7��Wo�c��B��c-�ޘ��%�S�d���.�$�뛐T���O��+ˣ��Gm�\S���a�U���/���
�K/~��RF˥KފC���_���0���U������RpB�C�����o��\<�v�+�J����\���y�@E�6Y� ߇'_�-v�^D��ܠ�*t,s� N� ����@���^�/�N��I�/f^��s��ے�') ��}@2e'�����10Ƙ�e�?c�:؉N�)vl����t�{�ۏ�D>���L^S�jh����sWoWFJ��y ��C�yˠ��yFv�|�w�8��'���*s�>���|���瀮�7���3���X Z�2f�U���� l" `..}oז����s��������ެ�'C�H����.�c�0������6�����V:�Ҩ���2{5���ة��j;���M��1Z�~�������� ��=�������H~c�MK��;T�P�''V��;":R��T���硩"BQ@����Y*i�lN�_�q�+�R��9���vQd��m,A�!|��ݫ�L�`�	�Pf��I�b�������$ ��KD\������S٦˨r�Z}0F�# /�h�F�z�M�)>/e�#'���]�����_�^���Q=絭j�J��7©�9�v+%@l���$��f3�L��-4~�*���P��Z.���T�N��VV'$�Jm�h�Ȼg$�Wg��gݓ������@����k����j����-�G�/����Ԝ�0�=��Ǖ@؅b׻j��z�!Z��U��\�/���-�s�}�P�+���?��<xdj(���T��z<9��������^ԨDN}Z�����E��!6o���m���0It:����0�JR��靳rEF3��^�^���� �H��}�;+��ϙ��O&��X�PHTYk���Qʸ��e+�g�E��Ԑ �����K�^��{c�Eq5��X`$����D�y��?���#E������P���n�J�O+��I*4��|J+��iR�4<��a"]Xj�ЋZ_Q�e9�A���t���8=�����^���2]���ݩ��\{���B28y��4"���9�OD�)b �@>ǎDr�0�nٟDz":���%ˏ���&���zUX\������ Q��& ����잚���4�t�U܉��<w43uŎ��� J_�U�\1�J)�Pr�j�+�8`h�|�s B! Uo2��CH.6�
������[�?��׿���K����(�Hv�D��k�򩆿�b��A�t+`|�3������p����`��U¤�����ĵx���^B@1�d P �e�3;i�fj�Ai�!w/���O{��g(V�^1n�X�6�D���_s^눛s�
��JT<���G~T�bYQY������5d��vbǢ-�w�R_��:ŏ�w�[��WӤ$�2��!���9�φ+�ٹ�<V�C�LN��9(�r��%Q�M=�Z�s���n���6������A?9�rr%>Ⱦ>��b�5���_�OX84�M]w�p>��E,[�"a0�)�P��)��<=,��"�|<t�;�j�;eB_R�G:N�D���(�^ i'um�B��<(�?t�{>E^�CMv,����)@G�Pu�W�;�g-��Aַ��r���L5SKuL��3;cٺ�ܸ��5��cA�dt�0��뭧�h^���|V�^��vjFݹ�Av�U3e/7�nw�[rAJ��_p��=O�FA������8h�n�h�~ �4%������ہ��]6��F:��7o���O���W�p�8W��IQƉ�);��yX��n7���E���ci��3���w|�W@7�}����6�4�9$�xNvNy o�V(n'��%��v��#EJe�݀���|���H�Y���%bg�ŎY�}�r�������nTYH�a��Q3�O�SIX�;�op���N���-��w�-at7_{2�&�U�
'c����Xpŏ���[�Z]":�T3K�	kxXd�˚�ٗu�;�:&���($��-����VB�t뻢犙:�Zw5i�(�ٛx8ľ��`q����M#F�a�/��ma.�q d m'�˯.�B��ۙ���i=��C7���s��xNߺ=���_I���ƕ�21����mRW�
7BZU�f�5���|�]��*ROv&�}�],�ji�$l�J3�����o+5L��f���^�/�$�AJT���f����n�e��A{�r��m{�@�:�G{+ego�+�&�hŇ�x���0ԁouJ휸E��s05Ȇť�JV�dT�o�w��~�J\Q.�e�a��	�
Q�'�6��S�w�!#sQy\4���Z��m�NB�ݲo%���ۖ��a(<_�
�ƍ�tp��-��� ��F.hŚ� ��=�'C� A��'=*���cF��4q�{4�Tht�q,�v{-1�v�s�����S�͘A��\\�$�5�_�GM�e�I��2��3iP���0�o0d���IP���"FxF�I�1����a���|)�F�(Te2���>���dy_��w�s�߁���r��9��&<6�^�jQ�hhҊr�b��X�Q�2#*I$
9�sv`��ud��b�?���ߦ�򚕗^��A�z��ׇΨM�R�	^X8U���e�'e`���v
b�cnj��Q��!� ����h�l1>�;����.v�p[^"�ru�TϚ`7��^H�Fv����@�6��8|1�������{q+�n����z���1`��dY��)ru�M�(f�!Fw��*����u7E��_kR,���o��t)C�Ƅ`��ɚ7�w/�Ƃ73����Brm�l�c$XN�%�rA͑n.8֚�<C��ZNgʿSα�	��0m���]E��T��Q2#�EJ_�0�y������Pv�bc0*���촨���n����6~?�H��a�QL��Ռ2��!�aEt���I���-�}�wc�v[/��v�	Yqn���D��y�w7�A[���P��L%�͵��9n��cfk�����dڴk%�^J!����A蠑��*�1;1�_ʷI<������W�{ԹpY��y�geHk����!�_c:\Ǉ�#�+Z��S�ĵ�T�" �_y���x�x^��?�@�%�j ;p`z�K���ֈ*���A���#�@sc@W���A��;��ԿiC<.;���vV���}^>���g�z��h{�p����5	�L��Vm��yl~�����0-�C/���{R��T��,�FD!0ݶRl���)��a�nwn
��#k;��NY>��]�X5H�ջ;Ӆ鿫�d6��%���S)G��=Aa��rB9ϓe@������4"��.��N����xt���lf¼�����b��@E�~���	�������P��\��!q�ݷ7��)�}o�69/�����Rm����#c�@�����W$�����:( �7yO��"�gk���f����Ì��?)SJ�\h���`$��МĴ�s&A�R#�L�x����p.��~�Jx�I�ӥ�Qh,Y���P�e�������Pl�vEeo{�=:��_F QZ8U����:?q�D������'�d���{���[��癳��s��r]-�*y�&���ߓ�x	�,�5���������j�}*��P�9aa$䍅x�C��E�l�sq��P�i��'�uD:3�����k���_.g�,04�01ӕ������	�����L�Ҝ�S��E���Wa�R�u��F��.M[:��ᠹ(f`�+��U-�������5XP�`���&AO�����}Ѳ�ؘ�rO�H�30������~xb��/����-�e}�|b���s�E�wM��K�Cg�����4�`c�_I���EDG�zS��������lC���`Z�Ml���`q�!N�J%�g�����E "Von�֑ ^�;t�����MP3�A��%
���Z�s)笢�o�Ӽ�);��-�y�Rv�]��jT&7�t�P�>7C{��[K/���g�������ܵC�����	k2�W�T,5�����>H��|�]�O����L8~QR2M1:/�g�d��僼���i:`GT�M\@F*���p�-�dC�.�3��)e4F 7o�{��0����w�(wp�x���J�D����!~���_r�0P�����j��x�o��*�s�O^ۘ8�e�I���I�U.4g#)�3���L5�TC����nU�pV@{|���I�\Vʼ�9!���I-�r|��%'L��qo�m��L�A�D"��Đ��އhA�V�� �{ ��r�L�Folړ�3�9b��[g��H�LKQ�kk�\�F���'t�[��\�sS����~\��2?cf���O����#>��h�S�v%��$N E��Qr���
��x��h�1$V+h���S$Z2�,�������:���{����W����p�kуw���tʁ�Ĕ��a,�lO ��W]��z$�'�ΰl9Ȓj>�~� ﾡ2�ڨa��x'Lޗa4����7�O�mַǯ�u1��h��3�Эke *�W[9�����j���RB���h�7]�0����������3'�Z��cʂ��6��5���l��I;$==�YQ���jO��U#�b��v_x&�h'2E��d*��֢�9ǟ�d�r�f����K��8F�\۵�~M�����Ͳ�A�-(��ء�I&�y˾Ӧ�3������D��JJ7L?(!@�c�. ����l��x,��2��<[A�1q���#�e�<&��:���0��AcTX�⥡�<C<`�M�lF7��|���O%�$Y˚���uP�������(z����sȁf�;�u�]KU�W>�D�qUؓ'�VW`Ä&7 �l��@��F֒��
v���\k)�C�+Gơ1j)�NpC5���9P?G��m4�f�� qJ�x��`T�[3�����z
m&�M!��c6�]�vTߑ+�i`�Z�F�i/�5�t���=s�&�gk%9�A"���{�r:��� ��p�[��[�:��k�5�w�<�M�XBR�U-��΋�҇�4�ğ�di�b�s��%�o�F�ּ�=ahR�U��T� ��[��Ћ"��ޗ/|�_Ѝ}i%�"���pI�˸҆�
ג!�뱅��@�1�S�n;ܞ��Ɲ��*}�ſ~�C���0����1dg���$�V�,1�5J���ݮ��"�v�c�%��v9�uUP4f�r״�͍̕~^^���f�-��/��{�tv?��^��3F����֝N�j5�Q��_A���b��-�.|�l�@��� �2��e27����fl[F�J��3�4z͠���!o%��1�8�$%��(���_f�\[ȚL�BN�-�Q���[O�j��=u��ׅJ��3\o ����3\�k�Wd�Q��W`���0�С�o�E��c�Sc���8h��:��ܲ�����Xk��.��Y=�J��&GB��w��ۡ���a�b�A�,���,�_����Lq��_`sQ�<���7�Ux�ᭀ\��M��u� ���c�.����Δ��x�t\�\�����u�"k%���D���Q���,��j���!�����yI��M�5^�ݽ�Վۯ���)
\d�%'�Fw�����s���� s��ѹlT�v�4�O��S��!�T��M�� �[�o~L�gy)"������h�5�aB�d`X�ݟ+�D�e�N�Mk�����X����^ �ύ��6�s	�s����b�c�������zrNFdW�إ�Q	�dnJ�p.HV��B��x�l�� �����b]Ԯ��#mY����P?d��C��v�D������0��B�._`�}��"���e9Qp̏15]�<�Il(|,�w����l��a������Y�����L�Rv�|�vԛ�4��k4�W4`;H=�,�W�!G*��3x���󟒈{��O]Y'�DM�d =P��%Prͬ@R�]���t�nT���Q�K#���.2�M=.�6Gj�׊���ܺ��~�w8 �
��=��|���񺎉���L9������r��sm�)�j���F���NiOS����@�����ʖ����w��Ż�����tgla?fH:f��j�,�$�/�nR�L(���I�d?�5U<d�]� C  nD�B=��;�g�<F��@	}ngE�8����������:Q�-����Z@!���>���	�F2[���C��8��WྃL2R�p9AY�������u;Ȏ��`��s�&�'�Q���,=s��^��Ձ��(�L�,���
��RTR9�,�	*�~h/�f�D�!P��4�.
��^���Í3�>�L nH!�pFvj�.F�a[4 [��
�0�+%%]v^� =uC9h|>j,ub�lh�_��f�U|�{�����Z�r�B	�׿0?���8����Lc���F'0�hn��}�!�ƵB:A�_hD�ql
���C����"j���)��8��n�w�=I�P�]n^*��O�Q����>!4}�uaI�"0e�i��涳z(����� ҔI_�2bȭ��A���/�?k���$�JӤƻ���p\À�!qB=�S�������sp��w ���ڡ�6���)�/�TI�2-�U��I�&29Y&4vÂ
�
Rt���Z�Y���d����Y�z7�)r�ಁ��>�Uf=z^�1�;���qwW	�2G�o!�_ L����oȡkaQW�d^�M�̈́
����(�	�)cG;s4_M���̻�}��b+6��s�V��$1߇W���ϐe۵�s%q;�ə��*�x�i�9>�qJ������S��$�m�c'd@.YW�g�����Д��C�	O�X��Q���,2���T���:U�~�o�	��Uw�m٣e��	��I51��p���ً����nDb �%�u�+K@�t�k˳E���Dl�+�o]Q���RX��,K�yl�����W�4~ۧ"��k �����h�C�<ِ��Yʖ>�4��;^���&v4=�A@�F�7]�FL�p����7	�Y����(�h��Tx���Z� x_�XkH�w�iŖ?�����/�J�����lc�5Vy`�?��_�8�H��)@��g�i�9��\�nZr?̶�}Jk{)��K���^ſ�@ɧ��8eS��H~� �0ho�Y�+��p���̯�g����f��T*��[GR�3�O�����QR�-�Y�B{� ��*609*| �G/'	���N�ȴH�/v+�mB�|Ը��G�N=}�/.��~��q�>+�\���-&�N
�!�;�E)�iՆk���,�E;H�������AS��`���MP�1gC(Ay��ĝ�F7��MR,�s<.V<i�����r
0J1�NeG������Wb'���΃�'z
c�ܵ�ÅB-.@��|�x�3�y��k�ow�G���&��w���v��d����};׏��n8Ho
��4,�^���R��!�a�R��P�O|�ǭk�۸��h�e^(F߉�2�m��Y�kL�)�7K���oJ�w���t�+�[L3�Hݦ��졝����r
Y�⵺�_*�i���R�M�(d�ꨪ�#b�7�����s~�
�6���.1���V��M,�f�Cq��!9���/"�(�,XIK�K-x��1�W���k_ӡ���od��-����'l�Zq�`�R��+3{�s��sa�psߕ긲�ʭJo���+��LȺ��WE�Q]g (���\����lQ��&�/�>�FEĀ���i��- ��5�ϣQ�j�f�(ژB����� ����v�ȑ;)X��E%��q3ौN]Ђv�8���@'t�13�-��{�E#b�8g��|�%��oh��p@��A��ŶI�JV� ;�pt������M��X��>rVpt�q0#��@Q��\�v_\,&|"���(S=K�{������z��PTH�Fw��v�!�p0q@��"�0�}dw`c��	O������!ē�X�4:{���S���.T�)��S_!�N�7�� 0Z豤W�1��N`w�K���/?*�%o��J7}��1U{��{l�J"���缱*�(s��jA�
d �("�������(�w�������ڏ����,>���6r��<�O�@.j68���༹B�_�&
��s�����d�\�]MXf�%H�-3���/�}��|��DZ�/���~e��qS\�9��l1��jsvh��*Iߛ�z5!�uY�6�����q�J�e�r�DGڄ�=UX�D'�E�u�E`E��X1it�	���Qm�B�np,YS���L鹊�l.k�M��t�}����iWm���y��p�&�ґ����.Z�F�T�|�7���RU2�����N�V;�-ݚi���`�8P��/�IM�]��N%3�g��F����=/U5@�@�"v���Z�E��H�O�W�����n�*-lU��8&\y�J��E7W�M����+�&o���� ?j#�Y"�-� �L���"��S��u@5�;lU�̖�9��)ߐqD|��ah?c�����?�{-�h�u����65mb� lEJ:� O~�^��ljw�����T��RQ����S��n&B1�h 9�e	xx��bu�`_�L�H<�3J��eC�NSzj:G/p�ɰn�͸:�V�7˯z�a����ծ�H%�����%������G>�y�ҁ�����O�9��ĩ�C9b��9�z�fU�}�M�uF�J�๺��N�eP����ߥ���C�1>��+ɘ��;�HC}���-�Z=RSh��yh��=|Q.���*�%��2(@5BK�S���R�wN�:�M��y�ͬأ+��ڲuÕ�Aaf�`{p��f����Ѳ1�w�0T?;/�	�wb?}��B�s�0�aA���(�,����s��m!��Չ�
|o�Y����?����:��g���-��a��b�`1�B姿���K�*/&�FY�j��mI�"�� ����我���]#3�o�S�*��V>�/�×
������d�:/ؙ�.�z
]TJ��pd���zB���?oQ����m�3�~���(�n��2��z�O���x�޷<���/iczP�Z���6��\2w���%(���e�ʯ��9���C�6Ǽ���#������,�S�[%�-S���2������Chf��
�#\��J�U!�4`ܡ���Q�@L�a�O�6}{x�Fо|���~G<@ւ>���nd�EH���_iC��by���K�A.�#���Go>P���G^o�]V!A2��~˽�z����{;��;�:�'����h����[�>,���E�g��gz��l�hrw�Q�/�NP���:�2�Jٿ[\<�:�ܾ���л�1b�#m��L�=��"��E�wSk���(��À�Ź��j����rXP��FZ���O1�BҌ"e"!��f5b�͉bhxzly�D��41�T�V]��2V�{��� �9��g��>�����UJ�#n9I�`<�oݓ#�;�\ cn%�Se�n����oߵ�(��S���%�0�Y$�_�/��y��UC��G���Pf�����W@4�� �� S?�{^��}�
R��%�����_z�Y�����%>˾�l$��\�W����/�!����'ڠu�	?��".	�k�㞴�b��{���Z��Y@�_�B&j&���X7-ަ��B{���}J���A���9g��3!o>�ޅ�sC�t��/}$1զ�ϲ�AZ��F+~I���z������	:�Y�L��\�@��&Oa�3�ٹ񋬨8MW��U��E�N�4Z"s:{�(���?ۚ��|�;�n=|�)]$T�?�v�oxg?b�Y��7�"�8�?ې��FYKS`��������jI:aQ�vn�V��W�9�TC��[��~��u��e�b��Ɋ�j\<B��G`X˄������h�A���5pU-��b��(?E�F��m��]R�>-үR�ɽ^S����`1Z~�ࣦ��7����o�:q�!&���Rf0�	�t��t'?t�uV��p<ҭ�*Dfֈ������{nT�y�L�tފ�!�`��9D:-����&��dᳲ�������\G҉��v�V��8USpS�39 �Ma֬���k5b�יcЮK1}P�(�~�(!�#F,D�3|uB%ğ��5( �6|��*Y��F�b�3���w�5�l��4UI��o�#�m��/�����Y����Ea��]���{5�b��ŕ�u]���ł�e��ފ`���|J��2� m��ge�]�t�ua(�!���68u�I��=���^�D�p�����"���۩�M��_;�ׇ�����������yΊ>��xh���!��r(0��٬�6bS��7�������ݍ��o��2���x�k'����˥����� ��:^ן�t�
GJ~Oxf}�r5׋�~�ͻ���@#�==�ی���ɴro�Zg)�����.Ak6�Ւ�`�I����fl�Mh<�h�J�A��Qd�Q>`Ҧ2q->
�?�xؿ���Rr���ә��� F\�@��|�$%cz�q����Kk3�>�����f�@�&����%P��R�_��w���&��JZ�;v�J�d�]ʑ���fL�wJ:�=�[�2B�\��g `1��6������c�{�#D��Y�6�J#c�	��11�/����zY��o2�ס]p�9�eK�X���·��`fd!���F�FF�ـ�H�6���7|A�Y�U2�L����b�by�v��"��&V���n�O���ǒQ�m��u��89ef;t��=o	x���ɼ���MaX�yT��$���H�n9w�q���d���{� ^c4���(���	(>��_�o���XGx�~{����3����@u6����D���3�p�>1���/c���N�a^�؝3��m�t#��$gw�=�u(ow c��5^��뾎��3�r�]Z%{�*�Ѧ��ˈ����3��d4��z
��j�5�}{�CNp���4� ���U�L��P\�����X��fcl�W���|��A_�m��+=�o�Ƕ2��ղ��k聄a��s�.}A_c���m�#�&1b�:���^{���a����b��KxǓ��ړ-å뿁�3{��i���h v���-�Uf�Ccz���^�x�k7�|I"�2k�ݻЉ�TG�J~t�<�������Re)kZ�5�֢ ��.�s�7�*����Y�o���#%�W���2P���Hu� ����D-�������_ʶ�V�b,Қ�K�K� c��@;�߈���宋��H5��<i�?K 3>�W�#�(}���g���	��:���
��J3v�͵	�? �B6i"�_qN�l�:0���^������1Bנ��`IOC�ke��=?b�y�f��.˨���.���3�S��y��6Z�,R�U��X/J`���4�սK��|���-�
x�dV=VI��7�`�`�N{(��������.Ǭg��d�l qD��a�z���x���nK32��T�"EZ�Td7�m���X�x��g�b
{QIX2�L��qw���~������մ�����p&��em�;�a��bÃ���D��mx��E^�����&�������� �_������T{�OY�SΫ֧?���d;�썑6�G�_�F��W�Y�p9�xJ��'?PH�M>���5�kPU�o�'{��
ė���C+фʺ��i`��Uԍ��F���_�3u� 2D"a���M,f����w]Ʈ�(?c�*�Of�:��a���-n�̓����8��?z\�B���l&:7�j�u��}��)O���'��"����X�T����^���$�AbE��3L6j\>���	Q�}���f�!��2l˷1��D6��`��x��tm���"������SV���P2���t�d!{�(\� t�N�mkm*��}�2�S"�c�R��$��g]KR����}ӕs���� ʒt�����q�������p���*����5ݱ��g����>��� =��jO�Ճ����w)>��B[r1�F��C�ּmB%:�&��a������G�y76"NcNT��沒$�e�W�i_�8V��
�F����<��NR��Kc
F�l��l�|�U����D=�O��-q���~C����%�w���2]d�|
F��� �Ʒ�q�SY�fY��ň�wa��Z٘��������OJ��X�j��ڧ�k��Dό���ߌ��畭r4P�ȡQ��jK�Q6J�������lOv��% �I�.:o
F
@��&(ݩ'���Ga���-Ѣ�
�DP���)n��p����pw���9s�X@�� ��fpQ�I�l��Mb�D��#G�a4OC|BV �Ϧ �*h�C" e�k�\��GI%�%�C�~���DYbx���{x�_U*���-��U�]�N��B0zqZ6}5��a?O����P���,~�yΖ���!�){�t��Xo��4��${���eU�H[��2v 
@��0:*�>��ːG8߰{/�Eh/o�	����x@)�4T�<��?
��eX���$/!ˢ�������V��W���� �L=�*�m���>��K#C`�'%��w0�ڑ�b՗�.��w�/��\ێ����׷���Lpf�U�^;ŕ	�w��'m^akDm�3�� S�����hKjI�4T'&�yB��S�g��ڋ�N	.���L[z�l��ԽI[}๸���\��M)��	kք�����̎y����u^3���%%���CF��V�^���*��UƉ$*a���C9�f��&�v.�g���l�@�����p���2X�9�٩��}YE	*,)O���"��H*�%	[.1�����O0���'�60T�-�H%9楍�I�v]G�����n�.� \9<�!V0vS��d�4�]wc^�{�c�LW�<%|P����HT��Ջ�^ٜ��[�/���(e3� ��u��K�>��tb�s~��s��o��P+�E��s���ɹ��?1��OH��1_Ϻ�������^bLk���K��9�� �Cf�w��2��`�=���ڛ ĵ��-�S,��Z�'T1�{-�z@yIIc�L�ۃ@������T����o��s���/��h�}���ş�i{\3�M����\��q��h1�¹�@߱�ҧ�)����^c�eԱ��-)�p�O��E�l�I�3���bPЋ|�"����Spɽ���9,��a���},Ai⻂���%=�'���CTַ
$�}G� �~�~�5_o �Ҧw��k2)�=)������$r��������� ̞@��*}*��$��@ ��g"��RP���98u���ڃP/�']"��*�;j�p΃���`s����|�ú�*U$���M��|e�ø��oD��LFK�$K��z�R�=x�䷉�j>��8��<���:���\�q)��]p�7$��(��P���	��D۰���P NW��g�C���A9ue|T�{hm�L�rj-A���;#�Q��0���lv�	Sr��U'�?�; j�ߦ���R�Z�~��p��eӸo�vƆ�H��L�����W\�gm�!aɝ!T#9>z�t�%��7��)F�S��UVӱ�J�Y�/��;H�'�U�o��c�B����1���C�f*m��k�4��E��^ ��;c 0�z_n�^�\�|��^ڇc;h�ƹl,zc�0�|�ܩ~�6E)t1P�����W	(6�4-YA�H��ze/��>�doR�6�ȼ�
O��SQ�|�IF�j^r�슴��Lih*��B!��L�= V���W�82H~�o��YU�)Z�~91\��VV��%�VɈ���jxa����ڢ��ed�.E2}�b��TF//E��=e��:~�%8!G���j�v�1�A��Uj��0pٗK���y���&S�7��s��e�H�������;c��E��ۨ��U}��Ȇ�.Y�S�����u��aZ�5�آ3��q���` P�������
�-�P��JJ������P)�쏯�,����	N艱�7�]�I�W���.����OF��V�c�(��l��N�!�*������۱E"-�a�yҺӎZ���TZ�l�6wG-O��/!�r���e힓g/[�����cfN�ydi�H��A(�@_�Q��؛�|[T��	��n�F�(쎇)��Ťw��H������P�����Z�v��l��ر��u6����ػd��9*\��
�G�9
FE���b�E���G_5�R�ܹܾ�u͹%�������̰o�+�>���5/T-�Tg��p*b�jyR�nq��O�Y4K��F��xU��;�8�9��	�& tK�&?�B�v����})a���hu�U �L'l�{\}��U���{��U�fiB�ƅt���Hl��ƣ9s!��`�����^_<xCi YM�B7�p�Ҡn�d:z˨��&�-�n�jT���c͕?n0c�%�����*��6�Ӷl>R762�����3���7v��[~L6?�*��)j���|�mnm�`�ax�z~X����]��f �c�r.����qv���v���5��%\)
�a��6�z��%}�WS?2q)��*��NA>���pS��d�T&Q��u��nO��QƊr�덮ѿ�|ԁ��"��dӗ<|�
�����}��^�?��TF{ ��q����A�+S�u��]�Tć�p{���v�`V�o��%G��b76��[�3R�s�}�dp��!H<����~�NrK��@�V�2W�Wfh��^VX�)nҋ;ڛ��[���}U �GX$�Kw�ei��� Θ~�Ծ����Gkr�L:�Y$�-�J�L��>>��śEjV�����Ȃ�k�D
���#�BH �,�a�[�EuaԨ��a~unt'*��w�..�sd�Ə��&�t�*�.�>Ȓ�R��n�.2kё]>��ɚ���K�a��wu%�̒u�ϸV