��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{�H|��6	x��:Rg�Jl��?�ʖ~f&�n�e��*�[.b�H�����;�FM�K�+�/Ȉ���Ҽ���}�.����~�|`�����Y~&�C eC_��N7�gAk�Fhe�v��\��Rr���7��t�������A��6��_�h%%:���e�ĹW�sQ�˱X����̅��1��#��ވ.�U@7��L{��j�q��C'D�gF�MԀ��Ur"k�(�m\I���~ݎ\�j������P�P�J����3ފ�D2Dƈ�����x�<�z�\�c�ĩ�E�:��t��ᝨ��H��Bh\U�XF���p����+�m����~%��+G90� ,����E����c�7��NӀ�AǫN�s�<�l��(�U
��s��@<�=��7��s�z�?��j�`��)ʻ\ ɮF)t޸(�.a`��jF��E.���tl%��=����"
�9�`-n	���TI�@�B�nL��]R8Ko���f�#���EP-4�����MpS}%���v{���k�>�T��Kk��,~�}��?LӀӜb�Է ��=ffc4>5��%0ӊ+�HR�\�\�ĸ��0A��ЖrY�\�"H&�r.|6"3h�I_�W-�/1��QY�8TPy3<N5ѫ�[���FW�'�3�~���딨ZH�D��2�іٖz��W��s��AO�6fa:�V�c��Ќ��#��lp��U& �*�Q^�!��,X�c@�+��M'�{�����:MB:���L~x���
n�0�C����1��3ё�u�4��q맂�-�q����k��JL�I��-UAf�ވsX�#���6�������Zv���q��Őr]9�_�/B�^�	G�n�],�-
Q�G"$Z���h��7J�d���Ւ�rK3�a��)]S��E{������^����[����݌�cSܸ�R:��F�>9��C�lZ�n���� 9�?S@�6f��J�i�=~���nZ4+�|!k�����f��mk���#h����<����v� x��~w���\i-��.��vG�+݊j����%/²a|�"B΀6(�=J�P��� N��l�ܔ� h�*��ň�P��Hw�0�$��V�7����+�&��-0vڮ0m����j�!�ZFv���L�En�!�w�lz�@۞�X��ׁqW��T�O�9v����$��N��U)X�[����֗��Ç� !�V�.�m� I�>�$���h|:D�b�N��$.�<d3��S^�W��_�YO�aҵ�׊-��;�i���æ�N�- 
�51�>A�r�~�JܧQr"�]s�H���&���vo�a����ե#�ZY'.�B㉮�/��h;��rE�<%P�6�aFѲ��m)  ������2R�h�O3τol9g�L��p�#���(@6�sN��g@��?�V!�#�"�'���_�S�l���,��ʾW������AR���M���MN�7p?�5��w�A�*�KNEL����C���> ��'���N�����*C��S!�P�s]|�H���(��������%�D��� Lf���"���!Rtzb���t�����x/�Q�����X5T�O��	���z�s�[�+����@����?����J�&��@/o(h�����V[��r�ޜ�Y������A+h�H�gH��5��#�����kTʳ@g�IG���w��]X�s��r@�+��抸���/‴� Lc�m��k尢�I�loΪ/_�	�t3/�jo�i�f�ƴ6�?��%*�+���RnR�qQ<�	LW�{Q`ަ�3)�	{�<���͘ 0�ޒ!�Ǣ<)'f
�`�"7h��"�F��1��4$��Ր��	�G,�ؚ/Na�5;a�h���5���n�b��� ����x`h|��H�R[�Ӏ	�6�:{��;(�x�乑Hn�NjH�|�\V,\�c�Ɖ(������)~R$a�Y���$�����J���9�R��~���?�S^��)&�f\t�h�t�.����p��������(u���j�&H�b:ݱժ��N�&_�q��	�@9�W��usm���8``㌘ۉQ,7오Q�M㔄��R���y=���> 9�#�Dv�ulk-��K�́y��WO'���?���0n_e
��4�S(lO\2