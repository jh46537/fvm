��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�;��I�0�y���Q�&H���I�q�TlA�<�ЗJd���� �P����@��	�d�?��ҧ�iw�MԼ�k���A	Dsd�M��T�wY���׏�1�M���H�e��-�BZD�V���ȫ(_㨟���"��M\5��"�J�g�<X.,mc:�'�A������:_�+�**Ẕ.Q�~�c�0aTdF�qME��t��7��x��V�?�`$�U��'"𩔠��������q�����H��\>Cɦ�C�x���5�g��#�[�PFL�3O����֝fc�;�t�í��ρ]Wo�sU2i�*~�)h����v�b�tTOJ��.�%Pp�5�T���i]!��I��<�>.k�u�2v�����L՜�e�+��iܾ�0�������B�d���̓MwD�D�L�;0�"V��GV�f�/ni/E��7�|P}�zbY2L�(�U�Q@�*��*}�A�z���k����I����W�S共T�4��FLd�uMU���OcӇj͍�H��h�B�^(u�G�����}�YTU��C��E������K�G(�I>ڬ���]�8uG��Gꓽ�ߤ �"w������Y��̶�zYs���ƀ!��c�BR'�����U�xD;J�����y���`>�n�����3܇be,t�,�&ZԺ5@yDjF8�I�N���޳V���}RNx���aKx�א�ol'��J����w�9 ����.s�ǿϒk����~Py�r��&!3��"��yxjw�N51<���-�%��̅��6k�o=�B�Y�"��I6�3צo��S��3�Vb"�g���b�/��Gxw��>��v���@��ƻ��$ J̐4�Zo��ɭ���c�#�{yՑ1ў�b=�*�:d�RCd\�|��9@x�$ڽ|F�i��~���=�����u`l4�r���^a�NUG�ߑ�ۦ���{�\}Jc��~��L�ң��E�+<5�|��n�Gƶ���DJD�")��?�AR���8
�
IY	��l��P`j��$NM��&�W�z��VKūqr�ٕ] ��_8z}Ă�<G.�2q���l������ً�O�6~�	0�}p\��"(������+8��M��Z'�'�|���+h<��{�ZC�{�0�`x�<
�0X{�T@�*E��H^g�IJ�	o�^dT�p�窌=�&u�/ǳ��jx��b�FݰTB�i�G���p�KW�؇��	�^� ��M��r-�y0be���w����W�uo�m(Qwq�&|3�Y��C��N��Ѕ�P��LX�������G�C�D>���vG��pY][���CGl`'^>�/@ܹ��
<U2�s9C�S݁���sr���D�� ��t)^�ch�Y�g�r:u��!��Ox�pA4�)V_$�+|,��H�����q�7M�Q��\�o�+{/�*���DK�C3������ބ���Wa���W��ͨ�D�ry��Qa�|5�Y*4�S�18�ȃ���3גY��Fy����Z�h���u�������'K�Rc��.��[����/�J��L^7���E:�*�����O�VM�th�B�D~a�+1��W�������e��c�VH.U;�81
F�
GR�D��l�
���Zu��?�OH��͔1�kG#�vK�noˈHq��#8�ņN����BӠʇC���.�� �N��{��	4��Ԛ���_�$�X�F���R�����B��&�:9"D,<�T#��~��D��a�f��*Sۋ�Ƒ��	q�T�?��E/ؔ�[$�" ���.�r�#��ct��ƚLdZs֜�$r������A���Dqy��"��"�&E�
vyGZ5E�vE�}���g�z�?9ـ5�꼤������H�\�DO�0���5�]r�������_t@̽���e�B�ej�5�4H^����`�m'��~�E�ٻ�85lբ�o�$Wq�`�T�Hg�{�֋#�t���M�_)ŤMỤ-�CҿdJ���ޤ9*MovCZ�_���_�Z�qP���x��������1��q�}�e�ǻ��c#|楑�ўո+&Ǧ����>��p�&~�W�	��O���g��DĝU.�3�w��\�[���ž��"���`-�':=a��w�Ű��E�K!����=�/w��������v�c�����W�N�� ��=����t�i(��'ސl؄O3ѩkB�0^����6SB�-Tg�R�����Ȍ#�	YY�^�A��X|b��8�3�â���Sm@nF�5u�<9�x��bb�d��an��|oe��7�͊��Ψƌ
�$I�w��E�wU���2�s����ѥahI3��+�ط�N�Q����r�� $kn��ǂ�c!�!���Y�Ļ�L�ӽp��L��1�5H]���������Cxq���B7H�w�8;�CoC�	���@)�l0�z؏!�u6��ۻ9���3�@��l�Ƕ>��U`�K�/Ar��.�M32�ݬޱ��'mCsܮ9ۉ�і�#��P3�u�����&(,g@dj7w�g�: �?>�~*t+1���!;zy�>�?��Y�:���n\k��wq�e�Z.G��I��ҘL�M�tqo��c�y� O�j�(��rB��!z��-��[���`,�=�bW��#U�س�{Ӟ��F�[�V��)l��{�x��P�Uw��� ����2a8:�7+jѭ�_Y��N,Iu���;��>.�L|a%n��,�)�4��-����_�@V�f�ipV5.H8��ete��x�I8�%3m
����:���a�%�7�'FDW{fp*_������z^0�(*4^
�4��3���w�Ӧ��r=�he�V#�ӭW�:��t!��c���$7���7�J/<ϓ�Ψ�#�F!T���-�cr�����+Sj��B��D&�SR��#¶�B��a��&q��YF}B�����bIJ���֒N���ȽW�̢9V@]h�����(DЭ��S��c��
�La��8�6�� C�G�����B�χ��'�.PN�cж'�T���w�4��6�k�N̦�'�%��]��KnM�l�o4�Ědjwʘ���ɻ2	��X���� ���2���ɦ��^�8��� �{����FJ �fj�:+b�㠨�$�Q-D���zK�=��C�CF���.�iv���m�DKJ.�o��0t�١�I�:��-]D�ȰC�m�����N=��׽^G#u��v#�B kj(�*s�.'����L��n��%�Qab�N�3I�NJ*����!�\W�J�
`X�wvA�b �Lo�����:9C_�� �锅��#?�h��}kW�h�}7KF�:�Mv��wJj��b�8��	��M���Ca�
�[�+P��3�1�Bb{B]g�v&���!�6\qA��}%n�sfX쿸
՛g��"q'Z7ՌD�=���H�ɼ2�ѱ̫?d�G�s��i^8�3"W&VS�f0�S2�(�% Rp�O�]	�ľ����6�)���M�+3U�N�ie�]J\��� 
z�cF�{�q5E�r��m��@���gt�����b�qo�$T�O�MT5���2�-��"�3���}�V��B�6�S�q�'�ĴT���݆&$�c��t��o2-v�^������T�[���U	db�r�)�!/�#h�l�N����Sp|Q�	����&�Vnu��Һ�D!#z���젾���L�@_ ��5�*�Ee��}H�%�^��Sq����֓ư�>���-��e�[��@��	�+Õ,�80�A����k�Ἃ���~2��[��qx�*+gj'"w��V�&�"�!Ct���D�;�� 7x��i]�AAF}�ɴ�c�!���&N�0F��طIr83�3�����@�_�4�Qi�7`{��X� ˻g�(�4(K�Q�SMjg�3A�_��&��*U�i��v��������D�9F����������2�|`�<bA8�_���r�Dȴ灔dn��^�#@0/��m��]q����d�<����@�L�����"z���v�!�)cuE�ü��Ӯ6��! a����q�``�0�A�U�o��"�����f�E�4�4c���th�k�ߠ��fr��u��c�ܐt7�BV+� E����Cqj����`��ơ3C�|��l��33@骻��E�i��[1����gZ��]��qq�I�����3�_~�G: �0�:��\���?
���$�Z{����l��H���j��Cn� ��D�҈��Y�/�8�y�a��1�<8���GA��\��΍������(O6_�d}6q>g�}+!\YgP�:���t�n��9o��-��!�uʞ
�]bJ���zx<����uaKõZs[j���c�g ��������L_�w&�n�ͽk���cU�>�ݞ��tQ��|�i_���X|��ܝ���Q0���(y���_Q�[�[���I��%]y���O����ߒDmEUտ�鐸�K��+���D�B����)� ^?��e$�}]"�ܠ��>9 L8�<Un1��/66��s���g�޵�P��N��
R�A�er֍8j� v ;�i�e���;�I��γ%h#$ ���J���ʼB(`	UR�狴6[p��S��s��)6�d��DgN��,{��~"5�}�\C���RkqǄ�S�����c�^V���C�}��|��3���Y�h]�,��4}e?hЍL�<�ʑ;��K�]����vpQ�>(Q�h*|�+���^æ��
�����I����I>9`���ȟ>,t8����������:u�Np�^�L�)Bâ"5��X��ô؟},(�Z甂ћGS ����t�|�Y�ʚK
�+�(
���;�[q�PU��.]�@Pq����sS�6�M~.��������7ܰm�7�F _=J=���!L�r��\+��n�&��P S�޸b���%�f�ق%j�p��tH��G�b>�S5�	P�@61
��I7=bq�9�k�:�3��{#�&��,��)i;E���>%ZK�fҮ���7����[[vKi�������� ��S?�b�2��W`7P��;�����B� !0NJ�_�(�>�����O������w;�j�!�_���=��rٖmz_1#�;b��E��i�G�5���ނ[���% � �e6lk���@���/�c�پB+��_ˈG� ��\�-zJ1x��_Y�\I\Y�z�̶g�]Fˉb6[ѥ(P/s�r*�ߚ�M�j-1=x���m�zި���t�e��Rt��^E0ܬ���t��ה��G�#����}����e�#��<���^�=���~_{9�.�F�Ɨ-!���xC|��S�.ILx"-(��gnµd_.3���7f{V�-_�_gJ�]�O���)�I����sn`�_��H䧚�1䲷k�j�����JX�֌���ys�]�aۋg��S�ɤ�BIu�1���>�j�H>V��l_v�(#�zI��"ӄ����SX��k)��A���Y�@�Nr��z�q�٣ZNݚ{s�>��W��c&ʡ����k	�j�߅W:y��uf�<�7x?◵N�h��J��?�>���;wrμ���P����h���=}s
�GE1�1����A
M�[��b������_�ݮ4$��Iu�1�IS&������Ot���_�&�)�X椷�Lj�6K���ޛx��J7�;+�<�Ug�O�'�Ű�>��$���9�Zز�a�?�d�п�k�Q�n||�N�׷��'f�-!^ǝ��'�i�Oa��T��8CcIBw�O���Sn?a���Q����V�!!%��_�J��YJ��M��^e�e^���v�V����ĝ^���*ݯqEy��OTG@8��y1+p>/7B�����H�M��hM�-f�P���K����ݵ�"�Hg}��ΰ�w�aw7?Q��4J-+W1rjsՊ�`�+�*�L���?Qh��(~�C]��h+���VD�,[�Lrf`��(�忡fu5/���,�/x�|��ؒ�1����=`'��zP��Gǧ�|��P�z�9��O���,00n;vyA�	Z+b���Jf���sT�P�d��ʽ�(>/*��Є�fe��>p1+�m�;��b��1Bv���쏓M��"Ep���ea�ti2�o3�c�#|��F
���j����B�~Q) L�Q��&B�s���%���Ui�{O�OF���sc~>>i&,��F!P�u�����c�K���d:���@�|��9�84er��!������_��u�3�,�6s�٨���?��?;.y�x��(���<�<�Tx�	w��۔8�����ӊ'X#��6���&��,p�sh��ΓF9���	��q@{Ih�'�S3e�\�X��3���}<��&	��xn�u��K��Y��O�T���h�d;VG���I�a��>�3\'�|��M�fH��"��Bs�_�<����:�۪m-с;Io�JC�e��