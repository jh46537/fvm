��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k{de���ӱ���!B��ρ��cb��c�>RW�V��*qn�����.�e�i��m�pm�G/�Ѓ����X'�w��6���Û"̧�/Z`G�2�p� ��0��C��"�	,�TƑ?ɂ�1�����
!������Z�}�or�[J3z��@^��G�.��_"��FӥN䝮�ib��eiK��9Sm���*��v��6�
hM\α
͇;�p�&���cJ�<'���P����2���kj0����#J���8k���-��2KU�?Aƙ,I�nL*p�$�ઁL�
�U��bZ�ɩ��pXl)ƹ��H�����̤�ػk�yL��p�pP�xWu�N2�?�f�Ҿ�ˎ�-��&{��?н�.]��δ[i�-a�*S�P�S�����,]�*s�(X�2T%��Н$zx^���uq=��*k��&�ݪ���*Q�����^p���k҇Y�����枀ъ��D��[/��es��1b��Qa��=/	�>u�T�7=�=���P#�}��Mج�$���2�T���;5�����S��	Y��v
�0v~M6���c�d��hQë�uGCv����'��~�>[%�w� ~�{Ѡ9v�2�'TJ��-��@���E ��c���W
ϢǦI?�
�l���[����m[��tu�������"p����M��+��s����}�{��D��|tV�uv�a�|T.��� �4	_K�5=m��
��i�:�y�s����fS�[7c:�=�z���9�/��p�r$�)�4v��3p����#t{!F��Z�H*�`n���*�ð�uKY��� �{i���]w�h�m�K��P����^��x����ղ[����$q��Z��������h�h��kO롟r1���wӡ���^49����5�1W��r`CS�0X&%�Dwk�D�l|<3ط���ZK�YGety�U�Ԣa�o"������	UUڤ��;%�@y�dT�Xw8��E�+���pVUy
V |.�5�l�cS>O��1�B�M�Kx���վ��������!7]OK@�'a��7.��I�'O��7�
������TASA|E��#��+$�*�R�Q)E���0o�Y���h!8�g��bO�@��h��o�h���l�·Y��t�Ջ/�&F�����0�灠�p��Gd���X��O��R tH��MdL�}���v��{�O͆;^Z�� �5��g-�XUZ��Fh�yX�c%��; �T�95���7���{H`�J����4^�>`�-��~H+��Ƀ�Ѩ�(���?��m0�~h�VX��lw2T"�+ƺ�Bx0▝�>�q���n��P/u����ݖs�B�D
�M�e��QN��f�#�m�"b�w9Oˆ&z�Pg�V^&A:_�$���C��!W�p)�����pI��Ҧ��z���`	i �zކ�TL�Y��i������p|on;��S�m-����[.Q�/���g����UW)�:<��t䒆+	*���f�r�[M���ҌCA���;vmM�t)8��&�W�xxZ�������� ��{``���4���!��w��0��06Y��M�Gl�=��dZC���6Yd���I::���g�"Sz�Q5�d��1�oZ�$I��8��i1)-�J�d���$��꟧vTp����DB"��޸ҥ4̞�:yͳ穏S����Ш�d�:�����]�gj�t����U�������FB���9�N������쀟\zz$���CLH�����%�A"��=�w9B�g�o��=x�+>�@��z��Q" �6�ä-n[�C�ch~��fn;�?����N�F�(�5���,��o�{����c�a�x��%��@�����W��~�RL񙕾�h8LĚ0`���4 #}��t�*����y%�hq��:���]�w)�n&V)�=x �j��k�p�Ǚ�*��i�Mp�b5�`����M��^�����n�X:GtByBuEn�t�Ȓr��i���R1%�n��?'�QΣo*�R�"������D�ؠ(�(����)}���jrc'3Ў�qs�wxX]8?�����Ζ���&���v�Dn��Z�]\{�#�ib?�r�����IO���唏x�%mfE���)�n!6�
����}�L8�P� �w*�S�z�u��ԏb�����w�S����Nv��L2l�H:�~J0�0��ʽ㽞b�T�b�NZj���v"׸���p <붠2�;!Hdأ@R6Ř�|$�d����v⯐c�?"��w��|���M'+_Ep��������i��Xꐹ����'s�L?7�-���U����s)���� }��9=�aS0[��ұU�`1.��?��+n-�XɄtf�F�$��� GW$�)/,hÂs�������)��LDef+����Z�N�En�ٹu�\��d�.�VZ���Z2���s5XeMjzG�iM��6��u#m����c�t|����z��Qy���]�o�[�����[/)�9oG�E|�h���n��im����/z��¿Y�v�癧�Q~�]���Ј�q4�?��=2��-���Y�}��%Ar�E�D7������?��qB$F}��+3Պ�,U1�>��ģ���;˵{Ɓ;n�$R∞8Q^�3��O~:�f%�3��5�ih{��.L�m�N�Sh�����<%���X�M���\ؚ�R>�%*E��^|m�8�d �y�g�Vj�b��{�1
����u=l蜟i�u>5��zՀ�B�5b_�B��g�8���'�i�����kypX���d�EQHy��Ɇ��c}ts�/�*�/\39g��ٿ�������8|Iq5b���a��<6�H�1'�#�
�Z�gk�wZqmY���7�=s�����le���iH��x�{ɚF��a�Y��9P�<g���f�;����r�۸2���$�ט`wE��@/�EC<�8��]��J���RP-
�`���{��1B�	���_��&_�x)�X����LX�=OՎ��^eL�v�cOfۣ��j�E&$j���-���A���E���N����/��a��t�����=������q��Jn����y�MT�[ih�a0F�} �{�G���ͣ�Kf��6��T[Ty55펺tiP�F���&5����Jަ�7�y�(��v_��n!��QZ�r��ΏHte��g#�N �c/����7��H^��@W0�Z(p2D������O��OF��,`MR�,%c�ns�L�:G��Od�+������A��I6@K��7��8�A[��Cg���{�*����Ro���^��R�0�.��,Ͱ��7�q��\m�d����5V�tr!}[̤����m���L�k_Qg?�ct�`���A�tҏ�	�t!g����������qN
lc=|)�KͬL*�f�����b5G��V҈����K)[��I���0�,O"#F.5�F�:��A
$���S}�x<��t]���¥b��K��{:��=�a/��}a'��Gp���:��oH,�Ǧj�7#on�-`;0�������1b<ro�Jx�j�mV47��"�C�/)�=��i��(����$1��\؎2�ŕ\�;6�M�F����"�:\��5F ۱��9�F�%�����tT)���?��.F�U��z �G-�� ��L|��։��3]zO�j���Sc�mrB6�17�ZT#d�]*���|5P��nj��bve3�=���Gs��ﭴ�>�F�=b�,��f��M�'�mWո4?/C�z����S�`��/�1��K`� qG�۟'.;�<@��@��>u�T����t@/8��E�52g�I���U�?�B�ZZP�vD6�Pd+���F�Ս�{�y��������U�,Gqf��h���Q �����f��!tӇ\2Rj-mZI��Χ �Xdqe��Ȓ�v�]��ΥR��J��yy�i�41_^|�U�W�+�tǗ�Z��M	�M9�Y��݇�5�s;�x��R|�����i!�����a�����l�@U�e�:�$�f�B�:������B~g�d>����W�����Ž9����6���"k����e0	�\�`�[d�5Fm�J˲;Q֬���W�V�&�x�b	��>�X-q��|㬧����f��B�(䖣��ܦ>AІ8�fa���(F@!�R��EH^MܕuCӾ��
>\���y���TR/�@��RsS�<�U� ��#����=���'�2ҷ�T�J9-ײ��d��3$�Ć��q�2SgP�s�&�k*����`��'Z�,l�[f��ۛ	&���/�P�����ʄA|#��jًc��S(:�,��*��T�y�:�����~�<����z"!�V��?�G'\�y��mӻg�};�lÐ̺��F����s���X8�9�k06��gR&�VE�V�����5�<�%�,"���M��s;��>���%�^6����r������*�=��[�I\AI���,o��μ�����#��Z���u^(W����e�p���z��)�心���B��0�>M<w��8v��wf]Ӛe+Δi����cM�.��Ɗ)���AIx5:`�t��94�1(T���ta[Ia�8 �M����1P��p�kt[��s#��MdK_�/��/���t���O�{T��Q�ӳ_���R�*�BC$�Ϻo(1&���ǲ$T�ָ<��j!Y