��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0����>�P@�:����j���dV�[J�e�˪���ؾ� ixc3�xz�S����}��������1��e_���O[�7��]����ؖ�m����dk[_+ �s��G�hq]oH'G-jP���yo!��@�w���h�n	y�O����?j����\m%!�O�W���iXƿ���-�S�]�:p��3�f��ղd�0N+5�愶N�	�8����a�Y�PS�t�1�[I��n��/uSg$o�%�眩��t���i�R5&��2����f�?�vA(Sv�AH�qB� W��FD]|��ő|����]�}(��N��hR�����=���G�E��N/��^-����
QSz%��s�Ҝ773b"�3
5�ˍ+=��U�'�`1��.!hu���v��%���T�؊�E���N���n��}���!SU	�~=���c�U#�T� ��"��触A`o�9OvV<���ș�Chu�|���A�b���,f|&0N�됪��I0M�~�Fh��"�C�<�h�
00�,�8(�����	j�t|b� �p!��]l��?�b�i����!��~�5Ur�٤�m�XF��렯�<v|g:A`O��T˵z�#�$ъ	'X�lu`կ.0s���6H�`�V~����"sT�H�<j�#Sx��{ǜ�����3�=�`��0X].� ��P^�B|�yO�t;ߡxg�!D��F���_�bp�!�P�A��ɪ��hhT:+ٙ�cr��3a�R{�8�]L��~{3�?���{4u/ƪ!��
A���~�1�����Hg���WH�)��[D�7�$a�s	����[v�1T=-�X��4��r7���/1�^��T�i�᫂�Y	A�u�g�"��]u��t<�'��� ���7O
�J��y�)�Ø��Y�������/��dieʾ�d�nNq�`��{���s���?��Kzr��S`�E��-'5��cF؈�3�3���:8V{��A`�t��� ��N��Gab�&�	��Jj$�D��BM�[��f��7�V�tL�����u�/����Y*W ?�;��|G�Ouda�
�f����Qv��-��F���y�.���:�%�p�3Mys�>Y�|Tz��]ԯ$dL��x`��y�C�{*��Y5��_��+;J�Ҿ��$n�`{�4�s��%j��g����]Gɔ��\��e�X��F���5��]���m�Cy�Ca�~�%B]��B��b96c3zP()է��!B� �"�-u�lk���E��I겠�����Ht"OXA��U�mJ#U�*7&c�����ޞ��(���_TM��:��Z.`�?"ǯ�����[���8��T�itu�~�A"2�/�՗*EI��-Hmɶ���9>tޑ��'�8��u��wʱUFx���ϙ2X����1=j�x��C���n$o� �9���y���Tؼ�E��(�b�D0��b��_xt<��i'�ڨt�{P��#pz	3�%�Ӭ���w�VS/�wo�����=�z�m�Gy�;[��43��- �F�:�ǻ�!��	�i�v9��su_�����(oI �G�:5!���{\��]"���哩q�7��5>��	� Ȥݚ��/�x�$@�l�|$7�d��/����y�`叓��Q_��uI#\L~`�g[��L��<Ѯ?xKAS���W�Ɍ�c��H���'��P(S��սz���V[�� ���=�
as!�*�z%��(�kOd�7lbh�7e"d%mr���s��?j=��$�x����|��)OE�j��O(:����x�Qxf`���J�5��EsIՀ��������y2��Qd�̷j���#Z@��*�+�NXbE{c��4osD'&�B"��r��9����\3�G���̼��Nkk�#��R���=X��i�#nf+}�y^J���w������DD~V���Ā05��<��>��A�je���-��� .
���rI�ٴ����̬���ʜ&�W��H$�4~[z����>��?/2��q��YX�cgw�gQp��'>z�1$(U��J�M@��̵P��&%�~�q�9�_^Y�|W4?]��R]��[m��8"K��Mѧ�Q�I'y�6��8ZP�2�,�e��̗��BP<�+����PJ1��j�'���3���e]3��}������1?m��^s�9�����~��TM#�5?��a�K�Mt��Q�Ky7��8ٶ�\�"@!���O'�qv�f���'uji��z�p��}�<��}��0̇չ�0����jit$���L��j�"�g�J�V۱!�84.�
E
��7����Iy�$��#��<z�~N"���?<3�b�h�t��'�j4�%$��=g�zH/s�q���ak ��wr�Qń���lc�>��O܇�������q��8��Y=Z0 Ѻ���
� �K�f5Ʉ�7L	�4g�vsX��C�0S;�?��Qy@���w�Ŷ>�g��=}�2-�\���Am&��k2q�g5d)�x�@wo�n��TW �>���E�_��dS�
�M��h�t��4��Fp������h��Ǚ���s=�l�1:�9�K}�y'&!O|s_~�x��)��`� ��q����qg�m��Q��̶@ci�\�ynV=���_��j��{z�E��/���[ỖO�bw����+����H� wH�9H4FR��Z�K�ۑ�㍠YӃ,5R+$�P�yϗ�2#}UD[�� t(]@���wW.�s� {}<`����?���2�]����`�M�%�:1�-np��ֳ�֩큃��=�ߑ��F m}4i�3B��	<��h���i>�T�@{��	���/�����&
�]��!L�kJ\"djn���[ r�8��)R�x0�WQ�9?K��c{T0G�S�Q��gZ�F��T[�j,^�33�X�8�NQA��)�Ǜ��2��S'LV!�!V�y�fA#����7�ʩ���@aVݒ���N���e�S�"^���Հ	l��C�ˍ>)ݏ�?��~Ϙ/�S��M�h!m�iPPL�z 6�.
L:�5�C6-f.�u�������L�1{Fjo+�UAŚZ�E���o}t��;�F� ��p
�H��\����f3����	��K�S��sXD�:98��*��VD,&�N^�R�{�K��}�\�ol�3��q�ǝ�΂[�����q@`k9NAg� ��,�o���2A��ɬy�.f�/N�q	x���?p\B��+f��:H�x������UAt�w�Ty���J	>�n@��vs��>�
�xǼ��0�2c�ּv��:�Ì�