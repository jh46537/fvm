��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�Gf�`x��*�=��	��,���9Rk����F��g�BGu���v6u���I=�  ���B0��+�I�G�F0�9���O��:�S.��h,A�.���}��&W��3^�m����:V��Ϊ'
�o�����"��X0���
��G�>ڈYh6$9��b3e����C��sT�ì�y?��}�D<;[TF�Cx��:Vp(\-X���,!.����5�G�^-JP�,�>J��ʘE ����x��\��'�X�Z��f_1��QE�Wk~�>&�.�������� ��kŬ�/Z��č�=��c�o�.��@[��1pR�!���:�畮�uS���΅�o3���>ǹ��oW�/S�Űxv���0/@��y��|vk���H�Y?xp鑔�9���BN�$��9�Ť`�&��3My9P�=y�7�&&$��`0Fمl
�_�7���w4@�piB:��E�(OqU=L=gLo�#��à��	�Kn�nM{^�8���(R�c�A�F��u҈1ZJ�������YWQ�#X�����߉�>�Mv-��(��������+�� �8�7#*e�P���5���威Åk�*����`b4d�����ȶ���������Ba��:BeuM�x�@4}��K5	������q���ŷ��A�"�� �Vfs����TxA7�8_JH�M�����oA���I�ZN�f��)����t��0A�L5�{�K���VB\��Q��+hؗ§��O��.]�ѵ���ľga6�8*̮4S��[�
G������-VV�F�XP�R~�sP8��J�D�=XBM�	����۷<5]u�r"�������1;�B�@��*`�s��¡l��
�{9@ɞ�����^}�ݻ�k�1"Yk�+zuq����!Rsi�W�ݖ1g�W#���1�O�藕��%�~��v�����i��	9
��5������2~m������1�3e��x')�/��{�iB�m�\'��%*+��-���!��2�ݍu%3�u\�Xi.mO��5a���K������t�0���D�[H �����d���4����A����2�}��<�]jA7l)u˟����t��
hs�%�t�}�C�u-���>��~R���{%���D�7��6ɆD�����߾��h��Qu'/ vqK�)���E-md��$/�ڼ?��p���G�@�^��IZM�\�ʝ_����.����|R9?<[�UP��z�w.���TCh�p��voI$Pc�(�P�?rX�<��Nk���~�Ki���^_�U?#gµ�c`qHZU�
Qu�ڊ�Kܲ�[h�'ůJ?,L����4�
�\��ZT������(��J��| ��h�����/��'�$�E=ʒ�:�P��IY�Щ�H{�!�����R��7�+�Ti��Ċoʉws�px!]�Jo�)H�����}8�H$7�i�u�6�m���1[�tt��q�7l��p){�a�T�d�]*�΄~o��L7�Cb��J��seE���?6M��R��sJ�.�K6J��p`>�诼6���X��H����Q�����@�v;ؐ��L�J������fv�B���,SQ��jꥬC��q.Ʊ`3��9t��h�!``����G��n���84���n��a�z��o�#��6��m��;I[=����K�[� ��u� ������C��OxC}�E}����>6�UOr���>6�aQ`�j#!!��@�K�ӗ�V��C�L��i�u��rF�3 c,��q.<K:�t����Ra�vz-��I��&n+�ע�ܸ.���w�U��i�R�X�(T�Fb@E��,��{��HQ���"4mbD�z�K�3�ʫ�r�f�s�M��]�'�UɆC���l,F�2<�L^��@/1�����q��h���ڄ	#�$�6I��t�E�އ�� Q����=Yǰ��I��uq�GĆ������S�C�{��5�.ɘ^'tyyURJ�Eo����y.�Jb:���|߆_�������Uu]�q���V�L&�aCZG�T,�Fļ�ご$��YU&wn�-hҬF2� �z��uU���쓨�-6:�����V�����Tvb���R�H�L@Fy�Zf�[��G�&�XD��c��GJ��a�����4�k>� ے�'�`G�qS�kM�i+I�� R�Y��.��Z����zTW4D���:/�_����{�MnK�w����/���쭮�r*�^I���ފ���m �њ�d���L�1�9e��젿=(��lx�"���������a���mp�.v<�|�c�zLE5� ڔ�"�@��9��>{�y�DbW���/�ls'��2`��i��m�fc��r|��/��W�G�}�k�><�񲤵M�Ò~��;37�����ש�[�)QUvT��é��.�n�u���y#l�t~��'�*���DZ�$l\��:j?��u�����8Q}�6ޡI��8=� ���w@����c�3��W��_�.
�h@���ŋ��y�D%�@��!����ou �zaQP�ӵoU� Π�C9*���58�n�[>KN�I��z���0vm,ʥ������=x̤�d�hB+m/�NH�+�)55J:L]���S�ѫS3q@ ��h�F�W&��F�"lo��E7�h�V1#-��<���A�s�H�L�+������ʝ���<����)B������@B� � �tA{\RYv��.?7�t9�x������\�`]7�\��޴쬠[!�6��3��E=� ����f�R���7D}�Vx�E�,�n*�'�}U��J��G��L��p=���#���Snj���y�H^��5���,�I�ُ\:���
�{��̽$��/t�v���7�\ܧ`30�i&��������-�"�E�G�i� �u�C����s���(h��5W��åX�����~ԴFW{�f�ۖ:ܞ�9�������5��1��d�҅� #J���Q
F�t����_��i{�����;�!�p�v�eL� ���{�f�C'ֿ:�c�@�]�� }Hj��i��qL��ͬ���_-��6V�U���b�o��Ik=1���������9� ���[? 罰�S3%{��w��\��[��۝-ɳ��"���=�#b Q^v���d�����'��:$�!L������헹�����l�M��+�k�5ʯ�?!�"6��lLEhz&R�S�d�e=o���Fl�'��uE���������F�59Q;N��ӳb��3�TlB2����tH�.�����]I������C�����0�Jx���34>�R_�����F��L[l? ��W>0)�>�U�r(�����Q��sw��J0�G+%d.�_d���b�P'�N��=O�P���92�ꩄ?�Rq!�Z�]j3��CB6��E ���DT
�[qP�	l�@�)��pwO���FGE(t��G��y1Yp>T�2����E���d�������/��֍��B��� �bf�S���26
_TA���f�-V��c7 �����k�ˊ��uו���bf\�ñbO9zU֙��,.��,,P_����u�v��n崂�+�Y�����kDÏ&�i������^h�݇j�����X��d�/��>ݲ��p?K��Az�i�Vh �� �����6���l�b6t6e"E�ii���/lK����8v��{M��j��v�ÂB���<�/�w>ka�_RJ�|��e�#)�eI����x�|�<��%�i(W�P�Y�eh %��눕�KC^l�PP�S%�`��pM)F4l�������fM����`���{�&m!f6�gg�K{֘��w��|���Ӯ�^�1i>�U~�}���2�{?b���3��i�!�Eo�ߒ�*�(��1��u%�S?�=+T���F�ZS˕7��`���A���lR�~�C���y4VqZ���w��ۄ/���l�_$ȓD��Ytl~���y������{��U���v¡�笅�T��k�ǌ�!^)a�cC��O���R�����pK�3D��^��cn ,�S�|�������>Lf^���4	�k0	`�3���� W�U�V��p�I�G�Z�Ru�B^�
�Y�Q���{�{AM�qYe�f,�|��ߜO.������7&ܿD7[�� ��"xI*~b�ʭ�GM����,�'�$�[z���PQ̒eT����18���X����e��fj?kA����J��/�œ��Y�a�k[Қ%J�%��,��q�r�lo��k�*����2S����L�e�ty�}90�*y倏���o-�e�U����e�]I=�j �4^�W��.����g$�V|�m�����S���� P��ÌO`t�g�/�׬i<�;ڳ� G���o�@ՒX`Wb��>��;s��S���Y)��B�c�� gZ�1)�Vt��B�'�\���|[ж�lN_��Q�7�]��V���+{��8�Z��6� f
��}A�MU��[YQ�X����p=_d�lk��a{������t�#�&7�v0�gL���&��G����WALG\�����17�$�جO.v��:1�Ֆ���?��L����:sr_�+7��]���>Թ+����jX&N2��B�cB���^�s"I,�,�_����Ж{�I7RZ��\4/9�?�(���t�����"��R�wWnW0E���Ⱦ���[��N?۹]:ٌ��
b�5ƕ�o�p���F4ZB�
��[nS�mA����	ydd=f�"�q�ɱ�[$\D�It}]7�����/5r\�<����"�Ǐ�y�H,��?]�	q
�]%���~�Rrsas��Ԙv@1R�ch�!_����d&<��<�_�����i\�1�U@
uCT��ox��1$�'�?�u�}��Y��d�:$d��Q9�I>��q�a�-��"j͑ۤ/�NSI�!=�Е�@����^=�:�,���)����O���>h��#R�V�+N�Q_��R����a���[ZVC��M���Q���i\���.�-z�i�3�,^����N�:?��vy�dWo�Lͫ"�'��Y˝���I�o���V-f��ѓ$6��뀏�)}���|/�t9[�qQ�[�,�樂# s�Gy��=u3C������HD�LPf���`��bp�O/qR�N��>[�[.�K��{ZK��ӯ��k������4�ƅ��T�'��#FT~���Jp�bwi_����O��M��Ri���̀F0���@6��-���B�Jɘ����v7b��Y�����4*%50��mi�7#��~�$����z��I�ޘ`iz"B��^ ��O�������ۖ�;	� iU+��K_pfyfL�:�9�=�3�]�ujϑ��0/6�qܼ��rL��mR�y�)SOP�HT*��1�<�5�~=|r57Q�
h�ቜ��8 J@Kj�,��D��y���ߋ��DO�6#�V� M��jĚ��;S�H��k���Y?���B�\�]�8�Y��(,z,�b�c�.�N��:�L��(U�P^0l���VZ��C����/�Ώ��|Ft5����Э�W��%���V��&�l�2d�8g�p���o�QY���y'�wX9Q�Z�	�����p't?� L5�y΀��}�q%�H��T$J)�cu��o��i����u؜����卐���a�}&�jM�!W�8�ܐ{�eBX��e�C�B��)�>i����]�U"���4�+��J�ola8��G�����O�β�",����ze�T�1�WIj��r�w��L^��Q,)>C��ѵ�l����@��}/�%2�Y���b��*�~RFe��.�K/�����S�V+��B��ӏ��b��%q	���	�Z��e!i5�[f�2�xW!�i��&�HK2��0nÕ<.h|b��%1�_��/+,��@:��Q�K�\?�ٍҎ�Nl��ܺ@�i_e�^�4�Z����
�_C��B�f��[|<�ꡮ;�2 �'S$���_#�8��@*����k�q7�-�IF��P �������pR�FoϼP��^Q}���r~|���0殾�%��		X37��)�^�����N&��ד�����;�M�pÆ�Vrs�p�t��a�
�n?TE�ϛa���+U����ZX�G$uj�zhѵ*���<)s�E4P�m����E��}R��I���eCF|�=�
1�̨�~jb2
��f�͠��X^�e����� �3݀hzh���j�C��/#�#�(�G���z���
Z_EA~��G�a�����%���(!A��kWV�������^;i)w�DW�k��`kb���)t�_)��5�E��Ee�tuH�X��6��i������v'�#X��-��@/��@���Vֽ �]	�ur����"��UzK���.��'�>��3�T����?��)�5�m	 Y8˯k��h�0��	����� ��Ys~X��3/��nf_7�`=s�t�1��^�Y"ؙ������:=���|���A$��OO�~9å� ��<�3��_N���@��Lk ݬ\��PXlɅa����Cr�أd��񗑎�G!��>pѤڕ=�W�B��i����B�	,�j>VE쒇C���\ѿ�f=	�O��"��߄h�m)X�BOn��2&0�|8����Ϲ�'��=
�!���>����_R�h�K4�����&�>�>�5�l�2o N��N��/��DY��dD4�P�Q���/*۔ ��!�ksWC7�-�������9ϊ�F$	=d�Z=��7�7	�N�#�ra+����Uq�3�k�7���˒�ʄ��3����GS"5y���k.^>8�%�a������ER,��A�U͛�6w,iBLV�	�e?O)8QX ,�p�Ǵ%Rf֘Tx-�Zeו�*�ڃhY�E5��F(�`�|�F�t�8�XL��V�}�S�́h�����������-��ϗ���)��fc5��w��hH� Ø��� ��G�4��<��w�=��������[p�6�x�q��UM�B�b�Cj�����;��db$�#Y<8�q9�f�bzJju:���=�-�8jI�Ъ蟼=��?������a��n�B���5uU҆��cc�@�=�!����t�,��;�˫˙��Εnڗ��l0�tYr�"���*2�V���L��j1/�}���9�^����7�ᷝ�1.:~�.�%�B�gzd�V�<��
s{L�5ؐpg��8�����ȣL�)�����Z��>�,*��R:	��6�=�Vջ�p�ƳՐ�F���1!����9m`��a���&�`�f�L��]��[����C'#D~��jr��gL��6���>_ /��E#g3S/�g݊{t�:%ȍ�b^17��|�`+k��q-��8�qj�ݧWO��/���;�0�	@}L.�=�v`�0��5p�o8�W��go}��s�<�H��^��Fġ�X��EfgZ+�P^p|""��zD1�`ɜ��3��ͮ�g��j-ϯ�T�I	�'dh�1C�M1<����,�L�(mi�@G���p6]��t�������ղN&��3 �k) w��Seh��Վ�]A���ޒȕ��)
�]����̥1����"f݈Q�����(��2��5� �j�NR�;ɫ�?߮�Se�_�_���HY��9>�Y�+�.�������a	�נ�!��	f0��|�s\�3�]Ԉ�%,�x���!�̟V�[����6�D� �,��J\�m+�0z��ZߟM�ae�]��be�v���/܎o��r?�Ҟ*ryV�@v�i�HM;I6"����-H��n͸8��>��K/�zQӅGeO܅%Z�}��,��°�"��Z$8���%&o��Y/ٕ,�oQ������C<�/�Pg��!u��	��<�FPr:�B�o���&6�^"��ޘc��Y��x��$o�7ф�/����3�-��	`�53R�P��zbZ��VA���]%�<���E�v^���9c95I�~GG�U"w0,�z�ڬ]�-Fs�&Q�O�s�\�
Z ��d?[���>{J�3/�B�����Q��.}�;ʔ1��t���WGj���ZF�;<693�mG����r���Q�Xm����I�UD�B�F��X�����3��u�E�;8#�G��N�ʠ;{�l��ʮEH�E�0��4?����)Z��˙�q���N4�5���H	B� 4+T���[FfB>�r�ssl2���+��E>�y�i]����t�x֕���X9V�q�$���@��u%W2/D�S��"W�m�{C�J���j����=[�<v��Y�� SV��o"1s_�\D������J$��}�E����k��0���c����ۼ�E�t�`�'bc�A�:n�s�9�NB��7�Z���h��Se��gr���wi2q��h��v-W��ޫ��[�h�8cCH���0	��V���E �����^�-)��;?���%P��&<[m��$[U"yWIH�}���V@5e3r��"}
���#��D4����,w��˙�W ,8L�����=\kgV�vuF��1ù�$�2��)���H�5Ϝʟsa���h�#2�UX��>d��F(���[�O��]�%^�o/q�욋񗴒�M�	���*_�p�O�{wV�Q���Xe��"�;`�2�4?�隔o���7>V��K�wf�p��Xt������1*ac���wAj�S�L\�T�{������`fJǶ�%�C{�;&�j�O޳E�3����;Ė)6é���P ���L�?��G�/�)�q,� 9�&��?o+��t-b8�Ut�/#��?����g/�g��j�����5��K����z�\�Ҽ�$K���Q
C�ߑ��!�K6�ֻq�ӥ�j?�sb�~�gO��<�����E�Q�1&�}r�@��n��U���L<��<`%�l@����]�Wa#��~x�>���� <�T�4� ����C�r3!r����9*Qǹ��D
)G��d)�w28&��C	���˦>��xj�F�!bd\X䑵��J]��i��aaEd��e�-h�K��_�y�[�$�^�Y��Rot��;g�[�垅;����+�\�U��i�N�Rq2uX��x��TA�q� �a*�!�C�+������dJ,������y�j�,���+��k��b�� ���z?��t�����+��Vhx�����<�L��"A[7�j�y�5`��Wh�^T,J�%�+�*ԓ�1�Ņ}�AOVe�G[�5 ��&�Ӱ{�ֆ������O3ж ���B^��:��#[&��ۮa�gN�f�[@�3YKy���@�H�~�;�E@̀�k�PX_>�VX>+�N�D�A���*������26�+pO�=���ɝ�<��!�t�V�5���S4�wqu�i��T�ʾj���sE�Y���� w�2�"��_��d�%j����K/o�d�a'A�T.��-8���Gr��LQ֞|�����I!9F���Vo�P�83�I�|���Uw}h��5{���Q�r=5��XY"j֬9$,��eY�� .�<D�5H�]��iL4gN�cbU� �9w�8+(B����q��t��QF�a)�N��- vPj�_*&��y9���@�r��D�����K]����:�}��x�ִ}��&�5f�+�kbKS8��L��A�:��Y�y/W�[.���_���F����5�0A������T�^s-��߫Hx&{����=�q&�O�'.t��} (��s����=�>8$L.8��<�����UqUY���pP�ۢ��l�ސm�*G�Lg��W`��&R0v#'U,1%�b.�❐�Ki	�e*�S�N��ʐt�f���?%�9�,7l�Ī��\%�i~���R�{3't��|Z���4��Y?vV�؏T�0Iܾʒ�I����o���!};�o�q�IM��:��n�S'����g��A������5ѣ�C�OV<]���W�[�Z���K�t����)L�%�jU��O��=� ����I��Mv)��ʌ�����PC�Y���.:���m��2��[�i��r�S�2�S�KXM���Y�D$�V��WS����?� Es�_����b�����ȕ�{е���o��V+:��q��_6�}w4�n���Us��@�N5�5q��4Q0�aV`3��AN�"e|$�ˑ�)�_=�<��lLO� ��4-L���[b^w�R�u.���H�v^6�z��ko�G8"]���U�0�����v�2Ζ,]P�!ze�{�9�p����~5���\����e<.��.�9����'GցxB����R:b�9`E�?r��&g0^�[.�׹R��΄HE|�S�R�{'��,~/	?�旄ɵ7������D�>�ݴ��>O���}�k&�l�m5fiP�gh �u�H��ab5틅:ٛ�;�3Y��+��MI�! LY��CȃŎ'^Aށ��Y�+6&�I/�9iWq��L����$��-U�1��RٛIG�kL�)�l�|�K$�+Q�ݔ������E�
E#�8�w2�Jǿ4Je�c��/t.1�2�����H-��oA=��Y7#���p5�	ߣ����]��*]H��q*�L	�^�^'<*�g��,��D_����r6NG���W����j�I38��ǺA� N�5�U����	����kc�t�`���NzDN����ŷb���4��1`)�y�u����lk�ӵLJ h�д��!�,Ov��T����i���[��7X�_���@(,��z�|b�<$��;D���o�	�f�*R�gE��-��ڙ�ز�Fv}�5�>��ޘ�ݜ�| ��*c�������d-���-Q��l�Ѹj�G���n�����n~�g��C@�g.W�͌�9a�L�o��۽��ė3*����+~v($h�;Qd��WX���wh2�$Y�	�Z��
�D&�KV]EWc�N�������؀h[���X���ز���`%��;����n�e��c}�R`�B��O�6};o�R<7۶�c����/,6�L����m�K�Y�>�Y���f�8�k}&�C�����9�����p	?��}k��˃)-��|��;��>q4��m�-����9|���B�Jqw�T�8����2�vh��9������1O���XɩA�"�����M���QäLs�����O�3���(��>= iӃ5:Ɛ���x���\Q�
iV�O�<L��K����n��b�M�N�ZꖠC�)��ؕWB	�Â�����UN`GX�9"�A=�Fr��R$*��J����)�BA�T���^�wb ΍6� ��(�%>_K'�k2��ʨ�k4��=	Qݑ��L\M��Bm�v̭g̱��&���5ӝ�V�t��1�t���89��!���p~�B�E8	-��y^���������F�V���5���F'i�À)Zϕ�o�6zJ��,���?Z�!�Z_+1�\�bV7��(�c�¿(PN����о�&_���"#R�L52��%��	��-;�.N��"\��2�s{|���0�jCP���쮐�N���� �S��u�K��>�o��q�saHń��MLm��s�X8�x��$C�U�d8�2{b�Hm8��r��w< �zL�!F� `l�'M�FF��� Y�ğ�s�_��jQ[*lh��_rJ	�0�Đ]hZ���^0�v��쇒O�$��q���`��7ߊ��S�N��N��'���x��
��B~�j���IKJ�ӥ�q�P]���;��+�lV4��EC���%o���X��A��]���Ş�b��ׂ��B�U�Je��w��'�0�|����t�*|�b����f����G鱗�����a�q�-4����Q�Y!p��Z\��ӛ�|���΄�dz�y��bz�8
�D��V�G��J
<�}������/����H-.N��.�j[��h�} �a�ȸ	ov�6S�b�cq),ھ�:�{����������}�0�0��\����nQ�PH�4��N�.��X�A�޿bcg�8�٧�Q�a܎'hf����>�K�0N-7��.L���fɣ!�.s;�Ĵ(ҧ�+$��W��̐��xF�n��#��~w�Һ*b�Ï<�}�Q��Y�14$�����k�9
��2!-4f�e:=N�Jě�6�~㨸�� 
�Fh�6L
E.���vtϫ��\���l��T�6�jۀ��Z��ܱ&
�p�OW{�Ht�aȇF����c+�a��|+��"�,QJjrG�k���/;��#��^���ۄ��d�R_*A+�S��a��ҵw�m��ޜp��T{��o[^��pց�nVZ����L/I�^�dz�@a��'�N�%/H�g&�G0����L|/�l8P`Rݗ��qT����Mh<n�� Xd1�����������;�"����r�����H��"G�p˫%{��[�4/�oe�~��x����2��K=���C�c%팛��-��v�h��(��K ��`N��/�@��9�R;?%�c��@R�]㙖� ԕMf^�������@7Ή":�2�ݿg�,:�O<�SYQN�Ý8��f���J�������g�֚�Z��
l�o
�'�vX���IJ��q�4�(�1E�֏���i��.�׮��u�&�� �ת"���5�-?.ev�I������_�rq��4S��)a1�{�dZ����9�����