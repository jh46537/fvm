��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e�i�h�N>��v,�lhZ~��Rc�	�]^%����<��C�'�������M���,�HB
�?T1�7����qڪ��w�N�8��%?��h�џY� }`0|�3��4L�����֦�`a{'��D�{5P�W����#��S���.n�]���u���\$�Qk�F{�z	#K�%�gs�F���Y�Q�
OLƭ���ZӞn��y���&�V�D��t�H�ry*�}���^��i���`��1t-Bim%�`Q��M�{��j�ȧ�oM�m�ڑ�+��o�6�l��y?1R�>�
�e���>�+���{3z㰟N1^w�����ݛ�+�7a5�������`��I���VI?���< .O98S:���'����m���~v��-�/�}5\�Q��k6�����HS���p{�H�8�2�1�\��9O'��K���u7��b���d����U sPචo�rڀ�mB� �OK3�]�����ΐ��Ć���5ӝW$I�01UMhx9]��d��}��w���B���������WQ��Z�c��LgтUmY��A7P�V�G������ԔTsn��Yx=��O��Z!c�Dw� Î���&�ꤒ�i�l�}NzG-w!ʢ̹#Ե����W��&�P��)U#.�_q4�_���"6όą��о�L��:/i��L�/��D�"ϟ�8� ���$��R!KD���������L^䨼�.��S|et�^�Bʿ���̽~'QE�ʄ�Kd�6��=��;��zM�G�g֌!�*. �ă6�W)�(�R[��\��b�_