��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�{���dʂ�V(��p���ha'�-���/E�1i�r>Z�@Y�_�p �vxm��˪X��~�AbZq�\+���n F�6u&����h������=�A`0���O��`z^=�sdE�����gu6*���n��#BŶ9��yM˭��t�Er�71K�ɘ��E�R)�u^�`�4��^)�dat���E��Ji� �y���7* �<fΰ)2k�龒�1��6��O0N�78������q����6�hО����"�����\ �54�ߺ�_���,���5Y�ɖ��9��h�x�d�I<w4g�s�E���֮B�`���<>7cf���[��hZ[��A���^a�H	(f�VY�7�i涇�:��+k \ݷ@CDNy�>�[�0a�m_ �9���yrា*�֣ȳs5Q�)5����aI�4��X��#I�6��|�ڤ�<�s�P�jg��zL�I���A2q��I�ˮ6�NA�[�����)V�c�	��:+�e]+j��ߥUεrꯚGC�~'I����9�\K�T��@к�	2���z~��'��B�0�Uk,B�CE3
����������z��LB��L�d
	�L[欜D3��pߙ^aC$���q��`�>��f �=����O~ۋY�JT^#?GѾV^G��Fj�ڠ��`���|U�K�{T@2G�u��oŉ����Gl���V�{�FIkE>�22��li�$����tV���,N0�^���s�+���ށ�K��BF�q��B�n3B�����S�0a{��b9	���p���M�U�?p�u]Fnq��B��r���W��*4� ARX���\O��8m`[F�~b�X�2 �6��v4R��:op�ȱ��o#�U})Nۑ�P��D+�@(~/j( *����%y.˨�L|�W\FR�� �^a+.��6�7��3���-{lk �M@���J;�xX�Op��w�4���eelU�������"��8� ��>�|2������ߚL$������*��=b+ʹ8H��y$X[�-e�9Dy���E驁E�7p	(/�����}���rQՕw(*���pD��p8~m="��|P��2�9R0|�l�K��b[�}B���VyY��HNy֦��G��R�ʹ�j��tM��U�Њ�ȃ>�M���V�"�-�禄�%�k�ޕ ����·�X�6Ce�m��Kڭ�Aj��R6���'ۋ�|p	\bF�u�h���?'�Mr��E���9idE���\Ŝfq3�b�wmY�&Z� 5� ���N���������4�nQ�F��^W ��@�N>'�	+��U�>�xB+���	�,[:׫��8Aؑ{��D�������Ƒ��:}Gә�7"�y���%C�:�Md|(��E�ar@��-|U�1��PtMA�"��Ag������k�::C�^��C6eN����n
c�q�������	7�蹎��yT;Dn:{���Q0�f���p�{�:��\�דh��3&����1N��<_��t)�b홅;RF<�u��'	�FSV`�*tU���,�k���J��å���HT����e��)f`�Z<]�q<�%�1�m�.��O꾦�O�$@���B"jy�?>a����\���g�AT8����2Ɵ��ve�B	A��,���[|(�v�@b�w_ɦ+rBF&?/FW=M��E{�P��ʭFg�7/�\rH n?@�-���c�:�� ���z}�<�Ȣܔh(���a���/�V[�?}\����P�u�D�	�W6���nU�~�G�9��jꐽ����D��2�րo��xnv���&˗�|�|��d-O��.N	H3s����fZ�H����ZƵ��H��	H�ƅ'�,�0�4��ڜ�-�Uk�0�L�f�zM��;w��+���F	ca0niߙ}�9��$�������h��l�m`h��l��u�D�Ψ��AoGMB���݌yտ��y�\#����H1���6@ޝ�2x�Q�r}nx�e�d�{�Q�*L��ґ%o�EQ%���b��2�E5rn.8��73fm����W΁?�̊�����%+gG�L~�Gw̱��X�H���z=���n��B�<�h	v}�<c�}����I�	i ����g��f<<�4��N�9K���U�6���p2#~�>2-�w����y�6��x�QC�|�	�Z�8��mX������1�UT�$A�����G��*^������:�i�"�����hu��"�d����9��a3;�A�?I���P��G�h) ���e����x`SU�G��@ƃ���\M���I=�&Y��%�G�0�73J*��Ε�<�(�!Ӡ�AX����c3�����(>sml~w�ʥc6v ��֪�`8΅NJb��X}7�3w�G�E�Ep�1	�D�ˉ��K7�8�(Б�}/dA�K
��bO��T�{3I�y��RB�H����	���O	��C�i�F��Vt�(??>��v�(��B4��n*��+��5Zą܄VPyr���L4K�����������{޿bP������
�����i�wC��]-��i���lli�}�<���	�2������%���Z��1Dͺw��CA�rT:�n�E2L�8���"�'Q����<P"߱>��>kNfN3|R�?�b�Ц�k���,h��'@���Ѧ�(�[�x_�N6���X���ߪp+*��y�-�B����y&3���69��&�}h��Ԟ9ٰ(�3d�F��;Z������#d'ڟ^j��
�D�`��&x�fԳւ�X�#��t�_�I�����xG��3EG�ܠ#"#G�b�����F�\�v����=�052�Ě��E0�6���9�e5���D�׾�Ffά=�wN��P�w�W=$���������xz��+AkIΝr��#ٛd�a}f�t�[�
�i������r@>Rh�!�% J��5g��Ī��o�ɰ����7����M�-�/��G�M���e�F����?#ˠ��������H�ܠ��t����ؚ�(����5��#&�E�����>���:x0V��Vc�g�|�m�՜󡏕&f|��Y"G�ΔrI34�y�p�39�>�(�K��i�*�OR��m�.��Cjw�k��e�S.������u���V?Y���76�_�)��a�k�m�u�째\�Hk��7�u��ص��,/�y��0��]�|��`� ��^�t�X��)�-��}1�(�s�����w���ȅ�+èH��uGq�oȖu�.|�u��1��G�9ZG�N���I�IOs��S����_�\�Uc{�(^;N�R�)��WĄa��~x\���A
�e�򾑑Ůl�R�;�"e�E��Rs�?}���9t�-���I-\3/�1����#YZ���0D�,e���M�Nx-=����:�Q���>��_��:2S����~^��4��K�1t�4_\��5D�D���L����*|;J5�L��s�x	�Fd��{����_)�u�SH�ڗ�t��wz�s�� ����g��1��Gl��&�?Hy_����)()�b��\�h�-L��S2����T]���|�.�xQ�Z�yx2]�d�����ƪ�Q������P2R��h�́��_@�-_�F8-׍��Y@������ֵf�(�o���6ڐ54���z0j�T�\���/�N�;�IV�?-�t�RD+C]�̖���u4V`���L�{&�L 
��aÇpI#���8�mZ�sO����SO8xu+��&9��xu �=����`�t �:��*Y�����,�H��,��&�g��m��֪�eo�t)�����p��j\%����, 0���ʛ:���5֞�0v�]�D*)�����oϮ'�RJC2W�����}�M�z��܄Lsi�[j�-�)K��k���0
48�Q��є��t>�1G�jXB?5��B2�'g�,,�-%�s����s���l�{]�(�֖�i9{�j�4Za����Ǹ������,���ߚ�T}�@��*9�����N<fg���w��%;�d�iC��|�7u���Q���؇���2u��n��(�Yiw��Z����Ӟ>�u�c��ss��'ړ|��:������d�tF�3� mD;�e�tee��j��+��p���8�p#p��4l9�@ʨ8;36�~m�|��� ��y�|�jlW��-���� j�$nT(��u����-�<�{�M(p���ȶN�Z
p)��+�nߟ���r:��^!;�kߧ��b~�U� �7\�pL/��*�J.D���P%���=,�N�%�YY==�Þ5�>��\��u�D��Jf��}բ �~EF���K��d����9�UH���F��5��n��k"oC�k� p���l%酇�EZNt�w�j�	���:;]��)Ǉ��"�A��X�әO������!m�fҺ$ x4Ks��i���?���m/!�,z�V2+�.1 ��9A���*l�=�ׁk�V�쪘���M8�����;(ϐ_��ўt,�Q��UY�0����J�Y�����O�F�����q��	`�I�
݇!w`�'|�U����}Mӈ_o�jx$�D�I=��x�ᇪ�I*��4�	l����������ݛd����ϱ��A��R[������ݎJ`�C�������Ӊ�v@�t�<v�D����=�GQ��JeH�I-��T��x����*V��9��5�T~_T�#�Z��09��TK�s�U|��8��{Ă��Xn�ps�'��:2L����"�͓��Nd�)d�!ˠE�'�7N�>nJ�>vb�%x"8ȅ���g	�,�o5�u�Cʠ��!�7#�����5���bg�1�@�ԙ�eo�z/80Xl
�d�	�t3M����p�W�����&�x~7�[�K*f6��u�CgH����Z^xfA�nx�q�<����CN�DWA�ly�$Hq��ހ����o�����w�����D[�.��5�S�"%�����{cI�2S�@8���Jȯ�X$�@(J.�4���N���7ag-^��X*��2�p���7�wԍ$ď$�c,�M�=����`�X�aj��N-m�l1��%,�aI�p��J�Ҳ��<,?���ݳ�`/�b�� ��h�K�b��K�}�Ug��})ެv��	!�$��e�G�T