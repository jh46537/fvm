��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egz7?���ص�-���q|���YvNH�#}�u*�����Q��H��ψ7K�B�l�J�Wz�R(=�ϓO\��7��8�G�_���5%�jP��z{���)��;���},�)d��ʐ�;�cpmW��W_�ɳ){Wi�F��ܾ��5��Bn��r$���4�Mf��PFMp�
۟�~o���ka�:D�'�����|�����#��|%�ݿ(lf3?sp �A����*Mʆ��^�C̥Is���A�Y��%�߷�ї�kD��>��逑%0{@?��:�C"�o4~���R0�0�Ab e;�x�.4�����@B��]�ʤ̭7�9���4���d�f��{�B����y�c�V^n؜F	
4e�`辁�r���bn��DD�F�wsݱ8%2��&��w��c����Ə�@�A�X+���+*ضk��2�� -Y�1s<��i��=�����C���^�s���mY��ȲM��<�"!�����xEvV�_��~�b�b�ApΚ�Zf2����P9 c�wT���zꅳ��C�E���p|j�~)C�#��N��W�Q4i�g��Ur�������?b��jsi����!RU�-��8lD?8Њ�������톀)�!J�<�I:��c�dREc6Xn<m%3j��V3�G:iS�짨�S�0��\����7�}�#�ܹx��K�X��=�����_5#�Kt2�!D�6z+j-lQA0!mH���&�Y�f���c>�,���m��$���nZ�z�k�1��y�C�lC�6��ج�{�D��Y$(��F$(��jH���u��V��R[|����6cW��5�y��%TY!:-��Z'����LOt��q���x-��4<"�>u�H[x���g�T6�~/g�z�>�'e�'������%���Q=�e��8�Լ4��(����J��H��4)���rYq�����/h*�2�0���|��TŇ�G���Z!W�]�{�w��5�!v��X��~f%:���� �EMذ	�N�K��T���1�n"�%���Щ
t��
d���0�ō��v���]b�P^
P6�f�pQ�	0��jBl��,�F��4���L�������8�\�S7����D�B},����O8�?��=�w���0�M�%�)���yMeRT�\C�6�n��\jb�P}�&&f�HE��lSt��mw��:ڸ���$���"``��iLY_���>��먹M��ă�X���U|����� ղ�ϔ�)�FZu����\�k4.@[𢁐&�-zF����S��m��NA����'WL	�E�}Pz�=�I�t�廗s�Q)�����Su�5#v��r��0�D5�A�o#�7aU>Y��l<�*z@�D��T���������������ƾ�~k"����tfUZu�Gl�Қ�\������U�����Mv+G��R�[O��υ�H����-���4݃ /Z�P��q�\�@N�cS7,��t�Ed������Ή�|e��^%�S?
�~6�UX���2�=ƜUd�����u[@9��a�ݤ�?	 \���05�o�y
��O�
��
.�P�$�WNb[KN���~�DF�S8;�1ޓ���nA�:�?��޳`'h��u���An�[��Q����!-�n)#�"�M,\F�m8p�U������l�O"���Z	ɊV?��O�c7��l/og��������7�}���y��zoV �
�c�[uO�g��tĭ��c��$��]}��M>�����,Z�\�`��E���;�T�f�{���+��J
"����$5m>�h��#\f�Y����8#�L�����Z��QN����tArlv�mԤ�K�j�QYE�� �ĵt}j�ŽG�;�4�!�rztV6�_�8�%�l7Ẍ�PMd���$�"0��~��@I�\�"Ġ�_>�mЅ�h)Q�bܻ��6�')ӝ |�+j0k8o�2��s��<�$y'�XԧB�?ĽZ�՟�T��t��G`~ƃ���$<�����b�Q=mj~�ѓFl x�=p}{߿�y��R�d��\ӯ m��K"J�]+�������HZ�ub��ċ�4~�m�g�Ĺ�7v�,�^�)����GAW��M�d��c(w�ئ� �1�/m{%����R�_'�O]��]��@�5��T��j.���!]n!�qr�0�f�0�l������Lm�R}����#qJ��i�?p����{�Zj̗V�����\��d��4�3_��ݞ��G/	XLaTJ�vk�Q(	 rHҳ���AW9��pc��)ef��h�_y��OC�/+4J��u�@G�)^#���^�z�ђſ�����&�ζ�X�L�'pvڠ��.�/el#0!]��X|�Pq���Z�Ui
�BZ�a� bd�/,��Gb\��U,a�����+9�GC��&P�7l��T<qVw���	і���������:�vYM���,wă�,@̈����1�?)Y%�o�M�a���إ���7���m�n�c����EFya"z�~EW�$�͊M@��VQ�~������9��H��v�>�U����������u�x�)?-C�j5T�1�x�	o;�g��FQi�1a�t >8��0�L�U�ir�n��i����܌ff8�k��O�]���#P1�n��i�_F~l*ƌ��s�m�a�NMTĄhSlF�����cԽio9�����U��-�H$	��}��V��!#ڛ�	_F|$	�K��<=T�R�rA�I�=����b����W��WDs���:��-[ӿ�[����2)~�)�V�^-����F�L�M�{��F�f����p�ԸP�%9�z��f�Z�w)Q��v���V $ʞ�������y�ȓc7AtH��\��T,E��#��§_]I�ñ�"l-���:��N2�l��fV/)��!>�3޷��(U��L�o�f�WStB�=]"!�/t.����<Sܯ}	1P��[dh�u��l�y�e>5$H�T�#ӻ�@�20r����|Ei����>H$����m���z�6�l�D=M \f
��䗨����Z�e��G.|���+a
l���w�P`}�1ʦG֖�t܂��k��f�N�MN�V	�Q)���4�+07hG�ֹ3L���ړ�j�ې0%��/^fD �1��&�+�"�[zxk8�m����lv�͵��ΘPG�o�b�#��տ�ߟ���m��Eo	�Lz�J�aT다���P���!N��E��B�-*'ySw�<��:�yb��ُ�3s!H�G�ý=t*�	��*��+�p����f��n������}����и��,ﹾD�;�#~�������Zn;]{�ll�g��x��y�5u ���a�v��^K�1�s�͗��-��X~;�>�ڨ'�U��6$E��@q�ݍ�W��� � 5�J�e5�M��{Q<MIT�wx*�ױҳ�T� �^��b�^�L�^6�PU�x�ޮM̤,�?��D4��^i��By-@]��d�Q�w4�ED9�&�[:�rb�PnE9��;Zy���m)4Kr	/@���ԭ��n�h� #��[����n��;MT����DJ*\Q)uk��d/u�t����h�"��x|"#���K�)�oMM^^U�h@�� ���=�?s5}�Eq�EY�x2}��tf�����k�2$�A ���q�����0�%�����:t�g}��
�g0'���1��6m�{�hf(��xW�\��v�� |��v�D�6O
��n�E%��VP��z0	V�1��z�s�1���)���ԯN��u�2F�'�����W�Uʮ+2l2Ҫ��k Eǀ�x_CO�"�Vu(��՛�(����M��
@n��w�GV#�J�\)*��]h}�&���T@g̛��&7�Rū�Ft�r��<�3���Ӛ��g�GdrUQHoC�H1�aw��S�2����&��i@1���p�s[����Sm�o�%���z�t�b>&p�<|0� �/�S� t�%�� ����m��i�3�Z�f��Vؼ�	SX2��W)���6<[�*��@������p�k0C����d����.� � ��^���yV��D�"'�u���#X7���/
/��\N[}��T���E3�I��k�s�l~��~o<<��6���1�l5K◛g�l�2a�W������W�<*��G\[z!�R:)�̔�(���8��zg�9����T�۸)����z�B�#�np�� l�qR�d3��܂d���)7��Ɯ!'�����N�g�X�?mΞ+:���եuI'�2���PM�ʣ��7��Q���.��#�D�~P=����;�?"+W�t�}:��M�q�2;n_��/�j�D�!b�/p����Y��e�����ǳ��D�$[��t�A�U����[���/VU���=P�D�p@�ya���GO��X���"7�
�!�ף�w�o�[���E�zr��x����"���]?��$u��P��1\�0>�?�>R�S9�O<BB�D�ȿDڂmZX�� �ք�m��Y���[�sRt<��Uq�J�Qf�ɂ��
b�9����y+^��r�� {�f0��*�7'WC��&!�ݏ���L����rP���=��2�6Ќo!\t�ÏJ��ww'�N�Y�����ϡ힫�����-��h�|Apr.JPv�}�������.�����Lf�  J�)�A~d|�,����p|�ܵ��O�����gA�y_ �z�%���2Ϗ��b��},�(V\����	��O�|�@Q�^"�1��1+�[�4��t_���TX�X<љ��4��H?9��P�Y-�9P��ʁe�E�S�T��d�l��<=�=æJ*V\ɡ�o�-%������4��yxW�/�}�	ɯ�J��m G���}�~�%h�`�����i6)S���F� �Ҥ��v����A
e��;}2J}`<l.�B� ]8|s�"j�.���3�Mla���
��GZ�:�p�)Е�xEl�h(D�+��#/�G��� �"^Ȼ��e��*��g�"g���oVR�0F @R"�E����T��@��5��W�Y� �ȸ�����~A�ߌ��p��Y�mZ��W'�:��P����c�����>��|�ٴ\��k�5 �|����o����͢����25c�����٨"qVoI�]c�)�?l����n�;<�o�Gg֚�<;\_�4s�V:!����u�*[���2�sY��І�)NT�[l��Jc�d]���8���B�|D~:r����=�R[Oը!�9I����fn~# 6��st��i�I�֋�(���d4���,�'�y���g����-�������Mu��]6����tEZ��2b����J�a�_�(�(�ЎT�y-~�}� ��}�T�'Q:9���)���oGSǱ�fw�Q���B���fne�SsSXOui���coq
�d�r��Ck(�R����+����d����ӄ�Ǐ��9tY��$e