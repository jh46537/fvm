��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9������t�qp/�{?I�0W�
�G3�u���0NάA&*"�p5} ��	||)E����g=��+*���4:7���UZ$|�N��ؾ�_��0ٻU]#r�XIޏE7-�,�m���"�A?tgH��Ÿ�F�4cC�� 6��Y�痯&g�oP3��+چ|���}�{���*nԽ�Z�x�2��}7bL�]^)_�Ǹ����B�ʟZ�����x�C(��i��������/���g�J��(��X��̦eⴡT���Մ�Խk�9I)�X1
�4Qf>ȟ���ux��v��L���ZE�W����K�a���~�CC�B�Ŗ��)��(���f6����7��O'�2����N}{�en��'�-V^���� tf�Wu�ѫy]�Jo�-��$��Ř�:�:��Mo�Xf��	���YW�.�+�%�Z⍨=3�?���J�@�?�4X�'�l͛��q�^�+E��^?C���(�-W'����Ǳ]�����7�'&_�������fHh۹D/X�-�F�|ƻ2n�k�F��^��uF�b�T�
��|,������b^���QG�^�hE��6�{ĒP!�A�p5��@��~>}��*���`.� tJ׌7ٔut�&���mU+��|��K��6Qu�)��?���_����1;~�z�s�AR�^a�B�a�l^��0�1s~lEt�Q���<9u�KJtV��_���ʨ�[O�=f�M95ƛU�����:�I�k %���E�Fm��0����Ż�G�TE(�f��<Ʌ�7S�������t�7��ɱ>,̆R�'w�w�>������V�2��eΠ��F�t�<�0���ͻ��U�jX
j:q���#R��� �p�@��e���;�,�[E�Ó�ڻ�Ty,c.��6M��:���;�s���Ӆ<��͍�]�����/��r M�<b;=D6�i=��t�(U�w�����˜o����<�ɦ9�|Y&�e��[�8�k�*a�s���@�0"L�X��
/��B;=0<w�DF�L>���&�NҸ� �
x0H����+�vƱ��(Ԇ�J�1�:�����q��8�h�OW�����|R;�//��ȕmG����^e��kV���J:�H]JKu��u��K�7��]6�Ԇ��F�
�>[���{���\+��,*��χ�4�� �0�[;��h���l��b����\������2���������7}���u�����C��ېc���cZD(�Τz�0XsjO���p�E��u#,����,��������@��2�o�'ϖ5ɠΉs��������P�V�P�����T5|�v�8�t�����#��u엝o�O(��e0�Y8-u�/�w򠬉k��9�q���O}��U�J�:l�W�e����`=S�5�p-$o��ۡ�ƃ_6�h�G�x��2Z?'�~��
�xû�.4����Qs�v��-�����-��e/��5w��� H/��[�!Sz�m�R�̶��ߋ�l��,c��7��\N����!�m���w;��O��[�"��Y�}�9��Lx*��̃]oEybr�\<�*�`#�}.�IxS��u�u�+�x��)#��-iÚG7�p(IS��c%ߡ3��ú��E�=Api�'ٝ�c�[#�/L���"�rF��{�F$�k^�a�"bN gΣ8�	�G!2�?S���܇�@��%�]���Y�Bİ�|��(�Ѥ���
�$G���� ��XmC�M�s, �Cm��VGo7�a�9��Jv��#�i���Zi���}�ߥHݝ��K,;(`h��<+B��M���&�A����f��Va��ur�M�
̬K�nm�L�a�mB�%�lE�΍�!�$�QJ�/��	�gbiuN
�R�m���R��DG�H�|x�q��ab:��d�g
Z���|{@ն��s���V�n��_��&�VF��Su�X�t_��O�8�[�:� э�����.#M�p�i�hS��4�My	*�Y�@Ź%�F]:�i���7��9<_�#�|^�g�f?���\rV��8�(�EִBR��K�`����@ڹхd��|�̨���������9�t��|M�m/ޯE�Zxe��q
I��D�h7�at����;pIr}|vσ���ۃH��q��W���D ^�Գ�?�l8����(C��|�&8�����M6�I~1��9��sד�7��Q�v�O���u R6����.SX�"~�f�>k$Y�*Hs�e�h��n�Wn4�k6��վ�ٔK�+P�� 5�G�}U߃U	�������l�ch�riHR,����cO��J��	�pN����+������M�j�V�.��G�~P~���h�+4���6�φ(�i����%=�Ñ)����C��D��p��>v�U��U�G�N���y��XG@u3C^͡�(�U*c��S��>m@��T�E��Q�`��H]�3
�1�P�%*��^��� !�}]Q��P�8����s_���'T?M�/��ޅ_���m�WS���������17&M%D�A�q��C�=��G�<
x��ߤ?�Vu�/�}]��3�jL������/�� a!���C)�k�Z/XS�5~��
�Լ-,l�|'�c�`�c�A�Dp l�_#m�18Sw֊d-#��8VM�Զ��ǒյR7�/�Oi�]�P>�rѩ�E�ʴh�D4h�9���Tf����Gܺ������UFn��-hM�%jf����M��{��^f��2�ޮ��M���