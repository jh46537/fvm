��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&ǲ��g�m��0�A�v�=F��X��sld*��31rZ�Y�X�(�PO��IF]e6���F~�Z 
*U�}ԢF�a_|h��Y*�Ԏk�����'棧�]���z0��2��е�D_�"����������w��)�nkڊ�ɫ\F�Np~˿;>�q�;����=}~���	&W	�	�Ǒ�M��[�*1��:p�g��F�0�?-	�:���C-�n��U��D�Z�I�
�!��glS�{ B�S:c���L�n�(ؗ���������k�B�"Ƨ�S��{;b��?=����q'��D��x,�^�f�OfxXK��]����C���>*�6����+ ���A��(I�!y
���n����!�L"�7���t�;�J���8����+JD�^aB�;��C
"��&;&{ō�$h�H��].&ˏ<4�S��~�c{w�o���O�WR;j^P3J�a�kf��F��&p��Bq���$�&�L��К�|��1��.I5U����s�$T=y��ё�X�Zک"�Heh4�'���-OV����!��}5���� ���gίP��@g�ZqU���Fw�Jc�yBl�~�ܝ����/��%x�6��\)L+ƛ0����� k�E~v����C ���)s�.�4���s�@m��w[����P;X���K�
齦�"���MޯD�1C�N�Z�� �^Uv��'�M�0>�|Z�=Ґ��N���i�A�T+��O�n:z�2�ZYӯ����<�$)6���t�_�|��*���ĭ���-l�����pծj~|�=�G���'vFl�w�s+��;��8r��J#���D��f�<�`��sJ[ ���	pv���~�ʙ�+w���֏��*��X���=��ҽ#Zy������5�`A��H�!?���Oʯ��n���c�ߙ�ts��d�Vn��x�Znʉ�v��돈/�T�d~�%��F3D�/6�Ϛ
��D���3�f�	}}E|�
��~�]��w�a�I���qZ�`G��(^O��Q������&��|�h5�A魩n2��>4[�?���ED;�������w��^��z�����L���ſ;N7B���{E��?��0]�X?}�	��t����o�$�$,)ΓbgC��d{�k��gk�0�W�D�w;*V�fO����JC��h�[���@Y����w`LU�����<�BB��U濹�G���!�*�|g�2��ңe�d��29�V�����b����f�נ�)У���4�?��p������	��4�a�4�3�H��ᮚ�&��A�4��;���n����G�4d����'�&tG2&?(�3�=-��U��_i�_l�n�Z��xn��*U�W��8��J�d��f�/�7�m�}e |���g���A����ƃ6��"��Ɏ!V�5���^Ri�>:t8� \�K4KK�]G��O��Yj�D�gx�E�f�����.���h?	��-�T�ZSա��c������N:�e��d}����S닅G�� e�-�"���|����3�(��P��:��wݐ���G;Rˠg6M̎����=�E����1�hdn��W9���\����>���H��()'0�]K�E��45EE�a�����_�0�})�u��8;�A��HG(Q�}_[A}���ō���p���:k�Ne+�pu��=g�e7�.D-	ִɲ��Qg녚8���>�����<t�7�r ����M��Rv}�88f�b��W Ψ1��d�����������T�bB�M.η#&HP�S����YB�d������U����)��Gq5̆�$��]��tR}g��}��c�IE�1^�y��XXD������j�~� p�4���gf�J"��%�=٦�&�w��m�b� ��Bު뱆nIUƝ�{�Li��l=�5/]�n���aǲ
g��ē"#m.�N���!���|�^�`L�|�c�t��5��n��_�+��C�9|M��f`�,�,���Z~����ª���M?�E8��ɐ�j%뒜)���~C�`�t�┣�O(!ۍ�6o���"���@�Q `��oĆ��8�7Czx��D���ѫO,�+��"�����[���`gq���_!�����L1<.��K��/���q��1݈塎��T�p�����,