��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�@V����B?:S���/��݀:6{�#��~"���w7��v�:�!�@'��e����A������W����xZ�ً*=.lK�@��΁��K��D~�~� �b�iR���f�V����B1R"1f��!��s:�c-�Ï�`��j씊�(����o�����0hr|&����p1��FVH�g�m)nό����V�5�m�1�i�8q<��V�_/�D��['zz�EU��>���h	X)9U*��)��Cv۠�)����>��~GF�4�%p36����ܡ�y5w�f�	�b���GS��3����~���YCӺ�k�ЗT'��7
���[�=�bT��}���Zԡ����7�X&�D%|�o�홈�7g8[N2���Ҽ`ne	�)�� �h3��b�4Sr$w�Y�xy�h��Ș\��}f��ݫ���p�r�����ԠSg]���o4Ic�$nÜ�)�/ �j�&*J��Q��<x�|��l�wd�ͭA�v\�z�Wh5�
���G�ecr��&$�z�Z�m�+Ᏹ�L,<��ߐ�K'��Y50�^|�#�'a����¢�AX���N �0�\�x�!��C
i
��kz�5�M��}�BjzE��ܔ{�ԄW�A�@)��a��]}�� @�Pe�ׯ�Sv�|Dd�h���u�ue�����"�93xt�Lf;�n8����8j.v%���|����������Q F`����ŵ�5���\��ι�3���ݪ���,����b�X�j�xy�����LM@������2�D'� Gv���X�R��� ?=ӽ�3t��yQ�ͤAɔ[&��;?�i&,腥>]�6M�]����TS꣛�j-�j����>�����݊N�<|A�Y�[7������0��B^o9m΀���?�8����{4*x�hP�OdGu1 ���c��,:��S�Z�E��²����ڧ��~Zn��.�]��e���1�H��L�$z*0�g�CB��p9�hU��Bkqu��2��W9�?O����b����i�L~��5M%X�B�(���ƃ��E�u�n��XSGM�v&�A;�7���Ş3H�m-5R#Wpٴ�%{}ϞD�֔7���=0���SۮWQ��z6�-�ǀ�ɺ��Ϸ˭Н[;,[%�NW�����chHp����4������5V��R���w��xs�du�cc2}q���:��;�+1Ir�WI���3��L��$Nۣ\`a6P�J��G�S�t(
����ʼS�G!��ه��-��>8e�2���a���)/A:U`�r���t&��itc�0�(�hN�Lp����D:f�ô��Eܝ3�v��U�#�������WT�"(|l�eɎ�^KWi�ff�ۭ�F®|ꒋ� �]>%4]D���[�uӐ��_��8��s���rq-�6h,7��Yv��4z�����V�$��j��������o=Y!o>~�΁��~D'C*D88AQ�Ͻ�8��5�H������/�C�D���\F�$s3�f7z�/5�B��� 樴��O���.�s�'VΩo!��p.���Ax���G!�m�{�z�L��K5\�y��;0nZ�e�������� 0�����Ϩ����!�e�+��Am8��)��'��EoUpZG*x��S�M?�F�G��V\ş̌�e��&3*��X�q� 4���9|n>��f����$��L0�@�﯍z_v2��m�8g���O��`���0�'��a{�~���;0��1_�{�L�4WE0s�, ]�[������:m
�+�G��� ]NXO��*���/�4j٘5�-M����U��z�Y�`�F;I����z��BO�B��][�'(��g��E���w���p���<a]mƆ��O�q2T������=��K����@$��a�՛~����j��v��wn�E�!�M-
J����K���((�񑂓܅��OCz���C9P�,��?��5^���#;;�4.l,�}�!�9���l�5�_�o<�w�]l�߿'dc����O�J7Js�A�h�v�����9�+���C��y`"a(��T{|"��7�(���Y���#)� .F��"	�C�/�uJ�k;!�g`LqA��h*��*�p!!X0&����ߐX��z'��m���3d���K߮E�~x����� ��)�%�O��Ӱ�)_iz�b�,e1J�Uǝ��Շ\>���[�>O*�;�~S�����c�$iL
/��N������:�O�h��M��;�ճ��ӂbk�v���W"yyf�2g�V�a��u�W�V�4Un<;C(υH�CLu_�o�A�׬��T���i�<V$�����Hau�K���� I5�?'r�i��-��B��9��Z�,�O�ir�B�9�ӓ�{�����G�#&2Ȥ<Y����=;Uy>�@Ch2Ş!l�QऔĄc[8c{9J{\Q;(0%���D[����`�׭P�H�Y{��V���b�!�] �Ӕ�W�xC�eI����ַ����6���F�Afێ��$;i�Z�ޫ�ɂ��ai�����#��~9E�~�r�4/5�8sP�Ibl0�Xr>>T,��\��JI&s��� ���y��p�@vy�e����E��ҵ��Xcln�=�a��	��-�
&�lW�����R��M���l�5����B������u'h��GeN(�������MɄ�w�/���|	� ՞�uu�6,cΰ �|��~Q�jP{8��֋��H�ړ��O�!=9$=���cp���jWL?��we��l2�M=�LM:���o�(���z�h�'Olf(��MR����ۓ��p9Uhp���1rՏuǸ{���Q��&*<�ǚ�:�z��Q��u���ຣ0�Ȗ:���t��8���.r ;��d�Wk�e��'����ؑZvU��ѣ���4ɤ��e�;U_���������0
�#9(��ab���'k�PTu-����3��{��+RH~T�s����Ț���S"րV3(���X��h��I���2@ށgݘ��,J���۷���ru�w�/FҚO��H�qpG
A�_D�<��
��1�\�db�"���]���>����QYw��*�_$72Q�6��9���\����o�[OT�� ��)	��>U+~��T�>��<�Lc+�U4U�@:�D���0���WI���*�+a.�m�A��'bT�y�R���DсF	V�]}��ަ�^J�.M�%Y�L�����g��)Fr^��\ȷ:��3�;�"�5�-b�JxQ���C�&F���L�q1�BO�	�!���i�s���y2���<���R�!Dҁ�:?[��l(��*P/��ض�%���ǁ�#�N��f�+�� ��m���C�|�l��� Pj��oV��Ѵᬸm$L����o�����Rz'{�{5��x��	~7�p΍��m$��^.-��
�=��^>0����i�Ď�Z�� 0,�6�1�:���p�	'(�HNQv�U8���r9bȟX�$�T���צ����iVpt����(��y�*��z���ЩY��FP����P�#y��z�R�g$�z�C����+��$y!ꍂ��|PN�p�9�L��^���rabKJ�' �R���h��J�"J�j���������_��)�5�m�2�X;S��6ҏ qa�m�`.s�x$��毤���R�eK���o&���s=3�TL���e�2= �MNCEժ�i���_�`�&������ @p=,o���m��"�����Ȧ�S/4π|��C�w����s�T�:�����M�SCs!����:rЌ5�R��-��]*����uW�� �)��ݻ�vFq�G%�=�_Jw�lǺp�����;a�z	+�D��J_�����p�L5o���ǔf��J7��@����:��5��vn����NE����� i���B��}��ʖ�iߙ(R�SmΗ�-� u�=� g٭��jO=R����O�Y*>/N�y����Nϼ��=��˪Og^�)��<��=i
�_BSc}O�����uZ�m(�d-�����{����B|�z◱��)��'|O�D��C����f��O���dYI��FZT4d۷܆+!)�G��4����S��燻��+Y��o��C�w5���2�CS�&<�4�~e�#;���b��a��P�r2����{����}N{�M�dMY�7�� O-�󛨗%zl�G_/�)��H�PS�:�R}�r8]1��(�
�zN�:��5�p����s�\f��#�p����;���bܵ�Z6�e@��d��A�p˂L�H�JU�7 ?�%!��Y�#˾�̗	K~���˚��y�Q��I3/a���C����o'�_U�ٜH�<z,/"4bA�&�xMwޗ���K�������h�v�z�'��M��h�ϠjY��V�A/KsQ�ɿ�ꓻ�fC :3���һ�P�m���j�g�XrY�HE&i� Da��PF���^�`e�m��Lx,�!��5�� s��;=������Q�:�Z�~N�<�%�����"!&�pV��`��Ev�[��)�����$���,�� �V����S��Q[��*�.�A��nM"@J�(���r���<.D&E�'�x���A>E�P����U<`t�.�yݖ'0"9�"!h��/0��M�B��_���U�n��`d p�wy�=X�VQ�-j���4�'�����X��YUqfX[��;c?�n���s�G��y�s;����q�sw�C5v3j��ۡP�W<�.l2r3���>M ���
�I�0t"(�G�:XE���?o��A!k_�}���-�����-vfW@~�/#����@�yɓ%����k:�� sI\���������>~�u����P�g��尫#��}�L唬�Hĝ���@�^���(˱_0ߎ�{� m#�+��bץL������[v>��`�E�1�r!�]G���Z��ނ9��^)��@\�ۻ�/��:�[8�e=��lJ9��S��Θ�~,�ZuH�;�p帘�>���A#��y�>	.`?��a�����5�)Q#�I����_v�"v �Ũ�<'��Ak��KF���ۀZ�����ঽFW2��go�׷�\�9)�|�y�:�RL��_ot����1l `��� =N�c�ǃP��lnq