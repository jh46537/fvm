��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�k��&��Bvx�s�!2����-	�C�o$���%��e]YC����td���bQTTn5��r���]��ו������`��r	��ڈ^�5Ng$�]��� ��ڷ$@��VEbs,��v��a1����UiYAY�֮�}"�ɛAJ����Լ�N�$��Q�Z�����I����\�9Z
zd7���<$�
4;���/xLUd���\�נ����{��?ҿ����8Iј8^�6Z�,z�7]��Uj|dӣ�����vE�����{�M>	�V���_~v���ܡYQ|{s�a(�lK����,�>T��3\���,e�US���c`b�()��+!�H�q�]����CV���F��^�~F1� ��+F�H7�IT�!�S�K�-��cW����=��8!EM;�X�ß�Z5���71��a:�CȻe�(�;N1;�Bi��[)�{��c��!��!��~x�|-U航��v<�J��@������iO�
k�ړ*��_ŴF|�U{n�8_�� g-��K@i��i��S��!(�|�b]�x,=�ޮ�XX��k��#G�LF��V63�
t��r�v#0�D�f�(:���.�W��7��N�K��j9���u�J��] -Ҭţ]3����ڎ��6s��vł0)���P>Td2�ZL���N��άb�cH��m�5�O�A�Y�����R��έ��c����3��q�i�q��+�d�i��%���a�|��N>X|"�?�W�ڄ��3:�f�m��Z��#>]9�, 3SK0���)kSlG��V��:��=����>�ޜ.2(�c�,�P����b]z�

t>V UkbK�f:[���ϖ,ENVG���Q�^:y�1E�A��cաCď^P�j�>�v��:��v��B܂p=|0�??����i��\��hL�(V�8J�S��L@:#�%=j$���@���P�Ģ�K^���T=��9��t��EU� 6��#ga	7E�9�	d��"�Y�\�ԇ�&zdϞB�B1�i���������+e�C����
[''>��%A��Ea�y�6�@j�$�N>�&�+���S�YN�q�@�2{L�o�U���/��B�Sb��W
���HA����ysH�0}U��iz7UO%=I^߉�N�`�s���	�i�eqI21���G�A6x�H	n�/�yv9�.8��a_��4��0��޶i�$ٿ��gN�~��#9�0*�&�����6��������3�F���k��x�=�EP��sտn��	i�o�#�J��^)=�:���M��J���?/�>���1���RЛŽ������"o̴��[ٽS�������v�������@ك
�&EL�\��;)�Q�	�u7Ps`�`�Ũt0�I���4/�h�/r�/U������������I?8�� R�Į��2I�@���n��iM�-U��֎���$�?\�iۏ��5@>�lb���^� ��A�q�aR!}5��<���r��8��粵��2����=�R���
�L) ��~��JU�C����qq]�����������e(���4�4~���meɽ�/y`�|����%F������O�cp����+�4���lZ�ű��i�'z��oK�=�m��ȿ���.5z���Ǹ?��,j�h�l��b=\���$����8�.y�	O/e
�#^>Z����?�p��\X9�]���x�|Ԋn��k��p���*�	K�2�!�0�~��i�.���B�s�����{�!o݂��p.2�jZ��5ԇ��7=����bd�C�?�9�=�5Z͕�Gn���)}�Hqr���J�U�[`���E�	��q�.p�(������A��lE�;�Č�ϼ�	��i�eZ�ie�C*�IO����|���E��� ��zT�Y~�@�w 4p�R��=}��@D,�}�O҇���m-I�D�vyȂ\y��z��S�`*��1���35�N�V�.���z��5ߕ<nF��#�o���/E���Q�b��j����|�ޠ�C��J,;��&��>�6���fF���+����e�# Ê_V��C��I�Z�����a�<�s۟��P�7����� �&@�ޗh�PF��=��'<�r����I��̜�>7��Y��ꅿ�5�����X8C�B?ܹ��9�*#��*�H��<�R�K��vca6��]B��W8��hm�P�}�d-�2"+i�d��H��P���GQ�(�E�����wM'^QV���"�q[&���	��>D��B�>���ʴ��ҩ`�n�ʬ+HV�$p��1�&�H]�S�V�?0�H>/?����ja��J(4y,�T^��E{���cI!���:,�.RF���3oYXg*��!,0����Y�zF����<a+�l�(4�>l����)�9��]�༈mv��h���ۇ��|]�b�tyR2�Y����O����8|g���"��a6�n���0��П�1��e$�p���Y�RhL9��Kj�<4��(l��4X�W�ܺ엨|����U����o�B�C�ȞrL��i���1�A(�g�=�U��mԽ��xh��H�[�6�cҽNR�}����f��L�]���c��e,�bH�;�
*��_���
��)�i�~�]!�-s\<sGű��'Oj��
-Z�	r�[�Tq�^_jZr�H"pź��L�*]��g��1+>tQ��<��6�-��Q9�1�����R_��Q��;� ����/_����I�ލ|��X�w�̦��*!����\�a�I���\�D�bx5�L[�k�g�z�r�!�2���>��b�	�6��!/DO8��7�t���B<�h���q0�`���V�mrh咋��@P�G}��`����P���`�]�( ���͸b��Hm��G��cq�$���37�ϣ��^`;�3!��R�%O{��"��CMffKr�.�M�7O�dH���W;���"&�6��F$H���)�^+�����1��3=sX1�X����O§�:�.�xh0���I�\b.���pC����h���܀Ȗb���O�b�b0��(	��y����Krw(}>[m;�mi_�Q�*`�*C[tJn�YO�vn��u#0��$WT _ k��=.�c�u6:����`z���@��p��v}w#�{�f�I�S)�Y��1��7��]@d���0G���V�?�w��,��+iixR<.5?�Κ�� r��DD�'���2�;Y���E'>.�Q�A
[�z��B�<���:��g��߬ý��X*t��w�ov�A
�%��#���`C#��D(nۘ����k$;{�6g��	��ֲ���{(����ߨ��j,>���7���
���~Ҳ����9�d�5O�LN�SӮX>�UY�C�dQ���14_+��$� �����Z�-)���P����m�|�Wց�Qg��Y�̇��]�x�fj��ڙ��7��ŕh1S��������$��)N�}'���������;TB��^�9۷z��5`b���r�D�鍭L�ۿ��S��~�!�1SNXCm.�ur�u�[_��6��z�j�JZ���<(I�Skdb�U��?�q�Z1�0.�ô��A�T��\J�įy�(;��^�Y�P4���li`�?�,#�k`	3�~��v��e�|z� ��hI�S��Lx�:ؐB��v��G�Cn���)4��Ѡ�iNU�T\;�����P9b��S�*��|�_�mi:e��Ⱦ0M�8઎;Y�����O���ɵ��sx4�����Guj.[�N�,\;�!����	ܰ=��)����n��O %5�39�f��V�*Ė��a$冁�0�+��3WH���$7�頭]�6+վ(E8�%� xb�j�¯�^��FO�v�"q[��)������}``��HJmj]_Ls��\�!-l� *�:���i �Ov��g|�-�e���68��3��HCܛAw�'�r2��ɢr�DE���Q����eߢk�X��]�J�~v������c�K/����-
�@� Y$�ax^ѧP�gl��'r���VX:������a!έ��_��D{�+v�Z���~舳o�hz7��ڹ!�c�6tnF�;uj,[�;<tŃOr���Q��ׂ�0qrWH�44�`%����zJ����C?��3G�XKC TSo��4��B�j!�ϟ��Q:�D6a�<��J��!�����L���(���h�K�)���wn6괊M���
!
M\��!����7Iڣ!� ]QWG�����7�P��w3%f����2�0�����,���o��KxP��/L�
���RaALc ?��#�����Gz�����C���������:�L�-�<��l Qh<�XW	��j�����ÂG�tf�Ĉ)��jF���`P*�#�'�PFO�,�/��y"�X��fsŢ�Vk"����w�"`4�+��TJ,11^�y���{�W�\js_c��g��D�R��^a~�V��ᐴv�;e���UB�m�mp�G7������UiS�x�|ý�}�	|-��,$�sc*�M�'���*���/f�ɹ���D�9L?ʳ1�g�j�|kLDy0�/ҩ^±v���;�h������N�Ck,��ԪN�tP4-Ϧ�!lj7U�T���L��)�|�`K$pr�g����l�?}+��[n.N;M�C�>34��#�{�Y�V;]���g�ٯ�"������w�|w��d���f5>͓��͐|��<T�u��7�&�M����04�6 t�+�8>)Ȅx��o��9	������b�.F���eU�Eؤ�{m}��X'�G���`m�W�)'���s��.�ʢ�\�g	���'����o�hƧ���PH��c-*-���h�G��+U�i�Ur�q�e�֓$��22A`��^�)�,��5�x-DV�W�%N0/����F��B�@pZ�)d���U��$��T��h<y�_	z��1!�`�If�=S�@8�����������ĮZ���l��L���J��$�/G��Sl\���C�T=&s�b�A����d�[�y���~Z���=�I��N<��]��9儿�c����㪿�kX�$�L^�%��٪�ӂ�&B���0��@a�l)�k
�z�^�����B����94��۠/�S��v��U%����Ȃu�>��ӌX��\���,TƤQq��(���i�EO�}_�Ė���#K��t���i���O ��Vtk��$��$�Cz�>zhj�1^�ڳe�]8��ǣ������D�o���H���}⮍dA*$֍&/�ĕ�D��7I��Ve��~��Z�~W�G���.܆������u3��O!H~���W�8�
��j�h�+E�����ˣSj> �}�JU�(Z���ԝ�4T�|y�KZ9cN����'!�L^�~�{�O�f�.�UyŖ0�M�sv3ڒH�4�Ѥ௞��M�|�
��3��V	�H�3rE�,6H�࿑�xE�������2��ݙ&?H��h�%V�rX	B���>��Q�>��k.�V�Įq�*���@���^PShѳ"�3HV�
�\K�6��<Z�b ����U��2
��'wJ�=��!�|�ʍxlD2Q�ItіR�{G����S(D���Rg���'�Ԅ�4l���X� ����_����"B��sgGI϶b�+F���yf�P�C�������{<����(%	Rw j��Ī���Ȝ��w�Q[:U�IDtf�k:ȳ�4�ʓ
$�w��U�;'�ml��-�z�St{o�F�n7��ߡ2��$�_�.)pa!�����mr�f�VR(�w�V���V����h��fhS�im��'o�h�[�W49��3{���i����Ou4�i��0D����B�CRү����a���6�c�`��~zvG:����c�y\o��pJRݽg�����8�74��(��u���4�;��\]���m�ƿ��0K�ת&�Yv���c�Iy=1��{EН{DX6��_�[Y��7�p���a����Q6��Z�g?B��g�	��G��I�E`ג��]ף27�7��I�
�p�F��K��k�t{�9��*���(���`��տ=���JX2���ⵥ'�?����0ƃB3���yMQ���zӥ�N����2�O.��vk���˅ͺ6�s'|��Ю��,N��*��u��}ps��o7x"�.$0Fq�>�o���ϚQ���+v���0>ͽ1���ةG�_W�[��ڲU����·�+�׊��U#��2J&�e� �YB4j0\7TJ����[�>dxWp��5��c{V���f�qG�"��cB�d�A�ˡ�[��Ք�$c��loּ{L�����mH(�ܻ��&NHW��W�H5P��q ;��'��^>�$`����$��7WLa����ښ_��5�*��a&!M���J���J��{�'=�Zx1%m>������a�Ub8���V���l��7`����x.�8�zM�8+������G�:_H3���	'0<�]��N`$�f>�OT�H/�(�ᔤ����c�o^/}h-w)s�s6ۯ�Si�o�r0��(���|�+i�|q/EQ[�x��~��$�j[�g��4S��s�d?�Xw��X�b��>��y/L�$�ҡ�+8�v�<��y7�"��aIF9���#�̭�>�� �Wm�C�,K��njd�SѮ�fY|�p����j����.*�\�
V�<9��IX�f}���c1��l��b�T�d{犢�WP�_����{��mFV,�m�	����X��������|�Y�&_��vH��Q��:���Q�D�k�6+b �4��&U�g<h�*ihR��T����~�F��] zUN����� 'R�.�٤O����{x2~���#$����U\Ɇ��1^������k�P��0|���E�M��W�U3f�J����tE%jכ��a�("�$ޭo����GPu�֠#,��6���c��j�M9:aX�Rt�K�g�!��#n�M �j>�G���({xOQ�ܻF"5��J�����
j��?_�j��M��P+��C;�i�Wͮ���Ʋnq��������Qa�$>�C�R0�}�Ȼ�N6�(��}���-�HM��� 袑��A��1�UP�KSM��y)ˁ�	�b�o���|P�1T�;�ݰ�@�,�����o��ayGO�*2s�� �z�����L&H�!��@q-T�:ʣ*�aX�Cm>-��
�_:z�^���7z���D�	R*�*�y�i<�G:�K�2�?�%�f�<���A	~8���SX��E�ӌ�����W\����p�9 �����v<oGTZ��.�t7-%�5��h4��D��'�M*�yu-�1u~�b|TʓF��Ώg����1z��[��Ћ�v/�V���N�eo}���T���~*#�:���Uص5N�ޥN�"C�}NhN�c4�0��!�VSح��|?M=vUZޙ|��?�GѾ�,�3��]R��n���nM�Pv)Q��^0$�9a��{�&�˪)w)��2m^eN歇(�l[���s`�vCǹ����p��Zm����Ҹ�<p'�{!0)\������ƹ:��`�U���e�st�$(��?�9�G�)o�S	Y��Չ�aA�<v����a��R�m:}R~0v���K��PS�WvX��*��EH>������OKK���$�I5�#�����C��q���m:sF{h�>z�72��+�µ>km� �&�Ju����3�N����ЁO�K=f�u�HHN*mV�%�2?��#�\R[�|���**@�N���e�(�h���+�>�;� ��Kjf��a��������;k��c�U�ZW�����ف�����Q���ɽ�/�X�IEN��t���6*�	[	���Vmpr�m<¡J�B�E���i�bXPNe��/�=��[�s���T����Ouo��|��� �n�9�+�f[X�PK�X�o�>�b���3���9-LiX�ghY22`�xp��*���l&����B��.Z�����r�j;���@�遴\����t�D��7�n:��ԛ���x�G�Z��#���*m�����)<E,�ƹ�|��.	��m���u��| ��B>\�k�X9���P�߇�(zP������ٸ��h�I��A9E��frף�;<�i~�%T/�&�[�b�ǂZ�~��M�S�z�)\p��)*��̭8��m��N�o�E,����V��B ��F���9��{)��RN��)�����	.#cPGO��eJ�@H��,3D���70�vy��~`�#Ӣ7@��(��7� �m��"K:�ڔh �U��$=�7#p��\~5'E��ꏈ�`�*�W�^ }�};��l������&h6�a���h%���G�,[��pFg���${�3�o/
�7�"\5��*4%��5���g�I�4���9�� �a��/ T���w�T�[�F�B��u;�)M�a_�Zjq�]bԯ&�2D.���#�\F��E�c�ԝƬ1I��X8��s)g˴�q�1OeZ��d�W`f��%M�a���\�+^O��N�I>��
�*�����_%0�7������yCn�$�d�R�*ź���k�B��5��s!�E"_�1'�@8�)ѳ/�o�D�W��
��0����vf�+]�)lϝ����97F%Km&VOm��42P�qi/jal�^EA� �O�O��D	v���ǌ9dK$W�GZ�鱠�D7�5�|đ{�$�]���&�updD�%C7p�&E�hyA�cn$�^� �;X�Q0�ڄ�p�L��߻��p%I����3���a�����ĳ>4C�w���'��3����l�}%�~�U�Y����FL���:)y=���V��C�qhѨ�����[��-/)���0���-�+�`K0���8���W^*X(�L�/{u��z�O���)Xk��U�ݗ���,x3�D�"� n��zL)޹6�� ��v���o���T�X�Mw�z�#��T?��M�թ#3�s�G��t�E�ò~��d�q�j�ap@&�G�$��y�7Nܬ:�RC\���9�O��J:w�Е��|�cngE�4�ч�gr���w�鴚��l��ڙ����v�K[���`WA���ot���L��H�U���e�ɳ��v�ϡ��iR%�4S����춘fP[�2�+�w��xPZ���%�>l�J=��H��>�im����y�����1����i��� T��M�+���QF�]Unh�����KNNW��h����W�c�wxc=�2B��A�G���.q�� ���AyxN=�K����)��(t�z�aG_��2y�s����+:vFz#/�����]p0��9d^5��Te+��u���Z"��ޣ��VA���X�{�yù��`$�'���>�+��YVrL�~N�����[+n}��ɽ�Zƨ��xe�^��>�VhW�."RN���eP��j�q���:�{t.%���l#���2H�|,r ��i�����M�`HOu{K���� �@Nvő��[)L��2�E.&W��H�ƴ��&!����<����L=�U�7�L�^��R�O��`1���a�Q4�l
Ɨ�|��B)m���N��CŃ;/�&s&�M\�H����m�o�Q��q��V�n3}cҟ����9�R��W'�����G$�R�Na]C7��g��G�w~uns��!�7���Ό���~k�W(G���&RM���jd�dF�B��Ϡ.e��&��B��	6�O��x+~�a#����b��=�
fS�"�6|��_�NH>^��Ⱥ9lL�w
���wfn���̇���	��wCA��_-���	����Ml�gIl�����)N�_����N��h��?���0&htC��0=8*��h�>������DM�Rbz��"k��w��:����U�e*���A�	��~��%��!�'Q{"E�K�Ũ
M݇���I�8'^�s��W����mǵ>;��$�ќsDF�^BQt'����c7���"���C�ϫ������S�Fy��ů���8G+��C�OC�﹕܋z��@l��qM�q�g~Ǎ�g�ǅ}cg&5I�5I��kغ�Yet�f�Q��L�B��}I6`�Шα�۟���]7�Z��}Ź��QP� N�F����g�S0*m�4������3}<w,mƋۼ{O�����Jf�5�P������n�O�(�޵�/���IW��
�$K"]R��PN����Y�x�����77�SL��o�.aZ߲xaݕZ֑��i1c)<p�u��$䪈���N@ﴱj/P�R�����3���5j?�5��g�q�f�n�l�)sC��/�r�r�%��쨚|������1���& �f��_-9�qB��*� |�/o�����,NF���]����/�/������G1�Њ�����! ;r�b`9��/��1T��!:pA�{
���b��_�6;�����2]�/�%��
)�96��5���!:�JW�bi�%vU�P*<�<�]+��^�w��H�f�r� ��l����k���x����M&���4G���k��>&O��G�I���㊣��X?t���p��&�H��*N��QkZY&~�
��?{-�WlNV=þ�'q�J�c��Ȼ੉�f{u��w䵠�b��M�Р:d)i�"�˭ַ��z���,Q�?Wo����o�"��7������I�e�OYo�0��5�����B!C�w��W��z%��H��x�*�1��9^Qz�B՚ۇ�j��6��"�g�}7��jԎ���3�������˔t*�i}EMG�Nj,mD޴J��{>=uEe�W]E�����z� �!�lѽBV$�VF9C{Vbe�yj�R�[�XR/�1=��ܞG�y[�\�@�/dMvwVT�X�GQ�8k@��8����N"���O���4�1�O�U��!_^.E���1%��*�������Ո�R۔\����4�c� @r��(�j��43���PTfVE��:���vv��a_է��.rD:ͶM?ץ�K��:�E�$=��m�_���E�G�B[9����yX\�;�U�"�r�RT^�f���lV7����g��	}�Qi^�F�D�8����	X�$���-������K�&���d�/m�3�a�h������^_ ���ې�t�Θ��No�	�ǭ�d8��^���8�6a,冷D#���̞])2�ǙNi
�z#���G(? y^�(2�g��O[!�u�Ɉ7��z��� ��#��$x4N�C<t[0�*'�4hw��M����O?�{$�ׯb�Qg:�����ٷ���O��8����&�N�`�%E�V����%wn|@����Y�s���޵%{�q��!�g0��4M�h(c�A'��͹7�T�y�݆�tx��H��1�k���kSIJ+j�F6Тg��Չ�`| �YD�O��?%"_o�)��t(�8ͤ7DW,�R/[�ԒCZ��d�#�3�	��� ]�\+�.cI4O9<��.�ɬŅ���lm�\����[k�R.c�(����BxUv�&ZX�P�G�Mzg|�e������jl�5�3:SJr<c�ǉ0��oJ)��f��}ɂh�}ȥj]�+�D[h�(�X����u;#sE"@n%1��b���J���ú��Ώc8������	�	��,j{�q�Č����-'�6�1��N�0P�eN�cw�|K�� �,i�7�/}N�	Y�=TϫY��R���91�WN�-5�������a#4�n�F+�sƩhg����G�>��:0��-	E�)"��ۧ3���	EBno]0�L H�@P�	`lc�*��P�x���<yw\�dI�8F�`�%'&�>����_�A�W�u/���hL�֓6A�I� �1J�0;�LMo8whA(��V�m?��s���˒��1�:w�,ʀ��:d�,�W9X��v�1������"�X}~z8�p�aȾ����p��p�/����s�Bf�@�@ב]�_ �a�]�هJ^[�x�+~k��[)o,�"�P��
��P��F����	��&455��
�D���oj��6$8��*�����;�%�+��w�tߓY�r�UW� Hj�/hI�ѤPk��B��9:򳽏Ϲ�̛Tcc���8��͆�yq����Y���ʡ��(r^�Җ���8����!��?��b�iJ���
6��`�\%��w�s��0
�%2�Y�[��@$n��OM@���[���4���Es�Q�p���x(g}�8�I�L:�(���\�d*�Z2�%�g���6�&p� ��Q�%7��#c(7���c����n�2��)!����m���ln������m���te���I�����Wg�
����\�L=@ԃo~:r��¹���M�
��t7FC�Dݑ`�"��9��1�HںE�p�:x���W*�zGx!�br_��8��>���)�3�g�����g���6��+�¦�䚈1�\�wt
HU��a�C�'Ⱥ�/����;�ڧ,�K�^�(Q���A��2�� �r��
{����~A� 6y�ch:���H�;+V�RN�
�(�W�*��zp���z����&1��N��_���e�IG�OV��w��/�����S �B�#
R8��@�
J�c(-F�]�Mm�֚��G�faC8�����C��wKk9�L7{H�����?�Ն^وa#E���η�2�½��D����MͿbo�o,s��Цm̟
�(�Lw�%�0OB2��צ�:�I]�յ�r֋���zJ��u@"�mOW�[�	��wA_���-�������w�u�bg&� ���˶�t|{;Xj�o�wm�c�luB@wK�k�q�j`����������bq�z*�%���ŵT��~o�����;�_�+�d{�b9Ea+&�!�'?e׷��|҇��)�h�j/�8$:8�^�_�6�r%r]��
�:��o�e���Я�X�u�ն��������t5������]i���5BX�x�oJ< "�+���!��f�