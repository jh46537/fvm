// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XrG0Zny390cl8SpYmrlhhsauxCPoux62Is85c6Zaras1IYICGuk9Y/SpZT2ko0k3
d9QkZCLlkaMVpOX+MirqBqB0WlJdQB5HQ9SaMRBUQyOAfP6ybY5BHClBSyXIqsyb
J+eOJTDDuMLgM4ISmChQN5sSjfQtPOwx9GJ2Ex1Ly6o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5872)
n9dz8aHaRZYPrbpXldxQP+6+OJSiRGxZ5BwS1V0iXg9xqpoPfM6odowYa4kop2s0
0teYQSPwlpydnBD6stq+CGUvbnGJq2+JAltnlAqJw3E/XdTn90sTbeva8A9PIzv1
BrqIw+ngZD5OylP5bWvrO2v7IzEXMdlPSzr+cFE1/BQ0/1znEBNrgiu/j6zcyQ6b
seIfHVOrUuplzMe5SU3RpPXnTSYisgAs7j3L6cc+HyCTjEhKg3prX3XToPMr6GXX
CB0Z1JLrRvUkVC51GMT1j2WeRRQv/PV8njpOqmf2FIJxlcDNCTZr5xj+Z3bArhxV
Wsz4bVCmZ0U7ytaoxpgmMNLTJ0KgG+WmYkVJm9Oq/vwKnsg6gmMcM8yZUxFrQlCk
q8Mba6DuCM9iPCZjfT6JIxRJRpn78LkIhm9rhg9+VztJGeg9ooYERyTaXwc0WHru
mGDQOJTak7KC1KEUaDbxY7NyCjBGo3ptehQhwQ6bFJPAjmYRIkP05vBnLdEVU1Vj
P7qa+8le6ZV1uwB6scApTUOzfQWudf8y6NdlxY3sUldFtUR94DEaV4eo/pfnMnu8
8rF5sDkVol92Jiej3BINd9K1IVwxMbciFlNMf4KCD4TKTI0GfMRifmF373VAyP5q
w85L3CCWt1mo8L0cwYrUVYJhLSffwryyDTYSzjZX6sqFLYNISQ5nsMu8vjWmviDD
N9ErKBm3Yu709dXjMT7q/Uqe6A5LtetifMhpBkadDaS90GC9bu0Y1QTKNYiMyI6P
k9a26mwBCUYPwxKCUHgy9njmGRa9W738dWamSjuruByhjd1m15cq6Ynkf/BeW21r
al0fMwtirqhhkXxqNgwE89CIshM2nk57cp8jnZyHLOwzokpvWMbTsSLkhGeuNv+a
r6g0RJX+THfzOgZjJ10wi3NFFjCSgleYE8+LSl9Z+1Rg7DzDLldUZbc2Rry9tVXb
dXb7hoE47G3iT0qBgUcnTKjaigIffRmwudhxeW8J93rCNex4LD7s1A95K7QtkG0Q
A7spsFQdJttBXIj9allaFpPW8eXiDWGLbYUa+78vo3OhtvbRVZmRtnbZ9GOI20Rh
9cUhBmFSXsGIVcAS72VujYBI9FdBwrDJ0plItggzTeyhOCzfIuzSHz7ZBMCMoUGo
kEv+WeEHJvwhJLWKXeJ4P18T8Vy35YpblRg55XyJG3sTPmjkBDTNIdju7JL82bn+
9NoESpjW5zmrxTTddQ8l9ClZ0kUKrW3of0VzSfk1n4lLXW9Ux1ScWQnbZCvJrJcH
75VBqp8iWXccpP6tRXGGBrZG7ReOVwCo2JsD+kBOEFLFN3JmiOWWO6nyUPli7wJd
m31fxsQZtkjjoRcAas+JAinuHk30mVbZpGV7IGeqIl2V7c4/LH5xcM9PoxRM7LIv
qoul8QHkkbGx11CINNmZSHxckon0xWMQ95yK4tTAPxvlOL8puXXblI/THoCpyHVg
U+Xa/iAz02UTGSO/qjFaXsZImwQq40B/iva8eu+BIgfIp0X7HXHypLYNTrfRc2RE
DSltnPnGkkP9Ad7HFHeIwle8xwoTQog8bX+cjI8NralRpYz5WVHtB+OiIDQrP0K1
off+udsSb2JV3oKL0iGC2tQ949vjHVtsR8pHEAXpLaaKmTeLoWHZtEqOqHXJ5/o8
yEnndlX/2X2ni455XppXBKfdM5jAl+w2XCYuCAigUCA36VxWImxtiiyQBYLnxehy
jafEif5SMF977oxhpARtt4zFq/CtQLwWoOxEe/NE1sKv21YQriMr9lybU0N8PZae
dNnMLBI/wvOx4C9T3WuKJgfaHuqSJadZXZRFyWIFqjTwJtbALnhmURL9fFpGdApy
W2hjJLpBuW5JpiJ2fIIc/kYv31qvxqYKN/gCkPPutstF5zqv1qWQifOvz37rRKVo
kZ62kta+YZvFAhGBWJqgTxKxaQr09s+xYbWT/uRIiv3vOpsV27VouxZleMmiufVV
BW3KFtvieWmY+ZaVA5BY27VzpTCks+tMjYs9uXUZZh14wNdiccKrnphcADO0iOsl
j3l8Mizptl2qCLR9jCXXjPqgH4jlGo3w+Wx+zQLSR6iKBJOLUiVjY6qD5nx8ePB4
sQwkoqHgz9dqYhkFqzbzOO/SI2h54jSOqGh+OgEG7VBpE2sagYy/RdlYZlEmbIZc
gA6dqGOhDCGePFayx7tEYryv9ODQXfPuMNytFjEt4+YtBGxe4JyipD5ALAnUbMfK
zOkxlCTvQt9zVD0bDkKmkmmVIoiO8ul5904U1dpC6koLFuuic5Cy2DGR7B1sBDtE
rSOUW7uJ4lSloPjhSgJ+fCqUqYnTweP+7MK5qPI4ePFrwBBr+itI4kJEyDGxMYkC
g1LJYRl0x8AvfQEp26EtKWHeeovgsf/JTXqQzIMg2JGVBFn2ge8+HZIr8kQaHPpA
eDp4x1mh2c6S0b/dUo/zpS8cO6ccpQJ4rOAPB1VD2jt1Eo1IwRY49PTsLu/h3d8/
rFKFEdL1siGvuDq418kcxD7aWLRgNNEVLYqLvqP0SFDRSY5alNeHK/Xb7o6GCyVj
7SeSjXP6IY+iG9/qsqA7CutT1o1Vy4xYDJhUTsvyFFhJkWzN9i+zz2fETzh9C3Zs
zADQk17pVKr34L9gb6aNUUZpPVash4lTmB6Aa6bvU0DOXFXaCf6+sMkPu+9OkGQy
itkUeWvwUSVK2UN2WoMtpTu4IeY4JBE/YjXE13843zW+IlV9Nrss9zSlv9q8n2yw
pNyKB/OX4SAuZxLCAuTa1n+7mk9gWetuQETjG2rCz4dLZTkupagN46z3LOb8manz
u230KNaNBObmSMrspQGDJtOO0xmACex73KvCGTcna1DE1cTgIzJz2rkTx3t37vPe
vFjkKBXBtu+UVy/kyv+jLbH7OJw3PQ2G2V2DgWu2pR8cQnfdeF3RZxZTmb0kUKsa
ziQK/ViVLYGmxHSqOaaSELnKFRMCZGIRNTCuPxF9wCgk2nsCp6y3/y3liGDnQmnz
k80KpuXkdyYgwZqnhNTSH1GF4EF6qdNXtThGY9ITqETS60IjHsRNy+vBWDeBeJi1
If8sujwLpA39V3LyY0EYZVmwp44QNtjG2ciakvH5ZugmdXv9dwHmiLieg/92FvDN
eJzPZtpeQ2/MwjE3qPJ0+L4IfR2RlnerRjmkl5ZowWvRMjiAXZHcnWv1z5Qv75jh
1YvRF5PMWBr2CUc5a87hz4H6rvWAk9QxYrAnutyzMIGuDFLPu/U+lGJp5HESDel/
wnrDTJB3FJ9ouhoOOINbCbiWxuOgCrkQ/2islKzqbvA3hmqteAKkFSC7ffGZyiAC
g9SlBNFS/gKlKeHKv1UsCbB1et+YliVQIIWy8eqR2ffxIKI+FKc1YUXC/EFkzLms
oyMCjQarR+wPaZ20K2GCl4dCodLTJkhOMfoKqolLNc5ZPNvoKiXFxknfmf2oVD0G
8ljxOdQEzQfAQa+c3Yf8gWyxOWcDBcaV8KYT56axoeQB8iAT+7qMtj4obxaLBEfs
S4gM7zB9egxHGOpVGzKNiAnLXtvl/0IOKMkhCUEVcHgVFgA1Le30J+0O3nKlx13h
mLwMp4KhUl6xdL3evIqSySbRovsPHZDMwVdIDHynLXxjdH0nBNTDAAKms1EPHUaY
aAJi189+w0WARvY1DdpIdHNGw5eum/NfeGHzBJAy3aWIiviGGsehOXgH+vnB414Y
n4HtHtmuxjLEaHRO3kn/Mr4gPqExyuVO3zSdZin8vkkJ7Dw70gPUKSt4O32vkOxI
ewnHHnd6wWgyFHZxIIZUMHleiEvtUpeftLcwJhtMjfoUVGraq9jAbWBqgdLzJy/t
QvNhOwxogTEdeBcaLyNcjowEBy7oJyMdz0vwehEC6FQSSqED+44YgOw4dWVi2Zho
TWvAmrtWcTf8s6fkVYM43ySa89r1G7m4nbgKmr+BDbpwy6/51CYbok7uqJHCJi0H
WulROwK/A271otkLfApaS4FAAaAbEneAsxKk4PlR68J+MZmTFuqmzVd+2eGR+ySg
oWN4/91sTOoV9Mb3uMRyYGDTHL2c4MnBQYpCiArYpUCinoKbnxVvjwSOFFBIF1o9
ilOrfiEtsCZkN6inPNEoXlnWSTSlprv75F7mLAu2NehAh2DWYqlXmV1IzU9oOaZ1
wsXTLt/bf/brVzvrFsQMlv4k7zZfRs9ZA1VviwE6c/Oxic7zdmqCAef1QMPiHPPS
pFi6iZa12mwi4n9Cw9BIyY8GEAKJhx14m7SwGvKv7nR842y03uBDfk/W2WGZZ1vE
AydQuv6QrFvlrswucLt6rRubJxjKUNFmK67hi8bBfEnoE5zUVQtH3/3DFp+XGWqh
kShrvQNKWYquiuscnZ50V99ZcgJB5qEpeS/+U/zifNj0W8G2TThNvLZl7iFSTKYa
SKhEMuu6NaE9ad4ZcfXL926ZxAvhSq6u18yyUGMqBMYZhNmMUeG2ivMDTDQbkXVn
nmIDo5+xr02L5qHKZL/Kedwc3syckW5nO3oDxoXRbsHDGgEvo2MkPvcw7cEG/8qO
NSCbTuXsFFyi83Pji6KIvlT7Mr8JHPoUqKLInPNFkkq/iQc/u+00VRruPc8MY27x
VKtesCeCIjuUpVQxmKR4qDif9KKDjM/6hcYd4amu6L1kWP+twmEPDDz6PHMhidl7
F3zzP9FQtfIWsbUHYiovGH9Wnt7uKiySe0elSP2RgKif5FSIQEF6XOjJuebW7OBa
Cr5HP3OdOSXX5jgqBPhbDdBAAhX906Dy1JsqYkDSCVHu8zuNKRjYhG56g+CSn7GP
mLW2Re6MWkelg7dSZZGcP/ga0pREFt2CH+0aNHXdaAcCREjXQouS2kCIRFVzaLzC
VGf9KLow2yGV6gIHLX4rsg4vnfSxpFimPoAlwH55LCt4SnyI1KQiwXTErlI+Lii5
iytaA89IMqvHQ2LF/mYUNRIr0yj8zBMvM6Ts9RkE/tQ7oX1zjCjXdBitsw9OlFaF
cBLyuqGG7jP8FMfU0IdYyNKE529tW69Mng4KtmOf5MUIgnI6OxmsozjC92EnlQrS
o7FORfvhfIl0XGi4Ke46urWuF1LTWiTzUaP2yIheyri8SNnljxvRDbbYDLrdOg8b
4Fzy4zcZKcn8o3pvz+NRTK3NpWqqQ9eHlCMXAzk0uKlgaH+MRQrKny0pDrX7qyzL
5dZReLxz120JcUKp5E8mXkYlBfH/5IjeGbSaR4ShHc4fm53YAjLpILCVyRakoteb
mIdD02xd7E+size04I5EqWKDxvLj6SCwZTDxr2B8YnlWUpXDogI4PliOelLWA0Rq
JWBjQbsKJmd8JbaSBCVGj7V/vOasiqqWR1JD2mlPmAVwMYahry5nxZDlKsXRlkyY
gROKxawB4v+fRwobl/ayH8YDHj/zrmi9itWBcApx5ZjxzrTTYrCQoJze2Z9rvrPd
OORWHyQ2glLHNaqEVyRhgPdQ6p3Pibey0UqFBab8yhAvzQbW/MDfqHx7G6Ej4Uey
NtCZSM97HSRpTSV/xPUeTKhsSzyIQyhk/SyV3zvYqvEpfb80uuQVXPbhky8fBZWf
ACKjUgIH0v0Iio1mdIRN6P7M6Uhti+2XhtnyDdjXuN/yMcu5/Hx9WIsSJ6BEpprE
WBxdPjD2ZZj63sx1rv3ZRXOQyEBNW86deXwGAydVXXlUWJ31BGXWOFxSGQL/shqa
KzvAb36PfYQICqci8J/y3YXzljgZRtvjFzPHby3z72gDOUUkGd/Ia3SOJno+Ep+w
6gl1dLBMWR6wfQwAWpnrUTxQ/IiAAm4EzS4RDSROTWgnvks4PRjRUtbSQgiGQ/jC
79gS2+/E34tO8I9/nyPMC4YgWWW3OuYmDwNEvtd8ieSOZNxcDYUQccOU4umIIKvK
ArN9m/LpPCAPXiI3fxEctChi0+CwxCff3nrukAOjRNJun/Wwre+Rbkcke/Z38oGa
89vH1cJHT4UCNpFXqvROaSBY3quEgZPajRIlFA8mz94g0Wji8Snct4BqNSbw0mEr
OQjdA1Eoyi4uJyJW3JfpfirdIphhHFhcfHEUrMTx0mUzTc4AZdghYC7VxM369/RK
otg+cxbK30Q2cffPC9m97F/uB6tIIyFGX4etCG669LdamBi5FWH0oagb05PbED93
JSCCLYom8wsfdNT9C4JBM18ExjLqOFuuGYIoobgcqfp9NfXRvdOrBXesPFGW7401
XU/Y9yprTLSKxRgPd0C987O/DG7ZSiwxC6bJnzCsK6vuZm65xfZG5o8EGOMn2che
aHQQ97T5rRkGEtZokoV+KtuUxAVlY1Dkka7sRy5uT+0W/+CwAyMYO3poLjOobk8o
qgXduWkOkZMb/v5N4x/dbnSDL6BVRqQ04+q8zetkBu6UPABddDBm5Re+uX5qZ3XP
mETAoqiwPPe4VlMIpO1t2r1l2r8V+BArOmR/SX80osp45a+EUcdRd9DLNZN/ZLwb
kmh3ZvNupa9ymXZHUEM/gsRfhpDMsfqppcVorxeIqYuKVplkuzqfeGNbxV10JgFX
zaSGy2rKKjmYHhBdx37OdyoKvH+naZm2GBxaqaVdUnGmYaSJb0qJpmgK9to1t7U1
dJUX1EG/d3llHlkBhnGP8mDjFqR0Q40/bDk+ff5+tvR7LhjtbOowUwOqTKFRSAsX
Qu7UJ/P43WNZ/pyy6Pi3d4LJ18c5KFZz+D5yd5NhnYEyF3S4KT/mDD9w7soCTKvf
OW8mRmPJVf8E8VtNVnZ9fB9nSpk6rhfKM4hHzXPYyK8go2/961WNziilE1EqC9mS
cQbNbNnWh8ndpVpIZeUOo1CIjyCeOaOlaeYXI+/yGWK074La3ffFp7PwIC1pl/mZ
z2Z1YrpVqFFaCl41DB8gry9C1ucooC9O91eB2i4iJz5jTQSd+TrL75KKo1JqBHk3
LucXN27ZJgJAshKqzdUHTKk4DlSOlIkl5mSmjlJJCn7AX0YHwc/Bp6Hk/16TLVLt
0eniBDiz/a1Y84n5vmpglVJ9Pv7y6Kzqe3XaR6wrZ9k2x0yQ4u/Fl1uMb58kH06U
3Z2Qzf4ctdedVDypqp91/igRQymTqvQ/btNtb+aRSy9T5oCyi6Iz4XYOBxlXd/Xr
F9QUCVJp8+FGeKyBSxixBz+ozMwzr/VMlrRQLhM54RLvdQEfKrcCFB6fFRfMrf/Q
Zph+p4rs8V//lj97Ej6LTafUA4zyEuJ5h9ro/mX/JV7Dgoqwxkk2L4iliin947/R
Er2LAN/5cqFzjW3OKc4PEYE0h7hH95TPgn1LCgBQ3aN7GJGCeNP842Mr68v3aH9J
6syhlJ6hTF769FyBvCTWcb3rTyK6BaLAuwDEgqmqZoaNOFdvxvBQICfpTRA6x9W8
VBhK5To8rD5aL2xTZ7gYfQ02so2dHAVooe5Bk96J4h0PqUhxsaO/PINNF/min1VI
7076Cz4pXkBWRGEQo6hdQSzV4/5DZY2S7KyXedYBzVudHmPvtstbVvNL2EXdPC/E
PKzLq6KY4SlLWyzA08yeOOAzROtIbpe8pmZrZxZ0cfYSnp9ES7mQ2nXn+5mHeydG
2sNVELmS5sqCD0R+6ZHAwi4CnVvCdkF95m7XXj9v/HRW3N/GwCj+yT3OXt2v+nx9
VTwk5o8Es5L4VDpCBkz9e3UWfEfaRyR/JjJBn3AX2by2csZSS/HJnTTchVV//zK5
dx0SQXLioeP3W7XEUrqbaUGzffiIh2bWdq+dLhpGAvJWGrOa7Ekq/zqFUXIRw5GF
G4MB4yqXmQ6fGfvnNHQImyHtOyHcJmjrc60lKk5U1vZx29SndS1Ofq4vj3xim48+
BpLYxV80vuV3aOsuO/VSgQ==
`pragma protect end_protected
