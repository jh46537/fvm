��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�����:��=3�J�r	=�� M@Q �:���!+��?kC6U�T/���&��	�bK����V��D�Db������V��yfʀIG�D�Cs㠆�.�`OI"��\��L'1dA_���%��:��c���'P���G��4BS�_VW�#�6����ZT�v�O�! Q1�fX�<o��3���x4��̢�!i}���IZ���C} ���ӣ��L�l�,��Z���#)GO2��ׁ0 ���_y��7�����m��n��tGo$�=x:�U���������3�YX�"}�ۋF1�0� �-3��{^Yt_-����W1�>_��M�-�����������&9�^�?�ʄ�BϦ�s�V�gW��ĉ�Y@B��9`wg������t�I���Y�<���A�T�L�Z5p�C3Y���D��N<�;�n6��y��S�s�ok��P�����������i~��()�8��Q��B�a��ٳă����T�4H�\�dRn�voj��~tO4G=��-���*~獷Ϡ�oisʽP�� �mGE�˰��=�s�e�/��yK��\������]�s=!d�-�IeQ�eY�u�d}D(�!M�C�Q�e�f�Fs���)���װ�s��Y&PXJ�#8[DI�	s�YN���\���ӣ]�>�ͮ�sFM�Ѫ����J��A�����&���i��(���R)Us��IӬ5�w��B��D}�m��4�-�|f�L���W]����" ���kY�'dcl[�f|W6k�	��B�(��%x��v�(�/�^%f��}�5b�bC�I�t�i�ւo<��h���O�a�A���>���[S��Ym�Dy��%�LM
-��!L�1��Du�/���X�Oi�� Nk��ݥ&���K�\�娧��؁��Ds����px���>�P�w�x��u�r�zVT\����JE�Ų.�G����G�����7dA�ŗ�5��Z[��]��"eR��j):��!�2�N�A�waO&�羛hT4i�����x���	�-O��م E�����AG!�z��Y��5�"�Bŉ]�,��>�~�۰�c
=��c�ajOyr,%䌪�r����A�d���8&��47��L]EѢ�o����F�ِ;��H��?"�+/��+e!EWng��5z4��໎ a�����̸�k=;���O���o���Z�|DS�5�F�sk�R��}���Bs�#q%�ѻ�J�߬�j���d�{�.->Ω�P^����B|$
��1
��tk`�d�K,��/���nAL���Ө��R���(������x��B�\Oz8u�)��'�ѻ9��s�M'�Fb���`��_j��Z��f�!Lb��Ӭ^�~El�ߴ,v�Ob}G)W�?��s�VX�(ԭO�%��ex��N_��u�͙��*�I���4ϝ��4��?�BXI0��d��a��-��`h8�삏��o;`�`�g>'���,:�;u��z��ƫ���+�Y�҉]d��nA�ǃ2V\0�ST|�!�e����=0�r�HF��W��|H�Wլ3��i��8���U:�q��a�k��?+D.�3./3�y�F��!�)�]�S������y�S����)�r/�
�h������.7X��g����G���4��qQ�Y�3��(m�1)������I��*W~F�k.�19��w�R�&���(*�h�ן�������{�a�.+$��6hT�ך�����{�+_�[��gf�M=��`�gJ�̂R���o<���{q�Չ4���r�Z ]��\:y�f�����F\,tL�i:�/�D!0�y�WD�-������NE�>��K�k�/����j�V	Z|7�) ���pW�^N�c8���PU!O�a���9,6F`��p�!�bu��h�f�|������/�x��~�����ʁ7�D���P�Z���=����%_ptk� �=�@�XzF�#9��6a���ۓ�,$q���>$!��˸%���� y�>M5�|�*�g#+�md6L�oy�)l����_�*�4��P�rO��ߌ|��af?o`)��>_"����^�:9���p<��V����T�k�,���|�Ŀ����~I�:k!�&"� xѪ�_^E�=@_�q]ǜ!����͝C���ʳ�W����6s�o�2��Y��;m }u�(u�B^!}UX�	A��?}��[T�b����uι�x(���$c?�������\:�XJ���>]�4+Ho\&��8���';gn*��U�t))���>���Iz�%t�H�͆�}�	����u�yo��+*t�u$C�]w����z���	�SK	\��[�0P�t�=��i�Ŋ[�+�!g�j�pN�+���TZ{�iv5��WS��Wb������c�� #I'�u
7�	���Y=���,��;��V�l����0Q�w�s��@wiF���l��3ik+�X�60S��@s�����z���.�����8u�{��,����j�x�g�w'��\P,��+�%�s�G�H�/ �YJ^��D����b8�|�Y�טQު~�Ew��5������+��W7͒����T�So����<51��76C�)T�����M�����j3�f�TF�X�r�ׅDScu�R�fλ�H)ʽT�� �Q	XX����:����6<n�1���q.�+�	��,��Λ�0�Z���h|@�B٘�.�K�A�}ϊޤ���ԧp(�!r�z�6�i]a�S@��(��	�x���W-]��Q�6n9��v�q�Y33�i� b�hS[���u!�~&�A�5y�ԡ�c�b�ܼn�E>|��Aj_x?Ђȗ�� <�5EN&~ZMz�������$5u��^��l�k&�%��K��8��%� ��9��+>�+��jZ�.j��G�;��P��rTK'��vk���W�ܰ&'��q���'ξ�����5��L����'�.!fK��?I8���AV�K�]�Vhk�����H����oi+�a5���Zdȋ�c���Y��/�����zgz��TG��Q`P��{TE�*M���w�b��X��m\�WuÉ���M"��X�[�S�^�Z?P8��݅~ ���U&�1�0���TVZ���Wo����_����>xK�p��o�8��t�{�l�����O���{����ڧ��b����N��A,�ΛL�Mл�-MgҞ��� �DΎ$�!�(Z��nޭc�m5NUB��ɷ@�q����5�������1iK�6�.�\����a�.�x�x������:8T�	��� q��	ԓ���
[ B%}!#���6������3Bҷ}!W/W��i5NGG�&�]��l
���q�2�o
��Z ����z��H��˪�s��874G���V��S���I&���y�А23��R���ꖈ�sFּ� 3�5�
dÄ)'���ov,�LL�1�T�zn�ǔZ�Y('���`!����-Qd�\W3����?$>�ݳ@$2,!a�)V)LX����H�9	9�2>#=b7�`J�r���pװ"���^���h�� n���W^��������?�"bR�RhB�&M�B0����3��fG�HP�{�	�$1݄V��܃��A�q�cI�"*�ˍ����e����I��{u"�*/E����R�h��=[��ŉ�b"��^n�K�+��)@%5��5���<��k�>���"���C|Uh�l����}�O��4�@`b�(�4��̐�خ��D���+����!��g��Wt�o��dnr�����2{Z<IԠ�GV;r�]����ːoqr���$L_��tu�R.�]]����ڏ��q`��ӟ��cl�c��#��x����9ژ8���kPe�r`������/���l�E����<\X��^(��q�U���i)��O-+2no�����Kf�|��s�`$�U�j&��./��?����������VU�H�v�~9g�k���l0��0��-8��(p T�y��`�$�T\d��cn�z��@!�]��$%e#g9���Z�f�����ڣQ��]_�RO�U����
Q֓-�*NF
�+���bЏu�\�R��QD8�\i
�K\�u�n��^�<��&���⚝�aJ�T��h)��J��$���/�,��K�uKY�c~'�e�"(� ���l+��Bx@%��ى���BU���I�b^���o�\�,�F���ݜTh̨��������?�
ex�u��J�N����찖f�*�slS�+�Ɓ��EE�~*~+q-�N�Ȭ�j	GǷ�GU���5�_�2�'��?'X��	x[���=֟�/��F��AƐ�IT;�4�\1p�Kx���K����6���}����1Zet@�� j��ɜ�b�L�";�pdƛ�(X�	K�
�1��5�-��0<�h�ԤD/c JŊ�.����C;|*�k��ڨ$��LǮ�����	��8�:�`�\�Yyz���Wv�P��f
?��)��ߡ�
�(�U�B�n_��G_b5i�l+��H���w�**9�֑��q��0o"��WnA�̱��(����AQ@�ڳ$4��J��! KGbp�4����)q���)Y�<�	�9��~�w���!���uf�g.�I'JN��CWa���r�Ό{@�q�@�?g �0??�Lh����+3BQ�G�3Ҩ��p�`h��XT��S��k�P�(����^�z���^~�D+l���^�$R����y��E������6��&o�6.��V�l`�����'9�Iޟ�	Rޙ;+�sER���B4�К3�Iq�Z�*j��ڳ���VT�_��'�
W��^ ��Xc��_4�+�{���~kƟ-(��R|��<�- ���HA��.�j���F��@P+�m0��t>y��7�ؒI�z��	A"��ݼ���̉����<��Z���m��/bND*э�u,$��6�t��=-�J�̻��g�J�b㚊w�C?��,���W&+�����H�ߡ��������Ĭ�]�K1ثɈp
�xh��(�E+���`qr ll��@i]�-؛?�7$�,��F��?UO@;�2��t_$�d;�\���|m|t�4=ŋ|�@�h�d.u>W�H �&\W�:��]u������H��t�����M��ovYȰxDlS.k�՝������z^����֟ݓs�\��ԗ:ov��my�ſ�"ț�������W[q�7�}���tD:����A�z�]�{�9��G�7���G���k��!f-�H&��~qU<�eu�,G���otb���Ϟl�s��x<E�;;��ݶiޞ�)��v�}���[�9�3\��g")'\~�I
�i僓�h�h��$Mn�e�).�TPf��ߠ��~�<��Lz��\9w{%-'��"W��	m��&#x�
D�D��z�����/6��n%�q-ʲ���/�5I��K?q�ǭ�2��u���+4�@�n��xXwD;a�Ӵw?��[�\oC{0F^�-&Dqqi�gJ?�@K'�xO����i�*Y{�?���f��0�[����*dt�d��Qlq1���<D���W��;Y��}�k
x��ɧ�AF�؅!
���O�P���z���ף��	�5���1!+y��Tr�=�W2��v�c5�_ɉ����6k�}��|��\(�n̨�eJe�lD�#^%�"9�d!a�vV��rEL�X�,���W@*�\?.��6������+(���g6c�f�c����w��ɻ�����s��(���d�:��������,�WR��Ҟ�*�E[
n�V��@��N�,>�K���A�K�����m�KX��8jn}���^`�@��,/��h�fYE�s�)|RAT�e-9��/E��vt����u؛����&��S�B�A��N6�Iʐ����Y|�r��~��z?���+����U�#$1v�dȍ��~�8����߆�{G�U`;�r��%���V����\;�j����*��s�/[_�� (���`$�)(1�M�t�:4$>�~��9o'O�u�֠��~���{0D�z�������,tpТe� ��4%0�cL�z��d�|9�C #ڎ�����!�:
�Q x� �f]�dO��~
�?�:����x		-���w��a!h�1<��B�6�F����㯂�� i��ߓ^9�4\��/M���Ns�/8�N���&�7%��%�w\�3�֍@�=�E�yL�4n2�`�z�����^�?Y�mpyin��ûP�"���G�-*�Ҁ��<�w�^��^�[�$�z5(��w�
@�L�/�0��C��1��r��wB�5�� w�K︌�$�;���J�
���t�M�v�4�&R�+qd��q4���Nul{M�I� �V)�I�����ܟԫ�"Ш�Z��"�7���π5R��vY�*uVk���p�x�'6�&�9��]��Y[d&��(�N.5�{ʟ�F!�w��cn%�\5~�9�$�7�w|�W�?G٥�L��g�%��f��M���(0���^0�j�H(���mV8�?��Y�FD}ݥ?J��-4a�=�lA�R�G���쬨����	�L�}r!�%H|Ϗ|�f���Y�i���^�oAs`���������!�0m躞1�q덄]ă�z2S`F�g�#�W�i�jE�T&��(�uI$�츫f,�K��M(�50
&8F�_�ӳy���C���qr��:�^� E砵c�eV������)C�P�(�hUf��JA G@Hi��t]�����e�9Y�pBl��UE��yte�����v�L._��U&�x��+��C���^����H�+;�X4��HN$ 5�6 �ߢ	�ļ��O]�� ����@����~�v���.<��cݜ����Z۴[�y����CJ��[�8�០��>j�eU| ����8���l��S�D�� Ŵ��` ��4�[)qF��͑�V��r�o��
��	�+)a^۩H���H�#�ˀ D�g!D��Į���%�@�jͳ��2�A�XHO���5���j	ݚdn'����jӳ4���4$�2To���>��p�4�����t�J�P\�"��)0��w���4�� ��{I�z��o�!��p�CL|פ�B�EfQEۛ����Y˒�g��<�Gn��u�1B�gT�n7�dw<?G^�%�P��X
<f{I��筸~e��GɰLA7���׺�G���B�i��🜌&�CS�L�O<��k�#,���nf)gW�y�O#=ٞ+I�E���
��6vޓ*�Z�dÔ$��#�9e��/�-�Ey�2)
���,���M�.�B1Hw,�z�RE4�����e�,�����>��'8±�2�=V�X�[��΂�u&hjR%��Q#,���XN��}�i>���*Br-y卭s9���"!��Z?X����3 k�O�ݙ�Z�-Ք�Й����	�5�l��>��f� �Fdܣ�e(+�*oW6�\e�� ����('q�m���8�
�s�%:V�G�^;�p<y�6�ܗ�E>��J��g����-7"���*/�=�)w�#����s���?�͝��\�kg���2û��Ξ�W������6�V> �X䨢j#���T���
��lGSH�;��`yO, ��9"Z��*���7p�z��	���+��z���-������1�f�!�lN}M\�O�8����g�PC��Kd�Wۆ������_O��2�<Sg��A�M�YX���+\R!�7/�VMr[��6\�PH��`��>�3ܬv�ѾJ��N�[����r�>.~0�2�*��Di����-���hM#� V wES���ℑe�큏%�	L�8��Ed�(�י�r���9�"a]H~�i��&�G�'FZC:$K�N.�Jk.Xw�oo��K=�xU�Qh�ݤ��m�w?t¡�3 �nk{N�au�j'*"Vnb�!�R@�x��F�t #_��4O���
�.�.<�P���r����r��ş���CN���2c锱@��� փ)��L0E%m9���/L�W�����&����~e���rC5"\�3
^����`�&��lF ��-���$D?�j����_c�ދ��<)䎣>c)L�2eR�hh���D���p�c����/��`{@ɸD�jZ�@�T=����*E�9�����1��я�$0�^�f��p[�kTv�&�xnEFA�<y��ƃt����Xy���8���=�[[��l����3dt}���~�m��i�l<,�w��?���9��z|cv!?���t!�0�e��#���)<X�j6~3<�C v ���B�F|k1M�6R9�A�̦Z�s)1�i���"��$VS��YA�����Vbcޕf%��id��o��	s7+��r���m9�b���gm�[ ^��D��Z8������%7�+��J����$)\�@��"`�s.א�4�	��K(�$�L��ᢐ�7l�V�z��b����P�N���#x}ʅߛ�xIp��L��cΡ���΁x��$�'#H����a&b�7/� ��3tn��FW�D���km:����)�!�3�ky吖�󦓖�Ʀ�$s���F˺���G�1�Jp3�Rgֻ,���B4'��^6�;���i7.R,��+D�j��4GXP�|r�ig�F�M6ZzD���hl�*Q&�\b)�S �>�Ka�il��7��h?��w��	����0��٭�I�޼ou}����ў����Q��ۚa������h�W�,-��څ�X:��1xu�b�ćX���@��U�� ���<џ�{U, �?�P�r�I��+$P˟��#��|������c&�pF� e椝]���fpǄX�5��Q/��V�U�.�pV+�rػ
 ,�w���B7Rݙ˧���ѹK�&7�F}�[����?��$����'�lK:Q��h^M��8�P���JSSjOYFG}�+Ce_;ڇ�ڕ��~c����L����E9X��'m��0}>2}T��yF�cH֖jn:��ϲ�۲����Y�t�T�&�a���|����,�x�
Z�S�hwpc����3X!�o���H��eC�Sl��}$�PHow�.|mx�5��A��J9��Ұv�4���w��Gx�`Ot�#��B a����b�w<؁�Yu�ߦr��SU�'-ζ���+|�y3Û����c������TTs��1:�U9B�����`�H6�x:�{�����ջFv���1�@OM�*��@Y�ۺ@ǣ���L/����." �~v��ΥK$�3 �6�ٷ�U��ԔN����П�O��MU1^�.2���էC��'sRji��ֽ��
���A�]��G �����e��K�P'��x;,�ي��Q���Z]~`��$��0�j�`E�S
��~����T�*�o�#'������T��L:�Xh�k*�D�>���.j���8b+m�Ä?�a�ۍr��c�4
@%�{�'�S�s�8�$eT����T����A��HP����\`�����a�B���l+S��a�����:��5H��V$%釃�e`�=�$��ީJn�[��]��	��������I�;ਚ�"P�A� �w5�㏻��@R32�2��߮����-f�G�_���؜U���Jc�඄��QC��|�cF��ؙB���������}w���=��k�]��C	x��������?b�R�L#����7�&�6-�3CY�W��6�[ޭw�ܢ��Y��'��^4y�GT�j�on������:F��V|.'xz�?�~����FJ�H*c��-Pα-`��W�n����ّ���q%��ۡ��y]�����D;�87ͬ����l��ӗ`��Rpd�Dܦ�n�
5G"]?R��l���.�{x��i+�V�wqt����Ŀ���������J��"�R�8�@��DTr�^��}�fl�{�8'�'�۲�\{[~8���_���+��kn���|��p�a��~�~�v���½,�"���J�
~�m��=��I���e�T�;���F1̑�]�E���ڽ���QSѴ�%�+��'_Kg&����H��G���p����ٮL�f��|�@p��92��?#��{ؠ�s��RiBz^^��*N� L$
��Ω@�DJ�3X��eO��Ϭ�⤌����n����r#
�������),�^��3hۢ�S5 ���61�Y^a>6c_�����Q1~[4&4���V���D�:��5ai���)_7g�NI����yB�4aڛe6Y�?{?'�w���,*:�R&�&��uc4&�Cy�X�jf<��
�J6`M����.�3(��Pkg!8F�O&E�@ڑ��G'K"]E����䑨��^O��9_��Z��Q��oǪ���Ѐ}�lu}��u �A�9x"k�!�Xi��p�R�?�p��B`�8s��%��PTT40��\�	����/=�/*���ft��?&i�#����Z�C�&Ckp���W�?w�䗿8H��R5co����]1�F��慘��5�$T�����K�ga����$,�_�	4�c'��"�.ޕ�L`R�N� 0h����_h�����ѷ  jp�NX��G٫̀w�1�����{�Q�}p~���P�C_���d���k#y~��S��6, �h�fj($�O�s�h�ARD���,F��<�d��`g>|B��xt����'1ŢO P����<
]!(�C8o��@� �|ެj6����*�;������Q�`$�����=#�y���E@��g��05��A{KlӱS��D��p3v�	޾|c���+8�2�A�������ەca�fx\�rW?Y�m�����oI$R�\½��1�Ҩ��7EmF��=�u�&���5�K��ť���1���WV�$�j�պ������O ld��\�WW '�
������y�#�`�ƺ��OD�@�ȼ9|� �1�N�*ڈ9�嶦g����2~�EXF�G<n���_t���k�a��N^]Z�ߥ�(����} Sǳ���i�>d��N$c .�����߄_��p �2���ޑn�Bn���G�p�O5�C{1�-:�<���W1�����ܔXiP/��H�s8y�*�������bֱ���]�@J,��f�÷��
����U]�c��J@k�ܦ�����ɤ�U�u^��xV5^�z��^���7���E�o�,ʺF�~��rO'_#/�Ӯ�5S#�*В���@�۵���ke����I���x��k�O��.C����j ���-jE��gI���!��/�'�o��1{D���aUI�`3��'&�ȥ�d��B�f�erdU����<\ xQ��W��&;S�=
�� :9���hR�
�Ȱ��V�y�3�2���u�pX�3�{�\KU����Sa��x�6��a�>�#p��������λ"��d�M��BI�!8Fc��s�o"����΂E�;������**�?$z��
"v+�Qg�4WJGj��D9�W~�(k���i�x���>�B�PAC�����«�T�+�r�)����s�E�+x�Z_I,�q��M���6����<.ի�%�_��q���v\K`Yp�yz)t2��l�6W4��˯�:�[�#T��[1�y�$ԇ��\苫�Jf���5%�SnV��ȝd�o�!��<E1��R�RN���"�D�t�#)&��^=*K�Iג�%���s����D�r�:��6�/W�!ڥV�sC	�U3I�d�R64{��`�l���ިd��g�0^�1�b��mia�t�K��G8Q�p4��;���7�h4
�V|R��`�7
#E��쳿&����ɝ�g�MW��"�ˁ}�7鳠qv~n���c��X�	��@�I�7\���Rϰ	��D$w��`�.�5�i'Y��������xE;�cɊy�6F�Heq.���_5B�y�1[]	���F!�)%R9����x^z�@�~n/Ϧ�)�(�� 8�z<�+��
=��z;p��8���z��U�������X������NXwD�Fk��kP d�?j7z�����b�z!��/�'���N���H_}���z=�=q^�4��"U�
"iy8�J���ann�P�L�ĥ&I������KƄ~��r�X�7^Ƙ�3?nZ����L՘��ӵx��q�v�|�2�c������}�F���N���B���^O\���:3���'>����RB%�;P��?�������e j�x����h9��s��&,�s��8U?�-�$�H���&̃L]b��2r����b���e��n�ŢY)|vd���H���MK����2hU��o (����N��>Fĵ���ϳ#����
.{����2h �{�7�?��zG!�t��%��7t��J(���\	i��:/�k)��1�
�t;���tQ���u�����`�Ū3[���݀���<n��sKc�q��^�
��I���;,�,(�x�q
���Դ�f{f���c�~X�Z�����r���)�G"z�tϯ$,}��nGc)��OX�b�g�����$�lݤ���`Ǔ��K���6���K�W�}�s�(��A)��x�1+�����K�&@Z]j"	�8���]+Ӳ��ĻH/�r���Wښ� �(�WZ�������֓�
��si��l4G3[����������Pe�S����#Fl7$<�C��p����z)&Fn��6����w���2�N'j0�/�Yc���z�YŭI��-��8��*[�V�ˏ��H�
�ⷀU6�K�A����Y�!wo��D�Xxz�@��y�&�� ��!]���Z�Q�~G��w�R�����	C����X�k�'�-@���{no~���������6�	OG8>j_�t^)d&>+���ԟ��7y@+452� +� L�\��'<̡�AJ��P����c���W`يϳ=Yc�G�
��\�"������D�Δ0��(��F�	G���6�Z�k��ҔX�W��AH^����p	�qi�>囊.�C��o�4d��
ն6��H�;D���ca�8�Cu7nn�3�	�Ƚ�R|x��8w�Q�)���shЏ���
PY�XH��Ij� �w�2z�