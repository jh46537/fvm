��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B� �⡐*��D�k�(ʸ;+.~/jը6���1�@�P.kZ��笩� �hC�צ�'� �.��%�x�WOL�^p^��L���Iv�shI ��>�{5u�����9!cDn^D�9�b�mp�r�|~f�l��j�5��od95�� б��P�a�f��>�l'�w?5!^il@^+�>L�a��*r��w�Ś�М�0�P�c�͏�B:�I$ZtE�Cd�T<�	!3JCǮ�8Գ�1��t��>o�<��������vY�s��R 諚�̪T����fo���)�a6��l�Y�A���toq8�rݢ�$:+�~�P��# ����dAe/���A��ӳf���|�K�F�!ϵC@w؊��)��ZG����Ǣ[M�iS���Er�S�����§md���k�sR��C�����u��촒�7%&�	�uD+Y�h�|�b>1��:�:��',d���g�~4jY�'�ڨ��5��@z����y�˽������/�'�Sո	<+	S��c[W��Ev�vU�0��.���ėX����U-�O�{�q1��|	"b�U��pUz��He6����Vlv\zq[� aA~��W�QF�5SK����v�_¸�����I�A�����ce����}%f�,㷉�ȟ�C��h>㼷�I
��7�)�e ��'(7�
\Pc����N���S����$�����6 �\��E�Jc�i>ԓ+���!k�l��r��Y�� ���4�ҩg�I��<�DO�z�B���B���i3b�}�׈�5�qd�B��Ъ�M?�����P��0c��(9���)?�\ho,�.ִ>��8<��7I����u�17�JB6BiUG�Xݷt+��s-���)��W���b��<�9B�(��T˥54m��
3q�ޖ�Lw��5$T���#6�j�hM�Q�����=6)3иE�;�"�@n1圈�%TI�;�S6�:`D���|�C��z�IVD�<G��W9���f��>��^�}�v�7H*�|�I�L֋i~8��5��
��W/T�w���|N�6��M��P��'e�;|��߳]��\��D匂O��w�2�.?�f&�-�<8�_bb�r��w�^�����lbub���l|}�<<�b�!��!�0�|6��������z]<|�'�|)0Xޢ���xb��e|�S���J�%_̂�]�3��l��0\ZΧ<�E�!'ZT���D$jw�x�a�����!�eM [��/���u�5_ؽ/�"%��`O�֖ʘ��o�,J[��$���N����>��Yף�}_��s�Ն�����j�5��6"�U�KXD��C�RP���p�Ę7`��zK���>���\�,(�U�^�(�a�l(	��Q;�{�o?C 6������$."��&=s�}�$o�}�XL�Pׇ/���AP�V34��vQ&	i�1z-�6d?`ZG�~�ƫOC�C	���Q1�p�h�1�}���%�SB0�����ʥ�K���Tk�b#�2>����*B�'G�`$3�{I!Ǘ�{`�݇2C�lM�����fN�˵��uC�J�Z��[WGJ�Y�IP�;��`�,,��L�M��n��	^V���P�e,�g�\��փ�LL?(�[�/�_7{�(+'�][����O�줌oDx�xwj+ g^��;��F�"l�_��K�Н:<q�e��O�F�v+������_����(��<}�R��ݕV�:�g�Ao_�~U�d "i�1nղB��~��n�aiΓ��`��Oڅ�ivpUd�y��Ԭm`���D��~eÕ�C�j�F�mDU�܉/ {~5�1�gyj�v�޹2@IR�_2k�U��c�q}���*��� '��?j0|<�"J�YWzZ�G���`v'�TBe��X���uN2�vR��=���b�xLW���eؚ��0�]"I�D�L_�̗��v$e��~}��n£|\�m�u��Ȼ�^Z���w��T�t$��������g�;�u��N�#�w�L�!�+���4e.��J����S�:��E)'���k0�&2�s���=#��F*R�Rp�b�՜\C?40Ԭf;��9�C/
+�j� k4��[VK��^�$:��Z��'*)�?�������.�� �G�������J��X��N!�Gl��6;���u�
�pv�lq�&�����XB�{ QC��S�iY��
�^��������h����N[��WM���B������ڒ�A���L����m�,���`C���P�مg31�ւ.�!]wJ������M{"d�s}��j�ߡf�Z�J_��˿7��Y@�R���ʪ|�w�:����DeXy������+w3�Ɋ���r\z��4U�󺒲�u{Տ�<��m�b�{�dԊb!��J��ۄ�GE��:�E�sX�ZM3�ؼ��XJ��u,��SG�X#�O/=i�qT������ǂ�i����/�ߓEE.�ge�۰٥���ﮕO�;:c}WQP^^1���8���<�$�σE��c)��%84�A9l���'�9�I�E��Mmft,���0]t 9�nO2h#�Y)c嚳�eNQ�Q��y��j�l�p�P�2����]m�G��gUC�"�d2��vʵ�����^���J��!Nx]:/�F�5���r����7kPwzDL�b+u�[�cg���+�i�ч~����x�1�Ȱ=Ǽ.0W�X��D�}����`7*�ef��T�L�_L��d���.+'��S`�-X~S�G��;t	YKzM[�V+Y�j���k�<#�g�#+˜��.olO}O߅�j����i�**C���b�WE$�)�w�i&T��c���W?F�htC
�2����¦5q����� pD��s�/��{͛����Z8�_`��TVW
Fj�B+���/����Tq~gQ!�t;MU2�Ll��}��0K�!R^L3C��B������k�A�oFk#����u�l��5�m,��I�g��Ѓ�"�T���t��=ז�seX~��U� @c���\t5T���b=E '	b�^P��NV�b��M]7���� �����6����$e=`v�+�l^��z}��e�Y�j��@��zƗ=��wx�[-l2e��;cǚo|��.V�5fa����Um�9��N�GD9�"7$h�aL��-�R�ȟ���w�LI5ԟ�NV	"l���$� ��U8���1�[X�eiH��Hl���		�A2�j11���"f�?����0�Z��|�z�ar:)ĵ�hQ�B�q�a>��DO�,#�
ær�\�aWn�O0'�\p����C�F��-
I�|5mH���Q��Z?�ħK�� S�_3}��Kummq��[�7u���F�ҡS^L��?�^��6�4�%�:�8������p��bZ�2�U �׵�7��Q�~�l�~��v�ckV �%U=�7В��HLm��:�a�z���l�/�5�Ηޘ��z�8�FB�� �����,^W�&�1��>Ά��un�0]F����&�,�7�%gB�N���-n23�����Z�S8]��c�F�����V���3�~q+tq�S-�/���DVC����l��c�d�����DW�f����5����HE��r'���nB1WY�|��I�i�]3"B�C|���O(Q�����"�:��ŕ��u����?�{>���:�� ���`���l]y�N�>����4���J�]�x�8fڏa���5���| �����X����O~���7�+�V��N&�D��ѫE��8�{��H{�iQZ����YΛ�� �a����Rj�9�~s!1�qG��>��|�>NkZ<oc2��u�W%oX��`<�����j�.��t��	�z���I���N�{:������9.�a�]� �uSc�eM��P�*�R����یm��>Z�Y�A[�Q:�����o�H�bU!cֿ�H"s�q���daVtW��ALw��Ϛ+*3z��Qז�-�AI��n4)$�a?�&�q��ү>�e�|·�A�ڊ��3�7�=�����>c0T��.j�a)o�����+�����/��Z�Ǌ�!a��}׼g$Y �7���R��s�~�R\�c����pW�`�i2�r��e�8�5��.P'�$�!��J �ɵ�+�wLs�]G���x<��<tb�NK���e'e��� �VRAa�g��8����"�	(.�����9ݠ��wT�����t�1��sJW��e����! �ڵ9АOY�>k��a� ��*%<'i>ƘO�q3�5s�L1:���W�hƋ����f�:�n���)J,�' l	h
!��m���eZ�"Ե�`��p����Q�LŢ{O޷���<�Co2��kB,��"��������u_镅�JҖ{��Ժ� a�{��}��p����i��B��g��X-sx}�Z&N&��2W6K�ל�F�3�1�N~8�]��u܎�s&��	�"IԒk���&�K��5�_�ЮQ��o�o���	�h��m>����L�QT5�}���4���v���D���wD,�Y_pfè�W�P:�4{(�s���G�i�����k,�<�轨�T�$˘*�w�$�\!(�߯=�5egn^a.邊�Ӝ�KB��JOO����.~�;+�̙+eoK���8Icgg��A�	C���OH�+���R��1�n�����de|�6�}ZC����"p�J��I˗v�X����+lIO7���P��@ԯeU��|z�P���Q)1�P ���-%_�g�I��O��n�i�NC����#�ĩc�o�_�Lc9��#r��Z�2�[�Jչ�D�6qWo N��o-����|�Y�?|�z
�fR��dz�W,�Ù@ �g�p[�9��I��cM���w����9�ߥ�N&����s�tEcUW�6�k�'�[h����ˍ�T��ea����H�54���xW|	��Ez�N�����yIs�T��G>�.QC1z̽,��~���$��#���P��n�Li�3,l�R�9`�^�G��I4b�|m
{M�u�x����t�5����֟G�MS�~��ˤ-%@�MÓn=�,*9��o[��c�m��?��쫀�E{.�)^�
��Jd�;d�@��d�Z���zh$]��/wT�@L�Yވ��3o$�P]7�����底���-���`�[F 5.[a�]�������uz6�])u-4�ꇨ؁�\B�ln�&'� �*����=y��z
g�����K��oXw��uǋ\�2���	V>q�&���v��A萴ZD��0F�>;��G�{t2�m���Z�k�)T*��Y��0����a©����b��,�t�`��K�f���\vө�$K~�%��Q����>p�,����\6�s�z��7�]E:t��2��/�~0�G$�pO\:N��+]At�HϪ�Þ�h/�i�w���[���O�J�����Hil�WAU��҇ȗ�)������rF��D�@�1?=�C珗�I*>�	u�t�+`�TlEǋ��KK�8�5iP.���D�Q�8	 '7Y��k�;�yF����]�f$c��@]9_IɺE�"r�τ���[��F5�R�g��-�J�������ó�pq�Y�NS��#j28B�Ag�kedɾA�$g��=×:
�J7%��퓥�V�!j�\h� �D�5nI�$N���\^ ��e�,�����ҌK	�B)�C� � ������E���,K1T� �%<RaT	��27p�ye�=�����.W�5o�`�O