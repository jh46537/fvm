��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�{���dʂ�V(��p�s�0ZI$G,Γ0a��Ȃ��Z�G�"�#	0��=�uw�N5�y�����o���zд��`%ȭ�1�2I.�(�Z�
T	�?������G�9�sY�(I��y��e'�f�O�'�C@�p�~���,���0�`<�ɿ?>�n`��!���+�۱J�y��7��S$�lD�G$�,[)��͟��s�M��W�C�Suy�ť����;oZ��ّq�r�	�@=�9{d�g���[���H;��.������S�dm�Oh$o��\vJM|u4�0�#��xq��r9�A�R���E8�rK���e�I�:3l�E�+�岻���2�c��ߏO,X�
Lʹ.�MN\+�
h��:�t^C�`C��xG�5w���1��H"�;ZKB�L	�ILG�U�Y�׺Bn�xz�o�����MĔ�k�X<��:]$"��-�p6�ձ��?[oM���	������æ)�v�[� +��S48�TC��O��"dl^ݑ�n�$[���y۴� ��*`y���m=aω��0�2�}n��=���n��Z��r.~s��j���`��`��%f�Ѳ~ ��[�
տ��0E��;V1���(`İg�z�cg�7��L�6!vfh�/�"�3�l' �04S|0(b6����<!ǟ1�^��'6��@@ǎ��I�c��/�]�_N��L9�]L��#͙V=�H�ch�2�Y����{�q��g)P^���V��|D4{%��P���� ����I���[nݴ܇\����7�����6�6���'y��V���gA�OQ���P���8[��<~�Ja�M1���{DQ�z��fO�5I�߇���vӴ8�����X�{��k��
�!��{�R�pwx����MwK,CZ(�9����)��l��@_&n��0mSe.�E\����g7��9)f6��&��b&LR�n��5 ������BpΦ$��u�������8�ߘ��i�v��#�ۓ�_�,��"����wg^�\�� ��V�n�{%��_��[D�Оa:��5������韛�B�-����Ȅ��U�$2N<+
���ɵvz��n�bY@ԡ��~@2�})�s�?��s�H#�� �4.�l',7�DD��?��ȩ�o��'���٥o�-�}�^MZ������2��� �G`QA���i�~��#(.�����r��KVHC�c@��ח�;�BP	����(��79Uf��p�H������g�Ac�l&��s�Põ�@�z]*�q��Oc���؉�n�r�A�,üoo�3π�%��_���jC\6� N\�y�lwq�]{���?�6�H�*�;Z�.�[3���q���,fag&�Yh˙׀�h(~�����fq� IH�H�r����G�4ԠM��b��)�����p[�B�/8�_~Vɍ%�.���(� Pw�Z�Zpr/��ƽ�̐��h�9�������G�qpăh�����<@�J���1��n�0�7��W8V���X�\a�7���x��.�l#�oE2�3���eɁ�L��0���"8�0�03=�KZ�$n��{�y���GTv�;��Ԧ�4�G7��@���7,	Z��!������=_;�tM}|�?�%Z��@ c����7ɢ��`!X�~�:���*}c�	�ɣ�|a'o+�"#%g�K�J+�k�e{9�l^�5��Y��ԝ<�'��'���H��v�v�j���ZC���� �V��Xv��.h4�h6�ES� �V,\�.�p�Hm ҿ�k,!��F!`�>��]	:��nq��L���`g�c�V�j(�7{�c[El� y�,�&�Ju����R�E���KˋF��EK�'[4<5��獦��uF|-,?}Ο�Mz.a��BF��!B�7j�gjB��%B~�4��1������n�|�����E���a�7����[5s,�M�i-�@�N,{��Y�i��������/��f����Ni�[�d��k4�"����%���`^��r���A}X3��? &Auw��$��w���p��h��錒/�S�謾8�WMJ��5��t�
��k�⾷�(��WI�Y)�fN�7jX��xz/�/�d�=���H��y�d�r���7�x��*��A��R�:�Q�î~x�]����v�TmYIL1-b	�[���M�t1.��k%76�1�	���_y/S�%�{���;�J�N���8�s��켍= ��8/w��福�ݣgq[\���6O�l��be�5ٌIk�{���hr�������LE�8n�B��h���W�Z�$L^?l���x �����L��W�x���CD~:�~����jj�/�^#qB�b�_�����(N�/jgy�}Ze��r���+�2��6Oo�	}y�?.�q�Sslſ�s�hJ��)S� f���x�.��\��׬�.�->ȄTN��^����R�V�=ؘW�_�ȞIU6���2��H��MUIx��&��-A���批`� R��M<�D[����5$�H� s�^;��9y�Kƿ���^��<in���|,s�Rj�x�d�~����NM��>�y{��h2ab _Ǖވb��IP2�C��(�j/��~&��
Q2�1<�I����`*�
X|jŤ��'�E��R�*N�%�2�=�V�5d��X᜘I�d64�� j!�i�5����yX�P������x\ �� ��r�(B�A<��Ћ���O:�!ō_�A�gV~��C!�НmTp:L"iZ S*[�,f�_��lLJ�p�P�3��B����сx�\yj�]ܯ�|b�oP�pŅ��,���#�Ń�
yn5���v�ԯ1	�4kSc���{�g�8_���e�����Y���{x���O���?��AGu9�Ҭ���A�ԫ�bL�n�/��V��^�*�=�2�b���'�ݱ@X���9_��/փF~}���8��w����HvWC��O���g�.�f����ɺ�?�n��(n�}5�[)p=QQ���7q����\1ZEq(�(�) �Q�9���#�b��k��i����4�����J&X:�?x��GS:r���(�i��O�[������u�����;#�D�)v�ΰh�>JOH0��
�8�E)t`pw 
�������P͜�h��2�Ey 8��d�,�l�k�Cd���{���Ӥ�
[R��>4�9O���?�v�й�ל[�>2���Ð�=�͂����Ttd�:W�B��5g��._���\�b4�T����+��Q� ��9HB|8b����G�:�ѐ�8�1=�k�P��M�����3vzo��6Z��0|�\7��R���QA��8+��'�y��T�o�a�JZ���W�>�[�Odӊ��b���P~$��<���oPDU��2j�n&���!���H���1���J*? t���jk^[��S$gA�Nu��>%�L2�k_)r���}�@<��=���Wu�=��-�Q����W%��Nd�o���	�}ܮ��ض'�~R)���E��؄�('�>^mX�C":��go>9����h�Oj1�y����,����-;9��8 g|"��]t`Ÿ���.�ל�@�[���#��ʚJ@�����ƑO�G�)�0P-�ln�i�Á.c�2J����yk�1��#��\*ϓ/5�Z-�M*�~��",���2�U�MUz�?�i���D8݄�K󎌮`(��?��a�����~&���^=?��$��D���4��	�u�@*����t�ыi���	��+*�R��|�^�t)���TJnZ��Hd�C�`��+��G�J/�ݗ��hzϐw��hlg�����]o�����5�K�$Oq�ͥ�N��s�f�|��r�Ӄ��-Н���Zh$�&l�Jw���a�ț��y�nǶȹz =��gp&~q%T��#=L�!�BP�bEOުd�Sm d;Cc�ow�%��g��>�j�
8I��e�9��]n����̪���P9ɓ�V��K�o�6�v���¶7�sM�?�@J���x�
��R`+2@4R�v~�QYn�LM��G�^��.g���+,��ص��0��G$r �.����2�� ��u+2�XƇ0����w��m��z��{>H��G4x7S��lo�J�7q_���X;�7��M�;�TU���j��$����r��N3�F3�-�̈́�>?`�	��J'�=���Xu���YI1�'��l�ϵHAz��#�wA�6��7���E���u��PC�"WUe�5q������R�s� ��nٽR�,DZ�!�"�f�Uęx9��,"����[*�?nht���@`���:$<����JDE�ے�ϫ��0����<��N�B��*���+ ��0P�S)}��'ߌQ���=�"p\�	`K�Ƞ0p�V@�`Y���.F�*a&h+��d����(	�^��R�W�ImF�����H��ؒ�����v㨝a���n9�mq䌢�1�,��ܴE�BSAr�*Půx�{�sᰬ
U<<2*L�꿳c	�8��x���Uqr:{D_���������D=�UN^��_�Q�^v�E9q���@	x��xʣ���l���A�W�6�O�\h"����TlU��g�eU7���A�9����R@� �4���f��x��h՜�����(���^�&~��
,�9%�q�Χ�� ��an�f����- W7�i4�*.�U���ɽE�i6]��g�Y@n���$e��(�(��?���#Y��7��m�������J�/�����
H�H0g��?p�����_�(��]��t�dŬEӞҋ&#`�ς@��YshE�4�� G����<�l_��Ǭ�5��{ �Բ�6?����W�z~_>f�S����bg*����9k��ˇ�� <�w�r�4-J�T9.�9Zz-g`Y5�7E�ҳ���+O0-����xcQ*����DZS�j@y��rl[�"�$�h����:�Ӱ�r�_�`��G��M,& ��	��L\6U��S"p�+ۉE~I�7B	��