��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@���C�X�-.c~cX:�,�B�Gq8z=����?�,��5Ι+rb�4L�M�6V�D�'2�99a���e�,W�YS���|�F1�W�*��KÜ�Q��j��:�i��'����p�B������#�R�a1��3�rjR�4��|�.���y�O�,��:J=�P��Xv(��Y�]�l���q���(w����N���[�����f��3�%&����v�'5?��و.E�y�+�֠�|���7��Z`Уk��߿x�p�[d�)_��
���q*�e>{�d��5:�n>Њ�(m�������3t1��@P��1+%��s٢��#�I�-0.Bvn��D���6���}7�2�Wi�.�%��J����O)����jе:@T�?���f�| �$�HD9��^�x���Z�'FA�G2�G%�X7\��Y��֐6,�����.@�� ���1�O��,�?�T
۟N}Џrŝlh?�}w�9t���H�a�FVP�RE^:�^����f���(��Hrİ�9�F�͑�x��;��	��>d�TF���̖tR'pȠ�N��l�=T����!�(����\Ϝ�s��Gƃ��p%;h������.��������-5~��Ę�xg<
=ǋQ��]����y`I�p���ô*y��)�)��o�z=�~}Y��ڶ�5e��(�{6z����10^>Ƣho��q�nȀ�O.�-z7KFG.�u0��F�Cz��<̟�����,��C�&	z��ah?��cWH̰%E;�i]��^�y͚H,ц=zV��B�R�����Y�?�Z8���94�L�L�Ի�ؑ��B��G�L��@��U�����;P9!��[�D�gp�b�G�/`�~˃���c(�k�mk\�}�;��b<7!���U�@���z����Q]A���!���P<��h'��8�|r	|��D��SSL3�N���dn5�:唓��U��oʢU�8�&�J����݆7�B���V(��:��ϻV;��&-,B�	ЈW`�~&@?s-���8��M~�L�+3��g2�e�7��"�Q�A�3�,).,cP}�S	�Ƽ#T�8�5?(l�n���Wʰ�⁠�]��U����n��~����3�j�C�����U�D��LkG��}�}3� q+��J�]��%��2��qg��O��N��6}�����\5���+��0�F]:�0��c�FhB����^���9O�{����|��PT�m�A(-^�
��vR\�u쳷n퓓�e��sĨ.˷#H3
����S�(��#@>X��;��w�_��ࠈ���x!�����?s�]�~X_qɇ�F�~�n��ר��~�����~pX`����kyS,"i�2�OX�6�<�>�-���"�sا*H`��؎F�8�ʐ�����1��U���ۿj?����`P�瑕><,��gH�U��SzGm���M��Yī�P�һ��>��p?O]�QDr����z��ta��L ��o"���'T&�mi�x�aa�"v��I�j�h�	�յ	�ED ��� ��/Tis����$�(.�q�g(���7�Bg���*��U!���KQ4��gu8��qb̶��zK��@d<�2�w�R��w˾�p�y"'�U%�B���kDw[2e��L����q	2�dϘ:*��]m�v�ϓ<���CBڭ��pK�-F��Q������d��t����X�^���(����aH���f�8,�ΎM�/�[�I��,�^������/���� p��m�G��+���: �Ξ�����8!�PJ�6�ǝ������u<���d
�Pf�t����5k�5�)��0�	K[�^��p?2�]V�7�4l*urO4G�'���|�n�}�'U��F�#1�Y�5Kp�yA�,��p�l�W��!����5�ҍ6����P�N�"4�k�ZC=�3��:����A�}��G8�n�W	�"*$�Yh&�����]�v�#;!S�%N^�c�� ���d3��2�XK�H� |��u��=���#ԍ��P�G�Ӳ��}���A~]a�	��uV�]B]b'�y2�����t�(EuUT�[�[����Œ�3���@u|����}_nMi�y����՗ ��,���l^���n�Q�|ϗU�D�FG���V�#RI�ڔi�$x�TP�@#W�t*<4ڍ�Ssv<�>�D��AM �ͬ��-;EH�e��%�T:e�C���@�uX�3 �#��O�Y+�����=�AC�lw-�%����5��U�3\4{�+Myd�6��'|�~Ѱ� �(�Q�D�T�;�H��L<L�dn�U�Za��JF������8��͋��1��7�nl_��^(PX�M~����f��IBWVk����Lܦ��5�t���!������}F����>œ��u�;��x�v� 6� UG𨜶�A��7i���S�K��[:^5�D����;�I"]s��$t�%d�Ƀ���0�ט[���k��T(I�����'�H!��Q(����K7vT+Dk�Ćpp�#2��Ő�-$���h��w����|R'���cj�L�;fU/��+���ƩX�s����<����9:�zh'
�S�~i�X7i��V,�4���c�|zV1��S��l��\@R���C{�v<��v�f���T7Y�j�\��G6�yi��$V�r����b�v��o�g�-v�����=�