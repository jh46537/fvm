��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�~��"yAfEi�)�����B
��۩C4JA?ϋ���n����g�ҕ8[���!�܅r(�=����UG�O((�K�`�0�t�s��hP�D)�w�xJ�[K_
�ԈYJ���LݷV�2�콷iF���}Kq�I�q��h���H�i���m�����-�bH1�)��Z�ٍ�jӰtr˥V�ڥ��L���|��qѷ�&GDq��ʻ<�����n �Ꝿ��d�T�\j.+�wH^E����C�]��b��`g���[~?Ӷ/�}3�oN��ѭc�2!	�PC������B�+q�z��*����� ��z^˥���ER�J��d �-+T��o�9��h�:V�%|�]�i�E�GJ��4�G�xn�XV�Gü�g�4�a�K����ѥZ5j#��T$3�"��!��K�jt�%�8��2�Rk�h�ﾃ�!�����rm���� AX#J)�%�G4�u5ح�4���<�uxعט�=琈�bO�vk���V=Ź���Z�
�b���,hAE��Z	��Vi��rWg�M���8��R��;��~��Y��0x�(�("ǠAR��<'2���i�		]�\�H%��'En|��.'4&�ϸ �a*�Sli�+z���`t���R��Jܟ6<�F��l����x�Dg.#�|��t03ٟ��U����Ob}���F�8%�#��|S�]cNr�qWX�O׬d"z8B��w��Uӯ��xR�l��n����|����n��P�3�g���?�� ����lT�*à�Vk�)cQ�c���9���hz�姭�r_��&����y`0t	�� 	��eA��p�e}3J���<	�#�Q��"�i�'6M��Dwyi�M(`�bʨ�c����S7���T�F�t���͋��u�
����oHL�ߧ��(Ex�x�(�o=��X�Q0*D�@IM�<+�T�2s&��)������ɞE�w����>���������y�0��Ȋ{=\�$�j��:�!�u�9��,�S@V[��������0��+�&Qy�M-�:�Ə�X�����O��@E�t��xn9X��� ^�g�M�N�v��;�K`�^9*Yi3O��A�<�<]<&�}*뮥�X�˦�t0���/����"��^zہma$��S�N<d�f�m���h��t�w5��h{������	�ᚶ�p$ @4+(F���Q�A��}~�*��#�+2�z�E/9�>��N���.I���q�]�^|*�1DО�]��j��w���Q��6JƑ�?�o���E$S�#I--A+a�Hf�9�����r�w��]B��ds�����n��������G2��x]�"�wz*�1�˔�놲�D����K�%�����0א�3X�W�����X����A�r�#��)��B���6�Y�8����x�d��HXx5���+ާ�q�/�0ӫ�`9����,���Z�ߑ����ߖ�#2�wP�є�b�@��~�a����[��Q%
g�'�(�
�ۍxu�����L�,e���� PP�{bٿ�������^.P�w�-��G�L[t��R�/�n[�#�L��$A��qԺu�y2�"�|]��{����$���A"(.�k�D�zyF�c�X8�:9r�,B��y�dާC���c¦eΑ�\�´0�0�Q�ܦ�^���J�n����o�G�v;�zM_������"�&6�]�#�s�԰p��D��RT 8 ��YZ��p���_/6��D���'[��a�
��Y�+0e\zz�2��T�[�c,E;�V}�k�.vcNk�"8�EL�,�T�%88#��J�;��Z�7�\�f΁��%���0+I��C�Is�=@9+������[����Iyp$���a5��/u{1G�� ��^s*����iӒ�{��BE����ɒ�[9-1��!�q��S�)����r�b�, WD�D!��:t{����ce���:$G��a���:�PG��݉>��]��`L��%Iҫ0��#���,��m���.�h@�65��݊����ؚzp1e��)��|�شE�3�խI6��\C��DL&d�^:�.�:������m�VqAps�h������j,E?{�۸�P^=�|��x���K����t�<J�9Tc���>D��o�W�#D�QSk�K��;�S7��fJÄT"><v��:,ы#v�~���ʘ���i������_����7��X��p�3T��k��7���j���k���vgzz1��;���y�4�_\��|��[c�SU�&�S���������f�5?�p�p��́s!���
�C��u��3�
P�đ�Ѱ� �|#��a��Ѯ%�䦘
l?&�\��Ki����#`*;�o� ��:Ư@�a�_����ͧ� �{��ހ�	|T�ah�HO^{Ter3����Ͷ`�hh���z�����|�׫"0�FOg���d���v����v��O�}G\�Ӹd����k����[.4��
^��"*�����j���2�G������YG����Q���9�"G��ƀ�5�2�x����󿁯��)6�(eô���$��N������cȧ0��P����C�R�}z�K�W�][�J{�|���{�F�En�7B,Q�b�~3��������F+Bv�a���u�+�q��JO%U�9�͠@��T����)h��6ݤ��T���҂d��z����\�+�l��-�.��V��A��oB��iK^�R����%����4���2o͞���/������Z��՘�!�*�����=ȝ�7��<��� �v"`h��[l8�I|����b�UƳҎk���R�	���H��$&����o>}.�v���z��,�?�E�`G#lԠ?EF�Aɠ��A���?/(���w<ioA-�������Q���N�����9�Y�Q���T���gD�wD������#��r#免����d	�xWU��'z�!�=���-ܥk}x�s"�h��]ۉ��.��h'���x���b�M��B���G-BT{��Yy9�<54�`Ƭ^�.�ϑ�~�n�-�	̞�F�k�=I�GjbG�|n�&݌�~�o)s��v����ȫ�d�.q?5Cv4QC�nR��v.S*��F�ʀ��rx$�!ҕ*w��%�*����ZP��#����q�=�y�߻g����U7�ILv�O���rxK�+�)ߑE���X̮*�^��|B׿b����7��Y�vW��l���)��@34��AAJ�J1D�'�;��W����1c�]��éS� .�q(�0m�Ϗ�قM9��K��Ҿ�~����;�����We���_��+z)>en�M���Y#Y�Ң��M[��6�c�Be�{]܍��]"�������P�~��7���zӦEi�s$=�b���H�3 �*3��	OPٷ�g�Д3wܗ߯n3:��d�8$~@��nRk/=8aR^vO�<!�ue�*7ޖ�z�r�V�� ��g�{�X�j��L5��jnѹf2��������+/��.��܁O���N�(�KO�O>A�l���b�mՂH���V��s2
�mk���O�E�Om�"�4�)x^�L&b4���}�����C��lϟ��K1�W��=L� �	����x �؞z�1z��I�����@��"�oy�1�֠�'1LM�����ʙĸ�vZK0��������+A���tc���	��\b�0�R�j�x���V���ڧlWZ��0�H�^�%��T5����s�~Z/�\���2�-�.�%%ϱ�u��.9���w��1PT���/��1΄���=�%n�����I��sc_(����NQ!�
F�.��i�lg�$�� �.(D�3�i����<w&$��� ������(}�˧Q��C[��#��J�4��՚o7�L�3�0��<y�����Y$�#fU��
T���	�(��*O<��(mAnV#� �S���������E8��8��X@ϙ�Zc{�\�lE��W�:����i�����۵�c���6��`R1=��T$����>T�8�}������ַ�L6������<E�GM|��D��<B;�����O"f87���b�FZP���M>���Z��4�{e?W��%E�����,(��`HC��88`\��l*�q�{"5��q{���L��=�G�U���:����٦z�
��X��ޱ�H����*9��zH�	��G6SOV%�-�?܊,����J^�K)�.Be���ǂ7n�o��A\@y�.�nr��C2m��'�&�a�����JcN9^' �F�%Y!H ���l����vJD��!:�q������4���^����Bha�r�<!uM@���7�.I ~�t��|��&���ã:�Hϯ�tSŴx�hNdA����<&�zE��H������h��K�xDh�a��@&�tLdRmI5@ez�m�^m1�c���\G��XCvLrΌ��cE6]�#8�h��bCr��T-��oU>�$��03-��ӵ�V����/�!g�heP�A����;{���3b�R�
�9_*�[P���Mr�����X�ڀ�3�?��hk��$p��!P�O%���O����/�~�������bҷאJߚc'�r���/3"KɕF���݈�e��4r�m��\Sf*�����t��(%-��'�n���^%��'ĪU��%�q=�I��3O�(�{�B�*-��%�̛hH�[����ά4��J���]|
��(g���E`������J�;���M�3(`^�Dsq[Yd��j�y2�\gCQP
��z̫}f 6"���qx��X�����1j�2*�g @�Mq���bq�5̼�@��ө��*���$�X#ȯ˫>"�2	π�Dn�J4����_ˡUW�q�a��ᷗ��}U:K!��Rl^�K,���1�>��J����x}6"pw-e����z�๡��HV!�G%���y j�5y��WM�_�K�%D�o�h9�c�p?�W>h�Ǽ&V�o�O��  w��G�	�X�����
�L�?��Tز�&�{slC���� '��}+n@��?	��;B4�HW�`�2gJ�f�"3�)�C��
�u҂��gbGn�g��/*wg�ӬX�p��R1 ��0M����<�ƿ�{2��q1�^��`�2���	���D��ܦ��3~�|�g$�Z�4}H�>}�>
��I��{K�ܺ�O��(�p���}H���X#(����`AaF�d�i���1Z�Ʊ�R粬�k��q7#���s�{� }jY.w��I�tb\{���B�w�� \ݖc�~/�]z7��%<�L�O{����(aC-�-az��O"@��ek�.%�EX��3�HÙ�A�N�i��hrĜY�B`��<@�խ�$���q���C٭%�(G���m�ۥt�;���kǮmƈ����?�%Sx�{�^�(���s@P n|#�޹�^���@Α���`���Ĩ w:�Uh���$�ڙ�}�@��z
�s��ěfH@�U�X���0�ԥ�%�J��vMm#J���L��iRx�{�ʧr���$��_~�( g	���]�lՊs���!Q,*�a��ᾷ����Qf>X��
���t���Ԏ�!"��S��پ��]:ɱ��hb31������[��3�&����9ybv,␧��w��WUk\��;��
��)�l�D���c�L��S��H�=�۔�Z5{���Q%d)��o��s/�/�#:{L�'���;Z}v�A@��OEd;i�U���عr׋����7l�.�r�.��ȓ�t���u��ŕl��Rd�\��m�
`r���c�x��y/_&��rYr� �j��\u�m9_�Œgs�QEk3|"���+⺣�� [�(6ƕ��;�/�z8�rzy���y�3��Ϟ��=J3�|��D�`ʉGҜJjt�؄�f�A�Z�����e)&_��z~�j&2典�x�3�l�De7��SFY_���n"�n�� ے����+��q�n3��3"��L&u�E�o�B�eZ6�h=�8v�J��F�s�2�m���~#�^@��h.��f��n���Ic�Z)��H��͆���qH(:h_�
	Ŷ��^N�̆�Թ���ce`3���lI�VZ��������M-Bc��Yuf�����}�x[ګ%�5<�+��)���l�g���"^��x�+[O�_cY^����������U���=�7F�U@3��<1����(`PÜ�}� ���¼TJ�	3��t8f
x뤖q��]	�ނ��������i� �L��TEf�z�vRB�`S�o=0]�of��e�A�}4&�C�R��pK����&�����R�%�X�ڷl�� `,���:aƦ��f͎7r�`�	��q��L������ز���^3���
	�n E����/��u'͕G�^�?�r�^�Hr	�F��^��X��$b�+V9@�ޗ�2�� ����A/,��9�Ss̜ڀf�o��F�m"e��'#�HnC�n�X맨֨������i���.�Ʀڱg8ů�E�P�b���x@Oqr��#��0�|�V��`�B���z[J���`vq�LxG���Z���BR��m�^_�yy�h�նɥȀg9��6Rg��H�; �`�^h�K�%�8��A�{�%��j!QC�P����RK�CE湦��8_����''Gos���5�곞L��Ɩ;��2�!@H��~>�5C�����&M(O����?$ʲw !�`����u-h>;�{��bI�ձ/�O�)r���� ��`HK�-�\4���" �Ⱦ>�v��5��#C�B��!}�<�]�|��o�f[�`��by�e+�'.�7S�Hx����#�=�~�͒sA�t�j+=+#/�w=����##�u�R���f�6.�:�>�v֑�S���k>��2R�9��
�EInASO�����%��o�85�e��12m#��16�����JM"�A��aA�-��2TB�.��f�~�KT��=�0��I�,��Q*iM��c�I��Աf��.#��i���>���Z�B�c���BҲ��o�%��kI����SKZ:Y����j���a)��V�]�TD�sg����Jτa��nJ0�t�W�7'�C�B=��'�V5K�i��'\VP��I.�9Zu'�.�M!xi��1ۗ	�ci���{)����XR����ygI��X#�ٍ^QuM|L�\D�;�8Y��E��*�V���f�D�"�;2�����_}~|�;ۃg�
�X��%Kj*�U���"5ﳴ2���ʉC��V���\�Pы��{Yڒ��}[�n`���o����w��W���;J�H%���yj?Cw]�)1�l7O#&���D�du�dO��);����T��Y-�Ao��ܟ؀Գ�=}��H��!ѹG˫�6���y3�Q����G��p� ����\�.�o��*�b�c��\	�Z�I��[�W�