��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-�L-.��ajF	h�1��CC�ӕ�S�����0���9y����@G��8����k���Ƅ����j+0�j�8b����[ɊYxh��4��i�t�!��+>��ʔ���W+���o=���L�i�1:��?�g-m�V!L�y�u�
��oN�l�ڎ�b%Q����2tujM����kMI��y�7��v�ZԻE��{^��>Z�lxH�IR���i*��j�=�se\��u����������Q���f�ݠm��k�8r�9J\8����TJ��X�P� ��Ԝ2�M�}�`�x������R�W#�T���J;�,��>]kx��QmU��vG��n8j�l���,�U��<%�c����hw�s$��gt�FQ�<�IyN���Y�	R�)Y�S�VfH���!��n9�����!��ִ�80�8�WS�si[��[���*uD
.-���,u����5�s��E�%V�8�����[�O�̵]!V�x�Mp˷νǮ��<0��4.�P�]30�-�&�5�n�P���GC�*6���vp�O��կ
D�#�BG��2ǽ�4d�I�;	r���)ij��\�L-���=�?��%�;{�Z�Y����I �:U��T�����dB�M�0Y��Eg���'�����e�!�?1����^�X�����6�C�)Xɻ4(h��7�.�b��V��%�}��^���T��/�<n�q~hP����|���V��z}�˴�8�L�`�d��}=�
~�Ƕ�`v�����~@�!�Q}!��^q�
�nj�:Mj�|b�@��9����!�A���ߑ��wC��i{0��$D�ڶw�����y0QP-��4������*X�$�H�	3���Z����	��0'_FFFo\9^I��,Z:�k��ϓ�]]\��]z�� tp9N5Ә_be�[\�S�6Ŗ���y��8�ƅ��qe8ٱB����S�5�|%ݱ�h!�F�0�D#}��*�,��܂)څ�p��t8�Q3��L�g8*"$pdY��iЩĲnj������_hYgz�$�Q��]WZ�+ѱ�%Pm������Ar��ܑ���kk���Jh`�	�-��p?����"�4f.94_I��F��h��;�����i�wғ8�M!<����I-�R ��4�F������''�3_��*��x��}h^乞��g��r/�Ŏ��"�����`���<"8D��qu@n�N��!�:Pf2�IW�=Y�9l��yP{��/���	����	MD�8z�{��)�?�i�K>BO�0y�9S��!��������}M�:�(��jL���z�+5��-ޚ��E�<��]���̿Y�}��i��_
b6k]��M$��\�lɐݏ�+����TF�h��֋a��ť�h��1���%����3U��-�]t���Hp����ڠ4u_Z�c���A�(��H�3EL	��p�g7** �4�J�k�0�:���m$�]��I���]:f�o�d�5�y�n,v��l�h>%���%nf�ǚE� &RX!S6�L��m����By-��O�sI>�O݇7w��z$����e�
V��_� �[���R��g��2�{���\g�jSN��a\�cRۤ�_ݠb���s�)� �g�b�8|\=9k�����z�m����B�R�EV��w+f"��zA��˪0]�X\ۛ'�N�.�]]�'�?�N.�N߫��x�a
#z��ލwUY��S�~D�	�o��>���ڻ:y
Il�-��N����
(���K;�2 �u*�	�w�����./�v�<*W�^�MAupH����?:�|U/h؀����:��QG6��&��11��L��pr"�/@s��"%�<!���h4����ħ̤�GQ��e��Vp�+p(o|C��M �
�����.��Y%s�N>�����]C�j���G��[i���L���fC=�P��K%��2 ���#�Չu�g���23a)�mԄ��A���Y���VI۝���@DP��]O�|'�!���]��og��@��nݞ���KxZM�0m����r��<�г}�h�ǅ�ll��p"�v��l�����~7���6�of�㼠9a��y���%P����E?��1���9�~��6���>H�q�� S�m��L�r�SQݖx����H�@A*1jT� �
E�̹������Ckk���J0%�72;��3"}|aZY�dNŚ�<9xDヰ����l�fl���KǕ)=1#�s	�1ݖO�I�U&�w��-i��]A^�~���?>4����%��Xx7�XM�7Q�b`v����'���n�~E��ye-r�?*�S`��G��<u1�����M[V�#zN��90�^�'^&^��6]���+4<!n�x��w���,�J����]��zi��&�]���ق��:vZ�U����Mɚ�����[�]����<��@���=�Yˣ}1S�g��IF���ha�l�#�z������H�ʗ��B)A��l�]d�������(��,�#��r1���c���״��Z�P���_6�z"莱�k/�Љ�HG�zCt�� �TA�^ɛ{*M<���E)nOJ޴���� ���,��'Ξ68^�M6��{����q�B�`9���p+v_.bLˠ)�p0*�������4;R��'E��Tn�;��5a�˲�zdv��0	�^���l* � y=`����]�,� ����G�m��L�y'��>@v�YH�l(m��<m�G�r��q�����:�n��G L��|g|8^�*����_�+�Rq��[�"xVb���?{-��[=`9q�?R�f���/�]�O�`�4.�io*4���S���+��F90g�J�LC ���,����pw�x<��&n���G��Ǻ�yQ��;ރ�����˥��Y��۞$����M��,��o(�m�J}�t���r�����d��+b��P���l����d3���=5?����ұ�	̂��s稏��i&!d��&��jO�7YVU�ʹ�=sl�%�_kS���k	��@�M~|Z(aY�
MщnZi[�H�y���B<���5��4�!Av�ր��҇q�hMu
cD' ��C�J�ʋ��f޴}>�����WF�/��9��S�5-�,���G�_�vl���>HR���u&!d]�{�j��O�h���7����wTt�Dà�r��}�� $ݓ�_��y'NO���ӥY����N#�"�5Yr����-c��_&�~\�,�l���-%�3��4�fRXV����C"J"��c��K3�~�ٛ|Uf�ٚ���ܩ�ޓ�.ͬl�:�q����B�m"xDݻ�$�7�_�S)�ɬ�U�XǶ��^VFu�D���x�v��YvS�٠ J��� ���Nz��+<�3��8�)}^E7,|��"޶ٓ5�'�A����|+fz�ky;�d�h"�0<�*�<һ.9����sP�.b[tS��ދ�;��U�w喛�K�:��V�Pr]�ks���rc�r\�b�0Zy�xS\��~�i���)k����f*�|�R&�`�K{�A��.��7/y�Jwn��{s���+����w�팥Tp$�8�	}豶���j���LZ��bՉ�*A���
|���ر�Q��t�z��7�ލ��δi��N�>�J�ձ�pkm��G,a�uߋl�̈G�qe��O�/�M�г\Y�s��̾��,���^�ʔ�T��~�����o�5]h�~`����	��e���LP'H~�Ys�O�"4F�M�:��lۣ<�;�?���s��{�1���l�6\n�Yȇ�h�͙�$�o�&N�g�H�>qTɈ#��ĝ:�aU*%vO�G���&�`��`��E5]���eߝ�P
I �N�&E�:�@n�,����|%x�!d��J��K�����Ҙ6bd;_�]�WX�� ���]W��4�g7Hb�ٻot&	kJ��D��Y&�.���9�<O��h���JS�F��*�ǫZ���I�������K�
��1��V6�T�U��*w>�%�
 �!}��gs���8��~Ξס���ʱ^� 0����ֺ�l�U@)��׀�{�Ҙv���<��i�w������#��(/D[f�6.^���l���(����z���',y-�M=3&��*,��L��*��2E�1Bm���.��\��b�%D둁տ+ZM|~��ݳ���$� A���_����k�/	z2��6�W&5�d�ǫpNؽ[M���(��S/�-AxZG�!>V��ٳʲ�.��>�0��XK�	��ԙ�D3J�ܝ;���K ��QzN��N�.�En�Ǔ�c핢E?<�K$�����Z���:�:�@ƣl�WqPޮ�nC;�Crq���
��K7���!��S�B7q��pK�ˉ��P+
��(QS�?���r�߲P&�<۶K�����ڄ��Q�*��Z
3����ua���7DwMg�&���^�	A�҅:���}������ikD���'�c�9s)'��"���<�ƓGՋ�&�U��F@��4��^����b�,qD�=�UqZ2��-�[�ߵ�(M���V����%n\mѶ��=FlwzJ���
��'��8G�w���B�\v�ɥ��d)6w_${>������9Z/ٮe
�-�ͨ�_p��X�ڬ������F;l���z�\�>@���h�XG�����D�\�+]�[<�Hwk�f\�^ŗП��e'ԣ?6��䛬�����~Xv��0Q�,|t��0g�\&����j�G�>�q�F����٨uIql����I2�^/^���� �`�@�M���5P�T^X��Z*��٩j(�k0I#���&�� gI���O�0���r? �]���qFQ��ssR�ӈ[�p��pf�?o���a�7FȈ+T���݃�$� ���y&�� �_��^oF�MV*�5E�(��8��]oJ��������;�i�=�!k�߄GV%�(����6n�m�f����;���Ӟ�ʂu�_� ��XbOk#}m�Gӈm��PY����t�)�"�����\��#��2v�s�jiYo�Q2��gis�*�"�Qh���~��'�,ֹm� 
���o\��{�WBKˌ@	z ����3�T<&�	��*$�Y���x�4^g<�y��Fy����,��2��D+��ZZ+	M�� ���8&[ j��ԩJ�H��5�.
��NY�L\n4�wM)�r�p���d\����e�@�����C(|�T~WXl,�~R���Am�l��!޶��y=�E��k	�c�fE��$�,�CL�R���9��?	�慐�m���"�v"r<Z�4�8��{���07e2�0a�8l�R�$8I�ԩ��W�H��%�&��STx
�Yd�t�S�oMg�+���I�H���?!�������d�h�=��ۼV��������7�j�;/)Un�"/[�`��K�� �QZW���B��Fw��ZzY!��w��"�S�`xMsKq�4p�
�l��rb!Z�Mf��g��&���Vm��hv,j��z�b���`%�e�R��H����k�V,xp�%Qc�+�2C͒�Af I֩w=թJ�;?}9q���ث���Whڂ9E{|�ا��]�;o�Zy���Ͳ�!�2Y�ϑ�}�ń���s-�&ׁ�7t�/�H��>=��-�����+��Ơ��Mow� ����XW��H���_ioQ�2��{mkL��	o(���x��5�J�I2%�[�ؐbu�Z#9�bBM@|�n�&=����&K&�<��4'~�Ii�B�o	U׏��A������$t���,�A��qև��2�@3� �� c/��REf!��������5��AF�c�z\�|e-���o�m�d�
3gF��]� �	:L���V�Q]9���a�9�|�_Mc�R�}�ڋ�<.���6ΛL�]Bd�|���ތ�\�E����B��-���Ǩ��ۇ�dx=�ؾ�w_@dWu$�z$�2-T��`t$9�w��c
�GF{PY<��Ӽ������!N��h���;&e����Р�w����v�h�ūp��A�����0����n@ȳi�0��6��1<U��\�v�������GB�GEA�;�N��ۗ�037��O �Iq�2%T���I@��
a�-�g��	WN@�I1Hʓ�d���J��o61�ð̙��q�'�R�8R�vq�rWe� V*��L/C�WT��H��6u�g��7�C��_��/�+;%�Yu�]��qxr3��Wo�\�o��&�c��c�
^"%����]�g3�����?�������k�b�G�S��Cٞep�n��P�M�w�~9�v�E8�a��`Y�? d�jFy�^��ֆt?��@�͇ڄMP������A�=ҳ��FI��e5�v#6:��6����]o����W���_��a~U*�0u�50�V�0>��v*���jg8���S���?J\���Py��e��Ԭ�~ �����}�pB{��M���7���Xv�� Qv�v���H��k��+J|P6�w���]
A�mɞ)���rr�p��ߨ:�T o%�ŒCm��FG�l��D���ٵ���/4�k
E�^��(Z'�KK���Q5E�;���(L�P�h�ɩ]���;J��F}���S�b.��锒0e�����_*aO�D��|4т��x���l����}�����-ݕ��	!�Av3Y�v>�h�����phה����mg�w�z�����2����r����s�8�9�BhE���︟w�C�$��c���W�|�Q�%;V����<Fi�h(�ˀX�]vs1�����O��M+�\,6蹠M�!��8���T�r�q��9T�@�t}��Ԛw�S��^��L��K=�O��p�~�Oؐ��fna������ۊյ� ���?�s�r���<��$&՛\��l�?��K/2���Z9�^9�����*�r�Y,��κ� 7�YC�ޭ�y�� H�67�מ���S��'b�7��Ľ��#S������ֈ�
�'wf5j���|kC'�w� ����Q,�� ] �Hdg��0�5Ko�'R&�=�gP@�{������t��<��Ux� cl��9J6��,^�F� �mҾ���șp��c%N5�a�D�3"��X�����Gf�)X��;��U�1���9��ʯ�n����'�E஡n��H��L��w����!m&7ɔfb��|�(�;���4�b�"�]�z�$~���P���:>��W�F�7�7�%P·��H�ؙڦ������Ab�K����P������{Gq�r}(bv�MW�\`���\չ�=����?����ٳ���Ad�	�$��1���Q)��ݜ[v�$�<�#n���[5��Xݺ9����%�� �� �|Q|�v��XhNI��J�kz驤��j�V����Bg�'��-1;�<��o�S������;��`<�D�a��y���0+��UBK���-T1L�]i/��ٝ����p��glK�z��W%�4�<$�Wg0G����d�o?����9\���§�I�N�4�2s'ぃ�Π	��	r���Q>��@�v���/שQo�%^-�}V`��or�`VkVJ�ێ�����Z�rrޗq���Rb�'`B��ŏ�'&I�LI�4dF�����pAɥQK��/�'��	�D4��']��A���\�5R 1���Ͻ6�l�c��4�6��PРp��t���؅�gM���H���oj'�|F�Y�tR���P~���΁u O6=J�B��T:�x4�3�����&������'�o�FB�9.�
)����=��<ա3ٛI/f�*zUֳ-����9�R���m��RA�x�������:eh��&����.z3Y�J����>p���=�G� co1((���T�W�X���\�ݝ*����(n�C�cܙ��$ASu�X!��2�z�(�S7��膈�{���o��xmF#뤷
8�v��]�C9��)��sw�2Ф�dx��7N�������q�_F�xR&�w��5��3��ȕ�1c52��]Q��Ud���ԉ�b$����z���OUH`�v��J�� �Y�=��'�<��O8R��	�����<���+;�m_��N�FU�X9�B.�,�J}�%�2Iw�~�ӮM�@�O�R8��^_��f7~�Y�\���,袂G�%PI�Y�W����i�>���_ѻ��R7��@��N���c�:����_� q�I��7���d}���U�-��G�2/ �&�L����e�3�����Vo*Kj���
{�7!"�_?�o���S�>��[_�!6ё�Zi�V�<7$6_M�1�QLƏ%�a�-#?�v��4�f?�g̱;��,wS�H�i�\�EE����x#٭R���6�#���I'���Z���0V"c;��+�eeo�8�W�FO��	+p6sd�/����
z�|�.û��U�y.n�Бmo��&�aR�"/6��L1�T�4Ot��n7,Z;��B�sK����s��VO����s:Oi�-C��|�8���a��[Y̰o��'���/��A�0<��	�TK��J��ϼ�cmnv�c���k�)A!��C!�y��bY-o�I~��� �o�GCb��͞�lY�\`v$5��G'8�< _�]2����qe-~{<�_	6���P|~�(m-�UQ��V�1ќE�f��k�|ѕ��4lc�H~�y"U1��t��V��麅>|���(3C�j_ch�~v�OE ��GiB�Ve��C���;K&�;��3�$����l-bqHeD$��j�h�/ee�jH����q������TI߯+�w�*�U6XȞ��s���<ʸ	&��ܸ�ʆ��jڴm��9)�$Kb���"�l)'��eQG�|!:qB@����/���8^�=5Z�pɈ�r�MƵ�
>aݭ�&�i{f6I'���J^ҽ��0�W���kI�[����M�;2�$�k���Ѹ�ג	b�>ށ�aP`)���ݨ_�*U*&h�ڬ&?]"D��Kb��Ku��'~PMs�k�XZ����=YݺQj��9�A�AQ��J���������y�m!Z��7œl�ٽN�}�z�l͑�4�$+JM�(zhZ��n^ȁ�"�g
L�ձ5��)�rV�%vA	����l��m�\{~��-r���Ȕ��܋Y�f��Q��bOOa%?F��?2r�5�W�U��JA*W��6�#�+ڎTO�{���=I��6�~M��Q�W��Lg?*CВ*ӱ��� ��#��1���4�	���{���+��M���&\	�A�̃���i�� �)���)���
4W��nV��
��3�x�m?'*�aټoe���@p�*�%|�i]7�U�"iG�nC�:؆���߈TՀD8����6���ꡪ�u%��� �©+�d�a�`�؎��C�2��	�)�T��'��jl�m�kp��;��	����RU���<oCk�d8�+au�U��qXE�]A!�m�Ǹ/Ø��?���e��Rl�|���Uk��0�9���WXom��OJM��;.�i )Xnq����ͼϐd2d�ܥ;B°$삥8"�*߸:x�=8�;�a�q$B�y�h�R]mǍB�� >��=�Փ2���a�>�Z�k�^9M���4��`)z�n��ɸ�,/�{�ݍ��_�ϻ��.�J�%=_jN1�V/%����:�5�����HT ����fG�G��|v��ua�5fR�Q6�X��Ѳ�uD�������ð�P6�y�	$l7ۧd��˜Zp�[�|��W�r�Ky7l�7c��o��r!������p��C]�c'�������3��=6���N�Z�&�8�jGƚ}/�w�y�Ց2���� F�p��8U6���yV�$�������-!M݋w!���R�5`T��m�1ۤ��~zSV�P����l����6on|�w�u�ֱ?�vR��j�H�#�h>����ul�6��-"à� �.o)T��Ty삗6�}����kkǵt�[��O�r�D�Y�`_�����7j�]��s&[�a�:�.�}��X� T~�W��x��A&����h��=�F8��تD5*W�&j������7���P�� ,�91E+g��W�X��zH�N[nU����u_�h���P]E��`��&x7*r��rk�UN
�cJ�C�*1��kU"iݙL�n/�1�¤�s�KB�&��Y�OG��_<0ܳ�S�*�P�g�������0��o¤�9sQ��±���M�S�^zOul�N�y*��u�'b�Ҩ�I�����3l�q��y7ݚ��e -QX{�@K���~�͠��T.��iAo� &�Rn;�O�C:j������y�,��X9��R~�F��16���ݦ�P���mq��n���u¸q���I!��2�8�s[��q���FL��ږUuw[k�=�Cb[f�]+���[�|$ �+uWBJW�i-uUA�B�\ڱA���W!a����!� b�M:p49�l@P쥚1�3]��6�a�ɔ�m_�1N>A��_s=n�+�w�~Q%�
�|��eab�Ut�BV[(������`�t+��ߥC��a���dɕ�ő�X�a�@�ᱮ�d����F��.)�BҲh�tā]0�nl!1]RBm�r_�y�7�BW��Ɉ-��u�!M����SH�!*Id����l�A|���/2��"k��Ջ��I��ะ4Ku9?I�ic:��֥��E�S���&�mi?z����:�F�/��rd)�>�$հAv{S?��ד;���CF�t�qۥʙ�Eϫ���V�c���9I�4@�Ӡo̅�����[�eL���~O�1�����m�9���1m���*9�a�~~�*;�MҐ�U���|�)՝9e�P"
^�*}xQ��@�'���<@�vl��&g�v�ΉZ#����4��	z������;	ǯ�������X�'��)���ֲ��MCI��~��$P��p���\�E�9�+���2k'��tĎ��SYw���W����M��L����*��^�H!Nq#������9x5��6M���XK�Vw�iF�ʯ�����}����Eʀ��N���K^�S���k�f>�m��\d6 3#��������8w�ۺv) �Ii�R���R�AR`�޽���\6<�'�� �bn�1�rK�HP��^�ّԲ���*�t6_�����9io_Ζ�r�aH���+AU%޹eY>0�Z���πl}�����~��h�A�ú?x6i@�&zf0�u  ���2TR2��M�,�ua
�j���Ů>���n�w{ٺ���j��]U��u��C a��l/��-�uUaQ�Goh%q��~K�C�At�bvD!Syy��4{�,%c�x�r~ {�9T?��A!�W�z�I��|����E�r���F"�P'!�|���-���k\6g}jAƶ?���	(�f^�P�<�����z�|d����b���}��J�..gke�á�]��/�߶����e�܇�{a�1X�e���.y26���G4x���qEd
v`Y5t��ŚP�.�ֹ7�����&3�����r�l�k�{�??X�#bg�C�5�2O�$�_��"���=k�x�o�Kt�A}!��{*@�������MK���
QO��ꯑ�D�l�2����#
m�����n*��|$=�\��6����J�A�9nnr8\�1#�����_�ĺ�Gz��d9񢋘�j��G�6�-/�jQO)�p�U��@rlqhuʐP���L�V��.&�"�J�T�Mw^H!����(^�M��hH˘򧻚h����~uk ���Ĩ������]!��y)̯��p��?ա��}���~�@�����'��%9���PvRe�G_'ZS5�D`��.s:��oX�D�r���7��,� ������}�����F�=<G�%S!7�8��b�G���R�3��E�w�~:܎DL�j,��' [���4��}(k݀0A�z�UX�btO3Y�C�N�Ü�$E0	�Z�Jtn���G`�e�-G�]�7�`�e�UZ��v~MG���7�sn{����QN��z�BE�"'(�~�g���|�c���M�z���`�Y��L7�SfZE�?��
,vgx�t�XJ
���E��9g%��D��P�^�T�~җ��l\��ҳ�q��[����B�U�+�^�=���I�q�� �,W]7�䭇#��
{�� n����Fk>����lj!��� f��AxTΡ�J�2��P�S�Y����DA�]�C|hd�0���3j��cgf�� @��I�X�p�8���{o�o#^sd&�Y2��MQ��;�Q�Y�� �d�l�D�r��!A,p��/�z;�:vdT�n�G� ꉂv�~;@�[#r�gD?���pO^�T�6Y���g��R��2�n6	S����I����/7���i�M�f�ҿ�J��9�=%fM�:o�$j� �1��k03Uv��O�Խ��ih?Κ�? �8a
�e��+E�H�V��0[N:r�^x���I�L���x��g$�i2l����+]����&?��Y�2�)9��I���ZzK3J�sgk�P�B h~o1�*e���M�X^�`��bri*�ν/�����|4	�V�l:U5��+N�y$�d����<L0���t�ǜ���	a�^�����ju�.?�x�f����k"�Piň4t&O�o�ޣ|J�U��)^�ƹ~�!p#js�q(&݆�1�]��0�m�l�ƈ���7w�h-����S�M�15'xx�3��]EKt-�τ��9���i[�pޮ�A��o0ܓ�*W�Gp� �Q��* �%)҂IAtc����=I�ud�&K��$jh��n���\��q&,��\���<��\?�\�	���Y�j�W�RW2
ɞSL������UK����}g���q���МB�b�� ���pN�w�)��,��/&�I3��MO�E�$z�����B#���)������H(�^
�^�l���rW$�F�sj~�tkl����oNdt��H���C6�NЇ�V�6\����"���FQ8�jXh g���h�@�B��~�]����*���מ�b��t���@��rϦ��l=�mPl��VA��w;<�:2u��5��yo������'��* �n��!�y���ȱ �\d!a�	��DIϙ7am�MI�L�[+#��Bb�q�ID��zP����/5��H� ��y~6�W��������������'����J{qЊ��@䃛s���/@x@�slĸ� *g�ׂ�Q=���p���sȠ��� )��M%��=����jx�E���c��doC�*��A�T^Y�{?�6t�-�"��9��R^~X��Y�i�h<k�e"�G�OZr�b�����aq�sSHX{͔�)&�ȯ(ޯb��M��u
֙��%T`�0hx�@����خ�S��m���:�m��^�*}ukPs���������d%�F3 =x�n�1���ET�Wm��7t���t��Ne*��� m�R�呰���b���{[�����,�ç�@h���8�ǵ���9Kh�d8��B�8�I�4s+���١�����h
�P^]���ٙF����1�W�dD��
:�/yy�]�@�G��)�N���mnk*����0��W˅������^�J�0�2�.Z0�0�
9�ڴ���#rNB�[	A�����y�1>H��!�b��1O�����u�*-����\���sC�a@.V�W� �i��0��q��}v�&�g�*-(Z2�sFi���5@����G.�+��m$��7��9�o�0O\� ����ڛG �I�{���{�7>Ύo���PHI��g��e;�� _�����0�ۮ�3�ϡ�p��.,ͭt&�ǰ`\���6��0�Hl����w�#Iғ� ���+g.̲7�f'��wҠ	!�L��g��y��k��Vw��D�;��~I6���D��oC�,��,��{�N!�#���]�7{ȏ�=Y������޿-o\=U����$3c���&�jm-JF�P�n'l��� �H�h��;���{�F���6\���fbo_W�'��e"��r y|X��b�	Q���(`�a�`�`y!c�ڬ\�T���?[
�����U&#W�cC�$*ṽ �ۯ��N~ݘ��-�ޚ�:������c�pd��`�e�+�fI-w6V��; `���w��wum�FU$� ��D�a:$O�kK�|U�vg����l�+lrS�IX�,#�F�N��&�78B֟�Ѥ�ًn�|л���Nx��0�G���?SQ�8���!��a�_*�O��u@poٖL��h�#��QΈ j�Q�nF�1�T^-���i!/<��S��vt9K'�-����q���[ڏ�&�	���$���?�[B$x�G���S�ޣ#����ZbLޞ��l��b�8���j�V��.�@#����:a���fwm��᩿
Y�Q�4~X�1�#�Ø�}o������,AB�(�tm�xu�25:<�'��H�����;�/
��e1�垹̂*t��^ߖ�A����a��D��7t�x������0��V������R�jfm8��w����}@w"[s��_�+eP�c%�I�!����"����ƌ�_��N(a�I����f��*�C%������t!�LJR�(qa ��@gP�z�H�̊e�R-��$7�.��n��G����5������D��({;�-��Pw��U?;]��$Ƣ�_�j`]É��Sm�MqB~��U�ŗ=j���o�o�I�Q�������N�Y��FG���/��{Т=�%>(�<�g�d�p<0s�	؈��� ͡�($7�e���E�*�O��Ob}�֡�zcp:2�8^��҄%+-:?�z	~=4)��v*����eU�ON�����F4V�Y��T���y�e_�䦝�ٝ�.}0���5�U��2��QMG"�p!�.�`o��hv�RC/�Ж�����ۖ>��+8���YMAf��)M�O�" �܉S�o�!_�0�,��엶�! �����sq���*�N~���{�������t���!��t=	��1@%qj��,T-�D0Q�@����PU�.?�w��io���1��gF3��(����!`Lz��b��֠F��Xq������͹p��:���(��{q�T ��5��t�I�=�ǽs�:����>1b�1�W)��S�#��������S��,�H�m���{i6(l�����[*?koqB��}!�`k�R��8�~W8�|�����JU%�26���Cȣ���p���@x�������Ԗ�W�p|{��x�{��B��WX2�Ж��j���f����U���4V��:�x >n_��0Ю);�6�j�]b����� e��;�V\����7�Ա����轁t�]J�w�qWm�����FV�t�����C�-#����؞�T���v�l�l�;�56^ө�5ގ��W�_B�d���T[S#�sN�Tz�)�l�j����X,+�W*�ا�+�R���Ҽ��mܽ���.
�d}����vp#Y���:|��k�{y���pAp�|�зH�F�THyI��`�DtV���ҕ�Uj9v�6�R!M��p� ���W>�<KFi�#3�j���uվ����~I�tO���ޅ�9�<u��oyxj�?�[+��R�.)�=H��(��Q�����L>��[9zC7�,z��J�T��\�����Rܦ�q�Tf��Dj#u	$Ph����t'Vw<���������G����R�B�B1�{����6��Ө���V^���d0OUM��x��'M��Q�_](H�U�v�Le�����'.�.x����k���$��,4޵G���h��	�Fc�����'fh��7}ěD=R�!!L%�Sb���Ũ<�	ֲ� �w�{�[g���膖�rd��5���r}��SVl`�P}#�xX�{�>��^��'�yM�3�Bg\_ŴωxC�%��U(�9h��E����26@R�6���Y�H}(��.��r������ƝID\'$9H��TL�R+D�r�&
� �����ʟ���R˦n��_�ԧ��kwa��A�dE�^���wq��*�tp� j6擄Mp�*�hG���y���J�z䙯U����5��:��
B0�A�IE]����+Y�~
�!q�޲�D�*�2�Zcް�������bS&d�y+߰p�����ۅl"����a]�p��l��3T{��Fǘ�Z?�x�����R_��)�a&�8��i��l����L��U��E��4N�r\����_������<Rb�,X���?��a�$�+�,jj'�.�R�@:%rvG�c�,�X��h���t~`��f%Bƅ!n�6�w�t ױOd@')��P��);��2N�������Lg�W�Al9��k�  �v��jk|��u��kG �?{�7qOB�l�s5D�ܿ{b�LJZw�W���.	�w�A��Yq)��E�g���*
���l?�dh܆����|\���P&��[���s�^H(��3����9~�>)`J�F�TE��Vv�ٗ�����_Q��J1�Q��� �?��g�ԭ�~$d����=�fq޶�?>S&q�z�n���r�!�dd�
|�`�ᗏ�f���&����������/.H�yt�w=��5�kO ���ߖ��a�������P.£�}���HPMB���ćFh��
�6�?#W��
Kz�9:�L�"dx!��0]4��y"��Q>��A�)�1Dg�a|hX�g$`ƶ|0��kY*[*�� ��C�FĴ��u\�Μ�6���=�޾���f*���V�����fSB��zj�? ��������1�GO͋q�Rvܮ;1��5!����$��J���X<�`�}�[��}��'9�.��ݭ��ɯ�h��-@���ڏDCn�(GN��׌k�\�]���ɧ����5)`T=�HO&��)AeiE+��;�IiG	d�f����Hbf�t%����k���g#������t���Q�ڍj�z���Lp�N�M���%�Q�d���%����lv���'O�-[W�I��f8"N[�-��w��	=��h!��	��7�Փ$'�$���c�������W����u���Rec��O�l��JړX�~ö#�����_�:�nm9n�B�L|�K>�pK�f2 
�2��T�gF�'���/2��K�ǼcV� (L�'6l<��1���\���}�uw���TS':5t4�b̂li��{����z]�g�e���HQ��<�=�n�ٮ%���5��B��`�8�6{b�1��ܙݠ�v�B�`]�"6�9�o�,�T�t�Y�Y�h���e|���H4)����Qm�d�;���є���s���PX����ΗXX�ݾt=�C����g}�����Ǜ��@�Q|�G�J�ܵ�~��S�s'�x^��;�}Qj��W�̷����\��'.
�Y;K#�@����'�oA�2�w�nt�x�?�����vn�mj+�v��zL|T/'�9S�V�|(��i]l��M�4"���F(��RSAF��7��&5�~?�fl�Fu�o�\.��I>t��|F�s�<'����0ݐ+�^t�r�c�.S��!ɬ��ͦU�DFD����.E=h��H�*'����[�׹d�܎��PY���E�hZF�zV�<�����5(�S��X�O0
�+��+���SӈP���ٹ���F 60U�\�y�F&͓�.��D�q�I#����MKI���dW����?�������0gu��9Zӵ��������lC�"P��_��ˍ��Cj-@X��}jG�"� ��}�M��Ex���r��40Y�Ơv�.(o��