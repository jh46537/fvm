��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�=���,1�jӛXT�d݂��ߦi˅����H�����C��X(dj��@�=��� i����&o�)EH��sz�)n4}��KC]��,���(�B�%���S�y�7/΋҄��[�,����h"� �I3s}���>5#7u��M���eAY�jb;ڶ;�?R����Ag�YP�аWSL<��~&��[��+� �#�T�w� �/#^�~jV:e��?s��ރ����ձ�8�{t̺��?4/x����th����+n�Ԣr��?ګWR�.��M槠gW�d�|��� ��P%�i�Zp9<\<��r��k��0�?H$T����v�wO�>ߔ���m�"�Cc{��f�	��%��̉���;�(^�,��R�L�pn#4-e���IT�~o��n�a��V2�=�P�Z�xL�žp~�񤜲 c-_��b|K{��`;�k�/�d�~B�Ȣ��+��Vp�F��6<
�c�V��'�:�� ^Ң�L�#H��g��e{�@�����BcTZa-��d��-�C����ʬ����n0����&~1�`�y�����z���`�1(�D���	`v���򇘲3qڬ:��"�.W���N�`,���+/T��V�Ř	�-��s�E�0�QK�|r����}@	����mw��	�M��Z�쪒���!�O�QI�Z��^��k��ש�
;�B�x(!��c��'�~�N>��y����H��V7��c��~-q��&41�4I�=�_�qc)0HV,�wKU��y�ɻ�(�9km�G���vd���1{PL�m��i��]�]�u"e�]t�~��/��Y�d)2�Zr���tֽl���z���TY[s�k}NY�m�� p%�y�#NS���xi��FJ��EaLfq�Po�#�lq�c˸�E19|/�o�,����UA{�p!|�2!s��[�|���V�|�6�k���W4�Z~h 륩�x�Q㺡Oق�8e
�1Z_����3x2C/���d���ҿqA���q�X���X\�=��I�e��X�I�����.p��]�}�RQh�9���jD�0���$o"��uk#t)
1&���,�"��(��ղ� ��Cm�M�-ͨ��~�GߦV�fb[���֏��� �0�qg_t	���l6C�e?R�9��w4fO*^��X,�F������a�\������`���g�L���"���,DՃf>��?'�#(b���+6P�����u	�[!@�Aj���J�~~�&��B1��㳡wiff��pq?#���;�-��u���K���%�x*h� &�F��E��˜�}����P�(��Y���g��	�綘�[���09X#~g�� 1�c���po#MP��g�o��w�mI���Tia�~�9@�gx�� ��`��g.�ŵ%k�Y�;��E��tLz�j��2��/��,W��J��	4a�^`��X���1
1���f�Aq%�-����]{h����q������(���B�<̄���#�����t�Z+�?u���d|��������>�^��7�]()r��������_G�n��!�
��l�� ̒���bs��W��/?�h��Z�N��)u�I�x]|7�H4Fr5����tS��ӭhZ}8�_]L�bAD2���r1Ê�z��Lh���3���G�N{%H-?����Eqg-�U��r�������5����M��n1��ġ�	�B��p����9�ެT�+��aLvݔMi�k5;=m����yRW��"�-D-R�Fإԩp�p,�FT���fa�(�D�ß�$��>�b��U#��^�^�b� �K�]Xڗ���bn����Pc��8;�ǉb�FY��2�����DL���2��(�5!��,���Z�!i�������Y+�	����1N�|u��o��)0� ���&�U��b,Ys���`�_��\������zB@Q0��N��5T^���m[���ȶR��"p��{�|���`y&�E<$pAt%�x
�p%���ɓ�����t�6u�����E���GƉ��>x��F�0/�h���3>�<��d��L.@��<�/�j@ˮ��NI��X��pLѶ��?2_��cӥ��-Y�"<Ҵ�2�N>�2p]�o�J�]l�J�46�PV ����jr�K��.�H܀o\�Rv��;=�F�V��hj����RG^ʊ	��6�C��	^�	Y��2�Ϗa9��'�-��&F�˹���2#ݍ:��̉�����<IJ %��>��v�P�N�↉��[��Gb���騣Cg�� �\��Q���wƻ
36,�3��U�?x��C7����KB}ܰ�ɿ$���MKS��+DG|�-�e��ճ�:��"v�<���G��l��TV���UI�5p�)��(8��Zw l����m���b�eD�����7��m�B����Wз��d�1�U�Ht�i�>�|�� �k���0>��=9M�h�<�Ƃ g�U/�|��KS5��� ֞W��>aI�I0WآT��.Pr��r=�~$�7حVX�]_t���xStP�5P�88U��Yβ�gM�9�{��� ���sUZB
��5��m�MGŎkM�Ga. 5Delw�*�&f�?��"l�:��p�ǳ�#

��﭂^�Z(�Ѽ�o!Q��ԟ���깪��C΀}&I��ظ�K5��10��zT�Ę�Mu��ð���Sd�3� ��eFh�*���Tۖ]��N����&
������4���Ca�a(@��|���0aB���+}�)��5�nC�Q:{ƭ�}ԕ���*�B���P����8��C����5�m:	��_5^[D��/�D����m@�L�ʘ�ī���#C�?�SQ+����6��&R��Mп�eB�1�;�*?~Ҕ�F/�R�y1�h�:2mUQ��(\"�Ǳ����v�B�JZ�� �=Vݕ�lLi	�-3�Tp�*���oG8�/n~Oڙ���y�BȷϨ��2�����}��{so�:��k95��k��K�]���/��B�u�i��C�V���֎�d�KW����>���s?�>��(����"�l�/Q��>��j�曤����$i���A}B��!��d��um\�Lul�_��ܜdND��w�d�o��ϑ�quhY��l�}�D�ݶ�Uks�|2��a��'��!;�(]�]/�h����)ݙ���h��&���:\�H�%��D��2Cܟ�:�eP�Q&�����!/����]t�k!F�"���cC8������U��~�q�phć�ڛ�rd*f �\����>�4Tq4��AS?@�ĚM㱈}9�Nl��,�N?l�LT�_b�4iƆt�q�(��ꦃ35 ���.�;�?���Ke���j��W(u,� �E.kHw�>U��c�9�`- ͦ�{�����8�?|����%�TF���܅�|p����kj�V	�DY���y�.�FH׃����l� ���<������m�.����l��P�=��D�݇rqu�	y���%=E' 	�V�9�W�*�k��E�;�_���~gu��'AF�֋� {SQb4�/s��Y���^��	�q 2\�|>&���W��RB���,��L��xE��xF�:�湼=�L�vuV\�B����[B�ck������#�m�Ue,�xʕ�8YE�`��I8�I�O������`��8ҙQ���PzGG8���Nw�U/�=P�}�g@Ӫ�I ڋ�u�
��ޑ�޻EwA��?�O3~*��e�8䎗�}�Bs�����0�,p/�G�U+2@Ps]�B�y��NP&�������8`8�=�>:�ٛ`"�!��/��s��W��;���"i8nMMH����>���*�o�%�%��ٔ���ky�m�-V"�1#(�:���۷֗̷ H;�NTm �џi3t�_�j�p<��C�4^5�U6zwtvM��QS0���]w,�~����5�A���HE�]�$E�5qUy�7:	r��q;��?ǋ�|}�
��x�oE��>B1�0)��w�?xH�J^?-�E ��@$8u�B;����,.	���ݪk{&����z0�wy>#���9[�2�2FV[�c�C�n8���əuL�	z
(�����3�Mv
S�����=8��.}y �f�w���ƽ���{���@�6��[\}�s̻��wK�G�+}��b	:]��4��R����RX��xH7�|��?#B�Y��q�Y��&�1�@N�z�����H�����g�Ub������&ķ̼Ua��%�L����T���G�����t�����yL��!T�x~߮��Ai���ԡ�'�Bh�!��΄�97����<|p�M6V�^t˷�M���N�P���9=�.���)��.��D��'ty���q����pZ�]e���vn���.�����k��Ι-�VI� ����6�U8��tb�͉���*@7n$ ��ǆ��7��
���=a�̶�s Ք*�g?���A�p�B�z�A{MN�ؑ�mF =۹m���y��v|-��FܖW��&N��r;�Gp؞4n]Q1������Ͳ�.�&F�@�*&Q���E]&lN[����r�G�EvZ#�g��ު���S��Z_ }]��ly��x{�T��D&�-�J ҠC���|���1"$����I�T>N@�6�1U>�VCj����wCX�>i�E_�KT� �@��]'w�N>��z�m���qВ��W�HE*,&� B���b�y��Hx��eM?[C^�\�w���i�x�j����6�6���q-q��W*;S��,!Y�y}�px�;�IW�g��(��}��F���Sr��[��h�{�����
�\��j��G���%ە��y�n���H��Q��h�u������m�R�������<�~�f|OKi��>-�1��c�M���[�-U�YD&���58�7 ����,��_�C͠8U���U�K
Z�d��W?9i���{�g��7���Q�A�\��7G���5d.�2NND�S��]惉�6Z����{�_K�9R����x��^c����'R�W*� 4I_Y�;��
e�H�C��i��@�Y�x�3�ӺW���anb,�Q�Te�;(Vyo��;h;�0`ի�_������1�2\�n���2�;d�뱟���>S�9������(%���>��/l_R�1��H�����bF]�0zP�����zd�b�z�Z['�Y/}=�Nk��a�ǣ��on4�%��w����9.�U��1H��u��-%����x�6��_�+ט7:���gPed$x��{'�����l��o��ZRt�j9
9A7��sG~`�m�&̭7�Rw����M_FJ�=�{2���-��[9W~�3Q���d��Ȇ;�R;� nz{� �@��Ͼq�$F~.~��ػ���
�ya� /Fs�}��=K�.�z$�#��-�	��0ww��!L��w�/�nt��i\��#E.H���$|����ȕ�!��r#.]�
��],�\p^��yƈ��ҽ��e���9��i`��|�>�s�f.�t�����l̃�!B�0**��Z�p�;��qe�,L]���l��yK�qt5���� s��Y�~�=�H�Yat5Gu�Iқ����u ��Z����� <��+,�J
�l�.y�nUVDS��J����gmo|���w��~NWk�S���j%�y�k��6�~-���GKj�%w�1�|���, �S�$�"lr�_�κrD���J�73��#E����r�d҃��T�+���t�����*n�͎�?�*ʹ#���ǔ��G��٤1=4��x��3�˨�7�:ay׬Ս��?�T[�E��K����]#u`@�'%.�u�HƳP���%Do��m�k~`�C/�w��c ��c�&O�h���<�s��ӷ���t��Jr������~��+Ζ[�� �c�5���^ٝ��Ekeh=��\�qב0"������&�}�ߋT���+'
j_�'�ς�a?����g.��|7b.}m�U�װE�hZ��13H���^�8vS��V	y�℣|o!���Zz}�KMȏet��������m���
����aل� G��x�'��,�����1	���q�*��>bG�%o�,Q�����%�W����=�+��9�w�]s�Ѝ���Q]~Zi(0 �yBL�
�������$�\�mxQ�yk����{�6��y����-n(�T�W4P�t9
�+o�-<۟����dS�u�x5��DSH�����1�����`��%����G�U���\�@Ȫme�o	� � x'�fލތ����V�.���Rg��\�Aiԅx3�K�C�T��L�� �`��� uT�Q<�������F�m�/4i:��k�ݢ	�$i�Q4ɛ�
�H~��	�G�T.Ε�Y���s0��F�����*��X���b�%��6���z�K��[���Z��1����%A�h� 6}�a_���BI�f���3`�_��JM�
ӻ��j?��؛\�&.ɔ�\6Z4�0��ww��a�� �P������?DAa1��C�.@��|܏ѷ<��u��ck��vy�-�����Xd��t