��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&6��i��N��j%�L;*�F��n��kO�͏ٜ�b_5�f_��p-qq�p)�B�&�!Z��T5ݻ�0��I�6g2�g3�s�6�X\�&�aW�
�ґ��0Ura	MO�LO�L�5ǝ��V�!X��|m��y�`|��-�����Q�9��0���wK��wB�=�LVȴ0�� �N�%_u�{��^n<��&_�v�pF�rwlV�OP�u�1��`~�l�Mji�^��-y-�R_�j��m+��5���恲v�5�.e�{�2��ka8�=pn'� ��^�8q(�TpR�`���$�s�g��HB�PߍՔ�罦��C�5MT(��)ą$y�W�Ts��ҤӒ����k�W���:���q�ޕF�+�������5K[�T���UH���|��lC2Z>��&����4�Y7���.����-��WP���[��	���4._��J�����A�K1w��u`/W�	�sȯ��߶Ϯ�Is���zσU�A�D"�!�G+ڈ�߆�G��b��d~/�z#�,���fR=����-u��Yj]Xy8I�~�!���@�!�>T9�>��6�-7B$8.X(�4����昑��?[8�i%��o������EAC�>��y�2��A��n�:r��7��l�K��.�O[%��i���:���.[�p����o���B�f����h�|�|���m�����(x�[fg��hؔ�,��w���7rC�ۿ�m�S�����3��*�)���b�{b���?�eۻ��	�2Z�ማ�
<�=�
����he"�	{r! -�)PW¬��P��Z��8޷����{��@����ߊ8�^E��t�ҽܥ�܂�U��~�z1)y@G�����٦��������]�ڨ�#��r��2�o�5\؆rH3�?M�����%Ǳ���0��a0������4�P�� gH����$�ЮA������w�zw<eʺ<�n�s�m����)��6����Ki�^��?f��~�>��ᴥq����|�շ7"2&���m@���p������N�u�'Bv���u��1w�ٷ�j�i�S�ϳ��M�o�쓻9R�!�G�2�r�^i��q�9�N�i�N��~�mV��)�igr����Px_����'��?8�zA)�?a�Ƣ�'��=l�[�fîƶn��ܫ�~�����(�_U1�������V����Љ��FZ��t1���zqz������Z4��ݍ���c.��4f�Ih1.�5@=q�.��U	3MEʉ���'��I(��r��pe�u�ﬔs06�$��'�bqC��\H$s���`�>H5FX�ip6�E���_螩�}k܁|����Ϻ�������+j��g_S�Α�F��43�uҀsLA�\�F|��vK�H��&/�g�����;(�����| ���k�V34� �޾��k�a�mo��u�yA��U�~ƚƈ�=�4}͸jE n��1������":�,����M�|�c�F`g��@���z6�&0�:\O���1��������ߊ�JK�/���b��-\$Jȍ���M�Cuv�woC�L̨�Q�#v��
�� �Qg�K�Pv.���4��kPoX�aE�	�����I���?뮮-,\�G>��ԆI	����A>D�0
o����J�s@��n�|���dwL6<E���פD��v>�^6S~�g��G��P4��e�rt���m|�]z^�T'JVx�!�"�\� ۖ��6l|_�5�Ʉ�L�7��X"ݬ�w-z��VIPn�v�v��;,��Hӏ��Fm[E4��I����о�:4ͫ�)�*���ٹQ��u��3bj�^Ƴ�<U�iv�.�:��
P�B�"GeNi�<}��}�kM\���U�u���=P�6&� y����Hv������Ω�*��,�5���&`��e��8rG��RvT��͎��I�ꏦ
�6�Z6��xFU���`�>-Y��6����?!�~���S�m�F0G�xrQ������$��=�Sqx��nvpb�x� �I,�0����/��6�4(�w|�&V�,����p���gK.��N;e+n�����ʟ�7���'�wB]�,�1���b�zc�y�>J��gޓ2���n�R?���S�fj����k�`�����'J���\��>r>�!i@]VNe���o�c�}�,�K�t=�[/T�~���*+L�v�ț�3.4n�)0�6�fG��MŜu�**pܕ�=�J\�<,&��t߾lY��AC�C?�4�Y�f�X�05��N�$��d?r���]|��-����)@6��μZv�V��B/i�V�jQ\�rcBG�E�0�3�b�� ����JL��(}��Ԇxc��X�F�)m�	���M�Ms��ZF(���� �E�:C��`l��ܮ��Z����U�#><�l9�P��
��r�>b��h�z���n�-g�lok�f��R��=��mvLk��T�>�[{ �h/"��z�6\���wZ_j@�qB�2��`ysO��&��AF�1.��>iǫcBE �J4���hM)ƴ�Smp�1-٨��UZ�1�$SH�]���w���	��n>�创�|ި;�V�j��;
�Ț����ļ��;I9�ނ�+ ��h��}���W;�z�f>�P�A1��8��Σ�X���/P�m����QD�Q�;��8�k�^YD�r:�ֵ���V;衮�>}��T6E���Y����56�,G3�xY6M�B�R�8d73���&�J�'|�p���O{�p؟-�q��
v	!�����{���U��Ҿ4��r��I��r@�=^�v����X�D̮�z-�K�y������1����k���8;=�2����֝��Ҥ�y��m�b?ud�Ы>/�Z,
�	�i
 ?9&�@=�)��W��[k^�h�$i+�����Яv�<RAR�q"%3�j�Y�Oq�;
����_xQ��U���c�9������<m�u�K;t�CݿS�!�o����
�+�U��[��*?ͯ�$��C�X����ƍ�j��LC�g���X�p&EJ�������۶zk�r�B��[Ty���v���M��R���j�p�CSVl90Z���@O�/�g��R�W�D�o�5�y���[LF�`�6̮S�َT�Z�S�g�W+K�t`w��'8�>������:�;>��߽Q�y��	���ek�I1D�4���V�6"� ��K�2n����np���-�%,�pN�XW�H���`��{���I�=��Ǿ�x��&�ߟYi���׎����y1>Ж�Қc�O���� ϲk��;d9ΛV�����u�����Ž]m�����>���ü�i�D��Ul��	efަ�?�,T��{�{{��!�	~�U�k8,{�9�F��h�<�