��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���c\�esR&{������o�T�e�Z�/��`%�����1�2��g\D"[ޏ�F�
܌�)�u�lg�h���T�Rfc��h��H��H�q���,�+��f,0NUf�ДB�
��䯦�ʒ[���ؚ�ޤ��fګH���3)h�l���F����2�78�^{	N��3��6�,Y>D��y�0��r�\���RC1��*�y�kM^ 1�r8X��<m���#���Z�y�\nJ��~�hl�z�Į��id���*��ǘE7�<���d2����_���w1����6|�pyǸO�Ű�#T�8GNr��0S��{1l�e���N�2���+�WZ�)�1�ĥW���_�1�Z�iV�p�GqRC	� �=g��{�U7I�DP,�Y���K{��F�M"j��'����X������m&�d6B��6V���[��4��9�_�Ϭ�@¢���s�7�b���wYN~��OF�N 7�%m�?�n�~�S�=js
�K�Э~v��O�l����� K|	I�d���p(ThE�k�<V�^��r��<�3�x8>��T3ykO3���f
���O�:o+c�W��Ƽ0��C���	����t���Z���>�8̎q�����Ah=�W��A�����A#����a򯓶޿Ф	iVn������آ�Sq�tHW�Pg�����]�MS��>	�����a��Ґ��&N�g�
����[�0W��i}W���Z��5'���ℛl�������-X��E��U��ɤ*ޒ��㿌�]�u<�ygrE!^�O�A�\K����ꕤ�h-�s�̌[w2�4��q����ۺ�(��5� 2)p�"~�
����4��4ŬKO�c~9hTQ����z����z
��G����~�@�5%B�J,E�Y���oJU4|�vI$iE��ю [&�S_#y`-z������+_�#�%�
�\%W���<�ir`��|p�>Gy�-��G��R�Z�����`��:��!3ʤ�M���wِ�y��� l��$��!1����j;�z�����«i���jc��e���-8!�_�u�}��!��>��w�A��{;3@]���g�d�!�-
 ��o>�I���d9��A�1�G���ږ1�y����[�:�^�O�r3�9��B�U�W9!H����k�n��K�߮|�z����
ל�J���I���0�.caF�Ű��˅���;����e�z!��[��-��˅���܍%O=t��>�S��� ��Dub�z����1���>����������ݨ���[�}�r��Bt3�� Z=��#��JQẓ���Vfx� �0��ށm��sm{����圄�[�do�U��,�.�j���e(:G�i�:y�g����������Cj*)���ۈ��R����Ь|���i8�xB�����!,�iS�>1/�}1P	�� �H��D{��>�љ����y����[bt6��L��%��/�t���^���{�w��>9�D�H@%'d��:�u�b�6�HdUȐ�>��]*�҄Q �N_�^�j4L|rdա�&�4p �e6�v��~���������9}\V�vgp�A�,�[�j��̖E>���1kղ�,�m��T�KHC�|c������[�ո��P�
K����L+C��5��C�t���:�*�����"��i&�2�4�e=4v��i�W�7o9�2H�REBA!ڱ�����-�ޅ�4�ZD�-A
�uJ>��86��A��φIG��]���
�K�=jj��_��LE�9���%e8�3�J�ڞ���r�K��Ivt?�J�*{�������8p��f@D~Oy�?FIz�M�BX���U�h��c���s��~$��x��ɟk9y����¤���E�"����!T�ڜ[�����:�J2�[�)B�@��F쳱����cx>�9�p�V�	5�w�mYJ&4���VTXQR4�+���؜p�~U�����dmDq���ѫ�4��Q�=��]^�':�҂�fcy�Aq��f��0�a48�Sl6Ĳ	���
�6۟FY��a�H���Y���+S}J[z�����:}��l1�i�^��#J��nΊ�y܍b���XD����Q�)��m�|.�%��{��0X�p���P;��n>o,�Jq�>���ɱ�^@�ԍ�����f>��J��5��E�����'��i�!�i\.%�����B<�	Ɯ��	�★&�8,����ʲؾ�C�m��%Bƹ��~�J���b����_7m`�S�X���G�c�o��C���C����U���dJY�?��Ơ�g��QS"�-ޯ�ע%_;2U�^�G����
�u��0��7�)(���X>�b�=;H9)r��۩����m��с�q���G�x7y�̡s#����� ���|�vo�E���]�R�5��Oi�WXn��Z(�LOd�	I�!v�#�� ?�B{Ь2+�����ו���T��`t�W��!4#��6m���N����h��,~� ��-��o����($�J�>l�i4-�٭4;C���[֕�(�������& }�q��)L<sܽ�d�=��S���!h�r����=�'&3=��d��+(��L�E�Pl(7��j�.�Y0���+��WI��� V��2���V�.����%�❇G~G�ɪD�cC���	��țvM�.[��Vb��~Cb�^�lfdXܤ^�.���ޘ�k��,^Z��["�u��;:������>}�'Dx�Tf�pۢ�ߪ�b6,Yh��5!4U�x˻F�O��Y\`t4�����b�x�81Q7�O��y �o�,��<��I��b0���"�+�ٷU�����&R��σ���7���V�#d5�Ѱ�K�_��?�HM���Id�+��D�kd�7�������~�47�T��0l2�r�ys��@7�m@k��=���S0����%w�i�Y����¬���6�\c��U�w�����1���z� {��0<�O6H�h�� 4�}���&l@e��.q2	���.�>W��P\�����4������l�{�s\�;tzLv�]��
��/Js&�iL.��]�L���r ��LK�3�!�M�#�n��@|h˯1�+1,#��' �!V"��e��똭��J�NyIp�r�_"�9��bk�*� � 9IyFo��s����T/�S*7��Jץ<מ�G�׸Ȓ��=��߁1x=�A0��x0A`{��; \��Z��h��[��o��va
n�\wl���	k,�?W��c�l!�� �+�����V�ҳ����iA_V[�C��=�r�,��ٰ���< I�W�8Tm�  �.�" E�3iE��X6��C��.@�I��
�!����럮�a�O�U,o� c߽Z�^����%�Vµ)��������)h�euXI����\7��(����`
o����<��p=j�W���~SK�pO:��!)hi� �Cy*]K����k�� rl�*;HF�27ŏ��5	ՁB1�����c`�� R�F��_�,����V,o
����XY��I$�>����Ii�NIύ`���[۝dp̌���|F5l�s3@�U���O�3���F.���Ɍ�F\d�>��;	$��X�^C�-eⲞ*��%:Ͽ���X�$�F�������#Y�6}W�tEa��2ϳ֘�-�P^D
:�4�矾 *���7_e��H�mN�i�G1�f^���$ҙ��;#���+�O֮���t" \���\��=nU��kn�?	>�p|�$������䁀�^�Z�CV���uWa]_F�d9���L�Y��@�.�s
2�Α�Ɔ���n�*����U��]U٨�5���l1*aP�Sf�}_���mUrܥ�=V�!5Ћ��ư���א>���F�*�ox����n`t]n@�-}�J�0,���Z�����|�x%�̪�9Y��8�?���<-�{fp�]ө�n��� h�W>�$��i,�v�	��P.��q������;Ԃ���\�6 �s h�|��V�yg�]��6$��3�>6Mj�Ot�?ײj�'�A�4��e<��1�gϝ��Dܝ�W)��ɇ=��mrk�u�zK�eo�*	7 ��-�5�>��/y�!|X$�Q&�,��=���yvt 
r�א��	ȰZd�(#v�Uޘ4���E����b�$������ �f�1�˖_o|��3o��rn���TΒ�<�P����X6�B��xxj��n(�!��<F����䁞���ѧ���-y���D9!?��Z��ް�|S^I{GFSz�Zf9��e��v�H|(F��LkF�.^BU�\� ǧ���������ڣ��y?����Q(���r�����'Tp�3�g�u�Z&������s�]bC��?r�3c�-��"X�9�z�p>򻇋�a��Ǝ᝝yZ���S���H`p�o^AkH	��[��R�:��S�kw����h7�'�I� �_�\	��А6ptC��|��?��a��:2B]�D1��Fp?�<��2�"��n�Տ}�ɀ�|z>��	�	��m�(b*
P�Ԁ{8��+��A����q�P�<,Զ�9�ã*O��S��
h��LC��+[�I'����M���e͋ly����M#9tɚdޔ�`l��ӁW��S��`����3��B�MAU%�(��[�f-�/k����/��a��=!�&���-�����|�eO� SRf�gD�z"�	�u%�u���e���
�H���p�IOķ���z�Y�h����s���$8$p�4����ˢ��k=����_3��RLQ�Y�6��+ڃ�Ke����̥U��5ߒ��!���D��6��B�"xD���H�@.�T��V%$v;����M���*��:�aDT%>{���LS�Նw�"�@�׋�-��D�ql�L�:1�D�jn��=Q��ċS�7{ݸz�#�M��v5�ʗ�M���b�}	�C�͇��q�u���s�H�釾<��j�E�߳@2�܏%5U
^YU�=U �ryc��.ih�K���&U?��d����?��i7�����?����i�ݝ�tA�O}�AM��c�!?�;ۭ�0&��*�h��1�I������f�M{���������v��,J�,O�պ�v_~��ѹ��+U0��| w�#[5F���e��fXu��=]��n��n�ʴ��+�4*�6�(�}R��G��p�i���T�m��d��!���ka��9�ӷZ�o�X �ٚ��Y��vj���J�X㙾��s�
��{ÿgJ]Q۞�9������M�2�2i�|*�:��5l�i~��@��(�$
���썎6q>|I�M7/O��^Wl\y�2t��7�.�?�_���5;��Xa�(��S�yܜ)�O��+b#�L�K�2>�!c���~p�?-2-#w�(~�ZPo؃)J��RC�洆|7��Θ ��#�	��h��u[ˬOeݏ@�FT�tC��Uu�MVe&MB¦1Ojw�Fmf{h���_�����<*�΄%`S�l�����E;�g���P���T�F��8��0l�R��׽Ѥ��x�u�u��5C�^�I���uL��^ M�վ�<��A:�E+�t� ���[��!'���H��3���-��lG�^r^d�m�����Ć��H` ۥ��R�0\�(�{�q���P����,Y4ٶ��
�{c���^d�,߇�<��f��C*��}�D�t�Br8s�b"Ū��~+(��"�2��g_H�������O�(�v]RC�=D
FcH�	��L�}*�{��G�z�#N,�_�@�P�f6�
�	�"r7�"S�d9�i����3t�%�"�Ʒ^�/l@�t�L�
�x�jU\��(�ٞM�	B�~�Yt�����Z`�J��{��+ aS8~�-��w^�)zT���xB��N��`��j��q��Btġ�߷�0�5�^��O-6��ܽc2�?�����3{��s$�O|)�v>��:Î=��	�%0f�=�r2�şʏe5Uщ�M�d����x�Hh��� ���N}��g�ZR����$d�#���%F�/�$��6����-�\�b��=����Z(@�2'}����:( �<�R��9S+�(	�gp	1ڣ���a�����xd�G�T��/Nv��=��3j�[�VJ(��)h��r�E'���.��)q{��>A�$�y�1�����8�o�z-3j�菼8J��I�S�������5��󰍎�Hg�1�6��� {ρ�y�>��Y�Ϣ�@;���=��DlNm��^b.�f�!����S}�/�H��P�k q�������	|�w,̴��<��ٳ���z/5����9�������m��ev;[Ҷ��R�_d����\��"�{0���^O���[a����X2�q9�+ޢ��өh�\R��՜�=�E\�fk|���Ҭv�Rj-���дA�?9��dw`��!:��Tz0d�KW�p���ϸ�:,�ȉ����[�ʺ����$C���t�;cg<��W��f0PC�/�-%sb��g3=��e��2���6���X�X��4=�Q~�7��O��n��Qn~�>�M��R�E���*�g�c�"KP�фpgЦ��Ɋ��(ș���%�w$[1�ZY�`��{;ؼb���S��+
�ӈM����B,ű���B7[%���_+]�,I8��o�*|O��kDps���4���ׄ�/�K2�Ԅ��.�#�d�����>ac�ŷ��T._F�bOj�Q���ͬ�pr�) ?w��vwɈ��z��$Y�#�YB&����I7��
R�{�z�TO�)̲�{��MJx 1[���н�l���@���������=�c��-�_U\�.j��&��`Ck8j���W� S�@��.4����+ǅ�s�n�4�3���D8���eGS�<]r�E}zIa�V*���H)��*��{�@�o4"�����xz]0��V�z�3��|8ŗ6�@��_Db1t��vf>�/Ř����q:��A(��w�6��tU�����S�b���,#����A�%b����}zoz4�2RڲZ�N0,��.?h��e��4#$����T��V�K�T���R騵
<g��:�^y��v�or���C�X)�u$�P?+s3/��OJ��l��q�}pvc!K��q�Y?�RR�4�^�n��-�6IT�4�$	��:'|�T*2���q�XHe� XM������5L*b��쭩N�(�@�s*E�Y�k&�al�]ta��S�{��Эkȑ8�X=j�bi��JORn_���1��LD�FEP
���A�a��~謸~���Ԋ>���`~��1#�� F7��U��*�ܻ�6.A�q�i�:��k"v�p�n�O��-,�7
a���Q�j��Ж��yY��rƀ�c?,�0
	a�?[?�dj� ����v	t�_F[��u��Q'�s��ڈ[�<����A� �1�?��rJ��̺?�GmQɅ���t��H`aʀ�")���aZF��Ld0�I�^�H8���q�� ��-��N��HP�D�p���������h�d��Ń��� {����Iƴ��xJ�s57�������<�,�V������[6��w�7N���h�]58v^D6.��:6G�f�
+���(��`�3�d���x��[1�/����G+�<(���Z��E"����Q�u��퍭.����~����ڴ��O����i��-Q�����>xĉG%���p�Y��Xǌ�D��_�ݡ#xKEK�d�~}�+����^g���<r���h���PBf�s ��~�D-��j}��v�HÛ_[xAvv�F������jPi�OX7������I���lNғ���&���h�'��>�����'C�� Z@�^u���7O��=(�h�=�Yg�ǝ�͂8k"G)��![E������N|�?�x���R0K�ӝ���BĹ�N)rqOD�[|}���ϊ77]��,5�A�4���u�-y��)SMnu1"{"5h"<'5)��JGee,��(+�v���o��� C#�zG���^W��.���Y�o�je�>�>+�>��&0f�������Pwg����ZqÚT�~U0���'��1���UJ�V��7�-�M��`j�����p�=��<���1��Q`Y|�+���
�i�oa��D��2��D}�&jm�.�}���Z;�E� ������*�1���Ɲ��h���	�C���;wIO-�1������k�TP|i&�Z;S�1��	��p��]WB���@�Up86
4Z��L��q)��T��+�E��[
��E��B�-�������V�$b��{J�6%�@�X�����6АX�.]D	�1��T�v'���W�'��0���=��э�����d��<���!P0|��˲�#���=�G\�G?�T�]����_Fs���)Li 5^���k�E�Z.�o$�م���C~���	�2����^�s��r�nuǺ�ǬYH ��޲X�<�'繩0�p@a��mK\uׁĝdE���i,u�Eq�*3��6�޼6Hy�{o}i)����b*�S)��gT�dJ���?���$x��t&�3[U��3�F�Dn� T�e��$��w�/�ui|sn� 7���C�sϭ/��R#�b]6ArT��&���d����2���H��
N����P�՞��-��Q��-��P۶���ɵDwآp��ր�Pz壵d�>G����+�`��D|������P J�_ �E�����)M/=����D��.L�ܗq���A	�dF�AQ����jE����ygc�z"��\���C063��G��(6����Xg�GA��w���F�
�y��I�1��\C��%o
N�Ž<���_�a�,�V����3�s:��a#A	�plX���\n쁍(Հ�I�W:�oΡ�q�֍xG(l
���)����ӣ�*�hP^��H����w���4L���&T���lizX�ک�řå��~�2jt{&��Í��7�j2�Q�z��?��P����ߎΞWx�wA �Ch��aJ,_���2���Q6ts��2��;�ޯ�I�yP����CZ?���I}�-6��N��M��.`.�hY���9g��2�l]y��F&M�����J�4��0��7<�Vc[����9��T�m��+����kO�n�ͷ��
V��ٟ�Rm[���&�	�`�4l�3#�n}��w�,���#b�X��ʺrدs�면Ľd�~��+�����lf��p�8�.�Ğ�����'�W &��j�myHXH?A���-n7c��19�r���{���d��E��������s@�f�]�HTǻq�#R�(R��������3wl.F�R��i��d��ٟ'�2�� fPX�� �O����w�=ׅ�����P��+»�c�c�C��K%�K,�۶i��TR�����(�&����^���(˴,T���XOK�ƾ�X���d8��-�R����^i���wU���I�6׳�i� _�fg�2��4j�n'q]Z��" ��,hj�w;ӄ��s�w��񍘰A=fU���/ɉO�L��?L�%�!	[�K�yR�Դ�$���(�	F]n?��e)n+��Wx���iF2ӿ,[ T�Xț�P�ç���I�N���n��'��*�x0S�^�oH��Ք����RP��x�i���������[���Vq�";�ClR%�>��Y�ץ��}	Svm����+��i��7��>�����u�}�C���}("k�j�pu�B�/P������0wm8�s»�	�"8.�ǺD���)��g}{:O��i�����]a����E��T&���ײ���%�1��9�����?h6y�z,�E�_������\�}^n|��N����6v����+����C��E���D�C0Z��PK����
@]9I���I�+2��x�	b�U��H��E���4��]�]�N�R��Y��ix�!���cU.�2�i�k�C�&j0=��"��Q7v���+�+:�L�.Rb �˻�Ph&*E�3�?�:����v�.GJ���"O�yH`�����%�����$R��\P���Y�6�B��x4]d���D-�\�Fon<�xۙ.�m�z��;}��������?��cr}Sl�N��4^G�>	Q�e�H٣/����C����⎀��ĥK����UJ���=�wS'��I1��}�6�|���33������~�����w����Tˎ�[����i�:�r�B�D&#?��Ł�� IxY�+��>+	��3�����wę�E���d��sč�6�	��b���䅡,Tyn�D��⎛����21��;`�>=����k��>�k��P6�Q!k���򫝎Fg� o
B&�n`�P��e ���ǲ:�cR�eġ�}�;�U�*��B��؊Q�(V�0^�� �*�WM�����a�u����4-���e� �g˄���\��[0�Oq�J�!�UX�P�;��ÙN�"������ٍgJ.{�Kk�i��H�9֜z�E朜!iw�_M��4��G��S�/g��\�V���Ĩf�%�ݥN_�����mm4��6~]��yIA|�9� ���ѝ�0�3`�p-p�h`���2��X�c��G��}��;���R��HG"��&�����a����� f����U��d��|� 5�����	�A��*M�3e\F�]=p$�L-)�;��0�NHz�p36�����A?���K��QR�b3<E��5����"2j*�Xj�EZ7u��u2��ڮ�0>s����38e�s�3��+uDk�:%w�ݡ�m�a�8�W�&o�@�q7��i����u�C�˥�����-��4�� �M���<��1$�<��`c��OiVW�孩�?Q�]�T2;/���Ys}ᒐzI�m��X��x��$^g#�+ݔBӤmA�ߋ^�D/ �W��"h�x7�>N�!kh�ǩ�#7����x���`z�|��j#����BK�fr �N�|e'��r#�u����Ҋ���F<0�3)�qB%s�PD���G�����\/k��ĂĮ�CR��s�O9�##%�v��o�a�vݑBFy@01��':�K�t�GJE/���tg�` \�z�%��L��Vk=�s�5<������V�@-�_������T�_2)�=��>���O>j�rsKv��!~k���B��uЛ2�N�h����yՌ�C�y�vtX�%�ݏ7�?$����[Z(�x�1lƦ�����Ex�DzdtG���$�ϩ00��5OX��!�z�i�h\�	E�epNp��)^5i�$��L�3���|�@Y�UK*+0k��QO*�Wň$�� �|��p3�:�aH%XB�����"e&����.�_|����
̙��np.o`�����Xp�ZYU��������A��ۭ�DVi�W��{�F�ZE�x���F�9v�phų�fRm ي+2"����8_*�}<օT����E�cEɹ�������}�š�nvK��<:0���5�w�c%%���I��=ɲ2��Vw�ߪ�R��vx�yo:E�%,�w�h;/���S�K�}�-��>D��ޡ
�r� �q�c	��{��)�t E^2q[ů�BL`��Nχ��BB��g��ͳ=�'�oVT�L�Qc���5�N��o��������w'��ċ�7�G%�X�Y�L�_l��.T�S�U����5䧛���J;#ȭ#����l �_�a��&�r|����sVn�í���x������X��Dܳ@�ҋ�Hr�/��� L(���m�����sy�Wc�*�^�m}�����J�b��w��pNU�|��9�ơb%+Y-z�7�D�
uԧJ��HF-&���&��%�3ޒaq^�?YY�!�	b �'p������0UŞ�C��nG1��D(���4�E�;ܰp4D���η�R4f(��l��r<��A~bB��z�[`[\��0��T��<��n<2����D��<\�@�'��(�+�����\�vnu����)y�%(�1�prS�N��K&�
�G�,����8�wV;d�Z<:أt�2����M��1��X4��R*=��&u.��ifթ<#�[9!��z�6m����vo�ã��*
{�:2"6Z�	���~-$-M�b��δX�۬��԰!�	��<l��������d�����5��<�4���2�W��Tj�(&�՞�hv�&�G��l?�F���e/��6��7�(n�i*���$�_��>�U�nmIU��e�v"���7,QN��"m��m��u5�J�2m���rv����9�е�x�D ^�a L]�"��塿�r�u�ت󠦱y�nV*���}w*��b�y�Y��n),
*��#+y�k���Wt21�pe�m���%�[�pL�������Q�M�R�gm���RH]*S�2-�<)�����_A��qBl�5����`���E-�)f_:��l��C�='��ZI��T�D����=6�3^��	�k�0X�����:�m�5-���P��|�zM[[ۚ+I�#)b��0r媋�t���?o�����M�=���R����F���[�Nf�͘WMR�$*C4c�W(�{���L���NVJr��Z7�X�C�lr*д4B
�j�S�O1��dU�?�r��(}՟ui���!�%W�U#�˘[�W��5�
7�d�,�i_.o2�@k=ٟr�� L�9%mp�+2������WO#e>����o>�Kb���0�S��`
�K{vN�1��3�;g�L��'zAč�ߟ��@{kI~&��;�j���Y��!M�?��Yٗv�
��e���?�HR��5�hJ"v�xgP���g��T�s^����fu��N�ZA��<4�_�!�(錟��;xs��6��i	�o�9�E����&��O��@�C��'g𛮽Ů��"�$W�W���S6�5/7k�-	X�GV_dU�����?�y���h�n��u�N��s���q��������24I���r܌K�IA��=���h�(�A�`�|{�u��{?�,gᴵ]��g�mJ�L��������η�~ ~�$�k�җ2*�W�:��x=y���܀L09�s� ��P���ǫdF,�id�_�	D,�8�(m.��P��W#�{>�y�D���3Z*D͸gY��0K��|ސ�p�{�=i)	a6�)Ժ�5�2��La��v��w�����'��1��c�g��A 9t�w�vНw��x��<��Hyl��m�9�_��F���6P� �ܲi������1���j��!MG�q�.'�V�u��Ŵ�!k^D�O�:V��
KES�c�<e��m���Ti
�L$ZdW���$WTWxVH��1�vV�z$��ʖ��(�Ҫ�b�1�����x�o���c�z�k�]-$��ߖE��;�US�_���Y��{��$}�N��oP7X6��0�v���DxY��p�D`��L4�S������dڧ��_�	%܅��{cRУ���2�L�]�R�](�jf�7����[Z�y��5��LW�<��z)ˊ��2�/��aV���_��KGȔ�lE{�o�v��v�LL���r�ޡ�.��t+�&�?��Э_c���^0�=���`4��\���۔��U�Ž��e��0@�B��-�~*�Y]��X�F��ŀ�^r�A��jZ�����`f=������m��S�;/�u��;���d��3�H!�y8Kө�,=ߩ�|��)���;�o�r��xAE�K�]��7���6���T-N>p�芆s���N��`Kʴ�$w[/�Z����A-��Ƈ����!U���߀I4��Z�/�~&�/}��GGK(3�nn��Cs��N\��P���0�G,��bH&>h��X^Eݧ7�d�:_��SM�����z�]�a�	�"�Y��D����Ũ�PU��<?k�VG*"P]�D�tx�L�'M��]$��ut�����z��C%/��J���ڗ��W��˪�6S.���U=�V�I�)w,V�3Ḿ	�"p��t�ZM���]�+r����%���E�N��M�?�p��Sۆ��}��H��dk3[�8�N��V}��+��0�>�����3��?bb�}�Uw��n[6۳V��U����F��)�2=_o�ƫV-�;[^W���/�Oo����1ץH����}!�V���$�xx����:�"^1�F�W��hDzn��Q�D]G�-���M����j�{y���BG�M��I�̾��Y���T�c�gb�Ql��g����3��J.o̓����A}o�h�v0�E�`�@�:{[o6r�/s�I!7u4��]o�3���ł(ވ�-���M2H�#>�!�V	�_�X{,�X�WU�t|)��W!�� ���,�&�KP^�k�h�/������sNo=�����b%K"�u�}*�Z>���/�m������d��r�X���B?W��Ũ@x"�����E�0�#m f���17I�gx6�7�� �G:�{� .���<���&57�1,�Db�-chT� 4�'��N�����S�P��g�c�58se%�D�3[r�1�K��mV| �Щ�,��\\Ȧ��z�̧#D�G:?�m��.hR��^
.L`����A�pF�}�d��������:֕���Ҳ����43C��e��$R��jB�R�۪g`�����2]9R�h�d��-x�m�q�cG��w�Α�_�⹅6ȆJ$Ǿ�hC�Zz��Y*���x���������A�sojP�k!:�SHwس[ �hm�^�'��[k�g�	���eH<G��>�?�-�o�2���+��^�A�ln�kɱ&[3�P�*��#u3�=>�0a���4<m�LzB�#��w�D��2<�B���4��,?̻��@c{�K�sX����<�r �>jT!|C�N��v�+Y0�HYk~�D�p��TR˯�^�"Vt ��i�hD�gq�0Np�*)ը�����bfs���W�Ű�$�;Qg�<hs4��B���l���J���g���1_R���^Ȃ� {�䔇��Vz#���U��M��8��fJ3�+���9�c�e/$�.T�e�z���er�)ڳ����>��$��ľ���*��wiew�����o��[��b*=���?b8�'f�0t'&wڙ�=�Ӛ�n N��{��{� N�W�w�����=�I�s�_�c�[��yE��zָ�n�b���*|b$�������eX\�=�B<�|��иN�*�ў�hD�����M!��&/��d���U�a�m�JT�y�!d�f�KH�pG���,�(�_������F�R30���	ȮRXb#�ċXtW�K���N�V�Y�0r���s����2�9���sj
����LS�F(���S�.�V�Q���Y$�"]�5u/�3�dc?5�.�����[�c7]��|O&x<�Wf�������:�VL�6f�i��q	�T8)ԛ"5I�K��+���j�����r�}/�HwZ1��,E^p��COJ�PL�����U?���Gh @��RPٖ� Bs�j�<V7L%-r`�e[U��j`[о�ޗ.�#�A�څ ��U��ŞB:�&LQ*�D�XOl�i̛9Cr(ph}W�K�y �;3�@M�B.p�Nw����G9�>,y�n�H�k�ȹD	�;I#	|47���t�!	l�蹥<��+*V<�q02��F���%�Ss�ދ���x��`3"�Öi{�l�����O/~��1x��a�������$'�ˀڟt���	L�����r�����뾖8
s����ح�9�6��r�rfD���s8�P6����	��#0�s�V��I(G��'O#ՍG`�]] ��R"?wG��k2� �QU򈡟K�������`NQ�Q���~"I,Z.���$/E�\xQ��p���><�i�=��"�� ��`7��Z_:(��&���.��p���I	g��V��t�(h[��U������YE3W+3�:hSK�̟�m�F�,��p�w//�xK�y�I�a�C�U�J����t2E&�Y�+��n�[��e^%Za��LT�ܱ�[�Ĺ�|�qv�Q��s�n��L�7�Їfm��f�/z�	���ׁG*���O�B\��+�{:6xe��8������&�\� �v�h�$ٵ rn>����л�D�t�L ��J����n�.'ꛌ��t��c�e�-SN�)T:�jFOY��:�E^I���NK������_�����3wvT ����9%_��=�P�RKˏ^������W8�0{?���V�ur�D�J�NR�N,�]�Ty�x�/匷���.mbYz�u@?.�Ѷ-��o��ddR�o��zb �2�f�W췘]����1#�_��#��ܚ��ۨ��s�2vm�������C���z&B�Y����3�FC��T�5(���_Q���Y���$�W��4Gy��O;n&RB�1�>>*�� 
��9�����]=	G�R�5n�\��a�8
7�ɺ"�^5o��.��,y�X D�):��dGVe�,0�uz�J8+��07�W������w]��*�'��,&"L6_���GM{�>�W4Y�{����o�Ŷv�%G�YX�'+�ہ����7�c[W�z���6��.aU�Nf��i�n�L:Kl���*F�[��J2Cd�lՊA�Ռxj��G�A�'��L�d{�.
������K��C�y"N�|:[�mJ�+8�<���
ӥ�9S�2�O+��.��Z�\o)���v�8�'����F�U=��P�ܢX0�IG�s��S�G�~��6�a ��-�1gB�w/�7i��j6L�o��C_4��Q܈<���h���l���]�iY!���&t�}T2鶓i�Q4�IO���sL��w����X�Qd��W
� ۲�D|Y���J.��.�B�P2�"mh��C�mu���f2�Dd�̝� �&>��}oʦ�h�@v�Pl�3^;�$�.��^Ȅ���9m�!=�ӠZ�~ׂT,�p"}���p�(���p��.(���j�����qm��k���W��,�����"�S��������M�F�B���0���i"�m�ˊ,�'����v?]�����/yB=��y�/q�s���4TT[�U�1R����w��zHc'@����]���3����6o��85�U'`�QXΊ��*�(o��"XBf|A�s/��o2���$�7@f
\�)U3��cD���u^+fUN)KD��E�v'�x���V�\�ߣA/�̻eu��:C�#��3�B~"N�*�F��|� ��Sy����=B��p�4�*Th�;9�'��o�aӷ|�~w�B�6t'�v���I��*<9�^(���z.�""����C!�ˌ{��uϔʾ&��N�)����	�������w�s��o�z��0:p�e(S즓�PN4�~����b�$��0���p!vϸ�U��|�I���P:�D#�+�#~������hǐ�iD��Z���/J,�� �.�M��	�c�>m#���BK����b��q�L�!Գ(m���#�n��q0^Z����[��,*������ݎ�=�%�)�fy�p��vn ���39$�}���R�*���}��]�� J0I����@���F���JY�/�C&^o]=ф�����ߠ/����88�xd*"���yV�5~���3U�YJ�֏��Z?�#������/ǓF�G��w��!X?,��8.@<+f�"��z�o���|�<�L���ޖ�N����k\�M�6�Y��aiOPM�q�ɖ}F���&8UC�T]Jě9�ڇ,����yx?� #����݉� x)*�9��gK���I+��x��hp�V��H�ȩR���=ım�߻y���n�s���z�+ `�
���!����M��E[�tLo=J��?=!���;(�^6 ���%(����nR��_PU�zx��%���4loy)�N��3i�F�8�V,-\��;�i���b���P+���ip��qp��U�R�����yi)������z~R�l��<m2Ch��`C��;����Tۍ�޿QN�Ks� @�/o����x�\�v���AC�C�z�6���FpЧ�Y�f�N��A�^��ώ��?�GM��-�>KY�q@�4��n�,�h#���fdyTZ��(�i�9�5Ul�0K:W���
$}�;/���a�ġN-]�H��t�s7*L�����ɥ*|���B7%�Ǖ�θ�z�T"ڊ�\�����C���O�@�H�5�'� 1�[��Z���<��ٟnC�?i��gI�P�s�ŋÔor���u0?��љC��\��L$ޒCZM��$��83�}A���n!Vq����xw#mr���`�p��#��Ӧ��l��,�L�9�A먭��q,Ί��P��T�az��
v�JU�(�*�A�r8C������D]W�]����^�н�6X��t'ɫم���G�69n���8�B�^�ݵjL�,�Σ��k!I'�z)�c'�}qa�g��у7CiJ&���2�QO�W(5�}�LB�*���l���8�