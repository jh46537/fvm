��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�k*b���f^��g�{uGf��*YO('��`.��7wۅ헒��
�C;;��Qn�������sVW`с��K���Jh�w݃�QKP���wcX����^\�N�A�A�UQp�c���n_lFgډ��,]��d3��z.��b_�����'�8@>J�A�I�=kv 5���
Gh��.	��V�����׾-��+ײ��	�M��:���|:[=�f� ]���s� ��aY�{AeN��'V���p�ܕ�Y+�b.59Nu��,��ZV�m�5��qӄ̻�o�܇X'�g��5��v�@�!�`��K���(d����%�!<a��]3�e��ն�3��(��Q�p�^>[��v�1-�*�� 6d��߭�����Q�ۡiu�Pzt4��fFE����D�8�XѪa�I�w����5RJ��ї��6��|z�Ju?�B��y����xw�+��jp}F��5��R�BgP$��W\~�C�O;;�#N<�WtU�جg�u�K _DN�JCv�/�-�c'�z��!{�R��"F��3�*�C��Hx<%7�yG%2ca��A:h�h�_�(����ʝ�r�;lxjXY�����A����⑚B l�YJ��Cf�� }̸�e}�h��SC$%�eT����?�#�뎩 �3��٭QDYX���zQD	���Zmz^���C]����p�E`�Pw}yH�>�CKu���:H�� �|�櫒$vX��1Ac:�<8��y�W�4]������V�U�+Iv�(�qd����z���t��a;���ܬGgk{�W���qY5�r�,�hK�|���S�ȇB��Ӭ��2j��
)�\����
6}�i��\�� �J��Ya����]\	�XB�N����bZ��$�;?��ǵ�H�:U�Z1�LW��=���{�e�WB���؇�:#{8�l�KͶ��/QZ�}s�ߋٟ 5fBßNe�ժ-��c$	ʋ�.t����h�E����)6����r:m�r��x��Q�	h�R�7�R�Y)��M!(�-gJ]]"J^�> ��V���c��d쏊�0ߗ�y�>���2��V�e}���]�oq��������D)V�yڈ�\��9Ft�2��rO��;Kk���jKm/�ѝs��EE'wf:j�k��:ե�/W��<���՚�`�ޱ��6J*T�����yS5�]+	�gPۢ&�}��q�f݁-A�y�їd�~=iP�@��ѩ��r<M3LnW2�chck����x���i{e�?��v��w�1�����=��(\���� �{1�
�N�pqX\��9t�b��_�I;��W��`4<y�#�ĔyO�J������\�Bޚ9e1S��q���<���������G��e)/ƪ�=Υ�4ď�@n���7���?
b1�.hT�l��th���.^)������U"�����)7`��1e@:D4w�Ԗ���L[��7�_ʸR�`�n>dd�EX��� _�ߣȠ��f�B�^�c��ifC�օ%��G���N��)��i��_��Y��
û���@�n�ũ�umiȓ�� f�hE-��z^�N��f�!�(���@s��*8���@�����,���q�U��)������n,�<i�P���o�	Y�����X �N7����"!�T�Z� n�%�