��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK���ʗ̹����#���)��*��:bE@�+��Q����}h���je��UAM�!�n!�z=��-x��bV���.�Uh��)lI�_�2s�籩��Fr6<��삥9/�ᑽ����g����w!�W�����eT�V��:	4G���N;��r�'٘{P��؆6�«��i{�k���P|C�W]�
�N�B��Oϴ��0��d��Mahtb�f�����:_�x�\*t̏�Z/����C�Hvr�@������`�rX��I4E�m�Y)x<���OjK�h���-��s;�j�Mh8���|�X�'n�9�ai���uC�sJ��Te�ա̦��"I� �1��:��x�]%����Õ�b���7��`� -0
��_r=�O�|��j$����y�����*�Q�P��Г���vM_�����i��g�/��7|��������$Fl��~T�1&͟?u��Ay�n��ִ�J����Љ��?k�SQ*X���t%j�f��������� �F�]$[�����ѾE;)��tK� �6�'�0�s��=�����O����DI��
�	�'a-[���^�PJ~`䖺[���(Ù;'X����֋���>a�)��e~R��V4@:�絶��C�EcN�2n���O�Tp���ff:Q1�n��8������=+P(�;��S#��wK�Cz�=��E����Y+Gkƚ�-�tާP�YP�cn����s��s�-�`.W�l�3&�[� z��	��K3-�P�:��Q�=n���Vp�����(�A��ynY/�����]T�2��]j���� �£����~l58�'ED)�_a���Ε�@,P�Y�w�~��S�ob�3�噂&A��N�l��{sS�$ l�E)��3U�4��J-�V��(�W���L��u�k�*�Tͦ@�Ow���77���].\�m����J�e�]��ǈmy������V���fj����(H���v����*Z��1�+�̶�n��wg�&��2�ނ �JcN&���c�v�������{�v��`�eh���9�_�����}���Q��kt<q��p�a
 ��RۂtAP���YvH��r����J"F\~����֪s(qU�d����`x������[��;3�h�~�p2��|1!I�>O\j�K���X@�[��l#N��C�w��,& ���B�`��ʜ6�#�e�.�ZTMr63�-G���i+Y�L�����<��-�Ǆ{n��A"λˁ��&V@ci8�щ>mCM���A%N&�鱇=/ N|c���Wg��W����A��9��3������#u�F�n�q�T������8�����4׫6c�v�k��~y�>�պ,=9���F��>��5��)q(���ΩH�GH�S77ԇ��C�����h�F廟��ˠ����{x,(HHG8��e��}h�+6�v���}��W���=�>)|	K,�n!���S$=4����m͌�}]�o��_Y�6s9b�sh7�p��#�V�r!~��B�l��U�0��"ǻfnp�i�M����n!�0`m��w�Xڽ*U��&�mD�(�߄���͒Jq{թ��{�� � ��^r�B�sC�3-����"�Vc$c��`�O�A}��ӖU&u��]`^�3�I�[��Tx��a,. �"�s}��MH�y��M}@��Ez7�����xI:�_I�E�̾�M��%�|�ϴv�1D�42g��Egk�?��?d�^V��B��q�$�C�r����/#e�R�c����R��Mv������Y�FYD�@-�Y�6^Q�B7s�T�R+�v�{�Fm�ȥ�5=�"��t�	2~�k�K:K4}�Z���Дr�rx{W�>M9��|�+��4@,a)�����웦�}��v��,ˆ�s��`@�M�v\���C!z@��s�R�ʢӂ�U!zؠ�kW��[��x�L����Ʀ簠�uS��ZK��T�&�B�.�{��Z�ԿB�z�֏"|��,�����	�c7���Đz	
��"����h� ������G9�~{%��X�`�.�4'���QyS��]gQ�������K�E�x���	#2�$X��#z-����2�����EK����$��U�6z��VZ��v�?A��;�M�x=����D�Ғ�L�F���E"���k�E��,�0ڵ��0���!�~T�	{�!Px w���YPq>��5��i�#��������3�����|�H4gѯ�P��!�M�j�|�|@O�j��X�j��4���1���u�X���d��;%������G�m?<�^(�C�Ob��(=��$�Q?���֬)tx�h���"&�z��IPo�Wz�r��#� �iKb�A<���vz��#�0�NZ�
�;����pFߑ�����˯����s���j�?���:�|n�������l�+L�.�k��Q��,�[n��}�(�M�9�����H	V}�x��d�哘�\�Tܶ���^���z���Z�b=~��� %�5������b4n�����$�ӫݫ�\I
1�����|���	��!������3�O��2YQ���	�S��{�,�1
�t�Нy=��Y��/	�|mmb��F��g����*�D��J�P�6	�j����w���gk5Z��@�xY$�b�0}�F�������tg�TD��i�m0pF��( �R��g����V�����4=�cnгܧ�P~:i��h�B��	�
��Qk�q�sS��\f�J��@*y9��}��OqO�J *�;��=�,I��	��W�U�X[�J�t�"��A��ugK��T���HU�iPu٣��a�V,.�B$���`ە��QcQ�F8�@}KG��19~�lʺM)��&�hm�h�	=�#���74b���@󬚳u^��/y�E�K$f�U5@�~È��t<�_�+��r%��e[и����4-�WogR�7X �_���򺏝����t=���	��O������JGP��]}�&_-�v��H��9�����c��������N?o�s�.6�>uT���f$�^+����(t�'ˑ�f�cƨS��"f2��g����e&�w�U�\�����(�E�<Ƒ���;�P=*`Qn/�5	S�I% _J�*�!/Ო���
�;�{���v��P�L�N��%��3O�����&
es���*���d���nF��³X�W蓯3W]��b�WK�Ɠ�t1q�G������(b�V�@��!,���n+�����\�������M�=u��c-�:�+��7Ӟek�y�7�%�F\S7>Ta��{b����M�� �k
C��"��ےO�n�Q��Ih�~�����VN&]��2������&Gcq�XqVgbI[\��E ���'E�yHgB��Aȇ �kcg?��OͅxY�K��9�!�z�|�4�nP�����p3^�c�O��1,�<ǲ+ �R�bT�|�
��K���(���
y����N�{��nD�&��.Kz.�����dxL��wM?zI'����Ge�6���MSQئ�a���9u��O�9\V#���,8?�8:įT3�l3sa�m��4
��b0��5�Ɓ�������4C,��I�y�����q�t�A�|��?߹������ly�c�N�0lek��2�Du����mկ+v�,�@�o` ����"͑����n:Ve�sȁ���_��gb�cE_��A�@~#�w��]y��
7Wо�YA5*���F@�1��=���f� BO��WG뢫���N?� ݂��7=˵��t����Ô���h��0���rZk������X \/_�@��W�J�����.}�?A6>L�)c*RJ]X~��-O'�g�2�R9�0�Ӻ�+Fi9¥��������|��*	DD"�|c�,�ۅ��e�;������@��a����yx��$�������+��p��Ӛ�6��ZK�
�����H��`["p���o�}��MX�G]e����eh�tN�t+�9�/-�	�bP��0�2y���e3"j��;����X��De��T���"B���GC(IC~Q� U���M�:R1�
�i���W��4!�:�0�7�EL���@��5�����7=}��.^���s����u���@�����ͨ`�D��p=fz���p\3Y��Q��l(��	>�V�s�e�Bذ\Rg��ϛ���~���a)�d�v6&�Ϡ�U�!��.�ǝ�mw��C��R�Ș��=��NN�N2H��`�W?v>�����'���hH S.���v�p[��܍N���z�QWM*]L�ŒHm1	;
���?>�g?ۑ��**P����9���L�)H����]��x�ado�O���5�� U�v�"@ߗ,tz��@�_�������Z�dU\��2�5��S�S5�|�ȋi�>
a�� �߯p\����L���"]|r����)
;�?v	��<g�Jj�?Ȣ<:����O�8��+J��wKV�i`���R¡�5�{�_�3���W�Ag'?�Jl������A�����[�K��	^\2E�Y9�
�A���bƐ6*��F��<(��6�9Cm��_dC�Ì���n���X��.�-.L��]��e�?���V=G8X� �ʡvVtmb�gRf�k�KW�x2�V�e�@s�0B@�]'�ϫM8Ax�k���V���s�J��ɩ���U�O��.=���p�8�= .�������7A�.�Y68�f8d�;�4Dc�s��\�[�I�.�n�V�b�M��U�6,����A�j�A<�}��z! ���QZkP���.;h;�p�2C=̺R@�i�b��x)���-Mc����z���e����(بTX�#G-�Ӽ��8��I��@#�P*�������U���4`��+���� �
z�Es��-����W x����惔ƺ` �8�CWp ���Q�+0���e�k�)5��S��R\�'�������x�����a���v�і�~~�ڰM�1�S�t"�9�#ɒ7���P�.a��5���m���� ,�lBU�c�E���O2�m9���/�w����Ma>��k�`��'���
�H� ��p��z��Q��T�l^s;L?v�c19T��C}\"k��\/����CQP�ZV�`�`��R6� XdR��K�,�-��M��Dw��<�۪���	�o�k�u#�y��9��7>�"�UK����e� ��9�ITNeHFO�w�T�=��\h�7�o�9���-�ʿK��&�d�PT���K�����_~��'�����+TK���������ك�����o�c����+���bH�����s�#��}=w'.�]O=#��� ^�3�Gê�>�����X���,�tɼI%�������]5p� b�$t�R�?��Z��Tz��PT�- E<����6�e�8�"h|���� ��6A<��D��cT���O�{�������KAJ�*��
�q��g��p[߽�H�gu0�Yt�W��/�K������Q���>w�WR��:ߜ��7�|��s�����r���x���!V�ɂ�C*d������4����⢜����6t�/���JI�0�����rO���w�qY�Jv	�՟��L�fř��N&�4Π�#*H]�ux;`)(��_hV��Z_���W+Q��5Z�)��-^�|>@!��W:��Se0�L�=�	���V)^�)െS��W=�8�0��+��p#<�T�=�K��.�ղ�L���Kr�Kx�jGc�,FV[�Ԝ���Q��k�n�@�I	V�}t�(�m��&���+`�^��S8۸���.%l�J�km7�!��_�EadEsy縢u`�d���гP�{��|�&l����i�qo�����T�>�x��"��'!�����콖�9)Z�ʹ�È���ն�4�{M�_Ǟ�k�fcCХK���eG:��SF��6�z�L�#F��p���9@� �&�)�7X������W��!��yJ;��lT���׊a��â�L �Z��ï�����k#28=i�j>�_����m���88&wx��}>c�����&s7��Br�g�n.�Q�13~ ���}�<n�?h!��5�F��հ����^͖�ۼZ"g����%{6w7��T�ߐҶ�N���%���1}�"��|Z���;�*�W��q2"ŗ��>3-)I�� | q&����}��c��,�%ii���B�p�2K���3!�>�r_Ix:�����Sr���O�������}��>��6E�(V���}�:yrдE�J���,̉��3����m@��o���k�˝�GoFz�ք���m4j7Hy`�D^<���䤡�e��b]�$n�����򂩔u�t�W���s��5��!V�\��`!Nxe~=�_�6N'�c�C� Qz�4Kq��X��ٲ��d���-A?�>���,��\�4k/xS:o��5%xIS϶핔�O�2A�,)`�ͳ�xI05��U�1;/R���i��Kv�c�
EC�����-f�����&��>_��D��F�戥��k�sDO�����(1��,A������;/%��B K(��0�|Jl5���~�
$h���CJx�Z��uxjj��wR���x�A�P��k��|�L�ǋ):S0 ���*_�FW�J;�E��A�м�e�~U<N�]�D�:em���j����<�+9���,+�3	�̞�А�CͅW���^f��9���e��l�=��8�;��͏��I���1s���~dJP�7		^7�pbt�V�ۉau�:sh���Dv���a�v��-R���h�1�;�����힧I@��Ə~�-Y�5�Ky�w:�ĺ+v����W��e�c':���-��b�h4��?���f�~��ܛ�����ÈC���+�^�?����o��0L��oW�B�v�#_���uTS ʩ�;��N����P�0�w+�ϰ
;�Y�qi"kf"$ �����f��?*��c��W/��<�3�0�����"Q������ވ����*x��~��;.��:��f"p�An�0P��7��B��Q:�5�dQ�� ���lkZ��������AV��7Wy�Tp�}ydE�@^d�@�}&�_4WO�)�5�!s�'o�Ht/�^]A i	��@�(�`)�r������ �U���9@9	Yeg'鼹2]臎<zd�5��P�E�3v��\��?����H���{�^���ql]�o�3"Y�n�P�b�R޴C�4�_���u�,�-�3��0���,̛`J9V=�q�ř��?��Z.l
���I"��� �S�B����"w5��=s���5���~�uS�JG��0t�kA�c���mԾf�C2�Px1&-j����؏���V��}���u�:�_o8����j~'���n%k�..a�%�1�pi���{��!�]��}���-*�o�hBى�>���r{7]R�k��:�Q��g��W'��W��\Ad(�X�/ ����C�,��
����ٚs<e�Q�|�ŽOѰ��Vo9�wb�?A���=�li��WԀF^���=����fu��xD�Xc��� k�MX&u(�mOy?�A��o/U���T9n��@m�����H0����J��Z��+�}EO���>����B�V���N���/&K�]���{���8|nA��ұ�P�]��x��Dɇ4�ubAU�R�����t�p�+?j����u;1��^�(�z���mD�F��w`*�]��9}�D�Ӝ�뀨��(��������)��inm�}XpSc�?}�*G�5�SDI�].�|�SR������&Π7~J�"L$�ѵpB��?�2�@���}�π�B��1/ޝt~e�+�pę	�k�현����z@�*8�M�G6@g���C�9�z�]�n��ZT����5�w]ٺ�o��Oŧݕ�@����;a�Lem��>�*����X0�6�s*WD���3;B
B?�lR�ry|����B5�)Uy溨h�Au�k�J�N��HKZ��}�I�[d� f�V��t_�4����8�x���؄��	Cǟ�u�RWN�պD�1�����D(�`#����Ec�˂B���ƞR5��K�=��0�^�� ͳ0UdY�i�����p�b,�Q�H��D	`��$�Q��&<5\!2-�v��X@���N��|ӆ��6Q�DAE~8�Dd�[�ו�7ϥ<��>?��D.du��w�`�e�$���z��/}/���������o���+h�%����d}��}������|)�j?aO��'������~k�1"��)�x���!*�+fŀ�\* �t���X��:��(d%� P)ՇZ����V$5��pb��(E���<<F��|9�*��%aZ���(��<,��F^er���OO���+e4�4�&�P�dc���})���&���\㩺�"�{'2�c*b�J�Ql�;�]}u�]�O������1",'fV%�����7���N��X5����s� YiZ	u���T7�i�= Q2����f�R����c��o`}����XtUT�FL�T���Ήm8N�+O�R�\YjLJ�h��*ƿ��˾��t��)�ƕ����Ca�ǵ�f!�g�e5��9�p���H01x�d�sK���3e�Z�j��۬����Qv?R)Z�Ҍ��P�j�:ކ�d�%�h��oeY������i�y55�_*c��ϯ?�Q)�OvA�E`D(�A1�6t0�X���3�[�Y ���R���5���2x�-e���"ޱ���Er��`��mAC�#1�ɍ�zTR��z1��r�7�O�8{4���G �4�	�+�I*�����x�f\OaUڐ`�F�[�[�BOV�7O[}�������f��� p�"�p��>rɺݨx�C5���Ĺ$���p��1���?� ��u��r�Vyd���)�T��*Z�e��lT=t����H�Ŝ��*��3�B$Fӆ�V���sű�̤�~m�L�~�_3y��c�8 y5��m�¶��pq����vv�;�9w���B����5��/T�L\����Q����"�x��3�*3ә�����UIF�c��4��"���^�W#2?,�!�X�b{�
@hs?�ñ���p�������"M@w3fq���+�9lb�.�_��T����ݟ�)���{���f�]IU�Ν�
�,�Ru슍����gj荒�/)��A.F~͙�� �&�>��A�������t�+�T=.��3-	�A|���+W*�o�j �<Ћ������l��_n?�J<z��V���
�A���u"r�Xą��8�o���C7u�4!��^`�G�Ji��<ܒ�0�@��0���Ha���L�q�K�	��OCD�pH�ߘ��b��N��.���+k���T��b��WU��A��D*�Ց�T@?ޫ5�\�3�tEr�j�K��!~y�m��w 	3��8�!����g��}�����am[r�e7F���([�,p��I��:'�!�X�A�Kq"�M�r��]��[���t�"�%X�Y5+���
B�ˮ�1�����6C{!;`�ܟatV���0�~۶B"��z���5⳽�Yr�6#�į/��� �+��^����j�����7�y}R���GdG��$�O��ȑ��HQFb�_ݹ��<�4��nၴ�9����@�����.T��'���z�?SCC�2C�c(��Y6�P S�ղ�M����n�%^E�M��WBʅ�Z
?�\%|��Wplle���gU���|%vF9�Y3�h:�Of��y�FV�STRp��%�MG��fV�?	������vv�f$Ǽa�V.���fR�k�i#v񜓜��_F}����7^�tя_Ԁ#��dP7e���4*��F�kw#��g~�=Jl��E6e�Rl�e<����/.	���h�fo�|��*s�g�Ա����H���Y8~�\o���I�b7Mw�H�_�ҁ��]9p�_�yA��j�uK��'�=w�;��-�T]L���f�e���V��5��;7�*�t*;W�"$��eE]7�G�*�U�'�E`8|0�lB���ˌ|D\���dI#gj"������㳯ɦ|Là��Y���6.ɕ&bX��S����{�S��49kȣf1�	x��,�����v�l�.u���rڣA`�����˓��1_'1�J�s ���sea:0���L�A@O��jĞ0�c<��C����һ̺��A)�p����G��\�/�	�]\F�#�������A�{����'�AƼ��hI���+-��y��Zç�
W��d�0�I�\Ovj�YtU[�P�;O�3��d����=�܀h�vC7��eC�����V1-;F�1)�;|��	������v��|A�3�X������G<{S����|e<���S�]Y������!z/�6`)uܰL[��9B��:�ق76ؘ_iGaz��0�.j�U$g>��9�l�_��5��8pӊ��f��c�]�Kc8	w"�mb����B"xI�yYm
3����H5m�^�WFT��C��6�8�u��p��o%Gz[���v��xjX�";#p�En#?w�3z��J���)�+kw�R�a�iQ2	��0���Ӷ��i��tɼ�q�P�����Q�W��{��å�0ڝ<8Ie�z�L�Jb�Q���tE�]v�\&{����3�:���^��u$>sL	t������@���'�0j�Q8��aY ��,����B�|�i ػ� ������y����]��5��"@�%�`�m̸���(��Զ52)�Ƿ�͘ ?��B<�Gj�B:��,�.C�+�8`���R��d/�y�fr*��e�Ij��Ls����@Xk�y���:��-Q�=�U�t����(1��+;~���M��VH���uG�"�Ȭ�E��A��tXby�:~���66E��@%�W�~E1�D7[a�/�ѽ��,Աo!n;�%jޚ�"��iJ����Թ�^���ɯ�w1�1�,PeV�Zd���5 	�=
�Z���Z�������Ѥ�RVӴ�F�U�bqnv��N��߻���s��v;�v�-nI�"f���.L&��/咮���ؐ�q����'x��8�q��mBƛ0�Ad!$n�M�1�)Q/9v�3�~���,
��!��4��B<L�>�E'��N0��r��6�?���xF�{�G��)���n�WuAld*��޹{��-$�ڸ�vr�6�s&���f�j�/Sv�� rZ�ĭ�g��FI5��XĦ����b{�xc5�D�e�ɬC'f�t�Y�{qǄ�ZDmq,5��LWj+Y{�b��U�B�t�f����F@��n&��֙.x���>�y��+1���b��U��L  ���R[}s���������IK��p(�w�ș��t��Nj�P�K̄��������qFp��Qd�B�K*2Y�!\����1��5Gp2[g3�2�Cp3���Ry�m�a���/I��t����y˄��ӜG��G����)����Іy6��ʥq^��9����w��HI��|$\~����V�m��ݒ�x����k�=�R�1!-ZF{ ��s���9�lp2�e'�FAP/k�5�9%BН���_Gm�V��X�M�ub�\�Bw�N�W�z`;g*�aG��ѡ�`�-S6?�Q޳D�u�ԕ�o����2�w�`��������j���IP���K�IZ�i�G7��QVGf��|!���ET��X�`��K��~�>�Ǡ�Z�9bjq�����R4�S�S~��> l?��4~��&�L���32D���^�)Z��s�nߒR��z��V�g��o@#��ޒ��)ڶ������Rf�������Z��VP9ٜE~��>�S�aH��J���k/��(��`�YE�8�8?��[y��.�*+1���"��o��v�b����@~��#��p䕚A ozb��͇�)��� K�����(
}��i��V���	���s�)`0[�2#�K���4Y��&L���w�)bo,���
���:-�j9P��b0�;8QF���]9�c�mm~H���'QG~�J}'��ƽ�=#Ȋ�ӌY�rP��  -��L�k��4��vC��0��|)?����-��E>|�9�cΧ7z��Ov}�����L�F���� ��R��l���m���-)�7ޝ/�w�HO���t����CQn�y���i�Y4q�kB�	v.��M�L��@D�+�X��~h�aQةz_���%��݀��	����A����.㔏��mY]��r�bh5Ī�z��|˖u5ApdI-1<FTq
���c��;���г�u�8ՀF�����S5I��2��0eu�g�c�"�4Z5'i���hĵK�'�g�<a�����|���a8��T��"Q:�4�"r�1h���y��M���7_���.�?�R6K�[{1ކt�[��e���FC�v2J�� �cXΓ��{��!�ǥ�.�aTEp3��|���^�,-�e�	NU}��뽸���]�+�r걧��F��%��ń�*o,���	S�_މH˷&D�IJ�N�%=V�5���=�������m!�^�VS�  Y�m���۹؅
���b4���9o��(��������������MS'3=2��˾�hNC NBE)�;+A8Fa-���P�ъ�+��w�!�?�"�e�/zMRm=�tjO�ڤʠ8l�^�kĿ�����1� i	ק2Ɇ
^�:��MpY_F��hf���f�?W������ ���+4��4�c��wz��*��+��oie��L���C�P�\�C{�*z��U���T�!w?�a�}�� ZY���b xl�:\b���#��9�^M�A���ؑ�x�l�Dv4AQd����[5/���|�qK���v�����8��``8�B�6$�!AoR�ު�]T���M�	ʠ)��m��QOZ� �^9?|~���󏽮N-ǔ{y�W.%�{��-�]ȇ��g%^D�*�ZD)��*�)��p�\e��ۃ�{���Q�g�l�6�T�Б�*�okd�*��;���FI���!���	 �M�V%�����т�O��}!��T�kg�_&��>兹lW	Og�����7�j�$q%f=���=��$�St�%4�w�w��_��$m����$���	�����Lk��\����Ϝ��p�9�=kH� w����\�k��׵�"�	��� �q��2e4-^[�����O���h�5���
��,2u>���$Ɖ6��l��Q�(N�/���]�0�e�B��x��F�.�Rć�3�قi��8ƨ-���i�v��g
7k,�±�	�.�4:|嫵҂��.�B�`��o�rXq|&.4�c�o`����e5�i�\��3���5D�Bn�c�(���������Fb`!�М/x�if!�f0���r<������[�PD�z΢izAI{m�9�N�m��,/^;�n��h6��V'�!�@g������[���Z�j�J"qR�����@�&��1Jx�$�=�t���(�doD�b�>����H�yX�Rۻv�6��of��ř��,��i���>ֺ�n�]G�"=j�k�cͨU��3%J�p���(N;�ґ�^��rBƲ�d�� !;����#�.����֤��!w���'�9�@��s������=.Gx�SyRf�$A76�����O�k����Y��h쭲7��i�w�.ȃ6z*��(�
=�C�7*PIģ�!��cd/V�zf染�
���IK^4|�Cu�\��p|D�.�Q�t"S`�S�ڮ�����6Xĥ�!QV��v��[�0]lR)<��*�8�<��h�"�#�<H�J}g����Y$v..��{n��![l�l+ؽ���,� d�J��!;^jDu��.+�cN�F!a|��eL��h.~�|�EyOn�XL�_ܻ��6z	�KBe��[i����z���x�Mg��x���Ēi2Q��������5<|n$%`�f�;�^���,�}/���VP�[٨�T2�˧�o��|��r}��MV��`9J�,�/�6	ܻ��wd:���$`��G;d�!9R�x��(6�ҿ�>��7�Y���5R�R|h����,�y��f��g'5=2V���GI����ҴF��KԒ+Zm��3�̷g��o����~���v�����[h������3�:�X�
�i3d�㽸BB����S�υv�c|l ��:�A��ŧi�xNX��f�X�2��U����|X�h�D�/�j%n��
���aN�;-J��y� ~�dv��<�$���x��m�7{r�������Ta���9������-a�'_���?��px�bك��1�r%�Ƙ:#vq,�R!�(8��(7�S*8[9�'�˷7���{�FNR�B�u�L#���� V�9Y�� �.m��l�s��8w����{ar�4d���H�|O��!΢l����&�����ҭ�&b���w����F�X���h@��(<9PO�j�[�6��2XiԲ}���f+E��~ ͦt������o��Z�3,8=��-[Xm�|Cxt~	7�~ՂaS@�UDwЖm��
g���g�"�Ʊ�(��͏R�I�e6-5�T`!}ۧɇ�9��'�&ϛ�[=��F+�����`�:^Ѭ.+�����g|����{�� 0�_��|�9�Z�+0!�p䋸|�\��ڣ�#��	��cI��ٟ�+Ư�'���ȾH��PPtϯ���|~oO��V�,T\��
γ��'"w��&��U�i.]�ƹHT���]���{h��)_�8��'	1Z�;buo��^�`�>�O(�YscP����3��D��P}�2v��~���l�D�L���t>!�b�� �2h�\�y�9x�EAsM��8���^��yB�x��EԣR5����e��b�o�zD!{K Kr��wp�4����Rz���c��G	E.�:�ṃ��*I�	�8�°�P_��0���
}�o�R�2��p�)���j��ɗ�{��X0u�6�	�|�#���ܡ��
,�o�E���Xà�� ��n
���4_��I<.Jh[�ӣW�������B���z\�q�J�J
���>p�[k���b#��/��q�n�1=;��BT��S����n�`���?��.%4P�:��*������X��`����E��_���~K�N�Yjm �̲9χ]`y��<�/��kt�������vB�j-:��*.���CB�J>3&ͨ�c�q�LĆ�8H��v/��t�%H�
hja#`i��y^����0d
�݉�(
�3z�w��Y���~�*Vp�^�&��|[׀���j�$$��ɡ����+r)��)�r�ꉿ׺� ��̐E�ᯤ'����/���_u{���HFv��t�w9at��6����N^��/}�=y�MbZ
+�u�ဍ�l�C.�0��K,nBm�V��e��Jf�^޶1��഑d�{<.��'D]�[S�5r�x�0
;��$]XƁ���f�qKl~��+6\I�)�n�?ͫ����=�^h3�M����IeP�p)�4�����U��v4u}�)���{6�H4N�����Dw�͵��1<�ž�_=�����@�rO�`T���������\L�� �Xb\��,�sCX�?LU�-t�nD����9Õ3Z�^��j%�¤�=�1���`ؐ6լ�줇���-4A��m���	�Br��4��͑�cd�:��łgeN�*rg��?�c5��ZAB�����B��N<�y�҈�.�,z;rw��}�Ǭ��rBYZ>��P��w�oe���3�nܬ���%�';���F�ӥ�"�;����3�{\�2��=�3���_�_B�l��6xT����}���$G���,e��T=�M�]�s�һd`�|�?�u�6��sXI�6��ɷ��?��:>G�cs��J_nqi㍾�=������&O/�'K�toסO��y	Qa��V��yLa=��p���FA���z�V�x'����Ǡ$�<��y�w�,:������0P�IŁJVL��>J��4��aF4���b�$T���a����sRU�B@���0\����bhCCF��\c�.���K!q�-�/�3�� I��:�]j�@��\�Z��U"��>�2 cGmE����5��(���*�]�2 X���s�\:�P;2�M1NT�����~�]5�vDb�g�q�^~�x�Ɋ_F'�C�j��ڌBmR�ix[׮3�d���@E3����z�m,�E�,��� $�F�.�EŃ��&,2�
�T1S	�� �q�?����ʒmg�袖 'c
K�]���j���b3��!$w�Fx����C��������#�^�$�I}����h��e�0G�L���F�|����"o���,|�8���$�����=J�ۦns�mn��m��Ǧ���ڢ�#��P�E��6K���;7�!\¡����+�F3I~��_�<�4$�L�WN˘�*�#[(|H����>�uĪ�n��KC �� A9�Ch� ת��,���.��i���kL �0����n=1!���]�	Z�Y���� ��oBXI����M�D�_�ab�]4�k.�� �ґ��G�E75I ]k�ǆD�f�+9�Ƴ��i�;bz�H�F�,�Q|������"��<�3EX��*�.v��ҋ�K98�<�fW> i���-$\}Ru�GB�!�q�u��u�%i�J��X�	�u+Bt��#}R������ZxM���N"K* ���x��.sE���w
|ywk�-̸�!��.���'l>�|R`'��p�n	��Y���஦�)�����x����q`��m���0�`,
�����&��ᮈ���Ul��wK�+%��6��_��5�D���FL�+,E�B�/u�=DQ�S&B�}�Q�Oɱ��SA#z��	%$��=�]�������+�>˴i&F�7�΁����Z0��VC�K��(r�Lܓ��.�� 
|%���ޭӒO8�91S�^�14���G^v���Z���K)���sN�S��S��c�m�Y���R�8o}ie�U����W�_��P�����ExT-[���#��?�@�uqG�mJ��fjRC|&4nk�#�n�q�
�E{*��5�5��bX/���<K��!�ڷe�T����MA�U��P۹���Q�ϊ`��k7ٸ$��E���o@��w#@W��>�z��fD����X+�Xs^���ւ��ݮ�H�� Q�Mɺ�/�J����xA�cQ�D�|�i��Ӎ'����t�m�®�D:>M�Ya�ʱ�3	zu�0e��}�~W?���E�H�N*ƢN�\�����L��ى���1i�M��ⴒ3�	ޮ��!�������J��"O��YH�����8���Fs¼d�y���d�'��ض ��1���Ϊ4V�4�#�^��]Pg���m��!��r��$���@�zH�9%�&ɖ�k�8�D���Ӷ;�� �R�$��ĸC�1��:� �i�:���տm�W@�"�w�_���-eq͠".@]P�s'4�C��Z�(^��K�#��+P��^İ���~����\���W�x��g�I��UU���J�<�sp
��'���n�:>`ܿH,:=�
[n�ҧ�G��e�6�4X1�R��U�x ��xo ǈ�Q���
o$wJ��oR`.�d�M�ǫ@j+gMq_5w����ȳ\��^��㜦M�G���G{�����׿s�S�#)���cY��+� �m�Z���]�a�	�x?J�5E�mH��*�>G�1_Җc
�=��p�I�F���0Wې��ʼ�o�N�����F�ߏB����kۛ�d�ٿ��E��I�/����
�� �;�j�}wְ�-�a����w���`^����1�`Tf���aJ�=g8�*�[||񦐁�	�&���]����x|��NM6��yu�ciF�c��]qq
���)������y�3��2�S�p���I��_�#E3_osq���%	o�
1޾�N�-{qk�:y� _
	����ť~+����CD2�v��pʲ����3������[(NJ4�sA���$���&��)�Nj�����o��D������g�����U����3"|f�F�Y�X54�|�5�^�~���[f.��g�w0i��Ѻk�.�?)����I�1��O�|�M���9^�X��|�u��Y��PZ���O(��w�_ 7+�t��W)n��*Q��,����tx�}���`P����襣]���Ɏ�&��2�#5��>}�8��Mf��m^|��]&\�)<f�3�|���Et$	7����ȗL�����7�nK��/3����f~��3W:G���2��N������\�a�.�
����;7�x�'"LT����=��/7��I�'2�g�j9oU50���h�چ�p>T5��LZ�쬴	�@�Y��.�,�[j�����'�/�&��(�X�A=L�ub�mؠ�Vӕ��n�3�]L4�bG�}�5h�Zi݅���/�g��F����V��ףX�+Zq�)��g��~� mqm�qQ/��� nCH�iT"G��B�c�(�w"L�h^�1�RZJ-6�J	e��W?`�]����$��5&��`@�p%�S��Ʊ�S��P��#rȇ̇�U�N���p����Fj:l���_G�U�FG�%��B��*� ��9^��7��ۆ��vo��t�[��Zdg�L��ֺ��ʋJ��BDl�.i(��ҟI����g\9iy�I�W����`o뤜vwK ��k���ᴿ�n�Vx�7	������#��e�&\��M�͏ৢ~���}6Hb.	���3TbJx�O�gO�<B��r�7փ�"���C8!�N��kQ��5z��x��Zm״%���hh�CV�Gg&��	2�b�S���g��p��]���C�^��gm�W(i�q
 M�C�v1{ |��~,�� w7g��ϹZ�Il;�tЛVm�8'ZV�g�}�\�|��y$[f�@���W2�;�]�:/�����v�ǂ�^�J�M�dy�\�>��kXM&Lcg�аH�4>�-��t�`��ӳz��c!�!y�lз):�&It|bX��a}��>?;��=2CF^�N��<+��'X��=��k,�M��������p{��U�����v?�����@b׋� �c�G��n�׼N�p-^��Ɯ��:`�Vo|^_��)��v�*��."M�Av��~Yrq��p�;g�..m�YUKј�2k57|7�޺6�]w�]h�i`��/2Rb��'����uN�jqd�["ܸ7��6(}�3�{0��([��g����7IY5��'^w褵�	?����cS��D���P�vY�)�V�C�����a�����e�d;��_�+�%G����8��7���>�1�]��ӵ�F s�"���
*�N�J{7��,#�B�;/��^q������UZەs�4� b���`-�@GIJ���SFӴ�R�p�<��<u�d=4u�j�6:p{��lMu[����e��Cey���*��G��f����w�jQ-Y|p'd�f!W��\BaE6��
��H�Y��_�,7�fY�<_ܦ��Eh�8Y�{:Е"Y�����6;�7��G�^�>=�����A��4�V�8����~@�w�~�si��Z�CM+HZ�ҍ�p:y��Z�o�In�
޺�{6�	���֞rg.I��A�"�@��hW�2�N~b�d��|`�,,x�?W�-���mPp��w�E�]&�E��ך1��2TxX���^��Hm�N:�83���?�x4�
���=���n"Ɖ���w+�jڕV�OQu�'=;��V������uޔ$�O�U7o{Y�������;Kܦ0׻���ĄK	ۤ�kl�� ��5l���ԥ��`�L�����ԶJ���v1=�b7�����"�`H��@�Z���"Q(�k�C?o��^�k�_z�s��9b�O��ɸ��FeE�'��F1���ٯ��}��善B�� *:��2�J��u�;D0�fQ�r�r�q#��5������S)��j���H��n���RL�ؖ��qPBf&.=ԛ���ưf#�0>Ц��w�����f�V���q�^!���z�$�e���v�UJ��ڋ��f��W�-�k:���>�q��ߵ��]�'PH��/���]c-F��"J�g>����՜ "�V�`%�/ش������%�l�if��c_d2���Ӱ�g'�]�)�R�.^ %S'1���f+d3j�i�j-d�� ��E�x;�sqc�E��z��8�=���tA�z�0Am�S�:G�oqJ�omGv�f���L����X���Ī��t�C>v$�ͶE��'7�1������Q�焞0��x��c �V�c��J�w4s7�=�}��+�}�>F�hF�l�e�mV�k�M��_kU�����*r�qnR��&�� �n��mq�Ѡ�m6�	l����M�s�R�����	��(a���q�7.M�p5�]�P�&�$`^C��D�"��Ni	��Ə�|I��2�j2�����=��4JԼ�Ѯ۱�ˈ�����ECz�a����]�lGTt㼰�����T����R���	���I�d�ApD��긎ۀ���'�ԙ$6�G F{��t�i��8��=9 W��B
�z�y�p�e�x�qҤm
�-�X�������i��֋��7XL4�,�Α�LGa뷒�܆�z}-@ړg��2bK+�p6ŗaA�T�<�m��ب�1�`>95��I�)kKmE���>�7���1�Ou(W���8wy�}>����x��v�=�fh'�H���i�r$�Fc>¿ �ƊZ,��Xy%�@���K�|�����>�5�L2�(o�o"���=�� �i��R׀�3��I9cjv>�:�M+��ذ������pN|�t ����,@`Y�wXЎS4��Ad>�Y>���t~�����=�O�ngX*��O�;�~��&�Fo(��2:e�Z��~�Rt7>�=wd$�g�/塨v�)��I�I1mG�􍄏m/�8�K��r�oƷtG]J�jT��/�Tt2���At/Gp���>N�.>T�b,�?��H7)��~��a����J��=�j�XW�L����)�%Q���K��V����GO���lw�.���R���= 庣m���+�dc�@�=(-E���N��ì?0 h�k�	����j�"��
d��^�*����x8�ȃǠ3�S=�V0�_���6�,'��u��<X1>��������F��F��;�=j���Z��~_[ۧ��G^�z�i_(�
�!��F��Z��(��I�f��vO�:aŷ ��"�|C:'z�
Q����s��-%3P�A�@�A������,L�ڙ���r�-u�m?��}�7o���L^���:i5��Ƌ�3�JM���G�DmT���f�i>Y���O�Y	ޑ�G,�1Ia�0���J�{[�{v��;�H�pc�(����S2b/���i���&�0j�b�◳�%{�3������JM�|��foWa>���x�ɨh,Ur��?�_;�gK��]k�+]�OS�۶�=�Dc�9vX�u���A�Ў�v!I��E\����=Gb��A<��� �a�(��ґ�A{��n�&���]q^����XݑZg������B��f2���_J�el{��N
H������G5�
�|��MD.&Y�P}ʲ��o�m7���prz��[����]����+�w��PMqn��Y� ��/DW�P�6�T㞑�>k9~Ґ�5L 
��h_�BUX9�كҟl���lFG&��=oh����`��)<J� ���2�T�^z?�������r��z��n.=P�h������%����9��Z� ;�A7̏�8u�`	�g��04P������BG��0�Z�5����Ж��k�t��@�[(��!��*?�Y<z� ��H���6�eW���H ڒI�����$G]�Bc���W��,'esf����`57Z#&KO �If��}�^�ʈ�O��:����M�J�¶U�D	�G��K�#dx�Ǿ뷥^lG�j�S�B�,e���Tf��4?�f��z�.��rk�f����p\��\���o����Yo�D���(�Dt����b��O�YD��+��ɑ7>�Q�Ѵ
�-%vU{�g�]�&36�5f(��������c?�+qPг��AC�l=߾�:��Z���h|�\�C�K�	M��Km�⺂*F���H��G�}@�s�AMԣ�獠���������C�Ya�Z%i~wdh�v��gKm\��
4af���:X���$����z�AzZ�_��w�[҅P�W��ۦq�=�4y�l�ҹ4�}1J�H�p���*�������긚Îa�8؃鬎k6��Ho��D�{��s1z��޵ۄ��m�Fx3��[#���?��d�f�xһ� Z�;S&m'��(k3>X�I�	�{,��Y�xq7y�;�@��j�K!N�������R�5��6Q�3��f|�[��Q��
G�6��D"����N,̙�����ǤP'�z:w��bG\wz4㜥�)�O5#&S�1�T�{Nj �`05��2O6�"A�,���r��2�? Ծ8 $N[���Z�U$271���(o��^�����'�5�7T�Y�o���v$^����l��[�0��R� d{h��|�4�41]���c��x	%�I����7�o����q��W1�&`8H�a��� �|�N����}b�1^���W����ޱU�')q��
)Z�A�õ��O��T@ԃ���ʿ���$&�S0��ՕM;��#H�L�ed�
7~?4�3l�	��,�����;k�ڂL]�vV,��6Y��b���vtmbʶ����^��H������Z�����{�b�����r,�L�^'�5	zu������Q�A�C�c�{$�wS8"Z;@�&�C���td������|L`��%�b�o�&�3�sE�Q�x�+�KK���Y��|^��;*\�r����y���Sf�^�A�`}�͘Y�֟��h�KN����G�z��F����pH���
Ґ�.3����G��O����m}Q'�LL�6� ��h��� �F�
�˕�b����Ŗ���2?�׹9���z!Z�)}�߽Y8;+�t�K�X\�NI�V��Yj�:N6�2�dg[��^-]�ӗ����d2�\�d	�wfE.�Lo/�Zn��支FJ���k����v����`�>i�j�L��W/L$��.�+�/�$y�!�ԞC=�����w,<����U���/�Ji�	����'J�mMӟq�e�M9S֠	�I�]<rZ��`���A c�M�FMRk"����BX��-(ԮY(���� �e�?�"���	T�+s��uh�M���-;�0���^�8��G���$d� **=�d͖".1�N��n{�)�$;j�WQ�^l3A<�Ob-����[�R��?����,����5�/���u��#Hkò�����c(�B�"�N�_:�VU*�P�*���+�(�qT���ݷN�E�a�L�)g���ԣr���|��p�^[v!�Zz��ݓ��t����m6w��������,�~G���[d��ޭFT�vY�ud&{ ;�8z�{�X�k[��GKc��)-����{D�u�q�,ts���t'�M]
I�$�֞y�1���ftp����p�\�4�������mՂ��')���W��@K�2��i�̚�q�l�7$��V�-h��|7͢���UԸ"��E5�lM�5�e�]��ڿ�����
"�4Pcי��9��p!��-]�*����d�I%w��������c%1�����=6��̓n�����$��h3�Gy���}x*�\QP�`c�k��v��Z������W��\p��V�!���K%`��.�F�Q�}���Q���̄+0CP��B�B��"R��)��N����U���~^�e����6�1Jj�b��,����	�6�)�s&���D���L�A�)�ǀ��^�?����6��T�����\/���%�>ֆ#��j��6\���)���:� ��-(t�k�����F��������[��v.kOh�ƶ$�R� #2�`8���d�����6�p�_���DN���hL���}���w�p ��8�W�BM�W��]9P�Nr3$o&�q�P���B���^,�Y i:l�o�A(�!-q��G�4i���[�M��nu���i�CqC)��R�����|�6�"�AEP\UzRQ*PE𲦰�����)g��5\�a�D�u�U�Ɗ_�gݽ4�T��:%���Z����m>�כ��ds</}��'��4Z�(�	,6iJ wˏn!!�A�'������@�9��D-ԃ�K��[�ύ��Hq6��㞢�P�k����h<ЙҖ�o��U��7�6�-;2�Ksr �΋fx�[��s�w���=�N�b���,	8� h��׎�1��?�b����V�	�6�w/�^n�ݍ���'�ٲ|L��>��FC&��hB4؁���64l̈[�'���֔�m�*��
a���D#�*<�!} �b�ވ���A��0�����nrpa��_�̚j-�lq�򘲑 �i&`0��MC�s���;�<��j4�4�YްF�����Yv���EX	�;|�?��Q��/�x*��4�S��%d\YK��@^�^���0�>�_�=�}�S�P�r������ʣ�����,���t�ht:���a�P���|2Fr�������� npT�^������F��q�"m�rV�.AyR����o�[��7����+���/~,ϙ����(��UJ�/�.��x'
n�E�$�e����Opwx���	e7��w�G��:�a}'�g��gnJ�x��s$�i��Q4^���y����Ѓj@��1���T���;w?h���m*8���FEQA�ILNu�Mi9G�E�w�'�/���)��k��nD����n�\���LH�rK�j�^L��oZeT�vt7��z�scV�����U,z���7p,(c��@�ņ0|^k�����qt���y���to���ل=�d�N������do��lB���PXer���Z�<b�N1m��$�Ñ�(�o��(�ݞ�1Q��c NO�+�q�IN�d/���>H/S�s%�.��e��Q���+Y�D�|�~���k�n:�M7��������\���JDFW��u9]A7��.����а�3Wat��9�Î,J��ȱ���������^��}[T�Wd�xQ�nB�� )�M�Cm�-��n�-T���yo�<�Hm��8ND�.	�*�����cH0l�[��.B�����WR����k�W�H�&\������4BXLO����ᅸ�n�R� be���_�yhE~��_��˻������X�FO�2�h#M����Kox}>�>-�N��:"�?�Xh�W��G����?�Qx]�3��_� �p��0w�x�)�a��`>�{c\�˦ ��$�R5^��{3ǈ�[�:?�&�=��h~E����'�#��g��+)�.Y�����s��[��ߦ��/�#��9\��`vְ����w鳕#r�iUiL��׃���@��L�[N4c�/+Up)֑Dr���n�߻q}���eG�ݕq���{�V%}�x[��:��j#�ɜ��<�Bx��˞Y������p�͏�! j��{��{�����RW�Wr٘���-��v~z��K�z��[ږ?]��[Y[���#�YJ�K1���N�x���[w���L]��*��sҊaݚ��<�l1�fh���^$Q��a����K��E�^}0�����܇�|i.6�^]�,��Y-M��(�*ް�w�eRF�5��~��˶�2�}H..�;~�W�H��؊�<Q��v��4}t#�ZP���!�T��CP.���\qg�L�����c������)����\:���;F��َ�����D�������y��3\���fz�)�`j���Z�BL^*�\����e�̸��+z/�s��a�W{>;A�OGE��_�F�ىzi�$Rd���A�Y�,��2��{G�� K�ZJ�G�aN&%����yu��6��2 (�)�?(�����1R��ʬ�C'���Z�a�}���Cgި��Sp��&�(�c�4k�H����Ѱ�T[�-�����d��
�;N�X!S��$W���ӯ�;��M�DC+��zR����V��5K'��y�:�A~���p�7�"ږ�m<.�^H�ooB9�8ܑ�|F�0�����O��� �c��7fJ�JN�����N�?E��*��x�y�cJ���"E��Lr�rJv����5X��2����r�5��l�;��i��X���O�A���[��k��^m��95S^�/���7)�f�_-�z��F�L�߼����S�C%@s�|Ƞ@e��u�Ӊ��љ�[p?�F�)͕��6��G'���"���N)���'�h����Z�&��8�1n������mɴ�U���}�;smYog��a���P)C����'$���}8��o�(h�a�x~>"j}�y�c�[v7F�@��*�y���5Z�j��\�'��i���ex�1��RU���άD�-�����ť)�<���V�k��%Z&f�3�+.vS�bF�5�
���w29v�������V����y�6v�/��)�V�����{�����I���ZƸA��q��ꎱ����i���s� 2oeX*aM��	�R !�=�y3%�R���pݹ19��=lJ?ev��n~w��D,��T��z�͏��AB��9F�˭o#eG߄gd���LQ\��ݛ
b0C=~s�ى4͙������B��;�Pr����\2��p�K*�&�:;U�rʓ `}O�xT���QJ�?d�8�(�CLsz�������Z�wPO�܊�GSE��fqѭ��te������O���$+�cc�g��>N�,)?|����JҩD��� �Rt?4\�+�T��FL.��hwycC�t�l���9?����ev��ׯ)�E�5�a4����*���}�,c�9�_��8-���j�^�D/~�:��������xF ���Qd�|�%����H��Ʈb��HG�����b�m,���#���x7���'"Ċ�!Wۤ�Z��%��^E�-^B�kfZ.��p���K)�fV��?IUe2�ʕ��^�e&!E���?�hln�����԰��{�ߩ/�g�W���:����D�s�߻�7's�hw�*+����n��_�if����&��@Z<�3&� B�#I�"�֑��I^<%u�V��~�=�
V`�B�֮����,����I�9�Шa�hed�C��l9E��qFOPKBD*|��D_�Y�{5�M��%�,���* Z�ҋ/����D�LL3��	��k�x.>�-8������ߒ��nP��/d�Cio�&ξ�#Rr?����T���Zpiܣ�FeS���e��u��<AZ�΁��G�-��id��_I{��тz�M_0��R0���#)�ƍ"+Vu[{B|j�h�G@�u�!d�/�τ
_M<���x�9����&5K���"�a��]j�T��q�d��,�#F����]�~s��rؐU�J�o�"�݂���ʨ�X���_�-o\���<�yX�v@��$B������D
����e�:'<��j��� -�-��:��h��~J�쫽�'�ڗA=���l�����R�1@�'��'0��~*o�kH����]w�UzT�'sL�t�Źm��)i%�T�xs�����ET�h3��l���fLe��vW�H�����k5��ۓu"��0-/�K��^4hF}E.6*��"�̤}��>�/��
� �;;/���ex��1�A�?���2�7��å?H{�g����d+Ƽ�h�9�0Xc��Z�̚���g&�xmF?>�w���(��}̖?��h��PγL�9�x�D�M��!�����n�@W�|7�	XI!�U�X��2ͬ��f����:�#�6Cp��!�,Y�o3�������zr��t����Y��x ������C��,eK�=�j��g��P�:�cZN�>�T��o;�� i�wdq=].s"Z�ʑ�Q��}�ƻ��/S{�Y�m����#�fL��sЎ�ܲ4i}{�����n�~��.8��V�Y�@�{`;�Ϣ�:� ���a�<W.�)8�x���]�cȶi����2M!�K�6D�� ���6�����&;8>pJOz=|�D��O�XOCDw4�9�ia_��n����]��FH5z�h�s�&��y�@�PxÿV3���Q�sG������s�"��ո���fA"Me�#��ĝ�5�g�XJ+��t���,��/�nH,*�Ϙ@�)y��?�ėI6��)5���UN�4W5n�����2����J߄<�,�zRtO��Z8��
��=�0
)�����q����$���� ��%4U�}a-~J��ty+��2½RX�s�:ė7�]�W�X���"e+�;��%�K���m'���{�"�h�V��T�
�~�V�=��w(�>r�.�'�H��~���\"�ûv�9rjA�|9�<c���-+{��=�c+���jUN��OY(�|�T$���d��ϖ]mҝ/�j��+/�vvZX�͏�@!�<�x85��������7��\�ɞ�=Ü�R�_��6塒�k����IXe��'����1k��}r(Cy��aZ�Bj����@f�xO�����w�翪Y>��P#S�Y�����--'�<����H�I�댯,-�� ]�z��2�n�y?����~�,�F��2��㞭��o׿�:��q��$���*���u�"&�l�I�b�����c��D��t�a[���t�sQ�*@W�� S��Z��E�Q����v��z`_��B�?��@�{�gn=.0ā�	�X����T�k =>�L�"
���/�$�ӌO��Ur9϶�I�+�����~�l�Xܾ��T%Z�����v~�wu��'H��ք!��1�]���ҮIw؇ ��Y��
�Aq��c���Oɤ�[�"H�Љ�����Ĺl��s`��m]:�	���Qi+�Ew�vC���_^�}�����*G��,� M�EO�w���1U�UI3'������m�F��/��lo)������`��c��-Ha�a�\��.^���w$V�b��6f:+�w�O�Z��qC�h����� X]���O����j����	�qK�S^A��z���9ĚZ��@�����u�/[{q��}5��ź�gr�Fc����v�|����nUP��Y%�#ֲBPee,�r��a�,�Ԝ	�s�����-������V�λ��g���c�����j[#"juɭ0�f~$�*�u(��39	�d�Ɵ`�5�d�D��(�z�$%u�dW��f9�x�~G�vK�-���ƈ�(9L�h����5ԏ35��"�=��+��V���؀�u�B��!HD���ߤ4�ٓPkR=���9 ޜ�p�N��M��	A�%ȓ3��g��ADsxOtjo���FW�>�j8��ˡ(�pNh��>�����xYBC���qH�v���@?`d��)t�T>Q-�A4��#4h��q�?L�V�q��qLN&+h�b!"~�5w���2G]�_v\���1z*��q�UHE[��mÊlr�����w@Q�:��
�"+���?t�h^�zvu�e軉�D��HЍ�WKȼq������[P��ؓ��y�Qfi�OJ,��)׆MAM���f�|�݁���D�tj���hx.��(Cf�����F0Î�]7�_�wC8�'�e���J��`J��>|�E
�Yg��j�;-��(�"�C�XZ�6��,�ÐT���@S��d%[f��2<ʶh�����!�5�Bg�jH��b	���w�©��	�Mx;�/�9)�SCK:B`w�m����Ґ�����I����^������M+m�U�ۨ�#�<	{�G���;s}��c`�~έ؟s@���A�λ�ȄmQ�@⡣I)q������BMN�8��*��V� ���C�=8�8h�`�|͞@U��c��8��W�)�j�8�<�2���M��I���<r����p>3�d���BW�	~�)D�������qX�B�,-��Z
+6���W�)N|
���J�������4
��͉������n��CW�,Ѩ�2��D΋U��-��n]`;�����yI��袆d�Br�+WA:5$��t]Y�>΁��9�3�Íj6��a��ɡ"WWR� X)�pЁn?"O5q{�Е=v?�ʍ0NF����9���+�O�4c��}ڈ�:�R�F�~]tX�QX\�5fG��3��{+*P�\Y}��#�N��� G��ٴ���7�"��ox'n�V!61�X�K%��c��(u�_� ��qlQb\M�s�2!2���$'�u�d��%�s9��ߌ�[�q�,��_���F/��������:}�99�*��5�4Ϥ�\|z���'��/�?��Rp���}�{��v����v�$�4Vn����'�K��Ln(�Z�A�m?v���bg�	.V;�����0����O�����-!�c��(��V���_���N}���IHq�����IS ����l���rn�(G�4Rr�����M�9�GVt��7���H�j��03�Q�md*�<.:&��C�DkAO��"y�7��Ŗ��O?�Q�v'�̂�HKt��D�q
j��e/�2�=��(Ȣ�ĿQ*2��oۼ���쁄rXO���"���%�ߵ�nA��Ϋ����O�SE1;/�N���Q�N�x�
�Lx
���ڏ�u�e"8dp5�{d|9(�6;k�\z��d/�R ��)Dsx׻�7L(�bk�:���D�w�ђ�h�{�<��+k�=wdY����4��s��Y��-��6Lt��@$��[�M��T�nIG`c�s��_� �&i�  7r0�;���� 6��r9_�Ƨ�Vܰ��K�e`5�ݻ�e�9�J�+5�y1��$o��	bQ���6�nJ����;���ꃐ]���`7$�Ə��NXV�9������+H<^��P�ܗ/�	cMy�Z2⨀��}�Ar�0��xܳ% �J9�B`���Í�h0�t������E3��"�$x�%��N��Lc��)�Ev)W����uk�OG�E�
b_;�W�2<�gQ*h��N?���MB�Zl�ZV���F��9m�0��ͯzO޼�����q������ ;� 0Ĺ���O9u|-lP�:ղ�UP��$�$��sآj��5�f�E�R�� �ʩ
H���p�5�����
,���_�bN�9�z���-f*+|Ԑ̀���������'6���5��n��t��44D��FI��W6��Ш7���i7���^��<n��?Z	|1�״���pZ�U��Y�L�1(���g |��p�̽N
�8�\��M<5ׇTAPۂDp%�G1/luJܡ��M��i�s�c�������c�SZۅvW�vS� ��������I=�3B����\���D�e��H���pl��� ϙ�X��V~��Ԗ�2���<�9�K^��F���i##��G��}*}�b�!i��t�W��Oj"4CC��מ��W5+��p��Bgx~SNv�IX�/{���~��V*����{-�}XZ�hq%O�k���h`����SK������Ճrm����e*�_�l%VU{��\Ҝ�����=/A@�S�>
'�Yt����=c̒Җ�릫s6m�!"\�*��3�vP|C&���%.�J��ʒs9v�n�?pif��y\��K�C,�
7��i��Ag�*E/ ��k�J��2�^`�};����J�H�Vԫ���T�����Ǚfרvɴ[`O�Mh�7}�N��G�C(�����>Uҗ���cT)�O+m	��)��msN��t�evʢ��:�nR���$z�*�V�
��;�����0�'d��D/���n�+p(���s�01��x�mL=��w���jdrCD��c�k�e+�n�lbP�;�[�@>Eɟ�͖�@չ��-'X�R	�6&5N���63v,m��9��g�dqw�"$T,�>�[��*�ݩ��}�/�N��I&P�Y�_�M�p埔?c�i��O�]�ܺ��n��5����02b�`���9�c*�~@b5Y��(X�� �;)�?�Е�eޠg@i8���<���BI���RUQ=�̉dq�8g?�|U��c���@���Nz��焽��)�oв���WJן��~�ylVZD~�;������}�Pa��B�֯6sT�⡞W�]�O�'�Hˋī/�1y�Gߟ`�Ѱ�dEk�Ơή�\��N�
`&܅Q��O��o4�S�w�Su(�_��M���b��k�ɣ<4�vkp�7T��������~��#����e=Q7c�n��Q�v5ػ:�1��M��=�/����ȩ�t���r��7���oJ�e� ZL�p�ɳ�L�?�b���@�A�&�m�i'ƴG�B��?� Y��p=�.wR��h,�^Ԕ�����e��E���7��-�A?�b?����Wʘe~��h-%HP��Ҷ~vt���/էe���rʷ�X�B��,���b�n��\5��}Z�E������\8r�b�f1Y�PB\�X������Q���B���ٮ�ϖp���ڽ$'���ȓ���ď�dm�	�J���J�(�S5��s�fNOX};���GJ�5��+����	��{Y��-�V�t�6�w�����"}��9o�]e���L\�7R	Pv9V�`�Lw.��]$2 �9D"d�]덗� ����5��<B�X� k�1��%��׹?����LL6'�vqRq�Iu�]�Y2`/Ei<��@U�5T�Fsv(���)�1����*54�5N�7�*O�P�В�!�� 7 �~)�ئ�ٴ���ItF\� \�4ɘǞ���X�V�:1e���&�e���o0B��-R՛�	�h��MZΪO~�����:��T(Ņ��.-�G�a�{�@9�7ą���Fr�}Ee��,�}���<=XN��׽4�-Q\��6�����^�*�	t�\�+GW|��d�9꒩4�+���4گ8�Ιq�D�vC=c{a87�&��Sl�TKL���l�����X-�@�n��	���Q$���NP\n�G�G��?n|�I!��s���@�*��m�𻩶��>�����`��Xr^k�_���.�b��*��Z�����ߪb�f�.��{��4j����u-}��8�1�[C��|�9t�&
WK8#��0BH�� ݂�\��} ��t�V�����S6?|_�:D^|I�s��J��`��K?}����m�d����
"/H��:-�$*<�߱�Z8�A7�Kj�f	�Z�eLM��!C�Y��@�}b�;:��䊘O;7}��T/(FB��u�w�b��~���Lv��p��5Քs\����oX�˶�ͮݶ������M"
�R��M0�b��E;V�	�U�~��O����_�,x*S�%���Ug]���H[2�&9����%TQiC\��{P�����=T���C���e�(]�:�Jt��VH�˭~��(>M;P�Q`�q̀��p��R0byOC������{,�i����m/�5l|FýiV���(��6�ie}DYj��F'��X�ӗ��6�ed����ؾ�=�~��l�7=�>�u�F�J�Ŕ-B�Vl黁�������F���u���'�`�V��km4F�E��wA9\;��t�8��d�.]���Ѝ#4͎&$N�1�XM�7*{Y==��˫�����3̋�"ޞ0E�z��#C�����C2�H� Q���ݞ*���b����r���^�8��H�Z�0 ���*��[����&�%c�G�@Bf��dt�����Z���ݡbx�֬�/E�������k�TS��-��5  ۶�ʝ���D�Z4gYN�:�T�3�Az��}��<8O����p��qZ�?��5��� ��^��T�+j�4y~V����~DK0�!�7�u�T��-�d���_����-ޥ��>.�K`y��*J��=��-(���מ@L>!SیuN�d� �U".h8JGr����z�s������i�L���Rwa�2��7��0����I�����KUI�s����K!P�)/q�&eՆ�w@?J �:8M�-��4��	�(�+*6��9b~�p]��EN�c
š�4+y:^:��T�dR�A��2�w%�YEK1[5���
�1)���i�Z��d��j���zuU�=;ߍ!���v�r(��7$:c����u !����:m፤�}:�1��! �+�qJK��շA �L�`�t�����M,m*��酚O5��:)�,}q��f�Ӿ�ܼ�2�S�=�4�E̠�[W?��v�7����8`ˆ��r+'�FR��U 2Xxf�jh}�7���M�׮��t$��d�9����>,]tuqd�w͸�|��sD�RLtER��Ł�3U���O���/s���q3C#��pw�K�ZD�1�i0��[�a=W����y�?�	>&[�$O;�A�|���·1V�W�1��ه��-g	���*�����K�>�oE[�9m��z�Z.ZP���������]V�.<�:z�8�6�\�u+�Z���ͥ�2鶒(زi3�@ R��B30��gi�:�"k%��������T=��-ATo�>u9��Y"s���n�̏�>���$Am�L�?؄g���E1�e8��MTF.���٨�_bĹ�A>�Y^�x�S�	荒g��gj_94'�k?�w�ɺ��&��>����bݬ"�4�U��pmϑ��pw�`�F����$)HGaw�3�oڰ�,�p&,ƃ'9���p=*j��K{�o.��	��$�q�M���yqӚa���$��h��M'��WM��i"L�U��a�v�h}-ޫ���t(�fX`�c���O?���`����9�䛺796&����ŗ�C�sp�5��RN}�U�i}���v�sQ�;�(7ge4��jOKf!ɜl
�B��Qo�2f�f[>�ENke�z1�F��,��t5p�J3W}��j�U@�k�+�ls�����8�-��-��,��X��PE'sa]�`����jW�-���/�W�2�l����vTQaT�.ݸ�(������V��/�v�vh��S�O �*�K:������@d����Wz �E��2[��0�jY��d}�"/>.�Q?��Nq0W�=S{Z�'�����*�H>T���(�&l2t˺��sr�� !��UR�B5�4s��	���5)����7h�k^t.ky�5x�*���p���z�*
��ERȄ���ZE3��">�x�]�mi+�l�2���<���\갨��4Xئ>���!A�;�0R����v���^1L�?��p��w>«�8�#�ɶ���bYΏ�v��h�g#�l�\9��k��9��b�K¹s�K(��+�;���B����ėb��f��@���&�\鍋p�u^y�.��ID��vG #�G/"?e�*�0���?5MY��z��{쳊'4���(4��j�ǳ�X�
�F���J]�0�̄���h��%+Vq���
ds���qE�!�7(Z�$��v���oB��G*�3S4���l�T�,���>�^!6��ᷣ�:J��Wcf��4�3Ϝ�E�.4]a�`����p$��e���q�v'.���L@�,8��任�H�qPc�����Sc���|�/�
��Pz���ɧv��������<�VP1W�7�1���7��\f�!v8��0|���j�+�����P�5k�sN�m �u��}�U�Ou�D��[̴d�Hp	ja���\s�K&��$�xy��XIj�����]3��d9e�i�g���1���pd����י��d!�������~b�m|�UG�v���Tx�v`������U�8h��ZκJ֭���J)�']?�^�%�
��yĵ(�:��S,�L)��?������M{�Lo8������W�$�aʊ�m���^��I4� <�@�l�1�GA��Q���;�x���uQ�dT�*av���K+k�ܥ^ҧ��[�/#�̊�0��t��էBì^�$ߔ1�y���|`ЄL'�~-_z��&���m�uS�xZ�\�=��BݔC �uv��>wxfpo��w:����u��N=d���0-(U�1���%����^RoY'�5꣸�%��1�$��Ы/��/�؝��Sejg�?1��jz),)\��LS�+d�j}'��Y��|��� �*�D��?ޮrӳ/�}��a:;@���lr�lamWqs��@U����<���=�ve͈�Jy4��c���:�Cd�f��{.n�O�;ZN�[ςHfv@%o6%�&�\
Ha�i:a~FX�a��~�GZ,8S/���)5��c� �'S2`o�dgNs��C܎�@6��*D�X>n�C�s<�܈�]�i~E=qa�[�@���Ѧ6�#Rg�"�#��Ћ�A���W6�#�/�6fo�zwuR ������#Է�39%}EJ��*.p�#�K��K���s��܍ss��1շ�0�n� �&�8)��z�=W��)Q3�8����o;�=r@f��Dld`b�s����k�go��R
е'Ju ���1g]Q���,�*{�l䗂47*��=ʬN��0��L�jȠVi�}��W��㛓��z����LќC�(�3��W�>`���s��<r��۞*2̝�eR�F���o��A�H�$?�>V0�(�E��"h$*ơ�}j�`�� �A\��+�C�ݱi�g���r���C$cU��hc�O�K�e��˃����O�ֱ�t�zs�����ޡp3i�c`8��M���'��c�:Ju�)��O�@�w��`p ��_'�}�E*"76������x�)dV�ӯJ�}yz|�
"�s���&���^��x[����`<?�B�vQ���̕z�� P�1�ں�`�t���sδ���Z�L�+*�B�㊏�SN/��E�!gkc�f2 .��5��}���5�*�Y��2Rx��T��(���1*��:)�����l�𽲙�z��:/17Z�̘�u��r�S4�� ��z�"Û4������u�if�_8����T�a�,U�۵�5�4�'������N���W�����*ur51C�sW�#�B��KSf��L���r:N�0�xSQ�y��}�����(%���5[Hsau# u���`�[7s�$�s��	�M��{�j�F)���:�����++��v[��������U뢙�0��g�Z�l�Ѧِ+�G�߀�D��������M���,Ȕ/�Ɩ�����d�w1H`�ʉM�cO��n�N�k��q�~�˫ ���@�����]�����x: ��_|�m"s�sk�R���x>�
x�D{\3���H�� gx0��O�Z���S�f��f6_�B�'^���£۟ęGx�&6�?����T���[�ࠧP���N�����J��۸B8���?�S�zʱ��z���).1ڬ�)��-=
����[��d	��;r�`S9��������^�nh�oi�Y�R{F6tD퍈�=��r�� 
j\K�#y���0ީ��5�19&���3(���s<�͵�ɆsXy��rt��
�Z!̯&�W�x�
�6�?��8��vj�3̋.�~������� &�+��®Ԏ� X��l����C�<�S�,�.Mpޯ`���`g|mz�w�)�d/+ Qu��|��L��sG�� ���>{�a\�=�$,�Q�(�o{�g�-Zhu��o̤A�X"TM�;����`i�I�y<f�}-�f�@C
�9�J�8�������l�=�#E�7
�j�Ƃ�C��L֧Y [J�`�h�20���1�[t��	�H�;qw�Q�ݰ�.$SK��W��y:�/�C���;����������P��r�>��)��	#�eWg
���V�ꐠk(9�f�?}����������,����d�0�}�P<�q˟���(&ͳ�]�U0\��#�B�~�7;��Ke\+��OZQ�F�(� �)ɭ�~�]?��Qȃ�����9J����p�#��VQ��г]t���e^I
�
�#�O�Dp>&�� E�����	:}�sk���S��RE5�p�&Ȣyi�A�R�VB��1o��`)5���i���R0Y�
�k\��VU>l9�Ɲ�*���������)f��:�csZ���Pz��$7�
�o��"K� ���*��$����?�:�|4�1��X9�aƾ}�E
�#^�P��Lo�U���;n?�')�QV>�t����U�Ӊ!���"��]�y/D��r�M�%dL�����'��贏�Ǭa�#�3c$�	�U1(�S���VJ�T��v����S#�t�d�������w��ե�o;,L�Y��t����q�d��������GM�2Nw�;<r�d��$�{��0��Ӧ5wT���(&��~҆��ƉtF�ۢ�<S�2�f�ʃ��y���U���9S
߰e��5���Ă�D��-&L�խ[��j����]ְ��P�T y�
���I��sb��n��T�&fVrW�V�_����w�� ���٘���ȥOp۞�b2~=;��5�c���t�Kܗ�D`��9*���׀��i���l�?��q)L��8����T����c�j�v,��a�a|�2:�k"�+�Ip���0�L��*C��@!� +a*(�ÖX9N���c��P\l�
�'C'?a�m�zd�m۷�ë?%8w��(t$�zTѰ������ݣ���%��{z����4�J&^��q9pC����m�^�Z4x-�H2�-PG���/�<�,�r�L@=�	X
i_�a��ҭ��p:?���V} E/�'ݧ�1��m=���2Yld ���!z\&R�������_UTOIL�]��1��t&Y��m0�xY�[�<GӼ��g�yދ���p1�r54U|��m���^�\+�ۮ)�������h�KF�#����q 	��v�����eQ�??c��@�D�\�C�c�F�q�od�\��j��U�q���8B%��H� �g��Y�QǎRVS_D�>`վ�-/�һ~���Ct�ϕ\%̙�!eXb��@��HBy����
��2@�0\�v������'dPRq�.냣3����t�q3��x����O5e���7E4�X�|�-T	�g�O�ӆ�yU{��b!Ŋ��=r�p������������,���4��W����YЈ�%rח������^���(W/�q��'�����o��i	mKmlҍ�nJ�:�&p�0zU�+aB4#]��9�)+R�dȧ�fvg>"�˵�<H-�U-��hB�3��[��L��xs��[yF!���">��m�Q,:�;�U��]8ӎ1(����տ>F�t�ࡪt�2�O��^�D�H�S����)H�] wWL�jK?3Bu�R1�T���rw�ݥ��4_9͟l��\�����W�1I�"�&��kA+�1sf�t��n\�s&I�ה�7���7�A}ƻ���0� B:d�:4�Q�;���Sb_����{B��&�̫�x����M�����#
eI�r���t6UC�ն��p!G���*�*��и5ɑ]#J��C���<��F(�PVh�5K�Ē��%��@�MMH%���D��Iq<4����ooK�O2S�	�_��mEXJ�RB<ex�P��*|kg�FW���Qi:�����E��C�5F/x�>�	����P'��v�T��c.ř��p��}%i���(�e�ϟ��u	i��S �ڒd�i�a�2YqO�z�� XX�F`P�X��'�3�a���4�W��SSe�8��ki�"�f��Ĉt$v��#p;p=?u�9z�����:��%R1�����)ÉVǆ��,Xe�3� G����{F��Π���kdch���#��D6j`���b��>�붤�hB�Z`�.3���4�?�SĈ/�AP[$"����q:P'�I��։x,�v�yw:2qX��Iw|F����z��o���z\��92��%�Lh��>�Du���B�[4lջ�.]݋�c7Q,�gC7U/gnF�ׅz��l��n����P}I-��`�s������YM�F �(G��ȷ�4��]���6C�A(�4耘�]g���w2&X��gu6h�L�GYi�6�m�@���уq��PM�U/
 �e�t��K7f͵هؿ�oH�O�.������@��;+Z�K���.Mp\��jjͭ)��.M�=�`�ۋu#2ȗ�m��4̸�D�_�i�^�,	��nªt�w���,lR���i�86ll��L�N��5�g�yB!Ց��D��&�@�aE�0T�������u�*���[���r��!�"�9�=�E�<�>&�d���C:$��q�L� R1�k��Øn��ZA�E�=!���4ܦѡ�쑰�T�g�@(Oc�K��" ���I�z}�%����!��X��0���"������D'# ��jg�� �U�$Y'�Q9�y�6/ب����,�;���H��&�k����N��M���ٜ�� i3�a�~G�.*~��p^�������	f����[[�{]����C��9����c�T��3bM&s>�/��
�u1[�s@�K�U����T�#����DWhڣ�鵌�wA�ු��-�V#��A"����T��W�ѯ�w�U��b��db����Ǟd'�@`�֮}�'g���Lv� �,�����P1�tu�Xy�u��]�a�pLY(��lsH�(H4f�}��X
�}BD���f����=�u��Df&�{1(o��e����,J�� y|݊���L��m�r�G���W����H7pt��>� l����H�tʆ�c�,R倅��M(@S����|���.��A5���4�>�p�D,�p������9��-0��@lƩ���tt�b�w�Qq�����B+y+S����ԋ	��;�8ٻ��Zbcn�w�Ĳ��qn�Q�Ɵd3ҁf~�΀('�1
�F4�Hv�\4���Yn�0G��q)YC��굽�BI)��Z��G{mҾ�U+��ʎ��:�3�g&��+q��0{�u
�����[�+���w��/08D)!,3?{6u�u��z�KFln���`��G#f���T��q��ޜ|��~�(KT�Q�Fi;1��WZ�QG'�ĶA=�i���=��u�3"�,�8��k�o��Ӻ|"W�%U�C��C�/���ܙ�0���ې�g�\��䨍^�sY�O!��#�N��5H���'r���Z�9�E}	r�ҷe�]Qe��#UM��nf^d���m�>��ή�X1d�kBp79���I�6xge�rw��S�����R��(%|�$7�������^�(H3|��9�a��E��-��ļ�i0��aZ�7�>�y� V�|ojJ��HOB�ʝܸ�ǐgգ��\m��Vg�&5d��5?^̀P(�2#��V,����*	mY)�85�-�82R<l�z��Еm6�� r�q	~����?C���!'�V�X sԃ�F��
C.��{IQǗ^��+wA��N'�Bh�:&��v��-�^^2�s��z��7�E��x����8�+
D0W0
��a��I`��Af����Ss����#�O�Uj����d/T�F_�\�Ō���k~�Mv����=�`�0��R�)�o�z�z�II�j��b�B��=�+���,e��n�[j�o�-o���(��h�G%iP��zg@��w:,�u6�j�0+��6��$�Dp��*�x�k�~)�!���Mj'1ݫ�����۬_���?`��{ =���j@��m��u���*O�x ����c�Z}N�!�8��Q��e՛ÓB�6�������a���r.�%#����?�%�7�MA�'�=��BA	]�-	��;C�]�xN�4�Hio=�c��m�}���Y.��r暋6~��w4�!m��2;�n&�!t��y���a
�!5�$��|@��v�֪���G��G��C���q	<��l��7��µpk��^��$�J	:s.tю(e��q��K����zj,$;8�����v���ȍ,�iС[��^���v����|�5d�3U���i]eP=G���U��4��/E?���cM1׻�o�ݑ'i��u{��M���by�v�M�ȶ*�$<3�4�5���r`P'�]��|����ߡ��/��޾o&G3}5�z34.K7��ΪjƀwU����2{���؆�mv7�0{(!�(ai>@��� 0�)��S,�Y�a,�:��~>e�#+T��W��˨�3����`e�'��JXC�d!}�PW:Րį���5坛A3h�ĨunH� �pF������3ݯ��5�M';f���Ʊ��F�W��G��k$��6i�_�ؑ3:ah�ɱ?.X���]X!j����"�yʺy3��ޣ����3U�&�ӭK�n.�e�EE�dnA�I�N?4I�'��p�,�x,�
��`g�/Ko`a8���g�nh7�CG[��C�4���p�� x�fnǝ���@}���g��r���H�z��nn],�R(ػw�LO�a�U�X���D����H�r���^���#q� ��ġ����1�h���*���(�Y�8��"�k�K��M|��>>_�z�t����ىJ8�	3��:TQ������Xz1�=\�o|xxZ�\���Y7���|�.��)�U�#��p�烒@㟼Z`k�c��xf���O��Iz�"
��<!Аw�'D���-!� �&��B�r|OYƿ�����v�#�fə��
�Z5]SY'�.�C�k^ऽH���k5fg.(l0�1d�h�][A��Uu���l�jiI	2?�*���t�})apwwBTf�/��\�gYiۘ]Qն+G�D�({�Qe�f�7��%�LP+�:�?K�O�nn���q����2/�s�𛼑݇=�P�h/O���-{_j�����i�x�x��)uy`v3���Z=��b_\���/H�?
��.>g������<n�d�,y�	9 �F�o|��=6~��nSAT�-a��;�Y�bY����/��(`��Sb��` 0��0��gTnJU�8 ع=ɓFqT�/�3��M��$2��	�*A���t2u�6h=%�~w���b�:[���Jv/����~�\�<=8x����f��x��/z8Q���&:��Ҏ�
#�%0a�-��n�VP�J�51C��2���\*@���
�jz�Ll�(l����1*�t��Y-��M}qn�?]u_M�MI*���$҉����Q�֋;�E�G�3�<�\2��>=�s5�`��C���!�R#^�	��"MX�qם�?��y�nfv�����r�L�[�o�4]�/��}�9C�l�oDͥ�zd*xť&v��g�ɑ؃�m��?s7;֢0Uᔊ�x&6Y�P�K�m+�z3����5��t(%3������S�_��|^����=Vou��\�����C��L�:��Cz�yz���G�34+Y���(5H�j �x�����ȋ��T24��Ä�������t4}��1�r<�U�Fp}����:\ÿ���W�U�ƴ$I}��Ate�T��@��� S�t�W�����$`VT�ovؕ�#��_�dp�a��H�����X�)���^�-v+�N��bKP1Ÿ'��m�o�k+�� ����$���U��V��~b:"�E��ݩ�jk�4����5� �q^����r���B��He���)`+�~�ߜ�]7ϋ�w��2t�Y�tk�r5on;�`�8�1����w�[��@n���́^o�$��5��b�u�%k�1�r?^��T�v1�3+ +�8��t9/�J|�&Ϧ�;)�@��۞b̈́벀������G�H���C®�զ88�6LtH&�m�G�ڏ*��=K5��U���@�Bs\�S)D�h��g*Q��N2"d�r�}ϙ�E��}~*�I��QdMC÷٬��3(ꍑj��v�e\�6
)�谱��&�~I:�)���L�Z��/�7��H��z�#h	����?�v����L�V5�����d�(Dү�Aы�T����M�����NW;����鹕��58��6�bD�=����~k���NpH<$���"�,!T�~��+��b��F���I��7�Kl�55@`|��;n��+�j�@��{�e���'fD�}r�{��<m�}[���Y�bӂ�4
�{m�̬9�w��e�$����G"r5��SZ{�2�D�o�&��R�
��%�{3��Z�edF��|����~�rCN��/��ƣj���?��o��	���b�k:j���?��c9pY8@�@iXh�����j�T#gg7I���li��Q�J9�DlҀ�=WiQ���U�m�����e�SZM�mSW:�M����SX�&� )�~w&K&��+F��%T����O��2^��\�^6�0#z�#3ǖ�����:w��d���a�RBI��1.��$�ҽ~�5t5��'+�+.�Mmt�qC	���Gӡ,�� �F|�lw)�j�_�fA��Ɇ�妆���C@]
��l�
�C���	����j�Iy���B�;8�/���o�'��b����O�n�ܑ6�S�X�1I�E)zq:����gD�fش2}Mډ���Ș;�wb2�q0, ��M��%\����'@�}����5�dZ܏"��	�,�X�9᣸jF`q�����-zV�z5�(�u�U��dt���~7&�*R��U)��RpEjgȧqf�sf� ��]#�ƽ1�Lhlp������#�O|ۢ�X����:��T�j���y��(<����|�G�p��@�%��+/Q���xJ,�Є��0����[�8�5Ј�@MJ۫b-�._��IFys�w���sO-���tֽ�a��gq�h���dr'���d��pnJ�q���Njq(�S�.�g��n������ �A^�=�1��B�$�������Ay�zgb��n���=�a�����!G�P����bJ4(���p�5��(�Ӹr<�ux�(��&��Á��L�9��e@(�i��N��\�������X��xSоə��� &���#�=%q�^B���2 �tL-jY,USTd�e��zQO�/7_���I��0�=����Z��(x��/u���u�N�v{��+�a�̓��k 2��`�٫�8�Y ]� �o9�m�l)�q{����$@|���3��K=�k7N R��&ƫ�?9�h�Q�[1Ճ��3��4��1x˅l:͵�9G���N��G�H��������܀�Y��
�����~܄0�`�£T�K�|2gg)L�9�t�_��)W����M��q����8���.��������f���:k��C��扝��=_OTk�l.Z_ƙ���]��3$@Ս��R�m�2l�?�,�0�%ͺ�j>�MM���{ґPnB�O�p��y�Z\A�qRj�ѻC���NE�-�Il�@�cq��G�ީ�S~5Y7I�SB����Pp䧐��7�	��g�&�l���k#~�K���j�=��֧�a{xF�1�$h~2�\(��:�:���!�h؏�B�\��K��D��mA�U���ɴ��f��G;]V����En�_L1���y�N�Z�������&:,g-�ƫj|�?Z��~.�D�d�$�T�t�/��5,%!��l�*Z�V�2�L�?U���@	�PM�:��m�A�Õ���Ƨ���x���h�U����m��"��]��׌�IWU ��= 4�' jF���e�V��f���a�)w�G�:�l��.`�-Ls�x��򓮡w;�w�^T��գ�"R����%,w����&��YF(�8�r"��s�J<ǲ�+�v���O��Qa^��QqV2VõJ���8? �����c��3��BB��;�VZ��Q��~��r���^�>���ſ��aK's�}�1@��;�4z!b�_��o_�/���f�N����)��@��z��I(f3k:�c,���W��+)���ٔU�J��V?i��K$m\omA?3-�zc�T���vSU��?�c���D��`�b��.2Pnܣ;�"����d��Y/B�U�Fbʣ���L�|����j#oh�zu鑞_W$��%O��,�{8����r���u�˘��UA�Sp0�m`�α�_�,�Ł9���h�=7PDr��jWv�S6�2(�|2�M/���#P)k	k/�,\�ZU' )~�˹j�,Z���{����������,7����L�\-�MF���[��*\�P��h&JZ��'�N"�UC��3�]��ϗj��]#f�n}
���T�D�猣�NF���l�3\�Q����6p6�A����좩<���P>�%��?��x�L�	F�H�uR�<L�Fi�%y5���m�U�sY
�Ӹ4��8|��C�A��/"d{o�б,*M]��-�0j�$��N#}�'S`�6���F�$�N8�t= �q����c��� �Mk떋<7y�v7�Wͮ����4���k��m@Qn|	w�TIan�1)�)�o�l��{+��er��f�F�gocGU����	��Qѯ�f|�
3������/�u�g*<�B�`r_D$'G���W85L��L����@�$z$�ŝ�#�*��Y~�r��L٭���5�}��K�����mx���H�P:����Y�G����0��v�3���΅6c�4<�&��7y�(C�/�=`)i&)�()�w5(��~av�,ϒS����c%=׽��p�e����wᔈ���E�I���-*��G�
K�>��ݟ��uV��ָ;_'�d)�#����j�kwI�x�9<!u���J��9��*��J}�{_���>�v,-���l��?�W���|\�X2�\���B��/�v���ks���B����io������a��ޕ٣S�u��	9	�s�_�pk�)�&�!��>Ȋe�>��*��S����!\�q�d���0�so�0&���oy��J��e��r��Ԣ'RU7o�ͻ���S�j��%�T#˒�(�/�U���w�c��E5�� �v	NO��mZ������nΏd�O��^��C���]өP�%��it��5�j=d*	��ey�]�W��D��Hm��6��c��"ni����R�\����YPdhK�v��e��|�BP
O���dt�򧱃,H�M˶�Bǅ�9��B�DY1��P$���a,�F���s�Hǫ�����V/GW[���	7��K-�?�a�1�`�����v��,^���{$�|@����Q��8se6`��
vި-��/�SՏ莣� 2�E�f	��X�v�LX���*,-�`a�E�
�����ıg�/+�,�[M���	����
e�����>�D��@
�Z���fN.�Ԟ�^ׄ�Y�q��ׅw�S@O�p�}�&�C�Ŕ<(A�c��1��a�9���]*�.�`��X&GD�)�/%^ޫ�c�a효TS9��6ŉY�'��x.��$��O.9�Z/�����b�#����M���3�spp�x������0����=Q>�ᙖ �����&[h���Ew%������68+�Ç��\aоK����GB�o�n��D�
շV��K+�]��ť�1����@��)��4<�D �	��4�a^2>鑅��@��4�D�L��ד�76,�魫*�U-�<]ڋ�=<����7���$�{wD-;\G�ယ;��߅3�7
���0i	���$��bb� �b#�ay
�K��(��s��Nobc�a+�I���%�����B�cl[)H��-%�lM�a�G{Y���r�p�����N3N�s ��-l���m��:T�%>[��ȃ	䨢�؛J+v�p-Y%�dv�g����OK���A7H�� 4S� SY�Ǘ��J��o�q���ǭ�c����!����g6�J�ɜ�H������Y�wg�����e��j��r�K=p[����Ʈ�Mɷ�m������īZ8M�'�,$pe-L�޶��>R#'9���K���W֘R?Tϗ��ϴ��G�M��e����)y����Y��M��tݵQ��_�,�<��6��c{��BvіgB�QG�fY:����"JX������:GR;��謽�d����,��MN���GA(sC���-.4��n���f�Evz1�r*R*��4*����ӥ]mP�EP��=$w��,ԇ79(����򩧕S���\ha[��� k{�����';������/bt]�]3wz������u^�Q�c��Q�� 4KS)NM�&9	�.�9�I��k�ϪC�"��W�s����_l��*7���ݚ�Q�aW/���^^��cY\�T��ݬ�Mt�8�'	Ї��I��q���q��zh0�}v�����9<��JM����3)��p�X��Q�!W+���>"�(��İ������Gj|����Q�5vqY!�D���=�}����!����輡��1t^�&U���q/��NQ��{�$��lC�6<[@ǈB�]a)l�H����F~3h���|����c�6�����d��#]9w��m"�dpS���A|Zp�כ��\z�w;t��>��I��2���a�ot�Aȫ
���P�ٰ~;F��BP�� �������K��~Qlfh�>�BU�I��M�������(����ɥ;�Q���I��P̃���hi�� `+�C�,����|*�A�;�i�fJ��o��4�����ao{��*?'���c�Ng�A�T�a��
����I��.�j�D_y�k���@���0̫}3j�o����wbj}�H�Wm�Wۋ���$%R���=��<�C�C^�C�]+/�V�[��:tU8�N�������4�6���2�,��ܸ�I����J,CN�t���6F�a�|O���*NH��������c	� {|�};H/j��Bc�N�e9���Y/�/k�k���N��(����d: m�-�ш?E�	�9���Qq�̄��j,Aם#����KnTUZa���+� ش.4[5o��y�J�,���]���K7�hF��qg�Q��`��2�n��w���� �#���#��`�b��o\<�y����!�RZ��a�[�J��U����v�e���.����N�&Qa��� I(�9t��(���3�Ճ�"��x�� �1����"fP��0.?����Ȏ)W7XV�����Z�]���|Ҳ���s��oE�p �1���90Ӯx�
(e���ޡ�|�1��@p�TR6��I�8I��IQ����ix���[�"���`795�	���r}���F�?��c���
��d��]�U�џV��Q�|?�U�Xϖ:j��gΆDq�ƣc�]nlD�{��0�s����P�t����������a|�c���$NC@?Ŝ�5�>���)��,�5Jz�{JG˵��C��ژ��~&�ݜ�<������xE�� R�qPRO��ћ]���L���(j����AJ����9R|�'��+�|�P�^�$�b��^���s��"�3��o����V�ݏ�[B���#N�Գ9���<��`�*���c�m�D��N��U�|�frG�����] ���D���!*�){��������e[�n-�y|��,�U�Y��&�[�+T3�z/e�(�t�u�d�g&��cE���f���Fq](�7X���@��V@Ȭªd���>�5��DC���\-KEM��sP-Ͷ�}�E��
D�Twa#p���\�)�d$��Z��úص�M놽BM�?t`���Rh��ŋ�y��|}�~n��M����M��|���O}М-��/kk��8��5L����G`�}�4�[H��Y�w���q�c���\��7�~v}Y��г�}�OXQ+���@i��� �R8fG���p���Spe5���⍨x#ֲyɤ|�Cѧ�u������f����<5������1��Bֈ'�ldaI�G-�'���i4�*(.v�:wڕ��։K\au��+u&m���\z��xN��2`�r�y@� �.2
�ģˑ(�E:2�2m\z��(��%�.�a_��|�h�6��b:��3Tl�g�+��DbP�F=ͻ
��Rl���hM�=!xnB-�f�P�����`R��B�[DD���'��o�/,m�ڙFM2����8j��f.'_i�fl��j��}N�?�) �4�-����I�*P�g<�;[vH���}��!�/��gt�nU�3�	�_k�^���������U����G�H�ePܕJ�}O���b�<�=���7����5W�
JcQ����0�Z�W�k�<J��犺�^)���dC���v�1�������V�Y�����t��MOl�v������vAV�?��П�/$l�"h>��=�B:���x�Z�5��Lc����C��i=��l�/�ă��6a��Y�/$���}����Ve�� �/�)uGv;@��I���[���-���T�˵�^��eWʀ�_��-��AE�X"ө���}�TFپL�d���s�k �E���H���k/z�L�~�Q2pi�$JB��7Xȉ���pܝ��� �r��r��"�sNEf��]��'Z,�����&W$ps�����:���d-�T.�P
�%Կ�ݬIx���{��f;����#]�]��i[���)t�f�C?�.*��e���]5�Sqr,st���o�WsV�e#�L
]�oCZs��ȷ����ɒ�:RA*XE�=30K�Aόzh��1��>:WFΆ3��2���|E*��l��AS��c���G�!��">� �4���8����Y��1��,��)j��'j:�mt�P~'F�= ������`��ɭR�"'b����79�vo�k�v��1B����B����f�	�O�n�� �ʳ�鎽���h��;��r�\�87�t��i��Y��Xe:�2(~4ߖ��{��T��.��l�m�����0�Э�-�/�7�,�2�V�2�;�=��b�=6.�&Ye3��W:�0R/�%�~�_ͳ>�#��;�q���6-�r4-�`卋B�j�w	) QIݦ�+�1z�=.�dms�"
���gm]A�ZY��d��w���&]�ʢ��ǉq�@����o�o����i�/�iW�=R��m���(=��e�����$F.����p��>��|`$��Y�;��U{���i(&x��ºj��9H���M�	v��;f���N��D���U�E2</��p��wq�p{��0�n�Y%a�<�JΐS�Gc8�q�o"�i3S�#϶Y^/*�Y}��|l`f~�*�hj�2y�#��i�_�l�E*��^c���
�TF�*,0=�aN�o#!ak���cp	[�u���|�D|�Uٗ��������f�w�Vl�ɰ�$�I���pt�gv��P��/��*��g�L~�8<J��П�d_�+����7n��ٸ�%���u9*�sw���{P��%˺�6�`@�pT¨{,��;Wߠ� "@D$;["���K�C�b�I��E�j/{瑓����ID̠�3�b�g.�
�`�:
�>je�Jʿ���z����ᆪ���H듢IiO�2�Y�E=v-t��D7�*���Mr���Q�ZV��=X��go���@��I�>����HDr�!htu�������[��G@��9�T	"�`��ã_���#�own�O�y#��1�{H�Ҽ�=A�r�ɯ�x��K��i�g2FY�� 1�K����p�������-t����/S�8��3���!�e窙dyz"���T�?�u@��d��`6��ߒ����;��V�;}"���u��ҥ�CGy������ʂX�Fa�e}�8��R����%V�c/�����X�7/�lG�<�9F��<>�O�K-����'�z��J�Ԋ����쐉ˇ�c��OiLV�3;2V�q�t��_ے>�������p!9��y^�aT�	A�a*Rf���-�����teG,+��*礇��	`(�v��z1��- X�1T���9����þ�@��W�.�SܤK�����n�8	U�����\8�G*QL���&9;�t��s�C{�� fE�Ƥ�[- �s�Hy������~���:��>hw���(�rr;*���"�4N5enR_q(�V��HA`n� ���BV��R�M:����y}3�Z����a����ӛ:3T��2�G��e��I_d�q<d\3�/� �}g�g�/�PR�h젌%�Ǘ�nQ$��~ޥ���%��D:�2��p���$~����x�'��ro&R�2N)J�5��z*���"q72�}*����	]m�fY���5�A���x��5�>]�2c��؃��;R�BՄ�j�(�|3n? �2L��-��c�n��cI1~�`r�_���(8�ujL�� �'�-���Ɵ�=w?��]�4�����T���W�mp�~9M����ωKP�*�p��R�E�\�O�=�=b�ߩ�I���O���~��h�+��n�H�|X��ڟ� �U0t쪬��������3�IHkȪ�E�q��e�kҀFA��\����J&��A�š�G�>��5_ts�ֱ�,��sIί (p���ss6���4k]�i>����n>�Ⱦ�	:c؍)&�4�f��G���rG�ʬ�&�#����k��ر���Έ���0Z�;��>����:���5~�����}�3T��5(�;E�Sk�WG_JL�2�s�ؔ����e����5��;/��ZWOm[%,?��G���3\ �lE�vTC�A��h���� ���iI�!�<�Y/�%�;:�k����0�ƃ,(�t��)�^yA>Ǉ���e���ֿ�I�0�U:3��C�@�ҹS�'wF
�`�o*��X|���J%}I\�ڱ��sf]����fL��\�&-�1N�cm��[wH>WX|a֗:�1G��a�we���%$@�t7s������[�^ ��	�YF��=�Nt@	Uw]�|]��۝Wn^��h��E��0B+P'�n�w�j`�m���Y�*Լ;�Tɯt��C&e�^9���/�jc}�����N�g��D�1��H����	�q�-`_��D\����^��6�������Tϗ�Z�E�Uk��"��J����L/ �.�s@Y-ꫦ9Ru#�xM��%�Vk�o��J2cW���V68�T7�Ivn���g�-;�P�.�+���sh�I|z53 �J���__��g�R�U�cPӯ�N�c[���?��cxiQy�p��h��-1��9P)�z�o��#h'x�P�.�QUs�S螑�a���E�&n�{������Rk�ڏM2��+�����HK�z>��P&�a��q�^(�Dɉ�j���}ho#��f+f@��Q�T�N�b�w�6��؆�T�Fy�_�uڔ��L�Lk��3��
�$�z�}�I0�Us��	lW,�wM�|�)$����F�b��^�X�ē�åS݈�76�H�~�(^Z���[&5!:.�V�Y�;��֞4��T��jq�S��	�0Ҥ#d_�/䞊���4����p�_���t5z2/`��Y�W��CW��^��N$�\VϦR�,Bj �t��DW�e��xpQ�Slmu���	|E��Aj���H��j^)n=�MUbS{�����<�[)�,@��GG�J9K�w㽏Yu��/�Mng���.d��=O�y
\��h�#��������:!���=O�y|`�t[ ��8�[���ڐtT~}c�� �Ѕ���:�e��%QL���Yv���A˶�=	���3^��h��F����
�;��8�W�Uv2��@�Q/j�VW����״�ۛs�`����=��ߜ��&���0#�#�>�.�&���O� m���M�rKo�WZ����J�πm:��BW�:޳�꧍&�n"�>1�����N��Csrp�NYY��1S$o9�}v�>�(Kތ�bQ�$_�d�ͷ/�ߤW?��E�4KϠr�����R�/ִ��2��cIE�M����7���{&j���(5����<�3���P��y{P��n~Mt���}�ϱ/�"�i�Y�J��o�ym�"h�>2��<:F6�>m]���!�m݊`��n=:yH2}��JZ���<y���L���%��?Lx�v����T��Yo7Ҩ􃨄��8��A��@�O	nS��2���)�u�i�>�vvh]u�vv6��t:���1��(A�u�7�	ѿ�{�C|�Y��譽������]
́CF� �S�������ٸ����3-W��n��0m��0���u�ö�TQ�a��d`R#񡦶�TqT�j���k�u�g�g�!D�E���µ��<�Z�u�T�C�p�Ҕ`'���������:b<��	8ތ8���Zt:3"FH���r�M�Ld=�k�+��y�����_�
|᳏5L��N)�HhFsAa���=Y��t�\�}b�I]_�����d��5km$�q�r��r�ݯ*G�m�k�17���X�%*4�$�sR$��?BBg�l�^8����	��r�Z#��H,��6�9_��	��Ӡ8�D��#+!����P�lXQJB�4Qh�P��epk� i�a[Vᶹ�{���S��t����t�Kt�6ܵ 	y��Cr�J���k��L�x�DS����[k���;WpM�>u�m��f��S� � uݞ+e0L���/R�$���K�+��٠�:ݣ[ʧ5g�q��O�l��6m�U���X�nqO'}�?E�.U�kwD �� `j�ݽ��Y]��J��^Ք���Ӯ�Y#�ʯv�K;�K�Z�n���5�&{x���Q��zO�G��[B��t��J��8l��U���,�L���N�=�907ۚ����"w���<7��i0�!ܸ��T�FW��M�Y�p�S��*��6&x+m��4R�C���	�I��9�Z2i����|���ג�oHqV��3�1n0ɨ^�X1��jpD�U��\�2d�۰J �O�?GX����C4���W<�,�s�$$;>������X�}��'�7G�wp�����(��2؞�F�r���.]Ȫ̦��'a��_�)Fz�.nI�q��Ԛ� 9���)i�Ci"yK�ꃢu����f��.�W�b������$*�6����[�B/�2y��*��"��T�5��O��iX�V�����0Q�c�3��߸7�I������#h]�1�	�P�|�*���M�u�F^P�&[#���g, 1E���<�o)��N��O82is��	��bj�)L�Ѡ�3X+d�!� u]=�WY�7\�P8yy��;\Dk���cR
=�6D� ��pL0�m?���-���Ϫ�Mm~�3�rM��4m~3��W�C�E�/�ИR��oS{>�hSf��ƀ���X�`��i�;����!���2�v�z����^i2"���c��<���F�#9{usRɔ\��J�IH�γT�bd�1b��08v�u3��pp	��|x�Mh��!>!�4h�~v�hXΰ�(��Z���D<�<zTRѓseY["�hr�@݃�5��F�M�������J�T���!]-���ٵ��3U�WAMQ�֨����	�Snᮌꜷ�r�}�@���r�フ�AVl��@�S��*ټKWi�5f�Z�<0tw�������w[Q�=�U�-��{��0�1$�*TA��F>h-:��Z1�0��7$��nE��{�Xd�% �uy�ie�T�����'��5�R_�
�oC�H�Oj� ���?o��퓊�bQL���`�B�n�^��i���	��y�m������bma��v�4 =t�ӊ1��Eq��g諾ͦ��HRX�}�a���E�a@j�2��f�<-0���h�W�>�xxM&��$��K����D�^|Y�g*��8h K�f�렘�	������$�Ǆ��Y�[���/ֿ[U�&�w�i���f��8DA3�8o�����z`jwU34�%�`���:r���,&G;�-�K��5F���Q[7(�2����́�<���V�������]���1�)!�V(��`*���Q�5�Fn�ܦ�![b���c��?��+��!����I�y��h���{@�"ӌ�BU4|��ϺN��p���k��%�QiM=���o�jM�7���.�p�Ѻ}�S[#��O��8x@f�&���腝���r��1v�P!f�y ��iX���Gc�f)�z�^��W=�$:Y���9��'�Z޴��x-o�he�A�m_'���O��� W�iHeS�B�F8��.��^�/$:h5"����.�Z�Q�b��a�sM�j���	Y�*�e(��I����.��b�9�2�m&��3F��8��Kmt֪���N�-Q���-��b��b�}~�q��"�"kJg�E��	X�	?��)��^�8���
��௡�-}���l{���q�jQ옧z=���)Ԕ=���z��i��c���W�d�� Iu�)��>/���:�w��Z/#�AS4�L�%k�a��Yct���e"&��PGĖ�g�=m�L����l1��%��_J�"�J��f�؃�� �|�{��gN�2�B�M���8U�񩰆&R�Q��n���qx�rJeiX l�����[6eE��F�c�ۘ���1!ͬ�3J�gS]A��3�p��2�"����e/� �޼ޢ#�����8���KYy�gs�6�6e��v�8-A��g ��\!P�O�4����s���s}�kē��M�
��	�%"���u	���|p�WKq�N��.�v�@��� H��@V�i���\4$l��.x�C�a�M��8�;����l�e�n��<^|	�^������6i?��G���FG�o���N,�Z�Ю�H���w33����w��.7�4ɽ�� �N���b��{7-G�� F�o�+͋[wr��~
����	�w����3Yg���$F�A���(�緦&����"�lx^\�H��U����S�0ǄdI�z��j�g-��u��8y��_�ů4��Qi]-�<Q���(0h���j!�Y��B�g�-y���T�(�'mt��"��/�f��9@2J_K���&W�ry+���)dlz�$���HJ=��O�&���n�4��'�Q�S��eg��*��4/�d���$�y W�6���>Eb����7���ը�W{���U���t��n�ĳBe�^���<�:�o�=g�H�?�r��]K*{�`��#e�
��5~QA��ϵ�o �F$�n��@� *�`.�԰����SE���10�<��
/�IZ�9SM0���HP+���C6H 3lu�=������ds\�ra����y,}�V�nอ��:��:� k���G>��~N~D ��:U<c��?���h�Wp�*a�E4 ƫ/.r��oȴGG�\%]mfLޒ"j���l�h�Sa��%�oOX��iX�s�i8��o����vZ��<x�F�@\��c���@��@�7=F��)�ɼv7��%��D�8���6�RA��̀���.$��%K�i�e�7td�}�܆h��!���y_Y|FH��7��@�v%0�E}$��#}��|BX����%/�ZR�Q���Q��O<��������&�@g��u\��g��J���<`H�5�@.�{����"[K�Ѭ#X�Yt�!���z�E����dx�B|"��4��,C�R��s��l[�_�W�Q��Җ �-�Z�LѤ+��L>������=�c���(Q���Zg@=��(����-����k���Q�'ti��<+{���s�2�Fgԁπ��o3��.��O �@�d(Y�Q��b��r)�I^s�I$<j�a��}jWW��:��9��&���7*���ў˵�H�Z��	;S���h=I?�g�G:bz���Y2%]�o	q��yppA�9(�УF��'S �o���BbH�72��$��>܂�FT��R֞<Ƿ��T��A����d&t�e���s5IS2�Yۭ��������˱�3J�����1Dg�ܵ<���bJ���H�������芵J����
�1���D�Znm�ɍ[��R����U�2[����ٹ�Y�sЁ�M�B��#�S-�AzxT=��ei�(�U��8����>5���H	G�̎ v�E�������1�4��#�h�e��b�ϻ���TUq
�8�[�I5i:��_�6���C�uܰ�˖�1D|^�/^��+�������ڨG�;v\����S�̿���
Q����R]f@��E�-=��/*s�J_�7OX��0���y��;�Ѽ�����_�{9����6�x�ؓ�����c�ғ]���K�w��ӕQ��|�d����Y�]͑'�/0����a��n�o��&@��~�T�<b�f��"�.��#�V�*���w7�?&"�&?��3�|ت���H ?�����C��n���_����E�V:rdl�99˅��7E�?�����'�49|��J�j|��
�!$�v0L��(?�bΨ�ǚ��'�;P&�2�*��@�1���	�������3K����"�O/���M�1%�d�*L���ҏ}�i�+e�c�����k��ެ���!���=��!�u�<�I��P@����#�:7ΖZ<�9
���Q^�ne��`�p�K��,��ZՑ����U�����͢;XV VZ�$�4�~�$��D�	��]��y�q��
v��&��X���Gʗ�{�i;H��b�&&�E��������p��S�t՗8�{���E�$.�^sro	̎�kxJ��z�g����`0�9��<�F���r{Yd�2@b��TM���C.� Qx�&��!�i
���&�{2Yp��~ܵ�5&P�}2��"{���b[�����!Ą�N��Y ��X~�9ua3�b^.�~<������ �D Z��BJ�e;��]Y�VT��҆���i�8n��ۓ��b2��}�����ɖi���O:��τ(��qsN�8�Y�����V,�{C�'d"��q�.� 8���<��tD�Jm�I�z��qьN�*{1+&��P뗊��~FEe3���,�?�c�G����4�ۦi[���Oܓ�N�c���C�?f3�,+�@1jq�n�"�����1N�b' �ڋ��ǋ���k3!�*�@)�q�`�Y��3�j�م)~��{n�Lrۙ��ۼ�2ķ��eS;7�(E��zQW��KO�Jm���|( 	IOy���� �'6�3鷝S���P�)�c��Uf/��������I�M���+ͳ��/8�,۶��.&j	����!����E��<�sN��K� ���bꋞ��<��c�<������
��Ǫ���/�Q�(�S/��x�R�&����gl��I��;h��o�d������&�NG����}� ?%���(��%*��0�@C����JO����J�iL�c����uT�t�X��@��n�!f���1���s��9��KO�`���1�p��L������yJ1 ����;2�~L�c�fG�3�:9'>$_�u?:
yNn֠�`]U�x���1�>)�p`�"���")�H`MʇJ��e�qʭɤ�6�D#���r�Lz�'����s"�Q�^��Nn§�
��V�7y����%�=�{��6:��i�L��r}qu4�H�go>���r���)m��?�H��͍�W�G�8 �xHoOc��C��쳨"�[�4���OS/�HߋP#�mg}s���n�4.�ś�9H<G�G'q��r;��v�Yn$�����]Eev^&У�-:��En�����C�)�R�v����4�2%v��:��!���gi<�(Sc�~)@9M�٥T�z�K�K<`�V<;?�~��iJ��}(�(}i��Qy-�q%��S�Y		6ls\w�."qG��}�ꫂ�"��#&S��tx���=�c���Y��HL�]�' ��Ob�]��a/b�g݉3.�[YϻXt�=3=� קqV���v^�u��o��C/����)*�8�v�F)��*�{�+�Ձ��RE��z�/��7�o%���/��0>q-��R R-x��j���H�χ��B*%~�z���DBO= @����:!�
��h	h�eJ��Ѩ�J�_����7�	v�LU�j���˩��*yqBm�����*@Ɇ�f
��q�����b��L)rոrS[t~v�͓��r�<���}ǭ�x� '�%��+<�}��Z<}�$����J�I�&mr���| �&IC��60�QM�'t��q���������y����ɾ =���=5�8���P���nۻq; ���hY����9�J�E���a�C�:�nh\��C�"^ct_2ړ�մwj򚊽���u���n:�'i�/��/R2j�;E�Nz�IC��d���K����&8�C��$B�w�:}� ��(�������)����p�0�&�D1��ڦ$����ۤӞ?捩�u��M��z��XO�b�O�M����vWT�q)���|331���l���s���ݩ2�K�-����Q�fk�N��<Y�X=P0#�␅�'+�RPF����G� y꥘�Y�4�;v��19<�쐿��<S^� ��m��-����ڛ�h%M��r�+�7��.�B�к׏L4e��n���C���\N-�k7����!�T+\��P~^�%? ��|�5�Ĕ�I�iU�z�ă����uE�V�k���,��$��n���%.>�<��ujЫoߋ�@� 2�f�W�_�{�n$2��=���a��8p�Ζl�g1F����H�Q��(���)1�#�/W��)u�����'>q�U;K�$�r����H�ѐ͙���T7��l8+S
Ղ��@PB��'�Y
h��&Q�'�d�A����ɑl�LN=�$�6bG�i������RІ�HyJ��=G�T�� ����7��46Z����Čk�V�&��e��	&%�ݧL®������c��5����e��2���ۺ�'F[�[y�Q>	L��uRV�u|X���d���8j���m�ʟ_��k�}�H?�Ċ��\��̈́G��1�2�6[#��DrF�Yt�-�wG?�cҍj���Rwlb�A����,Z_��;����X��=��^"AP'�����Y6?��P��P��O��ܨ_��e.B��e���T��uv�r���ry��k��_�`7,��4w���t�Ht���8�D��t�v;U;mrF9�����8j`!�n�����2�F��	���0���l��lsUk1�ϜFfi��)u�v�6������<S)���P�{v3-��ɲ���+t��Kw�����Y�m�̡.3��ot�e| ?��>X[����V�"�WY�DJ䝺�,��� :�a?~?2���`��1i��%:��k�J��I�}�Z�>�j�f	��h#7p+Ћ���.�! ���1�����g�*�N�O[�v�4fM���Uَu��"ݔYW)=3�3g��͏�Q�hH��U�6/<n4��e]}����H0P�M��3��G<V͋T���6��ҋ}`����i���9&ϛp}��,r�b��R���]Cc�⦂�%N�mh�}��5�E��c���L�v��u):���j:�Ή:�-�f9"I��Yb�!��ނgtwb����R�i�R~s(��H������J�+�Ω��vH����T�.�}k� ���<����~���(q-R�����p碓�t�����kr_�������붑eXy�@R���L��OJ)�S3�ǳ:�b�o׮b���v�����P-�5
���,>���5���9�Q��ӟ������p�Yt���Q�SQ�S�	�4l��1�E��-h5�2�VFЇ�5:��FY  ��>�5�!�¼�NnlzQ����Z1�����7)|���U0aH�`�E�	�3z4�q]]/��c'��_(G�N��ޝ@���B~��]]?��p^���Y���)	ˎ�-����|}�c�0�� ��K�0��zj���V^�!�֮�CV��l�	�$޿e�p��̈́u��@Z�~=�r;�!k�oCϒ�G/b�,��{!;�7�Rb��i��ݤ�v�=�u�֝�Ӝ�����Ħ��j��0�Q�JYG�.Eɳ}<d�����9�I���M?�~?��i@m�Ij�ʺfhhg�2>oK������ٚ�2I��vs~�8J�2GXa�`��JZ��	R�)��T5k���=�ڛ���޹��ȡ41�y[��v�CIg���uNM��*�,�:r���	�C�VC�c@>hz=#��_2��|éB�'�NȽT� g*[?P�HKq@"�	9y�����|�܃C%��H�=�P�ʰ�g��m���̔��Aj97�����<��W��ܾ�eC<e�]$a|7L��=�x��E��{�c �=�VE_��"��!��r��B3�wM�VN_��>�K�zr��>sp�`k-��CϏ�d��Q&;�B~���cn�]R��{ւ=L��{I��`ڗ�ކV�ԙ��O5`&'�cF���&y&o�G�Y�S:wM�cWb���:�T��>D9�H�{�X;���|�H]s]�����$,ySk} �I�6/&H������.�Xi�
33��"����I%׬�C��uwʘk^nOe�u�Yz�$.��'��T���?:�̷��vT Ŷ6ar���5�n8 D7R�-o|�� ��Ȱg���N�3��V$f������ �"�����J>�)��2��1C?rj�\���H.�^��@?�O!����!F��ޓż�-1�Խ���8��t�N5$��@�'���޲_K%C��b���0ҿANq�Kl1��A�"ǽ�lQ֢?9��lWt�ԋ����O��9�r �G���P�u!,�����{���T��'���xǞ�̀�][�>	��*ߦ����R�|��(���rm�z��uΊ��Ɛ��1�G-w�|J�-7l�:����,�����D���N5�tٮѯ���Ɣ�7�^��=�bgYk�k��.�����`u����#��kN�IĜ��/�Ae�aK6��I/HYu9τ���l��oL+钕�L�%MNǡ",�9,o3Q���=��U���v�Lt�4D2sU ��N�J��.��z��C�o3�@ۉ:�BP*�tyo�eK���?��sپo���Hl�����˺&�C���@���$:�<`��#���G帬�p���z`��( AN�޶�n��̿#y/�K��<2�5'aC��JF�w6P�1\�����I�S�ηd�(Z5�xl�63��� (j�_�5jK��k)P�,�)���:�R���,�|��D�CCtM�~�����x=�ӼaCV -��S����z� �%���/���ڪ{��D<�Õ�O��j�w�$��uL���)	���w:�X���q'���|*w������\`�����A����[�S��[8������Ê"�03��k�b��¦ڮo��Z���I�/U�vΈ@mw}f
%�*�2��{pJ��㩩��C��3���4UF�Y��WOCGK�	z�:��M�N��c��W�nCF2��4E�|�����Yj�����E�3.PFb]�M~;��5w9���#S���%M������T��&��@�����N���]�pɸ�9
������l"_�Z�H�DcI���;0���9�t���x�JómcI���W-Ó�)������ѥ�@e�܆����ʒٵ���?�:6r�ͺp��¤u�6�����OD�[���u ֐������!8Fc��w��ɏI'S��c���H�F�{���'#,���u�=�v.{?��Z}�e��q+<wE�%Q��^V��G%��W��|��LuB~�͹6Ú��yeX���߇Q�U� =�g�WfC5��=6?�	�K�z��gD�8`��V���9�6d�.y���u!�xu��<����2�`R�� �3�Fٓj��@S��d)E��<${Ֆf�}��_��Ⱥ�*�W]�6T�2dF�͸�j7�!�N��x=ؠ�֕�I��SA"�m:^�|�]1�ޚ�S����IY�E�L�0DB�&4㭧
�+������{;�<ӈ�ҝ���\	�%��Y0������|,���y8�k�n8"�o���#=>PY�T֨$+�Ug�@��>���RT��a��dD^���d�HmIU@>:��.�f/۱�&�Ϊ���-�[�3�^^���Ve�y�2 �߿(���]�
<����>���T�h��� mom�Q�/!�ϳ(6/� �O��w6 זX��H"��[�J�&�Nm[Jf����i����vM��*?]͍��؄P2d!X����"�D�%�H�\�K ��Eb{�yO�쮲؇h��V����Լ����r�:v t��{�ϝ�pI�(��y��������^�yQ�������,W��<�hM�����3	|���Oq@�9�q7��QiΩ-�ؑȒћ�����j�Ź�r�#&��*�����͔�޽J�#�a�j���A=�>NoG�*�F:���O���)іp�(��a8~��q2��k�-���s�M)�8ϤI�R�K���"�C,{T'1J�J2RV�ˆ��C���;&���2�@�(��#NF-��靗V	H��FT@nmw�I�w���\�"o�Z%y�9*<> �A��>΍�4�N6!�8����ծI��N:����G�$��bA���ö䶡�9�x��厹C`��~7��Pݔ����)؁�49~�e���F�o~#~�kj��}+������n���XTh�����dcXJ�Ȗ���̦�ۛ�9iB�]� b��7���f�>L�v���|R�0VQ�7�K�f���ѶB����dtR�%���p�)4�K̓�E�
�}D}��nB�Yʯ�Kf�V��MR����͔%�b3��%2q�|_Z���`�q���r��`%nT�j��ޫ;$�=��������X��~�3~μR�ѭ�?8ň{�ƞ�$��o.JӜ�� Kyu���k��.��C���T�d2�Z�;�c���5D7���z���u�H�/�ZU��(�9[E�S���k����hR���$7����TƇā�D��4�M�e��zoC�ܮ�,���gĘ	:<��"����w��/"���qaJ���y�=�B�ShE�HԢrPe���r���I��u��%94I((��6\C;[��1}��L��%ɒJ[UL4���1��1��AR{4s0�>�7\����1�Tk�x}�xݹM��&��Q��׭xo��l&�	����@�ԉ��v�� ��a�kŹ�4��(�.��}���՗6W�� ���w�et��s��91nN9)�=���ot�fʭ�P_��G��\�'�	��{ �+c38ߜ��7y<���W�t�g�u٩�-o�),�:pn�@A�o�X Ihރ-VZ��۴po<�|66A�Y�rҵ*� 
f��fj���3P����Sr�}���st�#m���H�DF�đq�rΟwoR�)Q:G8K�}�ڎ��i%� ��!���Pl�ٹdD�]F"����ԅ������J��b�cSwJ;Ks�i�ذ�+���*Y��t���,���2�����Y��-f~,��OivO׽��K��qե��u��� ����#(6�Z�`�rB����/�]7chBxOW� �Ã"��=7�v��#�LU���/n�m�E��j�2v�0��c��O8��mQ4��W��h�@E��yw��P��X"%�\�]Z�ER�m
�u��_���\I�\�h�:�D���fU�@��?/��Q?!�\�����_J�H�&���^�����6ypx$�H4��r\5���Y�?Հ���� %������V�8[�h�!��15��L)��OxĲ#N��duʍ؆b�ެ}�mX\i��R�1-����F����V����(U+�C���O�mKm�OR�6��L�?�8�m��c�OC%+�9����m�P����AtR�Hv��L���^��~d)�:�>̣A�)8���qu�Gu�'d���~���Jg
Zʞ\�z�ee���N��n�[��{������% {�x���#t{����ש��j�r�7��j�7��9�b^\+Z��C`kj=9M'��Y��z�4J�K�>nF��H����
���ұ,5�����`������iā<��i��-`�2�Z����,\_���Ҥ�%+��%�{��q~}@��3i�G��L���e(�q+F�{[U��q�qX-_����L,��蹯����v�z�^���� Ç�m��v��
H�~T� �|���6����<P���ҡ���0�α�������7�^�:̢�H�7&���uŜ!�|5���ri��8�i�uP�@��m�=�xjVwKi^�0��:6�R�Ia��F�D��[�W��{)"�l�0|Nj�#�&2	��ȧ��9U��}-�w�9���C\�8���LЎ�P�[��CI�z��(����o^�r�n���;N�f�)�:U�Ҟh�]r}<Ԟ5f��h{b�����%jј��v3�m��K/��j�\mh�2\˞s���<��z�n?����?� %4M���oL0_A]�������y1�Wy �u��H�ߓ�$�j�98� ����%rʩ,�V�&��f��0�}%i�}��u��-J�۟~ӥꭵ�iEΒ��Z:�� ��Mr�^�� �(.�l�V�y4n9�&��P��*�l��ŇY,+�7	Ǉ�Xl<��R3T 3.�B`J`�m�G���I�]��q�UO?�/6h-^)�f�T�u��ɪ���j?�CW]dHq��ͪ�묰)�Sl���U��s�H!�PƠ�:!b��	j6t����1�Fi���J:k�9g�F>ŗ���`�'�WV���B@~`Y��⛭Y��b}<�U ��?��q�&����q U��ba�xolP1�.�J-��9@F`p��}3����
õ�=�E�	˰T7�B��A؊��b�d$�H ����f:N�kG�Т�hf�7�~2!�<�%�k�W���R����v5��rٜ�	� p״��L�wA�̪7������y�+C�~�.�n/�� H��>K�L[�K�뉐�yj68?K�)���o�Eҕ�EUXy��X�f�3��m	b�Nʳ�!m�zh��X ��NM`k��~��Rp\�0����ٸ	�(��5������.���f�2�����K��G��G�I�X����&*�/�M���A���Ջ뀏d���|us�H���xh,�_WTE���������ux?�&�+)�)�%��� LY�a[�L��ċ�}?9%Zc�������g�Kn�˺&C�K:ʚ�ڽ"���9�9|7��7������4�P�'�X@A�]1_A��JP�<�j�ʬ�^Tu1��z{I��p���Ȓ��AV��*v���rc�sVr��؍lS�90�L8j^��ՃEo�z��
�0Q�#qgu�1�*6�"�jM�So�5<Cԫ7�hJ"E+��� vϡ�n�|!�۔J�$*|�����W��
�HAD�4�m�_ʖ}���F�w^(�K���{��m�����O.w��y��mx�D�`���%d#�ko9�#����QE�A�`���r�h��E!�VOӚ�ӗ�����%���S%�a�*�U�eP��^�>S�V���g���P?�'��9�ڇQ�=�����mzb��8mFj���4��S?#�J�J�0Y��	mL�z{թ�������� �2h'���<.ú�/���^%�y^��/;v*�:�Tv�	�y��\�3�,�A|�ǡ�0˓$�\����ڬ��C��ԣ��OY�Yْ��K�
����V�#�� ���Y�1�)�ib��d=`��T��F�=I��!ؚu��ٙ��nsz4N�:.?� ��v��r�.�=�r{ ��IM?����L ��ߋ��)����Oa��o����8� ����;(e����ĀQ�J�ã�v��ӛ��>ì&����S�߱�*%�;]c���/#�HZ�D@��r��&DM<���z�t/(��Z�a`<è>�4b*]ۭ�$�L�59��x(���4��>�Q碓	��H��l9\�H.d厑s��aT<_�Eˮh� ��S&X�&�p� �n�?�T������E*+��	��Z>�B�����ؾ�����C
c	�Un�6o������OD�f y4v�"��~�jQ(]-|�@�8TXv�u���uk��=X=C��V�i��]�䠱y�=�h40j;l=��<2��	��O�����V��W���6�0j���>P��f�&��/�做���plH&�rD�x�Q�|�H�5-f6����!,?-�?�iL"���.��=�^"�I��2 �O>�h�hj�QK�UR�g��i�|I:��m���
 Gs+��+���W��-���޽S��;�{a�\d"�Ց���uh܌m����Q�_	agI�>�m���'�i�E|(ѭMAO�W�j�܅kk��~U�P"P��Oo�^:M��8�"�+O�ip6+DIa*Q�Xsix��j:��zQ~M��S�Y��]W�&o�����X:��}��D}����I�8`���<��7�1�c׹�Ux~z�?&��|�����5>P}��Į{oK��;Q����3?ֲ�+���=m�:y�����N=���'7 K,G��IK����ׁ�&1�p6�e����gο~w��̳�>�ܣ�Bv��y�"t����8�-!���nAUUE��|I�k���B���A	D�m����awh����r&$�85�^X ��()k�Gƞ���J��߇��E�vo\Ǻ𶩿��g���2c}{lӉf��"��M]��xz�oM6Τrf�c���,��4]\�gP|��,���d��'2��x�K�\c��oO�58��V��깎P�,�r� �� E�:
k�:�~}�"�`f�����p�{~�}u��l^쓀�������]H�S�g5,��&h��\�PQ�T��W~�+D�r��(�kFK�e�ӇA��cY�S�I�$�Qz��WK	��wK ���f����S֕2�QW�^~�g�&E���g;�ƍ� l������A��NƌZ�/(�dzM�͟k)o9)da\=y�K!o����l:fz5@���|6�ϿY��K#�(���u�O:�}� �a}Ȕ8+�sݬQ�����HF�!**ݳK�xm�v��O����$@{,y�����<��w<-��t����;��������Se	|���-�O�2���pI^�����1��� H��T�2�}\bF̓�%RNl<Ʉ_ˢ��f��ŕF߅����>z�%�I?�M'L���������F�Y=�Œ�rƵ"�������1Q��9;zO�g���!-���hJh��j&�/�pZyE48���t�)F:R�C��Z�@nP�θt��������io��&k�m�w��[�P�.�?�3�s��Yoa�!�XU�q��3���_�%8��j;��Ѓv�:�)X�hg�p�fY���Qgh]�.�'[����ۦ/j	!�K����Z�:�Y�X����@�3�G����Dt���[W�?��`k�VaQL~�W�Xq��;�dg&~��Y�\K��=���BQzҞ��[3��d�Y�Ⱦ�.���ia	�q�
�s����ߵ��̐\�"FҨ�<�x�����ێ��x�:�m4	:�`�	�/��?�l�M�잆��WZs�k�0e;�3�g���XM���H3����FB�Jf��
�ն Sk��u�c�36ЭD7��+볃t��,RR@A~�:l�v}-ܫ�Vh���|h/(z�\��BY�nd�b�m��]\�e�x6��Ԫ*��Wr��V)����m+��5��,�tᣛ$��ލ��fQ��/��af�����o�P3O�x����+�����]���O���u����"�]����Y~����*��D�h��%T��)B�i�����?�,�>�������D�����1i�Y�LF%���CY�̀0��?/����9|�;v��@�EE@ܩ�)�'m�w�փ۬!�����HЭV^�*���&�m����޶��=pI�0�0}_,�S�Zk.���c[��/(��A)'.ġ�wP����8}�b?�)]�9���+�&�r�k�H��B��,kZv)��֑��I����k�^,�H��+�|s���-mVI��.��ٶ��o�M-��̊��xG3��Z�BD��&օy9wd�&pL� !�z���PuM��o����]M�*�y��Z��������5�1T�����{�W��rg�j��&k���V���!�v�����c�{�����~k;�Á�،�HF��Ҥ��f�E�ϔѰ���]���!BY���R������b���e�r5_�a��ǁ&��Ogwu�K`Y c�^�ѕ^zC{`���D)�E޲�1�����G�7=O�$��-� �5#�a���Kz�K]"T �%�A[��O��H3KDY2%Ntm�)�O�S�a[���'��y����/|�!�Ǆz}u�:�f�S��@pb_ԕ"A*Ŕ�$���vam>U�A<�.�-��sM������dHt�Pk�n$-[�̓�'%b��}X�kZ�b^�JV����M��p���3j�q+��f�K�OK�}2���ݕ4��x<l>Y�e�ɣ4����6"��3��Ujx�#�Xx���S�Ng(⋋�VW��ā�/�&N���q캔r�� �P��=�5���N���%L��Ʊ�|��:��,����-�1����u^=�����u(�d,�&H[s,�#e���0����}�F�7L\�X�w�g�����:ТI�O�j,�(��e�������n�U'��^�f}�w���.UzN\"̖��Y	�c�Z|����'�}��l,1!&��T廨K����p�V�	��@����c^9Ar	r~�uSϪ�����;�����	��x��j5_�v��H�oQ��O�"���srd�>%ݺ�1<��Y6x�
�9Ƕ�a�r�41H˅J3�������{��� +LP�oGa�V>�آU�C���]�4/�2��|�s;�U)4֗;i�M��.h��T|���c> �*��� _��?�A=���(4�}����C�K@h����l��~�M��R�Hm�1���w������6�t#8t,T���p�)��s���}I���#�'��N�^���T:�s]�G����F��C��,�g��h�m�Dը;��u��E�� u���F/c1�3Q�V�=���k�./7O��ǵY�,�`����S?�.�qq����pZ�|J�My�N�/�EcGı�q���λ���>B��{��<��3,��A��țS���A�l-C�^Jb�Ä�]�F<�ݪ8�XOʭG �T�!k�ם!��Zz��
,5uF�Fp��h�Ǹ&~���Y��~,*�7^68���+=u.Na��p�;|	a���X'$n�zqr-X0�O�N%nF}�;�_���ѵ��9�p~@��5Ʈ�<^Q�]i�����[�e��%��<�V�a���y^�C�`{;u�y�5���e}��{"�~���÷UӂiC{�+U��Hg�eV����Q�ϳJ�F����gۮ�=7�5�	����q�SBb���i`�fB�=����6�g2l���#�gu/q��\o��>wr;��4M�Zl�����+���[$g-Q	�����|N,����(M P�n`%�MC��ν/����Jc�4!��G3����<�~�9���eǨ��z�o3�����l�uIgT��.����Y� ͚_@Q*__�N$j�-7�t2�Z�����p�;-�V��`�O�6s����xR�J��3oh���t��UJ�ֺE���?=j6�6��g�G�ǳY5��&W�5rX���Q�b˳i��I	���EW�:9tq���7F�U�%��h��x̀�}_Ȼ�]�0�0�A����c��襏�]���� ��KKx����,x��abϤI�V�^ 4�^lx����Nz��(��Cզ#�;X�p�ɿ��nq�#�`]��5�=ԎT�w����fط���a���	�!���.8�J<�fy�aѺ�ȫ�F�K�~�ۣ;e�q�d㢿�������ڳAGꝵ=p74��ڳ�� �9<��Y�J�z-��P^yj�gI�H�S�$���!~�+�������'�M|����ӡ�iZ����|�R�7@�5j6�(�!%������y(���+x_k� *�c�ev1rLF�Lj���qY�B����6_t�8jEo�%�vSu�RT��,GZ�]8g%����<��?��M|��ӄ��~���p�ѠD�rB��_
9+	J�z���D�=��%���ݪ��N��o�Fu`���Vvi��ɭ
�T�\���hf	?CT&z���􏭁�Q`�%xpG�٤wm�F�7����u��@�ﮄ���`Ϋ(c�r$>k�`�\� R�����?�:3���C�cS�3�m����m�a?�ú`��QLz���rT�&[ѹ1O�+��3�yMۏ����zU>-E� ��1X��(���D��Y���d+8��M����$xa�.�RE���8�XІ���%�{`İ֩���22�S��Ld����a���l9�J6�-��OߌE�J���s�M�(����0n�a���zV���m+Mbb�th�Y_��P/�3��Ȣk��Ԡ�S��Nk��ݼcp����R��z�XG��'(ouw���.���X��@k�\tR�F*�4��u(1�;z���O�-�0
�bgV�HÁŐ�%�|�ZrUq�"y�i�v����<�Ȣ`>S��}>�"�@�"���Ӑq�;�5!W�!X7y����#���h#ô{v�Y�[�^܂���k�Nw�����Ǧ�q�«��w�����QΨ��5��Dm{�PG�����-��[���5�؉k l�-�l�!�l���y�����e�Kby����7�rrǏ���Y8��r�B��
�.m*;#� �C\ �����udu� ���ҁ��J���^�H\���!
{{8[r@_��[_8�M�z󺧧���,��O�.m�f�I�P3x�^��yԩ74v�@��P
���՘�f�V�d��t�ۧ7�.Z�B-����
D���|t�Z�{�A��V:��A ��~c,S����_#l��UJ��B��R�vS<�����������k����똕e]�Z>��ȃ�Fz���C7"�:�)ߑaP�s!�9��J�S"M5|�/~�y/���NEp2תp\�����Zƒ�ȈJW�>��lzg��1��ݡ��8;Ct3��x�a�$;�ij(�>S�xC#����;���OqK>;�)b<.�)�zi43��1��5�w�Z��~��_�N��)��L��_^ B`�'N�3���!J������Ez�䪏mR���;�/7�
�-f���N��K �[�e�fwO癨7��r�|��I�j'��Ց�y�;4<X���|;~�`��h��3�ht����.҄�ݘ�Š*�b�7_s���E�Hϕp��V��s��tuMmg��d2�Q=���C~jË���0�{l��_Q�H���e��Fq�\��SJS|�`(��ɉD��T*�d�
ɺ8��R��c��r�5�5���ہX�ʑpէ2�F���,�d�;��;y�������@c���nU��;I�^�����I��mo���m�+� (����A�n�x�x�u$�Яw�S�u��s�z�Ĭ���p�j�	!��~�ۛ4c�(��ͣ8�1q�����h4C�)A&dx�mb,ǿo����� <8X-���zQ��GPᷞ���)iz�n��<�k�j�S�OgKp9D3l��>ݐO���jX- �m��D��"�\g�z��Tl����[��I���OQ�bs5_��J�a�Rg/J��%���,�"~��e	��b��8��m1���tr�k�Z���Y�EG��%�L��ô�'&�a �X,lw���E*Py�
 �9\��gw��ޯ���I��@+�Ń�]b](�
����/`��>�C!����sKt�(��1�����qi��ft����\��Eh�U�nL���v�G�����XY���4�#{�$���]�����νm>�{���	�"ʟ��r�h9T@|TG��z.�S�:!���\I�Pj[�5�_T�>P�C#��D��O�RL��{$��Cګ��s�Of!b"nV�W��W���j<2�������l�lM7"�=U~$�lq�,�ߺ�+��X�Qô�_��Q�~5L����avf>Ka��iy�V�LWd��~\�b8�3Y�E��o�V�w�3�_3# ܆6I���LѲ^��n���F�(^`��gO����5��n���da/�i��'p.Z+�Ptr�@I�.��jR�
�������m/�r�i/����w�u}O��g,xq�_e^<UuX2H�݄��r��S�$��C�����Ҝ��K=��D@���*����fX�vvK|��T(G���>��hl�"�4�����A���z{ǃ���vT��O��!�M~����n�\�A���*qu�VX���ެ���5�τ��ɜL�bd�觝Z.�)���ը?<��0��Kx��8�؎�"��-��1�t�g��ȣ���>�x����-|���u9�q���z��Þ�_��o��e�tRFwm�Hr�Q��hv�L�C���(j64��\׵��@>�1��[映�킯B\���L'�W��$��Z��)k�u����ِ S��-iL�Kz��.�,!uh��S�z�����x�s�H�-ta� ���8�KfP�����z�${"J��24~j��'�Nx����7і��'o�41Lf[�dVX�U[��F;fIRO^���<}��$��&�Y�����YB1�mQT��Q�=Xt}-r� V���M2*w��6����p2�x-���a���:�G�#�,����w���s��k9��������ĘW(����-a˴J�������t����:�g^�߆`�Rk�h��,��2�q�'��[�q�����q#w�^�L�^>lH�+gE��+��ftb�>��IH�C��o����FM5Q�{c�Fa�H�E����5Ue�@YY�?�(��%_�쓸������O	����CpiGʃd��&)�$F��������x��T�����H,q����cC�8@�-�=�S2�^GM2%I�Ҝ��
M$�0=�oY&��m�d ��Y�n�K)6Damm����%��23u������]�^5/	��!r�}�w��8�`�X�b�}���6�x�N&��wH+H�4+��ƺ')a�s��� �2rSd�/� ��ƭ�輏�q��/�&�i�NH���xA���193Vk'�(b`̭�ٜDl�5�˳�Z<P9k!z��LG��g7���YK�V�0�E�Blڰ���mS�U=$��>��u�n��#;DX����OTЁ��C^�mX7�Ե�r��NsU��ܼ�!�f|}�rF�y͜�����J�U�2���0b5����m�����\��O.�_�^��PYk�o�:"n�nt[�!�a[�
�pb��%֯YFT������A-RX��qk�B�Δ�P�\#��9#D�TF�`��ūyZ�dWk��>ժ)���ڝV�N�_f:�
I4�4Wgl��<���"�_A��
�;A��S�FYo%��jKz�c�1ˍ�cbÕ�`��Jԛ�s�b��R�?����X�D��R�o�{��NߕMq�e�"���"�L��r���i����XbM,T�xPP�%��;7J���Nhg����ԇ-�E��9k&O���T6j`�v�T��J Ԣe��)���}U��3J����O&��T:�l�Ӻ#rq쾋[�XA�ʝ�#N-�ҥ�¸������,ʉ�.�/o��v*m�׮�vhv�'{%��(�F��ٲ�:��?���)���AV:������))�k��&vY`�mi��Z��u�ޭU��	��[���/��3r.��d�Z<�	�K�&�}�K\왛G�x�9�m�mZV��>���<ۣ8׫� H��+
|�;�[���N����2�����p�,;E-�+w�̍(��.�yz�:��"`Z�D���F�!���E����}y���Nl{�y����V�A�TX����m��f6�-K���6�����7N"��Ln0����P#�׫V;
]���i��a8Z�q��/i��)��k䕊A�33�3y�W��+�sB��u\ޤ+-!C�Ր���t��%���4�8�Lk�qм�\�n�6 󄀮1��K�β��%��"{���ß�m�N��j�43��F��y[��Û��R��ٗ�j,h��g��}��֕����z#н���a������ �+78B�Sz�+�ݷN=��w�0��*U�	lV]9�e����]����Ac�d��e���{$at��"��Z�!��My���g�da&�"n�9�	�M)��\Y�O���],�z_�`ʵK-ɒV͂��2 ��/";�s�d}8���프UZ���Wx�u�+	�.�- �KT��N��U*��'���!��4I�w�*���1o9f?��3U�-(#$q�~��uJ�1KI��ˋ��4�2I�j�5�,��X�hs�[n���8�A��{uy�;-1/57�&jK3��R�7�"��}5Qq-ШdP^>�N�v��1�$1A��p����肃��Å�n��B)X	�{��E��b�m�����5l{��71��4�O�U������i��ԇ�p<�d�a���ՔT½�#�N]���{*E�8�5��Kw�B�
��_���[�l7��%����$K0�f��#���y�8�����恿��S��q�1���qa�.|Gu@�2	��6-nI��D�a"�ڂIm�o�����"Ǽ$`��ڨ\6���#*�H\p��
��>Ѳ1��M�k�pi��&q;�3����L;���/��7/�y��H��t���pE����)`�I]�����҅_|j����+ͷ2rXÿ�f�s�{*+�+��2%����A�r4��(hŸ́w%Z������#�+�ԥ��h��OYo>��Ec[����ܥ�����Y<,��@���+�K����n���C��Gr`�c�:��|�|n��e�6����@@�f��3�sO�1H�� ���Ś�/�����6��K���*L�XK�6��%��<�H������Hʹ��!�IyF��K���Y��v�g�˿�W�#]=��G��GZ��f� �S���;�rƵ+N+9�+�MT�s���q��'�1�|󐈉m�%���w+2�y�G��6��\g�k����N��|L��ܢ �r �kzk7��=����j��0��=q�l����Od|h>ծ#�)���Ԯ�*�ݯ+����<����l�� S�խ��.��w�!���;�~e��֜���BM2<1�}��c�=
6��q
��\��YYf�<8��߯>?�B2��#�EԴ_�I��"9T�e��m�:y4rTd���R��<3
�`hI�K8��}�����E�ӕ�?��60!��j<�j�����s��M�N_���ɾr�/���K���Âu&��qļ���+�?��w���N_/�o���M���aǇ���S�p̢�{H֢4����崫�B�+�|��.���M`z����Q3|���֫	���ɺb��Σ+�n��T�N��aՁ4Bi���/{���ci+�P�0�9c�\��|�^Q��}�����\֋켘~l��֑�+�հ�m�t{乛�����a&�D���s�K!��7���Y�JĲ	dXV?)���R���aJ�Eצ���q��ԋ,as��0�D��+azr/���0�w�+�+���v-�S���R���E]����HG<��|sTvNy7�+^���������>>Ub#����C}S�f����]�:���X�:?��R�O���b��t �m����m��N`�o�����=���b{p���	B��~�sߥ�`%��oCː�ϣ��z�-�ʫ�U��%I�p6)�I�#k�񟶮�m9��k�]c���>ń����P�eo���Oa�� �>ӑPk�,��̯��͊���e��m�~m%�>[�Q�#�>����bK�Т`9V�.s��F�;W6��vg�%�KEpF�$�3|�3ҝ�<�X4��]�^k)t�Χt>�G?l>{���̏�O��r_lFPMd�E�$x����M��2�i��$B�t��-�B(PI8�b���7��]t�<��5�/����B:;�h�'>�=���wp��r��3�R�.;�-���<�
6���y�p�l��b���ן�����AX39s�=�aZ�G�d�h8m]��к�˒.@�4��<M�?�������F�_#����-y��6	���S]��\���]	�l���|�f�l�rv����(h�@, ����]�hVUż����P��CT�03�?�� ���O 0��i���ͤ�]���K6pĿV]�����	?T&6���{*��7;x5�*�d|+TGIw��n��)���R$�`ꔶ���t ��![&u�J��DT���f�����x���C�,@�r�?�j��[�˫4G��9~T$o<�� ��O�'Rd�V��a���Y�X6i�I�qP�,%���Jo��4>�II�M3�!Y~���� �*���#+]<U��lM����1d��T^_����X�`��&��Y��U�T=��h��:�s�Tu ��t&�A�G����^�ޫ��(W]��Ʈ�&D^AR��D����L�Ƒ9�#��'��:��y�-e Z�X36��}���zXH8qo�S}�R�m��APU�}kc��,�x9v\)$�^K��Ȏ̑0o�0/��t�Tb=B꘿v�tށuB���g��:b^]���zfV!�e��7x����&b	'2އv�K����5c���<B�x�l&���\̲>���O��ow��W1` h��ԥS��Z�R��8ot��T@K�@�Vg�M�@*�]���ȅ����&�G�����0#;�G� �4]_����rj�G��V�����dT�9a�틦�X2r�e�4��ٱ{��.��b8���uKl�)8�"2��g���&8�xf������%&E�Q:����W��-y^��Ba�o���>��J�
P���E  ��V�$�U�4A%f���D&����)�m,�E�$���Jt�0�Z�(�_�m��Zd��A���Z>���A��Ij~��"Icǿ��]t��[:�����w}D�鎜�~BudrRz���D����5�g�����?N.��I��s<��D�k� �cd�q�k��qM����jZ�n䗑��C0	����+D��yӪ��E��5�6#�]0��3����+�!���1ן3E���P����B1!�0����g��z}-:�C�d��s��ǢTsK](a�l�ОݤF�{[9`65���z�;o�׭崪)b�M�߉� ğ�ݓ����e�����Da�#����V"�=Z|�n��yߝ*�0��DYv@Q@h�����;������8/).��֠�h'| �!���+^��q<J��a�C!is
?�ne��0J���ȣUMNK�0��&?3o���{6���p�$�vk"H�D�\���3��hC����6�?�/֛��S��ث-{ �
`��¢A�>6aW�m��`�s�H�V۔S�Cu5�À��J��C�q�B�����rQ�6�o���M^��Ӷj/-w4�.O��g��x-���\�������d������j�Ә�0p�5��[dV���sk�>�o��/0�S`�����s\h��j�1��hڴGWs�si��h��4�ΧC`����w�ʪ�>6�N�\��&��5��r����!�:���J�p���>�@"�������)����_Gr"�^c}�{e�o@�J��;}��d�n8�d�VfA]���.���st�ϝ�½�u� :��.�E ����l�j�d��D�R��\���S��L���z�&�hX�R�@�z���?5�;Tc9����)�ͯ����o�pi0V��kzt�~�.,�Jo���� *v�Ge;�f0Ǉ_��;�����������L��H�=@Fy6����ɩ�qb�5mv��q��3U����O��(��rY�0�`�p#�����������͓y�'�� P��̧��v.��9�ɜ��#l�,�� �h��װ���<�*�GeqrsM1��_63�����T!m�ǅ}�/���ڃ�<!>o@h�2qȕy��P��5�!��u�uX���T�ؽ󔙫�����Y����
5U+|*����wv{��]�6I��I#� ��^RKN"S\&�!v�E��..����J�Vr�pc�� %����Lk?\� ����<������d���3�`�F�Gq��NwYo����r��H*ew��WMO�AiC��S�O���g��km�j8��ɸ���* ސ< B��vb���0�_n�\Z?�/�b�5!���[�Z�͆�zQ�a�����zO�'��\Y�Y�5~Y@�6IY]r��1�_�e�I�RS)�iI�g���"Cd�^�����j��#X2�"��! �4t��p-��l�-��̈��E��<�������½��4�k��I����vDjqv�yz���B	v+��f�l�x�
,��W�8򖄕����T��:Գ5��')Vm����<� �9*͒���8s��E�Z����^�`6��!��:B���ο!�U$��@ Գ�ɇ&��Y8u,�Z�vѝ�jCg�����oG���%"%���iAy4ӵ���W��vwׯ��.ds\��������C4�!�<�QS�ұ�����(1���Q��`�Y5�ئF�//����Sڋ�������v�/I��%�}��4��ޥ	2	��w���������M)�S:ȿ>n}�Ym|N��ǿ;��_#z�%b��.�U��dz`�� ��|O�,�g�����V>�B�P�x,�e��7ĉ�׻���!��@^x�GQYў�����KaE&�:{��݋�[;=T,�-������\-�À��ޚ0�[�7���������w���۳��?�"s)�
�r����\�\C�`�E��4���Zԉ|������r�"g\s�]�=�k��oBC�Sޞ0�q��M-4����RT�Y^o?6a�1����1~>�|�.8��p�����.�4}Z��hh���ͫ�m�i�{$kgzM��*�w7st���`i� ����H�\�1��a�F�epz�A�'�-�{w6TK���d��q2�l��G��r�VnrW�pÈ4i�W90�е��K\�;m�Vb!K,�a���a)���J�k�ƤEwZ��>�h�f&���34�8�!�Q%0
~3������d�M~+ܙZy�����<faP�ֹQvC"V��5�EUsD������jY����2%;��g���.�s��7�`Bc�n	@��(Z��{��LPY�[�&��a����������Q��\,!t+q��*f��F����-��:�Ԕ���v�3��0z�u�R�0$�'-@ٍ�[��!����� 5�'��F��P�b)�t��K���v��j	<rSY�u*�	g+Z�J�#\��,?��Y:�2�#ZP���#OA7y��6��w7�ʚlы�;;K#6�g�y���!��U'��/Z��]�b�4b��C�-)Ís(`� �c0G��ĝ���V�ۨ����*���'��s����x_�����ɫ�3"��<�P?T;`A���fV7��P�9v���(�O1w/�\h~��S�\� �
�gIY`'�)�>���#Y�//���^�`��:��_��Cٻjh�b�ð��Q��v�G�V����F��Ps�P��#~�t^��Sw#(�a�҄�TVzl�R�J�3y9�"�w'7�UaL�+�g���6إש`�GNx�#>���Lgg��}mŸ�=*qEEs��~Xo�{	B7��Δ|�5�D��e)G�,V�8��p5���� �0��ቿg]͵A�����|'����j�����u�w1;���(���ԕj���k�?��:���z��\��Cd�P';K'���S�'�`�_"�p�S;�����57dp��Ԫ�y� �v<S�ܤ�\�<_^<D�:���f����L��b�#��+{�ɳQB�f6(>ݧl�xM!6쳄e���^o)�,"c�QN�8PgMޓ����h�/��r������(�f�!C�*�V���w�a�@�,gˆ�J	H�
���#����rU��0>�(c�q��t��ξ"�S�|��=��u:bW�7p��vo���ZhZ���d��j�>��B4��j��nv3n\�F���»[�X�u����g�Hke� �� �X	���o��aωA�&QhIE���Ѧ7�%<��j���¾����I��Hc>>5��_�p6#�l�xk�.�ϛqLgFF�����
J�'�d�?�O���<�ztd5	�L:�rԂ-�5���c��\d%�����Cn�P�1m2����Ҹy�*����<��Xg��,�#�!���,e�h���zh�
N +�7���psS����R�ݫ�VT�&�-S4G ��u�
��'N�5ώ��,���9�ydmz���_�;��Y�RIR�+�	>��2�!�Q�/�t|��VѪ\Dר��\�X|R>2b��YQ �(�(bb�V��}��o��r7�2 B��r�&��cH�ˇ���8��Jo��'�R�����������k,R��O�^٘�P�Fj>'}��d��dp�����}��}F��㊐Q<�%��DiTm^Z.b�Ů5 ,zE%�ŏ�M(sg+Q�OC!Q{����	1���v6�tK��.�����m�c?��C���'��n����2�j��mM�#'�_��ژ �b�k>RK��v㩰<ң���o�T�ks4�(���|(���u���O4M ��<zm��=�#�r���� �cxl4���%uU�e%�;�|���\H?�K����(C&��	����-��(\��#b����
ae3
�[�����o˴f�{KZ'(B�\�hyJ�����'�RL����7��9�������0��m=f����^�HI�k�3R)��$������*D)�ğ�NvhB�m�c��YSӄc]3.��w@1���	���Łb�i�#���D��̲�	�99�󲚮�P�4hc�k��q��BTI|$�D`��dC���Ëk!R/�s\��v,\gܬ�I�t����EfG�La���8J��0_8w+�v��7lI����c��;}�>(����5��)
t������]`ј���qf6lkxGvV�@�ݭ� �&̾]R����0�N|~~���`D�"��%��X��|FD�;��=h�+����ʪ�b�9a~�v����������vX6X��'���_�Y��b2���V;ѓ���]�r��5�9�NH�Ս!L�Y���(�Ӝ��GL���B�Ίv*^w,�ޗr�z�Z��xڟ������U��	�
�^�q��;����s��85����#{"H�e״��&�JF-
�:��1X	@?�C�z�ȚK�'8���?�ۭr۶�UYO���9�?��z1.Q��4�G�r�m�G��Sb{�uX��y��.�1�`x[�g�ꂫ��ED+��&{��|�qV%T�Ure\'��S]D�ƥ2=N��@a'����0R!l���>s�)�웸O u����}t�E0�ʕ&;�"�$k�\�D��ڜB��=٣��}�J��|19_�pO���~(�9��9]��ƀ���5�&�H��l�7O%6+�r�sN�S��ǔ���:�p�`���V�*��D:Dt�C2��.��J �#8Sp�� U+���*-:����n1l��"?;�"`X��EZ�){-���Z��?��@c2�7���>��?Z����p XC���:E͚�̷[E�5ϛR�F}oƤ�z�NxJ��X�4�S�@����M�M�NGA�jM��ja�d;�;JNW�>�c��)�a?֚%Y��=�Ḃ���1�%���q�qW��=����j(���f'*e:��i����G�$���L�ɡ<�<��`��-Ss���!�J���w����Q0�
Qp�����*i^}C�7Og��k��z̨`0 ��J�ۓŏ�{����c��1���]�|��FF6=��sd�Q�۷��c���
������T:��x ��n(� �3�!�6^I�#�sk��6Zz�S֞��ν���&Px�݌�uvt�}.SϽc��(��hpɷ;~F�!A�t��,&H$��΢�m�bN���V鯶q.U�,�V�qP�?%�[�����j��\�:��6�#^V�>�:6>�?�3��K_�!��8^cG͚��]�\=��A�zjƖ�h�m�Q ������>#���r�Z�n�@c`R<[r�Jb�K!�י,y�U2Nc�!c��̏��!���a-�5�L�6F.�v��N͛�eVX�q�eG���:�}��~����������K�c0�V�5���z�fw���h���yNGQR�����v��Ζ\#�p�Y�U�q ���:�Z�
�g�j�@�u��̟RtK��+޾_���t1r	j�5̕*[�>���A �J۲ԣ]��j��=���/��W4�;�k���Mľ�lb�*�j���ک+�EÖ��:YW(�n�"�v� �$	�o�A?��ڔ��j^�&�:�+4�?�YA����N���T$@�GF��qIg�I���[`��q)�Y~ ΟyqH�
��Z�Ś�o�A�����7�wԨR&��iQ��E~��#���D���4c�=kX���M�5 e�&���!�(����sGZ�&�R{L����B!Q1�k��am=)�>Np����&V�J9U������,��/�k�=Ab���4��nVd-MÐu2Ț�^v�b}l8��"Y�=J�|����"6L����� Y$�ge��+�RJq��ik��ە�>n���^b':�ڴ3��+��u�9]��~o�Ռ�Je8�������f�����A���E�(n�t�;��z����I�+i3�u�F=9ZI6�@D%9��|O�C���$�r��������3�/i�<�>�%/Gp?�Vɷ�k"�����+9���
l��1��EU�cbf�km��:u1m�5��t	�`�]�L��8Sh��H���Q�_��phK��(*W��/�<�ͬ�e�2p/iKQ�F�WA��uO�`7}�=��V5�e��t�����ő]Ww�8ݍ������&p��#��Rl��)k_���7�b��w�.�{����1�Ʀ�G����l�3�d�2�5�J;R�T
�������2Hc5jTD���w�~o��]��'V��5{��札�P� �^�s��7��o�懲�	�A�z2�����X�N���Tr�=���T��yO�.��{��RK��R&m�@ű�E\����w ��Ŷ���j^I{���cRO�۴���\R`L��{v�aﲘ?��\���ő����8%�M�<�϶��A�Ev�t�%5�0��F�?QSaLr�l:�ݲ��a�"�a���C	�r+�}=��#�f�m�0٬DgΖ�Z&ީ.Q����Қ�`]�����}v����䞳Yi�d����ݔ�o���JV��~��rtG�іOR�ɞb�t	F�!�K[e����\�v�R87��5�e�_N�`rh���{y@�'�y�FP�����^�%�����������fh���Y�@bN��jw;K/��>cQCȫ�q��{���7Y�5��w����T&+4(T+]��#9�����m�@KT�vJk�Y櫥��.�Z�$�������o�`�;>�(��03��z7N�������/��d��a-��T�W]�Z��h%pwit�j_n�p��7�,O����s�q��;�:�)pE�j!�$���[�x��}g�/�r���\��l�-���Q�0��N�X����Kb_8.��'�f�a-΢Q.f�ѱ��S�AA��A^iLU]��T��6�L]�/�(p=���#Yڇy�ic�E�����)݅KY��g[V���p��FXcZ�������	�WLђ�
�T���*%�:$s��f�����@�;<S�c�%a�|�G1-��|FPĈ٩����nП���y�X��܁fnAM��j��!��J�)��U!����qb>�m�Bcud�=���U��^51�|Q u��B��JePL[�t��A�f�p���H�n9����"b�	)��u9h�����$��p�(ۣ���&I��^{)U�JIq,W5Zܖ�R��O�ꏑq��^O�F)W����	~/�<��g�
Be�f���ы�ĮAuG{�:���M���Ң�U�u�3�U`!�)�ś����p���	�\�̉m�����,k�֙�EN4����������n��7��Xi���������qf[�޹��=���o�C�W����XX�#$�����g��z�/=Q�Ih0�ƿ�Y2e���b��������<N>�y���LA���}�2	���S(N*�Lj6o�j�g5�g�ax��m���x�]��;?�z�0K����LO�o�Q�}����B��OV�`��q�ZW�1�����O�ځ���/vY��,E��Ҳ�nϒ��XcX��-�)%��ͥ�w�CQ*�<�uVs�%��q�RW��7;W��5T�V���w�Z=�J��Sk���.P�����`�'�L
۷��H�l�\��*:4�'�Z�Y*c���m[��� ��r���yq��F�K���$XШ � ��f/���/p�O��Y��1ᠦu3,��eP����C!�a�1�v�g����T+ֿ�Cy��%���A����s�+0ۙ��2O��J��v���I�B�?�k�����e*?
���� )�Y�S�ȿ],��[+���_8J���Q�X!8a��<�����`�l�m8���Fd�^ɬ�s#+��m�ܾ����`Za[�V� 3FI���j��P�ͅ+F1K Tx��PQ�_�eٱA��Z#8w�����=�ri6�8��Y�&����bB"�E��S)ږ�������b�\;���ҘW~;�hТaE�\���&�u6�,:��d1(*�r�V'�Am�_��9u��O(�?-�edؖ��JD���j��#d02�,���kT�:3T�O\�]3��ֹE�(�Y���5��c+S3#�ҹ�����ĕ?��9o[��hf�����?{�@|���Q��_�tl���hM�z�=��|7;H$􌆑MւV���^�=���A�T )	�7�a]��x�L���6�b��I��Zb��6�c�ǌ}��E�u��� ���B����i&�kAhs�t�L�ƒ���$͛��� ����V昤��w3O�I��$�:)s�$Q���Q��D�..�6�mհʲDy��d�,��娐�HJ;�a>)zƉ���0��Z�U�̮1n�4�-1�S�r�zg=Du@a�L��ƅ	�|`�?�G䲗��$��_o�(g��N��l�d� � �΍y�������I�n����#���9QU�\��G�N�1�l�L�o�xÿ)�Po�v �p�"���|%�'��L��'1`g:f)����_���s������W�"<���~��I���sP�;�����?�e��P�B���<]�0�*��Tǯ��4��T;�z���B�f�D�"bR!2���:��(i��Æْ���u2���n�|w�Rx�p�O������������5� |��,}�Å�VR���X!��-�p�n^{�H2{)�K�O󮌔z��y1���
��t�J~��DD��(��#ek�V �����˝$�s�k�X;�b��0��^zIƞg�˲A-ZGڎS�]�"7D]��&���^�tB�Fg����NY���F7�%���P?���*���T�&�(H��	7�w=�RO���TNx�g	+9�8JN`��}��=+ɒ��; ��l�D����3�|r�"��)��I�v��x���Π���X���5�簡n@�N]_�@@��E�@Ԝ�v^������O	�A������A��X�_�%NH�,�3�	�Z������t.ðp�Z�ςɺ�u#���G��\k�v��#��N��eI4!�O(�$��1�U)Q�i����Aq�x��
�C��� ����O�-�@l�v�V�m�W��m���r��&�m��EO��0^����ɓ��4�xƶ}A:]�ou^�@!t�'rE4�I������@��-����V�χ]���p��� i���P��8�:�+��q}�}�j4&�-�$�rV6Kh[@LH<� $�8���6ȺC��9��䆡�Cs�F�7�<Vm�"'Svy��~{��M�`+�R�<��m(��译;�����-V\�3q�8�9S��!�TJFK����4�A���+�$~��DUp�[ǈ%��ib�҉5bnL�1&�,�詰�X|K9��|eew���<�skc����*�q�x�ݞ�]��ef7�Q9(����w�@�N�eD�IYř(��o�*�l�b��߅^S�g����j��ھ���q#��v�钊Q�$1X�4'I`����K�pL,��M[�$���Q�$�ΜO-����@)�w�q���/4�O�Q*��x���R�����U�o�>r�N��4HO'�p*����'R/��p�<�*��g�X�OϺ[�fu�M	u�ߥ�m��>�*�x��!��S��3��p����|i= �^؅���{\2�u��̖-l�U=���7��3��}0��NjöQ���d~TR{�w��o���^�.�����J��QI�(Ox{��aq�8cM^{�b�dH�u+��5�E�� �Á\ �K�	������Bu>�Q6D�,��2 �D�aX�ޘ�8�5@�{��冥a�!~LG|Q���__ދ��'5r��O,1xPh]�rz;X Ja��GR]ҏ^��6l���"l2��}����̄K�{��e�vbN�����O��	h.B�-s��I6�R,2$��P������DA-�Ŗ������"V
Mv8�A`���5WI{��>����^�0�g"r�E�$����I��f�ٳqr4lH5�<]}�����M�L�~*�Z�r	���k�%]׾�-�g�q2���k�Zƀ]��@�H�}՝D�	/H���n:���$T�?֠"�����Y���Q5��b�\,�#�9U�!�Y�E��h��L`T�"���+�w9���*A?��6�IY�1�A��@]S-=B�DyK���|e~
ߗCr����D%� �Y�^�elnC_2 ����[��o�A֧Ou��V:���ʦ��<	~
B����AO����rrXo%/Ӆ5�1$"q�<0�{V������A��@Wx�ΑDY�'Ko�#6�~����^���&h+��?�����}g�@����'T[�?���]8���1�XK��_�6?ծħxy�7̚�֨����˥���3�$�?��	=�Mb Kfg �>���v�����;���F�d�Zw�D1,͍Z�-�����i�ȧį 祀:5��=��lX3/@�d1PN��rwQ��L��h�L$�I�j=2������.��;&�SG=L�Q�7�Fͩ[�cI���i��HbA1Myp�s>t��L@/�V��؀������>&�I<��DP������Va�ʅ���\��b]DI.]Y%�t����jHYFj e@�����U�ah�h�T�&�,il��Hw��y�⪖i�k�aF������Kr�{�A.L�;�uO�{���">n��Dk�S2_��tA���%6�,S�]K�����|��T�8*���j,���%�$��>�J��D�B���k��N,rU��]��(;�*��V<�X]�p:�wum�/z(�|kb�F�9��_ cV:��:��eE�+t��m��6��tF���/�
�:�I���E����!���(��r韚c$JsD�%H���[6�+�,�㛤$�V�u�G�7��M���'�џ�R�����-9en�:� V]�/�z0t��e���-�Xm���}�?��~w,Ov��M�WkN�'�V�Z �Ye�dg\?��j���k��aj�� 8�����AZx:MBY�^��L�1�)2� ��.�e&�*�̳�l����{��|k�.�b�Z$K��;br���4	|)��eQ�4,�GJo^F��Amf\�V1}z���э�h���z4b/Y��}噤��Ϳ��u$1=E�4�m87;����/�$���w�;�iXܒ�'�R]^���Y0��2R.����Y��d~�44�o����i�s��wa�&Q�'L��)H­��v�YQ��s���uE����G$�	pGȒ��*�\���Mb�nt�Ʌ�y����[�v�R� me�����\Č�g�� 長r�%t�_6�n���n�\]�:���e&�-��B.1�Ќk�(y0�t��
��T>��hD~�@^����>ر2pZ�Z���"��m}�ɘ{,E�|���j����]���)_�R�Yx�~�w�)�N?�{���^���P��H#�%FDF=�9�t�V�챎���������NQa�S�95�E�ӂi��枦}ׁ�xs6��\Q��e���h^d��+���w� �`~bpR��D�M
ox �J�pD��x�P�2�h�G/�rf^4mF��AU�M	nRzY�;��]J!�%���^5k��'i��ͦY�~>���4�<}Vၻ���ͮ���ׇ"��������{x�~ec뻟B�0�L���1Y�N@O���ZQsY��GI8�c�hݶs���9��&ƭ$e���֧"!zb�*�K6��b�2���dx�g8�Ѿ�D��,J��}?�{�������߻Ϲ�7ϦJ�7f�����r��jv�K�_AShM�K"���W����M�=N�{�ė�EoN˲#�ѡ�&�Iq���	���j=���4��4ygѡ�s������!�n���n�菁��G�.��A���@\�nj�#�&�Lm�"��E���y\L=�����P��R���6@�-y[�� 
��	���P��+'m��dW+��9[\VzN�Dz"��_悤b�50��tN"�}gT�h��X-S��޿�ʬ;:(Z�b���jA��g5-�&���Ib��'�\j�J���Y���m��튨�#�
[�=z��3`F�Sդgi |��p8�,'�p�W�u�t+{��ԹA�ţ�AGy�fԇ�c,�%��w���M�IԒ�����)5�����D~O,����E<Zq���y�	�4�������e���pF$�!Clt"�&/�BzV�j���9#�Y�~�#�����x5�~�kǂ�YP�Mϩ�Z�!����	���c`e�شf�c箎wyd*�b4�Bv_�#́y��`1��Y��A4���q�� �!q��`���h���Ntz��Ъ}d���gn%c�̉�5[I��YpZԮlgƻYx�H�TG������Q$Z�}�c�x�#�y\ ���C7����<���<"~ݝ��˔ҽI`���Bf����f�_�E��f���3+*I �T"\?vu��(I�i�^nD6��b�������RTb�>���ճs��@�^l'�\;~�x��	��(�o��g��͹�L��wϟ�_�Y�Q��wo|������n��˳�Û��(? ��(���e�-�dLϪ�(@��6}@�R�	����^;b*�#����:�x:��ZD/겏ꄈ/��g���-�>V�#��V�*��O��J/Q���C����q�)�pVSzw�����2�Nm,�$�k�x(�B�����yӱ� -�3�T�K�Ѕ�(�@�D�����.e�O[V���1Dj8��FQ'G��Uc�?<N��	�� l�޾�cM;�A�����-=�������I2���DK� @�kQ/�ڎ��(>~Y{V��~���m�b�&�'{��7��-�R�Qg�:F_��2�Ak� �1T�~`g�P=���,�S��%��,�I����+9��(N�B����������@�섍���sS)lHR�{M)�V�T����U�C=�xP���F��>0d$�ﯢ�+��޺��8Ь��L����|�k@�E�b|��w�N��uR-4�1��j�_�2�MA����(�=�d�߉�����eɇ?�w,��(��q۹oD�A;�WN��,��҉�<��$x���T0�����!�G�@�q�����p�ت�Y3:�~�Q7:�xr��B��ki�PgB��� ������.7�ly�u� �X�D�ݜg >�X��X�����c�K�
�i����-(�v�x�o��b�����g�Ù��F��Mkܝ��*}Â��r$� ��*Bk:ZVM`Kp���ZG0� 7�Lw�E
	ۥ�ʢ���
?Y�@���X�D8�� ��	F1H͋#h΅6�g]��AၫW��uYK���(P�x�)C��"O����XQ70E�QC]�g�eЗ��g:\���Sbj��Jړc=@����?0�k��z)�R�kn��Ӵi�n�ˌ�)�`�S,�"����:��.�*!)�A�їR����q�z���咃\�<"�i�&qJUu���f3<*8��Z��{�2u#��HƳ�$PXK�w�Ь��c�����Q��[P�z'ލ')�A�LE��W�s�����.$S��궯�/�������3{���[Z�����l��1��!�y���2�c���ު*�8�'�~�s��Ut�<�\��.��V�ܥ�c�� ���ݢ���z���3o��U42P��$�s25��>ۋDoZ�'�Vr�jsh��m�ŉ傖V����\�u�b礖���N�&�Ӹ�d/݆~ ��/�k��*����<��AݒjZ���܇Ep�a����*�p��<>��zc�A�Q
�A��81
�����r�$��\3U�IlT�2W�l�K���]�DP�V/ag*��ZG�}�X��c���`Iq�$o��G���(��{9zL��tDm�ߗ�W���. D�1'v .i�:��P!�J��W>\+��i�{հg�@g�P7�(�#\���`�$���5�tY���- ���ֈҳ���t���Ɠ��6����o�,Z�}�`y��T�DXE���
rcn�,�EJ�ܽ&B���Ok9�.G��eTr5�ݤи
���J~~��NG���e�v��J�2�'�^�m5��T-ˈ��
֏2�k=�t������]�v��4%@��Gl�0��A_����<r<BR4W
����d��o�/!�Z��>R6��`����i�2���k D/���_����p��V�<����Y�\'�5����j�l"�95�PsK�z�؉��l�9��
���bY�;,�<����v�Md�o����P�.�/��Z}�3C5ۃǕLZ�ݧm(0�e�1��<x�A����Q̌�Ҿ���Ѡ�![RBD�����L��?|Δ_z}u�-ЬB��D��%*x�4x8���R�8u&ː�l):��s�ߡ�?�L��A]>��2�����;��x"�΂�Z��6� �� �$���d�R$SP�d:�GWd��h<��a�U(��<7�7����E��~D?��)�cV�9V��J.(>F;:�	�s�	������YDƭAD�Ji<��1�p��{l`�}.����z��"բ�؛�T	�&���'�o������\�i{����G,�N���e꘿�8�x�����M�L��L���wV���+[.�M2�"�)����GoL�Jk9�<_�.\�,��[,E+���B[���Xְa�bZ`.g�ͿX�tֵh�9i�W��l��H�nh=���7�lG��_�6r�V��M.\��GX��$�h�OX�F������[\	��+��j�,��oS�l�)��1l�K�oD�:�G�C%DJtO~��4�	�"qE;�K�ӡ��	�=��y3�o)��i��Ʀ�Ƥs��DĺgM�!�~�C�4ƥ08l} ���5<��W��Gz)��=�?/���s�g�~9��ˏscU%�[��dg��3��&<�ݜ�9�q;��wB�� �RN[k*����¯s��)D1�D��xB��H�&�L��)�
�l%g:0ئ,9����#n�"gC�Z�8 mQ�Đ�&��!0�հ�C�{�M���Q=�AB�5�2fa?E��!�=mB[�����S~��_Yd!*��F�;�����2�.�*z��O�p�lsqpRս	�1� ���S&��銐֯y�N5��w��c&�$ւ&Y�ֹ�z{�1[�����h�:j�T��<����y�E��	;^�(B��i�U�&9a=	`!�D�/��^��[D\�x	4a�Ԃ�5OJtP'��0�C'�<P3��0�&��v���Lڣ�R�s^�rRC�wzQl��,5r�}W��y���gtE���cL6�n��zPD 1q��z�Fu���#^,���7S)���n�.I]5���e_������r�?�V���Ǖ��j�d�a�z_�E;��h{�j�e��{[RT;�ŇL郗hͤ!]���6}��Mo�'�%��#�a�t�c��Z��z�8<N������^9�fZJ�1p^S4A��da�XL3��)ն9���WZ��kY\� ��C�}W�Z�IU��'�ݗ������ iP�����_[a�����a$���F�8��.�+�jڿ�E]7���eX6cS'ƣ܂�;��u��{�3�|"�u�18Z6�HN`1��zE���?H":�a�W���j6�`��Z�cgR��RoI��=C?��̮�q�
8��M��m����P�@Et��j'&�-pa��p�NI,x��_���CHbih�>�SZ��#oc��E�5D����{�^s�-HdqZ΀ܒ�������~E�� 3a{��"��ߗw�:8��q@�b�TP��ӓ\C����K�7���U^����\@�~�B ��c�B�[? �ȑ$ ���m�M�����!-���M���G�v���w�@ݐ���4��}�NQ����BZ���N��-�>O!�tݽ�������^@��֡��+��-���k+�A:t�{�\!Y�xC���U[�*v��,��?������4c	b����t�
&��+���ω��;��m���	^��yy�Ԍ��tJ_|d�s��Gv�J�_��A[j+C)�~��fA��R���b�� c��?C���'wϯ|fm<\q���WoB���SqA)�[eL˘QV9�"ѽB�Y`>��E��B|�&�Ç�h���U�'?g�!��i�zy�I2ڐsD�6��ou�k}zD�O����W��R����b�����I��f}f$q�KܗZ��7g��]�]����P ����(tWi�$5�,&w>"�sh�C>	3֧�1�خ1� ��l�Ph�X^�ȴ�����јJSΗ|��V�k�Շ�j�U��^�s����o��mյ��,"�֟i
?&�~+G���_�I(�k�^3�zj���/�6'�r٫�w!�	$V9���D��P�t�����B�?M.K�Z� af�H����{�#s�09]�P�*��L���C!1(��-+c���8E"��KC��WXI��
���~��w��H��B7�_�� �h'�kk��������K#�i������_���̳.�D\FP�nx^�2dD#�r���G�j��~׀t;.���<Y�85�Tb�y,a>1��qC�[�"��Z�&3�g��S�GQ᫙�����s'������9L��\�o�VB}q�\Gա���F9�z����E��淺w0�<PO>��KEL�Ɣ�s�č���ǀ+��ƨ�֥?R�t7�dI�0�G��A��~�_��3����&�$%�M�<r��&Ev�!R�ڧ��\CS2	����y��K;�2�{�/~��
>Ξ&guV~�3��<���@��d���+�Z)���7a4a�"�H�$J�"�_���b�H�;�&(j�NgFLY���iF���/����6s��>�S����;���������y�ht@�յ��h�[ηn�I������Q,
��-C������XQ�! ��
u�(�VMQ����@�[F�.��IP[�S�p�E�~��?09? 4�?���
�������F�L'ȫ2���J����x�L�Hڥ���	 ��3>�Q�rk�3��SX@���|j��!%VԐr]D�L]Cp��M�w��*�:cb�x����&0*�@ڋy��"o�#1��$i��fR�v��~��������4%5#��'�����`���Ym���\��D7�l�_��N�iy?�����{���x[���B:���mZҒ�T�`�i�ͦ�m����Q��?J��ks�,5&3�8Q�
�rd�	2�h��y���2m6쀎�����v˂�N�-�J����jEz-@��q&W�l�a��?���P�p��?������.>S�I��lqd��Gm�9���"k�FDyMgu�XӜ��e@�t����l��Id�⁵/��G$��������֐H-YO�=Η c�|Xr0��FFA/@)�h��/��\;d#���6�V������
��R�1ޤL|X��s�F��R�V�!� ��q��|F���s����ȱ����:߲)J����� C���B�IU�`����L*M,G�~�y� �ai<��L�?^�:i�����@�t}<�b�5�	w��+`�uɎ�Դ���l�@�5OL]��k��,��s��է���mD[����?�AWW�uX�4���&O��F�ݨ�[��w��6����j�k�������!i]J���{P�"���ls'��T�B	,�H� ����#�Ǵ�77��|�[NEd��<T��Gx�M=㰓��Q_lK$�w��ĕ���h�t�1�.v�X�f��ZL��(��W�u�k��Z?o{<{5��v�i��6����X���!����!@F��x�է�K���l}Эk�GB��U�:1^�'��Xj��ml�O}��%e�<]O��A�s��2Pe&��Ѳ���ϊD/��܎[�e�b00��3<GN�~��O`�<&/���e3@���e!��h�o����ؚ���X��oڝݣ����G쇋=���7���VF��0IζJ�<�/�dQ�C}M� �����KTK�f�D���j{!\1�+\fj�yc>���߾9�L
d�7�]5��!%�f����&�o�~������4}i��w-�邒e԰J��-�q}`"�"V'#�Ll��htM[{��U�t�h�TrU�N�|�v����ݽ׈f���h�"�iB�<�B��w����~p�_����څ�'���/�
���d�V/�V���m����������i8mС@},8;����`�"x���/���/��|���ڴq u�M��}g6ިM
sW8��2������&b�,��`�o%0@�Y]+��*x���&Jb���D�Tv�k�o��շ��2�����	�n������2���{WY����m��QJ�����x5i�)��]⸡+r��6Y)V��>�<LCx\s��N�^�P�/?�X�"p�`*�C��=�+�̫�`��q߸#W���wf�E�`%�*�@��$�U:^\|�q�g�����m	W�ı% �z?�o�ރbz�GT��޵Z@.M!cBՐ�DA�"Y/���=��(���(ൾ#��|�?�n�$!q��F��h�+B(zƅ ��jB|<���3Jn�ס3������rzdf�יk,y�7?,��5OOdX��C�C�'����� 4��f�GW��LG�|�	\s��Bv����%�h��5݄ImO�NW�zy�=/�l��Ë��\Ox7&�U�;?�ןl�F�h��O<I잕����9�q7�o��PmwU#Z�3�W�������"T�0���9�+E�?p.GKe��uo/q>R�#mT����NFX�#����0�r���&�F~���RIʠg>S�t�4���"�-�x,��x(Abq������i;JEys�4�R�%�Z�7�\S����J@��Z&;���Sw�P��v\�M�4L�ͣ�4<K�I�e@�����)��4
���ÈPd�F��v�����=O�����S�M�{ �����}Ví��Q0��lW�Q$�zͨ��ʗNF�N�����|�#��}�VC��B�A�����:~�+wBo2�E^��Ե-�B��1�3� �%]���OF7!S�cҤ��#�q;�_��
��)ޏ���?�f�z�����GH�L�H/
ﮕ�������G�rQ�^���$C�r>+ ���N1G��~Z���1N�:?������vU����Old0bCDZ���"���������S�xx�l���Ö�r�%w�{N�rC��4��j�
����~P��[.a�n7U��s��.B����B�T4!�)����6�,_	����Ȋq���$�&�J\6�9����Gkm���-�	��#쌋F�E�~+��}#��f�_ۣ/���:V<TwqG�u�ؤ�����n�;���cm��� �Kd�Jp��'ˬ�����i)░+����o���^�l	�	1��'ǒ�^v
Ƴ�>מ�ä;�#��n�4M����;���3�"��w�3ȭ��c8)cl�',K/��6�G_�\�!�����u���L�9��j�MQE�.ή�XQX��y�zܧ��.
`��8�Q҃�@�ss����-�ް����,�h"#�(!o��I'�����"�3F.�h�!�qe,�K��2B�����2���[݌����b����a�#3 ��&e�pb�\G,�C�Uy�A��{���)�>�6��B�- lg�G���ڽ*�l���.�lM�Aa4=��RE\�sUF5�`̹�ڂN�}�z�k����=o�B#�%���G���)c)�
w�I�ߌC���u��<+�TU$}�`�"E��ce:�:T/��u��`p��X+�����45�����[��\eU#j^����u��!���ʋת�����pNt�<jdx�2h�7Clw�mf���vh$��2��~k���^�eT���k\F��
��ߡ�+�����a-���H\���-����	�8lC�/�׽�О�,�����:����ʢ��OEZ�\c]�ĚF�wL�U��T���pZ�c ;������z]N��Ѐɜ/�uR���B��2S'�(�l�f�k>��c���{J(����*-��u��� �d�\E���;�h�+9Ii�p�U8K$#��m*c��i�0�f����x���N�'��r[˻���sf�����) ���M�����DT�������T�D��D�[��E��g�_�J��i�p�u<h��_ւ��;�3v���i��0s��L�5Ì��8��'���I���Z��!:5��u+��>�g�6���GK�'9��+���7l�D*ʙd$�mT��j0ϓ'6�N*[[䆠�l�4.v1�D�e��f��ݓa�ׇ�}�$��+w�	Kn�@�(١>����L�����" E��Ԅ��.�$;��]��7p� ��oH�^o~y�.z�e�s�,ڎ�0I���JF�n���M
�ަ9��_:���J\T�~+��UTS��T(U�s�Gb�ij@�E�6��
G�4ˠ���Uq�����ҫ����z�\��ܚ�W��Y����^��'y`�Ѝ�:f%�, ̔ϰRY�ĞQ�x72o�+	���>ܰm��r`ҫOؓ��MAUdۤ}3�fS�Ֆb" �YAAsHe,:����<�s���]�z�"��&0;����Ļ�K+8R�m]bɨ�߲|�^��Ek���`%�@a[M�h���G�ot\dl�Uz�[u������k�8����q9��Y}¾�{gB�}B0"A~��~m>�_�(�����̸�]4�g9������0���#�6r�!j����6����H��>"�c,2��L�)%�˃o��~��S
��L�C֚&�� �1�O�B�lLf�(���r��.ܐ9�5�==D�.�#�ي����!kG�P_ڐ�����r�`�d�H�϶W�����8���$�qɕR&9�ľ)��j2��p�T�.�d|�U���8�J���v5�]�w�8tA5��:|l�Z��5�?��9N�I���EK���iUKk���KI�I���̣��D��@��<��|�FDt �~n�� �5$n���=�"<D}�x�i��I�LD(v�F�Z?_���	P�=�h�bj���	ޗƊ;2���͢�>,F�dVuD?E��K���𐫀�����() X�M_��
�籆����<�O��e���w�K�m���Xa��̜'�Y"'�+�?��FO�g�܀��tbۣpQx�%/.j0YI�;�_� ��r��Uq���Ђ9����G:�!m$`�l·�O�L[Z�	��(�5�̷����W��?~�nIDa�d�d�)���9��ɭTt���^oLM���jCc���(�<:^�~�F);���T��S�W�|���P��uo�sU?�!�n<�g���k@"܇�y�(�Di�>�w�����՞-�x������3b��-Bԁ*R }�@�Xܥԥ2��c�����l�N��n؅y�yT,�G���e5W�q���`�n	��?�������d�H�M|�'sF���pr��~���C!�D*���a�HZE5�e��T�v�s/
��GVp�,���N��-4��k�jԹ,z���zSpA0V�?/c�:J�|��q�L�8����x��S�SQ�h����:#��dhN��P]xo*M5��=�>=��2��׉X���\�S�Faf����(�aVM�����S03�3ĝf�^3So��6#�ҝ�1���J���e���ڈ�{è'k%A�i��g�08�jt�S��oy��Jf��J��#7�7�8�M,z�CB�=��a왐jb���ӛ�>Ǳ����ۭZ�8�UťD?@���?*d�9p�h�����=�NdS�0���ؾr�� z��G����hX���o��OX�Y�3�'����#�SoM���6"�U.k�Mמ�־�����O�Lv�1�R+�h�h�%"1�'E]YP�{dz� SD�9t"�mPu������1n���2g?��ǿwkP:�O�Ut���;����ͱR����-~���wю�U��l����\*�[aX�J�T�f̩W�^���y5$��镂T������[O饵����)L��l�=��Q@oj���B��"�$N���>_�b�A��4�̂�G"(7	��8��C�������r6�u�Xr�+��鵓X�%�ѭ����΅E��1k� '��ָ����L���C�s���C��k:�d�^��NDr�>��NwH����ܖ}��k��9.�^�����.�C�Q���'���)��gbY��lw����AGܤߞ�n��ȿɉ���<�	�৳�'�
�Z�a �~PK �L(��;X�fV��r���SQ�V�t���^@�w�Ѩi�7�T(��Iֆ���"}��*x>��|�gU�Fsk�E�8��n��
l��Wo.�%
�7R�Q��D�o"�2v�}|eN���^�����)��0H&�I��L�?���&o?��oD��N5-�`�~���`�u�8R8s�I)w���o�~w����K��t�'{�ʋd,�I�6(���;7J������7=�q�By�k_�o�	8�T 6hJGi�۰'ǫĮ�^Z/Jڸ~9&d�� ⛆HT*�D"�R
����&RR=]k��#���5Ɣ�-����|���i)�� �X��������m̹�r!��E�ܕ�tA�������L�I�;X��͛E� ���$�c���l�k]>d{M(�:��
�WT(���LݰT=G��m�fٕ�Fa�F�6��S��sU���jhps°�oU��/qB~��~׹0��8���W��]�ioF9�A���E��#Y�w�;�������ۡw���ߣm�
&�uC����/̚g5��B���j�U�hQA��A}Oo#mNy��X�%B�_~	�V]g�{Hl���M�������'�.>L3�����A��3'a��*����8Q���`�|V��E�GGhn�f=Eృ���S�:ĥ �-�i�b�]6�o�p`����	����$.[s�L0���Q�����$7�a����YB	I	�KJ��� �p�=w�X�|��8,�c���4$*.�oɃse�z��5@_��q$�g��r{�)�1 ����Y���R /�(|��,�V�Ќ>8�b\^Zb�V����w��E׾H�>�}u}#�z�(�_�9���y�'e�
.
p7��KA��[ڏ����d1#s�h*l��&��i��<kVp���~G��a+Β���T����Vȑ
�Bݾ��C�7�IP;@=�yx�t)s��
~���3�l�{���6O��9�l�o�U��\B�����l@�^��:�x��3kz3y��BU�e:E!�^��%x��SΨ��Y��\��y�S�b�̝���z�e~UB�o�ޖ�<H䇾��
D���Uu�
��2l�w��T9����t��.Aw�&����ڶI������F_J8G��GR<ҙ�5=:��bU� @��)Iz��!y�)^�7�DSٙ�p��Տ�+t��	��D8��}��iї��#�2m�b+n�B��F�c�
h&�����SE��Cc�T��d����x+�aT��s�4GE�0�@g�B�Klz�z@e��_����n�q��MS��s�Y�*�(�< ��-#��E��LՅ�{�_Y�_�<���m�N H���W�5�g1ܥ�t�t��y(o�Ͽ?�a@ȟD�1�I����	p����]a�|��|�x+D�l�=�r���߰`��^vR��3�Ȑ��2��¿��%�ng"����ז�2X��CS��c�¸���AD�!8Cճ쾿�Z������n�e����������m�ck?�3=�?��v[L�n���b�9�-�0���q��ߺ��c�p`��N@�o�u�ќS��� s��`�\�6Ze��ر��*we�+��w
l��1̃+�����X~+���U{b%�f
��o�(_�F�ዷk�eA.$ry��{0��O��c��|�[^�f\x��u�K��z.�!6L�K�>{zj`�`�zf����~561#8�Rp���9ܲ�.���}Х�ow���Jf�-�>�|���iY]�pN?�6b�םY�.S}%3xϵ���@��F���V-�v4�`	~(���1�{�4|y-=e� ��N{A�o��"xG[�+ֳ��ؚ_�m�n��⊎�&�\@� c�EX��Q~C?�z�ԑ3�B��sԊ���h;��x0O���V�F�
Gŏ4G2����P�P #]�?r�]{�M�S
�X��F�ʓI�G}�"m?)�NzGwV��z5Ru�+�����'�aii�)隇F�ۀ΅��Tb�T�&%�J�_�jJ���!fog�����Ϙ���SR�W�	no��WWJ5-0���C���RfR=��̰�(�}>¸��p�$�~��M�P�M-?�ET�~O2�jN�z��	�R?r��Ȟ)�Yg0�����f�b���LP�z�;ID��9���(���ܩE�ݙ��v<�7�����!�ôUA�*)l��T�ϔ�WZר��a&����C����v����h{ �p����ő<�O�;$���O��h���������Ɯ�
�f���Aä�އ����?��dq��)�VT��l�Fs�0d�ʳ��uPM�[� �V!r\����й _�-��\�w (���$R���Gď�g�-��2�l�$��^'uJ
�a֥���32Y�"�XV7�{�����X���3y�N������||u�3�G�C��Y��IG݊����[vL��!���TQ���
����Jv���:�G��ϻbx+<��_iׁ���Mq��'��C@�)P��j�7^ą�
s�8���Q Q1%�U#(�Y���-�
����B��!����{�'��z_�vJ�4�	Ws���L�Bh���>8��Ռ*z���o^��pފn�G�=�x�}Ma�ï g2F�=�S�(a�"�F,����n�H�;�o�w1�ͤ7S��W/ӌW�=Ԏ6p&�O�k�NI2�R�O!3+�tZ0׬�0]�vF'���?@����8����:`祱� -�9q�<�(���O�)kM�Zl9�����.�g�����Cs�-�1<B	jW�~l���$�5-+$	W�-�u��t]�AY�%�]�����b��V�2�BS��Z���7�+ހ�VD�x0ٍ�Lu���uP�p��M^RUhB�"!�.���kn�11D���s(�m2�{�C��!�R<��u��R�gd��,HyTD�5Yl�F�]��A��'y���g$$��zQ3�����)V^�)�E��)���j��5SW{n%5�.�ß5�����Ҟ�����>4X�l�x�4�%��:a��e�ޫ�7ve48�Z�?9�B�{5�5��o'�Ab ����Zg�=58HBX9WQ<%�>��ֺE�5lv�e�J��ˬ�v��?�5�[;j�G����
*uw'N�%e>��8p�eO'�mr�({��v��5+N���V��������}#mn}�8���{��vo�j�sO栲9���%he �/(Y1�p�ԉ�,��-�������-휵�7������x߶��Κ�j�1���fn`���o��aT��)�ߧ��f�=d�5[�����{��5O�v�`���T%S$��b0�g�5ee��r$R�?�rm�DRY1;c��*����uz���ަ������}��98�̗iSf������"m=�`��v0��p<�h�2&�?��R	�}:���f�(�b0$/��	he�	�ic��Z��z���M����Ւ�"o`�B[fݒ�� ��������U�}���[�~�g�<lX]�f���A�AS�f�u����@V4ߚjg.O'���lguCg�d#�#�<]�f�׈h�"1D'�g��6:q���t����������ᗸ*��{ҿ�zH1Kb։��Q/��1�Kb_��upɥ+�o�/4�X��b��v�XX��x�g��a�XOʵ�?�����ͪ�2n���s����S���x�"P!{~Ĺ���m]qXݣr� s�H泏?���������/ɽ��´�	7������8��`�x�;��fu`=�|���={������+=��i3<��� ���)����g�l��m�ߠ�eꌊ�`�(�b��lG!�FDM�>��x��==�����Y�>ՁeẶnd;{��@����c))�[V;��ұ֢Ʌ,� ˶�ztBk�?͍���������f#�g���3��:%ȤDk$�o���׀����k��G@���}7�������)�J��Ov�H�>ۘ�֑Jk�n!��O-�[
yX�YQ�&�1��q���ұ9����l��KtxX`C��=�����G��ųp����Hx�4u��a�� �O��?/��m_xK�2�ֶ�����TZ٭�o6E����:��<=��u5#ڪ�M��t!6,�:@�k�	H2|�>.����]���+�b�M�6�nȟ�)�#;��k��I�n*��.��βNo��"j+]F���d�/c�C�J[%i�w�{�m����k��(߳�$�� ��vS�pǖ��ˌ��E=I����jS��~�$�z���D�Մɶ��T��<��谧�`�n��ն$������\��i���3�g������G��D2�IX�g�f;��di���?�OJ�p-C�{�0�h�a<��R��ZM>z`IG��������rYP��͑��F:|Y�v�k�FK 
�S����|�c�{߅
���g�B��e����3�m�:�P	��
v����cmySp����rL�j�i��n���Zg]$���d�E�g�)�\��_8w�ׅ%p�59%ͤ���~{i;��J��a�B�*09��^��m�Ǽ/{��4�a����'���$P�eG�sc��uI>���^2�l.���t'�wGs��/<�w\M>�q���۪&-ɹ8����:�Gj���y�`�[������ݿ�Tw� G�ۓ�T�,4o��m����%��GҨl�mD�Dֹ��i���:��Aߺ7�]xf"?��J�d��o�mN혐64>��;0�Q\f��㷭ރ�c�z���"[Mn��[u:l��*	�%���UsD�i�����p�����`a�������э�6�f��ٶ�f�s:�c��&��O+/ڄ���6���=�g�])�@s5�(�!;��U �7���-y�8�Q�3&�����Z�&f���@���aOS5M4Q��*u�T��]2� �G�lN���q^�*4�/dI�\(��"2�����j�b:j��>��A>�y�oD]E.�H��o�x}�t���U�_|����pV��r�&�ݶ����c�D�|�b�K}����{C=[�3�O0�{�w�əe�oDL��A�҉��+S3,��P�l�f�0-�J;E%v�������7G���4B�g��KM�5�e>�P����)��o��s�!}2��&���J�Ɋ���)eh�eDz���	�@�ԍ̬m�9�$�d�)@ɰn�leEQ1[�������}�U�?Ir���0ՂIa��'�g��������.�'�B-�j]j�;�łɓ?r����i�M}%��n+4����f�}䐋8�#5�t�_8-0���D����2��L�~ֈ��2�gZB�!��Յ��r���s�F���>�yP�y�g5.���/����t�?�4�܁O�.9�0� ����k�F$*N���^�	ǫ��Pt(O�R�Y7�g'��� �s���ϬR,��W�bm3
�.�~����޷ �#��2��P O%65�A�`���XnrDd�;�gbP���6g���E� �_2�C-Fl�Ȕ�z����+���_Jt�ד��D�b%�YN���|ɱYJT4���c��m*V"���������o1�� �����2�! ��'��QS�%7dRG�KL�@c�#�Q����le�o�W�FەwM�6�T��.�\N�r+$���ͬ���%
�^�>r[0P��0-����b%-�o��nS����vM�3D?ȊX*{nc�pm�ܠ8�o$O�.ꉱ����<8p~�I$@�C�1j.j�.�n��ʐ�d��.��[�\�W`�ˡ@w���1��|����A8���Z�}h�7�Wt�!9��c"�\J�ٌ�?{�b,.�ؔ�Jc���Q xV��N��0��#�� ,���YOT�#-��M@�c�'JD����[��dx�c�U|��{�bV�0��~��&���(h��V���1�7�r�Iہ\����zLp�~m�eAcV����!27`ᜊ->��w������c�ҧE�sJ	�ǵzV�o�S��xl�&fuO�7�����	�LHY���Ni��vQ-B�,����u$�uJl��X��Z��%�Ք=V
�뙜�DoA�Vjv�e�yLx/�SCN�ՊJ�s/�m �T����x�r:������+lB��>���f�L��$�?��<�ʖJ���_�P�����o+�)�r���tʝz���_�fȝ���[���m���)�XU�$��>�N�+8e�Z
��u�(r{<5ޭ���鿸��}�&�����%ޢ��d���6�v���Ǥc4��v.�(fe��i�vG^��E�����
C����}&�K�v���+9`�T�o�����2��Z��ŻX�	��Dfk\k#h4c��Z��E�)y����`Ā"я���u�Y��+;���&i��U_��$%���9�<�Ǵ#��4 �T���#�L�^�i1��q�,@��UE5��X�����R�'I<(�e�x�ٽ BS���]�o�����
�kf�%x����F�N�T���w@���l,�X����YS�v�y������U>ZX��R�f�Hc�I�� B�b���m��sx���f�����(�C�0ռ��-)�Q��V�}��+KGŘ7���$]�R=n]U�I�v��x&��v�ob'�^G����ଢ*��P�O��#�>hHeK��$H����*��Y��Y�I�#X��>K�upS��8+q|L�����:����q�2Q�#��f�G�=���0$��Io�	��	m1�,���ī�tMV��Pmڬ���Q(�K[M��H���B�����3#S+ɲ�ݻn�ȭ���O: |b���h������Dm�?�a�4jv|�V����8B�ծ"*Gn���C��fس!��/���ꫩ���!�#�5�m�fܪ_��"3���_�K0YR�׮��Ĝ7G��<]��|�"���U��*�L�������[Ş����B��~���8i���T2/�??��U&�+�B��p_�m�#ˇ*5��ɘ�cOo�B>�E�E����tS�ȣ��h��bK'*L\yo���g	.�NkI�UӺP���|���^ߍ{��tF���L��>F��*�;EO%}G�����~p�{��������|V����S5���P�QC�_>V��3@��'�1�u����7��elь #(�-p�o`j���׫.��[�������3I�U8�:��t�~`�H& m�%Ì�oً�bD�������w��H�>8�-�'���6�j��_ܜ�qAMk��kax���0��H�7�|?�X�&�K�^��h���l<f���jQ*�1��o��P
�3������˽U�ss�A��ei���.�M�$LR�?�`�[�8k�Л ��_�2��l�ըB[$0���� 2fe,Q'wo��aL\���˽�]��&�{���6��I���z+�J�E@H+ۚlغ�QK�'�N�X��e*r�� Q:i����U�E��0@��pp��;����2�S���i)��@J����ڝxj#`�2��B7N}�]x�:���������}�nsl���
��F��aL �L�4� |�'��������\cji�R��^*AI`����ł|�O��b�|�o����X�S�F�:��_M��;���J���_��č����y�x���7��`@ ]�r׶	���!Q�E����I��k<�����7�	��%���(|���!*��c�yj���{
H�^�p�%p��G;�d%pl} ���_�� C�0��| ��g�N�`F����R�^���Ce�sj:�+>7��O�|���+>h�|
������B2��dٷ�$�%Dx^���0h\�����`�����Dn>�Y-��j"��3�i�H��oԃ�-X�W��5x|.�1�\Q�%x�l���X�o10kdSYdG\�m�1�T1��*8��`N�Hp���	Af#cc�����U�#W������Fv8��<9������:�aAi�Ѩqd�[-I,~�3i��Dj�����M�Z�&zN��x%W�����+���r�ҥ
@�s]13�?�9B,u܋=ʸ��>\��EN�n&��f�%��(��G?���R��9�r�ʿz���TQ_Z�~�]}��"V��}�l-��:���IS�B;;�H�9H3S���i���ˏ��/�.��S��Z '���E�cT4��%-@s0�=B&nR5�:�͋����J�v��h�j���Z��˺	�����5���ٹ}"����Y~�VK,U����z>�)�Qj�^w��:�2�����	��2LO�N�U >�)p��@�"4�>$m����'����[ԝ.50�i���\�A���`4�-���0G5�ɝ��l�
)^�K&F�N���-�A�4k�|�.?�2�9�̯*�e��`���4ߣ/�0|&��� mBQ�czsu��e�b��XN'y���f̘b.o�����������]�ܴJ��؇x�c�HIoR�j@��eJ�b3 j`�ɷ�@�(͔��=}��/X��<�'���f�3#�.�a�����g�:ڊC�Fp7u����r��š��ҋp��f��-�Mw/�mS6C�q@�����k�cЇ<JLf}oQv�$�F�cx�2�eG[�ǋS�Գz�S`�aM=��p؅&���#�Z�*\�?:[�ͨ��4����aq���� �@����d�w�C�e�^����]�JtSwS�������-�bK�����[�崚�k��n����Y$'-�-}}K�*Y� �w�a��� ci�e�-@d�I�cu�J�\�
ϗz�������?hW�F���Q��Ս��s���M�
g��j�i����>��W�$�cv��p���0��!�w[����_�|?\7z	�οӼ�����6�%����ʉv�}�	=���I��Ֆy� M��0e�6C
5n���&�u{N��Q�ǰ�u�4-��T��2O���ɏOd絩᷅�0����D�X�ψv11�~,�A�w�c%Io���v���eCk��F����$FѬ��Y�9SBFA���X���b�Q��_�"g�{f�@14�Ci�^���#7<�'2��/bl��6��#X���2��L�(�v]�N��߶+Z5A)�2��S�1�,-H�f�/��4ف_��t:98B�p7���p5#���W&B�Qr� �9���ϟ������R2ۢ�W��o[��hfĂ+���ͧy� �8��'��r�e��������:�V|@Ѻg��5��	�F�.�Z]��o�D��8[�ڕ*��~B�^����+��e�a�}oƧx������\HN��s`������#����s��_����4�	�-�f����짶�es9&H���RBY&o*����Q�`�Y5CZe����"��o��B��hk$��W�y>,e?�~ftM�-��g,lF:^�a��7�je�5mY�T�U������w��-�$�r-pGF�
f+�ڀM��҇���Ԕ�w���bC��
�-�䁽#���o�L8����8��c�r��埶�_G`!N���=1�d�A�����Jز��wm�g�Fm�خB@��n��G�s��^��DF6(�j�������K #@7���4�wʡNc�����=6�f���� ʽH(�싕���W��1\J����_ܾ<J��
���U>���3��`LT�F�Ț�Yʭ�:���t�Ҋ�N�oFT��V|\p1��t�`FbB�qb#��ꇫTe��M�L݄������O��-�� >��$���S�����#�PY=���Xl�����
�	���8� T�]��H=���~�`A��L�tn��3O�~���[�� �N�H6Q�%mb����|�ou��������j����3I\�ޏLf4A)b+wB\�dH�"*� e�7]�Gs��T��İv뢕�˻q$�C��9sM�ކ�hZ�)����9��/^T��ǫ���@�b(���8�a��0���B��BBo<p_T?^�w�t�0�l��5B�8Oy.�I�qc'N��e����#V���^��9z2��+�0����`��ǥ�pf�-]Tb�Y:6,�X4K~�����H���_z�4���B$jo�m�h�Q�'���i^��-�F�����huy6�Q�e�;���xt��s���f#cɼ@l �M��m�P1C:�)��Ұ@�w�p�Q���{��f�V�� �r��D��_����r�h���#>b�D����7��a���p����ͤ��;�wľ���G�֖	��Wd�kAf�oY��~q�x��ZǛg�ίz���5���2�a�<��g��w���+�5�E~�$��y�R{����Pִ��chO'vGo�g#�P5)_��38Q���@EIs:}T��YC"���ԛQ�m�ǁ6�.�y�_�H��;�1�x��#�S����<���N���܀��fӧ	�n�^���xAU��O���4��f�f��(�^c�j��.��3E
0��'Yĭ����� ��B,W�F�������y����$P����~�ނ"���Ȋ1��7~���BUd�d���Z��H�O8��vi|��S�wx $�@Z�pa�b�HJ1:K�w=-�:�>yѐv��+�+�A44���.�m���Z�׻��+�fc7�f�Xb^��޸x����s����"�<+���֓���Om)X?,T͑3ɯ}m��S,�_ᖉ���q$o����h�r�8P	��b����և=��4w@�?�}N�j�Ufu��^�:�ǥ�JLFs�6����̭��=|U�E� }�J����Ɇ������/O�O��i�L [�X�O1%�9������='~=�����V�c��J1��d0vp�:��Sg�E�h���ˎ�J�Hwe_ɛĘ�1o�z��&�:63��������|l���ͮ�5F�s��SV���,���n���s��٪��P��w��&g����F��m�e�x�v� ){MO�!lĐ$4(L�o�z�H4E^�������=�c���j\|��A���Ŭ���A�K�����*��#�0�Iֺx��To�\ܴ!A�_T�e�b���"� �%���õA&U�MYͷ�G��30����t���e��8����s'+|h;)Ζ/"H�gI����J�[,���w���`lgis��q�Oa�w$�S<L1�Z�C���xg *a��
�8�͑Hȋ�JC�C{.�Y�{�]H��l~ ��TW�Iu��pu�����t�A�J{|&��8�;E�?�2U8~��I	^N_����x��|��]�	M
�h�W�xK�a��o��*N�A��rO����e�q�a8cr��K�߮�^Nzc{�oH���8:�<����R��G�GY[_c�O��v��6j�*F*���a[bE���<.��=�O��`�Odo�ⷿ�e� 7�k�C$������@��eh����6�~�B>i�y^�����G����<���$�	>���B��.�L$.���WM̢�b��}�z{��q���t�M�82T�
"T������OZ���f�G�<;3��ؗ��x��o���q��~��d
+D��(�ō�y���gκDς/�q5,�  d�\wx�5{��+}���ta��K˨�b:�(��z�5T��1(^r�!�u$A��k9�P,vc$��ƊBLx`s&:M5�������*�'���|]����fcۢ�c��*��҆���[1$�����%����կ��;�����ʣuI���ֿ@���{��+
�%��\���g:����c���=bS�9w���[$o��_h���N*j����!�D�p�rnwWXv��%\fG�E�#����)@��y5�WP#hcv^�+2
��{@�����/
�s�ͅQ��:�jG1J���d��H����yl�ޜ�� ����n����_O�X7�]j�y��{6��������$Տ�؈�\D'o���{���|�8=ƒ�v�>�}�v�����RYg����~G�WD�w�������7
V@��R|�����S�!N���f� h������Kv�la=���i�fM���1�V���"G&m��{z��a"si�%���`�C��0?�7���s��f�3�ȍP��[�HS%r�)P#n�:� ��\\w�T��X%qԘ��3�v�C�å6��c{��?�㢓@P?�&��m��&%�]�B!k���4��?���8R���"���_��Va?t
q�lK�5��R�%���3��!�Ů��K�C�����c0X���2���"^����HM�6�*��p��$��%���q�ҡ��&Z�yUp�I�ٱ�"@�`O�1b�#n�g�R�&G^/ �I�0�܊b���".)�C7�%�w������СkAB۬{�c~U0��oT��ʘ%^�9��`ǻ$;�#Q�)rz��'����m��CW}Fevř<W�\w|'&=�P�G�N�=��H�Є���O����?�s�y�s8�"�^��rwn|r�:��Vb�V,I �RA����mF'���a���Ąsa��U �YB�h�<���I�[C�5��^v�Fҍ�A�&d�O��,!1��L\�"S�o��Bu2H0$ ���3�O�mT��ݔ�d�\�lP��
��;K�h�z����l������M%^	�Q�[�v��w�8�6�/e	<��J��.¸Q��&FU49e:�9~���i5�=��E���߮H��߮*�.�"'6~�<����@���m�Y��:�9�oƜOrʑG%���-�b�z)�Y@D�?��f�>4-BD۷Ys�	kA���"$"dvے�{ �S��K��2+���~�[�f�"5d��Fdh�d�p��W6}u7T��p~� P�Xb�VSQ��+�1��F���$�jM��-�(��c�3��t�0�Z�B��Z� �����q�VmG��w(%�@��J$	U��q�"K�Q�C� ���T����	��!B� ��E(�LOk��X�	�=i�� \e3�B7����?��R�~����=��k���t�Y1���W7��N��f˚�ޱ�t7�SX��lÜL�V���Z���0GТw�c�L'3U�OF����Ic�]�PFAN�,"�-��/�(ǹn�2V��9:X^�K�	�ʘ���e!*��%s߻�6�����0��`KH��Fp�v=�����M��s���G3�0�r��E�ԄckP�Ӹx��VlY�x��D�*�8�x!�ű �("G�CH��/��2�3ƝvS/N�]���}u'�H��jZ��W��oJ>��<Ė��p<�*$�h���;��>8��(���n���-�r�X��V:������S��]����]�]h����ʉ�L���ψ����d������2}C�5�P(Xܫq/�������@�&��S*f�,��1�v�x�4�\�)�n�'%��� �
�d��luT<�a��~�����Ȩ�ē�K�#T�%�xfk6�;H���&O�2֛6�{�Nb�x�B��J�S ��I�<����|A^_�Iv���	��������e/�!O�LR�U��K���RIK����$2E�~D��\�t�M��ѹZ��!8 ���-��}2�4�o�"𙉗���(�CJF7�Z���9�����Bl�4�j�\�4�K{%s��䓦����H⛫�)N�Cx|	@w�
�#��m%U���p��J� ��c>Da��Vm%�݁r��I�j��Ȝ��W��FB/o�H͖d_����j���y�Ҝ��ӃuS��Iͩ�B�΋��h ���Y�K�yqzO�@��롸j��jJ�`W$����Y7q9ԥM�R�H�ܜIx�^a��V����HB��5��ܨ��J��8Cv1P���B��&�e������T�@�����B+���x���v�/�d�(��Eha���O�����}2H2�OHF����gt9�dR�"֯,@.:A3<Z^��j �Y���� ��8�T}�"�5��+>G�J4��q���P�N9�m(x�a����w�G.�<[%�4(���e�-ӺЌ��&`g l)H@Ge8]�R��;�4uwm�I�8K�qWp����]�N|kõ��L���
�_E�2��ɗ�:W/�>�x���
�����D4��!3o(�LntC���Qto(�J&@^��c�V�o�
>�jːh�u�rS*�($B�>�������f%']a�%�AM����jl��ӂ7Q��glJY�qt�W�Y�Rn@G��z���k�$�l?YJɤ].�R>���k�eO�q�`�)O'x��ʭ���WO�x�윢�C�K�����=>�Ѿo��3HS��N�J�x������(��Pfa���~T{���h@նP"e({rV�=Z���9YoI��a������_�@������
p8X��O ��A���l� �ex�Bnc�J��G2�0���``	���Z��B��� �HK���GWtπ�rO�o�8��c?ZU&�w<�m�cJ��dO%�d�w�ӆi��.�1��6h98W��5w�X���o�o��pA�΀<�u��n��
��e?4ۍQ&���fR ���+@�5�X�p����H����QSK�Q�k+���>��(.�εc����-�Qƣ3ҧ��s\�ωB�¸�Ȁ�9R���߻&3/�r�H�ǵ/���4�Hy�bajf�[�1���� Iq���3��H3B~<�7�Zz���������O=hbA�e�q�.��@FT^-Q��9q�V��}���%V�[,���׬M����~����Ю)A�L���G��A/�na�̎����.���%(�:��ҽT�h�e���& Z��s��Ū&:#f�U�>�+̉*�Os�M!�t�w�EyE���i�/�VUg
�� ����ً�[���~C�{�IG[F6���1�9 3� ��Cr
�ќS�: �m�]�b8D2)��8�"�-U�s��^ �=},��J�i��j���y~�UO����&�`��F^/�	7�0nJ���+��B|�o����	�3�(��%���H�A��m	N���t�ٹ�����v�mGc�޴Bx�7|��#0j�-ngk�J�FLWe��,n�4��E/aJ�L*�i��a���)����<�������S%�r�z��,��Xki�6���d�I�?��e{�0<W�o�+�����>��,�azS�W��5�VE?����_�H[Q���MV��/??���pw��A�?q&gر�"���z�^��9O��"��M�����P��K�sL@eڒ���V��b�;�wOY��qR�G}T�<���Ф��J�L���I�t�i���G'�VmU�f�h�2�!���r���T���&w����d�|Qm��|2oȷ�0�D�"wǞ�������ڡ4�8��U�q��{*&�_c�wt-*�G�c����^0ìڡdJ��ۈO^�Zlk���Žw�E)|��mk�CUI�<<�$�^�$�6*j�=��Y*D�j��3[��4)\��XV��L���$��F;���WI�*�z�Q�#�8t��_Q\٭�%5 �AOR�By��PR����u���k/������'�Ktɩm�k^���ߠX�I������q@�ϳ��{T^�l�*2܆��k�[������D�^�=�>�q�N{��%��pڟ�g�U�,��n��n!�=�"X�8��鲄p���	Ƃ6����WKE��k쒡�,e����z���)Jĩqm�1�W&u�xr�^X�>��r�:¿a��:���|䵼h�HelIW~g�T�ʰ��E�I��fS�S�'��z�a�D!�����N$��.��r�~.��zl��ƳïIy�g�ؚ\l6_�����|�f(�Y�y�&�,��nb�$դ��-�MS.u�w�ο�8S��=*�X����]I:�lX�F��P>��c�Z�沭wp�;'�H�b�F+�8N��vD���C[jUQ����W���p��T�.n�}z�4in�Uy�I�.=�������̇C�T�e��ߔ�z/��*�hɓ�.8�$,M�}N&�t�I�i�b�E~�ȸ;.��L�pc"��a��ۻ{����Qs�QdQ��-�6΄������d#y�K�
: u�:h�y�G:�K��EgL��Q��z���ul�5I#�i�LB��)�6U�,��-�/;f
W�ŵ�r��.n<ҍ�
�o����ߞ�kOw���[1'ɘ���k��T&#�]�"��r�s�R��wz|��kl��6�e Q: ��3��m��A@�Y��ڈ�¡~D]��eY�ۧ�� �_�vs�`]�KUnZbA#�h[������V�Q�*c��3&W˟�����jT��D?!��#��������ZѮ@�!-���T�lNuIf���TЕ��[t{����߱�
ƳP��ql��v�FbS}mfj&ȒS�k;?<������&r��X/�"�=>�#�VU�Y�&$|']����|B����o P��˂�O%�t�~�P_��_y�2p"-57v�_5���'�+���,x	|o?Y�rsP��ߣa^�;����J<@�*I���!v;ć����ƥ��N=o��_"um2�ސB7G����Hj�
�X!�����U�u�踑�Շ���8
�(�/`��n��t僀�H�C���9��eR�=\2��ED�Ђ'nG�p$Vb���{����2u�x��n$*w�@��:O-��O�ziYB��C6�0A�CO���>������6���H/�Q+Bg_�����㖇�f��z�،���լ0�O�G�/:���U��@${�!N��,`�WX!/*q+�iQ��ߨ�3�o��o�E����T��L$�.7	F��0-�*�Rr3����0aOV>E�����8:ygr�㗏�#���&����<c����<�W��R��f�/��(O�:�
��BgX��^�-��$� �KrG�aN��t������i�"�#��� HFBɬ�Yњ�Y�݅�ڟUs٭FL�>�g��8��]�#(E�qh�c:G�`�L�*�+��7�j۔��p� ,ܘUT^�C/�:�L��<�Xg�W���hD�ϸ��N�6��%��|&+/���	;�]J�Ր��\)�Z�Zd�lnlxo	uAT�@-<�C��$	_Hs�&LL	���M`�ô5���a�7�@�.�N�J�
�GNr0c9K3vQG�.�p�b�NL��K�7�T�L<�j��E�r�>d���N�ۑ�`��ȡ��cْ�Y�
��.�[��wI���bǁ\K��}���' ���a��ͯ��5Bgeד�l���D����-)o��¬�H���`�wzCC�.��ּķ��љ�>�l��/G,�0��L<�Z�qQ��۟75,bU���Fԛ%����8���#�ծP���6L��J>���mq����rP#k1qB��$�/�̓���1�r� E��3���!I�L��<����-+Ʀ��%ڋ
'�qʢ�Pza�K��|�χj���ѾL�+$ȡQV^*j�(�]�Mp�)��N��O��l�6��;�^L��Y��4�B���W� }6�� ܺ9+�ǶŎH�V�Ʊh����mS��r9�E�\��	�8��a�����_.�&�\�׎���M��S9[/`ش�X=']�/�����{*�%5�tZ)���F���2Ƽi7��F�Nߓ�,�/oIйz7��2�\���{�;Q��*�W'��%�7Hr���������Ͼt����%���߆���i�'f��͙Ӑ<x����B�e��j
̫xP�Հ*�y�a���Ԩ6����L����7~¼5�*)sX������bH����7�W:��$c�%](1Ӵ\�M
�p�z��!��]k3s�wD�Z���h>t��7f2~�JXʟC���	���/(��Q�gV��)��񢤈�/���eν�U�uP��R�\^�O<E�z�E�}�Z}����k��W�j��u7Τ��*�p�CW��|�]���u�K�ڱ��-@�g>��2R���&�n��V�6�K�W0�P��&�0ڽ�!e�tUo�b����6�US��$N胐�ʧV�
�K���3Ud��CAG�M�A:p�"+n���n�E0~3R�u��a�g�0+$� M����v[X�7�w�_������N�J�⺋,Ĕ��mƓ�@4���SV$��ׄp&E�~��*����@�Z�5@@6М����[�S󤼞zr�G��P�	�S1��9x��I]^�!D�_F�� �[x[ �x���[z���
1 ?7�Al�u�t��ȱ 5�g�T�u��s���K[�X_�ޥ5 b#i=r��
�a>oZ4ci$�y���t4�NMm��I2G0$U��ʷ4����gvN<���4�E�k�Jy%m�nl��&���:�%��W�Z^
�!'uVսM�@��||�F���F��r�=��<;=sM��j�]��#ɨ4Q9�č,�9V��};EUc�2!DS������C���h���[}Z�aKK|�3��s�m�tԷ�����"})e������kF������x���V��|�oV�99D?�S�:�O�ū
 �E�DzE��9y� ����;p3c��!JN6dsa.�8�ȱ^|�Gz'P���_��+bg�:�΃�g�jm�KJ��y�TZ�K��q�/�-��� � s������h���c<��꽖��Q?*ЯdN�|o(�ݰ��/��7ܦV���t�w�������a�W6{o�@tb��rb��{��NCuzd�p|�qj�F{�	��#�C�7���~b��Z�PTf�j8R������!Eޣ�K�m�S�rW��M�|�?TW">�i�U�	ʽ��H�_`�!~�����*�|&��x.5nc����Z!��ړ{������6u�=%�ԆR����	�h��@��%0IG���q7j6�qn�Y��mE��Q�m���YIo�u�EKe���[V����t!��d]�������
�>)y���K3n-�hz�O�\{��
���1����E)���t���d`匎e�j���ŦǏ<|�w)�{��C��g��'����c����6+5{�HJ:~ˇ���&��eM=h��xp�j�ڵ4yM5��)�ڮvq��8	���м�ύ/K�i1�.\VZ�lq��:�Q�6�}�o�[N�zg��sˮ�h��Vt�iTـZ�O�@�r������I��6�] ��p���-�%$��8�tr�v�E-g�m�hGYO�QL��!$e�m������XS�b�Q%��踺��ͣģ�1K�W��%�{�S×��4/	ﳩ\� !���_��8�i.�x�"%�M�Jj�����,���w�E��܈Q~"W��sRR�n��2������Q�7Q���0�����
2�<&q�x�!?�z%�1���2��p�ۯ�d�L휖�9P�#Â*�)V���B�����گ�VB�<�z�V�2��O��%XU"�>�#�|$��}��bMQ���~@qv+���)Aۛ�oWx��u��;5�r,�Vw�@/9Se_�a�'0����@���g���g$�g�~	Y'��>�M��<��Y0sA��c��ͦ�l�����7�mʲ�:m��5i�~D�D5��֖�go6���<�qǥ�r�����것`.ԑ����X�R�Yhw���*��C����"�3�F8;�VQ�]�qdvn7��e�Y���孋
���������#/?h^�Q+J��Ezzn��W+����JO���2H/�a�,���!7��p,�:>s����=��H���*�*_��{=?���̑h��|�6�sic��y��SE�ÊS��S��D ��� �w�g�f�D�ƹU@��y�$���#s��]��0yS�k���^�Xd��͝CW���d8:�ڲ��{�&��W�8OV���_�Hވ���(!rsБT�a M��9�{~�~��9���5�:�ȿ�d�ap .F2��y�����	��� 
��~�GԭG�p��M�t�>����-��z�����d�����R�v���<���[��������D����ۯZ���ErC��1��Ĥ)0��[	ݡB��`OM>Ȭ�X��h�*�Zn`W�ۿ�I0�	K��������	#�,��Sy�ϟ7�wљj 4F8Dy]�K�����|Y��������z���������w	|0nk�S_���)�N�ǵ�]DS���^Tb�D�� i���=(���p�K���e���} ���M(Y-��sm>d����s@i�C�Rf��W�)ϩ��kd��]�$[Zj�^��ĆA�UGX�)!C,���99��FL�E	���%�n����V(�ꏴX�h.�.h!�}Y8'=�4"A�q�J�T
��59溚ث����K���y��]�ZK�����ppx?��sx�ԧ"��A�VvM�PX�W�_ܸ(��&~.��մh�NSO��+�z�)\;��-�Y��0�l��h����P�g�L��uY�6Cl�ks�A���cR�S�W������k���"�	�7ǅ[�!�>�I�
�]�������y�TY~[��%�Ur�IHJ^�jo�@G�?L��٩$δ��S⬶��R"ؿ��:��B�����+�,������-��n⽇C|�I�!��4�����h��pM�#���)�7Q�'N#+��DT�����uI.h�E&��W~��(�Hi��!Z�e{�"���
b�'�<��Dm�֗��vp]��)N�����r�m\��#�f��"ѯ�Jؖ��)}���D+������"��5@Do
F�`؁\g��E�D��B�NR�{
�#���(���f�b2!@ඥESr`y%���.��0I��Z�%D�F@���O��CA#��a�A�=96y��R�H{���u�V����T.W����k,�h�}"�I�����Er.k���/ژ�s�7��^�r:��X?P��UQ�����$�A��GU�z�	�����B NgL��FW�&�����|WcA+��5�vJ)(��a��8��7�JE��DR��-{[�p
x�*���Q����+�B)ėoaᓓ�Sz��ᴃ�Yh*7���!{M���3�z�x������#�����gX��1~tWl�#o?Qp ��R�vP�	VC.Fח�?�C��⭚�29Hz���q���͍EH��%B��^b����f�@�g<�魶u�˹�I�2�q7C0=���Xb�H��D]U�B�ģ�����e�Mg�4D�Z�:�g\b���=��SP��CW$���p�`#��MK������̭�K�Y�[�uݵ���O�h���{鍇�����|/a��0!�uWҀ�2ϯ�a�������~d��s ]c�ٿ�-vI?޶C���6T�=����{�X��d�U>�ܩ)	2�����V�p 4k�Vu�G���o��'����M0��r�ڃ�G�X�L��Xm�tu�z�a�Y� M�
���b��*��ڴ�zj�.Y����HSQ\����(�8�dQ{�Cpu��^�k��c�՝�e���"-F���7q�-��L��Q<��=�:n���$hY��P�������G�,�eZ{�ᯨ֜���.�)�[���+l��Q����q�'?UWf��3�i�'b�n�n�o_�D�8��	r�����t�^C:���/cƑdG?8�������~`�[������p|���)��
�R�������߁���s�3���l��F��{��=���DS���(I��}�EG�c~��s��u����0(�P�Щڳ�����Dpٸ	D[�7�S�I�*�����&�6����^��e�0�^<�����sV3�8��̋임hs�$� ,*;k�HQ5<1\�!5��Z�ү�Y�e���gt���YDArd�~�ǥ'/e����̈́�0����#4K�G�d��H+m��'*�e���j���M3h����I!�MCD���H.ͱ�} ��d���ҷ�bj��FV�\F�f��n��������h�Z��sĜX��a���F��>�Փ!�}�r����h�^�1��N�khl�oy�H�Z�f]o'�㑪�[��m�'��1��_�4ߛL  �I������-wH� n�!ږ29̧�SI<?�F}w��-ؾ�s����\Ëu^v��\�����&�h�f�naKh�^��m<r��r��:�:��h��۵��^[*�u���o�D�PFXY��:��;�u,�B~{
}�'�n�� W�UX�T�#T�D��M��1�E����«:�¸I��t�)	�"�;gi[݀ƞ�H5B?�A{,�nN +���d�G��C���u�&��>��_HM}�=�����(�j��_�ƶ2{-��b}�O/F�N�i?�Y;�|{�0k��1Õ9j���\8$U�va�ܣ0��e�ځ]QEw�8�1 �j0E��v5��d]׸q��IX���3��q�O(�fY4Np��HK�tɯ����0����K����B�e&����K٭s]������	��{��&gY+�����;>1�ʶ���2�O���<c���e�>�Q�mX��{;�M�r�zߴ��iʹ�w]l��6��:�Ա�1�)�#b��<�˒�r�Eჭ������Թ�J8D��r���^-�76 RQ�l������e
�ᰰЇ<�������!Rm.d���؞�Mb�)�М���<����Ma�A���A!C���q�tȩu���^�"΁]W^h��,�D��S���\b7�V�kwK����F�vQ&��tE�uv�@Ƅ��S(�`(p#�K�α���C<���=ǀ�K���a���B�O	r��5d�W�o|�h�ٝ�´��\���p�G�?=j����n�?�a�:֊KzV}��l�kl��~��ʽ��p�p+�����ʱ$z�&� O���
!��L�4A�HI�yh� k�cI)D���H� ?*��. !�Ɩn+��S��:]Gs���=��	:\Q��b�����&��F��=#v��������X�� d��w��;��3���3�>�(T`Z���V�*�X���PĀd���ܿ�S�y�~ǛNP��� �����3�ę��.�P�˩5�Z.g�fL��L�KPͪ�����؋\�<-'Nt��\���VԚ!i��Im*�! ��m�=/­�bZF@�3�=擀�[9zD���(E��Z�3q�Ç�U�v
v�H=����;K��.��,�o)&G���	�q�tx�I�R�����#1��q�w�!��7�Yy���K�W�Hv�X5YS�� ��T��e�,�뻸�BH��y��Z,G~����_t5v�s���s���}�P�EZ��W�h�����
p����qF5] �Z#f�s	}����{l!*0�S􏝆G-�r~�ط�2�K�L�(=��>/�g��*ǁd��:+�9�B0Ä�Ex��2k�`"^/��N�I��&�.�1/�T�I�]4'��ʱ��1����I#{�Fu��J7��M#(�RR���%G�|b��!����N�
��7����fm����2��
���U��Ǥj��H��S(؀ڰ�Zq϶M#�w��|�Tkn���X���	� �Y?�M�?K](���sbQ����� �Z��$�T/���k	U�Z���;��K2�i�[�M�?��E�'8��`�D?kN "k���^�0����	�Q�&��:�-��c}����v�'O��5�	���f��:m(�f �W�8�Z��y��(l��d)\��qɰ���*<R��zw��9qT�H$�c�{+��ZC߰aF-b@]ۮ�I�O�X9���<.t���c2X��t����F �j��w�k�r{b#�l�=+,����'�����֍q�G�_3��&z��
�/<m��I�1N�E oY`���s%�Ϩ��1}ق��V9?���D$�6F��Z6�i�����s�./l�5��U��gާrЄ�ɠX�`b������-e�U�1�K�y��9aFw*�m]bC���S���}�����]��9��$�9F��B��9���p��"]]	�N�KR��]5[��&�/=6��Pq�"�5R!�;��� �ú�Y�YZ}��ߤ�oK��hx=b�o{/ty,kT_�ݻ$�#�q(RY�z�ˣ����^�GF�.z ��NyjguUU��N�Wn��HD�3�ݱ陟���Yf�cek ��o�����PR�:1�a�2�g-J��]sG���K[�^8���2���)FP8��[��dv��׎$�9��4!{"����r��f$����108#��B��$��e���3�r�u��0H�Ң��*���މ���u*��/��9�S����N������d�x
VUȀxq����Y�`Y�M�
.�LJ��ۄ�<�`�z��̗+[�RM}@h"G�$�!���1��tFv1�=	��镂���L��j�GB�TQ��B�����j��yn��0ōݝþ=��c^�I�_�&��,b��"}-���¯�b�U�;e�M��d5�'K�Sk\�����l��i��lK�T|A�L_ш�
v�\�FH^%��q�t��=��7ENCհ`��k,��ك���ZkS||{١��Q W�)���#�8~��b�jj�	� �f'PF�E���b�(+�w�8�$/v�{.�o���D��DDu:�4�x�؇�0x�x�.��ȦI�AN8�?H�Hň����R���嘠w�isE#g�CB�,,ڌ3�j���s�� p�-č�Qj�����_j�[A��	"�E�;#�y�Iӵ�h�Pu�����������ӽ]�&U�550�FQb�l��+a�����kd(��k�܇(����7)�N-�� �Pw�*2���a�;��	��C�ه���{Y�4��_~�ƨ��~��p�j
�[��w\f�mB=�>W�-�];�u�^%	[% �U���T�ۥP��&&Xo:��Yގ���ƎU��r�Q*vd�'.y���qa�.�C�>��w#M��s��	woX~�;O���g2����y��Q%�������ۄ�b'<-���@���R��r��e����3|�}����Z8���u ���<�^�It�c*93ڮ$�&
[4wC�ãkF��w�2��N0��ө���:�4�2�uc�t�B�ƫ2hVM55$�������)�H I���j�6�O����yi؛���?*+�{��\��[l�qQ���Ë����ɜ�Tta�9lj�Ś�h�"'<fYW�Xu�Z?׃*�5��ˣ;�� 8�ܦ`��*��N�K���������o.LXx�x�����.FX������>Η7$|ێNT%D-����6��5՝�!��cU�WS�c��|}v2ڥ��q��NTY/ױ2*�YȞV�RW��6��۰�ţZ_k�'C�$�]7<SrB���WZ`�p�N,��pߛ�������� E�z��#����!@�������߬��A���c�����Vq��~�!�m�?��S䡱e&��s�a&�D
����.�(� dLA��Zp�����e"+�	��p�++�=9TG����l�B�"ӓ%1_�=:���6wc,~��ǉT�d.�@�+I�py����](b�h }�����	����/��樏����ϧpi-����y���j����"���Q9+E��d)�6�	��'����π+���H#�4���"N0#3�s,��_�M?����5�����	>���;�Y�q8"�%��jl�����iˬ9��l%�����%�q��
M��C�o�g�%N��/!�t�=����l4=�_�J��~�xB�H���1qnL%� Q�9��,��?��;�ꩴu�aL�,�4	�� �^?ji�x���U��pQ���%Yx�X�ɘ��ҙ]��-��j�Ј	���%�T���B~�Z
>}x��.��8l���]�Gi�_�ē��ᯭ"�3a��I����r�����vD��BrU��\�3�va�� 3�M��UX�����HԬ�{��#����O�x	������q�g6#Z�z���yG����z�;(���r��CE��>8)��ͺ���"ْ˹5��h�E�>�c-�i�(��Q�tkQ�76�#Td2W7nn�����	/�| Vx�Sv�c@�ͼ��t��p�����~�"��'�X�4v�"�9�+s���PL� 6���W�p�p�؍�,����H8J;�~b��8b�������Vøk�|atx��=�O|�w  ���VE���6�>e|E���3��d��JWt����A|Yn�uvrǤw��>���^�h?)�b��j�W�U�y�į���;�u�L�31iı�f���n;��璳���#�6�N�,��%�S	!�_�+��f!�D�Q=:ńsЬ��0G�\�8����a��n�c�0=�T�x�T�W]o	�!:�gFX�{K��+��.w�����8Q����<�(����X�x�ʈ��}�Y:�l��%��Q=�x��3;u`6_�<��l�☴@��O#�KLp��K��O�_�A^(��p�ʁ*��a�uX�j��M�Z��خ����8am-H��Z�߰h��-��̱?�b�:xV�e���B���]H�6��CF��w_�v�NL��=�	lR�>��8�[��Ŕ[�p����ٚշ6��>͙j��.u���a?�+zW.�)ȅ�/����|��p�L~d�}(ל n�����-rw��
sD��*�]┬��@Ѣ��	<e��u�� �|�P��	���[y�"f3sr�����qU)4eHS�	J$��lI��̿�H���9���X���ԈS�H��I��,7���J�5c�t��8 �Bu'��ـ�D'��8pw�ވ���B�v���W~hRӌ�ђ��x�P�F�DO�֪�����P�֑+ovuD/�����#������/�$j�a�'(R�����ց�{��|�������|x>�`k�
p8y~� �{�_g��ˊʬ`¶{}^l�A�������!���1�,����� �e��0yZ3ڞ��������rh�� ����=���&�i�����u�h�@ף���Sr�+�<���*6�_ B5���<�d>���,��[�������Y�ɵ�#�_���T
���T�=�CH�"jU�6�vl�eN6_k鏬45�[b�Ɇ���+DIr���h!��=m-J���B���͜Fa��&#�C_"Ů ��t�خ��y��D���K<�٢/mH0�ǥP�ᬅ{�i�B��]�?�n�
�����
V���c��F�x����8���"]��4֩Ķ�f*�t�~!��U}���I��Ȋ���5�f��'d��+�sK*���<�c�u�;LS(S@h9�B�&�G\3`?9�&�S ŨL�l(7%PV�Ͱ����s�ҡ���B�M���W�¸��{]W�"f�ɜMX&^������F��See��?�����үd�tm�Z ��O�b�|��|�mz���e�ǥ!�amW+خn�)��סǉ���;6 #���2R����ȉ8z�w�}a9�]�,A�2��>c���)@�&W��U��.����