// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jpAh14dHRopv0nKiITfYDBPo+fX5dNSQuiAG7Kn9IMFvncSjhdczsfUTHaI4BeX0
O+W5Bp74ELUzbq+Oh4HlansC26MOuJnBe6kPZ/TeEdrivtFo8FsBf3+xrOu3Xz08
IzINMs8QTB894s09YsjpTPf34GKj24Dg8BZ4nACimmw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12784)
lzDPngM0Td6hiu8fNOi9FpXQj4eYqnOzhyNESUbn7MT8wYaQuz57XHoM8bO6mWrR
ulrY74L03rJ5Ku38UI/GXVM1hfKvm7m/dnPKpfUqPz1v1639k7kEuK7MX0uP6hHP
o8PCxYd9YroayO2NeLO1Ak2hhmIQ5o/KTiZmqpVOGNcwhEi9th/xI2nvg8/LV0pO
XgFv2fnaf3MLtgvsE22WLmNIlu56j3LAEQqDfTNmawJmVZqVBiOD+LpjmFS43kix
PJu5mWTl3B3+MR1uhP8kxuYrYZc365uKWr79xkH1xlFbGHf68x5L9enZQ/fOrc+r
UMvXGM1sGOQeB9w+bvOCpRKIA9Jg2YQuH66p/aHOJdJdcGpQsguNTgsZjSut/aUT
xuRM5dcBSrxZgHKmYxlCWAbhpjHptc7I7X2cftFuXiC6Jv9WkowWfWuUhtJ1k3lR
VzU1Bae4axfAqsCUfo8qqH6vmOtwVJFSB1hR/JtbMDgzAjUBcAT2FyLrEhQmWrdW
WQ5fNo1QRzwBHO4GF+OrVqqImodY5iHF12HcIaKZhOTHL0z0S9wpkvWivv7rBGVn
HIIKOpgK8VK6pFE1ZhIJzclw5QzIsW2zSJT9uWVs4QLGI5e3iW/ZKcHNDjzZKN5t
W14tp1YfvJfhT7RWwHdO/64W8RjKFyz/lN/xXXAT1Lma5STrAAjuXP9aALflOKMK
kknY4x8Oi19qaiMk+pTytQJrluDIQgVl749g3IB6NKhzPfUCZ/2KaRRXG0RPW/fH
aXKISqRg73qleoaLXv380EsBeHDIFGpaEp2L/Gvp5xm3HIwII3aSalHlbug9RJIB
yE5pV5HOk9El50j3RjYfXVDIzDql+FplCmul5I+RfnagEVSuCtgfFGTd9+xBjcP2
yG5umkUwxyNZrUU9CiCd0J4KC0Za+2M3jvrsRsQ1uk1bVo3HC4h5fm4UVw8D3/yj
lLlkMJL39rI8qKtsHt/wE2pvf/61Dyu4YbaS1S7KIico1NwEJqVsAGK0Dma0vkEz
2bG33vRickFnHUkUYIAOFNWFPy3xMmYCh0V+kvpgm9eZlimmSRpxiRscJqmTNes2
/dxNHP0dpNRTZsK6y0YO4w4v0SbrgF52DTv/VUms5rLETjE0c65AonEMWg4XlotU
becw/V5Q0cHIVH/nO513qVMb/q4v45qxcLnHcVJgt+kLXjlyaPz0iucGRebxO5xb
WbLYzqJFSAoSTSSW61IpnhqlR/0TJ+D8GyyMZ0mL9szEJw0cG/uwa6v2l/OEYQQ1
Ypl82OfWdnNjha3lMn7KwkIsv+RDUWnSaqanXaL9ViwO0usjFJl/dLW/vKfsNW3j
DN601elJhs/WWtEfuMPu1ibjNfIC5p/s/CD5vPpy3t1jkok4RKSVV5p3gqE40YWh
u2J9lvCIDbkaQjcJXJPUP1We8mU77b0TvGk6CA/oepu9HVGDvkWyTnWVCi41eTSM
u8y00DG9b1ZU47Fi46ACS7HY4ZEXV6pxWyGPl5oWdz5kJminzr2w8M2MxCAbitmn
M/GHKbUIPZwRS5FYaPKy36HYRZkdud9YuGPH6J7GcNEcDIGnXJhuWS4p3k1Tfsb4
JqFl+MjIR/0lO5qSeGlj6wzejlThaDP6V33xdYpSht1xCbuzozyaXfYEj49WA+WJ
I2cbH5dzHB2QzK17YeljfEGcGeKOIgi5hYMjoqHpJdrAVsCt8VnSR8ctJa1JeuNr
MD1Wvt6Kom99U7G2ZRM6QqaTm7a4+W4ClHdJAzRMfXp6e44nKKgUx78xJrDJt+b7
7QnIsDWS/B/2AoHJmc0WtjsDjZ0370yzYucHsItoVn4gZufvoWrLBFbwxM4pCkk4
JEjSolfH9mGk/nzhMfdeCUjXVqfqURm/QGUNTQKFAZ4XRVFqEs1KkBRd1ZFf4kzx
0xdxUE+VkEF1SLa3jfkQZSM7IZr3uAElrEb1528DF72VfM1KPsdVUQp5MNloopFJ
kjUQv1LD0TL7SI3/Qd9RV/9QOECAfcomxjpOmCcqiVeDOrJ73Q6bjnDFWIqYvSi6
/JOesZoGLOy0JXufYYnsBeAnz8dcUR3rFkY2PlGwjTpmbDHTypFIipJ0AG4ts6ig
NBy0kdsnVejwcmz3y8XK0YdrpbR70CWlE74UhPiqUzOl/bnN1cdgEE5XOeK/t/Ht
nCxdYmgtTjIOKKC2AYwG6pdtgJaLWZROiT9V6/OJ6MR2orluqKsb3C5JAMzhhsIJ
RbQfhbywlBjm2mjrHbkPF6yVWTfIenmTpAFSnT0Sb3FJofEhjqxatzboMZJFuQg2
3ZIXI3vYrSFpvfkyRnNntEipAVhaaq/kNIVBByb0pBdGZ1DT3ZXsZOCMMDOg6B5M
tFzDSIuWKcL5OEFG1e6UtQcQP8DQpvWVzQrzcpzPfaevXKlO2/Hign6JaNNXlGBm
K2aB2YY32ARjC9qb5hWlr2DgfKcyequ1E53HGZyD8Dqdavod7OMNUv/+ew4uE0RO
7f94mK9k/a6J3efirJvMRiPP+UZfF6M8v/69qvqydFh+QDvUozYi/MaOO6liyB2I
T/Y5Nlb/uNAGtZZj6Jpa0FH9UcWCccJxcnblUv5KdPnpmVMj5+H3QQWv2nw9H7eb
WpqmXc9urcmm94j2yi3+Eh4s4v9XpYusx30Wz0i/SQJ4UFty4TPJMPejaTb3ibFj
VvyVU5kaavFAwOld8sEcwS4H+c9LG4tpC10EFtGI9C9a07AEpZ7lq3YDOUtVbpzr
AHSDcZhGVg2sQgfTy+vljAEGk9mXv6sMOKe6+V2NtbMfjImHbUESk9rDxb3r29r4
1XOf0X3bY1OVsHzXFvMHit8Ue9j0sq6+nMqlQHKf6jSW+5qs5dtLMttwQeZXL4z3
yx5ZLJY0InfDzgk+mxXtaaAawRwnlKqxmNYO39zkNFhqvIHhB8BTdwtx+YfLFsD4
Dasfn5ziFI0emMJfoRv8d3nuRsysVOWfyqrfZ2uv4syUZGMq1CasrKBIaA5I+Y64
n00QzVzxKtlqTBtP8QqPH61s4ZzOeb+wVcdtngFno09XhG9h67KFcbeKuJwwvbex
VupDvdBcfiK6Sw5nX5smLJz4ffioCqUdWAERRkp8iv7SAq0A5WV7EXhZbIaTkK76
fZf24fgDlZnuHW2aV8HIIvpgv3nkoBge/NctYekCqIaTxbfj7RM4l9clzdKsHF84
S44LGxYbUJyxvyI5/YId9cl0VoUlrsHq/aFVbkvO01Q0R5P37mEyzoLBO2VKbWWi
VQANriXOYY3MKQllAIKu9WTeHyBssmBv82yKwQaaQ7DIZwyb5O8TeR0qbHVGwhqe
tBd7w8vR3wuOVkScfLx6vzJakRPeo35jw8sWNoIYYd2jAMKGbN/etlpbzT7+VI7h
AlIgSVUk7Q1fHxhD6/cN1DnCtxSeJBIaFJLrPbfwLjd4JiqFY1qT8lKJ6KTb3YGE
KxLjadtrEZuRDgtETIzomy88/xr9uB8nmR0cJ4I9WQDxLs/3pMjPvESsiiZmAyLr
dEelpyANsJfaoAvlU2k53ZVUPEM9Tnv8RwIlVdBdoBQ/tYCTDZMX00bH7Qnz84RN
9mTmhkNTjmXHVPaDPTiMWeQp5cQq6MlWnaYrzpR4lfWn9CKw+bElYf8xAZBbJXYf
mA0ImFhDen0YkNccwVM93gR/94DOTsijmeo6NwW1uzoFrpIREL1p+kzjulkpaa2X
YLAxMIBbIZ/7/1T1fknKA8W2cXpNUDseogAdjxcGIGGSeUMRX4RTM5isGbpPTglf
VxYsk4uYteVdZoAAwpQFyui4HM3D+4eHyfA40RloQcseaJONa3dy5PYfZjYodrUQ
9Uft+oQxkg0HhrfKk2zUR0bGxsX6NSr4cqlgY7h/yln3M1FG6kwkkbPL0slG4vZb
UzVwo86wdmyWQrIVyvyrOYsM5LxL0u2qPT5y0b0PRqsI2XfMJVtPGlPBAgTimyw6
j6vYXmbeoWpZdAEI4mnLKGM9ZIsv6ugg1haZpYe4Df4U2VXphxQDjvzRvlDgpJPm
dMR9uLcQeToHtu9Rs2iJC535/HawL/WgTxOB7R9pgMTfvkZb6JB5HAssjxPnRaBI
Krc/7ls8hybLqLyw4hclVEJclePQ4YFnU4vo3Bu3fV7ZSS+35eDZX5N3uVsZdPdF
9SIikWj8V3/Waj5OqNpLmnRQWMaEfVFKdeDv3rYRdxZV03MgQuFGPi+DPkY5IeBv
A4yB3nufF7P1nOJRTMfTn1FFrAxbmT6362FlNmwMm5QmnmDyFBeej85SwoLaIM19
qwQLzSRNC/RnesRY24olVC+7CzFG1EDy0Z8orhZxH04lBntLglarOk04n3zSRU5d
WdxJGYODxVyCoP//+1mFR0PpKFuuOmqEEg+kDY6hgsHcSrlrX2du4iAYdDxvCWp7
/omDqAuOD+Y9zIwjuD7+maRYmKvbH9/ZfnBooRZfnZHA1KOGlGVGrE3v5dTm9NB8
lZWT44Jbx1hUcmZSyVG+cY9+mSWfi7CfchQSfNHoCIwjrZ/1Z3PEFollyCNFwH6S
fGlNWKnBwH6yYTC/CS4CWfsx9e2JfOaIEsUqd9DQDrOTvCgu/Fq7zd8bKxZnBl64
rnCdwsQ6GExF+b6n5XCPHVx3KD9ciemidd+9s1hRkwZMoAuh1pWBYp7cm6KAd2su
2Nzqfxu3FtSviTMRl99T2u6uSHu3132hfJP2uy1dJIMGO9gI1Y8SXVpWGy6Sfa1n
igUzPgczDpMDOspiMdqL9oKZQtXEw0UoTojujlqYYNdNyRUO3fQ1nH6yvhePPsNt
kUQFqgdst50HsGkx17pi8MRYBGImoJP35K7WzSE2EPwF+eJ/8hUzxnXeakSF0F8W
dTncNwOUu7wrB9b5oGp9z8usm+uhBglwYRYg0J0yFPZBvlF9jxZxS3jvmjXufb6y
vnW85edoBgKE71s9hao4xzLVIpk1NR5vlIb/lbHWk1ItrHFQclCRwEeNsqUD9UhZ
2/CYF6FPmvzZ9bqBnR3yCYeI/eXghtXnwh4H94OHDqC6QwabuN21lKTFtrudeSLx
Rgfiy9doKB9A55PBCjS5Gl7xTodw44BxG5GiE0x5JJxbUmLxNoq83evHzow6giIj
OeFupoZBtDgTeH1kmwQbzdbWIar9CJTNjG067JEdQ4XuKJDqqjOZNk26eFKEcgcB
ZD20ZTzU3gW+mVtBzd9sKbt/d4Z5hK1zpw8GVI7R5eRrsLica1DNS39S+NrWspxp
uRJuHhYoSCMJZvxTH0EdRuqrBHhhL0ziz8VLuImomCaicZloSNGdafNVBAy/kU2z
abOJ7DuDEHvKZPRdFiQZvv7KImW8QUJaiHf/6Xai233EKkCdEhAs8L1mpl/zxS3T
sapwLACwtFzintsNqZeEKi8CDZPlM8bG/eOMFNiFqdV/oS37pUikF/SBeodgf6Wb
luX6jRB42WtoHpoISpO4HmEvCg43XrmuW/iMZLgc3hWfDoa+cGax5RQFt7vFeAqx
IzS+U5EeUDjo9YOpF6X2exNj3ezg65ZHLrqIyEjORRCpkCSLhVHXKs9M7287HsOG
umiu2sjMbcWP7qQFUKphw0zVw4BO5xj4XuxvWRdO1Udsje5gxHgpf5hpJdslEX/s
45rE5oD3At1Q5hBd9kbl5XaEkgXJrsF+pPdTEaRdDHokIagyP0yh66hGFZQuHD4M
VYd+JWbdhoK27yI0j8ybkgxCAaKZ2hHUZ304Ac/YPbVoZdH7dd/YQY9+EeDqip0G
3oon6CT91jm2cMtSK0WjDpEa6WlysFEZjzmsNIZyjRJnzKQB4OC/aZpkSp5g27Tz
miCFt3J43/msqH8ZzwzWWHMhGsZr8TaglY0mo4eyRzFZTXXqs7iLn7z2+043n4c3
DCKN6FvNnulR3prV4k8Rurelg4R6vFG/gyiQcz2mUGUbWWjCGz/MICEYKlwwlN9r
RqTDMeYfKNAXalh/cbnTiCq10PgkTT6UBjnNcqvbV0GxNEl6bmBIITIYzd0RvAD0
O+7WXkLBtNs4LGAFSVrfsFVcu1EGk8Img5hD6nEWZhx9gYCFoSwWlWM7RFJ2oJrK
DvvW9CnqcJcSYSBBaL2VMS7dv/+DUsxr39duI7/4jTm/LjbiatX1zL/TeH+prFMd
p27er+Rk+cnwkNNseXH7wiTVlhM9LouG68EHUfcI8WL9xnF5OZmFgp3qUEG6JMNg
7UZeRO0bP19gkzUFZSKawmJidxqI/P/01v/d9aebbRtX6tL3mFtbK6yHNvd92cbc
n9B7FNkao25mAxSorwz0KPBHuQzAcKIRzTcs2ptsbww8X5kRECB6QYWIX/OnM5+S
fh3xbOGhwuYmIioIOVnh9p6yEJELskgYko/vp3mZEuKU8lvUN4WYV2rTU6VIFCRn
AOKoR4LfwXYbZwPQBJdydm3r19wKN5egj4V37I7UZtoe2XT5mqhpi6VdJizSbDa3
K7pmwu0bLO+8qHsvZVX8KE3iCY06lAQhb73VaM/p55Xm8sKdpF735dzGnHTwhXOW
mlt9lCEOgXoFTMkkdwcNSMu6GDGloxb7sh+LcOsE/rorJCBUecenouBa+qu8UoyH
zAf8ADiEoTo8uTOaM3DyqOp8lrea0NJWEXpWt5MtBVrQKIWT6+2f1YQ1bgoYOHWf
o5CsEG61Yby/1ISn2iU8LweCcLK9Vu8iPMyX5ZfP2DoYvavza47J26DPvRxaNGqS
h771ZV6DymdWElI2Jae38XoKPr9XUGKnHBhQ0EVF+1xf8a/DEcyBh/gysUZLtO8T
JCVdmpV0WSx+uFIFYNGaJSYy+4pYjshMYNVAEs2S62fY3Ne1rEg2gaeJXahCboyD
4KkSTaeWz5+p67VpSH7BKsYhrwZWRyrjPYkzi2pfo6N7BaepNyVFZ8XNEEUHgc/U
X8E4+QCE1yCSdot17isu/9UEStyeb7fPXHQoOeLz85t5dIvF2jcb8gKu5hsjVDi6
rOyS3SfIFCUtvoTmCwhiNG/V1hxBvCiuFTZGUP6Ap6o2RJMH9+lp1h8V4wV0Dj4p
ZS8BGBObvkmYIKFLbHrwgBJiAZtpBDFedXHHNPK2LLxf+LZ2Cm9qEyw6xxUdqSRe
b3TWvrpxthZyZ8YIb0Nk/tRcdyEFe4Pzga42ZMgoxgSATa7LwyVHPkMU+IuTdtFV
coIwgh9Bs4/3R2Ry4PEHTXYD2TNZcmLI1AfyEjzJNf+5URZeCRZZSZlw6NjBQWXW
/qgSPSNuWUEKhlew17vVe1LbHtIZcXMELBpLUzGn10y+u+wAsXvx4LDHZMQSG+P/
GQt7PbciDfCDrhqohDSMMVyxxN8/DzmqY15bjHyNzZ6YCKUX1xYnIubLOndYFJUK
cCKDKdobaagbXI594nT4iSWAXKjQrXAmYCsHVxEW9I4Ot5/Wc7tRZGtdND7dok8t
i7bU+GlkETeI27/WcUpfQ5CYOybtKxv+DB2K38ZBfkauqixjEnhb35XNmqDrQ7Z7
vI8AhQUeJAqnEOR/ECmaVzFP3hrQVed7yXhkMoq33cleCIjvmRlyfrDCpP7Uw1gH
1xnRU9AcVhMCRqNtLDh2qIABpihSci7k2+xZ/pSKjQScVjOtC8IO0zUwNdIjlcat
A92UyYhoxHt25/lLx6kjR7mPEs7FEId/+ejEMF80OVoOGnuYD18nTBHJt8Le3+1p
RpEdzqqle+LufdJ5d55umUozXvW6II6a0H2HQ0trFx6Gh/rivXtSopEIRXIRVjs+
kGGh71Z7SRpBMbhAAdVGe9vVfVPoo8OrxWQJ1akbDxNs5lKWWCyFrDEqJvX2I9s9
dfEiXSK1QeUPPTdH6ZKhNR3Fvm5ZWabBMdufLiA+CyekuqFCv3UciqBKrmTp+rjh
VGAmIwOCl5choUz5AyHz4lwdic57JmPq8I6sPCTPiirhKkBkUjY9Y5eA7h+q1CEl
4ziqJb4zvuVGnhCDNZ6E/mss2SYlCHpPNjbzDTW6+MixuTtaxtfzs91zqeLH6his
bYyvU9Abzrp8xYN9pCpLWi9+M4w9HeYmTL1dyze0DzJr2BYyjnOgTv/3Sq3BGVax
6UGY+FTPVUupkPgP/rYftiX+OFFk9bTqiDhWbiddxpeV66dwCxaTUibCIaSKYnWr
mFuhISY1/+ljUi05I22JAc1DFZmSVmiYN/Hlzx64nM0L2IOOncfKufIm2LaibKqT
rEcHAdJdABwKZk1snOS9In1Fe8OxrZt9InGmqboFMrt8hu16M0l6OJbL3LrN1kLH
DrovzOmAiaueH7zWq+uytIbWvNVeMXAcADpVFFEkCHrb2PGCJ9mcN0AyQrWCQkYA
9qZunBgBjIQch7IDNhzLU4rZrUwEq2ym6/pWmtx+9mD52nnMfzJm2xW90VBDtJc3
sQkzpHSxPtYQfK4wkRUF5TbxsKno4gswAL6Y3gFORuQ3PxR4maS3S5ayCidlrABa
PeG2yLe22wCB/RTYzbnjJzmXiU3ITYiQX8fZ19Zn2jYoXqWd6+XynnDXja4Vpi1D
/SSsn21lgg7j6GoOw4LDufxuy9zeZPOHGh4NaKn/RRQTzKThID89oMXT6AaQY1tI
Osgszqd3SIq8UQQp7MP6r0jfaf/jE8VwMO/OK+VH4qsMgdGqb8AFNCz6X+eY59B6
w7+rzUXY1cTSsXB79ltVv36+2DKM5d2L69S5k+t6Zvb16KIvmfSyjqF2bkENEMjk
akMfW5Y+nDuCSEgRMRQ8rc5M3n2Ta6n1GO6pOVvbznNe9xnH6/+OTZXyqLU570hm
RqQMZHDA/l1o50ZfZqL/xi+oHaFJBaEq3LD0roiiaWKF+fMRtO/H+7u7kGE8Irdy
biYimZrazMvfqkaOw8sl5/sVLrHR8utW9vJpWLdTogjLVXeaWsMLz35AjIqYRTkN
gOngmVZAcV7FoaINCsRgVux9WRV/iEjC+pBXbBraRhJhz9HWxoSO80ctJs6OTy/+
GVcgiOPsqdOYvoXxcX7FfiGic9Zc2iL8E6CF3ckPAaTx5PMBHlbw86TVaUs9/ZqS
JrP0Upcx+AqibrxeO3K6mgPA3n0rxas3+7hGUroVVT1lUuPsvOPEe/IcTLCDzgiL
niYK8ntBECuDSgyDneMbgzouE42G3vmDCEx17Q93Aashh/HOxxY4rQt5QeiKGqUS
CcO3uOE+rgO1Ma5Cg0UKsNpTNrWoLjI1xMFh/zgiHYw8Ht9m6VFi8hqspkKPAStg
+sHRm8L+IObenQZzkVtvwwcuz08bwL9eNicLmk72RPd79W1EerO1zlul3m8TN5xQ
pbeIuifD7zQbIV5pZaUCx4+dDWiTV+hYItWEkMmmnS2V9Qs7IyjUQ6JYphcFdINq
p6/iROQA+l+vFK44+ytDJANbasHEfyrnIlzvEEzz5ixB4jGGinzPt6g1Q5xCTElu
2M2PY65FNj+iRmtGWhD1oVWGTfqU0SNHEw9PxUE/6OEB3w3i1T47w9QQeLbQZy2n
gitzhZnvxbA+7r+jOBqoxsSqNELkKY2mciVM6VE1u6g0w/tGwkM5H+czgKm5gW1J
8AOr8K1nHvLjfU6ktgAzN/NRl13WH3qCsGk+qWPrbcUTMWJfgZx3NWJshuooQJsm
6JMdVYpzbX0XDdnBwwsS4E0HVUFB4ksojdEwNOaW2d6xpeyfVnFRJ76ZzcdRj6iw
1BMf3j5TkIRtQSZZnB+BmQiplFxh6ILitSw1qUPcvm6ZAcLphR12vXhJSeO5ys70
4swag2dzJedZ1LzXBcvBmEQRShNLodi3LDhgZedxflV52ZZmN53KwKjV3BRGJGyp
8dAuwLVIabO7IA6w6/FzZo8VhuDgstlBAEIzlP5MmjW6rOm07Ca6gT9aWAxzsQBV
A0AqVtxc97V6+Nr0V2LOeEfMzWTZLsRYFnwXY464WwwVCwuG1mJ+uNlOeu0Y+hGv
Arj/EGpWdvoNGygh5O6Oue3hItdlV3QuZ70cEoko7EpyPL5d5283yq0AQm15YdoK
YVbSOxkOEs40UBkZaDY7il9IvtkqmMogEoZJQSUoeE+VHHgpMxQ3meRM4bjhTUuc
AykGthPH/b2QN/QqgzN5OUKREUCzwimN5NzjZjZDKrkAONqQRQKrOa7vl0ErF+0p
+S6u4LRfCv6ABezweCMb28TNiqBEM1AP8vNtdZGU8aNt8ztBaEEQ9gboLceAti5w
EVAdpJGEfvPdWcMlM7H9VdR8lnFS6anv7dHGqxv0cPUCsiDHpwIRDEkRGX6UM5/S
O9Ln03IpHK+cq15Pqqd0CrR7QOX+ZsyK+P/R1o8SFIYxhUN9rtkksHvLCSK/yWrz
XShMwn6IPKM0UAAtvOMY49Ek9yarj96JZqCH8eQC13mO1ryC24u8zuY9oPMP2i02
l0fVV+1akTCXPbiefcriPVmFmeex1O5ntPnmCRCJzJIjLsYIr5qWeIoKjTQ8IUhj
NfmWsnypsXyRnWTppxw4GC+5U2QHdMTHpUIDnlDEF3CYOY6Ap0U1ST+W9N11Ixyr
8Vsn9XJh/MyJd8MpJHca1F+fjM1eK9hKX1y7RNggDBf/ay9WvqilDPgZgqkz9+Zs
7yRxWx1wDzXyFXtjMXsvE2czjGVzTvxOqkjf4LygLp5ghp6B8jntAskhUg4QT9rK
SSClsbj7/yEmC/KXinMZ3Mf4RjfEwrEDl7fKRgsapqZV6GcssYHaAFZWF5ZcxqBg
E3N6A6AYrg0+CdH/AZi/k4qdjXIlVxfhsYJbDGtFmO0wmUOSgRVUK+SBrVThaTK2
Uj8DIUV8uVtvLgklCb6NQjMraZzYZ/TAmSXF2nqbN4lVFmtOICDMj1HYRA3U5umR
clk607xgMQz3GDQ2QDK0gyfauWzWXQ65ZXsznk8rUquazFn5g6BAfKnNyVtY28rt
iJstCgmREr98jnDt0E4NWbecAi7uifUsS3f751aDhQAE+Lh3LT52ZCj9uNxpPrlU
RoqonBEppfG1Ui/cPqTNGDs7D7RKhkEv8BjXM4XFF/alUlnuBTycSxsnlA1O+vuZ
l+Xeng0jyQkte2zgNrNL9NMO+If0cd6XPbKM7a4ucgNe3X6U1g735DbrAakJ8TEA
KnSwiaIWEYT5LjqBHUpZ88diLnq3sqhVF9vkIB7eB3R8YIqMmoWoAt3G/p0dfmrV
4qJWr6Vx7bZBq2AeaI91eRoP2suh9FKj9zeFBwyYahDxlh1aBxhYPuHUg2F2eS11
NBFwF73JnEkE/mgUFPNdObiB5cQwmKfoE7yvJf6HpjqmFsc5zKh0c++YO7x7ArCj
Y7yDGlEfGAq+hkFZi7Nrtmp8EBfzIxIQtV4Z3fbGaBa+VTJ07KiLy+wmPAwZ58Dr
dX6DmEo9Gtl82tieYgemiJFANKmbPn+Axiyjc1NFY8M4/K8ROochjuDtuTlYuPG3
sVtQQk/uaPDCr2DESFAmAhCnpkM/QT8NauxYo16Uv6DuGeRH0ryzzzz2cfJOjC06
Nil/t4BBhE7kYsoQwngGTLPF8i3sDNlIMMvobX8AxSYcwe01p2XYktOy2vWlCfX8
1fZZpOMhUFOunEfWAlaDbRsfVpOq7uanMNR50eM+QuIu8zvwwxBAb35pYJPPWVgk
WP9COhip+rkDvHvw5d+0haK6dQwViUeq9E5CSaZjvKbGk3374pV6jDrIQdaIzRK3
pEAeuJu3wRZqhjJ/0IQmbgPDGBy1PwLGUqJG8DKDXk/0Bsn/rLv7Ft8iU7Af/CGN
w+hLRKWkDypNNL5RhhcdkbcCNNhVjoO6sbrx59t0183ItTX+rB5SYt4nrAB7uSqz
AgfrqnDGBeJf+CsLM7T68ZsoS8to1CMAbu34by3/to7t+bn+2UatsesqZE8z1QeU
qSB2Fg6BFDHmip2SwDD9a5PqraAmI7lAWkKYRVo05RohscolDp0oaFE8dW7Rfzh5
umlMJuJLJpAp0y+QSF6hSlS30UjZzAVOUjZz/kkdha3bNEgfGy+S/61+pp0Cc8L8
yGL85wLUDVftT298hzkjGTBNwRnvyXgOTPaR7kJoD0rvjlci/ONORQGNYhCSaZ+n
IzamQKLT5skgkKEZkY70vf/55FDwlBCg/b9KFaPiKkSSnJ87WFZusR6MTFJnNAzj
BRd+wnuYNgMbrVkPA2a2APPsAYaT/G1LgofTsbxwXv82lM4egge4iGOdPLk/qlXn
HOniG549gFtCrDxa/SxPUzWxjBgWE1WmbAAB+2qVOaRFGqE45cLq1fP/UNxBEQRd
OmeQho7FL4aAcO6BbF00B/BpdB5MgFfuZttgWBY9niyGaGdAUmu/PiOYWvUX2Vhd
2Oa/ufVT3GEVej/lT92a43Ly0Vsm+UioRhbLfk0uWn/dY5fOQ3RzBPATWCMjFGQi
LJYmlsatPPG+ILCCFv+hB85+1uh4xG8xzADvGu4Di40NvIcjJZ8oxurUDxmU9WVL
d/lH4xHjGAmG80xJaN6Yh8eXxk2TYFm7nopOTR7ArI8q9F/n2n7yNmOLjv+zajtb
iqhZyYKjOVXRFptH6kDEpZgiEAjn58TLoTVok50eIijEMPacsPWBqxQ6MKRG3mip
V4lR1Xgj++Y9PTWCjfpVDDa1PZw7pzpiZzXheTYTv3Qf77hXI4renyvzr/VQk+aR
owNJu8D0MVb9jHAVm4fyVRs8rbjK3b2khe2hqpneFUlQl6FbtNqSV/e8mZBcsDdF
pBDI4IjCyNsw7HGLavKLQ2ePCB3psU8o4r+lC2mxrhbuVCU5Pst5Q1dP4EpwkGi+
3USJeeX8akHkWAYeAYgof7Io2uvvJ3F5OTF0lfKSOKRHoJ8c/2O+SfNaR2VwUPLW
Ceii9ry8JVtlNr0xC+K23cq5Esm5qsvS5KAlWsgY6b3i9hqLP2MpQOgLW5/mu90Z
CoF5OK3O0PPHFSD/ptuxPcAHbDNvkXXH6iZFV0RSyFVUilFLVZHtTDHZH+wej47z
D1xO83bhEiFZSw5iBpG459GSPacy8gjk4V0z5s2+wWiG5N0ab2I7IH3shhd1mC7q
rFEVKdt68tqYHBJcGaMutfGSaw1zDoExqAWl2dbPe+ev0SxA8a4p3Kq4/CpXGdNK
j3Mu6PJ4m6ijdqyMMt5IIvxqGiRl54MVwbMRChoaMXIO6XyF9wMWQupsB193uTmX
AVysLezlZI5lf1MZvtTvbeJQEubFrcGK7KYgVzQS8zsjDpBDr2O4OIpAl+6FUaxh
/UP/N9ZF0GZQotLy/0x54byggFR0d/V4Pa0sCz/DcV2SO03ZblUKcPfz4mI2ou4x
rSf3u4CsXayPEo0Yoi1NLXLIaDMuxY0kqz/bEzrYx1Of0j8XCScukWCNMwRPImOc
cTVOHhgOIiNuJdWdAQI93RFDpRqyRXpH7EIMrbw8nE2O49BAikwTGnOMmqD1uWx0
gS9JJutW+rUnKvCmF1GGPFClcyrmdQ8FQOiLD7hlt0BMAIFcvNmICkr+WZkyXvyx
b7VhOCa1VxhJa6ZYva21EThBf8nRe2BjuCV0GnUxCXLt+/tEoOPybwcQI60OzxO7
RLJHNmzIYoUFQYsbKAPh12bxYIv2i1bLZbu+m+4TzJ8R/hCuXfGlsIedzIC9j0GF
excov+ARV/amKUzF/TsuB83Y0mihreseTpqlvjKj0/WiHmAgXOcPVrHYhOXx7/x3
A2xap3nuhwvqR4oEQ5L1/R/6Y8Ftv4Gdz+VcI4m5220wDyPpaXhOaKIke0eIenRQ
hwNAkqydRStPy7qkq6STH5VfbaIHQvdvViPYbIe8L82aCpLDzN7k0L3FoiPgGyXX
V8us+dSykg68/jrMq6saNicPtLUPfHxZy5wuxT17xoow/nwsbZeF3RQmIRH0Z0oW
Mq7KJjwHg3qNJy4ia/Ji/tA0yZXF5HduOaks5Edi1oMQds55hrxk4JArclPzOQrp
LDf3oQqoonMGV38pu0PAwINADNtXl/NXkLtkGCRWtF1cL1OVnV/ijUtcF6weQ4iT
pCkk6iLoa3Zw0cb5smRR0mjhM6ptZUUe60c+zTuEXB+m/hy3vw1qJpHEO0nKhbq4
AWg8mPbBlHmHsi2zjlR3i4qNx4QW9X1XOb4e7va8IGF6ouAD4iOJKe1Wr7Fgu5T9
iJOdETNCaKAga6BuGlVFpVf5/iABhES+CTUDiInSrbdN0A7jMJ4xlxMCSXDKGdBB
UJqvcVf9rtC1qD+Q2bzqStr+zRBLu9xeWFKiMC34aZbrhCMWfMOCOPLz+50BxGja
nfLua5ZzRtEbP7a6fydyHNUM8EU2COk14IBo5iBlkn8xja49jmrUHhqKfTMxvcm9
AG5PjKFgeiLXbneuDcSA4tsVO+TmhwHBq9890+ba+c3FPcg5UgIkt4FIJ3w588C+
NxXbO6lkFMY3weBXL5EIAybIWFbfwbP1Zkfz+i1GyWVemzk+ZYU1jjTddcPbBnA4
GciftZ00q9lMXvy6FcW/S0qKgENGylEQpQtS0GQEAbld2wpoOlWkVR+1gSFNFTCT
ACCt6+kfe4A6EYL3M7kLJu+MQCWGUiGw8f61eK/159vXS1DGUlLrK3LPrAiFXyDp
ez1hlweHmiaZzFYzOgASIDEyKs2GuyKCXwJ97IiCMubClmLVKUkSVclFlkm1JlrZ
o0X6VoM0MRMjrj+R/KRd1jXLl108v+6wqEzOBAvDKY3cgpC6b/E/pSH4pWSLBsv0
9iocTS3aAg7XauUfh/5uraevfBPoZJjen0VucF6OmXeSva5XyucpHXT3QRfRj5Ok
bwA4lIAT6sKF2FiUwzF3olahe0bAwI1lp3/fovXNV9LT/W9f03wad8jhbvHsVLac
+I9JI1WAGJkKqe027kMISVkmG4EPUCib4+TYFn/a5IMAc+tH0mormZinRjMoSHv9
lTrKJgj3Nb8UsWr0jFzQkd+ShM1FhSF9DqTFOut9OZTArRH7I+BKxy59d5ZVpjkt
+HMvBFzLuiByU7/r2el4B2zWitE39rzGcLCYUe924ob5PB3zuP2UnEPqse6j0/cP
OVZ/fXASF2BgvTxv3AfM3V36rW5VORxPRqbqHcxkUqXhkQqqHyW2dJcNVA7z41j5
QdwoHzBSoLclXQHAYYvThC3CJjN26/+rCwlDuTZVk7GTUKPcUE4+hPNMgKMbaQxn
HVDKV2PLzfxuI9eI8W1/g5ygkCyanqIoNjTyqib+0m4Ph8DvrltbahLTHw0ecbmg
l4Ty5ss8O1ccouq1ursKfXTQ//e0ThZycTAfKnjnzxFIy7z/MdFH0ob4U8Pzv6BN
KCjwFt0d1aEbfW5sjtERY/D9059nVCpc6k9Xz9KsPwvfCLbJbydpAh0QI5oRZHg/
jOnh9kQNgble0ypjJie1W5y+u94wDd+ec+YtaIl0SjW3uJEvgcB1I9UuK1Ue1yYt
xrX4CunNVzZj1yU0iIo5Ih1yOlx0aP/k62TOzx5cyL/JRNCc1Exrg6KybaT++npc
pisZ8GIyGAPz8VacqBlnKikTjkQYxHlcY94QMPLNh3cPtIDOIdXfJfXgHzu5EcK0
VDAeKJRZgvo0TtFIpp8l3w0SKQStXjs+jt2rHwIfkbfKlXTA5CrO+ekEEyJaq3wR
vJFPcEpGF3BMG+IH4bduJpWLbBJixbD1O7hYR8wMvdJ3v+tgTc6zCYyvuIlOl2Dx
zzp5Z7UpR2XiMWLv2TgL/FJfx/pqASKo3shxBZQDlwlq7iDsAxR8s5OTHJrYA2Hi
Xj8p9kU6lM1CNtkq5BOYHqqRJ1pvG10B49g4lUEfxsAtlfI1hEQIZNcFa/FSVRGQ
8MDguenY2xyl1mFzbnL/a2Uwbnq/5cGfx03n4f4Y6nwm8a7H0UWExgcin/AVM1/Y
T9RVwbU0vQ+HwBn19SKQcobo+YweH6Aqcqyf+1JmaB+at3NdNJoTwGccnSBDbZJJ
TFLg4bnDJ4/Buz8iUFThefB4KYZvayCzTLHpCLdNchzY0EvvdJjKGKHFkdm3IMi0
xkuN2EmYLCAF6iiPnru4SQ6Zi3uAL7npp1W0slMwpjLTSS3k0RvO7JJOIumunThm
COnj8+pntcRD3eb8YyymuCsNzZhuqfEpIYEpJYBLisj6olNJY0IZIaOMTxlPBn3i
d5HGWoGl0NyMsSMHAq6izrbxAvhDG2P9X4aS72bdmauTZndVU9+lmt244d22FeCs
M5OY8/jPGwHQ+J69tHSGxHgTue6wdg8DM8fW3ChA+epAJnxzdcb93fEoXIGS2NYX
KQwrjpDPKi20gyOl62KnXQeQCMQkaxqw6+ZBXyit5qhbLA1xVYAwVBt6YuI8fq9q
3uwue+KylYXMM1j27oUYhij0dpRTs09GhotpleBsrkwD3KaBotGe83kW//Tj1Lqe
zqg+fNmXKK2L2gg8fKGfLfH4QFYt+z5/B89QYAyzavp+C27kcM+mR8EGG9KANfsg
/HbrvjFm/hMNrP3oKsWK4/PnstWkttfqJavKgIfTnC09Qq5Yko6vt5ApZ1Pufzp9
OxYZrfxJzj4Ov3lx3fZGCUh++PtGNJIkTjWrs4ZxSTdO3P8eBADTw10pRHExr6Ec
/WxK2OXJO1YxZ46gxNHZOSiRjMDdd61DaDELN+wrb/x2pdhml6ipKmOOXwQdgE+/
q7CD1eLPSFIccRgUHFzcnOt4bE9WByTMJxD6Ew34ywzeEx5Mi0sK1jH4RgIpxzuo
wswRa3Bw9sWRKBwCWoHX/jodQusw/RHdjwg2g9nr9wGdDTdMjqUsVI3xfeOuZTe6
8/MUEcqXq+rHrcgX9stxe5ZXBUeHmKyQhcj9U8gHrGFsZh0pJ1blYYFo6FKXmU2a
O1teCe7kDy5Zv+bzYey7GmyMddfoY5Xm56xE0QfPdeiroy+QRoiBtA6SCrhCok41
1pd4jn0LRKyEI7dZoP3WiqFk+3tjsm2o/L5Z/9sHvxGgsU7/DbI8Cb2D/mVx5t41
PfSWdWuqLtlXceq5F7brNnpiGstyNGpmbigtBFul6xkKO5Ci3jXH+NgTLzOPQipy
Fppv59v38t9XvcT+yYuUJm/LPiqgf9MxUwNXzklyOeshn51ARM+DbghOZpCvxzZL
BAykxnvfEQikZumv30/LZw==
`pragma protect end_protected
