��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"�� $Wժ��Lg�7!	����I 쀸f5=�����c���n��w8n��`<sM�u�p�m�8ku�8"�֗��Ǳ��@Ϛ�����S��D��LĆ��j&5֠��n���H>�|F}�����U+���4Ȗ�p��l3��B�q��~�R!�)�ʦo
/f~�c!q%vn�.7���UF���QY����%��;S(�J�5l¸�H<�Λ�<~��'V���4�Û�氛
� bV@d��]foG�����1� 9�/�����X#;�3��;�����+'�Z�S���5N�)���G�i�7�hlȾqm����($L���ڀj�RT�nQ)ɢ콬N�uD�f}�agN���v���X������X}��q�Y���~y��G���B�u<�
-誴��Ǝ�����c����I���z��E�t��B�1i�!I�M�{굥�.2D�&��SsHRǺݩ���ۗ��+/J*4Z���;����+L�Jyck<�H�o�P	��:�q�m�^��I@�i��0.:�����ܣvC�q�L�I(rVu��0�)P�&�"�W|Ny7���Sjl�y�%��鎈�B�^������ �('�}�@�/���x� nR(EU�Z·�H5o{�]q�[M�" @���M��z���JF�~B�꼅�P�:R��7��z����:��>+���x��_Y�3�&�ڂ;�&�f��1@O̐�Mv9{��/����Y���o&$�9��Q _�J�6$_�LF�%����Z8-�)ɫ�����L�Ź`<��x��<gq4ԣ(ě�S"C�%hIh�m0�s���9,��xTۗ����q/C���6M�uF���8V:����e�?
�I���/H��%c���I���7	ɔ�u��(c7�_n���'(�:J�C�Z��ؐ�Ţ��	�%�ԝh���6����)}��a�n��������7�����) !�yٚ튛������fi�)�
��u���:����Jh���T��7���C�ѻ�p�\ͤ=|�%������ϋ�v]?���)�}4���:��`{*g��m�4��wy1��k���:��O��Fihl��5��ܠ�ț�9� �=��U�5��u}v�AR*�kG������#���Į���
R8��x�E�,�?{%fG"0�)�v&��|�R�L=}���
��|���Y�`!r����Os+J�����y�e@`���;��s��]���k�V�_���j�Q��O�,F�7|t�F,�֤����DԋQ,����mzd��as����������t:nC2�
;�\��������7��ʓD����U:�uC��~<6ׯ���i̥��X�l��?Iv�[�=�傠��eZ�獦�����Q��̞<�<W��&^��'f5�"�O�
���1R_����Lnl�{b1�1%i�d�[���CI8�񀹱9�d2��;A�3�gQA7C���-��b��}��Ǖm�=���D��G�,;�V�3���҅��f1�Y�󐱱�J2�i�l�J�J���4�2)�˴���X��2��<e��3�5�N�~�:۸�s`����<	�'g��