��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{�ףe��	�A`�������K���R�y����R��ꘔ4�Do��g]�v�f
g3s�ޠ��rC��u�B&$ش��^?�~�=���[���>{x��D.8/�^�_AM��	-�^��~����)�~Rِ����^���� �}̟D�!�P����v9����0E�-�i�zo����x4z&]�_N�t�>f�|���3T9>�.%ﮩ�<X嫹q�ǲ� �賴J d���lݵ���"\[�2���@K���V�ؑW��a��?�d����1�����'ɥ8�H�˰�naN�a\^�Iү(Zj�f�|.c�����6W}"��e�ȳ�|�d4P+�*���T������"�Y�bv��6hym���N;ӡD鑴w��S��0����c����cI޷�� ec#]@�;%�eO���' ˪?;f؁��-$��ܬ����\��)���)�-ۂ�_�F�R}�����/�6��LM��P��X�`�A�0M���Y�|6���s�`��=�K`�a�)l�u���� q�]-nv�ƶ�����&c֒y\-84.���	�S"X�@�.��
}����>Լ�1wq@�Ø>0x�ӫ��A�e��B��4�p��1��d�1�(p>�7q��rjݐs�TMԑ�ץ6o��J�-���#d��՘҈��x��$���>-��ӭ(˼���}`V}�~���Q�m�C]��j>[�\��;.W�Fj-+2΂�1�� G��d��?�!`M�QH�r�pƺ�S�{ 5���*i-��g~�S`gl�d�퇝`{�W;��Q��24Sz�9_u�e�t�����jF;]��B�ώ��N6��2�����#��*![��5j�{��9x �����$u���5vȕ���E��va����
��_��%| ��o��+���sPhGNh�"�A<>��X�x��+�D֝�6�Ū�!ي�(��-�Վ~�]��YC5�SZ2C��r�eɧ?}x��RSr&�rc�{��x��N��<g����[e��e���XC��n��́]�N��Č�S�H?#��5��v-�vi��2�G�"W�m��@�e%�DE[���<V'}ۅx�Z@7XL���CM�|�!�e�\飯�;�*4��������~�ڤ�*�6^F���Ah��)(P�A�O����|�L2](�X
���@��9[t��8�~J��=�X��+���Ox�%�Ҡz&�^��{s��5�,�.>������*?V��W�?��:s����Y�~��輫+Y�*���Ū������S�����L�j�s#�U���(,bݪ�Ş��'��]"�!�٩}<������#���^V]Vi WIT'ֶ۟[����u���-|���J�4��ۺ������n���
^M�5G��4�.F��װ j]_���On6�y=�?�qe��i[�������n^�"�`�0��o+�?��ōȫ������xv'��'{�*��I�=OQ;$�}g��20�n�Q��C�?8f�S�i�*c28M�9�U,]��d}:���2�	(��C�h�&�װ6�h��fp�K����*2�=�
/'T�J�g�D���Il���oQ��t��8��j�|��a��׶����6`\��R��e��f��s2ӝ�s���`T˪r�].����n�����\�Ⴡ�]���uz�Ȋ�BW�a-��Q���o?zQ�a��<���:Y�8�k�b�����4�bRU$ ��e�@+�&B��Gy��1�Tz�������T_��V�p�u���ƹMz;�;�@׍���JzJ�81!l��Ec�����b��
��kN��qXIT͏�kF�k�-=L���~��AG���)��+�Y�R4����3��^ǽH�!��M�e؊�-���9r`*����k������ft�D��T ��6A��(�ZB�� .��0����k-U�ZE�'+�k�\�>��1����A_�La�VFw�W-�Q���(�A��1�[r�3���H4�G�f�����V�wm+
/8���Y�v/���0gʒ�9��R�x��U�㪆�`RV3��!�����nݍ<E�w-'r�7��m�4\Ådݍ�^bT�=1�¹]9�"'�­��Mb�|��9n�1����l�򳰂�N�����7A�QcV�_@��}�iַX���]��Ϯ�|p�~���>���m����>���;T��M����Oj�"��]��N' ���������KvM�ި����^�Xu4�x�¯���A�Fv��B�j%pd`mǃth���ѕ�4�ağ��O8\%��xsu�}�G]��Fw�:D7똙�K³Mr7��|o1��W�#�b�Q��,��7���ED�$V��u4lG����PK����?��y��=���7�&�5~bs�q������j�����v-ui+_�c1�ƕ/����b��45���Gs�3r�}7&�/*߆& �dp���+�T�)���HnaI�1�=�r�r(xN�]f�R| o����Yw(��goJ]B)���c"j@��h�&�p1�n��&~9�E�}��I��B�%r�5M���Vd��Gڃ��^W��E�&��T Yj�U��Q�S����p�htR��U��f�o��͎����4�v�q�O���koiI�C^�ᶞ�3Ć��=-2<n�β��0��$2��9���>í�*���X3\��ZT�i\���'���/t�Y&�<�Y��