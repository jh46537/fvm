��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}��������r�MX"@�����s���(�)���t1�㿃�JV:�Ni2��߀�ϢB0X����E�m_J��Ì[��l�(�B����
�e�p�W�5��,��D�Kj�ώ�T�����QR��@�����s8��H�>N-�(����T̶��	�/���4-��3�)�1��H����Lg�iH�;�'�Y�N���#����r��O_�Q���+���b��sQ��3D�U{=*�h����S5�p��]�~<r]����b#j	[�і=���k;��@�� ��W��t���<���F�̧
F"ᅮ� L�?-м�+7*P8�NN��j���F5�0q�%T_�F�6p
�$(��X���vѼ,�3L��K�#�+�����j`�j)^��ы�5��U��Le.,�n����(y�=P��׬�|l��-�i�)�CH%���C㩣��9��Ne�x�s�3�H"C/7�p_�L-�s.\.��59���^�V�L�@��q#�[_L�{ﲆ�k>��"���q1��K5u��W���a=�2��&�9m�G�n5��L��-�G�_���a���U�ޮ8�iE�E*g!H�oi<�y�u�W�J�`���(�:Bi}����u��~���Y6DRh��W� -�Ġ���1Z1�6������)�!?��Tl������Bm�Q+>t�n)���/���Ѡ���HBƜ��7n��0���+31��4?[�d|�lqſ[��t��Ғ�ѿ����a��Ⱦ!7��Y\�N��	��[�h0�P&�<"S_p�##� ���'�V��x���۬��ȷ�= J�cdZaD��t�����s��	�!*��L��Y" Ҁ]���a\cg�W���e��A�8���M(y�2�p_2��"l+PSB�֑�ߛ<�YHz��!�$�!����[+Q��٬�b��D|�љ����4�7?����Ķ�8�������S69�J��J�MYĚq�H|Եx7�mꊠ�W��냐:��{+P2�܊I�q��vAH}5�#�7�t:=!4�D����=.z����EE�:�ۛ�O��ӆb:i��CC��JH2H��~򢂌��L�����?�I9���h�
?��6�h��ǐ[{Ɩ���ؖc޵<Xz��|�D��1�.�U��,�����*#�؛��lִļ��u�)���(�`ī�,�M�]��G7���k��TH��8j�:������<vK��)1d��r�� 'h��@5��]���W�9[��)O�G'& >�3�C�eu�T�6�s��-�����J�c9��m�k�MݍH�4��Ɉ��k^�E��ZFB����O�yW���b\+����g��0���t�ٳz�t9Mh���әx���4�eM=�A
������o�u��"^�,K��ښ�! ����0�!2��͛�*�*�B���5�0��y������k|�A�Ƶ	K����/�ݠ�m�R���A�n�m��.��ȅ��M����a)3"��&���E����'�	��Ղ�&�nɝ3���c����/�ѹ�S�d��A�x�3v���r�L��f�XJl���5��`#��l�XK�?9p��w�ؒM�s�Ŷ�+�@
�9'���?��ѠU�k����ݦc��o�\����&�{e��dV��ݡ���.���͏p5\��	=ֱl6��F~ΌW�yOk!��'�)�ɓU����^�+��Ɣ�FW.��Oi��M���^����.��	;296���/��W���yP�S�*��ٛb��9y8)MJ	����L������$�I��$���k��V��4������O�
f��5=�����-������
fڪ`,��0u��p���V���Q�*]�zх��*�Vt3��e�C����мY�����P�>QpIYƔ�����C�o�e�C[�/PI�q�,jɀ-��ʓhr#õ
�����vo�(�)���;=n
_j;$ԧ:�B�N��d��k��~�zA�,�-)WO
�}h�u`�2�VF�/�T�S��o$X���UZ	IX�tg ��}y8
��}K���Ӈ���5����?zm��;.�Ueu��j"�0k����Sk�2׳�������\u�o��L�{��*[n��;�=�$�$�F�G#3(bR��m�%�#r��ú�@M��ﰶ*;�t�!ή��ӳR�eܗ2� �3[� _P�ɴ�yȑ�>pd�qC�%���F��KMo���l�>@��JǓ|,S���OP��c��84]��K�Jij���C3��?~��A�G�w�*�E���S��kFj$�#(y��JŴ��ɢn�2�/u.e�NDnGmK�����b�'b �90۴���s]^X�������0gK�լa��IG����-��#�y�k U���������ۓ<�f��W�=0��n���<;-�M�K�HH�`�{p���;�6�&r�]�o�Y�p{����3t��gũ��TGaٿ��X��%�5��Q�d�|7�5[L��ޥEX�oՔi��V�����a����=��y����x��!pU�4��k�*�N~��&�>a:��_�P�ZF���SLǲ�D��y*{RN7g����6�T�ƛO�V��+%چ����N u��#�s���!%�}e�-�������G^`�mL�Ro��cM��1��#6	=6jf2i4[b'+
}S)��}����)F
K��搓c%�����q�]��?O%�%�/��-	�ޠ�Ղ��g�2�N�(�@��_>���P��~V�(6n�V���nZ|�%�N�x?>�n&"ŕ3S7/n��p�0���3 �b=c�aYߗ#�5��pE��=2��`��1̓T��Wq�a�I�C����`�1�W:5�qZ�Qw+\�Y<>, ���I��ڳ���J�֥Uh��&.�`��&�a�0��x_'XCM)���>��Q�Ba�+P�*�o�)�?��ث#p��H!	� _�X�������s���*<.s��=����@��|���~�cR���[���'�s �dT5{�j�S?�<�	-�ڳ��i�}c� [����-���L��v�a2X���y����t�����Ct�tޘ���|ŧ�J�[��sܒ9G	QP�U��6���)��0���6����T���W�p ���T�ἸJ|���ܔ� E����B���%|*�ԅqg;����g-؅l�
����q�����5��G�՗�ހf:4�ڋ�ȗq/,E��]8���5��Ε��6|t��h�8#�]y�͔�׬����7�M<�=O���l� *�eT�TI\�e��:��ز�q�(������֣���gw�\C�耴�݌)������t�SL�r��Do��Y��ܟdugTN�	GNx��ͦDѤ5�%�\��d
�11\e��|����'p�>�˝�>�Ǡ�g"�y,g5a�ޜ�&��ݠ�5�X����y
��ˉX'Q�f�*�]�w�G��n#�&����Q�+L��EDA֨H����-����p
0�{�����#�s�5y��e��k�Dm�69k���)sh>��W~a���.�Lcd[�T{{�����SI�7�y�4w �X�o
�0�g�఩�����ٝG[i2񱵆^I�0��� ���k��ӻ	C��U)$X8X������+n�˰"�\���0 ��
�P[.)������V9Y�7;ޕ��-_T�^8� ͮ@���*'��0l���`@������>��h?�6%��'�aKB���;�E44����B�MKW1<���q��n|D�8��[C������f�9����v��@nP�&UƂ6�X�>�j_�������R��K�g<7���Q\�쎝k�ށ*hrx��R�J�ڳ�0�i
�=�^�-���+N���ڕ�Ԁ16�B�����5g��M���-��T�]MXG=�@r�?f�lTR�����F���ͼ	$�/�� �<�9�<�ykKH�Й����|?�R�2C��[�x>�1���r�8&��}�^A!�xԑu�?�8���� ���RA,����1�rn�c��pBTB�x��1�4���>�/�؎�_���c�������z
�t˿U�9��̨mÚ�;�����5��}T����)G�=�T��E�o��PXFk��NW�� g�߫������KLSʳd�`�W�!uR�A�?�SƂTsx��v$�Ac�[tUHV��,Y.�o�W��������M��;^Q?2{��!O��y}���q8gi&݁X3�teʦB��ͬ�Wq_�3�)dܻ��w�H���J ���~@d;U��xw�v<A�;��at�}�?��
�J76	��!c]���tO�Ve��Pm��ɚ����̓K��j�C���o;}�Ko�B�竃��y�p�jrK�Ƴ?��H��~��QB�<������<i+�`%9^{�[�b�qYfa���Y��{$�p!��:y96׶л7�ՁI5k�,�S|6q��!�0T�Z�C�jѼ�@S���_�=l-�F�Hz_�ރ&r�{����q���0	>w#��,�mh��R�{���f��̠�WT��D�n��-�ۓ]���/�;}�$�Em��<D=��[*Uˤ��6��x&��"�T��Y�5�Iz� 4�h<�ϭX��^ k�ړ�p��҈�F�34��E|���{�������
݄W�p*U�,.�.���_�ڿ�s�B�È�ơ��֞��\j/�R��ew,��^\�ض�}��ٍ��.������
��4;��:,�q02G$��U���Օ�`㨿CO��ڳ�7��Bz��y�W>�Ԛ;WZp�p3<��dns	�"]�e��	1j�eKBG������w��8L�`��H~�VqA/��E�ԣ���8<�N-�.?����tDJZ�wdR�w/-��k"p1��E��Y���"�,�H5�Q�	,ல��A�$K�JZUZϷ�Ț���4�넍*N���2�☸�z�x���4���NpY�϶*�"z��4X3��kJ"`�*���E=���r��Q�ҏ��qg_��d�o������ʅ�U�=���Q�+O�^����2��;�9��G���l� �@Sf�0�|b�ϡ�)�{r���zo������֤T�5���L&��lN��[8bV��l>�KG��쐤!"���IG��ԣl|l�$S��H��T�Bj��X��d�X;[5�~�z4#)�23=U�a:fO�5�3>��c�,�J���:�	^0�l���=MZ�p�Ja�%�}����G`%�ٽ�8�  o;j���Oy[�3#�졹���1p���i%Ϻ�*m�˽i�V����|~΅ûr_:�����Y�K<��=mB�������"C��1�c�q�k����>���T�[d
���;�Ae����d��,5	�OwA����_DW&��ĝ���fd��A�r8u�14
{O���&?�?d2Q��I����"��L��ݿ��=/jUAv�3�[�B�y�U3��b��+�(o"�����q_�No���Z����f��J7ݭ�`����d��2�bS�������]���k��zE���h��E�g:3{�L�3��H&�U��L��q�*����'���6����Rʒ�f���4�^�LO�վ�Ԣ;��B�����A�c伸��)�=&UV�w��n��1�)|@��J*l��ml��C���?���O�p0�n�~�����euE /�Tc�3#-R�'�N�����>8#A=9Ud���,bt��bbڛh}ӲxyF0/�N{;��)�����Q�Ս��4c�8s�����<�˾����g��T�U��)#I��ѳ��<D=�z�}�	�vO_\�Y�QD=DW��r���h!�]�hȎ����;�,�y��!�Һ�R_�g�=x���B��w��s���=����rZ��(LC�ˍ���]ی������+ehP9�e�a,B_j=�̄����(���l-y��M���$]*pv�t������V�Z��#)�u�Q.�v^{s�ן{�����b��8����ϕ��J�p��e���M(`�&kOx���F�.�3dT>��l��R���x��$*��Eҍ+��xHN��({�Af��M�#���_0��C]�#�b�䊱�@��'�� x��O��a�Rm�v2^� i�|zl��'�6�:�#�.d�яY"W��M�#K��)7��ܞa�Z&b���&B�-��]�ԙ�Z؋EJE���3�#��B���+t�f�~�߯Fd��c�s1Eo��>����y�E3	��(B�Y���=��@N��Ja���bެ2�7:@�Y~�1�M1�J����跉�y/����-�B"�W�:�[5,�8�E�ku�����f��L8���	V���FH�e-;���c�����()�w�*�q r��J�)	:o�}��3�KȲ+	_�kh�������4Y�ť+x32+(�h�����j䗓�A�
=C�f��-?N;����
�oy�xT�O���q���W���`H���8b�Y����[�Q(L�� ���3�Ģ��i�R�o�RŌ�_kP܎��)��cgIƓ}T��a��TF�Pg�R>���GbIN���lQ#��M��h�}*0���ٱ& �X�so��na����P��U�.�
p:���NE��M�r�4��*%�MO��.��7���ٲ����a�����kgԳeW�+w��j������{
j'r�܄r8ǥ��;��3s�jo=6��tύO'9��E���`&�^"���b'WՖ)t4�RI9��Fm��	�`��׈�e'��_.�dor�C�b|6�=T�1���x-�[���z�*���[��=:�Yz��'�J(�Ђ�p��F۽}xix��mk`�;�,7�,��g�qR��)4�럾�P<+8��p�zy����y� g6��`�ao��l[�F�s�*�B�[Bk��Ȋ8ww:�փ'�QG�W�}���X�A�3��� �����ݶ��x�
ϗqC�<���J�(�Q-������Xhs�އ!�h�8ǣj�T�'47ť|R��j���$�� �&�fb�d�����T�ep����	��X�A�p�!9�ڱ�-��WLU�����Б�c�Y��B���~��E-Rd�J�kw9�6A�b8�0�hW-c��8%Ά�Os�pS���kOEHm�ġ���6��$�B�k����&_��g��m����=�.����rq$:�u\P������� o�`z��8������i�����3�_D���фH�cx;���rj�c_�vU�jc-��C� ��^�Q�c��8�S���&2ӝ����Ӂ����sf+9x8�z�8-P'�^{�t��ˣӬPw�=s	��e\ g`׶�9�(�����3�B��=a�ι�n5ʜ�s�g,�~��f*4V,+�#L��?�����	!%a�߉��ШE���I'��~��i&������&�����R.K�qn�g���Y0���&(^o.6=uɎ_��p�#��7�F��C���"�yNj�
e�`������Y����S���a"ʡI�4��=-�U��i��K�=��to������⋿D�/���jW,b�>��K�C��zZE6c
���B�'^b��2h�Q-}JY��;����<v�l�����hGJ�4�c'�&I[t��-m��I�V�{'#�����@_�w=���
��A"�g�Z�h�v�j��	,�7s���ޑ���B�����z�Л5a�UYq�`Ҋ�p	GgMʆ@��/������<���V#��U��95`dW�a2���c?9Q�#Q�.���0�|`���9��i&�+'_9�(}���?���;V�u�h�3%�c��rӚ�k��s*�;�D� Ta��˗oɬ �>l�����TON���G?�æ�DI�\�<��v�\�\�p�@�<�+E�$h�k��GF��%b{=?(C�9�Ϙ$_���.la�p,%�Ew!�6�)^�69�X60c�����EO3}�P��*��kT������jw�/���hn���� ��M1jz�!����y��e��N`mmx��d��@�?�2��%���b�m��Y2vxS���)��9d*B�v�x|@9��t����Iwv���ˊn���%(}�/J�.�L�Q����'#�^�����\u�nFoD��6�*Dy��n<x��/y��isB�&���ԁ���:�[3l���+k7�KeQ�4�x��%A��X��J�����8�1�\C.a���%����w����u3=ep��]Vf,�<<��H���˚��R���Th�ia��b,� '�<
��"��R^��K�L��O���!̝�7֬��sW��"�v��Z��U����pF\�<ΨD���.8�^Y�1	.�lέ&��;���;�����r��[&�^�J�?d�G!}�X��k�Uڽ�� A��M�*����Jp)ߦ��$�x�t]k|(
�mG�/YW�j���S���d�E�yұc�]�AJ.������<�x���C�yL�K#���	���-�؜�� 0V<GE!�mu34)p<���|{�.�����������~����K�K"R�&IU΍$��|a��}��Vǟ�"�ISD^�d�4�C[6���v`C>0��p\U� <��CE;� 5�>�����tWR�^8��l�b<Ã'Xx"����d~Z��L�:�k���p��B��d&bQ:��0��.TLJ:/����V�,�'`�]�.���m$w��>�@��O����bH����Hf{,<�I8�p��d����r�9�e���}�W�kո��^.��=�M��m�r�����7I�^��{�n+�\l���!AJ,"/xz
��	6y�r��H��֏�ȃtO���՜vu�r�����L�(且������Ғh`��F ȮE�3�!>t��1��E�u�]O�x�L�Zji�q��f�Gȟ���p��)�k3�ߧO^��7�i�@k̕T�UhHE����ZA.�}C�FVX�ś��v(������:<c(%u����6Y�,������D(L�b�!����(O].R���]&��Kv��PTL�8L��� r�m6�C�2�+>2�ɫK���~M���?5�P*�l0�!��PE��m@�xG�0����Ho�Y��4������!n��R[��J�����x�Jͽ�^�+�1�w�@X�Q��ލb�����i뺍��o��N�c�Y׻����!�"� )䡹y�C2��oF|�/�x����fY�$��A:�4^���ʔp�j�m�W����%ɷy�|�A�e�l+h�o'	쇵�
��"�Y�o�ʺH�-�,��oG�S���>�	��]�6���b(bVո��$�K��+Mi`$h�����.C�4G�������X��D##��T!��B�'�+���[����gD�h�)G)�ȊR�Q�"���qI8-�؉i>��W����6���3��)�4\�������%���7��s>f�V��8��Pn�7�A��Q�B�s�kB܃7y�Q)Q������*C����Bۑ�kKB�$�$E�Wʩ��
.q�D͎�L����9ל(�o�j�ǘ��Ro����p_ґ��_��G���H9��:~_T��و�a�4�{�C@�g���U�qIv�/�L�)�\q*	�a����+ϜF�<��-�"U0�����Y�Wh."6܉�%��/z�ł���VX��P��Q0�Ԥv1�h�=zI�-R�s�4����{�@{�P̡��z8-ZU�"7<"
���]��M�A�R�ui��H�7\S 딈T�Mz����g�Yd8yi. F����GA4���m
O����Fe=ɷ�V���)�'h����bD�6��L�T�����*���b�v�l���̽��YQwg{�@+��L��:v��/���M_!&.h��j�?���4O���{��p a$�����Q��Gt�N�uU�r�>H��c�J�p~ ���r��P�|����£ݫ��ה�n�KM��<�J�7k���z�|AJ�7�Q�~{2��In�Y�}�"���������.�7Z�+��1z��V��V^m�4���dHIᢺ
�-N�ד��Ozh�rv�V��#~G��N�ޖusS��k�BR��e�I)��∬E\��JT1�0̅E�Q<2	60�{������Q�K�S[%N�p���E��in�&�.j�-E��6��.L�<� ��V4l-���e�1�rz��t_sk�̒��_�`7���X�tq�/�M��F�_�ofNV�*�%�o�HY5�p�Dk�
@\���ͩ�<��>��6g�=��Hdm[P�	��g�E�S�v��zو�o����.�C������EQ�r�{�s�b*^O��[�,-ou�*<�N&�l·��Ȗ��_�Fh��[P�%�c���N�`�8���1WIވPx��e��a�xL�)��M�;uL��x��G�Q��e}7�2�
��H遪{��޵is��hQr�0�� S�k���V9���><���ޛգPVW�J��F/.��Ƌ].?Le�f����V.لj���P+�Ғ���$r��*[�У�>5����'��[��>�����>�[�21�2Y�a���Zk���egO�	�)G�I�?�וi�W���֞9�m#IȊ��F\��tH��y!���	�L�TQcN�֮~t�uA��#۳Dn�v�Ւ��a��L��r��j�8-]�����d���bUc{�h�D��',��3;��֎.!,ʌ��(�}ͪ��HF����TuP�T;��yv��*���W�iE��Yʁ�Dq&���}�7�?��5�
���\u!>Qب�2�M�=�w�/fX "�f�Z5�ٛL_��,�I�����4���H�
vv?I����W_I���lk����G$,�Lf���1t�ɠ��bh�KB������/�!"uoM^1gP��&��θ�V>x^�;	?�:1H�i��.��w������� LitZ� 
�h�����<J�V�����#�I	�G�mV�#�G&(������p/��o�3��i2��.#k�EU���E���b�N�U�,� ;�8�A��A����²�y�Q:�K�������q���뷧'�����CG���G�d	.��F��m_&�9�4��2C�"'��5�s�!���X-�|a�	���O�?��;zjC9��>�q�,�1eH����Mj�u�P�k� h$��d5�J��óXY���FLNG�b��U�y
8�ӸD�(��c=O�+i9�v9)�}��&������p�W��Lv,��?�͌G�r�]�Ռ/�b���SelX	N�� |R���Wگ��-�S?;!k��?�~����yB�G(�~op��F�yY�Vad�ġ���ȱǜD���y��;A��T��%��)�����d�&D�T�N�D���7�qv'P$�S.`����NDe���J$�Ӻ0�O=������e���E����j$z�S,w�2���9u��#n��+�5�$�N�Z�ҟ�����Đ��ӓ��X^(�`TX�2�8��0�><�{�ڣ�;��OY<̫z��������`z;�,I�|���f��<�*(/����t`��o+r�ӵ��Ɯ��B�!�6|8R����CMv���g��	�3��H���0Z��fy�A���(yŞ�ŝ�T�G=\�&d�G�ת�6��p��W�rb��4����1��7���&�ç0�O]����v##��l=�Ԩ3��V�Q���f��ܤ���JZ��i3�]Y׹�P���XŽn����=s*9��%<q���m�� �����;I�T������}FF> ����t+D�3�7�@�գ\�@�n���g�SG��t6PL�"�i'�בh&�F]�}`�j-2�CN���7N(G� ���/��;�'��4����&�|�ޅ�bk�nRY� O�v�q�5���:k�}M��<yc\z0����=�OU�y��g)z��$)� 5�n]`̑�L�&�$�:V����޷�����h��������7�� ��i�#��t�T"oл	Ojш������qt�M������E���U|�C��yD����U.7�1�N_���t\���Ǐ�_���/oO����8�6v�͌m���OS|訄E�Ƚ[�e͏<�~l*QroT9��ܶ|J3A�� @yX�yI2e�魑o�ga�MB�Z��a�%N9`ӂ����~+�i���3Ͷ�o�V�wxE8Ἂn��ɠc�]&km�<��m�iC��@�����Ѐ�����4<	���s����&�pRV+F��OY��N��-3ȠSY� .�	�S� �|	�/޺ �ԳH#!$b�s	~�ژd�f�C��MlŻ܏��^}\ᗏH���)�5E�D����<724"��]��F8 ��dvFO������,�	��v�)լ�p+�-�r�hrcyi3ė�9@����Z.���D�?���[� � �8L6�=�m���tҷHr�s�9�T�J�1:��_#X���������@��7�~��/���n�>	%d�՝^5������a+��1	2�����P.{��0@8֢N�O��j�C��.��
�^��af��#]�0�c^����7�HJ۳9�Vo�f�AVDA0����?������d$r�U������Ub�-GÊ���$Z`���L��ΗɩZڊ�s1f��|Îb�j 
ԼK�/��Vo�mu߅Y��8�r[󛱂��3Vp=!��#��">�Z����i	�����Ի,�\0΂X�܃���[=�A K0A��9iF���q���<*i����]e:�����T��x���� ��c3��yV�A��ߥ���?���pŦ� ��+���	�6�~��v���7�(X�/3?� ����ӭ�_vq}�|�(n�b�k���Y��".E�h��1$N��3r��Tl-wI�(SW?E������g�_z��d��`���ӻ�?Q�5�}h�m|�2���;���4�W7�����`�*���O!Zu�P�Lp,HmX3��Q�HB>!��pV4�.�n�Za��(P>Sl�)�9]|���,�u�8�#�����{��:�Ӫ��ȫ��kq<1���k��d�*��q&ũ���/��_YV1d��bN��%}ץ�x��S/@�2O��"Q,#����NJ�&��Ҫ��1B��[8��5	���3�gk�,	� ^|����n�s%���SZi��zE�ͪ�,��)L��a���묬������
��v�<�s1�A>�@RI"֋��Mm?0��̧�VU�f��ȝ&�sv�Pg��؃1��{Mw�,���q����J'�6RF��5 F��;X+�VqҌ;d= t�Pzܫ���C
Y��7������(Q��$��}ka�M�����~^#?��?��q�y���H�z�4�x ���Y��'ъ����DFn:a��/�t[so�!(���d�&�����5�"��ҕ�#_x�p;�� -C�!��)�2��ɨ��0e�a�>��wkiq�9����W�=�g���)��T�^7�&��K��M[�u=��ֻJ5A�ǈ-ZIՇb�9R>��I�D?��V�6��>��v�l�%|E�2q0��Km��h�IH���e�1(&��*��K)��.���8n�@t>C�?`��o����̹�w�Od�B��SP�y���gp�s���#���[������l��a�T�H��!8X�z�T��e�d��9���S�'`�9Q� icQB	
��9�T�������DX�u�@S4�/ŞS�N�c,��C���)X��%-��TsI``b����B��1��b����qS�d;6�yK���w(�ڠ�jY�KxP�F�3�Q��%��
t�L$�2ڇKo}�಑��w�B��x�~ �)s�X���E�wN5�.��|1^%o�L{!�I�Pp)[����Ɩ���Mj��I ��}�����2J/����w�
wJ�� ΃Q����!W 1ɵaγ��0��(IuofX�(Q��.K/�$��f�|�}����du����	
���g�r�H[��nMy�� ��?��u����/��>ӛ�C�6�:����/��G/�=l�׵Q�(�>�ޛ�;5; �?���QAcl��0c������˖[x��&�+.�s�ƪRI���'*^M^�`�4#�[1B߰!�6YA�I�' {�ơ�՞ڂ	m�S�=�^��[���5̐�4����K��dv��o�<�OgjT�\�TKa��$��b��8�9�V�w�I�$��C<~��ٺ�_�3�G�KZ��6����4�5݇�����7/ߏ�V %���0����{�1Cu��q�"s�'|a�K�Dv�y�L$S��k��^i@�꼶?�ݑ�A��{�3 &:����o�#|����&vt$Ѿ�L�gБ��|]��4�w���#�C���������|r��AL��	�m�&n�n�
�t�sԏ����"�fߕ�<2�b�SDݰ��2��6���~�� �Zs�5�ܧ�����>��	c qD_��aiD�l�m��ҟ�NXk�t������Ʃ�gI<��6�&�u{~$aKdx���Y�w�H��ݴ�>T�qhQ�;�M�ysb�wo�O�-!���q"a��1bM
��;7�H�0�+F��s]K��ߋ�;8�ٝ�<��0���w/����v���9�A��̖?/f�:���	F�$���Ħ�G�8��0I��;�`�Pt���sS�ꪓ.�!>r���%�qڅt�z�nEU��޷5c���������ɕ`��ݞ	��z"&�^����~zʄ�� >߂Uȷ��)��B���`�2/q�:���:�I��L<�o�A�|� �Z�=A;�aR�	��¯�Y�fS?�^%�A�)�zNs�ad^sqj�q>�AZ�� Tk'�\��H���s������H������*|�B����/�1+�*%�[պ�#��c5�,wݟ:��R�5e���� ,��`��'�}�̴� �>��L;�������b�>�֫���_��U��fxY�uƃs�,��h� ���K�e@�����VKY���6�(E��vdg��ٚ�e:�֦<��(�g�m�0'�~5�F����1~���d�L��0�k�Z4Fl�9�Wj�38�x���3��Z�I��3,;���q�t�{�R����7{��1�Q�ǿd�#��dP���KO	#�OAC�e eJ��V��A��Q-���bR=W�g��7���� �#�b�	{�.����,Y�\]�`�Aͪ�	mLZCg==�X��R�agH�N3�TFEo�B��#u��h`e�De��ϋ	�ϊ�0�}�a�X���(�1�?��.�B�UEx0��C&�#��T�)Ϡ�d�ּ?�����DRy����8@��F�;�L�H���wmC���e"\\χ��Vrz��э�5��7�ߗP�]���JMA	.hG���)�'sw�
��8����^i�)�$���܆���q���#��}�s�.2�����F/�_�d�e�g�9�3��j4����U��Y�p~��UvuY�U,R�!��#�I6��ic3�R�9-<ȶd���T�!s�K�&�����Iv2Me��`5O�����eFy�3O�N���M�$��ٴo���]4=���w)�u�(O ��M!�E7c!u�x�!Co >Ug�O�$ 0�<��*H����ݿ�6��x�ߡ���LN��b43�xY��?|���e�5v�8�س���"@VW��N��A��[�N4, �������
�̉�3����0�29s�������tr�!gu}�9q��/����F�9��m�/� @ݺ�8���P0���.��<Z��8(@�-
��#]άg$#��\����r�2��T:l$I�����tר����^wA����k (���qB�A��G����d��Pl��4y�����ؔ�m�V���.��)��I��$�2����{V�ؠ}�GX�5��u+�tȀ�|MHviQXu��+�D�ڌ}�fX�O���I��'����A�;Hj�qT�x�#�+��N;_�,��)/�u
H���ˤ]��Ǝ.|��JA�3����D �"� ���#E6b����ŕ�b4�݉���z\�/E�9ro6�OɆF���v��w�z0B@�n{J4���Ӿ��2�X��<jO�-�mj��	Ȇ�+��h��6nΪ�����
�#��R�H��)����h��z3��U1�`�-��U��)�Mq�}�oO5;�]��b��N��A�awA+Wiډ�),	ζ�R+qO9�o?�<�;�?0r�R��7�a�zCk�!`t)���/_��.X�����3��N�z��#�6�N)�4bF��H��v���ۥ�IC�l��Չ�\�v��z9���Q���� �y�:�V��Ð/���n�z��9������i3%zٵݙ���#�HC_��Zب��d��\7^,�vL3+鴇�ae��G�6�x7v�|T����aRR�	��D\���yMY?��3�~71z�'��_	�c5��l�@a�o�>���RC ş3Ǩ+'�r*<ᓑ�)�c��5��M��:KV�qF�r�D���H|�0*�r�S�U���5� �b`Ν`�r��E�A+�h^��Ē���5gE$0����8^v����}�a���fi�eP۶��?	�z����YD�!�ߗޱ����N� ���V�W���R�V ��]�)� ]��B�g��i��J�)~"���#�=>�x�����Gt\�CG�s���z�p���F�e��)�z�t�Y"-'���hu�C/��0�n-�ٞ�nt��_���|Y_�5��|�#�u���ӸK�N�hb����� 3'p�p��`���&pB�nlN9�W�@|�a�7�m"�$�W{El��L�Ϙ��X���_1ӕxi�u񍦴!J��"<�/�d�q1c��;��:"��>qX�zs�CW-��×�
���~�{�5,6_f��4������Y�k��)V3�i+VキO+���Ȫ��I=���{��Խ�u���Z8`�{;��>��-�ЪnH3v�C�O��}�z�w�G���K�9"����a�~&�o���{S7!���J0������.=#Yb�.���ɸ�������<u�����;[�-]M0�J:�HH)X��H��v��+�=�b D�#��m1:
#�(�	\ܛI��+)�a�g��'�����&�qn�[�ѧ�o<`�n�5π͵�}Y��Őx^+5��cPQ����~����z'F�l�o�%��r�Y$)EI���j:����r��ՈV�m����Fe��T��
�d'�x�a�4e�����D��$�V��m2�`�ZƂ�A_��g����`�ws�ų%|X�/�v����u��SO.����%�4����gW8��q��(�:�?0A^�����y��<Y�v��"l��-Iߎp|�S�p�a��V�R�[�d�������
$�Y� 6�h=0m�t[z�+�@~zRB4c��E���b������u>�c�ɨQ+�P.��;�5
�xܺR�.�e̹���e�y4{82�H/��>]��1��9�O�F ~���O��*�Z͔+%��9ƮL[�*��h�U`�(�u����4���<J�AQ�:�jv*k!G'K�"�ĺ}� �$�!��n������<�������1��"�@B�@�ԞE��@x��
�P��3�����{,t͎f4.�x��^ ���0;fA�D@IO��Y볯�����o�1P�W�P�)�@���r�'A:��bm���l�9��Q��l5&4߱�A(0w_�]�~��?Z�v�G��B�����c�p�'~K�z~e����գ���%�cR\/Mԫ~�%��p+��C�vq%� 3ǁB&���уO�d�~�o�x�d����?���u���)i��Is!�V�k�hz5��s����p�S-��������pc)�<'QQRdow�7\� ՘Fo*�F��E�ZUJGAI��������H6\�$Z$�?���� ]!ʢ�@o̾	�W�"�xv��Y+���[�p�,��XɦTĉ���8,:�|L�B�#s]��^H;��MuKe���)͛�J����C������ߐ����T���;��C5&��j�����K;���$g�7��j��,��4*3�{���
���J����t=�j0��|P�e�@=Ly��<��ڿ�IW#��g -<���7�jÄJ�?�R#G�hz4�4Q(HOY��oc "]�:v���)�@���Nâ@�t����Jq ����e5���(���]�s��Z�N�6lЯSR�~N��rY4'�^3ֱ�x��s,�.h�!du�RЛփ�و�\�Fm�͠�ϫ�L�In���%c�+yG�uנ�KǮw�*�ώ�A8�'�^~g��g�{i�
�4$����B��^���7��u��e(�=U��ζG�*� ���,����gb���{44(2y2�Q�WH)NP�Ž�aq�h�H]�ͳ����=�qO�p  �? �|��+��+(v߻�'j�2�k�T�� ����i���[-���S���^B�[e��zQo�RJH�v)�t����975� �d���S�A�;࣑�
�A�d��F�+H�_|� T����QV�2�|.Q��O��,sKY׌p'�3�	*����^��y}OR�[a|orW��
r�X^LbDBQ�<�[������uD�v��H�㳉�Xv��u�ie�;��Q����	�BH��H���u^��o���ԣ��ƿ���M7� c�XPV�
m!�H�~���AV]ӗx&,�Q������h}��y4;D<�00\����5��|`@!2n��g�����U��U%ﭤ	�Q��%�� ED�q4��ެ�6��v֬RK�N���C �~%8��s�?LA�Q�9타��C�	��u�&�}qP2��w��GQ	�1RCq����d���<׿ė8E�@���;�L���������-��K��;���A�Ci`2򙠨 �L��UYq'0����{�è^��G�2�[o�X�J%�W�D�=	�웋#�QW+�� �0���'m1���x����A_�哐���r�M��9���:�up�9*G�b�#��!aa
gn3� ���� .�]���U�~�+0P��@8F��P	����|L��ę6� (�� Tʏ��'�*�ԙ-vL���a)�{���8�J�%D:{�,�|���ТM)����&t�����9����e�~b@��I%�W��@�C7Q�����|Sr��6����~'��������Qs���(���aA�'p7��~�G�e�a��t���/����k8î>a�,@DE~[�"%� l��Ԍ�"߼a����v.�#��,�{�]ъY�}�: P"�v	^儬��.����&�؃����ڄ����Sh�@cM��P��apY8i��jsOf���%봜G�������Guo*>�pk���I��j5L[5�UA���.-7���!!A$��g�M
~����]��P��u	 X˕G~�PǪ�z_����C��:)!����J�w?`;Y�z2�=t#�_lT��gcDS�:T�2͊`9Di����_�RK��3����M'�p���[�^ѥP# P��"OAR�&
�X�!b�o}��+M�	��i�`�٧�/�bV$����D�G}��@`��s���4��etq��Z�ޘ�ue�F����R�wї��1�q	��$�U�d?����T*J�Y4a�Fv�t�zh�d��޷m��U���S]�й6�@~���� ��U�[%k�1�L�	z�5��y-��Yh����|��a�DbV씴鬁��_�$�=�f�@f�}��?/-^X�F�X/�P��"}�i�s�ޏ�Q��̇�;������Z����5�M0���^���Pu����G�7k�&�zn��\�0p��ϗG@�1��Y�r��2���4Կ�+��Ϻ�O��t~>7�S�����/,�$����(�P�M��K�P���d�j����J���V���YJ�8�~L��.���8���*ǰל� �5��$��R&�W!��T
$_pB���v�y�R��+mL�D4��8�-��dIz��=Rm�;X[��+��v�w��K�Z,�}�1�L����ο�j@��JI%�nE�����T"�!��9["F���W`�34D����X���@J�p|���J>����!����a�?%)��7|��g�U/�B�0"K�{�N�Βp�J�S��ˡɫI�U�P���`��ʲ*�)�	U7��LlM�u���&��}=ߢ��f,&[p�jo@�k�����気����h�%���t� �%2�[��X%��z3 !�c.��`|<���~�Sәj��S6=]j���w�sX87}��wOA�ߘ�Q����Ҡ���NRV[$�<��v.�`fu�Œ)]0�=�H$F
)�w��҅Ϳ�������!$�S.Y�Stmn���͵n&�DF���Mn�H4���_;�uRfhr.*�f*h�i5��;��o���o@[�b���؂F��<ד>��l��T{���&�ԥ����]��!D�=L����88	�p)��m\]�X��@�?��z���9k�>oC�!��B+FZ�Cġ��~ݹ���?�@sW��n6LS>��_n��1��O��Rbf�i��>�/�f����J�qR��KҁL]����̕�r>}�C�kރ� Ӹ��U�����9:w�5�2�D��O+��P�]� �`�-����p߯���`��'�Z��E�ȸ��WBP���j.d_��x�]4/��� q�/�]6�A�{X�=~�VgJ*.�#ǘ_� r�W���,�Bw}%����W�<�7l����-]Q%�|-2t���p��a#T���73�������k[>�;=*c�ǯ�X�e9P���P�?AKE��&OP�b ��'�WK,Guŕ�H�dI�]�x�%m^����d$3����6
��=j_I_��nR:��ֿӴ���-�Y�}M�C�@����}U
M4̩H�i�k��ܴ�`���V��1g�d;r��۾ܵ�|
f��#&��s1�T�^�\��C�Y� ѭ!&���)�>�WΏ�_�N�Y������u�����	� mq�(�7�:��kS8PO�$$����9�z��r˵�S�ׂ:�H�u�d�G��=b
g~�I�p+��w��2j��+V�	[�;A5/j��f��!����f�e@�!.Jv�c���q�nq/�i��."� ߖ�d��IQ�9Y�s�%d���Ea_�-ӳG._��8h����V�E�}���3�d�Z���Sߧw�錖�J.߼Q�����!Ow�
��:�wy�K��д}$����9L<���
5Wmj�vU{v>DT����q�w�^V!}?G��ܺF�g� {d�*JO�y��0I���	��M��ڐ���&kU0l�,�8�w�1�';��<5�ڊ��:������B?hK�s�\\[���Y�oI#�3�={��z%[���D�=���T�EF:m�
�P6���Q��k����.����1
<��)i�t��g��.���<Ҋ	��~��p�E���g���ٞȌƔ��D����X��=��NIX�.��S>���o��J�G���D3o����nn08@.�s�]X*$nV�_7@{,�Uҿeu@�Z��rc���
{�9]K ��s/-p���k�X<X
��W�n�u.���
9sQ���󰖲�y�cp|$�� ��&=�`��p��@�P�?V�&�y��,�?��w�O�������ޱ��Ω���7�`~߱��Qt����kbb!}][A��Yt�C���b��A�kt�{V��&���"���tB��w��: �����\@��(j�g)nL��o���sڭm�M��j�g��P<���EC�.wm���p�̥lҷp8�ދ�s�M��u��j6Ԗ"�s��ht�{pH1UW>�O�y�l��#J,qc��#�VS }r�%]lú�yu^��k�V.]����k��uΌC�(��Y.S��9	�i�
�h�YBAx��=�	���)d�!�
c��"Ņe� �����w
jPl����A�N>�|�ވy ��Qͥ�b>`�F��g�m��t;끧��ǂhXė�i���(n�(�dD�˓c��t� �K'Kt��R���{�,�jj~����\*{�N�������؄�O(���K�U���GG9~%m���T��`�P
睊�bk�l��8�<i/^��Q��|��,R���]����3C�Ak��կ!Bg8\(_��n �ecb��[�<
����L�] >�0GAc����ν���D�>* h}�\
��rAe�~FE�%>v3���(o�S)v԰C�����_C�k���� !ѝ����	M/(T�����	����00�B��.�f�X�"�꣡d{X�p�����W`�\��[GF�y5��0	�?q������[V�����m�����7��4�Z�(m�&vA!�KBzTT��z\LR;z��=*2���9M�k�l����J}��+��$VZsw+�RF����LE�*�o����&k�����=�eQ��q(mx�v�1?�i���!MQY��~^���ـ-���'I#R�sM��#�фy�-j��zt���ٖ��D�@E�ƒ.�q��W?�!��@q���+i\^������P���^O��E�']��Z�:g���1�*��< ���̹�@(3y�?���R�h�� \t��@m�F�9��r�T���9����C�P�B)��n!�|V��&�_x��g�E��3o�m����Qg�fϼFM���������6��0��lNك���iER�&����i�g0#j��Z�!}	kv���� �bpMa�c�|��L��T-�bd�����5���2�wbG�'�䥅�'��)� ���<�U�|�]S��Ia$<�N��3�JR�|P^�gA��	�ΐ:`ڊ�@���i�Mj�C��.͐Ǔ����@�$��Chr���#�U_O`�+żED�	ǐ�G$|и�s������&&��>�(��j�E �2K�7���.0��iC_�Ӂ[�a;��G��b�F9�w��T��;�jgǎ�͞(�����V�gJ෌�>�uZ2�������� ��*3&�J�)��l���Q�,@8*:d�h���B��.�k�.�Q��-���zi��9���"��/l�g��-�y}��#�Rf7[��s�#(�3^�H���{4��K8��\9�<�$�T'b�m�_٫P}�_�6zsI�iq���Y�F6�c����e�p��h�Y��"ڂ�$�������"b{	״h������7��E��q��DL��������e��O"�%$Y�}P��ָu��@�Nr���q�%Ynf��������#�wKU=�i�}�����X�b�C�$�}|d�<�^I��(�)��d뗒�I~ʧ#dD�e�#N��ë'��Z��W�Q[��gaX�Sb�.�iGJ0X�{X�_>4�s�Zbk%|Qc�+�]�p�s���Y�uj�^G2�밈�������㩱Tr�T�K=��yo!�wS��n��d����(|���ZW�����%=OѤ�"��ʶP&!\�{��	s�l�?�k�cc�+"2G	J_Iȅ��z���O�����g�UzJ����U��&�Y{#po� �HMՑ������C���I���NIud�GbX��9=���c֒����4�`��ڛ~�ltëh���ǹ�S��չ���n�*$v�9B��
A��G秅��L���m'�;����P@y卵aU ��-Awv�k��;�(}#W�t���l ��5� �����1�Z�ޤ"J�1�F8�׈�#�\�|�#fۨ�2�F�!�I?m�	a`�Y���O�E�뻆��<qdӳ��Ǖ�&�E<�N%1�� j�GT�D����޶�����&T��ґ��h�y,�^�%��	$��JZ��Fr{�2��7q�Ɗ�R�aՔ%5j���6�| ]r��Wu\��J�[��S�C<���2,FRɼ����a�5�j�vP@��%F*�=do�e�cA��/#�%S�����_��
C3�yM��ߢ�6���= G�(��Ed��D#��8o�?���j�v�x�Ό5��e�t�ٺ�G���
5�.��:���?����i΀]϶�JWjk�ʰ�Y�p��bV6�GC������"�р?Tg��;��~ �l^�^;`F�>��F!��͒��R�mv[�3L`%��M�2șD��bC|�\���$�Ȇ��[������V��-�ǮPGk
V $�'muhH6~
p,&��B�=`Ҟ��}j�����.��h��		�VY��(y����}����5����y@w�ڍ�W�~����.@�O�Ox��ŷ\��d�]�����4�r�����RGj��c����E4��)G��?m��,:o_�c,����z�Rq����P?��@Wɠ�(��l�SS��?Fu��)n������H��p�)�>�6�m���?��Ga�;�DE ; �^h9�rH$p8���ʐO�;~H��\E#���Ậ��w�����B,o�\�Td�~���$���Z���$��,^R$R��Vo�@[aŠ�4m|&��6O�6��\C2�f����E�М&f5:G[���SJ�=���(C�֑'l���a�3u q�Ȁ��&���4��d��\��F�EzY��f�,���y���Sx��$��/���tFT�Z�� QWZ[�u��4��Z�B��B�\ x�ژ�E�%��;%���i��{w��+'^X�g��"�N�>�-?�[�
u�o���J��z��^���0y_>@�ٍak��N�IZ�ֶ���Nx&�/�0��8��$8)Zf��0�Ĝ%u����1�����U�1%c�$�ܾ��A�hW�&�UJE�+�]M1+N���,�[���qʠP�@H���3h�Cd��Ҁ�Џ�|�E"��?r�{@�$h�3�	���8.W���� ��-~_�8[���������b{��� >!m.?�A:SD7�u���a��17�p9@=�����5R����=d+l��6�똩~��6zp-8�&_�j�l"�� ��6����טn޷�W��	�P���T��;����E "$����E<�����lk�5濏��O774B%8��X�n;d{�,Ohk�	�4��X=�2����]�C�C���L��$²�Ty%u�U��n�$�~Wh��h��w�ﰮa�)�P��c�"N~Zx���pHn8��T�M"z��݆�U���oY�rd�f�aQ!�+Յ��Iq��������`�]��Y�ȱ�W/3ߍ�&�lZ?�F�]�z=�^��w(�Y�6���۹X���=�D_�h��~de������е��<�v��e=O�_��id7����:Ir-o���a%�2�wA�I�,�+�RH����Y�}q����?2�+|{2`�A��5�6����c]2ww�`O�n�KkWV��`���:?lm☄Yj'�/F�p�֫�g���紒���m������o&��dC4��MD5*���<�g^x|�}�Z��C氀<��5�J����|��붜��~uŻ{)bC�)f)%���ˉA٩
����^Q4Ϗ�1S��A-lV�#⦩�^)�	n�l[�x�8�,;�,U�B
0>K���A����4K�z` :Ӳ�UMǘ�]������|�� *�2BI������O�P"��Z�ɽPF�jz7�è0��[U]6�"
�.>k3�F��6�/��)R;Y��?�%�-yJ�[��G:ؤ��N��mo��͌�� �-{.8b��=�&�S�u'B�)^#U�!��?'�i��	�QQg��&+��8���9GBÓ'�跸+@�'����]<��ͱ��Zy1C�#�q��]z��B��|`�D�=�eY��@w5VW΅*�?�a�Q���מca�N�����J�D�w�!/��s3�����v��YF�%l�-[�.\�.��C�
����`]�}+���t�^K3N�e1�h�{�*�Wiq�^��V<1��F�ROj�؀t��+�x�׉��dqt�.�şP�ق�K�ז��~����XR��g�&�J���z���9��A�9�p���B��ꁍ��^���qṔŁk��=Tml����\�Quc��Q��=���3�^�?t�>��O�|YZK�I��!�1�z�]
�ʅخ�_g֩D�ϳ�o~N��}T����i�O� ��ٜM�t��~|�nv���<�y��s#�+B��������� ��梠���u�s��b���ѽ4�ja���蹐�^�/z7�����I�m�ѵ��qE/�.f4K;>���K r��x5S�A̶�o�*���楤b�F=���18��HTx&l����*��+�����Gl��\�ŋYLLL|�/�!3�o2�ju7v �F���������i��Q�}u���q���vϕ�aQP�"?�w��]/�l����H��l��zxrpQ�7���a�V�L�&���u��k>�-�U�[(��Q��:�%)=����;�8U�K�|B�@Z�W=h��F�𐵢����7�m<5�����;^�D����?�<��Rd}ҕ�i3t@ |