��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^��,�~{�q�E��	YjpA������2o&�0���c�LڄX?�i��+�#��7J�n北�����J��kƧ�6���+{E�b��pڢ v�U��4��WL`d%�Zx�Һ�|�N2L�\����-�1s����#�+��l��"����1,h�'� ��a��I�k����^	w��G�Z��k(\H�9���# \����5AA�f��~o�ItMi������)Mn���e�4eӜ�^�����[)�F�0�?��~��w(-�f�sS��c��7����3��/��ֲm=o@=0�*QR��$�Ym*2�ծ>"�j��MZ�)є���8���'.��]����Ai��b$'�c�]7�a&���S���,�'1�O�U2�"�7�;@�医�.G��C^K�F]���_�3ϸsN���ј��`a3mWQ����UJ��|���9�~�4�3vf�b��aw��_��nm'M������-Z|��0,t�f��06D�@A&�[�\��Y��*H���闚�����D��z{���x�( �t� 3��ŮC]o�G��?�g�,�0so6]�h45��ZۥS>f@�0/+��e74�h�D �����D��������T�/�R �(J��CE'�b}	S�6��Ӷ�� t��@�1?KK<��]�b�@^���Z z8L/�0�`c�ER%Ƿn�ڵ���a
�o�g�;�Ql$�����>W�Z��4�\�
�#��� M�`��P�ǿ�R�`��)h|�FWJ�?2��+���yE�Lc��TR�~0�	B�-"�Hi�?D�����-�a���+���RXd2�0�p��A��m����cU�opVlO�9_3/���Qh�6�*r�ɒ�6���s�Z��^���k�EOo�������\|�M9�Un�yd����G�%��!�.bP+����V��S�IS�����:o��_AF�3݇��1:ʧ�cAd�l�`��%����6���4߹��*Ꭷ&�g�~�oJ�1���~�7�g�#��rOp?���J*��/��DNꔨй�p�j(���"���N.
`�3`���G�M�_��Qz#�l��B9�U���O�g$9��m����nwO��,�?�	�#�0q�c��g4�����z�a�H�o֫?�©���*m.�����/x¨��Q�c���}�9x`��y;�::ϱ�g8��<d���"Q^:�v�_�wJ�z�%�a�鯴0٠���ݻ����Q�;����¢Ys�[�o�:�{K���k���Qv1WF^?����ŉr:�����)6�8�$�,@�tyN�J��F%;~Ӵ˔qrY (�.�h�,�����$�!2�]䞹E�+y�}Ԑ�o��F�K�v�q�Q5��x1~�xѧ�7$cT%f����$�pc��㚯a�HF�P˜�?$sk�)�;��/�a����i�����~@_�Tr��f�4X\�}l�_4�*;�,�6�]����6	���8}�ơj���H����Z_�����i�$�g�;Y�~� ���蟭c�1�j��m�0��6���b�eʃ������NE��k�~�dC��F����%��:�@����{��O�9�d����<�(~n����7C�l����,A���.�lzb��Wa�5>i�i.��+V�[��V�zf���"�"���>����aP�x���P��/����u5l� ӾY^R8�������������7	�@�J�ùQ���p�+:YQ
�d��3Y��ɩ8~f�*����8R��ן�>͸N�V|�܎��E�tԿC�G~%?l�i2�Q���?
�Q�ו{�#�<R]��d��s�O5G���{�,(jSDGB�O7�jS?	��?r�5�D�oPq˯���?dǝ��}��z����9����!,�`�R�Ξ�إ�^_L�YS�d9�>>�
�:�������g��oקs�0���'ᷙ�X���R��J2�C�ޠhZ���Q5�5��*�r��.�kt��c��E�:P��, �n�vRO��XᛞX��3��N�alo]9$r@�:q�b���r�Z�9nE7�Y��h�n����|:�Γ� d"",��D�A����E�n����I�i�i/�+}�$9Z���Eg����H ޏ��ܯ��i-WN��[���h���n�cHw1Y��R�1�W@5$��__��7���S�n9�y��cBY+긋�>׏?�G��S�s��G͗+ή>+��+�=�-S� �;¸�Zu�9e{�/���� ��oc�2�7��ٷ©pK��${��K��U�?z�%�=5W��X������j6���O���~$.�S9��aJ�gɆ������5���(��`>�#ײE "~��rR��O�\�
�<h4E�`�wf�'뙢f�ٚʳ�&*B�8Ǻޝ]"�8�&��Ƭ/s�]���
Č��H��^��o���'J��L~�}�O$-����"�����w�ɟ�\��e
��o#x�a&��}�|$�B�@�c7�O�r�la��+���b�<?њ�[�j��n-ޢ�{x	�t[����k^�ӳet�r%��j�ͻ��ǯ0�+h7h�~�֜��M����