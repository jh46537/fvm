��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{MEi$ �:r������]	��+�N�L��+\?�w�hp��ۙV��<���>��2E���~,�3]DQ�8��3�z,���a8C�ʼÚ�?u���E���52d'�ȭؒ���R9}�"#���dC��nLu�2?�%�Hb� ���l�.��ܮP�ʘn����`'�X�R�D��;R��Rʜ��M�c��9�{ ��-T�o�����(���(��3.��հ���B�p:��&@�=��l2o��:ē�&y;�Ui��?'���1D��r���&��O�h��e�7L���� ��{�Mv��4�O�������}.�*���� �lH��@���5��	�rv<7ih����9:�֔:B�Z��_�_�����bn'b甥W���*�
�̽ X��&ԞJi��Sب񯇴DNM+H��a.p�7o*����G�	X}H&�{Zf�d��J8`���}�{���X��P_&�^p�{����U�
�C>�z/Z�>����y7�D;�#��k[5�XԺ�&V��ޣ7�gbBl/'�M��E�>�mt�-��i�6�5�5�b���~���+���<��1�Nj�|�+?���(����ϴ���� 6��I�8�uE���1#��0�(߉3�8�V�T| �+�x������(�D�]��;b�����ZF����ɵ�rk�Zc-�{�y�d�$���7i��P�L��e�m����X ���vS*��Z��%FI�! 䳳V,
$���6�Đ��Y^�~�-�q��oݰ��"d9o���Z�5$�[oG�~����_�����.0Ԫ	�z�p��s�jT�-�.%*����dU*UC�w��Q���iJ�#.�}Xr/@���Y�\ػ6o�!$�C�j6�*-�⋝��������A�G��h*=�^�Ѐ�ן=�͍�(�Iu�*,th؊������⿥��M�$A� ׎iIu3%c�%h� ".7�B�(���W����,�)%�����s�d�	��u�l��\���U$U��e���D�6�T��^'
�YĎ_%PQͤ^���0�Y#���2�pq��c y��;.�iYЉss-:���=�Q3��wk����qx>��E�M��zB*Z�����C�${"�����V�s+���A��D�.� `o������X��|pO��� � �zO6��T+9����`����\�ML�~a���*"��)ꕤ����i��&9��7>���j!.��ʹ�5 a��V.��ަ���T��-R���w��.U�!��;g�VC$��1�=K�{(�H^�mn�A�d�)������HZ���5eTx�,���[�em|x"t��V@o�,��L�җ�*�Z)���H�6�PUg��Yߙp�'�Ձ\N��z�76ZAÇ�����@l�ε^=���]���lH���]�_yCˮ{	����U��t}�4�&�$��@�Qל�a"C��{��N�;��0܊/f�����u~����]�%�%�-� k|ɩ�Ϥ7��5�%N��7g��x��Dv�n?�a��Χ�K�Ç�����>���On��cG}�?8�n�������lk������n�'31B��:רb��k��b̗���a8C�>���P��S	^6OM�,�72�����o�~`��Y��OĮ8^r-$~s�+b��v�藐�ȉ������Nk�"L�"\�q��ɂE_�	DK�y��Ī�'Mk(Eo
y��򁊗&[-��m�DE8��+w�4��S������d�E�<�����d`�/��T���ݔ����O�Ad>����h<��&���34���awpt]�qC����&X�L0�\}��iGx�v!�LsG��Ȕ�m�E�����:��V^T���$�@:�k�{��bl��D'L6�Mz-��`&��p��U���BLDz��H�Y�f\�a`�XK�d ���?��5��#
?AL�2�y@9Lr�m{:yc�8�;�ۨ�J*D�����T�9�]�T)�'�[)�>}UMD��'S���q0"\��5!t3Z�Sw�^08%u8t2�^�Mc�� m\����f�� �~j�zY���2T<��wٖ>�/M�z�Ekߎo�Y
�b��|�כ��:9��