��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c����}����ٛ�!"!�lvVS׿mi.�
NO�4ʣ�k@�0�A�����d��%����g��g��/����
�>�l�@��YST7f�
�W:�f.��<|<�(9��(>ʴ��o��q!V��l�z���!'
�j�3��Z� ��Z��*��n��De̤�%��vK���'�9���U��k��(;�0H����
��8>�by�U$8B�z���I;R��Z#g�%��b�L�vE���
5HI��+��S�<�0�ݗ$����D�˂��];��|���;�P4�1��ݤ�tқ>�c����p�=&��>U���S/IJ9 ��s�k<Y��mk�O�	%��純c�g��[��5��ȡOM�
�������Ơ�zɸO9NƄ߮)��o�
���d	x�$��EN���e���s�B��\{�;%A���<&vz���F����tH7�ɬҷ�`�����
���n>����(
��Y6��J���媪 ���=�qs���0��9
V�D�*t9�M�6m.�[t�^s�)h�7j���θ�`�E�� �B�鈩�#ٖ�9!�ƍZ�:�J/'�v�P��d��H�e�7��dA��a�^�LH����^s˷�к�f/��0�!�cb��mo
��]i���� ��n}�탇?|M�������M^2�#���avf:S�_��3P����=���qL��������-X��X?�2�
���r���O��tA�.���<��q�jW�Ȓ�|3��|��u�����96!�Jv��Ё�%0)=,�Q��Rh���&�3,�ѿeW��L�臡(�a9$x�_ e��"�P�[��LBC��V��`���bJ)0&�Ѩ����jЬ�i��N��^���D���p�Ú_��z~�Z2���`�w�l����z?)�J�l��h��0��z���*�i���e<�e����٭[v|Z��9_�6`2�.��P�Z�HQң]��5� ���?bڛ�L�Պx�ǪM�9����
1��86���&��A�u����h��ohӪp}�z��T��iY�����_�S� }�R�6f���G#Tt8��UO�U�B�MŔ,~�\V1&Q�����!�2aʉ�dPu%{�f%]��l�N���Y5�q&f��mR�w7��յ���N��/�N+s|w�?�䴒3�Z��7,���-=V\�z�,PVˢ�Scq]C��>�ߣ�N�8g�Ʒ��q�������P�yjr��G_qD	�	�� 2����td���90Ϯ](`!��4o�S���2��Zү
Z:���{�t?\vpD��dg��M��/s��"�Ѷ����e$N��TM0�|Є1t�ΰV�EC7���z��-�e!�s�Q�����.�:6��U�i�*m�Y��\o�kct���h��Q�t|!��3σmf���Hq#1�HM>.���aj��YabP�N#��UfW����JZ��`�#�i
�����]�� ���tH��gf�2�G��C�Z�SH����v������p�{��fZ�v��D�x$�|��H��*�
��Z�5֣g���Z��_z(�.���W�@��Q�qlɭ����_�*�"l����>��Sҙ��� q��Ig��$!�a	�|T�z���Ϳ�)	�������3�	� �Fф�����ط4}�q�XtG._��ue�hV
�ט��cO������h]���W����,�A��ǋvb'^5�S�[`6�`��a|�)��[�'�	��Ď�'�ar����ܮt�B��x2n��Fr�V���?74s(	��ǐ����7.��eW=ڴ�ɍ����k\�i��j8b�nAd��Às\�>�Jp����M�=T�i:;���K�kpi������F�<T">�Ő+��A���-����q�&O?T�$ Mi��48�e�¥�P��r�$�*��O���q�r;%d�&�c���s�\���;�@���U:�d������K,��(�e�И�M��8�5�ڐ�l����ywD52�c'm�@���n+��]W��b*ٍ����;���(f��;��k���-�1uğҹIó��\��W�G�����5�F��I����|� �`��{���Ow8�;%�"�C��&�����KÆ��g���o>'ݑ ���?KF��G�va� ��L��'C���޶�j<}�S�*��jK�� |�-�?"�c�r�d2\�K��ЛN\�0\C�9���������e�V���ߎ��!�NaL��e]��h&�)UD�y��� ���!<nM�r,�!�����E��@�V��ꩼ'�9��}��%*|�UDv�#qe�[g�1T�w���,�hV���>7���
��y��M, |o�r�Ч
����n�s��q��E���O���!�@R��~�����i��B��)!!�4DS��\��+�}���ST���*xz/��%`U��sN.EF��k������X�H+�
2�9f�'�M/xϫ�31 +q�\g�0x-���1O�O����9U|t���;c��m�[n=$P���EmLf��l�.������}���1�P5���2�HF�Œ2f���TW�񲂕Q�&r�������;�î��=��[i���,	����J�]N�݆��� (?�c�܃*c���BÕw�aQ��\�P�i<Ե���������?��&�ǟ(���N��^�l��,oo�(��O�b�D�?%���b~r|�	��*A=��5;Otx���HIN��m�̊�����X�;9�A����'��@�!�7q���&�Ɂ��� ܔƌ��۞�� ��%$7h"x4����Rej�E�b|�e��
IĠΊ�0p�_0��&�@X��*>���\U��_�3��Kӂ�ӣ�a��C�"��o�]}�����E$�^~�N��y���b0�(�7%
�&ĩ�cf����dKN�;���un�	�:�~��*���U��@���fJ�~8@B�`Z�!�y&���42����8�Ǘ@6�8�����μ�g��n��t������<����U���0��G 9�k-/ElӘ�~R�7㏘|I�M�	�\��qU�?�0+Ͽ����iGu8Z��o%-�D��yK�&!�γg�����Ef:����Ď�;C�M�`��kԖ�1���7;� Z��|�44Λ-��$�kz=��"+ ���-RgX���9>R���"�#����g�g(�_1��_5�p���w�l~��T8~�(�fe
x`��o����`��r;�bjRE���:��|R]�?��a��܅o��^a�Җ�����r��M�Aqq#"����E=��'$�?/Ȁ��*��!���I�o�	��	 �.T�?��X���>��;igᩣ��#e%>����ѵ٧ei�[�Zc�D�}h}�h'��\��}��iC���X�rs2��$FoM�/>�$��`�j��l��퉌����P�W�v51O.�8m�@�tᦪ)~�#M�n�Z)'�gJ��.�m�a)��FZ�K~;q�Y6��K���u%4��:�'�3����d��zi����v!���0�^�ڮ�
	���'ՉE���+UDI5��U�� 2�	Y�[?8����Bk;�T�A�DWݹ�A�T�	��jbl�4��Y�"d� �Y9�ַ�#ц�[���0�=OLl�p�p2�,
��+�*y��3��Bߖ�3�T�d}���U\�i��[�1�n��f���e���>�m�4k��s�SE�#}�U�@<`�	x�xs>�>���lی��8q��,,ٓ��9�Nш�$6s}�9�k���X=#����:I�?��z�(Ӱ��tj��z*�<���ݮ&J��8`�����^X��pv}��9�B��m��|�v���7»6UB�2��	
��K�HN�]�"ړ�U��ՠ߅�jI`���M%1R+�B�;_���NJQE������^���kO\W#l�����0��,�'�� <`���)d����L�y��&�2	�gFFz�P�b���u~�k�3[��j�Q��z�ϼ�p���G��s�|z?�+�j%�y�'�ĕ{�6��2nBL�f�r3��<:����xG%�blQ���.�aΕ��7Qo�3V�\�d7Kc�Z����6|=���rA�3M4���~����0o��;]Lw]�	Z��g38)[���;��$&4a3%�Hޥ��+"�����qл߽�'a�*��8�gRS��rv=�L���Y�k)%�~�>PC�8i��B�������M���6O�����;m���i��/�İ�yݳ� �2���Am�w�l���U
k�OI�p�s�}�DR��2iY��w�XB�{'gO#����~m-G~}���l��-����-��u�������I�{�������E�	�����w���۱��<���'w��¯;��S���"9r����aQ�Ѵ���󉹈ݡȧ�툘��\Ƿ���2`�J��ip�����ґ�Em�Pvlh��|<��BE5إ_��#/�i�������m��bn��D�Ʒ$��w�b@�w\9�e��>B��`�c��R���~kX"ΐ�Tژ&�A$z�BF�ݍON|�J D�G�@��B�o�߃�UH���"[-Ȋ���� |�JҬ-V ��ϊZcJ�Sb��J�!UԸ�����P_���҈Ϗz�rؾG�b����>���e�B
��Y�<}d�9�%��\R/���H\�_B�\��V�`�$J(|���p$�c����l՚�Yb�M^�d-�5�7e=�~�������p�"	a�Q&�Y�),(h��]���f�MWEFF(Q�g0{��6�����M���3������%�Vb���%�	å���r�T$>�h�]��U�6f��BFB;�>]6`|a1��s9���5�A���5��_�@-s"ǂz���X��:�El�A�xȢ*u��j����~��߷��n��Ā�h��v��I#eR��A���^���N�Ao��F��t8m���n�TPFL0�⽃���W�?H�E,���.��c�o�XA�5�}9�$O9R�d�T��q�Dw����ש:�ZX���\�iR��