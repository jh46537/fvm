��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,�������_^�6�3�@�RU:(�3�ݵ���_��+Z�&ژI{�-��*����=cM�G�* K�M��;ȩk7�d�9?Qj�뻞[Ur/�Y�MG���^DQ��-�`u6O)�A ��r>{����UW�EG���i��ay�ݽ�� �F%bW��6J��5&D�:�P=�w���е�}�r�I�v<�-�$�>�����d���`��&��k�ӈI��0������T��S�!�x
y�_���5־ўX��
 ��7v�+}BC]�FV
��g���G��S*�d�,q�f4��2����b�t>&������Pf��tzY�@)�(�p[;JN�uؑ)���E�<.y��_�ǻ̘���Ԏ�0�
�,g�Mb�<c�w1Y�4�
���Y�`�L�~��
�ᬅ5͵C�?ZVHh͜�s
�w�q�BF�޶M�:w�N��I��z؉ NDK���^�������~��������
�3n.;�Z���b��
�:	����7(�Ϸ�b5��=��ƸT��7)T�<� ��轛��>ZW��`��y`~��ܫ�"�jPQ�
�w_�W/��ɬ��.ǭ�ۻ�d
�d��%�q&��{z*�8ȷܺ/q��{��:�*����sGl0x����\��D}0�kj���mq&�1NZ^��*���	p���� ��&���W�p��x����w�5�G3�(&O*:,%�e�^����GH�V�A8�	�,SO�C4�Z���z��E���1�Tgzۉ���P����a��
	t��8��ߙy���5�B�g'�~lj9�� *�S[�ƎP�T�n��$���@�4������t96��G�ڥ;P�#D>U9�`�?Y`�A*}�L���W�e.w&�#���j�"���"7�<�O;��̇����vK+��cb���x��c�!�h	b�_��}a�Z�mzH��mu�c�[��]'i,�V�]��t��H�yF5[ �㧗����9�xFf_Yh#pJ�ޑ�F&6����������G4��2Ɨ��iLE�=r�)�r�;S�R�͐�#x8�Q��-�����C�g��S���)8�	0\{���̦[��(��bW9�\��3S[PC�~���XҬ�_tϫ�z|\�C���(g�Jw��e�>�6����D�p�u�'Ts�뿮s� �uS,�2
Hq�5zX��ƺ����[,f��q�G�K��#���P�ɝ����M�p#$�+t���~;|F}�u�^>�ّu63��q��1�+���̡#;����@o�i�"�i�J���?��Q���?Q&�������<)Q��Yn2y �1����<ۉ'��cs4�9?_�UO0�ۮ�ܾCYTΕ& 2�h�.J���^�9n�����|��vm�C�*y���m�o�˷�7C�Eq9�ǎqP����V�7�����^F�ے9�{%"E�:>��\����Xk@Kp����TA�d�c��������J�����<1E	�i5���Œ�`�R柲vL"o{��;�m�������&\��ZcC�gpk�n�:^Zg �%�M�a�"�.�ol����Ԃ�0�^xϷ���Z�� _0Z'/Jf��b{����Q��z49�[ ��S����ǏA�;
�:���iF���Ȃ��B��7SO�@Y�*X+Y���gƧ���%�GO(kԭKt���إ��U&�bӵ�$�������9�����ϔ�l{+���sJ'���r�h�A3�6�B�]�#uݴ�2�x�I-��3ba�d`�c*I��^T�>Mٜ�!(�������#���e�ZS	c���%'\F� $4�~�rgCbMnv��Ly�/��1f*O�E�mDܯ�işߊz,��=��O��a��#T�Q�+f�������}���l�4޼��ͅK׸F�l�z����,�X��Vo/����p|Pt4F���F�W ��ҋ���B����=� ;�Y��a��1K=�E !��cI�[��ۼ�`B�n�\�]�h�S0�.*����b֙���<V~q�����=L���|1U��j�M$T����$kMU9��0���w|�S�N�NX�h��,�؍��Hl� �[ۼW܊��OR��w�D��I\3�9��
H.���mw"H�Ѓ��7�Ef|/R^�نh�gXu��< �/D0�k��n��K���O9ڛ
$�Q������eiv_����^�jep]�Ò���]����(�Qd\�`��B�F4z��j 
��2��� �%�9+�K^����FV����I"�+H�Y��-j�>ijx:�]`Y�*�����DC�=c'����*Tm�4#�-
h�i'������ͩm��3�T�;Q��`��{(�P�ɷ�u��%oy��@(fލ�q-H���s3�BGT���Z7mq*eb������#?\~77�pv�)N邏ˍ��n0x9yi�cv�:@�Q�/)sZC	9K�Yc,�K��ø�	�)�!�6���X�ƽ����3�?��-l�vXC���l$/�9)����k���b��@�ږo ����2g��_�Fbm����1v��amP��R���$��^{�g�^�7���(ѹ^�3j���z^98�������c0���OR-��T?�Y�Gg/ۤ别34��fhWE�o���T�7�_�Xx(���|6@�\���ćk\���ȹ-��B	��Z1g�Y�l"K�R�.�׮��j1M��]L��ÓK�����xG��^|�P�H��q)�D2VO��~�����V�e���v��4I�U�U�Shn�z�U�D��o!̈́��Te��I��ˈ�<�Ee�� BUG�ί��g�l�@-�Cd��b51�ub񯈍���0���g���R�#}.?w�s#e1H0�hT�gF~�=���RőlfvI�>y{U��-s*-�����	(�5b,P�3��&	o���V��ˇV� =��g)�a�QD:�?��M�\TfbZ���p߆�/kG��!� �Y)������/ݥ��u&�k���,�K������@u���2�G���&�0�1�d��2�X��翅ha3G�X�muWHY��*V�\���l�]E�(�"S8t5����&��=Σ��)��������	���tB�3�x����������64l
�:�,�cqb�-"��euF��O����y��#�l�.W���!���Z��8��n��������7@b��y��{Ӛ׺�FRNM#:(�����/��[�=5���]g�z������n�2ư�x�'ٲtP��`���R���M&��T}�,�?rr��$�4�s���;cɦGǩ�����"TM֢���UyL���fA���r�Ft�"�Iu���Q�C�T,u�.T��ٱ֭��ۏN��:��Ӛ�]���K�I�c�j�^�Z
�M��I~�ɚN3�TF���8-�l��@��N\�p�~���"�ĲX��ZM��E_��m��/�Dd>�5���O ���j�{-}��z�/����q�>�Pka�M�"� �7�݅R�;M��k��i�����l�V��$j�w����6�9��Ab�ԍ�V��х����iu��� +n�N��G{@��������f�	�&��;���6�R�IVL�'��{��T�/ٸ�żw����V8�?Z4RSը��IX�.F�M1��7f�O�M���'2|�1�Rw 8Vnb�Hh XK��/)~�Q0`
�A2��E5����=���2?�(����d("rsB�2G��ԓב���=؜{9ҹ���o+,�#b(,#�8: m7 aT��bD��O7giE�\,��|��/�mk�}fF�ߓ�#��aG~�oֱ7�̾��l�n��Q6Ѻ������eljG��v�dV`��w�B�z���'B4wA������T�V�[XnݛY~� -��YԤ�1U{��6qtmQ�� ��a��h�:V�=pێl깁O���t�%�����o���P�:���c4�E3!'���Y�Yi&�`��;����v)�/��x������,��)8�lndyFs�t"�l�����J���BN���i�e�{� \�4w�O�kK��iUt��:+�2&Ȅ'����z��&����-;�Ț.��~�6�;�E����W۸��΍��n��X�.��&�^U��	�k5
�N�(��ڭ�����/cQ8�Dth�\��h��fvs�2iۮ� v�p��4��?��!�!�o ��b�Q��) &A}5��d�G���"��� ��	਼����v��Tg�W��x�^D�u��Wd��K����P�H�e�R��\9ۨ47��Yn���ϒ|��{|F�A�t�h�a�m�j�_����p��-8O��0�	7N�R!�v�-��.a�w��΁Z��}�MC�����X��SZ;w��� �8�m�%5I)���AC�+��5��|����%��I_�Gg�8ూ$��C�%�E�:gh�T�R2���4�h��錿��/�(lQ��51̻W	0��1N���`I���/f�cِ��$��� ��A�E_H?��iV���?��؋�ձ�vn�LaBrm�͗dK�SW��M2�����;��u��h�n��zz����kVɬ"�g���TC���s�7�c<q��^�}	��� 7,�)T	�4`��c~9~܇u$񗹖�7��3��`�-�߅��Y���QKD�w�F��У�j�QP`Utq���q��2���h�V�,4ϛ%�)�{�g�m���i2�ێ��`pO�ڞ�h�����x�B�Ԉ��xw���lU�\��lUu�޵�_��UnT��0b�[���`ݫ��\#��^�;D��o§\�!#' q�{���� �Xm5dW�s5�	Q�kQ*<�P�f#������l«���c�!��tg��O5�������_�y4�L�kJ�E�P����P��.��k�Xua�m��ڳIGU��{�*�R�3��J�i�xs�X���zd���I|��N���gf���xI���q�gt�V� �^+��� z�M�g5wDX�FKWeo�ݲ���3~�� e��(��V��LFFd�y�[��nR>�&�����UkF�I��'���A�h3��H��]��Έ��9����z;�e,_1����$ȟ B���Ty^7Y���x[�Oqi��a�G�Ȕ���I��s�Ԉ<fZ/�h��B���5*�����p�R��,��G�B�%��~HiZ�u��J�z|K �Q��Ʈ.c�=��д��<Ǽ��u�h�@�ʐޥ�Wa���֤��j�A��F�`u��>.{l�O��D�݃k��u��i�tߪsJI��X�S������CZ���`}����֍6#��^�0Bŧw�����]ц,5dh���/��Q2�!��u�c�E�3��E fR��z�ۺK��j��������d�S����ƍ�+�mf:-��(��Om����$�])�mMfaT���_H��gj��^\�.�ɮϸ�ƿbKB� :��\�q�9"&���������[隈��T7�5���"�#Y��ŀ�����1��=�[�$&̴o"�h�4���Jjv/;ÃC�W�Rx�։�|YCO��5De��;V�(PzsػD9��리��Z�pڼ4#87����{�6y���Ș8���\�c��>��p]͠�`=5o����>Z'ٸu(��,A��%�l�>�֝��X���(x�Ο|���n
= N� v�����h�(;�6HV	�\�B��80�m2x|�-��L�@o'Ҟo%�Ɛ����B��
�W�#���[hP���$'~�gS�8�9.����qW{P��U7�_~�d��S�wZ�)�/�P�
,�]�	����W,`ˢ�̴�"{%"x,8w�*�0���1"]�@�QW����0��U��vXL8�
N����mP��H��1?���z�7�!���~�᧌���D�O�H�1]�#ȳ���CR�2��O��b��6.1��"��ꁼXn=
����ۆ���<�+�A��9�u���`X�d�`C�g§y
*l~d�����b��xs��
���j@p�������i�c}�\zU��{���uj���w_Uq�	�%.h��X�%g�H��)��.ܨr��8N֫]���g�+�(�� ���@�D!O~)�2�9g��pP
(����#�)��M����E>�e wt-3��d��-�@���`4+oF�cO"�1Q|L?���<��q��ΰ��J��7�����+g���#9���Bb(!� ^_����Q���)q+Bm�g��!�@�*���9�1���!��N/1�h�������f���\xu�����^� ��
.0�+r^H��1�E�8�d�ML �>���)�L��/
�, ?�;|A�.} $�H���#����$	������lJ}�k�V�=�f��ջ`����Z���;��n��#�vz
��1��`K�MVsE�w��yY���������to���[�m]��{�$쀜�R'�i��f�`)k�\wk��)j���<���h�O� �@���&�*���\��}9/7_F��遇�`JIS����ї���46$G�DQ�O3{�U;�ET���B�.�P�uy�J�.�����ߕ�]+��Ӂ5��ѳ�%N�R�aC�X���}�������9>;�֌M��!.��$s���5�Hh��F�=J�wcTFU����` Or%\"��&���r'J�	�y[m*���^�.��fȯ�럹s{<�g��B�nQ]Q3���^��}�~�5���A�F��
���\����Jq�@^�D)D/8a$�F��P����?�<)�M�H�W��+ȅ�Fz@7�o�|oᯫ{�>�$(�=��*�m��Liɠ)��U�H�SU�p�(b�}.R,��\P"�k���7�y���1=3-�Fa�P/f�c�l��z����*\}U�]N��rw�*fB�� �N^���Gu�(<~5N�KXx�|3Y��"	xٺ]����ѥ��?&�6T82��q�Af�t���$q�Έ3 �̥$Y��,���T�D����kگq;�CX�a�������`	E:-��\aE�ܗ�̖ �,�J/���`跪.г�V;=�� [��9�:���ᨈyے�`N�l�N����m���;,�~��1��0,�e���9�Q?V�)���q)𳒬D��fF:l`Q�g��B�֙�B�����).�#"s��y�O�I5��f�(�F��B��g�T�tí�q7���oh��T�^�oh.�|��2��АPf�h�P�~L�a�j�&�*,tl������F$�vA�s�uA	�*ݼ��SY�n=�>G��Ҁ�J^:�H+JÕ_��c�CF�3�Y�9���(O�!Z�A�������"��e�Ug�z�9J�[��r_H[��a��?RZU7��V�]�d����x���ۈ�M&~-��jP�ج1�[�8�T�҈+�\�d�h����YM}	��s~�+j��N+��0AF�R�}f�׵4p� d��[o	Q�&۴��.|-nI{c4�;�g'�`1HzO��l�Sb���R�����O=�@xc�m�3��Dy]�׻��x)�f�w%��$p��~x�����U!�Q�Nbg����WYin{M/p���7[أ�j�j�x��b�Q���ǉ��N�y��k=��ar���2���j�`t�na��7�$���T=$Q�����L��U�S�1e4T�[jWcnᯔ�B�L݉���7;ݣ%Z}B�,a��U�A�������>���J_V7��*�7��':L�JO��=���qt�_���?(�U͠��*6�Igʉ��9f�=R���-��M���M�w����x�[ݶ<��ß��J��B�G�1��ϱ}�E�zf\�:���APG(;�{QW�b9�`u�7!:�H�eIh[�5��?N�!�������XG"����P'�7��0��7� ^e>� ,w�]��^3:�%��6F�J���憒y��GSA�-�=�l�Z~K��Z��W�x-�Kv�!��Ce38�v��G��n���ɾ��J�"��e���տ'Mv?�P��(X�|��~v�Sc�Z�ڟ��Z�Y�I�v�z[���-�L��81�d���c)� �<p�>���v(`��n�Nv����̒�An���Zb]Ɓ̱�d�iD�F���H�OX�-�4�[d^>�9���F$�L|��2����W׳���v����L�'�23����V����Z7�WHD��0�2W�8;J�-��˻M�M$�3� ߲Bvj�8;�/o�p��� �aC��K�$�.N�������J;�%�*�E�SS�1��)h�|�{"��١�$�t�q����9����L	p��@��H����8�JE ��H�+�������8~�H6��2�n�y2Q�sW�#$��42!,r#��D��2���O؂�?��T��\�7*w�䔈���s ?�;߸d���o����e�}��*\�����#����	��uQ���fub��v���Y�#ޠ`bNș�@n$�����S?�w��%�؇��E���b*g
՟�<�\�%�)l�@�htv���$zԪ��>{jy��uؐ,`��[�@\Z�|y�j.r��c����!;���ek�E$�(��f4�˯�K�%���60�=2c�cz�t�u=֋��vz�b���u���'r�5�?����{�n��@���V��ҟe�W'�\�j�U�'��t�/�5|Ic]4������Cw��R&���a�Cgv%l!s�O��@]�_
㜁I�y[) V�W�-fI�;��c(zؐ`a�6dz�p��*��Q�[�b5��Ւe`ׁ�o$��ΘK�d��v�l��6��izрS���,x~��x.�����<6�����C�j��H��Rn���ӏoG6�(ԍ�!�W8�1G��)�5��/3�W+�B�n2z����$��b��Q���Ӈ���>y���@w�����7:&��Vi����bq�U��Z@�DԎ�	�8����*-I���8+?��+
D[z�u�9��0
��`i�����$���Z���ᜮzQ�83�ǖ���@��G0��7�t��5�!�p��̔'4�$��,G���䥻S�oR�2�`#�����zb�zӛ�6�jw0�fdoG���T��i��f��;����~MԏHe
��9k����5-	�Q�U_�.�L7?D�X �@���o��8�ڜbF0k�|q�U�2u��X�����J�kt�x%�0��Y��+�f�h3J�8u�E�k�^�d8�L�aQ�����A3زޱ����/db�^�Y�`�S~�6��దKoL\�L<r��j�5�1�@���M�n��{R�����W��J�Б�Z���g=�?ȕu?���֙V�����Q�g�=����~�+`�[��:ʕ8�S[���|����	}&����4�D}��Kt�_��YR~�U�L�t�1B�V�oXi̷�y�U^��#��Qb|+�.�3J̏���ִ�r��mrPt�z����,�
�^��7q��WV���F���[�6��ؼNǍ�pʂ�?��7A�����p�����]~dޮ5�i��٤�.H'�2��X3���w E��HpA
�C}��3��s_(wk*J!w��w���6t������I�tDD���r_�:�%7��@��j{"C�b������b�5И�9�(�X��.���B+���=R��8���&� �	LJv���X$�w�?�]�=)N �3!�ZEܤ`�3R[�!�n��*��)���\��Q7q:�������̷k�h�y�dL�ײ ��;�2�e�(2ɹ�7�O��Y���K��A6�0��&v�t�[i�s��i��t�_���c�J!��"g���Jμ��f��o�wr�.|���dPguJ�b��1��9����,�������� ,`C���}�I������M9�
9(�3���N�uB'KJ�q<ZG����p�A>*X��0X����^+�zь!���o���-*�a�k�?o��Ҭ:�4nBn��Ng��t�þ�4����JI�H@�f�C�J�`	�AT�4kH����)�f���������H����֙Q�y��P@mZ�d�gܜ3	�xr�Fv-j!ub`��D7V+��*o��VMf~�xbA���Jl��hz�2l�D���(��]�b��+~�����f��ď��1����l�e�|��������*L�W�fJ�~�%���Rά1Y�n�:���)8,�*����Y̛����ta?͔����T����F*y��+��,��̀� ���<F{�1��A�i�@����%��%��Fߗ낸����%j;����}i{�����9�j�f