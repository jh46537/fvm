��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�=���,1�jӛXT�d݂��V�k
��&sq��s�Ԁ��8�N�r(x�xI�\�jw�.v8&k����sqXk .*g�1�,��΄:~��춟4"}gjj�	�D&�*�;��tlj��8��9M��h�"��u;�p�r�뢺)��6s� ���c��hO�1�s4p���!��|D�㈴��d���/�6����)G8�����fAHm[�?ME �c��VPG��]v]��=]0�*o��1WE&%��Y��;��MΛ�p��X���Y����T�m)�t��a��a���66��s�F�1��M�S�[k7�ٔs��$�\��Z��kV��������*��y0�7����-��d�)�� R�!�`dS�����}�,�C�:��%����Tb�� p�B�D�`z@�i�dZ�b3��'x��
_�`��+���f��9���w��о�R����U�@8�1SVĿ�4J�GĊ�]9��Lǭ��r�4?�2J��IRQ�3?wԘ�C^}0���r�r[3n%��Mz��+(X�^��>?:��oc��޷�(r�ǂP"Z^��������v�CW�E�#�\3������@�C�+Z�<zcn0��ԭ9f2/,��(��d�&��k�G�w�1��B�G���N���*hR���L����i���Du�~�U�
-ȇgO�ki?$���)��#7������+w�'b7\=��i��>?z�S���H~*?͹L��hk����~���a�FX�{b?G�6B@�Q�_��k^�<7�{�hj��L�W� ��B��P�C���l�(G��:�|�պ�Kd"�ΰH�� �b!<���΀�R�RZZ�ؖ�̠,�6�>,r7W����y��9f�G�K�4S�(W
�^9[7�!�6��P?)k��b��X��z���S��t]/_!��G�6�O��w؈o>�î��mi��8ڽ!0���L-���mK�Q���y~.m�ׂ�3��u���+@'���W|̔a	�{�&�����B)޽`�]��,�|�jх�i�;p==T ��F��O��I��-j�Ĕ&��HK7��Z.���at:�ٛ��;��g_K�?�\��GtA7 ���	4�}N�$��������en�Jv�W49��..���ׇ�X�2�/��#(,�%?��A*���̆���:���Ym������5�_� /� :�>�V�Y�4S`�� sk�VY�"�=�t!����$q��<��d?J��B|���������@�=�!�w�:�}��"[�:Dt������.���821��f��2�?���&R�iPl_ �@t�6<�����x$g\��e�2X|�B����1X��kZ��Z7�w5JD'�޻Go>#�Q�G����X�h��! ή�W�D�2i�9�2KyI-��9n[�{e�.��HRZ=Aר`�� �0[����u�6�u��r�5�UJ���~�!���^E�m^W�S�����VHC�P<x@1�\);ٻZ皣\q8 �4xތ���-ԍ%e���N}��G�,�e�Hb�Sw\�9��uǚ��������-����w4b����,��0!��[�{MK�
��{�k>�?�
�����֡���1�w���[!L�ƮI��{��	���d�8��g�6荃��g����߫��*�x���
`S�������Oపq��(����k��8����X����?!����J�t����9@��&�)�*W9�:Ya�Y_��Cb���$�Αa��M*�-*>�+h2�E�-}�f���*�)MIX��Ԡ��Ֆ~��\~��9�.�x�F�?ӯ�D�W��BA(+�Ί*�Á�AҬ�d�D>VP��>���mN�p�KI�$;��?���`rӉ���U�$�9�u�O�M�DV4�D� �$����]?�aZ(��Gf2�5�"�PhP�c�����e~�JB�#�Y���XB%P#a�6�'�®En�	B((G+H����^l�K�
2w�t��h}�C\��\��c+p���R�nwΉ��u�~������;�5�A��lbw�&a�2Y8Z(Ũ�_>Y0#�!�N�9Q[Ó��+ʇT0�yE�8�zy���ب�a9f2�xI{#+r��V��:`0�:�A�A��B��vM8&�f�����E�y��7C!"��'j>���`����5CcM~�����L��?���NN������V�>����)I�$�Q�Ηt����I�6�&� !YNq5���
��/*xPM͊H,Z�&��t�FH�>(u��K�`���X�1T�?�����5'!2���� ��ޜ��� N���
�O�x@Ɖ���´ j���?�j�����O4V;o�\��AP�â����E�.�v������q������>D���b9��\�P�^K��Yź����>�)��7@_'EA������R�en�U�����Rv�51c��S���y�?����`F'w�R�]����k�IW��b掸8�}����6^+��f0�=���Ǳ��3W�(��j�A6U� V���0q�NW��C}�a�;6���O��)���ₒ⢡�$��-�7�uj�"A�6dyhedR �L;���)��K����aj�&��AR7�:��C0��6t���bQ�.i�:����ɏ�7�"��@Ke
�(q[]Z�@���e�2���q�Q��V�	��_.���kqs����?�ӵ;��x��I��.��Jt~not]Ȃ3�)VZM����||N$�+# �կ5�[�{�&�a2|��<����YU��&�n�%wsɕ�_�X� p�c_���L�ﻰ�l�x��~HIoAN�����W�W?Q��7��'�!�U�v�8�A&�7Nk(�h��(�$������jq���*�ص�2��4N��Z4Ӕ Cy�U���x������`8��[��A?`���,M�	- sP�_38�ͱ7=��w�B0^T[�/�&�f[�iK��"ǅ@"���øK�M����/#��磆���"�~��K���Oa�jR\P:����V�y2��ߝ�߯!85̆bT.W����&zB��Y�]�ͤ�7z���/�;�gM��R��j�)Ƀ��
.s�Ϩ��\��0���(2d�~��B���9$�!�`���Đ>q���4G��r�|em�Ӆ��(y�`�R��d�u�VU&˗�w�����:)7`�.T@�����K�X�c���ʕ�sjd�����`���=�nB�188&4�
q<�A�Y���,(碴�9�aq�EI���.��U5��f+<Q�))�������7��zӿ2�x��x�6Z����S�2��feԷ���¼����#����}�{�k��N���倦*k�Ba�	ܡ�^	A�������1�7�T�y�����F���*P��6�Ĭ��	����5�0����yn�ԡd�j�ߍ��
Q�!�Lu����ű��Ry�iV�B�b����O���O�l'�9)$"?~��M�V���L���<��D���c%]7���p鱡�L9�s�\����+��f�0y�1%)��F�D�L�M�YG ����[��#U7 �k�;hf��7k<bC�\6/bem���n�
|ۀ.��R�3�À�ӜRܸ�%�Hs<�GU��}��Ϝ���bg���_��<�'Enyv!8=(f^q��-�QIy.�`�R�Խ�.���Yf�@�h�w��D�ԝ0tS|ȏ���]H}K��^a@�
E���x�ZałSD*�1��^ۄT�ѫ�4c�r�z6���A��R8&����k;���*���8n�lf�)3 f�~����v��	�~^_��h�d� �
�8�Wj,�S�[u,��\�s�v�c�2�y�V2#v�N��/>g�7E�	�s��s�-�Ԟ���̼O� F!�¢���$��U�J�h�bg�cRP�B�H�z�!ݽ�f��oJ��>�>s��*������䠰(�Z��o���^�[Z=���]���ե�ж� ^n��8���v��X�j�DAM��]��3�Lq~�] g����/Z�4�'h�)TcIa�L ך��uK��h���D�]5��)8�g�y��TG/��������(
7��F:ST��f��"�lv�09C��LK�=����F�v'1��5�f����.@�&1we�/�ݵJk���W�$��p}���^�iAE�����;l��Lf��?����Xj���@d�$)�`�V'c��Y�]��cjg�G�&��a�~'�B3���SDg) �gO�N�%���:h-X�1��Wm����Oa�C��s=����+���мQs�ɧ�u�#V"�${t�tޓQ3W�Բ��k�%��V������W�>���~Nё6c�{)R��6M��L(��$G�>im��Ox[���
{UA� /���A�������`��dM�e9�NQ��,ƭ�.��	a�,�����k�=��m��t���{��H!:�s�2T�	����ς��qܼhmԴ̇4��N~�pԪ�^���"r]u���V����3���h��m⚤�.�3g60�Y�g�7s;��Ql��A�B{X�X%������������
�*� nx��_5$�{
B~��X��?���6؄�����aOu���J�Wh2���9�/Zɢ
�D�Q�ˌ�X����W�T��0�3�aa�EJ����v���FT��K�+�üɞ&� �=�>|��FI�C�DeGP~Z��d���	O��^B*�q�;�yB!h�,�"��Ql�&��?��I(/�8���!�}?L�JI>��G��٫;~��h�^��t�v=���u~\W�2&�M�֛Bs��'Ѩ��~1�A��b���7��L��X٨ڷ�>7��NnC݃��x�r�	+0��T�y�+�%o���4��S�t!��h0B����7X��ǣ�#N&���A�z�pI��e[��Y�!ܪ(\�}��#(ڟ��q