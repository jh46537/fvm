��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7]�s��^TC#�yM�g,�%kڅHе6��&E��1M�?��z���bkk'ɝ'�y#�O?��A��,�ޛ�t�B�7O�e0;L	I嬔���=�\]"��]{��~�ĵ�����SOUAEo�s<tnj�I��vj���Q¯�$��I��q��o�6�͋u>t��-\���g��n����B����{1V�У�S;���#��k4'�	�(�WA�wU-�}�nH��\S�kr{֦u��&>�-v���]A,����c�BꠟV�$[�Zi~\�b�H��w�ג[$��T�TQ;�F\X2�#3H��ɮ�8p?������؈ٳ<T���+� ���M�%	Q��:�^����;�p��^4��u
Y^���9��0Ԇ�M�yeg�	1<W����G[�T�w�IR�d���W�L�o���H����iK{b��3ߧ����t�^�9�.�p�!�+m��������a����� O�Mٔ�m��t�{�7��]Ű�օhK���/�f���ߓXh��;�|�Q����v�׉�^���(�l��f�*ۓ�h�}7fe�ܽ���Q�G�Y}��O�=�l��ξ��D�?�2�C���:�yo�/�,ީ� �Uy��J��Zh�'$�� ���Y[^��M�j@��]r�&��}nP�k{�sƦ�V��b7K{~���+�����q@d�M�i@�+�^L�U���~�_$J�rc�ϴI�ʈ��]!���.J�b��O]�$f�~+D��Q:�4��|��H�SZ^��`���R�e2
���a��7f�������9�Զ��^+�+6�<�kp0��w�� �w������w��"�e�8���ǐ�`f��O�u���E�)�`�&�
�O��
7�8�H ͢Sn��1���aY�ь[����iWG�EQ0�C�(�l�G3�tۀ����l�1��m�O}���wيV<�f��q��%�����F�����3E��RR?�JKwy�*$�e�h� "�6Z����[\��ߧ�N��ά�ޭ�+�^������ST�p���Dś��%��]�`����ȸ���I.�����P�Z����8�ȏ!�/�=*&�cs[���bVհ&� �lMX%dI�I�ϰ�Φ{�o#��C�z�b�_
tF7�[3x\Gy�psĜN�n�`Hl,���3+�VcmM:\p���d�b�B���.l�Ͻ0F>�ϸs��O�Q�< ���[���dp~o��(�W��L���&������P��. Z�Y�Q �'v��[I$l�}����_d�r����n�Я�4��哉��vJy�8�d�쏍�7ez{�a�k�N˰Δ����Q)�נe������2- .X�EP��۳!L�n��1}'k�mY!\��_�3=�{9�~f��K��?�]��y��	W�4���W$�V�Q�2��x�ZM�:�i�AΓ����2_}���#���(�ТV�5\�[���V�=�{t�!���Ѐ��A�m�$����0�J����{sKM{5%֗�{��-�C�ny�71茡��tSll�R��!� K�#鄛E�'jq�Z/��˗����ݻ�ȍ4��MQZ4�]_ �M��@�V�Cx�=f�P�p.����|�͚C[{�Ǭ���Un[�?B���v�н"��_���Sd��>Z��]�.�=Bo	����?:B�����y��Zanv���霯����m2��~�To� �"�n
}��j������p��0��!���`��6澲7�J��l�J��%9ux�O�~�VK+�O�\�X-9�n�q��t�g�4���X���Xln3���[���X��3|�Θ���s��~����ֶ;�����S/P��(�@��l]^`�;�����hIPU�Yc]2�!5z����IZԵ�����R/!kԓ�ݟ��Kl���F�-�d��o���33���ܤ��Q�|lF��֕��D��3�`�����P"N�x�S5"e����bP�h�~<BC	��-�g�`+�����et�s<�%� ��g!
h���R�'@����|�>�-D�m/dTu��?ϣ�W	@�)�G��O֙Q���d��A�a>mb�ک~�� �E�ϱB$	lT��1��7��$�_� e��U��"�d�2>[(-+ ��@���ͭ�A��8��U+I�J����������*b�Q/rn��D��Kb���>��p�M� �\P�}ȱe\
��ׁ�'	�2~3���6c̥�����$������� m-c��
u��G��x���]eD���;$e�p�2�,%��DAe˟�KP�N����MO�p!��l�s����K"0�t/�ޫ�Wh�V1�cH+��v1���lAoc�b� Pz6�+g����J~�X������� ��6p�١���z<�i8{���o�:��m�it����E��(����������\-�x��ar��%���S�}�ݎ��6CE��Ȍ����r� �z��#�/٫���t���\=t?��K/��E��������A�,o�f���eQ*�F�d�A=���=�2Ou��{B�J1�H�a�x5�7����Zl3�
|ݠ%�S�τ߮5o�D{Nb{g����D�����<Yޠ�ɒ��ø�ْDiORR0�,"�U,@��x��YJ�'~��'��:�R0�`�1ã�<��970��D�S�?m��n��9O��ݐo�bk슭�����
��d1� �WE(���D~����M	���b�%�,y[��,�4�5�8�U$����wV�f�o��&�Ѿ#�;�uf��Dt�9�7記�>;���=XQ��&��-Y]0*��K�@N��8�9~��G�ԭ��rz�*�ܹ�_5B6N�#L�6�?[�����#��N���$��[і��t�Hۋg��$$������]�&��4U��M��.��}o}�a�U�X���X����Ծ9s	�_.�`��|Ǡ�W����ٗ�pmx_�t����ʲƠT��&��,��ԜS��}��>R�k��&�Wzp#d������D/�o��6��<,+��ԡ�I�pe] 2Ls7K�����<[	��e��(Q���X$�²5e��s��$��k;͘HJ���xϑ�b�rH(�*��=$��hǾH�CЫbT[�>N�d�p�f?��ɒU��{�SBL���Ksb�$dq�A�;�U�V�w� �y(�}�u�xg����F�߅?��[�.���
��n�Њ)m�&�:�֛�l�8w3n+Ӳ=TƂ�,�� ��T��{N�4P�+�`#Tʀ6@đP�|������$�P�9*�S�Zfnm��|��`#c1{�m�H7���~�����I�@�wA��gÉ�@����V�$z`|�e���h����nd�cW�2�~Ǔ>{]�*P� S7��Yn��WP�P��%��k}S�l����	:�kE�y��l8�4�A�%�x>}���Rݴ�������ʩ(���//��Zz����\��� ��%�G�&el{�`�`C''��<%��-PA��p�گ�$x�(V*Wr�ڲ��Q��N�z���9��0�0}��4��zp1K"��? ���]`� �4I Uo��IÒ�N���\G�ͳ�]@��ut�:�b�D�eL��	��E���*�P�VRT���7��}�^��ب�`�NǼAd$�7T*�b��^k��Tq1ŉ�ߐS�{�(o���Gz�H��o�8UGn�������.��m���[Y-A�!n50
�g��
ڵ}�21DVpf�s6�	zv��]M���	�ߙ�I��Yȩ�ER��%,�uz��r:�	����;$�-&Ĕq�r���H�= Ĝ��BN��v�q��1�&tWp�2}�L��a�u`$�1TL0�<��'��hE���AV@� $1��B�|�r]÷��1S1�	���=��E�M�K,e�j���8Q*�A�)��Ӽ�*�t�4��V�aQ-)�lwFD�D�ux�Y�*T����0&[ ,�ѝ�������7M��u��dI{=�N9�y}��e�`����!���1��O��M�rz�Ul�����>QJn土��7�!w��ǳqס2	�`VE3/�>���To-��k�R��"t(xa^c_C�Y{�q��#��	�C�����O�0Go�w+��'�F,��՘ș�<܉��q�
%n���o�"ʣ����{�m7?D)�s���+V�GVj���F���M�u���a�-:8B�>�5{�S�0&tE2�n8����E�R�86��6p=�� 5I�_��'�~�����:���%�_ke��H�n(��1cه�Y���L�Ec΢��^�Ҡ �� J��x:�>�ϩ�� ^�]�j'�m�K�m��/�3��Ģ��3얈��+����J�XO6.}�Փ���ʶܡ��+��AH�\��#{�CL�ؒ��U"�(��|U��7n�[�������A+�\��kޚ �_���H��NBL�c��oM������A�=�&�88�u�jnV}��v�ݠ�]63~^�a����dJ�	��ATR��K�@^�_B&�>;��H����?�䱜��&�A��uy�D�����'ϖ�s,���09y�A��9��3�:����$������� �}�J������'�y����O�Y��#��{���z���ъ�ҕ�/�F=썐���!�M%�,��YEk��c�L�9��U�����+G+G��=���Z#�H"��^�Tؒ�t?j����0s�-���>L�}��ä́�C���#��F��
7����\
�oer����N��ފ��#1
b�Ҁ�M�=�]�K����R�T�����z͈��a�Š7�0�7vKJ�����^K��D����1�~��)�ܯs�Q�ܗ���G-h~{��0�v�Ʉ$Ջ:� �
�X��ɮ��_�k�f(E��m-�VMJ��/@MT�7��ԞM������I�r
B��A��O�F?���N͏5���#%i?i�a���������ܓ�q"�x1��ʩPi�T�ZϫC�� 	�=uW��ӘڮfV���d�$�"Z�y�Y��
}G�6