��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw���Q5��x㛼9������6���*|7��?��1� $���"R� 6���*�p�+s��s����k��Y��?�:���1���O�^N}3L�qE5%�Bw��h@�6q`�_�9�y�\��z?��nf�h̅�1[��- w�0��PS���`�S���O,�H���@�����l����Y@��n29���U�����2������ߍ*'��6�z��;$�T���� �B*�$炨��龈XN�g���A=�b�x�b[�	|I|y�� ��:��UH̆��kW/r������&6T��EY�C��{>7*�,�u��.Z��0j�=m�	Xg�*�_�}<An�4..��-|p!�3&T���oj	׺c����zvĄ��\W�΢�R�%�}���8���'�p�)rO�$g��In�>���Y�3S���?M�U�(g����(�\Af�GE���0���6��v�;�p&�����#R=�D@�l���h�j����}N.Xj�c�)<F��x����C���6�j���ZKffE}���S��%�Q<!�t2��&#�|/,!�l;/�ej_�H�����{���v�^U;���nD>z�]�w8����8�1�VL�1�#WWP���^y�.9.Փ��?��݃����J^ �)�W���H���b���e��T�3�R\ ��։�[!⓺ge4}�L<�����uv=!��P)�4��iZ����YN+kG �>�u	Ľ�m��W���wF���XX�%����T��z]��նWx�-2^��/�Tʀ��!� cc�ì�C�c�Rf�j�)VlF-���.ӡRJ�zDU�y�͸�c�rDC[��tdf�e����@$6�b*m���,��;�GDa4�I��)��h����2f��փ�F��� �1=����`���"��VL�4ɲ,��#�f�ixz��a�;qEkϧUC����q��B��W�v���
J���P'������K�zn�āZ�5c�|?���2��3���܉n"����#���Y��_�
j��t�����������־��z�*@M]�����j��D6��_/�P�<,���5s�P'<w"G̍έ��[%��,,1�/� �P�^���}��os�5b����4Ի��2�V����Q���g����D�:���Gt�,�*�t�f�3Q?���|M����W}X�<�	4���DR	5����*��tZ!�&�7�3W���x�cӞצ3�-�gY��H���cT�J�ʛ���&���O��n�(�j���� {�d���\8@��`"U�?KPu\��(�;�uOΘuƟ���[W�'��$�'wtU�AT����P���%ﯲ-�T��NE�����ۏ2��K��-�LU�w}�m�D�N�P)��J��������B�0�ʉ�"��6�F����[�����̱�<@������6g��'`�O�M���'L�2M��E��9f�b��D��A�����"��M�	�P=�ǚ"X�1���}� .�"���ٺ�����z] �Cp�Q�[ƫ�I[���R���h��$�9s�4h0B�]po����,�{�ugFe��J	Ii�/LjKL�k�����ڗ���sbUFU�l�Y��ʏԊhB��?�w�����!�J�9���/�9�!7�4�����s��n������z������;*��z�NYN[)��*��ԟ��T��z5��>��&[!�U�3����P��[d,V�Z``@ke;tEŏ�ˆEF��uk�Ͱ�x��x����3��[F�!��ެ'���p뫇�F���1�)`��$G9-S��M��f�d�����l�>Y�������O��TV�	]S֘���a8�N`d�r���bAsn��V��,�P����\�C)�V)>��=���1�`=�Ӝ��𐹙x6��*G�:S�bT��F��;m�V�J
S����!�e?��֕y��	��W��!j6��B�{/�xdJD��]S�'Y��r��Ƚ4멽S�WW��-����Z��[f\-��7���4�v4u�ٿv��r6����s�}|`�,��e"4�f�n����NҶ�⃯�W��rQ]b2f�g��-e�<��MD��5�O�i��7H�U$�˽��C���%�H-�,fL�C����!LZ�R�[�Za�i2��t=��E1��U_�0�u����,狯ji�~�9�`D��Y��M[�eL=(z�Uy�O:npfr
��?.��1uB�ǓY��TJ����B�� 9�X���sq��TG�@��7'?���sxѩZ>ų۲V6ί���^�ۙ�����k¢77��.9����u+u�<L� ��� �LñY�H1�ؿ���6��[�SG¢0r���\im�RÅ��ٻ���i=����!4�o-G�`(`������O,�G�{<���3 ,���_3���RZk�MR����?M��V��%n���**��C� ��I���Pv�j�E�����o�Z��TX�ݵ(p�\Rf�{X���1�����N���UZn���'����I�?�I�y\̡>#��M���4Co��cUA�`<�+<]�T��\,ȍ��	9����\�w	h��D��Qõj�*}����pprX	��b{����|��!��/�dX�bsD��S�#q�M�n�U���g��G���E��?�r����rC�[���)����t�o��f�z�g_~s+Qyɒ�>�M#w��9���~��B��q�q����3~a�ċ�J7vg�H�]�m=	%�<���5���3��N�
l/�{�.�>_؋U��rv�P�
�:��ѕ��Baiq��ԣ]��W���!���i.�Z1X�G��r6}t�����Ӱ�M���c�w�E�.�Pٰ��L��s�LH��o	�'4﫼Q��I�!��@�?yu�"������!���LtWS�qע�B{���ٞ��Ν���ٲ�Dl�U�A��B�ym��u�H�~���l�j��P��i,��Zs�ѢvGo�!Jާ�=�A�9����n5�̈S�>�y3~j�:->�B.�	l����s�y�[�4��/��'M�}]���*U1J�5��)-ӊh{� 0֮�I7T����u���#����R��Y��y�3^�H!�� �: �����!���&�㹴�
)#����l���X~.�t3��� ��V�wh��I�pѱ#�9���R�:y�UG`�{$I���m�����N_�v��@	���n
�-3Cq�����ew�^PP3;.;��V|±§���K��VK�ZQuF`]�������G���i�#��m�#��P�N����ԞS���"�(���`'n�Wz*&��N����$��
O�obݑ��uqT���}�qooR5��\�!Y00h(ڭ�54�K7%W�ؔ���kɶ�-cuM�pt�y/�:!�~��������R�Tc���j{c})"b��vvר�����W�9�Du��٬���^�~@K�+Y^�����+�kQO��]3B��jy�1��k�w3?�o� \[S�k�5�jf9�޺:�;�T"�	��7����2rStز;l��	�����55�#j�R ̨�Eu�eO����'"��~�Ȇ��`#�4d�\��"m���I���@�	���
�'�}B�0I���L�2��'�"!AD���O�~��3�Ȟ9+��W`��B�RR,��Q}�N"��<N����Ya�N�8�����2�+zE��0B����\83��ڕ1�k�Z#�@��L\y�n�Su7&{�5N0Gl��!K�p[�h]�2]��q��:<)_Lk���w;��¥{,�ᯤ�+�0��B��]�>�+����M�M<�=B�'}Z"�ߙhO�R��*D�n>��|'>�y�?�k��NB�
V�M�L��H^�D	�A�Y�>Ж��@�9��Ɯ��f9���Ǽ����+�Vu�_�@!p{�'e]�R�Ą6���I��B����`%	kE�"�Rx�O����R����w�=3�v��	���V�W��\"���R�7��O��HE���ۇ�����oL���g����dW�fg1�6�w�o�����_��1�a�5�uQ�1�;�Ǣn��7���O�����������&���� x@У�D�$Z��V.	a�6�D��v��@����q��.���:'�61�e7����� Q�z��quʭ3�Y��;݊�U:ƽ{�S��F�����ÚAs�yc�<�|��§!$L�7�FQ#�b���2qX����c�؎4:��>:v_YD4�5S��``މ����V���z��ߝ�� Y��,�2��	m5�
�@�E��)*1|�ǌ�1�(ؿ`���N���� N�v�F�jkF��7օ��p��y~���A}���{$�'n[�G7ZvI�1>�����iFz�\���2�T��=��'��^c��A6AJ?�hx�Z1����?�n*b�ڶ��?稲[١XԐz"d�-�s��xDfH���S!�W*ǋ��-JH���B$�h)��+}wd�^�c#��iE��Y�����R&d�'wi��5���yr�����Q1�NI
�����Gg�l,^7l�[�>����7�M�R?��I��{9��!��P�>�kŎm��̘���e�_P&,��+��H��
 %�4AW�Z�%C��F��ċ���D#*Z��5�"�
�!������娗�>��oC��/�uC���������5��ߞ.C�Y��.3�����:h�{��#�O?	�dh.e2��@=6*��G��m�8�����A� ����!�Ƕ8D��C<�4
�)���/]�d��]��Ňk�}�����mK�#:"�4#��0Kڴ��ѐ����{�u�{Д�)�O�O�|y��
�d�9��;���RPˢ����_n�}PR�Y�hc����m�1+���eǴv��Gvtb~�g�'C}�	 ضag�p�ڼI璶j(^�^ȕ`Q�y�q��Z�(�{"U6$�F������g"����1w��R�)�g���D!y��"AtC���������&��G��LP����.}c������ͯ�0����i.r�����R�Vv7��L�?�����Odr� \��ѹp��*s�]�#��$��[*�
U"B�D��T&џE�u��$P}�c�_��"� �E��4r���~1�Ƙ
��2V�6���n�s�l���<ς�3-������QU�Ls�{���np+�� d�`^�ϊ��3����<��c�n��3�썫!����;�'��v�����;�=�D���)���ݲ��'2�znO���)>-F�CS��5���E�EX�F�#]����$�q�i�T�Ȭ'�s�M5��
�x'��F��WkL�sp^��f,b�"�p[�ީr�=�y�qާp{Q�
���%}TsRI^�5�x�2�m@^��q,�B���s���%�=f�����?t�8����P�b��gJ��&�����uw�7D@��g�D&�����-�۾�34�M�#w������������^�49CnOѾy��"S��^d*��A VFQe3VLūE��RY�p�|^���%��es��_��_�փ6Kq"5��+o��߳�͛X�����ד��|]�Ƒ�%a�bV~<�i�e!'2��{4���5+�@�V��O�de�M2 Ͳ���NĒ�&��<��v����
�7�ߛ\}��"�Q��yb������J�\V��V0�_L����v��j�� �p�/��X"�9�&��5$�51�Hdj�i���gZ����ߓL�^�)�2�2�s��2:qi`"��I��c
�=>]�4��0����.H��z�i�PЂ,�{1є�uAi�6�j������x7;�/�yc���;z(:����W!���JP����J���Y(�yw��H�R4����^���-���p�����z���ŝEjْO(�� "Coh� "E����D�̗��r�E�Պ�[����r�m�J��c���!=�ڻU9��:����,��汇�l�+7|�����'���u�mg��&^��|�Pң�l8�M�ZW6�����@1 �Oݴ4�e��b�xՐ��x��b���ý0~�<�o� ��Cm�w)��>Γ�"�e=��$�%���H�CtU�L�Q�ڥ>��]� e���"ۆ�p�f��ԇ��=���C	���6�.�!��	�as���bU�2�7���/��c+�PH���m<�����PzV+�+S&����h��о�2sƴ�����V\~��o�dבHu�}ύ����B��TMC�Q�4X�7X�k7�cՙv0J�6�|��&�t�^y��;O�s��p��z�}�r@P>��K4���h���c��oʨ��\��9�́���T~d:]5|J�?c�A��&�����(�������8�[����P�(�,Ǯ"CٚVGsZU��*Z�.s�!�"_J�>)/���TP,���Xm��W�(\�������ч�~�(C�/���*`��؁��(̌ϊ�7�e�x�Ƹ�>�t=�LH8����mԱ��;�'�=�x�q��y���(am�w)6�S��<��OHʣ:@�%r�j����V.�-��;qC�����i�Y��}c.=��PP�4�^.� �BK�'Q�k���[��Tn�=k%��<�L���r Hoa���xzQܤ�[G�T�KKR�G�,s��9�hig� ����m�B��!!]tI¯����/�o9|�r�ER@z+��I�,� �k�t��`�'&�s���`W5O���_�c�T�ge���?�Y���m�ܐCY�QH��ī55Pہ��|R@����YQ�z�!�|l@\�>�Jq�;���3q�Dff�N�{ChO�<������ 3�u^;�f_uj�8Kmk�֝�N�����t�`�֖;��e%�w0� z�7��}=��ܴ�UYFO�Y~�ٍ13G����,�t��N�`��5�`�Ƅ��o��X�	 ��L~T���$�E��%��U�;O��G�G�"��!=��Xr��M�{t��
�!?S�0���,Ƴ�l�żȔSDg� A=����b>��%���e�.�ĺ�#g#���>w��dc2l���c6шv�δ|��������(�ECA���c�+,�sY��	Pa�U"��"p��[;�ty���K�~�"��F��W��[�G3��v��� g� �ω=С�$|�n�������Y���*1��C���y��eҴ�k�:oI�}��Q�;� �����yH.�s�XM��a^J�1�[S�e�\"��x��>����@�E��b�5�!�%��8��쮃�F���l�Z�S0$���ذ�&� ���(�Զ��1��<�t�@�a���Å�����lܥ����4:YTn�غ9�q:�ርnS��EU?0�A�CE�h�~����|3D���h�&�}��>�<�'h���y%��'e`w�!�i�{�އ6N����b���zp���&7�'75�.k6�!���L٠���d{P���>���B�mTj�}��|`���D��憱��n� #�m���:&yW]�f�<���YO��l;����~"��8b�s���p �[��[#O�C�yh��l���<ov�ʱ��۱�Ɨ�H�\-`&Z*N�fŸ��TJ���a���y���Z�!�M'Q6�Ha��+�����E����
��K�df���D��B���B�I��$�Db�ǿ����0> ^��\����.e������jw�O�}@"��^��Un�n������ΡԠ.�p2K%�;\�t9�D�0g�s��RծL��ca��UZ=\����Y��F�$ `ӥ�CVs�kp�I��0i�p�UB�����a�!@���K��⢼��\(�&���b��$�Jf94Ϩ��*bHA��yb��@������'�� �E���%�g�麌�+��EA��3�92�Uw�s�u�ҟy����W����E>5U�M+_ۑk5��Dr��~≰�u-Q�1�i<C�`�1��"{�BTΐ��oF�=k(���gz�&8�t	���ʹ��$7�+�L���@~s�x��Yv��H���n�tG�#���v4M��Sz�@CX��R���b�q�ǲ��6<;��'�C��N!�k1W�'�X�R\��?>=.!$C7n�� ���fy�j��և
��u��D��}��v�"��ϓdؕ	D���Qph���r�S���8�F#��0.�Y�ـ���IBQ:a-�.?�ٻ�p?��:8	h���Rb�&f\��1U ��{O�c6�V�P��P�7�njo��殜��r.�,�9n������o@��#�"������[���Y��W%�$�|��ba?��k��>�C�^᭢�5�j!h �%V*r�,�Ka�"���\x,�� ���c���Լq�j{a���: W���mo�F%'A6�#��u�ԗ�+ܶ����ِ찃��){��&lJ�+i�HK�.�Y��T=���F#0̼xY1�ı��<�,����*MS�c�����I���b��=�U)�BOQ�]�2�3�|��oGh@��U�79y#�c��#��o�x��ʮ�6@ɸF���b�^- ,M�"v5�@�#�ؿYk�m:�l����#��]ŗǂ�-_��yI���^��+��;����1�>����6k�Ā�~��!|�=v�1����8��[�(�C��BՏ�߲�bnV$�����Q�=��'�}��F෗b]��@�n[=�:]�B
s����7��I���y>0���%2��ޘ4;z_��,'��Cq�z;!��#�����~b��~R�q��u�+
�cL��{21˳$��&{��l>yZ*���A�H��O����h=�-�����bAC�d�-�?���0^�>����G����9�x�ѵ-<�Cx���E����Pd�����7�p�z��]�M�k������'�ǢLG?�j5��}�r+��"�0/` �ۺq���4�~	���⹇����YE�w��H�-�{����:W�W��PVɕ�-H��+�:�QS(�oӑB���ͫG�M����sArzOaO=b��{��]�x���rD�Β��"B/A&O���,����p��P�G7{�jp5��[�B�I��XC��Ԓ"��� B���1t����L8���	��4H����9	:K���	k�b�ow�vʹ�{ژ�B��3RH�whN��k��ہ`�ꎏ�X1ӯ�p���w���L`N/��z\%����3�V.3}��*���4���r�&��Ƨ��|6�W �~zM?������|v�R ���q����G�ȩ⌥�sˆ�.'5���;���f}ě�FӉ0P5�����)J���G����py �R0UF�ӵ���v��Y��S ��-����V ݝ���4=&*��f���ir�����U�%��a���h%4A��	�/��ʺo�틐n�ͥ��{.O�?��',3Q��.�!,�D�Z��)����+x�.}�N��`��t�Y���>�ݦ�Ln�HI�^��;�[C��6�`��J*�^���_R�^�=F��bM�J��P�w*λD�2���YTN\o��'C��Y�0(�+��vf�I>��q�J��2tF��'][%#���-�2H�R�����n+ ��X>�X�H��O�N�f9����!�P���u C������)lf�@]�;��S����/V�ʏ��](BӠU��f�f�H7S��3��k�e6���B�}�~Ƹ������Ql (�`8�`���%�z�^��y��tmN�j����"�q��8J֞�#b����gy$A��۝hv��(�]9>�&�ϱ��c�[�Qa���L��1V�=b��=<�bv��);_�]+<o'TK�O�$�c�쀡�KOLJ�Fb��Y���}+�e�적�\8	2]S�90LJ��No]�_֒��Z+�:�D�ƕ[���"D��ZW鉾��[u'>�_�=���	��J^� ��{���� 9�	'�mO�/�tW�R��E�w6�z<�l��T5অ���oۃTt��Cj��IP�	�]�\^��r9�ʦ�,������7�g�H�_���7WKe��0qN�c>�*�2o��̡:k~�zgy�%&
,�9��+Q�>�]�܅'��P
�nҋ\� � ��k(;����8�vc:@�1��� ���u��ۨ;f�ө?��F����J*��{ ���Ry�w"�z�C�2u������Ɛg��ٷ$��B^��:d�Q�l����ò��X��d�����=�z��2��y��cz��;b�����&�����S�5�P\����t��{�_�[+Ai^ԍ����B��8��Ke/J�e���V^�<���?�4�!�a�3�`D����ݖ�9���9�&����˓��hf��6����		�wu>Y�5q�+E�w�K�0��+�J/x���"��N��) ��sm�m�`u:�����ST���o�(Ķ�~�N�!ߡ��Dg��%$yk8j�z���i�����<�`�(�����A�ˀz�GU��c����`➱�r����jѧ�;�x'/,�@��4�Zr[�L�C�u���N$�8�U�{�G�L��O����A��;�6VOP�$�t�w�\��ؽ4�Ur=e�N�~Ͼ�n�������ͰX;%�സľ����>"mkDNd{�)��b�N�ف/<5̶<��{��� }c����/�*��\(j��(XA��*&��#���M�/����#�H�t�� 6�������F� J !'י�g���D<(`��<"���R���@1�^��_�0���{�W^If���Q��굣����X^�bd�[(����'h5'5��~\��\0`�My-mkG�XP�e{^�vU_� ��
�">Y�ע�B"A435'��*/�d�29Vu���b���22n���U�-b*;>r���FdM������+y;����@� �o�C��
���ޭ��A ,�lKZC6r͊y)���s1&F޳h�k%0�p����yQ�ܚ�I�y�s&>�5�֚�����ĭA}Z�Q����r���������A!�M�Rs]�JH9��}��r��P�Wy�DL��!PHy"�K�̤�R��g��؛XB�cS�b2�$�,���䯟��Cr{���:����R�p餳����
a���%mf*��7�` �*������!/�^�M��d��b,Q�zqrn���x'y�*N�����I��	cD��qE�{婾.�|/��� ���I���i��<%TָK���[�9�� .�o�z"%�壛LQ�'3Z7�|��H�{�V���,��?PA]HP@���v�bϕw_�Z�*B�O����⿎��K���\K�}���6 #$�vH鶺R|16���|ED��� ���d;�R�m+��6����V��f�U1VAB�H�%@��*� ��f��,�W����Hd����q���4�R�y��LH�z�O�-��j7�-0�����?("��ă�G��zE0��ź��'��|�`O��(�{�Fr��YtY�G�F9 ��m"������a��s�=R������}�+r��
�Zc��~[s�v�W VO�v-Ì��v�2�L�
-v��v)���T˥����g֡A���SQ
UϟN��U��
�;,�-Ҷ��}���4���`��!��>G�i��!��O6��^
�;D��o%a�,���Wa��X&Jy�ইH�m�eō��W_�Jb��Z
g�l��#��a�8xu�D�Z���	�M�ݵ�
�+HY�M�$3BVX6���Z�R�f���_���/0��<O�l�^1d��ʰ$N(ӷ!�B�{l�0�0� %3�U�g��������A_&,�qҡ;���z����g[/ڔ|�cQ�vj�
3.ˉp
���T�� ��j�m�`T��Z`���π�{���&�����W�@N�"�䕩~�o�@�l�=�aȲ	q��̺�/w�}7���Ӊ�iښ�xj��2������su�K��=&0~��<>� ���q�+!/��y�(,�Л;�g�!0'wj��vPV�;����:Db�㺋q����kNP�s��x�!�}��[�GH=�I�2ߕ&	Ji���o�Wp�r��H��~�J��������ڊg�:�ֆ>M[(��=��*�vN�ں�(K����H���D�B��]�7r	h���=�q�� �*!�n^&�� �4Lr�U�H>ѷ>Ď�M�~v�J l�Ldy��n�,��~��3 _mÐ�-�_^e���P��fm��)-�k�p�p[�P��6��Oۊ�W7���!�`йI���Z���k��+�k��"_�w'��:� ����e4ʋ-& �JFxPh�9v=������	Z��w�$/��g!�݋5g&/Z����q�ԩs�]?h]��AR$m�΁X7���|�hLM,�H�Z�:�5�Z�7���*����<Fqd�$҃��ۦ���EHl�jC�������wz�E�&�5���̉fQ�8-�����i/���S�9�R0%��+��N�3"�0=�+l����Y�q)�N�+\�Ȃ����(zSq�ONK%�x��LC��M�#�������H��1�5H87��_��#����++ux�L����BQ�'�f��q�d_ 9?������n
T�Cv�x��?�Oٙ��J̆�(��U|f�����!���	��pà��ɱiR W�y����$}�K�c ���C�����׀��v�/�X�RPYm�Ɛ�ixK�h���m ! D2�~N��
mS�q���d-��E���g��A:QvR*X��f#LqRާ(���|���\R)^R<jɽщT���f	�_z�G�6[�㪏3�q)b�e����:���tKi��pM�f �I^n}���bL���ϸ�;N��I45t�d��M8�j���FSs"ݣn�I������@Z���KM�@�XB�:���hO�]�J��P�����av����^��ٞ�G��'|c;Wd���{r%���)�����r���#��@53,��#�C�	u,�������%v���6���7��Vh�o��HV��	�1�QPu�%��#�x�sV���γ�s��:^"#��v�.�C��7���׼��2�͗G}�]4J'cO^��np�����5j�Gx��3��N�pP$d/��Z"@�6iw����9��"���#�}��"��L�@�Z�E�؀��5���<�J6Z�M�2�W�6���>g&�U��[���x��N���@�P�3��\?8Ģ+&�2�*��ft�����LP�~͋;��̀ ��KQ��ؒ.�!s���zt���� ���+�M(�Z�М�a��oӘA���o�κ;�mW��o���/���Fzp�f��I�V��_xs g�����u~��^��o2�v�l"�nP�8qmx&�r����t�"�BK���}S��*���Ґ�a��4�$<yHˑߥ3�_����mdK6B�Q(����e^�R��W�D�ܿ��W����e��)�x���uc��A�������s|Ɋ���Ő��\>���I�ʯ����T��E��".�xr�ﭫ����9[��͸�8���b�|_���tf	)����~�ʴ�ڞ�H��y���5n���ʛ������V�z��.�}r��2<�Zhu�%<p]����I�,Z C���N�B�Q���A��2�t��0��$���8��J����2�ŷ
ӵ�� ��)��ys%�� 2����J����2k�6;��&�Y�+߾:X��rB��	���M0TؕT��q�4��|v�hÇ�_t��'<ı��α�����d�s����,�u����b�������o]�(,�� ��3Z�G<�H���RKZ��=��ݻ��2�h���S��K�������KO[���-Ϣ�U��T���gK<9i.�۫���߃Y�4�b��5��^�.E:x���U��~is�"w���*�_*syy�����kx��L��f�y|]EB]z��5�Rx)����-����ڜ<Vt2��$-�~��$�̅Q!�$���n�*5��u�q�5�8b6���_խ�o͠�n|����h��z�V��p���-�6O�:~�ߐ�\}g����]��k3���lPزLNMbƼ�bn��Cvh	<gd�|Utnp���#P�D��t6ls�=J?��qg}�d����j[�!&�]���!�	��2%��,��s�zd������U�<�\�9����1-_oT��(P;��n������m��t):}����J��x���8w���W/d�-�3�8�k��Yd2RT���"���j��,�B5��$4���B�Y	P�iJa�����lOD�;`�՟��32�7�h7F��xR��Ou��ݱp�f�Pp��Q���9|��*�-���둂��&����0u����L�~n�UYeJ���Ǫ�P��WK	^��J�6�1֗c:�eh<�x �nI�����~�C؅����2ǒk����(��V0>��!8�^e���*�pH!�-�`*��A}w��x�כ|���d	�^��9~�`�j~A�s�}��v�w�	x�u瘳���?g���i��9r-H�pk!A�zN�W�ӍjI_ʯ�W�赤`�;�}J��^4�6��n)2�6���޻bn�VgO;��T�c��`ܰ,����UB�ԛ� ][O�� �'���8��8����W7
b�OG��_�l^�	#'������Sm�����:�oɹ^T�u��Ʈ�q_b[Q���ߦ���PV '�L�b�L�b�������u�$��LDL�RX�%�*浩S�y{;�6�/��`O��O��u�P�Mާ
(lni}�kq]���ydل�M-J'�e�`�K�H��MR�I�+�w[VYW�伆tr[�x�s?u���@�U�6�b%�1!̡O��7R��15!���8�⻿M_��@�s�l����HV���2 ���Ds@�[䙁6���J���'(����h&��ǧ�U��r��Gny�C�M�Hl�a���_/��~�&UQ�X`���i8i�I�Z$��I�,$�+AhЁ�?eJ��)���ұ�I���/VAb6�|S��0t]*n�r��=->�ޑ���vJ��0{o}�PL���M�{����T��}��6��ݻ�dg���Dr;5�8�5c�,xe�)u�64R��c�pw4��u!�wX���[�t���8-bvn�Nĺ����y���N�����!)��ˀ8�6R��.d|*�i8)�`Mo5;�Q�3{X�|��I�vG��b��9Yx�ܿ_��Ԙ!�4|끮��
t�-b�!қ9ƪo*��I��y���b�]��99��B'�'��y7�qP���"�"�2w=ȼf�$ƇT`�Ȇ�Pb-��'�a�J�!��@F� hQ鼬k��������}s08��	K��W�R����T�B��L�[�H���/��5�T�C�q��XkY3���zv�f�d�Dni���A>��M�V��V'BL�Ls>t�
�g�����L�����Z-�ޗ���ƇT �+�97 ��줾!0�1iA1w��͂7P��5r.�eIol��{�W�0�
#�p�� �'_L	+�v�C_�I�E���ɌEJ�ʌ�M4�to��>T���S左oM�&17�I�2�����z�0O~��۾��HD�^���Μ��&��;�u���L/�waB}�-�q�����n��oC^,m� d[�Ha�K���@8�˷���%�����g8�ˎ�T�b�PM��,v �n��C�Cx����&ɰ�Ь�l񚲀��ʍ�h]�r*��?]�=���Ҍ���& ��q�A��_o�OI���@��c����i\)��a�4I���C�w����	�>:|����Li�e!��ar�W�D >m�s��x�y�C���t��,ϳ��&�m�Qn�z��D�"/Ĥ��ς8�?���>�̮c�u�x �_E��};�pÉI������Ip ��$�m]�A��N��/m�C���$��2C�E4�����'�"��=�d,�Q�Fě�R�$q�'*1��E�|Е��>t�͜f$uxt�Ӡ���������1��mToM�h�a7��=�.��T�������J� ��~Fc-25A���E�h�if9�]B�7�rE��&/ť��%З,U�J�H�DW��������撙�)�ō��ͱ#�6��"�v]~�]�����z�޳r���8'N�!s&9MP�GnD[��I�m���(��*B���^�Y�oI��*��y���q�g~�F�2z21�T=q����;{�����T�E:�j���?����w�jLP!X�;|�Ű��4Zo�K�O�A�KPv�i'�j�=���谆��t2�an}�$gr��\�dk[�0%館���k>N��d�Wf4����@R�s��&�ҹmP�FbX���-��UU��-j#�6L���~�3>
��|g�YY��/�P�R�O�2�ݛ�OA��fH�+<Rc�J���.�b�Ȭ�}����c������Ş��E�O 3��z�����Gw�̻j%�QY�ga`�&ױD�ܠ�
*��*[?'�]p	%?eE�������i+��� �����``��6�`��u}�&H��3����	�=$�5[�L��(�����R�zg��J𴲗ث�Vf���mW�:��
#tm����h=
�N��B6>!�p��?	��7rD9�0��߫s�E{�N�|&�S���~�ο�Zܕ-Qs��Z��oM�UA�v�=H�r熞��E_�+h���5~��縷uv�{����&0�g�F[a���Z��Jᢓ,!��tLj��uɹ]4�d΋�1�7̾T�V����|�
�ӎL�}ۿ�䭷B#a�_`�>�L����_�CٟG���I$S���t���v���w5����K�}�r"ļx�.��'�
d�r�ZJ?=R�,s��_h�Rp���I�>����:mA@��s\hW�ٮ�c���IK��A*�Pq���J�qN�wM��1�4��1,#�����J�o֤�ܬ�,y[�q~�'/�E�A;"=Y�h�#��`z�"�4�'4E�a&���KH�#J�7���Ю�&�+�b�����At�%�]iV���1�\;U���ۏc�og�B�²��!�2fg�)�/3����G���q�Ο�*��%t�*9_dӻ͈gru ^�O�e\S��2x�D&I��6�ۣ::����:�D������/�m�\�*���(�]r;i���1��
�1r���������b`��8��6n^�N�b��qc'E��s�P���FҨ���oAȘ�0$��S��{,�1q���A8C6���H���*��۪�]�ң��M�) 9!�;��Ve�3�d�Z_Y����A]UX�`�|�.҇��(�sef.nb�)������	c]��o>@
��M�^��LB��b��	X���}+I|��R����H���}�Hޯ3��z�]#<������1%��솘s�Bpuk��d\��V��A�64�Q\�Y�kbR�;����L^٧2>��ϐ�d$�	}Y=�;�MK/�`�2��@���ǹ�Y�'Ϻt��0 ډ%� ����.g�)ub�E�0��D~���F�N�C�I��|㋻��a��k1��a���pX�6-��ũ^�N����W:�Ȫt.��ܩ�R=�t��G�Q7�8��=D�En���>!��� �c�OVj�rr����c� ����$�`��U5)����ҏP�����c!��ӽ�`��N��a�.T�@ws	�����b��H����/��t��q��a��-�b 򡧗P�����?�!�*�Хo�aA�&{ÊD���V�S�U��.$��F{�`�M$�s����������DR_�ı� ˵D�@�$�[�7�b2��MIX��G��Ӈ�{3�3hq��}�G��8l�cTr׀�^�ɢ�Jg��p( 41�L�Նτ�H����=�<�3��j�/G�3Yi��=��H&�������U��Q+�h4�k�&�t2��sH&h?7����u��C-�{;��!��|�����
��yb<�mn�,P#Y3vGU�$S(]9�ޡa��|�ƴ�=�j	(3\��!�vB�u
�̀B	_���aQzQp����2��0��n������7ʬ��A��I�qC��&Ñ���nm�N���'n�ei�>��#��cz��z�\,��Z6R.�/I�~��o�H���-���08 A���,܍l�����Y쩊�'E��z��9k����l�D����ܽ͸�`������k,����x�����i\����޼lS�Qw��(�W��o���K�6��8���4�vpr�O�98.�*%�@C��z�Z��#������ˇ4�#L%F� �R|��l#�=q�Zn��w{�.`�~+��Z���B-��Pd	5*�1ˑ��9��z�J3a5	k@�&ʂ��c�[*��ST20	z@P89;�ΓQ\1C�Wxq���]<)${	0C;x?�����!=�^$k�.v�����6tCk��޸���AN<[jɥ�-�-�H#2s��'�=��uK�/"n8���5�F
��:]m�X㶠��U��$�Ӂ�?J4NQD�3�=(����1a��wl�G�B��1��'��X&�|C�s>��y���}5"JE]ep_���M9i-R�f��� u�z��ǗTO����bv'̜�?��S�&�[���)ew�����X���>��'�$;k%�LJB�_1�7�5Ћ�G�\��Wk�Z��mo�(G}�+Ͼ�*6K��-:�#H�s�My�^� G�����DՑ�{�jS{|�� \�kH��Ԉ�ۇ�W����;���G�4�8N���ĵE��e��gRl�	����dQ��@ P��c3@�O�B�`�͌�]}��7Υ��e�_ۄ̣V}��Ҫ�t�	��v�����A�v=G7�^+����}�,Sis��~C9���ؙ��4���g�@�PD�t��cS�oy��zf��N�"M�!�l�8x���o������)�zl��G�
ϻ�����wE�t�=��h���g�7L��f�����^G4~����2R&A�j��X�0���@���yt|q],!J*��$�ktb+������F<m��F���e���v��1v����Ŷ|$���3Ĺ0 �B����im�S��[�뷪���v������ŝ����1pK���Ȕ�J��-�[��ڋ�������n��ߩ�N�C��{Q!\�A`�C�^X9�f��%���g��]�F��W}w��rpn�v�C�`��6�j����/��z-O߱��ڏ)Ƒo����<�܌݋PN�R^a�a�%��(��>*�kՓM�ϴ����^@�s������Zz�����'�(xpW{�p��JT�d�+C
|D��f�j��������B�/f��zK�%P]G#�j�̯S��/ҁ��W3W���X�˾�cp�W"��b�ίh��+K��e�l�$9�嶞����=q��/�?Nydpp.[C�+�?���Y�z��vXga�����u2�ͯ����D:H��#���&C`y@��pz�p�fRԭ�g(/�f��X�"v�*�S�%ݺ�b0�a�B�ȏ`�+��ܷ	ҡ��<\8o�ٜ���25q="����'�Ae����ԧ�����0���R�&�F���xML�L<��'d7��
La`맊F/ʩ���Kx���g���1�Xb+0�����^Ҥ��_]R@�n- �8w�&C[��C�� �{S�eТ��w^;���(7�;��.	;�����<�P�||���w�K`UId�o�wO�*/fw'�����]���!Z�G�;~�#b��)���C�10�Bg�i�݈�<�u�H�&�,�ظ���(;�\�>_FĨ���M�	+���
I�6 �v��ukW��L
9����T+���ڠ�k��b��3Hh8�$�`�����l��G>�)��s�Y��%�Ӣ?�f�n��`��$[���� -9���۬o���NY�F��P�}�e@k�*�-�wV���k��aL�D�w�4�b���t���^v,�RŞ˛��fˢ��i����%gNBr�&��S_��~r�6��e- pr�i�O��VX	N�{����Ae��������<ܥ�@n�x>eY3Q�K�#C�G�%V����yK��|�'��{�R�m�E�+K�}��:����{�E���SC}�- ĘgӏR��օg��ju��#�ػ�y� -B��=���b�#�An>b���M8G�����:�����eTS���TDS�|��R��5)�D4i{�l����F���=�s���~p�I����ct����Y�5nb$���6�����fr�凢�$I��<Ԅ�{�����7��K鯆���pz���f����0M�
qm�˞�a����m�r��II���&��F@�G��P�cn�I� i8\����UP��+�5���[�d�C��]�T;ǒ�#����v��t�!�C8H�G��~V�p{��:Fu�rFK;j������/��̑[�f2(�8xy0ߑ/�����9AeGG���	�Z���>��
�}!ٓ+d�4#�,������eHs�P�K�?��FGh!T~��t���Y����Tڜ���� �G}Cx�&����0y���<Q��ý���l��A4�`��b ��R$ÔJ��i�3v6Y������R�������1��}b��3\j�$Nw�-r�_��ᔙG2��1-�=:�i]U2{�`Y�A��j!��B�mo̯&Ѝ.��,��I@�o�P{a�L7�a^'��z� 8js�����cTt;ث�@��xcZ�S��'��'�Dȝ!	��5�%��w�J,�W�S�9ί����I��s��l.��6:jwۄ���)\a�E�1�M�9������
��s���,ю+h�7O���,颞-�!v�D��Q�d2��9�|x$���vo�bhq���3��h�PՃ9?]�PJ��y�%�ܢ��I]|se�(��<��à�8pYW����6OG���٩�����en��ω^	-�- ��.�k�K�$�]�R�fNNsW�Q��������⥱��\+F�[�FM��ۈ�皤�v����!�G�clS���V��!������~3�B�H-�i'��~F�Z4��2,�f�	�=+����ш�M�2L�y�gs_�Sjgw-B.�d�I�c��]��!�[$��J����JU��{U���ܙIh����1&��V�T��&��r(ӏi]\-�X8
/k�5e)&j��&�� ������I�ij
Q��>�
�|�����_#���
��t�4�2��N�C��T���I�1�3,IJ?�Ho������M�vU�F�f~.M��Qab$�!oX��S�:'���j	�&�]��^��\Aޥ������>���TZ^ �5��%�Y{��lƗ��	��4�XxMz��s������󚭅��}FJX�n"��hJh������*]��r�v]F�p��,(��)6�	���NB����J���9�̴�;��rDzs� ��j�5v���3[�1�ء��(�d�O�/�!d����7�8�o����O�3���Ǿ?M�|A���3��)F� �y|,ۘ8�v؉X��o6����S�I��9cػ"��j�w�^�O��7����Ƙ��J�j���IK�v`��0WI b�Q4�D�{V*NsS�۪�cxC�V%����;���,Q��	��X���B�pj;�1�����;7U���= �d�5F��AY�ց���P\���,�[�b�������<�Rp�du5}��G8�̩��G/Ϲ��q1<���]�� �jUq�|�.�=U�RI#�Z�H~N�E�����6��*��OT�bY��ۈڕ72E��f��D7#E��:Z,-At�����4�����*�����"q��c��/��ŃM(�m��Ėb��zj�Z3�8A��̇3��F��/o��o���kix��ؙ��E-'�|m�[l��T<����Ɠ������N���r���w7��ƪ���iK-�Yݤ��w"%Mǈ�� ����<X7�ݹZ��3%~x#?�E�{��V��=F�1
�߮������u;&����-PR����6�9�􋛲*qr��x��xd����ؔ��G,��#O�&G";5��CȾ#���G%+�����}W��z�N�������U��t�gj/�n��QI+�C
#M�.��Y�o��:����+�`ɝUeK��p�ĕ�3}WCg���
�V�f{W`��/��ٽ��;O�g_��XȄ��Z��?]�g�{@N#٪�^0ޞ�S'��Bh�9M��j��*�7�5��Eԡ����c�s��W	Hf����M�Ҕ3��~�����cJ�t���	)��*.vRz7�4�T�nX�H9��K��߁c���y}��(V&�c�Cx/i����/���QNwp�Jt4�58�bE�ʒ�o�ʮxe�{��|^A��)�0��y�h��$ ���_��F�_�¶��~ȫf� �89ǯ{w!8���?m{ɍ��kwk�6�C������
I�]_�
A
�&�?5*xGY6]��K#7o���Kcv������D�#$��q{N��m_�aS�Br�z_|�@MZ�Xc6��Lj
b�T� R�2��|+֕�Up�:�<[��g���a	���e��MI���4�c�1�6����	p2QM|�U2h�d���;:B�X��7���x����˳���� 츿R'Q|�f�\_�P��<O8��E��a�K{[ !$@��yxޟz#���^���vBV���?tiī���#X(w6Wj�R���;��v�D�5�1�Ě�
��ND6)&����g@w�T@�%h.�*oS��[��12:#4H��-藫���CْƖ2���$�̶��jρ�-�I8L~��Ҏ�嗹a69���͸W��ѽ�H���J1�� ��ȍO�^�M�Rn��v�Z��o�.	�^�_�VRG�SO�9'|���~.�\l����[P�겆��P���s��O�ƀ%��Q(n�#Ζ-C�U0��'Y�g������\�W��rK �L��ڀ��@Ė��z)8�]�K�v��BFt����&�L��K'U�	:�w�>�DX�<u��MM�hE��Z:i ��fQ!6��7&����a\5��K������ ��4%�z`���Z@L���B�_��ex?���eY�*e�����K��Q��s���b��Ix)^MX!��_�":�q��?���֒�q���}�6����8ha�(lSݴ��L:U���"��X ƈ:�TA�.��P�j����s�Ħ���O��Q���3���j���_9./ҺU�:4�h�!�%�����~)T�nߋXE���59B������ ���+Su/?/Q�|� HZb�HƐ���;ǔ$1�, R=�|F=���_CD%\�D#�����hG�j�3!T�`���a�9�������]���L�/>�d���kp/ÿ��w]���rt���k�QMS�w]{�ܯ�Y�Z��y ��p�E��m��v[p/�����C��W6�a>g�����e��61��ڗ��w�zM!����4��n*�	�ʋ�%gʥ���<Q�ޥ�Ǆ&���YR�M��S EN V�����jAӆ�@;u����-�f�?J�;Y9��U�-���`�64��͂�q�`�x>"�	�c�����F�#D���|�a:�� Տ�vuSM%�Ef��J��V>@O�X�w��J�@��]�v�WB<��9OȎM�a�*Xs�2A W��e-,Z��>��ZZݞv�.�W�۸�'�V��o��n�j���E�^�_ ���O�b8�'dO)�����L�
j�ͣ3�����JO6jg\�˳�ID��V̠��]�w�KN0��6�b��6��`pŁ2|$��
�ҠR�l�˞`�Co%p�����ܲ��>��ӗ�y�U1U@�s�� |
��;.�Q�xY_��W��Ӈ�c�s�-�r�K q�����g���P	G�{��Ho8�@���N�&�?�D�v=�[F� ��VĐ��\O.H�?^�����*�q�>�B��_�ve�$M��Z6�1;Q�q�pB���aL�*�SǪ2��K�~�?���ۨ�#�J����qou�k�B��`��C��>��aܰ<@��y>n�A�bO�P�l��{�;ʏMH@�^3�T�yI�
�&��ЋroΤ��R�&���j���]�O�^[��2�9��G�M�W8)��Һk��-�G�i�Ot��twV�̌��%ߋ�l�ϲ64"�$o^df�.����G��o�B�w��<)W?��+�����c�P�9�-.��D�z5��8��<88F�T�R�D[ ,q �s���&u��O_��q�-����+u$�؋N�e�ɿ�j�$�S&ő)��E/?���U?�]���J<�T����PX�f��5ƀ!��K-u�����	�Ē7���y�WC~�O�1�n��������IT���a�A�-)���q �xTU��x_<:�	�5�T%�FZ��ܢ�<})b���;�9�M)���c��u^��M�!ܩH���@Q~��m���%G���"��˗����ɔ����|��S?ӿ����q",z�?`ݜR;X����ۅg��Y���m�V@e�I�s6�sk	��^��/��Q@'х,,�B�g�W	+���F�8�� &'+}&��/��#Qp�Y]:Lk��`P^-���s��v��i�,/����I$��%�t��c���
����\鋽����\� vX�S�$�O�\�/V�}��"�����wF����~#h\�aԨ�g&%P��Ϲ� �s��D���]t���>�E��z#6ȫ��0��P��wO o���#�,{�����.���I.�k��r��+"�}!�@��N�r�(+"sn�����%��;�;���bz�������c��c��6�'$ͦ	b� ��4rU�)��w%('5�t5�7N7I֮rVS�#w[8*��'4��MO�����/�-SB��t���1��Q���I�c�j�	�m�Qj$u���r�=��[=7��ZM�6���{����A�8��NU(o޲
�40�^�<j�w���/�x�F�;�G�x������( �}�b�R9Dmt��-eI��4Qlǅ�#Ur�E�� o*ܰV���Do�3�U�H�N��b\�������N�����~:�-N�JИy�c̝�zt�kأ��V��軟���O�Q�lpӁ��Y+��h��.����� #�FY�g�UL��&y����:�i�'a���JҪ�;S�/ن��u�{qF�Ф*�
HX�����`�"I�h�Hf�7۪��u�X�=&����~X����.��e���~��*��qN��	�����<� �р��ͼ��ir
?�-*�oa/ ��r�rK�[͚�2#�q�O�m���.(@�3�:��L�FZ���j�H�`���e��\YV[�!�Q	�͖�>�V��q`��Qٓ�C���i���6�8qz�i�ɴ��gP�������ת������W�B ?��1��UI��|"6�a�5Wec�#�)o��+@5>��{�w�e��m�U���6q�}=�R{����:��
-Lz+j�˯�cBeP���� q��@#��t ��Ԓ?����XR�H@S��k�㷛[a�B���U�:6�����o!Dc��B�<tL0�ghL��"ެ�s.�C7�pW�@Vctf���q���q��Ұ��G�j�8�,+l��9��p�l����h�_+}�&0��m��d\3���\�۬.6�ڌ9	ؓ-VU�<E�%�V�ܡ~.`�r��fɏ,kn�h��W|r�q�A����u�w��R��o����(�l�d/�������HJ�@�� ���� �����H�E=T�.�_
#����g�tA�殐%��1�)��{�,�*�ѝ�M!]ƒ���3���IXc�?�s�Z�5h��qOr�TR��gБ�i��~#�['N�׮}O�s�e?X����.��'x!<�&w��y��č9\���M�V0��t��5�oةH���_�n��Y(1tF��+!!�=�c��F�K�U�q�Q��)��C���3���b��9D��Rkэ�N�����6̴��;���P�W3�3������RuL��V�/������,�طWY�W�~0h
�$5�B{VT���0k�=x���s�8c�+�l�6N��hα�����k߁6C����t��Z,�Qg�~�h���5:f�5�t�kx�^��������D{ȅz*�v*�����/V��p`߂�'A�E3?�Z�jk"@�֘��Ӎr�ι=��C%��!G�Ѧg��+����zh#;��w���
�y��9�>��3%�6e����&J��%��̃���d�^I����>��c }=��\�v+�b9לUk�MU�P%�#���Hlx���R��eq1� s[��g[tU�MM�M���K&�6F�MI.��~�(w�"��B��5D�=��>�k�ɭ�=KN�k��5GKȡ�Ӭ"���X-t��y�NbM�/S-+��4��E���9`|�K�
�;�1��7c ��?~��eǿ����z�H
~-�t��6��zgG�fO���uj�S
�#*�dx�4�m��1��C)�oJUb�w��E�Qg�����&Ý��	����[�1QM�@}�S3��*�O��L��ނ�!�+�6y���=��X�d����%�K��)��P���U�
mx+�2��2d���)8�e���ng{�5�~���]��x+f�K��M!TNХ�/��j:��>Sڹ�p
��yʅ�3�_��E>E�_ ��p��?��-��+?�� �orf�7N�V�X�C�J(X���Om���?,�db�<h���a���Rm���bCJ'���h.���y2VfY�Z��������M.�O���e��r^�O$!�P����T�W�ߖ���U�l���o��6�jk��&�PNE�O�XK�ߘoX����x �h4ܓ3V��e�B�A��&S�h�q����Az������5S;�Z$ة>2py�完�T��6~ �[+3�g
���DsQ0�����JiL�ɻ<z4abM܈՞(ڮy� �a~�8β�K�Q������Q���5H�l�x�r��v`��f�o���t��'����C����5m� P����� �����������sȏ����j+1c�������q�UI��[�#1���w퍫e3R�g��>���dc�X�E�xm�ٱ��� RwӪ3#�}����2�A����톲�Dp�g-bU�?ʗpx�0���Q����*�_��q���Qp{�:Q���>���k�I��{ V�?6@(� �lr6��	r;���<�pwJ�Q&�I>ܘr~��E~q���+����5�+��ꘋ �v;�~� ,:d�*�oم
�3��>ɹ�.IE��K�f�7�A�o�C�A�"�휶]�<.7|��K�܈R  �&�]��O�紒ƾ �����5u�����~|�Rz$K��U���k�G3s7�~Rs�j����7+B���w�����V[�S�	1x���Et�Ɠ6��s�]�]���U3�2�bj�,��CGN�����!c��6P�SC�b�}�o(=m��2��8��g�h3�Tr��uu'��9y�t�G�=��T	
P�Nڿ#��_J�9�9�5��-�A����b�e��=̉U;7���bG�:0>`p�>������\f�!N8�p)���,Z��\����E��\r�a�͔8F�l���)"F��)�K��Y+�o�+CQ�:�����ԔS�����xy�ũQ<�	��{M�|P��7MWB�Ij�3E����XTF����it2Ue{�~�ƅ�s{I^%�{Z���:�h��Z7� �X��v8'��VY�)IILT�D��>aeD�Q���'p_�5֢���4{�ɄGGfe��s4vi/3]�r��v�M�tN��Pp��Ш�т��u�a�:k��p��M���S�z��@�;j�״xf�ې�_Xq4�z�����g�W��.�uMUf�n�/@�k��,"����ͦL$�ǲ�_���]E�cn���۾�o5�Лe��=1ה�fժ�>Y|�.8r�O����7h\W�m��Y�*iu�@ED�
�GMP�Ƌv�R�z��[�7�7�'����y_���q3�Q�\?�!�ɖ:O�F�VZQ��9n�wV*�]�����߉��v@�P��pK]u�kMD�<��{@���J�@��I��h�d���ba�$F�<e_���_�tΜ�'~�K�`(D8��'�%Ա}�����y��$�z5!ph����1`I*A���r^@P�[0ت}O��К*�X�n��^�,f�!,io$8�ki�g/MΞ��b��vE��I'���L�u�T�����1��t����_NL���qe�Az��Y,�?�!���f��ўq�y�h+I��������Y��Xҹ����[���w�]� �7��r��ObA��Zޖ������YV�?�SN���~��*aƈi���);��"If�m�L�@�#^!/s�T1��]��f0!��a��ym������h�����Q����Tin��ĺ����rf�����	A�]�\AlK�;�m�	�V�W,҂�>��Z]0[��) t��u7���6��_ Ldˑk,`C_8E��M�hJC+��ў��P'��I������eL�����d���U�)�t�A��@���m"���D@�%��v��H�����&h4��f���TC�����K3�z�̲�Y�HWRr��
A��4�C�a���"ng�]I9�UV=������n�n��7�-�i1�^��-��x�d�����vƧ#�
P�N=?��1���hӚ,ϗ��XJI�Ģ�SWmqQa�6r��9��E=�2�L$��)`"%Pz��E���j#�"��t�|�v)�����\�p<%Y�ǄCZ��pv���e폘{�t�Z$ݴtX�����̭��V+�ʱc����C�d�������ĸI�Q��0�B�Q��op?���4��Y�Y��/;�ҶqA�*�Ӈ?���	��g�RG��
�}#�O��� �C����Be�̡���ž�?0 �::�)�Zh�A�2�rY�)�^��#)M|[������O. ?��&7C�����`�u����Q(,�jM�$��/�o�����v���В�|�W��۳�8�G��1�am	�z?��D��E���Eף��(ܿ�3J��[e0���i�5�R��w��9��WV�p1�N:;�H{a���H7�ާ]�y�˳m�������p<�a@�<����,�~����!-䡑�WF��řs�~���0{d ��?lb�Р��Ⱥ같�mh�b��y,�$�֛c� ֹ�R��M�N�X<��6>^Q��n�RR��S������ݦ�O�O�>��[TQ��~&ֆC�����y9�u���`�0taKn/�V��'��!�W�r9�17_C�j��{^��|u2��&,m��9sv�Pء�Oɚ�g��l�R��n'������ gv{ڗ`Ay���p�S��-H�MǏ�z�k�L`���1L9�҂z�����N2Уb'T��ޙ����� :��C�	��,�<n@xh~S�4xw��r���I���(.����\\_���{�,�Cچ�/�'�4-�s c���-?���p���D��y�.b+�S�\H"�!Q:�=O�@�fx��$�!�kjb�֑�?I-�`_4�>|m��s�~��B�ou�*�+�)�X�KH6k��ô!�[]0���Lm5�!(�Ǖ�_�n������ng�8��׹�מ?�v�v"4�5ӧ��pI����ف�ZL���E������-���.v��8�� aj�Q\�O�-vH�����A�F�D�M�ߙ�&�L�w��-Q�e��\��G��p��>'`�����q���Y;�hN�S,�r
k����IG#�@�0g֑��9iJ{tiX/�/�(�҆�D�]��#T]U���IY����M���o�����bc��>d��aۗ��谷8zA��Qh%�m�v���g��B_Ϫn�4I��_����n��A��]��S��8��!�w?
�UJ�+לTb���ɖn�r�n�g��is5 >��X{?Uߖ�T�����%*�#�V.�#��� �({�wܐ;�8e�d>f��`�H8�5��U��^t�f��Đ�Ɏ]�Z��
l�t��F�"���\����0��дu%K���� ���t��:��1l<�C�*��l������.HA��Bvt92j���w3N�Wl�堸0V���L������"�&�/��T�DT�<ު�W���M�uX2����f�Ċc[�����?��:�b�򲞻Q��4y�~`�}�����2؝!����GO�P�E��c�E9��99�5�9065��ٝ�ڋ@W�������~v�P���'49�R4�G�h�e/�F<�3���)h����j	��`�Ǥ2��wí���hy����B��Hz�,U�+�oOة'P���ε�G�0��b߃R�u���[����@PB��X.��P��_ٵ�AC�!�j��*�)xJ�.���|�T����A��I;�����FN��e��@]p
�I���[�~��}L+p��O����$���L3,Q�/�D���nr�5F��s}��x����l�c�s^D]�pԁQ�'�5�J:˷P���J[Gn���&P���F���q?��%,n�/n0ۅ�q��|��32��A t����+�����x�]by�E�� ̀��ዜ��l�S�
~��m�&t6غĒQ<)��h���ƺ+0G=m0Ƥ�<��[��Sv�i���NKx�$������\v;�=����ܰ���H�[����EZ��3�eW��yn�G�k\�k��H�3 �P��Z��yhQxr�*JF0o��o���V~�()zf,.� �������z�G\�?Ţ�����V��ǱUA�*����M��e�8 �G(/U/�m^U��qZ2\�yJ�"��;ؚF)>�x�Ct�m�������;��Ify�"��eX3(��zy�F)���ڤ��[/�
�mʺ��o�M;�0�@h��~�S�\|*���D�pz���U=�R����$�s���Xֽ�(Q�4d�>:*g�7�)^��iR�}��q1�j&e�D-g�H.���Z��`�b��R3��v?>.�j�T��t��f�f5NIi&�	�\; �X&.rO,*)�^sj�"$�O�vQ���Z�r�?xƀ[����|��&�̥P&n�������{�P�a�,#���8��J�F�_v�G'��7�˄�Z��g�5z���)}0�/i��*jvzx�0l�����-�'?*�d�e�Qt�W���0�[�xc	�|)]x7�!@N.���5J�ߌW���cl����+�FI����Y���'�:ت\�Ad��o�[t�v��%�Xy��Vǲ�:5����w��x>�Y��{�6��"]%Z�N�Z[�e��� V���r��`'<j��e�O�4�M��w�#�<� ����;$@�5
�~[ۧ�şH��!�H��&:��y��dB���|	��h��HJY�����>�3>O����*��̅�s��r�e�7�DD���=E{n�b�Z�����z��ϋ &�`ZTj �5�;x�{�Y%aȇH1�5�be���(����ξ2V��g:h#�^UU�D$�ha�4�Ԗ�R*�W+�m�Z�ʤ2_�ː�����ʎ����W�2��䎉T0(��T�iV ����|����Y�:StO�#.�ܰ���uW�YҘpQ� ;9�����$@��q}��.�:W��\�!X�|*��m��FM��ma�~	ܲV
x��-Z����t���&���녠N���wF��W�h�'a¬p���̫wŢ؆��(t���m	Q��Xfw�PA�����ox%���b{Z�S��;�!^�{����3K(u]�6������a�q"�����1��'�\�(��D�
sM���lXұ$�,@��oWܲ�xx�qu���4*�p������2||�P��hO6��L�3��K~��cTwJ�	�>��=�\: ��w�=���f߁����&iuZ���%���~��T��ؖ��nX4�R��_���.&9o��Ne�q����?����y^�tp�&&�+o��"�6M������4�Έ��#�lvf�FR# ��}]R;Ŋg�jGGq��
:q��8:7��fj���0��_��=fD��C-���W�27����B[7�z��,�tk�p�5*u�}c�87+�t����o��s��C�ݴ b��Z;<������������9AI
���.��V��̌����Y�ﲄ�~<��F����O=��Kv��͇�J3����0r�5]F�+I9�7]X�¤I�]T���UL�
���ϡ�I�(,�K�m@K��Z
È���me�=��2����[4�d��|6��� �J3���(�Ћ3bjs�3�1F��P��Gh�ݙ��V���,�NoS�ri��ƈ������I"�sR*�;ٲ'K�t��b8sr��G�h!G�!C
���q�v�S���d>m	����dh����F��z4T8�q8W.�;B�Љ���3C��fg��q��i��v�:cQ�٢��
�o�7m��w7���bwx!�G���&v��PZ�G	������>�?*����D{H��/['�^&C��)X�����(�0+��u!XU��_�t�$�yN���Z�b��q�^�A���:O5���4�mz������%�#h�pհy�9w�AE؊&�AkR/1(�cdn'�H����=���� 5�C�b��ȑ�9�u.�k0�Y�+�J���vߑ_1�D�e�����!D$=����ɍ2����e�BqL�P��Ĉ*��Q1嵫�g��$�neߣ'��U��Gh#���R��@�������p�m	הt��|�=�
���B ��6�c6~���������kB@pz�?Ʀa� }��J%���2K|�����ڛ���W�_�TIY��|��_� �q�ܾ�N_.�����+,��R:G8��jC#(i.R��2H��3�J#�J�88�L$� �f�-�,{���g���%�V8�]�u,ߋ�#�m�5lq�qDB3�� �x�ITZz[B"�f��E5�w�w�L�kp|�s����X�ݍi���d���X�~���./!펼��:�a7�֕ݝ˩�����ȭ�]���ߎ�oI�Dn�U!�����e�k�%Q�T��5x7�q�!�xv.������i=2BE��g.�1��br4��Y�g�񟯺�a����u`k5���o���x$Xk�EV������?��4����67C�_O������}�?C���Su)�g'��b�S��^�B0-Ů�vQ4���Z����	hs�^B8���ĕK�t<�K|kE���zCB-�{�o�*?�e��qX �~+���T�3ԁ��x#5�b�Ұ]i��k;b,�4C����~� �J�Y_��V�T�ʍ�~�Z�����D-8��xI̮B$ۦ3m=�ߕ'�?�V͗
xe����E��c{��h��/�.$?�k%DV�!�5t�P>�Cu��Q���1P���qMM��
D�����H�$ ��=O�����:Lm����~�T���}m�\� H�VE��wl�L�9�8�"֮�E6���U�x]Dyy���:�A�����Nݑ&��%�P��.�໩А��3��I��.��\g�v�c0���*L�[l��V��f�6znń���,A�_ c K"���s.]!6x�h����&}Fב������S�P���PZՁ<o(�U��",<��-��ߑ"g�5;we�p�2���Ӽ|���m�Q��P>V`֠��#��6��%��%D48�Y��y��v6 ��YH�s_[���-¢���W������m��O���z�o���6k9R��
�tB:&a���tZa0�jb0:����2c��:r8�tE�Κ��e� ;]�{a3]�|r�+)���7_��g"�nz=	ݭ�nNʩ����==/����`iR���� ,�@�%-��>��T�>�QΫzqN�g�͔�m��/��`��5�i��{,<=��Ә@
i�fDM�����<=T���f��8R�)�V�ߵA9�s�4�p���4���|e�;�M�{�أ=�rZTq#��⇳uitş3�){�`i��-���y~fS��BA؛�� � o��l��J2OcĽ��y����:y��Z��!��s�i��k�:0�1��Ú�7D��a��^c��c��1�l^L["R���'������i����y1���P}WB�K�r�z;ރ�r'�r����s����2g�n-̀7�(s7c�Z���9�WW��9�4[�	g���Yt��r�Y�흎{?{��PȨ7���;���������^_�E��KG���z�[.�"��y�XaR"�ҵlQC��hƪ;=5�IWr�w5%t+^wm���+�m�n�}&MT��\��
� �7�}l�Vq���fC�C����ڝ�F?߉dP�D�4�S�������Ub���� ÜL.l]�}����{f{pm��Q�,�,h��}$ �<�xs'l ��3f��{±v� &$�n�54��r���e���\�g���$;s���@�NUk=��bb�p��m�dŬ�C�N��k�b0Z��{\5��W'�/��$,'���ɶWi�f����&ԥ(7���΂գ}Y`c�W�qŒe�O��K2�=?m�f�;@����{ ��$�Έ3���gz�=W��s&4A��G��O��EIo��>�??��]�MH�7��V��F!DB[rv�(>��8O|���Q�%����c"��OH$���@�����S�p����j�V^\��ϵ�(���gc�l�ޅ�i�����6�1l,�䒱��(s��Xug�(�N+A@~�}�=w�Y?V�}�I����������<Ƒ�Nt�f@��u�@�v��M3�y۽d:���	c�!���_r��m��s��`�B����0ˆ��R�k��I~�/�rVߟ�M�
��y��*��'����1�A�ہ�`����s4�s�w�y��6�.��$4p��܌�e�lζ�8u��^�NW�L���t8�}�"@�|��Ƞ��3
��4e��l���d��`(�/k*^�W׽Y ��Q���8�vk4Ǐ�'9�OK�:��Ӻ�~�tL�o���"��SLa�!N�)���=GC� �1��ʩ��D}�͗��SP��/k��>�����m�P7�yI;����{@ղL��1��������YQ/�K��o��Wgc=$T�/�Lɴ�M����K��H�v�.�R^:�2�u��2���REa�M��o�5�ct�Sn�ޠ�5�*��* 7ݹ6;����*"���;�(�C�݌b�'����Z-o��$�i����~:���c��Ǿ]H�r���%VN�������y�*���L��!,+����<9�6����|�\�j�c9EZ���B���[�Z�E���n�{a�D��ۻ��랭�Tq�ޙ�DF�ׄ��
|ɐ�;9�E�ߵ�C�3�=�V�=����G�\������+Twu�WR�z�ޅl�'�*}Fi�6�H���T	Mօb��[�5��wyuD����S�5�4�M��)�e�K�= ]��6�5>t<����GZa��Tq���q�/��f�%�nW|�H��`h噰�Ju�qWi�4"4���6jupLE�&�W�ms`�I8c������+RR�RU��>d�sO�2񍘴�/Sz�7�/���²p_�[;�5������w����c�<'�&���YޞP[�&���^�uNђ���~��5$��Sf�f�x"�T<���D�(v���k!�{YS{IɝD�l?�c����S0�sQ�R�/�YKh/�-�?M`eʁ��&�t���Xݴ[	���7��^��W���W!���m��k�Mj�4m�V5�پۀ��Y^���96b�+�C�U(�w�s�Oб�������ؖ0׻A:_X?�^O�o�-�Vq!z1�u {Q0����mr?��;�C��?i�_���|m}��ˬ�P�x#�(�����E�<!Ӽ�x:��2|���O����/:��5�/Y(�RQ�͡���H>d��k�j&&#�_(\�)�	�xW!���(�������*g;e&��|Tw��[�4�7�9��C�6Vr��v�h����XU��4���tMHD?R�&��N����uwV\���=�	��% �O8=�a8ב����l{sXT��~����Ф"��;�xz�q}ØP�0 
��2�H����L�U!Xdz`�s��p[�J�6q��o?k��#]����x�BY��\tLɅ�;��-L�X����F�]��tZ8��� �	0L�̜
-�=5d�X��\a��%T�ҞX�	�����.j�'��q��#lN&�	��4�i)oIW���^fO?N��dĿ�G��-�O�Ԟ#���Sj�a�Ӄ���ϟ�����ۂ`
vt7G�;�Z��t�$�5�|���	�cNG��k����F5�mp����5��Б�s�3�@��INf��!�X[�5`C�-� �܁�q�	-Х�h��&&r���Dk(�[V[JV���7�3�D����b<�,������>���d~E.��Y��N{��9�h`j� ?�A/	z��٤ɏC@Q��ja�?T�Z��F~I��Y#��c���=�P2��T�z㯎 ^�an��,��r!��� oM �r^:�M]э�Cl?1�/�q�w�B:�O���+���|>��q"'���4���㐠��_j����E��Kp��g4�'0҄�-����:}��Z#���@�@B� �P]�����k
Mad�^7�T>�y?ո�>�|V8��i)�a�Onv���S�3YP��k9��an��b��D�(�L���Х����L!�IH�}���l�������s�#Un�C��^���nX���1����+��a�Z�ŕ��<�N�*]0�����Yz�ߨ�e*M���6Ye���� ���@/���+�Z��\d� #�������Njx�#�9F�v"�g�������ݸ\�4x�K��-�q���1�$��������`&��������!+b%�`)��]��ڳk~Ƕ<��߱��L"��6�!��Պ����I,��V��8�O꣱_��.9�^�����t3�GL5�$ȣ�	WR�=b�BQG�k��9]���Hy���� �aw,3�]&N�~F��y5�D�N��/E���3�g���"��l����l�@��Q	B.��jan�&Z-�q%�csd�A]��Ez�~]eϊ ����l�k��1E=%�J�<ղ�&o��ɔ@>b�m�� ^^x��l�a��oV�<s�O<�H L��
�Lo���x9-&7:��Q,4��R�lT����8�-����v2�u�B�h��I�.�Ǻ���dM?����s���s������#6+j~%n��Mc�,9x`kjU{����U:?��Ge�>>|*�N?A����C5/h�e,��3�NZ���XI��1�K<�9Y�� �E�ȋ-d�>k�{�CM��-A�i�>p�ǵKx��o��i��� ���j�9�EɘM��'�ԴH-!����k���t�Y����E����p��Zu��5<��J��M����+g(�����@���Ի;k���t"Z��D-AѪ�k�!���9�Fb����A5-ubLY�)�O������׻j�a��3Н��~��q��>l5=F��usSlR��T��|���OE���"G��6�r�^Ͱ���@1���+t� �L���g�>o�cT0�"2�S``<ql(>\��fIy�h�)�][�1��2:K���Zgƭ~�6�����3k'1"�(Z�:�@�[⩖���:=$d�����d`v�B>�hAɀ����JzoH ���S�軩�4̧קɪ�/��Ø�-N�7��p��tQ�k#�ŲA�h=����Ap����7���LLPOYnW��tD;���'���$�.�U(f2j�?����.hEof�o�JsШ+cW}kM1�C,�f��2�C3��tg?�6��RN��f���ft���u�=�K�8I�=�q��˿��+�ѽ8�)%��-�E���W�q/�����d&C@�wg�}��Ze��P�w-Jne(�Z$�n�󵫎��6K����B~�óNc*/����\�i�͖�W)��T��yg�8��\�
O �΀^����Co[��"m�u�*��Eצ�2ϋ�x��E:�g��ݠ��6Qqۘ���@��rb��"u1M���?Bv��rj0��V�.�0�a���X�=��L�E@ڸ�K�a}A��I�-�<	�+�v�3"����Ȧo���8��ɝ���5�J@/V��^x<5��teFn���@�|�X,��,�d��o����$^7�Y�I��x�y(�nn&>�B���U�DHQr(�^�2��]��mO�P��. k����
���\ff��P�T��4*�ͽ��t�����W+���;��p����F_�����2���:x]N�hEH?��I�Z�%�g�1Y���v�<�|����)-/��?�{p$ �W��h�dJ�`���k��(C˪\���?�7��ULD�&3N`w�:����i\\^p��ݑVn�Fax�J�yi�C�wF��ԉ_���v>�A�:�1�M��׏U?�UDLY��P����R6~cJx�L郉�>���b����$�9~/�K �a�$$��)�C7��+4�,�bP��K(VJ3��o!�)
v���hs��/�%�N�W�d�bL0�v �Lb���gTp���x�j���a���(�!W>l�W$��h�"	N��m��m.��y��"��4P�BL��x�[J�逞Y�F;�G�U��&��f!Lk�S�ay�墯�`�Z����3oQ���	��>����a\G��믪����{-y�����b�I�M�Şܓ)��d�,��+�*�v��	��r �l�����wH��D6���k�Q}t�ۜ����F��.Qf�_��ˬˌi���J�0�Id�d-N� 7G�׍�*����RH�rZ�#�a#9V?]m¹�S�:���Fs�C(� �E�Q@<�N���3�H'Y4X�*�OGl�=xY1�KpF��M%���0;\3c�!��[��T*q���x\��"���T��p{�G��jX��� �[�M�2��(ߖ{Rw2��Lq&�)�J���YC�w� �7�[�@�[��G�C�x[�2��Jo����LPw���q4~݊q�����G�����|����6�b/�	��`a�� �����Ɓ�&�+����0Z6��჻�ȥYA=-.�1���5E�ፃ,�C{M!���������4H�f�?u�.�|}�i-Xv�M��{ݡ�z�u	%�t��S>d4ӝ�c�e]V������Ẁ�a�g�uC���]A���[`(�-���T�I�l����(=�$ ��=�O����j[��vF��=F"C��ov��cY<�d���yf�x|(N��+)���Rp�JG����7G�@)K�aP�w�D�����_�P��M$��<3mQ?��[t�B�ؐ�缬�ߤz$�Gzo��d+y���S��\���������<�Z����|;�lEv�vf��Һ���D�������tU�_l�Z���)5�*U`̏�ֆr�7#u��5rst�Ϗ�����Qh��[����(4-��wԍ��[=���C�"�	qߣئ���\R����IB�@���>��1�y���k��Q����Ex|��fk�ʶ2��?ev���2d`ug�C%Th�Ю|�]�Vha]֕6�� ���E�cw̌?cTMNr�	��$�1�{1;o��Kƣ������T�(�h߶�s]�>L(}`���2_��~l������lNϾ�҇Ou�R��C��rD��{O�K.{Lę��,�q��ξ��V��%�Z�y�6��#^!�����#�D��=�w�=�-<�"W�'�p╭2|�j#��]��������D5	�_p���k|� ��\����̐bo9LR��� 5�"q(�x�jR0���.M���eA�k�TC)�Ѽ��_f���k,�������.�n!��VҧER��f�^�h���������,���5[��8�t{�n{�|v���L��j��`G!�v��ҕ[B0-������hr���}o!�w�h��r�l�v������w��Ӏ�9�!q��5#�"����ZE�%E���mT]�?rcs��fv#�F,�G��х�T�v�2���eh#���:��X�
M�q�r�ǋF�L��+L8E��8]H V�E���~<�
N�dൖж�ǃ1�D�Q寳����W�s�1��G[�(R`���NI�"(��t��P�;������������bMQ������g��_֏{��}����WT���J� t��n�z���ﲛ5��{ ��mg�<LP?~bm�9�<4-g�D�����<��0F S&��ϡ��S/��$��;h-�ǚ�s��������!PT��=�X�r!nQ�d��7� �,���
A����\ye�5�?'/�1k;?'1����B�:+3e��=R-��bH'�	W��K���-�+�� ��IF�=9ޚ4��m+�~҉"�Y�T(�k�i���邽����O�$�.�b�.i���	����I?�	��f ���>OX�C^n*+-�m$����t�]،���r�v��t܊h��:dz��o���fV!d���h�?t��v*ګPu��u���',c%������o�7	�%�� 9Q�9x�blg�R�V���Fo�\-�
k���n���@D,tM.uzOV��ڛ�f��Ջʒ�]�%������~[A�{8_�������J;~|�e� ��>h5c-C��(-�{q���kڃQ������q!1yUn"����ls�K�ތgFw��θ�^���Yb���V�T�vgK;ͨ���J�<�N&cS-��� Ǫ�(�Ϣ�|��R�_��sK}	y��'��A��Ӧf�J�^c�q<�t��h�B���ݜ�y�ʫ������e��#'b�=(g���������p������N�|�!B�P��c���ޯ��s:q�4'�kf®c8�fYaHYeOL[�du��y���L�]k�j"�"�������z!dڷX��kA�#��t����p*�#O���ͪ�5��Z�q�h�p�w����z�5R��)++@t�ro����ʖB�[���?���ʔj�̮p��iP�J��Ou֋f���R�_�pj���z�2��MJ�/˄⡸�w�<I��b��A��M�:��:�\W	�� ^Df��3j���=s���v鱃�~� �E�@"��9|�B>��s0����e�����ȓUn��#t~��^��9r\�Q1q�%5=�^���u.uL�C��b]��ݽL)̺և<dș�`f��B�����`9j�,AT���=�"g�9	�R��?A�c�n��b�p��/=iW�P����5y����US��鹾������t��t5*$�5)j����V���x�VWN��&Ĉ�Q��+�X8��`�
��;�>�lJO���=���u!��b�F�m�or�=���,���A����g�\Cy����1��+�;f8R4~r�N'�������PZ�q�Q�e��
 ����tI<�~V3kk�K������7�XbH�f��nml�H@�P1���)p�d�ow�lx�F�#8�6j���7Z�c���_�x�f��*1K�Y3�4�~f[�vKq(�3��"�s$W�߶O?M�����슥,��k B^��=Ԙ+>\�ԣR���H���y\���Y�Ƥ�ӈp��>�J%�xVb�)�ߜF�|��f�+��:.yy��iE���,��u.5O�_���ܢ�����8%Čo
��|hk���o���5]1W[��k�������@u*x�:M{�,�x�$gg�l9R|.�5j�}t�r{(H-�.�W�X��Ô�2�!��?N���[���8�L�c�xaa9R��GB��̐zC��H�o����U�4VҌ��^�{���FL�M���1�G�ﶝ���QV��Օux��EW�ԧS*�4�k݆�s��}I*7P��������¨+���x��͛��+�H�>7k��u�D������a_�l����r��d�����|EZ�����r�D����;�՜�?K��1�ta�ͬ��I�mjb�ĸR�!]��>_��U�H �rk�e���J7'�?+�*��s������k�_�,⹺݋��`υ�7΁�����t�ug��6��y%h��+��ԋ�q�r�-ֽk��@�@�����w��p*����.x�ϞN�te�ۇ3������*�W��:Yr+⮍'��K�7���*���R*0�ÇH�K��8r����'�1,!��9��%d4f�������I^�i��)��M���!��פ����R[2w4�t^�-�=��lD_��s�R��闩`���� � �����%+�냧�i�g3�xŔkuy�\)�D�0��5�&-��~+H���W��μ4�srZq�X�����^���_��ωu��y�Z�:�W�_j����T�=fn(�W�U�P]Ѱ|�,2�L#��!N�ъ��v!�0eH4�;�.�%���/1SV�^�u�U���TР���VP���w�N��;��B��LjS�Bt?� |�:�k� ��^�m;b������ĺA�P��Kq惭~Z�X:�B[����{��6�8�`��>(ڳv��lc���K���'�����Z��ޞ#HS�z�'��$;�%ɸ��H����j��܈]�Tx?}?�7ǲx�s�.<S��FE�Q�nd�?`���u��cIOj:߸\Br-�*�hE2/�����p��r�r�+;C�.�a9��,�� N:@��m�u�fr���&�Ԗ�GͱeO��R����F/���3d��r�۠������~6���Tn ��ါ���B��,���w�L�F޾�lf���@V��؈���M�N���~�9�.rgjqT(�M�T`�-��RP���9"'�VɊJa��d1)yqQ�X�v����`l��*�8=���>��+���z�>#v^�f�>z� R�utϓxb�ږ h����xӻ��o�C��*{���ě_:���Z� ��l:E�(|9��k����@��n����d���>�p��؞��V�^�� ̫_�����nYd?c����7A���J�O�ծ"M�j"8f¬lʵ��)�߃��qU�6^��K���������'���~� țێf�)7�{�Z�W����M6֥󮏊���b3����1�T�榤QN��\�/�,
���ϐ�1���a�6������=��P�B�L�_�����ʪ�i�!/L�hQU$Z�{��s\a���a88���_ /LF1�Y��\N��� x�:���5�Jz4�p�/�^r�c��2[�נP��0���҆M���g�L�@��Mpw�ž��<bm�������3���jiWHln���}/"��M�gR����f#R���`��#�	")�%" ���J&�EiL�h��LͅH��m$D=�8�?w�
�SR��>��fj�%�C-˶#	�׻��{$��K����B\]u`)=�  �R�sr��-KZ&w�=�������<�a�c+���$��л��-z����<�ʑ����[�m�����^iv����[t��k8U�.���f�̦p���Tԣ�^p!���:1��T��o�Ce���� �l���� Pw-�;�T�9Z�z^^��x�ZV��'��d���Q_�ȕol���)ٝ����y����7bV��ϨF�DaXҡq��A���?�)��>��:�P�آ�z�.K�OW��*��H��6f)��ܫ1�S�-�"+��c�j�� :9��s$��6d�/̡9_�<%�P5�=���A�ɧ�cJAh����Y�a�~��}=���EF���H�I�W�@̫bB;LLA�։���ຐmU���d>>Ҽ�'-�Ð�^Avr�W����}W)��q��/f#S�D�9>�L���A>�FB�vB����G���xA�S�:�rC_�ĺ�V|��FG�^=���!�}�(�~���(�c6���;�,fOg��7��I�����ߧoB�}���Y�6�mlv�������&F�;3Z��M�%��8�d�I�9b.=}=^O�2'#@� C�Qmd��b}�y25�4wM�����x2�g뛾����?&m}b#�3�\q�����|jF�f<��RQ{~,�_<R�s�.4~�(C!x�.i�s�jĎ���D䬗&$ �*��g4Q(�����Ю��$�g5��	m����9:�.\���Q�'g�� �u ��ۡ��{�L�*���V���������~�k��vÜ��5�vJ9�NL��!��V{f���pQkOf&���֘.�Lw�<�`�Wu�j$�ᗱ����I�X�Q��Re,�n@����Y��W��%�|�3rbǲ]���l�%�&�	i/����VƳ\���6�?.	?�?C�PHz��S��V) ?��}�]���V$@�#Ϣ�c��ľ����VX���KL�oձ�I�����5t��İ���zݳ�,���7x���Z[�����Ԇ�22�&5�:.�	@1t��]��{�A��zh{��f�K���5����UxIy�{����A�.{�����{\�I�߄3[.�U�a"�"du���Λ�G�y�8���l��DW�3�WV��LHF��z������%��c�X�ç���~S�B���l��#%�h��t�6r��7���4� �8�.t���E9�4j�S(3@�j1�h���/Rގ�)�H�N~�X�H������e����MB@��M��l|�"-1	�Uk��1i�iA|�Ik��Q"��_�+����_5�P.0�����)�C��'(F�}
����⿍��J��%bd'�"aD1L�	)>^�?)̶JFwX�Q��Ib�@�A��sy\mo!��`�X�ұ᫛�yF%[R��Mυ�2�1ZS��MP��/�T`by	�;.�췚9��^��!�E���Ȟ?�JK�@�����8�dh�ޫs�M?@ ���gJf��t�r��o�޵ۥ:��@ �wH?,��QZ��|	����
C���^�'�h��%��=�$Z��5���e�T,;a�_0�2�;\Lp�I���"��O��Z.�I���/Y�"_����Q��|����a�m(�:�E���Y�]\�����A�ɚE�ʕp�"�&[�Z
9�7��N,���m?�m}��m�N�R��/��������'���ж����\Ri��2�r��8@^a����>���I���࡙�c\�ɂYvlw �`�^a��j�����i;g%i����KaSNL�)m���&@XC̨�&z�k�_v���"1�U���ڈ��ސ����?<�����gs�jD�o��\��}�Ѓg��|��"�_`ܚK�)��@/� D^ԛ�5b	��y�6��U�U�U�V�[m1��-�#bl2�Uw��>��M��p`��Zo�[��Z*��v�0CJ��t��G|�d�e�7�O\��Ѻ�
�| ��g���XkL�F�n���9�s�L�]B��Ds\�����wG'���8�U?��w~F��>W������J�Z�7�,�{��TQ��M>dnaNh������	��0�������Ctq��&��v#0��=
��������ܞ��g߰`	�ۄi����bu���Rm�e�&��j�Ʊ�4`1ޞŪ���Em�z �� V���i�C**� ;<���p��לó_{"p9��F�1&�x9I�g�1���ZB9S����
��rt�"-�u�^�]��Q���c=�p!Oퟓ-�'D�.n�^���'��nBQ�U@*�Y�iU��W䊼\���"Y0������!:K���Ѩ���R2U��b���C�><����Pn�B�����~��s�
\I�^�2�Й�`�N05G��&��t�����#���6(��5���|W�F�Y��$�ݛ@�b����ڣ�	4��Y3sw*�/�?ǝa�]���|��d�9�z�+^V�!�LI���6��9o���I�ğ[���ʜ)��Dz	�<=�-?4��K�O̶���O�-���ƜYZ�r!�Wqj�ՉcW��=Hn��r4��h`oB��B��8�����CsR����k��F�KJ �k�{�2���)�; �<����X�:�
���n5D�K���3%�jMc,s�b`P	7{}Z�I��j����cǏUL�)��
"�� �S+���#m�����݇���ߵ�̥E�*����R��7}�Jom������v��w�����:�v*�%�b ��^{��0x����Ɨ�`�~��:v,g�MDI�7yW���gm�[f$�ub���tF�r�\���&}n��}e�鐆��l���t/lS�o<R|k�������cQ����~E�`���e��O�_��{G�^�;_������X�u�C����_˳z��k�է��!�ǰ��:�&6��Ǥ���D&`_.z�O��M��t��Oݟ(�~��ɺ&��TuLc�Ė਌�ǎK�v��[&�#d@�{"�~�E�b�=V�(���%�= 뮇tm�,%mx��G��"�dl`��ƀq������a� J����6 ��07ML߲�Ɲ�@`~��U(��5�f`����v��D����<��o]M}/�!�� `qy+�L҄�B^:ۨc��uU�k��~>,q��G��D��H�6�'��ڔ}����,x���,�b]+�!�np���\����ǟ���P,&�0�ҴAF��!v���[scye�.t���E�� G�G�	O�ۆ ��Vx���'�Q��[x½�h��]ʓZwA;� ��
��3�&k�녂j�|��h�N�ݒ��T��'�u��p�C�L�*V�1���tRd����{�Q�-�У��O�X/<�:ws3=d=T�@�c4�x�[��j� ��	J	t�8O���y:�vOM,���=�%v�af�[�����Y�F��H�W㲨S˧�P�m=�F	�����/_�Hk��
mr ��_{A�D�L]Z���͂��J�KG�Fx:W\�>�kcF�b��9�tV8��*!����Ε���)�@�Pno�Ý�����'�Ĩ�ٝ���9m��ӧ\%V|�l�����>HN��֔�/S�쀈��b��۵���<Ƒ/��XT�Uq,aң�i�����J��!�m(����.$��S�B��S�*y�l+S�  ��axv!�����>�̓I�ֲ�r�-x}���T���VZ`1xfm[�S�l�YA�(��1�t��ƥ1?�7���c�bmgB\:��L��=��֒g�����Bx�q���I;�ڒ���\�&�Y7�;N�p��1t���Ldw|�W�Z̽�k��ȸ�sع�0�r���ss?�wI����h�m�v���e`�0��g��G �g�<�&z	����eSV31�#>�'k{O����V��`^d9��m�)$䣣�q��EF�jϵ��I�����4�e����4���CF�"UѠ��麋��7���qa�)���$�C����`����k|�Qp�����ƿ��NÅ�T�F�v���5Y �1j���0O� P�m�}���>b<�	��R!���a;�,˕���q	�ܺ�@!�r�́P���ɟL�5;P����qu?Q8���!7�nS�-��y��e��ʼ��zi�L�.8k�Ec �0��6���T|� ������];��������E��p"�4W�q���Iݵ[2��&���W�-�����[R���_va��=q�x��y��
E"��!��Hy#���5Κ�Q�\�)c�IG�L~�!߰�}rϰ<�>L�@Bh>H'�Hߦ:����t�p6�Y  w�^7�O�K�(Je�f�S��Sȏz-I�����> mEpɴI
���ʮ�z JK�7S�o�dL�^��LA��%΅ʜ)ŤH������h&}�����F�,lG�8�`�Q��^�!懨��_��9�*qP@+��Ol�{�h*_�-��V�"��7�=R�#��>S��-� ��<3L���af����"&F?�s�Mڑ�����m�,��lc��裉�&�S���&�'o�����t�ؘ�	����3\���̖�!�XTpG2�d���Sb�Q�^�=�˲���:d���,@�>ST�����~}��h�YN����}W��a/.���O�Ƃz�Tf�`"��&?��,*�_y��Ft��d���s5ah�������S�<��oq�P�d��<����I��i��ܔsշl7e�O!�{���n����n��D��[�֣n��2��S:�6Z����_� H���ѐ�����^ŚX͜��fͷ0(�K�Ӱ9��x�C޷�Ų�W���\f����<��ʺ�Y�����P��U��9z��E�zd��'̙����w���8�-����-��\C��i�����*���;�E{{��T	h	��V.|�4Iq0t�¦���Bs�c�^�*1��Mt|3�R�+e޲Y�x���Hq��!�d9y��{_���Èi�Xh�	j�)A��ÒoJȋ��y4���R1��g�xuN:������p�I��"g[��3�6
����yGP��C!�����V�����uS�͐���jzQ&+�DV:k���r�H1� �Ĥ�C�6�� 	�}��WS֚l0HyT%���jޙ�\��
\�/TD�q�9�d(���h�쇺<�G�7L`�a��&��Z��:��"��_���'���+��\?�>�P��/�?��άIu�[��M���h��tpݗ��Y���\g�-�Rc:A=����+ր���o8,\��,�v]����IJN������ȱ���T���<�l$�i�U�}C&���Y�B�,�yl���&.M�k;�篥�ϯc���F��h�TU
�T��,	t4�1���ȩЌH��6Հ�OI����o%��4�,���r����s��f^j\du�G��)�/��g�ßB�g2�	�5�£��6�Lx�����+`h����k�6���Ƴ?�Q����ݯiـƬ!1�阎=L�;�D�!%Ƽ�00g'h�ʹ7��a]~�^�]���S ��㝑��@�_�dM!��J���Y�������e�8����(�k���0���O:&W�6T@���C�����z��W!��\����1ݦe �Ww��,���o��s������D���'VQ{�Q~%	ڜB×�skQ1�%*������B����҈h ���鰂��EH��#/^/�ի��H�����g�Bf(�e�i�M��V��@�`�NթFkџ'�����m�����s�2u��N�O��b��=�����h��f���܂ �A]��4ܘ�vL0@s?�&H4/ke�+\�H,�~wم�`�@<��v�^��;=��Pr��D@���	�X9�p=�9�CX����Z�T7�>�yh���4�5yA���oM�B�:Ć��ǏM�/B���=�����6p��Q!���tK"I�m�)�D�D�}�&1��z��u�_=��1��F��	��4{"�bt�ݕ�)Sl�|�x���J��H!�
ʭM�[-�oDĉ~�����jq!�3�|f�s*�($�)��,�XA�K<-��h^z��I�u�8<�e�ՕN���S�̽�4̔�"xl��_��b��T,7f?btmR$^˴4Λ�݊?�����y������i4�iD�?�@��}�9�e�!����ޣ?*�}�I�▘*��b�1�"�C�x9L)OoK���AZ� ^�X����إ|���� �����#k&Rc,?��En 8zE@���q��(�f���|� M%k#�s&K����r!��n~�̿P@�`��0H�!���uUw;\���<�q&��=�����	'��������B�� #��%��]
u����#�B��%�F�)�`:k�Y�x�ܖ�J
5�?x}�N�F' �I�6��h]��)N�u @��T����xċ����/�E�E@d�XJ�.,�eJ�.hX>�ߢV-5�\�Į��XAl��x��Daf6�h��>�/5��a����z����~ԶL�/l"_c���?9_�rl��LTs*��o�Ry���m���;|�Ё��R��I�٦��^�2�ͼ
�{����?].�_�qZ�6��M����S�����B�RO_�g(�nmh���5�i�o;h	���	ߤ�A��#����Gc�{r�"X�m%�a��O����C�j��}漁��=�p�I|w����-Cg?n.a��xi�	�/4�yZ�l�z�I!�3@�T"z����,Fj��%ⰵ�w0G
�	�Il�"��Z�h�Y[v��+�v��u�Y.���Dr���.%��P�VW-噜v����K�ZZw��5��}�)[~����5�F��w�� ,?��ۥwI7�GtKV>�O�}N�^��� 㳛�[!��:x3���e�jDMǮ��ǚ&U{�j��2�<Ot�����#�[o�/�h��':n�("/f��O�#:�N3j�\���ߕ1��~��xl�P��ݶ���/	�/Nz���@L��`@rˢZ�J/T(�l+���$~=�mm!]1IY�Dm��,p��W��!��X�_Rn�:.�i��)ŲVIu�pR۰�"?���
`��6o�D��X�}I��&3�?y��3�8 �T���(62M:њ:�r�]�j���۞����vx�!���_��H�Js�&_W6 !�����"O,�h���K;���K@
����_U�;L�uF���¤����N�ϴ��ϧ������o3�.����8i�⳨C�0�fF�Hy��*����gD�]��!��� ���������v�L�jF�[q|+���Bc#̖։t���3C&�Jh3͆x��h����w4r�-��UL���F:gK{Q?D�,�m�I�8���UY�?��c�ԘږB�+����5�����
��
��T���Y�^�A2����t�U�ڌ'a��2���a��TbN�얛�OQ~xP���0ҧ&���Cw�V�ϣ�k��1Ɇ��;�0�$.6�J���U;N��X��g F�4�{��sFZ	�=�o����{��m͔���|��}z�qsLCH.��W�|��m�`{��E~�lV&��������"��R@�>i���&L3�=n�\�������fM�AI6�v��/})PIѬ����v�n���Kki!�h��8
���܈Qt���t����U|n �7���k��E �O�tCy �j�>Po�#��1�O�j��|�	�RG}q��A�u��򟈄7Y�\����mB�R�3M�^n����6��Ы�ߘ��%��Ii��^�*y8�
�LQ�.5�	��x-U�� ��#U&�J����"��&_����u.93����Ǻ�J��N|v��Q7y�����\{=�-�'�>䡇nU����ߴ�VÊCt���3N�x5�����Q�HS�����і��&ԗu?'=��s��"(�������J��z�D$�c%/�T�;ER�Z�# 5�0����t16nQ��M�!�0���F�՝�#�^����ñf�J,�b���`:/���"Y�Q:?�N���k��IȎ���ȞqzȠ�&f��<�<�G�;)������U����d|f�fTL}�G^�*ð�J�g�P��mh���"�&�1,0�ɫt�T�D��b^�h	���e���p��B�M�FM7<�B�u
9P��PcC�*V �A3*�^jt�C�7����Ժ�q�&�����³�옉Ba(�
�w�x��3f�����l̼+�ؤ��P�HQ��<�%չm��X�+E5�3��կ�\xOx0��Jx�w�y
FU+�uO���k���׏�^�>������O֎h���D�`k�{�o�Dw�5�h3l��s4y�4�嫭��F�9��q]�!�΁���c�z=�s��*Xr6$�\�v>��5u9�u;14�޹i��:p�M� 󘶢d5"�]��۶=�9>��DaO����C�Hҟ�I���6��( PN'-=v�vqB�oM'���	h�`���_�0���&�C�`�~g��fG]؎� ��XYu�P�ocU�X��Z��M����kⲆ%N���i����iW����j�����}��Eϧ2��!�X]3��0�`B!��;�0�g_F)�ƘG���A�V3b��;|����ꇚ �
�&$t��άa�ӊ^ƃF�k6ޤ�A��  )��(*3aV*�ܭ�4��1[��e�s�@kÃ�\,��p�n���B_��;������
��lp{��;_m�։Y䦶<
�t.�Ǫ�τ1�rJb���F�=����vI\)�[tG��3��r{������/W���=���.b�z�F"�p>]w ��M��l���ʨqa	WÄ��%E㘕��o9�!Wt���I7I�g�	�~u��>:���"�x��ӷ�!ȵ���g�EkQ��>�Q��L��5���L�òO��	K��h���@��נ��XǊe����EXi@z�z�+�� F{p'�~�
L�Ѥpɫj��ΰ�n�,+��$I��@6���D�Њƴ.��t�V(�[>��qG���R,ͅq�g���F]�ބٸiT�v/8w��3�0@Ӣ/N�3=�W�`>�Vw����(D�J!Tu%�/�M6e��g����]���i2"�.�n����ȿ�e)os��#t�HSϷ��ոը2���*VP��=���#�C9H���d���{ �YtDlË�~�P?O�[vUF*h�.�c���1,({j����N����+�}�jalm`������5�9q3�,�a�Ȧ,�R��@?�rmMz��v_5��-o�I�vp@��ʴ��5���SSE�Llh�����8�P�ܬt�s�ꔧx_�BF0�6!��LB��^w�K'�<H���;�Q~�hx���s��Ԓ?A��fznx�]uUs�X/%�����X(�5[l �Ob�9S5EY�)Ӻf�5���'��d�[�U�Z�����J�Nu���l��$�hS���S���^�j���i������<(�k���c�)��<��h�V$�3�շ�����Lܓ���/�U��2z�^�朙�[�MX:��=o��`��.�q�3�c�F��Z�OPJ�Qi���ӟ��+W�Y$�Q$���O�n�4�L�+X��o�ʀ�J9c�3���=�*���M�����Ss�SD	��'�\
�&�g��zE��
K���d/"sbS>��E�븂���ŢfR�3��GX�G�����p��8�H�&b􆧩�Ĭr,w0mƜ2�uDz�,
E�¶��{��՝�F���L�<} �B��掱n��w`)����t�{�>n0J� &�/��C}G�qę�E�!ɻ]i1�r"_ �d	ډ5l�0�¯���	��� `v	����9�2w$N�i���~����s�Nݯ���ˆ� �-dBX¸��!������ٚn�	�\Sv����`��3�W�8�Y����kY5���{�rP�X�{��o�0xS�W,o��`h��UI.��MWl���#\�J�m;*���1>8��Q>����Kj�����7.J���T�����؅2�xZ@��gKX���s��N$X�a�������b���ZM�]�{��]^���2����F�se�F�����s ;z-�o{�����>����X�7Ps�ޔ���[���#��������&Q�O*�s`�J�Y	}��1>�Qq�7Y��~��R62�&q�l��29��E��ŦzO}�X��Z@X�n�t��$dG�DH�_�M�~c�P�4� �{'(E&��\�x��*	ȷ;�8����������w����4Ծ�΂+����Sϲ�R��ɓ�>U�K����+�{H��L�a���b�� ���>�b䲦l9 -��-�B��c���Sg��\���*�.��W��J�V|-���Y�S��K9� �(㻰.��cZ����WNt�n�L@Do��9��K���+Q�����J�ڭ�����lqoe2��	�k��V)gU����L�F~*p��}�[��V.�8� �����XT��K#��솷�%�_A�s0(QI�(���F���`����%�\H�)����:U�0g;CVTkF8��3���&�����pt���V��÷�N*C*j/mRf��0Z��*��Bi-o�|�rm�z�]�K6��$�l��4R
;�Z4�Ѓ���<=�N�j�0(}G/�Ӫ�T!vl<;��u�i�FE]�u������v��?��V��}_�SN���r��ٍ�Y�3B!_�r6���p���Y�,5}���ǺGǞ��(_���W�M<���)t����O�3�	�#��;9,�Ϡ����O^\�D���~�kE��xp*d�U��C��^�l�
f��X�����݇Ȳ�"����J�� B�S�I���'����=��{�	��]�	8c���oVY,8�缊��Б�����Ū�a$��~8�'W=B�U�k{�~^R=$�!ʏ��$h�4���~t��(Z�U�LJ寧�$˪�&�����UiA0G1�ށ��0{雑��v�N^WW"��G��~�V�ƸK���n��A��i��M��3��x�@2ҥGs��&p��ܫLB�ۦ���0dd�I+W/��d.n��3����/I{#�&��Rt��2���R�̨����X���ힼAx���@Ì�`q�)��AS��.�HeM
��Ij?�B@Km~��,�"�	# �R����{ ���ԍPR*�O�;�>󱮌Je��q3�#I!<
�*�73���#���>�� ��4\:�Q�S��¦!�9�4+��d��2u*8'��
�X�IU&�'��k�Y��(���������zN\�;�ؘ=�{g�ÀC�r��k``ɀ�e1�U3�-���OV�v��_l��xl�n+�̷������cQ]�b��~e�c�8����kp`ul��4��5�>���a���#�[�m��1�F�,"1�͓���9do,`��;�Ta��>M�b;�~����爜����+8pu�Ъ�?��A�-�/�z���TZg�=�T4��bB[�)���\D�ܚܡLS�:�"�7�!4)#�a�P�U�ͺ�HSGD�a��k�gWTC�ʧ�8f7�P���x��9}��,��EH"#ﶏB���*�i;�,��qw@��Ŭ'���]�)�s�2�*;�-�{���Ǎ� g�1���>�n:�7��̃������4�93�1�)���N<Mh���Z���{�ηH���o>&�2��ćL���+4R�x��9��x�(?l4��w����&�x�Q3�{=��:4�[������q�-��1��θ'e ��c��>�D�-C�/c.�	R�Hy��'1�ᡇ~�"D�i n��ga�sZ��x0�]�.��o����B
T��S�����(��=�1a���|#��E��L^����S%3Y����yWBD���&J��,���_�ٷ�e��m*���	�Z:�t_0��@��I���c.y?e�\ẃeW=p�LN�j�(t���Q���l8���sWaE�}G� �ck�����D�s�}�79�qUn����z��	lZ�1G񁂩�Gn�n����L� ���� ޽� ��G�DSa(FU�(���~�:��*�I�`�&p�x��#�+[�p��/*	�[�7Qa��1�v�]�����*!�f|cV�_A���ߓZ{�#��t�4�xu8��⩦|�Ǹ	S�X�H�b��`P8`�-2��.�G��A�����]F�z����*������������)��(��� �MǇz�~�5�F��<�}rk�yګṍٻ[A�>��p&- � w	d����P�}�6)�����l͡��o.��;D��~��/��{-�[ueM���:��3
���cH�A��8KP(qx=}�\ɻ3�v�=
]d����(	\�1b���ar���΋����6��:�~�//��6�����
RIw�=��;�AyW�b���$t�S���`�k�.���<��ms���Z_�8��ܗ��0X�A��~�������Zڡ��~C�,]W̗5��^��r
>f�Z��b���Ѱժ�a����D��ߡ���g�����dՔ�UW�Q�:��:P�r�<%q��ߍ�v2��V�/�c�~��٧��(z�Sj�a�H�ٳ	�~��l.lQU?�C�K�<�'c��Uq����J{����µ�w9P*HK�g�1��C�!k{%vB��;�,�ƲN�}-�7t�5��*�
�u �)���!-���hl؂�IKَ���^�j�,Y������j|/�F�����hƢ�t��W4휐Pl�b�����1�	w�w���G�FQ�k���s�������+u� c
���g� ����w�(������Vp�B�}����������R�"�p:��-�g$��Ʀ���?���Չba9���/�fSYaF�hh��WA���bfyN���LB
?���4������W�j���gP_�1� ��M�S`t?d.7��� '2��hǶ�-Y��gvl��U��sH�H0�l!��[�7=H�7�4��uB�ێ+l�2����	6����G�e�<m�!������QrU�	�&�I 7a����t�x)]w��������+��p���ܥ�K���[aɩ�3�'W�����|z�_�`���/��̹�1h�0_�=��ũH��
���$��S
�E|�q�f?Eҁ��V�]m��%5��_m����4@�j�k��{z"e�8^�11�(��wq0������-S�8�܄��S~M5\��ʩ�-~P�V&
����n1�n�/3��ڜ�����d���k�^���x��nԶ��͇Ah�Z-X{�&�$j�S���	c80��� �0"Y��=9�+p�Y:�,��j�+GY�*�_3����,�z�����ϐ����R9փ��Xe�o*vh��:�>�d��۫��}��3;�gA������]�g�����<!��;��?��p����$ �Tj��즣I(�o��>�@sKӆ�"R����@2j^���6#�G�a-oP��u��܋�����b4-�nx�-A��d&�j<��a8�u1N � =z��;�X~MH�U8k<56<�T"dBƊK8Z[`�n#	��x@=�G$��)'�
��k��>�}W�Ҁ?��>[�6%�H�O�2uu��~�� L��G����Q�s��o�m'����K���_nB�ĸuv������߂qq�ec��9��ogv�0��lG����DX��_��XuJ�Cb3a��Y��.(g��\)�ƚ'��-j�"j���̜͸�Mb[\�i�4xM����2sw���?m����O1�X�� �������s��n�\B��d�B�qL�H�0���\��V)c����ң�:Iw����f]�,�Y��R�^��������|���u�p�_�K�u	s�{I!D�"��uD����"�.k��,l+%ۈ0E4���^�MMY��-��ސ:��R���p������o��'�A殈�<P���+B d��{��g �������t�)��h��It'kJ�򗼃����F�\�ǛO�D��B2��J�	哒��	�QO����T�UjӜ�#+��E��D�2�SJne�� %����	��U[|a󆘻��+E(���(D�G��iQ����In�-�g��G.�c.��g�7t��&P�d�()�����zN� =��`i�8��L�^�������n|��b	򌷇ϖ᝝;sdӝ���r9��Ǉ��/�[��$���אx�A���z)�S��oz����|�v�1�%��kň���?��������$���)��~x,2�E^C�� �F����Ƈ1�6��[�X��� �zu{g��QI�ƪ�,Pd���>l5�;�ݵ���E��n8`�Ҁ��`�%4�h�*�j+'%Z|�����6�����²@���`�4��T�4��>�a`(��)W�B ����3\�4��OX���q��X�A�f��˕����:��>���E�S�
�<]5��Н��W�P���f'��W�?� r��;{�"r�!�O�Hi>t�8����Aq?7^p9�b`�v<c��(�J���ԥ�Q���Ft�c`�^V�fg�j�YE%D��w�>��y;θ��I	JS�z�\�g�5�1�Ԟ�^��`�ؽA!��}�Hn�S����SM�VJg{Z}�8O[m��+*�ʰ�-(H���M�k(�'��r�A��9�u���$E
��5oZ*&&23�j��)��0*:�<���&�����{�N�� �!�D���z��*Xn�N��5��n:S��&zW�HȵN�I�C��ZYڱQD	��矐�?`�A�cV9`�w'i�л���J���>P����qS�DXM"�؎�r�:xPjf�mקV <�b>�oN�g����������/��3���K�9JgH{M̛(�"V	w��~A�I��-'�S\�G�B�l�wX���Y]�\��l�s������H���B�5�B'!G-�AJ6��޳���3� L�^�#]h�#��%J��cHbek�(p�sZf�p�}�A�U���N���]{��葉� 蒧NF$۳tW�h�ΞyK���TK�:@���U~Ԕ�X���{^F�n܋�Ub���v(:'N���05��,jQ-�x��NXm���G��M9	����h��B9�.��#�
�Ӻ�y��D	ox0��P��hu	�"������ B�`���O�Ͷ���V��9����A�j����$Ρ�
#/>�q�:P�^T�Pϴ�g/��q��>�(1���Í����$�,�S� vC&�U
�4X�B2�~ZA��~����%G��T�Q��u��
u�tf�K�\�坃�;�RE�_,3�<9,�Ёq@�q݊ۏg���.�}6��,H�oMN���%@c�H�p~���(YNt�Z�-�`�=bRغmk��1�v�����|3��r�^֬3��vsBz�ə_�Q�Ų��ΑJ�?���?V�ɇ+)~@��y�Fa����;���[��H��Z����J�Nc���3�Qc�A�=��2�=,4U�9�o9��ܬ�b�^UL��$هS2E���tK����~�h^��Q
�f�}����}��OP�G�],��~�>*b�V@R��Z�"���N�f��9���4�X�+��L1N��u��됏�/<@�-����g2r3�D\\{H��?�TE�xɻ�b�k�2�ɥB���
%�6��~q��3k����Xv�����M$���Q��|���������'�w/��a�{2�����1�ә1���J�rI�����m̏���S y����_�w� ��8K���ǉ%mM��-�B[�؍M)��!9�����y/=q5�r=�v��w]*7a�ҸLy��<��MҐ�&�(�(h�o)�ܿ��W	6�S�����Ir��qp������%��3d�dWh7��ԾTB[nd�]�/o�=���2�!2�q������XK뎓�T�Ƚ/��f�P��7R&18�;Z��Ŗ¥�nJ�\Vs���쳎��ks\�P&EwA��e��nXk�'��v���%��Y�x��`�=7U=����Q�M��A ������*���_�ʑ`==��/MQI2�k=��j��<jF�k4tk�{B�����e�Ko�e`J��>�ԃ�Y� ׬��(��T�w�!�_$f���WC��pD�O���(�6J��`�������r6�<�RK�!:�sY����=6�!|�i1�Y����l+�1�e��/PG�s��V�q.�RD�pkB�����%a�r�$�5Ct�[l���Wp�WUS�Kg�G; ά$��?������1_���s�Zɬ�F&�%6��i�~������-�ױ�z����4p�P��9���L5%J�3FU�M�v�(�jaW����6fQń����-�~M����YC�J��Q����AB�u�U�ō�p�Ilʷ�@��v/7�|�8e��QF_�ξ�4<�	�t<�`�7��pJȌ�J^�K��fEDʟ�S7�:P�p���TK-ٿjO��0�� ܁0"�����TW�˧
%����r<9(g�t�`Z�A�b�Uc�ʃ��u:\�;���`���Jw��{F�� G�X#�������ed�q��ҥ��Hvn	����w�S����%�eݗJ�x�WzH�����rP�)l�}�%�@r	�&�V>�c"g/���Y��y�:+�5�����LE���2�E���'fF�� �K��x\�Ա!ɷ _�hW�R�&�"��X]y�1�ŭӆ�� af������5�����<F���Q�\8��4>NN?��X<��� �qf]N�Q��F��)�эS�虤y}7zb��I9��� �{�{��^=$�/�#	`k�*`��4��)��0?4���[Z�*�v�J��y�	��^@��T�\���#�VhS�+����A�z�
�>(�zmhy_�i�:���n�����H�(IO'/.��e�3w�j�ΚfPQ��AF�!s����guDQ+D_-�AgD��eܗ����8 �����KҺ�_/e�|��|�M�!��f�Q�u�P[NN �����I<Hg��*=�(���O�A����'S�� ���*�`� �uh�|Cw�cK�Wa��y%��"��ڣd�qf4C�c��0@�"ď�H~�茡��g������j��dL:���MV60w��ɇ�m�'��N�o���"!��9-�P�4LZ������Q���^p�!җ�;˶�,�3��tt'q2H&�M�յ�|�'Y;jVh
#ͨ��۰���:�T��8dRM�E�pkk�7�;��>�Z�$w
c�-�8D�f�����)>�u�n�rhR��K��e'�Y	���&�М�1����Z�E��V0m$`E���䛋M6��CS�]�8��nP�)��	����B�[��SQx�ya�H��L��BlWژ�+D��v���8��$�+��V�^�Hi<$	�;Bm��֮�5--ݜc��������vM����gG���f�|9Ԕ��h�$/4Ѣ��x�iF�t�%�\ކ ]-ao%S�q+ �Õ�xh�M|��G�o�.S��
��'��T=[Rl�ՊC�ถ���w.���-K��`n��y�zxV�R�7�'?��V�������i�&,#�2���a��޺e�*3k��,b�j�VLZ��u�2��U4�� ����Ξ1;��cF�ԯ>��1ߍ����L�_� ��4S
�Q�
��;a�:*��O�q�{�ρ���-��!��'�	�l7�L�vc��ie8�
u3��C��������0�|�'X���
t�	`�m��EDt�%�(�t��yF�Q�q���$-���r��4�s��u%��T=3Y$~W�˷��odˌ��E���W����3��c.~M �و�H%� ��Q��]<[4cYs_�g�,��%�k��S*?��?j���L�"2���=����t'/�>:>~�����'S�U��P:,o_r�K �)IX4#:'��=T�ç�՞21�p6����w�%G���@���Lq��m�N��Y�֖%�D�.�� ���&��%�)�du������[,aŗ�C<�g�rι��/t��aJ �����������4VD4ޕN��	=�J��G��;0SY4���鷞e�INT��Y���U&�(����[a���v��%'U��`����y�.o$W�����i�tm>{y�B��c�~R�jz���s�M׮�m�[I��o�R`����NUC�~��Oq�!^%�5�d�����y�R]>�_���+���T�Elk��
nw2u�gx��/x�\�ڮ������)�$� ٺ ye*��s
x�}�d^��'���a~N�֭�\V���>�%ӹv���5���<X|H��挶e4�R��l��v�V�P�!?hE�HK�����P��ő��!�Jg?%���4���%h��7k)#��)G`��� 鵎��u����7x�_��{�_�}��1E> ̝t����{�ۅ����Ӆ��UB�c�3I�H�׶���'n��$�O��F���UX�7�K���K��]�i�4@����f]g{upM^٨z�f"#3i��0D�S���ΉI�ε����1`^�3����[^�ק�6��	�>0�a��������Jem@CO�5�zU�Z�;�!^��Iы<ʗ�Ƣ�'��C�2q��q�}(r8��Q�{�������B�����y�����p��U�\`q ����dݸ�R�`e�)�zJ��<����� ��+D]n�$|�{G�^Y˖a#?Z���A|���Y�'\\�{Iݞ��{��?����~���5�y]���B��Xl���`�(�mnM;�B���ҿZ� �㧯���M�%vM�È��U���ٵȄ�s���I<q|R��Xv��z�9��8?�g��%r�Ț�u��;�hkI�����RZ_����~6������-�_A�����6�pCo�y��0=f�? �ΰP���`���Wi���$�ՋG������o>�{�^�������<�)�kȟ
������-s��t��%:�9�pk�O~�)��O���?�Ή�tƄ���:����^T)��,�/�ih��D�_����@���l�A.����w()3+h��ðyP���ME	����書#�Q��7�X��ָy�3!&�_��F��^�BD���v#�vi���5��V�(�#�p�"Ml�OH�,{]?0��q�4�#+8� ��`�#�l�c�kT�U���?��!��y���,���B�-�iA�@�6�V�7w�򂫂��J�:`�Ý=�b�ѝ�x�cb�Uͽ�Yڌ����*�k}�嚉�x�V�h륅8N>b�Y��u���&Mg�x��,�H64Ĳ�i�>h�޶��y|��Br��#�|	�p�����:t�v�\)��f���_f�j	t>���ܯs�_(e��3� ȴ��d��X@����\� ��^?�+,�th�«5U��\�q�,�p�����zq|�U��b��ے֡���e�Gl<>î�˥DCU���XԦ�k���������~Ug���ю@3�Pb��o�Ԁ�_����7�IŜ_������)r�osh���z��fF��񗍎�Qp"DJ�|�b���;�ж�����s��Y����8 �:	 mt�������tLl�����ϛXÞ���+x�wW^���p����d~�.��l�G�#��z�ǣ\�-���[���qRז��U��`y��o&é�-�D6qu�5Q�-�:�����&�.Z{�3���B.�Yu�Ftf�}�Rv��g~zsA��L�/դ��!�E,�;�����"�Ϋ�2z״v4�|�|_��[��pz��R����Fph�/������wkO�S3�������:��_��ٽ_�����+߀>';=G�#�~C�z62&{H��V��T����Gv��Am3MC�I���)}<� 4��jE��i�0x���t;�@�g�����'�v�7S��I߁A��T��"E9̂u��s¯���|�(��Y����B��9�0�����9_�(�xrM|���Ř�E@�W�i�>ϔ�ʷ"�t��pB�J��//F���_����G������f�J�
�&�s�6�e���w�mD����Z�٥z���~O�W��r�|��7H����gfev���D��W�b�>�U�ټ)I�N��F��{؏p��J 3�s$(�0ʲ�u=�'��~��p��!	�2��XDCs(�ZO�mj�5�e!4��-�_��8i�k�͉i�:��C��� j�q0>>!�HbG�~fӝLQnu1�k�(�,���4o�~	-�zГSf<(��p9H����L{�k��)Q\�{l��ƌ����<�1l:�z�}<}>(�Fޔ41�]��k�)�0��Ӵ�Ͼr�1���_���$ɣi���3�bF�껐ڳ�eG�`���^�n�f�	���t�3��d�ƀ�� � 
�Ɖ��Ԓ@�� �O��gR�*�ħX�_q�m�'�`��ײ3�J��9�B�_��6�z�`�PF�+�X&f��3orl��/#j����_Kwk֥�hNaG�$Pg��w!����>�X�LӋl:3F��/fR*�W]���b�ظ�xB�/-O��`�eu�/���6���"hy; (#�t� �0�ȸ����0'-wo]�\�Omd�L�p.��4	�)+�L,@)9��-���)%hA.R���8m�t�Fm����ھ�ɺ�~Pأ����Q9����>[��^T�Y
2��O�/����P�:�=�����e��J��E�No�i�	�����WOطɑ��0��P���=��,y��C��I^�D\�fj,��=s����B�%H�1B��?���>�j?�D�̍(!��8[v��$Ũ߭ d�u���2�p�X��D�T����E7������f���%ۍ�U��������P�e�#aL��fA6���82h5�1MQi�Ӻ�@��\�|��J�Ƒ4����QYZ8��P	�����7QS��ON��{M^/B�**�����`]�����p�_�o.����������3Y�N��ě�U{򉱍��eA��'�@�&�����L���y�UÖ?6C<��Pl �b�^�,9%_������;��8�r#��T���%+OP�H@�j�w����B��r=�'�k���z�E���%%��v�;����&&*>+lC��"{�aFb�D-�L�X��ˣ}��Aז�����>2�ZN�3[*� KT��M��i�N &�m�+A,�_�w�t>�v�r�|����(��rPO��x陒�f�ǜ�C?p����%ӗ�d��瀨��V�r�+�"$�Ws�����~r�օ�f[�O�)!N3�xn�	�Μqhg��6:��7�K�	#:�Qڃ��#+r׸P�~.w�w=��cde�[[}o������t�9Q�f�vY�-�N�.��Uʹ�l�J�}� 4��C��G������*JD|=�C���Le-�"؂�\�.��_�bFi��rj�yg�E	�x#��4������ɲ���|#�M���h4��5�p�9����	�j(����E��NG�϶�g�\�`�/��}c:���#kM�7�>0�nSt_���b
'�SJ�;1��M�2P%3�Eu/.��o����ϲ�Zn��JR�Y#���>t� ��X��ݔv;BW'�����s�ǩM����ۗ�(����HI�6S2�`��gT��>}U�>�Qo�G/�8��7���Rd�@�hӱ�0��W�OWO��o�Q�ws�]��D30V�2�x���Ә΅1ǘ1��G4{it��F"IP���rȤ)��}��~!�7���5�=]����h^E�S��<S#�ޱ[�5Z����lz�d�T�P�p��-�F�%��	� L�R����kJ�G؁��9|�P�_����8)�������;���'���a�ֻ�ZB.]�Y�[�ᧈc�M��K�ś��,L�Q�^rлA�x�Ҕ���SqRW\�:�|���W��dN䏕�q���A�0�v�T!�NZS�b��HZA�CP�Zv��g ��y=���G(''���77�G+U70�bq@A����<z:�&Q4�T�e�؆����P���Lu(V@;�(4I͍bı��V�y|�_|�!�E�_9�UK���)w�u��,�<�ًMC���I�54DcǑ �	�g������vb�o1,�� ��ɺn-p��<��?�<��B�8����a{��<���6
�ir�F*�=����A�ۖ�I�N�4���uRl���X������W7��0V#�i�J�miL��s���Z�s��L��ذ0��'Ւ��}g�b�c����p-�g�^{{��Ԭ�!eYE+�]��M��v:��չ��C�u�N��-d���J�|~+�K��L�YM��;^I�� �z��(b73J��۟t�gN{���f�ɐSnչ>耘�������8.�#'�^�V�f�Ur�}T�/}ū�,g�/�#��d�e~�;&-��Oy��̤MWKJ�'g)���+�`��ݯ�L�5ٌ�}��Qm�Z!����ۡ��wC�4f}�TF�w澣����q���Z�|�!��/�Kί.5��r��R2ZN�E\�q���9i�o[ ��NP�P�����O���vD� �e65ۈ'gU��lP�l:ɬ��J���Y&Eٍb�e�ؠԉ��~��R�J�n�r���v�c;\�j�K����
�ޱ��PT?T
��G k����>nd8y�"�LߗdUduD��D�w)�'9z�
�d�6�M�%�G}
p�c�d�Ay�	ǌ�ƫe���[�?�3���S�	�'����W�؟�+�F��㸆+pk�4A� ��Ap���|#Up&}���x���g�g��%菀lm!¸;�b���[�/:��*숔O�2jFk�]5b/��4��n?=�����z#2{|�����a�x�b�pj�	:�܁D��Ж���Or�������L��9�d)�M�(�H����6P(r�nx�&	�����,���=�_t��ߍڷjd�,ex�՝R8c��nu� �l������Ū�ѧh����A#l���q��v^IE�:�C��'t��2v��A����dRo�x}����O��E����ߚ�Dv��ߚ��֟*���R��
�mÿ�p�h�i�?T<2�[�*�~2~�:P�!�;϶R�<B�6����׫UpVoN[��;�a��X��m��0��)��= ���M@t{�P�S)���OC��ৼ��� ���ŵ��	Śg�5Ӆ=zΠ��``��ۦ�)�{��_	#��@����U�+$?p,���}Kêf����Gϖ�a ��Ź�5 �"f�$���u`�%����/TFP]�%��$�<;JN,��9�#���f�!H2u2}ыА��7+ܧÖ�GcÅ7�5��� h��}e����x�����\y��S3!)��܍t7H�j�J2N��z�xC��@� с��^=���e�2�G^�����K �˦�<U��h��8Y�n�� )F{�8�-���0-#��v����;��_�wNPMp~�=�9�"&�f���O�,b�.	��2�T�֓����^�ްe@׶�J�e\���y�sӕ ��~%T �q�=��*�}��񍁷L;D�ѧ�G�����Rxb�XQ#�g�5�ˀ�w��LF�'��0~
E���@.���X[���=�3qMߎ{���"���-+��~�۔�n��.3��Ѐ�5e���RfB+����M�P�}ڑJ��� ����9������E𜞧L��L�Zv{u	�bB�Ov�vX��L�g���a�@�j��d�6�4�_1&N�b�s��3&>?��ճ�[+hݥK&'��{U෋ݖs�D���v��:ĕ,=��6Mr)_�WL&M�����dn`~��#f�ƜWpT�]gO~�6��Bxo�57���㦹�j�ɷ���(R����	Z��+S�v�~�U Q�m�Q�ȴ@�
�D:�N�^�L��F7ߨ�*������N�h�E���R�2�}|-[�*�ӕ�����:�������E3����$ȟy�H(��0�I�.�;����� ��$="F��
\9p����Ǌ��4[�@X�v���R�	$D�a�VcPVvj���d�|U'��_��с~�6_��q&A�%m���ҥ�s�:�D�QN � W�da}���v+�]5��5�:�ҋnC<y� ]��\;�L}a�i;�KOp�p;���Ga�~��`�LlƦ�S�Q��Y��M�
�E�r��9'�!N���ۙ��K� -(���w$t�y�<�Cc�bNAUӖ�eX�9x4Q;�hL�9ٖ��5q�����m5)5�4��v�̫�N��岣�n�[<�p
Q���+�?���6��QIW����b�L7�I�Y���"&�zb~����S��\8�D��X#a[g��B]52C'�h�n@�x����SW0[wNh�7��b�s&����4
J� ;��mV=ܒ{�nҩ�b�u�$D2�L�\}�^���&���uv�k�;���RJj���XX��q݃N���IY�{9!�=/����=�2�H�'|+�z�>P3!���H����|
���ݷ�Vz�K�镕�
�}eJ�|E�Tj�Q�xǢņ�-�kfNR%�'��%.���~��nIX�!��7RkeYQ{�ځRB�ė5��!�y��b�����^�@R�hD���4������R&0Ć�Z�W$2C��*���v�ѝ&i�׸m�<!��R�u@�D��^%�@GFT$3dJo��|$��a%�}#Ԃ��j�Uq9�OTT���Eg�[s��P�;,� �<������7R�p��H�#�G���o�dD�������]z���j�*@p���<�W��q���L����Рʟ-���hdd9SO!�GLo�H�%Jl>�-����)5��w�&������}4�Rrp��*w��ě��a���KF4���0� 7CZ��.��A1�Z�ϩ���3�c!H�-
�l=�.8�!�\[p��H+'���?@����W`�4�H�B;�O8�Zh�IT!Y�O�;���|�LL���I�F�1T�<����q���w��$jL�7RдL�y�
bҷ�\���?������=�vK��r�G�8�=�Q��$UM,S�9���3m2�z]:����M�|��m̭q:В|$��-Dѝ��8��Iſ9d��r�ȉ�E���gt3���_��x��;�@��?�y�r��L?�S|
^h 2�
9H5�&슀�O��= LT}�<��Ű}�d�0�YJ!�q���'��=��;:�oL�  
�Q�=@�����qZ���o[㩑,�5��>����z1��dw�����6�BJ�s�Zن(���2j��E�oH<Q;�%���o�bcx�7sa�+����'4�G�t�z������I���G�dq����Y	y���(�q���2�ԓ���8^��TT&)LX<l<�L�`��Vv$7��v��ݤ|�!X?4���	��뢷˳N�R{�aS�>uӠw�9Ij�m�SX/�`&�HuH_)�t�R2�C	�?�f� �,��ˁ�8���>�Ly]`R���X���WՎrG���!�e�����q߿�p8�*ԑ=��������Z�wp�9�v�c�Z#79s-��\®����^h�	B��C̛��Wڛ�Z�8���=���>�5�fM�3���ڲ��M�,Ɔ������	����䊛v���Sq��M�����M�YЈ,H��\��\��f2�-���
�d�In�Υ����-Q�${ؖo���P
�������wep�k�s������X�@�M�F� ��#���H��_�j��1x�o"I�=���R���d%#Ё��~O� ɟ�g��ZL��HJY�=�.U9�5aE���#?���v,V1�'*����k*�b�]:t6����mk����,�h�[ԕۿ�f~�b^��P�=l�<�,+C��NS���[�����yB���� と��N�l;����*��]�3�T�&p�ʇ�����^W*�2�2��v����B5z@�TJ���b�y���K��W;��wmћo�|��r����>�_J��>u<�n�7r�_sV	+�R�������.Ť���=��"��	щP�D7��ԔFA�jF}2��{�l�<H��u��TѸm�b���\�v�d�qW_��a�[��Kڣ�r��̉�1s�4m�_D��J��<��T����إ8�y��ܮ����!Y8��'(�n-2��b�}i$xo'��d���w�2��x&���'�ڏr��l����F���&�9��}c1N���ڧ�J��Ey�]+l�C	�02�g��ƺ�vH��^�n�G�E�cu��2����y`�_���E2�=y�h��.�?W��QY�j�7;���Z�c�8��U�e��+�,�z�����C��KU�>��DqB�:��4��g �����u4v~��O�L�e�-��^���+(%��d��2hMMXV�=�	�{/�լ��L�����;)�"�4p	YZ� s�Дs�;���(�������p˶y�{��i�ל|��X��\�O�g�Ix*t�Z�P����ۊ� ��1��P�x;�q���n��8�.�	���E�g\�'(�^&};��Q"��M�*4�g�U85<��O�dOA���
����G��lu�Y���W�A>c�8��U�_O1�;�⇸����r	��Ko�́	~�(7�V�%�z)v&���n��7�Fo������O�Bڎ�����Lg����|Y�"��P�D�@}��0��J+_���b47�c�x��!���%	��p�����VI��Bܳ�)t&�%
]��:v�6ёA� �_!|�Z��tX��oXg�إ(�)2%b|'��MOHRr5%Ӊ��[�qJ5yCͩZ���ߑ�V�B��M9�O6�7����,�����S�+�����JucL�U��J!�8���<C8�*t��p �P5��hOS�e>F�n{(-0Ip�K��1�G�A,�)�3��4�=������<3���L(�<������
�>�ݓT.6���K����~�8R\&~}�OP#���ۡ�#	�+�Fb�T։�����.�>�(Զ�_�:�r�Z�)l���s�mE��,|HL�	���-��X�Fi�O�g���߁[|čz-g��>��ܯ}������r�rj_��#Z I긩�^n�剀T�T?�2�o�x���E`(��s����0���II=(����X��^�1Ic@"�M_Q���Z-������rU(d��0C�t���3�y��=���^��F���90/*��G��xX!�NB�aB��!d[��F�!NR�̛gh��K�;���2�mͻ Sb��q��Kr�I8�%2fl�`5�,���g���gO�N�ZV��R]i��ŏ�?O�X;�'u^9l)-_^p1@���)�j�F�n�,z��<7Fы�+�NG_i�gu"�d�������%�ݱ�x�����e��yG� ��n�����7%�z(�.� 5hw�!7F������V*�Pn���V�}�~�p��''����8i�r��}�?�����b����e��C͆2�[A-��R�d���P|�Q�f�;���S�aS�^��	�)�>���$���Q������bн2��+�酖����!ޥ=(y[>Z� G�ħ5����-Kn-��[�*���4�R!q�Xb�J7�ٟ-T�H�z /����H�{�]N8�[s�d��1�Z'�EP�X�cf��lR�|��p�l-���Q����? دobm�_���W�-��7E��d�lWύi�We�I�}=�O��N\�+���Y����w,�o�GtE"�����Mȇ�k,�^9��KE��[y;�I�Q^�ߡ�}����?X���9�!����C��� �(�m��@E�\y[l��+��:�L����ii\�{�ڽ#�"��Iq�M�[N���r#�􎙀Ģ�Y=��&	�A��w��r|�0.e�2_��C�u��L\p,A`���)Δ�-�D��~
4:bo��yT�����sr��E��ˏ
���.�~�����������fî=C����G�UKt`��kn��������2y)�s�a
�,�ځ� ��)�f Ϭ�kHx�5���t�ҍ��c{���S-�k��4���|��D�!?���������GmP\7S�Ek���'k��dsq���6��8��O�0E<��-[�k�mf�N����͌�(Cf���H�&yO�n�dtj��C	�"ך]��	9ډ�0�D:���-�f�m��yg����Cb:fd�{lz�����A��56oB�!��)&��q��(���F�L�@l��Ӯ��Knl��><ݱ&g�?SҜ��[x��k�<�ƷM]�c��.7��H�cy�✈�A��sx�=�9u�Nm���)tA���*+ ��C�#��s�Gq��w�~&w��V���:�w�T��Ұ��.za�8\[��hD���{��&��gr�U�{6Yp[�"К|�fM#Gc�}#]3��|���{1!��d���CYB.�%�;=-V�X#�!���#Z~2X���*�)>7�2�N�dm�Sz��?%0 ����i��#.�ӽ(�0�����\Hj�V�Y��#Ը�zF�.�<�d5%�a =�r�I$N,��q�m��4QS���<�پ�u:l���{J�u���1O����BM�jd^o�`{ S^ʜ�5>�{�%�8�rz�i�ِ4�����.��v�Qv�;��*�TՇ�Sj���7	jt��&'���z J�,��B��"	[��Ň'da!77q�z�����)K��#�W�g�<6�[ �󒵩�=�V 4�E3@^�+�X��2q2���b,�pԄ�����q;0��#z���z��M��Ew�C����9����e^e��x�Q�V�����拷QԮ5!]�(�P���K�l�Iw�81^
}�娐�݁	 ��I]�A��i=5��6?��l�f��_\C���ۏ}���[Z��&�����9f���v!�!F.����HÌ�)	���]q�6��g���f���'#l��߰���5��L���K5vrr��=]�#52D�p���ڸ֥�e��p�<�Ǔ	�?6�z�c�z��*�}�rE�>7�@���f�d+~�UW����pu���1��g}ϲ���CA�Er�"� ��
���a%��_c&?=�Q�iY�K��]3O#��0=^.���-�}�J�e���&�S�uy��UnJ�X�eY�;�+� ��3�g���&�fh�
�����S��#%4Q~�x�\W���v��VC}�	��5nwQ7�l�=0ӎ�c��,�*|B8�I��ϖ��>&�qcX���A`}�J@G��Zc$�6�__h�0����.�!��y�*w4��v�UQ
�,j��λ#���U��O��b��f��&�-�y��>���LVju��d=���ǁ�r�MQ�����K��,\�]f�%ޏ�ʹi�/�i�}F��Rܶ	Iy�W�����{=a�i�����{=���)>圝2L"xdu�EB��rz�����Z�U��%4	P�� d8�XN�w�{���I-�1��q���}d�&_�;���-�2ЍB4�!N��E�-f@�r�!Ǘ���U�[�Y���İ�m�<�L��ݐ�ѠgCN���{���bB>GP�x�|9^��%(��%⸎0X�ٴ�b�tg�V��R ��7+86�!WX�z���9�"�c.�"�T`�����}a�Ċ�3[�;��
��)r�Wи�A�V&�.�V�u���8�����8�ӖWa#
�����2�n��R�nr���2�9's&++͖�K!<,���w���9D������O��=	�j���*���ب�#��e��9fA������)d�ðB]�Ua�؊�xэ�w�j��u���;3��$��"<Zi�SMe���E�d�k\_�-E���	�;����m��La��H6��)��12�� `��3�)�[i���mB�9�:�t{� ��x���������6��PNK&�3R=T}��e��X�]%0��*�!-�����8Ӱ�&�x�'��y@E)�A���=-[�P������~��h����Y��/oԭ"���ɀ�S���;��{O=N����$&���ߖ���z�K��]�������� 9oL�R��,���]�RG	A�r���Ǳ�ڴ�Y�j	5 =!��h��^�);����|��/����]�{�t��[;X�svo��b*Qz^P:�����3 �YΜ5���kq]����4�+[ �����p���5Ӿ�Ȩ�v1�EBZ�Cx�r�sF����e��R](CI�d���e�j��2m�`��z�㸵~#��t�Da��J]_E�6�����S�D�sa����Ķ6J5U�dx�����{L|j+	Ϥ�ML*s�yc���x�d�XVSi��KVN���q��
9�c���$�M_��=-%���lV�V"��k}R�ݗJx�p�4 ��b���'y�IY�+�w2S�w|���K��~�$P	ɢ�S*xZ���f�� ;g����{&�>�Ŋ.�CM��I�>�.�uݾy��3��M�X���:%�p��s}�U�t}r>3� �x2 <vˬH�\�\� G5,�]�����r.� ~"��|`�:)UN�B�}�������_��
�Y��wl��"�p�Mf����F�.�#
	aN7�ł�gm��&�v�:�<n�=\�X+�#��*�	4�o�� �`S�M-��pBT9U�D��|Z+��1�e�h�����h��X��!>p_t��<��Jb��]��^?gN�G�U�N��2&�:�\�b�+��G��kvጠy�s#�Pa�P����6��3���1t��?Az��~ f����T�8����^��ڮ��2gXގj�j�xB��5�tZj'6�����|B�d�f� #p?X��oШyTWL�4��e����(��*��j��w�`j���s�;LRP-�*�����]��������y�ܴ���ku5�c��Oh�ǃ���&N��:��:��Ou����5x���Y?X�y"\��$(��`"�p����?P���S����#�?Ra��mQig�lhe�j��T���2����u�R�X�ѕ�j�lA$�"d�\}��\j-90"弳��S����_J�U�G���zlDv��K:�od'�v��[��h�	?uXi㗘p��O��q���@|ҽ�*b�&����Z�>�p'�v� Oz�R;w6NOz�ƪ�Ai5����ۢY#�@��3�n��Ւ�	�0�}y���/}L��O6RT�l� kmY m}L�Y=ʙd�f��Sӷͤ�ەg cc�@%�a�b6�v� �֚�\��lmƽ]�%m �֚Ru0��p�cbԑ_6���NM7�c��{�|uwf��7X�d�{������`���KQW$��A.��6��ج���-��R�p>�Ń�ti��+��BmXv����~�s��fo�"��N@\Ǟ�}Y�;}�YS���)�M��K/�v���7`�>�_�$g���VDh��)��ҳ��d2+�UR���Y)ܚ���ӒoW�Q���ŉ O�������?E�f��aȤ.�� R���tX�J�p�,��(U2�}��N�P�T)a��XZ��e>3l�A�mC����+t�#�������}U_� 0(��`�_��woz�7��`����g��^�-����'��q�2�B���ȃߢI��'��2�$�S�7οu:6���:����R7��W�1t����t��ȡ���(g���u��w��,�Κ`���Eai��]C�JDf:�pȂ�k���Nx�Mة����g��ػ}�b���TMA�*��܊s��|���������&G�5]c�'� y�?b&��Ȁ:��:q�_�g�c�F�q:[x�{�h�O�O�ɑt��/_#�����ע���8�X�b5Xi*<KH��[M�j�C����S�.��S'�g4�9�: �s�4E	�d�{O9Om����cW��wm}��}�3O72cxU� |�Wqa��'?�ߕ��@�7H=�qo���	��]������ԛ|8A~+(���i����ر��Z2�_����n li����SG/����.M(D��X�S���N␀(xw��:}���}T���/o��D��
�Q�G� )|��s�y����;4Q<�o-y�p@`�>�j��Ɵ�fu�8j�x����F�\%�_e�5�����>ARξ��O��B%�۵��DF������c�#�=�:�*.�ⓥ�f�H�X���-S��D�4�(~�"�C��� �B��0�Ĝ�hT�v��U�����C�UZ��I�S]��@�9ë&����IS[�7xr�p����{���
Ι�[���Y5,����k��`)3��t�����g'�e/�rO��Fl���>.C]²~�O�����V/����+����qu�o1������+k\]�mb��,��@5f+S����������=���P�դ{É���+�����)�|:z�����#��!��A���=�7�B�R�#����c�V���Q@\<\�{�d}��s�
uV�}�˺uP~dJl#���/YM�E�;��ev�@���Vd����� ֺ��c8�Jl�m>�TxD��A���)�0�&_P|�Qā��	��}@x�i>V���ϣA5Xɵ���\ԭ�"j[�j��
S�AH�f(����A��qo�%;�?���:��gͿB!������4�xo�^KO�
����{zsn0�w���y�,�$p.!y��Ĺ�
����ц���n�BA��sX����{y�(�YK�F2�E���m\��I�Lx&�r��قOK��m;W���{H0��p嵳3/{"��5�:�"��T��q �qw�� �+�j��ҕ�ҦX��,[�a"�V���x�VqpEE�:��fH��	Q���t>3jN��P�q�7F�$�:�w��X�}{.�Y��M�����`R�]ƙj@��|���I��5ϑ�~\Y��]��Ex�/�g|�� OHg��8GR?��v�^�I�46*1�G��ʛ�ʌ,�5�?T>�9r��-s�����
�Xy��%p\��Jl�;��(6V��n-�;_�.����d|�Z��[ߣ�Z������'K��5vف�dߤ�/!\s�Fv��)0��c�M��8=��c^�I�Χꅯ�a����}�y?"ae�{����f|tu�ԝ/��Q� �@�;<�x����/��#���#��\�\�]�(�{�&����ؕL>/l�A����62����ͷC��������x�fܘ�����qq;tB�O=&�:�c��:�"����0�����1O�d�{��T�Im	jU��BΗ �>_���sq[d�^@���d�:���ڳ(�oڍ�q�9�~�
�o�b�m<@E�c.I�F�q��RX�q�fG��@������n���$E�%B�D[=ػ�-��#o�g�0�`�o��z���,��s~D��b�fo�,����o̓�Fِ>)y��]�ƨl�1F<�����W��Mr�X����(�n��R*C	���6�9g=��b�,���?v��cc= �܉�T�,$��1�hMb���>v�% D��x/��¥I���ڢ٣cu-�_���s��3+=ƴ��T/��a1aށ�7�%�;���
������MQ�ĭYD�c�z�(�*&�>Q�,ꔓ�>���iCe�u\�/�/�EЫT�N�����Ν�V�4�.�(e��2엎'�`/)Z"4�WNg�Mw05���ݸ<6\��ܨn�Ѯ�$�u���B%h��	�����Y	X"&��?��ዙ_�׈�/顾�L����!ԊB��<Ri�� ��C~����۵����V.Z6�!��C�AD_��o��f��6n�q���n��R�CK����_����@���1l�f�:�5�(nmK��y��c︂����@cw�s����������,0�r��pF���u-7E���}f|[ �}�<�� Ad�{_��Kf��U1��A�]���pzϾ���EM��N�{�9��f�7]ؑK#
镉�R�����6&����A�#'�}r,k�-?��ڶĚ.Rc���]�*���iI"RF.O����S=K��bm�e�Y�A"Z��X�J����X�
�S��u.�:G h���p��2j��C�zg�SX�"�e��ĈZ���a��[��q��o� h�ۇ���k)߰����1�F�3��(�qƅW�*�ߌ���Ͷ���8� ���-�`.�ց�e$�и�-._׽#��4X[��� $�V��P�E�����2Tdz�YamB�v�:��M��ׯ!A��UM,�t!�P�aV�ŔO @2�"�0%,_��hM�Z����5�=K����=���B�vķk�F׽B�,M���z.ZV3U��5z=��(��BmM����q��[PzV��Ae:���,�˅�}��u�uT�C��R&X�>	��l{�%������2ϲ��l\)fmY�.�z���.�����W� ��X 
�U��OF@ث��s[�fKvU��+%y� E�19����*�x�3o�U��t,�����`Lj�ҵ�}�l�B������P/�{*�[���d���DlhL��NqP�=k_�ơ�����0�=��� ����r�����0|j�8�2��Պ����76��'ɢ�O��uΨd��	s�1VLs�t��&����'D,���-�V859+I�A��N�`��9.	���`�u�T@_��P�w��<;D���[������S�t��)CP�����t�AEe�uƇ��ļ��X
L��as�^��K�O�J(��i�"��i�7x�����g�7W���/��O�(��RqK��s��r��-�� �Ƙ���KW���$6o�ȕ�܋��y_���+�:��K��E�4ɬ�Ӓ;�4A����&	d� �$-� �$�ʰ4x����4������ɷa8k�J���W>�,c�\�^�y��[)��^�z�[r`De|~��1�Y�5���I�9n�Y��7a�?�f=�]I��Z>f����7����%�֎O�2���%*�t�K�������>դѤ��ޖ���)�6���=5�����}:�-�8�Z蘔�wcɣGP�7�;���Sy��2��ߧE9�M@O,T�Im�%�=z� f7F�SY0@���T9{���&(X���I�熡.f�;1�Wp2Ӿ�K�X�]�������s�v��Q�<8[p���_��7�	[�T��z��f��L��6?�����T���J)M�(D��3ࠛ*�G�F|�8��i�j���7׍�`�j#���K�[U?��8�{]��̶9iu����P�"h�Fkl ����*����TX��*���(��>x�\-9`6m):B���i�rI�&���B:��$.��߄3����
�Yj�����������y���|�K�z2��P��k�br���ȋ��Z�E�<=�^�ت�)6y  k�W�O�D��g������0>�&���0Տ�[�&v��%����:h����OM����/�'@�2k�l���^�IO�g�kС:X�ЮO�14��Oh26�k�H��ڣ�oT(�����*3O��wdx*��dR FG,�yi���Co�/��X�4$�+�����1늕!��eJ��g����cH`���$xm�%�ԃh�[������[Ƀpr����:������6Cڄ�3��^e��Eha����� �Ģק�zѫ:�4���
�?�\kV�{�^��S\���R䨔���O>����ا7�3d�� y���E=��&tf*&L�S�-v�ce�b_��=�]����k�N2��t�~;�����}����	�?��+��3:�_ĸ6 &M��m�]^p;�˙�R�<r|�E�Ɖ�]�Bks��N��@r�u��,��uGJ�Ί�ٗ�����?a�2"�����)�L��T���|ņ�������ݍ��rR��:�������1j�3s�(�1�xҐ������-M0���k�j��K h�`F�pe�J��ۦm�K� ��	hʉ3=�zT -�O$��$�2��iB���.�ր��0��>2"ʡϲx��Yu����D{���[��@#���|O(f��]6�nY��K�Wʍs2/��NE��;+�R6�~�S�˩e��o� ��Z��m
[�R�!r	0��J@BtR����t��j������p&�����I��
,�}Ӡ�'��]�f�2��.ߥ� )�&9��uޖ��U���9|@x��<̂��ȵ��k>�C�	�+~U�(D��s�t�9kQ+i}��)�1�^u�-�6r�[�cbY��ڌAQ��m-���yj����q�����S�%!��_%�X$���r�槷����M���x7j�Ҋ�Kߏ�ʏ���ne��Ya��hn���6�uDc�� ��a�J=�^Rc>ʡ���̍>����y�Շ���M3!���
�����V�_��O/���B��M�N-��)����d����!�!Q�ko����mb ���k#�AF@Z�|䍀�W;u�I�\���~��:eP���eh�/�(���l��eG����PsIfC֦/5o�~���8TO~�T��x�%�.���+Z�f�y����d���	*�H&�*W?
+��J�ӑ=�N�(����j�G�����g=3�]����t'IC�a��m��_����<�A\�m�>��D%e>�n�=�J�*	��p��k�4�k���UA�2`�Lhԇ̘�#_��KX%U���gXp{N���g&�뤋bB�)$���p�����N��9Q�H�X�H�8䪄w Z��,����,A�Z+Hrg�a��H�Ƴ�8M�[d�mq�ΖrZ�� �z�|O�3)?1F����gҢ�Igkc��������Fȋ�5.��b�{����{�V5���t8ƭ��/���o�3mY��)g�-��C��ϓ��i����H�|VA�<6n�BZ��Pe8Yf~���1pt�f��Q�?�"3	|���(b�5�d��T�U�Ӵ�;]Srɽx	2����I��WYbq��(�P2�[$� �9ޙעq�=Ii#B����#.{R�s>	~�Y ��M���`X�8u�Mu��h��;Άkt|Ζ���4���ͤݖ�8�p�&�ni�Q-��_Z�Xp:w�R�
?�� E��
.h�ya����t��y���0�M���]��k��>ʈ�*BS �AV��dE�c@�xC#�&�,O|�&a|by��>�����Xt3���kG�.��]�79<���点p�S�{���������7�Ș�ױ{�K�1hF���g?��λ����5�{=s����r��3Z��J!���Ft�7N�2]]l.���6�1��Qw�J���u0�|s��
�Ykn��7_���I
�r+>ߓ�P�\������0����6���O$|f-��,�v��a	��K��*)f��K%�b?��vI?>�J���cs�g��hB����e�&|3$�G���f�������Pb��t���N����~B���w�X;u+N�/�Y0�B:���7�A'�B�g�@	��]���Pt��z����+`�C����v-ǥH�m
f�t���j"Z�r� �.Fge��)�8�؝�&���?ܾ��3�s�h7�T��Ѹ�ݐZ��ُ���f 2d���.v���W���T@)���#�r�5ZK�
�󈧞�#7�No2=�l�CG��������~%��`����a˔�����A�c�U~��#v��7���k�Լ���bg�6�K�~�ܗU��+yNd���0uq����^S�]���l��ï-; ۡ~����[$������ᆻ��-�3*�*G��uQe�.�JA�=��Y�7)Ġ̪\��Bmh�D��W���L��<����b���P�Y��|���S�Lվ�dU��3�lc;�����O$
��W~�{�i��4�g�靻���E)��X#"a��0P�Ɋ0�[�=;D���-}'$"�г���^�n�Vk �0��T���
��q�{��=x��<��r��鄟�Q�9JA~��ɪ�'p��pi�s�Lt2y\"��#W���9%�F4?eP��9�$� p,2���i=	��tTM{t����([`/�/���y�vc�������;k�{˓0`f1v�nBض�5�TP�	 �� �(2�f��uJ�BxɖuZY���Q+A۪�~�n������jOƲk�S���*�� [2��-�	�e$��ܗ@r��	���]j��]�r���R��.% ��G�p��c��NJХr?�lۤ�-��##E�<s��o*�P�:;@z�:�^Ȋ�E@�Y ���a�\v���*�b�K"J�&���Ɂ�
�s&����sO�`=OS>���y�Ko�f��Zvi�U�R��ݍ�A��p���B���=�[�"�z*�X��=�@�`/�y
F�ˉ��,	|'7j��X%rv�V���)��	`�#������L/R�c�g.El�V����Q/o�Ěto��d)z�K�e14��J*����0��
���KlZ��7	���zW ����]�?��=��d-�(l�|@��c��vb�n�V�/ؙ!q(�+Ư���X�l��f��4��=]���)l~W����]������U���Ǜ�m^8#\h�tZkJ@���FOT�#r��<ҙ�����vN���X0��m�3�}�։�����AD����/��x�m��fa�: �
P�o�;!k/D���1Bʮ={ݫ_F�|E�	�&Dl iX?��┏ܥ�l�՘%�N_�Ҽ	q�Io+]����2�K�@.��)(;�	�e�A��{����C"��H)@�~�J?	�s!8��T��҅e[����c��Ky�D"W�G�� 	���L|����r����匮����@@\����ă��U�f,v�I��ow]��B�rJZ��&������!U�q�)�ɞ]� wJ=%Մ���ǧE�3�j�����r��m��3%�F�V�\�rBGa� d�����3ռ��K�Z"8�KK9�М��c20��~o��1�h3�{R�xś%�u
lё�{�N'�^��T�0A,qO�!��"� �ٴ$�wNMnΚ&8�4�3�;�E&�����C]��7��#M�=�� ��d�~o�[\_�>��T#�3�#�<\m������bK���A�E^R�N?����p&��4 6�qT���!m{)�88����@k�G+�Ϫ����j��� ^_��i���;��2��E��-��:^��v���% � 6H���i�tF~I����-�K���O�O��r���v�,��B�Z�����xի8W߬�8F�߃��z�TS��P,����L�{�t�$����)�%:��}F����B$'��c�u��o�S��^��*�z���e��	wF�$��	�����a'۳�#�!!6'�}A<NI?y���1���'S�I������tg&]N��� ?x����ÉDbl��一��eحd�/IcE5k�y��d���!�N����Sʿz�ѹ
{ƈ{�cH�Z�3]4��� �Ǟ��ݾ
��Yf	bI_������?}-S��v��OE���41Б�/�˞���0��y��Y����03�B�ʮ�!^��INk2�^�HH�~������ID��Ȇ�,���V��ɣܲ>��\b�C*k̚dǞj�bWT�Ng���*rI�/`	,9
�vX�Ž)���~6Pk�b	ΊZ����tE��I��&�^CI;�$�;�G�q`��=F���G�c�I��0��-�_2b��9�
{�s/Nk�o�@��K��6q��LZ���!��\�>�&����6����|;��7�LqQ�#�ݢl��NK]آ��ɡ��zp>�4W� V3�h��9|v9g���8�-�����p0��s�|��x@�7��h"�A� ��@ڕ���yô_z뙒�E��P��A�F~����ʫ8'}L��z�5�h�ƞ<���鶰R�;�v�0A/!U]~���,}#],������r��>b���.hO<��{������
�^d����{!�ao �w5(u� ����)���siGZ�����t�B>Cp�
b�mC�v�n[�1�s���{{U?��=��;��0������)t�Y���	�>��GkZ�ibGY�zE�����գ�����.��-���9}Bc��u%�w���x"
��ao��
[��❼/sl��l:P��� H�;j��~:e�_�IG���}���E%Gl; �I��l�
H$����H���Z��@�KP��`�9s�9�d�4t�M����1�n��u[��QΙH�y���
�AzШk��tK��`�i����L�7��Lչ�xi��EǾ���J���X�1O���4��XJ*���.!���N�'��t6���)�@�?���w5_Q`A_��P���6��N`WcPf�S��c잳���3�`�� ٬�x��x������>�dK7��=R�����7=�l[i�r�ʛ�5�[kZ�mJ�7�0�HPa5����>�,1���U�&�P�$59 �N��2z�K����ՙ:<���²�h�Ռ������D/�	E520�B�iÎ�W����':Z}�ǎ�/�0�i��<����D�G��5p������(�~-Rkp)F�������;���veVj;Ѐ)[���Z 2?�DL?�}�R�����d�-!�EW�e�L��GR&���d�5���j��GdLm�|L���6J6�"��oij��W[��č=��R[~J�[�PQNʕ�������W������9I��:���t��sh�!���(I~ˌ�ұ�ҩE&N�O�h�Ơ���V�r׺;�o��l��Ht�n-;��i���tE*kESә;�f�>W{_2���z�ŕ{���Ga9�:�k�%��?��i�k�4�lP��Ǹ,�$���N�弔��B�9�����6�YDc�reis��Y��fZ�4�2��jDc����P֬����3!ڙ�1��.��P�?9��{���J�K�u��(R�=�ũI˘�K4I	E��&�Wt��/����{�;�H�)&��;��M���CLi�Hd���D��q#�Y��M~ʻ�D��[}/��2����m��J��"�=]{�=�v\��-��������զM1c�$��� ��k#��'r��U�Z��"�SO�q+�+T�&,�K��]d(�P���$�p���[���?{|¨�����lbՀ��*p��g���X��Z��
�OOyR�ÑO|+�b��` OHC����}K�Z�:&�*�I�C�N̝U�eZ�_�l��H(Ԕ�W��s��3�BD��f~:hU�����շ�Q�G-eA�"	$�����D��E-�;�d\�K��>]A��g�E��g֗��P�V�a�f6@�<���8���@�0��H���!t7B�<�Y�mt��wq����p���ҍ-��=;����^�ت��	eH�oH���x����"�ݟ7o��V5/��I�|zך�Fӣ-u�	M���s��x�Sc^�	J8�@�4f������ܯڔ����HἬ�i:Ŭ����LW���M�쁕6O���8bT�)҈��0߶�"k �f��2$9p�k1!�]��6�#2�;WW�m��
��>����`�i[=�����s�dǥ�)�LQ��a$�̜>	�z�il���;1"�?���D�Q��h�P�n*PtQyf_/���900�Ƚ�j������"������V�e���M��p�Ե����HwS�%Sשb�����Ft������/+d�ȑ��\�\��a	
r�Z � 2��f k�"_k���+J+���njkH�f&��ؠ�$�}rB�~C�jb.����0�*B�ܖ���yN�������BWҽI  �yj4u�B���-�5�l���ɏCe�M���X���"���kx)�(�t�E��}�� 5��������f<�Nnq����Z�@#1�|{�͈lb.��/m���L�e^qÌ���͗e�e� .���h�09(��ɂ�7��V�R�9 x�l<��Md����ͱ����T*�G�߻�!� ��G��Sk͇o�gr� �|O�:0C��X��棺x^���qU�Ŧ�P�e_l�5HOvɰvmL�iGz}>�g1��s�+�&��Dn���M1�JӰ�**���ȗ:<�iif�6~�}�y2sl���W��{:ƹ!�~���h.�4\�#`$;8�6�pc�9� Cx&i�T���뉹��"|H�N
�Fj�����t�����vd&Q��7�/@�rV,��4��`�g��j����@� �k���\��b8�Q��<�����l����)������4�Q����Q͎,p0��Я@.iUs�L����u�i��E��2���˒d��
s�6IBܕ~�bK>����y���1�@�׋+���,�u:s��*�e�: 	�������w�Xֱ�������KV���<��U�|jظ���ܿfW�����aV��Oڅm!�Di\��t�""QX������q (��U�f�h��V.ģ|��^�2+e�'8D���:��4M/c�,���*�"�H������a�$�nր�;o�gӬG��*R;���v�x�~~��P���J���b�	�d1�����->eej��ᡞH�8���!��Rh֎ElUe���E����M��V�aayhĵ�� �j�G�o
��o�X�W�lB_L���NW0(�/p8�d�VX~3K����&f{h	����ۻ��}���؅	��x7:d�8��w��O4�[���2>�Vv7��������Q�5o^\?$є��`�P��~@�m�U~���F
���w�_ ��,�u�~Q+C��N{�<u�^SDU��t��n��Eo�Y�go�lx
kK+msevH'��4�_��&"�ty}q$fČK��#模)�-��e
sQ_�G����g��V��Mt(M]��0~�§^���G}��;���p9;���,1���@� �'b��$�J_'ʏ���H(5S�F<���W�U|���;NR��M#�`WN��pP��!!�����'����Ա| �g�F\,������
����Y��,���
�̜��K߄Zf�-C���Öh�,����!����_Q��b�g������[b��/�u�?����K�!�����75���Kq���d����S1�u��<GA���os=�	X4ӇQ���;�57�m��__���r�T�W~����\��hJ�aD�
{]M�vN��������F�q�{t�u�̈́Ą��V�.[4�_C���)�1�o��h�?�l�q�����:�M���*���|�[��8�y1ۼQ'��Q�Tx����X*�]�<�ff�2l����=�+�����D�U0�6h~W��sU��93��/��w�� T�!�ĖK�uORplBla�y�����~�2y��Sԙ�hF�Pe�<u"Tc���LU���j��5�U'g|ߚ^w���^��7�*���W��a��r>�,a(]�a �-�I�D~��T� F�I��4xA�Y��Pc�C������*�HY�<Ր�\�h*��z���,�Ѿ(y��C�����wlg/�W�F�؜��n��f��'����S�-����8]�O:g�V� @����?s�
��؃�&�NE(#��f?W�ꘙ\!zMR� �M_��+º�� �tv�ٕc܌M#-���EN�ƔPD�����&n��p�R3�j�W�ѬjB |X��B��_�.x��p�������i��k�xM1�@[p��>�#�����v���.�S�{��p�gD�d���N]z>An5����+ŧMCS?��#�^UQ�j(�ӝn�pn�$������7�D!�A�d��Y����%�-z����8�J��캥�8� ����kpe/'�9��nw%i��j]{A]`��k���%�6j�yr�94#"��r���-����!�
	 �������g���5��J���F�2.�	hn	e$���[֫=7oa Uz�Vֿ��I���ۦ���ƝGl��%Z�Y�����p�-�c�������eH��˺v�}d	�O�m�.���㑑&�v
:d)����ƪH)�l�����(1s"��� c��G.�������l+ɗ8�Lfz�b�Kga�T	�������*Ϗ/VoEB�L�)�GU�!:�f�;lt���T��҆Mt��n+��ɑMe��;/l��"Y�i:��ã�fp'�@N͠RIg�
�c�H��eͿ}�(���0�y�h��O4�i^ݢ��N�Β�����eo�Q�r�0����@vv�h����l�&KU2�W��������Z��D6�>^[���p�d�͗GCh�!on�����d���R�:^�uqW#b+���U���!�<އ�O!V�@L԰O&���&��=3���s\:��s�V� @��iE�u��N�a�l��ab������ ��;�b��^��W�
(�@��g�q�w�j* � >��!��'�B��� }��J��m�]�~�l��n����D���N֕��g�PU)�l� JK��� 6��j�UC���T8��-���$��!�'z�V�;!�q&ס��`�z,���̻r�mWF��t����sS�/#��Lm$�?���=��b��k�w�\��u������KDשV0��ZZ\��v,w;����~C���0ϒ�b���V��]}ĬJ;����Q|�G΁78;҉���$Lj��.��؏�������F>*f�	wP���e�/��U��jTam�筢��"���֡o��2��\(��6o�u��o'�R�zflJJ� ��d�9lLO|3��E�wpU��}jJ#��j�F�@ ����nW���E�%*��R���h���=�4{j�r)���d���S�������{Ź�2���#��%tb����9q���3In��ER�9M�!�<%EK�$)U�M��8k?ؚL�7w�m*d��p7��I�ޗ|<yV��]��Q�q��ى&6��տ_PZ6��&�H9xh��b�֫K�'2>q^H�2���-U�����Ms����p�/���or	��V}3{��	����{��d�/��s����rj�!�{ũ��n�����ܞ��kc��{�.Mnǹ'��yp�����L����H�����Q�Ṑ���{�ky�'5Ʌ��U����za��r[�3uYK� �����v��C\#2WhV�J��v!q�^H1��K��m�;ͱ9�0�/tɂ��ݫO�w�w|B���pف�e�>˔�d��Nw){v&V�|Y��,r�/��G��3#˂�������Q]d O. ����i�R�������&�m�0x5R�U�Mc1��,No�ƫeⵟ�	��5��\�|J6(���K���AeV�����c}������j�q^Ή��77.�r�j�3p�8��
	�戇�{��<H���O)6�C�����m�`j,a�q�8F/���=����Y#-2#�-��D�4/�H|r��ƪk�>-�S\.�R+4��?~�K@�+n���"R��Y[���$�ݑ���|�'",v�Ė+D�M����+��c�:�G�N[�4�$�k	��츆���Aq4[ʤ-
�NK�{�ՑП���?7�����yd-t���o��'�}W?Ҙʂ�7�6������+[RN�$�8:�K��������E�l1�bk!�|���M�j~�,����\������z[t� |���{�2a�b�����-����X���&��Vwo����,���'�n���"��#�7�<t�^���)4)��{A���?{lX[3G��O ��3-�����f[H����x�:E�Z������@��F1@�o�c�����A��O}y�����یOc���+5dp��A�_|N�O1�1�(����-���{�r�;f�H��P{���N�|3CM )�#:\���꼺Ʌ
�O|�;E������@�9iWA�)���C.7Q�6�*OhF�!9տ�>�	���u�y�x2Y�|ul�#!6�~x$W͌c�%S�FZML[Za�\}��$c>�9�՟�zeg �7�gL/��&�	��W,uC�)���_Tv>�		��$T�B=�q� �	-W���c��>�S�n����6�]�r(]��ۃX�ql3�F]6���Gڢ����GPP?K��)��U����B*�W�������2���Y]9���=Tw�v��[xp���[�n�+a���2k��'�'0"$���mWFpWhJݨ����~�1����bH�L�o%8ev���j �u��|��zVE���q���IfV��G	��t!x�o9�w#�ʖ�d�'�� +�Y��T���lIM�g��b�MC��LC�PK³�`W
���n���@��5pY�CL&�!�fB��:���7�;uJ$s��n�n�>����մ&�����.�Y5��B�\��uū���a��e��� _�w=��*V<;F�TҚ[�i0+�ޖ�(�d�#�قi� `NP��8	��k�h�)c"�XS��i��+u����5��1R�#]Nx�)
�������S�w������e|���x�:��Kʧ�e�c�t�m-5?>{��mY�6�z�y�v�^ZT�N��������e�.����{���p{��(r=/��h�/�"���݃rA)O8�j]z����fH�e��i�9x�������-���x��ZMrvNə>:?쒝��H��u�����x�o��K5�`"����ZL�n��sb+KoΜ*b�w;���^?�.|����n����F[0�^���^&���Qe�"�x�Y}�Jr/.V���/�ګW^�"!�D)6d7�@ ��1�Y��)25��O?� �o���N��b"�HY硋��=�����vb��(&�K�\���p�P�hЎX7�Z��4V/]������$^ba�%�� Zg� `��l�����3)%YC��w� �9�߷0�� ����
I�:�d�	Ȟ���z��!����f�J
a���ܸ�kΨ<$է�'ɥ֚=�^絗���GN�td:��;���|��+)7P�$�ڙJ�(kX��� ��[{?���Щ����s��/9���t*V!��i6�Y�݊�A8O=���ǉ���;
���nR���|�e��ww��w�V��S+?H�J�����I�fY��k%f�a��������.�^} �B�p�R���ˢ�m�W��ݮ?�vzv�B�����&�bT����u��=�;�e�2?�Ԗi �O�xyX�pc�c�q�<X���x`7�ҝ��n��ZI�^�>$�޼��cs���O=��
j`�]8JdL�s��4����G�?�s��H	��>_�{�597H�n�1���\�w�D�[+�R>v���V��o �ʬK�#�ˢ�yōj0n�=�II����ҏ����{�f�g���j`G���b�.#QR�iia��,QDG�Vx�UP ��l%��ZZ��-W�@�S�$������9�]�����+R|�܃�o~k��u.{����dB�9Œ�4��s`E�Lhjp�7cmޝ�1:���7�d�D!�Q@��
�-��L5�/�^Šb�������[���8���C���[r��� VP�u%&���C�(Ƈ�h� �#7���5>��#�@��e<�g�,'��W��GqNF1\�	k��;*�bk��Qa�퍰XL�YW�s]�^��$_3
�����W������r�Ŵ���$��
��u_��P5�Sa���E��m۫��A}`�r���'��� �?���m��d~K���D��(5{wC"Hv��� ���2�Q�<v�x������^�薼���c&t#��Gk&޽$�j��k��k3�yc\E1R�R��bbW����r�K{5�~�V�qeG��h*�:���rçi,"�?��־��k;ڵ�{h/d�T��\¨п��*��),P�g�A���w;z���h��ˇ����$[�?����F�0�	�ak#�9�VZą�{*��\��ES�=P���̚u��I� Z��R��/�;���qJH{bÄS2����������\qa0t����h�����|r^r�)�+�~P��&͒��W���{�:�p��a
�>�W�)��H��31t�ޖ-���1ۭo�A�͗�x�<K�Ox�㯁rC��4�cT�+N�0 _]�&�y�wrea c��V�D��ڐA�-i�����*���ۢ�p���
��_*�%����C��z��� FԾo���R���h�Ӝ���V%>�o�Q�<5r�DR�� J��ûlA��=�[�C��Ò�����n�W��N.�=�Iw��>ĖPM"�%��]�\���:���F�4.ٽ����ʞ���8�=���� 
*�_��
]I*͒���6�v�vV2nH�\�%�2����j�>��� ��&�ı�8>NH���|��O���	�<���IH�I����S���N�N�����_qބ�v���=�f��ޥ�(mMz���
�
.W�\4T��pa�RaT! A��'r\dA��P�딣h�,9�B�C���9��K�wΫ��Գ!��:�B�{$
.�8�~�����V��,�3��j�p{rp�Q/��G1�+�G��$���E_`�%�'��֗�G���3���v$�iZ�7�k�Q}��K��6��w�ɧjG
�݉F��`��_�I����p���.]b)�����=o*ur��U�Xl+�����L�v��ϑ�M#�r�smI��hފ��<�Hm.�T���;��C�*i�rJo��8V7Ǫ��\��*�)	���PO����j��'��{�L�$K������V^pA�'���c!�m$�)��(�!�W�����E���!��p��t�G�����������;�ɢ?�U�G*K�v�=c��lP3'd�H������cC;)�zO�yA��^�.�M�t\���+�=�|H�w�G��5bB�@z�ٯ�	Ǆ��D(L�v��KH����b��{�z��C�)�k�G2��t]Uz�g�Ϙ�v{�ũ�w�hjr����*��/��iz@C��d�c�+CN�b�P�J�qbǥ��y��[@(\�d��j�P���_����*س��[�w<�ݤu���Q�n�&��?�m*}f�����H�jly���.�i�OK�t���#��!'RWE�����_�Z
��<��M���Q蠭5%��B�z�Q��ɰ��7΍lͅ��&���an5ǆ��Nm����ZkGT�(������?{'�uF^���x!�L!#9
�k��0�zBo��(%��X[_��:J�M���T����<|-��6���<�g���=��C\w�yFISO�*̽����s����ْ��;��/�S�d�%���g���1��B
1N|�sK�H#�A�rNTN酝��Ƈ\
QP6�l��n�gC�v`dP��b~L�D8&�뮰��)�k��w���3G"��1�Em���ϑCc�~��qC���L��w�q���Nӈ��u1��|�-�KY�N�j�4d��"�	��$�P �4�>.�!���BIznM|�����5׉��	�<7�vƨæY�Y/�P̥���8&�m�(U��l��{�ٕ�?�+�Q�(�}��������$m�ӈ�~'���YS��P�Q��[7�<G����_ff���9-6��l�����x���xJ2z������f�5_mC��s=��j)Jr�m��8F��|��ԅ�ܚO}B��y m��h����%Ӽ�Cv�5?ikO���M��5ƈ��e�Ej������ޢt[��2�gN��͑��\"�P��.�PDܳ�?i��4�e1~���ub�`�4�:����'�G�u�	u�
Y��&�g,"�#P�Ķ�^���Z��=����4��m���g"��q~���
G������f8$��������P={	^C4/V��d�-����j�&�͂~�/�/wsa���Y(mԵ4z�b�����6��I�cI��f�̨��^=�����XD�
O�}��Y5F�s�D��ۺ��	Y�N+�ߖ8HM�(��JP\���r�gGd�h6I�����	�& ����X�Ǜa�G 
���Ug���DK��2�}�]���g�*k�3�e��n�;���#�'�ċ��F��y;�Ǆtڍ-NG��"rr��g��lk=�r^`Qfxw� �����R¹����z���W��T��m�ɂ��#��¥9׼�B3�|�sUPW&�����Ҧ4ă�Y�
�ć!����4zU"��ȕ���Ֆ�K�Q�F�ש]2�4w�^��aql�w�(�I|X���7���1� �v� �5	�Qfˌ��F6P	�wM�?��ssw����Ȍ7.�5N��\]�5r_�2R
i4 ��n�ʏ��b$��D���)%\�e#���:Y9*���a�O��,\�R��>d
*�G�=�cD���I�o�ޮҴ���Oe�� ��`��i�p�~������3����4Fg~R~�x�̡Џ��{`�ˌջ��F
��$ ��	��-�ua����SZ]n�<1Æ+�	�m�Z�P�\��"�*mNj Cw�=���I�.�N0�N�:�����%�8笶�hDyfEP5�u17yD�8Ϋ�p(?&R	1�r`<�آ��-B�Fd;ãό�9�yy�0�02�Y�|�݃�����g�բ8��� &	h����@-��L䜟�>LR,������1�E%襕����d	?y	EGB+W���D����SN=���ut[���q��C�p2�T��Hf���C�Dp/�'8(䊫h�<���3�C��u��"1t�$N���w�����t/͖����i�}[^
<�KE���8:=��� Q����t�b(̥
�//6c�u���?a�`�	���j6W�C��le��J*LLdݕ��I"5^m5뫁�n��Nh�P�#���k���-?�&�x�ZXQ 8�z��B�F>�-���n��(����l��9�ʃ����ğEP>��#K���.���{��֗���A��/�F�@�(��u��l^w)l�|����0�;�´�LSӪ%KW���nY�f� �3�z�m�~>��.0Oft�=��p�!�ղ�Ag1F�e{>��1�&{����@����$�6Z���.!��[Yr�c�\Ч�ʲ���q�s�t��t@��f0P�.L>YV�
�cx�WU%�FHȡ^���3�e.�MO_Wdi�uR�Ȕ�f' �l�䋜s�&C��F����(�^�Fc
q��E`����3���ОD�r�^�.L�|��t9�|6������+�����d}�z���X�^������;}���0J;��TOG�p����!e�a��l.��
�t�Oxl(~�G�����S���G�^O���mk�_#��i�/�L�M�IӦ#���������&>9�|O�Rr��v��[�޺�����Z&	�,��|�:�Ɛ5*�@)�W�x�8�=U0c�*��q������h2�uߝvS�0��+n1��?%�D=t>�7�)�޾�qH�%���)ק?�cق�Pq�;ڠ_k�0(�9�^�/n���)6W�sri��G�CKvĪJ?n7`��QQ�Q犗��8��̎%�Ļ��A�h�q�\-�*������H�d���?Y�$�g��n��Z�Ooɍ�65,r|?�<��hh����+���#t�� �m�Y��x ���z�p�Y?e=���)�,Ov�J��[�$�Jߟ���{�y� IKy "��L�f���vEBbP���Y�ܻcR\%C��H$)EL k�?���|�� �L���������4�b�>��Һ��o��֓=���CWO@B}��j�.��h�Z���ˎ�R����me3��n�0�t^��.���1�,�g�d�ưџ��｟��}#/�]�xQsW4�A�z܆WM��,/�&��	V!��&c_�%��j���iq��_p0I�������r�jl*z�
F�RƳ$�]@�3G�x�:1̂�������Xۜ?U���'�X.��78��#�U���q�Oo���+oz�V�*а�C���E>�ǔF�!+DPxP �*�#����Q]rD/w|8H�^�v��؉��T�	s�¸X8c3���Tl�;�u��a�0[Q���6��\� u��FA:���n@#wH3qɳ�h¼xC�]/;��9nG��`���<�nh���.��<ME&��l����z�s���kg�v�}x�^=v�ޣ��̾?�$rx�v����ۯ&���=��X��&U�e`��2�oUF�p���m���C΃���6��1�)��#v�b��cO��/���@5��;�HUIn���9ԒIk���r��71'� �g������mUD�}Jz5(+3 !�!�d�)��<\17�:К(Q�5%ӫ�f��E'}�a-t?��\϶FC2�fm�$��~Ը������r�-�y�b�g�܆x�E
&fC���M迈�0�J�y����,��%&o����:�ֳs���K�6�M �BuI��L��ܷ�6wM�3�\��Gy8z���V�e�y�TW��W��vwj��6e�_s/�;)rO{R��)�S��[�U���QЎݫ�����J*�Wd-�٬�6��v���^��d[	N�(���MR��h��Tְ�02���j�s|{�:��dI���T+ ]�2<i]r���sM�Pw���с�Y�����d��e����i��G�E�B.c2�$/��(r8!rI�FP|ٟ��C�`���w +�6iR���6��8>����H�	��.�񌖹��ܔ����!Z��v*���-7r?n�kT��C�������g���P�[tީ��¶*+2{Ƀ���Y�
�U��
���m�2�U[�f� �b���E����,�h��G�� ̀��������Ɇ�:)�[5n�	--��2�4s�(O�Q�/{����Yo� p�}�3����V��,`���= ��]�_��U8e�*7�@`;���_Q##�$3��4�چ�*yߋQ��9}���/�/����&����fK�����K7��xs��p�#��*������'U"~����@@�d�8��{�ɯb�X�<�R��I���96K�B{K��Ǝ�AD���Y�
���4�>(�}T�ձF��D �)e]�k�(���5��5s�����|W����r�B�������v�A���2�ٕ��3L�z��0J�Y��i�E�``巇3�ڷd�}.n�����tY���Rxi���71V�ys�Ϥ	�q��F��y�>�����(��A�*O[�$:�l �IH�� T������h�Q����"ހ!�ޕ'��m$}8\Ș�w�|����ؙ����D�7m�Aoz10�؝"p���Upf�D���b�Ð�KVʁ��Q%0(��R�_aoT���*h��H��l��DS�(���-b7>�W��/5���&z�o��>��*"iF�J�|
��]'��y2i��*Ȣ��|���0�i����}#��qR�^�������n4�OR_9�ǩ/tj�
����Û,]�����FVw�����V� ���)!a�\��9�H샒��4�n�<r_��<g�VX儊�_�}��R�-b�6o
����rbN,v������R�K���}Tk�Rz�gU���>�7��I|;�6�7��at�!Jt6lwX���i�ցi��+�ʟ���2���T��k���)n,���,�����<u�,��R)㧵�mR��+R�V��}����ۯ��u�( ����/X�.o�Aw:s٣�d[���2T��Q�X���P�9��Q�SSs?���rK7]?Bq]�9��'�NϢE�9d۵�)~3�D�bs	��Q����c\H�(����,�˃^�,��U���!!@;3���l�Ez|���X�T�?n3:�s����A�p�.��fY�LQ��nv�s�Ia6m�����7�EI�L�|�k-���&yKf�{�c���P��͈=6%u�����L��FP����ҳذ�z*��4�!0g���Q:`���!�/�+&��E燫=�'�]b׹��mQ����^��fs����UK���4�3����\�����T-&u�p��� 6�s�&ǒ�*9{���K�ǯ1���C}=�=��x�Θ�%-(�{�}aϼ����U�Us�6<����t�сV!q!:�*�g������FO��̔�h������w�� (��a/)�sFC
��ᅤ�"�)�J��[�޵>��H�2?��q�T�jn����ȸE���&�0I��[EP�kG��	���W��R!&j}��rǏX�*����(�bjHA�2�I��G�}�� �7Xݿ2�0�y�V��Z��rRH�y-��!7���yyF^��"�k�n��Mc�v����=��5�y�
�H���aȹr���i(��y*�x;K Bt�A#���E���Ĩ(��˃]����Ι7�TaKQ�7�E_+G�˙-r�VX��P�4�i3���-�2��϶?�r�H�z�/�rE	����(�����Еm�%��3#��Ԯ��z�fe�.�W�5�D��M]d���Y��<��)r�r�]4�:棂O��O�+����s��1t1uA�w�9F-&as�� 6�I?~��.:l^OlI�Q	�2��]����DUu]S���r�آ�'+�;E��#���O�=?���rӮ�����?A;���D�	�~���O�y��U ���ۙd\X�Ig��EC��rQo�0�
k���� ��zg��E^��G��~#N>��z��O����}/�N����YXh��N:ʙ�����	m�*�V���^H%8�a�e��=���Ж��ƅ7��@���Dٜ��W���Ξ7(x�t�w��1��Čq��Yv�������WD��TЍU��#�� ACdԻ��7���::�W�����C����v�h���K��$(Sr���^[�p�����U#�|i�u��B����F\§���fȉ�,�ۀ���W��Mief=v�U->G��~�Q�4@���[����j�T�/V��QL�U�DL���i\=��A�s�{��&�§��>���*v{�@�U���\���.�s��k3��[����A+���S�强�,/^[�s|�R>FO�����R��XEt�x\���b��ﳗ��J�1�\�^�����_v�^�LJx-@���N�����
�!���O��\@p���E�3�[��p�e3��I
��}iP%��J.�7���6�٤��$�J.�eF{$�w�=)�LI������L%\{���r 3�Vr��U֬�ʰ@9�����x3���lYD�?�ʑ�f ��;�h��� K�	|�����RP�������6��#]��;}5��o�I���Y0�����zZz�~��3y 0͇� ����n�#�}�,oaˣ��<��C@���[���E+�`�<Ve�9��>�ؚ���D7s�Z [�����Peֽq�'��a� M�X)Y�];5z.�?d�f��6�j���
r�>��䒉�֧ʵ����
LZ��_��B�m_&e�wm�q+����o%�Qat��w�tބ<��{�9n�y���"j&�����|Z�\���W@7�cF�x����k�[p����m�a�uͭ6c� +�'K��K �8V˔���P�Z0N�]�7��*"M��j���:xOv6�K~�s����+�	��L���R��$�m�S��8�7�"%��Ǧю��$��,�\m=l���?��ڛE�#N5vPJB���,�^$��liڵ��:�*���&/�c�5[�5�`u�A���y�m��,C������J����6e�B~�>xyW�	69��e�B�rK��{ۨ]ĥ�aj�-�td��!����������ֻ�i*R��L{%q��U6]�^�wF_���"+F������O��Vr���=K�
����	�w�S�	�^��ԙ��>w�7-�vP'�6-c�:_�7NiaeDA�D���U����S�'��5�������kG�[1 �53gJ!J"@g�P֪6�۩#���m��nӪ��%zS�-�P�!�瓂�|�#�zi�q9�/�-��"��?u2��[��a�S,b���rpR��쌍q���S�CG�z��dU<���\�X��&'1fm�-@e��N��I:�E����U��#S�4p ����ZoXÇ��yh������L8��N[GyH1����.0؁�C��=⎉(�.'Wh��B�@LO��=�F�X<'ĕ���D� �!���j���>1�������?dw�T�Oz�=<��{f�&\���s�((��p1k����H�޳�6��2�F�ދ$��[K�Bk�f��W�y�s�ӥF��F���P՗�����ֲ{近�(�t�Di+=�RAؑ�f��e�܂g8]����{�A�K�lfҥ#���Tn�X�̆5=�:#��\hso���yg��<^Ł�ޙԅ�a���.�5��gi>UP�-��fe^pM����V�H��j|�ڑ�>X/��Ae�s� ��Ը��?�p�I�kɒ�mǒ�dp��<����A��&��F�2=�h�k�7
 KD8]��kX
�/K6�!^؎��C��G��2"�c��= ɺ�>�oӦ�#LE���!*.~S1����C����bI�D�H�ia�2�2X����*D��]��y��x�^_� �i�a^�����C?Tx���/EQ%υ,NY�OST�u��z�1_����W��x(N����uUE���mo�����]��t�A4�?rfӓ>��f0�#�3X�Yf^]�ðDޝM�e�6L���|%��ơC@��U�w�qS���BXà;�xGӳ��uL�V�T�T;Wʗ���(7{���J�g�P/�{:��"Џ)_�X9rxeob
o�ځ�C�q�mĮ��@�.QY�#�'���8��k���['���Z*�k��Q*˷���'<�/}�qc��$�������'��JVj�I�c�+c�]���Srr�Y.�MS �*�: Q�if�F��H'L��U�u�ᎈd`/��w�:_�s�����Y�UZ�=��aF
�'�I�f��20)\���6������6�Qq4���D����gw�9C�ΰU�3�wlp@��	A��C
�v�)�ي�'9�4�?!U�5"�~D�eG:J̡6u5���,^��B	�����J�4"E�pR+A�`%�u�HGt��'��Mۧ+�)u�eu��־`�5�M3�oM50�C�x"	1�n�y�~�8�ho�=�bﭞ�H��-��>�w�"S�ikm�(���c/"������m�K��XKd�{N�P{��#�'��{�~c����� j&��e$�_�O�l�IȔ������בڙ�v<�<5[�a�=3��=ⷜ�eR� *:��No��Y�pE�)3�9��������Kc^q�+E�l�mCgX�!���R$����YWy��kͻ:?'���i����sby�:&10��7��Ie"�5�A*b�L���@��g�yvQ�{QҐQ�7?������(�쏬���:����:���÷���.m�i֥(��薇�'Y^��B6����Hr�cF8�Z$D�4n��E$�e�?����a�2�1����@YHh�lVX�����Ư������[�h�:���vQǂ �}D�e\?�4[��_�1�-@�I˰��/ ���z�JT%!��x��oC�by��}�ep*ng��� B�������fē%�O�Lo�]@���a�_<fY.KJ jo~IY��	e+��������:�b�*�{�$Ŗ��$FM��Yl�"��:u�E�Ǯ������N�{������Y�Q�vAp(�(H��N�P@��1L�E�ሣ���l^x�/���I:�	Q��ȑ�j�=$~�Fi,�;_���HQ3����= ���&�YV�΀��Nf�wd� ���M-Bu�R���

�Rq,��F��0e��� �[D��0,8��O�'�_��Imu���@�0Z+w��h��	�~2�$�:m����Hp��1��c���߃�䭟2mcԽC��S}6Jd��������O0� �B�]�����Qm�B����L)4O�d�<�c�6V�2ȡ�4��LM %��Uó]��6E&��be��Q~��'��P5�rJ.'5t�<s2�*��j�,������Ɉ:���tz���OF��݊�,wyY�v	����������aC߼��ԥR�X�W�U����3�z��ߌ�7��3�x����XsJN+6���2V����
��2�9��q�ǇB�����E�8z����Gͷg�S��q��/R��N~(����|��:�p5�=M�0r�i1qFU|\�-ƽeh׍�wn6d���&N�˾��Q}ތ��G���D�V��0���4�\Q�u�$�0$GwM��Y.�Z,�oT���X$yڤ�"�E����M���(�8�-�v����m���_NO��Yp�C3GZ�P�?��\��_&����=��P'�J�<%6�o���]��|���o¿Ʀ;���R�.j�(�Ik���ʹ�v�w�#�S4��h�����X
9K<LIn;�'�����H[E�	�i+�]M[|Q�+NSjj�#e��Sh8}�ɋ�`��E!��`�O�'?0�  g|���d!h��<7�A���Џ���߅A7[��-M�3��G�JAb���:�p��ib�P,f��a�shiZ}R�)�MR�.��ͥXP��=Y�#i
G	�F_�&pϕ@�қ��2�ԓ�+��H���,�v���ٖj��d �Eb��"V��@�o�?9��%�RAE��z{rNW|�A�����2��iz�m�*�p�7��~��=�J/x�_F�\VO���U�mq��iCg��Ԝ���/�|�c���(�n�Fo�֙��][{$*�p�d�����{�4�,�n�1��&b����t	i:�e�k���$� K�
�_�W*5���� �ǷF _�Per�m5��ᾲ�^\uu�e��C��6v��R� 9�J��1����L̅����۳�*�.K�779L�~tJM������H���G�a+{ B�T��!����b�����E�}!���tRr�!�����b���rj����X���u�,6�{R�6~�ɾ��Y*��q6R�����L�һ�c.�'�g����MUzq��m=��7p��ƴ4�^�dB�j}�a3ƈ��=��8X�,А�7nN>i�����'��W�:��z������M{�'Ӛ�!�ԡ\m��UGŒۃ�B�yk(`XS�(8J�L���n�#�+�8U��5h5?�-�6�	�)����WZs�hD�1Z���J��.�O)�:e�گ��1���}�D��Ņ5#����>�)f�C%?��N�����iŕ�$2fu<��i>C�X�'���7�۶��Y��6*��*��<mJE���5f��1��d�k���j�8/����fC3EN��pN��Mz��JL��
dj��Iw��B͌5]Q+c���,ޓ�1�ih��� �7K���-��=�Y�d .�$�h�������c\W��rf`~"Vֈ�=��j9Z��Mv{.�0?�W ��ǯ�f��(�qm���PDA=�@�Fx�Zˌ��{�QUc^k�{��"��GMJs�X�♻`��Y�z�H|�����U��~�a������w�3Lx�$s]-ID��S�51�H�Z���D],����Gɏ���@���[j���7!З�spl��~
�nSb�{7co��ࢅ�KT���atX�v ��s�]��(tT�����lj���fd0��.�sqx�T�S��45.R*��2(|��G@�bpXE
��3b#�����r�^F����*�S���H��!�{��b� -�K��Hj�@��,��2[Xu����5>v�7�0B�{R�SY�)��;�Q���	q5�M�D�Y�p�WA�:eE��&��ă� "M�pM��S˷N<G�G����%�uD�(��(LhЌ���ivKe���dQr��; ����E��(Q|&F��\Dtx���r� u;�xcB=����#��ҩ����1an�U��n~���6��7"&��Qٳ�(h��|Z�{��B��%�!�gmGCsHO�����)M�>q��Y�U��F)m>����s�p~��ޕ�ல����<B�L!=Ē�~���:x}��dc�ߟ`2�o�� �
����1�ktO|�������+�/B"�k�j��ٹ�	׵�s[��'z�F�"�0�uG�X��3��^��m\�A���v��I�]�<D�e��n����(�)0'��\Ej8�V
Y�7�x�ֈx�>�R�-�Oyʿ����$d���wJf�[��Oz�����b7�@�z�Lk����{��򄺨�W��P0{}�P�>�r"M1���a�6�r,��1��']D<e�V�:��K����W�V1��e8�K���-��	u|��ŵ�.�I.��7>���ܫ��(J*bJ���~f��a�8����ؼYk%j,�p/}"T�*pv��2ɢ�o}�B)�x��֯I	��VJ�[��)���;�{9A�
�@�VJ�nٛ-���u���?�S��T%S
0�-b �M�E��lA���S����!F������־��������K�X��Q}p�/й��
譈̋-->Bf�E��Ri �c�J�1��]a�D^�X`������ևd�E	az����D��ϑ7螧��*�tfȺ�%�JJ=A'������
�Ԕ��<��H�M7��q�����,D?3H�N�([|�:X���x�0C�n<�F����ofi	��L���Ў��<wD:*�@'��R}��y�~��*�G�X,��������AD�Q��Y.5�bF�\�~=O��:W{�_|��y�a���6��}����܃]������R�hӺ�贖z��gSs�@~L����������1����^�B=�l��q�c�!d�f��A	� \�h��(-���x&�Z�%�C�olܢQڤzT[�]}�#���L����Ֆ�:#��6V����r	2��B��å3ۿ���K�C��;�����W�<�WJ��5"��e�~}�ݵb=A��S����#I�/?���gz����n?<*���5GC[՟Cr��'~�_�`sL��1p��Q����_���4T� ��'}ݔ��4te�Pʺ��!�֌���X��%A��'z�x�"8~0�ko�|��<�LHak�z�	��D�@��
ʤQ7rs�=���I�'c|h����k����Ͳ_�D?oUb�����ĉ1k��$�,����ޤC�L�[�9a1? �=����4A��y���Q��v��U�3&��M��޽ক����ڀڨ�D�ʇij��GC���a,�>�����yEH�ta��D�
��7\����0��o̠�����J@Z$l����q����KX��`n� ��h�XZk��@%�N����K-��.�e�V;��p���~�6�%��R��!x�8�d9߉]��C4�&-^����\�3	P	��8�*�I�IK���z{껋��qc��_B�̩�8�A���e��&������K��٘?�@�n�dN�\�����]V�	g�t!
Á-����!\�Mm0>bg�ݾ���Nu����H<�6��?����,ۚ�95�n�Z]�m� @ڱJ{�_?���4raVO�W�=Yh-��O�1���]n��¾:܊���}����a�3@WKև�H��is�3��BI	��v�qh�����;ʡ�&{q�����M���x�U�Lfr��M�5�Y�M{��Ψ)�y���"j�?yc��8�|5sD�k�y�nKA̓и��S֦}��[i�\���u(*����tU��B�iȽY�$Z����E��P)>�"Љ{�d0�$�<�u<a��=�!�yD��_�q��n��V��n��ܱlzq�U炊o��]녹rkx��5p�_�f!�3b���� ����iv�N<K���^���@�Z K�x.�3Z�i9������r�	x�-zT
*��/n���s�KӍW��D�$m�^Ɗ$-(�S�֚me��ۧ��MgжMHu���((�A��J��k��q��w_ַؐ�8�:[d��EVЩ꣊��	>R&����5~�g̊�c�����)�\Q6zD�Z{S ?��n�;'6�ΠƱ�kr���z�	P�:�l����#]�L؂����~�T+	�2�a�0DVءaځ�Ci�z�Ն	�k\������B7��lf@����U1T#v���s�u�~���cӟ�<�b�!�5`� �аȪ	���,�P*+শ�	IԒ����u����.��O�&��/��;�7��qb9��m0#��:�黃�x/<��RJ���FD����sیvmp&s@É�H;���6�Xmm;���X!B��~t�%�DL\T���=�{h�!4E�J��f���k��@��_^��a��q[Q#���ٮ
{+�cmb7D�}�G7c
?��ls�)Z�p��(G�~���z�s� �ri��bRH4��}�Ȭ�3��ɛ�ݔHRA��*XP����^�ڬ˶~Vr���7[�|h"���#E�J�'�KY<|کP�ሂ�:3�j�lMa�'�Y�����Z��QG��Q�ʻF���H�w@�G�Q������S������,�9lrJLW!����l@�!�xH��+�M�;H@��3��p�"< ��>�n���T���g���?��=���!;�_L�?9�4�~���^G��j�����v���L��Q?�<0?��aȚ�{��iA���<�_916�Q����*i��D���8�A��yz�v[�5����!���a�OQe��8�0��u�]�[:H�-v��|���0�u�e8���ᦼL��gkQ4U�,#EO{K�����ȂKhs�(W��4FP^�MN��
W�^�}��svad�toʉ/DP��y鏼j��[�}�t�dS�ʖ�[<V}D>6)*�UYd%�����Rɼ]�� �B,����e��S6"�H=^D�y�"X�B	+�}E/ړn��-ɖ��AW*	�}��w(���#IR`]����h���,\��۵[�{��E[��P��	��t���"h��Rcog��������a�V�`O롵�z��=�,��Dcs�ˋ�[˫�}6��=���H\���%~�������i6ϴ'C�2�>U�*���{5 ������r�gM7��4;f�s*��|Fm�qCq���z5Z�(,�fa���3�]d����T@ܽQ�?��B�T�)}?�Ru����s��#���qj[H�9r)G����C�u#�/��8;��jiW6�_�<J5_�U�;x��H�̄Q'��$=�E#�.ű�R7�G��)e�
���z�dg@�Z)Ǿ
9n0�/�n�yS�§<A� `�_���
vq��z6�;Ns5��pY�#�%�����U�@ADK�j;�ǆn6����I����*�'�DQ�/��T�6�s�dNSƼT~�:�G����؀\nih%�!֩1T��&A���v:�~�ݓؒ9�R0�2������
?[o#��ʂ���i���m�>���`$�Da�jי޺ҩq��H����f�<��?6�*}��'"��*1!o�K4	7��ݎ��ڪv��6ՐzZ���m���X5e����m.�m�f�)s��YBJ�a�W
n�{j�Z���RZ9'�jy	9��i���#�h���
�c򒭓���؂(�Q,�����yA�B���>U���A]>49nRp+��CN�uMX��w��#)� �> *_E�`��I��y��SP�,9�w�P ���?�ZA�d��r�.���x�
[�ckb�7�M�w�XI@�k�)	L��oR��1_���@3+�6�P�M�����Q��#��uA�n�h��]��\�r��O��}r���4��5����������]G��(<G}m�<ȐIj���wX���������O_,�ㅒ�.�T��2�G���z��y�˳_�4u>10�t%�Gz�瞏q�4��E�����6�YU�f%�\����2�#3%c2-��u��kC��gw�湡��G�p/�������9	\$B;?(g5��K]�J�$e�OX��ۀc��Y��1s&��	4B��d[���)�%=<��5ē�T2�� ���x՚?�Ǣ��ǰ$���=�h�R�!O�Jm��aG¢u���'4�����kg߲�D���W��`)!��-�px�e�һ\��Gl���۔�C'e��vg���X�(��Q����i5U꫘���Jm�]Vm�[C,�	X����.�J�Y����A�l���p|Xi���5>w^j@���a�(;e�c9o��͜X���A��߅N�2VC÷�-�-v�����E���u��-�li:����"o'!¯KZ ����9#;�Qu|+ؙbp`��i'��p$�Ʀ9k1�
v�F�K���1�ww�ţ`��%�
�l:�/��f��PO5EO�6�׭T����
| �40$���C�!�x]p):ъ#cn�����{!�'�Ӄ��֚eb�Pk1����"����6əq'�*��"�OԇouO�U�}B�g@M=;ɠ�n06�P�����+�0%��{I=�t���+���{���+�)�B[ܗ��j�=Z�Y@ ����y�@�'$�s �l�]�^�Z��l+�H��d�p��c��Iѻ�k�19��ٱ"�������XFkf9�iŭ8o$#f��%#�B[(�V�������N�ܥ�hw���r���R�\�[
f��;����K	)��1@����Vr��҅��T�E�ǰI65Y�4��i��#N� �ffX�f$Őژc����f��K�������(m"���f�j6F1dW��.���P��W\�g,V0����{�'\��¥�Ro<�S��~:]�j}�g�*B�E��*^�Hw��"GR��t�Q?�'�2� �u��}ܹ.��q�&ͅ��g�"�(û�<�eH���.��S�P^�� ���w/O!���D䯾��ᇄխ^N)��S�7�D�Ea^�IZ~��j� �.�g�g� l����@�X=�����xx)ۂEH��?�p|8�l��8�]<�d~Ne�E��C^3 d��{�:�������׶j��ǈ��ܸG	����\���Wx.��������$��K��Zp�ư�cV�/��D�B
�I���!�`*d���/�/�WUUɒI-�9�n����_ND`�9^��Xjqt;"(���+	mU}2�C1ZO�K��	��G�V����&Kl�fW'^j���dP��w ��!������V�l��TZu��_�d}�Á���/���E�z���Fp��d%��7�}��j��}�/M��j�DNmg}���� }� l���:�ʴk�N���bZ/��{CB���F.���!*HI,{^�	b�n�镯�:��4��/te�p�m���}�@���NqM}�V	4����8 ߋ=�\�o�Ku?�i��y���n�`�S�C��j�j����ĕzfMs����G�r1�ť��VԷg��E^A�qe�uhR���ʱ�Y�,mپ�"��q�w�1�ҙ@��j=��>��Z,`��8Y������`6�������&�&���J�`��0��FX��cv�B����8��Ոnxk4�N�$�5JU8�ɞ��r�D:]3f$<֥{ȷ|��-�8<�-ld�"����a&E3��g|}eY}��7�P̮�5��]�8xkq���
��a0L��������K��j����d����4�x������U��H�&��]���7�I�+���������M��3]�� �9yY�x?��f�R ����'���
�� 
�Z����v`r�>�,�Y.�=TT��$��B	s����ŴW7�Tهu�?覨Y���WEO>X����<~u�#ק�G���� ��>6�Zn�l�*���dysQ<}FS���?Mh�/��W�M٩�،m�c��m��hDXÚ�	%?;����i��H���TcK��֧�N�"[Ӎ�����j��&x�
"���5t��RX�wb>�f8�� �ʬ�ȏ�;�Ua�C����tK*
e�O��B.�|����9�#*'�T����|{�ρ�X�Lwk�$�2�-�͢Ucg>$��?��55�I�i����U���� ��ap���?�R�[�Y���,I�/�ջY�u-�_�؝yKM��"�jf5�,��ݜ�皧�����z^`���È��(nC��"M�Ӡ���{=;����Z;�B�/��Z���]R}}�p{o��$��, �_���ڟ����9�?�Q�8���`�2Y��U����������N�a�ּ"fV�� g�ߊI��4�|�e�?W��4���L��uy�X���h5�j��4�D[�c��.��L#�c!;���OӅoi5�ʮ���Au�+��_
�� 6*FHǩ�ǰM�ץ���
>�,"[ ���/���OwX�A���*�p���L[ܨ��=#xK��k#(�:�05��s���_�wc>����)�1��O�J;w����im:�Y�O§�"(D��߱����=��+(n��3�&�����COX�|5��#���!6N\�MCۮ}�N�+K^�2G�d*��R:���T�r�+7��zWO+Uk�h̅���5Ǣq�_�>�-@�i�5ı�o^��S�\��7j̪4��@8s�7=�I��x��)�g��M4�;�%�8;<	L}�Oa���xe[���t<��n�«��V�`�OAR��	_��h�f���@D6��t�8��4?I����5� ۈ����
�]��IM��B8N��6�L�ۻ�p���I�
�y�+���c�NkwK��WDVBG��s�BH��#o�'�E��˻$�
~���gѐA������2�1�ם}�A�Gy(:�_�Wfg_�~۬��=W�"�_�A	*�4A��X]��^�����_A�^#�be���U>�u�$��2�.}jND�S��GBԱN���1:s�դn>-u��-M�Q���]֘��s)���-����~¨C���ӟ�\l9pr��:��f��2��g(��6}i�גW񤛼��[ �^#��m1Ù6N��HBT���v��]����[����h%*�T^8�9ͮ�*�f�{:��QbLi.�K*Ao����7K��b4J	a�5�r��7�LF��nrzi:�r_d��-?�-���� �#H6�~� V�Y�Uh.;�-�U����]FY˃���⃃N��Q!1s,�[^|������Q;��[4_�F(*���K'-Ќ�� ������Mx��o�u�>T�
�_�Vu>c�O7 �	�w��Z~�z�=H}�ܡ�;3��,����y߬��H����	�G���Q��� Ҋ���k�u!q�./�՚\މb�!Ŏ�A��UH| ʱ����q�-Hr����71L��T�Za+�r2j���CYU�iM  � ��2�H@�^�������>���&$L;�-��}.e���e7�B�t������}4E�W���K��xX'n�<*�C`
)/Ō�!@A6vL�����ߥ։�=Q:��`d�W�����iU�>�x:�
ղ�:%��(ߧ�j2)i9�`A_g�%�	��~w��ڹ��N�N�S��i¯I��F)<����~4��0���/���(&�3�S�9)��V����2��1�C޺��f�Uh��3?�'����x�9z�{Xd����� 7k���!�?��d�����4�Qz�Xф��1�9>�f���
�!�ȥ�����i�������˩���t�����ͩذGy\�,�[�_^`Jn'��ӈ� !�b�X��t��W�����0/�|Y��֯���f+���_xo=s
�
�?����f�"C�مF�L�۬�'��z�����r�_9w�=l�)?X�'���2���]X�R��Wa��p�M�9�p��OD�6Y�zT���,�
?1�:�fL�by
���?�q�VM 	&E���d�~���Q2#��mhЏ�1D.>�U/��������A%+�ah��p�>�+�Gm�55�򧪽��<�����QX�n'��R
cw�����7pn S~^)��':~�ȡ�1r]�F�����ʻ���a?A��N*6t�Q�X�!3NY�$W�ؤ��AG�p�)a�f�2�b�V�����nS�?<�,�5Y�6��քR�ҖV(�Q�㱃c��RAǓ>Ճ�ݓ3o�~��
__�R�LD
z��u�,��C�;ެO��e�>�R�V&�n} R��9�)��A`�=Á:���%}�]��O3�.�Z��?�o0�f)6���ي�4�o���y��$�K��sÍ��]�Yd_CJ��ǵo�xs-?�׷���p�����~nm��LMBN�gėzƠ�aѾ4�|���K�k�����+�̞+&��g �s��}%N�a�,��0�wb��tA~�[QH�IP��d&����*�TٻT
�Gb�(�)���q�28�ϼq ���K��V��Gԏ��h�^���� h�P䛡W�ˣ��_��p�A|3˹�w ����Kf.Z��h���g}H�Eץ��7�YHYxQ�0�sZ;̔A��Q��:(ݚù�#�Kh� �d�h(Ƒ���qw'����p}�H��Rf��w��u'Ñ���2F#�7B�fK�͢����@���N�酁��S*P�}�/�P��`�#*U-�}A�g��b�6K���$#�DÌ�:s�_��Y(9ǕO}�ea�Q�(�$I\戏��t���?��J�}n�Q.W�Gt"�.��B��6�0�N封1�!--�]���D�˥qr�0'�&��-�ǟf���`]~��7��޽R
��AW�s�k��M|\d�G������Fk�]+N�39q3�I�����z�/�"�	'�?~�DgڏsV#Rb��� �m���[��b>�G_R��GFOlS.V\��	W
`:�lg��\Xچ�-����њ@�f���p��A��иU+j
\�.�v�RԾ�������"S�>�N1�'�m��S��Y�&=�J����d�4#Z��(ΕWY�v���G�!��N�i�y��r��/9�T�S!7����	J�MA���������z�}�B�{#b�Qo�A3�ja@ �Z����&x�p3h�oKԘ��8r���e�S��^�ʉw���3�� d��A��hr�����6v����Ӌg��SN��fY��;<İ��Iwf��.��KD�0Z<[�9��Y6��g��Ms�s!�[R�4`G�ӝ]zڛp��CJ}��w��oЏ�]>��i�@_�%�R�.c[�dht�G���`q﨔P�ce.\x�*4K���"����
��8�9�����±Jx87$�K;�$�S~�t�:���N�dy��37 ������0ǌ�~�Aw S�1]H���.=�$0�1��W}�0�o���!ف?���M� QJ�s6w3��������>��i¬�+���T���2���)6j�[L×@�E�m{�jn������/\Ħ{�?+�T�j��S�s��w�L^�qI�<4
�!�[��C������k7Dv��e�?�$�5���۠���y�	�l?��ab�ӗg��XC�>�	�g=�h����%�uv?,mYze�l��i�*A�F��+��MDٵa�&��7��C���%t��tMs���l�.�H�? v�[�(aM C'M^v���O3A��ʾ�3�=d��M@��JC��S�,�\�r��x�@E�$�9r�)�	�'�\�Be����H�Z��}�3t�ǵ��-*(e�2�B
��o�����J������lx��F�����SD;C�^O0Hq�����r�_Y��I=W0��Sy��V���t�9
b;�a�a����_��� ���fo��b~�!��D�Ҷȅ���H�̋��0	1����Y�\�n���>��s��58Iy��rq.d�bF��x�X��${Epc�o4���Cij[��9���9D_Ʊ���� ���FZ�21�O��{	Tnb��$�bFu�M�Qj6c��?�.!�ς�����د��di�c���m2j������^H��7����@]JH�
�:� ���]�.	�1�Z!O?�W\��Ϛ`p��߉��2C�y�+�L��A���N�&:!�@��P37������ԋD�#X������*O��?!���GB��v�	�ㅛ�'�}u<�5ZQ�C���"ٖf��U�"��TN���)������v
F��&��&�a"C$�7̉��ô}�SoVF@�tlx�������H-�+��X����u@�$`�f",���p��?;��ۅ��o<n�<�9�8�;Qgn�V��B�Z�v��o�̓>���1>
�+� �����s��1�R;�S��j5�Kވb�G�J���Y�S�F����`�̐F�(B�&��,��J�˺6 L��r�Kо$P2���UNΎ�E�O��~�2�/JyHAjȥLhTO�����y":q-#�kٛ��9I�H���]��9��B=o�`u!�֐�NS�� �4:%�6밲|�Gћh �X��Da��&�-�*Ҍ1KN-`�Mp4݄�P��Tǝ��?u��� ~7���W`H#��E��G�:I�
Z��.�Zu�x�)6\L�~�3?=�D�N�E�j�|���m]T�oaB�. M��tc��;���
�bo�S3�̾�e��K�}R�H�g,���{����w|J��?7~�NO�������1��;<Xo!������T���V�}�'HI��)~��,���δJ�~��+~�#��|-����+/EL7f�\�������w�b @tė0L0=�<��_�-�(q��Ñ
���除<R	x�l�A9�{����Gv��Z)��pdЌ��s����N�cDgJq{��|DϒyL ����쑇Q�CS��"��oȘ%��ć���H�O����4�Ɯ��f��mD�j�"F��:�7!����E�r�nD��s)��~5�^�|Z�ob�{�Y�z� NIbQַI�J�|�r�e�7~�v�8<=��T;��p{���3I�M��8�/��q5:�utSn�R\y�wˡ�c��)]�Ka��x#+��@`uC����u.f���m^�D���6%���z�"�ً^�I	-�Ӌ�r<%Z�������ܵ�|s��t��D�>#�k��y� U��Է[�:��IEU��lMO�Q��ϩnd�WK��З����hB`�N���H܁_On.j6�S�� �Հ��l�̪o>n�h�*SݤA���J���d���w�]T�I��<")�+��`����2`ޒh;�F���7ޞ�{d�a.e��Ї���Md�u�6o:����z��v�e$�L!.J�`�pi4^��"$ƈ#=��Ǐg�w���2�[������dT`���K"�f�����7vC8��� <�C��q�I4��9F�P���񔑯t��[O�7YムE�'�eUg����|X��O��� p�fQ��x�5�f'@m���H�%����ղ��e;ed����/�*^���>S>=b�R�+��Y�Rﶪ-`i�`��.1��%]��0��W^1��[�A <�$H�4YI�+��I��c2��.�X;#�j#w�f#��m�����ȉ��̜X㷷돨�g��թ�Ϥ=4���/�z��1�P�؊%���J��m��f�E�+�c]2cWa������4b�T��:�]�/�?�����B��ݛ���\^t�!�����]�v!n0<d۩Θ�ڛ��}� 5UcѶ�H|�\�Cx� �q����P�a���8�7Z	)s'��"�=��3�����}* @�T���Q��L���a�o�0�4�~w�dSҡ�௱��nt�\�]��6w��B�!���睾&F+*�G���#���\�y���~q����5GY
����G� c��Zgq��H�1����=���	��bgf�X���v�@_|�	�e&��Lnȗ/	�=��� ()��&��`Ny���=wA6<�ѝ���c�7��5����Q�:.�s���#6ǡ_TE�h��m��kC�#Oç�D�mR�lY���!k��u&h?l���>{P��H��fc��Iw����5����@,���'�ToW ����F�w�!�DW��I0β�AZ�&�M�\�(*����'-	���lO�1>���s����[����<�o{^�]����7FL�s>u}�����.E9 �GieF!��*$�V�Z�%�֐�W_^|�G.)OB~0�A���i�����P�d*~�m����2�:�M�%iG�v &�7��n�BvK���5	���B������@([}��g��j;��N�=�ѫ;z�=/�\�����&E�Pߗ�D�QXSE���$8w��i3����E�t�۶���l���r���m�G��|Cu���w��EM���Ơuk�gx��k��.�ܗ������0~rӥF�8dd��z��,vd���G�<0#��h����9��H]�Q��q��
[�P}$�����+��e�m��C$�l��<L�`���dcb~�|_���G�s��X���������Y�X-����-�v���b] ��	E��T�~��?Ng%8 OgFg�D��T�Y��W�u�z�j�މB��qa�K/�â��Y������|��ky��y�q~�
��Qj!I3� ���z��A��r`��r���m�-�P�i��T�QU����$&�"��]�<��O�������젢�Mќz���ά� ��E�\�䑖*^_�v'�u��U�A����P���O�`������T�֨�V-.�O�/5*����,O�����pR��(�#w��������5
�z��)����vX��X��o�JPWd����,�%%�����;J�+�2^��G�&��dq�;��k'��;M���z�H�F�n���r��9�
�}b����'ߊ�vj�y����p�;�ܵ<�>Z$����]vD�j�	K�-���U$�;�G'`=�T��}�X�m-n��Qe��5�61��fM���B�|х���R!<`ѕ<Bڅ��vV�z��ِH!�ԑB�jI������n.��T֌��//A���:�t4� �9��^�ǐY��#Q-FS���/��pss]G�k�A<���2���"��7������j�{O�e�32@)0��~G�+w3��_bb�v.�?���Q���aZ�Dϭ%1qq����%N����<�xb�K�>���)U��ۢj����i�P�T�0%]�X�tyl�����/\��(�I��-���ԡ�ЂĈ��ڮFF�����g����!�o���ܢ^řYԡ�.8}��UYl_�A�R��eτ���|;�U˯ӻ�&�WN�B���n�'Y���,�L�oǩ�Q)��^{�P������ݷ\��V�%)UX�f?vq�\.��'�������l%W?���gdT>l	D�GLD�+�aWk@JQz���Ô� D"��;��Kճ���{|�Q��e��޽�%�,���2ZHʡ+`�bQT�f��*Ƞ�����I���ǫ8����Bf�1bi5��fh���*�ɵ*��s�݇gޭSC�;��W}�2�����#'+(��Ů���Q7rh���� g�&��@Uk���C�;)��kG��2{]�zO��l�������}!���Į�"�K,��K�F�^fLR�j�.~��Sey�4%�ݠV-�_�ņZ�����]���#v�뇋��-o7lt�`	��PrE����� ����}�ϏkT���[��=�lt�KM|f[��
>�bE�V^]+\E��Џ�Y	`�<A�S�,���BQI�2��0�`u\�"OO����FN��Y�Í���ԇW���2l����@�,΁7��y����B,�Ft@eR�o�y6�d�o��)��^=�`��I=����܅�M�\N�X��y�/:P�)c(��!�b��<��E:���O���׊ǜ2H����QY��M��|��ZZXR�v��Ʈ[c/_A��%�mD�z���!�7�W���:zh	����:�k9C�8}����ӧBN��H�� ���b��G�21�{W-/H럣��vG� w�K^�li�ա����Kh0-��X�:27dV ���'�����Q�>��-���-���ĵ�K���~}(�t���������-B��(�l�}oj�
!�B�Sŀ�,�Xڭ�\̓f/q0�e��ϐ�l�G��A�aZ�Ǒv|C 5���8�<A�E8S�\_�P����к���*�ݷݷ�����qK��^�"��~@�'�& ��K�^��+��o���u�%-W���#\	_}ɔ�;gm��
�7�V%�
��,��2��"G��i0��0[AI��)��l�`�O�O'
X��۫F��������q(���a=�a�)��qo�aB�*u�v�}����ԅ���h492V�*�����]��T�ܼEU^��r��	т����:*�"7\S��ݩ�*=�K���Y�#]�aeԡ��ܨoLc���3H{�0��صP
�4��+C���mgO*�l� �k-
{����XR��m>r�ҸΠ���l����_��/�O��dJ�8?E���6|,�h�5��6��ŒY������Im����q�#ɗ�M�)�(1}����H��A��G���9���&���$���9AM���%��E��|�"~ެ���'���BĆ�n�@���(�6��b�h�`�Qv�b�ύV�U5�;��5s&�I��/l�!�y�Vﶈ[?o �<�a�r���rS�Q���Gn2�x�%N=
�|S����P�Sj�M����E|����b&<M=��A;��p�����ݮЇH��gAQ#�]9P9ʠ�u+G�:����b�����}M�}��i�/�K�]�:�W<��i}!b)�>��ƫ���-�g�������^�}��SHXڈ��`�抒�a�������JsoIKN�����z��e���K�M �*�{�{��wM��촙XY8�}sجI�UZƟ��T��n���ࠣ����c��O�~pJ��d�!�F�\�yC��_� ��ֵ���ˏ�$�b�j��j(Ϲ��\����[:�B6V���Q�iI��$k�b��R�k4TCٌ����[EW��.z]�I���@���y���t_0!['5��-!����+�e�"�)	�GN�c[�q]��}��}K���܋W�9"_;��m�*�u4r����O%ݕ,�h9�8�ƕE��0���0l���ʿ�(�7}����[� +����s^g�euO�Ǭ�@���a������:�����*���@�.�M�ô��)�����Ģ��[�c�x�!΋���+A���я�0���p����s ��9+~K�g�5�(����>Jd�gR* n����S�K~�� +{x$����.��,q(2��y�F�� >��q��n��U{­P6�Peo�����߸�7<I̪Ep�S���rJk��m� ('b�Qko��}�N����!��_�Q	#[�s���doЙ��C�k{�CP���Qʓ�X�A�u��t���rks|C���C������{���6���#��~��ZUc/�:t�ݍ�M����OF>��$B�܌ƶ%�8SV��_�̈8�¹��/����.����c�W��C��0�i�t���
D�=�w&��;���m�h�+ ��u�<�c�Wr�uy�XB��~-�M����7��2����wi�Sb�.~�k�scA4ɮ�%%i�O`D�Q��:�]�8�b�r�{�d_���+�8��Y��0�@�|��?E�����������p��p��@�F�0l���D/���L������0��GÁ���\��w�zW��&�ui֭�j�~p�����6���ƺ!��sm��Wrq�R�O�>�&K��qt����z�+R�Y�f����1?�Y��M�_<Hp��/�8�!KUNa���1ĴR`�˿�{G!7[*.#�o��		����Ϋ��ɗ�>ו�$Z[jė32�T^~�sl�����94�7�<p#Y�%&,����|͎[vZ�]	���`�x1s�������a��� �x���N�cr���9�N� ��o����:ѬBU����z'fr���iRpvw�(�z��|In:���_
�v��bqY��a�]1��C�7p>fz��w7���N&�}�'��2�I �
������t��@������gV�q�D7���V�vm����6[��!��������wf�Ѭ�1�L�H.��i�M�2wx�� M�� �%�⽔bk}�]���-c��;��Uś}��i���<p��*2�35�
Sa�Z�Q�в�%P�a�["'�X��S�W���G�`���:�&|��>e�Jw%�n�\)x���C��������ʰ�7dko����#��.ȪZ�{g�u��:��įzx�WO M��,?��/�K��Z~�^𲲀Rz�צp-��~��)��0���%�WG�|��C*�ơ��nX����6��'+��(=t#]/�����2<�����<L{���n`=�����3�T�iI��7x�|s%f��4���5�:�ыl��k�Zc�V�u\�>�����n����s����?#W����Oq���ԅ{�n����c��)y&h�r��%�]!��@��ߪKKCC����{�d��K��'#�*��mZ��?E�� �a/V�a�W]�Z|�x�drl�#˖c=x)I��`s���3��c��G��V��K�ZԺG̏�v��Fsxc|\�篿�F?��y�)5H��rk����o���"�*;笝�����4l�����> 0"�w�tտ�`o%�;���{��4�ܿ\j��V�vJMz�����ω��Iyp�t���g(�6�t?%AR�v�Q��5�7��2��;ɮލ`�?�a\`w�����s�'�J��HǳP��gNԝ5�`�2f;U�i�-o���k�PN������_R�+/���N�!є۟p���ɠ�2V��Z)r��\t�r�n��)���v�6۳LHʕ E`gV{99�I�j-(CK��~U�v�@�;�}���GfERҞ�b�͸�{��>���&8G��5��G�yw��
�Z"`��;`G�%�k��7ƫQl��)g�����):b����Kt��8��7h�~p�M4���¡u��x��Ɖ ��k֯�i�٤�Vj�,W6J��	�h�j3+���y�e���u�;�u�0��[�^��� ����Cgp
T��(���� ��5�*��pĝ��″������g���n�DfULuWP�vZ�*텄 ���i��]��-�ŽP%� �"?�VJ��q��W��_�qx�Ϧ����a�]н�HP�ԑQ�J����l��jԙX���b�.eDW �� 
�TgQ�I�r��׶�)E�Q6�ܪS�7��`�q�Y��nT�1���
�통)�_G�J�K��g1��+�����	��3@�-��]_�������X��i2m�9t�(��H��<0�Gݦ��s�pw���i8��P�<�R�8�.�VY3�gD��gV���J�H�JۨنN�@������Kנ�Bp�66_s�X�����I,�ij4=�&s�v<Px?(V=̛&Q�,"U�
X{��<�U?)m�N!)�f1���x������"c�;��jT7����!�4��x��In�A���C;��\Lٍ`�~��D��^aY����c���+�P��"���sxC��p��fe��y/o~C�M�yh����������(�2�,#ȃA^��P���#����F_�e�?�?/��2H`�~凅��(�\gX&m6��o�|��K�v�{|��(�#~����Q���?���L&��3x�D1�jɕ�0���3�ȳ��Y}�$I #x0�)�)e��rͿ�&����E�������0E��Ɵ1���!4Kt�:��2�����OK��_�`�
�B�HB.�p��P��0+���ou�����ʦ1}ь�EJ��Ǚ��@J9<F�����oN����ǳҘmwBܦݚ�?������e��~��X���B�?���9[zn0�ov{t�!�V0H��m�q^� ����`���m[E4��q��Ә�T�"�ͣ��hqH�|�Qպ؟��=�)���>l �=�J���XTK��< �¦x��o���2RL7@��!k�U�Yd�&W��sJ�l�U�$�в$
��w�%�ġI���+��O�Rm)%:��#�+SD���V#�%O�|�&c	pR��tF��9G���{ 
��3V� +��ǚ�|(�~�ʂ��(m�AVSkK6��'I�
q���дi�?�).o�on�ɿz&m��N�(<���xX�H�{;i��M%UUe�)�&�	Z��TRb)��S��i�+E�����`�߀�˯^�G	ZD�*J��}��lXy��I�R
Y�_����MnR��^�-6���{���(�30��Wp�sÅ����VV�����Rq�Y�BH�Iyo[a�>:�˿I�SxB��
������A!��R2� UQ�kfڏ�Bz�rߍ��̺ b���Iu�<a �5h�(A�U��Ӯ�Lp8X�Jr���'���kΡL��N�"M%�}��?��Ow�ОXnM3�����̲~߄zW����p��^^�)��.,S�:��AȀ=��t�5��\k�MÊS}$�@��5�E�v|�%4'��$��wh@x�
k���91�`�2S��6���KS��E]$���=M�
�ih�/wG٨oMy��U,6�;��\���3���ȴႱ��4�in�{��zq��eɘ�MsSM����[�T�Ό������WIV��-��l�N	��8����� 
����d��&��I�%�)�g���k���h~�G$�65�f]�N���+�*��]y���|w��s	��1c׭҉���f�@7��W��ծy��X�A*B#a�t�E���#�
���?���6��D���6�/GS@�S� ��`��[�{6��g�p�ö.�;4z?�̢��
�f&?d6�0���5���@�w}�L�Q��Fp?=gf>Tf��+�&�zN�� ��>��N�9vB�[]�n�֗`�z-Yvg���8��֕nG�W���aH������i
�o�B㕡Hձ�)xw9OJ�z�\�)2{)'"+�ƣ���=�i�v�8)˘����r�����OE���y���Yd�-���D��%Ո�G쌹��F�3����6 S�wJ�O����5'is�䏨�Y:��d�c��ed��C��V�6>�d@����>j��ۑ������Eغ �7_\g5-[7}��?�T�`hYnT�=�q�9��C�X�Ƈy捹?�� ���(g�ߘ*Q/�,���i��J���:^�ig���>T��\��Q������\��QV�m����伸�#$��:#�}�f��Q�X��04e�u,�W �$/v�I�8�F �*=$:i��pstA���T�"j��ӎ�Ht���#����~X��n�7����kr�V�j�Ӈ�R�P.����_��Q>�'9��g���5�Z|���;יdQz����\mqn=Tp��vɧ���.�8��Y͓յ�>9꼡ߵȤ��C^��[�Ŷ���9S��ha:�~��l<󷝸l(��� ^JD���E�8�������k�gX�24�У�V���̳ծSIq���?���t�[�3Ӿ���7�E�bkaV�����^wB�yJ:1�u���1ǭsܮ �֋���N��m�m��+�F38�S1d���5���dg�~�(@Y���#ϧe��i�j���Ⱦi	b6��Ǉ���[͛�o�T�>0?�К��=�� Ο�K1WTF�o�l��o'cf����)_���2�G^m"X��t��^����h�5<&Ж��~w]�_f�7�ח4�^7�aVyI��Yx����d߱��	���ݓm�������,Y}� ���� zT�U���!�jb�?�������˱����m�NUĀ�Lj��]�"� M9�s8�?2A����~o���Bu�*
�@��e�o������ b�k��>9�;(�����l#?��p��X���Z �O�Z�
�Tt�O:L�4I�$���+P��8�:F2��rukW�=	7�<R��u�/��7�?�KssƫD`s��xޞvbN��B�An(�@|�p~�i���b�k�9�=;��ڔ�F�o�q��mye��4-��!�`����f��-��<��vXZscpf15�xT��ȅ(+�D�اa_QF4b�Et��^N��n/_ʳ�Ir����?ﲥ�j+�'L�B��f{vN��^�����zR�X������w5�?j�Ҙ��r�
̼L���)s���!��Th�"F"*B���T����F�]`�S��mn9���}�=_����<��e"fX3��j'<A��VB�r`��^L�J���S-��P�~�+/�z�y#��1�;3J��f�������Q��֡ӑ�s�O.|��_�M���`їd�o��x|E;���!��9�M�W����sI��|�w�I��S.�wyُ�V��Nt�܄�5t������՞��A"'�����b�<}��,�Z"!T�J��P���~0���)�I�CT���!:����W�  9N2
�<�1���Ƭ(�<s5��=�պ����	�el;?��J]�E�C=�B�P3�q�}ƨ�W�β(g�踕]a�~#���w�@[O���[�UJuJ};3<) �W�E4!�z��K[�E����,� �#�K�P�QyUV����Z-HN�}f���vM3tͨM�0�ާ(V׭!�	�D���S38�7+���(��'�"�;��������fS��d6ps㭠V����7�?�Nћ��ue��I~�j���=+�^�@��;�2���_]{�v7�s71n�!��)#
Vt�'L�t�@��{XS���WaH`Ɇ,ծ��3?Q-��
��Rr?�;���ؓ/sF�G��di��hՒ��|L�p�)}�Gv@C҈�CV_7���iY�n��N�����v!c�oc��۝� ;1l��8�L �y��2]i���Խ�O��.��8��fT*6�YA�Ͽ������ �j���9����hW.�f2Of���e��:��l>�y-ҍ����Y��h������F=�n�jW�o�� ����d�J���}�xGyk�g��;�3�V�� �w׷� ��(h1�	<o�N��<l�oj6�V͵CM�\-+�%���CbR�37��S�N��5�r
�Xl&}���|�G�Q���̎	�=ԑٯ[���3��N, �<8aP������VA(���$ص�c�	��s��aX��(�����=��ъ[ز%rZ�m<�tU'oO��n���\�˘������D�!wc8	´���(��̯����o����:bt9�\��:+�ܑ�Af����V��+�� ײ�us�R�<��aP>5�@�)�F���e����(	�P�.;=rMւ����\�p�D��h��� �$��� {5�FB�[Ω����M ��6�*��Z&2KY�|ﭹ�_h/t`��(�(*��m��h�;��nڢ��@ࡆ69R6@�������O�ɶ��.&�Y��f���������g6��.]�Yƥ�t7ȎNT�Lr�ع���C�Iٟ��n�������l&��@��2zgg!�?R���ȑ?y�UX:�P��W�-��`|#`r?Ţ��;5@.'���ޘM?9Cmyh��-���G<Q-�4ó�/�n�DRKkir�j��繚a[(��k�_m��C��r�&���&��<`�����M��_
a�4H.B�����=W��,;�So���5��o
��lG+�d|���
Wg����	��e�E$\�>Lț ��Pt������%+{B�<�������{U��eq+/�X��Xo_���-��_y1�o�xe9��g��\a�|ƃ��v����h�t�Q-����ΟSg���b��9N�$Nb��p�x����Z���pbJٲ�T�v-�-��y��e�V�(D��Q&޲�s�n�X�댍6#��n�">:�𾪄�9Q�����v��V��D�oW�����nEC�������շ�o5�q@��6"��5i��-��i��m��FH��������BZ�l9і��Iw��?ɥ�1'��sӆ�L26��i�	�bS������Bu�z%���E�,�HL��{Cᯞ�3�V���I;|L�[���/o<��^����S!�fto՛��N�ɮ2h1��p_Uvy �(;��`�:V�����ܠC���?�4X�3b����F��lH�\J�|���6YW!��6�}P����;�g�=`\t�J�}-��8x�޿�7�;�(bfp�'ZPC���;�lB��x8𼭢�H����(�!�Ӭ�!����/ i�;�b-�E�j=̷�(qiчW��j�
�����K�d��⮫�/�"=4���mɏ*���=$�Ey���m��(��wR�)kt�N>����s&���J��p���<��:zO�kNc��暃���S����h�#Rߙ�7G��$D�%��� �`�u{|��	�q�=w�~���'D�l��;g��I	�#���꽢���.��
�H��j0�a�}' �VX�J�64h�D�B�ag��HN@�r�t&����r-Mѭ�zGJ��61>��;h�--oP��>�O��vD9��e
�=�����R�q'C���
���g��Tt�����MezY�Y� }z�?-��r��JO�(�_�����l�/i=�VB!$^j�c+K��M�%dً�7D����7�F��H��!ik��l�����e7�̄��Y">�eR�:;&*j!�Z�5�']��%N���"j�����)��S�$���9_ٗ���&5�kQ�lWEx�g��_L��#'|��@��2<HC�@v���҈�+Î�EB�Ĩ���.�0�������c��D�P��!��UP�4����~-��&"�ӡ���&rM��b�10+��x������ꀆ����~P Z9b��Y �u����q�cV�~s�?u
�Vt59%��/�'ZR{���E86�A>-[���ޱ���������iF&Z̸�/Ya퇇K��` -��O�ŸE��e��F%���_�~8CP�B\)��-�?i��+��f>[��4	�A���ޗ��,��ɧq�ZA:�vGX��c��e�%��-8�Ui��Ö���@�_�/n���o%^��S�Zu������hg��W��n���S�wJ�Y""ܪmY��W	dappGx%>��ͥ�Ko�>��0G��k3��,�`-��vۼ�0�|Ҍ�4��ui���t�G�9��J1e��(B���!,L�T�/�x��gVIH��}���y���n�P��θ_���~n�~p6M�FՂT�2�T���zJ��(� q�<�V���]��ˊ��c;_�ֽ��&�O���u�������h��`�$l���B��8�L�Ma�,��p�5�[��[;�&(�7�7v��CF����WI���&�X��_$jZ��v�ve%v�"=��Q1I&i�b��/4n%��[:'�sk��{	)�pg|�'��2�I��	�f�5=�Հ��/6M8L��8��*�~V�H,�8�eq]e�p�n#X�A^�+*b�{@�	S�R�-��: �kU�A[�n�np�!�R�;Pj��%Zf,���	�J���g&J����]`�Q���[�P/~��m��&�BmƂ.�oۛ�a�KL�'5H"��v�ϛot�5'��в��F��ƕje��*�7;��;k�b<��@j�=%;;��XOj��j��;o�aa!�p̪��XgQ`.^̌h��z!� H>�����wl�[�f9��ϰ_��Y�����'�zB�W0���;щ���>Kyp�k���QJ�a���MI�o�ʈ��+b������j���/H],$|g�X���-@ 
o�XU��@��Yv�42أN��IS� �}0�G[��������mI��D��i���z]�=�_�� �O������ ����6{�u�k5�* ֹ���Y�����W�܌b�g,��_'�\e8��/�-QL��,9@5���W����=-�.G
Z9=�z�)[�߷�����r�pa�h�8g3��̀X�R{������ ���S��(��U�9��C�����o&Q�6"Hrzud��3�H\Zݤ�>+��u���#�Qe��]���>%����e��f:�z��Z�/\��� �	� ]�Q�/a�Ux�W-β� ����q��;��-=��e�$�Db�^���������'��.��_'2c'FZq�2�sn2u���k����v���i��Lc+P=
"��{�� +O���0e6���q�L`6�V�k<}߄������t
I��^���f��<	#!D�M�2q�8wT��DXYwѵ����ѹ��� ~��J��<}�`߬R�	U����Xk1S�CTNq�Ƈ�<~L܇E�l|.�?|�{�k�5��03��&c�uI9��!�kS��i�@P�����ܶ��'w�e=a>m�YL����\#b���D��#�I@��Ni���u���K�C �q?�C��`��͋�*s��;�?/?t��V}�^��GwA���+�^3��Ǟ�f���@�I�ֲ�Hǉh3���/���8��?���__77L#feF�LF�s�������f7�iEk�&������"S%y	�����\�_�'�!��߆��ʢ�,2����ڐ����Q�bp��7Q!�usIq��;�W�iIW���ˋŢG1�[-��hD�e����M-&�W�-D��
!pM�^Tiزr6y�LO��ck���ʦ��J����[:�?a��a��iS~��<$V�#���"����\�MX�Ь���4w7Rw<sb^�"��C����w�-�2ܨ�F6�J�i��A;N�&\,�|!Ʋ��u�E_ Mm��K��S�`�	K�M�Z�"��A���k�ݚ�%FDD�s�3Z��2�WL�v����]�}��}q��F��!��o���%��7����g*)��ڍV�|�%�7�P��%�$�?$X�¤eݳꓐQps�b��,*�j�v��'y��c筧?w��e��;�ܽYF=뙍rVF Y�
��<��fuV�%K\���Uv@rA}ՎB�(�}!�)o7fZTA�q�ѩ�=�8a�^5"��6�������Ar�f~jz�+р2�nY��em�&�)�������A�B��uC��~����`�� ���s�"���K�#��.��nIǊ�'ߙ}�QJ�k�Ƒm.��#��m����j��-�Ș�Wg�Z�΂���BɻT(������q���hk� �Y��XCC�9K�)!����él��!7[I��n5g����0����2o��N��E~-=�Juc؜6s|
�����N�s�nJ��H^��g������kH�s���M��
:519�)������CQJh��M�
G��I(d}�`��|�����PlvxA"������G��ap��zB�P�A��v8��KW �0aF�As�\��NҤ�4 ލ�:��+%�8	�g����Uc��/�f���`��ښ�/�HF��o�ݶbs� A��|~Ӛz,��@5C�yr���<�ʚQe�J�U�#C��~-)���j�h��.�	;���n^�E.�=q��X҉�R��|uM|Щ���K��)�8�hx6Ř!��˲i���0��$�ݐ��4k�%5��� ���_�6TɟR��ʝ��f\��� X�?�	+�����`<"�ا&�u�64�({����?��d�����!�����F >�( ����Ag]tj���4�Ƚ��0uh�*S��]L��	(pｸ�, �ᕿ�O�IY��D�H��@�!# �n�ZK�T�H/��Y���]�r�I�tz�E�ݠ���2M�ۏfY�M_�����tX���w�@p �Q�F�A�r�B�3��#�ӿ�H:�M=<j���"��v�7�2:H}�3T��co�>g	-Z��p%R3j�7R�k(���t^I���Ő	$`ȕE�q�!G �{����Zk�Vc�F�#LOk5u��xy��U��Y���MndF
����O�8����_��]"Xx}l���k�@	��B�n9���@�a�Aճ����5������[�mi�w�Q�l�dhӥ�q�Z�\��*��q�ND9WhvZ-!1��d�.c�c_�Ĭ�2��;o�e��� �L�ܨ[Jԩf�A�q(MD(�<��|f�����_� n8���{ĿH��Q;?Y�> �?ma�:0��H��
,�&��P0d�X�#��i���p��m�W����&h���0V�v,�!����"?r�!�*��<I���I���������%NA;�I���o,!^�.|�w�j�g�������oƿGP��.�`K����c� ������E5
8�t&�,}��\��PB��(V�;NBP~o}�dhy������ݥ���.b����#�,�c�ba"T.�ϳ�v8&�����u�ٍ��5��ʸY7���0���c3s��=6�Y��:�'a��4���\;�a�J�Υ�r����q,R$���I'�H�/�ȳ��r̙	�ʣ���{ĭ�	_�=����%,����mھ�=�=[:B�+�Yt�6��{�sw����������`����kw]�H�-'#sb�<���>2�1�.��� |80zñ9�C�:��.)��"�%ٛS�?�	K(�L<�}�pPX5�T#�>[ם��m�l��ۯ�ۆ�Oc.y�>= ��02�6Ye�e����r�N�5"��<�Ğ��y��uY� 1���nÄ{��Ȯ�~v���kME\2�t@���B�)�J�G���3Kw�~]��l�9��y����W�Ԏ����� {5���oN�u8��M�E�y%��=�.��� ;Rٮ���.e��O�Z£nÿF�GD	� ]WA�'�Ξo�Cy��{(����=]�|����oq'��dk������e��y������T��dexC��Z'��ם>��!�k��62x04���W����'j�����u�r��r�CR�d��Sc�5��C���xL�n�g�>���i���� ��J��#��K�3x>�(rGC�	�4�6�(b�rۣ��Jx��0���-=T@�ͽ$�!Y�Z�,�wH�b0ܣ�� �*5��g�s}�%8�T�����l����s������b�r�˄n��=�Zh�+� �*Ѻ���w�S��
��0]L�	�NBWBN����!Q^¦�Q޺mp@K [d�:�8����/&�n�������� ٠��~��D=��*�2�ʷ�ʅ�e�~�n�J�N/�ĩF���NG������cd ��������vF=��.���j��t�!�J�_hP�k;w����4�4��L~����	�����3{�pE-�;G{�n���u#Y��N%�����q]@\���u�+��.Yv�0X�^z�g����%�'�@a�T0��F��,��3��wp��{3Z��!��<��"t��G8 O�F������,\t���H!ذPC��S�������Ϯ�cX� �GZzͦtο�8����Ѣ��8v�����#i��wV�����؀�~mt�t�ud�o��Zw�е��&3��(��0+��A�X$�wo�ۋS�D��nDt�0S��*���à1ZC)NW	8Ie'��E�^����e�Z���n?Fz� �I��8�O���1��q�tı����� η�[��_?�2l%�CSS}.[��=�]�]V��dfR��X�����QH����{!'m�;pF�`� ��Ⱥfq]b���2�V]��*[� +�Oa�>h�O~B�]�DC�06����Oni6�O\j019�G���od���`G�I|����	p%Y��Dؗ��L'��I�P5Bķ�~<�0���㥋p�ǭ���3�n�y'U��
>��)-z@��n�r)�v��<K��.aϒ���g)��,jAFu\E�����0�
C��E%]�d��w����lM
}�o0��X�x� 
��(�Z��z��2�z
�~c��x�L����i{F +��$0���b�/~�/�J�����'�>�9D����h"���3�@Ũ��wr���?λ ���d�7���+/��EBJ%=�G��D�� M��۩��G��f���X��q����XQ{ws����,�e:�T
vY2 
,�:�R@��)U��C���Ǽ����UZ�ЕɽY8'�:X. �F�^���=���^����=���X��0W�aW .Yj�&M_�w�;�l�ː\��)!L�������<��Cń�w	Mf��m�f�:f�AP��.���D-`��e�P����.�j��5Z�H�W-i�0��
�U>�Ӷ�5�����D�f�{�qV޵ΰ�Lx�$b�?����:����M4TY��t�Dĩ�$U3gP��9�N��8=�m�ۦ}�j���{i��mO�@y��պr�0�7j����+����+�.�ѻ=��L��@�<���t~s�̈��F��(9-�'���J�O�.-È�F�X���.cY����f�1պ�N�wHMӎ�z�g���(
�-�<��i��\"xs[	�Yt��A!��e�%1�9�e�����ɪ}�hn�D�X�����)I�9�"bk�tY�A�#���/�9+C�Qb�,�*�I~�5�_|�kvk�޺�W@	�Mk&�:>�9_�$�M����LD����L�����n����}�y�4����1��5;�Ұ�S�4;
R��f��O6�'Ҵy_o�Be�Z4 
n�^9����!%�5Ho04t� P��蕁�׾s8垦jpP��]���^�������*�'�ڔ�7�9�=��n���Y+>A��/�f�G�p��̄����ϕ�В�m����yM�R_鹘���Y~�	'Ȥ��_�I�[4c`	� �hZ��ݱ�Pw6��q8�)pG���$�77ЇO7���k�Ly��lA��6߈"+,YP��y�0+'��o�xsd(�'Y�Z����:?>z�\c/ԗ�_��=�0���<����
� �bv�mU 8�\A��y����M����>v �,��70�M�~���?��Q�����o�EA�bԙ3�RE1�ˠ�I�V&��C��E~��>t;�{�oU���y��LX[��6}Vj�/v��XC$#M�̄)��Յ{/��`��B���%M�g=76Ω%����e
֎)�eo�Y���@�`�U�<1	�J6s�ʈ����9�*�o6��wm:�w�t��f[�mP���Ʈ���U*��\�Q~^�'��w9�J/�*�Ah����z��\29Y\�2?F�l��jW�ә�$I�m�Y�"�N�γ;�=��t�=�R�7	��WN?4\�Cc%��H����L��L�{bn���bi/?H�A݆���GZ7f���Z��u�~�<��A�(ҝ����k+�L�����s�3�R�N�f���/["��uİ��p' @\����okսZ1[Drګ��v�\�X�EUE��~��� �;a0�G�F���,�G��LxO.G��p��Ik� G {�5�s_�L�ynq���)��I� �l�:�X�y!/�՝�$qcU��(73T���)\9� -�ߥ��w���d����Ed�$�w��ٿ
�i�������4�!ͺ���'GI����;��:S��X|���%����U4�Ӻ���Y�
k�����(���=���x����r�Q�;�{̯[��$���5OPԡ�+D��K!~�(���`�B���-EC�
���h�J�#�ݸ&���J�(�?�"��#^�&u�d�j��7�k%��2���oazH�ҵ��
�t,�+�>E��k�<�qY��q����a��Vpqۏ�ɉ���"f�B�Y�er�L(T�.)Ţ�@X���㕚��E�`:���fbe���4�G[�������*S7JO�R`
n^��&�K栘�:'�BM����VN�d8�
W�b��Oe�  
�������%��.Ё��&Qc��Q�)�2����"���]t��J���Z�RN?�@#�axV�h��H%&I�#��{�L<�Q>��l�c���6�k��ГC�.��Y*F��#S���1t�|}j�E�BE�TP|�D����W7Ib�WHC���&g��b�\���d�,yU%�ґ��1��ya���"hM�e6穵�v��V�r��ٿʬW�N����;�M��<?�g������t Ɓ3c���ʲ�9�_��ո��^�B�#��/.�׾�Y�p��L��%��Ø/εpu����<��R���W�[['=�=�6#�����ِOxу�K�1��6����f\>����Dd��D��<�Ev;^|?�zQ��.�ӄ��mc���p�B]H�>$K�`fm	Q^��u�� ���~xy>��D9o����rl�~��o=&x���up:�y� �E2R0�}$ELS��:� U_a�B�����6�𠇹9��~l>�8�@ϲa�h��4�c5����1��{�h��޽3��6v���+�z���ӞUu傄�h����i!@�N/L���n^�K��X=ˉ�ٳU��R^��bʇ>��=��T��p�x#��fGP�e������5�������	?y�4�ᗟv,��o` B��X�yV�LY{c��얮k�ݨ�
$����� mhaXS~K��&������a���^�ͱa^�(V�[��*�Lo �OC-��[S>�Ƹk�R#T�xx�|���֐�͡#oSw�&�F�3.����aOɒ]~�z+iG��B�N3\��'k�g�mx7�_D���0���)����A`.��T�w.��G"ZwV('�6:�M�O�pu���Kby��ǫ��&���u�w\�W�⏋�3vCq��f�/�"x$[¬l�/������ꀉ�'�*���[:�t��;�㌓,���b�I;�����Γ���G!�S��d�������$��I<�gQaV`��Q����{6 ��pdλ�v&8x:��м��i��8&��&IuX�y����"�t'��~�F��ί��I8� ����}�p���k���xTG;oRMT3bQ'۰�~�����3���g����F� �ɧ���%��]Z
�1P\��X�v*8
>$ �hN��k�&�E�௟��!Խ8�j�dk�c|�7�����iu�.u�k�+g@{�����f?�����&��Uko�Y��>�K����(�Q	[��q��� UA:��o\$���7���I.I��t�
�,"��+b��6+����Wl��\�w6�n򧸃`��(�_�}�]J�W �7q�0%C�QN.S���YE?���'M]71I�p��ܞj��4���s��^yQ�F5;^ʵN����Ou�S��d+�Z1�����K�󊠼�;��mm���������O����>�4U������ �g���"\��j�5aő���	��?�nsʭ�H_i������q��*0����H6�Ҙ����^�!�<H0��N���W�1��p���
n��;b&;��e�/����h*�V+�F����d�����&��u�Q�g�~" ǘ>BxR�dP��4��b�*�ן|1~����<�M�J��W����m庆:v��5_����+�r��q��ķ�����.�%�R��-���*F�`v 	�Pܽ�&�y�]v˨�yNץ�M̽¬��8�է*$�����U}w�9�`X\`���dj�����B¦����/�5�Ïu�:�gѰ��]ր�a������+1c2LX��h��-D���u˓S��հB���|��+[?x(s�+>�L�h���'O��B�F���U/����^��0�9Z/���:�w�A�Rao'ס���p E�!<J��g���3x�h
���@(B���?�~���9J�C��+A�smZ B�4OG��QdD��hA�d�\�ߒ���ֲ'
��m�dD5M��Y�2�~�0�B���*G�ݫ�D uh�&`���#�&a=e���-�u�B�Ƙg�f�iǯ���.��@��ǖ2����V>���ßD���P�W��i)��i�7}������#�t�����C�����W'&R��>�/���-��	-���ʮ�tp�������>��(��&ra�!#
�29Ds�Vx'x�p� �v�2��2_�d&��!����كL+xx�M��s�-��	����KR�!�|��5?	�{����ao��t?�@�iU&2 �6/����cD��7r��!�|�3j�~Ք��)�M�M�[��Q"̃�)�I�ŏD�;���;_a�!�q^�;:#.ӄX�������A�͑�a�D޷��)������i֟�>��A�j���c3�����u�n�>_s�l�P����ԚZ���;GJ����%(>LU�^�w�oߴ��Z����j���Ì�q_�:�ؔ�W�צ����cC�a3[0d&]z�?*5."���q�20�/1O�ɤp2��w�P��������O�o�8�c�j��tʳX�S���~�XrN���=�Pjd�|��.��ٷ>>\��2ܭ��q!
&�Ǹ����T Ʌ,>�V���36PJu6�$i���
l������kS#�C�p@�T���w���v�|���/D^9���e�p�PG���	ZQ�;��ik`=τ��H�0]���=2��Ik��D�1���5NP��38Vn��,��Ư g���i��<~�>z�$����Q��ѻ1�UR�s�����R�&����^i�U�d��l�*`��t��|�DӰo$�ы~��[�І�fSGv��e~�CQʜ�Fp�äq|ƒ�۫é<��9Ս���ئ;ߔ�
i� l�M�"�� `���*7ć �Âm�*ZK�
�g��G
��1r�y��r����D!����o�z����F^�����Z= ��$h��)0�j��W��$�*�
䫟�c��S)�P��w	��;.�H��<��l��ԛ��tv}�̷�Κ�#B4k)��l�[�0W�~f�㸭ky�����<j\	%2<�ܝl�̃뚏�a����H(b+9"؝{ ?y"pH���]��=0E���\��1�v=t�u�|4n*��n��)�I��YR��;C��Rͭ���4$"�_h�Po�� ʈjv�e��H,���^7qp���z�a��*���v�]�;��E�T(�I��2$#C�'�B��KL�/��̙�҈��>H73�� á�!���Z[�pk��^��B-�_�f�eF��`��}����9��h�`�BG��q�t"���U[�Ӊ���S����I�b@E��k$��c�P��W�I/O�������B�f|�\×����,`�y�U����
vW�8>�Z��������+?���N��)���Cˏ�g�dS68�_zl��e��,���%q�c@����q�F8�K��j8�ci�v�������mfG��8�@�>��� �jA@!��_1ƼA	����,q�,|̛4b��tS��v�/�m���M�0O�v�Wv��cǊ�P箞Սf�x���L���Z F�u���q�\ye���qi��I"�xy�_���n�vѪm��n�P�����7C��\�)g�<fՋp�0xp%=��Eu���%��dЖ�ѱ��Ns\Ѥ].3��M��`��� >A����êObG�;͆��XŖ]i8{��Z)���ҳ�����|cYZ����ew�w&=<�@�U9���i��Eӛ,P�F	�=�M��4P@�4�4F�3j�,�J�M�d�95~�p3��#Ԅ�'��n��Gj�_��/z�m�U�KQ�z��'�(;\���6Y�=,��4����#V�2Ls;u��}<1L�o��ʨ�E���=��r�1�J�0°�e>���(8�	�U�8��⺬�`_F���A,�~&�TC�
�ҭ�2%��kG�����*]`���Ts�=r��	t̉H�;�SA)8�Z�?Y���Z���:���m;w 3�.H�7μ�gb
�g!��jO�5ש�P��0�_< JEWp�P5ɴ�D���sO���;�Eό����Q5��6��(G�̴󆥪S�3T<͒Vn"��鎿YBa#���\�9Q���A�uu8 �fDH�����R߅̦
yvy:Kq��"V�V�8������j^vQ�>�>��� x�(�̷��R)�hZ�������2��z�HS5�O�� ����7Y�t�%�P�,KVC��ຌ�_�0��!k���U�����G��c@-�.KW���{��籴�1w�:1�nA�(]�D~T�z�Oyk��w�R�S@���6O0^TԠ:b Y�H��S��Z�и�����Q���^F�����nxu}���1�	�q\�6M�2ԿAS7���#UAo������gȗ�~Ar�EJ��!G�����i�c`[�������6�RA��òpvT���VX2��ݏY/�M�1�29��m�85��H^���k)���6�����G�EZT �����<ݿ^���яB��)�X�ux��,8Q�`9OO)��t��� ��O�G�^�O�y7�\=�c|�17��̟�(���D~��{r�������z�;u�4��|$8��қ3��N��/Ł8��a�F1�%��(�������	���6v���k�rB��@n~$��n��ܤ2��x�(����C�M������jQ�q�#�����/o.�IG���;���|)��X<����L�MC�D���L�a�(4V��1H�����r�l��3a�m��N�xJ��/��7�cKK?��jS�����z֝�|�X��Y��	Gy��I�)�8`�	cɾ%Z�~�\x��/$��}73��W�C�r�"�VLqz�#8&���0ACͷ��w�?1�>|��D�9k�f��7W�qc��k�
��EjG���;���A��Eyv#!i�&��R�hvI�1��٫�A��"�Э�I�YZ��Ǎb��7�u4�xN�"��Kɘ+�l!E�V�4��9NeP,�0���S��z��'y�������6�z��=��=����o�}��u�O~�#���#ʂ��Z��:�He�d��SЙ��@1�Q"�mގg\S"���.��H�
��N�>�!I���ܮ�'�U�Y�xu�Wa�K�XZq3.>c�����f\���68-�! ���:�<�W�'�7L��
9��Y��y�n����d]�$�e�3l����c�J���Ju)�o��Tj�8��y����h/`���fb�qggH��+a@����M��ANQ�V���@�Nt����?����J��H����m��"1γ�����ߑi�W*s�����s��ė��Ĝ�,�@�w������h)Q�A��B���TºQ��+�)�����Eۭ���~�ܸ�e�5��M���ڡ�����v���P	�c;��^��"�LR�H������YW��&S��PY���.�goE�^����?�c+v�̀>��d�����#�!�G&�n�H��!��=r��f��{�d4�q}�-� +  6V5�k��bnbx�K7���R*���Vm�?5t��+b#Gd9;��;{�&0^���g��7��Xm�q��#NB#����l� ��뷮�9� �Z� �h���܂F��+�gSd��hQ	��&����h�z��#���VA+�Ψ'y��TB������5��'S�.\����eZe.`=M��8�Z8͟c��sl�s�4
����P �j��E��v������]y�>wb�;��" ��$u��MgPG�	H�e��vG�wc�oj/f�Ԋ���[�ߖzf����<UfuRТl¬ ��9���/�i�DT!�b1��-���X��N��_N��n��k��h��� כ��)�z&c:����D妚["��F�Z�.�]rf�(�C�-{��{����.	���f�����z����}�v���h���C&X0�'�R��AտܥCHzCq�$
e1P
`"�:X��"�J�>�6�u[��"��:	�q��Co��+q��kk �V�5�"o8G���"A3�F)�;�y1��(o������ڭ\�-��#�!�q�&�n?XÕuV}~4��^���G�I��������؛�*�<sjo	��5���	\@�`Lh�u���F>����"V�m@��DN�6������=�aET�.�TJ .���5E�2R�xF����K�s8u��[/�H�	m�C��͢r-��wD�Kcc�T��8-Q����t~N��J��9�5�l���j��$�@����Z�R� �4���p�_�&���9 ����8�]y�o,��R�^j��8�cDc��G�7�+K۪5�2�yDn[�%~I�(��� 	o�Z��6P;*6nZа��X��A��IZ��0�H��O5�e���0N��}�3����'"��Qx6��L�Z��s��|�7Bh}"�[�9蔦M_�y�P�dy���`�f�(�J��^��v ����mT� V7�$�d1�����~���E�mJ!��v�5�k��zy��ۨ?�C	����B�{��Rp<L�?�44����k:��H	�<K�
��:�R�e����9y_�4��AV_�V��d���-f�H��Aa�bV���Te {�t}Zt��'�3�[���ѧ��ɍW6��ϖ�,5��v� �F)-�4����0��p�L�O�1{*�o(�<�~�p�<G�TuKG���?2S�$R�q7��V�_b�W�V�����Y+�1�����p#���`I�ʬ�b�,����#ك�E���O�S��7����
zy�%Ӊ�{A�>ic�0ʿ}�W��@�z쮗ȳɈ�E�XD��^2���������Č����A���J��{*��ө�hۮ��W� V2��2��9�ͦJ1
��&t �\j�Pg�ƨ`X|�O��Uǵ8�����M��qan�N�_t%M�l�%���a>�멢�ѱ!l�X���K�!��hH����g�$̎��,#�g�k^w���D[�������?�Џ
.ɻWvD�L�rp�������`h�-������d��Oh��2b���QҖC=��e	���W�̻L�櫪�xV���O�߉�R���	^�����/�����~�����J��9��K0���+�^"u���9�j!�c';-��{� ���ѧ��pB�nT#�1��x�l��eO!���s�qIyS� ���sP�PMoo%i��[ocd> �zoM���;G��/�gR,�c�:}H�$�D��v���챞K��-���+Y�������?�����g6:���X�\A������.�|U�s^F��}��y�E���:v�U����3������t��0H'�� _��P@9R�Fފ*$Q��
B�y�$,��C5�
�G���'�վ�.�2��6l��\��������ļ�V��!�R�����ne?󹒌������**r[�$ ao!��3�A��hJm���B	�Ħ]�df�I�zb�����:K�es�~(��S��������Q�k%���^�a���ۧ���ӱ�b���M�ıG�횡ҥ����УK��h�
#M[k���5�K�4��n�,�"�ؕ�A ��?��� e	��~�V������U�ƿ�p캰u�������E�}��>��5'�fϫ���h:�f4:�.�-���F34:.y��p�_1�ߣ|���������3�<�BQ�Uw� �*��p�|�HU��� %���h�8�a-�Kb'�<d4�m���]m({�y�]�lf�[.\�%�V����/�ar����'���H�C˳��ۀ{���5�'� )l�<`���n-ݣ.���#"�ʹ��
F���'?�4:h��Hl��骁��М��Z����ѿ��׬�^�uX����D�W��\����h�)�-���ouD7e/�5���B��a4�a����r#OzJ�����-vo�p����R�k(����a��R����(+�e���ӿ�9���:,G
�.�m ���lg�]�|�l����˃�Q�b�J�
�Iv�}�|���s6H'DZ��a_�ؾm� ^ۼ��?x����&�����_�����
�A����}�1�ښJ^U���K
���?��ێ��%�.~-�������.��ϐ��y�\�DX�?�
���ᝋ�Yn�����L%�Xt�SB�\��H�
BƂ�����|��C�����q)�����!X���9 �)������%K t�-���R;"� v�Ԏ��)�S"��<O���}~H0�\��Hx\
���#�R��]-A�@Ԏ�kpIX:o������)'I3`'�mp~2������?挞���{��=��y�{%.���,@8.���/�O9��VTf M�!p��Hj�}�X�|�����-'\�͆�Cz�^{]!Kx%��ע�+�D;;�{��XLW��U?`1dz�W����@�o��_�W�x����&>�˿^R�dK��d�7v�'"^y��n)sSMԂ�b���b�J��}����_Z!���x}Q�͏'��b�[N���O9�i�c�
���ڍ���r{��U����%T9ȥ�I��e1�����8�*<�rB�SO5ul���c����fl�(���4H��$bȩ2*c�Vŕ0��E�'\[>����.�I�a[.^�.���HpnEu��3���N������x��W�t� �I��o-YRY��Yc?�苠)!OOo��Eb)�j
®Η��Se����,�W�i�p���;�����T#�&����>J?o?0#��w������h�F�H{��Y6$w�m���������<]?э��vq�������J_[5'���Ǔ)bN;�-Hp_�����L���ͅ�iv�n/k�A란��)-����P�Y;_F��@ռ�{��0�ut@]nE?�X��⟦[��f��l~L,mέ`&��-^�Ѣm��A�>��lP� m�cW���:����e�Y>�%9i������\;m/u�Tg�Q��Bz
���h.�CK�����,X��T�Fs�!t���%�@���~���`���)��S��1+/����b���>��#BbI`��[��E�G�WJ]�(bi��+���D�۶{1��l��ʸ����E��#�8��t#C�Qu�p���V�?/-��e��zj���~cQ�F���8����2w���O�ϵ�y�|6�s'�!9^�{�c`���YK}P�����z�ց����j�<��X�|_��T4:-�qȸ�?A�k�����b2�p{���	��E�!@�
��B�&A�o6�a��2���T����B����T����meb�*���4�)D�l�_ĨIڐ�]�M�V��"Z�#4�*^�RE��?�Ǡ�B��_�o������\-|�PE$ޟ�I���2�%#���>94��HȹYx�\V���g{|��F1�R�%u�eќ"�X�v%���N�{4��<ސ�`Pf�T���Ƨ*2���کi;�Gt�q*��
��1<����I��Q�q��[Cߞ
�ٺI������3�(x��SS�������� h��Fi`}?�4F̈��D�����O�'�2v��Ǉ�+������BK c�K�U^�ߠ��E'X�2,d��<�@��.>������ ����J�a�Ո�c?)"S�K�|�h�K��y#����<���n=�7��sK޻1��+~�
�@�1�T���;���db��A�d*�P�P.�X.mP�d	d ��A�n�-6^=��W:Y5����t7�����a��$�8��Eص�ta�G�Z��b�/fPP���Kp.�0Q��GsV���&&XA`2I��`)�H�"G0�"��w=]��l�'���d�Ij�2;�7�T�E(�n���U{	�`��6Xy�G��w":�W� �S�Z4�75X�FWM\~�S=D-y��ʬ�
�uo+���z�"������b[k��oԕ%�A��������(M3��&���?x��������nD/8��=޿��8
�r���wg[�u���T8'���|��C�Gi5��mL�q���d-.=I����D	�&�ܚ�(L����b���R�eܮ�' [^���IТS����#�8�,����bEI��(���m����(�Lh79Ε�h��RVq�C��r?�R�MI�m����I�7�Ħ�k���Ÿ���ռiy��DP?�0�` ��>_vе�2�j�^�țL����*H��������.�s m�:~�!�N�N�e8�`�.-,�[�2�q����1Pw����� ��y���ߝ�L�i='s�~k~L畗��XA�Nw���V]��0��Zej	S&���8�ܑ�17_�E��@GM��S��V5 �,2sk�CЎ�y��DA�P��*/Q���W��.6��ܣ�m��IC_1B�',J�~WS�9���v'�6�J S�p��ȫ�Nd�C+�U)�3�0qB.B-,��`y��~��Y�AAfH$1҇�W��X�RU��	6Yw��&���zr\�!��BG ��ɢ�։��aj�vu$��8v�:'q[��y���Ft7�เ��2�*�l��'+�/�0�ԅG�r����J�_$嗨���
�[�?X,��7O�"�it�{�Ϣ������}�0S֔J�8ex�u����3�$c��։ԡ���xD���@�ԽΨ������귫�6�;щ�-�//z}L�]�.h]��k� ,#����� �9Y��P�h�_\yD��x�HC!��q?5r�-�Vc\¼���uf,��acY(A��y�K:u����˻P�]����!�S]��^=Ѯ�ufđ�o�� �K\��gӜ��c�M��Lto�O��M��m�g�'�*IZ_0���LS-��sT0+Ye<��$��یC'e��?��k
�l�ٴ�!�Hlq�*�j�L#3i�(y�3��X�E��`�s'h�b�Ll.=��2� ړ�ЦwqN  �_�U��C��菱#Wi
	�ɹ�X�hlFH"���a� ]��Z��2�D�5_! U)��AI^�<=��_棓t:n��(���
X:��GM>�wD{]wv�s)���6,v�	[W�O~�;L�wk��wݮ�*��+�i+�@�}��_��#�w� >�H��K�zN�R[2BO%tH�w) �L�Y2��Q��_x�8ˑ��8H��q�E܀��w���#H}��_���o-��B5=�'�'W���`���u1�T!1ߞR^�8��\�Z���Z��(�?�dS�]տ)��L����"�f���UYp3����VЈ9T3���dhv|��{M��g;�D��Hx�ե���8�>����p2���EU�n��B/��t�Aۑap94�`UL��F���Ru�0�T��}���Y��X����j^p4&۰ߡ3��B����WO".D���)<C*}$��9�%r`�z�t(7�14�PƏؒ���X��i�K���g��3y�sGv}��Hw��\��v�@�
H��ѧ Z~���_�Z|4�Hv-#!�#��D��ħsQ���A�}�����Yt������d>��9}���r�0�:d�r9$�R�/j����.ݚ���#�E����^O�-�,�����=�����Q*�t��������!#g�-��&��C|�TX�4���:��w9�A�5�7�a�-���3%��u��	�'y�z��Jk�:c�Qˁ�>e��tQBq،����(��[�
� ��H9�%��<���04�lM[-}E<��W�vd���Aq����kym�`W�vFO���;�~�k'g�Oi.�칦�*��¡�SA~:R톧E��$��HԶ�]�y�t`��g,`d��\�z\�*G�3
}���dQ�_d�\v�D�G���'_�c�n���Nq3^X�PYrJ3���#�h$�����!� �͟��(ST7�@�?�Ϸ9�F����#��.ž�ؿ6I��y�T�w�[EDa��iU�E�4�s���km�h���I0��:��ѽa�ݗ��9W�C��c� !�5P��I�����D~s��F>��$��.m*�Ǟ�+�-���������b�,�Q&5�n�|:�V�1;��ĵ��Se���a��QI�_�|����7�D{̚��GI����R���S¯93*�����Z�sul�w�Y��\��(!2�:�=��'�XV�Yn�$�~�U�
�I�z����쀧�a�_�lE��+�ЙpsN	y�y^W��9�
i�>�\���43r�*�M{�F-p��]ooĝ♰֞�.D���}8�E�9v3��7�;�A�&4��@�� a��a���e$�'�Fyk~��Ӣ��8��Wf�7V��X����-��Ҹ���@���G��E�=����ڋ5Q}3Y�]Swԑք��0E��i�D�c��ߑ��V��E�,�wy�N��$�d<:ey=�%�Eq����`S�lq'��:��SKs�޺!-�x�M{��D1&Jϕ'�ζ�,����KD���R�q�"}������E���+�ɡ�q?L�ۺ'�"1�"����~$X����E�?u�R~T6d\/��$9�͵��V5O��,�㬯򲺿�*��nvȣ�Q�3��Lؕ��c����t�z�1n�>@��ջ�P�y6����|��Tjj�N�A�����
��f��'�y6ڳ �)��Ɵ�(-��Cs5����ƫD��t�zo�">)B@���0��HI���o���(j�Cͻ�p���N�ɔi���S�& �d�wst�}�3/����H�&�4@`\�el����c����ĜO���zv9ë9��VX�lU��2.8�h�4G��=����%�4�r�%։�Z0�"�ڭ��i�A��z���>�\��܂�g�~�����$8u�g��Z~�������9W5��IGt{�.����(���A>&9�~ҥ�f�����})�hN%�ɟ#"9Um^6����i�����B��z�X^�m{I&ڟ�����W��pv ��Ca�m��yz��(��ֶ��Q�
[��� I@J�B�����w����b�����>	��1Y�[9���i�R7�q�yf*m���J ,{�%�S����B�����E��~�k�M��sm=�C�»���wT�q�R�����[XK7ڮ������"�����2ϕ��1���G5<5anX�R(["�I�ׁBw쬇��'���ȩ�,ֽ5ءYԺ��[�_�)`�ݬG�v��'��7*���P�?̤ݽ�B.�6˘(yzF)��2ͩn�n���(H2J��S$�S������' ����w��3�"LI���*��OM�t� ��F�ݵ~)�$}ȥ3<�۰����m>j&��aI����Ġ���Z��3��8*c�w�j1kn�I�H�;Fԡ�*c����K�/H2��x��ߦ�`QxL<L�cZ�����˼�T���a� Hw ��^����\�	,�-?ϝL!f�� 	��,���O�sPuq8,QyH�H��V��c1z+a�Wƈ���$�x0S��ϱ2;
^��\�Jf�`'X=3��cS׎�Uou���
XJ��1�Do o���)�����`#3�j)���au� k��m�@���vt*=6�Ok;H�z�6������6��Bs���H9E���L�6�l���V$ſ�QO���l��Fq��^�5�P�V[V�r���(�[��e@��=5��T%�GP�蘎�u�0�b�a%��n�� !'<�@N-V�� ���g2_�1����r�+���D%���7F:����ח>���W�+��U"�7��lq?"����?�����Ii��9����2�t+���,y��4�2GVoC��3J�g�������z�v�w@n�4:�X��+Гr��qE�@DK�O>>rk�cZO�=8�X���l�P����Ҫ��Wdڸt[M$7V������W�H~5�v�� �P��BAQ�yXe��`�<��ܪ�tķ����\!�a`.����������|p�|�!V˾���o8�9q���2�=�z�%�j�T?`�G��
8�=�^zz�G�ӟVx����p�y��}-IR�e�S��#H�>oƏ1K�~�����R	-��$qÎ:$?����Xo���&��v��o���?x7Y3ʫ��8���w��ӯbY#����f&�E�����9	�0{�b!�@�~ԇn�^��u��8"��տD�E/d������z:�Ӄ�y�{�� |�d�(��Q�)�'u���Q���G��%����A��D�2��>����yi�0�ʞ8K�h[����\1(39XJ*B���9쓢�J��U�xM���Hy|]�<���x�ਸ%ͦj
{[9]��|��0"���&\9���q�g�^�ej��������}�����-��=i�D ��^�G���Cx+��dGk���r������0�(mjZv���
�ץ�2S�J�iT��� �ߌm�f-���e��.<����(�"9'3�� (�K�A�����R�g���	H�b��T��F�*\�ٚ�t��_��)�F$�*�`���C�	�vנ��oMz�lS������v\	MV Hv���]�:!"��\�� �s���{eEO��f��8�0�30l�n0G�����U�Z���5�{�7�W�@Ni/�cj?Xw����r�$bɕe���D_�ke�q�J��;S�.��+��"|8ɑ*�1�[��n��ѓ�P��;���?� �KPZ�ik�9+;p�#���;�_h�^�_1lὤ�_ze�Σ�d0�6nMnz�A���j��UT���{<-�f�[����k	���_�QM�_}$��U�m̻��Ed�v�ɻXfvDkK�E��cZp�\����5�li&�ð�K���LE��ڔ���-��ݲu����j�fT��t��ߴ�����x"}1�%_a�#nC��l�:�\6G�0��Y��ĉ�1V^;��q��1"��6��bE�����n�{�P�J	,����El���+��p#+�f�����rz �w�)Onv6�x�� � G�*��@ m]�=+g^:i�d#���IZ���USvA��M&`x#�P�G� ΖK��,��_�{a�����t��G��Ik{����߾
s^c*b�d'y����YR0ۜDjZ�DwM���ß���_pvI�"R���q���w`˵R��l@���k�?���5;��k�����S���2�7��oUxN�;d���Щ���&7�U$��L�3Wy�&�r�b� k������"1����g��HZ�d6% ,��3��֋���HR��
4�ey�9�V���b��]O�a��W�e�#�C�f�m�M��]Fj��W �y5���/S�����ԠlH������Y��C�G׾������;�b	��(ݞ�\�x�p �kyyLVj�	��u# �<7�g���4�)��!�s���;7}7����%��Nx�o/�=-�©H.Fm�{�+}��_KGF|�E:#xi��l�x�&�5B�k��������6TWy�'&?�>�b!|����D3�]<�xҸ��MA\',e�|	�F��f�t
t!�,�j��3E�+�D��'oJH�����4� ��S�VSd§�_m{�5d�Ι�k-��3����2�>�`�q�� d�I����Cv�Q5~���I귦OH��=~u�0.�_ˊ�6�|�ҢEc�����Q��#n��Vkg�a3Zz��"E��gY5�f#��@N>�*p�׉'CL�}����F��,�%0�X�787ki$�_���g�`���(ey�}���psи��9�;vMd���^�-���p����TOI�b:����T�3���Sی9M
gү_���#é��Ǌ�q"��ƹ}m���Ϫ�E2�hmEU
���<jMP��9��ח�/_�Ŕ��q��Eꖳ�S���)���K]̽7��bbt�{�!Ĳ��������£F��O~$ ��l��� �v��Ej��Ѷ g��D��.6��&��6U�ؕ���h)w�H3�2ww,�a��:�E��<���oܣ_-�H�o����l�4�@J�����wK7�G��XI���e3�H��={�� RS4o�ɽA������@.�^T!��3vh�-�Fr�<<�{n�"�F���T�U$�`�
�O P�a�xx�e_�(�y#�_W������O���p�z��>Z;^DWr�q��U��E��KW6�]ub��SE����cR�!g�<Ȋ�>\�}K��!+@���3��Ul�rcO���(ZϹU�7H��iL�(�0�a��h�{;�N֦���)�O�77����/������A���KQ�}�M�	J�\-j�T�M��>�.D\�bW�fda ���M��ꀖ�~Ҝ��\}�O�"r�D��핣]�
��x.�md���9��C� O	�{QQ��~M.8\-')���jI�ʦ�I�v�ܟ�T�sB,��	�:WKS]0k�n������B�Ї��z..�D����h�.���t��ѐ!.�Cl��L4��k�A]�I��4~S]�á�*�Z��6��	F� ����ow�%ln�f\���h��D�X�&� ��8�|K�� �8\�7�࿪��X�����?'%��(�Z
����K(8��¤p���D����YX����O�zg��bF��՟�}^@px5�p�!|�q'��vo���F�[�k(�Zr �=(���!,�d��U�ӥ��*���G����'�TPR|��#���ZySA�d�ͻ���\Sf��eIh��-�t��x̌s����˯�Ʊ��)ѫ�Hϩ~K�^�_X/mRM�.A�ɤf�5��o7s�M�ea��l��"��b��N�I�%x�0л���$ �q�O2cz��>�z͂$�`.@�W��i��Gh����sQ�zGe'�2R}�dL5���y�>�	�pH�|��ڦؼ�"�/:AHX�Q�ni�4�@��S�m�Ɯ�6>7�S��{̵���{��dю#�zW�k�b�ٜ�}� z/şb�o�b'ĚR���b����ɣ5��4��I��p'�h�����L�j�un��S�,$�6��̳wO|{�
�r����T�Ξ0�0u��D��LM�V�>?-�]i��+u��Pқ�sV��(�|BJ��MyY�z�Y2u}���S
]���Ju��a����3X�[��d�J���Je'��U��f�_:�W0(�Zh���������z�5H�4�M]� XE��M?o���`ȫ��S����#�*�b����sZ���LB�hh�~v�H$=�P����7g��~7�+=!��Ou)���&�X��i��Up�I���񝷻��j�{v� ���ݟ5r�O�ѭ����e=։P�<"���,K«^���9��ǰׇ�7W�
�&��>���<��
��Bׁ�XDr[�9�l���̗���<YC����'O�.U�hu&�SդM ���GW@Eöqm����h�숵��މ&�$��Ѭ������.��io��n[ �e���h���'_�P�I���D���<��\�cґĆ�%YX{Fk��;l�VL��8ix�R50g���&����tO�K@��S'�; ��*��O���7���@4��h���R��E��f�V�kS~����ҭ�чFEʺ���j*D�pX�V���E�F��*O �i��� �p��v�{?+s�#��:\�q�����v���`H6^�L!�_�Nb�4|V�tS�8�aC���s?[�0tI��ѧ(������x��#�2�$K�m;��}�B�e^�Z���O]VΤS�� �b��`$6�Cu��Hk���h)6�)s�Q����b<�\z�l���	�a�xB B.kԺ`��\/���|B��_b�c���Ah�*���2�������f�gsZ`���w*���<��wd��v�ҹ^p�S���t>h1�����rz�[���;��{�2�E�j���bu� ��A-��G�Y�~k8���:�l�+���Fg�_As? =��
N~R�$S��\��Y����3;�;����Z�:��]6 5���S�BJ�Ģ������5vߙo�m���������YE�7�ۿ��E�F�Ģ��Ǒ?��j����:B���XE���̱~`B2a�qK�1��_9�����Ts��������K����g��<\�=Ӝk�g���q���}O^o�`�i	���#����UW"G
^z��GMD�$0-�$����h1M�8�����bMw_���2��`~3|�@�tf�pk�󂔆Bd� $����+$��_�ɶ?���m�~�HSJ!�ܥp	��Hx�`T�"��>g�0���W]AC�gIޘ7��^����%��� ��B�	��л'���{>�����������˾@It $��Ϧ���/�9S���������}��X�5Jw���a���8����`����񛚋4�zh�X&�����~�C��ɵԺp��V�1��ŘDu��&���)5Z�#%g�s����[�Q�˕�CΘT�:3�.4�[�����$�o[�q�H*h-r�>'���杋̬,����� =ܱ|Ӝ'����Y疤܁"*o�}Z�vwss�� 6�Y	��W��u/�~D��gfg��w',�`y�ue�Ԟ�b� -A�	{\�0'�Zý��� \�`��Ǩ��LW��<f��9�F����+wi�!�Z�B�c�J���xIف�/M�fm6�7�YxM�&\�]������4ua���&����m\Gmq�\?�ݥ`"�˵��UM�_�"N�ֿM\�C;�#�������z
����4�� ������%�(1T�����
�2�/�f����f���@Zu&H�(n!E	U0ec���O� �ޢ3QZjن&�b�zM���(E!��HhQ"�.��Wd%�����9�![}㡶S �.˪
3��&�1�.�-��e7���Z��LI�}��g��9d�v#���/(��VW���qm����/�vb�i�eu�8�u�r��6?�EP�ݮ����||b���{,�Jv�5����v�ԝ��i�|Z�I�r<�,�DqǛ`s��Fj����@bl<���h���A��J�ږ�:���\H���^sɆ���t���v�὿��h�X��⁊,�ȌV��]�O�}{��!�sI��=1��e%���7/́�~���8=�Y}�a=�_��&{\�>O���}�܏��΄��gz�UY��egyMog�FB�����=���$�e�G ��jАGD���o-%�u���N��n��Ǒtz�ù߮�^�?��,f�"81b_���:�@Z�E���o$gf՘$���}���S���T)Q�S���<��=�%���ت�4�$F�!m����-�g�T]�ѭy���Xn��'��=��x�q]�a�Z�*�<}��Ĺ9�>�ˎJQ�*�Ò$������e��$	�5�Uލ1��y��0��Qs+�X�t9t�Uƌ�qtO!ʠ ��a��S�����0��LdV C)ǿ;|��Xޤ���vC-���E^=�Q��A�ٜ��*T�O�j�y�J����-���'k�ئE���_&��D�3������)_���V��d�����oC�&I4��=6[�ua�U����h�&��J�V�(���LDL�a��z�!��Ձ�q����Y�RP��s�����vJ�\1���P���X�� kr���<.~+h.��0�\8��X�Q\7q*��O02�$�sQO�]X�3��[�-RH�(��.o��/���nŜ���ccdtL���#H��̜�m�A��(�&�x�o�6�#nƧ2R�IB�^��:���Z�5�֓%�a0�[''�D��i�q�Z��F�!�q)�u0���ci}XeR�*�hu��h�Y+w�#=�U��MْCW�o���0}*�9��#���473�h��~m���i9}����[5L<���V�Z���߯wϯ���'L[S>��6�v�/P����Ǵ��>�Q��H�+����H&�5=�(�9��[�ٯ8�n�U����kP@g��,79J���_�����%ۂ_L�R�x@��I���� Ɛ%v���}uGB�_UeH�F��	��g��o�9Њ���o��W]�^v�/���L�?�d��}��fp�R��-���٪��@�J@E������P�]S��/��ᯱi� �vy��!�Dt�K���܇� J.��f��!X�ưw0���L�C�3��H���m09s-��K��h�C0���c�*&H�wR�wv|{S��P�Th{Fw�n�ܪ�#H(�"�gCK`�׈G�����p�4���֭;�߱��w�l�QWN����Dހ��Ƶ��d#��Ӻ��_nj�G�]b�b"��	 �S�}�p4-��i����_X �ż�|Z�Ϻ���އلl��t7�0t��k�L�9����f�I�s{!#RT��Tg4Û���&�S���u(�XL��)��*�y��>�"	>��WY���'ޢ�*�DaBJI�g��Ac& ���������г-��Yc�ƾ�10���b����20�y^m#�WK���V	��,a�)��%*s�8|qKs�<���g�Qn��v���_^6����K!�!,w3�u�L1��	��pc6�6�4U��;y@��d�
V��Yҵ����d��X����
 �l��p�����l,��1�|�Y�M��b�_��3A�za��i,~��&O�m��ܸ�&4q��O�Rk�)�>�t�d���1��TCS�tݘ�d��x�WF��5#%�J&h��LN�5nsųn���4����Uk+��Asٸ�l�o�^�����G��O�6�����}�3��0�όߨ�%��<����L��!����G�����]�($\���Pi��B((����U�k0dpifry������~�;�d�[�8�_�Z�a���K����8k�6��	��ڨ���V� ud�t�ִ-̣�VkO+�����k��jM��\���Wކ��)�sA
�5"@��7*��+�*�YNz�Lg��m�
�žU��Le�駓�m���U��vB]�$�����[�S����ݠm��9����.�1��m�;b��1����o�CdDRq �X��:�;�,ȸ(�#�a2�i֏�.=�aG�JR���s��g{���Pw(d�1������D��� �у�~K��ң#'V�%�6! k�Fʼ�d�	�`��{���V5b����Z��*~����z,^ܞw kd)l���y����%pc���3(��Ԉ)3�߇oC�s������w�q%z�M�W?��M�BG�K䧪�X
���w��V���W(~��j�����ĥ����ø�9�[fw{���>��0���*�w��w�[�#Gr�!�g�T��W���3��F�X/g�?7����v�W����O�`�����U���:;�O��[��G9z������'��:�h.%��}������E>�&��S�t@he��1'b�w�� ���X�(�1 %_��m\��[���p�J����e�l�b�%�/B�BN��A��(��^�<X�y���J�r�pT@��ݵ��D�+�@k�QH5�_�́�`"ǜ�P��W}�0�J�Oz4vs�ɫty���K7��j4�;>:3Ro�&ϊV<���j���h��}|&�n%�3��o�k�d�~5Ȥ��4Д�j��KҖuk�7�������IB�B4<0��K[��2�E�4���ߴ����k⃠`�z�}kM��t�&�y.F���C�9��W3���:>#��M=�����ƲH�j��	�9&��� ��$�KM��n�p�~�m<��j�ͳc��3#�6����ɗ,��� ��7kҭ��R�؞�:k�	��璱Gs��O�I�O�B�L�2,?��j�D�����0U?]����� [(���z�e��\�O����k��w2��%Sq SּCU�s���ϣ�� �*dK}F�P�6��ڹ�i�l�|��Gt @TR���9{GH��{�0���͍������Zq����0O���߭tʪ�5�;����#��i)E1Ә��M�ߥ�����"�U��ܡ�]�yM�_A�O���;��}��]�?]a!�u+	솛8�`<�=gr�IM�8ª��nq��L2�?�Y�ğ��I�����^c�x@�3-h��1�܋�g�i��KD�]H/�Ug�W1ŒVpF½q8�`��@�ỲFB*�pO�[Ӕ��j�,��z)˥9���#q��C`��l���=�k��1��r�%����$��oC�V�Vi�����*B��i �"(c�]�l��'s�d�P@�rvUܰ��1Xw���t�E�D3�O�R���_�Y
և���q	T���ы�}�ъ����_����(�����f�l�X��OΖ�{ 3F�%?�&Ryn RR��LH5	!��f�I�&���O�H"'�5b��N���TJS��}wD�����cW���@(ڸ̚b�M\���ѿ�����Yu��ۡ��0��LW������u�On#Q>,h"V0õ�L����@(��}6;)y�'�Z?�F��|^Wq�6�+Ǚ��ŵ��� �^¬2�w�	0[��Q�998�f�N��gc��J������/��,rv�/1}-t��$X��gb ����>��P��Ռ���X1�{O�S��:��>���Lo,�X�?�߶���+�*
�	��h�×W� �T��YI��*O�z���e4Fɹ;�5��Y�M*�S��JI��4 `�狎i�Hǽ�p��Ed?�� Ƕ4D�J:L%�`@(E>i�]����bU�z9�mg{�k�B�03e����\]a<�.���st��A�3oD�?��<#���"�[��x	ѻ�����;.�x�3�Mt����E���	�a�;��YI�I/XJ���PA�g��m��^���V�ze]���3�2.�����c�>Ǳ����m�F�J��:�y3�XS��k|+�o�u暋��}h`��i��IS$��O>m�bm����|�(duVJq0��wy@�m8}����"�@��\�37���Z��I{v��~>K˛I��H�ϏI&�#����I�{|-��C���]���B�Y���*��Քhۀ,R�mp�A�R'�F�����yK�{��a0c��P���Q�:�0t}��^ٱR����t�R���5<{2�䴝M\��L��+���҅j�2���P�8�� L�a�/��1�ܫ�5�����%�|I�X��_,/�F��<���cwڣ;�H��3g4֧�	�ɬySrN�r�$+'���⬷�<���2d��H��2�&��0��Ycf�p����:�]C��m_��;�&�@�q�&w����OƝ�;�3&�u�@��n3>qe��X`��J晹?�1��酒�����D���
��j1�	l���xI`��,��ʐ�bх��W��m'�	g����Yf��$q���ߧݻ+��W�O[��ݮЂ���J�gy�B�x[W�0?E��.�N�ЖD�7v�:�G���`�w�owqgrP�zn@;���˴�����r,D|V�Q�%-���=&�eYf���_V"�_�7����r��qn��qA,n֯%Ln���e�]��8��Z�F�����b@.����Xm���J%��5�r#�H�<_���+k�t	A��]�lCE�ҷ���h�On�[mb��cTuK�X|�?���Х�%L@�e��)�V�Kb���GbbC{�V�X�T�R\J�$3s}�oU|1�d�	H��R���I%��ǩ�Gؑ�8�C`׆a%�����z/�����'׈@lTJ� Xg�6�]���rZ�$&� �a��Cr5s�h�G	�Pe<zY��}�(Z�n [F�?
<�ה�K���J0 9?V}�I،����sN�`N��I��7H�����%�a�B�����c��JEcvZ~��8�b��W���g�e���l)@j�\���<�i2@t8�g
�x��,��,���\�q`�@DXi�vW�����3�.3v��:��6y�	����a������m�����+ʌ�2��<��+�
J��vK�@k�
�/嬟Km �9!��J�~�|U576�����<O#�$��Y�օ�ay�=䄝j�k;�6�e�BI�bt8޸ϖ�^���-\�Kզ�Ԫe~�S�	0�7<۱5UXo����;�U��2�WT,<����h[k�{a��V5�����-��)��3�_������I̻�B����]��Đg�HO���:c[�͕�b@ ��T
�QN��H�J���_.%��� ¾���S7`0���{��u ]y�E����fk�B����^�:��,���?��̗���Ä�bM��I>OV]r�/×,bx]w4	��N.Ï�x�D�a�����䛇`�T�Bc蜶�8��^�48�e�O�j�J֗3��%#k���O&� �Y<%ߝ�Z�h�/�}zf�u��\ڀ�ސ�F�%Bz~F��-5:����$�h�L�n2�{�iιܯj�z�-� ��Yr�A�ҧ ܒ̳V �m����C���n*2�M�o��,��hg9[�g��ɽw��B|��&��ǟz>o'�����(�Kk����!*P���c��	�'f�W@w���%�F!�+�P�ړ��پ��JL\t������P[�+5���(��j ��v��o~J�Fd-ٍiPXe�jp�9�S�h�̋��sK/��M��.:�m�ӢT�����^�G�2�O�T�!�[�D�QW���`��Du�ǪC��@[����(%C�8��f�86D�
��N�͐Z5�^�"�L�� ���H/��%��?���ӧJ(m�y䒋0G��'���B��ݡf��B�v)�:-0�j�/%7BZ2��ا�H@�8�Y/VS�qF���B����]�_��u
��fd�O��s�A"	�@4Ej龲�c��&+Џ�g�Zji(Z�l���`����pY��)��	`y�%N�T�X7��O�C?���pc\�q:���r�cLIm��b����`����Hh��E�qe'�t�*ѡQ9'�x���2�MD����3���U��Չ2�ͦ��hȊ�LG����y����"%띵�l���FX��r��$��֡Y��L�j�[/�$V���|
��3����U.u���S�7����l���(Fw��`����~��w�؀�*vM ���k|Z�FT8[_�{��@[�B�ӕ���^�4�zӼB��2��k�:�Y����I6L�8�<Q)��?�܄ ٜ���,K�2���ه�T��gj���i�;Xh\�d���@|{υo�7}<�%.����뫶0�"�F9�a��y���m��jwKI��o�J��
��r�*~�L>���m3,�#�E!�����rd�!,�1��N[��u1�.��5��U%���3oṈ��q�zY�Nj�2͛g��w��Z"We��W�� �Z�5jZ�-������Gf7ϗ��-yo��@sI-֫XT�KJdDpMji���)u��a]�5�`T����,�K����3�ن�(w��c8�Y�s00�['"�kٷ�^!�'IJ�^�7-�Er/~4���Y����nO�`��Sm�ǀʯ^#y�@��.E�����i�b�	�$]��J�U�W�Z��Bj��)� ��G[L%��2H<��"s'���p�w�c�(W_{J#Z[�5Rʤ֧��Ӑ��
ظ�"����t�t�����.g_��|;�I���n�y�s�9�P1�4��i44p������kr�>��8S���BS}�:�G	���O�t�=4I��3��ՅUi=2��\�ˊnx�f6�R	#���{�:^Yn2���d�&�J����:��C��C�,k���G��m_װ�=�=�6�JU�`�p}�ˡC(�a%�I:��T�����F��� ���.�Z�d�"
���0j��� h�?�C7���ݟ�#���R���c d�\/�L�E��8�)*9��u�{Z: ���7ŔIV��4�5B���d�~׳8�]�tNJ	M�-�����,m]!��uWi&��^�qa8|K���(�rM#�@!N��=>��T�	a��@w�(�#
���}��X�Kưt�kt�q�H+S�hˊ��A�GkT�75̮0�A�C����n��MK���'?��������S��m=
�qK˄�l�����-�lF�����{�e;$�}�;��?o��}+p�qLˑ��ǵ�R��x�70�y���(�b���&�3i?��"9���v���y�� wnF�q���`��^�,.@�B34�."��HXz�Y�f�H{`���fȃHL)ke�z��������V�=��������x��4#s^p8�P9~�{�2����Pv̭�auw�LQ3� ��p���ʲД��y���(#+ٸ��Y�"�pjQ����G�z��cH7hC�xp�O�{Ȓ��B���= �VRQ����ᭌ�E�b�#��x˽E�t��H��o����^�����j
��Fm�����D�4T���U�5_�6���Fb�Ǡ�U6&��|f�O}��O�A� �>�YE�i�Fv�X$��P�Xo�u��J#Q-}%\ݿrH�������^�]�;-I�����#�����&�)c?gkJ�k
R�^^U?��+Z��yf{��4p�]�G�#1���TƢQ�5��.}?�J��Wy��޹Q��	U��a�������Ӕj�����/��fgbE��R�HI`bޫn�>�2:d��E����K'�����o�TG����D��L <�T�j�
�0�:�R?�8�߃�ГC����9hpg�<�as�,�<�N:�f��t��u�x��������L�_eɓ�l�8`��퓋9���դ��R�;E?[z���$�fa<Ѫ�ж-�[����qL�7�4���Y�0*؀ ��o%�K���Y��T`ac�x���ڗK���eP� B����r+"5�BŠ�Gk��V�dd�::~�����6r����T����<�;�,�qV�\�Hg�ݲ�ի�H���/�<��.��e����l��Z���@�h��e�T3��̒=�I����+r�o3)W"7�^���t�����zĆ�ׇMQ�&'k�z)rI�Ly���d�UHQ�b��N.��Uw ��7��O��'³�������.�h`�-j'6�k��*=P�ܬ�;c7�`P-)��Qڹ���-���aN��FW44��,���h��:VZiM��9�(�KT�71�1 �\kR&]0�i�Ƽ�:}AN���Q��
��4�ɗ߉~�{�7ҩ\��K0��/6����7� �^M9�j�+�ž��H�查�9Ö�đ)'i�0��˓�z���i�fi.�/K���ov;�X�Պ+�3��R>��e.�e7��R��H�[b̏Gk����{�s}L��c7����R���e�>�nmvB>9�Z�8yn(��%9'��kT$�<��6�rE�:w�!��4��lQ���`�Kl�#��QL�
���!��A�zw9s�_�<���(������� �>��P��
�#S+
�;��x]q���w��&/���tQ}��w��I�K5�}����"�M�Nvb�F��͸&��1��.ђ����(���b����HX�C�K,����f�z^��Nhu;�r�� A�l��e��(�'K�1��o^���2������,�?�8z��=�Ķ_��U??.�,@K��cH���� M�C����h�F�,~@�p��8�5������n�!�� �^G�׮̇qalR{��R��I�r�&l��uVa�W��ߤ���q��>�0����en`��25AY�&d��]��_�&�:��O��^Y�T����d�mS�*�^АO�S�{�"F�4�Y�m�?�3B��E,�L �}��p�I.?6⪩�����1�EeN���g:�0@�,h���.�@��Zu�A��>�##�o4f̄h���5:����������n��틻	�x,˽�$\.�/�qX<��M����_�6J�\U�Y�:dx7���|��p�����#1���n�;|�fey��m<ծ��&������-"��8��!5su�lH�|�\r��p̉�_8�G�S*t����^n-K�chU�vn ��'��	�gj#Х�|��X��E��M�x����NKES%�}��U)nt9�������.�wi?�/F7����)ѫ�L!e-:ruw�b30\��7������J��lǁ���S���p޾'6������d�1��M�H��j�m����3�����͞����R{*�|�Fv�R�3d�o���	��+�9ݡ��+�?o�ᚒw�K*����J	<���Y�����9~������J��4_�1����gl�����
�������Nq��ޛ@ȩA�|�!�ć2��م�2�	G��	. ��A��u�5�e��35s3�e@��mD���r�����5�[�eZ4��!�\67G��M� 3ӈi�հ�T��RK���c�H��Fk�F]3s�������s������>e�=o�}�-���TX�
hV��'x"�f��M��xmt�F��Zp�3Gggh�_��Hq����zZ\~��H^�t4F�ĸ�F=W�,�
 ����Mt����F�Y%gئ!�{�'s���_0up�ݺWG�\���R�}3�
B��OX��� ���rM����s�N���	�7q�\��pˣ�X�7��u�(�֓�fx.�W���Zy�/+�T�����f3�re�ʭ�q��P�l��b�YяaX4{8�a*{�a���Eސ�z�<nQj�����;��R3�?��|C��u�2�7�K�v/�����۰6�F�5��0�t�TX@���v�֊��.F���Zz�
�f�h����`���\8]ݫ478.��v���F�?�faU��H��u��z�>`5�O�M�\��fr�mA���gT�(� ���+h�b��q�5\� t�H!��([�:����j�G��,���_v����Xb�23��Nl}����Ed�C�wS�I#1��[o�>|�]�g�~�4�
y��󺛬����(A��5w����:<�N��H*<M
�R@\XΒv��X
\��
�d���b3��w���X>m4��L+�
_�,ׄ�X!+J�n>��ь=V�j���24ǁK���
Ӗ�d��g������DW�A%圐�� Ӑ�;�<�������|�k���&��D���?���@0x�Yf�5s}�U�R����1g5�F�O4�b�qp�� pT)������tϣ,8'���j��fN��.���b-p8���^����mq �:$��"�Q�;�d
���_�C��攚J�r��@�L˂�L�,��� �M��>&�l3���8\THP�/�ʻ"�����r��һ�0�?����#�hg3Y�bӪE�����{�<��j��g]���F�4�m	(��l[�|9����o���E�x�ߵmG;\�Y���Xak	C_�N�?��V�߂�B�y\Q��78%�*�+Wpc��vo����ـ����]&�Pt(�+�V�&��H/(��o����DYio�l�J{� ���^
�޺6��;p��1��m0eZ�ɐy�~f�^=�Ǔ稴����ӄ�c$[蝶�S'��@�9%��w����%�+�e&�8ݙ8��n�����Hl�����?�-Q�6p�����_j !�h�]���"�|�>U��c&�gf��D���y���2ձ_�l��ou��@����������ƐH]X�	�+���/�H�Wom���b\�a�%Є�^�+*9�r���x��P$����rU�n������;~�W����2�A��BE����GwD�"P�ц�4i�B�4��~�%�#��q�z�m�R=�͈ t+*o��0�6a�=���0ƿ���#�Т'i���F�u��NIS@�̯���Ի��C�dH�SK/VÛ����~��z�/=���̔���D@�`��L���`�r�����`-��	�Q��C�G8V��מ��&����Vz4�s)I�Gs�XF��p�N����\������yj��~�і�W��;'�ܳ&*]<�>y��+�1�4'�9�c�>�� $�]����I���X���~qR�G�i��&(*���5	H����sLzS7��)~�P��n�	1'U�ኁ�D�4�do�G���R���I�`sK�j ���jTv`i���2�t�ͩ��&Ƨ�l�'�B����*�g��w�H��f]�%f3�������йC���L ҪnU���F���-)�4�i�,T\�3�tb���Ž{�K��� ��2��_��i^5�n�0,���^���c�=Ԭ����-�R�=�� ��/n�܎h+�J��z4��&~!�"�u�����gI �S���i!�輝��ԑsh���J�G�N�|��#_5�0U�1j��=���\�G��K}ES��\��m�J�^��A��;b]o4`�Pi�D$�8�ЎGn?����E� X3���.��@-X��u�<m*�$�I�N��p���HE�k���	��Nd��g�"K,z��w��u<���p���-��#������ˉLhWC��V,���3}V�]���Y��£ν���5϶��Y��j���9�2Q��_۾f1�&#��9G��V9r�V<wq�+������zc0X_����4�xX��'P��ݍ���QiPFx��骳�u/
��G���E����r��b�QpטL��5�yoq��(��+�6 ��ssd�uG���c�E/���@tA��9�A�Y�hY)g�����0l�@Z�h�?<���l٥�	FT���G�¶hw0	#f,�f��_XG�:"}ׄa���c��S`����>Y���̈���tW
�eŬ�+�>~I�k�3l��|���e��߂e~Ț��a�:���r'v>)�S�b����f�	D�H�����ɱ`T�ԝ�󈝡�?%�b���jM���:T�겗-��J�>��+XS����&�St'�!��R�m���B1�b9G�uɦ��K�9���àj�3TF�Y���y��ų<��o�@���wa{$x�ȁxb���1��-P}��NQ���nCjF�����%#Δ'���Mh�1����l�t-T_��S���'C$�a*� aw�q��P B�]|H�0��~����ص �B��?P�j��.�`qb��Ǵ��L��[�Wa�@I�W����oa�W��A��a��˾��o���N�C��Wq�E��PCf�¶�K�O�
L@�Ĭ6*x�Cvg�I��_�U+@V40'�HqT_1�</�bժ*t�� i��t��p����L����Y�.@.�fg"�2�����i��\���0ݹ�i��s��z�8���
���U����^=@�O�	j�+��W���:bL��ݴ���x�Y\��(��CB{�yb�7Mq���ȏ���s�~E�<�{i�l�t��fS�;B�#����I0Y6��@��s��ܖS�Ⱥ^����r��4\������U���@e��4�u/j�w�O|yG�8aj��Ӓ��À	�m�Woo�醺\:�F�
��~����l�T[Fk�Sw;��2/q���������h|͡*礌��멽��-E9ߐ���:У����(E��۫s;��E�8u�ql#�EE�Z��aP�� ��F1��e8��z�T��ͧ8�0埗��c����(n�J�;��5�^���c�@.o��4cs�L-t��]���i�~3��%���]i�jQ�� ٍh���_��d����ѧLf��^E��dP�xP�p�R4gf�b�6�@:c�Ȫ�Q�9�v߱6g�d�\���P9p�x�޿!�c	�����,�P���wC���&RI���c|`�����j�ܮD��� ��~�9����<���t����_.��Hy�渟�ȯ�����&n��]ȒwOь���N�c*��ӽ�Tq�[ ��#����k`���T���ؙe�¼Q=�z�}��C!�!i���c={$|0u�.x]\7�U����%[��8�y1�!�K����2v�)v��߄��>�.�!�U�_�����2��t�'�絃���*�k|��j�\����";A�Ļ	8�v���f,Nm�����M���O�cQ�|a%� �%��:���7g��R�Ⱦ<�ժ����(t~�"������U-�Y)9�)����jœU��"��.px-����V��ޛē|}\��A���*&-�
��P"�G�:�������C��Hj+D%�S��1����0p���� B:����ukVg�C�:��%�����}	��&�g�0�Ds`,ѯ0�Pa����1�pIJ��MFAɷ��<:�F	h8���1@N���^�N�L�s��j��d�J`r���N����33��Ѡ���H���Y��ʟ��QKR@���g^.c8��8��"%F��h�fOaX�w�����vwPf���o��	�~;�l�+�c�����$�����(�y�`Q=�D�L3@_ڴ�,�i�O.b�t�4�آ���.�@\3���8,��}g�Fصy�!�&�h9M���q�t�T�m�����.>�߰oB���v�,�V�8��J:���Թ���nH�Ox�l����Ȏ���Շ;p4� H�R�B�3l����+��E��.�I՜��}��ן��c �%������ƭ�A:��S�j��2'��3!�i��>*�C�Ge��pH�W�x����M o	��\3�t�	m���M"�:�;%������ܺym�N!�2=�E����}���Cv2<Ϲ�� 35�UHok2.0i�dckx�mjB�P�3�SYC�pSI�&��t��V�-LS1�Á$;��7�l����3���!���~���¿vc�1f�
J���X�S���QI��]�O��+�����?�~�&�o(�i�f3`�v���D�X�f��̝t���]��#Z�%z�h�D�� xsʹm����P�G%@@q��,)b�J�^�^!|U9�Eo��VL�,�K�s��X}V�����J�ǂx`�����n԰Ͳ�o��.�<�kG�a���G!�kIj<mH&����Nh�&�g��A!�r[��xj7��j�L�N"=���Q9	T�a����'��@pŠmY���,T�-���ǚT��kMe�Y��M>��,���Fp�g���uP]�2Pu�	^�3�Ȏw���pn�:o�s|:ԧiSX���;D�of���+1�M):j�(��G��Yq�dpۯ�X9K]Y+o�N׉c���/Z�:s�/n�a�
$��?Dt�RP`.���� ��EI�|�;�'v�%�(�U�>��G+�-����܊UF����}�O����/g+�6��_�Ɨ�/h�r��TTz8�pN���Ahy�O��\����u3���0��iTD�Y�sJ�NOA��o�N�
x!^��J���y�o�zs�J����X
*��Pg��{W,&����#c\8@�����(� �P���>��>��iNp���&�r��e\jK��R�c`�O�4+"�{[�!��r}\�s�nyIӽ3��٦���߯s�UN�����v�%�F��׫�f�:"p�"[�E�PEGd�q�9��o��Yx_.��S뚘��o��2
��W�j�k��t�z��vhuxU�_���(��H���
�4M嬁��+=��e	��[_P���?�iq*㟕`k��o��Y��Uu�yE���4K�#d�������hvv��vly���QsR��+�I`f�&!P�����M���1�Gr���d�)��"eAE�y��Hm�
ըﴶ����`��I�~p��a(o��Że����Gpɉra�[(��n,1����s�~܎���h��Gjvnn��Ǽ�r�������w�;Mk�sE��n4�<)�>�.�Ы-�2�����)Ȟ��x�e�������Aj�8m�R����ف���o���!��|0��1�L<�3��
5͉o�F"��fc��]%\^���Ƹ�Q�F�c�6�\Rr<�5J��iAQy��밞�HY�B}{�����	h��WWM`�bAS�`��Z:]�"+�%���c�s��ݠ��<�(�Ŝt��M�d֚�1�fD1�+��-~�
MT ?�O��Ѩ�i^��QVL3}&�/t��	zq�ϣ�1	����(/0"rN�	n�r��#g(�+�o��5���؁}���Լ�D�x��`H\��h��g�2;{O9��Ӛ��S p)O��J-5�C4*[ۊ['��?�,��b���b� tHs�ˠkÿ�P�$rH���������Dc���W��#R�\H�'>�I-xCp�5����^�C����Ό�A=;�Q�\땅�R��;=E)������ʟ+C�o���E�4��v(lB��i�54P&*�|���y�t8t���E�hX�Q�p�k�����_���ʔ�Uy�ي#2?s��2S��5 cK�:�D�k���Þ�A&dF��\�	� y Z�=؎�gr�n����7�P�N�F��؀;�����}ҼȒ 1$��������ycl( �pUޜ���Og�ϧ6MX(��RQEk�F�=��o&����-���K�|N�o������$ �Cg��sT���U̩��Z�(ì�n��Ѕ�b��A����QIctw�����@}?���g��`�*�����cy����������#v.a���!�g�����C��:Y�Q| ��b� ��;S�8e�����ӱ�(�Y��!7.�pޥa"VQ1W��P���$0�����ǥY�x�]ֹ�@�# hBj'I�S��5x�%c|��z��^h&D��?G��m
6g�f!Wi(���-dddmP�:ڿ|-���e5��}`h)��U�Ǹ����qf��;�ZV:��u���>Л-N�^�+?�IbpT�T�p��2h0wu�W�����J|���� X3xD'y}�[�nN��p��Ee��;��:F�A�����'���ר'}=�1�R�4@�Y��|��m�e�ed!����#����uRm�>J�e��"r��"}`�r�q��q����$xE�Q�(�s�Xa�N�����O fb��h�&�4�5�����?SJ����b=y$�걓`@��ft4��܁�E|� gT�ʺ����2bY9��6G��Lc��X��O��+V�
Ǯ��lk]  �eT�9�?ڮ5t}>�����*5��!�i3�L;��X_�=!��t|�Q�14���Hʶ�O��3=0��1.�W��ں|B�g�p����f����SB,)� ��Y��H������ 蘛d/�8��iu��pj~ �%6+%�~6'w��U��Q=�
��4,9����`�`b��}9%V<�@�7��z���)��W��W��"�=�>s�$Y�ă1��a�f��DiQ{d���|�� ���愗�՜#����]�ɧk�vz#WN�D�;%�v@P�"��m���&�:o�����2�������7W�bv��z`��맲�,�z�ĵD�Y52	�����%��}���a��8}i$H��H'!Ó����;�����K�="�%b���� iH�C��}"��Fn��ڏ��fc�aA��J��Cg!�Bӏ�gX^���)�b]��Z�
$���/���$�J�L.7A��}9�H�O0th��/��{��# %,�t�;�?Y���.���K�R�b�P���cp�y�0M�������S(�%W�!B�Ϻw�g/�u�=_{�r�I��;fqJR��u��N�\�N�A�IW�"Wբqc$��E�q%1׬�m��M4��n��/Cz�Y=��O��#q��������q�Yge�l\%3��Ϙ�Ŷ������]*^sՎ�R�Ht��q�ɡQoK�I��2��R�[�!l:��~��v0��G\Q(wxУh��z�v1�XZq�"|0����z�/�'��J�E�	��j�Z�R���rb�,�f�;��AQ�Q���ԕ�j1?C��J�g��@G�iO�I�����q��:�\�\��wjѱ+�15�G,#�~�д�$¥���y��q%�6\���>��hV���HEt/b�x��GQ@��}ޠ!��/�*��k[�\�J3�ػ��o����Z"�("pe�M:�a��{� ��z� �������BL�U�񬊴��Ŧ0V���4�Sw��[-�9�a��r��_<�������7͏��Ln�ރ�y�y�6����{�E4'���ElÀ����>šu�B���|��i��w>��X@��mg�?����]��&Ƭp
,1ds�����K�U��=9o��'p��)�[xT	�%o\���j�r"(F���"N���D,� 
��8�n�a\
?�p�T���vU�?�� �h�:��ꡕ4�7Ή�/B8^�1�76B���64!�d70���iv�1A�Q4���a<ȳ`��Й�����ƙ鲧7+M2e�E���Ȯ�˲���7��z�3l$XP����}Sq|]N�����J���e)�|�������:OϜ	wp ���SK��	%[�db+����E���C`�/),$5�WF77���������PY�㔈���ܥdhHJ�(�xK����y��Gx�Xg?���q��7;��q�(@d�r�7�Dg5}j�������)�V���u{>�����n�εK�ia=�R ��}�H�ʃ<��ގE������rɚ��@�#�~��WԊ_��Q�{?�m����I	I��vB�Q�V�CO���������H��ޓ3�$�Sȴ�` ���~�{�d�r�W�E������J{�:C$h#aMQ�ys��������IY��$T�pf������vdf�qrW��y���v_��BkU,s�]|�A�"��nJ�PqS�d'3���?��0?
�oI���%���ղ��n��?(c�a4ib`,�x���Ju

;����V���P]�zZ���Mqa�_�"����=���*	�ل>�:ȯ��q=�յM!Z�=}�?ǌؖr�-[[�
�Nȃ8k��������.����dr��M��|�B�l#����n^%6Nb��	G�+1'�^Nj���#O�}7I�Z�0�U"Ykb
e=���R��~�lgX������J�f�m��� ۷<����r�$&�P{�S�

�-/U&�s~����~����������|���#���5�4�1�Z��G�ܑD�����?�<X��Kd�wa~��s]��Ө��A���Br��y\Q��0��,F���;�����i��B���ьH]�?j����&G�Z]��{��� 8�4@T���#_:��ߗ��M�F��l���D���7(=����zLt
������_�/{�][�+�'_�X�1�v��7����ou-�)Y��!�H��ɮ��R	��%Yg<�m��E��(V�M2Z�� SG:`fw��5+^OO�4�����~�<���"d�} "�%A|��|$3��5�ާl� ��2RL���\��m���M���tY����p���I��{|�Q�BҦH6	wsr������_Zy9y�|gй�Su����J��Jސ?��B|���}�Q��p�y����V6�F��24K��`
�B,~M���y��:<J[��y��E�68�Ns��b�<R��L x�����e.[s�v;Sz�&J֌���b#�Z3DĔI!����t%���6ீ���%
�v��2Za?��*���i�#�t��b.�Qƹ�u)��l�Q%���3�Y�Ŕ���ӣ���줍�ҽ��(��P��f%��i�.>����:|�9�z�l1��.�=��!@Y�j(baS�@����@�!8���.��Y3�5Z<���_]ކ9	��4CW>�G���dE�8�ߕ^���UÅ,Q��Q��9V*���&�H4��^Ti����a����c)\���;��׊���V���ߴN��kFқ8*����y����;Y
��Q��O��r�d��I�a���S�M��A�u0K������˗Ռ&�uR�T�I�4�w?@�"Tw�]_y�h���q��F�<��F2L53�Of���^\�V��Vqw�� h(jى4�pHl�����4��?!vѯ���v�v����۝��>���D�``�*D9-e_�j����1�^pd��ip�IU`IV����NGM&����;={��W2v!�Yd4�@yhA���Ut�ģ'D_�ߒ�1��]2%�i��nw3}-<c�bc��E�χygr1�Z��	˺�]�ցT�Nz9n9]2�X�!�s��-�'j��̃�J�ߊo��=RSs%�z�5o���pQ����W�n7�̎%�%�K��5c+[�'�!rT�/����eCV��hi�+%g��U����8�_:e��OQ� ����9�ubb������la�*��$w&���z���<(֕G�מ^�N������,R�����,���cy�1=`'���oF�6��Z��n0�C �A��JЦ��8b�O�[ `�D�]�������j�[=�t��7X{C��7�L���M�r�����J�\8�ߖ-V�Y����?9���y���[5U�z!��8p���s�`�x�Ĺ��+L'�ܵ4�6Q��9ch-��ᢍ� �%����� 5Ob��7\��[�T$>��wVΕ}���I� ���a���I5��� �|��$��	�D�Ãt�2`XR܉���'c/o�������6�@Rb�Ƀ�}����#���ֳA~� ФFj]w`h6A#K��0|<˿'ko2G�ݺ������8�R��lJ�p�t�Fx�7�)�,u�պ���M��F�EQmZd�s�7<���fk}�<�!�q 6�b�OcD��Gᩩ��+~D�K��yh>��g�_
*:B�i�������l=.� �?��ݯ�>4�6Ζ��ʉ���j�}6؁�"T>�L���u�A+5�5(���(������b�6n�
�4\�5B��p@A˧�"��oȤ��p��58⽿~�r��6��;��<�]3ANi{��x;#X��3��-�	4f/]U+�� quF�$=�q>��@���r���Pa�� Ӟ��<�osu�mi�4��tm��	���E���4N�ÈCK��!������j}����3�a3�����=
 fD��>{ ��7�l��@ާ!km؛���
@*%��7$  %��d�G�V�9O%|�8��2	m6������ӢX6�l��-rA�(+y��A�!	���QKJ➸�0�� _BQ�+T9��_0\�t�R?t�-.M֗ik.��ާ˚Uu�ޓ���F|�m�u�?a}?��'�'7��¿�A1C�����'5���q�3�^��p�߱����O�LZ<���w`������B��7��"g��E]&�α���v)m�^����������m���p'�=M;w�9B�)��$�[�k��2�À� �?�p��@_�(@V�$���1�r��m����t��*�=�D����5	K��%t-�������Z|o�Fɸ)�Π�3&�a���ܰ0�D�M�jeԧ7/��~_�	��kE��x��$���)�!ޣ�o��QS0d'_A�[��M$nSo�}��!��K+/;d����[Lz�*��!˭�w�;fOM;���.Y�~:��l���!�7;~54���Ϡ ����̽�*I�:�H���&������\hO��c�P���ީ�5�רh�	��4�M�^�W(/�³&z�w@����|�E��_i*�?Ű��%�Rx����4�Ϩ��h	�f�b&��;k±��"}l�^�a^��C>���`�K�MK��<'�k�ӥ�,��`a8Вg͎���<�vm�>��`����Z1L����"�&|Ͳ1.��A�6�D�ܪ"Ϗt�nx$-/��})Í�H��J.o���i����}�Hc-jZ53�NС�	�ők��>e#�R��I�¢���pPϰ�c�e�p�C��U�%Igm{ɺ\�$E� ć�M��Z�C�g�?�S�R'����� l$�@pֳ����w�I�6ӨOq�f'�Վ���4�$�f�|���0g_�>7�>��$�\b�ڡ8���o�Zq*�t<�U�u�3Y�����K
����2#U���.R?��,��}u���;z����@�e��8�nFj��JY�>�[��`7mW�O��Vm8�	���Z���t�!߱E��n�V����X�+�F-�*΁�P�^�'��6s��g�A6=*�OL̇�=�?�L���#�Et� �څ�Ԡ��W*�[a<ɉ[���P-��Ѳ.Iu�C�!e?��
�jdnXGq'�^C�s�^Q~z�J�jqy�+ϙ���v�Ȇ��a�s2ui�I����{�	�D>��lw���%����|��)S�Kʒ��?*H���}�<$k�	�U�h�=��H���A�mI�z�TْH��%�.��U�%��!�.�aJt{���TGXWDo�	��Ip�x!�B�X���%�S�l��9S�u�`��N�F6�5���ћ>����m�>��`X�N�$n�j����/�+�,����6��wo�a���S�����ϼ�k��<���V�+$&���Ksa�#N-锸16��2I�C��.�K�Ai��w���7�>�s%�J:	-��S~��������cC�$D����i�[���0�w�|�r�r9(�b�/������v� b^z�D_q-n���|R��ɂ���OV����X��g�n+����&��LdNG\��JmzG��aO�Z���NM��U�ɵ�8��mۊ
w
��,�F'^KSb&��W��@6�ER��s �����^Dr�-݄�O_��9!cQ�SP :���E��J�'?�/�FE��8'�Q�����2��%tRy1�y:����05�4q����h�!�X���j��$5x�Adw̌�V��|a��H��I)|`�J$���Z���Y�f�`����#�깡 �a̶o� �/���s�`j���v�bi�9��. �����4��W�� �P��9�Xu~6b�ؘ��-�z���k�Nr�?$j��)U��a�R�vǏ-�Td�3 :�B��jɡ�Z1�e{4Q���d�A��/A��f2M+�*�9���_A����/�hϓ�WVG{��_׺v6�WF��8Ob�C8_�%赵g�uL�	��2(b����,��V�HՎԣ��:�/���j��'�!��"�Y)t�V���=��d4��Bׄ�����S�P	��u),;Q6�;��r�Cb���{̭S�-��mFߗ��������@�3��nٿǕ-���`=�Dl4�-7�M� _�3usz��RX�3��1�<�I?�[�A��'��:~��M_\z1#�� ��'���K璦r��;1O씡J�\V����gc0��f��0��鲲��w�>��_ ������[��6��Q�_V��C�M.��,�I��Vv�� �c�g�2�����\8�2^ڐj�5�5��nրZr9/pR�{�vO��x_�U(k��/�Ƕ��N��� ���l ���~Y2��4c�;�������#Dpe���O��jL�!7��uƗ�P�{9n�p��Eչ��F`L�Xr5v�EF��\��ҟ��"��{�?�a�1��p��3׹:����i3��=O���t�jEw�����3t���噀�R$��P	Ei��=���k�,~D$�vd����<+���m)��:��Zm�&ނ�a�"�%g�C�.O��r�����Va�RŖ�f����̃Â��,1����Nذړ*/��I-Ϯ���T�����[1NDk��8�s{h�l+��RV�w��,�S��M�]�.����c��Z�t\�,w��Y��~����Մ� ���47�o�Q}/5K}�����M�O/�zI�iQ�a�%�I���"�/bSR��J�pTVsfc�A��^=D���@ U���q�gp�9��B{')<�6�ӻy��*[۩�"�MB���-���H �G�����2mK ��w�l�������4=ʜ�����%��/E�<>,��eɱEx�N��SLOs���_	OUu�ߦ9�N��|�g�L3�ɍ*D�N��`��1��֤�n�
�>-����MN�uU���x0@��- "{$ע�w*���'�+G�Q������Pρ���|� �;eH��V���yQ�2�z��%u�� E�d�5g �#ˌ��L#��*���2c�3�^��PC�[⺔�@w@b�-x��^����slG���GMFc��@�z���]K/&3r����yz��;��9�x"��l:�Y��,���.���A���%��`�L�N�5�3��?���^c�=��JP��Ao[�Ҏ��b�*��[�)oX9�UJT��;n�y�<A�8�'��#��]�k�u�|�5��Zߨa2ɰ��I�|(�QH�qN��VwArׇ��;1N�cPױ��bp2�	B����-.[��_��l""p��q]�ǹP<�p���Z�ޟ;��}0/ ��r�`\O���.����sk:�>}'<<����� �I�s篦:����r(�����x`�q9���m:����Ee���5�?�qֆ)���M�yFW�6���L�,lq`�6~m�|1��K��{�>�<=ɷOl��Td�����a�IS�#��1@�)��q�}z���c:�"b�ks/�q��n�)�HU���y���dJx$��9X�ҾB$A�%-��l mËS�6���iK�*��̌��c~9���<`����Kx�rb��3$X�@�k#���2�3R�d�V���}����e�!��U��X��_)K��+�eC@��=�:����?����{+`�RY��������<���$�����~|2��\��Pl�e�%��$a�����U���z"_����������{x���J�v������-������0DӅ�g��O��:��<|�v2c�Z?�{͊mMϺ����_��5iWNO�ͫ�j����a=1qc�V���zOZ��>�U�IW��(he2�2�lK��Gc7ۍ|�t"���.�ҁ����q�����I��K>-�w�?2@Mn�pz�F	��+���v�f��`'�����8 ����L���='3����9�73�M{+HĂE0��r2���m�s&4���Of��OÑ�����2;a���G�:c�1WD|�5>尾��p�Ez1��W��w.����JS�h�1��!4L}�	�g�e	����j�z�(��kJ��f�����?#���4.��6ȵ��4 �${����A���%��2;rV�`��%�9![�z/�ʁ=BW'�R���?!wC��Ul,�\�7n��[�W ����x��5�`�θ�,N�^<M+a�M�Ã*�(��Z��CU�9ұ}V]��\�H�ݲ���BA.s�RE���p��>� �}7#+�N��t5FOL'���%cӼt��mg���/��y������c�X0�]o�\��DVG��	[ri���i
���e�Lb�f_��
�<�e4F#g��k��,(8^y�e�x���>��4U뙌�a�3�'��7�m
���J�Vɡ�b�[����sYЈO^�ZGR͚,�MV�~D{0P
2Uv�%���n�S����T��f�R��� j$��88�J�z4$����x���Q��,����@�X� ����K(J�7Y.i�W0�X����g+��ޱ߳,ޕ(��x�b��`��TN7:��@���j����W>�;��X�Ä�r����\;�k8���E|�|o���8���8^W�dحZ|���WQ8޺���M��s���JɃ�%|��^�G�h�Ym�̜���,��m� f�{D4S*g�JD��d�_a��j�2��Ѽ�9�5��߄��Pw��wĊԅU�?���%Vމw�o���!0��ܘI��ˇ;�)�NX�`����G���]Y�C�;���*�P�}�X:%�+��Z\�a�Yإױ��h���gXiv ���[�f��o/�)\�(E���3ޗ��R�m/����b�jn%h�I�v1������|�ɄP�E�iw��o�^#�u��iq�~��J,?�N׊�E�	���HB�\Le�h��]�	�։'`�翮�M�QbwCO���2_f\p����j�qh���^mLe�K��:-�!���Q^ˉ�K��stU�Xj@��k��	�#,��m�N�fx�!Z�I~2�-t���/���"�#��7B�i����.��m�T�ڑ�"Ol:�7��)6j�"�SYU�Y���t8�a�|�=ڎd�O�e-�4X$��5�Zp~jl �c6��[�R ��X+�
��)|���밤�a�#aP�	�D��bF�DX&]#8����h��iW�3S�=��o"��+�_YVJ�w7]1�-�Z�����]I�{I���n�7���yNz�1���b{%�;H�5�F��3�aB:��K�	cZa!�����i�\&�A�@������"�LWc����.��H����Kq�I����$����O_"����J�¦�~���Z��������;�/��~B6����L/���
�TY	gM�h�̝7�������ocR������&������h�hQ}����3g��Ժ������Ǵ\
����e�/X���z��@o�4%�T�2(~���v"K���%|��*np���4�,Ma�������#��v �&e�����RQ�������{~[�@Ѧ�ϣ�V�|_��k)ovn��Or����Ȉ������g��>T1�;�������'D����������W�MKq:��G8�&�+ ��u����v�qپ���tg_̗�GrF���V=�D�G�v?�̛6L�e��JEnu��6Ƃ��{�Ӥy��2�sIy?	_��־�WQ��L��ɚ���'��{�f��iƋi�����s��%7K����^��|��\��_v�L���q��@7�K8\nFFv��ȴ��Gֳ�x;��K�!���Tt[rj��)��@W�¼Y�Ǆ�������ȵEp�~�l��j�.B�A���/n�Ҍ�t\��iA?a+5vyY��VZU49x|�2�+�=k� \��X��� Ӓ>����B+p�6�9�J��c�pA��Ҙ��J3��&e��-����8��-�*��&�Bff]aK����y��|ߛf�vaT��vy��
ː!��W��>�Ct̺~���d�xB�+k�Fǡh�i����Hv89&�G��u�j�ײ�������Nr��ߴ"�
*����������ٞF���RkHli��z�
/f������>�a-��P��>:�̬7�J�Z�i�.&j:"}斴������h�^V�t:��c4�<��:F+�.�:�?Zx�KR��=���E��n���<�		G�( *s�{My�>��Z�sq�P1qOWI^^��`>�`�����MX4�j���;�GFgA����I�*����|�~.�]c��i�4�OO�˙9z��CXև�ɾP	�\��D���+��#��_>��豤wP��Vy�k�����9�E�]����З7��T%�f%X�[�F���)��5ЙҼh&7xD��$Ǣt��>7��7-�\@[:@�?�+����b����o�{���D<Ck��B��Yd�]ۯ�ǌ=p�\��2��qVg�򄱄Ǩ��G�g[�f.$e�+iGG��#`�ç�U��YQ��ڶ�<�����}_^�L��We!��������mմBp�fī
t�9��>G.�l�σ�T$�U�2�� ���b�j��2�S�����92O��j�b�t�\oET�f�SH����_���'y~h�ui-�Ӆ�*���ѶY#��qԾiSOr\�*4���u���.�|����<�G�n�i��*[��Q�?ce*�,��R��P1K=��y0� �3��+!ߍ�����is�Y3K���av1dҰ�e_��Ț�6U)�]�o�?�{�⼑�j�m��y�r/[�"�_R̦�>5��5vT�� #.zJ���h;j#�uƸ�����ns1dn�Q<��t�r.�J�������{%�a4^V@��B�)��UQY.�`��rZs���g
X�ߦ�Y��/iMM�%&v�}�_�B0��-�T��թ\|t�f8rCj/+�!���G�4 ��R:9�3�����CPZ�L�;gڔ�OS���lDI`���R�n�
�N¦���76|�4�;DG��pNy��T==���=�d��U���>��ǽ�0�qZK�;�r�~=�s��Yv��z:Ɋ���^X�%�㩻xp����ՒN����2��YS�i�������n�7�<�i��z�9�,��LHg���.n��d�r4)�z�՗W�� $��Zjv�}�*�Gp��� ��tr�I��:;2Fc Ic�Cvn�2N�ǐj��+%Z����K�����*E�аLM���M6�7�#W����F�o�x@C�bW�KN��@ۢ~J�T�C�ܕ�z����ۖ�S֙H7�X�������B����[�B�h��=��|�m]Yk&Wm�ln����@^��N�����*��p�7�����+�g�$���e��G���tf����	�c��l���=���a��zu�K ��ukH�����定� V��m]|�Z�heP.�?��@��VL�Vr�_!v��Ӏ����x%h+��J��	Qoa��!��<��	S��p^�bm�{'|[�Y������Y�)�v�G�[H7O�{��0���9�ڥ�ݥi@nLk�BG��Dȩ�0������ ]v���v�z��W�1'M\)�M��H{?��H2"�pʯ5T		���G�yl�(������q����G��G~��R��m�OCe;� 6��3�F_�;�1,%��s	}m�>�C{��98o���8�0r~l��ď������!�Ѫ$�$ulL��>��ĳaS���҂���'�̃�CSd/P�N8"&�.`I�J7�y�?��)aF�z*�3�冀�W��.��所 ����aH�8^vf��V؟
NI�]i_��f؁��@;r�I�C���D��7��7�ѥhW
�)c��ʂ?P�#����V&�����7�]�-���?�[�u�gK'JN�R��r��M�wC���7�}@��y�" H|#y�D���^
�Q��I�ӈY!��MQ=�����S�?���e2/�|Wپֳv�n�!K軳��WL$6� ���i��֠���$��I>���/
�6I��QϏO�<��L��kg48isK�wU@���3"�+���(�c�g�c\���?&n�j�\gSM�X��2k9�-�u��W�{?��Sb��[��bp��7�lY�����݀���<f���R�@������@�����z��_�ny;g�!m_Us���/�cN��2|��Qjލ�1$9%
�:�nR�v��|fn!U�~\��`�Κ3E
RԠ-�x�ih�@H|��la��퍪8����>Q6:4�br�q<4�_�qUػ��{��ع�d'�R�BK�jw��9���n���R�<?,�f�����2���hϤ�T2;�
�lRq2���u��YC?����`W�R�wN<��N�@���^�� ?�@-.�؛>l�L0S���+n`�T]>�Dx����Q|����`J��պ��wx�d�ڮ|&��L`W�lDV0��]�}�&%�g0�>�~��L���"ÿ^u��c�X����n�f�X���6ƻ���� ��?r���9��j���FX�s���;�R��:  X55%K
Կ���>=���Ɯ:�i"}�p�Ë�y!a&�S�p��V}#H��"9b�S)��L���LB" �	Ki|#}��,���Q�<��c��o\T�S�F�����M+*A4<މ��ɞj��Z��%�R�J\��S#u��	}������:K�]i�{��v�����a�Y�iT�[���x�챍��t�H�xY�e�,��n�J�:#�tÆ_�I�R凷��#V��?���!��Pd&�Z�]I~�@�Gw�z��?,䆮D��G����O�|��������Y�=W[�>ЫB5i;F�H�Z�A�3+�O�e�ɳ��*���m���=���f�Fyە��x���p)�̍�q�2���b��*X.Q�/ֹ�xF�GS��Ǭ��܊n�T�b������q'V����J����E;[�U<���U�c��{��F�DWv�p"8�@���9�O3E�!�Gk�7��X�ĺ`B�(T�mE��YB���	�B��,�ݠ 7����vNjx��_cZ����g	� >�jTZ��3s4��!�u�	���p};��+�[�~'�cPF�T�|į�_>;����J�^����k�Y!��J�|x��D,�KrR`���{�P�+���w�}W����V�1(yE��BLc�P��Oqy����~��՚�7�Z)m��;�]�_����-ȷA�L����Λ՜��s
bl��.�[��~Խ��G�Cv�p��,1^��j>�	%kU�bx)���)~w�Wb�'޼�ے��eM��@6���Eu��iÀX�����cr��9W��	-�W3�������o~��QH�*PS�|Rb��]��5��a�_��A���a럪@�L�2_Y�)��Z+�<[P*^�R�U��FMUzLp��xcOs�!�f����9��5�����=us����g],�|=Nc?U�N��������=\�Iv�=�aY�".��N�ѽ_V����W��� קPP��
���A0U���k��Ҧ��F-�	pWlT��־�C{y�_�=�
���u�[�ql�iy����!�זI� G��k��g�9^�(��s�t0Ψ|"��ڔy��o�Ǻ�1��r��g�;�&�J^ǐ����2K�_Za�M���"�M�����i�-��Wc�����p���1��JD����jTF�%u5À9r��[�=U6�\VA�Wq���0jZz��/�#��)���E�+��K�&�Tf�����P���+�=a�xܸ�V1�?�A֑^��y��^�AM��7p��8��i^ބ��1.ujX\P(�O�89e�[��6��fפz[|5�K8qXa)��N&��W����P5�?��kb��s� W��|��o�Uo��Dv�7��g�����8ա��7��/���@���$ߦ�Z�U|�Ж�sR���/�3�^g%/r#+"��SL�V�}�o�ȅ��܂�tS1��y�������W7?bk�����*��_1�C�3�ZI�FؗsX^'�I�!��EY��DwZ�
�(��k��P�ُ޶���Hp��^qL�=�к��X�"�Xy8�'A��+ԟhn�䜤�����(�ȯm^tahZ�h��BRxTHڵ��2֥���nH�!��Us��!lZA��������s~���� .�Mt�f�#���P|}�P��/���}�1�R�]�c�f�}DCl����^gC�H,y��dX�p�1�5v�־���DF�t��0��E,�m��KUI �Is0OT|�@��-a?v�ѩ�y��>8�p���������!^��[`�Eg�:���k�z�JLj+,4]��]#�����Sy�=e��2�5X�_,�O�5��3��Q��XWH֪����W
H�ړ�Zk3 ���A
���:�iwpH����TQP����C��Ͱ�\�+~Zw-j�z�>���2��g!Z�%1���T��S,��(iՑK�]��:��t=�Q7���V�K�о2�
x1�!xp
����:gR�od�J�t�6 �%���E��e���XOn�*Ǔ��l��@��ul�iw��^5��������7���3.���:�[w��Qtn
ܴ񭖣���D���{�&1�S����fSF��!%k���)j|D���7�_٨j{Á$(���BK�QL"��\��7\��U֢�yT�+3���@;�EJL�6F���}�Ye�Mq��`����EtP<!
��Ь��Jq�@��Bm�!��Ss���Y��r��j�a�����Z��ە.�=7@���F:���[S�+��'C�����v��M�2�v�S��h��Vö��w	��D��x�ۧ�ԉ't�&��8��
��|��BZt?� 4QR1#+nG��>�)l@�O�1�U3�$�g�	���,��J���KI���� g��_���h��[���	T姕�2G��S�mc��~c�ȼB�U/��z[ �O�?��{wj�+����3C�ER�7��o1�7�!l7z
I	oP)�KMG���M"( �~��z�����-k�����Xl��ߡ�;�B^�4�>F��g�Ќ E�F��-J��pBKq������u�nUs��CRΡ�l��=�sWĶX���U��0Yi�����D=�#� '��C�)�$ً��OD��dBi��f�D`���Te����.Cf0^4�I=������I���0z|� ń�w�nEl��l��7�m�z�|�Û�Ǜf��_	
ul�og�; ��N�=�$qPGo��K��E/��Cs�e\I�R�I'����&�O̍\t��?:g�-����8�l�gdK�߆
�|��hൿV������e*ֺ9�����4�Lz��bm���)�{c��&E������.$��$|֥���V�G##��z��2R��rb���|�<�Z�>�F��1�9��t��y��W_�٣�ܥs��;�;�G���MV��Zv]��&:���7v}6 `��n���̘znkm������)1L>�c��#�>�A��IAd}s��T4x�ر��W��x��hpN*<�u��<�<k�Έ"�31���ͫ:a�E	��+& :��
ZA�Ώ/�*K}�D���P^.~��J�d?{;�z���w:>Q^^_��t�C;/O�+�|	�t�
w��gvOv�D�T�Q�`�5�@Ϳ,bˋ�b$����R#p3�LJ��l0T*W��/�GM��`[��:���ˉ����0^���o�`�En^��q{F�/����^����	�k�'��w�p�ۤ���b(��K�bQ��O
׫��c�+������@���2����uP޳70ί���ay�+g���3��[���&���(�T���<M���8���Gfj�9'>��\�KE�������FM3ѵ���;����b�^*�t��ɀO����Knljd8�6�u?�}��-��GK?	_����t����y]�#��tۧ(�ɗ��y�V ��r�KR�'�0��.�m�<�+ʌ-�B��*���G_�g_*J#��v�<z�.&C]Ȩ �m�p^��A}�f���s�K���Q��ߘ|6 W��R���$=2�0,w���/ݡ�a��(wn=�s�ޚGk�FY
7�ճCk+:	g��s�&o�V������ZXmc�'¥����\���J��OQ���ATiLy���Mn��Fݑ���HGN������"@�:�6�Яf6Ā��l�s)�s$D2C#���铰?n��J���̚K�?>4%�?�^��l�N�N�i�.�R�hv��m�)�A��V��`]wȲ�\��g�c(�\��RR`����&����i��x9n�� �����J)�#�۠t'2��-�Á�Ψ����t�[�+�"�{�u�4��g����~p�ٹ��v��3l�a�۹�������ۏ��Wח��Z��������M��^Evr�&���!�I�ۻ���+�N%%p�(,ϫ����?�>�g�׶$�Z%"�^�̏C8М�EM��0�w�?g�a$�!Ĕ:��t�f��<��^�}����������Ժ�F�.��<aV.��g��<D�+k��D���>d�щU`alQ��DÓF|��f�g�=��M�K���ˏ����)u���F"Ѳ��.�;_�F�P0e�;2��랤]p�ֱ'�F���_e�2+(V�R��	����ԕ�Mm߼��v/�4o|?�d��Y�]��ƣ�z� ܗ�2_�*Ə!��	2#^0�lg�/�E����)V�s(o4�J��I�Q�T2��_���V�Ǧ�"=	ye�x�`r}L^�|�)����e�y�8�D�(1S*���}.B����|�?å�"ؼ.J�"��ja�޹�ѓ���dd��0�� O��u��sv}��}�I��)�yXѓ�z�]��(�Q��M$]��_n�f�΋��	��(C=��i$�>l�ʚ�'��$�/:��Z�#�Xv�k}L�d>QL���C6�\��)�߬��ި0˫���l�����iͲJ}�D<ߏxqzA?d���ɧ`QK9z�e������Uj~��$����6��s60�c7jޏΞ�Iu>1J���)x[_�RaŌr�p�7��I���x�~s�ޛ#Y�:|��B_�,�Y�	�����'�����ЁD1�r@),�!L?=��t�@3����I���۸̔���TɴW>H/y_b�����:�x���C��O��T E��$`��V�3�+�^�����N� '�`?h���r���
@d3:��]�1J�J[�����,k�J�:nAS�����{K��ʌ)���9�So��-�2�qyx���.Y �{(¦�T�H��Va��%�>4^l`��'��,E�ŬO�R1��}]�Cցq�N*�~!n��>`j]}����{���IlB���E�w �p#G{7��]8A���Ы\ډ��y��ouz\�7ՌW�*D��U>\ڮ�L4SQ�8@ii�����Lf�C*�j�*��JW�|�&m��������R+��Ve���a�t��?c5��"�z��Ӫ��������f���L/V�&��t��I�*�ca����e6�3�uOQk����`����e��"�.+?q���"~�:5`1S���ʢ���5���?9Q-;\�BF�,PI,�=�'���J3�'7�
�[Lw��������;*�w#:���(Q�|V�7���}��"��nR���䰚�D>�٣DFoK�w��(H��to.N�նh�y~�3���씋�)4�V?	�&3����`�2�5W�uY�Sh=4z�ڑ��W  ����'�!WCxq����Iժg��98ֵ?�VK�p��?ss����S���d�!hA�A	�Z�$���N	����R� Oǀ�Q<�ӽ���P��?�z�<1���W/��ʮ��'MUt:/��J/E�
Q�
 ��VH;���{��Pn�fת?AgβF�?��{������k`�1����?`@�jn��c���沰 �&�A��v���b~ժ�r��0<yֱ�˓�Mϥ'�s��M��4�̇+A�cL8U����zRSHQ����D���
�{���ǢH'����v#M �ON�����f&.�}z�O�x�Uв��*���W����b��5���N��"K�׻����Q�(����^ 4W�>t_���U�g�k]��Is$��߯r껞ר}�À�f+���ZHc�����۬,SOt
ۿ	��1�>�Mx�s�g� =��뒪O;3��˷�ϯK�맪�Z����A�9���H���	^E�4D�Z�C���|Ǖ��YH(�\%��OZ����Ӭ�s��8}F&#ય�"��j˻d��?�9�r��v�5��|XMۍ#��E�̃�#WUO��"�Q�^���>2;��;�M~3�{u�lu-�%!9����Q�P��U�X���k���G�ã2h��V<�bMy����JZJDR	F ������w�@�a�����V�w�D��"1�:'�CA�O�<BrF����(J������eHbbd�:��я�� D�	9?�/�0��kFa�����C�1 ��.�S��M�8� F�x���~�|���ቁ�LJ���l����K��,���_���9�q��b/��
���u#�O���ɷ@O��u��BD#Qo��9����xNf�+sI�#���D��]w0�p�uC..��Zz��� |���Օ�R	�Y��d�o�A�E�w,$)�+7����A3}��E����ٓLᚋ�X�j	�R���u��� ��	�_*�mΐ��{�����������ܷ�E�8;�Z2��*qIk5���S��g� w��n�����O	`��x���Er~����ihF*��(f�C�>�1>�~|eh�o���R �&O�Mj"�Ҷ��ظU_H7����Yk��2��N~o�ӑ��L�.��p�ر��l�m�F�m1��a��f���cMY���ᣣ�;$Mz�[O ���Ԅ�ߞ��?=�Ʊw�m�*1��)x�x�ko�Z�:m�圾e�����O��DNjI7�N2O.�Pj͏��*�U���@{����y�*ڥ��ւ{�5,D3-л����"��n)QQWq��U���e`�	�S���\8�c�R�,e��{U��[@���ec{���
�