// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:29 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G3hZuXs68rNu6cUdMTckkyCtbsKvqWSUtS3Knr9U7NuxRtdpiYHpYwWquo4p1jZa
B+qwv4Sc2HxZatNcS4djr6xTPdbUArsj59B4rww3WZZXqPnu/yjokj+PzkJzZhsP
u9SvGbQxeZac5W3QNsArdxFdH1G5ZmssgvlQywShoFo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6704)
tQ54Ug9aq1a4PbRW5zieQQhyxr/ziXpWgxz7L0a0LJZhuh4rhNESWsqaby7e0ehG
9ObO7T9WEZsIfPdiKsvVsvYO+RuQJ1c1+EijI2f0Jfcjtb4ZUfezri7xMzpvbui+
gDoZ+AxtDdDuypDjodUZeSY0zB8HblbaJ6rYrusvJLju+xTUzQdYv56wJBEeWlkP
CHUosZkfaDr3OHoBqcLIS/DQp/3NJJQQCzOd8YSNoGhFER0Q2Rg7kMZD2Ph2CqQ1
Ivnd4lO7KbRnI1R217ptSXScocl8dzRPxdYHuP78RyeID+FUzSlaV/NT0xgL7MQv
FqUyxJgUMIB/SuNr0gpm/afHZuFaARkSNZpTxN+90k/Nqt/y3ci1RJWW3UbZ7xYC
GvEhI9bhVlCQM53WSMl5KSy13N/0/qcfia4K2S7xuQk5hCEauOeVcwe0KDRr7Rm6
WsnEqIzArN9GJI633U7X3iwVZ1pwtd0o2rD7+8zdnWtF5Er30ZRRtnH1izZSsA+l
Sj46XoUH5TeOGKOqB1GAtcyzppQdA6sTv/IZa3370PD6aupYrQgjDuE02OU1SxI2
uCW5DbbPaBj5R0Qt7zSO6Uqa/TIyFGf5UgtuIr6L1cf5Wltpzphcsfv3o3dm8eM3
LZHsenAnyGYbArdzTk98KqviftZDU3Ee34zSi47mz5ggCmiH1FiJ2+n9l6eHl4u1
HoI113tdGoddu0DRX11J01MRsM3nVbDi03tDvtSruQpvwOeNyFn+fkhEVnou44/B
TqO94JKJZ87iBjpTBiA5tqqsf/P2jespUIp+t2dx6f8hU6xYycc8B/7QwVvxZdbH
tU161Q/TcUEoQFdconPdgKo0CE0/tEga1wuyrORf8RIl7+jVYxQpEtKKr9qg7O/i
JVmz+aTR1S0jrKYiyixJaz94df15eh8xtsqSV0TLtcf0xuMmG3cn6gwbwAGzKPwe
fOn5kqIDJMatb5/avj3uyQ9kRokJS2d/LCPe0GRNJAt49vbvH26yThI+ujRe/AVD
UbwGnWcj12c5RQ9dRtvytRiVGp57z7QtRvGCo4uv966epdUPywmv4fcrQ4hrJXuC
xgWny91BTe8C5pkpr3ZNXwpFGh3gYEyxUoNx0BAp4IAYub4TAxzu+L93bb7VenWh
yQjD80QZjKBU00M8FCo/AvXf7DBrByxE36fED2+ck8dXS+kW9sWPcLbMkPJFVnw8
6fFJ0FDmdjUXrx7bIzOZLiESMngetQ4Pl48mUB1flru45aTZqXs3LZfWWjLksMOg
JJPSlk1esBsaycIDBjuFyQ6vd32O9i1dZQIov1/3J6rA5LzytVfLD6ck51jHU2xC
e1XpeA8p9C4Hc5RBaW2V6h2zh7XKzvN+WaxADAM7Y9DV8bbqFTGLtsFEW/vzKqIF
met9+GqNdJnOB3084/D8OO4EqDNw4BP6HfnB+7knjTX5L49xNpdhqmMhQv3M7w0b
UcJ0H2iXr7UAF3O/rOkspTXZMkitOw8EuyoN5CqwH1/qTr3++4+5D0RDYblw4OJf
kmo+1cGeu4P7R3Fc7bDJEewDMae+5AjcrAh7fuSsdL0dDDmIBSEfPz8f5SXf3bHY
GAVtr1ZMhPAGyuhNWWKQQI7oEEq68wISXIsM+AStViZqeOW1h2ldl9QdGZZfHmGk
KmQyy2LjdZzXR8fgD5EJZQfVB0K1U1w4PnfDxOq1g/pR3hWW7Chr5y5BumhqNcnY
EXCpXKlyMGc1ND5wihRq+UkqSqHtpv2fJrYoeGwTVh1hKg55YG1Ah19aIIVLJnFc
oysYfDnRs15JK36GEtQcITeoOhZD607jDp+klqTmOaKx8JkNeTcihazxnH5Ziv0y
KVjYpYtFPvqxweF7OLa/qs2e7o35YOwc+5ObLATffCcw6fOg9yr/uPeiNGyQhTlJ
+uIWNKdpsqVCRzpCnAzIIM0rnnKz3vPDyypRCvqV20b8m2KZRbNfCUN2zA4VSzwo
or5z9WxUhHVMJ2ORusfc+guOw65stqVN4GYn7uDhz2um/Oh3aQmyFP3c8+8ipCxB
eCOH9MwwA5wxxvDlyvgJS2u3/lim7LH94+ZmO07g+lo5kRubTcVy0GRRb2dp/0AE
bMCCcJkAkYX9hjdlxnrVM1mlKlb9TH/hkE7aXaHWM6cEelBzQQo9BSpFv3u6BHjD
BxTf4fQifEVZNTEiiHoIL9xeZ+x6ACvYMZJkoAbfn3/TRHM9dhTVNhe5yTB16cZG
wfAQWXCeolU7kUBue2edxtMeuEv3sg0tsDe0VBDEj0okLKdMW95mi2paRCm6nqSM
IzRDC/VDh2OPJFDxogwRPWhz5aK18Ey39L0Rnz7IcZLaD0ml/02bwGJ3o1nnZrEe
Jw3LR9VJGJ5QxUeAg2Bby+QQYlLQksMPA8TDmI6tMaAhPMxmt2VFTsVJpNZHgyYr
OzPWFL5iY6DdqPoNfRJz9Dx84sGnhcgHGG1lyBoamf1pQaRxJ84QXHsvRMlKYRkm
hNgJE0hwFpVB0yHBUGxjO/8otkMeMwnlUIzHUsKi3BiOMx9IpV/0HxFy7Thb+grR
hpHFq8VFSTHTjIvjHnh5rr+j09nNToNq+JZO45M5ckY/YTbJVd2vH+uXMUlNU/bu
OCCRfQ9f7YXJ7sVpPyQLOdFZETvnJ9Oe+3I16peUBaDZBWdc69iASoCNPxxNHFp6
adCXxabG9hLZx4z4xZgXkHvReoAmZZkXLdBoZFGUDwwrSyDScfo0CaRQaLHuR0oR
ENpXmbicVP061S9Wc3V+HWVD5PClxW76sdqn4Nb7wYf+xu6u4q7kbwDPd23Ym92C
IB34WPM70sm1ue/ipnSpuqEDPAEVU3PpPSDAVuI2XBdCWrzKok60jduKsaaJTuLC
fWC5VOvlvVkfKgFSouj027jcqdLEn/L5AKn26GKYAT81yCuW7mYmIO2MeSigT/W/
08WWR8zepVTuLu8C5f7CKscspokXvdlaKCIIZOpcWEWoTYCO07qjxEU2POQywtvt
6QO7aZ2FtYq39H/Q7YiiYar9RyZ/g5sgUKZkyRpM5NEq9U42GleHhp5X8ah6ejPh
OILlhGBRGchzsT8Q11g2BqfywTFmREWoHY1xyHXYkq+7gHrVYe3Rf9CbU+UlRuQE
a71ukAo+Uy6vjGadk4MBcFbgXGDF9t8vCgonfBguKEzohn4zKOeLBTmR266fQsBx
gGsGWbPOdbvdxd8ByGk6Dr03P1LB8kYin5ooTjQimRZ0AbUip4DcF8B9uBzR34G5
dhhkz1F6Jq5yIqLIBOFIHGdPwOfgXdbJzVkGXazPwGjylzbtDRoH3Dlbrp6TLU8R
ieuHQ+K5hApDszAK/NWtZvIqy5xNdVmZTsaisDw44huC9irZGOyExbZIf5AZ4gd3
656P/a+mXDSk0IYOE4p67J9iVZwFZkMwaj7NQTB45E2lH6LAgznjidz0Gzg7TUUA
wEztPH3nZkPxvflXN+XtyPmTSPWC147bIRPpFOJ4gIwYYC0gGFSjavwACwm+KuaF
dKJ/HehCW6EM5hL2cKBi8lWo+CeUKT7oChdU5aApleS+ls806mnrWqMTfK1YV0IB
pcYJ8sbIjHzQ/t+ObFO3SxGuYO0k2KVuI6msQp1WqFZbe1JuXlnbRcUgZ5AXAkd9
gaU6MuTeSjNo+dvha3Wh+1tZ7SNlkZAguK/n+9JCMpcDEI0JH6OpLg58Er0Us4Yi
b9sQzER4Dbtwd6P9f0doVRXd1gah6mvDoZZs66ma370cIv2YvxlakssEzYnPUzz2
Q+Dc06Y5KsrdcFusSkm1lb89gJ1fUSZA75lAQMeqXka9ko6cVOFrRQYA9fw6otwW
CWt8L3R9/exDSG+b6HMaTv8g+tJSQnBz2ms6otqom1PWJcM5ghI847O0O8LJUll8
zWdKgeNw/oFr+xPJ4Bz1AOrJtkI36bn+6ZJmhDQDJrBdaTtHrtBOqNM9dUmKVZTe
JPN7Z7b2O+LmhgEZnaI7ly+blkgkL1/ZU/b+r9nCdIu88DFjKO1ZdSKpJCbpswg1
weEdJIlVswHBZO2radDRmlT1jvXALBVpXSRypc8jFCtpN1CTnE3E8o/QKxdvJcyq
F/N0CyngrjWxkjT2C7o9Z4vhORmKEcObIkfydNmx0B6ECCWFB7FihOrjjcu3CS7L
cdgoh044gVcYrFihVE5rrWhQqqKHkLp19p/7sMStLGGgKxyIFOugJRHBTXYSqSY4
tJ2/dIQC60KGjnLsyB1wQJxY1ibwI7lctYx22xHLuW3/c+LW9L0azz15d/q9IAN9
ALJmee/cxZ8Q37Z4PyQawtakYe0yrxNRc6AYdU3QDBmadiIAmF+17E73YnuB5ddR
fC4ezVFT3bkJUmGk0XTz9KCO2HfZh5bbWN+QlwsX+ik31IRfEiqn7MkFhQP736Dn
D69spJVwzE0iZXrXmkfWqO4/25bwAEuA1PqYXY/pZ4bUbMd/lYvsGkITcTx3J+pW
CLwNfkr1hDlm5F9Mw8yObp6jEGeK0nF6SccfQ30ebs4ldKsIPcOOm3t3pl6hI6I+
t13vR/9wl6kig6k+Fc+GPzxjA4s/XqiAAiXHUWy2j1aViSckzgGOCNOWPjVm0Y5k
q87zvkunft8yZ6pN6IWZ0OFk+6c60riOqaiHppkYLn85a79TLLCn3IHxgKelj2oi
xOPJ+SJeQKPCy2NAOzO7R2s0ZV04jEbKcUWUx982VE67c0E+c9bUQg7stw6HluKR
ikSugRqMVYR5nHB3zcN8+fNFnvgVqgPzhrZjMwgrf9tBeRecbHSv4tEtVHzwG/H/
yvAAg59YgIDOZT40SiQw5UnzYcoOFY3ZffHKURU9tVYHn0yd5NgQzSYp+W8fjBky
qhSqUAHvtizkNPJFGP3FIAgHxeGZUELqvT49AF40LdsKDunHmGzYv+w0PxRoobE5
xSDeOtn6UysZiMXQJF72aMkd7XmlX8j6KsTDww58zq7W7PHNFbc5cl17tu6KQJF2
Gtojq8SUN3FvGaIg5DWZ1dZun/0c0x9ESxIkYtT9CsAnUHQr0Sj9vCeML8zQUV1H
oU7EL1l+a5D5vCoBNm/RwhO39iDljVk9HsgOnBKlfaRcCwei2j8r9AQlmV/PIFqb
NoSZ0LSCqdFjg4OrKCeqSH0hPmTovs1w8qehNxLZ/oJ5E9XE0Y4s1r/SOx7zXzLw
b03FONUxnPULA9twsV/1GMed7OGXLqrLJzdQ5+Sb6HB7mwTij36vru0f8IZ9RQNF
24pf69uhp38KgP452WFK3fJIg3J9TkTybqZsFFKWCnXPWV71NEejbweJgfPAVuXu
OF+VtnAYtlBMgxqb1fizz48xLnmq+XA1h2xuIuzBA1pmg6YXLUM604NKgXINVbpn
7utef2pBuE8MPpAddn6Z4C0gryWSXAhn8O8zIjnmWCFKXOcK/fXH1Ql2DHzwsawr
ltOaEstNw8PUQip14vTGuHIWuNxfAVqtYzQ9KDJvPF09b4Pib9JKf0kty5Z/Vpvf
WnHWNxKpKS8iW4ReoxwHOV3tngVhzLkdMejY4icFe3O/DQfWkpsozmISpWyaU4ii
l/2mXvS/mYa8yCZHnp0cUN/hkh5dXRkFlMW+xoSfImpJNccGzThTVs7jkT0Kb2KS
+5MNBw9avev5WmX6Ez/m30FA1HzRdlYFoI3siT4lW30iulalDXIZ/QVTMcCcQG9Y
lvVZ2m9qqYfSwvx7iXwJs6GUXq1D+EAufey370KGsZAzvJ4Cp6c+8TRU2Vf+P1bd
Stc10EgbQi96pvQWG8trGklBM5FL7GmGtlNaOJQUL79SsL3tDXS5vb6uoF2QgCTY
HNPT8u+PbYRQ9tU3WIMcm1zzW1RfYYN0fGqc8YS+7zPwak9Leh2pkJInwIyeRzxa
xZSwDTF5gIUULRh72UuoGBJIRa1Rp/fSa7Atqjqe3K6P24eXTee5pZa8lPe81GnJ
A7/ZHnmC3Fxw9zxLWh4ZqtJxWocY3omk7YLJUdGhKHuZLGQTH8ZOPA4Mf+pPDK7R
oscsH/AUqMqz3VFZKVKRiQsf3eCwcU1UC9hkjgtYTlBmsN3YrarfKdaSO8rQXbKX
wGsi/ua8ZAoOumhzztA52LrbeXOD5woOttoQD2583/hVd5bm2JzadeY5hlhE73+Y
fL1FnTliNRZw+Oqdeq2G7uWm4HICEXe4p0iOyLKuPo3l1eGjsT+1ccdaMtQtYU+l
x7GxAKs9qtP2LrDennTXaOFB0VIgYc3Ejh581ueObcPKWo+tS1v/XaJghiTaQ2r6
1FbcpkkF3hOHMwqcoqjBCg9jLgD9kUYJXF1JzqMiv+1tgmmEaBfR0KgJXD0LyVgP
ciT9HkIqTSRRF57Jbj7QSTIM6Xuavfj9RjJU+HUGImGYburpcjM1nGgI71PCHVZe
pnwHN/awPJV0MTinokeUeyQs+/3kX0xC2T3n2sRFFqtokiffCEQd1USvZWTkrOQN
bSjgnoYC8MwY/hsE+oAfSC3TxHNTHrTABSzvCV5fqy3bKim5FeQLbY70dVPhJQdi
Xb1qpH+icplVwJOoEDF+VmlKt2a9oTt757fuWGW2p61J5Gew0VXR3rXgUcGo5BuV
KprFWfSA04gt+q57YcKkQS6eycpPPI1kr/NKk3Em2O0RYkcGtmxs+AERNQHOD7JK
w29rWVvpZA+jrJ3q2QQl5+44J8kzkzw4O1TGQQEWhRR2kler61WU2QWUNOFzyQ9p
uX3nkInxWqH/WXyPITnHYI/EM0Fp7yNPHPMjeCANZQz6z50Ob886T2v157mFCyUf
VrmVxFviIJzQcsfOa8lZ5WY82Iu17PpZfk6GXZCL7qC4glxtAqmZHf5Xs+GukjNZ
xuTVwBe7IwVnQCmjHvu9W9/20FIvOq9Gmhm11jXj8TY6j7zGjLzimg5byRdh7n5C
Gxd+KxqbC8BgE0uQqKvgNQrV6E/aTkFggCBK+H6QjCgeHwwb6lmtUT0VgPFjOX4V
SDAk72JfTY6xoYaX/bkVxNj6I8E2MjBQAu7eTP1zp3qTxGsDvG/7FQ4EqCV78SrW
hBzs2csdudVHpBz4uHDVdCC2/whgDMZTf5Hi/LRgr3fjql2YCMu1uX43czrfFq2M
qUuflEOec5izSgGllw9XJ2d0dkT9jcHfl+lLOtydvg4/Zm0yLUH/+V6eL6ANxp++
aMjtkuxzj59d80Lf1Pbydbqjrz80LPA2+Wv4cQUV101jk9uJLjLPIdOZlgHZkUp6
N+C1gqPchNZoE+Br1KHee2UWGK2KZrabSwtJJw2gIEFxuXoEEG9whsVP/WLdGx/z
U4Zw+rRm3Yyoyf1XID1kcyphgkujE70DlRqEluRgFuey5FVrnO+8mN472/ivcTKf
YTokOrEo2pCmQnL4ZSU+jHQ/mzhserLW2iOdXVmwa1lF3rbIL2pW5p//AMsiIdot
D1Fhmd6iM5F7zWwO4eaxD3hAB+EG3GT2CAfv+RdAYh/GaMItPLLbocL8DrDugoBy
sduBSpN8obBKW1dxpMSIVGe6bfGUCTw9gTVN/imFRn3KEg8F1b4kUXtRpcy3tEaJ
quqZFUjEh5frAt6p2yAVo47NMfdtGu1Svqfjrx7GG2bHzTD8DvvJNqoNiaLTBrfH
3HBQOZRcsSjydZwHYRTxUxwe1KYPeHU5W9tfb7/uyBPfEUU57efceyOVqFN2rhSy
6Tu3mdUGe7h7NwG20lW3lfATZ2D76U39bFt5Se+Zk5Oc56jgHH0/d9ydf/z03Auh
hw0sgV94fy7mr3lFjhd+1rBzJbEErOcyit6gwzueBvDLpjYQc7tBwAT/sw4dG/Zv
+BzofowZBJaY3QIXfVpYs9iVPOPnDEf2XuL1svQV0i4Ik7AZKSsRUTljrOu1bUkk
qX7izrpLF27LHcrUFP998GBnuv31jxDnIFP05XN6v/JPyEF7E0koQdBcRSBkUDHq
0sJ6Adt+o1AYpc6cUui88u5hJ6ZIzHIXMBs3e2Rixr0jMVsQ7IilZJBMWI86+i+B
g4HaM8bh1eH6nvkhaRvbNI4bxnMDGN7d8xHZO6TkSSGH3e3DLGsG2I4M/pUUKJva
7F9ZFvJt44BFenI04KiDCjDSO2QG31P6zSwPClIaFOojsDx3wXeuGtCj9bu9CarU
x+4ti6gjS8VBMB2DWDoX1wYf1/pZ6Y3iMp9r3QyLDhX96LOZ3V4+Pc3W6uicE1YR
iwGd8yQC+JaJNSl/Lfwcw5MgVHRVNHvgcW3QhxCOs2+9lyh4vD9e1VVC/ePUvGZC
nZENGWGfjjmhNy6IXpPQdPEVAsr7JpZUhfEdfFAv+Aj0jJB/nnt95jUX2RDvVL5d
F6TmBCdBimuhaPcVgpZ+U6+qUaZ7cSRK1fVFDhxosgUZMtm7I4sdUJYmh52dDqR5
ij8yr3vFtkVGPOuPNehaNh8TNOli7/PYshR/GQ7aaCFUSEsqYVgKq3VNmL5v2CL5
Rm0sVSCxF9lUadc8N04JRrrDBTNsjl+w5kgWy56Egmvyiy7u9dy5RJ61F4SY1sNc
+jb2SzOfdQv5q0MRyxV4NoR6rILL5pu8g5TZOX+OH+h/1FfmYtsztbyKl4UxETJu
/nnZCMFNiZckooT1h8JrtOQOR43FlGzGXMpluIA8hgfVZlLH0tcZf87pu8vINPGZ
oystzwu3DOHAgf0mPRhGolDvF+8IE7tyROYMxJOJnyItUG3iFlMTqkGYGm6PErlj
PCQ8KhQPszSglfwZCDJNM7pEtadVdSmoBg/GAJWq0o3urBftDi6j5dwH9FbzNhsB
Q1BP0zlUROgrm/A9Hye6GqnzkWuADRNcnl0W5KJ+HA0xuTXiUUf+ivLTQwsIIcrv
y7EjQ9bfYBXFX2/aXP+oHBQiSYrqcRDVY9ji1a7Dlz2iS4HYPP6I0swJ9n6GyZNk
8Smn2F70MyizgHvsM/ApTBU2Qyz6m+Y/LjL5/nVqwEc=
`pragma protect end_protected
