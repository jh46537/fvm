��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�����jA����'J��V-�@m��Yx�W����A�.�ƋB8/dq�4z
�7�LJ��e���OM���L��{�`s���[���z~2Qu6�Ѹ �5�7Y4��ڄ �d$��*wP�-��������G��S��4����x6����[�u�s.��/��j�GE��r������ܐ�-(ZhG�( 3LnC?y��|e����Ϭtl��.B�$�یV����T9H��8�EA
�C��f� xKO�E,lx��'#C�����Pi25����0W�\T��L����^�n'�k��������g�-�$�����h �2r8��9�"WH�I񈴁��D_q�'r�Q
�bͰ�pYT���oz����N���H�>0<��F}(SK� �P�k�v�B��- ���9�b�$i*NT$� ݊m��չ#���%Y�	�&g�(��J�"�3j�b"��JěI��r~~�u.ވ�H����]����׀��o�3a,
J��ί��T�Θb�\�m��c�@�ڏ�p�����m��O;�ޛΚ.1n�������FA>e� �o!uFڋW�k�s�c��Z��c4�h�����O��2�VH���=�v[�G9�h��������:�aX�����@,�S�ãCU��=	?��C}�c/1�����C�j׋o�{��kXӄck�cp]]=�,,�����1�D�f��P���k��`6'�Ǜ=c�NyAuhWTaL`� U#�����-�gE�(�����"Ie���ͨ38$��ŧG6f�@SH�l����D���;�]e��Q��#������B&���(�zA�zc�Q��ZR���y�F�.�>�[<Hi-���0�c��F���W^q4���ۑ��u�/g���da�_�h�|l�uh��E�.d��ƪ�:�oE�Ч]�;����d�u�ֳ��NŽc������?�'<JW絴�*�T��o.+�o��3d�Y��r����+�#G2�o�u�r�M�e7�Z��q!�]�*����޴*���L��*a_)t1	Q
 u��]����.Z�+�07T ��a�H�_`�|Q��D}�������A�ؤVqe$ᰭ�/���bD$x'3�jZ��YӛԨ�!1f��v
�?r���.lr+��z%qm�0��P�ٽw$����OGbp�\�ܥ�������9q��抰������J7�J�g��,pC�2c�薼���V��h�gIHC]"�x5��u������������A��5EO����Ͱ�����4�R=�ޣ���V�*�����꓂{��u ���	�0Z|�)i���t;�4C��������;���'#G5X�ӈ���f�=7C��y��ew�DKGo�����!����^�-���w�p��1AE�kK8�����Uzc�4��q�������J��뚠W���!���M�qz7"�L���8[X��VAd���,�ڳ��#_�#�ʟ�ңf��	)!z/���?��d����Ņ��P%����|�s#`�1��T�cP�S���^�ѡ�Q�{�4����;�ȩ �~1�U딟�5p��flv�tX8DPJ��*�� ��]ҭ1J$,Rɚ�%�.�ˋ�- 3�5����rG�nkz��$,�u���\S��3	��OA'�tG��p63���2=�Ѕ��y���&��|�U��*A9!�Z#�Q
�}F��W����s�q`_�8��M�3��T�j��w��sՅu+8,�-F#"���%�x��N>�!��-�$���k��������x^W38�(�6�'6�� @��%�]Oc�m��<��@�=l|Н��4�� �x�����8*�Q ٤C�7e������IÙ��Pv�Ӭ�,�;U���S䄞��쯭؊:�aX���%B�A�p1�}* ��*�I�;b��k���2:�;T���CQ�!��uJ�jZ81� "���؏6F�����F.p���~���"(�8�:C;�%Xu<�ԋX ��k�*���!_lZL�~l$�����1�Q���"�|��@��&D��HhO�������5*{8�;�P��~ߘ�8�pڹ$43�7-�[s���ٽP�Ԩ�j�A֔씧6�(6��żO�?-t<�������mU�zŜ�S�A*ܽ�6�|�
<o���$ICD ����������ɣ�}�=(�WiWҿ��]z�� G'�������`��*v�6�S V���9��+Q�>�®�����k�[�����l.(����5T5˸�McU~V�ܩhq�[����Y����ī>h�p�zY���q��GP=n)��h�h�G#��["�����ƅN�����H	Q*�+��k@���0�N�"���L���%���_cæ��@���-E�pؓ�[4���C��$���|�3������ȎFp�v�6h��R�]*=����� ��x��p��9���2����\?,F|58���?s3@tu�F�U��pIU�HTfR:.h��>����=_S�g<�^|����QFr�	��Y�E��-8�r�ŨN���k`��=k��W]�g��	�;t6\O&�E���,o��[o	-v�q9�H[A'��/l;k��)��G B�r4��%.��:�u����������i�b����� g�s�vaiI'|�ӽ��cwT�һn~�n��/��Zʏ�Gњ�m7 ��O���^�� �E
��TPXF���=��8%C)�;�J~�I�������F�y[R)�BR#eM �>}zod>&���=�_�ߗ���e� ��ʵ�j�\�?2 (��4�����h�D:�,4���k���3��1&*^�8���1�h�sJ3?4B�e%�|���rb+�р>Ӓ�<D[N��`6�����Z��c�g2�17��N�@Z$����C6��ύ��GUʇm��^}�9r�1ȍB�79�}U�_�P����F�[2�]Y2�}5%ܯ`��f���~ʠ��Z*Í�����Ώ���h�ں�*�M��>w�P�h�/so���r}{zW/J��}�&V��%y:S�l�WOA*��������5$eϚ�n��Y3���39,ʐfX<���|σ�1�f�U~��i��O	W0��T�\�ّ֐��*�8��굞QHG^�5l�c�*��]$[�W�-��z�]Mi�"B�^��u���_��æ�����a|ف�aF�̜�x��9q��t���K�]�pjt���>����!�S!�E%jd��2u^���Gm�;6��qQ$�[$#7��B݌��+�oGy$2�^�<� �Y�W��V�R�������q��o��Xʩ��Z�ȂG�]����rk]*���6d�o_j���À+!��d*�߉Ka=f�>��$(�!f��9��\����n�̀�D����>���&eyCT��V��� �63�6E�@�΍��&�:6?�ۈ-�[���1����4�I�L\�%���h��wx�a�/q�ϏH�^ٴ�N��峸�:(�D��7s_�O�8˦d-�FErV|��OPԞ�n�5�Ѵ �>c��0��̽��,x�o�R_��չ�p
}׮üz/�Z�é����|��SR�0�N	�c5$Z��3��ά�9�eCB������#�Qά��&��{��!LHnE]D��x�R�&��@E#�Ɯ�W�̋G�-���GI���z��I�ʢ3���!_��\k��z��Q��ݓ��Y��"�ϭWH�XH��	2����n���d��_DM������;	��l�&�&��س� ��
,�X�c1I�&$a%lU�9s���h�vUfYJ��q�4�L�asm��;��8��~װSb�6P��k����ķAJ�-���qy�����'�'d`�L�
�oO��KOV��/`gJ�ó�i1�	�ǂ�r�<M`ܱ�d6�^%t���5�v�F��8��r�]������͗Z�f�dP��s���=t��IF�/w`(o��[�� �R����=2X��a�4?�'Cq�6�w��U壛�����f��O��m{7?fo��a�/�l�Q��mm������6�=�Yi���iU�N;��il�X�W.����o��c�H\Gƃ�:���D����}nt<d���~AC��b�uR���e�xϕ[Yl��pq��0�.�W*�����ut�
/�v���L��|8���g�r8qH7\�	ڑ����j6����m޺ŋAn�u�"�edP�i>�3���i,���H���˅�;��A_�SK� �We�W��m�W���9L�w�����ΰ%S�jӛ5./I<�:A1�p�޷]%��2�GFZϟ�qL��j�	�եp��k�ޑN�v�S;����ۉL�z]�����觫^x��aś�A>k�x/,�:q�1@���&��mн�a<��Գ0e�
���RL}�����l���DM���K�q�鮿!r�0pŏZZu�Z١G���_����H�\����_1�LS֝<�螅�����lˎ}��(�RYԓ#`���0�7�b��<�ښ3��/d�6(�x�a}�U��V񆪒9Lﶽ#��?��ΌHV�xS���q��T:h�x�qX�����~#�]ߋ#X����P�B|�$^�@-^�9*�9#��0��fIϔ�p#(B
��P �ER�|�H ���5l5f5�8�A�W�j4�:����j�6Yj�t���.fVڮ
4�A����%��l��k�xyc-X	W�*&4I˄c3Rlb-ay�O��W�� ��V�S��Do;�~1�=�N�Ȉ��!�I���Y�z^*2���S�G_���x�J��'2��ƛ�����,J	"�-�z1�޵)�k&b^@}�j��1�6�n�RÀTl������U��$���G\�ey�,a�.(��{���yz]�/&��^�X�wk�&4�ݸ!��@��IuyEF�� �7H��\�J���fE�
X-1a�j�fis\��g�=*m���|>�ՖC�n@�u덲�ӛTwE�t��Ryg�n������{�#o�%�艹ͭ��5SϷ�0ld����Fז�b�uVC�h����Ο�{l�i3�Gx��/��w��/�ad<7EýyD/��h�FBgC&K������2�mi�����:��]!�;'%��o���D9�f��D֡᧏ɘg_5�;�,A�z�-�M���ș���
甇fs�����6ui��}Ȣ���!D�k~�E� �XF@ �	>_İO��������V��&ΖF�"�Nij=�Z1�XV	ʹ��������+m+A`Dp��c��O�?ݾ�t����!��
��}��Q��d7�'�S��D�'cE&r��g�-/�w�Œ�=��3  ދ�gޣ���'!�D�^p�!��T3i9u"kl����i�LEa(���RFͪcI�\�QJ�5�0�����S��[�H]�0����97�pe�N|�+Ձ�-�F���X] z#�B�T�oi�}��VU`�x��_�/��Ng���9�j�G:�.k��QWqz4���n�pߔ�(�1�D�g�S`�G�N�9�.I_�8b�[�p=�k��إ3E��ydB�;~/ݨ�κm�(K��h�������jM��Pn֕�cSD��=o?Wm[�$�sM�����o�Pyi}F{��[?I�M�y �wʧ:Y8���?��ЌL�e�U���o��%8��)��}�#i�#Sޘ���^!��������j��ו���4�1&����)oT�O�#s�òIh
7o>+����11='|���t�"��XO/X���6:q��8;�|$8'�
�����k���酒�C��|��/6��>�K��w2�Ys~�Qf ��7�Cgۛ��"HM�E�i��^���b��Y�=ܓ'��W�9�T��ּhPF��^�	R�;L�_���s�ߣ\��W�\B<*@�ߧc�~~��D̀/z���n��d�m��pA�~C:�,8�1Nr9I�U<:�[?�R[�#�l)5�	?���k�XЁG��9��Hï��g�p\��-5�}�]Z����:�oR �8j�1x!� ���we�W�h� �Rm.�>d)o�[yPG�b5��w����1W��F:��/�wt#hŃk}|�5����"�4"��'=�~��:��i}1"v��O�p���*��"����������ۺW��%������/b�9��r<���B�����53_�[IN��i���#�Sv�17�!��r�����ʍ�/��Y0]�>�c?!3�7��to�$�,�s	78�E��vI{`����x�S�2,�_�5�Y{�I�m���ch�+,����/���J �"ڟ]����iӢ�E�QF�4Ky�J������ �6r'��W�(h�5�ѷ�W��y`��"Hh
Q
�
*�֫��l��2l�vS-֐�d����I��Z5&��n�S�Pǳ��bf2�~��������Wo�Y��&�j�*��pz{���V��Є�݅\~��!n	�pJf�m �s�@~�$�dʋ'm,u^.6�={���ȡK//��C�����i�o��8�x�hk���bh ��wU��{X!�U��_*ѐ�e���{Ʊ�?�2t,!`5����w ~&�q~���㟪�ơ�j���~���OK]�	Ƞ/ω�TV!Wϒ����/��5��?ٹ���D�=�4���H�y���DV��DW��&�7�z.z1:�0waq��"j���"��lU.JxRΊ,���:��?�}�06�˟�,z�6r��\���r�����#��8��)��T�-N�Ā���� P���[(����ΰqC_�ԚO��i��S���'�k|�#�2�����f@�Lڸ�[\0����ρ�C����j:��<�{LQ���O��[�F����k��@�D�ۅP�UP�FW|��_%�ӓ:Ȏ��;�![�ݎ;_�J�Q������U7�/��ɞ疣��P~1���O)?��N8�,�E��{�73j]8