��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]ǂ��O��˰�	JL��Guy6A;��%��:Ԩg�P-fǤwA?����u�n=|cc�j�/���\6[_�����l=d�m�VQM�v���Vhb�7U¤��:*ˁI�5�\�oC�����h��U�-E����;tr!��&�гf�p���$�a3���%�'�G�x˘
���� (���_2<���`|���؁��%j1_Ιs�ʐ8��I�q��l��"�a��Z�V=�^���1���A����2϶�[��ygB�XJwya^*���k�E��h�^-s�p�!󤌡C����a�TK�y6������	ˢ�{��`�g��p�go~a�B���p�z�ޯ�i?����ۻH����ߏ���=V$�tpw�~�	�Į;9 �
�����u��|����.̍���#�o�u�a�D��q�[�y��uӑ��u�2