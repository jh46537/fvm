��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<���Xz���f~6>���꠼�Y�Nx��<�y�����笵�)$=a�ԏ�s.6�/�y�h�]_���m�ix^yl�[�I��/�Ϩ�X�7V]!?A
��-"���|KED_Ύ�t5��9
�;c���a$��
���W����Q�u�HG:�w�ְ2h:�	)����G[_0�lwEt�� ��[k)K��>b'��m���4ijR�����^*{�@�l�ӗ�tBi�zp�Ծ�>ztӰ���2`S����6��o�X?���+r]��geиpD⢎P��J��~	/5yt[l%�d����L�5V�S�'3��k���p�hf|��~�#?��\;�a+>}{KJ{�z�$ɧ��=C�u"�\�{��A��yĦ�O�*�N{��xɷ!q���x9�xƩ��q��W�rƖ�@��ۚEx"XyoY(��(��P��׭($c�+O=��	}�P�F�+}�׋rƷ֭eU~�?޸Ku�E��R�9�^�Kɡ9<��!�y��v��e\��*�yv=�M�*Eju/��1X*�"��P����$~�f�̹����R�h��VJ��/dF`@!'�I=���2������֚s�">6Q�����JOgN�hԦ�*6������] � �=��!�V�H�h�[����v]vkL|ƿ!I	����L2���N