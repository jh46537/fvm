��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�����jA����'J��At�JD��>�dtW����.��E�?8AҰOU��d�%���0{f\k��(PO�s��@�h��u��	=�o�l�s$߰��3Tvqz���^*M��*�\J��.6 �C\	�ڍ^��y��e�U ~"���^���#���`��gvuc��ޙ�b`�ӯ����Kru��"�l&�8�_�8DH�XIC;G�Z�^�%8j>@�gl4}���|XC��{Փ��՛����4�cw:����_��x�$Ұ���\s	2�:� S��:��w�H��h Ώ��pG���@�j���s&��v����Vl3�e�b�a$�ZQ��x�|A0:�&�;���ő���2�����Ο��Z�P��Vv�g�]=-Y�T���e��+��F]x�7�E��@��S�QH�=݀f��w����E�̓H�bP.5�η���9DW��$���i�9.g���(�g`�sa���ۓ�QNu4�a�B�&�b�)�?�ڠ�!�VEr�Gr��a�x�dh � (П&69�nw)$��y5u*;��r�N�m	���2����orڲ�|�_V8݉MY]0x�c��[�<%���tF+��h���<8��Q@�����X�y~�v-ZΙ�Ew3����_18��� 7�U���Ӆv�����B(P��i����u�߼$���̼+��c�m�7��vR�{�4ݞ![�ZU_�n�u>5��� '8�X��M��)� c�1���fI���F��l��������\�^PEn4(A�s��eY�I
��0�;;�*�B�p��,�sԶg�1�S	l��.�;���o)m��]Y��AIp��1��2MQ=���Z ��:ϟ7�;��A����"-hȠ>����*�a�����=��w�K3[�[]���5Pȋ�	���Q�Č|L�@��8B�U��* �n��ߖ��;���|����E^���on�� ʽS����AyrH �Mjg��O74�'��iODh�m���9�°�U]����֐�6��åi�'KBI�u���1�N�S�;����r�$�����E7kI��G�~XEkif�T�����{�H^+�1�_�D��=�mt�z��,n�-&Ǭ9%���B}Չ8*��rm���Ѹ�2�0��8�k^=�����C��:���u�û����[RB:���ծ��E��k�Y�V{{�@��}��>� ����&+�`��6�o��Z�T�D���׬�z��'�z;�֌`Zr�h%��A��?:�_����X���hR�"ݴ��t��V:�&@�Ip���Q�/K�e���n�;���oH���$���jd��3�i�'yM��ސ���%tҖ9�
��G���H��i���I����~(l*ߛ�6��b���p���^��_���>Q�� �x��9�r*{��9�S8n�ۀO���o��H���-!�3WKJ�ߦ��,l[6;�-)��,��޵�p7^�� �9h�h�4bF��tS��R����Q0֮��璘���UT%��?4��Q@�_2��k�����ͤo�l�H�_���o�hT��q޹D��g�������*��x�(?ۛ�$��UIasK�h�1_S^z�[��D~�u�F��`?k���7�u0`�8�����ˡ�&��t�8
�.�L��y�.� ���*6�_��V������"W�fTl�i�� �T>wl5��{���5�	�	)��褥�TCe�ӒǤx���V���Ӿ���d���e���>b�s���)Ԁ'n S�W㓮/�[i Y�)�}Cq�Z�԰*s��M��Sd�$�D�@h��J<��h��x�S��ґ����F��؝z^z�eۖ]}3AD� 0I�ݵϏ����`Ǡ��P��'���w���	_��N�$�����A!0
���4����0:���&@%�!(��QD��~e�Yg`JH-Z�ܭ6	Po�)_�^������V�\Bح�H�^�e��[�R�A��>b�����|e�>��
�;���pBs\�w��j��9ծ4�^D�C��+~F�Xu�|�	da�>Wx\�:(#saep9/A�x���S+Ѻ哯ʈ������H�����Ro��~���xևrϞ{S味_�xB#����;ޕO�Uq��}ͯ]o�-d����H�v����2U4�9�I	�g��;3��A��6���k�#n��@;�X~=�56�y����T�����g��(>�	p�O%�d��B���E�`ei3����y�|�����ݦ��Uygr>鼍F��9���!�"��ϳ�G��"���uVm���
>b�l�m��(���S$��nC�=Kڈ�4F��C|�K��a���Ȥh�G|.]��wF�͆�4����}��\� �p&1���`�6N�0!C\�k�����
?�l�cD�s���/4