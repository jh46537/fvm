��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�}`jV5	Ңf�G|.UTC��!U�Db��6Wr9���zZB��0/ūa��\d�LSp2ժ�R�mH����h+��Qߑ+��/o�,�il���̢�ڴ�����tY�+�6B4��B_����X�����;�=�>p�)�<N^�y�Rt���g�$��IYdqIl3����3�	�O�����
N[�SB܁�m�:�%g�-��j=�b�qN�zg�i�D���Q�u��=딋lX�'p %o�)׌h^.g11��dۄ뗒8�G-�a�$�|�I@�Cx��u]|K���ž�\9hs��uW��I���PuŌ�� ��sR\e��ϛ}��;q���vs��[��8y�;Z~8�
���@�iѣ�����o�^��������֛���jt��.r�?�_)�b:o�;�
�Ag����N���]�BB+l�$7��'e��·�o �0�1�XhJ� ���l73����%m�
���欷
��o4�~���[ly���3��oe0�,��d���t�u�
s�g��]�7C�5��]���r��;���Y�����q��H�m���C�0��6��;���ж�Y'��d��Y`<�&>�����%�-mE�E�T|�P\���X8�����ӟ�x?�!�:} bG!#E[��o��z=��:��Α�s� ����K
-�\-��j�m�ԲUk���.���M��N�G��X\���R�a�w�<(~E]F���& )~��z��s�g@m��o5��qyL�S>8�b���z[�8�nJ|��q  w���׳�%��2HR��N�'\-M�u����J�`�T|�³i�m �涞g�sų��iÄ�$����һ����Ֆ$H�@e�}V��t���c5��H���/�nH�%hoo֨��9��l�d�noF�sK�?�o���5��/�!�hӜV��	.9Z>��C8y:�=����@�4�����[ �q^�U��H�uFlc�ȫ�9�R<���#8�e�����{��G�����b �\���3���Ohͤ:RR�n`�#�@S>�a�����
�I���H#�nY�>
th��D���d�3G�z�RN�ɕ�������h=�H^؜�%��w!B��ޭ���j�&YA�nO]O����"��Bܳ� ��s�cP��yYy�{���D��2o7�_�ت��nYY�Si�,�d#Ă���>S�S)R"R띱{�O6D������(
��C���6�2Α2�xۂ'���R��:+�V�'�8��
o9��[6��h#�f�:��,�2�	�(�I�{0�vB��<�Q7�.f*����K%����ӲͶ���������u�;�e��C�7qW)r��Z�F
8���vn4�@#�4
 �5���m�|�9>��S.���zj`�v��%��sИG��HY�rݾVa�߼Вp`Q�25�-�<�Z�w'F�B�c��΄d���l+�`a�>5σ��� Iˇ�OUi0f��ܬ�t�`#�,�j)�����b3Ks�� ���K�Fk��R�ʺ�l�"��w�5 ��������=���0j"��P�:�@6�Q+֙�R��[L� �_o�8)a;�u��@�C�����7�(�wgw,��vA#9p��q�Iv�	p�[��%�ݏi����[��͈o	2#)z������a8!��h&G�w���Xf	L"D_t1�\T���B��ID��T,�������8t-P�W��L�ao|�����Ȯ����Q�-ૄu�|l��v����|�2N�gY�D8��lo,�|�6J����n��RN�D�#���ؽB.M���f�S�At^x@Ueή�v:�v�0¤���rK�gX񳭚�<�l�i��Z2���7Z�8�(���|ˤ�uX-b�|L��HER�X�!���>�j���o-�=fg����^s8�y;k����&���9��P�x�����0Z��\R|H���c�T%�\a��tP���N�5.�����>>�U���wл/W����!�3ѩ�%?58��2
�_���T��K؄����Y���ߴ;S��+�K*��n�_M"�&Q`-�8L�.����<dr@t}8U��)�pT�VOy~���!A��2��%"���Z0Y�|KQ�zG�u��9�e��}��.�	�(j?TOT{M�??V1i��hOm�?�pg����s5BH*_�mnj�9|Aj`�ؔ�������B�*'E~����5m�������y��H/��P8]����'��F�ӈ*��a^o7R��6
0ȋ�Ѵ��D={G�J�����*�qs��?�<d����R�%�qA~F
�{��o�K�+��f��a?R��{��9U�֙EM�f�T�i=�Q� qW�z}MB���-�w��j�k�AB�Zs]�[)�AZ��4UWj^�_wj� �ssh���#72X� ������H��MZG���	zx��\�,q<�H]�}Igݴt���rk��V=ݪ��Ò@ �+kV�/|#�SX���	ߘ��r�l8��f�Zރ���p��RC��f�1�؞O6Ϳ
e�l����A��{�������Y�{� �c!F���8.��,�|oO'Զ���&�r[F�I�Iaͭ�ږ�͗��&�J�(�*ϒ\�򻞌x�#'ל���o�Ǣo�%Α��þ%���3��
x�K)}�r�+qp
��6Q�����[:Z���fP�jH���5ب��o�_L�Yam�s��)ѐ�̻r��׃䡝�x��_0e�Q��� z&�
㎇�S��l�:���a�"���FA�w�E��l��W�
�3.'���$]B6���Y��PcGC�e��Q��OM2�U-�+K�~���-Rzk�B�Z��Ag"͡$˩�3��� �1b6�[0)�ƤK�a(�+q�8��WU��)���_�%�Ł�������	_�\WH!�	�SpY��/��x�A�*@�M������������	�~�{��NR��朩���L���������c��)�ÍR�(�S���a���2��G2��=!/��B�}.4�Eh�s",�h��K�&�����~�Ŝn��Nd�1�T����zzD�H?7X�̙���@&�7�d�;5@�nG�6ʢ�&2��/��;�.]�V�ZM�ŵi�:kA���d	���j��:�)�1țhG_ ����^��5��^`������׫�h��t[�&�7�-���XQzH0��JW���N8	�U��F"R�c��b���D�a�Z
���r��9����ű:?�7G;O���zː����#���5� '����l%�Us�<���&^�߮�D�0(z��Q��]�����hW�T��4�kI�F�:BމYx�t8Cu�M�������o��B�W�Jw�+ܩz�ҍ�-D@@��Gp���ί�/-:���N��$1T��m�4lsW_%�Z�̑{៉{�x/�8�Vb�Mʘ��E'��u��״&�yƁ�BHȋ\��~����l���b��X�X��2�t�Ke��Y��.����_[��W:�͑���1��5��ٛ�l�2���zO*/ �a�B�h����OY����x}"`�J TYnh��]&r����yȽX�皵�'�J���*�.�4�&���=Qp��M�ͣƳA(X/���J{Ո��S�,��>}5e�ǎ�f��Z����Ǻ��<ڑ`"g�#S[�4湜rA���%(؅cB#���vG�h�Y��|�d1��R�����1ۺ˾�T(띂��c�W X�A�S�甒���b>��L�J	�/+:�O�'���\��2��j3	� *"]��v��y�yk����r���`�B���M��ɝ���ƠS6U
�N(���N!��Z���g�0X�a�ڌ~������������*��� b���޻��L9rܹs���22T�&;�bfX����e�ܳ
%�~��ua����}�9�ʫ���m�`�9q����L��]��j�T���q���v@zy�Y��L���	���@�D��̺!��#{�9[��C���m��X25���L����E�G~*%|��U��fq����x�>�58Ƚ�T�#ܲjz�XXN�L�e�5cR��3��H@�$���O�C@'2�\"{ ?v�����uC�C��==@�2��>H���)��P�%ޟ��a�,��D�X�K��~�ZTP9DE�V���r�L������x
ו���E-��ǵ���o�"`^� .�`ڹ�/t�kS�3�l���*�땻BZ�����I&�F<��� \�$1-�?!V�jnY�U���^����9�*��F��Ė��q>뽹������ �V�[��P����ҝ%�޴�)ր�??��}10��/��FF%@��I�}�3�`$"�R߰�=�A�ZU%��ZH��&��k���gs����W�R�Z���O_-�.w�݄?�[zba�`Xz�O%sF%l�J=�"��Izq�8�jH���
�v�p`�z���?��Uˈ� � �pc�a�ˀ��ڀ0;E���fW*�@&&f�_�	���a�zN�m�0Bʹ�kub��YH�Rа����x%��]�d���:��#U�����]nk.���ؾ8 �TF�c�a���M�g�c<�j?�9]2<����O��'�q���৪>�XR�C��i"�'q�?����/gB/�M}��Ǡ���^7�+ِōA����ݾ��������
*Zj����.k�[�D����Ck�x�E�lr����)�%�,P�KX*<��n��h"��a�\���)�: �� �1nY=�q`��{�ܷ��N���\�eIa4����r�!�|�Q�j�(�$8�<��I��9��6tq'ي��̯w|O~7ngaX�\�Qt_�������4�0���Q��:�婔i��-�O��~�j>
��~e��)�q,!�+�R=���_��p�ф?@�a�c��c��F7�ׇg�Wx�&�N螚���_lY1�=�4��l�Òy�h#e�L�H��_|�����'����J��񴲨�"��<�췲H�
I����gDCP�39E��]���po��7gӭ� 9k��LmY7>�wKc���5��˳�c�l�k�)�^N�1��+J�J��qRZ��
��1/ѓ$��a	��2�
Z% ��{.��������@�O�����R3j.�v�u1��|8�)���f󆴷*�75�O��M�j���
�xG�|7q���Ђ�k�X<�/C{�]��ReP�eJ=k�U��;A�o�LB[/Ѩl�$H�U�V���|Y��M�z��� �;&�Ly���Q��xN)��� �[�~Mc�+Xl�h԰hi-��3��U|UH�6�wNe��6��M󳌏Gþ�'{�����C����&XGIG|ab/7ln���f��P�����jG��監��ѝ��W|����%�6j ��!���ڋ�
^��N����h1�S��6�{c^�x����˩����Q��s|CM���ڤ*�e�g��CO�h�}2%)#m�6��U��]	��ND�/�R��a������z�!o�٪i�Eq#����(	�^��F �S\�	���o��<�V����8��V�&���<YG�؛��e��x�ۀ¨�_��-���&w��ɪ�=;5���Ў��-i>BH	�影y�Ӝ��ׇ���q�{���bRb�5BgzP;��s0�c��m�������Cn��(���8�i�G�5W����=L�_���_�����?jV��H�R.��#)�]�
��s��Z�� �h��29�,��E�{d���/�u��F��RE�����Q�&z^b�ZVO�'��3�b�.�֗��Ew�6\�'RP����Wb3� �k(�N��Y}��t��1C��Yej�:3�"i��:�Z�E1bm�����_l�1`��i����%AC�DO����'���^G+�����$�%X��/�N��z�봷�sU�j�����ރ�����"����=���Gz��6����썒+������	otd[Y�Jw��(O��(؁��ևv*x��+�':���O�n4��C}��]�,��!���[��X
]-�=B�-O5M�艹{]�]��e���s찛[;�ZxO���ƿX�6���p��||��R�V�C\twz��*��V�<���e�ל�b�3��*P$l_��4m��"��2;F����g�)8���b�Q��g�+�~�܃H*��`��5XLGFYr���mY���7s�3�J�Wto�6�3}�ͳ�8Yu���4!~�?�l2��F�)�G��r'Sܓ���f;}� td����R�����KT�����E�/��C��E�^&&7��
��Ê_c��۳�o�
�+/�S��U��	�b�S j�mK�*K!vx�S����Noۢ��l���o�l�S+V��� ��j*����&XPN����xnx��E"�ҋ��u�HO�#���B¡#��;���%�u�|�d�N {�:�׵��L(7$e��]p�~{�74}��"q����;�a���By-?��H�����V�H2~�w~�,-{���(9�a/M�Oy��y�;� 8𡎶�G�C���|�P�g»0�Ĭ�d�X
Oq�ė���Or� YWLje�zK�;�$a�I1[.� ����I�(������+O�>K���A*ڻ�v��3YB���	`ⓢR8O"�Z|w����.��}j�?rZ��LFZ44r��*~<�I�z�����2��`b
oQ�$&��}Dq;�f���܋�'����&ږ�`@Lm��S�����'^�I�����Z��ѵ^��K	����o�����ochnH�?�%z��r��١v�A��t�!�+=/T�<���P7g �a����;����rAw��#rs::�!��%h�ưd+pߛ#y4:o����Vt�o`�7�H ��m9�g)w�۳��m���1cm�B��6��?��ݰ���ebL#���� ��d�ג�k���[l�?�#�����ݨ*(�oB��,�|��P���J�r0Z��o7K��z}�����tG�Iow�n2ъ���Ds�`��
��!UX��A�m��A���]����9�ڕ�Tv��E5��ǫ���F�T.,+���u9��F�k�s��:ͫ��'�U4orSr|D���LI���nw�)��?E4�|R!�}6�i��ߨnG��� ��x��׀�F�_����G�@����)-���@��l����/�&�;A6����?tfiCh�CQ
��Q�V��_�嗉�~0�{w��ᰄY��Ѵ��2*v�db601� n�(M��$�wI��1C�Ɗ�+�_�9�;�e05�a�T�������%��	��QVQD8�����l���
*�P胁{n{�=��Q�������:/ظ�U�>���f;��DgZg�ѻ=�h0�r��2o,��>�ة�x������<׭Lv5��줢b_E�P�;v*���D���{�H�f�̂�,I�!.�h�|��q����tQ���q����Bß�i�sJ����eKQ�Zk�>�U��T6RȄ���lK@��G14�`>w���V��K�<s�R���?R�	z����o������R�ў��CW"�9�/ܾ��v�	���V#݅�%��T��p�����yލ��sb���f�f�W:��	W��[\+���lq�d0�k�*���"q��5p�G#y96�C�R��2N�%���<K���BO˙�NP<A�Qm��޹��'�S�h:�1y��w?2QS����gI��v%1�*u��`�㡦��!/[��wp���?
�Db��w�\
��j�ꁪW�vtQ$����lׂK4�W�*J�u�:�m*�C���݈i��t���f�^j1N� ����fB_��h�J������πk%І�r&=����ӓO�N���<d:8�\Sp�Ϊ���C-�Ͼ���2[�Xg�cp�eL����-��qy��	�[8W��&�=�����PEZod������E��A|��O�n'$=�{Z�)]q%������Q� ���D�
���a;���J��`�&�u4P���H"��.�`QF���E�T	�s�.�3|����T�)?V	K�!z?/o-դ�Z���<�k�+pt�_#�y�8�TR�Fhfz
J���<��\V?��>�����~���`�o�gd�񣞿�}��Kv��b��e�Oʫ�p��%����x@.T/��˥xJ�6������d 	&�:�њsi�P1��<\��0��X��t�։�kQ�b�"-�@
�Ldv�ΐ��vT�rU�Ho���IG�-7]�T�?`AϠ?Ig���U[0����&����:Ο�{�ܒ���5�V�Wx����a�N����G2-ڧ����b��k�Ѿ�w�%d%�?gw��.b��J�;�Ku���T���J|�N�]��t����=3�P��4OHn�;ou��D�*�(=�΁x�l��N �fO?D�Wő���1�XdK�P�GL�ǋ�A\�����M�s���LK+�n��+�h9�na%G��E�"�f���<��i0 �Rded�"���2��_6P7� L�s\���,�gV����rY�$g^S]���ݮ3�ysY!"G���"�Mm��_�Hjض�s�/�C].2���7�����$�9�?q4����s#�_Q�*��Ф@)Y���$�*���!��*v�E��,�ٯjx��3���7!�/���%��P$E�fnP�����2�6&�s�O�n��}�d=��Vw��-��y���[E����3u~�\I��tC��z̘�����1+ō�z04s�e9�S�+�1��g�d���>O���kG%��$������h(J�k�ܼ'�%�xI����I)��j=S`��l?�)�,>K�h��LX�문˝����O����2���cf�˞qb���&&�oH��t|�h2i�r�"�Nh��i\�6��/v���h��[7l�Q2 �cy\���V�jK�+�u>��V}��lzY��y�*�ރ�"
�uSs�BI�"YŅ��ʩ#*_����\B���gj']H�v�����x�m�GC�'M��Ć�뭁{�M�HI�v��Gb�n."Uq����9e�"�7g���z�倧������_-e�Y}7K\	Sɮ�߷�aW�*�q�� n����O͔�EsT��6�iV2��ш/�>[ɛ�T< 3���.Y�j��sM?�l^_�e�θ�����*>�FI���"�(R�96�k�A.�V��2MA�)1�L����	_�T����Ux09�)��I�Sޭ�}ş&��7Jlq���k���@�4��]�����X�X�Շ�]�X�Rx�̭s�q���.�h~�U�](=���SHX��!�9.��A����<�Ԝ�~a19��h�sN�
ĺ��6g�O���b�{��3x5*"ގo��J-2�������Uy���ӳ�_G��i=k�I}ѩ���0e�L�j��������7S2T�k�7� 5ۖf��e� iF�O1�rIs�D7@��g����:��&�Or-�qnGL�仁�YJ-��m�ys������a@�3�D�qԶ ��Km���ߟ2S!�tb�6o����s�0E2s�]p	��AMG��j$u��=@�!�L��#�z�M�<cc��V �+�ZӜ�F�{��#0����g��m-�e�2��l]n$�F��!�mO��qӍr�9kB�������c�ւ��?o	�lF�V�Q��5�_?q���@X,$��{-Qb�
�ZPv�N$/���8���S��f�374x��oy�7�睃_��vu^������ȏn�xV�;�2f��9?���ڞ,6�T��.�t=���q��ky���pg7淸��țC�k��t�M��o��9CX�R��|�.E�o�Gx�4���7�&t��Z�t#8�3$�޵w$8ӄ�OG54�?4�.9��þ ��:��l�\�
�H���߂u(���k���b�m%o�[���b��$j*!f�z���=�TŜF�d�>]�1�z2*n�/�L��˕��ے�a<���4�l����#ҕ�?�}��Nߍp�)��<���^�ǚUl#��bGx#���J�ɓ�oAAI9�SNhC���6#�;��u�AQ�!�s۷`��E=�c�P���<p�"��z�qt�P-M���1ƙ[�:vt�Q� p.���lA�m��gX��@`��P7�t�5	:ٶyH6����Э]�!�a���L"�B]���}ig�*��ei�M�վU9 �\����bݺ��x�b�ٞ9p#��'5o	����ͥ��
g�p���Sy~��e~^}bY��U�_�޳�E��rNB�GE"�����T%�`�����3ﬤM<-$t��9��v�ގ^懝� �j�(��S���z7lYxe)���,3�������Kqec� 1E-��V�X5��u�!�u�Mָoz���Q *�%�Q#�ף	T'j-A�gь�m=�m����\���u�xo�6|�Z`KmV�d���/�ͳ���{�� 2W3��}�ԥ7�\�Rt��;�d�7�|t;�z�W�؆������5�GƆh=]��;�}%�-.y�f�^���m��f��m�}�q;�e�@���蓹f�i��HK�-�_��-���`7��;�
��Ч�}��A�S
c�i'��dֱd�-��#F���O���̑��� M
���ϘY�`.�m�R�#V���pKۈ����8;u�U�M����;���ȃ;�4WƧuZ�_�|������Kв!,�0C4^M�U��A�y����`,B#j|�>چ)����D�,�E|sU��ӆ�:`ן���;��%V��;5�v�	�l���x��?�>O��JNc�H�H��S�-��+(w���Ǹ�4�(���)�P�G����Ͽg���T���zJlRS��
�1	�f���ܕ�S?��䰸�i�F�>�h�M+I:}̵J,ތ�]�2�C�hK���A�6��BsC�
���\\�B�r�|��|r,GWBViy{���x S��3��8�d��4�.����,��;ָ��vG��ܗ7z�n~ƭAt���~���M�V<��_��*�
�>}�N�����#� [~����~Mu���4৛|��X¤�%�0��N���0��4Q��MS}����Z�����=�$S������+�V����y��^Zr)Z�^��(G����!}�-�d(���w��h�ߏ�~`��%g�]�	�>r�4ozt��!]��V����I�̭qv*A�,t*����V��9�%r������T��s	�A:�E��7���zn�=�wM�5pvHTB�ۨ�{.��o!�LeO����W9�:��>{�X�}ѩ�a�L�~$�7o/�k�9��\�=����,���V'"���6(QǾ�_Hz�&��*5���=^º���D4��;r��9Z<\ Gx��H,��膖/�@�k�/��)�-��0�j�2T�Et>�bK��1P�}��7U����.��v=�������0#h_Eժ�~<��xR�8�O`5��!$�dԛ��� �$gT�Pԯlj���5_��I��w$�bqk�G����)O �^j���G&a\��ߜ0���#Z�|3�n�C�x'ٲ��Z�kSE��ɕ]B:E�O�_���#Uà�=�95v s�R������`!Ώ.�s�g$Zϻ#��X ��8q����Xg��(/5�ؓ*�G�h�q-c��}�/�`L��&�&����#8����u�2��>�Z,0�.*6#O<�[R��=�c*������J�@*�e�_Q���TKd�4�=C.�%M��?9?�w7�P�)���Q���/�gx�u8U��:�va&����2�	�sU[M��@�I����V��I��C�f�<�Dm�dzw6�Y��ʨ����#7�ڬ�Q�)�]h��4Y�~������Z?`7�U�2�8Ei!�	>:'L*�VR�z�7����>���"Q�D+c ��P(N3]�v3�m�!{��l�8����D�!�o� J��
�'�?�rxQ�����is5����E���3��@��K���"G|&bQ�@ ��n	c��Q<��B5����Y��O�;�g-� ��� ywO�r��Be���i^�ƍ.�,�Zs����y�|�x��6�rd�� �Ńն��Kш��8�G7��i��Fa�5"�I*�T��Pp�q�v�ʖ�Q�7r���T��t,�×J�밧�.�(��딾=��x�n7z!��w �N�c[�}"�8k���f|3n��0;��PR�6���R�����/3�%А QgM� 4��N�t��4�����!Q�����S�5mc"�Q���o����X��Ƭ��:�
(�Ze���E�К�u��KF���L1_�Zv"P�Փ]W%,N�F�����:�d�@�)��.v)hf�8*x�߿��CYݤ�Ň)	��;H�/��E�]0GX0�,�_����V-�䚿�����b��j�u���q�6��P��C7b�ಧ�؞��������q���Y�2�]s��55���`]�Y/s�����<��} �,��c��yٵ�T|�Mɂ��7�k�F�\�[*�V�����n�g�5[B�R��M�/Bj�s7I��C"jo���Yd����S"G���l�d���w�e2��W���MΌ#�����Ͼ��� ,w������ �_$�����5�W�����(�ܞ94��u�Ϸ9G��VjSCk��OpT�T��<��2=�.t��4����պ��^�-9
l��"���f��[��s�_��9����9�F�R��D����u�4�N�+l�v��R-���ĉ�� ����5�p�嗹��=�����l�"Nl��������.wO��u�U�+�f����
�D������k<��BB �emZ�#j���]�L�����i���
��e���	��7�g&6|vݾ������w^C��� q�Q��z�Ok�2_�39|NF���-%ʮ�Lq��I\��$����&şsh;��5D�~^鮵�M��F&V��Dx:ow.w��jn�B̰iPH]��툡�����oln�$*Ss������ʸuċ
�-�=;���6z_C���g�C��f&)Jn�&�����0����:����f�򍔀8�m'=�B��JP�֔�y��y@6�����Ml�*�
��Q�4d��z�����~~W�n��}�޾Q{������9D��5Mk fHgP@�'8�����}���{�`��tg�����0~���V|"��o�<Z
�CB(�UҜV%��F�/�R]_���F��~��x�8MLi���4]5�#-f2�˛�V�-�A4bM��� �+�Xx���u�M��dzp�@�e�Iݘ�a�I�NQ�FOnb��e��*�[
�^M?� �P;��L��Xzf��1��Ǖ���^{�H9Ƕ�ߥǕ�P̏)i�XQ�l%��|��������2A�w�z��i�3#�"��z���b��SU�29��nF��t��}UMy{e0;���/��Q�U��x+S�6>`g(��R��Sڝ���J�HPxFR�݁hK�H���4�9���3	�@�귭y�]�ɿv��Fn�Tp�*|�m�>�@�ɯ�4�	�<��Y[g��-��H9�\ 0�[��N��+���Ա���$B��޻�E�"���|yg�� ��t��pN!�;ڴݣY9���e��Z��������I�ȸ;��N�L~����"W��Y1+���!�!��L�"Ѭ$�k��m��3|��{Q�s��FB<���j�Ӱ�ڋ&�Ph�p�J��t|3�'6ED��!y����At�������Fq����GNJ����[,�)�����6}�5w��v�.����'�jc�I朐��h�����c�����:^ 'ִ�ѝX֦�
��\Pb�r&Yc�V�=�d��D@��(��9U>�pכb8��m���;��E����8�z���>(��97n���-�L�]��5� �����#k;�w���?�I6ڀx��/���s>�>�z=�O�W���c�zNkͥ[��s%��ǧ?6	����E�N������G�d���:!���K:�AT{P�N�A�B�b��RT�{)a��ͧ��v"�)����}h6��V�:�+w�y ���1�~�L�A#q(�g��R�A���Fw]�Ѕ���(^�{k$�I���X�zr���7��r���7��b�� y��4ӡt ���P��0L��a�����鐦�V弭F��}�)���	b�Q�O�nQ�=����w�IfSҒR9�h{/
�֫���0�A��Q�*2��M<�"#�K0�?bb3;'�3��W�]���y_�@��B�?k��A� ��Yz:���B9�� ����f-9�ʱ*�R���~y�N��Ҧ���He�aI<�j��,���G�>R�D���z��ҳ��(e6-��0��_�Р��� ܀�ɕAs3�
\��
-{�h�/d��BhG�Ha	-*��W_d�-|y?����$H^φ���_����+ԧ!xΔ0�|���� �����L�d$Z�6#��fd�-[���moc�길"����;��T�hw��xd��Pp�ty�]���ػ�,%����?��d,.�Mk�9ܩ�1M�q:%�7��n�;�ִ��ܾk{_!�y����hV�?�ku��;�G��&24��
IwϾ?��1��
6�H��4�d����y/N�������Z!Xzc�X���%�(�sm� ��\`L:1Ձ+�i-���
@�nLeZb�l_;�Ɓ@�L�e��9' �t��'=�<<�����jY=�t��\A�唊����C� �l:X��֚��|���3��)]G{q�n�* �U�r$�y���/��������k��D@��(J�&$- q��Ft���˥2ʞ���%��"%�J./S�ˢ�֠Q_+����P}ٰ(��RJ���d�*�byr��	��C*V9H�0E�y�\Wx�/Ő���S	*���X�W�BV�����<�|�R���Z&�:�D��ʜ4�����=6K=����wA�`(<�.?�|�WN,�`�<�K�Y�����o0�����I�Ïs�C-3�������m�l��t����r�V���*� �:4�ci�|�,��u29�m�NMjϧ�-��n�%n��w����(k-v����]x��~�{�P"�#�nd{4�l���}t}��z9�d���9�\�)��-4 "�1G���p���F�Z�,�W�.��U쏹����x��(_�n���_���g�9S�>�+"2|7ܣ�H-���Y$6�(E��89b�2o����vv:�1���p"\7#���bq�yk���q�NLQ�OPD,�H`����bȑ�%�:�f���ޮ��6&�~�=+84G"Ɇ�����J�l�ԃ؍��F��˃Z�E7���R]t��V����)��9��Aŝ�0�80��B�N�f�T.���׍���/�ѢS�7u�5������2�Y���>{cΐ˼�lU�$��o�������Σ���#%%�h��z^|d�����Q�ڛ�z���q�/^	�2��
K��v����!1��5�('p��b�����Έ�}1��73������t��̟z}�Q���C >j�6J�K3�)���'�e[ǰ�n�+�u�%.l���r�zr�v���	�f#�P�{�5��������OR�qlc����4`�յڔ2�����6�Xqh��͟��U�
=��*�<��)._B��@�Q��z��bW��k̒���]$�b "3�T/fa�S使�Y�V?����.�g�	|W���[)�L�>i� �7(���ٔ�#�y���4UOiHg���׳��j��tqe�o�?���CЯ+�7؈+�Ό��Կ�d�(D]9����7P�x��� @�PbH�vm�&۔`�J��w�n��)��l�R{����X�ΨK|>.�^�$�D��6����9jgp=ё���Fk�cPu��������yRЮn!��bյ�-S����5B�2oz`>�a�Zv�*�评�H6ˇp�!e<(1��r�6GC��i�W�Ҥ�I�X=^u�5:6���Qq R��V=ߗg|=���J+�ur]�b�3���j@�9���K��d�N/n��z�]��I
��rRB}�O��GN_>���]�#�YdU/��q�N,;����=d�V��g�'.���3��"]~!���`�< ��`�
��`�ue��Rj� J3��b~�����{P_ϭe����E�.k�>h�Z(;�"�״�ӻg��_�_�ga���O>X��E5;G�����:Y:�G2���
,���)���i�Oi���v��g=�2H<��I�d=�z(��T����/i��`z��8�'q�iU���J�E̳tW�P9�����}�����v�P����:wo��[x�z?י,7�8�z�4B�x��d*C�"؍��v�۹B꯱M*�	nɸF	���L��v>m�ː����ҥY$d��#Fʊ먘��FuB���d!�����1 A�v�7����+��Հ���}�]��E�|�_x�����a?	A�����������R��Ѡb`�h�8 DB!|�7�EM�S{�'�v�b����?��9�!I !�綥��}����v~�Y�{ncx=�kq0Y,�/ V�u�>D���0���	ȇ��?��2�T\e�ymN�q�^�U���Y��Y�4F�8�P����0�#��r�D,��ŧ��D֖���]�+�
��⥬ȩ��_�P�EA��l����ufPx��&�Jz�U�$�'"�m
��9O1�K���'f��%z��]r2{2��s�����j��U�	�D����.3����IeP0K��f�Ma��g[`���Bsup�<�>aW��?{ʧ!�gw�g��w\�:�3*@�f7�����<N�­ީ��bFFA���:�~&`E���	y%�N�]��vȣu+�ϝ�T�S��7X�����a V�,[ oo��»��<5il)�ƾ�@a�E�2Qf�ϵJE.Z3�I�������h�m�̽�ӕ��J~X&1��zK߼�׬�*w^�-�h4��ֳ����Y%��������N�|��Cf�sZ�U�~/�Mʊ�;zZ���ظ�M��><_�a�E�&ߵ��*��BB#�����aS�z�K�^&�l*�\�S(�2�����Y������%h�	�:o���N';CG`	gB��ј&��T3�a����������I�=QCDS�Ztp*f3TC��{�c%��vfo�cӜ�Ƥ��O�dX< ���ew� ���΋���%����"��5����G�AT� uq�ChF���&���ܭ���޽zy�Y)痪N�g��H8[�`!�+U�%�t4�
2-F�a�?��
`�ڵ*�Ͽ��(�?w���F_It(�^�ɜp'��1yH���1o�$߃�_DZ��p����W{s��\Ox�`*W�ϊb(�`�[2����A�7'~\>	���<	���`?2�#Ǣ|pk��p��>�(l/|+��zn&������{��Dzt[��j��>Dx��w�+x�eMݔ�s~��Ki�gIJ"qJ��;��p+lȫ.�29h��{�PKT[��������|eڣ�Z�X8]�Oqmb���3����1l���Vm�o��Z�PW������w��	��8B���A�M�]�P�QK��M���-S��G������׷��������l��hC7���c���W�8랊u��Y���Rm#��)��ΒM�՜�ٵ��n��q:��/�ڷĺ��W��IY�05>Ɖ�p1�'�D���D��]b�&���PL��X/ �c���L=�Y��Te<]=�t~�sӴ��='�^8��"ߥI��ܤf��SDm�N;W�r�W4l_�v��}���X��gX�����>�	z��a5۾"�Zj��Ð �S������SCl��ǲ�@|oQ�@�KgnU��xT�N���R7�v��/$�+��৓����ܞ̏���p���J��y+��'(���k���e�Hvt&9��R	IMڛn�k���/��y��+'����4���yU�]p �g�%��S3n&e��HC��Eve'�������C0�܎����sI��X�	zKKt芓��c׌�_C���u
`�Ǯ����dz��Fշ���Z�욤���H4~��m��;�����B$�u�����\s����8x<��Ş�[�>���.�!����P3�7.��n5ת`�6	xni�S�
\?2�����>�	����f&+��99���,��!>V��ᙝ�ڞ�aM�|Dc6B����6IIWŞ��-��MD5������Z�E�-Lx�Ր��$Z����"�}P2�X1:%�j�SE�r��Fl*�IPV�V�����9�Z���)�f�˶�p��r�jl�A��=eH�S}o��.��
�H�t���M��2gc�ҽJ:�#k�������ZEu�zSӌ^L�؏19ۜa5��n�]ۈ���j���S˧��z��9jIj�-�*wg^��D��Ȃ1��g�@d���Y���Đ�m����i��/|���Wڵ�脂�\�w�N'����k���� ��TR>^���.����el7�_6t�(�h` D�&�������$W]c ��q���Z{D�?�њ�x��^��>,�q��Q܁��*�8���Y4if���#_��۱|�O@)[�5��ʳ�0cz�:��L'`��	+Z��z���)��D��l�.�-Բ)x�o���m�,D����a��+���[�y��i�w�/��Y�d��ɑ���ھwsZ\(����K�� 9�s�z�֏Z�劥g���xe؞��e���	{}�3��_� K�����
]�O��I��C�E�)$쯇��~�X��qE��������W��;GԈvM�Ĝq�G��T"�	F@�t¡q�o;�^a^iLa}��l�`5J����l�l�����*~�g�.�ae�E>�'^�����c���)��Խ9�ԋ(Z��x�sBW�8�D�$��-�B]P�f�Rmd�8抻b��yIl������<`�����L���Q@���~-�a�
�o���������d.iKgR�uIV�Ý�t����~���y3���U2rTϡ��=�_P}��'1�"a����cƏ�X���ZY����34�|^�%��3�k86��#9����A��Mc�>&|���3��k�?��#�������$
U�Q������Y4C��d��vY������^��?^�fP�Q�@�\*�jC��U�RG*�+��~���X?���Ox|�⁏�r���!9�^�oHF�/v2�؂͏�G� �>/m܎��>�����Iha����>lwr��PfQ]����NΜ��`o�(�N ��~'���"��B�Ɠ��u|i����D��
�����d����^�M���C��ۻ1+*�
L0�Z�x��	\�/՚��EG����;Oڼ}nÈ�2p�������9{nF��O{�a�抁��!�
�AH��tx�w�%� OsA�8Ӽ�� 3��{)�dR�����f���ߔAQ	������Q ��sI;y7�0vN	~6d���!?b���]��5K�L� ��в�,j�~T!����D��B�� ��)��I�����L)~r��Xۄ>hI��_L!v�<r&bu�2s��Nr��<�F:ė�
����'��+���IXX @ħ)4{Ht;NTN'w�苞�r��z���HE%�FL6�Ҹ^���ε�_���4��b�[tc���E�҉��"5l��m�*e[lX���6@��Wh��f��LM�i���^%,��'7�Ԍn�%⳿�tV��G�T?�;w�q�ȣ�ouó�#!�Ht���.7�!��,26�?��5Ȁ�L�B���<�An�.���)j��kiC%����_��}+(�Sr�ob0~ݠF ZRL���{��A�����āL5_�`�F�+k2��+�B�KaP��a�	�Xcr���*�Rj��k߹���M�"�|!���	^]�J0��-�tY���f#l,[G����Z�5FmI�X��j��r�^z����8P��Uy���/�L&����BOΝZ�K,?t̻�v����`��m���d�y�����c��xO��1Hx�2����N��y�sd��b�2��x��/�4J�w��6����`�o���*�7|[uѸ&�.����C�XS�����7h�c��X?mkwY��6�?�\o{d�y�0UA
ρ�(�cb%��s���c���7(@~ur�s���>~'*�Q(�G �`�9J8Ɣ��^U�XA,����)�q��cA�T�wi]����������ʪSl51E�p�K�0�M��o�)��?�DkH�1\�o�--|��n���F%�l{����p����_Y�>��>�9���ow��.������6��~f��&{:�%/n�yqhcO�T����~k5U�N�dh�?d�*G,��l�?��T_���)T�y�P�1|١׶9�ʭ�_�4z|#���?ׁ�s�/�[1��I1��yՌ0��EHܱ���Ab�������O�x}�+WPܴJַGI62�n�A�Y��Z�>���\[��N�S=����9I�]0@�+p�7��&���d
,�r`��s�� ���>��j��v��*j�4������W�M�7<�-�ף�=:��Yw������~K}�=�=�a�"��k����ڃ5���J�sӑ�d[��T.o.^�C{e:D�$�C2���-4�Z�
�h.K
��K�l8�?�t����g���+���y����c__�W48��ϗ�S�+u?����L�$ك�k_3o��q��� �y�w�1�4i�]i��& �;&9���S{9p�-�L-��C��Imt�eǐG/Y����>%d�t���C{�Gb��Ż�rN������oQ�y7]��D��3%PS��	(#����1~iEL!��ܺ0\޶�"\��b�V(@2�HS=v/K�cA@����R�zʟ��z�(]��7�V::�,Ȏ�a- E
��E�d��WK׫5�2#��O�wY�T�%���r�'n� ��k>�Om9N��ZD��;:d�fcjH$9�Јt�|�p<�����\	��89�t�
0�A8r�P�U��ե�kz=�f�\�^ش�IR��B�gH����V�h��R\�P�g��IO�`��a�6k�	����au��c5��jpx�(26����ԭ�K��5lf.h��s��7K��ltݪ@��1*���?�ጝ�S���0�ȸ�xW�(U��	�� �Vi�O��|�3�2&xgG�J�&��LJF�gC�o��ק�rp�U�� ���fE�2@#9�$��JuqR�<���>�\������q��]�{>t��1~J=���Ǥ�(�=
��3��Z�:����RɑK{L�������N��5㢑���X$�����ZB�Y�s�/��%�=�efO����	|�<��|f��m�M���2���3��d8�3�oQ,-Y�<����*Vب܄Oep6��UA$*��*�G���i��3��.�e\À�L�xtR�]u��������v���mh�ì�q �X� _�U%�5{ɧ5�Y�
��9t�zϮl�U�o�}�D]�>y5=WS×� g��.�H�[���h��`G�F�I o1lPA�$�t��&�汶ӆn$o�[�D5Te�d�,.�?_\0U?"�P�H��&�YX���%g7�)�����9 �	E[)
!Ď�!L%���GW�䚕��w.�������In���yYT�qC1�-�Xb���E��!9����䌰H��5bBi�9'7��?�6GO~%����[�����O�p�#+ ��"p��O��e��/z�Z�-�(h�/�������7�d��	�_`���*�k�����HOe��}	��`���M�K�3X8����{?�U���`L���=rT$����!�MvG��E�^��TW�}u���C�����&NKp��Fh�WA��b�_{�Fl�X̼��&UKo�����a���6�X�C&�'��տ��v���v&��%J����]�
	�v��*s�LV�ջK'�8m%��uj�[E��y�*eQxC��VS(�H��v�xn��eѮ��B'A1�w�LWz�ɋ���jZ�hnw��x���ct.`2��b&c2o�3�9.�t�ݟ_¥b��4��M1�]��!#d9���כ���� �r��mT��a\B��E`=�>��yEC��0AMV��Xƃ���G|S����hc?�[�V1�W&D��<���/ɏ<����wNw�SW�8��p��_+���̫�=�ӌҞ��,Ji�Nf�u�5ܝ0=8wÀ6�N�\/��f8��%�AkTkB%1@�H��bb�N���J���%�@��6�S�$��3rc-F=�$��9Y���y��ڿ]� ��[� k��B%���<+�/2v�ؑ��q���a�/������7��X��n�*� R��}ZS��B�K1r�n ¬�'��۰��C+�ji��9�W��T�1�"J_��y8e�[O3�*��s�i�C����r�	/aۿ�0��8 S��z*�7\|']�	�����~��{t)��|�~P q��m���8�V�=RQC���ҥ�;̀j���L���ӓ"I���}�._�3؟��p�5{D�9�3)jk��.W����x�o�������q��bZ���#��$�tf.�(��,}��*�j���.�j>�'��iyw�-�N��i����摧�f��U�[�jg�D�+�+�� kf#��/8�&�{�Wd�S�(y�)!� 22�"�����n�d�v����
;��&�(尃 d���&4(��b��3b1���j�^��"L������!��1���Uˌ@�/RqZ����7�)���镩z�B�~1Uz����s���"���a�ED{<d�,�8s�	�8׀&9޼Y��*;J�`�n��L��8�&���%x��;�b��vP��	|D�����������������%�٬�M�� ��ӫ���DC/7��֟�F
?��W]:�T"#��G�or�~��B�ϼ4��5�ڨX�8��{u�8������	�"ǯ���p�h_(~͋���Y�(4�U�h��E=6sGH�]G�N�@�.�4(��;��T^������M�� �t �������V�Jf���~_�Q�͊.��C�t I8�W�j�E���(�a�aˠ�̣��T����\1Y]�����&�����怱���,�F�ɭ\��c���S��V����������ǲ'�xF�#�����dJ�)l�I�8�Sh�����ē��H�!��0����u��)4)����SPtҜ����v�z��[u�@E�i][�!�9I�N����V9�~�|�7�:��%I�ɹ,85.QH|礸c�+ܽV;s)�J�c�W��+�n�E�X|����b�zy�h����a�ु�a�X�2\z�+O
v�f�-��iU�]�.r�F�	-�R�@�?��$ڡ�����v�eXv�݂@Cz>�iws�����iU�@
�xp6@�I��(ͳ���^�=qgHa�UA����~Q][V��m��aܷ�߁L��$�]���4$�z�Uh���Y�\�N��5�$���yw\��"~�*){�!['</N��]|'fsV�V�ɹ�q���z�R)ۻ��Y���̝�l#�Y�U��v���O����̈����n)�����0UCi��ʢ�������F:K&�u�6��3�A����i�P����b�2�Cz������z;�Mk���f��Wc�.�-�i6�o�4�`�"OX5��7}��Oר�'�6��>����5���$�"�A���ah����Ě�<�:9m�0��5�z��|�ir�K[��TQ~h�	P�(V'>��ܕ���|�eޙ� ���8�6��[+(���2Yƃ�" O���^�.-:J���K�`u��d���v*�;�p�d���w�b)n���b_"�ZC��_{Z�a�<�Ҧ~�J:�/6���������-ءzמ��Y��B{�sB(C���10z����0(G+Q5�v�&os���e7#ͪ�l�\e��dS����]WN¬F���̟��2��rx�GE�j�I��e�����bL���ի�<aLB�fHP#��.j�8lŧ7������x��''�n͞�͡v�פmŘ�Ui�u�H� :S���3��gaI�?Í�]9���:튈kw����F�2@xb�I�̉����T�P���PB�#��#k�����&�tx$���Mb���nq��<��Ɍ�4��u=��� :������V�9VS�8���R
\D{y�m����e���!��a
`�D='�5�}�{���Vx0��/�����0����I/Q������2�F'��<��:4��A��`v�=�MD�K����A��R@䩳e�D��ی[�P�;�X�c6��Bx�%�%G�����k����1xc����ю�|�v���|���\% by��3�N�(7v���t1Ԉ��ÁLI�$��yL�����;��ؗ��ғȤ��w�-Q�ף*��Ζ��ء�3+�G��ya:��+glW@w,�T�cjf|�h+��h�LzNf�{�]_V��/nƎ^Q���+i�DF�A��g
�.��/��\��y�*�������ڠ�)�� ��C���_bLH`��cL�k��.��7e�������[���C?���{S����� �|̔�I��rR&P�x!��?�ȴ*�kfz;�2���V�o���=�i��So�C½���3Am��
>���>x������㴭���컾�����g�{*ϖv�1�X>u���a�3נq૧h�&�=�fN���YPb���?3)x=��3��X��D�e�v/6[����F������o����>
5���+;
2���U������Y�؃sn�)R�[k�L�p����J���X۰x�>�c�4�J1P�<'�1�hd�K�-��Żم���T�����\�TO�������J-*��_��±�qb�� \i)�,e]����<��!�3���/į��g�����KG� �	V�S2z�^�z���s87��I��L��GI0X���w��ą7*�Cge5 ��%`����H�2%iśD�7Ɛ�ڣs�56���&Go�g�q3�t��M����\AR����!�X�m�KϠ.d��m�bv���1���@p�U�>�2���h+�O��mݻ��¾w�
c�K#t����+�N�p4�� y�ha$Q����5{5ޱ�{�пǧ�<���A��T�:PR�]��2�y2��x|
���k��~����iH���I������jPF���l��?'�⡗�>,�i�!�N�a�`;� �Pv�r�Iբ�r��0�~0�]��������ϰ�����6`���Ru�G8����ˉ�g13��I��?
�H�ՀJZsor�ġ�P�����G*����H� � u�H�3y�i@p����.f�� Ƶ��}����k�>"�F�N'ϥaVAz�*8�H ���7d�R��C��*�ȑٜ���<2o�_���JCu����8����Os@�* M|��O�I�52��#�:cOe���}yD�[lw ����3�0&�?R�b���P�����~����ӶL�(�0R���Φe��r�.Q�SQ� �ݤkj�J^�>���}͙��6�A���@��5���q���ޢ*ۥR��^�9xXUF�2�Ӻ���&�5����%)!��hrfJl���A#$�C����?Vُf�sW��-Tf7���V��Rc����ܗ1Sez�̐��t2�=w!�f�]JmGxĘ���P�� ��W�Y݂'E�l�F�s�:�,��6F���!Mk��B��w���R��d���@�XϺIa_Я3�5�BF��*���#��7�����Ppu&Z�$D�ߞ���F���I�����^+���?�8y�1����vl!{�|ڻ�E���e��N��6��hL��.C�IF/I�~��!
�x7��c(���e�Ch-�g����M~��~�0�H,����LW���*c��Z����Y��0S�cQ�t�h�����������Z���uc� �G�wn����[��V�T��K�$�f0��8۸3���}Y�n��z s�:g�H�
V7����
��H}<F�dL�Y�d��Fw�[B���^4�E�-�w�lMء�'5'��M����;�#���5�+<ER%�������� [��,!�F��e}�g,������*<ݞev�qz�PPAW�4:3R<y�8�V��h�R�}�C�� Z�.��KN�w���l܈��rOemn��oH��=*�xa�����9Oh��ׁ�Į*����^�"��s��ӴD����A,�X�L&"������n���݋0��z�Z�������h�^*��uq	80f/�{��-n,�����چ���*U6ql���X.�=��)(���<�B��Xm��!Q�io�9e�Xb�s�+�1����מ�\9<d�[��f�Xx|������)������k�[��I����
�f�?�+L��'�"�q�
2L����,�5ǾA�i�z�p�)0�fd����OF���?��Yp�eyV��	�ܦ��mb�4��Y|���_��x�rTTb&�Tc����{DO�S����>����y�*ŭ�#����¬��|�{a��!"?"�sQ��</M��r7��¶������O��A��[�Hil�GwP����E�`0��Q�o�`������c�-Jk��tJ�y��5�=���:Oi�s�6r�9���?����qPc����a}+��%륶b���+����)ږ�I�K\)=�|pт���}��?� (��|��#G#��x3(�I5���-���������C$w���JQd� �g8X�X�-�u�h&���jwx��k���q����{����'A�{�b
0mMw.�������7m��]/������Ã?ﮦ�M���kj���}\��hZtI@_�u���G�u;m�Hr�t���{� Ρ[�j ���P,�5e���ot1e�7����?��*�����v�q4�*��:<��*,����$�{��Y��قe���D�;W�C��횕]n�Č���Xf�n�\���zS*��'�e��<��FY�}�[��[�S�E�Y��*�k9HS?�.o-ȁ!�)�I.=���b��������9u�ܤ
}ù*�XB�k�����~9 Ccu>]Z7B�����N>����G�q�p��hYSe�~6�aG_&��e�Y*d��O�+��^+Ml@�����OQt�������䯞
h���Z�����le�9�n$���6@����mѓ) �|��I2�>�7�������B���J�
��G7�@���w��7�(�]iT�l�?�3��@���������l90��TH��P���`p��ݾ��5�.#˷Z����}��pSӬ),�a]�nz N��9�F��T�n
�����2+t���$o�C�-yP�J���Z�=�[���q�^ʴ)/�e����=��+���b�0�e����׫���c�Fg)��#�2��[x��S�A4�*�!\,f��^�̉._J��O�p��l	,HC{!ni��D���MTY��X!�:��	���\�:	�54cf~���V���������u�/���o�����5����RP i^�W+eɌ~y8[T���g�mGʌ����%96��R�2V�(?6��P��=<8&��?�Y����2����<-���f�)�V����|���֒e�`3e\�椸B�ÄAۑgآ����i����˖�Z1�������UqxM�Q'�q����K�7�B�*�K/Ÿ`smB���F<����A�!�}dN�\q+d���^����~��a[��*IfR8�S��a��~uWCR��, �c+~SDF�.k�&ql��h�'�|/Ĥ�:���^�0�j$XQ�.9�"�%����3*$˖��c�Մ-��O�`�*��}\��
���	� J�ý����{b	:����<T���3�����f}9i�-GE�����+��M�P֜���'��2��̞��� -!����{����!r���R_Dֽt��p���U� >r:8F�X�$q��,�K7/B�'�W�s9u�:�/�j�s�h..,���i`��םr�2�f�@s
��M[JP����:G�F�%��iB3.�FJ�'���aKC�KZ�B�*�q�)<'"�1)���:�?=�v�jz�I����-��k��?h3�`s� �r�����p�Zq#!Vao!���o\\��1}�*�/�#���-��`'xn�+.t� ���JD��ӆK�s�Lk;�X�\*��7�8�&�=�R��:@Xt�c��50Y���ܾzi3�X�jJ^O�mt&]���Y,�U�y��-��$�����c2{K���sν)F�=�T�RJa»��b��k��ɇU���U�I�q�h�8��N�9jLs��96[��Kb��u��{��M���2� �K%w�T���봋�9}2Mg�����6��˘a��q �ԑN����#J~�GIC(�T������ﲉ��m+�e�b�\��U;o�u$�?��Dte�C,���Ae�@5R_s���3���yQY��:��A�������w�2��]��͎��)b&N��ݡ�\(��Wo)hA��L؅{���g�Wu����	7�+�QE6Oi����T��T�x��ᰗ��Z���l���UdJ����2�ee�a�]��.�� Ь�u�ڔn�@��;$eQ���"v��g�F��1��@�φ�-9/ �d%T���� �0�)�h*;���49��h}��z�W1��S����@i2ϱ�9�&0ή7���1	��*ð�up���c� �0fa���#�WH�"�	 *yo8��!�X�����yU`�u�ŭM����7�wG�I�ᅟ&O^��A\>������v=�"����W�6�������:}�d� 췃��T���ib��!s�\4�w=[��=��:����ȯ�=	q+U���&��G�L����5�b �g�J�,�
�`M��C���&�ȶg���kv��8�2E�d�:#q ��: �C�}i�ކ ����:Ϧ����v���y��t[���S�0���_�Q�l�H���i>CD+\��2\�����w�X �;c:=��=�Y3t]���u|�C�d����ԬN%)_UJb`�[)Yqç�i]�=y�?��� (%�5R$�@���S�>T&@��j�1���O�ň�� ;�,�a��z�Q�a\o�A��򻧵�WA�F=�8��=,3�i�D�~��3��7C�v���A���u�9x $W�|`z�x	�Rk�mp��� �w���}B�^�5����z��8��ba���e˹Vȍl��A[�L�U�v� ��$��.PuG#��q�#�w��$$�����m�џ�Xf=�>Bd��'���5��G�?!�]�c����}Q��L3�����ɩl �x�9g��;�wP^��A���4*Ei��e���Z�Ė�ueKc�7j�FA^��_���L�Q�?Z�FO;�B��k�m�S���2bꐜ@�"��S�4U�ǒ�o�B�yĄ{��U�K�;!rz�1�bv��h����0g�����qC��ζ�@�?Ռj�R��dW�W3�X{.6Q;^E�`�.�B@�4�������'{n �G�(�7���0�s7�l�<D�p�U������`����Q3��?�B�4m�\��k7�GWFF^	I��Y����IiLT�g2{�X���*�Q���U�U%�3��������$��*���`������=�n�L�9������
�j�a��Ep���$�zY��o��N�%3��	j�y���&=<p�B[3|�5�N�i�뭥=��8��R��j�h/����5���rq�9V5��K��A��$�����珖LR����ՈCqu���]�c}��]ƌ��~�/�2/��>��q�����Nj>��/[h���	L�D�����9�[�v3��t�ݛ:x��]�X�f┓F�,���S8��U�[�y��=V��*�5�����++�-S�ԭ-zB��H�g���%���[Ui�t���7��#���bж�UD{x��s�z&�|����W���������е��I�>���
{����q���/:�\��.:<����hs�:��c��?���?U�U����R�`�, <cy��#�T��+k�z�����%t/�S��fnЩ�Ǫ����R��Ϯ��Ɛ��Rh����F���*���7� 9W;�s��ǻ�G(~�^�[��8�N��|D�B\h0$I<?���`�C	]�����h�<��8Q���f"���]g<�Q8m�mK�W��ne4V�΅�M���r�2�*3����L�?	���4�[��f�w�^�#��$#�$��uϥh�S��4q�bV|�_t�B�'��
�%��J�y�!��Q��u���&�I������������d�||S�����!W��Pk�1�A��D���Vo�:�%I���qA(�"��gS)��2h8)�`�1c	æY$��@"z8?`o9�L|������nc��D{��M�@����G��#_�s;8h��rƬ֭�|Ĥeza�U(��t�x� lU�D
��.15��ej'3��y���g��1sf`L*��p0/���!0���>i�x0���#h''��>�h�Ȱ��=^2ޠ=�֏[@Gt�t�TwSb�a�#gI[��IElX<���ɭ����arX��Z��[�#�;�ypj��',�y�zöB~��fWs:#
��b�e��Q��WTl�L�k�_A��jЇx;�Q�oXP���o�p���ͷ���7[���n��� 9,$5��E�退f�9s�9j*E��RoD̓���|i��Kp�#��� D�%8'����*�}�{r�oR(�c�d l�7�����X�U��/(>��"��scoF!i�Y9�,���鼈�H�ɋ���%�'�և!���yy|	��f�/�z.`�$D�SG���W�Y�eW�F�b$��=Z�o^��#ü͡B>�Q�?1W��l菉�3���h�}��8׬�P����|�F��
ws�Ge.L�7���ɣ���
��hkK�%����9���,�%݆��c~4�d�x��6���W�ͅ4�F����'��r�8Μj�R d�����ʬT��ǰpH�H
����/�]ĸW;�/o��u��f=����R����+�+a=�z�,����J29k��t�Ġ��K�2�"Mx��j�ȣ�!d��5����G8H��W1U����٦vJ<�K�.�z�Ϊ���HH�xX����$R7r��ǔؓ�x�W��^}E�_p)����ġ�=��bx�m$���F�r�q1�}!�zx�Ԝ�p��᱅���B*{�qs��
����m��Í4/�Y1��m'r���P�/~���ޟ@1�[�K�Dꝱk�L*�I�A%�ދ�}��!gE�6@0�9kG�(ǝ2��AY�)��:�	�I�yI������
��4!��wh�ҟF����	#/��m8�c±ɔ��_8|�a�(�am����JQK����yi�a�!�r� ����l��9¡kٽ
�
��j���F>�Ë��	�`M5�U��T�x�\��A��^2�o�s3��l_�B�3Fw��ٮ���{i,P���p[!�GKhI>�-4뒍��a}��� �A��� ���fN�Bܾ��ι�H*_+^���oU��ϋ��-������5�G�>��:�&�\\}X�Ex�F�t�A���p�G���UMV�!�HJ4ˀ�d s���.��vs��2 D�_�=OH���nU�ya@��$�ؿ��MO��!̮; g>Ð�a �W��o^����	ne��MN�,� �?�G�0:ETh�Tß`��(U��u$nw.˓ѧԂ��cR&�iVw�l�	��n����hf	!����J�{+�i-�qx�%�q�H�(!��>Z&�}�M��/�'gr��� �s�Z
�+0x�O���>�K` 
H�D0(cw��);3Ah��<e}��G�}�ʟI���񁕁.υ@�D}������oHU�
ro-߅����tۧ⾘_0���as�V��P�_������������7�p~ "۔�Lt��[io�����6�lkϪ�[JP6��T�2ᅲ����:��F&0F�2S&��R3Ӡ�S��P)e�L��C$�qa}ق���!���#,)��9@��XAu�~�,`��)Ӈ?�s��c]y�U���9�^Ԃ�-!��q ����Pˢ/g�`ː�t���l�}�]!2�&>$n�7�;e�*�u+$���(o�V#[Ǐ$��V��V�*�y�K��Go��Z1\r��� ���}p��8�i|�g>^#���@�:���=��N~�s��ܯeIa���F��e��G�y4
��t�����G�˭��~�'�|C��d#��|�W�?�����c��&���O �3�1��5gV^�J�@������T���M�4�N6T����@��]P��Ѽ\�!��d0�2�炢>�B�S(lܘ�u�<իs�6����Eq���3���Gy�>iW��>�{M��~�Rt���8�
���}�nP@q@FTeVOD���0˵@|���Y#�G>�5�R��q}�vr�8%}j�_u!�p*���Cg�z60$��Z#+��p(��R�(��;��H�˹|�D]�.�0^ke�)��v��L:'�su����ɦ6�ܽ��`o�1�@��5U��%J�Q�`��F�����(���=��S�dn�}j�V���Tb�4���k%���o�"�{���$ި����2�Y��Kr7 ��#p� L� s�9���e������\e�F*>F��^�f�֖�R����^��lU�֊�������5�}�y:��r���L��c:>U��AH�,�#m���C����ǝj)r*F7r$0T~�qT��n0��i��UA��5Aw�Q`�/:��߇�X 42��_�+I�J��F��+�B>��>��n��8$$�u���"ŭ
l���?���C��~rRDZd1 B)�?�#(��<���A�Kv^p|�{Ħ�7�I����^p��!V�����P~�������9�#6�)&�e��tQBS���戴��z��/��Ȣ�~�X��n�_�]Ŗ�#@���&�����eEz�w�����~2vy?o5�W
A�@b-	U����D�f�K����:�mkN���G#��������C�c��SN)eكB�d���_��U$��<9�8�8Na-R�!%Ll��+/`�`ĲV��(̯�Ow"�g�ꝏ��|D@�¼��urY�p� ��2a��ʧ�Z��)��W�L>�Φ��狟�I'��\����Z��̠�'�l�=p=�8�C�L;���5wڍx�G&�7}A?��ƃyl�xW����x� Z�"�!�'«���O���VLb �ԑg#�Jd����f1C����:��H��g�8Ѷ�i5���X|��d]ŰIj:��y36ȝb+�~%Kk�m�Jc�9������(���-`f#6"JkN�8��X�C~[f2��P�[�="}� P��'��T���Y��S�ZQL��K�3�b�t����a�51�����T�c5z�N�c`���kgz
bA������rUAp��a$9Z�*5*��C�U�� �ջ~���L*ߝ빝	F�+�T���=#t�"��`��(h���=:X"ێ��z$_�oI�� ��۽
[��	8π��,��������gX��s`�5_��NP��<Xt.<��k�i��7���f�ܷ��Ԩ؞l]]j��F�(%`2e�s��ɺ�(��apE��,R;��#)�����%(m����;�qb�|=�2�-+Nl>�=YZ��H�B�Utc��X��Aݚ!T�^�z���q�A��mtS�Vk.I�ӊ�(�M)R�b��L�_hYW��b��$�U`�>q�@ƀx(ċˑEp���;�H�I�T~
.B5Z����yõ�i�H�QW�>ՐI�G��kd��淜յ�P]=�mף�s��=����[C@��S�ן�������>�3�D*\d՗&���H�X	�f��-Я�����f�ps�= �ܘށW.ٮ���4? DķH%���s҅��3���3��V�*��ߢK�H=�5om�z�<��4�`��H�v��ke�Y����IV))UU�O^@�Nh�G���5�7��C�:*ڗu��N	ʑ-|��>�i���deB� �����$\���ɬm%t�лa�f����:�e��^U��M���{_���~��8EPU��G~U��A��J`h��� ��#���������v�n=X�7~&��eU'��G)U�(��"�Ւ����BJ\M���"4	#�V�� �kd�N��gV��B�Ĥ%��ݩA���Lk�R˥�|��ん1��@s'ZGDR�r�l�c�۵iv�d1��;�,��@�sf������uZ��� u�؁�%��]x��{P肒��(dE���� 逤ʙ��ĸ�l��o�w��sk�rw���.�F��As�^ܗ�E'=�(�sG��zj1.T99��3w!��	[H�#�W3
x��Q_g6�Z���X�'�[(����H��("RDS�8ls:����"�|�qy�_T��[�^�x���\�ߗ��2��Q{��ㆥ(��a�'`�R.� Y�vl̆���퀴h�8V\�E_�+���E$y�Tx`�"W:�;
b��������Y�A�ǯ�o�5Gl	)CZ>36��e<jl�ש�߭n^(�2N�.��$�V\�3å�����״A��,���֚��:MX��b;kB�M;XIP-�a>�@��e��z�ӊ�"�sf�L�}�|'���w���=J�t�_�q8�ś	���L_4A�����	'����W�l5�Y/Ȗ�Ћ[��wv�U�F�U�vjأ"qK3�����7@'�K��]���QH�b�w;�t�oz�]�Z�g ��Ti��mo���]�M�q�#D{ZMK�[T$=&�n�c<�|m�=?�	�7��2S{\&��O�K"LGӦo�^]1A�G���r�9�pO� ��`����k��*���Y\�*�=�r���m����Js��TDU�C�tqWq�X��$����'w�$ w�cWŪ��id������=�Ey� z���"tR�@�@�b�/�VԴ7�\���������FU�g��268��D^EZ�yP���E�sR�ޣ0b-��e�3vY�S�z��c�V�0Kx���B|�q"�6�M=�/V|큙��Jqz['�#�>�KZ�F�v$	����n��4� z#ZQH���[߸d��l%ᳵ2���8��,�"�&:v�1X�|rL�,<�m[X�S�s��^�"j�Ɇ� L8,�
�Y|�W	e�g�3_�����^�U��GELHt��=g��O�hn�I�b ڃ�E�I�d�iN�S��G�pc2&��m���`���<�UY����)ҘS=x�v����P�}�e5VwF��x�qA��ɾ;�;���md"�{s}�ޏN��9b��)�+����"`�!>���.��s�Nup I���v����-�-X	K���B������Z
������aV�I]U��2K�<��r���^�V�2�Ř<�U#���2 ͪ�Ӳw^�q��sԎ���%�T���,�)L�*�	�ż*#:n��:��$���踩m_&1DR�G�n�������>j,���	�԰�P�mO�o�>���Z.��R�2އ�$�{��5(�������%�c� ͪjp�]����}���rE^sqPK Y�~��ą8�C�r�X�c:E���&F�E1e�/�fS����=S�Ř�3�������g%���[���O5���޳0�
����N�E��͸	����U�$Q&�r9ᜩ�0��������mtq���i�BT1��Sy�쁌�
n��cD:ĝ?�0��D�~%%h���kS��$�ձ�7u~��Q��|؂d&��.��
�Ž����Ca�ASe��ȋ�ʣg���/l�����Ɣ0�U'QEN䎘-#�+V�k ��1:&P �g%D��o���\���ౠ�ǑӨK ��ƌ��殳ATD���^
L�_X�Ď�s��̨��n	�@��K$ǀ�i=Cd�}<�3�GD�ƕ�RK��&% 3WX���,b]a $׮�Sł,֡*��9J3��x��󤺙�$��k�B�=X�� �c�`����5R����o�ލ+�I��!�9��ƙ?Nq������E�� )nZ9�fG6��&��s���a�?�2�D�S��='ێ�:V(*��k�� �ɩ@�L���Q�B���'+�A�������O�3�Lk2Szt��O�p��XژX@��׺4���� (�|�����~�`���P=���2pQ(��K�����wA��Yo9x��0��)�@b,h�S��&���-����i������l�=!cq�P���U�5і%�=�����K���v�Ww}���=�Yh�;�ČV�E�2#L!��K7"��/ަ�P�p��	�YcH5ܽ
����d�g�8޼"�' q�
�l��:?��׶�d5��?��N��r������G��n�^!q�G6W%M g�����.���'h�+,�o�	g~�7��ϱc�Ro�(r'������=_��R��N�`[�.k���_�� _�īr�i������;qsY�gA, �BX^�P��  ���]f�)2���Vgz��\����Ρ>ڧC����{��w�R�T��9=���F�fM/$	��Y��������RU��q>E�6r���5���bN���8�UA|p���}��p�&�_����Y�<:�S`�O�w����o��r��(�M�y�A7� L���Pc�����,k�P=ߚn,��0��.+8�ol%���t�ȴ����|{$�����s��u��0	�����r�%�K�������bM
)_��p�~��0?O��ǧ�[���[�z�X��G�\1gb9�\�A�QPr� ����2��B�f[�����V,hH`��bk�tr���Ö)L>���LT_׆��w�c����T�K�Ջ[df�o��k�gs��'��B7?��:����*@'���ﷇ�����,�{ɪrS�i\�wO�1�uL4+e������ͩZ�sp�ю���\�~%5�Z0�$4q%v4%��DK��K
�C'��U�coERۏ�h�ZiJ%�?���C���	�����i���V�Y�y�*1� ЧvN���/�����b�ɷ6U\r���C�lo#g�.$�}��wH���y�ҫ�O+����Y����7���1�����v�/>jM�]t$�D�޳���ˍp
�H��8�;�2I�՝_z �̸G[&�	j�^�uPT��0BK��PO�	[AsYyS����O�j�9��f���JchG�P~l�*Z�lz�,�����ᩬ+Z��<g��0�+�&�p�f/��j��mM~������5W�0�}��݌�羞��	1*\��!W�o���8fiо�w�t^����&s��J��ԓվV
������=\��}��J���������t��}HA ��V��VEH&�[/VX�� �qNC�_Nޒ�t@B�g-�Ԛ��οj��<�=	R���9.��d]kkR�5l.�������
�0�����--zx0�(�d/n���D����3��}&��
w���aڼ 鸁+�ƿ����Dl��	s$�"�����L�q��D<�����'�y��3+�M�b��!ff�����9O;�汮��'fk� 
���x����D��yޮ�K��v�_0x�!]Y� �Ѱ��q�4#V��0U�q��C��,���fe�ARGf�ʾ1�iZ��')CG�9�(�V�ً��xg�a�]�^�@
���=�~������m>)���ZaNgݣz
0�꜂t�{���Gvm6��ۢ�<�1[��UY�e� �<I�{ �A�����ӲT�����M����Uj��0��+��=��љ}s�kұ�o��������w�f}���|�r/�m��Y7��Z{ى�J-2�����'}� ���Z����"S+ܩ���lG��iW�<4[�\��Ic\'a��?���X��̷���ҿPs��LPNa��g�,���ēHh���̉v)cPeZa<�'gƆE�U�c�]ڹ涏:���3lc���0������ 1�?_`^U2�bö��Z��h(�9�!%2��W�Q�w�������]�d���!��A�K~C/b沴�礸d���b��iu���ؑ�:/h(��\n�k۱�x��?��w���t;�s�c]�N�j+�t�Ff] ���
UJ]��ՑX\����u|C�h����]���Ǫ��׻�� �Ntb��/��G�����b>^w/Yg�E,�4�=��6�v�ᆉM����n|�Zcg�Ej�(�x�vx���4
���B��]�=r#\4��X)ۜj�j����g��r�<�7?�㓧��%/F$�TZt�����{�p�戁x�;���Rz������ Uڃ����?m\�
�I��V_&��ۺ#��1��_��]�[���k�� XoX�7d���Y!/t�7c��c*.�2+K�Ch�<���_0-��<({�_��.�/���Q z�o���Dnդ9��s޻�SYUZ�]p�w��]�'������	!ox��i��ٰ�\�5T8�h����'��X��_�Bk
�O�.5����'���Ѱ�8�ޡ�����
h����C�Y���0��Gʻ�B��U���[ �����+�Aӌm���@�1�kt�[���=�0��W|��ԂV��u��.��niӧ���m�gjd�r�eм賧7j�̪�8If�M�	�V�x�����և�,����K��6��g�����q_5�ZҜk����_�&E�=A�i�f�׵yJ���l��o�N�>����X�\��na&��3�m���E�v(�hf�f6�\�2l�C�>�
#.��O��Y�(i��K����]db�A8�����}zNǊ|ict�ex�n+���s��������U
���L�"n��zM���O�uJm�&=��>F����i~�����KL������?e�3����^?�Q�4j��)i;�<R�4��}G�K�a�(�#���K�.��t�=^)�ap�g�VX�Z��N��O�:��V@'1�s����VRњb��@{NE{�G%�t�tJ��;�g�,@#3�W�$�|���i�9�e���|�`���֚�⑱ԅS���w�G[�_��	H%��)�!�m:ݹ��G+L�������0�z��q0:�PEx�*��==:���MĿV'��b�Ϻ�ɩ���clM|\�}���[|#���%�%hy��U3>gW��q�4���-(ե�J�H��ԃ����Ie��*�,�J L�٘\�W�M�tK���Н�W��w�,r_%<�6`1�u��W1͌6��$[�zuJ���/jZ��)��|$Ū�4:}4��yP����v��n�!�3�A� I�C�
����G