// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B06zisFOTMVzTRXlFR89ZFstGAWlCozPakSaLoj5gZUvWgigeafd5DfS/3SScqnb
FinZmPc6eXOD4Cyoa4hu6KOyhKRHMe1nNErFIvJb9NNLG9SCSiUtcle5etkuBQCY
TgAw1vtHSAh9gsUhV+QMv3qEBEO6K+cgN7SB4cfipG4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 128720)
wbmmGQbVlLYHzf5d0bV6kIEf+IPVobG2MhJt3eo6zGKFuI6gBWDZVHJBxrm6ilb7
oyT23vGrkQwvLo2wzpSutbMz+yRPuNwYYyR2vrrfWd2vmGM/sjeujpDp9b2XFLiu
IfvOVBqv5kjBFGZ5WksraQZRoELxHq9HQiS05UOpXl3o+ed6t28Nct69XNDcr5u7
0MpgY8dDilOSndvJ53+fCuvPFWF7AFTE1Og984tlxkYPCeLopZDoQfWYATBd8dp1
ljRKWbztv0N4m3DBreYYOFzDFd06iOZ52bItZ4pEcXqma6e6quH0I16qgKmvnrpd
4SpfgSHI+D1D0HXtnxXuUUKF0Q7IJw+TSm3UgAV7blFX/ReRUJ+yzuC5T74idaH9
PQn8Hbvnp+yB3c6aX0KJg+YSg4PvtuR6/HNGb3BZrmiF48NqgMsGLyMwd7YOMMrH
eH72u2vZTPPDWwD0Awe5/VpwSUI9jgsv3Lv4ppkblW9o6w2DQ3zKwYEKLpW5R/th
zUgAcR3iuUvhwWDUqew6mcaq71baQIXneD6hvKbPvjme/+BLlniy28asBu2Xu2zC
OjQdU5GZgIk+0s/1aRoYLU51kCugmT64c0XiuM6oZZiHUopijb1+Ltjra8WPSoGC
NrpdcZMXni3aRZJRe1V3Z9L77WGp+lfn/MDYJGElFi2xhACnafWJ2TX4gt90sIXf
tHBROMGVXa170I3SALdtzXY2N0rzs9URocbBZPQmsUsnTq++GJfgQmHzixZaFt5Z
l6tmL90acC/r4CrXqsGOTO7KtTj6l/+Y2LQBqHLXyiR3gG2DBKJ7Z/v3Duj0khE3
LQAy1ENHqtA9ETtsIxJlmG4KXikMckIb6Wfswgh0zEKtJnrF6WxrVCulyKYg++SM
0pl6hvRVGXrKdxUm9np+xvAbSgg1iRwhrgXGcjHJahoDZQw4D+WhPgqKq+BvLZd8
JXub/VAh/fz/3+NZUSn40+1G/Th7iz5zSs03XMuzouwA7Bh6a1KtjvGP/4QGVe2a
IH5anmA6GYFxLwiipCF4k4cQGArnjrbUebZggZ+pufnI6KsYzlyFiVi7VkXm/rHy
91K09xCSG2hyOnf/vnQmwomYtwqqMK+pLXeDUQdR0DsLLeK7UA0tGS1o87hk7tgK
7WVOVrnaSwhuDEIL2dpApl5kWjeAFGOF33O/CWTl6JfdDfQkCwaTYVyZ53VnI+66
xcBwXspyLLjsiLk0jemES+LCt+KoaRygfTjlqLIIHh06g1C9XKIMItIPsrqHEB3F
jJm7E/028Wxh4tZAxwweur3KtKnoozsFEwsxPzItgart/I3S+aGNZKrcDLYGXffn
+3+jQdgNyay/bbAUKqx81WrNofuDelnC0R421P33ALuM3qSo34mM0vvV43t7Jh5l
Pv95aGsB8TbRRuKgocN4QjGN47eos8CU2P0R3l4AX6x6zyqNFqjIsooiKvc5mj1i
nO2QDGaweNQ+Jb02wukt6hGs6fIFM0G6MzH7cnmqqWed2PnJLWsGqLPV3vjL32Nj
IL86PmNKJPfPivzZN5f0I/2euHpx/acPky4RrDbOFSrf9O+eAjPwpXr6uWeeW0YQ
tzNQYSJyOYA+jsn5uxbcbu56J0DE7MlawRavCFMWv6OAtjutHIqstizoFPVKTF5Q
ik35fHy3DumninMrHeQn/RIZoFKg57RyRkukRr21ADKmTTfolVofsdu03Gbu1I6s
rwmQjjvvOMQ4xTzfBDc8CKCZYaJUWtMwKrwWX88ZwexPVDZaLxipE7aapIQzUyjK
XWVTnJIKkzOcXUJqjUDgzRIjRMme3YdRkZlkDVNtJLLN/pIcVsL38FFijMU1oF1J
EAQ3+lMLkKlIAh+76MEwzra3mbMG/8h3m7+TQiHgkXxNyYj5sLL6WFGxI66rsA/m
KkNg75WC9Jrh26HxXOlQA9f1LKO8jz33+58p94Dao0JyBa0RI3jLx/oT3nsv/J1d
2TFMnNZO4/pkqfWE1Stq9tGBkjRYSGQc2FXvHTrczwGcruWPp79SpCl8GIeEzkUq
8DDmZCEUgMV8qVlp4ek5Mw+Sg1wb/TZC/3pXf+in+v0rz6Nu4vkqLa5x0y6McIL5
1n+2zpkoePTSa5npv8H58lV+J0mF7seFAtmYi2a9N7Jx9HznQKQd+M6xhMzBviT6
/pyqDx8YfhATfY5k29vajIu40zulT1+E9mFDLr7SMq+tEqwFxub+qJvV18ros4uK
AH9wredrmtZ5fyKhdYODpjIEz2fCfKyZzHhEEf0KMS1zD6lWWm1eqOAzGBoVgW21
Nf+jpkandNtgH3wwoX3xHs8JF9PawYkM11qULpzg1ysK1hnr3k++DUqRsmXvzAQm
6W2MnEOmOHKofu4RE1UMG5oXYmqGdue2cBNTVDv+zE4jrPLwqghmVFxJQVGg9kDV
fYXqn1loD51IgvwqTNz36jxMa/O5PAMdOb4w9neXLw4HOa4KGrUfeqNuSPWWG1Nt
te6XZGXCld/vd93MveU2nuoX7cJi3dynvsM4ZPQeCfIDuOIzW1oFhgL2f4o+cTib
m9BoZKLQRiVVMf0j5XuY1tNc7+KQqO9N9VFwuvcUOOUna7Cdq5hhpjFwY0VCkP+1
M9r0ohPkbpLUnulMFmzcsIG1HhOcWz+f9dyo/H5664+VZvU5WIqWxOrBCPRc3LMA
9atUSt/mBR0VKAyBuMutA5VCMuYAmdBAfnLkhrAji7QRv1OVbCl8qevH7XFLaqpc
xWUq6pckwyFburIfphi6MiLLjiFxfp6H4wdENb4SPBrsAzGS/d1l30Yc6ASX8XoY
mZgFwo2PDUn6HqbUvfAxHdrc10SgNYUf2JzXtFqDMvla6zmUNp+Vov6YHscT8A+C
FwuuMJyojF5PVpp5niIrlaxENCpdKL4iJnlugJoqFs6zjUd3PlvV+skaXPQtRnHy
9qxeEaHtNoVbg5fGU8IBX/xiDjbwLPrmXXP7HttZ6zyt+teqXCMNcaFSioLSPMyZ
DCvOTsKwPlCXteB7zxc6UJHLnzF6LBRyC0Y4pM0uEY1V65nEPVW3XNVsNYewnxkp
4sqq26cXcCoCfymYdQotPLucwrryempiMklhJ0G1Ld4uqXiK/dUVBmrBvU+6rpU7
nR9md3EUOg+WkgPtPXCtXXurkjzcquig1+jWyjptt7m/GrNUf92gm0YqjnOAG0Ij
vr82w4Qa7pOMX93xkcVxMAXxkG5axCDGHSuEGenO33WnhZECoVQE2cPFJLlRSzP4
R6qapYjH681mss55kT1YHkQDWfHqB9QDj3aJKY0KIn42YfbzbiEZbR1UuPfZ5mgN
oBCSpdXb7/9pu5UahesQ78pHZr5QqO2ZO93KKzotHEHuB+Kqy9MRTKf27Xjbzad8
ATb+Q4X7Y6NZRDArlbA2n+dp8/Zjm7lFkMcXQ6glxAeoN05TFv4/5MnAFVGYM5jv
6ai2TdZuvpBNI59LXXVHHUUqbzqQb96fHf7OTEbDGlPFlU68WOIau1hD1pXwv9C3
wbdIOtR+ntVJiuzs5TzxDVJ7OnxsUS0u1RgiiaC8Wd/jugSgctmtexBBsfl39Soo
c9wBC0RD/yZwRGDV3SaPykIfy+vEpSJ1jQtdW3rgFhQt9HPxO8UjTH0fURScdztb
W3r4ecVdDatOXi/4RLnRmcsJOve+Q8/MXVEn0Fy7Yp5z1IYdDTcD4VgXTrpd0Ulf
Gn2Ih917yuT+mlxpck+OAuoPU6bbyBJC+IcdOPo8i0Nb1XuDnbVOSfJxYPhtlT61
dFMvRaWGmDzq5AjgG4WRwTgxtPVLZzWvRKa4MC7h6jQaQehrMGPw9nhiuvo3EXf3
By7cIG3M0HJRzOF3UF6z1go9H2UqlmEIciezMzdcgimcPoTm9JgtL8M0kB5LmdM7
ml9tR/asm5FR4FR5lJ/PbmrCTWBsbw6Z5xKnGLuPDkQhuOgqrKZ8n863WaoRQk2g
tqySBZ+vD1XycMlkYngHoY6nl33PYjnLkWqQ0K6iz2y+PIpcqw1XuupMDwr2ZAk0
RPj0p2n3WUUT4Dg2RDBA6A/qbGl+pqAKdSixZcNiD+l+aEz0NUShuNmcLmOGwmDQ
p0bUq837rW878j1lZoDfvPkC1EHhb5eojyYA0H+d7IHS+qisPIMKrdGHU4nEvlwT
t97+EPxSnkxzuFTgpWnbV/nw5TY54hSeJ5mQbPQMV47cMlA1hMqozUVROWWjcJqq
WeHb4a49tI4y4fA+wdwWP7EnnXik3nSvp7KNoHg0wT8Ccd7t3XfFW/ppEB0SlUUj
hK7GjXdxq9uAEV9gJ0Coew7JF6ITEcgyblIVWmW+MNsbvBKOD6MJc2huVrXjpadD
KKVNvOWimBkSWAXd2XTn7M8lhLftuYc6hzrl3ZqUPqabUi+vZdeg5PjxNE0CX9Ef
UzY9uZIgifmUNySqeDBZfTbw/NDHKMJPOigBgUnqSi5984G6aGixD/0fHY+YtNS8
I6flShLxTs7S6XVaUdJh7auz9axoDPOE06/6RMlTtF4Rh3FQSJAay/7A3lQ+ZYbW
4IvTyqI1r9aJrhRQKjtdDNkrviESvgcf/2eiNinO5OOOY6Pk/a9w/4QVjx7w+7yG
PysTJCRH20AJLNKfynWcsXn5tnYWQyVaDhipN/TyXenJHdghZzRyYS4hy5le7jBq
RvvE0Gls4bKaV7ogCjmi8dRGa2oR0Nvee0XXJloB+etBu6poLncnBlm7V6SCcNoE
DPJqzRs2ivs5MX2oFhFqNFcu22PIbvfL1ZWHrs+cWx6mWo6abVkXMHK21W29rcPP
ZmNDCYLriigVXHeEkCg7b2rXl5iyYbZWLSHuyrcJU2yHBpSdPVMUWFEcDv/YQPjG
snpQlMMqUlPlAMJLx2Qa983RHoGJOsjOl0jkpHjYV8Xn7Ch9wfpd+pCEKLCqFpyp
rrhiNo9TJ0sBUlqgTaFRzBHdYH3lar3M+iPICsWM8cvR0q2bF5IqQCSO8jkZsiKH
/j1tfJ2PkoD6f9on8QGY8Urp0kMFuJGfndWHyO3ROlIGwT3Hnw6tRctquz9hi9MW
vMvviTdmK6KGXKq7n2k3q/TCe+Nhr3Sb6My4lj4KIGEyb+i4GM5j1BBEmhuU6Hcd
bYCJhQ93T/S1CT1CM7DdK0EoABw+1JEzVOvl5MlonfGAfCWd30d/4MyprBslClRs
qCudUbkbVrdsxlwl5XULX9XpQRY4NMzeKljJbzlVIh38JOdFHMUWdeNWCMtFWuHH
3l7ZVqYGOhh6nB5qRKk645fgF4D7Ni9TUV7UwWvpocXK82bv00yOxboXeEz14oEH
b67rxhYHV0zf+Vwz4VjZcSEISXu4DcJzN7/IffRxuCLS7LwiesGMrDnkT4usPhre
NFsVAvyndfPcUgxZPiKWyHI10Cahpp03pkfaaSxBBYAXpxcciOBgvnCQOV04BS7T
tH3IanqBwS9FMvZ9t171foy+FfynNV+9E/1aa+DD6RRzndhzPN7i8gG6VYbZ3mjr
p05gT2VTbXskJALa2A34Ni4on5ga6YCZS57VCBTWpvEyEZ6rhXjzdFRZHkbOrxdF
iso0B3ObJWP3WBInAj81r7jb+1rZW/9jxbSRrEmiKC2KM6Mr3ZIkpCxDshvbxgRz
ogqOPzkFxgIV4o3nX4TfNJyRU25F93fT3lwtrqHxyxbVcXX/2yqQVzgM7QSgl1k9
0Q3zvLIDIRWCXRfm0y/Gm3Pmt5s2RZXfz+T8RtV4KLNRMxZvyGbJD26+8b1yHYA6
B7JsK7Qdy/fRd8Z2BLu+Wqp8SuuIYYJDi4Kh8aOHKvRZO3IDZGIBFn8Y7c2USxgO
XZbl9rmspBRxeg0uqPBLJvB5k/1v2cEDY/ZwQSUTk4pA2QcBBxLOPvYwDn++ExuQ
14fRA/Um3R95EavFNAphdoCXbRLUScsHZZ9bIA+9+CwNPD3UPEISD+ahB2UGRmg+
zyy7yKs4Fhmi9xp2UKgpJUyFtxn40U1WeK6YogzW7BWJFLv5iMEUlWfEHBHXeYUg
OGgYkg/tr+mEP+y5igpKFuug/BzRcR3mQZ1Qn9Q+XkwDfoEomKme2vFhiNKq+GNP
7kSXAnhwuU0cvEoeWuGaG8CSC+CnPTc3LxvQS5/8xlxYiwrLZkW1uWWobbl93nsi
EC6UjcY71VyesjSLfFSlDL/ogAVqq4YLmus2ASCWS1FjnfZavow+krvtjY5PP85O
Nr2rBSaLjllI7YZPpLo42dZ5uFiEyKIYttrwIZxHa39AE3Kd620NRBttJyYIZkhm
vNlZ3+UdypzyJZ1xz+xbsKhFC+HMpjJ6C3f38T8R8ajbDIpDn/thJp8W/T9g+jMf
D3+tobj/LANA6RHE1xuBp1QJMW9x/XU/GqaaBB0qgd2jSVuveylJLSCMOl4izk7+
yzO2E6AgdTSFV0OLYdCYiNUCO8LwyZWL9nBPHub272BlQ5Fsg7jUUYoa9N6YZ7vz
xo1Ofk5qkwZd8C15MMABSGhdM1mv8MrTWcy9srtCvKbOFdupfiRt/TcnMzFdMNLT
/ZRMQTXH51r3Oq1a+vLptSVDCgZQ8m3tqWu3K12CNljOWfnfCFqNoM5jdzlsmYku
9H9NgUa5utAJlOoiGDsG2UaayxqkRcaQXUO4njU96DCtc1+7JR4Eggmv3gj5VDjU
PrtW9T6rx6LGzmHQmzKYDsLLGrNnyUQ0hOH/Y8s1qIzKLxRlFfCYZXL0y7c3hkqo
Fb87/cfpCMWZ134o1wsWcVT1yTLHjB8O9LA0m4dld0M/ACIvnA8Edai535CSGjyX
EBCyVMPa8K9zTh3V/qBHHextfMeKmxspLgvNMMNL3VlC8X+8wso5Irum/n9ZfXCt
J9j5R70GIzrsB2PFEVGzVSWp3DXv1B/B+eWt0KOfW1gQMBLlR2mATtDh1h+Wtu6i
yNgT0HmyZQ4Mn7x6HT5hjFM03iydNaTVP4DLA8TgRXMuMdB8WetQxN4LUaqSRUri
plU/N0F9iVl7pbpprRXMjO3AyZQyB59Sop0po9bOmlEuEAWrPVpev+sN2J/8aNbq
zVsJi7mz9kr+juWDkzdcP9nFFWmEmmih1CQKGY10pBAzkv814LecK6/nVJFsUA5o
jmuKJqU54GuPUNbSu5usWmf8r9vAL8UkjqQrpZg9D26r0g6KTrFkpgh/WS+e+NJi
w1twNqnDSn+ucEnXItm+RqUhM56J29NBMpIq/XeOtV24gnYmQpjBKVCw5wxqqtU7
hsi3/8mITd+LUbMG2fTdbYwY8V6GoSJi68qSekCN5IQB0D7nXkDApzBub5mYWTNf
kTPJwo2xGpd1El66qb2IuOHb69/ThckOPWL+1WR77t/AlQbnpclzWPauXs2a2la8
qXgV9viXMeMB0NBTWk6Yh3OVxSOejCG4hf2KoYsF/u9isIF5b9tomvbcJG4piPyB
C/nJzN681UIUeTiktCNHqE2MHRYjYf9SZ6i0DuEA37pxHzHrIwmRogfRDYj8IFeq
885CmfSDsd/GZ72D6weNXeS1AwO/KgY7n9n2n4tvVc/S1+WC0VsJHiag1qJWGvHV
UyEU8n4dRRLeMrdDcBpb7TOVlG5YhCygkHDooI2CG8Wv5F5PfSTFFcarSI8iNs9S
XJuID7JPR3xuRWEz/9i7Wx6opRGPigQBN8auZlc6sOHRO/Lw119RDqYA5LqUr0Rn
0C6GhOOYj98MP5aIVytFsPGLyy80gNyEhECvBxPiRm9Q2G6jOMG9pX+F7dodkK8r
5abPxTsWo1Ofbi04Me3mOL77go5dKhpuUC9D69sfj+GrB/rAME0CFDQYEC99BFvh
Mk813EWUFbN3+Zb262+hP9MlmMRpbBTZXyTNL9Ov50oe2XkwQPhsm5DkS1FUW2lD
9SfJuXVaWlEFZvjyUwER14VyKLpcjgP/O7x0fTonL+Mv2YVny6flHTurkC98Baeh
GGsDCdxMG/bAlwPJig8wkRlF9YlBEw0poOUCmvCqyYedi/YERUv32Jsh2BNLV8ia
QcoqGsbeo4imIH0zWyncYtSnu+ADMeH3AGxwIh98RDwgewEmIBrmBQU0N8V46JNz
KTvN4tzFAYnZAGmtbvzZ8JFWUIhS95MUzhg1GooIQ0Y0DYWvVoMQr5DKSJHb1lqI
0vsBmDvmXxTzpUFxjDd9ZPoCSZLphicuELo/lZKzkyxLCqkUGMmAj6jHNjWZoV+m
sIo7rLRcmCMttEnliyC1j49fhDDsS4MahDtmNWpmDo+pRwg97PyQVLSoUKuCnYJB
O4dzNlbRoQOp410mYS1ycrAEiC7DUF7pHIblvYMWt3fqk1xu3lE/w8XqRtQNXW9F
Qe8Lki5UfWCk2nj1rB6pdkzB6zRnU0ymVvB44G+4OSUeIeFZ92VQJgT6/bh+Xvqe
UZ7UY2dZ+OXby8VemdmA9CL3Df7pVxtN7KBu5FRTBvIlXBTnN6fh7Y6UOZdbF4Fg
NSANZrRj6DUExZPluVKC/zk/85FvpntMjTXed56MRebuTQ+8/GLAmolNrBK1MPRq
0bdMyocObXq07PtXOawnLhCUTnqcmGjrWlrT9OveIGLOgiJolT9z9/dYDt8V9NaF
G0P6mLBVYmbd6WqoGf2Mqt2stf8Af0JuftT+MgpZanjL5JQaWFy9vh2czQcA4LT8
OMgfqkIeS9IfRpFls+OSsw2Z7bU+yKZFWJM0cIyQnf06d9HL0ACufD4AxXlquEPN
bdLaI6A+tU+laEWGVZCkiovOwNi1TUfk7TYGj3UBG+TQA4E8X6K1rItuAunLLu1y
gX//IP5XvMv0na01N2S11iPpUKgSKxzrbBJ62mdUAIE58kYMEuWUrRP+p5Vjdz8/
dG2iLhlGUL+PPB2VZklEIUB1svR9YV5AsFyr/zOwsHdc4d9uCk9Lo0kXkqapK62w
dnOYgSwShIccDQkLWy0lY5tpeHknHoN4XLfcFZmpIEkkHFmHcvL1Rm8sM2E4kOGS
JtjA87wQUWbib73PcmVPfW+XPGwA/ynjrF3+xT45y3RkC/YToBTkbOVVuSkfVuhC
h4VU/c5zUcA9w+zKk27G4MlrQ+/SD5QT7+WCzHlNUOxtt/6X8KN44gurWgEo55Vi
59yphX7cKg6JYYOOyp4U+4IULYdGVKBj90eUaqhoormDEVQaC6cxffRKk1KZVR/L
mcYiKPLqnBgUXH8rCwi4ANytujH4hwZ0zbXdSvlCZijXHJOfNlIaaVhM0D57qij5
sqg45S6VdyIlmJgLu9RIf5NL2/SBINufUdpqYtxt8D5HMGc2Bk5232Vr17MFw5lE
1iH76T7Tuzay0zNEKHnfyKMPUxvOWl2va8FBnRvkGI3YU9YqnQT5poKPUwlx0auI
N0SCWNkf/hP/DgkfbZ1/AvoOekKDkF04D9KyH0NRL74EPAE49mC3Ar++igwCUiQN
Vi7f7p72xYeRUTW3uxzKGkwddrRGHGBUr4mdxpTuWzgg89eIPiIUHs6wNY7KwkC3
D88SBtPWdsEVkeDE3uPc2m5Yc1nk3CGBumFvk7z5MwO4XlPzhDOGhwKdiJ/ss9K4
/HpQF3PUeEjcmEaPBphrLzCYgcl1Qsg5Ol5Mznj+m9kh7dsFBTeILUQugZLKBG8R
EgmzrDod4s2+OpFv1o/bf2XiyDdVMAkFrmf3rO3YJi2f8a3NqHdpifwIESfFzlwk
LqYIEehHqlsEI/d+6eXJC1sE6pVV5MxTduQrsLFsEHgEcdy5MMuJhl9RRS6A2qJS
gdcZ2smdJuD6jf8j61R1JVYu7DqAaUU1TdCoiygmHckf3qkP0LmhaA9Y+7/SuNON
V7W0LMfmDGSI7nAtYIn77L0fKMUOjwDUbKKlsTpQyWxJJs9/58ndCIQDd8MfjNeU
eacT5uILle97MYlGoqJmtQ1iSmgPar8M17ZiC392UZGTg4wcIB247/AUkQ+0li64
u3yWlGjPIYi/w9ovXHd0igaUsNEGxnx8V0Jwe54fbKgWnvWnWyirtvSr3/12WzAz
Kr2nmUPQDAXchSShsgffA7zTwSl/zeZnsGceYQRkk6cm6CBnUf8wfXxdVenpXoKM
t4rzoDrL40ZdzX+Czf5Bth9SaQkWJh+6mB0Ao1FDqT7qg7BUMKQ3iqX+VHfHOhMg
cdesLWqyfgEZarzdjyNQiOZUG0B1dFYJ8r+fQPYdVx9I8eOJVlPWcazOrxOr9tYd
PReuLsXg5jvWN9XhQQRYVUFkHBdGvV+GVY/YNClPHpIW0HjoKqzYdFnhZSWb8DHW
JDZb05koTgzb9JAJ9o38Y+BAYHVXVSYd8bO6YVe1PusxLzvwAI+iZ7nNEquEJxAO
Pdm6W6jxmg77Ng/1AlWj6uU5B+BH8qJK635RPisRTH+g5vtlex+L+mZ8/8Ay1jCY
k+Xvny5PrDCykZxdebLTnVibtbcreSna8xtemoN180Qbb7wuZxe9ZGQ+WYY3FO+s
HCqyi74JzUVy+R2R4W6z+H+RkNX5s28v0FwZj8lnz5CfjmPAP1SglCbcDB7/5wqO
20kqWe2T7LEzw4F7wxRy7Or1EIFjWj1+binvOebJLpFyPSpu2dCMn2KUCkoYSz3q
fxUGpUtGB8EGOete8kSYlVjdOPdDpboStldVhI3YOSRWOXimE8VsDIwEBNk+hO8J
dw9oRU5iZ4V217VipeE+HKPkImZnB3Vq4ppWqd66kEJ18usgY/4/6KFC+7ZoRJKx
UaqB6jXlAwdq+nQMhACCHYBoQpIrJpqFmSp8HzwmSIIa5FRDF8i+aTc+Wp3SFdVB
qS85Hv7IuMviGABsDiiatkfKc7Duopy/bi/dqrNPapvRCSH839VwvlLedR0vluCu
c8fsGkW1F6iJT8Lap/Q86cfMZN4BqXAO9fS7tCuPRXDtnO+YoT/S3N1AWF23q4aj
QWX968tW5c5vDBRRKaBNo02XWOax2uGzYpOXonC6b+I3zjfciAa5shOG2Zq5LP5h
nuJbN+zUXKsyw08hd9woO5CKfyE216pF7IjHLlMM++iwdw8JVF0u0c0tdgVZwTaY
+jW7bSwOFjgFHQusEkrENJRrVSeO9H5TcvDMteKUHU3iR0sE8DuZxIBXpQNnxfig
aGbpr9nRsFs8lnEwBDurIh+a8lXbskR5Q118640Pr8yzPkkzVdidpzKWurtOdhSK
gxPRLgxGyFSrbo0dGpQcUpJeC2LjK3yzhp8o+anQ5WcLeNEEO131RRQyQxx8RpMm
DZXd3Qs8XIxXqCz4t6NtZOyXZzSF3JPwn3zf7tFOmY8c7tBh6jkX/uY6e2A7SJr0
rz2FfU2kRg4TtSuQlNiwZc+NvytJT4zUJlm+KfoNaa+Nkg7srTYN8bhROMs0D+hg
T9zCW5HUoB38tL1wpII2WkyiIi72FWU4+28Gr7C9gfCMUsdcbjbMz3T5MDcsM8Yw
HZgkttDcUFO08tB/hu66eZlMpMJUfsjHmk4l9jasNMLb9z3z/SAAJOu/2cn/NtRk
RZGdEJmb9f3S3Z65MmFMNxLG7s2FcW/rUdxIlSPbHEsOaqpTrGrt/tqdrfC225a4
wq7P1s9VBOYhtBrPyha1dnsUFuDgyGH7ZrG1uwXWzb7LM805ESMGRFka4FbsAwG4
KvaKYeITNnzOU2pYqqPOYqmQ6gUGCu9yJRvcVzkoFIN9iew8ffROP9XJqr+ReSxB
UxpfVdBpvxdBz0nwWsD2PSyYjzN68agHF6RTKC0rXxJ5M2tGJimKMafIlCC3Z+KW
Bob6RZ8gdMM2U+S580x4O0I/6fw2AHOtf+FQqfRQ7bLaI2jwaQ39kvNF+QzqILhW
FPNNs1IASLb6n4FzAyxSersShgzi15xMSB7mnb7DR2cKZxyt7GBDRoHGagF09p1t
7mukK2FgXjxRYxlZEQiZBaR/5UZS74ICKpyR6Y43IzqauJOIKKT2FYCg/l81wY7R
8+H8a2kc+iVOd00pMC/sUk5b7mRoZnTycXrRA4v1/8Mx0GkSmWF19Z/tfckrY1Q0
LVWizMB2PPf3Idcvx+0cWBeYg3gN+te0ipzILU9kECvp9ukckF5Vn9o/VwHZKMTe
gLcBCRhLr0B3QI7gTDZhZ7jfMqOuEpVa9Qz+Cc1svW/Vz1Y2oMVg10jB8+od+dqs
W43lcg7hyKmXPCA7eftx1Q7GpAVtjk+fZ+TeXyWPFcBPxtxSg6CNaHvc+Ozi9m6z
NiU0HlMZnT+eAXBjHDxB2lxmDxZuqMP56Jv00L14ArxC4HC8YVXI7o8cQ6JwxnYp
avUQ+L9IPh2AoH9wYgQM6yTNFNuBDLhps6gHYv71ZS3PD8YOlmn3yS67NXWzsia1
XLGNGE3JYh46I8W1dEP+h4jpoCGaOHqBtytcmNvXiU3w5Tge9Nhcz7sj9/pZ5/9r
vALNFagSDcp7aMw1Ly35iJLpYfJw4YASfkPqqkYEpYEnYr9O3ne9yScS+BG0Ezjq
nIuxe2KvzYUTmGr/5CHW1kvIUpV1uqzuo54+xSi3vFlVgBjkaFCBnZKbW9m4rdWq
v6KUDkKkScsDlKGSvOmP2pMFR6618UWxUJ7V2PjTiWzVaV1lCD950vURK9fsVZ8A
sC8B9q7eY7a+RWAGvN4oSlgItSqcDYiDPrpFlhRb1Uw2i98u+FHJiMemm0p5u/Po
g6Vh/Xysu0HSvdVJhZu2IsyYXCiSli2pKvYMiIjc9dizR+55+dpQ+sb++uqHGOlk
zFgh2AUZvrw1V5yomcH3LwuZeYHDCFPqvjQ8h/ep2BoXqTUeOspCvFhr38LWP9qq
vp5Rf4/UDBHS+5rd0u+IGSEeKaSeYb0m34j9x1n3jHujOtTliLxfwEaj3izd7LSg
OBinrMumSoYCGELB1B+imKemVbyNOeAvv/QgNYO6+vTm+RoGHuvcfMEvqQkvQIIY
F62Ij5UqcsgFudMYrzSNvSv6+5KXmItO3Qcw1skz0FmkZViFFU7DKojXuUacu71u
bsuu9atySRYrnq0vQ0+a8edlqb3IF0oLOCcVQDEEnP5PQhO66x3cmAIL4TdIxl+B
7LWuyPGObRRmGvWKodRWWVJcLXtdiQFNtBO5/YYVDhl1ctLquqZiaoNoPq4X6VUb
jEsbAbyqi0oHhFbMJ+4YhiLoqboS0N+5rWa7PLbllfaIKtmOTW2hsTzyMTN+V4O/
94FbE/VrAo/I2nODfYr3k27fQaHv0k6jmHfeF9v+y+zI9jr6fkHlddjc+ZsCMF6o
wXa40RjzKPXrNmZ0qICZg9z8bxFDftg3TGz115smJZ4xqk4Y3HYXoCSQwC8zAy84
HZd2QCACggEJK/St7E413qkZ+6mjenmDV98UL1m8n7ddVTNpVWvqSDAf1KTuGTPn
SVty8BH+4K0HxkaXGcfS8MstDLTRXPrlhXk0219Gt3GzCe2225t/r9W6C8pEMLyr
pevvbKmw19EWEI+31ntvWYYLPzhwDuPynqVCCk1xCCJ4D+qKyG2og0Zrt61ZZsvS
2AnjXu4i8tn5gnOtns0njpqAlvc42SuMkoAPWNRX/B6rGGvqiLxwlYRXecL23z6w
n8Za9nFkmDy3bUadISD9OL6TxuChNpUNcgGl8MN5MJ2cwR2SXa4MlOA1EhWP5LqQ
CjHIAfrvzEx2mfpsH+32KVO31crgccreOe1Kv74G3v/2rV7uujThSBVhGHy8VeMI
J/W8+LPFts0cGMza0Nwl65lNYat9DEVpw5/RZVIP9zgjA4Xy5LWE2sCvPyVhQtNW
0aAe7kw/8riVt2enVl31hfQDmE9jz3OIqGS7WDlPHBPiDtK8VqYJfoQn8xqhsyhz
ksG0M5+6E6UXaeDe4XQ5255YhUkwvtu7GUr8/RughHEsqMxTvRhT/kQ3jEtawgjw
6ZcEwGByl3rVmxDSv8D+P6zlcgEPTUJ94V+jTaD0hHpv+9tQQeVbkvWgQ0KTkzsY
sjgl3Qdx+WTpYCSIxJhLspRoIL8efIR9VN+hPQekJq6sI/HZq+6qpg0cfIvAurUM
3G9ObmxMnI0tWErKUE9ePz2GUVEsKhkA8yeJslFB1jAlFIKDfzFfdHT3Ki8GvH6R
lXHlIbsgAxRWYMODGasp4OYDNUtbN3mizJiofgFDMfvOysaUqVuFabbjsUU9wdE2
HypczbQLWrCyk2yZy46a6V20LryxMVvSBV4+DvOHfyNDelZchsHmOksr+DovsTfh
86OLyCPgy+hdNzBT6q8KvdU+yw5YBlSpzHi2axWdhsulkBdEBAl5n0CDxt1VvvbV
12QOOOOgh17zdLdq21y+EPNI3OALTwPoKz8ZmEVzofjfoZEmTwJ8NnPu1/cN+QOD
Ap02RKZo4uRuFFOWgPDz/dlnhSlg6Ijv4KaYpTOhYj0JoDMUFHny+X4tT9WqEdhW
q4TC9TtFK0c5YhDDn++sT13fYurCsJMCC6SRu7JlOEfNtR4qI6/n/n1lSymWxhF8
DZQc1yTNFBU2rfVlYqywpPHk0m46mBJKjmEIQcAND9qsM+zZpcyl4ZlF+TYFzR23
357slTX9TT+IoX27Wr5pj6iAyx8v3okSv/sNqRdOiqfD9KchnDarhTT98F6atJLZ
cN72ohgdm525LKTE6qCGuixkqu/JvqRezLrjsTvIAp1eCJBw4iEQD8r4tmxUpdfI
uMy0RJCMgDXtmS80p8lvB+jufr6rpMFAWulmRoQ4MkkPALOg+ZwSOMdnjrsaWuHH
yaSVUaVvgE5qARIcu1nlo4P7f498As6wbuop64nMQkh2F9blD1Qq6MP6wIXaB18Y
Hq+hM7Vw6fWpRvC3hLrsmzTSTmdpciAo0fkW1l/6Xr3YhELxwG5qbByPdOCWinnl
84kgFsMEzPtUjXgU6LUFAmlEjDV6DGLKf7hQbTIjpI/qYsqpoh54g7pPSfN6N3mu
s0r1Y2Os2GYTL/45VuP9VLw1e+xuYKJC5oz2PP6WgnUjjsO911zp1jkCfcCASdp0
Hr3lxcJ/MKTOFcbqg2QAvWsSSo+WQ1sCZjN9FVdZq54kjgnjSm69vmBE0RxH5KNv
qi30SC39dQts7uS5y2OfL879208/pjiUfs3ChlqYjD5d9Kd8/AG5NF0SoLmdIVO/
0scQ05f+Mv47vGX5vqD+LJ9NlGPPmbv/CW2qTg0sKzS92RT+n5LBPdDit2aRhw6C
uLpStYcWZrgcuScE/wV2fomYySW52hkdtjXSqNftFaWH85I6inMymoN3S5FOuh9z
9n5pb2+VNrMmDO4OWdFBpBzKsXPrZX7j3FH/pbfJO5SCMqSKWBBXRWNLPvBtt+Oa
MPyQeYBWLbpPUdOfE8rX/lj2UeRo96eg+QmJNC+YLzCOf/5hkwTjBQSxIvbuc/Ko
bwM9SauAfpsIx3C5a/3SlGuS3bJrOEVHaBIZV9ZHngDmks2AGCaQu2iMI5fsdBgS
bgbjL2AcFIQFg511+Oq1NtT0KD/YlYGMQbngqjWtsikjbwG6UYY/OZ8FZD7lBO4N
PI5Amw5WDmey1WV4/50V1jiRYorbfwoFMlqvvlBZ5QmiKaCTdtxBe9rfEIP+vy7S
zByTWF+A9t0rb2tfCA/GrRtu+8mkrlCsi6lbwyh3SGb/5Ab7u1AzHpptmyUOTXjq
vX3jognD+xnYsST5ILmwVDYCfwTOXlD1kK1cHmTfxxaX+bMcx3SWOq5kN3vpz/XF
Lut+6BA6Vq4XCboJlvH/G9PtVTvbg3A/GVQ9YBqd+IriHPDb7EpxmOEv8M3vy7Oc
1aVeME5mRSw/e77OsbzsohPz2xZkEyFqC6Krleb6aJLFMv9qnywAAPSbVMkwIMA2
EYY4RwcZefCyqlKSfU1B/ZhuNVlxijFpWukR0egDdD73HLaeLWct5hjyiwqUjoPg
hYHvyeeRT1v+5mvOnysxIEFF1V35N/IkDCggSLY6xg8wgKnYl4LkIWLamcUyZQXR
FeRVgUBqgnMJkZgNLIwEnMCCyK9ag8/pQUQhgVCTaqrSTMUVlutWd40Lr9rTJQye
axYkDSzfqySm3qlMCORDL8YS0R/atqbAFKuRL3rcY/Kzelcnjk0UFZLIypM6VTuv
TcOJ4A7Pqj6BNcwXsxXE8o/HS96TVJGpPbMl9/8C6Sy97x/Z8a3hl99xNNIyMTlP
Xjpc4FIf8DK+TuH9loB0cS14mA1HIl+LVY1ma6IgZE27S6wsU7vRkrkxaWP2hYvs
H8wGSyIvFdqo9Zta5/GgOdetxx3dRhmaVyD6dk4v8h3K8G1QLeN38yG7Gu2/+zY1
rdobR5PJv8+oQesQf5DLZh2yjhj+Y/xI+KCbck/YCWDq1EyGyZAPxNAWkjMfpLEV
TgHzI3HPJerbhQ9ydhfysIh/Ngto+2vYcQBEmA4M1Ri2ka/gdEJxmjFfcg4CSpzu
SOx4WzHKcIesTJ63EdJXPdYxVPoLK4avn9YT/XLiJps7cVkOndMGi/OjufzTokVY
Iy8EG9Uzcvb1m9u+NWhkZNfowRmmzlsv5UVS6X6DNJhW/KRJk8LaVxsf5BKvxMWy
GJmuAGWWp8A6XCUUGQ64/amZc5Y8rK03pTO1WQCSFHDp9sKdjN+Ububyf/OMLnvy
6NZ74kVg6J3v4mllllA0pKFYWgNST5/cc6oWwkkCMxdsP2rA1vjvsN7osG6j/+Iv
I6ExaHfkiHyPIH+7COYdXkxS0Wbe8I26B8vUxMJRPj1DpNfT+6h8dOGzy9Dqxv14
ZBmOLJAIn1wME5hcQCp9EXsHdqcduEWOfwtu26IpojIJQoC3J/os0TOEbUnGZxie
veKT/p6Unb8SakMHYSswYFFKPUik+4a4MTt7D9fEiAAsGeeylXfgFUiYRaWO6jot
W+lrblxbobk8qfF+cBWop9nQQ/rGy4JtFBdiD3dWXbOhATCkZw3o8R5c1k36UgPp
cvK1rUGiFedVwTqxj0z2EohJ71QfYhkBeOHV4zBIVazYLypwUz/NRtDAfVIor1vA
oIo2p4bQ+lkN2IXqDauX6v1ExEfVO1WRewrAitRWoqoZFKdsxlkfXPbZAtXK0nke
8wOVsjMiBoKg9InAz1Ot1K/A6kmfTHdvVpyaUDamKYTpBbIKhzmiSwxLGE8oOuMx
IoiIGRqfjInt1hP6yNiz7bXh/ySjaYiLL+AJtGUqObcSBNuopzWHP0H2Xm7OF0LR
VaX8N0cTRN6nqYgpZ0lCNNiYoPswIIBdJiN8ImWe5GfR8fPXFRK0SGi1ZHBP75Ha
wkUM3yqhr1qYhdBvcn28EV1fAXZibV1HhdPKCs0z+jZDDtSwu6lmUQfGavBOZWTy
VGXBClFzKtoSr0mUSHtcAWs7jETRcvKUpUgcVL7EpYmdvYpaXPbvMNRiOnBXj7C7
E1D9fQZ2flGm1xRzgvah+L1JW8MOrrTP1o2hdbZvHHA9cxXR4P+zLXxnCXQYheS+
PpCqeQ6xNzqykNhhp5idp/Rt3tgaZR742DHaOLTxmOFa+XCMV9szsEnAoZAegAP6
JM2T8IvEQooGwWN6IyNbZqLimqa08fmJzwyzCq8Dmcz+ryG5A+w7GZxwrv3KxBuz
61MgOimULpnHEEaxQVqtvKPc1m+kum/6md+HZCU7ToFgnREtBUPmvMCIUoYBRSmq
gmcceORqBvC0BCWZ4gTgFq5cOirCD0+sL7ecjISmB0tnJL8v/Z1mzJaEcLnEFZ0p
8yVRlGZjJNN8SoxFgh3B8UwBx59hLd/O+sFRLmkOybGsoqZOIeqBATBu0vJrvp93
DHaS9p36zX4Q7oRXCdIp0cngZ1MAZvo4aKVOoKeXDFrfy0t2a5apFtfUQW1PPCYf
q6TBHlIx+a+l5MNpIRMmPt9q3Ats2pEZ7guSLQ2J45jCZEYMa+fOU9ErlCC4brhq
+THJnJw+Zt8j0wdeF23+8DSnUVGXnY4Fj2qf2mmn62xb/WS3JKe5JzBrvNg+5k1e
TTB0sFb3XQBEAGH4CyFfczXtHJDGuotpUsdr19lJrn0LQzDklpEJqYTt81czkN2W
3sJiFZTPV+y4msioC99BcJmFCn1c2ePM1RNyT7HHYW0+p8RGyG7mP40zt2fuBIWR
DOzxzXTpl1Nm6kKDgMahtSBQZJqACAJ/STXT1FVRhsvlZz0l5DOYCwFffDx8D2hB
GREOK9cZtE2g80NG+VqIcNrMKy9QikGXaZtx3YqNzH1wUWuVd2tMSJAi3IWyDDyw
ZMl98nDGk0tdMzpjFPgZtFexRGMG9opk+yrelbAd6fCrkCOXcnu8MDfuJiDbBomi
Qlv+5jFP8phfMcLLsgVqr3jwo3oPZBW9HmKcHtiN6TaVBBiJXraEHHyTeUNBlsV6
WJa1CqniJEo8LwW3sj88w7vlZ+gFmSbGlJPvQjXDmSXDe/B7Sdkbz7n69CMQKfls
ye3gE2ZZYmnrOabuaMrHSriDYkPiwjQm2aZLIu4n0QkdldfMI/tIJrmZHwrXAq4x
Fnpi7+YOCc9Qa9JBCistT85fyAqIxyoiqpvejeVQN5ibebomgB+psMSON7xpHbiY
B+UO9VabWloPqlhux7a4uIn92TSEP6xKJDTMjXYoDdLalEc+A4VPsUdGpFJvqqfv
rz4pQm5gFvQBCfxygE0nAgRTxcO07ODFzGmlbQ6KpBp74faF1X+ki/OpN6zxaHCf
Qx4ykGjloDP3mgfOplNURJS2uoFHLWnrQEhMAX5kuDjiLhvieOzD1/y9f+l2Cwbq
c4XAd7x6AvBKur+T8U/rG5nKUmgZHECMl/8MQsGtRSsZjr3M1CMVVXdpslY+IjKg
MShNTwmYCmE5tzWR+W4E/1T7aicRB67+GtfLbq+NmUT3mijmXwKk5SeCmmftq2T2
RoK6AezxLPJ7NnddKoGZEd9O7LGzrl9lj186e4Bja7M1S4ZLxg161ZIQRsyA+chb
EjbcWpAKLxiQu2O8+pbUuGy89RjFhQZ453SAzkml1+RsScCmfKMy4K0nh/YKhdPg
dY7aEjPw6FYi6sr90HZzDRquCfrvKSDOIo8W6pHrzceOScMkCQsvPzVjq5UqaVaI
EY8CN6XcB6oiCGPEH93MkA/7VwUlzRdd7Rebej5bGtSPeOSKTXvdBq2RLPi+BQDW
n3WS4UVrLVmmgLXa7GpOdUmIZ0ggPIqvpD7YgXdZKcYmyZgcIrWIpj0leKfyw2S2
c2C6pGT9kUNn9OE5YYpfxHMRx+3mydzANdeii+BaiPbSjaO0Wrmfl1SCgIljSN8X
upWXlC+MWj6rIO6347gqd4YDthtiiGNFCLbSdNO3FBaqc+gAWQQUvk33JyHMQNGL
ZfdWcKfehH6CYZb0gpZOOx7Hs3Fv25mJtbSXTIxKALsUHNFVQ4bKyiTITdmkE9ap
5YfMCi1t5kjhcQxSzxO+tlzvuHXEKNQ3JxgFrUm+d2bF5FIljygmKiim2cKEZDEm
0ssmXIVgJfggUSvKlarKMLnrkdZHCD3pakMsd+G2YfPVTkjjSJjfVU/2sqIi7sLl
+v2caHd6LUdqX2hy7yQYnz3rdk/2+o70nmXWgywDzChOSEJPSmzu+Tm2qUDH7JzQ
XJC39RRsdT6Z2XQwoXGF2MfEufdAxMutwYlUuGbl5qx/2Fva/1nylA+H5xKqi30k
03+FOkO1XyoA6srQywXg41OMZVVKwmkUWzJ9tZA/ua7Clbwr2X74v6oD1aXKN9d1
WZvO4UCDmFCBPcvKQKUyIgBhTe2gT6J4sU1ajBVg493I7MLAeCohfMuGh4aSSSy4
Ghh3/3FM4V5WoLS4z8oFkp0NFN9i0K9OwjAPbYl9kY5HheQbKKi2AHD+6M4ngROR
FwwrSJhKRqE5XawzGr3qc3yRvktKM6hzeT8XXwwq1eYEUs7gSBTAzo/0jHRMK5AR
CLrJm+j1GRmjAQQGWe6iEHkrP5PWEuL5e95wgqHLtUWtGmSS6YuhI5mxNvwVQJrE
YtQhWtcQmhX7bAm6UFznehhYiq04WGisa28cL0F+UNN2r61Sc1cZScScE7K63zLr
wLRwyCaaY+COt/GKHWcmedTHyA7plBqn5Uj3DAemnx4UFYkWTVcX19IYNvfg+FaH
e5wiQ6b/fueH3MGLuoN1aFb668lHOJwb9F718lLYbGUAeWRUtRgKxzJZA59r1iX/
IU2plY0TFAjr4p9Q4v4Q/XElFMPTGTxqS1+t3qorUJ2CKTCuCVz/if4050fpdDB5
XoZ/WZHWBCiKRA7fkdBKNrBoHlYlKyyHw2TlMlGw9OD4dFwHoaaszcj1yYSIEWHP
Fq10TuU1gw3HunW0IBZjI5CJeZIx9f2bINrtRz6iDkmw9nNRDmc9mVP+wbYRfHhM
8b3VrqkPXy9vRop/roIpkDwd+6+cLwSA5ig2bdnNPbDAv17AhUX/kNRK9AJoCjXt
DXim/M7zGJKsbr3x5t/E0UAJXIi11ENMCfv331ukns5hOY0JrGfRzVUx1vwe/T82
oK4wJvaG9oFzHtjLfaYL7dPPCrs8o6p64OguFpHgmGUwbi3N1KSYUCcSVApP9dQc
pluuyq0/XrZuX051PCoNQMxYpPpGjNNuQ9VsfVzpoV1uCWtf9TbLWrzX+/luM/6O
rfXr1xSoZJhQ81bd8LSRxylhF0CcORgjARTaDl9ngUMdzp0KIcYZkaNkxZ7QwQzw
alljVX4ahuebJFjqawo17enhmHm1+KakmQTPDXOeDx5psmX6N52IwHhdrzuUeWkE
+NIkO+6YbfkE7DBwv8Q40Z4m7dES1lJkAxSsIytyzfEMi5sGFnFHmb/FcKasjCoY
LhN/H/Iw8e3SVHSMn8EtRUP1cLjujnJjqf1Y8k4Q4b6D/9GBH01XBhNzCT8jB1L7
QeYTTvRmGgJQk1NTGxwGEu3p4e+gaTK0Lb/GZqK0NUSgbkpc1z4VguyHcsp8+s2t
N74WcbUiVANlph4KVG0LxAQtMFZFfcnbv/TYckOmhVHqgIUDJPhF8sA0cn7hIrgK
TkvdP6PnU7BD0eGRaXOGXNBQFSLFUZOoRCsY6oeuLtRdhe/lxjPEW7iTdNKRolKZ
8QntN8sxlSWlV4oZI1An/fXJvzjAK4s+Wnzpn+cn0kJGTQZnU3ubmJ1zyjyLzsl1
Md7rWLIQnx+7ts+BBGEBoOQd/FnT4OrMF4km0jrFIbmOu48Eb3HG0yMy501lLdb/
GgTtde7YwQEIK/4gFI08/2yAt7ulnGKdMCrmjQr17khqZ9yJB8xIMkhLqGHcqBwj
T8ldBZBnvMrvMW2D5W5ZVSfU40Nh3JlIsiACdH3RT0Fz8pPHyRkftJH7/94xyEXJ
bWW1DQYy97A/HJp6bF1MsRzhFf2GKPrSA/2ejaQwwNbgtjTs3Hi516BWcKpbTCpz
QhOv7d8VWWgtwL3lv2HcZn7e7YSz/1GREgJ6X8DNPvw7Gdgam5NmDyCV7GFnfaMd
DQsjFQtnfTYxlnirVaOzthtQCjCS7DYlrgh2bD9IuTx6f9JmKrrt6kjSiayhyDVG
vmg56kYCQwOugSpfyQ26AkYQoju4PG2a6nkcH7uTLeMhuHSBjt6BpYufdOGfEYHt
P/UQkGh7nQyFjHyIXDJisjNAu14E+/aQnDu0qUGh/yoZRmAd0Gnt9moD8Ifx+xUG
trEz32JFqmjl5l22WnwWinjpSi3YYGWTiACzW1ngkb4ZS5N49XNmXX5Cy/5+UUVY
P42d3bZU+BtbfW2GzauCaqxp2lQlSUsf4jiIiEdWynYzOOzGU53waZU3ipz7/LT5
wzjich66r49qquVtm1kAj1j4XXaa9hgkasn/JbCNYuDrdDnXu9kypDNrHB486UZn
rTtPND/mfcipSwtIj6LGdXCHNipttqWFMRcTO2Ux3MFxuH3eaw3Il8oBWh1odt0H
rmz8TM7oZv5YXuTTHoHj2YpRo6zCXF/C5TWBR1TOc2D5FymPkDElLS+C6K8NCznV
at32lDZG78J0xIpDVQwV6u5182JiwOAmVtAAXNCkGQC5+tAV3nlFzKI/pU6Xod2D
Sq1UHajLYBp8KU1uCNd6pjTbvsJh5GEW4zO/m1tE62obvh6aGlNgzceiT43+rrdE
tnwQGygOAWB6S4UF/Y3tIXezFFcv2+lEX8Wozil+VBOmurYMwh2WLeh7Cxl5lPIO
XHeN5DUNsuN0ciMLQ158/WrcQrzrRcj6IVqzd2GtPe5nCG8UgBDrQS663XT9QM7K
FQ7gWrZW3YA56c/j221GVDLzKG9Qvx0HbOw6GPfyIpROXQfSgD3W2cgCFJxoAYot
1gbDFGHpktkiJ7zRZZqp8g0CeMDWru8MWKmaHudfu1Fy+Lo+ASdNVY1TtaPSOi2z
Wpvuis7fvAFPWGEtSSmUHSPVmXocvEjX1E3CbnVW+EV3bEnmxv6JOdzVN58KGNI0
0sGR+uS38Msu96W9wbwTG/MLmFcK6Uog4qZdFl6dg45PWOa92qbag3YO8HR0jXTN
nLeGqyiLciqSrgwmuQkA2n9jvADBBAymJYHp+SnTS3/d6SeNl59Oqe0oiTs9pK4u
ODC+dZXcmiDe2lMTyM6zp5ofrlC3zIWkbXPEkmxE1tOSAvmTcW5qlyI5d2PWOwnm
lC/sPWvFIqxPawa5zG4sW3nzp29PSN5iHIeRW7w6b3fbBcTZseV1AzaeAWyUBbO2
vSQdKifFNE9n/CfoLjtgOEylykXZjSq0AWwNCiOg6PEC3eEJIXeRw/V7v5hA36bi
CI5cnJMxVfMXDgO8YOIUeye1+n+yUuyZ6zcdhYXZ4ACzALRmiiWxFTnSXJius4RI
4+2QnGEl1jM3d8Qsn3DmXBe/PXa2sxJmprvzBJKt1S1gBfrgnK/OzV2AtwWH4+a9
c1CLndaFldjEW4QGV9f70nbXBEWmJOKgiVjU9ylTsfRqpTGTS/0zAg/tFvtUMBEm
DTH3a6SEH6aFkOA0GWAWz5gs/BEWe+n5pdZ9B3gV8YMHLKWj02tsIyssrjywYi5w
dkQfkRDZ8ErmJ/z2Y4jXaCY3EQnJ3P9rdma/E3ZCzHX0fC3RXeWJ/Ib0SduGEA4n
sqQOMt+5Y8fY5JXdpRV9oVTEUU5gj20fw0kA6u1LQ4SWq5tk6LKVjb3QewG9S4HW
jJQuu4zf4WUXghZ6JRbKOJwEBf0fFDbveN1FVv58xfvUk0y/mmjZahNXXlQSqk9B
BCNUkapQgkBYvNeWqGljAOBrRQQNx+UT6MxQklUK6yPen8JAJ4O2QN2OxhucftZx
lGKFGMU6N35O6OHsIN+nMRpYp6umARQrhjn+fuJvTuDHCc/kcgS4BCCVuRqYcgv2
jWFR0GH2CI0oBgkXtYLtxFKoMtAHlMGH9X6CDOypK0Aiveq7+fA0H6cLICfpz5st
unZik3mIWx5rNnqUGcp8yHZlVzcCOk3qvieYnP4zO/qXNP4TdYL/kvbZiuSdJhmY
+iq3WQMypxpxlRZiojOgYf3pDX43/qIam87OqELRyw6ouVixy1A5XqjduXb1dLqL
WMXGnE3gSYZJBsAA0JIQNa0y5tEDTB/52KJat7vCoL7kOMwT9xRXMtIIOqvjHc33
9eG+ybztvqeGr86EN49iDC1b1Jm+09yGlkY4NrXhO/ccMx5iYf8lkk4irTg43I8/
mzz6kFkD/Tg5UHonMATsZjSIqTRUBsRiXhcJw9bYnX283rq+9vfhIXhlsZyRIKrI
y03NdZdd9ygK849yWhYv1K4vm3j56KntXd1oDi7D2MoQCVduwAgUzPoCpFfwdrVN
Sbb9NbYfp5wsWB+IuTH5LXrU0vl3BdHngjPYSa3LMDmiakR8NPNHnLSZ2mWzXxS3
SAXlT7YwP5ZEf+D4fHOOhc9dpyGHuOGNacRHf4J0Ex0ud4750uM0CjPXhkb/Ciag
SbyqnX/iTij5v9GpUc7UxJEswK57qUzmTE7pM/8l8cKXEq2KxJZUev1O9OmBewjB
oD7MgwFx7V8QZNS+89F6UK98dcyPhN04nDRUtJCXUxxhBjOmJRY+Nt4NCw93Kgj0
bAYLD8AaMHbKHzsNu5tAymA73Q0qlNMil7cOqRrLU9bO70Ekfq2cdg5Z0/iSCMGL
xUpFHF4NCXIm8oMhIeKsdVK1uKM9HZx8Lf73QqJakLK0rvIsHJMvZPXBjDwgQ9el
et3XhHkcZjMC4mukdntaPA1uOzxUXHzRDdLHLPj8tpiFaijhzQJvaMylubs18V38
jUmRc6MKzygztfp119aCEPzs1wtDWpa6tnklv1MXRSpN8jBAjCpvfI1d2bf85Wgl
oiD+07F19xaNghYlu5Pbw6EbKOZWasQyT60UhnOZZeR2aOIBAA/IgFSJ9GffVlNO
6eR/5itsT+J7BC2Nrv6KLRPmc/LRrHxBXWL3GJ0TTSqQwEdQBs5kCiEYHdIZjJ6N
R5nVSuVh2ycssWD50Mb2iy0K/YVQ8eQ1TLXFYLy1ljH7A/HXiiORQV7Aay+vg7qb
q8bHkvXvOs3tMT7PvQz7AXzioMI9YRG/5ybullkeNDHGnFmqEmnILnqV4uRbqvzC
PBhLF3GRlRtATzB/EMUn9CeoYhGRaAoHIKfvwHGbZZaeaGFhhuRXfHJg9ls4ZLKI
9p/4vs05yzddeGl/AW8hbfszYuPmGrjuFDwK1+NQeL9XaGTMcUWagW5GbDE9qukM
sAMLVuFIx079z85Ipc/GS1S7yf6wXiqcdL6Tu/VVGBtUpyjCjnclTSpWk+IWU8hJ
nl2b34zGKnPIGqg3yGP/3QpIO8ad6dQowWycUNgORcvvI65QAZ+vFMxTDvRgsTV7
tIHmzfqPlhIOBGy33m35yIi+YTpNniCPQKf1tOqwBnNuLZE5JdxXj/tvfE244sKN
m/bJxvNryDMvn9SUlgAbUBq6/aoCAmI6QvP9FObWwpn8dYxu2tN062ACgla8H0g+
Y5lOg64x93PjUF1LL7/AC+hvVClw5zPk2OoZ3eTp2sZNfbOek3o0a1bU7mayaoIq
tCstbh2r2vD8HcDonxhCo9CiQLapbh+krCaxW6zdjI7yWPqHnAGTeNB0QGLFlbLL
x4lnn4t4XnQ6QO6gVmbbvA8sFW5yJG06mzC/5/vqTB7NQ3qJmAUQs38HHCDAwhFV
CEFnETf3X0AvF/ZS7TN6GB56r2hFdF0DeuTdQJoVTPS5IPq5JlfyZbOc3/+0m4be
Sj0J2OzTzI4c0MDoAmCOn0vYH2M+i3/gS27nFz7qAo/NCJxPaLxuC5SatwOIHtff
ReDiIxgIFI9uz9vEOnebBlNNdldZx5XVLwc40Qqt4u+f4sVIcytPDw7NesvlOH2r
GtPF5n2wSDbI+ni3NhiVSeUTEPLGjkmwA/2zK2SwfANshHNwlkuCC4RafeVYVypr
9M3MTMiwH0IMEw8Ek2jQ8uRhj2+ogtixMo1/EcYJPICKlaJbfMLTNLkpFjXhxtS4
dG5gxTSVStg/uEgjfes1VOYiWVLhfn16c5yRQArKCN1Xb01aVBynYCBAtL8tBGHD
1P7Rwge+0VgZeJh8m6PZRUktn79Y9MBaj/+s5TDfEQQgpQ1fh6kd+D37T0NWOffb
qkjhrjPJVuA4Bf7/J4Pr00R+Vf3hzTAvfSE4iOg4eG5lsoSzfa1llN0DVVD9GbTB
LJJtkdDzURmOJO8ViHdQQFeWmzmmaANAOzG5eaaovitKwesYsEXBt8z88/lo3dUQ
OZ5VcmkTiq+Y/vlrsLe5qS2Lr2/s23ux/UszL6ffHThVtyALPgQiG7bR87PSSJm5
64D02m3Wak0a+Obp9MP6SrPEMjEBx6sVr1uMORgfpCNcqbN7Yt4YtNCHZ/rlpCQm
uNNt8e1CXMug4TsMs+xY7W7focLUqAshpOQaXQql8Z3faepXqYts7BFOPRV5OcjI
c1jejqT++nA58DXJoxi7Ml0poqHLbU99a9nXdApXXZYhZ4YCe7+dGP38DgPa3GSo
oNnuG3OdIrRVflJVhs0dKf1UrT59KTkcPe1r/k0DKRRUY9A2r9MF4KwPLSVCU7yO
VTQtCwHAnfVo+KPGcPEwl/pTfGWGXvUal5cIcswZD+uXz78InSAxEE6HPu8Tlw+V
VexUessjcDnrsIcix+YngTeeJT1/59LZeG+WJaztGV6l5Wp3BLT3L0Xrw6SpaZpL
9xDibPUcX+t7lKqn4Em7qBlXYh3eEte9njU7qUo92GkJZMYP1LQMG6xBvFu9pTm9
vuIBALWq+txa07Pi7P+7cvK3ICRtl7JyVKZajoBdwEgPlkPsK36wl1GA1HhwA2Pr
aQ5MewN2AbEg7uu7U3JdjsW8QATbKjqa0nr1k46QYG1voydg+ImhHoLn/eHYbmLn
RvsiXUYCIwLss0TWDpvAKfsXTTVqnzvbCIvfoqFQSrfWUcvaCvMXyPbrxfhy8euu
slIdPEaKbgN52rqZUO3GUwYAfq0QsPuyUkstp6VNneK6+NYBwp/wssegUczOOxbE
wPi8oCd9uuJqygVymzXDiic/FJv0bbIgviRAvjum+gajUhyj0CQO4SGQ2P3jP5q5
ypVAgGGcXE8C9fRv/jzcY43/UFx3qovZW0LlwEaBN36XgULoNPJ7giS2b0p2nmFL
kGI4Pw894tBHfdLUq43+dLnESQ5Ug5a47unP+0qngwZoreD0+z4UguQjblpJ3Ltp
w9E05JO6RJYZhGvTB8jWOTS344LBnjhUfwJeVeu3WqW3M8GmuUq1/y18yNOyDvJC
rTTKI4XNhhMgI3uTh/SgfMyMGUCtHbMdq5YE+U9o+ZTLWm7GprhQMDTOUtziKXy6
WOwRIdn2+GNjZbk2/ClUMiC48iHbH7aV2KPWIKEOXd5ymGjTVbg4/YhJijP0UF38
NvOTz7sTQKvB71b5OrYj+vbIxmQE5zzlNJWjRZuTSXlbp4Viwa1xlzstQPPvOxss
TRtdo9OoHNuSR9203Va6AVxy3seFi9u9T5i5/JqMMxqqaIS7a5ZSPeEmb6QPSOpM
1Yu+uIq1e6WbZt18+QP/i+Zj8xgeRJwtB3LlnM7RYdDDAvXiQrr6ftb1+qGygEka
K2Z/memwsicvzfuque1BHwf5Sf47AE0zJz9SnnerNMzSDze+9iLrNl2ci1o/gslN
boYojwPjy0XJdhMBVKzikwQJ/Z8AgPxcOM+WgxhYeMPLQHq/VNVmy6eUdUPd3hM5
KsmQ+DUiFPx0eB6cSqmpkixzp1RPyvH2sf5Vh86GfhR05XjLm+cnQVAOT5HHjv+U
zKWN1NK/zqeyGsKCBI7HgbW+nDazTJpnetxKgIGShQXNqPTpxt74sEU9uJivxZdW
U6LRfkJaMKENnl26lS3R93AAhAJQ3usTpXdr3n177a7NWD9us7QVkcy2J39Nmn6X
uXn7oILtkRIo8kbKq53qVG6yYTMWyHZwEhvMJywMcqFAmrlmkdW/zH8G6dOnflU7
qzlp15wE75Lae7mFIiCziA04XmI0GlF5FDYfzI1mvVGD4/fkIjICUyQIQXR0CCcV
95bAyfadUSs+9WvKyeZWnaP7v9bKOe3dVhFn2yX1cGw6m5RFKrzBD/orlVPEiD9t
MnJTS1mlwOzmKNNKEEBFlT1tTRsaNzjvBcP6DruI4DA1co79KvCNa0aUcHPpYX2C
RZyFWGukyg9djGZGluoSujmiqOkAyKrX7Qa9YmcBDb+oQo0+FBGFPxwA564qfuSa
60TkrtQryQtPVoj1zb+x6fqSfXzD9e9izuPABv6fj2YrzWAPFCK5DsmGRZclu+yK
Iz5YJoSSdrH0BLFPGovbkzqKyinNQu7XwsBQtIFBQ3I6D2qawlwxzIFWxfFh9KXW
K4g+/MsLbVundFTAgCNi1jpFQdDWObesZISjnZi86rtb5r/txGUldDwULv3YcRUW
whnaCbNEe4CB8sDD617u1NXh/hcZlnddJJ1giiLIyWmVbMWOUE0hJOXe5McZ//TK
3qT5eTLxlmPLwiXFfyW6tunvHlEkGxFUx8nscuN0+Wj+WPMlIqXb5RR2GywWCLRV
iypvcwgRL+Ay/dQXsIOTB2tLLUQ0vFurNgRbgd4gFcw2XohB0JJfBEtUJ4jDQosa
LeGWcS/9ZqYFutrHsSYS6c9N5tKmR/0DVWcf9AUY9roArJ3c+Nlsy9Mqh0odB1Iv
n5VxBlZLJ4WKULsSkCwxubA7boNOmfj4WsaF29xugjD71zbxYR9iJbGNh+kRVqgB
F0S+DvoVXIDdXu3atPKaHgnD+kvNrQsfgEkfX1VQvxjUoFjfVqEc3ZCREckUHHQV
r2jqiDvjAPO1M0YsZbsbdbgCBhHx3tFQtxID3QYiSQiOqDUKX3/F9rMqRQqqG9FP
fZbcOCnjILlUpz+bz6AjaahfS9mM7S5X2ayiG/s0y/dtzjaJqY760ETJI89qLn6p
N0SexdBPZaHuo/vDYy2yPrpFbjDHNwpUtOrz/5IzAg6b9onP8bPCmekiawUwdxz5
CTGC37oFf5mdXTtKsI1EvhEKIkbJnJRR0W/lZOi13gI9gV35KeISrNjrPaL5FJVY
QZSqcOsbFzTjMXXvS6w0/Nchgxa62ghDlLV9yxSwz7x1dBAI6Od8IHR2fCoI2jlw
qoMgcpWA38KgTgiXhLTVSA8a4WXxa1BkH6fP/LomWk7FpwfO8W62vvG+124QALaE
GwXwIRR3hnA7Nb/GZwT19FxuigTCRXTpuj3cHyb7pPY5tm1ZxykfvKcuTVsgoJA2
LtoCK3U8FGmWrVXlBMid5ZcyILbSn2RxjncLuGau4dQtky+tTVYFa/8uLIDGUlXP
0fPB2ajEoujJXXYzATPg2yTtldzpfpLkLLF9dZexgDtjAqYJncXrP6PqfEJrkLvZ
fXgan/FW2caZkivwNnaooM4M3SmPFXkyXBTcqUVmFm8ZfcV8kysC9k4QfoaruIjK
xcQIGCZLh9OTj8mWX85wo3XNs8/GqRy5aMJl1DJTRe9C+a/l9T3kVecmRLoKK1DM
/MM7ogbcyCe2ThRANGExh2HP1J/tg7AF1mOjlQcZD9rSAFJmAk2OUFx3afVi8W0s
5Cyoom3FwMLHi6STUA4ExamUt/xvGb20dtiNBleErx30EacTNl1PG7AFMNuRrr2L
07LprV+nkd1zxBQMz98Tw4O9GOD7GYECiDeLhWjc6cRuod2QshXg2yCvqe9GCC3v
WSD4pE0Yat+Hmkd/rKqIAHbpceNuasV51KN9OcHxeVOnGZUaSM8nEuceMqcbmmxw
7v+3LGWFKaxlXTRH5BUwwaqN+znRMpQXTa4Wd5nA0kIbIivIo3/r0znVOj5/eZ5Q
Xm7GpAXLh+iX6VKoHSnEe1DD72ih9tk7X6mi3PAMLmMGUotcc/gZfWR6R2NG8e2c
rV3op7HO2V8eV++wtmGlioHjexmu+Mq7JUxJF6ivxqK68lZf7obAdJ94NwQnobWt
JrgNuC8c3bwPkDxZQwuHRh6KuCuHFTBCAHWfjxrwoniyw7YnZtxVu0oQU0/zJz0G
xmypYRCbY/9elE2tV2ppxFXyCPdylVS1o/C2ypepTBcKgexxJRuye7ZtFeIXUqdx
yRsNHF7+s9By29zVa+RUk2G6st3y0/4Sj1AQQwVuaUQKERITLejjM0uRJWy5KQle
msYyJXT4DiDIPhwMIAmYH/bXBUX4qGmsOvZoMypeybM833aCvjuPIu7TJKoE/85k
KmWzb/YJSlTxT/43/KnHvYRLlUBOlAP+4pq+veTStu/7qWNv9MPn4n1YGiAGOcgG
YL6A0bU0n+tGMZXJ3urIG1Wl2i9/1RYiLn1CievIAtU/Osdc8IAREGyAJHu8VgXO
mxDSGmOZ06etnm9299UiG8NmjvxZb7+G4MbRVs5yXFU2KK/SoouB/N4HBYW8VmcS
v9KZDyymyzP6kYnEqWLis4rE0i8DoEQCG51hh47p1QttENDP3lXW7U8gaU/oM/lj
GlAaRRQTgyEXUQp2r2YJl7/GEhuDnU4B8iNCK3Z3NCR2+J1p3pzK/Yv9moJxb88n
rltIh3k/TipEZPcaLiFfzxcFFA60xHjsb0ay/kl5OLUhyI1tJeK8DTcpKugxfG+f
vvfICZNi67EthLt7oK0TejzYM+92TQdInWX87PQwaKQeG6p02MdGIw5dmi46/8zN
3hxAB2iErfrLk/0lM3dR8jrjNtWg65ddqZWTV4/I3e1fi30I1YfkBM3DAQNo+9GV
bDvJ8nxdvRo7Mr8fVGqAOYSYZNEK5peXZLIWCzAIGbF0ZZ9hRFRXAWsUY2xTxDYU
lpIp4/2OVUuUuVCuW7nOprh75gHeWklZcxiYwuxg2P3QIdF92cDFs0ZHQ3GPuI5W
T1AYXyT4HWtBEGpe81JIEk+Mwyo3V9e7lvRUdW0BeB3jxGDyJ9G67+p001bO1gRX
WXhKf0bCUJNoQXoCb15AOUmi7e2MjVZEWYaLlVTnrn5bBlOve2GlyHlI1vKWkJ3P
PMd8S05/jSe0mc6DQX17qD7KWLebgLzNCefCKu50Z2AIJv0MBTSz/jHqrcdnM3uB
fLG5UGwmPIRortHEvfiepAIJ6POdbB8U0zvNoa+A3GuLGpGspziSwRkM+6j4qnGR
nrwTvikzJMTAPBrwN+j2FVibd6l6OINZbGnlI08c15wf0lsQGZrLqjjYpk69NCbU
vbDJzh5j2Tya+/OTrszCBtPSYXZtmwIclVZbe+C/3p7UN9IXOfz2mFPluAW4kFht
yGuJ0ZNlgBbNU/MOh6ZnzM+LKyWtKdLSuHjh3DgiCyCBELAjkGGJ7xnj4cGe5u7D
Sd7h1rElEKRMenq09+179D9HWABCB+5WziyWoWb5nG/taBIZwGVDlbFoxKzHrGyK
ZjSL75cvi4PB0v+ibbHgtWnMrxVrlo2T+IAcuqTezEZe3iDpV0Bf4+k8YIi3EeEB
OuhCv+8kmF5JvwPM0XamMC64i6oOuRABLwJ2K7uLrv5GOGD5oJpZU/SXLHsFlcvp
A3v9DJzMwGU/Ox1lD3OHPsbxu472+uWmPREFMkT+Tezf2/7elr5dHjbEIjgEpVoQ
3vg16Bp+aVLha5qgrE6w1Zu0iH9vpfPahSplhvIvkm1LVFql5ZfN2r1iUSqVJeob
rtmOmTGb21kl3B74mZH+QYM681K81ZqXRmJsHbdEaPUXcaSTkCMiWVuyj9mwAH7Z
RFgLyqsYtLNDLKgypOqtTzY1quFQVxLUKbWG2p/l4CnXxviTyF7IIMB0IDxsYrBo
+4lNKeUcl1Yka9gCvIAY3/XrqWWO2d/H0+ItAMBb+b8A0s4RYv6OpWS37w5wfrom
X77Ut4qTumJCeohvMsMGjUeCXjRjV29vxmCLkdqYS3ds56rsIxLlrHHyb5+36ywu
LNuy4XVIrJAKNWgm9HHz2OdfUtjNC2M6kQSA11bKoIfvJs1a4wvvdvOpYgluJksn
Pp0BGzqUPwciW3ncG11W3RWtZCtqJBn06vVmQ/xrC03GbBzCMfv/D+p4DHWqm87U
oZu7rNVUEVao7QJFbsA1VU8rQoYWryywEsvd4pezr5B0/7fFNX7ssYiC4itz6OLa
AVAVKv/Xt9zlZOexzHxNbsaW+fIpuu3zUk1F9kTVUf1E93NcobDMheo5fqffnqKG
rIt6q/7KyptSDkR/rOJ1fcknw4wKDNI3aA0gKkOnWGCUuXd27PCwqqDnRkuVumdN
H9C8fOqazUMXqF1tsN5HHTiYgYPSXRZSEYGKTI/9sdx90n7hzhpJkrtXggk9WPn2
JDR1TLU2NsOT7VcG7CTiWWvfmVvso3leceDB2mGF2bEiN+qUgwucJeQF5pcoZC5Z
1ZGeN2ZzuMMdrfmfJWCS5Df984ndcYZ80fWLJueLG6Wdhnh7CannB64ahDH8UaLJ
LNJqCQVPfxGlvK0vNFGOjHxD7wxifvU50Epk9TRGrWyi32gT6ur0YI0S5ePc0RpZ
JKNo2wsSEmUdtThkPlV9uxUODW8//H4Phd8goPQYRSePPFrVfyxhTWpfrCH3sa7J
FS1GjWMmTR3xeBd50oWhAbnDg+8V0mY7pvl9J5zLg3Gt3mXi9YSDGWsw6OqcgdEe
WiIMSmtSpX/QYUAFvtA1ojwQkWYcPyHlTQohldRk0+jlGaYOncLPPGxkyxBuC9VY
oVRSn74Xh8E9Ye1GwwK6bRsrdM4dAcTft45wbTUN5zHo1KH5VqC892CTuBEDTlaa
nZm8fGHyzUjljhS/wx+/H0+gnIoa5E0Xt1NxtecnkhK797XL34jQrDixvhVoW+gz
MYMYJncZVx/IV4r/YFLjuM6NbPwYzFA7l/hrk7oOzmKkpwG5yBn7g19bOfGuPcX/
5nP2pw+j2IukX8EIojfKemrBpgjbF5TIfShcKPlOwVySeLUVN8QppeGqzf9Rg1eK
faib1xIjYn8ts7tEOAy+VpVtZx0E9r6Bs2R8p6RikhLipLXtGDWuarqfrNU5T8Dx
PknsACjy5DPtEfpLAZhFrLwvIII/B3iQ1XEvjJQVrdaIMniGK3JG8nue4CAua903
jhcj0kq1yf3Nal3k+6C4utORaqokUyJtliPlE/UKrvPwfPQrRwaQXgROrRVtEw1s
XDgEbRCFs5vfPqmeYkfcKBjx46Tj7a+iyOfYYBPBf42py0jXRUM+7TS++oY4FLsS
iFSXtD2t7Qh//ccvzWKR3c1wUnKfq8zNUj7I6wEcBHb5R8PIxqgUuLxkEVCPG3WF
uT4gHaufAXfukeiG77mHN31TYgS6D9WL9lBXeVYwKKZz963cMl3R4HRf42izttMg
DkmGOIm1+pDNeou1L77gCcS+3U9USk2yYp03D+MrHgUtDxYtAtA6zCS+5SZ7KM79
fDcrU8sksJxWC+BSmEw5tJk8POWgTRSEkOwSgCN+GZ2Aol0tCQ6iFAc40iS+j1jl
FJlZ38W01OT80qKzp9/7EWm8403PY33D4EW23U3GXie5HZhwBehsH2FBLUBAkJhZ
3RG0eBuBARAepJzfzI2XZejSzcZ/5sqqL0ZDjbV/xAJ/y/htQZY19PrW2IqAIu4a
6LqoOPzDelY/JqpwErFsB6fiFZH58qsFOIEjIxeeGE4LOzQqW8Drd4iDNaZoTKVb
GbNOSmQsLKX2dJeiZof118yG2k8JgvA+MhV7rQECwgPAbjZFNUHtY+otiu38emzE
NE0Q9WekjBnKrtgDjzq0daZxebqu2JKTAWrhjdfoMiBoOIG4IX9S7UihWVYNtASm
s2QcXQIWPG04eXnzDxAxZb4M9UDyJU5JUhKLU9/2KT+u50cl7I33DJ+Sy1V00bk0
h7S9kzPsyTm1E6X0jIoueGCPkAVARYr2hzSOLiISPNPiM8FdlMsrwkx0IYCRvQRm
JHnkZ+FPkenYXWntoiwaX7EKNtdQhw3d25+IVPN9boBtIO721txE4yFbBDIhn8zU
UEVDTxdWvafw2lVUP7sqzc0z/r3JgXmoaXyrsvFYOB3Bj15xv49l8n7fA+lb74sI
mRsy+PCE2R3Yh1Xq334BAW8TmLtIk1VhKMqM6fJZRQxlqhS2HaJqRmpvI3TVpHrd
dAUOkb6b3FBkvmOFVX6ky+vgn5FzmBUJZdTZtPbDIL1xVOyMhUmapwNU/9z2MW58
X0GD0NtxDNtJEyDakfQYUDIpsEbGj6RLFYPfHjLSIrZzcr7gwqg3SqCEO3TNg62q
9UvVLUNnqpJx1JzRkzoXhHyl85/ruQ9Z6fdN8diEFdGt+cOxkcPDPYFnDkKFkcv/
bV6CkZWrlSp2tp06UyfYv40xt9bOCURrTURLF8mO4lyV4h1/uL6XSxC9Xsy7104V
yRHBmQz69M2hgm52Z2jlODXdHBJ85VJk4xCpnU46X7Df2+PATLTyUrZI4h2k1gRj
vJ3eVt6EKTJ/cO6/O/LPmo3JjhAc4iJbmZJWMN7qgZ9maQ3CTeEULu/+vIaUTtnq
oS9whvyM/88yfb3XTSqNw4xw63HHuzMbq85nxKhjt2A4wJlSAZpIHftiU3QjA5K4
/Zjc6R3Xg1J71VDae+TtWJoJWyTzEL4E1yZ/MZwBfP0Jvw+k9DuuEUGzScd1jW6l
v+REoETt7NDhWZy86AfI/uC4tqR5LXD6iOzXUfdzx9DjcRKKRmB3xMR3TMHJgL23
ohJtW0yPcvr511fiaEzFQqGjTOeh8BPrg2B8CMovMwQOgRItXatVpThMu4+TBfG9
KfnklHeHf9pv9iSb7E9rZcvJ6hX0T2QmkFs/ucyvTRUIkIpCmAHNHSKYlT/ix5qx
6tj6jeP0sf9RPVarqckAuKE4NLfASs2XD69tcOVD4cCOSHuzJ0QAciKO/xhK5sZT
SIJ2XyzKmW6zozVg9olJZf2MNzBH/Q7zm552UAYbGLNMnfoPhmLkeKjP2ZqEVamo
fqP2UUwO1n+YRl/mM7YUL+kRmDcYIm3jl6QOOip3PZ01gj8bFpZfidB/GhWzO/Cm
7UgT3aVuOzQ7xTrqdGTzv2B1DeOmkx//byADUtrI9fHKzUxT43TLaWbgj81vGZkf
8HQVzPynN0zZ7k1GqIpyyVu6tDwXBJLQo0xxEPa0U3tjm5Qw9M4VTnkjlDSu3aDf
noER786GIr7fGL3QbbP6J9MjPEqR3ZAdMiVloAlriNdRnOM/APQzmSb6esutHG7y
e5SGwW2pu+UMMEylhAKf6Rv2erT3h/pPW09JOBgVNJtHioyR3TE7TJGee8Rg3b5u
/oR2QryQUk0uHL0Q+/gLquCdWGzn3/YjOb0gHjULOCBKjWsY1LVHU56zG+nk6BOH
URkavhQawrYOG39qy+xqcDAPPa9vFOYU8a/O1dbs6JnoaN6VUVFRB4CtPmBN+1LY
FjIvA1sTCJj4G9M9vQa77TFyVs1/eub9+VCg6QgEWkDUMZbxyd7HGxK2duYSHN+j
H4KbeGJwvoWCaVx4CQ8lTrtLvAZjJ9LFgoiS9jWCOLGfQaVYhoWlQr+D/K63xlIz
Ldvp5/XwPp+24xl+WHAEbSxCUx6IH2kE9RO1/n8GrRzAeoYQ7AcPQyp3itB9vD0S
t5/e6p9rSBayip0qSFD5rj+vRkjbqLwvVGB5lAFibH42qvMHkPY3GllHvJCRgzzD
MU6UAQcTRLY53gTP8UfFXqI7SEEba6GyPDzejWUllz8iyJLgrhxbjwNxcgI1z3m3
LIw5augM0VY4fpfH6o8lL1/3g+1aAZsaz6PeRxJKyzqzZwWk9nMa1TzNPawhVSYK
CvtiyV0bDBZmz5tPZrtiQGDj770ffb2HpLTmf/HndJzO9m8PVUNW53mBe2mdGyNz
6Xareyy/lrh9FOg3S88x4UV3MSA49sa83R4LaCJDCwnUuUpIk/akEMH14DVvDtiv
fiPdbEPGM3nRpoPYsgyzHQBVX/UMkvrdtO0xmlzwD1RZtzrc4mVVqYPG/rwn8zlp
shVqhsyNTXC7srBljBIxyNoCpNadfFHNXwalF3C+idqXFP3VT41KoHktOznpdxXK
jiR+aCNAkYz9creSh9q9RJ2FPWL7+BW1lxi6+bslvG47L3KuAiSm13HpnSsN359m
uwdrpuj+sjJwVTAa93yEFwmHpjkFuSmlqhgzntxb5GTJQlx3B4ODhafDVsckTp6F
DNSk6PIYusb02ZFbTU9mov0usDmxFe6cKLXyNK2Swmv8n5gK5rSfvUjok3ytzLC3
kxBdZhYyhZDveN8LQ1hSM/lXFjIww66cIoRrE5p4F0QoxKp0znkobBARfb8BkhEB
8VyiwNycfXKOwL4y8cKbk65Lb+jemCdZPhLfEmDCUTol2Xn/M1Izg0gBH8Up4qj9
y99Xs1uwDfHAaIr8EDfE8j8Jptf8m1B+i/tLPS5bHDWIIYjW8w704r4WZxIR0KcI
yEI/M4P725zmvhoj5PMCEZk8NoL6ztslzGnRVAa1X3d2RIW6l9mhC0Q8q/mXp3MU
5nQDqiMEMsJ57MU6O37PcK5IFRObqxYYvBOfuq5B3gm7Kq9nFZGoUQoxsx0DeHUw
mn92pAk4uQZ3Esut+XOkVLtbV27FutX+r1dzQd/fCwsmpkygpYfFzdUYPLxtcmHn
9Z0r3P/w4NYJ20aIXUmFwbHSYJ4a4DOxU/PyhzMWfhPWSaSpYlspw5TIkqaMdWNw
HZAetorS912QFjnUoJoD+JoHU0f/q7fUB9kCdJTToqSqRBGSmFm15nFz9P37egGw
XJiJdB0AQvPF4NdyAAYyh2a98hxmyzkXyirxYjpONnr5KwqIihBZAnzKSjWgi0Li
Hqj3vKgnOkmhH2bYC/s4n3j0UAce4HH7of+OcQ46Zmi8LJZ9WXChOnrixIGE1VoC
/jAXRTZrjesxjsf9OzgcpVcIKyTN4p23C86AEf6gbuE3OR/TXr7tNUfsu0EdUkfK
kjuFCTKnBTGEDu+HMe2bQxhHFQgeRqXsb1hF4+V1vFw62DLGcdSFZbmlhV5JrMto
kVl6pG/mWeIUg3YkoEzANW2jA3Kop0ueEn4okYFSzNrXEYl6GFce5XQMgud3oUG8
5bdH6d9D2g8yiOgVWWeEOKoSOQh0fyPTqhgZYNvXuY0C0wUNawo+zU6dIys9fR32
lyGjM2yzIf7EJ1JjOd7SiWIGcf+/JVstw+pu/zBe2p/381aUm+xRgPogDsiAYGU8
pvVdiUo8SjA0gRpGQPEweTJyiMqwi6MziIR9UpUvRfHCa6nc0s9NBTac3QieCn1e
48ntVvCb+pkF84VMgGr6PrBC2ts9TO7SB17y4wpTShvZO8cZ7yGov0cYCFkLU9Fe
zQMdvb72pmMUObLV5PW5uu59bHlcbrdJR4R58owXPim0/OwAb3x2lwHZgyBgyBHw
AN8SeoEk9HVOXYQU7NPqAdwunboP4UO0ndaZmoTmWYQTr9Xh8h+fRaVvUzRClgVZ
wCt4XkH+VPsuqjY5CjbfhIYjoi3TyI01hEaZetExnmyEi0iuepnjWLjrxdiaAGn0
PQyF4i1pYaLTiasbecoMkcAnYBl7/YEldEehJCfuWVsYoY6nwe8Fs+Uh0gnbwmet
FamPPEeI4e7EdoGkvXAljUfIEuynaKfK/YjfKL+v1K+Hp6LPIPbYCbVFjd0fllNW
U3HNTcHukdVCj1VaLOi/DMF8CIp0wIe3GJZRWp7vZhO12HrTZnZSClhqJvAQpz1F
0/62oeuea+RnEXJttyzK+FTmin46f/yB4iUDRvLicONCIRYgxzX06gkm0tdTpOls
3tQ6DM0TVxQbIHDdUW/E6esIcxoqXp+gmDWfT+13RFx+dGAV0dc4GlZx53CAnJSn
uPcxujb7qNoJ+jY+Iey2+apsu/DOlXceBSR22WlHsQIb83hQxNalWm1CSby8jNOh
gQmI8jyohu3HK7l5maijFR7wzHrjg4tOhyMObXeJcPjjapj5nMb/L80GboSe6+N2
IiVyF5V5fNAvQUNOgIjmf1jXIg/TfRSOgd0MGiOg9LXDXPgKbMNynqSzReL+va2g
VchOFey4f5w8MCOrVGY9cnGGgGRuke1Tl2D+XbxkNM/9Fp3iiVA9z98ZY3xW/hcq
2wCPMg3HfTQxxJ6YJ860XwsacHmzQ+CN/2o9qYsEmuVpYnc0q4stwHXtETbBxxg5
b7HnnzUJmwT0jsgh7DB3LLlG3bRS3tGzT7UgJonfnlxnSJAZzk8Eb/tGPrHwLsqX
VGbSaR+tmrLQtb1xSv2A4QDFi46oPO2Lk1BGIQyhj9Meh7WuO6L25yn4uvjmtlve
euznRxcBFth143z2n+/jOFyIWYjLR9wWMy9uQ26O7xJ3vSdHugpj8FPSQ5x57v+O
hJwkTaM007cW57j0WnIONFXseveJQfG7lp7jUvFhQ/r+txrsFy9mTGU1F6xkKwyT
zwjZY5dqo4e4G5IKDVfVmU5jnt36CDnhSJBizMoU6rCHnugw+QRvBzFXEcb6Hizf
1l2ccTmxjS6qx4Yc4Em+6EZE1C7RWWlgt3bQyOg5WuO5wpxvRMwRhyEODChEY1mj
FiI8fW9yS1hUPfTsmqdXgqn2Emzlzpibc/FJypuFRSoAKL5jRlYp+NCL2UAHSZXA
pO4VcgcxhFygjkwzD0bSuTr2+Bd1S1Ad/Afzyrw5cwNuKfctOMgoZFGBDKL0qPLH
VzglM3npPnsR3a6+lK0okGGFnIpaMfpAsGR7L7wMS6Lc5/UZDRAgnfhTj4ofn25S
Fjq7uCiWDjaGYgoNOVMikT9nq4nGvFoyqh5vkPM7sgKUkhwTkZwsWmoCQ4aQeJWj
zkY+bFB2I9nD17fea9b0fFYHUZ6XSx9C89x0BcEVdFG2zBn33uD9OuIdO5KrOo+g
pTn8ZVNcf25oIz4mrL31fOWbjlNntUlSg1Pw2En1mGzvcOHbRWw0IBqgrGcUk5HH
VneZFIvIF6voaXjUKgdiID+ZV5afeFsgHIgGM/6UEtyXhGnUE/k+ORmfTNyuFNrf
iXTqVWgWobmMktu3FfXz6kZhErH16GRrUICg8w/+ue272TUlmwC2uiej/rTw/D3N
WVLgYENKEGPCRvVYp76jJ5ihvT7E9XWsxo00a13gHEfhFSHYBJyC6EPQzbaoZrKu
nklFJSR4NoP7D/bwHju2ZC0kyy0AYnmMszqY1s+BE7d9jvDcsZBYvd3DYihvnJCf
miTuaNnDRh3MSQcX+X78EqVQWMhYj0hIje7ERheFxKPoOyfnAC5cp1ngfpSvjqGF
WTud97zezuXnSfcAF9EQlYpmMkv0lHIs69DXDTPfvWuebwKboJvDwtCYjdO12KWY
G1pho41GbrZ7EprYMl59DMEwTbiQWwsowEDGgw++sS15R+J56Z6nHyh2DmI29ar8
7l4RGTyxgFVr5RutlxXSggYo+WS+9etEv93LvgMpNJ1IJEmJ/djsyREDps8bMU+j
s9w44eCCGiQivc2vROKjelqyhrjJExtkB+LHKh49HCputZ9sgzsz5paEltBnJhYo
8BhiXF1W3srINYYCS/AFX2ZWnxTFD6Z97CD+8A029HpFaxcbIbkcCh6VLourE3oK
YZrgGulPHQz+t3VyD+g4IxH8WLz/vG2q/fmBvT95cmgQH3wPZBcPghQqFFEu43ZA
DLDALcKbOSicKhJGKEPLtTOvo+WGIDOzM+mfHnBFkQ6ygmng11DHctZjAVJlCW0F
kN6iXu16oaZxjK5DHxj7po8a1CctI4G0m7nyPZaQNP13ddcnJR6Bw96WQmseTZbr
MHagYbLpYXJozYtcYt5Z3wqwVjvD3z60kMFuEUGTYfQgYLQAsJfZybhCB77S1w0G
2O3/TF80Nc0h8ILwSgW7U7hmT3rimcexhgj/CJXtgp8Z4p7eB8/TkvtxmZOLDOXW
u3vFDFKWwmZ9DIRiIj5T6/5cRwmuMg+FRG7qa82A4MLtIUbQQY3OYrL7mx8pKFLO
/awa+s1hE4yaOSh0l5OCCCnJCsc7zH2LsBt5pOHb+zr+rPEo3d/yJTx2ZSlYmkaJ
RtKa9u6zfWOnVG9fiFAJMhVZAIvSE85KuV3LhcDR20rifd4gH1sSfHDjK32p0ygT
wKO3hAAPbZfPc2WL12ENJ2FnmmjNRnajO4nuiGq/sgmGGALQuu5CxZ7Bo04Rlqn/
1IPpO9jINSM2Rr75NZ9EGLTr4g+w/gNtp4S157zgdCyV5zVX+lrGBurXt2YE8k+4
qpM4DCgUubLQn5C0rBNcVAhoh+SGXemzpsZm5rNbx9ags8eEkVvbYmEJkcGFIKnX
ppkuhR0tqsntJY6lcujvqo43lcGHnBGyQwwibx+EdF7atBBNSrxW6X7ps1IGnY+r
gPRkCYDBcK6bz6sJF/sUVMaUiBAvGi6O32UGG+u1h/OmbJ6Ftb7XiMlWbv5bu1DH
56cycWJj0tR8pSABTyN9tSoHG+QUdHK5L1Y1HNZMFxbVnPwjgQI8ghm9WRiklXxn
L0QJNWM0E8rK/A85P3qYx1jZsQNAmOXGZegxiZyWuvEr8YnnBOlUs+oNKpTJ89g0
VLpAJ75lQIaS6q4imo6gJASbIClqxPA2lNLG5pm3RKrJHh4xtGGDaFqIQcwzGPoV
epVKmoSG4yvXV1s+v1HXpKfj551hpF3kSxSwl2N/eA3taXcs3pVSEOBelwt5GsH1
sFqKl/MS4dNsO/W0HI0MflovbnkLj3qYFP4HsKg79mhH8K4VOd/4UsEYkcpaKR/x
V6egmSQUtbZcTengh94kGyof6RcHCKbaCwI7ome+G/SctPl2Z3ZxvvD8Gn5z9eSg
i4hm1jZZewt0UndQvVDmaHklsMquIICMi25SsQFr6mLHafqhsNhGDymn5T5ACNV6
/uUG/kIXjESmX5GrksXYCepjNSaTxfj4e/DueWA5Z/3B61+/YIH2yUEYG1sbHJCI
C964SO5bgUBzLJfxs8bcb3ksN4fQHNpcT58TikzVrjfMDa4iobjxFqbfxz4nUcfZ
gNCR4YaSf/f4r8JpfUXwW3iHOWYD9z9XqS3EX6pOeqQZ0TeFN2jSgDjAR+D6AVvU
rbut2cAjJ502YdNzf9lVvkZvzv0ZEcPvgL0TjBPh09+hZFik+p+HHtvN6IrTmWFx
7IdbgtoC9tU5IMh0Aamy/hM837TRcbSTKLMsiJUotkgbm33qp5nTjX47oTDi4zm6
SQBxl+vVCMcMJWytWmHxyHjgC/pP6WTvMUQ3FStZn0pAKBDQgN0GnLW7PJHsSn67
Y9ejdRiwt2UoMmc7JZQ7JpcOFQ8fDXH7OQcsU9YpJnMBe+o9j1xdXpflDVCcA0wU
cWSFkkLN1KuhXnkqID6iKFm9pBp/2+oj+l7ka73t5sAvX1wQV6Xfm7p8zR2g6p3W
FBjctpezDVTnq3Z7taoGeStW7fBAZqxjGvMqPkk0moCussBGYZnoPlE44T05aA50
Nu59qrYxZghtA0F5JuvFMt0b0o5pqgrV0BcmFJBWp2mTDRFh0Doqs904huhs7IYz
tiqtk5KwDu6gJhFmmqarNx9tpzCaIYNAREqf0lrL0hVEKS3oX7aTTtBcAGJ0vFkj
xomFc4WTRPfWJqr6B02C7yV+08SdEeDMQteSfWgdxW6uKKPyICHYmiodKzZ0+XoI
cSIlpW4SVbAjsEJE5e7Fh/m2Q7KTvL67/+BC4EWmTVDnwYntWLlfL1Ngjbe9sA0C
v+6Hzpn7AxayLqdwM+Ps5PQGk6Mvp2oeFMNa06nW1CbFj8BrolDihSC7lmNLJRZ8
uNQ0G5kdgqVcsmbVVyNygLn5W6JQ3uP3Qpw+bPyNjDFT1cxo0f6/j+xZo86jYB2j
M/UwmuPqM6K+wmBz5FeVYuykCYxPucMxeYbC3RUuevjPxC+GzIb+XoO6i97E/iRp
pQfJaXeq6kAX+lXN09OninNHAhSs5+Ll7a3cPewsE/XwBZQHZWRa0kFo5QcRJrWZ
h4PylyoVI9ICLmWP0objRopmlJ88jD8ITC8/oTUO6vG1XoOJXxESRZJG9m/PwooX
Q4AN4Azym22hQZjflSPBwsNncL/spgWvx4a3s30z8rI3TuUvwzZwBkk+ZXvrBREd
4W5yNLJrx+mArnbSzQbRDwQGsyJE4Iz4/WU58WUxm9d7H+gnjZWXhiStNOVr7QsI
CTNTphWCDyA/VFXtq0DR2zF6DeGVM+S/6EMT7IE+1ZsWUXkG6RMx5phvmtJiSnES
mOXlKPhmFgSbApRwHBRooa03mA14rRfmWqzCZQFDdX953YvUZnMQ/Ur92Y4Ocehv
2IRXInOMnyssglW4s5EzIO9oAM//BjkXetnBFafGoyVFVV7jVQ0zy3Zlre5fCMFj
MhypkMzDu5h//6ZuCP1vHh+I9ehm8Hgdd6h0Hu6xWiaHosrrAEE2fLMd/78U8EkV
DX/xAz7jy70TvCC+/stYArOwxlI8E6RZ1K2j1M0k+QwmiZnA+ZvPQfWTn34XhCA8
c1DdgbuwNIIDODeXm5tBQ3og08NQq5+88fvcksquefvNsu9P7CpiEOzcpozjssbE
/hT1u2KV0ycSbbkuNTC42Wb4AKm/kaX92ZXdjaMZLpjs8ebxiv/ixZ/pKJPzh7Jv
T8WnL/WxJbd3FdG0+3E4EFtfHDaCUer0Zoe2+csNfGiqObHgKHkcx0MTiMm5Jap0
GywKJnvdomie62gcOAWCxPR3PsNdR8deJKUP9cuELYmvTZEd6/vRNog31dGcpIJf
PTQkpnyboLicofWEBaxQu7qijp53B38b9PsiL2gBWEU2MuDMXHuyOc0AaqftxbKJ
ToePncUfrMk5GBO8DkwpObGTkJIi8xyUShx3E5Zfb2yska3RGyceoOezxSY/smcT
1hbnY3U/Z3FQx9TfW6liGIDJIWswPrcwyVLB0P6LOxDwW/gdzXU6yV6n9i4IHgAb
67dzjFJ7Dlsz3snVARe/xosYjwCvUU2CWkKcZyidzceVJYJjUyAQlWDH9eaGA4Jg
ggvef/BBfrTYCIoppCWgZqHbqzXY8w6TWMlY/RI8NkBQMrebJD5FMJiLvn1REbF9
EKuSZTRAVDurXqb0y/J16WUiMDvi6f9ZcRJ0Z1A5qoDMCWgzZZTch6GCXXghYi8h
7QBBaCMHQLi2pSTfoE+ADuxB2N6mx9ZcT3vnqpC6v2hVEXChonQ720uKvr+iJE7G
2HEI7xiLGs56tvESDL5C/bLVgKb3+2FKev0wWxIJpcQA3n3XtLaMQhV//fLLIyiU
3Sg6LB5hxlClCc22uK27d2OruhC7vdfmhf5DiraLmg2sFlnOzTF+T0Ebaigs9Umw
Obon/oxBMas1poQasvyD67pKAjb6UYAabh65s6szy5w0KjoKI8hNO3hgq7NMKaqZ
L9OoHdzsOAzPhsVqibyJKOVQxPexqxD3gpQCQGoKgwdDOdnij8al3FdwsSsh63p+
wCkL6PK6otMY6l6lMWR2vzeFyL+QHsso6c9S0Vs05hh/at1h60h9u4Wd0W6CrxDc
7dDBCxtFVtdP5NC8a5KXzwoik6oEchMGt3dYekWIOmF3KEhjf45AKvRipRVOaBhm
L9xz7hOzEItgqjOBBt2gpcPUnALBP4psoGSozchV72VX+zrYM4OOxBcdvKRrPo+R
5Z4zHx4AwCEkx2Yp2DJWBeFa08HOUYBFTJs7pESDogxBbC7OGhZst99hPKKi9I6t
KBEXcavvj1unvjtjX1ETTSb9JeKaCexTGCwZPoBC26WnVg25dwQdTxxBJWGiHVH+
I+iiYI0/vwMYZJPUGyJq61j3MLrC3fpMS22Dq2v34+XRSlE0eTYYA7VGwKQ1RI4a
kuepsMy4amKfG2qTfUBuuo0dPJZHU4YC+x0I7rcor6h3tmB9oJBO/bog1qhCGMwZ
8SToWmoBUM8Qf2vaXYgPxN6YL4pFRxb8SdaLrgBdRAV2R72d7vwOwvoyQDmr/LRY
73izRWB5myvOd2aeCtrhdPrrIwmono238fLdtXQngml7yiM0hHwAE/libTsVvY3H
xsOrSzbpG2vynTjFz5nZsDfM6wmyxP7TLJR0ZjZo0yf4mo86aLqV7CWJNGDfqOGe
8/htygMW49Oim+Shf1B002reb0I2yoX0vrlWnd/sUL88pr1NcXWIkV2F6bGgoXUJ
do1Y80E41R4DqX5p8ocqldWWcRHf9s1eXPO4E4BhHCQiCvINoHFfdDnV0t0T9Z1f
ne5vm/GoZdDbMwpSVRTFrVeq8C0K13XNFP5Qvo9aDdDkw9ELNSjECt/Xrj4+0fo3
QszFRuOjHlEvhu3NYt3LgZ7VZ6MhbfpFG9UNiw++izsN3NPdeGOoZUAeUUj3F++x
0wZ4vDlwfC7vbj/1lkfvEN2YMctWz2w1nBi8Vej6h7hY3EFNqU9hGNwkV4gt9Cm7
weXVwe/uW+ol6KXrDDdzEa7/TO+HNkmy2F8/lJzvAZJPei1h7IILuWhXfgr/aLwA
ky2hPqIHWpUaFU0tJciZx5MNSFX0MG5EuX6giw1ROXh4anvJ2fwZ/xuxKhkg9Vai
CMRZH1JJKfxXhBUlJu7roi+W1juUEolF8HxPSz8q/pi/mZw7NHqEnvKCIXoQ5tES
CNPZefdVtO/2WnqCXl4aVPiga77FQoTg+yJbQDdGWfOqD0xw7DL34RM5NA+P2pTV
Iugj53Pn97Q1Y0ugag2SlVl4Lq2erK7UIhPBoTeULaExxUmzv7+1c5XIjC05qpm0
aWiV7D4VczyZm6QY8dbeW4/V8lRY6dGi3ICLv2rvZ4s6n//fYDBKYeNaM0+yCfsD
3lrxhwaTlsJgGjRmd+kv10FEskv/0fxSPju2PZ4rxGCcwYatHUZnVTuDH1Po1G/B
F+TaHYi0lsLvf/7tE+bJZwswOnCylQvKmyOcwuytXkgOMuNHMhfHXiCtjfCVsvZ2
RPtDLdECnfuiY5stEKHRGRsnijhzdGejpNYawmdBKrX7tvYmUYgrvl/T/MfhQLrr
JKs5QXNNV6BUtneOKTA8lP1s9jhEupkQ+EVrOoAOiJG00UcNaqC0N93OSezb0T/Y
8RSPqwxShor4JQRgO9tbeS1ugTdNSE2KR2MeGur6DNGvDS3Rdqz6nQSCDU9pyEHd
vRM3EE1jnpzgoqMEEpfsxeRAtGt/EHpS+T9gNlQWO9b+9vldKKKaeMbogaei2yOd
tg+aTa0hz/k3vmyG7w2tw/Ii72/N2jUyNvR+eP1KNynU0/kjChQXIygZGMylPnvy
a4b0mhE2LEqtSvumhnbRPg1dH9DO/y4ud2hETppVsx2Q35oUAKgSi+9rUNJ58sVJ
4QQ+LdEebS8uCi2/zbsuj/oEPsszfMh/dva5nF1cVGYCVFdlG/uKb/slVKgmtrNv
AmVy/FK26GJtSYnduJ1PhFoB5A2PdN1bS9E0cj0adSe6NeubGN5m0fLiK4vidGMw
7f6uv4wCCjZ7j/9bfYV1E/+1YMVdM8CnU2dCctDciuZsDH48kkEB/MscY9WBVqj+
4PqoJILcGiLkLWVXiOWjfG5GTPLKsPj9hyca2U/MW18NqHfRx79fxgMnFOoxF+yO
Eei1/QhSOhdZuXZOTLFWm9rgia6mZ8fSBvqiGhWz9kBCRG1/y6X8ecUOU6AeJpr7
tVxKIVQvdoFT3X8TjBqyQsbzIxYyjf+v4pj13HLVfaRPduY6+lDfh8E80ykmvUrR
8UtUMuA1W35tN8YuGEsXBiePWKtgeqsyiXeeu4/h4+6bqOT+4Na8eGa6PqXoOHoN
CzcCf5yC8w3v/f+ROEayZ9K7BnHoNFmR4RwnAmfSSuacsjyTE7l1liI3S0Xh/u6k
wAei48XTr4Nf2uV0Pb/v7RlcPX8S4CbPkj2Np+lp/x/EZLzRyjQ5yNeX0kU/sxhs
GgRrepzjJPIWQw8y2ZlHf2liWVxc2Ab6MpyVYyycoAs+D6BNjQ3A/7PjcI3PuVU3
7Wde09kCaArLYdieWBiZtKoSJeJLMzvUay0A/BeJB1DRevbWubl5jx4N4O75BH7a
UyOp2f9k7qLAvu/Giseix7x2sF9UEnS/PlR7QDwWE0wLecLwR+6Vq9Joz4GNVsYk
xWSwnnPxto7a9NoN7A7KxopmpBCMp+/xpdQFnmiK8TkmTjoRhRApdEEXjrvK6AQm
ERu2Fyj2/ik+BTMLlAFEOgObs3DBT6STdns30xexuOJLTq42D1ryxkNl8/VNuut/
giWwPo59fj3SZVWNyvr8WD20EbZshWoKlHJt4hFqrIJ14HMt0zVsuMTA/XnWJ/Ty
o+SkKRn+eHsSTL3bwLaGXXKmvae92HWyeCHhMss2/D9TwKZVgXwbLgwWEs+O66DL
x4zgQgSrUEVkbn+vdd2GlATX1l+fsknqSlGrISgq4jfAlfPLDouJal68HLX4pKgo
VC1Egrdsw41jTHDibeMUWtp5YpYH+ux2PllpVFFADMth4gHjbzi5XAgq8OsbT+1W
bRRoFVp4JHL3qM76A56w7JzTDsY3J5XPbQJjBGrJkEA2u8LivgBr0yIJqTAFqal1
aHswURuhitCuGbivHW9p9MV1YEFr01z6yaS66cqr67qJKnXU1XWUSvjWchV0bMfI
8Sy76MBJJqTUNPt7fh9jR7l/0X9DMXxhAZYHuF160ea5xahOYZAUIEBypukMdfOS
tK0kepF3ApKtFTcDC7udg2qHKakU1k3Nc82ikT0peSWDiyqFKzRa+e6F/tFlE9jc
0HEIckOoRpWrSGsfoCDJZhFigDkEugs7RPuW/TKsSCSA6iSGY6YFp1hPOX85vs4R
9Ps/wG8gvhQbmFuHI0ywwX1EUTKdGuAYepcHxQ0uXxvbZ9E/4f7qpEjohaTkNdlZ
W9+HUQUxsOPkhRLWHBP5CDcW+TlehWb/BieqmJswNQ46Hen2Ap6UqYFMcJs7Lb65
ySn5M7tV8j6nFKCKFq+KgzGiGsTPh3WfwnBSBQ7RTpLffuvdiqb4OMuubgiUmY1Q
YdMwdd6wQHP3NXxKmTY4jTnOGIzapVmlV0+3eDFTfiZirbbVUlHjzod9kcgfdHBA
Igwlp5OtPFzGQv+kjzxRHqG5uXtE8GomX6iQAXRMQs0/gEqvF+7DPTTXTzPiOooe
znPHd2ttQpxsB2uBA/lBsZT/0saGA18+Aw5j1FGIvr3a9rx0DB2aHq7ry12wch8N
yFqPCK/Ux+9x4zKR7SEurJm4NVOcHNIPLrA6tnuQkxnZ4Wt/siGYDNRFlkJQc9jv
9dR4t/W/lQ2bQYas27hyYqEoSnt6av+sKwkk04aY+zX/H9zqbZmON5mzWjhxWVEV
Cok8/APyf+nfQzE7hzRrrdl/PmGGFUXF6jv+eRolT9GhuHm9Cr3S9v9wUsko3G35
swmr+GjIQBwCAlOBWi0EguUxcjbUA5Wms8ABPLDj4vLy3W3pwKOsdbGqm2YeG+bg
8MzWuy6ZxctiuIxbSV/3x06dQ1VWhDaxu0Nq0x6z+aqCvCH+30gkmGdC1d+nN+Up
nm704bTUdkYdlXk+P+spL4B6qVG3IHUkLY9thdDNc+nG7ABo4T9hFdq6bp1rv1bu
TK8BHRpx1cllGCOwo0WG2K1K1C6wBEGxNa2R2k1Fz9NcGO4TpMjHNWUezpljVnot
Qaee4HL5E0zAOW4PtU5xvIMs6JuiTxQ5G7OddiluNfl2GsavaCbhMC//NVmlRAak
oh14TCPYu0n65OQagpfR0O+0+asPETdGpisUsY4gQizb0WV4JoJVMFumXh0VxNVU
Sk1XSx9/1s1uX4IIJfTFbywH66wym3XoHiofXcymQE1ZiZNbl8axRhy6CrBdjw4B
f2AEqP5PDEtovVrzW3sk5FA+ryW/JO8wHtD8/WFk/vVVaFMBHkrBfaSebZe4EfL2
y+XmUzyNtauk4YAEogAH4/lnzvBAOJ2GaD3IPWjpopsHqnMcKBkHqGiIMi+6lrac
h7nJ0x5dzrsavh6tHYfx8ESbQrp07QUNaFLhsXf5c+EfLvOAaCnwtZHGIAb5UBzi
XdWAzm3bNW1vgXIWZbZ9QfVaIUE10MbBhBgmnh7f7zgJ+mAqIqiaWHBdYbTdErXW
M3+mJQYyb/BWCFJgCsJRfVH7IuVxPZAge8J84KlRMCKE76dVWVajAFpeLDowITha
1FiKeQGobwL+vmdXVbW1v0b1wL1HH9yg2PDSb3Hpf35e97XqGc5TcTDALmfUyKPd
sf6tTZy+/mO+v/ubQII4XLyARexLn0XuTLM3mg5NaKcvqvhW8eJguhpw/HqRwmk5
k2i8Pp3arrtIhgZ9BHBZ79H67Zl/Ym8xYuJmLhU6pEXkpa10YQWDR8uBiAD2tqMV
0sZGHHPSqGNfS4URTTR9TlOC2zJlRntLIVaYkkE93v0DBvZSegu//fYsEu2VMyZs
8K8rVyXbHMv4IXamMtpWK/lUVq0a6GoYTTOxr0hyA6Xnt6XdFRXDU60eH1AWoZss
/jA09Uv2hvr0Krda9bXWFV1niGu7xvU/0PE3ZTZyMpZyUC3sTAK/RFfEohLnBxqB
d1u0U4IPJ/lKZUuMu/md5AWWqTu0sTbQJ5+sEoGcxLpOkax9U9dyu3kjhMMQBp/n
OhaRK8VbW43KNdHWyAxTnIbawsgsfD3Ll9wIgSTBgVY++n+j/DAZ7V7AdQF2mEhM
/DDsubPPgHaLQN4Th+fM/0wsABBl231Z8RUMmCYV05VVtx+KpZD0KcOF300c4Kaa
pEP9szJwHJYR/do3oLaBka0mH5BQS6wW7TfnLwWAqzVrh5cGWaeIWVqCf3U2kk67
xwnN/jqGFWEIhBSBjlbP9CwGy3b9XHOoLxUfyEeHqE6SshMX9+/zIzX7EZxHgIG7
867Owv1COHMi2qTo7qg9qhfrgFO5U4vTLPECTEbvjWtTczjsMRLhJ4spl4+Bg1pX
3+HZqrqink6+MggexPucV+IGvYVmM5S1vdo43peklTUI8mOt8pgfHKOe1M+TknDf
LHXnT2gDN/Mtp0sTQbewanG/xnCNGiXiOpG+T+b3aCcdT0tSyEWItRh9thcfu+2e
QsqJd5igGddpDGLoOwJwITCA2+Iu7pjg3WMMXe4WafK2lF8kcRjvBChGANbyR4aY
S5Kqvt+7sUl7QV+tgfQFhQ1LqnrFKsXGEgsKeqQs5ZilqU1xbxn8xtsPSD0q1BqA
GIpjugSZId4iDl39JIrLEnvaViSaK4uDETkLxzykO2CpWpD46Hw4MaTsnaS7kftr
73nDmTZYJb597Rf0zoTGtw2qGh1YFCEEkaSa1ujU8XRLHWW49Fz0kf4JdyXDzSeJ
JV5jpU+YXiyUQcT71takbAy6y09HISEwBufmonnZaYF1my2ypUg2gZiovr07Dqyx
zT3Wq+6vljfRg9T71FzhnK6E8iedcxuQxbHnWPrUPBW595Dtfud/ymTMikhL+/gz
KeS8eiftkO+EqsI1lYAv6MovzSR/9EHDs1sx9wFIh1NQq8Loda4vU4aSgL8cG2hc
mr0/OtmOhGYwc0SgltBQRbMXYAa376vTKC8uoE6chJq2qWfeftNCo/EEYOvKshN2
Rh/+IPxSnoRCkoiwj93jJBp4Z5HOHo9ECKUystKh7e/Jk8zne/tqk0INz1OsXyKf
VTaPehN/sNSjEFskDBC0WhEYJHMYgvznYDlsRs2+7WTJ1YPp6R4Oyq6W0QDngpLj
9kiL1BQXzVenCOgsgIrWZuBUwAjjoxCXoYxpEMzDebe4CcpmzeRoHTaAGs5lne9s
MxxVcjHJ5ZX/6Pwt2NQpSUWH7IsZgXDG5vzLNrGLm7AXm8sYpMMRQHDdQqINxJ3r
Owz9Voh+i3jsqQC6LHWLYIJPU3SO3lnSd0ShyZ5kcEEpQJC7SXf2503o2BJ4CorI
N4mL64VbT3tbgKeiUXcbFxi/RJ7cFYswRT+GZalQPFj/uOqPq6JP+EjvMZDdfLGX
IwbjTrEMhF5zhC6VVDEctcNmh2hYNhIIaCQ47EDo0oOCrtYaqf6ZIORynuXZFmti
1ef3u73aDP/LREYWCMxho+i5p895N7M1lIhGf9+m5VTCRNY2IpFiMv5Td+a3gPoJ
aoPrQLe+lTF+UxBpGa0Nu/endQJKCEu/3UDKhl8pAcAaNkkihl1rNLyS15g1SxU2
4kfH8PufWNs0oc8W49PPxlfGT9wNTgXPHjd0T+TuX6WwlDN3ZSGHEfAl9gX1E0Gf
VelJhdaP3TvU13kajKvdPjJbO1aDftrBwF3tfRlkJdySX86HGsb8HFWReILuams6
q90e7Pg91/zAO/g1Gbhy31NWsd2h0GJfEsr1xOitC8TkW6Nk1xt/BTQ4iLYyxMH4
Z1dmbreKHT0+nIsqzrjTLxmpyvEuMmOmflPCKOekYhmaTm9E8sUc7fIZP6VltF8S
Prp5FZHaM7x2FN+/7I2v/Zt0rjBfoXXlJ4El2aqF4tirZzN9KMbuKRVzycBrMq13
yQdFffBj3efIaDwXIQ5KI/UXo5dwZEkwQiJ4FenN4c31NYzvz0M8y6e3HKVBYgJG
0YkiPVsZOYdOr0e4D69xFUYkNqXF6os+3jotKfAESQBmcA69N3NOJm/gpfvLQ1nt
uLaaGmzrKJPOW98PnYbMm+uoTwflwV8DyoDjFUU983KeVctVk/8vvDCbzx9kriZT
AhbsY8dqKukJ391pnwHYnOfjV2AQF0FgkIXARZjJmI+WlcP3gyJCrwJSJZR4FFYv
cDQJVS0PLSSiLAsxBl4rxhV1DCIgHuNaI0mZmuXvsIfL/3qjyUzY/OH9sIseUlk6
+pV1Sj/Fz5rRrOKlRUbXC7rg4zO4U/QONKYEh1gX5y5fstXeb+pQVQQsYE8/w2fo
uzUseB12MOIjDXp/6l7MXS0cIFZPCOjsIbAws0/LOJmlPLspIwtSKc/+504l2tVA
pI12gFRqbh3SRtdqvtLNj+DOEUe8o10agriiTWAtJ91zckVUNsMiQN7/4NEAokrq
8bZWlZAtUbYttozUkY2biUWXoQyXu8SirniWLVJKrIKzJdBTK/nkcd+2TOL4A/LP
sANJ/c+EMK2DhwZB29svhgW8Ao/qHNYLuljampdEk8vF2jmc03Q6HvSZbOlAU9ir
QGgico7MDXJ9AR7j0S9iaHfUvwX75nxFDKNIdqAcAvgZz8n34IP868zllTbKbaOj
oL1Cu+rhlq6yVhFt9KT44zo9KLuXdTr34v08rOcMuTx4I/RYSOSu9KqXoHijlPgm
zZ+THWFfpv230x4SnhoLUeoKiMcZy1c1/ZQZJIB7rjcYydOOqTlZsb20wrGg7j8E
oxPqFU51bVv+D7gj3y71U/uqvqSJbEutSFFwsPSJD8u+awZZoa3QU8I1WsnjH3ZK
+AKLic6C0cHxhsvNhutasvz8GWkwUBuKGPlQiXHwYARHoc3tFFADnYwuLs+YEdeS
9RG1Xj0P6f2k8ZUxNWm83iCAqAqobGAsZ1AXf9j42JVwod0XBME5jiR2ca0BQb2R
FVOaSlPxUJTcVL8qm8jc8A0ZG9yGlMT+Fqfeu/5C9vn+UyxYVvxNAsdRN/l798Bu
U2Y9ylkfQQliSUwXKdpUb/9EccJE26hlVHH2uAAo1MBj+FSLqR32imxHNdc29qhi
DlOzjL2Bq3Bdqt9Sipv7CBFNu6QCLm/Z3jl5fRKVh/LuoL+VxKu4Knyb8LJq2m9R
QBhAXHy/8G0FtnV4rewPVUG1Y4FuL5e8akU/OGkR9Gd7KK2kgjG5XM2ljfa0JDR+
jyEizB6NAMelpVPyE3ZN2xyiKpDXRNTUMiHckebuTWKz9t8NU2pwA+xpMFK4yUPo
yOieumkAeuLDUGaX0MqnLFVUJYLqd2LR0HdYKgpWpp1K8N9g7A2l+uGnA82jZroU
xpNPJwhAAz5NnrtG42E+T9odXlBuQwJGtTYF8bctmTlTdPZuH7472r95KNZ5lzcv
zXzWjmgxC8JO5maXX6utnwsKpqZ3yjYjua9++I78pMkl6vFgw05bFgncwYnv/YMD
81GYxmGlmVD1/J/avBAxxvt5V+g/lchmCqJvBMNvjGaHgCBSV0SbB/LmanlGqDYk
zn5pSlWdv5j214Y3+iSGPBVjopjiQ8+JQ5UnFGrL0GMlYmYXgWnc5Vd//tsunQIi
BIk+VNUdcTPAU9oAnQlr9cOjka9Zo+m9rJpYBle4dhKI0l0HYRIw8DiH5LuroFmS
+Li6ekPdH2JfNGlPeCjou8mul+2Jc2wQVYF8oUPYezfcynkoUCzt+GxG5lSCStsY
v+Fgt3daVOMGi0E4NvafRHDjr+Mrw8PeTQVZwaN1jNnTetwYPribEDHORFnjIcsC
mYL0jCN3KZZ4Hk8835KoYPOc4MsPsTMhPiQeHJE3ApO4pdrhjagN53I/0EvIYHWY
HXRchv+BJMiiwTPOKNzEsBbCRkVDrIs5V9Ry2zshFO0/T8G51o8WAN06uyXpfV5j
MGTXQ2Q5zgTEfSCLRFeW9i+OM/dQJmkEPWaCOu4b9cSXf6cGfysfzDp3uh5RDyD4
OKs/lJwng1DAqrZjkr1kILUE034tCJiZArCnrkQXcmLls7sFAmFfOmQZJqZj8cuA
KnIBj6qC7tK+hVM98dIiHzBvzeR/0nl0P6qns2mv2vF909KpkCa4zVPKokQDqj16
rE7P4J1tui3ZzUW3NuUxOqIVGlL//e3rF4K9/rnIZ3R5oplZ47zkKF44R4QY9YfV
dRmkXRx/9rA/7r+HmLTN7EQwGxfv3mGoFlO8l48kJ5pzitEQ3O2cGeJJE5dvFIa3
mi3M/d4wibuLQln7/upUB9kvwbMGnpQ1ku2AOZKPJJkLtlXpCAwNw0pYZjGk52g7
RQTrT92zWjqypWSRCu3LVgh4d/fo5fDOP/6MRkzfpUNxzaZO5OtTFt8y38UHsggn
ZjvL3EQyLRr5MeRf0SnnAhO0zkhIMUroYULSL0/Uv8sBzE40E1cAMwYki198mLyg
j2+GbQ3PSYeJF7hZDWanFBbH3TaKPoMX0XKRkUEfDsvhFnUXjnlsUr1QCl8q1xVj
rv8zzUKmTyx2+QZF973SHTljOmncUEuftSBVEsG1wNl5PeThD8nEEstugHAW+2aP
bncrz0++TCFNa6FpgglI20lOepdeBFtNR6hgOzFn5TpdmG5nS+zWFeofOhraGW8K
PZoKuacEnhhFhdmyuYcXImknFRcxoSAcs7ytbv+MLrvnViHrBCzly2XEzrQRqZC5
6RYkfXs7/+SZBemGOuAAdanHwiKuvROEILsNKUy7EdBOnhOCAsSxGkWC279iiXXR
MICH+jFkktJjWehkafJ+5a9nfrqgXTbSCo2lyogXBjjz3WGR7obku3kpZopWL9Iv
LjtsJUAa3f9JFLkEx/k+VYFRbpLeX4sFMeiFAXgrpkzLLtsA9DEPCMUDCx9jGgjL
9F69Mp2iFBbZKdmre1lteFSVtk/nsS9HSSTbmVLLzMeARBpA8B7VLlobTw/wz2rX
mgueo5Vd68GtkvoKYnAA7RMaHxfer8L/HsRIipUiw4Jf5DjutmnQER0Ka33is6dV
qqaM/kUQ04ASKi+S6PSCPBrZZFcQ/hh3KjFpetxd4w8cckPBKBJRO6ZAcU4ebBCD
IL50UBnohjrNYvypb+HXA4ESaY+HAMJq5FO3GAJB3kwt9z7Cmjm9wrTVye7/CkLi
iZZyW477fDKzubHuZms9AJpJ385vuYIXGFWR1e/9hQtace7Y29+f9q3e3CmHr8Ew
hQ+QFnNlljUDnnOokOA2n85aDE6FBCRtoVISikv+B4XTAtXi1S0aCuuO4Z2EOIYn
Oc6ugvIInN/J198dV04cPmRMMghfDH28wwWct//S5tDvWKEfW7WoIsBfmhtvQPp/
3I+FzT+9UMRR/HqQRS4s+SiRa2/fo1sQpR+yE5zHbKjNMQC6dpV0q3Ggoizt1lm/
lfoTMs88C9BUJKTbrKGRvDW7+D1iC3QYrtkIUFtrPh6fGnbT4e/LQzyzY20szO+U
nvq6mTmcaV+Hx1A+LxmBkSA39Rg0rUF157NgIQPSY4Lf9Zg+ASkenU+2q1t7nDI3
e6NQF5ShpX2WOqRKk6OYVC6VBHxy+qNsgNJCSQghvJs7AEWbinMVVqgBNviVIz0M
8wnF2b1jzdBqs91/G/fm+IQyka/hGocw4wFc0p4MpelfV4oId+ltToeeF7Z7+vDO
m/7wa0Tuz2O2QJd/8/IvUpGgsZceBEtZJISVKGRs2fTI/T1qLS0rl2NNJVFi8MRv
c2S6yqLz5Z6mUPqEGIT7CAZbPsGXegd7yScbutok5QpcmBw1f8MFOs2PEr9e7+oX
TisrZPC6bUA42J+4b4kZqhDRbjEp1SCqgN0JSZv0SstOlubjhLvXy0rp2QoqVudh
U3u9hSiaBr0UlXO0RbiBnYlZ5fx+zabzW7xOJ2wsJsa4GJOPOPXCv6js3YdvS3kP
4ndRedAx2hOzQExLSUYIHQ6VwmtMM/vJgiGXepcEfNl19VpUHBtKaAvGO26PRhBb
9eGnY+FG63h6gP4FYVPPynFKf5eAai46WJZ6F/673kZH/z6YhWeEVgZI5neZB9lF
pTVgypWGA5cFcqBOh4tPP5jyr5Guv+qKl9wr5s8yZqiPjDfRD3Yq4rF95sK080/r
TKjR0jdRJBrAKHdr/FvwMzAVDrkgxVZYqXgE6Sc2jpO6BpLULWVqLGByQZzljoF+
QhammHkT04t7Fn88sJf7A6d42JEDVhtbrdjPNEcuzEJlG+paTZgNkdhYOXWvoXQd
W1j5AofgnQGaRmszKE4utE6QWnQrbf0T5n93oTUVErykLtOs81cf0+Y8O3o4f0Hr
kC4fx4S4cprSvfUPXQXWyCxz5YG16eUAU/SSi3V11SCFmv5zHgQzJ/gEPYJxXVML
hMM8vSeExQxtTAmH7Cp5GFAg6CyPPvfNA6/6llCVOE36skgDJ0g0DKMPSqUenXLn
1+qD6GvnSCDXO3ipXAEBAOAQOOfwAN0ldsobON5JeWl1BtA/6tuUwaBz+ApB9tEu
fMmhrxmOfRnaar8U6z6+guNSBpU6I0hWsm/e0uPdvnySDMiu+2nHa/Fj9kepCn+/
Gd0Hn/ob5A+I8Ucz4hlEwOKZPpU1R05S6mlJ6mdOdRX7KPXqCoAhlgL6hiJYDiLz
G7ZEFhjoUVlVn6JTK6RU30k/zR6EZV2mxYItbgmgcx7/wSw5TQp/Bimwsy8SysrS
XIiV4uh8HowSZkjzfk9/NRs3fj5xlYoWeiqL8FBH0CkpnDwVB9VHYZKbquYex97f
XhkZJKKUqpnI6VRL99v+NrLYTdz8QdBw///ooQlX7futpHKlsguAkvAk+rKoUos6
ZiYIryX970rPa1h6LrfXsExpAFDwxyVZySuUb3Rtgnk2HnoUVK5sVRrbQA/mVxPd
djWxNIyjhNUuQNM+UsnyOZ9RfQnkat0bG5cD2HmJWRWjDSlIj4+SiMkjWeZdR5Yc
cSXpXz62R8hETsEdN7iPYBqKUT0fXtcTC6XiyIlryca2sVc0jxGEHR+/1eYzyefB
4fEURMiRIdd+8M8/QnlVJXGVrSckL3pFayXm6MEJlE1g4FOMYiVzpylgaR/Vw1CN
uS6OYNA5EWflfw72IfgxW5KPkk7SgDdol0pcqC26Jwl6hdG7bOuWYDj2Co0p+uH3
0Jyd4I34P30CZsvXaGpJv9rQD9PJ+8XJ61PGIR0Fca7DnNczH0DGz3chMTa6OBkv
nOSIsAPA3gc4pYUdjXMVBN+DMYBV238t5KOOfE/fYfksekAh+Dq6xQnv6QKto8Lu
RVTTb3E3M4pff1vqGXyPChELjMokiD2/yPVqtjWYTnLZLAZwYQnM+TjxvmzmCQCY
DgxrYI5KNlJixSZPCGIPvGGSrp2/RNskVXp+gZY8Jp/B3fuNeB6qPdLZj1JB6wMo
TynTfXzwQycj4VTUPRfvQfKjvRVlL7LBsYvhtCEs35fvaoYn3nZOQKijqkjW/eq3
EqNN3lTSVpbUlrK+bIErwwRxj0UozPxFYCVqvYHtWdjOu+dsEcpKxvUd0GmJcJJf
9ZyJvk5KqP8wqQZD3p48bvhryLLexYsk3ABpS0r7RfdwwxS09bg9FEMMW6Gr6IpU
qOjh8/tfn+fP4bBprydPcc6CIurUuPZM7Oy61RaKdZDpQsq3gykkE2RRen+meaij
waUo26LVFoSSYXMyk5hrWDEYGXL6Pb+8QtdUZc2x+JO8+utAm7sDqu+nsEuY1uK1
FL5pIdItfjricsKsVkup3jA4mmOqZm6Jgksxbemncurz7LuMnPUUWp9MGc2kSF29
7l5mDSeOSuZBw6l5bCtwqKzQziIaNg5env5yDazQiAQAKuYc3ooYiYhnbvL+mjQm
o+UkJU1l1rJgj8OqlIx4pMrEqxHBB1TLWdiWKTNJGXWGHuHpu4kP5PT+wE22QkLa
2sE+5v1fWK0LymLQR5wDlH0LUe7kc4AVEoboCzhG8Zr45bAF3CE5hEAjQ0eZBQL+
y0A9cB2K66FI50RFQTyv9y69J8pLKOrIBoLO8dHSq2+fNhOfsuME/J9lhOPVAgUm
PD83rrHgG7cRs0rMmvSH3JCHDftLejyi7ttK1/l8+xwBwBov/aebJJZZSYtoQNai
p/CQ0xHgOWtCzw1udxUtViciluRl9F+HEZ10+SCQyjt8VKv+WW3PcyqoQQYqdF8V
8mioWUcnHDXcGlN+qzfwm62WVEH73dPy/K4FtZjK932Xhk3IS+tcFPsIL0ToTIB1
daMSA3rhaYwM0Jp7kX0x8SxCOce8tmaeL+FdsiFk+HPaoavFyerrNw63aUcd3nP7
Jur2iWfZoXScXvgDazJggVSviABGyOJcUKRfF5ZXdofRUNsIVxI6AdU7jj7HyCaL
4k+YHoFjZrOs1pYayMC9mzQfHfP3vGaLO71I8L8VtI8IeUibamcLEyGQYQtYAw0a
bjD2TO4nnXYif5BRa3bqCu+Ldk1+R7Mc7bmNEsF7bwWSV70Ly3rIwDLaYiHH+wLr
QA8egR2Cn5xkFW0oyyAFooC88QtTDzIU6fdlAAElluF6zQOnX528i6d42SXcepYQ
W38FMzUS/0xkeCYk59hhvDvnM/iF/WLKwOAcEF7UkU8Mu6YBUVY2/jW3mBPGFMTE
21tH2GKNnQQfHrwmacjpl+cGkrVnk6hsLuJdb0+2EZgv165K/WwuuQ8y0S/QKlUL
EbtFd1OhzXFVXIsMTDXukhAB8LmSFGHXz/SpPLEWWXwDFltIMr1bn6H4dJAOwWRu
xtC0Lpe6T7HkMN1jVsp8x8PeEc/+SF6OxxTKhYICIgYIiXE59YadA0HrGRLpgb9J
N4bhhJcZuJMOwCdK57JDAvbFOUMnVYY8di9t4aPwue1LsippaX48gnueDTqna66p
Umv2ZGX7SPg2Y3NiJTqtriXWRsc80NMt3IAWqFRUHV1D7Ra5q5axEA0BwklnaMHa
YqrfTPED2ZPkiCnB/l6mqavpD+OmboxFKG7+TGWIFoCJWXafsheIOka5zXSzeDWs
W6+1hFvICdxn1692a+37vurmds06j7FTsw4HLyFxD9/xX2QxYtE/dDonhAuxyTIq
Egu1nf9Y84DjwZ/vufTpvlStmLW1vPqPXqI0d0TbXHZlwSufIjumvz593ELmZO5z
ASONyQAUdGajRw/8K2/ru/qncKtusrbyiXhF2BY3BVXF099IBAIONSrEZ2VcjOjK
m3uwVWSBdF6y8ihdMpDvpRXauE1qxj9uIAQs9KJMqER1T+OxnJ3dn8jt+hQdfyAP
MpsPe8gVJIDzrvRAn3SVufCtRiaJPtNRoGpss54u4dMipDp6Vk/EHA6z1h82pcAF
UB5enb8upqh97TuWQP6c+Qx0lPtOHC+kLwGN2Cv2zaJn3UlA4b7T12y9BIunyjgz
rPQxas5RNVhMFyn4uvs4kK3SMHpU2NhfbKWlUs4o8cvErxesS/6B5k31bIXwWmlK
f0ifKTbQWzmwklUZftJxyEcpXRflfaDQnBABXQHOrRU6tRHUXFYQi2SxVI2JoUKu
tRJw27OV8Nnq3IMkgamTdcnJabY4I5WW+zMKjXrg/6VsZxS3jUgXrosqhH3x05uu
nX7ES4eLi7fueHoTG4cjZFsbcLd4n5I78LKprkJBqy88Nvb44bnFCyZ7F9LeVfM/
LKfw1KlHNNWP8MoHUOnvRIbgoUEeWvxPZIo9hAh6L/6DkDjW61cei1NHeibdUKgM
MABF3JppVUg63HwAcAF31z5YumIhzUe1kfNMOGAaPX/O2GzLgu6QMr0K7XYaC1Bh
S/L0/rSBWrhHGQoA2QY9r9eeaB1o6TV5FZXk9FJU0Ig6LPARM8nr73aZFnEkL/qq
cJ58gxuFBcFMxyUwnUfZulQAeC60GiiVxgk963PlHAnCgqfJ4urtiDUQjrlCV3J3
Q3V1pWVIaEbPWsKGy824IVFJ8fqntQBXRK+Barr0TWUWZbZKwAcvStL6vmuQXTm0
LUYp4Dcp3eKnwQHGb34DipfNeVyTXurkUZXzq7B97EtT9/PHn125PIraqu5IhBIe
MhxkBU37wcdK4L/6PCIC8jP8wmWx1L7BSoP/nc2Pw6fDK+yaGRwlcRtdpNag2n89
lTatJgeCmFcwkS2QdLUi/nwN6tc2oGeHd/7+OGoFaFthP0qnxHCNHLpFI9XbO+Bk
rmeJtPmiQvkvLcNUAvPiEGKI2IqkPqlKcgY1z4fUbtQ7bRNPaXFsPk07Lp6ZtgHY
oFcEMfYwFyBh/wW0MigTzpZbgPaqemV6heDiLxWrTotY8nN0gPRSFKJSqmjWGGOX
FxFR/Ohl7aDr1OwCi597Chm9Hb3A3q2YELW00g+sJTe5mhyouByi/XBULjiQu/Gb
pOnXDJLWYuap9TsVuDuyWtGUv1S2ApccgxgsXSP3iGcgrpB5LAih1BcQeF9bsxeM
yMp3E/bdSsmRb4Cs+4IhpDD7MnWiP+auzIf3MVeeDPqPaPLNroDdAublrxweodlw
/RGI+A2MGk9GIDtSVBfGyl/LMFm37aWk4L9QFqaGtjdvuoAgbehvfmA6+1dFCH6Z
Ys3/A3+Ee4cCFoSpXED6Qsv4hjbGQ9Cy7Q3p/Wt/CRLbv7yX4EVY5lPLzYS4cTle
iAEjBzoZHIlM5AEOHxs+xVWIa4snDSKLgHbo66cdCGJjkWchme9gSfZtbBH+F3wz
SSJiT84aMH9X7fvVtY6ayDw2WhC5S196cc0GxIay2Ekxq5QSjH4yKXb9wjEPuNhI
AnpoYXMdoq5xXpoQUHAQw50TsrJ78KmTXoFEsgkydbQBf6H2fg53fZ9QGJ5R4Xmn
aWlnHpde2JNnBVBKOVLxkQ+sa/rfcAglMt+OxC+h+M4soq+r2/eox0V4EKBCdhbA
413DDzqwBua5AGaqYMR4Iz37b5+VOpm9WjdP4rnH3Y/xHzeXHU4NCQsoVX9BNHPR
hJheoefN6gKAKHenGZVRJYW1WQU+yP4IeKgz2oGLBE1TOo1OhvhA9Z1qLJEfzZUE
7B6HfBfyOFe9Kj5fhgjZSkpY/npI8Ep3PSyBbPpSzBn0tusukfbiCDqV0gXJAcDb
KKr/6h8MQhmr6+IFzWpUxkpypATLhdXeQH+uCRPt7InZ0Kiqxzb99L7n3MAdW2aD
/83WTUApIYQuxSDUz92HT1RLJuj6VLj926lCjov2VuZFSJjU1pxjYbvLecq8UQNo
ebXnINccWHPU9JlEWGVOjU81I92H6nv/ODwpoVdhjgqLebTEFqkxvp31CsNVA+JK
/QwrsrVpaYfCwM0ikhcbUnTpfQrVnmD6zh9Kd/hdaugvPxCS0C8ju5T0w1aLIlU8
z9qLp/zhu1XtWm9W8Bq1Sd64JfvJoyfo0VUfWLuQv0LB9pRKIlfdnrfkCCcGcR6k
FLHZOC99aqfZSMi3I9TSAqnPlbFF/OApvfjfv04AOcYITJuJ5yM4yhHLZ+rVrSS0
HOfFi/AMIlTSogKMT+CTIe+47nFQlNeAfGY5HTR227aAXt3j5PjfjVcaqha9dAXm
o4bBS3E+4ypqCk00t8aAaKUh9BclTeCKeYLdzDRdxqg+JJHNQmNTGKH+eiDbGpbY
g/whrZhAxqJJFHvfnECSSuYlioOZ4Ny17ZIAwUQv42vWg36flolF3ytvb5M/9nMY
EKOhB5bdptLzzS37CSqwGr6cRv9ENiJZLAjnwjo+2BXdP6tZlkbrTnikgaMjWvAT
qPGN/6krOSfvcmbtjUrBYgMBjogjHZD/tpnXLlbOzATTWj+rHbr8rhOCNiGeTaYE
rwQIJM+2dNpqW4rcj/eyWS6D3YSMze6llCDS+usdQEOB5WNs7PcK8FgOkAyRp2a1
p/p2xjM55S0bYxsx1moKhpKAgne6PqaOgINdz7zWZyeiJoWgJk1L5ZosruDDLz62
5IeTv1DurNe3XDMqG0/YxNoTwEWlcGtJhCQ7YKKc8cQb3rYb6QQvd0E78PdyRDuT
X4Yi/UBjgLeiCqE/uuMcW5nhlak0/mcQaaaq1UX/B+VXkbP6pHFEj2Qu29wlyb2E
f0f2Ri2zV/NQ4VuBIT6o4YyYqOSpVAOCNGbCtGzP8wuSqW1KfIuL0kjEwG8Bin8I
lGX0lK/5BuaK+P0uHMIpXannBv7wyJQTsg9SOrlZRWByXZw6x2mrnO4qGAIlmovR
7u7uZFmXid1mLdP12TyTNjAAkyb9qVB2gkwNq0Tn4qlPa42rJV5R/W+NUvzpzqkS
v4ks3mwXPbrOjQ1HB/DxW21aoFhECtpB3ApRA4cN+gTj90AHLWIiC4/K30i+xsZM
4GCswPXFFU3KczFyjIodhrE1jB9tHXM3WZkeDjiUYQWVseEfUAtq6gw3te4CiOm1
Q5mZLflI3g8XGwYhEBDQtismKDC8Wp2X5yAIo2iI9SySwbWiL5Tuk8GmWEj8uu6c
PiU3+xw0Yq7hK9BFTf2UlvVrj1/y0MFTqGkjxkJUqlgbBcca6ePGbFLolvo8ZHJC
josvPkQKMYhinQHASlD9N98jq5bC4EBbg883CupMSUKfpwtuCrENGafsouWxaj4R
D0EZHZCLB1PDXChBrGpbABgXi6AGCR8TZo5DoDNn+W8bV9e4y8aXaDciLKyDxlNP
E3v935njvY6XRrnHCHujPGlx3NkTv+mpBZkFBRpYknFABPh/Z3ks06z1T25SBjUF
HNbrxvBAyzO5xkfHRu0GMA05obpVH4JcbHvpeOsV2yktMUT6xoGJ6UiWC2XMaiCN
Mjn8c7yUz+D3o0a+Pt9GqDTMa+IEm6GbbX5tZUKQCAX0iWGHWQ1pnr8saHHYsdgI
FNRYtfl6XWM55PlNa5BVvES41V3mptDOI6+NUv3+O8DqYRdxyKWud5LigX+VYpEe
rPPTWpr7RK+ftf5i+CscTKV0rmM9a08xzAtsSudOeDZ+V0h/H7M7RA88xWBHJrmP
XO2yhlIRx426BSe87Iji7uWi1QnGfwrT0gmIVaguOk5ChyzV+tVe097Wmjc3Xe+9
03olrzFbqzAOqI4HT1HI6/fSBWrOdkGjGa97En6MbBGuFjAQwaWjnFoVMhPiKNBn
5VALdjOzzt5yisRoe9oXgbEwe4n6UQ7D4td5cJ09QuKPCutACYfVXuaLqu6vYMNT
YZT7ku+rJY4xXyDE2jOJ5hvdaPEO/0Vqlua3+JKLpXJPMZlnhKe9O0zaMhEMoaNm
Z7Jg+6GepssFVk1McecB2O7NUolE0S6wWfo8wTyZqbJ8KeNAJLZllj0nqoztC7Oo
FannU9AotDRNBt87ColrD4Y7HHWCp0i9l9rGpJrNSe2Sx1vFTZSFzGe4g5ES7DER
/gV0XiZuw1AkJ7ck0eOdEJhJvh7th6cGUsOgKYxxtY/JoJzhk3xkJgFus4liJeQ2
KOo5E671tNTMMNV85/kMUNcY6phJe4amIFgj6iHsInz+upi0u4q6ughSy/VB3yzz
jS/VKGj1iy5LquvuOGAA1ibSBghVXwjSkz8xYX9MuiDEyuGort66YQwLxJ8b6sY8
az/QEDT9oF8JXZLLeDkT8UhjmxnW/9pDPGWIcCqSfRjivAt2t+PIS6BkBuCx1uNo
AxmLCUHY6gMjRSktwF2mnnOXtAXKtQ9yI8qgTlYnkWwTq61VVlqeE5SANoQXYNw8
HxPY6Q0/ZGRMSsLtyE7KitFgKGE7F4BeVWkkqmUgEpzlvXYy1nn7UB3UY6VFCwAM
bb/nqD93Ev8k3g3AhneFx+kAA4mxSaaSAE4Mglb8dP4bi5dPX2+oEv9El4Gsh5su
wRGjkC15swiLqPYKEgJFOMA+TgQ4lNeOIzarqujxvGGfON4ngPHIj4awlkIgE3nT
/GTOligtporAS0jAlwUyaXR1I2axbWV+Wz6b6QAKOspgtbVbXORMFMsgLjU2urf6
g4BGcCCN4iejlL+MneE6ffWXldZjrQCpxlG/H9S/cn+nCwYXowznd2HGaq3j6CxZ
S5YEkRzczAhvFiAjo7WXm0gXVHy7RXS0m2IK0NfP8RZEbFH1aC3g0jhC7i94RsDd
1hj2EoPILdC6OrFXpBnWn2fSugMuIbgaetL0FLLNztAJqCyN1SSgMn6DR9y2E0rS
vFDOgxV5QnCr2qHmj24sFQ+RZKf6UW6aWJxzKr6ym0zDyh78aDJjxBB0xKDQzpVf
Wpo0cEDeEQ0UEdrqQVKZP/uGvgHVOFj7VRGk03d1SK0gxjpWlxmfOfNC+SWkc3pG
FwFqxnnu5Z356DIQMffMKy2gLK1zkANVMJMSQJwp51j2GAEy6iSVZfObqdTfy7h2
m+u0zb7qlYm3KwdLLaCqGsPxLrwxQtaG14//SYjZDQAfLsadSjSr5NVygjCzW52m
PzL4IbFQwYPSKMNce4oIacDvD5yqua2B7hK5/D10IPGuyIc/Wv4b0FeKn3+bzcRv
tsLFPnuqLQSpVdON/S1471wTR5up4nA2fzfZzFW4ZoAwqIoZ/P6/THW6T1fC8Z9+
udL2lvOy2hxawjN8iBn3te111i6DuaxeAkSRlfn5P3xLPb0RNRBu/2SUjgucFag8
09oQPu64KpAK2yBis/bqNcIslgEs88FGH4LhbpS5S+ADRJAD+Mp3BcFLe/pYpmxH
MFla5GbTxwi7bzcwSQTJh1ZMYokX1WhBwQgMOtmIWXqIR6MVfSwRfcJ7DeMVCw36
IxNIguYvyQCQSG/dlLT6os62zmfyLibgbjYLFDQVZ/YA3q80Kx5dSvzx2V+i1Lxh
9IE88XB0FugtYdZbrl0UcEaSGZ2GPUS4e/6BilHhW2N5LFDzfzAW7SgSMqd2r8yh
9vTL5q+rNQcGzoZMRFJ5VNZP1sqdPWs+rBTzzEhicwXz2AI31XoXfZLE3669n2wd
g+UFRKBaY7JjoMLBfUAZR2NXUuIl5Asp5rbik27w74EnbRkEL66Nz1MNCawPHXqo
ssO3vcDkllwJYB8NnA3L0k5/O4PrBfuGsmZjpyhj74K7U1YXpA7os9K3Y/+a7YQw
dHn+3j0scuWe0I5aqKXT2ctybPD8ucnfELAIkYjolKDAPx4+qGcYhMNT7iGn6PKy
3RhCZyZ2CEg44MB4pIi8IaCo0VUbKzvhHolG+EZozqTuQckdS8kxjgMNyZXeJ6kL
6eLU5aabV1l2g6d9uzEz/Z9aBUifuVZZTktJXop89tQqcADcdQcwC4uZaOd+qq/p
yMjX5jdcnWDhS90IWI1jYLjR2X/12441lcPtMQzvY6o+T7BODXCU4RTkvczepbK2
gmiZobrYI8bz+Xk9zyymlaPAL/9HYXHtxMJjUWTV1AyKGaBlBvhMClChO8FKIqWK
NILSozEJPTs44ab62RgDT1PmzMGE55NUbWPTh8TLJinLCuBwkjWRw5RCbYz8krSP
iIJcxEhdwsZ+65iJI2M71Dadr9ZMcAG4/1faE/zcMUjZBMGHRS/KLZJ2ThQBt9Ba
xkEj496fTW3QxnHyJtRlocGxLfQVJQgt7NK0h1x9DGUl8e78Bu4Oo0Jwn/37rrOb
IJNWEd+cNhn4RCMPh43Ah0uh2felByvrmmorCnrTFUG0oBbRW/wNo/0rFdLKvSpM
giTcuwYHc7egSDP/SVSv4pQk18aicLHvzYhg1cRynAIF4UAtGmKmPyNqRM+CNe/L
jfxrwNDp0zbhr3HXifGsfEXXYvZbSse1UvJIWHyBKsqt2cf7oXRA8qvYRSTrHoEq
kxupDVLcSPXc5oPRAt1zhRqso3jKHH1GNhSGiZ2bNiTJIuB2UefkrDusIisL2I7h
UreAUTFjJZZi8r91v4Y56JdHo4rra+QTLn5/h+G63EBkkFScUYG6ZsDdyKppnfT1
Mbpu2PFi6eQyph4FCgfuSBgHuScdIL8ocUw3rLuzQZD84ONk+EBofHP1Frhe0TdF
8LSphvdaB7brFLgjDtokJhIS2g2Tqi5G0fw7wuwm8E22AGLQRqaSBSKEFDdT4e3R
S9RwXoya2DXq0ZS2sY671FwVf7pon3DUFuCd8DjBsgXq5zA+LL8JB9xTG61ZhWjh
88bnrI1zSbDFlZJflomx2ODI14A965BtzAe4i7ovGEJ9OKhTacmObB76Y/Auziju
niPIvZ8vWfwv7CKiEepaWnCOir1CPhf9HMZ5AkNYuAs9grU/Uw5HrRHqk/zM9RUF
SR0aJDdy10I38xy/bLTiaZIdlkPAbqAg+P8z6H9dttJnNSdFY007ChmV5Zacd1jm
J2OpKMzEvgxk4972cyGlV96m0EFlpvpn4vk4pElT6sM7EXECVUl/fiFnQu0TALa2
kda2Rc9uZ7usnYqVSe6LGetpXq2K7X1xj7RbD9g0VT8ormYH954efDYv+I0httKR
nLjVCSCZlQlVW6A3K3E65qguqdH4rTYKCCnk6TVHmwTt26N80bqLpijyZisa0QTX
Y6+h4XjTYH2FWXU68PQXFYcnCEPv1Ph6DLUWJ6n0kGaVas8msQIr4XMQk3xmKrEs
d5Z614CVxER7oXR1TkGAejrv0ApcD8Ya8AVHJ2OUQLVKxk54L9VZqI1fDltgoMbs
khjqZOVzCHd0ZpGjB6LWZwiIGHhWLnHb1yLHtw5G4vWPQ0pv9O7SzouItzJFCFAT
/hGB5m/KI6qLfnrp3FIZE+dAByxQtrQND3GyE74DD3N0Nr/HtCJkcds8mQgXoBCG
EqPLNcNDTVQ/m2FEuLNMI31zD146xof/LGUpCeRv6fZ6Nyci5Y4peWPAlSd1BNmh
T249AhqckpbypKvQj5ZuUQqYsaogTXHNpD/7FiR+ejmJHZE2uD/gcINK3olkktMf
jVfRvcF0yQJ5VXGzC0U1WihwScuxw0SOLBc4va4MRWbrEKJ1tA3eGM92rnBzE9tT
iXAOQzIzgNGhdu+JQXzfBn6PEFCN42wCHThvEF5c/yYUiZNUWXleB0K19zXEV95+
QCXlFnHh0C3PkNFKNGOGEdcFLBoU+6t/8Yp4w9ToIU1V74A1leUKS1f1YYrZIdPz
yop6HDrKuEsTFwMJzukUYYFR6hiDVb/X01YLrvEhHZ6hfklJjqbuQr/uHCqLhlox
L0VHx3vdCuvFYAsuFDKHns+D540Is7Bqx57n/Xc7HIYnLJ5jWcX5UciD6b2H4OAw
rPZ5Q+YtAXe72LVq8cH93GWpD3owXzVVHkyYuvxYhmkjMO5wCQLrQZyD8wmE5qbl
e1V0jvjBcJhW0REmqD6QDWVMT1Mtxtacgak85I7mqNFImy6NCvSXFO5CrQ7ng0Go
/y8z3dUJfSLYBg/o3Q6AN9IqUcpuvtEA/U0RBoxmpjWgbLaFScpoptHAAa488nn9
b0uIpa0D+DqZ8L9hXg9pBF+A/E63VcO/eQ8Z+qK3GAzL4Czi3lIRGA9z6qGv45EK
kyO6uok3cJtbboKusLqZW1rMoY+kt6nhjmoA6LDfNZ7ehBPErjADHbb60TvU/VN3
gMwanlOCC8bMJAQ5HLZ+Z+++9Oo5cXjdbaOjITr9griHZbQgyO+KJuWzXNuy79CY
XLGgG8ZdxWst/OAUU9T0tOs8SYyhXcyOb/ut3Rr2Ti+HJLwLTjTSzSl6OuUmJdIy
zH3ZowfE7Gh/Emm3g3bsPBBOEHBE9WHzS07HJZ8MZ1yd6Mf7NrAYH4A0Icr8YQOr
7T+5D38NreCXiKXpE7c8yAacbR6iuoomFpyjdYNsyfSsPq3yCYX+eh7KMzo+kkEI
JxPlt6IiMjXVsbDXZ4UXeGYNbrejUTckvfPY+smgeOtPPf/UivHjeZh+lFUm354m
GpxPaOGTtvMMR74NxKVW1tZ+wxPhSxTwADQ/5XThfypdlsEymjI7r/WZrIkyl1bQ
gnq0IEV49ePkLfHTxsXYnMfGu0e9+j5yfJweUPdjrPzu7hjE6lCJl0x+GsquqTt+
MNGbpmPvKmokZmSVzODHaua5kgKCd7dXtD55T4VQ7kycMcMubs0xoR5yXu+J5lqQ
zVPOY/Bs/DbDPWFrQAPcrQU533TeNe1bE0kTHYlymzbNovGJrZwuObdydfjxdH8D
xYaEhn0FUmyr9m8ZjClehKSHENZWEMWK4CYwtgbGCw4jI0YBStzSQi1q1g64B1JD
TTfSOYpMghqlFtDC1fz1v6qralESGSOkWlSVFNUWtCUQHqNNhgFVu8GpBjLnm8Er
a5/A+VPhUajlTw1pXut6vOu/R3dCrYOKz+w/ROn5QYXyN6Jyd6HIM61UGs0SK2UN
9lxEHHz4SUicnkY/qDKZqxvBvHQEXuOFh7LSL3MJy9yWmSY6udrwM+X8lVabUEHW
lLAk6WpKR6pl4FcSlep8a6MFoiRJAyrs7gEbdnRQMNlnc3xYlO5oIGFX2l0HVJWR
9bqdWPZAFAkMd0a78+eq08Zph+QIVt7dnrINMk978Id2/8jiTgaEuP1PZJ2pIsOr
JJRN+e1cUWoO2IJoI6laMMnM3zjLz4sQshLcHZU1YqRgfz+kYUmf2Q11Ycs0T06N
S8QMGqGb1HuNCM2LyzlLbHYDckMmeBXqkVhs3Tdtm45mK/WmoOSpdPpzj63Ec2rn
SMYxCJHPwYLtjM1gujyK3HlChO5qpmL2muj7KgUgxEkTEmmSB+Igkl2TivQvA1aj
MzBMYCErNgTkr77jw/YpU2haGaDuXZgOPlwTNu4Ns/YVgVSLOuaywUZ8E58582yB
IPwBI4EhS2uHc3IAn9+d4Xs6T2MCGPa/k4rDIiIMq7K++YwCkpJpdQ4xMETNqyUr
guONnMOsXQMnMcMJWlMYkLw0s6IBeDjpKtfRnbnk5Bvtid+1C71NwvsL8zK3PJO0
CmhjDE7g5aIUGl/9nuZzV6MQ0HBDn8sUlFaJygD4JRu4pAi/jTlHb3lwM2cZAvKh
ACfmTwU8dhZdQA2NjY+XeTZqTqnMARiHFioPSG6DlhAv/GYPcfXxcVvk2myzI3cW
DqRBy9MPCuSy+rVSYIfCj2pXVXKceqTPSkD3iX3djXRMFbXIR8EUusqdjYm1cuoh
hC5mV+ZNyqkOIyiUqdmz4AZxVuMK2MzeEUAaQOb1PAN5cHmNSjbWFFxsAjnbckWD
5MvCgwxTR5JJt4KoiGTInU858FxYdFIhokRA89ZYeIGdQsZu2wxj+VQij96FVlEt
TxthIKTGvrKlUjWmLl/eAaTkeEkh07C2xHytHgsxqd6PkdyhgYQY3VttdCf/HGiV
hJ45SDEKRphxKNL4Q0MohSpYbYy3SfHsJMVwV2ST6kqLC8tO9at+aGYeHUQ/t/Sn
hpeijOmCCePG4XFeIs8XcE1+1lPfU0Kn9kNAy9HIvSUp559MJIF81RkCqVD2bLzx
K+yWSHAecnmsa5blphICYQEBPCnTdfvLGT+eErrJiQ5YdXESULXW2WdlBJhWnPC6
hu/BcqXT9AkNj8B9nGtdIYU8PkNW652nzHOyKT7pBu06J29COWYNgf/q+ifbcBQl
svmFEkWshj3Gq9M3PocAETtRAcdoR8TXQcJALemO5Mo53pnzo7HqwFwm4egZ7yYu
WBmO/x9KADm1mh/OyiYM8hYtdeq4H+Wolw1h3QWQTqVN6VxAffaI7pyZ/FTgeSlC
oLAvJfRVPySgk/2KR6ByR1mg41plhSRa67YhrR21TlO9LibtXnurJvl8UeiwdxsA
LLX10a3n9xrNswqpvgSj1YjX7IgL9AyApGXimuV1Sm2oQ+83NySW6Qfo6Z+0bGOk
qkLIFgKCdVrlOoTHmVZMjaY+G827J4w2RmC7iAYL3LmiVOV7FQcY0ugZZqpB27b6
7JVl6ymLv6y199lQJyk9RIidNImQ0Q5TyHGRjqZycN8RInPOUML1O9bC3Zuj0ZET
umMshpBhMRtpcXz7G+0OfhnSIqb3q18A3K7oRYOB+aeXX1Vud6GE+lhj6BG4RUQo
z5hlzw9eQjDQ48c3jIOB/rzcgkVWb1/Q17h/+WVRvOWG20fAouZQSM2D2f/NtAvd
zPXC9kXW6qFsLITO/0xvRXF3djziLyOexhqtOgc8JV6S5cqON0QyxU7QoyoJI16O
zcJD9tD7qFN9aLJz66dx4Z/03zVKduxbzKUKR1dUXphwbDVSTKg9iWCmfl4gYKaN
3rx6r0+Yrnk9gbOmdYC5h7WrdNpaoQwt2NyjqYigCiCAPd6TmmavRMw4m5ArZWM/
y9yQDbUK4dNytYtYsK4QfnmWbG5GcRVsnbWWFvvcmGgoCMdzlDzjcv7GT59PjIW0
6xkxWYErujUnu1trBRENH55lEk+YxUaxs6MS99clURtiOdt3k7I8VIRCs/QRRUVe
8Drqygf+iyAOaL/jo+bXjnsZLohadA8e7EcbDJKkL5pgmeHbqEGmNPq5LmlA/pwb
/0+yhptwFk6OseLG9+ySrRk+YnZ+i/AcH3yFtSUG4Eq7pEGS6K8feeRo+gW5MFOZ
ib/Q9DIsC/Higu8FDqy40IhDC9j2K0tajlGjsH3nrvGpcN3/GBg83gggizN9H0Is
p38B00R+aSPrDkpOEFeEu+2lnibtNHNKXU45DCvKCU0EEH4Ibq6nSM8s9CGYwltX
EwdLFI5LUGZGew354IK1rTlLVGw9nLfHHzWIQKn7Rj+cAnIuQ4bGPnSubMElIYvl
hlbVCOC4l8S3DGJ9Ou3qE2kX+wTleZFcbEbm64e9bqtt4PTBUq8l1fRpLerFrP37
yuzuphhWZMB2kBSXFBI0C8TVJUNyZRZIVEeZJTty0cuBGE4I4LiMUHhbeqk6SWlv
jDLqbofbA0LriHOEvips/+1dYjYdqfhaIfMM11NvY8Go1OrmljdfCfNCPbx0LjqN
77oLQAYIgp7HWEsdcCoglekY94YWd8BixjhghzJiK/tyaUGOYt1Ad5pv8j9pTm9e
II9rKkKfSCXCCsiLzA0HavpXHpdNOBsTKzmVZIy4VGEzJUywAUgj29qkAR3tP3uk
YFkkbnk6m0K4xxX62C71GPMfrvkLpbh2vyjtvkAgYxGfnE8JAfIw/QLumHuz9K40
MTgipTpOlq31e2OWMaeQLsL2yhW483486TwrUnKv2vorI4WWVY9zB8cQxRrKM+Hk
x6/FPpRGEsCy6ObyOXQJ4yOXMOYjhrUZe5aB9hVRlRbjudq0jCM+O7dBGnukEwvN
xsosgMAXJsL1+gLwnNgQjji5rJVUOk7nEW4PR+dr+RRs9T0VsQiYARgKpGdhiNx8
/uJ7UKO7Efaag/hn26w1oHtQqjtkJtCtIHH3uOCnHKrgC/AUoEL7PzAxtfSJM8cW
DQ13Zbqro/ZsDvnSTV9RpUmamk6LTIPmsEY465ShQ79WzUF9/nEqODITGPyqvbhO
FtuVGQOQm+s7LD3TqolYcoP9Rrh966ZuUcvXW9Y4UZv/WbJPcui1kD4M4QAPQbNX
sIRh/iVBKpRjolp/aMTYrB34gmhgbXNzMB4tTqA8OXWiiiWSj+s6Zd4mLHgSnBiN
yxu/Tu0ZjMiyOB/lFigrasRGxEgYETV9RIQdN9l+28MuJ0CGfBTWwAMd1lkojSu5
UIvdSmOaDc446xf3MI18PcFXaPzqVkMkds7xHk3DWbB17tT+DehjnIhgeZ3B6ehq
LEeOvxJIJW3c1jd1VGoy7DYYzv4uPCGGoyN4iQDgujMKisUYHQ01+c8phE+MI479
d1oYxqatfvqJqNnw2AeB/FVP5oOs5X97AYvgUiCW59f+oM6RBG1iHPl2A7aiGbex
MzBgzc03DKM6m7It2ex/Fj+Zp73mSPNLAGdjHhXS6OQBDFrH8Q6DlBrOIJKv1ojg
L1qQ/Ubuau46oxmExfI0VU5a2W8n15gA92pfViZXMGJ+R55ILFX95rPuAgnrkaC3
iYw2BTw4sFLjikGfC1ssJMVjV8gX9aiKGQcbuJCvWm/Qf8hj3pElFfG56yFwsbH0
F9N7HB3+G2lq3qDdvWBl3FSyjOJ7r815XAtsTLE8AFrKDpOddS43p537PCmOPaEw
JtPz61gZrGgY4Uuo872xfQSygZ97eKgJT4iij4Z413mkv445C9EyJJq+XEv0xviO
9dLkZimhYQql3lt0A+jghG9WwsZq57uuCXVxI+NyyF7bocEbTJKjA7Ek8ef1xf7D
4ifdTE/hUIA+NhAYLoRq4h+Gh1LhuhW7pRCxy2R0LCDMRVymLqs5QeiLck95xmmL
4KChCk6YsgD8VxASHrWP2T37w5b6NRMlUdbWZ3bg2i3I/CPEeTpaZOoM2HzCU5wk
O/YBEFEnrF8TsSINKtGYg4QvANQRTrbkadbX6fvf0bCvl52jC/SECXlB80wer/gJ
QjJRw7CzsFw4n80F16yZ2L1oM1P1rgNAOm/+vUSfGrtcBpwDKAThlBp6/we6hh8/
eHYrdC/Lq7nHsSF+bGKh8gvuKmpdhKZmB7TRm97LoiY2BPQZqoK5X6tkIGB7sf3v
Adhou3DiHmhulX7m5FlEN5UEm8HFsdqdAee5yimOuQI5CHbQj3gW/aERTfNNEJeM
bRklW3jSUG8bP4r/Ij5nwNO/4NtDE+1yHGFZGs4WeeUHm+XLi7eC6xcSyhFU/+U7
WG+0Ay83mcs4XUSD8H2aObrMBp4rrbR4WMeMM52aU7Nkt5MBb4bLVMB5iw77L3AC
Cg62+ip5eKRCcvDNcqAlUaLlcRGm1o3JL+iWXVvO2ROiJLo3jC8UctQd/D1+/1Ey
9hK91oYhSS/nWSpxdponLzavy/oeIMTWXDStmS9iG14UZBFI8XGyMKtDG42H0R34
n33FPZD8myJQ63uCnTsk+5LSFt2LadI+i1/PmAw3kU5p5klR3y+yrmhuYwW6jI0U
6XuVyiMUz4lbEz94dV9BbSyh1UPT1MePjZ67I4kKF1SOWtuPSW2Z5+IHchwpLA2Z
TcmY5uDN/ngOBAW1AoQA1gu7CeTOCcsRadm+TZwO1kou/g4sZ3z540rjvSM23q63
bXy/pU+t8l/H3HCk7+46ZhDcXN5I6p2hC/DLA8IrFpmB/+8hYWYV+Cu+GSyPlcg7
SYGdVsQHc8hQdVGXIlw5c6lGcr1MQ7stJ6tH65oACyFWk2T2tlGlzGww4cwjLIV8
UbEoVPKZbzNdo6V4JMGTs1BxMzKKjN9JoUx7y/4f6j2ROL6urf23WuSKJ3oLBmDv
z7Z3cLN/7rUWRlgJtYPvzSptydIqDqlav0A44g5L4jfSs3TyLMhLqBi8YVB2Sjj/
NLQNA1nGf1V/wLttTwo6ib8YdQu69J5G1eLsYc4w2HtUcKbXCxSrh3UNO3K4xJPI
i5ffdWbG5T9iAI/RRjYUAINis3t5jsRbkE7dZ7Qu27/k+dyASJRgCovP5pBI6XgB
fK8VlGoz78jnjr9Ea7hjGV3F9gyARCG88ZrSPtlRC+y3DfLbUHQbm6FHtICyzawW
olrUURI5NCLd0iXR0f8oe/JIjxhNSGFEBZl49tUwQ6VebYu1F8ZAyQZi1uR3QqGV
bHaq/cTVwevznpFjmSE9KysYrTMthz9O8PJ9Q75BqGEmeKlwNw0yRCTLjlZ8ASDq
ofJ9UDE0085iQGs4PtAy57O0rc2TOAFDzq/77ShmylVpF9kJOcWpIzg3nAaBLukq
tV9iIXDuGV3QDpCb8YyzQofqt0EY2t5qw1uW9cfJT48qg2mtqKS/e5O/DO+gmhQe
ckPbSit1hwYWqB5QLER/2TF+iYs9Ty1SU9P/G9F5y3NftTtDP6iLflukv0S/NbAf
4X5r9zvE9SLZ0cRTigJhzxJI3BmnEJHUX2phRg0WM73ExOKy5B8xdbfkX5mFfKR/
JROqdar052eEEn+uxbW+uM2Eqp81yQSy9frZ7EBNB9hxCNo/1M9UHDG52HNcDsbN
1z/6RlSbQ8KwufxksOOXYE+nUMA2CSsiAfGaf8FL6Jo9EBU30aJTzS7H4P9ZNuug
AvrsJHEsKCHuh+p0VdPi/SFdQ9wyyPvOMta52uPGb34gO9vyiYkOmsOJxEIeWOtT
MBui4QN4PvfYreZB77Xb9BLaMn9fN3P0up1hg4KyiDba2m0nVYegSplboCR0RpAR
NnPzWUl9OrZyoOKzKtMSA6xu/1WebJZ1zZsrmk8+RWfrIg3gdERq1OfaxMPiiwg5
UfuqyKp32nzSpFUlHb63/yXEvtZTubLU+jZkJOoCH7NbSawEai7Pl1GTFgWmPlyF
429Vo6fdLQlBkhNRHISsNaftuulC3oeZ1ir71Ubc8dO/PvzaLLclkvwNdkqmSVlO
Mt2LtsUwMQy2fj8wOCfziCsk2j8rzKIccYM/e3TdiVLQnkNzW93Z9sBp8w3Hcmpl
COFsklo8aUNZ5Yw+DhSgwkltJ5uqjET1EOHNm26tIZ67JCijnQTjCSkfQeBp/gwd
02kF98Q6iuEzns8xY88A46sBlKD24xjLPer5sekNcmH9gr1VvRlp7SUjIndCcuwS
gBh/BePI0bhOcVXQlK8TsH5mWoD3UeBgpST0U9hZj1M6hG3lZbSlIvKNt7URtlxV
K7yQ1UF0QVA/ZBbz2WJduc9qujigOCX00C92hFO6Dl57xVxq+2zaxxabX/J/6N3Q
6iEQ0/PMQzBPJ5T/o4cLBHzsl9kxOW1hfe6tjnJHQr+HzhCLvnj5ibALmvfMiUiy
d7S8ipKIeJ0hSMIoeQ5GRBbJrFjsIaosSIkGOXgg/KtSUm2cj+Cdb6JHL4pszkJ5
rAdPBam11skW36/t1ExFWT2qVmFclxnkByduGC6CCNmM0620mwAJ25tpH4MOAovs
qkRwLT2d2iaqyD5YKBYIQInsLDnfvTCD+YEt56PsqW55EckGex6OFLKEsIppyZAG
mqe7JUwvfnCOIpUc2+wTcAHgQFClfinRrBivaPhlNGLnYOl//qIxu/+hFB92+jLV
1Fe0QHYgCVrlVGFPYArCoPni/70MWRpFvShVIJ87Gm5s+9VP07GvTfom0cZ4EYJB
XoT6ueOJHb2l03XWw0jyyYj32mH1bbM4IHguuvCJ6JZjgXUX29bYg6Ic2DRhb0+0
y/JXT0spOdrhgZJzepktBqHhZ4DaceUXJ/dq7gv2oMX+FzfbD7whgzeTLTPai1ce
6d29yNyBDrrz8q4dQFmORNMtXQorq4bg9H0pbUFV487xNqBZzZMVo5YZe8rlHfB8
cqPMKdxPzthqa+T+8xwKPx/10txwSs3mKALZ2Bck3KpVKmunx3kGsfJXsxtFF8fi
ZTm9j6rHBP7Gf69ktTVuSukOUQHSaMGW7k1R9pKFlxlHeHV9tAngvaN6PZw8sF/O
nOS5s6gxyIBYfXqQni9GhYnIg56wUH1OLOAsxC0rqgZ+OKAuUp3MZ+e9OgUWs29J
7HjRyzbrcxRjC+3IEsInT49E4F4v6HkG09UyY5lax4JlNoeKyx8LkVn7sxK0AQYD
QYVOlcjCb09m2GLvHAwdsvqt4Rj3bUWaNfIB0OhgCo3/MtQCh2gCDG+Dok0mT39S
PPiXuqmQayPKV39gb+ssLeFPeixDHwBWg+HbYrfR1Cn76Xz4oT5zCUY8MWyW4CUT
troMYQIuUTKJUN+2Mdh9g/w0HGFrHLu6lg77XsyqJx+S80rLvBTJZ6a30bAtLVCJ
sKnFRPpUdf5GHf2/AKDostVs1rvvElHGIKI3pF+djrH5Nn4A2SCBmERmBIPUoQX9
fp8rCafhzT69CEthrqQ4NXnWHcQ2qQzKtPWJSycOA2wJJzxAnAhxUfy8gEc4Hz9s
Bra68UKuNcDnMB/uA2Kr7kSrxQZkXLo5AB43u1AjPF7A1mXbOSVdba5NfnE04yxo
jeTnAXNRg+eDkNfQviFob8P8iink5HJDn5IUlLT7pwblxIWaSXsjgHWp65N71wn4
0XJ0YSP6hiF0AK/SOHgL9p0/6yxfiVnGxvmOzdz7oXmCLSy/AnJ+nV+cv8nzGPkO
07bYrolWJfSaaiJYwaLk9ng61GAwnKXSd5SPATBA6qMzBcDkyhGLiY18eTWMPL+g
mE/N0zAbcbUbk5aDw6eT1bVSZrAGd04Mt4/kHjyI6HrRjrq4nsp4SQh3yhQKDWZX
aKF3EpTbBlJJRVoXGjZcgqUc3j01pMxM+wIs5Z8CLhgR04QJguY/g019AtsARk83
xzJmskXGmVk81R41LlrQywypwIDVyqoHAOWYzSebxbEkckQoB8y0319pZwwdzFta
blSbRHkfcqdH/FfTESxClNR2bh/W/GE69Mh5hmUtTrI9gq4a/DP9HcF05Zp8FQ3w
2ctAyqYjScK5e439loAKwAVVE24yhXLYebnsDZ9eMKitOk/vAXUu3PdTFwss6PiS
ayel51wT6Jp+qnZUB2WSbMFq5OxjO1cXrJHMDr3VifvbvXJs/r1U53hFCRymX6Zm
4fcLH3b3j92rp/tDw3mDQQUg4bajQRGBC4c+7AdLru8xmVtjq+ub6HTZhnYEzU7H
3VMhN3KivsA2QML/dYiavCVBun9myDaJARUjfWfL1+bds+fNi7JQGwWg2drOhmAO
hyiG2be65uA7KDS1O57gkt9KkbxItWa8oux/39XQ2amUncq3nbk8ggPo+d/G6UcA
UlfmQ1xEMqf4gED11LXMP5rQECGDFXlDfc6MHQ0GUK2a8rLLelpVoiuqlt0OQJNQ
V+5/lFqmKdnYg/+8sMdQHcAJD9Cia6/ouXw0Tt1uzuOLgpKU8UL6bV6K7XUIisFs
wzs+po376cl0cv5UxA2Ga1l+HJqLCzC66WBegyH3GfCvQ2Qy6Y+6vX3Zml5PC0UP
qLWK4V4sP8mNztuD+YNtOPe6VCLOmEFEqCCrPfbzHIOaYztBOdwrj0JyxL7U81oT
ScvsM7Mfl7zghn/WBqnkOr2M93wPRspiy7OBmLng6KeCI8Y/faOCIUtrXH2f3EkK
lK7ZEiI7tBrYPeUule8G5peDdFGXMUB8PXfBQDITfXiy6tngJiuQ5pcTj8mBa3Nx
BnKGIkyfPHBczB+yKqSOhGpw3nUJMifNPGPZk43DmJQ7RVzVVGv2HSNgoKZvzHmq
9hu1dDLiZpDDz6wBPYdUBUf8z/pFkJdFTcGU5eRU/h/Xj1agIMqVNriJ1OyJCFVu
GmkzBvEfWPwJGsTiyj7S4ixuiJgfHW4yjzWaVzANWiCvi3Rm+BONRe5gW6egXZ47
ohQiHmeL8Ap/I3zt04VuYEi1gvEwzmipFl/Av2YfHF93bhrsGHX3WrTFyyA7iALf
nNMOPX1+tE1F+9zBQDleR+7kaAeOCrEZ00nlv/sfAyNBCzo1tTPVr5h9SNgEVPhC
/CnC03lFbZt79F7YNOPUMLzNCpOs84bBZhCpfSLiPQ4rwIUSwb/mddxOtz9xz4j+
pr+uZ5LmqSQBOB+oGCxBuo6oXg7ZpFWQUlcW+nvQvSPn5FeE8uRNlvs9uSBHTaQ9
hHGA0oWkwRIlr22Qnm9A/zJlkZKpiT6RfzIZbkFI4lT5TdhJWSm0fimiXGT+guma
sF8DCimJ0wDQnsC38ik7f297rp/51kCYYUwUgspvTD9pRxBAVFCheCPch9NfoVP/
XOAIuHs/Jf/OiNDZB9p6ujnOGZ7oSEOlcWnuHSPdrireX7WDcPBmA6YdIxfSAM+f
vfdnE+QzzzC8E4pz1bQ6g+2iy83rjzEYLRJO4uOoW4MgnnddIv3pxjhmT8+uAvks
JYRobMB2InEx3b6RBruJuCz/KDf98cTn3dcKzqxFinmE23pEBNgchNSDXkNQjQZb
joy2IBohZ9d3UGY4HhrKRMp1DCEjYn5UpxQcCb0W9ubtlj5B+0frS84be77noGzE
NEV/wdL781dSiln+r/7TJCe/H1GAHEcP7zDfCHp2GO/QCA7u5vhJ0VV4oXmw+ffP
T1zw7gJAhCE1O/xaVsVs3st4RMHvDI9mYwpTqix3zRhDf5WGm9K+bq/JkTF/Q0Ib
rUmF/0A8vjo4/ZGVqpA2UKlaQoHzpXt1ioF6/PXsTuLHxa4sL7DKr+KF74Rd9VDW
y+4VYbXRbrdY7UpwXlhQnNeYA5ZFo6Ijgf+qqxpy5iJiNUUNYwOL7DSN8Jx/1vZV
9+NGYTvXwBLFHKxJl7ggz11ybisCgDZElHWLtT7EM8gNdWdJTGKWS3q+OaV41/RP
erq8AGcHbDeGFFCe7G37E+IKkdpHq6KXHDWCXJG6eS2R9F8MhNGHA5402Y35zZvb
pRe1lIJqt44/L/ta5NqqHZk2DnFc4C3R/exL8c60W1vB4qDvOmkfnQvH/P9cy6J7
F1rqFch7uFf3xbh5qGYcFHOadoxYzYCW6zYsSx34JcrQCbdOd3kQM17Qt3OZeOOm
Q35F/rGRyKXE4OeJbjHiDLx+vaAgzj+SPEKYqRBHTkW5M0Ve/p3aGQPqUqjWS+xI
aNHjYtAdhXwyOgrVCN76/AnSunKnm1gIgL283mVgmywDhSQ0BPjQkgYDYk2edBVe
zFFWccdFTG9wLFXB63cdTLHm+1M1D4ICKEkdCGCkwD+c/W3fccgT0Tk7FqNmlSp7
pwqSnV6VbQRocNYBOmMpwrSx7raW1gYmJHv8uYzzTsgQXuS6Nlory2SPizQMcaty
5u3z0YzBeUJByUbvBz7bfYBejx4FII525zJsj15qKGpFRoC7d5ugrGo40qRyzWND
Amo4J2lQJS9Iyi3fexzwq+dHBwRr2drCHezWUxt0uRsmbRolcme3NLzCIrzn0dM7
FWiQ0Y0M+OTLR0KL2cP+0imuFs5poY6JC0rTm37xRlSAwhD1+YlVm62I6tPO/c5u
Cl6ai6/y8hUAstGs6sQvDJ+C64XWwdQ+SNm98ryZEApHkNokeSfagTfXO2Uof9oD
IPJBotWct6wqOnuMLfcRi0xFV9FUD82P4CdrBgbiZjtJYSMb9qtLNRch1KwCQKHF
WrUjWn8zcuWt+Mmfy808+bCFt/ElWbBgf6JU7dGlPxged+p4CEO5DPBYmDKUecFZ
hWUleJvByJ+xyM3odR5GkJjAdsyVJWWiO2Ps6RaW0PG4EtpoB5JxJEhNEPIeOp/d
WYn0hfD0WicpdhC3xQti5PiYUjkHtHMChzO4ud0jiaMO1TXhy3sYpysxTpkr8tZ1
9a52lfogo11FWpR4JAliaA+uItXlakvWq/p5RLlqeiJCEuUw5RBNjFvWoOTJEBzV
kjeCzWAYMelvBwQED+j7J9FbseJmnZxa7cL3HLVNfKda4/NhluAifd+EsG8yVNfh
V091ZDfhfInqUMTLSIf00FPneRqwgGypdnYaUiTnI6d7NAXR6C9Qg15p6clxyFf6
P2iYJ3wuFGWa3s/9exAziQXyOfCvW9D+xIixLVhE0W9/o/CYYkIidsH3+CHz+is6
fwkoop1wCVx15pqnjLiwgSwJynfh7TPlZ1r6x+6BVue5PlN5RUURtvRjbIriQhtf
LL0Xh0N2FxHJJvDQj88ytq9vnbZYBnYYxqCKQdI3TGANI9jb8N1rXd29a5c+yBqW
fWJEPq4p8/F9DuKvD8aSy4eyvYk2994L9H2TzdsI6AdLX7USs2cEeME5RWYBQaWV
Lpf0bVA9i1SN7TRcdRujh6XsKf1I1sP1MgUgt4Z0IKhAg2JFhub5a8XnUwFmqPoa
NqyB3P6fCJWcVZhs+nSL28tZBFqN14pMAj0gCy2EoUS3YP1fH4E+nK8jfMj70FrT
W6G2eRRo0wQybxkAtQQ07d+gHr2f+nwTxZf89fmfF707QeKSb3hwrpvZ8Q23xdou
Xyk7AhfpXPTsTHyu2ST7UcRfQ719he6JDcIaJtXvqB7RCDmDCOJ7flgX6xk06HxJ
0+cf4+jLCk07p2s+6fokSOE5ivemn744LyGBAT1swi5YIe8TQi5uAj5Iw7vXzxqk
11J01LTUAjqmwM3eT/+O4mw34UAjCLkGo7CiieDa2F8DdPUv1e7pSxpO1pvvVHuf
cu7Q4dVvLJZ4iZXcDBsKqhy7Gjc0WEQYJokAw5yOaxebwAic3Vop4L0UnwEFLRn8
2inKN8sVCWiZSkjxh5ftBEf/vjGQVIRupX0hAyXzu0kq6vBAWBVNZ6pLKC/u5DmH
/sFvEJBBmnpYYufhQ5d77UNCVwGQ1cogWbmm8GqscoSGrkO1MZI2F7Lf35xKj29n
Te8EIpHYOg36uNmY4+xrofta8yIXKBLFzaGh3YOBY9TDNLr0iuVWkzD/SI/U+Z5m
uBXHXBPLT+u8DX/tqBdQ3rCdWzNHf3XvWQg0q/dAanP4R0NujlmH+u+4rddqt9GW
8G9y8wcAQXx65j1QIGLiaxNUG+1ztpFVwUJfiFyrSDbr9qA5NZ81IL7DIsNhEOYF
somav/x57d7O4j62kHTTU4EAotRxwh30rrFoKoC+6nSOfvIyYAys4oLnlfZYLHJO
Y08DdkDbLNSdvL1fzftrY6dItlmpbFCaKnf8bbHtAsFwO6FQpXjIxnPCvt1N9miV
mINQ6YWMDAjvN4/l+BM8MXXYtu1KYkBK72ecOue8oXucah2ObReu4RVZY7sH12MH
vE0LymOqc76VHPNTfSueVP2w/a5ESN1mYAJqXS30hh5ULIel5ifSXWnMx6qOSmHI
2JL4bZrRGyHP7wo7iQNBlVC+vFag+0FRveh88VcMUPyHcuTR+ylB5vmtERo+csfA
ZBHz0VT+L8Zp0Lz000xT6ScdALqZ5e/VFjrFqx/F6imZBmW7/B8ludhoSI5A8Tpd
O3s/l8BbPskfzjATMEmtZD8x4H4LrdnndxY3Zk9y/f1ia7MsSCVfWpYq2GfKzejW
1/W3X/NAZ+okb9hxR1V+tgo/QTCMKs18Wdj1ZdTdL0/5VmHGWfRFxVsmb6PmnTyN
EFbSqOCQHHGO5Qnm/rQ6GJzczv9e+hp0hAgE8PRBI+uCpBb1qgMbuN8nP2AaUKM2
64VABv0kodIQahEDXkqUe+n5oxTGdJeU/TAdTnjsXur0wjCJ+KBpsIx+5p5QvBlV
HSrxoTcxdgw78nELSL3W0fDUXKVrp+E4ReY69mZpZcEzzO4pSmWUKmjuWxyjCNAo
aZh7b9AmMhHPiVAuy5Z6SXvUkb7jkg2J52BGqpmWiAjjIyj233NV+TynQ13KHTGh
4IscDEV4k8qmdtcQuCY2zT3KhBRraCeNAcH/c4Dv9ko/HVYKKukHtWxY+80c7rRQ
zGhnM+Xp3ABtGK28vOaHSYG7J7mWeAc2/AWJbAj96EZU4LfFf0V9c7NMO8D5RKRr
WlGaN8kuS343elTx2eLHxCETnl/+rBzQMP068KstbsCDdoo0GhgFi0Qf/+OJdhTa
7BxEwF4cpHuaWjgjNr3OUKr9OwGKre7fe4HBAL2ZosXib3dtmbL+7uiGZIoV1Fyw
PK7mZr52Gqtx7xCKe5JCrMCx3UL6hB5oafS99br3FoFbxUANAGqcLV9zFzYj5Hd8
vNcJwy5gh4274IW3TjFp7qFg09FCcyxewPVzKvZBI3QseN2TM3ZiYpkNSh0bb7im
6qwNktrhkqqhXwRCQCbeXmRW3+ShL0pz+GACL6roiFjAndrn6FeX3AcCaTfNTlQ8
dJN4E4o/WqF/49DOAgh+W2IyC6dC2Kyl/PUTXBzTndlsVSS64afhD4/W0vx0AO0q
sjQhNlBseF8xhzaB4nT4d/TrDbXSeB4/Kx7eo0HvqY9ax1ADmkryJubWXLBX9/b/
ygmvRgnfFMp3KA8RL2oukJ18oGQ759ASD9fskffmb0dGu73PULOLj1OvsZZNyQOU
MQFvFKNFwiAvDHNrJmZkS75GkxY23HXedFfo1PK9Ud9hVrDQd7/7INWLf6J27hA8
hvoRe3ZDLtmmxMYsS1eak14ZMyJLUmYyGSkVCEs/bD3oyvzi1lvowMmR8xqS08ok
+fce2DpvbYPIl2tuR00EpNwew+cFEmuKP4YmaJi68tLDj+Y5/gk34hDghqIdlQyB
pY7rdb5HIEMyHCG1Gi8gu7QQP2u1uj9jpQ1bwU5j+h0EVLGX7FI3LCwhoAz3wx+y
SBOI2tSly5Y5AmRwf8GEU3OWsC4sf7d3EgjXDq3orQaNA8zeCuFvtz3xQssO3fv9
QvEs9cICffFoYuEtMHMaKUET7bSEhRvb6IzhEYtrdlefufiiRTPvafgm0URweDQs
9UpkRocZvXz6hD65y4/adZY8T+zfHKgXEVMAPYf+9tFVuT4kJnqBVs/vbUdgQ49W
K7hnzjWHPHSUcfunymQ4Vfe95dfdL60rFTvhWLidTx2/yWAkgvntjWEcGfoIcRnK
O1lkr0CUNwglIvq69iry5kMBhKceCNwHAY9l/K+Jkr6uPl7+Z3BpSXhC8o6HnSnK
KjC4uwMpXr+JWVZKXCR5FoOJGpiO6xVWyVIPTP8mO/RtHVB1PgpB3g5qGXa+cW4x
Tfwreov/xQm36dedyA3ww/eVLHipqm7syDxDCMPNdEPknhCNzYtjFKDEwuasD1ED
bjooVXa8KBlJI5KN2nfxDnnt+XENVXgESmBVhDLSD42HM40cK5l4hN4VturgtDc5
HKJkKLvMtJjQWsFdftddjyp+qjMlGzEsEEfpGaagaJGn6IikHjW7uIBnnaLv04Lj
wyoJFtd08YrCU7fL66jy08hvY3nmCZI2//GX3kyP/zh59rsPp7iCnQzvvavXK3kQ
pWl3HJZpX8xPl6+TDYxU7BDIJiUphfIL30GYYCNUhs2H/H6OiZHVvL1MC8LSI8H5
7BA6D3ybSkbAn/p6UUixPOGaK6YyF6wpS23nGm6An8N7KaDU4X06ymYjJ30cnv5M
/NpzomsKzTvTpWkGZz8Ci5OiGycsrj/3EoZI1fqoC9dWJLVe8wE3vTSBayXclk08
tnHDdc+qBbU1oAeuVrmmUyha2ty6JkiUpIIckaKjYSoSNIAJuCsRuyn0DNSDIZUz
NeLW5jlfB7oL63Uhe80YMN+zA1hwI2YWAG634yt8BZLwcaB12kApt9oJSdrbyk2G
fXhIwEMaeUG+/avCxW1nIh4J0wt7Fiv11GrsUVe9KZO2XcWEsAo0T36DoQKgnjJL
NdEQKIdhuXwIm8CXQGO+1pazxXCrYn0rFS72mY5Po4Nvra4UPDy0Sx7vO/UJd8U4
rGWfxiHndgz+Q0+D1m+pmieGGs9LbNPI0q+Qg/tYfr67QlCHo8tLImp/cj04/TJ2
Lp5IL6/C5NLSTvXT4bBmMOvpwIcCgo8fJ+WqkzICc6CrVyQ1j84CNonuhASrlW4M
GD8jxhwYP/4990g2Z7ZdGBRZf+7rLmbJq+TM5Pm7V8LUGLtsNEhU/R2sFSmidlG4
x4I8Vd/xaf6tU0tBxRRxK+1hCFhFqV2BUxBws2NJXrh7NbO72Jdkx+D2fTrjNmMQ
PPH32oMXeJmmlLcyHO+Nk0PSpOxMzSl8INGEMJVj7PBGgXLVnTOs0Kz6gnxUUQ1J
/+S16W0qKXNHdImRPSz7aSKAkFWi/ejvJ/HtIGnnxyD/oCaR1WLHVFJyRtPQkhBy
8fCODTRVo0u6O8TXXRiu6M8ZFyyjgrzVzRwIJL4ZraIScfDDKsQhVacVkUiT5cIB
xoRiEhJkwRWiZq3c1c1duurkliQ6fVkRBOwqcSd1Bq0wHlj4R8NACJdXJYbjrvoh
qHCKW8r9qworqcXUU1REtVDUBIEfF+lgrp8ozlP/WlnoP5qVRHNZWFbjh/ihWBWR
FjXX2hTbd4HNXi8J67w4g6Umi4KRgfMA6fJLo5gmd0lPn7EblZG/w5ciqp2eAeNQ
YWa4RJ7ubSBItBzYAv6FpORMsvhRAcMlQS3ixBmb6kbu6V1VODRemAJbTDezD1G6
zCDJezArZqR6hybABPwHv8SqEApZH/6bNJwuP2xTVF8DhPs0u4SQb7OvRz28AEFz
4s1tAviXkjzmVl5eLoe7Katy+2IVtj0grQOedFhmLzdBpV4gpE3CSqeSV7FYaxvo
0sJTRGoBMUVOUV7hgM24bYFFynhz8TrQyohgcxzcZBJyhVUZJwC1ITdkVyGi750W
urpEXijLNUn+FgVTHQpxJjbOiaVnPCpES1OlzBKA5j84Jy73Efu8B4JeXPxHoZZf
qDfWyPK/pO6kRXyDBTDmLmVc0AoIJ7oOTc6cqsBqxbvJ9hovlEQgKwwYZcyaFkGh
19t/WaA5f4v+CVLx610dhPUfd+vuOwmPp+07XBx6Ua+LvhVgyU4mxDf6RymO8BZb
U2tzUG7QsADw4gn/o1dmlFfB8HFx7i/vcDWeK4+i/huUywpZwBdi491OaDvN7Tz7
5WRIRI1xat7ver7YZ4MTkRlJP7w4f/YcChnllV5IEsEE46QkettlGM+ITOLF1RT/
itoR6oLSYHQ/ka+aW5x/ocOcTnlXAhmI8y6cGuaF+AUeivBl0TX95246461bWg4N
O63ilZ1clFImT+59n75CLHLl3pcUNScZAQ6JhrDYr0JoGFTZDwYj7kBQ0T0eX3z0
iOVs4WsZ6Nofr/UvlbV8HJVTPPQZLcBXK7sE6NqXQKMMgqo/PVCnhoDjBwmyEAcZ
GK481kSRmYLljFTmXMzlmkZLRqW9R7VkwDZZNSa+7u4fMwY8J/0cldbjjz5didJb
JjeGFuxtF5P74y3sfhrx1ksJpaz4Dwtth2RcXQWOoAkw8wHFKhbnpR3OwutfyVd0
0F+UOh3/38A5SGd9sZ1RFIkbu0ju+SHTHMRF5Fyg+SYoG92hOvgkB3dK8cXDvYPd
HXKDS3G3C8oQMMYmIeci/H/sW88+ijSzh7X9CZn8za8KhEuaW1CGqbILz0XZ8VNn
9dVJw4iOk22UiYshmLfWmJ1Lk17exMqYxhq6ac9cg4mCxjAihE2HtzrrDyj72nYw
zujLo+lqRVyWuQD9Uxr5+VpR6N2OOMOlsJJi0KjntruZZlg7/tti0PF2UgVGbnCs
5YXqMIqFo8rT2ggXOWPIQBkMbF9YjPxeZR5YJO5Y7dLCipkDsJtPr4lWi5N6duhb
EOztHKsTMw6kKoZ+c8i/tSOKslzREbipUnBvjK++oQB4uVV99Mxaewmip5Rwe4wK
LeCl2xZC2MaG+8HxI505247nmmY9lQz+iE0qYfe6jlUjwOPtiNA5JMNRaNwojhV2
F/p3LtfqdmTE5Rr5ZaCTKgl1AioE9T0y7pLGWwmJDcavtUiACF7nSUiKlRhH3OHs
yUhNnkIrcIZKtxtI+JW3nHBdgO/mc41b0zaLebzSWLhR4nOrd58oBTgG1Imk6U4z
i7rgwgcvhpIfX89o+bD9PsARVxIjyPODtUTepjhJ0PMvGfmOD2ZSb8tRyTxYEJBK
N1gtbRmtA4zFHi/yI/oDOQgkGmLoGxPqwpd2a/ZzFGKXSn497ouY+vqjabCtRxzu
nDSehKioOSH5VEqY71/8+nUf36tevY0tu+OT7DXFvoWOeNCUQxM0aC/v4+p6Fdmc
lraAcQ5QhzumjW4zT1KeG8Oub+InnN8zrP2HABu4ShhMwEe9wKorK337vQQzEvM/
5iHQ3V0C5f3aKyASLAxPwIctfQfVZieiTI83zq2PxRZQlb3y7jljZbQvaKFUlOLD
uXjxKHLyxjWvVjhimDqyEQS3Vuw1We0VZJfSm06wHn1KEPl6Wkn37QId0ed6pk1m
pXgI6anGg1HPS+hOsAjrLh5B/RdrVtaZGVS5szPO6q8yVgRNdg0G2ETAL4e/WD6i
H23E2Cj6vdyJvMDYpssTXO83eryy0B+dipBviXl4qBEJlJ9qZu+Fr4eaDOY0TKvQ
Z1vXt7SseQ+R/2i3H46ajHVotBFu/pN3rzi8/ON3A1J4UOh8OmWcDVubY7hre+a0
Xxc6rnt/lLstqfIjuEA8/psl3wCfMCJ209//qZBWV/3f+PysfjmZ7WeXwfV8SWLv
8NdkDgTQCkHCSD2i8L/jDzexxp2ihKHQmOdS/wjL6YYatHHLa/e6mIsyDepm+Hhb
4sDX8TNjD7bZf9yK6/DwQq3Kwv6xFKvHsBtXUrb+Ec6fCuxHYKoQWNBzUxkI7pQU
D+FUd2+G+nkZFj79jW6pL3EwbDwM0E/DuW6/CqqBN+3pqCFl8NG4ath+d/wUk1Fw
IAO+MPJnxwXqTIm+ctTS5C+Gxwj+IKyGglHEqJO/GaacjkRUNEm816+nSx1ENnUi
Ds6bq+UsWdLudWYzbj8oPreSMBUI6AhISkUUuod96c+3n1QTIabJsmkQ8XQ0Gac3
m+9j66kxoCTkRlXnku+Wgdhxy2vGGQk2bgG+xIebf4l1QYnaCrghJX0JSn6RGGzp
WAI5/HZ2Orkg/bY4lzroUVH5x2n3X5xptqb3Uz7I+X2CeX+Jd08Hly0rSgynBTm4
Os5iQy0IXVnsNUXqPzemW1ILPW5uUMym/QHXUu1Ie+WUEgWR8SvTYQRpWFzoe+GE
ImIdr4pbJM1MGEyyysmct+kQrdGxb8FEob79QMtBESjIGJ1J3QgpiUtOfit05F52
akfhvWjXi/AO5NLBGFB0SYwF/j9YQLy4JfJ+Ov9CWmHgPuD7Amz4hLo1lSphDJHQ
N3YcuLDffqQvsJsSZLuLIdc+TvzLhnJYhkO0R3OGSjmrl38dXkJh6NrJ3f1UG/C6
7Ho4zfFPwtiaWtS3BuOijkLrTWyyzTlx+qJlQmHOInCq4sXAC3U8k4Dw4j/o/WTL
CVPPTx7SHos3as72/4OdNy8hwy89l8Jzkre2xZoaHOthDZwiMA4iGpTcfyZCKB5V
+TgW2COVbEYnU4imSp637weK6brxIzHPJl9jRZgycQ2uP057S9Qgz312mwKljEAg
AgyI8THTdfyaQZrrCJvy0IoBeYmlpigv8ZpCprYOeK5zbkfcMba9gFxR84B1Mh9A
Fu802dYrDZ3ra5w7+Vj8uz7d6PsjWIPP+Da+LYYkAyJ/DeQc/di1Ki0yEcVn/xq6
lyh0QRW1G6Lsdc7SbonkJx4reyC+8j0XqwzE3noc1LeOjaCHQUqia/y8ij7WQcYt
VKMKiYoK0MlrYMA1SyVbuvs8T6Ss0hKaewfxQiL4h6yA/4d53b1yeJEWoygPWxwb
Sv2z1Oo8m4LFt3rphJL0UrBBmHuD8KUFb5xU/ckYp5lVcFgbGdzNYF1QBye7dgPw
hHCbBHCb2XCJ7GoIdH+aLyfej/4VPR0rxqluuI8uqGYV/ZNnv/O7A7AGx/wvd8Hi
WttotSnbuAjLWPxM71r8HpMXhBFYGHcQsyfRC4d7gwjh/Eqs4yoHk5OHH7RbNokv
C2E2BnRKd5TfE1sKOkSMnuUhEdy5A9ZFVmkjKN/f4YOo1V2ZVuNttzVha8K+DO4n
xje1iu6U5ZtRAL5jtq6nLe5uDUCAs5ak7S3AnnaQuT6YZkqTIZFJ79+l3TwuF7Ji
gLGKoOHTVZH2eOXnBYn2vW9YVhhPAnvgerh6BwaiVX9BdTkdm8q1U21jrafhaG/l
MvTnC0JjyA02Ly0Pu1Uwv64nu4UfrIw6iW4fBSDNZrDQVzMz/MmOR4kPgC+/ZVxj
3uZRs6V51aO+62VHFNiyHhwLVCoSYXZASWDs54FljjE/8A83llrjntx+99gA05nD
jYe3oJQwqXfQjeF9eY4Ke31nZ/N8ttpTqVS3Y3U4Lx+aXwBrs1CHtXOPr0FPuVv0
2K7GQPP5/bDy54Y9P6r+369QagoovCJuLYdDMbv/fJVN+eQ38ke7aLO5UHD8Tkss
V2QPvm85kQM8+z2U97I1+wLJt5PL1pE8U1wiNaSN8F2aaUruh23exU9YpppD9IhX
BcvMPRdC0pYFxhTiC9iNxsIdW5+IN8hNq5JV0djmnq0AZUAVBduSer8FJ5clq8Hn
NZW1mOUXRtA2vTYug+P5BB2ysnvf9KuyUzCRZc7bOJng/uVeUCLiJAcm8XE9hYtR
c2MxIQ4G6rUp8RfEhwi5JRDwF8Iv9oJak9fHnKraET7PP/6YVLhARdOPtUGw16xA
IRtAMAzcGRDqYjWloCQjIOaBuoSUrvHiMDxeWS15IOPL7qg0FOqqqH0NTrHYKKQS
7jEx4XKpACCTXF682oLZNtxcJRAbX1mVIb86mzDGBW5Bg7N9T9NApE+jT1hR1P0L
to+LKJMUavw/GqKnYt6cmQEvVvYlR+l4I2YaOKpKFWdscD51n3lImhgnXYJicpu/
lXiTqEQ5EFIoGF1G/nFpSuRo8r44QKAvvNxsa3U21JbRQA67t0TCA5HJ4KdoZo8F
2XF445lLStAZb4WajUKv7mmSveg6oVsZ1OHrtBjIhLu36Wkwsdadwf51cNZP8RX9
/Sw0cyx57BKATyiiaE4c73/gle0Tbz6Fx2cuDT6zXHa4/907JnQUYJLY8jrUH7bZ
NBYlR2Py8h5eo0SytV5mH8q+TNqN+gGYdUBJIZrBuWGMERoy3FPrfKfFZkCIwTgf
pV/+W57gNwHxrw4hYwd7DEgGSjodw2G9VSWzl7gZko8OJNOFMBAjlaMSko59c7fO
qqAZpWeJ75sFSJNf2Vqydj3oWusVA3hgugQZc5ZDxCLzjkmyVI4xNMvDCeI0aSaN
MK5cdW8Xx/vk0T+nGygxMJbPP5WtTeQNnt/AkGPCAImSVGOA18I6cXbWApbMRx8S
h7IiLQvNT7iNQPI1eqUZRHhcAQ6JpqkIPNmwhlDSU4RIgN5x/+eh/ltRg97nywCP
wIfbGgTTGvjojQ+NrLmcodDvbZHd7eJK+uHRcPCFd3YKzxl2wuO7izljPvmAIA9r
f/Ync2kdKRpVmfS/i0Zja5dQgIA+kL387obBABCJzHtOh/3RhoyiJWEwnIf6c+er
APF2dCh62zTkRhsdSJLQCsGcvi80wKVw8jeSt2hIRd0NvOUy48Ss6xnkvCQ//IXk
nCmViWvZ1i3HFyDyWmEQLul/boE1vIaENdo8CWFeXNp0v5jCalZWLjYkbVd2ogE9
YAL0BwmuTzbj1wWEwCBVqfFTmUo1p9/Ax0w5tUZ7dbraPj1XTgT3myZvu3L9twKX
2qnhmo6u6yfKkjcfwHsZMWMAyp0MZl94nZqr5WX0RG5/V2mmmWtmNqXNT8MDubDy
x9+4HkiSWvZO13W9BeLWIgh+aQqvcnwZd5NX8HJWKoT4A/6TwHNTnLDBENuLs2DR
O6VWwth6O1Zk4TWMzlqIuS0yy2ild+QMQmOsA15RV3MGkzmTSJg3FUA/qUeEK+Ia
OnHUJ2jhD0ssfqIy91pxvpHX2L0+hFbvaXPk7cksmlalHxS//J3lHvNNeK0TASN/
ffhSDEibj0dHo8ZJ0n1baI3fc08UHJimxBuvKhsUUTZjo172/abO1RNyP0B2yDcB
5kvzVXqp34ZUuXwC14w0p2+rElNT2o+vZhIQmPNjr5ZiOIw9GUAvjDtf2TEMlSj7
WCUF478pb/mtFt41wLe9f+MyFg/dSfVhKIlbcgEUQjk9iMIteEd937gQdqeTZPZl
rk7OIfs9Stgv/D4j2DUh6sz4grcVdRnhZ3udOpneGq7QJW1V9rNk5ez0VhC0Qjc/
K7CdANIax6sAqU1+VRh2T+TdXtk6cYiqY7YIpEKdNfTwsi+QddgALdBa+3Q4S5rq
1oCtMls7wqFENWqMYE7qj7XuhcogNd6PfCZcVM5zjBd5SaQ4N/G+HGFWIVG7B3SO
2eWx81KGFXY+qymVej7qvjjcLD1vRi2Q6V+zdhnRxUiw9VeXaEpzGKO1kS92FhfR
gXNKPyOaav+7B8SDshaVdDmb/QkRaLuhxJkERru88iessZ40nZbAs0XCo9OzBQcy
zIDx3PS1+Hp2P8BjdNX6X8ERPsm2cfxTfamnfiupBsk4mrH/o95Nw/t4n/saoCTH
t1+5cy433StjUtBwDvIST1p94FP1+3m3qxlC9DsO20+HHOwBqv1j0Nyh8m1uxBJo
QwUGcE5b+GEu6x+Mw7qrH+YP5Erjwqq2vQBM+tsJdesmj+URyBENf52Za+zn/Dkr
X2E4Vcgl2w3+UNPsyGoDwuHnLqwdNb7ZlOK0R0LAfNyzfT4osu/VUdWQqM0PmBxq
Yth3J7hI+nMPeIl4MmCtCAjpxdKZHQ+3E3Tx6AIjjlEzXG9Qli2l0TiQjzi+fiTF
6WIEUO82OJBsCdA6G5OtAcGDSZut1SCCcsHbXVOtXCgQIQ8wDyuhg6KpuQDVcM/I
GDcVpRealZ9cI9B1s31t2twa48XGXpfFnrB/dl8qGE2tO9j96miod2sSNKxJ0rqm
oXXbPEa0C8z90mn3AsoMCEaIVb7gO+/si+N9rKa4Hnp31C02odwrzLbIPyGEDsV8
3DgUtywli3Ei9GdilEsJllhLN/vAUddPUi/gyxcYYpJ3Mfv+KwGSOO5AgUqHzXHU
JxbxqWm91oXvRiXBOqg9ANqQCxZ8OXTSVippfdcqESUmt7v8H2Lm70knlG+su84l
dbnC+uGy4PJf94s3dIMukG4GmjlSEKa9SoYmaT/g490VAke8LltCsyfHQk7dYWLD
CJWMusJDiDsiQ5hU4WPM1xPFDompjVyWsE/6CaE0+qfvWgd2LoypxgYdROwwBI4r
WrtJF3AEGVwK8EmmL4CRtORyFOvhDaCXqceEu04PjQQBG9FeQLmUx1+F8LzS+8hH
GpPzsG2tH4vY+N+Gx+CCs6nU8zJw1jZYplqPFnRdVXzqlMDVpox/vfPM3jaxC9ic
cx/VE180R3reY9hhU0cHxyuug7Lh/fyjnXBVhhEogdRKkjRbTT+fNxKZ7XZ7NY6O
T2NXTdUN/W7SVSNwkTTp9AUSULgBm8f4FczlBIDgMmWgTRYNgccsqkMcHVeyM4PN
DeY0TP6X1CsZalmhtH5cvrzs3gCumspQf7zm3M8JFpJbYNqtfSgQwC9OdAIE2HsC
fdV69Zq0TDO8fa9YRYrnuCrmeLsJ4Lsrac614Jf2/jSafE22wd9abJSRNy0+Bh71
UqHTsRNOwqbXOXQgSUVaChP0zr1r2hXzo9oVD6g0soBEX0yuCx6TdENirT/t0fqb
ByTXaGr8lDO6OGtHnkEPGq+bpWfUIJYnEX8bc8CJQcOBn4ThHAPwBHNOrZByMCGR
jRut6bh+atalv0tdfS3Kcgec0JagjstvRMHFSVrAWLfSSI04nQhRDcs+QJee+pnK
+xtM6Pu5KDl4sGiMqojwnQgJZtltLeMnyff06ZLUmL62wv9wNGVBDeJ0Ahg/qU8U
jTvxv9s/bdteCBR7dnNoRtbrP16qabNrcttUhCdbONXW6QEdGfLwcAWI3i7W9y9A
pdNGwOjPH9FNm1SoVlCvbZc/4kqJE4XMHGHgOjMNEXfxWLGrv3QW8oQylqaQv5Tx
L5QBInkkggGeHG/eFKx7JiHW3HZbHjEhKacYVAjM0Z0S1+afdGYh+O7p67B6acUB
1JX1JJS+VNWGkujnTyjEZCEyqjAmdwOKTt1C9FVGGa3TgdDIyw4kCXhzg2zTRENs
u2S+uAVQOcQU2oyDLavtENa+NUDg+uqX9epgAFbCoeXnw++Kxs9xSaKGXFjWi2hm
fyliuj0qTvTxmZ9QYBJhQpfXS5gKSne2thor1hArHT0W1KLOMX/rgl+3C1qOSRei
kRGcA8Y1/3bOaXwcknFBMVTKJlqLMcMk56/lUpy0H63jwu5lRGjOiYkep2s0MyjH
Fduvq7Z2etEDidtINEjoS9kJXz8aymZi28AtiKysrE/udYz8nB2NdauKvkR0JFk6
TcJkkx15VMnp9Uh4AFkf5jY5C2TbbL+OEzGg0ZrsZsoOqYO/tTnZxPZb3itqoiCZ
2xqXUvYhHTkTEQ7mmoc0pjj1KsXV+vQDM0ljpBykdTegL75NP4M+wkeGAxOa5nbp
14VT/JYVt5YnHWOXTpVBF1X4Md8FrrSkeITpLFdssScXZZVCBUoDhhP+RqYEpXVe
a7XqDXeDDlk9RJBbfncVKd1rHoW5/wlZLdMoSeP6ZFM61/0TL1bMDRGOPxdYLD30
ZTc7ZO4V1A7LfiQFe2hItfeaX8ZTCe5NXA1Hfyc1rvwsA7uVsqe5ZSfZJ/slPEOJ
09tbg5KDAjg2KYkSMpMLXRcg5aSwFs1dekteO5FsEN15ZY3OQnsU6JQcKnBA7dgB
Gev5OjOxxcGg7Pn1cQ8oklSUfNpKGL5Y0dyiirJwBj7luT7nU0XHgeBj6dO/DDFw
+0jmMQQzHInGmrXTHC7hNrKrnaZ7hYSN9gIXZmVzjxWqlYCHnmhG6m+Cf4QHryF0
yUWXC3qvRJJjgF9wnYEcdYKrsyB/3JFybAjF3YeXHwq6J7o/nDWeieAuyp/uRZ/y
pNrd1RJneOPD/sQsenZJa8OzPVdYFVyOhMCHT3D3oXLl++JdvFkC+Ge4Qg1M6Gnr
BEXvvyL2tQbml3mZPIznhVXBaxuvnQ0rcWJ7SUdw/x9GBGKjao5C2xuhjlpXVsBT
rNe5CC6T94ZrhW+bW010zC0ejbRmPNqRjKEdWY7NkCL8uL9a2nmaXpgGC/tOdrDE
hjyr6knqJKZcAvY8kiHRwn4bm9Ibau5o/RmqOH+B6Vkdc/E8H6iaG2kmlJ1ZPlhi
E1sEx6wbl7ac3XZ38j8+gBl+GxVospx/sdoszN4YqADaf1t/BAsMGqpLZZuqc37U
PnpZRlZwAYVwPuVTvSZEmrdgU/NMkqiiOEnO50D6ZWNQOkboXHNVO9OyHrG8Eu45
9IYqkbB3vGAtJlrgDoBRPPJz+Nbzj8wcuDb85n75zeFRGWGm+NnULZAf2eEySXv0
qo360ZNw2g2AMFTVIKO1hOuuuxqXbzD89fFhYTxiowV7z0jEfNzTyIQ2+CwNYJO+
TGst1p9BUtdL9eIur9QD+qOjnrA5DMsX4mDn4knW1U+CeyhVHuq9KyKjQfI4Lve8
UTB/OTrWDSVkuTpk6ngg8K5Dfdpl5LLbtX7/HdmLMQNd4SmJGORGTCKS3UqXlRHo
CpmI/KjaiY5UM/Uaryy3EWOU912OPpS6kk9ww8mkCVv0rYWiFToXaVyQq+ko4gNo
C4u7AYqESM4DBiqSbL7C5mNpiCXn2OA77BmoWKLGOygadkMGImI9IRDVtb/3+01J
fO1EMBf3lvwrsHXfeD9sw09Sj1juQ+1wI/+vWtenR5BpDuMrv1J43SeI/tR18H4v
yXu8kEx5uzMRl0+Etht3igjNhjef+6sV99KSxiLo0lyUifn0WyLNvEf1Egofd5d4
7bhGc2YX/lqE2vLScn6REQv331683wGzZno3ImLAtd/tsVNDGTnfW0SYnSR6d7Jv
P/6py1kWTEpESiDkOTYo9t1O4gu3AaYrT+um41mdIMiof9mDWuiZt6GPlPQL/NVD
uAEyyTl6QeqcOquLLQp/QgIhdLfje4lSwQum78QIEPSvOPggrz6Nm3h31EiTiPEV
mWPx1qLryr4xjfCe6Chyt/fwJUQ52WkFpOBkEPMzaeKekC5Dwx6d1fLT8dmPq/lw
to80JD7HB5oBqVOFAh7f7yHXjo6+2A5s1HncFdsaLQ7MklGogeO27Hqv+iEFzOBr
bgVAFuQ5esUeeEi+M1rXInOmjLwtSG9qsV1TtimgVGFL4efeIPmwMAmBz0dv3TMx
nf8YWs2mSIHhixepmD5SAlSPQpFTSB7CnhVoCOvfs51CsFl1KM+XOdfdJRt6LV9G
7uCUxE/0TQI13Izi/pomgdESlV2hQmAd/6w9HGxZYzTY7/wgeUa2HBsMOzS4Rl8E
UnYMf3WdtzbsK+shjw1J44JwkceLF1RtU2F293oI9h28cOEyzlT3RXikZXp5Dz2f
qTVqfy82vC/RFy2CJadbewbhm4DShZXmdHdq97w+6PNQG9Aew9rUiAhGnGFsHY6l
IryIc4ErRUn00m5hVq9Z0bfE2sfeCbOXzpuakuSsrENXd13Ka1VbWbfC+C9TVfXA
joWup7eBkfVBA6W0yN90pDm1o/1oHvg1WqmnB5FYkKWQ14Gatxr5k8Yfd44RQtk6
EZfArMoBdTXZ3L+xW3ef3E1TI3eeX23ecgXC8STlyUGdzhGonza33Qu9wEMMaVDP
M0QWHNZYZxXmbsrXTu8WJpg8wEiI9Cn4LmhdUPx6qK42bbaDuIx+Hv5jdqRAg5a8
AnEvoZTiE0iWf5onlVjf3AhdB2OnJ5As4ctuWkIe6Cb7DtAIHHrpu8SibW5j0dD/
u9iY6XR9BLbk8TjT520WMaFweMVCU9fNPbmSrO3JTtfP0EqmEFjQTySDe4jSZPZl
/ck30EY5PLreTkfaoLnPrmzCvHHkjAk6bzf/WQ1/o7L6NIUkRJu8a9kfZfatbVs1
A2sZm1pHuWc0hksBaNLzmGtpiaB1DO+d6epZi8xnOzbEPX67K0+VqlpoRBO9Hs1z
pTlW3ty2HpL+uaxXkTBMU8O0DTVS9Q8h2SBg8zLr7arm0Q82puYx4w0VwRHBS34+
VICh+OPpAsxNuFDP/CVks22TZZ67akJdJyArcz3cOJuTl96AviVyfDae7l63eAyg
vVouKpemGk8GGfKqTjYvFDTHZ/mJdmEUlUBZjZFiOqsgOmNnmh66hgaKgmIqFVRG
TXUSV3BdyT2tLtYzWJ8ZOI5LOcClJv9qYRIb546vfePopWJVma6aWuMh7KZeYYIP
AjlAEEIbzVRygsObsrbTDjDivulsmdQagLPCici7/dZG8yzpkHLVQN3Nez1vIKJW
reTxCF2lvPBK2MBGG9n5pUUkldYDVP6g3LKngAEgsteV4gqriNvD4MiqVDFem3cP
0AA1b7tNEIVc1xcQMqkZlL2K4W91Y8PJxWu6wS/YFqtd2hr+b4Whb9DSwEKEUum6
CzcVEbqwN6uIJUQL3Ufs4wwOYOT3YGEV4D38rwE9aX+lpWpmlU2HO4lephECJQtK
cNZ1OnyYPAS8ZqsdWsnPrmUf2NhWbu+DQaP9s0IsPvdT5rkjfXWF13/wB+ZyMeO0
FmA/BgrndT7UrLCEaK2qho2O8hFblkRK9kv0B0E5Tm1r1Bz/4ff4fN2TZ8d1MuHi
0Mc4djv19dIE7Gbd8UJOWIFOYAVOQWgrLxGhSW7KfcneWVz/1W2VPzNVoLddlN4Z
sBMpKvAQjIaUjjBo5ZvUVH595gni61Na4PXhTjaXd6cRXnFX6caQZcd76Z6GBn0a
E2/ks4zD/uiqIlviwhVpc08VmdXgW5rR2mtFW806QABajldCHTACo2uEugQ+Q8Wd
qV0lMrg7+J/RXi8ty+fX8sMFfZu7mlXs5fOLeCyDItAzoQ6BkWO3AjZpH58pNfhi
KHJVf3x3qP8zn1JOZk8k6aARXmtShqY9HJwp/uIWB02sZpeCY/c0PCW5O5ia9Hdj
FNcXcHrFA1mThHszcE8T1xkkcjP8Kue1utEFnDsMs/Af4RTNrPpFi5pFqXC+36W4
kjO0/mENB8CLKTfWeFaxgpufaXVux6YzNCoUZFk/6p90UQNbcjdwyNZjbA4NcRBG
wU82uJijbFQ8C2S3EX+qhHZKV3yMBkur22oGzRXVzucCdZbb95uRPTWKBLK9h3zg
52mc/MfPES8iF/3uiRUFbL0ifmmC6LhOWk7dHCFc9V8907VDDQDsCCLYNee3V5SM
r8usyOWAx8Q24d2dW5UNN1s1ld2TN1/LjQ8dNHLAdvdzNo/x8AX1M3WImMKi0NUx
MztH+67Ob1AOq9/mmllYvQ0u2QmDxcWLJJNWDIKiZ+qtRD528De4zXUnz/bP3odv
by7GCesqF4l7rA4v/l8H+xWKrAKsSPYljWjDl/fVHCQXJGrDUFRNQCzuSWs569Jk
edw+PgeeFoalDzbS+IM2e2VwkdfFtBymsOhZeEqawH5ztXxC75e6jcojOQwWx+IU
lFb1diCghCBGpEMICQoQNHqwamDkZQvyr78QXzIRMueYJyzsQYDXA+Eo4cr3+Efk
U1oJQw0SsrwPXG64WX+CNcrwNlLkXGC8O6+RNdkDGsCyITlqhHVqwjA9yTZEvCee
6laG66BxQM2O98bfGpCjwhzxrNJHFuB6nraFVOadIK/3ssUS7UWry8cUfYknkpoP
KstUA8kv/qKM3S99UkyRDaMw2UyeInftq3SzCGi3yWVv927ZZEyxmpDuKEs5tEJG
/c21m2Y9o6S2eHemlUoindimB0cqeQ0ijecRzrlyC6XG7vgFoFUToLQQmBcaFswp
csOvDIoMLf/DHkeu6inGJmmwjA3bunLSkMpSLxG+FjLfiBgE3ZXI8Od1P3q36VTv
FIPMBPFGq2T1Pdm6r6dPf9ffyqSe8JDU0iFInwSh9QH2izyxfDOEde7DqA3Nvz6f
/XKpS6iVK+ilMlXi3vZ01yQcXTC4y/q+OsJmcx7M7ocHG22MXZHEb20LWac8SYl/
34ozrUNLv7BIGaWHIDOeX1zyxP3WlT+nq4NAcXG7GNqXB6JvIHPFU2+civ+4It3j
qiZ1jPz0SmkKLIgsnGsniSGAKLRgA7m591bMJRccK4u+wO2OLR0nMRf7axL+EZJr
aaulPLo7xt845B00DLWVbZTY440tekVhujRQMXdUBGwtTGPWi1dj+Vtkuf33CYTB
bkHkkUH4/dV6kZfbKrF7R4KqOxsOqSHHW/C2ZFCsCBSLT1SPrWntU2WAYoLRnXa1
IFyFj268xRrRMJKkG/SvtdQMSBbnaNE5/L1ieXFhZR9oiTBImJoWN+krwKZSZMay
rLefdwZqLt4F9g8uyUuMpT5UwPU6W5XY4Z9Imd29cGyQbCQdI318cDbN/qAOyyfy
0C0JD+ZW+U/PVZv3D8fGPlWkVVV4Vxn31UqdyeM78a8pB9V0SH79TLuyJ2wap6aD
+kCK6r+4qxo9ode+n/ejtyXEwCrH395KRKip9hJod6obQxqO0UBTcVTat93kF03d
e6pKvyfyn7NCI9DYeHGqRevSXkgOrOsURWQhWLkXXZ/SRrh9ZLpBB9gkWGVfet4B
I1aFmqJy8r+IAVj90EwlZ6lC4fTkAth5uK9g8i382BXJCdFpce8nuKA94XXzHs9g
+g+EmdPheu3ZNDIvKR+qEnu7bONeJTyn5aNh4bqB2VXhmWeixXAFuMhwxVqdKvY1
KesTo7HoCUJp/TnNQrNHxKWQ8U/3K/PtZqePCj8U8YEiOGBeproZp4LlwlOjUycn
2A5bmFcNTOWNdxkyBikWPZN+sp6RQU/5pdZiwI1hZtjKDcHoH5CVphx2hQSR/hjs
069eKxBIDNf62ofHJb8wB0RJOEfPeP22d+evsI1/fUDnRsurPceEqRp3Ni4lVJGE
ftiblrCdB4U7FfRyk5cIt4riXRM+gGFtJHKjhVIXM+uFUQD61oNFk+HuPrASzfAn
9SOKscptjpwzsWPrEmGIEvvrt1wZubY7BFb1jrJW6C5ZvUsm1DJyTwlZDKqKGKzX
xXQsi1kh3hSRK0E/tUcHIg9MJsmKUpG4eSZE7tSlb3v4qt8/jZlONy2uJiXb8bHX
GGmyOQpdwQlgaUsKEWIj+/QQCCkLBiD9p+KBNVVpyoRaUDkahFO4p37pb1590jgB
IDZ7rlhiYxiktaqRPMrqtZIPqEkJVF25F6hAgZxrSgllCmekBBI4WzbQXEy9LdUt
LH+tqLyLffzStBfqDG14NbxEli5TyVWOk8guxSZJn3wRLFzYe6m/ptRpiFeoRY6B
nArNmsoljSSumF77aVbLP6neLc1GbWHuzddEwUXgfJRZf7YvdpEDRkK+N6kqbgCG
xfHdXyQUnHEzmcuolQWQ0GCy91Dt3vUEDRWIZ0CtSMzMQFW1LPPOeRrFLt0QkMV3
noNJI4H/GYg1d0R+1luXMO0O/AfycdHUueayBSsBuSq/d2FsmMVOyDpGrY/Huck3
epVrvrO9LeAffKCP5sUeSOwCkbFMNbGEuqcNekAHEY1ma5F9zH5P5zClbuH+tzUE
f90827eLWKqQ1vUPhbBIhMrx0ijCXzSz1rc7NbMDqVioRgLVroMgGSY/Tq+cOW0S
y9s6+9PtZrb4C2wlj+W5QIA5qK3ySk6W+DfwIWPUNI+/YjOuT/xqTxMtR9oxK1uy
vux2O5Rf+nwSEmY1D+vVY41UUxB7fYMzm6ZfosNVliS3vi5YGRngToLauYKl7KFX
d8Bc+WCD/QAee+6Z2oOXl49acrQIWX6mmCphxiN4k56SLaXz0Br2S7Zn4hg6jYwI
3ZkMIh+m6TPSL9ro/N9sFUwTqZKAHruHrMlUzhvpF76gg8XQfZffoV6nvysAEmHx
X+V8hY93CEKAxjLkezb1h3u+yU9oME/2DkIDrKsD8i+09oZrCi83haLRQEsFtLd4
7lX1vLFXwltCZW1TwJSk9cQAOElKmzYEe4s2Fdl82cCnWxYL5mClZIcV/EhnKQ4j
ykvMOTiejZI7nr/5B47l+8TwiOt2F1MjQ2smJNwEfDCLJIlfwNz58mYSO5Wi5imp
u4QKCl8+1O22gFCMxrRCuy4w9a1m5A3m87BLUZYVYGLU2n+PFMR+6VK5IYYxeMxp
ho0VQUpGrfStwwUK/gMCyq5EpNkSwavoGsBiSdco0FXHg+F/tMHJkLB8X1zkx534
rOjA4FQPgBkhBCgTV6QXqV8AjpyybiRUY10NavcD6EGoO22PG6DS4V0INyIvuX4A
dCvCiOSH9wlA/NUASQwcAytq3fzxBXX1BddFGf5bkKaPEcFStjs+brVgBMTbK5O7
yRJEeFCGnCImxsjpP45xqXqGuCwFMRtj6uvjwo/RF7kXr+m1+OkmMMOx6faAeY6N
X7YpDwcgttD6Rm4f3TXNBtdEueRtV6ZSQ8vJnYuAEvoilbPTOg6EWzn1MijAt2fM
wl+XL7yvjRKq0e9pKF1+rBzqIoy5Xcwz5fgnMca0YflZFBXX9zgw5w9tPbJ/7yWD
yK0ZtTSqlV+SFj/V0T79qc2oaw2d7cR9NSvQPNypfZBvATIZzLGVyjKrbCls1hR7
g2xikHhTgNWOROBzIU2Lz1FNiRLUWsGX9KvGgkypgUmG72FdbTAleQvhZPwXp7ra
5gNfonXvUVSSisI88Ca2fcpG7GplUhxaBzyoJUPmWeqUI3jAwpJFIP1DtxkSUJO4
M1GZFMyWRhTrB6T3mkjcpUzAIgDIOadl31oUyrfXAJtr+M5j3s8apkQFaT/WMDw/
+a2klpiznzA59UjrH0RCmyXCVrLInDfbTELI+JLtqTPeeFUuMPQVfPLRrVgbyKwm
RVsrV6IdiHcgd1i6BDsoip9hZAmvYHVsC0tl6ac0PVVtTtqKav68Z08+h+5RNnWn
tqayIldMg2Q7Rc7wuT16Pzt8FNwScg3+Q8PjFIdTI2dJ07Mt/HbPSHLwpdz/wT+t
SSdk5FjB9BBMLwp16UB0Lh870y6OlXwMrsNTIDC4IbcOkNJM81iIjIr7XjbTVy/f
nAP8LE/a2QZQoNjn1Xam+wZb8lyz6wad7K2tkc19y5W3dsi7GiJCVNuBw3w69dMQ
7amY8IoFacLiPULcHWIB2Lq5tZ8N8miPBiUNcza4OKoyM+uNEW9blAc6GliTlCZP
95NCgD2Um6rlh+z+amDkM0/fNrswbUw5cUtINaGSErSx06UuBVvVt480kFwIadaj
B8ywMng6x80UgXUU9Iii+wepQG31mH4H+jYYPQ3FWlkRHVCnZeo/kpYzQjz3Cpcc
zu4Z5YiWK5ylvyWS9EX8GQpg9/st90QH8uLKDHO6efS5S3pQXXXLRmTaw1HuyMZW
a1Q+gLpShjOGSLb6yQYanv3/eveKjZJiYdZcR22pnAm21DZpgZLczQaOPC/aKX0I
/J32CkMUKv+Ci3VnOhIAPPe4wC1nMDM5Zw3T2WneoQkOOs36EofUl+HQmOs8j51N
Od9EC3FrzZxQGWZGw2NOAy0ctWFiToFt3LJnP24xeLdp9QQpa327AKMETN502m0y
hDV9rR4ZRVgeA6Me0P8G0pO1dG3oFLVQiTKX93q3108bPym0zHxoFsna/BbsFEnI
J6EAeTWocEhwUOg35qOXm4Q1AMUUsZl54sZlF8z6UfdVk9wpxPUA4UscuslLTN8k
hMYbzl7cg89TvlUPC+vj5VO63JTA1pvkgo2BC8ic+5T/GnQ/t/atgIBqJOPaFyKB
t1LNZCSkIB01VvqU2YJ6L4SFOp/AkRkTDTJ3bMb7SQ/9T37gQ8N6ZuhbChLeEw9B
VqnefuCDZRdRRVGSuZyGfAcY56VAudbWmdIXLQgMIMMMcIPflrrteQS3cnL6m3Hm
XO8KZBitJ/KOp4IKO0Xl1d04WpAEwn/9xeUpRCTUkcQua3IXJxa0p3x0JA54vXOg
pxuiBbATkP/BACz7g2lFcHaO/3W7RgW3AxiCoYGkPl4LheOI5pCvN7w8RhrBm3A3
ppbszh425eOV1sU1WtPzKjdNma8eeczP4M5txbv3IVGuZrZF62N2OCbD5wHR7VIi
76GYxdMmpxp0nXv2tYrCSDF/Tol9NNk4jc2jBkY2pD5qcCFc67e4/gOcQblt6TjL
Qbn4Qjx3lyMlqYV+wmQKfDqoonTNiQvSVavqXCHIQzuTqHNZQ+7FvwIS3sC4CjNa
O/xk8C8l2SgKmorhm5DE5ZCGajqr7sAJTuLIxnNUVqGE9digOE3+A3JKPbQCIm48
43aoNzM8TZ48uZGL3TtYaWjdGs2uRArUMq+4eW7f2X7sN+OVj+TA6hOb+lD8G+DK
GddLIS+wZXzZnjYRBOy56f0x9EyN9f8+nFF/HMKSJrtWNHIQ7vRAlBvL+FcaW7M0
5uz3YU5emTGfNDm4m5aHkRfonnq/XVif2W9UyfHJsu6byF0s4yAu1lM7k3edUyH7
GNMdWV4T+0G42GtrM73eMzVvfnao2zQfkWAKmkspSqX4/1YuyEb5lRFYsvnIl3hq
4n+yNgXYZj0Iz4tFcJFu3UC+SpfK1Ia6b6y3BsJLcZw63Wg7Os3q4C7BV53eajbk
piLb9Xv9lqFIIC7S/jDb8/Z+82SBh+D6uBX1hGyWPziUGct1/zgQ9BlBbvvgqDCI
Xy5hBlTuZFsK4NASkn99eyWjnxJZjxbjcCVeaKE97NzasfqcSQAM26T+xOGid4o5
mIq3Oab59teCFt/Iwub2r10KEx4plWaMrCyEDkw1kL3E9t1subEGX01fqGJwlXdy
ACC+9le/AqjwUaPBcVxVSJE/4g+wnSAbgCaZD1bz860abWz4IHJeLmjet/58RghT
B4Mi/sTFZpzlGxqBlHFGBzZfXY6aEMHmyq16gFwvpGcSRIPp0vDK79XIsuW+uxHy
EUFOGUyi8zlPJ6uonxnY6QXY6BL9aKGTLW/A6gxGl+7TiTxplfAG3lkLCFBfnUhQ
kc/nwHG3bFuwv3UhYG1qOx4zn4lOUkpmO4sSe2R0EgBaT8wVUYIl7yA9t2qevqXQ
XQCD6eE2EvNUaRKIRjJtZeavulJ/b49WZKNoNUNmsF0lgn9HeiD9jyF1WHbSmUfp
OS8n2voi1w3oXrtWAelB+jwZRIZgovPTWT6K6EydQ1Lpr4K/aUCgOrVW7/dKeL5I
LHQbVFEqqPVpuM9bch3GwQ0IMhc0vtFy6pSb2nf1I5mgJyVjwhWyJe5YXtR/PdbW
9P5DWSHD5MXHJUmGPuh63Njaptx2C/O0Ff7ZfgsOMVlc3o7xasGMplckRvY6GzQb
3oM+3CHR/gjXuZgA26JHaT5Tk9R+kPJHKIYdAnkj5AjveBPvPQqqR4FHsjY9lvGQ
RrswFZLCnpizPDr/2CBiYHYYS+x5nlTsrNKGYP9cTg/rBlet2pA8TbuOHhk37Sx0
2SJ6Inpy/FQkH0kKjGcSgUaBVi8YTIiMBUsbU14WTWiheLxnicOIIVRgYAEyAht4
IT6bYAbJWuxkaD4agL0lNyv8dPAtMYJ1rV4WmevXKMhx8GdkEBGjvjPEmQNaFnp7
lgORbA5LDSPU5kN6laPT+BdcPb9uiOT3hQPiOiKC+RRRr3A8eioIMkwl75ta0JPP
zZrPFHX1OWg5/d2NzFB22TRr0xKuRm77NFTiacCjXfir1Wzds9KSvt3FanniksIi
DdNooojQr8TVXxWc1V3Ra2Hg8DrG2/MgyEBZ6aPddLVUJ4slapGyYg2vIK0b9rs/
LxyEi2lTHsyAj5zh8voWC9UIQCe6AEvldU82eKnMwCdrltJROXBIo/RhfLFl3UTL
7x4GWQKqHOmHnYQcTcVTt4T9V/jAEqKHOJDDsDrUZbcKbyPNevFfOGI/BQwNLzBR
/P0srIHLAiEBAJvHzELDMXjF5hFrSoTUZbJ+cuc666MqeZ02luwEGCrKl3D+SLO5
/2u31ajXV/6se9IA5+u1ch4wEdGiVEx3JiWOY1c4oCFjCtnaOEhjuvPRts0Ax5nD
xSgI2T70f/Aa2NisorFVLDeRGnioplXYrCTBP3CjrUEpTJrBVcTxQo/JZ3QJgPnH
7LhDveYF24Y5KGmO7C9r8aui2Zvo+MVPMTw9KL02iwmo7dew9oX9bzJIhoUzX8bP
nJmYU8c/kueqUkSW3Tvt2XhSuMbJYTzyAfH7enk0JUaizeQYP6hx3jj2U/d6Wvg8
c+AE6a244rT4uHJ0DSCs1f6ijRVN2djD7zBfoNlOe84S1bCM516WbywmGrSKmCUn
NlUXo8gmqE3TD7y2yD2zEFNuvlfYMaOBWuw9KcyrwdrM7WI/14HBzRRHtzP7WZUE
qP9CQR1NaShVWEHecg1AKEUHC4ik13p/bT2nEnbtvLl4FVGfSDjaGV6j/QDU83/S
jFi6/A1mabsib4Sx+ufhPaEVQNVjJtOt/Q2Odibrne/W1rG2FKnS/WUOEwG02Bsb
+64p8GEX0okBcjLz2ePSmwUJ6+JtkUeXp1+SZs80ehIjoiNlwQ8uFWTtItjHlewC
5dk9e/V6mhlvE4q6qnEomXbIWIofDiSBM0pRchAy3+LgfGTs3dW75tMlGqvc5/3Z
30KZHPZ93FhLnRETZSyXjWHWVIShly7viP5w+HEVTlt7Y2wXMLIgNZWfgdnGyIib
wm/BdrTe5qa8Pl2QsKCh/MJHuRfa4sIreeonRYCkUJcQHgq/OpubNXSBBx1QkQVI
PWaHoOpG7jwzt38CZW/+RPt+eorqiW4io150JaC/X/euAw9Irvn59tinbk6qrKef
sPESzWhOTcZuPgA22F6VhBKkdsZ2WMRZOGk51UBYYOFTOXTKfebKpAcZt9GCSnEM
+yXFOlaG391V+ULI24JE3/IRbPZK8El3yGnJPlR67rXQlNke84pCCeguymszYMF/
YbtGpy4VYwlCyzHDQ/4EDqQ+XvI8Y+JEHNFkL8aE1WjtmhRPyeKMKK2ghykHnWl+
8mBK4DHjttKyQuAKCmGT4+rammWh+R+OUh7peujtcMgNuSRo5LIubkspgMeaWsyR
Amxg9tUcM5vCnn8gHeT0B3a7ZJH6vzAIIQ3S9q34UTXVexd77j8ttbRraCBnfYIL
UaY2ulAsOQXok7LmL9sFLnHX181ECvr5rDsuppmihV0CjIFzd38Vi6diTelvDr4r
gkJHwBHpiakJj+R2/CXSETc1VJvDHmcuVyX5xtqZSG0RcpSIe1/1JZ3LO49cp7E5
GtmkhhiERObXlz5BjVlKKOiaSMXOHLOXC1hGIvxeYHfW2cHEMZygX40iQ40+FfFO
HYLGTqhw8/t7SFyy+I6Fz7TsZZXW4J/E1HHkquuIBO8cjl/4D+3mmiTbMnty9DUR
4crbLn7KB08ZwXfX8pY3eMJ2yYKmdbM8o3+CdeaYJcW7vC8jPOiQ1cuNf6t9tcAz
y62fqkt0ZDIsLVxsVHEPomDp27NC4MDZlGPjJH8ZXayQU64GTmgVyQoaHIVxpGw2
HChyazEMeJb32WipB9w6yzWsFubMfPk/wZOVFpS3y7NS4Fl/xoke1tMkuOzbvAvU
q8TwXa/lHOaqTIghKqtCGZh0XNHcspGzdG4ofulSlkJTaAyZdXMdhEQJzbzeCjDH
nvrkxaQBuO2xsJkd/OuxcHQo7wHZ3dp1VgkBX5YXqPe/ikD8yfKGyqVghMXWeOhV
7FfcYO3RI3EUwhD5O9SwgWihMqWHW9LBKra5ZTNNFhPQ5XXHvNlATzj2l/wuW8WC
gPzKBtGxa1XtI9vXh/FmGFxQn2yZfYXvYh6M9LqEibcLba16lILdkLQlbid9Q30p
qUuAzZ7zmhYdiyUzmg2zDWpzS1uAK0jZGD8H7G9zOCJORxFU2KiVzuzdwqnZe+QU
2MYmEqsqFldK56ONhz0OyM4TBckMnME6c1zKfplBLGsal+9YOKdCNzCtyE1e7uvz
fpp8B08TQTZALslVsw9Wbgvm1+BZgSTdrZbBZZHUx3mxVMi4gZW6hwxUT1m2EXDJ
7rccQV2aZCyZVvBpm7ovMmWerFLQKX8fdobFvLy2hvI3legfSAVuxiVpHhSQEdSS
jLBLfkxLSDOHbQKC0yO6qqfLGM/SskjmukLmKKjHNfzaVp+7UNIq4wYl3U2HzCqm
hOx/fZ3X49sD9zqFo6YBoIunwJVBPL7HRhDvu6CJ+MtS8FY2hkHm4GSULWOAp2WJ
vYFTNstfA8AQffg3E4+Gfs0kEvz8nYh1OBSH2o7z3q+yHdIrhRVprJrkf7zhFZQ7
OzfKKbbrCsSp/6blQBDxSdgIQdZ2Ge4j7VXBVnDeJtEpmxxrMdfERpEEm5bdRwyh
grK7IitPxFpINfmfksbbJHOg/L5DKnQOhC9js2KvehGXScIN9mp56EvjAKqlVKav
g+JZ6hBtZS+mO8rXZ/CLzlbiwX6s/KD9pRkjYA1pF06BLxnBAdY15EL05zcMhB/W
IL7zVq3kxoD6dKBv81Ep0Low6S2gZisRr+X/CxKsSSQUrYb8DgkYv4JSKn0TdURF
OHZ01+CsGdU1nUPzEiRDvSZj8sKx7/gJKsSd7hvosM7uiz4rON4bl+wnQe0flEtm
j2F/otk/N0ZlbckoXZCiwxm6stQdUyzfd9SMj0J/TGGqUC36vO2mOJubX6vPOAzX
eqeY2yMfkhvwfHZ+Iu/gAnP2e9+8KimTQdYqWc+4kOBaUrkHa1oZIdiX2FWy6yzy
PE1bSh0IReAFDs+TX3kF7RRyQfRwLnTO2BO5nz5sbcDImhl1nVu2zD+whY8GaAno
6/SS92kMHCRqwYElJMVNKXmA7OAK93ezr1/9RW4rlqAk/E+adV7GYo/+FCrmj958
kfLK2P51GvklVO5J4O5RnbBv9PNil/0KjpIllYgp9KQii0r26tFNJA51oR3e2w4U
dKlNj0xMSLm1xp/FLzLdwggkV1kkPR057ILxmP4i/7Qju1Jxr3zTih9da2i+wscW
sddmZd84b2QWwAbhUwFaQ0zhFvlubf4kgAhtVMQdvRdnSvcRkoUk7FbGw2PhcHp/
uUcxegSwzpmRdn9MsTxGjGGr7YC5G3A5kBy9NbJG6r/94xkOrlM+Muc/V8IkdEs2
gjkgrOY2uBEqst7KaAnVf+R6OQWi8e5IIJ8PQF2Nr11UjBjekIn4PpBNx/3h8y8G
AOEecduj6ukZXL2tuNeafbrf2+qMX/oQqBLHdUpr24LpYd1xDfxWn1bqjI6qOt2+
iBIZ3AyvjJ6/WDEkkGaUYNaBZhSOm9qH2JtM1o4TWr8R9iKlYtIFYABzz77rSNRX
IDlng6Ud2Apdw5OhDV+y+zVvCKAoeZwuWAxmLiJ+PhcW0m9/3Hli30dStLnTQm3c
ROKYvgU6x11h5RGYqNo4Q8igFOxJXJ6EMnqkeDUz9+H2uWLoRFC9bHvCUVIBHFiS
YH7u5cUxCjDP02O/r+ohl4lF7mu/U6wPRkhXDW6JsJHbGn52Bs7CUL0VX8b5rQMR
PioA2C9P8N1xFSCijN1CLhiZ7cNUIQvMTuf+lq6kAHdMhczfZA7cTaJOWE48u7xH
tpcV/rI0W/lhFTRpUUOvFmb4j7g3UaLr7mQ4o1nstRokxCPjnHCL5VrVl1SpRqpF
vLKdxptxuYfdba0FUITVdkZeKSh5uiLk+N2iHq/y4YlTANOkjlFp/9X8jkZ4wEzk
GCWCGYmbAsBs7ltjRPS0nQluqvSai4bl/H/e+ZD5M5BXXCEzRqqRIPiCru3wJVp/
M14WKHjfnN92rbZ+jNtXRRm6eL2c4p+tZi9LyTrzq4I38qjLMHedaUGAgzIC1VQr
SCY2WjiLBdnwJOHTLTSgY7ig/2NUKsbExM4Cs4Bcne3EEXBTamFo/1WyxTiA2otw
7nC5IyirKJ5OPj0l1FJmeyFenkQKylySQySaxChSTt7MALJMJgJieg6SzmSc5buC
CAv/VOG5HBrq7/Z2KYFHoIFMrnfA9ikcYRfpYTynfd/Zz9wYNF4rFNZW0kHDcvl4
jCVhxxIRZ7YGHmI1psT46owR8euxl6ewnCDjQB24GlbH8HUE6IMosrRJDf22mU/2
qHFjWAV9BS9mJ3OLUeg2/95DZoJJ4O9Oq2EyoaT4oRnfzk7006cQLL+S9k+hQ4Nc
Fyrks0C0p0cx7nXjDD64+Zb0vcthvRBnYcfwcyGRVAVYUtaMlmeaJjvzCIZmNwAn
blCCYj8U/2g72gx699LdNn5ITrASbhhV4YmpzCHm4Z8buIp2mUpzV55w43xfMCvw
MuWh5y5qky4kKjWjAK+4wWHpV+WsM5cDWTxUKYM+QkwPJmWtRNihE3HVgwdQocQ+
YNrJtLZjse/Mx/arRyCdSLqLwvASVD3iitasMeTW7dQVfm4H0X+y2FG4biu7GQmN
klsXUrTdWWDvEro++iMUAAbbYSEJKLxy+uYhfV6JD9KesmnY9YKxmRZFAfgZbNZK
s7KH6FJDVn43xp5HRSnypKTxYiRJ8FC9+taZD+8/FgU4z6uiWSChZLQgKLWiCMll
5q8F8lTZRR4eDqL8X1/sjwY8IjcpAEUAJ59Us5zm+xMwEPg11JC0A85fnwuSxtxH
zlt1DK+GztPBN2jTaKoz5dItoVGQXYl0lat3BSXabpfZYa3yVXkBu60AcxA3dJFm
xDCAWMtW9WObTIJRvKoYufPwzNCDk74xrPqhStxSZs9w48w9ErNxBWBxJPk8hEy3
gxAFP/uovnIrY34ImzlMn1naLSTkfZYQ8GFIJyQ8b6EB5rTaev9aURuOd3jks07l
BLYEeLSDl6+kYmlgbh1QssdqNA7kct4R8+6nM4Do5ZMkBkP7p4FOjlki3fie6haS
rBCWvjOIHuOsQpwn3o3TG/PHTRTLbnCxXlGZMcy0f8eyGZ1SyBWHtwP1Q9VOn8G8
fYz5smxOHpXqen2vkcLFx5Ua8wnm9MTDLPW3cF+J6DOH2mVciS/pmJXxiaScf5oh
7s4BOHNuaUShYHxRkPkYpXLPqv+DBkMMV4pxakARZxiY79GGOE4idyGhSKji+LhD
S6LKTw7Zq+bDEXZTKlTqNrZZOh/JEV1bsgYUxAoLFmNhnrtJGFEHBA39g3MDQFlY
KTnIEvHSiyam1H9kogaecVrmI480N6M6qucHtJT/YTaRRU8+p23AV05QyXqWw+I7
ABM9ZPO7JGn3BxQ6qij7CXvec6Q45ZN2GHukJPVt+W9pKS/uGLiPkfY6uLuIgzFU
WWFU+ydcaNt0yFGnQkpr4WGoMIwl+p2rurBPDtK1jysJuXeOlUdhEPsGQA78jus8
ymZ1L9mi7td4TrKmzRCeLoFAbcJc6PPmWFkWt4yMbfT56v8eMbI2GnHBh/zl6tSu
hrrA9B+gOiSqpGkHMImoWVVnNPmHlMtmQc8BOJm6c9cL5YZMGscxA6t4vrKV4AMo
FJ+opem3mfIhylhCHuhrl8LM6P3BqPbbdQLjrtjtZa268AznUGNHRWsoUHcbHYHz
PsKa8VeP54SWRrbznUxsYxTLatBEbaZbnOIO3DHV7OUEP4qbwpTYeH2+WjdeVHp6
xAMGTxDskgwPc8NabMNRqWj+krqYRvvoWbcbbYsYYgHUUc1oK8piC2aXqXpSnBAI
38rrOYhaUf5lZYFnsORleTAlomApzU9l3dogw9x9RFgp1l2c895rQ6yWJHZw1tGq
7E2jmFD00Swx/TVgBzT+YrCLSfxk1EfB86TeKYuOcYScucu3jjwpqkfiOuefD3w7
wEMs2gV7CAwbv+dUvIEl7LK9MJgFKWqk+vIX48fopEdEVyRnLQYDRZHmdjzLWeiH
YKRByFA2aQp8bnt885I21kHbETjLPpZXhXoVsvFoR/tdDa6c2sw2NhD4bSJVH0SC
oheyZqd2zWu9mCcygTMk9wZckvZe3vIEGqULep1IHz5HMQiQJzo7ht2Bk4zFsRlP
0bfoEiMWBKvKWkg+rgBVwXKAJaHosbCB6HO/rXr6BkEnJyqQa0EXWk232Botah/D
3gcYSRx5CH+z5QGjNYFvuCUTa4syZBo4SxOQbO2O+r1mayjF6cn/+TOk3qxwMxiL
jHvU4kiuwfDV3LT4ursW26+IB0tcDiVO82cQ3WgtNnpzr7vjNRFYLQxLs6Tgj8+g
WHn2OSEFlkqFQ2g1YGJW+0aYcvNtHrUpieXRPZb9Di67OhLHCf7FMpkyJAtt6doi
SL72mz96JxZGarM6ICoYASbALSv2SqSYmzKyzQ9GouLL7djyvOdQFmYLunIYBP5H
KfJIuiFMMLDB9Yi6G9H897yrx7SQigk/owLFd8MIOlfK7tZH+8Nrl528xmBA462S
YpKByYObmdDBmYME/rubYtzD988l73kS03/F7FAJpSd3mgU3Elqet29GmDeKeeGg
NgKFJLytUtwSEeezyBNBJ7kwXrzPOBgoPuPawXO21VYUi9z9XyFELy6p8t3hsV92
5u5Rjbw29rqX/VEEEe/uE15P827p1nERm76isgOSsbgiC9b1w/i/FVlVROZIttfZ
VRKZeTeqwfBnAHQH6bAlAfr+qFFltzxBO/4pCxDiE9QnFVt77WrxQlQmlT/kgsLN
9nheXED0hLXzvMM+BnuGjC9Bw4nDdQM0YST49MqieLNA6sFlq7EU7F2lxnJq9o+U
HoejFkCit4ajx9RKmhVudyg83gxTcRUTFIycdovqn83pdaOtYnrlwNmMF5pW+BQY
iqRbxiwJ5g5dSsLOLyF1hos309PtY7f55Aa23ijtcHhGpZ/z8Iht7O7w+7YLtK4Z
fElxiv3CZL8nZkRl7t2ZIqdPFYZL9RqCq7YZK9nM592EoDKZ6ASrZurXPQuQNmy3
Gvlroxt3qIuvnGktCJpImLMQCYO88IXOzsPwqFHaHAWCYpZrjvqkfj1EbqDg1XzZ
Eg0NJ5lPOoroNsDAeygdVS6G4eTFsQf5uXOUfQ2sDE0aFXcZ4aBYzjaccJN3hKc5
qw8WV1oEeX6DDqz4DsD90bdaH7oOm0uz99Q+6kjwOcyvGop8RIp93TwtzqI09PVX
7xUa4ZYqGHafIvSe22oZ3oBEEfHIxd32GN+XKD9otvl/gu2zEcOOP6ke70JOLuLb
hqReMrjwBlgp1Sv2fa/2YU4EY7ztBk5Lp/gro/odtHrwoHGisJy82wt4QqyZqh5w
bUIulXMzieoX4Uh9zpH4AYE0WSArMACYT8DoCeoVlqSuk0If0KtGhcioqO2F1cIf
fABmdXeJUItUeps3a1ULSHyEafUBSwAKTqpcIANCt+3nPD+mn+mLTZtpQsAUSFgN
evKvRqpltvD2hAN+wYt+Lemc8jFbQJjtyxJZp6Ir3FI6znEwulEzDeCftaLpHRR2
plRwFidSQ581rS/dv5sLYS0Qh1FgGG69PZw2Pde7Ja6Cxb/Yo0Yupm5lj+en9Jqi
Y1gWCAbdEEgfFf63SrkobNP4g36PsiQ+9FZT8gYTq1E3RMdN5wSPiFaKBvtNj5am
h2sM6jN2U7Oda5x4E93rAzkU+CgzrmMkuQthoxZuSOm+63FCVzX1Qsm6DVUYZf5g
w1743pON2pm4qRQRpjby/Q6gOjqAnsklg3mB/6ePAYmZ25rQnjfZ3mp2+AQXazJg
tWpr6wfPf49fb++0TGv/MMriJu8eWQ8yNiO+ZRUIbelKioQ4uqSuqMptcG09NoRU
6ThYG6lc43jGo8AyiFDiwljC8O6K/kwQP14yMseSzZ/dXPWhpOTSQyGRHLzTISoK
jTDe/Pqwu3xEUOwUMj2TRrAxSclcX0A+Tp59NWiNpwVGvhHu//qWZ1ASamp1ijKA
hxMOwpMiOBIgpQF35Aj3X05juwQWpsKfv60yhb8XeJgDU4GvEcjsz+AZRsST3IZP
jAxxY1ZaFuDdzQvIuEHKLTEPpWKmLI4iVfUHNpOiam+TUx24AMhyH8n+EOdbRc/W
YFNWa4swV93sF4pitsFggTWPwueE+cnVfD/ow5vjjrqORB5lhZ09AgrWt3qH0DaW
U4aXGqiyD6OzeDg9ERNj8TgRg1Cli2tFFfpQJb9tSFYRKvSx/p4A/Lsp3Q3IyKB4
hxVdPa4+O7SqtjBuCHrcQyyD5fiRVthbu7p/jKKG5iZJ4Vuq3lDZ+vwbZ/MXBbAw
Ennm720g7cxxIg7BdcJnrvqY0Xl/M+GwMgHm6k0qYpCMxzkEIvXCA2jBUzloLfQd
wcp6OsGAqzSrOzj7f7xwp75NQ7NnGseUY/euPE5o7gD6+J+Nmz18N1K3wa9eHU6R
SnV7vfq8LBzzRIq9FeKG6qWy6a7S8DvKDDaMmvuBtJeUTn9rkRSMwEkbYJU7Xw5l
enKzMOLfaRtBB7vPPv48rv951dXYBpnUfGsJRFdanKDoPVJa0w5inxYOOTIEGLiF
TTJTPElUhQqIevQdPlsS7WKMt1dUeOA83iWZ8BCB+UCDl66W5Cb8aqIsAxlxtqXT
ZBCDUBKdvSN6Do4raS77PxOe7C3WoCsVkEXB81W0TGHS/sU/6fzGfPmXTNCKcY//
5uxPhbPJTBQHH8YbaVSylGzLGuLlo8282VaIUigjknFFQQcCHvn6lnEmab5Csh/q
8x6clQKegWt1geR5Z9zWwI7MenoxMcQp9bm9p3zfwyLk77CzRaaeQGtanHhRZgI1
mE7INuk6LZm58elk+tp3/bY5rAeTulw/eZhnGMkAGW8aTKusBvktuZKUU+TG1XTp
xsI4ZBt1XUKb+hotpXUGyA8y1uNWhSYr7wEVc+rvh0qcTqDMdAk6/OzB+7Rn86Xd
0dVmtMjFi0PJXylbfTN+9ODG1SKnybK52FJGKrk6PXWsx+RHCInCm7qxumRIOYaf
rt9U/H2TivSPYLyYqx5vqaR3gRcFp6unvu94t48i6/SI8UONyj+Ht+NCqSbWKCZR
YSjmKsNa91GEjO+9arfi4RBDQsbQACjyrpFgWjXMwnm8o4HkCZmJ02k1DMja1Muk
34BHxrVX61aGRIcWgZ83M9ZKpRJMzZh34OJDC5H0JWeJ9Nl6qKE7sG/U8iExCLK1
YJEn1Y80sNLXnAhlVfidk2/bPE/rWYp846UDwHK/JXFDYxOMeuue3JOFYfVtxILJ
OFFkg6QM180dhUU63ZV9Fb+BFVK+kJ4Bfd2oO7TyQeVr2tcsxjGfZFPk7IebJkVM
BKEXosIW/PIS0jYHcQzAhIH6MoVpY/O3QSP5w46THOMF+yxq4NFtyMn7kUvGCHzI
Z5SDVxRhstOoXTNFlG36Sl30plmP7GqrsmPCqJrmJYmRQcTsjuBmIfVm5nWsAcK9
e7gqn7UCStvMbp1QZkPPhFWKZwCkfIxE6CLDB6zVdgcYNpJnKY709Cweu6USWY3L
qjZNGa86VMrX2AY68dJHrj8EGa0GlLjkg0rocYL1rV+G7tZnqdI5wmlQ9kjlSPV7
ArZYQXPf9OB2P0XHsQqG580E4M/6FKIIoWWexmLeWl14CBcdqD5QRtY+aDbrz0dF
2V6L5arNW/I1va+G23gOvSGkN7Nyo3B1igKq6jAZrCcx8ozkCEeCEaGpxTCLaFRK
2L2NZARcNT3JBkoTIiTKFiEG9t4lxbXgURkBj2s7iQotobxuoSd9KefGPlaJyMMP
3aK/lNQAsXJePqpWGS4bMWUhFfkvIvlzV3l9hKWOkEapQHrRNBuGbgtZJ6b2fQ46
XDSSO3u4G6hFKRV3p3d3FoVT/hQzCHECx8pvqAzzr48yQFPcQrT5Eyw9Y6QJg+ZT
hrpEYrL+2z6eoktxauVoblrZkS/ohYz9zPrCIGfdUsPipJYX5XnWRitO1ABQpG4v
8eqQFeG1JEhtAFmg+9smobov4uKyYtxBHG3WDPHth9Ub73Ub5dSbFG6/XX6MibpA
ShY8S3L0sCtF/9+I/QN3jDN3dY3PMlmHIgSeCx3XjaOT6viV+o6aF1sLDwHSDMNU
HfzvhJ3vFXCgAyCVNwaWmaS35GYoADx9nIm8bvVw4ZJ0ObLZtaNTapxCwdavSiSa
cOOQRYZariLj6cZtHN+4qFFt4bAplF6UFMKSvaWNWl5eDz/lRT5SorGl8LGFA3YH
WGHXZtqbWHFcfSR9ehV2mILCrJ60SYm8tCG+JWgFYHN80qcKY6Yrd1GIq9CmHHJ1
CWKTmDzkj1w2hAWaWQ9l73ZAlh45dsfc8PTLX4q6BPA1pSWX3kR9NkoBR9ZHpGSY
F9f8JQe4r42UeSqa5W/lg6uWJ45KvvQYm7EBcP1WFOU5LRH0lwrVo+cYHqHL1+og
Kt/56dZOZQ35QDvkzV9uywT08/qLyG8UenlIsxMxYIhAAtsIf2RTUqjWh/OSpPVz
yxpyaGkazqMw42r69VEfZib2odU4iX2cLq4PKnOmd1UfXzhvkIgA3WlcdEuT2ZF8
EM9Q+/TkZwH7yc4jL9oWbMvKGx0EHOqcmIYCNfaKZBTJBxrq1UyL54xipSOvL+Wu
mbY4lYaBSERpS790rZrmP4uE6K0w6T/akTGnWisNNWzmxXm6oAS0E0IIIOSPhiYl
jrfE+9gMVEWZ98SvV6AQTSQvrqsKCqL909+8B/udv746VIrbkY9mlUVLg68S+0q8
ctkx9PEVM5S59KsMMcXX0zctzWg669hkeAMxZa+6Ea/3fRtVHcf25bI4zZ6bjEeX
Dngs1Gk5YRpm9ILADy7FwPN38GRlsCnpEHeLeQIzEK4BVGkreR4RxKtHEwu+kf+N
ouiVGDLvLFZNX3oDsLGh9ZwyfqmQ81BfSszJ6LgCO9HcetxSk9xM3h9iLp2jtUO1
L7R/NWPDF0JGn/cqiNrbC1i2Zfv/rLx/IkggJfWf99eeFU8i/OctP/tS1HXgY2VV
Kq/nn3Yo+rfnr9TAVt357bPW72bSBRbZ6NtxBnr0n5DLGCKPW1b7wA08wMzk58/K
YcBAnm9xzUMkWdCl8E/Yj/Hfqdk/Z0dqi/4OcFZgmek1M/rEeCz/3J5EjH1Khd11
XuR9OF4teCsrWYc1sgtMEMKiCAZIPzeBweWYEJhN13JWVvvX0pmHDzgu/WGEprr+
zxQNfJE5TN8ZuiudaV69Wtxl3SeAIkwXTaQMRJo/DuuL1JLVnolX9mvs+9WsE3wD
tsR+W4Jvy83uNCsjieYn5AyJ8a2m1RoaODGsMMeoH1NM2Ej4O/I4nWgprVJdNXD0
e76JnkSpMvOGT9rJsYq+dNadAWwwJ4+IfvbzwwXDK+YsLetAS1dLbglExqUn1oBE
PrH/2Ll7jaiRyf1kfaWTk7vnPMtv/n6qF3onRZbpVo5oXDp55nm0KPhQFKsAB7VM
CgXTaBhkZSVzrGEUIJHF/7QU5jw4J5wkSI8xmRAFT6EkR5jkxQTIeaHWT2G713WT
8scLjXeJFWI4QAQTlQ7AUGJ3b+nTE4CNaFparA4Ps5ENjPJpbnBEIUe9/yna2Uz9
yIiLYNp8yjNAscDT2q7jrp2J1mwkQqglaRWIWGoaWPH9522MRO6xxdknn/PLFIQt
9KPalwxWB4UqtaeJ9b+AdKK+fqt3eRUWOYp4D9BFgK9dyJN+eJzsDJPQmmXjJ6+s
GG7nPfrrRGj+nD9Ze1tzvuseItqcbS3gVm6zc79CYJf0Da8oLEKUO3CskPoeL8wx
o4HpFNBHXuFdBPTXe31AtZKUYFWifc+7fiYONDudE3mOHpbhnsPMla4+JecUQto+
kE+Y3bs/7PHhylnq9JqAtkZkZkWAz62ucfe3G4qytWNW76IQhNFG92L44MXNojQj
djBzVth5V/7cOWJMEd3jxx62cAetrTqhTKn0eQTgyLaA/K+Hq5N7dj08mfseV+c+
/70poNsIYkLIl9UK0AQSSBH+FvDYNHqN1dJdcEIln71d0skTJWPdhsx8IiXMhljb
jaISZ6X5YO2HmR48bMt003qoLfE8ab4HGy/CYcvlktY7QWyN0qnRmI9hhf4+2/Nl
tjQwcpt5QGczgaT7BnKVNozvmV2gsMJa++sU1MySzUShgU2oT74Mbjg1JtHHMdg4
1atS6NKCMWLfy73Go68gCIN785fKwwG7DbofPCxuHlyRkSR4ybAZNYJdHgIH01AR
ud0dNCkOKqWPSITYcDdhb72Xep4HEU4HKjXchcvKOgo/MMtmNN+ecHl7AaDhYgjA
ynDZm/myfpD8+D6CIhbSzdj1vR7jgcLGWXh+JOHS1LSjkpVz/ymjCKc2ZPA+OKI+
WyLvd+mX0GdLjK7XedAPHh2tGbksiZ4YmSxiR5OACFMgGvihOPZ4eJymv6TuOgQH
KTrOCJV+VNsn9w9v7FrAe5lywieqmFn5wuZIuW1WfWUWLYR+L3FMsJj+eandL070
acJaWZi24fLaWsHxbmZtPrb90rLYR82I2vKC3vOMdYptX1dZ9QxQ+kXacr9dlkbs
+i3E5tKv98/h+oM008LAGIZrw2m7c9hg71iJoETu34B4BAkM/w60D+SWRFVoy2k7
WeO1mV8LIQQaReIMhU6W5+iuY0BI29yjs6U6QyNFYsXqigVI8gBsJv1+/BSR8O+c
Tk0UfWE2DWWg7e1/f3wq4Y1hHYZU0OVFAaeu32dmwEGRVuWGK5aJOFVQmFhnHeZA
zPn3iLgFeOAXbRU1B7VZ4FraGova8pTCai8dcmvYB1SBMqln8eFdJog/3XO4RL0b
5GIk7ChpjhvcHBbUUmLQBFpgCKoESKRP2cAcQYk4rIgg6a7G1XHzbzOewX3tzKWg
9o/lrhtBto4vGq+YEZxvcdGW+DosVDvtRcI7IldWvRx4xNHMPD5/uyoEwYLA2gbF
eMGoBPup1emAEemJzrUf4jOPKMXnVAfRTDr/75Y83KY1pIWvNuL3Koh/UkIsq8vX
GOiXeZN8hegz/I60nNwNEt5UfTUuG9tt1jTd5Iw1ZFsMxH+ElBInP4GzxcdZnuOT
NXUfKcPO79uo8vgmbwYfYbb4iBXJVjQAC28az11l7bjAB3MWCh2HwSMAsNZkMzcl
4fodaXhpnpuzK+rIDMC3rYPZzDwHMA2u725gai124IZOSS8mf5HkFALiVepjhXww
nINM6SfJvLlyOUp9nkApwX4AsSOqKjvIucG340jJLA2iFPRAZEsjfaY/In/QLL8X
Z/tEPSVfqQb7tkH5+cDFAsAt7ZsANfvXQu34pE32CvdV1m/XwdSgXx8mLWzOEusq
wm2KdX9/4kHAnSBwuFywWg8t4830XxZzXUZIkJ/gEVgMRC6tMz9T0L3JKqjCWXWY
QkBWzVXKdEVi9APpcCRqjQe0TG//z5YqCDK88eCCWtBMNmvHPfqoYspyax6n9UoJ
XF9BXZQRwR9QyrYtEsv0PrGwG0ba9M527quoK17nC+LvQvBlF2XwZMPzExoipkT5
JPcgoXg3THQ+KES6oPPtGxXt5gfKGIMtEqvRxbRY52+1DPg/GE1ae2dsPwpy+mAV
BDC91Ey80CleI1NHYMdJ5qq77WJcxcMjrQjfRpXEadVpEH/FkNcPal9vX+PQlpMC
LkuZcMeCxcChEUlOCfzpDxNDQ/BUEnD6z0lk8xf2bQNvaZ+IGUjtFYINrjUBOou/
TeIWLNCOHHRhv6SDbTvTpX3Rhgm2+S+gcGv7NZUbXNU1ObbXnXeOUhllxy3JB4g2
B9j9YA8Qok4VSoG1gWXjyM9ZlWPUqvl63kCKWYOD2KAki6NHD5zzLpEUgi/nAUXh
fcWVNNTv++xV6KAhwqn2jffVcLRbqKA2sqJF8DBgqqbigWK8LGaxOtyMMJopHHJs
XPNVg4KxKBYaWFpNrF3rpz2/YO1o9JJSmHmS64Ov9moWspnjeJMHTsy7H/oAdQ9p
dAWAc8lGVyhY9iGOBJZ3zaS2hcdBxBEjvh5eXDTayyqd14NLghRGvIZOc1jalqqH
zkaHjlZt7phT3STUbb6+2UkGAfIAEA1dXPcxl2F6rlEqyE2P3AbBPmaPapHaQjlD
eqe10xj5/NTS0hhIdb5+zpwKQdqxAUwtdMxHZO+JAR7NxyWcFaoaqzKNIcs18jEu
ResbPljMq3Agkl8Cg8Ycg1L7cLo6J/7u6d4YF73Qqcb1pFusbjRKURscWXo/sFqm
AgR2OnJhbhfbDS7463eJNno/MRYpw6qQJU7SAQ6fC+SHj3BMil/0KhzQZQtYqNae
J3KL8L1P6uzbyOPVKQ11BuGJLhYtNctScBKTU51ytBfEep+RXzSAujuWTHinwO6t
sRRrZgTfYgQcw5yo2YC9OSK4BhopovUsFCrdDG1pBsRnjVF4xQBHRMKEiy9R9Mp1
8pEcuQnkV/vqrTgAKiRkeOX7QhcuPJLJ8KNAyA4dnxjJjjWdvkrUP74wPJpSGt8Z
gnfbtHl6xgRuioMej5pM+MifACpvve5Ko7YX5GvHzm6sQeKNq+BSioeJGXM6riGA
fP2P6FEFKuwQJNRBgGpjMRKSYvNbGV3HaM6wJDPXqjkx00eHyx9EkHMD+5PgLCyq
ItdA3CyB3/zGxY2VRMjw6pvlkSF8nqY+mMDS3q7x/nD3wpD7Ze8KsZhBkRPfJHTl
ikXP3Rnw7uZthDNdIIowzhZD1ICAELgG27XudHVa9jeDWTzkaMTbrjgyBLY6MBbO
HBz3XjjZiAh2P/QFEYOpWhpy+uZqDQwnBDPMfybX9wlpg804m6xpgPD8nUUbRAfc
vIEOVSUDMXDoDLrg83O5nda4J4SyDQVn6WXkGu3/pYOLj/c/wJHCfCjwP5ee+14p
YH1CR0MYvXH8aWGulnZ3RfRxqKixpL33o0bC2CkI3j+xUSZsTvU3HSZ8ZmR+Yy/M
53FKFmMbhoIRHvgLoRHaJrgy/xayt8z82stPpdJrbVlLQC3gQudbR4eRXFAS4cpl
uRb5lRZyunc35GbV9WBkJlgv+YjJYljHzjw+AyZDdKwM/jaAiOQZDzMvJIkwjSh0
LrbN8DJvCDfI+o4EiAAvvxckDQaXS7bDbubCk3DVPqMa1iV5twmL9r6jtRg1s8k+
xfFm1TVSAzwmV/tBwo6YNcrJANCEMlqBMCBlu0gBOnGHs1JUzbNq1OwoTmWppHcq
0sgr9M4Icx3bo9h80ur+6U980CNw76LxMF9YgAWBowlL7pt4xznZAz9a29UrI7Y4
IsYSc5/1Tnxm/OKPbuQwFgwOEGCSCyzKMl6IIpMWEJ0o7vdy+zohglC/qW6TGmz5
N5JHaXfpaEMoapsUidlJkyGE3HTZB1jNjgc+9y3Nay2WrfpjiJdMMzX7+M95oPq+
QOlmL1eylPgwQ3q9810+cdfF3+yCF2hpSgaQ/afcmXpLoClg48bikNhD8r3eoTII
r0ittao37db8kWignAbsqxbLYxLqd04TJyYCgFzYf9IMSETZn9XzT7NFBPGYFOk0
rVi9tsLApDQlA4/WNFikpJb2c7EsUfmOg5LCYQctlLYZFMIogT0ymlZZFJafjnYH
hQbRKRPClQmvN7+G+FRDKcUngusbh2CZ4N1zSCM/E7E6LxL0ZZqXmz1mKX3bCIf7
GYqLSv3p3fsM0MmIWhUilfMkbxOQeRRpnl1HbepgD+KR6vFOmiADe+sOPBjHgqEe
9/vBMvFrB7loaSgXEqtoWIYEMdgeA0gyDnbPuihiJ+nlRw+iCVvsDxsYRcmDC5IT
imvNjFigZ40n+LLINXzbA0E3kTz2wbj7q4hNBiPUN0eDTnduA0fnYpyGMQcUfvy6
7iJ5q/e+roGHZ9dJoC+rpxP9JBUrcjJLVYCR05n58ZLNnu92Uk27SNdCoBGTMFtS
ciZlYcawVG0mkWdWkG5cG5xjvcom0gbug6iPVGw/owG5auOzBTfoLyumj6HoGOQd
BNle/WQcft+QNvx3NBcnMu8qYuvFpYKJj1kbdqTwwc6xZuVPvWQdA9IDtppyHur4
G57NSYFpKkN6j3e1q4g0eZ+TG0yywgzO5tJKwufZs8ZQq+MJzT9vGZvbqjo+jdzQ
UfcM2tRosDW+COT4cOUebROz35x+Ik840Mh8WA4GhWMAexyBznHKX7uDCInBDOQH
qCWBIE0igvr1BtcwIY6Ni55HRSdSNfNf7MvpM8BMWo1yvgnHDkMvAjtBzPEIhVTr
dmoiU+3kOlbbqcaA355J3zUYvJlK49LT6WpamhyvAGnbj8hGk1qxSh/LQicMpw5o
6tyaTDhvoHBA74I5O1RIInu84CcafI6JC0/gKaCZBLFqD3wefyADAgrBd/JKYNvk
D8z6N+8L9o6VZv8enJD2G4YcHmYczpa+WlF8m0xDFG3s6mIKLQt1y8dNz1+H1HtG
73FeSjp2l3ZJ9OqcFCC0/GF6EhrE430qUs0qfUOD7mgBX1d08PdDsxoVz0LZiXGt
1mFouRPkVYzJe6I1qcIpI1gssETaq5jxQ3XJRwyAtA94fZnzEJ+FXujqn2tDJ4jc
51rt71RpBTdo5KwSayfk16uLGSNvTYMvofstm3xXzQxKR5TtWeFLSqg063EFBy8O
rFQ0frdlQImAldQjAsoMRUfHAQEoh8zCY/A3AOp7QTMY1WGmaBAiqNK/3bAidqQ7
b5Q5f5nv0WvqBjuhm1tkLh9rOdou6TCfKwrr5kSTAxnS7bnpiLFQCr3S8WpY9vdr
e7eVZODhaVYDyvXG3telnYQe5pk944zfkX7Md57nvy4XfIqczc019/U27lwJSgI/
WJV1+Ij9AS07V4I/iQBJYHGnrvxjLl5XLyXr3tqCqCA+s12NWzV/dKsO7TJpckVp
q1mI+DkcTntsCUSxa4JlAH70Q3Y5+nL3XkPrlLGs0mL1UzSLGhPqvIwdfGzAtx7K
/6e9PMsmHlMiou21192u1xy1MGzjKeLfKCm0/Mw0Gn1aFs5k9RRzUICFx9Pn76Xp
oPXFRnDMVE9ud8htL+Pu1L3LiFWjnlI8sXkJS9dHSpPw9HAsHB4UpHd9zRaoH+Qk
oURPQ9bU7QZfnVXrgwmggraVUbLINpubeMTWRmgPIata/duS51yRcCQMu7V1nsdn
yJLm/Hsw8IRRXVIVGrueIJy/YUBtqcyCheXVnemX70RpVs0UFeHgFjQsxYIijW75
dv9Qh4v+fRnTM5KVld5wAkqMewLswmS6NxE7LAHzkviewiGrXQfn6NT/6ffAhE+T
lSim4caKfLEs4Dgf9HebsAvV33PTgy36W9kTQ1aagEiN9f1ZQ6nsIltw0QDh5TVd
/0VHjjgklZ9sghCBhq1DbzFSmXyBk+9LmWFB34lRGI94W37woSS1okKIAGPM3Vdm
BFWX8j/sjquyp7aJp/O0gpwlV9MYnFoFz9bP7sJHQBbVnVuDCVbbN8aL5n5OcZHe
Buze/bLKNcRHwfsq8OS1MK2IImr0DqC12dPNtM/TkZgT+z25P2dMueK25mQgI9IX
B5oV2SFobZDnwXBp1wk6J62t+p965FBqyEGR/FhWlzyBq5WrFR60IDBEE4aDM61Q
qfjxdyM4fVW3OB2PoG9ENk3BKrOuWGSz9/tnC7suh6eh1Wg7dQXa/AFZo5T/F1Lm
gU/5CBNFoNcAXa6NeVnBLd2N7vsrNEAkmwaEu6IJDeTYEDY2zIwOqZC4PyRfIzEy
RDIj8qF58SRliVzgraL88BgSy0b4qyXEXyBXXkxd8z70k75me/7LDBQMm959PPMW
LJ+jAkB0Gf0Q+nyXxjUcNT7gxgWfZIAEoKLX3PAWc2dF/2o4PDH6jJYJqcovQ3EA
c4GdBlqmZYDTyMMjv0mui9vaVr3UBMTAuTlGmeSDQ6XHC6FUbCekcpRfzX/LRrTL
/AgavTlMyPxnw6ghbpSRrJLWwpA6hnDSNlPuqZy1ZQEPLCohYXJ1lychiHQgc8cW
Q3bzyXMtFyhhYbhAhLt/yX+yVdDEDXOqjmK5vEbXWxC0gpK/WdJ/BPMIjq4dA+Ix
6mW8d90chQ3dk+j4+iZscl1q/fA3P4KhOyvGi/0aRC7A8l73MFUJLJEXxHhUsgGA
BGcS6KpCuy4qm4h23eRFpWHRnl/r/oGGCjBdN+35Mf2ODa/O0rNY9WaGocXynTTG
kdNsKZL43QMmWhNT96luS0BlKnqSjHhY99fxI0cF0n7nSJMmVpAh3hV9o8K1GuCF
3TByRR+5RagDBEmYGvUXP0Q9LHSQTB0QvJZdXCW0mw5jRJg3SRry7gOtiTTovwk0
Iq7ZyUl5RHwShU/OFMW1PDXHLXeFB80UQQP2DBYIFtd7yc6of54otxwTGn84VBCk
FWJvhdxbdqZiLmtPFFgqm3UXhTwVSnnYdBcuyC+gAS25CLbegPxDXDwmW4QpF9Qp
dEig81AwTZzK9EtPlzzEGnmgkCg+mr23xrJ/Iy3pp2UFOk2e5QP0vsWdDlVDIwb8
BQSeVooOH5V8uB7WqoCOrqnz/d8qEkOon/P1uJSETulUXICOBs/B8kclGvJUA+cy
/3HiiVHkokpsaOaQN0yrsSjq3EFlmVbN8sAfTWwt75P8Lc9Lbmn5f0wGRIu3OYG+
NqgyQKek3deLewCL0Yve7UwruuRpSje3rwjEvlKCO0TpPr5t+33KG96y3ebO6CFv
6+7xDb4Z0yFvk9QUAPgAB1XWd86C03Rlg/84rrIquiSoIZ15LJvpIHSZJ6FjMEl8
/2bPcrd2J0qI4Hs3m8I6V3kyJ9MvvdzK+yv0McuzEKz9WMkEF+oJ/gItXgPU3Mc+
JJcwy6xuR6zX4Xn8JwXNj8BAsDT/RH6jd3urwk0vsuvlOBrEen84KvU+aiGR0rnp
j93u771S4i7t6KnAdpsxBHAIYznMrxu7tYHwMjif6sPLyApD6WucikNa6ct309hb
kqJecsoirto55rosVyTDUTz5p9X78DGtAUYS7LcKK7MyTiMXimp2lyupwu2spIpi
xkITrWbxfSto/XqY1P6X7uMET6t8Tl8D+nURpVjhXE3qkOmU/CQgab14bTHe2VCh
J4cc5h9k7+k0zx0GC6lrQWg5ujBpluJgzUl8Vyog4waSqRhn5UgKjAVLcucUfTi9
RrJf6dsdDJo2R4dmYVAn0g7G+3USeyNWiPfffojTU1CL3TAJzJbpSEG310iu/vcH
kIwTijfGFqpHjnHS2nHLMytRwqoFRU/Do9Cu7J8n9OWnfcKGv4/DjXRGDR0e3Qif
sIDfNZN7ymExkrMxQ0ZJSZ/CnFwp9jYLxnayWeFYE3CLrNKnaRcA5Kz/5YoVj20S
FENrDBob1rH+W3GGTXGvEikALnkYZubB6TDPi3v4J39KRQVIKIWpRyibHLd4pNQy
zIdRctHCIDmio52OHXXOyHVleZz8Mn3Mw8x82CXf1AFmFGjue/XHvuBZVMRYxkDC
lNGC5sHiU6UmbqasWYzCYtr/V9Y+0NhI1dF02rUL1oWGTjHlk3Cyb3wZPVI5Mwzj
+e7ohIZiPWdFyBOrThS+yOOGhUD1yYmkuEDmCX6p2EevpfV+n9s96l3aY42aNnCj
Y3zMbHk4DnbbRN0ptiOuVXwjG4Ar87cZrcoDbzRsU21o8Dcf5pwEwFREsjUa4Bba
2GkshGVBaUIqsBSRFGeF+OZmgwBm2JIHeqxNM3gCCETddBDvZQRmsNWqSgIgEhc/
VL26yALmr2fXWUBx/dcdcUT3AJaDTwe0N8tHkILTWfmLVtmJc4z0oH6tcGFPSvwo
pPCiMqadcZ3vveUhyjmL1svuBl/K9og1TfMP18New/dVoVWp7czfFqx7HCBMn8Yj
ywyWcR+oehsj324VjXEPMEY1Bqy+VtkhLFM66ov5uD7gcHq/hxZ8hqeV+BIPv3lP
8GwhBSfHLj18Yv+JaoQGbvZ0ZXOIbb8OkuA9aK4GGeUAzHGcJg1nOLKyw6v4MrJs
z7ExQlibGjZakefZz3rI49CA8JpdNk+3RccE3/aG9WCMejCYCI9N9Ktbp2cW4xYH
Nr3te3LqmQ+1+IMTjmEmeseIE3cmBlq3hS/w3J7H1QjoHUh/WijaHDdlNfvmgAfb
lOsa7t7Diz7N60zkY4zNdeQL5wmeOfNLRY8k+BQjFxyIi8co1Y6WL+SvCARJeiAg
TQwv4ZbFfHujSoqrzoya5JStmHnIVzYKMxgJEyGB5wSbX24Jk9jpzB9Um45YhY9+
FZj4iv3+f9Tl0F/h3WBEJPqm4+1/mRqMt/62gq3iBzOZ0jjpF8XY4sy8UK6qlBgc
pSZ/6CU4QzUczF59MFe1ISQy/EjxtG+bf2EuzTQ7icmErBCxlKwqme1n8y9l2IJC
8rAlR7FgDITiHtkVHiKzRrY7CcEdmikB1/wNz1uAV29a0rY9zaqacHDdF6I/aPdS
7nFcMLont3I+4mi1SQ4N/EWgeOEFnRSOlxIXuaEPmv9U0YO9PJ58hcMolDH6lbtm
w+4Zcf3k93VtPZFUe7YUfTlmrQeZpLVyzzV1gydo9xxHHDtsWz+3TmBjc8d+q72x
jNYqVmUiTQoX2IjNjd5kAMgmJSZ6ILNn/Db8vYgdybQCETqQqnOB4XdkA4ooQgaH
oRyhrkKOJ4jwmmbsHbBP2ZX0bP4BBzkZeBAZ5gWnNG+yeARAPaGXgAjHVyTEmO6p
OaAvBp1fi4ge6jyUrVajXuuuqRPJxeSu0Mw1Qo6v9W97xw7g/KWbpsqzaVbCCLTw
vT96aTfJGHsTptJAHDHvwZAr1jSpvEekkGoVK3NiZ8Y1/9hT1SNPhazs2hFZsfdx
SoTesp89Q8tOznx6bMPdcumjkPkueeJwPlII45B/FLXtexoX019xYqIc5nV3kxKz
P0f1qPK0dJeidgAD9Nd7AcE4LDMtGJmD79Hi7QL9qAavuXhhqQz0goZMoL6xadpq
PLjevFyL1rEaMn73FuHb3M0AGgIzzVPN3C9L751CBA0sYMWhWIEAJYFcqmd8eqRR
Jqmq13PJ+u4/WGSrgC0TZ1X3UsAy99gqm4C6xpvfUo7yH42of6wcBBpiUnuIUoCx
1X2ITq8A6kcf0YmOuciZCZYyJpO+bwa7He4PwDb+8COS2Z3nHRWELiMefT4pLOnt
8/Cx73VGNCcWt5NcvJN0lYHaPybNEa1uMQa09nphP3faIXu6xQaCSL7MONkbrOA8
kZF9s5vrWUl+Fi+ES2LT4JpNF4ZkogeQgOQAHsijND8ShzfIgbji4b+ee8MdVD0h
PCDvy0xVqWslVS6DHrcHUNQwS6TyrQLNJpQgypxvkVi/35GSdDaOPusrLPYatm+w
kUkBnbu1+90ze+Se+r5DWySVDAu34Ufe3iHAxRfbsInhbtsOW6463iqhnja6+MkM
E2pwR8uUUY6k5UXDXy6T5FgVYfZBu/xUYX6Hw1ShMQRbA/9JGLAXFr8RbzocMfJQ
3lOZNNGp1plWbxMvSI7ef2Z8xrRXCUdNHz0Z6AV+FTfxV7f2ZPxIiU3dvR5vFrei
rdm8YzofBiMOuGEzeLCDigNVoQ5ni29vsMcsSWKJFwQFQu5QLlJVgytwYmsRmPg0
2N9nFcrzbE+l8sC6ab4lA+QopQXryB6y3MXL2WGTZ+MeZ4ZB1syJaMkBd83oM5pG
tzN5utEQ9FSmZb/LTzmA9g9MQVzAKYC6DNdSNrwpFW6v8ZYAM3VrwzkziRAuWluf
pTOi87fG98Per65UFNkJLgCd6Ttl32XmsOGvlDjr9nNpfcUiPHMpIGN81YgnnjYk
l5U8otqESrogzuNk44xlaeR4SNvyWUOcOBXna+pcKb6xPsAyQQ47g5N5M9ww2Ics
VM5/y+MRH/JYwiGKldoao2qpRAqOgDyhAq4Zji8VJfcwgHwBAcJLajiAZbh05DA1
HeRyIwf85QJN+XZgX9IEcRu4HPDkeUg214eTQIcz3w/GQT/zyoisL3Y+i7gz2eVQ
hR/MX78Jz0FYaByY/Auk0mSDosaBuxmQfjRz+LD5VdJhtQU9PA7UlcaaF5kdpvgA
WZwIcHjUS3c94esfkU8dK8UtfrMtKrFRVhKcy0R2Unhlb3xjY1dqCtK5POuGstfl
f5RSFHLv4kZXH+fwShzjqBMb5zvHtcFoa598Hg+vFPWifaXJ0CRbsDlpjNs/C3dU
FkOJoJDlKeJ/b1xEMMjlw82eqjFm9hluLcR3Ea1Z5rCiCxLCb75nVFerQzWiPct7
D6mpzmfFw8prZpq3KFG9BA6+E4DmdQiE4imqUyhezQExbeljsyuL9DBWkGXmy/LA
X6a5oVkO9ZwgVG+++bXm3MLJMao1FvsElHj6xg71mmHpuKAp7qqQueTeve9MuYZx
hH5f0C3dh2seEUivTqHwc+zGmO3DzGzRugH9z9JhocVIvrbrwtQRcaV89JerFkbc
FLBYkSM7fRoFA0v4UzubtFMWbZtY6nUkslLDQ0DpINF2kv79BzdTQpBycHi3LQ7g
KPN9dU37wgaTr4aXghZHrI54Jqzbw4oArSQslrVq9u8UbZS9GsWXAMlb7SFIIlg1
cNp1SrMmd+T03bLa7xVyrAZhb0qNiy+qGReLDnGp4l3g8Z4k6zwX+Z9RXjqQCa1v
IyxPLrOIQHPkGceFGjdC0pvgHJm3njzpur5/FCBYgWLf71o3dg1nLA8MIKMHbrO+
l0bqBo+sJXhPTVwp7wauxh05E/PK2qG9Jyr0dQI9E8V8ziwunpwRd0fAigPKkkwg
QmfnhRrrINwACkytlwP0wftY/mmNOj6o0ckYIQkGThvKKnOgTUEXnZ/xiNNFVpsp
8Y9kv6WngHmTwBaFGoxYXEKc9Eb3MnMHkKC9o+aGjb8ttRKIQ2jQCjsJHC+aeoo7
eMrJc9yWTM5ygpBUaLzlKv4XfjkXBCrYhEnqmRBO54cU2FcD/hicN3DGaEaXHhdb
sxAPrasFHj2c+yZocjB7jv0zjNH+2Vch++y6gtTv+hGDEpFMZoAY15T97X+CsJ3M
VgH/na1W0l2n2vNtWtrJYnixJI+/nzIGvdVvk/Sxc08qgqY/fbZAYAUPoG8qn3dO
Dv1D8ot7Qx5GkErEg15dG1Kvm+Qrd5CKLF3BxUyUMiZV2zIQxNrakVmFzHwNhL7A
Y2V1B14CopDMI0uNVFuBQgiwpJEBEEl3O/+Ka16XNYjD57sfsrQBktL/LBtN/x9v
iJoYQOrT0G5Q8k+QYbcilNy7eOd3XRpSHKc7krUdaEhhP7h+G8gPE06EUB/4i2aT
Sfh+dipTkfQt8PJoAeGLXwowwP9Det67LOvBB1AyxNFNkDny+tAJNOUPrNUJXiXD
G1oek7Hh2zr2YgzJJST/nh5cgEJLjqnF9a40PBz/S3ZcZTIF4qt7v7fBHgwU1+ps
ZZgxcW9Vk0u4Jw23H/xAz9XZAvSZIurk8s6M+ssi6Ukh3XzoxQ0XnbEmkTNDMQe3
JLysGiqHwj/67vjL9HlCId6R1JuswC5NDjKaa1ekEv/W3SuDteCvtpet+9Fd2Dww
RB/GHMraO4aZto0rWXv3R/hb5ZPiJZjkJGPOEnRJnA5wfjmysJNuEOshb/yXvm4K
RIXQ6TT2hdHmx7Whdb1caTPzbNKk475AlMdaqMZmILbX+tIzSIvxg9XPgmbORsFI
m3F/lIKs78bemI4KVomQRsAT6071mO+jUQ9bovjJ3aGinzagbifCvVsFWoRDMt/t
cCAaJK8VdT2gjnypMgrK9aS+E66Xv5NhADj7Iw4wLite2t6MVo9BTZyQLlzf8g8P
uWaCVYtd4YDE9Kk5AgT33ckrsn/YJttC2Qya7Sl33oAuOgoynDdGgZ7pmMwxMBUU
+MJdAJAjTSD4HZCRaWN5Z0K3t27faW0st0wK7rM+tclkjm3+ASoH6y4EyUleWChP
E64GiIFpgP+nS6mVdJnvGHFXi7VQ4SAOkm2X58SZtgmWrF5AGyecAycJzdMvDSmX
+SeGuEdFg4pkItpwV9EM3XHgzg7/TGmybXhy9koCvN+o1qXXk+uDz4JoKYXNgb0h
4jLayf72gVNigFg0RI9mj21tbxr2QC/0a47tBoYa4OB2qh37GUZdFb6ETwS2rQqZ
ivkZcko3VYuFX1LuQKdPK6zZGr6+XalrDZb97XvnbazOXkLdCGnxdN6y03Cd858d
4tGfObKOc/rUQguNeWwZm2X3e8cRU6qUvBlw7qv1lPSC3bFdnQ9MomlVUYVdJ+d7
HH4mOUxFu3DRfC4Hxhjp8zd2crBaG/uxoJmDGe0VRM2/qz0ARa+vqSyBPoGThgcF
SwVaz9D+X3Icb1dOrH52U3tTIeSeK8XMm93FfwPNnpaChXdiufztgaVbOp76wEMD
38+OxE9GNpjOdIxSbmA+zvo9Oe84KICg2htKFqjd+MAGQepLzMLSuOIlrqvAWXxQ
ndwHHOcylPmsvYAU71b5jBKcrRGTvCm53OnntbOD2Ok5CfkA1VZj6KbVlF5Ofrqg
aAFU/LeYYGJpj4qz+qbGwaLoWoOcNFM4fPn/ooHW8cIXn/MvTVxrE2cJlEP+dhiT
6ly9sCl2R7Zge6q3wr14dJN4V1tHfmtvgA+OTzfyNGQwlCMhATK5ANetIP9lPjEH
5u8F1Fha5BMA9ZJudsABRJWzPur7AWTx8B4RgQCPD5Mr3GXWvaK5Ws811yXGBDeC
JxXgjF6o7304UqrfW3zSF/qI6cYAtWFPXbxrQAhNEFp4J2ymHNDhfDU1OoBQvmyS
NxW7inOXk9DkFS7L5EDkVLzatNUzaJaSoItw2nUx4QY/M2cjdmyNLIelmJxG+B7G
b/3XrmGRMpyVjyGm89MUStkIFQuj6sAM2n/n/ieQyQ20BtIJzFPBAI7tKLwx/9xX
yNkQtATY7DoZL/OaRbv2FEeAZGp2TQs3wdH9DR44zBlU4LCrgBKNPZRs8TGISy8l
dRlcdz9VmI3PwJioMl4sx1R9EnlxI/724gYJNMAaJwXU/ZhZasbewW91fHJ66VLB
n71FlG0o8pL5sapalkpTmAYWb3iKhb7p8vJCAfp3cWzBbYciTDi+RngFaDSoC9LI
kfGOSmVfEReGX99kQLBolvICHusmx4EXkZtF/kDFeGUMrsEOmlD9EAtm/DHZOSq9
tZsNIrSQVcmWKzYQ1GVl7GZTyWYdKbWxF6wH6G3eHwURisraLnEjJ3F3raSH7HZZ
6IusaMjKf37r5jFSuQOEZy19Ue1HP6Otgr6FtQWWltfhLaWiuuay8Mrr3c4G1yoY
MXgokJQLv/6t8uKNfSeYpUHTuM3z4oIekg5C6AMKSqwf23B8j9sCBLdPl1QYgdKv
51Ue8DS3Fn65Pp9GAWrIL0Fdvetd7iaLfLMYu7dcLXFQJADQrwPMIMroFyE6yP9P
HS3y+Ti44ZXMJXDFfBkjbzfIAv7NSY3SFrhs3UBub80AanvkNIZE+WK6+f92/yPg
3F6hXi2WpTan0wk4NprFaG6B1ela2nImXczIqdwqzyitxAVu7z5BHw4jyRwo3Cld
MT5piEQOI7Q41W2gi+ad7KvDM45kW3h7YVLxBUdvANzvCXqzozUIii1VfmOJJ+ST
KBSdyzypAyr6nOZrqhbVn6/I8tlhJOF5KeJXcjVCfVKQm1ip57VY+s122j3ES7aN
x873+a+qRDU/4Rr+mM156KvImW10Y48mJCnzTM5oeq5PCqvOeQFE+eBxeTUy+S90
mw2RY6tfrcNm14qNkqxTKs2dlhziO1OLbqnCz2wUj5tDPJ+t2Q7QrR8gwoYTTkEE
hfEDCX06RmUTsJlh66yDbZsAuepUuPSmyeCJff1K3GxlEHsWBzGABdPbFihATKxl
VBL8k6hdS+n8jnfhNGBUaMRz6a77mJHnfRgA3EgCghXSe8Kykxj2Ki3Uzvl2vLa8
27rUOYpuzvTkKx2VyEHAL0Czv+gP3gPlwW/bpE5fkW1c/K5UZMzWfVe6AGutY41+
O1eVxcrhiCi7ABRuLMyfGVFYOSE/Hdw5fUtTrwg51wRH+m7OKqJ7UanhkU9yUGey
wz5OEMHyqRNt23WpksZ/TdUcVQkB91K5P2Y2+sfk7imlyHCbVKWTghUIMoJmK8bt
5Jq8wI7bin0O1xFvN4jqyIgYY1FFUOjEjKq69/9jIIwmcx39XhpBzHZw3lELhB2X
v1lMVGedlyVbBmHlTI4OBUGRexit7QLAR3iZMjhnmaKMkvdoWM2Si979LSDZJsBm
zIa+3m01qHOPfROJbuqzKx8nBMsPFxjP5qNifFv7TFmcanvemWZ6LPRWEwrEc7vW
ZiFPS4KbC47ThLScVGrORVDbeWqXBGWhJtpfFngcpTwucWCShcDeZzF3sqiyJXjB
yTLzT722/vnwI6pmIs5L5HXsExSjkNaV1Z17rrinA2dCnTUShjlfOvgHX13rplbO
Y+s2pKF6DNmFn7JlWZ3c2EbQMmFyulCImLK2q0zpPp//BopPszbGDpKch5Uhgt39
nFVLi2a5lIZKM8Kpbg46xpNwyNAf9VsXKG25XvDt3hsAdJ0WGn3SAPAk5v/QR6at
ITmofyeAuiMpjYsnz2NsJmF8Gex49ky38EMkRz/jqrAKRvDufZCe1cz1cBfqq4KN
tAsD0mZGH3Vs0tgIPdQvFitby2k/G3Jbvr3WFN0H/TV9/G2Z0585almhcjdp2lUr
Te8EKVAlyNaJA3X1zITPwFytc0P84PAWWl8LzjbQF9KtlTnFIp4mvfPPIB0JLzzg
6//TOQniXhx5bftevPhu2cGbM+Crr1yJ1JzSK8NdX8z0pK46Uj+/zCIac0TBiiZj
xiZQimQEfRaOJ+qtvCKTB8LjUaJUh5aX5AnlvJjfuGMY1mDevENZIe/jrmTxKn1Y
RGmojH9YCcbG+3wq9eA7B3xdTL9Dlf8mkICl20L5YLRlKu6EzypkwcShdJCUSNRO
TIrJgpf2TCAnMSzC+tAhbiwfPzqPisx7+B3qX0xmt6G8IcKk1p7kLmmQYD+LTolm
Oc5sx2O11vemr46aB/jLUHHgRKoqV1zKhYxEU9t/l0+87fVxC9k38e1EO/nXFgv+
TnlhoGwpDe/21kPhRhV8Xr0ahjeNJpMWDnkMIriwXOl2AiqRiyQR8sPvFFsWJA/1
eWAVMpI2MtpU2apyNr/Bf3pQWRJYiAQXl4j21uP+0U/9NkVXw1xU+lXfe0EduDWZ
iu1y+uOmLylyT2GKDSlR52acug/5W5yyBcETPiM1BZ0B5oBP4seGXFecTmTt81c+
katFVw2Uk7GwySmL1bOZtTiK0cgw9qlLC8P0ivY4P2ZMPLjBI3tOhlvWrc/4cRBy
Z0z5TC7sC3dW1uIMG/SkNV4hKWz3Y27lj3lFCRQia86ZFrRhcsRMuB8yx2wA3bJL
x6iCSkGEuFzaLDjHvRK8h6o21zcxuzBMElGTt7ADkJ2vjBNRxw4JhpReiMn4wr/G
HPpq9r37OB/94MY8qm8NkNi/yMzPoyF1slu1AGviWUBpocRHYbY8UoPY+RmC60sR
4TM+Ie1Ft0b3RPoukekryR5qebYzDyJv9Mhqm0GkZZ54GAk6lhDDMGxQ+FnJKqPG
ArlGE7X8VVpvTZtN4xW95iNdS49woZGWi6mkvYRAnkMhNTw1tWop0/tNhoLDFIDj
6oFCU5pyBYegjvrNW7vtSoTHDkgQeSlpYJtH0SOejAtLqs9UrGc1M//t/Q0LR6Tl
tRO9QondM3tnbC/Q15l5+0wI9929tzY1HHXJI2YXx2BMWfY/VOmBMQ53X9SujC9H
bVyAwQf/tNnrTDJajHtm/vP+2HQnz9OTOhRBwsTRDYlvMqJRtlxzLIBg0NvSe5I6
i9UpKc96yV2nfTPGuolNGaVohYRPRFhIh1T76OmPvWdmb1BA2e8IYKigtz5GODLn
21hW4I14jDha5A7mu+qg7KMsF+0arpfjc2vYC9pl4EmlRQxh30MmEt4ItM4OcAi3
Q3I+oijIhc599GSwmu8heIcAY8+nCg7ZOQDVfUQcwFYgc7O5qimtWWXBXclTHa0K
ktvi2m+IgxB7Y61/qiFVqSbl2Oc+D6j9gwTcchREmDguMegynzdwoiKio1/5KZqv
PPDKpqSsWw1MV/DRu1TWUPeH1ATxlR7O9SrPIp6A44ALpTbxe7EXKpWnt4blfkk9
bFktQnSR9+VI5UJ59UDJkiiireOIl3QGzCfDBK3JxUR4Epm2T0tCU/8Exu30cR3m
xz6JC6UhCBwfLaDry+vcdtZM0vUfi60qqC7G+cYp0zZny+e+S/0kHf14Pbno4VYc
6hKBNLJvLxHaGNBzi9CnZxA7qo9oUFBs00Qy3kV9ecIn6KK4T2tHp4teoYr0Nm5x
ZA+VHiJRudkVZVDvULsNVyPmkYS54UlnsvTAAsBC9PBdO1XuogKVbQ/rK81jnqRp
t6g46czu2St+0SOXqhxuBq1UzBaNJ3ajOUetribacDf6qFS/h64QLOt3mnteHF+D
05e09FU92nHfzITxkyNXVCbzo/J7BBJ7/KrvxnLydHrPSS41pbA4TlIUcEyyqZXg
bDJhKdjtIKEBXwubBZeGUAEfKzey26FW3/AUeUUnqpcZLA8sT6n8pl0SMPHRoCsq
yqPUaWpvJOOnqtI+GR2YEY4d0p//CbphKohiepJWr1hreA8sHj1zRHxzSqgXd0Dz
S72ZGaiEIxhOkDFFtPtL71eq73QDG4F54mGHybIw9efD6y8jP36Rv0MBArLIqaGF
Xd7SmBaB3HEOGnPDPDCKRVe+X195AEq4JAAbsfqXc6qc9NZolzMFm3OjigdD/hkj
vNElRYnyIq7kbYQkypvDLhQ1+Q5hy8nfBDz/KmqnrZsF/8P2um+brApTEK6snDmS
O7xXZ1+uh20Cl6PmwFQ8U/wTYHlTCtEwtiT6i+AovfMqsi2B4nilhNGbYHjTZZYK
FuxJv4TwFTNDZqZNHr1487eMXH7dyv3oEbbXZWXakL+QtZ7AXVxHwVi4LK3Q36zW
2OXBKQQbA4LsP6FwOi7F4huQh1k/jWYWxH8VogaxqnbQ2fiWiN9nhuEIF6th1GRF
WDcEOwVCTrXgkya76hPDWX7yLWQycS9LRRmAzj6IehPhx7KETHLDLZoZJZssDK1c
SoPEuTy64Ana1YQQym/5bzZZx0JL1OSc3zaZIsWdGmy/60N+aTEam9/8gCIIt/kj
mkyn+8qOM0jfGYslUMRqqSw8xgmCqCBTHAALdwoFqKblr5u0lVmrXHXJDKpLMiWN
7enYhPa1xsKw7fwONTP8uSCptcfZ5XZZBMNzUD5Wa+VNvebIhC4VF9GxvUv45k7V
mNLFUWJCUj3jIA+lBsardPnZl83p+2qjxkTH2thGc0zBkHdeDaFnz+Y7VB2n5jqF
Xd8lgGZU/jQJXO0gwojzGy8HVME9Q4rru3YL3WEqos1vsTUkCR16vg9cHH+FGorf
3XjTGBJ7+MY5QYclXTeitiVmWhTvt9w72Px5z0OBlSOB9k5QyZG+Dm/D/oTIAnzQ
rLc5STdSX8TJOy5hShha8sLryu601NDjna+SUa6jKDPRquYBadMw2pQwzwHJe8U+
Zia5HPwUW1s3tHp3iZVuGIPG4V/kUBjXcI4lrjaLVLJlGUdMOT9PjWsPmw2B97om
7AY5QdzOZfkmUV3DIMqYa+/eTZwlHve1tQfakh2C8TT65P1SFFxwu9bpE5pOm6bT
5jqVjMbk/kllTY8SVR6PUK+BiRWqYHAyV/vJMf9NDrlV9ODFlQAoYk0RAy82uFcc
YOqemx+S6AgCTWbVD3+R8H9ZsWQw+JNyhwM/tu25EkVYd2JBbiCFjHAI95VU67lM
1fHVbaUUI1m+P6nixsD8MAGk/vaTdjRDJbNzskxFt2uUs5KUgX2MMmyK82lu05HM
9GGYek42w3BcrbciyT03Qks0ZcDrd1ebbBtwQ0UY24UHRmg4fZhdri2LogVWIFX9
oUCEjSq9SCTc6lFRiMad4rwnWvZ759jGo9Yc7WvcmXC2wD/vb+oqyPTmIU7NIU1n
WyAVfAEo/Y1Fo3pvfPBnnb7lqLLGjc9nkf1pB6uTLaIxaDciNqTgzYONziykSjQX
j5Xv49gIGchJG/IivTobpVmwoP20lAYVFEt/QBH3gCeaZ3TN0z73bsFcnh19JFs+
6IvKcw/CrPFdI0XpwHzKHPkzob+mPW6LLj+ti4bcwZcpqVbZe7TjpKVS/Kwy7dmg
h4QhXsA0GP7jW8GwICr5F63jJocnrbGhDeiUe+JFiyIqi+6MuFXWoImJA6BOniez
Y9wEQDj+hDgzsxBQfDndBcsmKyLAZFxgdFbdcFWLWjYp1Q9vTTm6a4AuOWVUXLs3
/CCPYJI8Lt/tqKmREqekkJ9SZ98EPo98aHtpQao0qH3OATeyeRYAKuSm8x/ZgRcU
mQKYA6LfSjf4dxhPbN1pkxgplCjZwyVyGRh0LEBnyNTNXDL6DENPYJwxny0/crL9
84KeD00rCgxQLiincDMbLj4BSM8qzQ+ANMT+uZu8oAJxq8jZnXus7vbAOBW43ZH0
BrsKKxklMg9W9T6IX40zgMhK5QxzWhYlkrKgwPQFaM6m1ZL3SQmUQgRL/uMdydfY
YTjG6K+grpn5bxxk4r3kyZjD4mC7ZgOBvzsvBetxpdtCBy05y/9or9ynYeEcGP2J
DdHk8t1kzXeSVI8zmZi8MeMnfnZ1khcVK+Q4brxigK3TRJAvfsjlJF/l/V6G161D
flQtbw6xoC3E4m6NZZtsHvf1k4YVWPgpn4/TD1D8SLArJdwR4aeU1AL9fb3kmHC6
tn6zt6766iRsnREc+EvprAT5UtevHLTQXQ84iExb/vMCkhDLD/IKxMRmwl+sqE6S
RkwLACM5VrRwHVCNIZV/mLEK96q32IXP86Ap1LviVV1mP2rLGxjdhVfca87i7dOV
4E6LQZXoyp1bL7j9jw/gZtmVa3Z+773rh1FKt1+XzKSAs8TaHUPfvFXZY2+SLctb
1qKx637keO3zdcHYoggLmbTYCW0s9A5WFd4hoIABLeJ/B0yw4WhDATU97z9531YL
AUdEi8YAWYdBldhjOqrwshKtI9A4LExKZYnMWAG7ElLbXcVxp4BBaPPJipX9G1aZ
SLAY8BKRb0PAPhDM/b9lDyop/MwElqwFEjNFgMkD5cavtqzKZFmo4dpIm0ZtZeXV
rjmsZoaobSZqS0VHT+k0XfNkWyZU/MbHQongZqEheh2G2CKuKAsXIsWzxeeqrdnD
+P+7qfmSHkOWPDQZM9s3gRr41MzG/iwo5tumEopJwH61ltrdLxh0vg/PZFvNMLLg
Yhs9MItPvSt9qZMtXIuEOPeSFHRasncEPjlDidRiKmEIcBoDslPq+10vp6jjRxNs
cIt/ovWE6v74xU2tURs5/kaKpwiGw30I02LRHynsr9OX3ZrfE+6pX+RT1UF2YWEA
cWMpLqT3CXrM4/bHcY++3ZhJWfbr2a18xRuYBqqTrfrbpwPx4svzBbIBftlOP9ln
Gx60PkQMQ93939KH0VR70nfifLEMpxUfsIjpq2bHzwOyPq4Qi6/FXFyK/o0MzBLG
dI9rLJzWBv3RYVMdLG3gPcB/WcQeWnN1DxB4hI3FmVT/u3mp+ZN8ROHn3ZEkEh2i
LahsosHp6W/N4K4ZT9FcJDGNJ0Was40BsAkH01Ao4SdwTI9us1dwyWHfq25O8qZ4
71t4FfyZAmNDcphW4a/yB9K7rL7hsxncdWGwMDF1/fJP7zxQ9GRz8Y198c+kmIx2
J1+lcXUC7L7JLS8oKFjko6vc8j36cmZvEgjz4D2OCXw6U+82pxVK/6wrI+edtDDw
WuTOqlGKBzjn9df6d/nFsPmHQgrl488Q68MSu7YzLIw6x/NW7TM76Gv6pVaKYCvO
C2Yb9J7BCOpjW4/J6ixsy5vzEGE/vhbrJ6k11t6sgJSgXzU+V0/p1uTWZx8DNuAT
CDZ0cUXNn6L4Alid6iHWAChZuMalOVcGnHK9Qt0c6rQoPFDewY2BycG3A+q1POJH
gSX5mZn8GW2wIpsaRomK5COb875o4mahnb27lptkQqSSDC4PLBcURfass8++4eEg
H1CiWDnQzHehrkKh5valR5kaeEU13XLE6XrvwwEoIh4u3MxIoZAqenHX9BDVMaC5
SymOYnQVLsEcBZ6ufCiZmy8gAHuRlEXe5IgTb7qlZ9/iX67JYZbMZSymHdlV3rbt
wyPCwNNTAmwZeP2mSLmEA49T1f7wrQAI+eAytT9Si+0QT/Up6V2dXHYMCdt5t23C
FXzUowGKglgEEfbQN4+8u7D4HOLtat0vclwveYuEbamQEdg+5jL2TtA73F0I3rI3
+vkVpD31bzGR5XP74/bhnWZwc9lzaJedMjOgv4ChtUy86wtxsTOgTJC0WgjBlLy6
YNVlYsZCqtjONbdsSAYTJ42khdXfB0qarbqry6ekhC5gJZQd65kacfzky/uGe7ie
63xvQagnUvzTbg90mO6KKtsmamTNZTHy/0dXoPqxnvIwwSbYQN/4v41nYR4Z/aa2
buaMU8h4yLZ4pHIxGvBkVWLfCIP3We+ss4stoRRVUzZPWTpnmhmJDF4B+6J+ulSn
B2JQfTK2gTq+L8Fy4nNkJUxfXbyyJ3B8mEqXX98uV+g4hvZeV6n5jtYiKy2KG0fe
3VFPqTBHYfmGlfEa9zyO+aiOSEo6SPK73OMPgfY84Q/DsNj61l9sSqufCCGA4rog
osK71EChNLu/iwFSnt7bHOJZKsm170JVkhCuuORQj9ax1/ndYq/jX41kqzua2msy
3Fk0QpQxmoZjyhHaUmerU1IUbj+nda90/N16XoB/oAK1E+L2wAeqdxp51Cb9AuKe
i93H1n7yJ17qtz5AiP+Sex46jk8ENqr0igVWG2wGKZrHGiKtNJNVUdJEWmg5v5e4
wmMtTdv9qjaLJz/gxMdMjdvmc0+ZLZzjtnlMJAr5TC/CymcGj4yVONcw6PAOsCcI
t0cxhUD6US9wg+hFtx3djvBw7OXzkpX5FlevAF5X5d2IuNtnN2TXYxNapF6fDALW
vrnt0lbA7I6+9/MlXkAYA3w/9ZB+KqNF9/UQI5/7cfb4tOJ4J18j6vuKbzxogSB0
rCHSAqRsuWsX+eERxQBXm5RH9p5JqZcFoSJ1Nb81CRExYKU1/x0ZdPpURK/RQgab
mDkef49/nwCqaGd0PB5FBxKeeAN+3cNuyxTv7Cwlu6PFswEcU+uVzI7ea9rdxCrO
ezsXcjiHFuJmjOUgvjuLU3OFKlDDXJvUqmp4PJrMQD5JRxjD0AU7ZCGIjR+JBkuS
sPWLXKRqEUk24TQNagShDZRQeW5uWI/82x+MneaaWgQu6nr/qRZ6mHkabP+HWe29
hAoT1BRT/VRH+kZVc3pRpeEdSxqhucDWFUmuykmYbMMFNzLsWMZdtgbHHXciy0+5
W3SDGKDjzdoDH55q9RuzjE4V0v9roxQ/uwByQZayxre5K7IOBtRxEbGbdgybu5Pk
eGmWSvr8pnLYGaf0gXqsihfFc9lSXVOeTMrS/wSJgvvDTNyaYnWpoGYtifOluI7k
pHiI44RypImSBwp0mEvmbF9tBDzYYk86YqGaPN+qfKotCUtmWILumX2JhjMufAaw
Ro8QGvMRJNJFG/qbNPd7dizCWvl84wfviPqGHv7bf+mdfM9rrEFWLFItmvuo0jai
h5iTbX4jGli7GKbhHR4SNhjzIEZk9AX0BDLBiiecDZRAiivZqNz8aUiKrIeFdAAS
m2+s+2wcWPWqw/FvLh5RtrP8OVHhnr5NvnoJhQJWVOeVu7Z+v1Uyng7Hp+0J9gP8
9Y29e3zcr/THMQlGatv8aDMMl3kE7Z2tHiOdubjxDnRkPFX/ZGvAza/CjLkKxihk
9iGyN/zSi2Jz8xK+fmWEVVNrGW8ETYc+iFlsVcnd0IcINp5PcI3X27n2cfsNMpU4
HVEq2viVqVk1zfgUFyIaU/NkaTDvKxnimzD1PJAh21t4ic7pEIP1Tzh8uLBcfbad
aEN+nWGvjTw1wSOcyXWVSuxsNqBtyFxl57Z1KTJ9/Hjz71w8tQC93vbO1LcLotaP
x4ZQfwbkfOv5+hAE3YuYGe4PRwAYkps9ywN0NQAiqu9l8FsBl/BYPIrMCJtCSp5H
1myPaDN4nLDhdC05DccRgsQIvWNCyZySQ9GC/hctkSc5yhMSWKgF77U/jBMM5HIZ
1HDWIblGvlPpG/Ad1FAzEiimH74KDgi8BhzEXDpQK7MwPdqdD7Y6A9hnDMPjdrEr
Khs/O1b20gSSYYLhzevOlUm27O7qd19gNLfSIwbH06lxy8JCoLkQQFQFCdklFv+U
7krH6cFN/ZiB7B3G/TaS/S7f23dmZzRhvuV3lguwVadp/n6SBarzhvLIJlUbsePf
qDHQI6n4d24woUaLpNj23IaEBhdWnItByatQE5Gw7LNtiM2m1pmiXctKuRZcxTgA
ctA+ogiXKBfp97qkYPuQ8K0SfHbL7kVjTrNs4xw3t+xtpwag0ZGmQaI5yNK/M7PW
t/LqulMn7b7R3W8i6xMBEQ4kWdy9lVgzgMxDjcOj6rPShyoOu2nNsYCq2ZCKm2tl
vxvm6dbqxznoYihQnnGBRTf4DQWH5AQlUGTrNv+nsjzLYXCC3jhde4hlDVUYP3Or
9b1prW8sIM+JmzmfCDEPR9tQdm77bgh4+aSMDqXgjQVXiS8hxJ7wZtFqp4FwaDDK
ewd7fP8YMbMjpOO4pqAgaeWMKqAs4No5wAJ+uenoXvKhvJuEfFJm4geK1QXRDpcP
zp+sM9Nfz5ypftWpbydJOMwVVw29Xtp0U8zIdgzfqzPcCAifsQoRbcahIlitUNUr
m6KPmiBsL3xHc2RrL8mGKjJD7+Hjq33msEJb11JOPXD9UdQLww0MDZ9EDCAhqmoj
rYZN+ixwUp8uILL6Lz0d1q+HvJrFO9a+3R3P4bsVTpU7MlqxVlyJDBhjtCYQOj7w
8Y3EaMQwdHNyCXi+Q6gp3PB0bWRhpNClrNtlUj7VPE8+1beKHD47Ny8zP8+WuIIk
SPpaKAdWdgJCYKFjwW0PPn6jpzUAs842miNxM9Eq0cCfgMBquwLqwNHSSa0IDxfs
7V+jJW2BUMtW/M5t7rcRE4yILwJuRMPDNW9uQNGCYF32npeOIRSdfjsjoluaosqt
54y3pwkvjQns/cGSpkmUlyItHl9ovXCw1yb9jHu5Pq4jNIn//4++eQMuLdf0Uq68
dCzGMQE9NGEyjayNXN1xngeAPN8Hz9+pE5C2A0jd/YJFNfB/aaL1Vo0LdTAdd8tX
J6Wp6wDIU987Dk6xaPH+4OYeJyupL37LDRuhuHmv4ei3LwXLV0BlifoAqAjnCJN1
yKlF8NflNEHAKdbiUp2r/rOgXeQFm7oBA5wsgy9hqDkcxJ29ehFFxJEZr8ta8vCt
5KUxEVvxjwu4wPXc1FMJT19exsQEivbf5oi4h1/fsSXoZmwAxA1JCyiffJzi1rv3
1FBpwYjIaEo67xIzPqu3LbMo13UbyuAq82Gbq/1YzXgE7+PCzHEBP1wvkPyYniaG
Ke6VeWo9kKLdSno6dYSx7oBQQ8Y3CsLP+czjxFox8ehhKF0qgaN89ogBQi9ykCYW
VIpihX9S9UT1v8ZJyaVo/1VX7zQV78i8+wOHXiXSSYGGtWKyy/svAsUZYvmcuKwg
s7kjVkVpFOKxefGlArjazdkBWJxWyFJaqF0/oqAEy0mrkbijcROzGxtG4PLSuKRn
kV0BoTuNoC9vsxbt0+vOR+Z9FkxXHNGj27mZcAyZDQrumfDY5k2l+3RwnXLjpuA5
esbj5keUGr/a1CWTCZyTVYChOE723vXbJATokTrtrgUIgjFxJHFzIi0J6YHs7UZk
f120FE1+nFfMwsIk4NJ/7fWcRB/Qgu8ARMEa4yGeavqiubOnpgR12V3mu8QIs07M
BJdEvnHdL542AHPeyclzGL8pzzzZAQCPrTiYbQhAsgE4y749pLcPF/JnjuyuwAm2
jdNdHbQBIec7UlXHpz0X9iz3immAGiuN5zF0RDNaJPU99YKfp9O83cNEaIufjb4S
x3BHCEcaZGbwtqU9xcKZInsibzGYhp+VQPs/LTx0Bt9YeeadFM4PnEaSKFa1/JmR
qJ2E7saX57TBiiSSKxXaJ4yUWL186CFLEji+zIxAuIXb4ZAgWoTfKhlKx3ffaLTI
tO6c8+p3psj/RZNNeYn5z2KAbTuEDtx2hh1Spo55mGUzmdqVA0vh+OKqd/SotDAy
hU5ZGKXlqGVJwR2RpY4mE6wIyED3XrnoNt1uon43EExhMXhSx2ar9SU0BuyKOMjo
guLHCdkTndnFPS+Mc01yacLPZKCfCJLVhhFXfWb3X15/d3p0jFI/M9dcgnSq+e2n
icewiCnFb5qWJQe+9p02xypODwOYgFMPzKx5ttHEWzwqZ9ih+4wSMp4tq7IKjn9V
Qp+0V5zvmL7FK7aHYnlpKGeYJJFzPCi4sf1nyuaHRkzHlA4MPlqYH9mREq9jKuan
CO4FEQ6qZUqxf0GfoNfeZsdyXdSpEwsc5jnS343biNynw4+VsQYMTLpAI2KX1EeH
mGf3E4OLeQW1kM598yBUCg8sDOxLrEer8dW7ESec+pE0GRQ0Dgk+J1IcdIQ/vyyN
FIG1yukf71Ihpof1FDi1cyYT4NeALE5l1Ui35dOvoO4gqVbS9Gd6y6cNFXjxzV+Z
yfLEoDGSc5l5GKyg8QMGvDK7TLq/bmM2Fd1Up/9WKSTgoYj3aAsxpTeg5m2DA4wd
2VlREUFUNPRcfBgdvG6wuDS4EP+aJM42a6nhX+4X0a+zuIbXVhSv47ONTQ1VXj+f
+wfnztnRp79z3R+b2fcmHQKa6UxMBOxH6oPyi5vm4nYQiH5nL+yH7AJVAFoLOL9b
EZ12WXB5YCYMRagJ1JCFmOkE0L+N/UbIv8gsVTfAZYhHnQ2q3RgSMSWV2bLk/4Hm
t/p22aVMPGa7IwjoHt+NFT2xP9tTICEg+0MfzC4bYtXIzjxLZwqoTCSPiXogWIx2
wi2XDYUaGNiBF5+fqdp+1YxVZ9ZSkJy1tOd9oIBFe99bKy713cciThdUYi+50n2Q
sZ3+yyS8vVz15vYYqB261EJo49lrcijljHbJTdfvEHv1kkVp10GQXBj5swk9fAX2
jE37+KhAWQCgpyLTREOUzMslg/+nDDDwjrnu+OiImwS+RUXEWcRh0cYBQv48HTfS
9d498f9oz3tqjmABlaL3zi2lJg2EnMTdmhBZHHiblSOjskY61AWD6mqYxHpBDQIW
6S7D3Vg1aLqNH3pY7I3UExqRRiBf6gKuofpkkc7FYn5qtQgugeHRlGTZuEbXDMln
xE21eZ7zr3xw4jJaR4FW/fd5PzepS4yIUWrwLLcnY5MTtqpuGmtYaFRcM5Sx01jk
aP6fuk+LnxtviPGAQGas/AqEZ9P04FLMqiHX9VditvApylwrbGCILzEcwsA1/TaB
vTOLLGarkDUokrMcOmlUezwNHHdesehDSg7NiWUE8vznTt+LQmv+I3msWwRJOktM
uX+YB2X4sEM2gI9TFdIEenMXdIav+1Gggso44uTjF3JtEehvWIXKuk9zdmnq2Q46
akGyl0lOlh3Tpk6nuB0IgLjOLOOBKr3RcqDc18sf6F0dReZPqtOvlNHf97opB63j
cjuRolXcmkPEf+APO1PwFf46VpixijqjQ+a/AygKHMJAQgT5g66qNexSX1ELrF+a
LgoaDzkkYhm0fwc+hWbbq0s99niWQ6at4qgxwMkKDirpYH/8nnnEvMtyaYZJPcAY
882Rmh9r51a15kUXEWbOVauMntzKB2cNZI2zsN+eoi4u8V0/eaXPtKPib1USJqyn
ag7Ycu+dcI5fnOv/zqFxE5Yxizd3MAtYs6+OXUsGpkqIvUa8PiPZxCtYMltgQbPD
eFrJ7+7uWwVSJHOOM71GJ60Z2HSTSuXiIOSj6Ke8zY9ns65y/K0pe2hBkEsIIGJv
WbqS4rONL+KDHnzG8ycERnFZ4nsh1sRwdOLBesvH8QpUTo7NSQw0KETf4YkKUO4O
u1eHlPyZpLb9XnbNnEn+AH03rKWi0f+oc3zUTYlGjKXlfHPqYaYsxUoLbe0KY6t7
yL//S4M3uMxswe6iCIj9ziMtL5KmUFg/+xHBE4r5gLvzNM9Syf79QpgF1ZbYis95
k0CrVUDVy9V5EwFiwO4/Akv/uikbddN5twFWxEprgYkLGfxeJqYkfDNogkkHdS2c
3TXDxvrS3BxmqMBs8qtO6L7lpkx/6GRq5LQORzxbDmP9zgj3rgN7T7bDs5cA/PXk
Tk3HeDAJ37ZdSyGIEhccYbMXRJ8JYHQaw5dfwA6Vkrinvt845Sq9zIXaLi6EHB9r
z6k1GYX1HUWox8mQ/mQIfMJA3/CGPJJ9+9cTILpjEV3J51P/4WrZ6Urf+6f8BbdZ
VcfcAMX3C67kfrcuKvWnLZ7cbplDsCYnO9sH6q7K4Jqvj1wwNkL75+Wl0EJoVODw
mdESwZBT/7Mtt+sb4cXw8AMCAkMllhrSni+JtuvBgBC2kyXyXAGVLEB8ubdxxkWQ
+/qSvDyVSHLR78jckr/QdAw9/ksuGyegkT8/nuZDedGlgx8JwzA4nIoxjV81qckO
hao5dAxFANbcMA6JEgqIvTmr0EZDQEqljrBl0Nrh0OsuialMUKasfH0CzTB1KD3A
yycsieT9smXlTQsRnZ0CHKdgvnRHSoH3TyCHPkTbC0PbJs1cUNBr1Cd3Ux6y59cD
BQKI5Eh9YCO7NAD/7Q3yupYYX0TWfcmMf1qMzHNILVUltSfO8G0TgHf/a015f1hx
4ltNj4jhMMQsENe6y85hXnzMjCWwDyL6VyMyOw6bt2dZ6tSKkhdE14T0Q8Yv862a
gFH0psmO5kOGBi7imEd7XZFN+Q+9yZT+C7t6vhWdTKjyM6o7mTSQOIADPm8Z4a1M
fgv+yUBVVOsdVeGs6Zgn/Zr5NWCyeVQlcGxKW/eAnyYTHBlGu6klR+gs14YvsGZ3
aQehfW99GyffUkHgu0o8ARTMIZ2nwls+whmsgT0kThHygtOdWnZIOpfclWOH3xJ1
9JquWVg9fOLAlOjhc8r92+XVnd2E8fT0PBRhUXjtfoCKiGwwxOUEV+6OmIM+Ui8a
NTS6n/MtLHTMYliTFxOedZbYrWULKzDK41rKwIdAVBG7A8pPkaatRT/2JYKjB6G2
3u22RJjTINLAwp4RfZ1k35k6FXC0lavw2y0+tTFszkMWp9XvmyIqcjg5ShpCEzMv
OunvZjReqwGM1wk+dwJOT9umXCl/rxIMkmgJ8UydjrIZ8Bak5DnYjHj/E9UCy6Tr
nbA+F1TjxcHGqGExd1u0j+E8OpoK+uyU1FMmy1F0iuDRDue6/FdI2qyuPhFeptCO
MF2ynADSF50OVOHcK3rELro7tvNTPrU9JVwprLWgcPM5n/Qnk8fdyFChUKVF9M6j
MOnY+84bfNVxjsGqlBRT3zIH1AReEGc2S6EJfu8QteV75jOwrR1sYCOsrwr1pXZV
JnyjbIrWtta+GtGvpWm6SrgTZqgUN0+pFg3FrYOMx2nm+GVf9FES1BkzdoPb1xis
inbjBmzgESBKfZF1+rGefxmMk6lEIvYaMsxVva0eP0m/13y0BDfEtuRxeI++H9BZ
7hp0BiT+SC+3fVO377WpBXw6R5oqHxzXz/s3eZYOnkKEuLFMTBZop6QFVDeGjEcC
cVuKHO0C4Auv8utoacoAZaW8mDFMXnRW146lgjoEWC4HQG7r/xl4stpPSmplyviL
ey85fNy9bZl29XfzKYgUms0rNuaY2YdoHcTeFJ5nSjWkl1Dxzj/K07q4eNoI451C
ZWdjA9hDwoBxfk7SmxuvQ34JDuBM2zVqjgXZIUIF5ECesrh9Akimze58jY3h1QvS
pNlxR1BaeiiUGaSTUvEGvHdEmUDjdNdm/FDC/hz9cs/6OJbDx+QCe0QUVwrBDuHT
D7gQHnLAZzhX8hWx4NThdb4UeeevcbDmm8ta2ifI1kaRQYEkwVbXSKK8b8zC+cQj
b+7aJd5IbT8i+UP3h2Gp2Mbcwd5OJUdbBqG22bBQ1nuJHoMptAFRbD8ZTQUxElSZ
MO3eYu4pCQYSWHs9195BshudpvLQ2ZrBcQWzQY0azp9d8q7fNTePIIRUQEvDBVnz
6i7HAbCZl9oVDRnIRLiEszDQKbPABIUR3LoAnPKYLL+R29J34iiuDLXZl5PaqRoB
iVh8aCO8PJKlyK7ovDtoWJXAM9LBlCgVGLEWGZHTbYRVIB1D/G2UAITJyPt30b2i
YU4wpUMyaSCfcgqeIrdnNBcJAZK/YS6P/Yv4TaMS5iAcC6k4OuwQfqyeK7kL14bu
1oo9EHylwoCocA+48U3APFqaRsLdqENuZtgoz7JQhKMMCoaWVXAtYOu33qz0m0UO
GkxTfP/+mdASat3OTwz7OSkYfJ7vyjsYlLE092H22LgXE3iLEwqRy5TY3ZbUHdxF
E5yWb2CHzxRwnfhuhPUlgVdu1yaUjZLuG5hmXxOiwjYmXgGkz7aYbPdTNPCoKP+T
WZOEN0Nq9n/wXYmGkGU7+qO6rKte6RaIrjTTbjbG6JnOSJvkhVpFx8CoXTDHI72v
azdaHl4L4IdXWmA7RvKOxfx/RQ7y4g2oHeVvE3iSl4e3WA7Q9yKgrHlLlhC9zNjd
91r4ar0+Zr2o88idf3WKwLCEKuFpneE8D1K+Hrx9DGNXBFOUJc1Uac8YxDDC6b6S
PFjBdvcV/qbfHeSH9l9+7OWuEdvebeXs6NTqThRQ8Tuq6GmWzndQpAT9kr9P6ro2
5BavpXvwTMPu7jawxzJBPE/v5j9dgN+xH9tArd+NKZJuTA/57aRnv52AJHra/Fff
0DApI6AydJz4CRWD7xQCdlhsvz18H4ftyj13U9N6lC9wdQpQRei34819FM0QrB2W
AhcQ1KFYlpOcHirXYt1GcsYvUBDrN1nPSV9/BNQitul5qoHvXQ4u4urDUAw8aBlX
GjFN8MKzwbVAgnew9pKKG7zjfNP/ApGN9qZxqb20jk9vW6fV5Gr/S1ZdWqsuFdwH
nMNRmOyplDHGrZ/49lRHaMZx20H0nWkwTnVaQkFhCXo2ZhqwlcsHsl1iaHKP31/k
K8RGpjYF3J1K+QslHfEfSOy6qdBNq/Ar/ShHmAKJmkPsuGFfg8MLc0cgOeIiPaPQ
or1h1RKBw55Scw6mzF0S2z+wqebsqCuyFlCVH4epLkodsCOT1EAalkAYdx0ODPm5
vCdaKbZhyNFC0uvTKrNdkPmh4Zl80HLM3L1NSBXe2VlFJLQgeAXoOkdWbmnzD+Nr
OPU9BfmUOWJ7kA/VlzdL618VUb9yzLRBTjZtZX6EKvaR2oSU6FByTtHZA6w4llMF
kiz8iwlST69cwdahm/h/OOL2mSVidVAAXN8eKbZNzpmx9kBbgXaQ/aevlMxFZMNT
QoSHnFkBVZ7G/3MfUKOZZ2aURZB4SvwwypahYC0ahJHgMAoBzdtCV4mh5Y9LcGas
2EG4rKcCqBVmZgmTnIEirhdZg7pF9XtLC8oBuAL/UTxq2z+DkMImlmDwalYZXE1G
0uYyFgUtrNah5rSSvf/qd2GQFYsWkUNwJOgb6PVuAqaXo416UI+tNAVjJ2pibtag
nYbF9FIBU5SUj84lyF+1uxwbrUJNOCEJTe6WLhO7Fx3M0qZSkHc26p2/8o7HfIIN
4drs39gFW1bhYB0AqR69RuraWsxMYjrwnN17T0ar4vktBv8qpc3iIGcDbcwnczAm
ArU10NprVk/ozGDStX7yd3F7FBovfr0VFTZ9NEknrifeD7D9bkceZCvzsUS3Pmxv
c26e+MZA0fgVNAQiCwY8rcldtXH0rCceR1TbYtd2pvsVS6SjvtS7BY5SMEVRxCyc
uCqy7ZvFL3vT7LTwfplnhC9oNzVAt7iZRwGuzNM05gTMw59+S/QwMHKrwE+WDhK1
PnNykR50D2q9OZSYH9/RFZ2dq0o4cX4UFcYYNTJetP4nWhAKRQfxs+x9hUHdG5c0
oYr+++BIyUOOQQccpRZBbew7ENWZkhbmhq5z/DYBKMf4EAIf3GDU8n1RHMtNtkf2
7/fC1acPXGBLmJmfpBNk04MqAYhXewTAit3yUh3ysueMD8JuzDv1t79FKQS6yu5R
0cJr6ivNbirsFYAabj4VxRTJPzGBa1fHTaFq8fNqLmlGhC+E/vxYER0/l46xzNrp
JhBRya0y8joSJVkdDSK+iE5J0otxhmwATfDV8Xrp4MbEhEgF9Uu8S9PmjF0L/MJY
Fs9bi6hY+w63jn61rj2NPPHM3eip89zLuBX9T5iMMoqWx/1V0oCCJz5ecya1tFIl
k0NrZ89Zu1TQChw1ncAFUDKKR5/5//o2sSuu+FW+tEo1kJt133bKTn6rVqJz4LCj
UKNSqSwvJzFXP6LtHpUGIYBMfQWBpVhv8QcuK/Gew8ocwOkWPzZPkxMDpoMTSaIf
27Cab1FwNjVKsr6GgSGqc8U+DQagwAmwKOzcN8K7Fv8HELwqqMaewAh/xZcgw8UU
yJ1gcEmpQGhVkFhZjmgvovAccidFon1Fr1vsh46IKYEEcnuXD87MmSk2iD7KpuaH
XAQqCIHilNEWYBqhLAqavjtz3QpsPU/1CtjMG59V60PU7rFLOdXL63bpJW5fBmTi
09GKee6tKHANELcG6hU4grn3dCNGZcxTPhF1kaoY8aspdv1alLi91SCzalMFDBEt
nlOrs6To82UI5y1bXgoXteWt1q4TxkMTz+/W5ywGdp7/u5CimKj4KB0d4Wb3N4sU
UTqsMRG6G3G0Tgy3/DladzuSVB2k1b7SLAC6zEhvz/RXHntMSCNGQk2Q1VXOHMwf
w6PxBQB07iuKCcHjIDsX09pg+bsVSTCfduPuwwCpiwFeedsmBPxNI4lcb4GsXYPj
DFYYbCKKyTdHViiDQIGX91jgxna/XYfhMqrtM9qSr+X+ZnsPUm5w+N2z9vaKOim1
M70XypHovDzWZjVFGmS7fBp8LjifvZZkTqn69X7+xGhxtGov8mnhPao/yL/5VYZa
sAMR2EBUeNHVR88Fae77dkmw4CvXZS/no2hm26McBmpzMeQsDN2LiGqSqTlRA6fl
Yp1ZWJk+oIfOHTx+XGjgRUzPDd5W4X+0vwb+Ua3ZxiWZsiYrqEh2+WmQaDdZP0yP
7EsfYTM3jG/LKVOWrD75pRG1aKzPCJ/N/IVSosoQsDxZxF/9DGN0yj03lr3BjP9j
ywAZK5JIG7gGpL1JBFZserhHcEP4wLjabKD/EQMKMFt523vxEah3b3to5C+OoF+K
xnw81oHr7E9ACChdctKw93AaH2ghGnF/EfOJ7Or7DlC6YzeeBZT/bNEdoAfRY8WU
GXpyxg/NN1riBtqAQAQFql5gh8zhiETFzyZlHN6VVjxGFNlIYIw5Uu4N6D4xj5/X
gH4jj7molJZvC0XJk2FLJafMajloOc66dC03jJwvX0/REFkHspJCkABRx9cKYNPo
xjvkhusa4kG03IQpuyunVwu65+NObD1PZ1kghckM+y2Bf/itr0D0KdDVmlfBcLHj
dKI1atlmQJ8ma8LTetVIg9G/RbnsyJUIqZhbsBy2oQC4PDokhrwxQaAX9aWtuih+
koniyzPweWOyw3ulWp6/bso/wLYJ555kM/i5nwcp0Uw99bo/8iGVT9IIjM8bBRY9
nj7w+H1om6iRwLABtA4KxAR4JPIqgG37fCAjLg6OvJxvOPcs5TjJpv7NwiuWAxo8
KlNhuxM/Tx32Y68HPZocxWOZNkK/uD4T5Y/kE3dZd8W2XA37kb1ftjKkR1nRDB47
MU/UF2/vRyRxqABX/qBJj4I5IONQsJXLlZuSmnT3BOelysf3Te77CUO3Ex05PhWa
ZWEIV68fK4CTK8/EdLERG4kDYBEv5FWnzyrcjUzEsy5dX+wpb/WqjbXTlVuDLqf+
cqwp+OgQxR3e5ptJkCrAy2UPRzTVc6cM54jIRCPfgtv0I7j7tgo2ToaOgbyeBiE2
N9pKoUhqaVH2fAzoTwZHeFRox3JeU+2jV0dIJe8psEstoG4nM8DdLudsbHrNovHW
L8VuWFSjFt4PvWGBB9HdR/rC/itw4OPA7Y8ghQxOhKb0y1ikjnfkSJ0FmdVaf38J
lS0RvVHf2W9RJzBRie5RMqRjXSf+UUUToVyrCJTpKC9u5SViQt5OPw2ttFf5wP2L
5FxWWSu8Do8dtLHjJ9XCvmKV6fX3XZc1SZgJykQyWOqHayL6CPSSafrVtpLHQKhy
C83VjraSs1faE61NA41SIHxP9A0Kc5pKjh+DzEi+JKpNuxMcLNte7rR441pzQx16
CG76i+2HnlgrWRpIgoidZtxiBxAEXwNXH7f5KjtfK7a8zQCAmSZ6EdvDMpmzR3r8
vVwB8NNGl9qNI0TqnXyth1vwT85cwaYwKVeTSHTC1RX8vw1HgF/R66FxDHY1KyB6
KArSl52k4BNYpN+oJQ0qhtdJN2t3VeTld/r1Keope37F47bY9xiOQcdMKOvMb7s1
+0t7A875oNmi55KllGuUSHq5i35O2JbND8tkOuEohJV6Id2qHVjia97ftBgZLZZ0
+spPMd0yGTNLrNmCysK+46vDFLXJNWWgAQ2KMYnzw+AOzvZCs/CBC/Mo6w6R1kcp
VAgbVfn99Ui0dasFlscAAy3N5zi3mFc3uIadcARR/pseOJTiGAaSHP51klsveYQG
hEqb1+uMWVRAXp49A3t/j3CMwfZQmXyvsTqCv3Rum3cToCla6q6kj8uBOnaoOtB+
IgLfmRSwZi/MJB5GkJhukb0N+tjOGFQuAh45ZbksE2ROfa7TQ6+srbph260/uQXl
71D9EyZc9sTgDrbZMbMSMv3dye4FZ1+Kz7ixkIbRXtIzkLofPhY85x7EB4JqIR8S
fXHDeXArKkDzDSzH9FAy9Tk0PX5YwGHJOiEwl2pMRDXfIJWxAiKqiTxDd9k0G3zC
610wUUbuLeW2yBNbSuYYdmS0ZgqEcZcOgrFQgOceThIp9x6Cx4/P6WmqyNygYS+q
2FRVnnyZJn3eAIquVNQqxcQoeier1huW5i/fDwD5mTwkXg6VEpQGog90oakdkta7
hkd9PaxMCFbgmcDjhJ4jimw5xMW5XSXQkIuegFp5vfU4CR9CLHwzUYSjz+a89D1c
/buzRk/2NdCGAeWBSb85zyXqqh/WCo6xXl++WYf0AHO8l2JHqpHdGVCOi+YX3CoN
+TKIuFY5KlTEc3gWtW2qhm/B5mk4f3Yu2kBSRr3EqpFl38S42k43ZnuPs4wl8Krt
AAIrLoAVti9B4dtfQyTJVxwevCOSZNsRxLfXoX+nu4UN7HDqy8zlhlSkTNGIIgkD
vdTd6/jR0AIradd/C/HziD9jjNCisARTlledVl0CkIKYSLE8V+k6iWdL4X1pxm91
9UX2yOwn+uGKV9K9848sM4bepjqglDpwhYOZOWP1ib+Zv0bdV3ymy5/4mi8wYv0z
40wtXR8V974vXCFMLjmE7I+pwhnuojQMuOKtJqUmzpWYB221sWhzdNG+SnJt2R3z
XN8NYoGiO4Mhvld+yJ/2z6Gz7GI4Na54y5dznAmvGt29A6H1oI8RQ4zkolIbQPf6
FazKXaqc+cSEnbBP3vZ1SLC95DVsRVovTl5GWaShHfou4hrx3fGgohdcx9zfIOan
h77UGSjtoe9z6k5ISuHpBg6ZdnQxogdpTG1NVLSJH3h7JiHIi/gU6BidrmHZ42Di
t7g7oK4Oys44wE6SrF3kclBO2yFXwChyqZohQBfRWegt+OL44Qj0UbVCAoepZHsB
ThkElztFCZzQeZhGTls2/6Jhhgs9hNZ6Sq9AiOmqWQTqfS2xMBtnNCjvkEAy9LiK
+o4c4KRWikDu8NB8B/NQBBrfOQy5/fUsd6u2H4I2kU7EYLhU5xa8lz3Wynz823K6
MTnQ6n+XNgWjtfpc1lSfdYEMl4B0yr9ceQnL9oI2bWTa/c6vb0b+UsSuv9q+e3Yh
5vTejsvewbtmoOaS9JSTjqCZJEx2RtriAKVsukaE9K2ToB2PR/zNgBIAg7uOsUEV
fGyLrJNAic7MP5mCk837iNS9qK/fMZMyB6SqCDhTLWqaCJfmIRsRcakbZ8b0VIWL
L2FYXJOG4uzcH53szm3RMgaSLZURpbcFVWdFIyWBknbkOIb23x6LqjiRhGCyjyI2
5jd7a4WVV3cVjezB7r3NJvDKl+2OSEevcGK1CCRT70GQhaD5WqMptH9DVOfkhLkr
8r15tVuSA9jv+wGsoZ0COPAcENZJI9kjMCChlssrqjXSFa2SN3T67eKhFpWYWVHq
FD8Kf6ygX7t44ZwVIY+ctk9ZFHc93y8n5HwRqJQSlViYiWkyM7Nadfc5JEwq5dqY
9muwoJQV69693LuL6dLs1S8/J08P8BtK3AUcOWfx0UJcyae0YqnUYJsUMNGjB+pS
ubIfiGnjCwuTRRkOwauR7oOEjYP7iufqQV4HYLDQDRRXqgzidzA6rEE8/y0BaQaF
VqwzhbNHOYISkbbTPAR1x1hoq6PqQb2YJH4UKULbSfcu7NmazKcGrlUqiMQQmW3z
yOa2MexXK0s6O9GQAy74ye6ikGVF+KhUrU+2/mQefcTCuYCYo88s5syXLl2ufrlL
Mm2hor3FtUIj+EpGQ6o93Q4WKWowkqAWGKvpNv2KSnDR9aIfL3IuJbk5pUtm9Ga8
SNgv6CJPoCU6y2K5NmQzf3iUfiPgOzuVWVdCK2C7ST5XLCF8ZnnPqV9lFDbvWpAO
Fu8Jr4SXz4HL9PNoazVlcVOOUp/dsQwvBvQU+fGe7DwiOZF0bEuDU6gI9M3qVT9Y
+t9y7jahkI2hcxJfzfDenjVqldhwuD2LSwOYPFvOfMMPAUMRByEUaemAP+QkaVLq
CpFxufgNbI9m15XTqLYbAQRwSWXy24kOxjIXUU0u+/mGRMIKHDj6NGkW27Ek3jCp
a8S/VH+i2hmGvTdnPWu2pMTsWbmQy+wKASgQOf2rZdpK16Ak6H/3BULq42TR7IiB
tsuJdaYPUgCcILyiDe24Y3A8uNnmtAPk/B6YjHp5JF9WzlHV4puFDIEbuaUOqhgc
+qQHl8qx/0ugkxokQ/JHVr3hKZFx9d1JN5dZSndCy+abM6uo/fF6yi0QInbIa/dD
11+nKR1ZXSbsZSSAIK8o1hTcQ91dpjuEiX9Qy9QA/OkJEyOFinco1j5hXBhCgKrP
8QxrDYkKGubUUHhv7gFU8vUrt/ZZlWb9olYXK1ZPwzn7OyTgE5Gm1+QlOrY0Qryc
S3V24cjXND4vIb7hzecwY/Btth++peFtNZKBmGmfY4Nveglcfj03P9MqmsCVFBcj
pUm+qio3jLqoPgPNCRP21F6TuaC2zn6QMgotwdQmBy0FDDZlaIB3Xrj3zecnWq3R
QCxSGnxGpmvXGCOhSKIDo22CDJhV8LSbcL4anHhk+NMv71yxhpFd/PL0ZOmBbjen
JVeLObE2MgodebuI1/HxLqHlLjiCg8/frUqrsqZKRdoIvVMiYYZCdM0K4sy3pb3n
VJSbXroel6k7vmlNZvi3dC1FcDzcqz8Mb2DTCS1LP0Jw5eaufMvH6uQI7MvZCeBo
zhUlC2vGqqhPeGBqETxj139jNP/rUzH9pJrHtjVV3R8Yq1NqCwrvYKm3Kol3s0PA
CXCcrNm0o+GXLI81UsrZR27tecIHG4cxbhrySkcofssODkFjyx4DJhFbDGYLVToj
9rKuVJRwTEecddP/TLnonplJ42/OQpDKTvu7bvOpGDMggTD3x7nM3My289xlZSkW
x7bEPsfjthZmUxNxm1CaTNMpSuiQbF2wr7w4kfLWXXwVZH/Py8/lB1inqwnPO4WD
YdfW60wkib4mpyxujlRRuAUshyxiZUGIpcesuwwSpXw9uru0ve+3Sp2OLaB/ZAnu
ep/Uq9z1yd1UeHJ9o7TATq/JNTwC4d0QJfHEMKpbUVZ7OSYP2Zo/g5RrCBq4FeqW
2cih9j/dWbHnj3T2mXYT/5/n5MbVawUOESrvZ+BW12MwKyoqSDIyv4SCJPFHlwUs
oHbVonc2r6jO2KWU1Tn+6SI/R8APQKD7azZ6XwghF+jMl9EMH0KH0N6ZxzyhcvfG
E5GdnZd0fgW+Q/1og8h7Zof08l+E68V8Aii//il/j6bZIs3Wr2Ouf3dw33k5//uN
U99UbvvAOKVlxWpxyA4IrlwA+9eXfbsxW4fkLH/VtF9qw03W+PCimtIBhM4h6++G
stp87hF6CrwmoXoa6uJeRNJUs9EaTbIwZq5WaF3sdqQ3HyCMQpl7cruyMwUE884z
WAQ5s6lvQ3sOIBfYTKaP880USMb63XKgtVyXdwaczCgu0kBzUx5dl+Jxzcb5hz5e
6TE80dAkTep2sEi3CFN2hEtuYnQ2aqVsI6JyrqFLcqSFebpOjfCTcsWWxw7uHWKM
PknErofdxYECsoZ5GYSjRS6SQBVeHBFM8dEtlUUqyteW36LWBVXi8UoEva9R7yxI
CKxjRMuiIz7CiEr2HbrYewxV00X1vHo7zOiAv4rEGcLhZ4Qw4sIjFLEbQOSd/64b
B35DSL9SjEJNU34LtBcMz6unOMXnK+ZxP+ZKeou96N/bKYuF1ZK+uRX+Y1JPAmFt
7Aq6dFj5fsOGMP5KXC1JsYu5iuPvi0d5UnL73BHvUbWZwu/eRbBr1F+B2Ld5Ko+d
+gir51Ziz9U+U7hKcQlKpWB4zMVWi98DS7TfOt1Vb9tR079FgFCS1w3TMALjmqcC
Ewg62Q1GmtAo7fhTzWolwBQEjUmYVKTux1TG47K6BliGIScxCO0YprVqcI0sQCcR
VToa7AJXtpH7YVx9kgjb1Oetom/nbnU0je7rqAwV6fDMQJT1PMHjpQQ69JUMBKe0
fFV6YjN2/lCQfvAk8pYRaI5PVawSJlIUpLQZMnJgmZxUMfHkV+82/zhWhv7/M7tI
7mzajaE/NvMMGjGN5l2koEmpmt0+qgvex72IetT24hjJJ521qozaUb2xq+WE88Tn
LMa5B4hGJ3VG+LG5GpiWNNPB9HsFxC5fzkzfkQTTrFNhA02arveZY0CdYoyk0xDY
SCRBf0huQr5V4EkJG1ajx3yY/k5k4b3/cxnzRsYXzTPkY2AjbhPcm7uV7DYOwBuP
ZF4Rqaj+lB7DS4/Z/8WN4ER3xe0DEUZbHN57D6UhfKm2D1W7c1Xp1oFQWX/TRFv7
TRMOx61phA7M3zqOLkb3M1q/iNX++mvXw+cRwU+lyHMYikTyRxBxPg+XifUNGl7c
GhFbfRA80eN9TG+hLN1WXKHWZP5TXHGw8PtV6pGudt/KDQCj7JUeGvbGUmpQZaGJ
X0JzQZkIgveOvYLbISIc/5GLnhmQaPxBb6hKFzCiHcURqiIywfOJe5GyHRDfdk70
N5Q1oQCFV3JA5fRVDHSasdpfEZDtsJdBeP1H9rx7fV9m1IiBK5kRFJbMFgmMA74N
gpswEJdaI8udCni3WFuRM5R8XzM0L9KdMumQ8mK+zFL2XuYRJzYXnlzCjVl60FGf
urgnYO8c46GKYj3sLO33cwYydENd0RQFEtp2kosmauiQqRUiWarQhosqhRtf0bcB
RWyrceTPAxMcfxWGOzEYWomRQ37QjOO6gChGUHqcCx3qzuupfgxW9nIbCeXyY/G4
u98LM5oYOwZqSLXvnOJZ1GnJHsbPPqFi4+iKxSXrljk5spyO+tlbs7I82gaxlYNU
88cstpH6M4iHJ66s4M2x06Rd4TdXKgNKwPeY1mF891byeMsVf18GuYDqlLCvSAlb
mpgr5lyurGEn16Fludh8Pxhy9q3gTgs3wraWz85WK4QSpg1gP3ksXKoNNcR2dxC3
vvJkbZ02zeBcEbisLa0C1Rd5aNAR7FEfE4TdRb4V0234MhPL+ueocMXfzhX79HDu
rSl2+EBaqIlwMwv1bgL+vLyNGC6xqs4jc4XEDqAX97n7u6tFDO9VsftcPW2yfZUw
abHyaFLHW9LL/61Pksf/7UyW79+w8mzNHffZ0yiN6g2+gCOYk1OnKhxQ5GR/5WdD
aGjHS5KLj7Cdty9qYsABMVqPJVjiLVpb+VRVOhCxuSftfs+qoZA40Ms9zwihzYgG
sfUXA8nzbbcmP5TpMUmmy00OQ2ww8IRqQVZ9/s7LDfP8yfrkAtQZF5WhBtyEbhFV
dSJ4ovjRb3IG5cP/o7mfv5yRBhx24sH+thrVA19e+bVlzaDmdDXedlT34IxwnjH4
sdfSJqE1N/BaKTHNbURQ5tkwYZ2Eo5/PQn7Noeq8UwZfkLY0/RB+rIbm1sFcWHV+
sdjMw2+JozE45jnVMn9is01GfD49Rhi8y7me3BtFbiH5ZV4jwMy/F83dklAMuf4m
1jBxFblTHFhPKS1azarxTzRCRTNg9qwpNd9VaGOZgvuw3oDGdbEwyKiGuHHKKyLg
tsEkc1/6V6IXrl+dyPpnNN8sPULKWtbIHjapXbcTryxn0L73US+HqHPaaDvOQeZO
c39Mx9KVZt9YcRlN1cZcsLSW7wdHUl1gkj+dziOspFJuFE3DGyXrVaMW0P2m7gbn
esWS5nmTwjAKuig4reWYnQ31exB7WHJSaDRdL8IetfzWH5wdzd7DgfN5f1Pzdb4J
58/rS/z3jeHehxI/V+PA+uU8eZXGeYTlkHiAMEOGTam73uwWNxCw2OV4fhyzBbQO
IGw/N+EVTYRcjx4GqESDhCLDxFEvD+mZFfWcN1/oLToq7U2Zinin58eNx1IboCta
9023GOkK+GahDUWKbhV/ynbSuY7qLaYTYKoQf18BDiIuZ/l1RexUkKTjb+KK5zYN
hoiXJsaq+GekwZMbWX4P89Cu+HirwKVvWsy35uQVaQOBXHCbWEqa+Uge2h5IElT4
N7IzvnDR5p4ycdDQ/xAdb7hFpF8j1xiy2aMvSK6+vDAP/PqH7OPHrml9/mMHfm9P
7XUNnbqNSD31+VbUIQEoLB0c0k2TFWMRhvXLdHQtiHwpzjUhYZuYusS71zfD+uOC
kPhEEVb0uLcqXT7f46WCMLL1+OsOOCoBebCrDjLenc5RMarkSFv7sg544DY3uD5U
Xt8k+bh7Fs/WZLR4YHluVy24LVgmv8/DvxfDojNao5wfqp3tW4XzwufJTk32EzZE
V+DGNF+aED/kpdb2hbiuo+TSVgFGU1OyR1qkwPxI7uEA2uT6IcHB+u9JRzz3US7D
/Hq8YEA61WwOyt4G6f6bpc7PsNugwrq1q9MtMvfSjc3kLhxI8Qh3L52zQwkoUMyh
QHwExcrSbSZ73FDbccxcDjeNh0hEXK2QVgLEzjdZMMxUkizGnBTHVIo6LY9AzerK
LPc54nol9L3K+5ezZazrTkxtVgPd02olASwSfO5FO56xJGEx/C/0TNvyzjiSQ9O6
yp2lzebIaQXLyAuC+7umUhcEwkTcAu/rsyfZPCLuunP8bJh0bwB92Gz88u32XE7K
YUbEeqJc9IW5tFXKuou6VTJR+7LNIWvvIhTYgZJVKcRoKEy8A1QNg/NOwdSHda9Y
/ytU7By+AZSrLudxkxbTIqdVx1kmEO0ihHgPHh2R9tsAitx+rmPyY81EvjvAfQgQ
2CvjYj1LOVKiwUQnBpcWmMS+k6Lx2GnnjFGmRRoH5LxELdO46Cv9tWFdZ7F9xHnd
tOgnYcHfoY4TOFv8AYS762kK1RVzhoFNQf55rV4T8Dgek3qF31zMKxE8XTg17lMi
J56CXa3R3if0BmUF1i6wuo2Scho3aDCYlBkNtB93B6+o7n3O+L6tfB1l7+dYJ/LQ
T/4n5HUGy4nbVymDUnK1c2z/WUuo5Mb2eDxM02OGaMP8605fs8vuOBCjEMemRZxq
JOmh2OOHhFl6v9sBknxAptijASFmPcKjiTGeg4VIE8GVwtgKHOHk0mGvpBFMM4VY
wR/xZF0cYvptPVU1kp5P8D6ei/di6uBX6F6P9bbKU6F+xFSmA+pdR8K6kWRKY0Xo
S8k2K7ftnCjcJ06oQUeOl97yq+2OuBxZ5pfkorR2Hp4N4sqleLRRQMk7pfrTStDb
u/bqJWEWNegvNVBXZuKHDcMf85GDbkeHYSI9UDvnzwqDqD2/yM1uT0ciigfEldgJ
IwfLmZESKQaT7dbeihRKECgSzZEuWQKBbdt4ObYrsHieohXVYRVi3ibPjZiyT9Mt
7oXDHzEIG5JRBI91uWWDQ2ZP+nZ2hSLZw0QK7GEeDSj8t4+XfgPuUShTdgwoL32K
gNOMSh4WwcU1fUVDZOGOMhxLVywp5lXQsELVIoL1CLYQ/sN6xl6kl5fSGPxMTi22
uvxxNvNIY2WwP87wWHA74o9apY0PIKn03EEg7ZTGyzKN2fVYm8CIobJtQ3NOVUEp
AnxDZFhV+3S/uEBrHgTBWZia95O4ZI7c05ff0FKZCS2IIM8uLsOgytPgWcEIengn
+8w+YOTy2dRRfc+oijlifNFWGrawv/59JUntBH3fhZZx7PpK6ngfRUUKuJNDHp4x
1hnR3VFWtJXEak0n/Ghx02pvgbCtFwJUOQhxkSiH9xYGdo+bPHeaS+mI31mvf+1f
UO1WXJgW2PJ7h5p1hwWDRlS1tmTZ6U3ON/pqnpF8rcfVOmgSNGjrRlWMc0obcV0Z
JtwVU894EZMTHiyggUOaVuFgrKEOQ6gBn4RYnYene1z0c43ATPhmF4Lwkluczkdk
e5DGU8qUNbKaCLMv5XDivqP3JNcA46CelKtySjmPUDCuF/ZXmWc0jOihYSJ4rJ/y
jx+OVo7l3nLVPQnmi7OeGu4nW+F6314wdBnBtx2C6c6RbOB17hlqc6jkPwEdccVS
IGNWLhkP30OvobFhlU4PLBB0ybMHNpFmBBfdEvEc/uhJGBz35VCsK7JTQsz+SvjM
J1+1hjbPXRx5SW6t6bGfZGYuLzHFFfZrHChUrvpUPjVg2Dez6hMkfF9QI9GF95u2
9qxwvgwjZZFO5KRpQHj+c1LI4bYLybG/CSglFILn/Qi+vmUsjF4f1C/nz9osFjF0
pJ7WydOBuExZaz2m7Oxclbm3HDQA10Uptsggj4lESvdrC+awp8MWveitDKvjzz51
yayL7+CDwsAUHsiLyiWnW1bpCrYzZVQ2b+WimbP+HxIWtGl8JGcn5Bk3G2SnrazL
RxfEZoElqJ0iaWb9JrLsIcHI/HIFffOOepKQ98fgT6kMRv3uJWxiVcU6WP43Dfz4
Lp0Jq03Dfh9UZ91q87tZhIBOx21/2CJFZESikJ3hRFUQxXz2s5Ek746tzTzVBqRD
9kvfFsZcINmFrh3I3KDWj7Jv1Ydd5KqUtFbMFcoiriHoKnQIgimSPCA+MhplBqYP
tSItozOMhRKAYrmwBxBwKuFpNog8nQOaGG0H7njLyB6rARoezyJR/EaqFkZvO/HK
2G9Y8XCJMsjeBi1FWMDcPu2K0Uw9c4POUdSkiuQ2dztd2lCQUIGpTy+9LSotbVVd
P9ECQLnsECEvtxfP9HL89OvBjTnRJXfpaHefyhDaBkXQAlKJuB4UC4GRHdpogl26
vS6OY4Yd1UfcTyGA5f17chQI1DTZDzdzVPszSHs+rBfAoeT6oFyDG1JbjOX3tMKt
nOrtb24I0RO7FxD/P/9rLmsLHaKXN4+lqrwgxroh/6KwIJMZCI9Q9em77ZNRAlNN
HQtNnJOXTH1RNDm3QoAC7fjFTHWRgO1Y0ky7t6vY6Gle4EOLdEd5Ywf2Ol6TTkSQ
yyKWs9zma75tuSfKvZns4R9zkQL7mbjimNlqz2zzCKzrqXxdVGmbJ7bQg+qHpx+3
qgvXISbuk3JTsPB+e4I24QwsOCey9ocDDCwm2BfxISeu7CmJNKLE/Rmspv/cDh2A
LwKYDs0AbO/iVPlMY8qgvndaocSRUx0yFH0dy0VMfH/fLVtZxZ8P7M/qfVyi7bx/
78aOnWWNGDvk1V97X8kCmb2a18N/EbqTAEWfjua3hiXKejJL8MEBKqmxft8i+ca2
wz5koAEHCCV5UuX0xAcIjwA6AxcPm4SZ+KSRIGkvjS9869aQRv/2WyagbIop4msZ
hygVwUjhRigxHh55XIefH5iWWpOi4M9smy7eIsDfdk7t2u/G06D3FHItbwBm572k
7QcPSElqAJjah7vJ1hAGaSIbKX19YokfD9A54M8ogyj2JcPghxcBPXS4ak8hrNCv
8xP4X9egXTC0dWWZT3ISP3Jjji+QI+FCe64HGvhAb4yWK7d97iS3WIUH0yuij9cy
evNSRFjtShnFzVIEf/faDNpiuDEf2lUg6YDLioCfHqimMd5TKia901MO4kjoznLv
Dl+mI3oFYM4DVNdtbpo6viwiEEJmooykBHrIXklLE7QHCCMCsqzO74uTeHtK2hOp
Zl6mlLnBbUf0UkbQNTuBilMaLMJWGCNX2bcZHpoWjQy3zaJ8iwPjztAX8/Q8p3ff
QW2NjWtj+p3XhwdrA3AA50k5OxDifVu0YzMjUwVkm0x/SzHRgVD3pBtjODoJ1zLo
UDL3ZVUuJ1fbpa43/wdQVNGVFDfjBfoMTFTUiBF5kzP3CHjV3H9INZYd1Q/7/rvz
x1nggDtrbAt4JxWSeLDpfMS6MaHnVuoIQDqxovZH6dUSR+r7dbgFwLda+k+ICeAZ
00j0uDPDdAVHSsD2OdbbhN4k4DboNFtaTOSSzEjzHGPj8w1SuJ2f9PYt7qIdy0NP
Nr5xOb3AZi+rmAjw9gBRnpvBgGB3sPgsxlZO/DTcAtAbVSOmAC4RmV1CkPuvr3D7
IwUXvdePjDFp6YD92jcghuSxtKekfzGMz/y5KlTHkj6nCRalvbo4ZjznAhh5rAX2
yQRWE+OC+xHEquE3fdfZBrsYgkgW88b0v3SH6y+jY+HoOFI5OiaMYAjHNVVHrfwA
K4PGQGIRmsay/8gUoTVd5vtxbDbvKHNCbN7KlM/gTcOqCZx9c1NfbG2SNkBEveMC
Y9/S376boDz2iGPxEaF3XuURt4tDE+XeaiNhkvsXSpwB7VRGHUEMqotyomVV5hNI
9iUUPTfbYYDPBORpp2KWfCeHoj73WrNILcZwcNZYXOxs4CiCZYDuaw10kWUPHdPv
rU8s7GQsVRC6XwpU3SyT12c8Mv8sj/ipzKepYw9qc6/3OtqtvVlXGC+9ITrxPDoI
m1wazyf52EP6awN1TMm9LlqfjoLpdQx57p4q3ujalzLJAzUrH3aBEmS7mCPHiDvs
dYSHNAzGmpRTo5ZuGEy8rjMJ9LXayNzPQ+u7pWr+oB0uDKHh+95ldQakeQoTYcEv
mXCW68yn4kbwa/tJ4qSB3OasiYS2DsFCPm7kPsbMEyz1Njr7u0UL9NmxstYwLw1I
iItbKdp09/3lI6pd/5901++ucPt3+fa6QftHHip730PhA7vJnwVeMHi7NmoxLR1h
CKpWGWcPhwCLWeDG4jI0cKx/N/qrDZqMuGKabx/YqvurB8GAzrs+dSDEzVUtWsj6
28FQC/KVt0eGdoQtcmbW7L898WOqxaVFOlrTqH5KqV/ymdPVthkESElBXyzKelcW
VeyIG7Ns4HN8TZZs3kBNdYtw3RZagFqQtxXkLlFMJCdieH0pDN4GMx+zKBZsXhun
YDfM6Y73koQct7kAA4t5BZx2kOVnDCb1sc1jHaZAcjuIKYn3RNwU1MG0+w29Nn7b
9OvvNAAJeWZI50f37Z8yBaz1KWecinw6MrBD0UGK/nxPbNGtTD8b4btRbPW9E/RB
O4QkuB/HlkomVmrLB9/51konXtbY5gxmtZCtzQQ3oo9S4TFnUrs5LAczzJkdnj3N
GpEya1vVgtqds4IXSZKLQLflhLW34suxBjXPgh03YMx5jU8LAxBvUxO8UH1vA9pk
BTMRzGX/TSxnxUThmTtsfEi/8/VtgauZKTTnzlYGpuF3g+AdnQpkKj9xxe0pFXWJ
KRcDJrpvD9PbNV+mf+v5sGZCfzNhlOHjuQQm3z0NU/1SI9fbj9rfLjttidrgbaRR
Zrg8jx8JQCcbwQRMXdY7xZ+odRwxWybfGMuFyJy9LSans3nRLQSwNn4HyTXtEc54
XjVntn8GWffFgmRVpyoDeRRFOGf6OUqo8+vro/jaxNu6Or3rHYWgT4wDviQB1BX7
GcH7AQPuWXVAHTvBjQMXQagcPVK0JTksBn2m6PgEt0F7cbL5h9hnB7iV7BOkD3GW
uLxNoD/JMPImMTx17lrIZkIzYyypixI475tPJGjwIZByKpm11Og2zP97w0uCb1wP
GNsu/Gt5GU0wF+Hy9/RIjwtIS9YlVHwyFSJ7G4jV7cnGevj4fnlbS44kAHkMEdM6
iRkAcIEbkH4dE5kESlBKr4kH0Q6Zx2oDIBo72E/8xiyfI3KuB4VV73EE0FYzvep2
7fR4Dz61F13b+j2jaY9smRZv4uRmxti/14OzEfXUzcpOGD5j3VQTeaCouU5htYWV
zUM9Qw4jd+OM4JLtVBYojQfZlk2w5GYPqeAbBp5VWtz/GZ19eL4hibShWWqf5DNc
EKEpxoQHUfC/lQbiMQEPxK4C0zFroeTLGn/MJiPyukQPL2M3lVf/hTbEL4UCfeXC
B86xVvg7j/pBcxEcW/+M0UpPd96hEDosCRO0JMKI0DxSJunK1e8cK8fljmBnxOxK
D7b4U0dCKJc/AkspJKDYGH8QyLEu/mk6PiTOarmrVSgHFgmcCGwGrig5ioJ6zTXW
kMTUasF0m338GE5ScdpxufvmZ1XmsrCOw5S+MAC2k/mgrAAPdPiswgkZSRlfUxJl
cHdrbj0aU0eVdrCji4MgNvOw5NwNH3mn3H4yF7mAnxeJibjY0/ssKYPNfP1JG+g1
lez+35XNvWtPpaEeVOMb2WDhoiAuMNkUXldRSXUr4UyFFIN3kkU6oKDDxSr3s5kY
s/eqAQVEcUlxCNddHysfE4NVyXoUfE4npzbYEM6vpeHYht/XoCEkSuHrpafWw8EO
saB62HasnOFo0EG4RrFXWfvpl+fyI9Q8OsFduP/UIqJoi97vwjQ85KAWHFtqs9FJ
wUIgB5Igs8c1VESS/wx5yqPmUlItQvz+SBJSDgCquApkV12okIsNnpVNRjzuVyXO
1I5uOc8jxBX29376tuVVmHHmvqr+ChqjGkxbwPWRqyHPe3EJl0hrbA3qbXe1j4x+
ME2nDhksEfRBLEokdNeHoLFu1suBMwfd+EMynJCuhGsP/sm8u46eGWoJVwvHklk9
Z64l0y5GkDUVX7wvImIHWABWjycHkNUiEjX3cntMnfY2sPhpt49e2zl0WTnwgCwh
s8aUt4eom+ZP6As7AncqQxmFAnCcytkLjGPsYRrjWxTwP4+4a7TMYywC8gaNloyc
vPbQvLD1UufSOcu+1+qkYi7+nMSgakbph4Mdhlji0y1NluHqWbnPLNPXZPdmEiO+
6hOI6VTVcHZhiyXfyaP/HVP202orXZA1T/mTWNLBtzLXQsmyk3wxElCVSWWXwHYq
pHxhtGjRIw4mMFZyosSEZko659OgBDaD/jMHgxUdZ8ctLKcRLadPMpBi0thJPXCH
ZfHZsSYT7DqKBHITkr8tK1/KeDsljIzKEjyldCTtPV95OSEIhXQ1XpsmZm0BJ7Qj
q7UmbeuNf5bVFjmFVtO4t1Mxym0ogSlVR+bXxQTl9ZeMr5PA6gxSmeXyl7QIAPAF
AxRe3RgZtZt/ldoGq79K4DH6Y9meoymcsYywRUNvUrOgV63epTj5fKSw4Kc5ELWS
1V/yCrpNOZlmmNd/AXqURStbyYcv5a8GWazqiFZX4GGPKZ+QIrDsSTZ3EQSDCdf0
50tBwb6VpLPBNWorz6HTT/m0VnvtNi4zXuf69XnACjqEoqkbcEBBF5v3ea7/7276
a2cLRuI6aak9oRETXrQwEwFoWQMncihE9P+Z14mk/MNT2XVLaaf/QtuNliHedN7p
yLW6ZbTYd/vK+BZEAyR7pconj0u5wPHzs+zHM/ayw6/CbPu2BIAnojrtvIAoDOcP
VBIQbp5wfFqTfEaik+6OD2usvFBfsAC+lj4gNzJN79jPg7sfi/EW4PtXNH72ooVq
IhgipmHxdQpF5dQ7zvHcluQ5leRH/fdAj3G0eHkjAFWGpO3bGIVe/L+4oO4fallZ
WPRIhPxw0bmiQRQN5YYinhLkr87m99BeguozFSQTxuLz+1VcsJI0rajjqSD3BeuN
4IE6js951wkEbyaBN3Ek2NAVKbBKNtFb7H0MAi6y+2EmTf/keRkmpEhHvSO1Sx1q
UWHkiXcGPKobRmVYuqw5vx23Z1UxGz7PICYdKe2A19w9YAzMexpkKMczS55icg8T
HOJOsm4b4JsZ50yJrocfLdrytK+vza51XPAERxw9KhZ2THSp9maWoBgDRk7a4tsp
k06NlD6kiZgWJS526xn8PjUrJg9cC77RZulG1W9xkGy4FSjXrmN5kVMx84nETH7b
O07dJ015WktuP8JGyVjRLgg3Py1hLCjKoZ4VtMPh17TBRlmLDOO/Gjzzc9rPEd2z
N8MkhHw3yHHjW3iYvFz2fdn1XC4eqUWMQhw2F7P5FLy1NSCE/4NnMmUsjzj38eWt
a35+uDXNrn81lZKQBePX1TG5KXOrrpLFHA6k3dUtx/hrlr/rRIfShleUkojztwwI
Vib5iV8n5A/8YCMLbzdxV67xdh01SYsMFgv9lDcSC5haRaDB3bA+AuCCzIVV6jIB
fd5XxkMhrwv7XZm6aBH/gUBmX6wxZyq0hcXgEu4Ms66FIaZFliwvsrDLjGH1go3J
VUE0GZtJKSy0VxW2RlRwLH+LmTjRRGFHiTwqDQ2yBpp3umk8uCK7TVMlh4fTYIOa
BmgSU9sdETCbKyDwVFQBPP3F3jw+sBfP/3/V+m6lkAF3fsYwQKlHlWne2BMqafz/
L7K30Eh2owwHor3qx5FYElOTIx+2qhaLpDzAQmSR4Gi374OGlKV0ux8hsRiLYUrS
r/wIh331h9cV0dzCAQzuiZ66tKFjNgFSwnl03pX55IEBsF8I4f0YDAtrFwYzJuJk
/MghCVB9w0nGuZ4dkcmmMLWaVUatqnVE99IA2Iybzj0VHQ43A+ek/5sNXYSHNsBI
OKHOMrBd4v/OtpMMGWJVgTftT0wC90vchi0oOLIjBVz+zH0+2iT7g3Yx8l/mHmuD
/mrzL/m6CPtJX+7FU1uuPNnVcuyIVundJWM8e250oMln2+s1Y3OuTqS8GpPYc0PH
hB5cO3c1TX/DASks0Vikre9kuCr67fE+OilybDbekgRJrvPfRosfb5M80lCj0aVo
/66IOj8cHZrYUmAvTI+EutkAYNkHPNsP+UT26jnJIpZypoFm4gwM8zXFyaqgX8Iu
+jswyiSQQYBrS8Imov+6UlpHoCc80WS+DFoL97ZdAtX+lLZ+kf8TN1TYu9UMQdyx
pXCUg7gnr95Tog7KpB4GR0J83wE1n/E8CckfhaedPFxoy1iMA/bZCk8G3WbQwAYA
ARpZEw9EKSk5pn3LCK/2R9r3aLw0GZjDbSO4PXPAkbhsfJaKDITR5UxNvnCcOimU
TV1Uqcyb5IyPu6L/cM3I03SC+d1fVQCWS3uAc+4zb4s6dARyUuaZeI0A5/Zl4Tch
Qp1p1MRyVoiIPNe/ZT60x+xhFueyIKXlwuVE5bPUs5OpGtmfc7pgdvXF+XsWgitS
0ZNBxz7X5HsJarp55+eiQK7mWkig8tQtlfIBR+P3VUHi7dZHJPM4C4KzSsDfpcF7
C2GTB5ve4qBsVodCu+SLlPdRpUNPZWFTQp9O6EMu/BmweYHDUhakJ/EZdY+bF+1k
P68GSfMTcyPJlogKsOyVrwGdt5h8gjPrjEXSlHSOiEdG6JWw4yfws9b/4jYelfW4
79kl9BKnZds+q3y85NiBpnqrbX60B9cMqLRDziY6ZkSTzHm9I1yHfNDWPuJqxoKh
AWWfaJ3Mg55o1RN8gBwmHU573h9E1Eeia283QOM2IWPv2d/gdNqHHXQ+vnvtEKCH
TU2Aa+AEsnbvVJvNfg8a4fHbzQrsHwno88Xo97lbqjr+vQA+lhEBkvhCU7Cr5/Ts
4AaCn6pzRRIJbTqnL4+ZJLt7IMYs2TRo9r80TgRJ+XCau6Zu5xs4rkRn3LtaDimx
Q7xKHFk8e0Pl0cJgIXhQ3pmSINqJUFwNIsN7OWddByutt2ecOUllRaP6w7Fy72KC
SxnoNShXDFVtuue+8gIR8nln9HrghzQX5YVKuFGF2CT+2rW9/RJ9nXOkxque5Uj9
RBpVPw6E5K6p3RH3fJapf1NnKQ+dxUqN4WNMTXHmhZrFlC80D60xvUBexXdFa5bF
ApsmcpCoBfNaMVAIerFxuoZFx6imyXTDznimZkr9QOwdbb1ke+H1BBiXNxR9IQcC
uyC8koIXJTN84XMQC+uri/tATV3C5NVFO/j0G8Htv1FyaaDnYFXsrC0L3jQlHxZo
r1Q4dQ8TXYzfiV05IDeO+XQuM0Ird/V8RjsG7UPC7jFVs51cc67dTYoCDRawC+Cf
Wk1XhtA+7qANNScaOCktX0TAkq2N2w/DgQ5mL2S2g3ka/NGXT+EZz7MuXaAiqmz8
Dfe1Gq67wc+Yd54hQ5XzrMZ1dO1oM1U/UFbexwDTcD5HNZ0HRcPFb9FoRfpCfN2Y
tbj+XBQ82qCBjdRV0RGOzMQuHCDfbez16IEuw7+gpnHLiIxEe+Kf2gu4xAD49uq0
dBVv0rIq37yehxg53pmO8Brgg4sIa0ncBUIPKxmlaZ9u38zQqhhAemGfdWwWOV+R
NDYCfe71iG+SVNN3/cM3iZjXi0QnUUJEX+RUaNwt/VF9mfDWsoCVYYvyPNhO6qQM
MMcd7LtlPGMLlZBCcwtQcFxjkylV747b7jRBoARbmko09ZKOJnJtAPhm7c4UZC+4
Du4VQmeOlEniXqEWCfx9kT3zPWOv9BA1iaEt0ccKGPeTP7chexOk10Xj1sbbfKb1
pb+NtN0TwEYruGtta+Q2jMuQKCgI34bBHURt9qdfl8dFe6Ot16u9Q1D1B1j0hD1f
7hrXNmqCH/sszIK7As5SGowCjCkGF7hmPavBGPoXEk/jXXScbq0hLx9V8uKbjfqF
/2bwlloICpRSqTs/0DJmsrebjIoLbATVtFt6NOJ+lcS/U8u/R8p2wrStI/miJTpd
5swFsj2OP/FF1gDQRPkoY4/rw7uBqr0oBoVdVKamtJjwC0OK5wbfpUffv6dLUfPm
armV20D5unPBq0eV/PCMBP9axB253Ae8j7yMm0941Jx/JPWTW1Y/3ZC5zzgP7Slm
JRxVYVcAs0Ax+TxowWfiki+Y6mz1urebaHK33o2FnP6BhXDk/y+HB+QyV5rpHAzd
nFIujmtzgunFqQ7kbFmfbn53dFJGKDk++MF9YUPPGOTC62B1kEmj0gKw+ITLDUCV
l8VZUCMask8GCEcvUAdL2VSnFcIb6TogbI/rU+1sVBXjvLuqxv5xFmtrU8hWi87J
CeeWbYBf6YraZB0ebUMFyxKRHzoKRiyxuCNw+cKR9lTAzKZcxk2BobpA9k7/nWkV
zOb6+BDmScOS6oSWEDvU6fwvCTMrsEovxOuSrBZOFJcJsp2WkZaJS4DIfM/0yAlb
jAOTtcWF3R0vnR99cjs3FIXSwzJISrzjp3DqHxhzIBZq1LarkS8dM/6QN+I3hiYd
N+l/181uOxz3JDvMPtikn9+MXZn9+mhnGvaPJyL+njKgBw0mcTMdQilo+uU2QRsF
6tkpHYooLWhVeNlqLNkEbCJce+m6nkhU/6T4TcyhbqXluveDJcjEN24rVT6UEMG7
lnKk6xlHRsYB5d6T8lN+aDKzTjiRs5FL86L+3EtCdb7j4yTaYxh6qR7TceAqutN6
5nK6ZUMfejJXg4P8XUIl0mjrerDOXjpQYNaCnwM097iGIsPi6eu1E6ZvNW+uJZrB
UbhLIyKz4CjV0P010yuVrtKXi1Ps/PxjVx0UZR6nZhu2TUUrq3EExkn2Ct3ViF4X
1bkYAaT/+tRPhpEpQ/iYibbW5T2YRQATmZp5Cfc4gu0l4WCpQCtfv2hGhGZ1MLMF
3KM+7SIGKpHLJuii48asEWfZjoEjljDIOIX2zE2Bp7ckDDYFo+Vpc9pI0buRyplj
rx44d7les/qD4SQzGsGcOh+XCG7jaCov+nmsOZd+naMRcseXUd9WwbteTiuAckiy
ePPhVKUJRBj89E6NS7Nc87TVRoDUVWkRRLsyF5M1u3E2391rkMb9JzoXa3xBbq5J
nbqlVK3/Ty1W46JpOoNfLykwKK3EOCsZ2PcS+YuwTWV4al/ltk6BgUj8f3sj9FME
pBITWEjCeG84uFyTS0u7Rp8laJpaVz96qllFNftuIHZmf+VMIMCuPJpIwEGbmczQ
+HO4i1nSiBzdgsiCsjr3FQjovUrsCVnoWgQv7FEK3Xnv5UQHaq0JytL45cRhfMx6
8h1S4QGGdAV3CSykD7KEr1EOBCcuIDMLMhzPqZ3FY67PuZ8NHiqHCCkqZMEzj50s
ZqQNSLxvHsYzjKgFzKM0x29WY7Bd1Ro+QALd4PU7xl6bS7r6qOFjwBemm//vq/q6
7iowagGPeN8TL2ThWteINsHyaJ6bMuWmDHmFRVRPvlnCyEuPdtJsdA007Um+I6g4
bcmS9BX2QkWD8VAbFFpZHP20LCQaefVHaXlt5BN+Ejf9aRgIEkfoGWADPie0vnoC
zEKvlf3dYGr5NEp91vA6raGuQBLdMwh5qLiq8pMYaLtHXBns5pAnwD75FcVUAed4
uw/FM1ut7Ov4dqLwcTr4U3Hl/WNArTwgTVEDhJFyQ0HiVcYRi/u1I+O7TazFrDqo
LcsSMjWFAy22IgW+3Ij9iH6h05fMC6uCaTypJvcHCm4iGBu1Hu7XsV/h1vrKCK8g
M70Q5xl5P2j0HPQzIl3O1K1uboTTrjlTRJP4RpNSogI5V39ENONl+PDFl/i/Je2J
k4636IW24AlhvDYKmCJ/8Rid0Lu46/4BYiUnoJZ8oB7Olyss4n4VpqZzIpWkdXGY
NneeK4Bdcc/BK53aGb1lAx9mirp/FdD96WlBPVqx5blLBZMHRQ8dnzSYYQvT2U8a
qjSFsJLnPZ3NB2fLeVJ/tc1osjKaxDL6NkgwmrJMN8Cv6bsPw6FvxZuSAyvjwMh+
+sxZZJnmW+1bNrn3gEYXezv1UxQGXelQvZQcIsqaPKVKSI4vQ+vzf4eqo0wL0wZA
4Q0LOn6odb6EATjA5NLKzWlIvH73vNu5nMTyy6jPuxNQyua+V8GVdj8/qC8BTPM9
86FANAyFnINPZl9o0Dhh+MqgDihlB3PpSccXe2co+Vmqu30x+F+/dGt4BvvIbpds
X1GBRZb0uXyrXcovHpXxe3zGkHDk0i8TBQMJHyf+n/l9r1BMeIfYFQypm+xCswsz
pTWmQDqUnff5hZNy/ZqZ2T+A7UajnbUaIatjpiQ8WbffH5Va4czJiKed7sXYHiR1
CYistvo+5acSADIkr8gPkiJr3csAVZwzHSxfFBbEpJ0TKC1BZB5NiDUW/L3m022C
KW0Re1eGa3WTsZAcEj4qv1mKs0hqWNjpMEQ/8k1AhFQxiyxGI+Es2kXx/t6Pw9kN
f9qJAH1vRoXjg6iBz/BjQ0RY0rDywtIwwfOI+7cUlJmk0NyBZNGEpphrQus8l0V6
eQfsjanbClJ10YVVg4VoiIsyzEUlHzs2TbcwgtzIZ4VPjCMgDzmcTDaybmhb1bCC
Qwvb3ydiKGguseHaRgC2+XamkR7/PLtzL2Uq/LKNsPltLvQodcp7F/4kfe9GfSEj
tcZuYOUN9mH766Pj/SeKCAk29lM4FyrLJPsMC9F83WLoha2JaVrKyROARHGkAGPe
X9qghORfYfFZ0cIhhEFm/naVATTPjazVep+XVV1l3faCTVphmD3hRmqle+3Z7KCI
Tk1B+usKhFmXF6OVWWvRiQL/ywDH7vNbwrbvuZvOb5j9Z4smibl4yg55cZpwl9Nn
KQtd8c1/MvBcPF5jcJSnQdCKM8rlc8NHGMnP6TvIQdbUwGNShoMhu7xoZVNLDng9
3qs+3NSi+V/mkzE1hEbhJZYdwFRMW0S9QiqmVlxqpOZn96ZaVsnhJCNcef29uOWr
J5VaRFyeqUcX/sbJeCIMvMxKCZNDDubZROcXeSgIxYF6gmAloeg45IQuPtSKe+dG
aDmRvcCe6FwyVTvpjupJAeDzDzMV6DxUUdAt6YzZWDmFqJCkMygPFChcZ/Xm91Ru
mPD5XHMtHWdkStcM7u1Fbct9JH4ciws5+JDmLxnyfQEX3XLY/5Q/ZKkYG6GO4Af/
Iyb3aqY3x1G5+5O8BBiBhh2a3cKjBm28Us0j4egd9LExb2T3TeVstgtbVEBdFaCA
8OoWWNiFvpunsEDBGfcN2lOijkg/+b9FRYo1Qw555KArB4WiA8ASza7IaGCWxcc1
nR6tD5DkWveAMfoNeMXZlTL5KRfAc7aMgbQmUPednQzQxKhIR1tsemMFrS10BRAW
QhPG0SOZ5QgiQYioPxVtYmWgCJxkmZpPjzGJEdHQzmVSRnQAJesOT4ddM86NzO52
3tryy11XAeWjoGcUfl+UEuvfCD3wRiBjcGfMYVdYLytjgT7kJO6a6evYJz1xqcme
e2vpDHgs+yUze6vE1csD54pwl/DvwJkX3/msyPtUvBV67gcHKx6GBPPB2/qIDnea
AIg4McJihxOBK0n/rOfKl+PAbN+WYgbH+NekDJW0HkpaJq/XS8q/Upgf8barwT7+
11a/bOzohQn+vuU1WTCCESJjZ1Y/mRWjP0jrEIcZ7ljbHD6AMVHR552V6EFHpMLO
ezWaMv3rD7DfJJXqm9uISnjyc6eZZOHea9nMiaShRIoWWbwh4DbQ5fV4AzqtZiFx
GbgxCniwvLB+YenmBxI5iBZWM47t4jAOz27Hsku7HFiaz9RIGpDuz3G++hpk6Rwc
+AUJQ/0P+UTGRyRLe2IyDLELg0WD9tREV/wl6ONfrgYbcjcDGC5TRDFls89y4dj8
VdoQMlbNqttH5aR83kIq4PF/D5d3RtuEE7zlM4lDUyLKtOKj/H7zlsJTltECKYJ/
R1Q3uve2IC8fkjSi++sidqvqsBCfWtRQt8OGyJi4QIuF6Zp7bil45nvDMgnvgeqN
JsmvZ8uChuE9+B39/45JcQLIr1IuUCzfOmaqJlyttOMtug7aG/g6QinLMBIlP1wQ
YVIDzCehKfycP+iJSdpuA6kguuhGVWjXSLGQm/vb8zALlpxWX/jeoTkTM2yLuvIl
sG/fPlOtJ3OxxczFIxEsJjTlYbjVHUavqbZ2C2V+u8powsBL8nSqtVWHhGnpFF1S
2xpfxAScq7fWKBvlaLE+vHXzndTZg0GG7ZGLGfYHKqLjmhR0DPFhpHT2FdDwnesd
JG2258OLBiQEI4mIujOQHuSTGKonh4ak+p8kqBhx8kkiWeivWflRvHltVNjGtYMM
lmrtlF2Bu3VVmH2k6/FtjSuvwVs4cwt2bMyA8pWb+2p47XmInPAPZuyeleoNPAgS
+KNQ3p6O7rF/t4D+Pss7fm/52pXl3TxncTb9GF+s/N79gy5/FvlIxwfKQocf3vCb
mqsD1aRBGkFdnZ5mmDRbhTlbFJvDV68036zxlRTm7BtPJmn9JvDg+S7tDYSZyKqf
dwCxNBDjOrhWluHsu31Q1khSZrfeIyvCtSWsJDVdzjG2WgoS6Ce+FVA/LYFJQmRS
6/qOVXaOGIHdxIZ1bBA3wJB3yDqRhsSuYQDKU4XaQwrfAspy3mEHBpWPN7iy6K1z
WdBKtl4ZUOemQDUiJQY1MdDZerDRATtRT2dTml6yCsNYJddlggFnqDYvUILSR7Qs
QhP70f2Ekrdyu3+HA1FnzylKiplVvazTKBsKi6NuMDikjMFz9MvmGTSEPYw+UKkJ
goM76l3zn6Z7nn12hrPn8b/qplCCegL9iskR8zv5jcGQGokvzueP5VDRoNMCpZRK
KSuncJWGh4IdHXu6QQpzGOVQjcHxguwN6Wy6oZDntHsqqvKb/g7C8bSdanuFjRRv
ZxKe7zrRbe6q1+NKa5mXTqUDLgsewhHfXvckTJsntNnBB5pPoG18IQSzacbm+K14
VzbREtnHdiXaDCEyZMhR5OEqregkRgzy1C9stKs3DDCfNhyjlql0V1PgnojJu+6K
RTF31FvjDjblgjaJvTfLuYFhUBi8tRHFDfOz7hWlCz9Xxqqy42u30uUNd1vkl5yl
gI59HbR5eGw3wrKkJ4+IZ0B8VAwU5Kxdx3/z/D3u3y8zOdYAB0I8hFnATcbv6gLp
Bfx+3YtO13pkPM1I8xj3tLj34k9Mn0/1AuGhBqoeKFhp7GqNywHM2Ay42KPCGCJ0
2jNJ/XiDm4RJS9OCATJidOv59VxjHXJNYrgcwPFRx4tAfhnrQLqwr+vbsnT8TA/M
KyJ5YUjx5ibN0b4WYjDkkTfVFNaT/RJF+570CgfNq/llG31LJgE+wMvT/rlJEpVt
ZTMQAeRyqX/HWg25s38oxcGJ1CCCdwVfNBY9uMLc9BIKtkEGB5MCIK+uSeA269nE
9WIUI6CxpCK1dUghnCXWaAYNYxI2p15uCyxzcOmrtiOTgW4KKvGelCb7v0Cvggel
aIFqdmK0sKd96uelfXSAPUFkcZvVls6LVbI0pdgAhQCz4F8g4fNyPRTk3j35Z4H2
NgpK0kLZwJFUzvFdXKuDUoRbTem+JMOM+OxsugQnN7+9d0fuJoqcwa6kO1q4EL/y
dswQ8AGHPBOOy+6HTUmOpfOR8M9ohOBdOR7FfQl+pnTW9eW1UllBPyDNPQ48qAOI
48B5o+RGmLAhc6alQcmthKoEVWkz/LdaYgokZBc/egWuf3V+yxaK+aOtqefDF4gu
oWuuMYKEvkknj7h6v/TJNPkqD9aoOeyn9Tc9bdaGDoX9EU5a0rUiW3xkL2R4rXyU
CaCBhr5D3YYASw4R6QU6zclDHdBXdQo84slkpEZIGzQ3mEsqzr8zdRJw6ASpC+xY
9ePyO+DYzxfIoccfGI28mpYoef5a86jYKlmVk+wBUspRTNnsn+cFN9UYQOq4acke
ksg4N92zNErc4BM+Ov26+W/+MUbACrDkYFijPkuXz1FRa9AXQsIdD/d8qV3F4OxB
FonT6Y6HEvgLVkfzTh18dLR9GD/aIxG7zYzOJwwX4Q3TZNYxzwbpRcUhx64wdDsh
462e5CrRmAt15aGMl27fuAMpYOxfeSs97LHitEJ5SOFZK09+FM2MpGn0ueOwF1PL
y7UIuC0+v7UAyQRFTwIBvdw3IP755yrgjuS9tiGEIprCjT3Bp2OYEgZGL6zcf1L8
lLFV3mCxdn72q27R8JbRC6YgcIFooVhyn9wpsINccQx1YtG176N1Q+MM/fC5p+mN
9+d0diZDZB8NoBrUgX9zIaT9W2C7WHASF/s+l1QZ8n0TGKEOyxQX5OqAjRqlm4e5
+c4On8KRt7yaTpDwhSppU2IgdALauF6W2W5HpjMYp7bebBqgcPxnXCoduloi5qF7
BvvoIz0X6P/xARYq9+46wi7m15tgOAmMNLCIP989V9wHWXOdt7BxEQ8/wW5Ao+/D
/JKR77vlv9roIlcqtxqhdv+ZfmeLqXGyNK2HezohM9C5Bm4QmW90L5hzDQS8OfsE
6tAeUaKFqMCzRlF9ApCn1PwOiit91bmiVxXFmmk4XtQyoqOs++44OtqCsZZuqQhZ
xrb5ncI2QmJJAYtlJi9S0H/hIzHApxEvhxmS6GFNlZX/nvP67N7GpDNQb3nlBd4u
3fuIo10oJXQZaGN6hFjxxSF2x3J2hxtrTXgAy9uwAqeOMw0cRODaMsGNpkhMXN8A
danRWBbH9iEAaqdLHUg6XlYG1FILaIQY3Fon82u1ToKjVfQgfzGrH5YET7sfMSbm
G1nDxOHOVV8PooMpLnxeWKd2iKW2hUlT5+lEfB4dYTC0WGowoIAC+c32FMS+B2tZ
XpsTFc5DTQPZVQhR13u7DkUzYbKbnFYcHJzJkKwBcZHKaPc1HcvegqAuoCwAbdrd
0mnJlWIg3p/P0JATjsj4Vuq5zTlDNwFMOvEXst3WDbbo2iqJADsieyyJkqj1f+F/
5xcvY4lddSjDrVg38ScXEaXe7TbEOfEQPku+Z6gQ9kDHtaD+PGZhCw2G5W1nxRAR
gY4jiAKkj5CnoN9Rgvmj2R6mQP5lUqZAerYZiOBK9nnkdOk6j4AG6tlDMab34FX3
v+VwAP/Ezye8hXnhn7muy2cb9/jZYVfqC7fZ9Ec8WWTPPEdAxpbWUuxWiW7ltF7L
eSqHDNyzl7mj3IzhXZ0/fXChl7nKgRWOM3pcdVRauEroAInrHLMKm+XbTutbRd5u
CxrrdIY9wcsZCqeLiHIDWiBRQ/52z/X5X1xZpG2zgrlbxATqSDWeULnsfTgPlhJx
1QuiFNAlSfpE3m52RRpFlEgcfeTEsSLfplKfRwNG70kD7m3b4sjhpbFKimKxVTez
DSwRDqD6ef4QAROWGnwJQA3t109IewsMEl7oyMSk5UpoZra1p8wOnmUKDb0K85XK
dvgrK/g3B8/K0EKB7xWcmzNs87HEQ3Y4nSYZRg42+9udB1eRhVqBXZ8hpqKnZDWK
ZJ9sUeXEpzDAVEdGHoyXZKZCoSrVKW7JVZ4Gl/F12Q24W78ypMCD9eG41e5ndr7k
3gWImLAaIaEGPW2e37jHpC+UpGPdaxZC9uPJ2cKDxKbJClNVODHOdGV5QfROP8NY
QAO09VfQ2mBATzI1yZRhOJe2BCn5fhouQn09iqloTPi4UAbzEG8JDTdkNGBy8dd6
tFTIYpcRofOf+G0QquVEtP2TBQh5ha9A5i3iq/y5wFDE8MRFfY+2NNBa+oYDTrlV
SbpmEZf3GqyA5KS90YH2EKNRnpbDoaWldRClCgc/0Sx6Rja927xQasKdBhRRbARa
RjitT9ygx+mXPx7RdS4+sCzmG+SAkj7ne02zlWqc06JBnhjowLoiW8h2a/fPZekK
9GX63TcpknimgM64KYeN85+fLoBjWmScSqbrCfj9dE+aWpgJ3If5HD6it910U0Ks
v45fu8GWwDL0VbseRkVaxgirfxVWdDMDba1jSJ31t7kse3rJNM3zFmkJ4YpSXnrc
Xjr9PclAWEWHVfGsnWmshd29IVV7pPISeiC1WDepvUstyeCP+FXCbguvuVMTcGgj
MXzaG5vLagcBG0kBCCK/IsIXa2V9FQajnEyS7oCz5jfBsy4dR6hpjx6a/VF3zW06
wQJa/koYAH6uNVCweya3ndY9tvmxgqofT5f5PW/DwZoXnjT1I6vFw4Da9SAOuic7
rxR1EoUnm7UJsM+6JJRvKgyjSC9yI1Nyp6Q9e9T6L65PkkTjy+7r23jsuS+lpzrc
JC6HerHP7iiWeYAxP6n3tpemmcFuY6fucs2iROBKM+dYb4Ob21m99MnLOqaihUkU
2RI0wUQznOmm+nEXK/OOk/dhITAgB8PeCmJDo8Rb5K44If05GNKJCXrfwrF+UkMY
g8TJxJtIwrR6ssAjzTzLw6UXYWY3Ax1XdcsiNgF0Sp5J+EkHPLg7fFt4ptPT81RW
GwhpDPI1zSp9XLFpOb+kFRUxZyZRdTspkcuKGS4ECHvJMulnKTGOdSNcSHToxZ6/
7yjYeGdjdj6+aCyrK6HYjE0ngQeQUT30cQaoYQri1BbUjKnW2mCrAFOBJwceaAbJ
u3km+fE/AwPZpCEl78Ea9RJrBeVLzc9bJ2jR+3ea7c1tvs8IeZz6w3hD6VWpJMhT
0TRngnoqQqhQscwoEm2Gv5haiNMJa5Rf4yEAORGJpIsfrOd5oUJ6cKfNTHRdFRe1
xb7i11/nQO0KM6g3kzlLcgrzOOTPupAX1cpcxeDeoJtPRZBMDk1xDIlNqMNMJsAa
LQdTbNDs0uGqo9/lfHyci/A98u0ygP1FZKAH1hQkPZrBKRVzWZXO8GRpYZGuHu2c
ZBlmfAlV/5imgQSzoU4LVI0xvPJoojBydcieH1vetHPE1o6iML64iRs3H/KS03Xc
7Tm7DMV5y4stpFPn3WfdKDel/ez5XTI39dBOcYEnCc8PrfVIOaXNNgq/Kyw+5GyG
BoyZoc6u1NOSSBO6k4+TuU7pqHjyO+B0DA4MuPSikjB2jgizMDAnvOA74YzYGGR2
GZckWDI24WpZhIlnJ0QxjWxUxwWHG9xm6wBgcd1v0LOgmoGYq+ZVYV9i95jm/VVw
PjJnM5NeLmRJrBu/Fg0r9DJGRyFAxLN8JkutJ2s6FcyBzZAClZJhdC2sLeQigXCl
l+HaSkHB3qT3FaLZdU6IKLIwKlmWb6+DDPRfmRfjvPErME4+MvuqD/b6CVaQntmv
Rp/zeJqEUA7wZDznv2H9FdmXRhUJfvKFDzeYgthimirzlifZdgRLSynqqsUO9fa1
Jx4b7sOQOHxLBuH84k1qHLIzhBA6897kFFP++KhrFtkQCAGtOTxuXmzjtDNSiaUo
2HxRojUyGPi9zlcSKyELNJjitZLDSyg5ZL4cE7cXuUZ05PQcORx4N3P3MTtXuvky
Q9hq/l6MEESpC7sT4NGQLVF6oO/mLU2feL0/7/bn0TrvSdO5q8MkaN9na2H3buCv
JNuiNfoCW3TPtN9oeh+sz8oVyr5VRoAO+W9Cvsyz+uXlYsoou7xym2lHFm9knJA/
HhW97X3f2NheM3rq5z6zmtyRYKcOM91dBLo4McN4sWK1OgCxM+Lrd8mjqt0sYgnz
NyQ4i/mMXHQQYWVAqQBuEWA4EAwbnFp9V+/MTluEtEQgjkf8T1O4tAqVYoh8pGHg
ox4qbOBwhqHX5Olu2wUUbKdFNQtngRnHn8BKIB7eFdGmVI+Mnv8RgqDEQ+7ozMlx
Pwz957dsUNT8oOxTRJRDmd8m5XT0dzAlqeW50PbpHHgAt8yui8VbblxS9aMyczhL
Jr1Aie+Z1k9EzqiEBAgu1P28jCVXq6go8Z9hpShh3nRhF4Vn6vT3FPDzZQp9NpCc
ZFottZIfaTr2VKid6zWtIjc9zLAc5whEech4ldUTIjsBatPEwPn03reohRP1qg9r
kBXhV0EvyUI+mL9fINS6T7Rw98iRRhyFA0WqGyoCv2AEacn2/V14srBz2JuP6b1w
FIjatJukEtrQsZU/SSTfJWNg7DAT2TNg/wGa8FCnstaCvLqLycLVHpjOXsAQXdbR
s/3XYE4n7gj+h+HM5dwPdvv8701jezFdEH49lg9KpbnUliDrGNlnjVgcY83nNBpk
6Mkxm7noX2ak0Uwh2M+a8hVRzXm4ap0eQ879PBvMy2gtBMDomAmJh0WAYMsSaSTF
pVkxHbMWVMqgAkPWx7vLBuZBeXv4O9dv4XLb11Z9j8rLWVHPhT2xggcGtOKyCpnL
EAZBrJsnHLYBnQmlqOVAuxN2Jp1GXg02cownynx2+z7jIhYEQxhdj2CNtbel//LJ
sLNiSdcdrK8YHuOfB+Ohi548taAV5flAmFmipOgJi+fsFudjsugCyjghPWKAPtMF
mPCoinwUVn8wfBFCJPjGtKuAlVWrlRYkO6wUqUpLCPJUQ8dFchPlMdX//unNxg16
LkkPdYYXzie8mfMR8+RpQvn/XYtd2sThtRIngJ9V+W7CZvSQDVF4LB2gv8NCa37/
Bd7mPuKMOQZinZtMaoq8P9H6wHOCLwhmMDtyfZca76n4XQq/w20dDBpQ/oQa0AmY
X3ckYMZQ1hRYYoIV5KL5Dbn+LhFoWjGG9PSEsdBZtka2qiIZ3cPjZbe3C5K6QUB/
ocLsBC+9kJMpvYxtB82ukLDet4N/Vv6oJp4DYLl9l1Gv8TArhqhx1vQhrXrseNA2
jipePy8+KQotV5S4sixU80XQWONdSB295rw2DAp5/Pv6lHLOqqjM5F/419w07pTu
A0s62l2XXmA/HKzNKyK3SOEk4SUGMl9M9SDNcwwAoxWVCz0F9a/m917JwfmfLD1X
mHE2pZkOa970yRrOx37Z1Dk9bPGDu3XSTanFWGi+vKIHMsNsn5zeJFLx7vpkzGRf
PMAfNds9nIJLitSNwD9iNeBkI6N6r/fSSpcaXBlhk3aenXMgLhE9BpmiEaXGCW/t
6qLaK3UNFGasDgGYZ8Qfw7+7wsz8OoWpHSpD9VpFF0reZ5XxTpCsiksOTh67HBll
nkpNWnUmsnlfvykZaU0slOEDmI7QI+g9eRWfvkFp2wFdmQ1oK+oYPo7F/ctRcHks
qy2aczTPz14WxS6RgjZLBAN2Z0EhN6m3mvzNUaQTn0o0+40vLwM7CmTmHZqt6J48
qPzK6+WcMWc+LgITsCedWaYsK3w80fnbKFFte5aySWXJ14lIixdHmEEh3BBx4zT+
saVsOc7rx7nZfWALbrRyDuwqfsC8IC62zLNTW/vZTOW+Qbw/BSBh9cdbc1e/DULi
WXX9nPhPHnQ7g5OmBgCZfJgeRicuPFaUtkoIrk9bcsW2dRnYAspzOlVqVJMQ5JGy
vcsc87THKD73d9fLiGMnAxntVC22zxfV32hQLbulqRwrM2gFhulBARNKuOjZDiGN
iyL8sR4prZaPh38a7RWdvUBCVjj+oOYDiS5T4RT2ePh4E9fBEH56olAn4M2dQDrP
NFoBpK5uzyY5B0eh563uT4wkSxcJSstzRBV+EHo1rAI=
`pragma protect end_protected
