// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KWoey4+Z7scILCYt9pGk65nGc3prRdGdVbpiiDkY/5BG3dLFBwDEGu4LsEwrcHnk
Rnc31JQld1YTd/94GSSF174UgYAeyMiUpvzTAwDfEWScMIsejm4J2gi4jwGkwnIK
Bfv+K9gPZU02jVe4OPPdLjZvmS5vA32+9kcmYrPT064=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5200)
sDZHGSCbEn7lkHfRhs3Lg32nNM/UpG02ym+JtAr1hIsHYuw7QNGB63uNjq/p6lvY
logYWXoFdH6wBbu/C789f3hQLpBCX/qAde4P5pdRW049Hy0H9cLVATrmnEf7O+Uk
Vb7KW2Ey+mysZEbvVef2tcFsxQVo0qmRkOn4E39S/YBAW3kTqG9RzqdeGbccCXbf
2rUaI5U2DkUVcrV3JE1Ag3Dgvyz2f0hRluEaLh7eVYQ1ELwMJLAPRRsREINh4/Ns
n8XAUhBz9nQIow9u15nkXK6RUFtonM6xmWg/iq8C78zZmzojSMGxH7BUlvgZxOIz
ip0VL+FMEG9RxCCdBe0g+EALHcOYqUh9CK9dgDN7bwOV3I2Z4JMUd8PGj5Pow3Kq
NJKT4X1cdeveZ1P/Utor6YaoGv+afADSDRfbYHiNFLI1r7WIpKy0zf8JxtRKGoQC
2CaITr61PLbawaG63HFAxioBP87S07/QuA1AdQoWFfAlyohO5bN0G3KYnOtkIVX5
TmunWzeT7Zoe2i1Bxdxrvr3isFSvbroNR4+/HEUBTmDZ65qp1RAMo90o9Ig+cQ8i
sq9ZJVM8Glp1Ye7uyagehR+DuT4xjEnTBK/Hq6G9znkSBjE1IkAhFTUZZcwImk/W
3ECNKg8sH1zhRCBJBoce0zgbfVrrx+qnkxJx3KXDD+OOD3tcFnuynQwMMPYCxXaf
YJW/3sP5d9KL8rlm/ZR7paNcfR3NA6vKibsIJ9uH6SXatiwxbXKXRlFoBd6aya3X
2It2ptVXc0mBIEOxGUA2YO8v3PG/qijLQoqb/+/4mHm2vx+zGdKU+KxAPAmO0QfY
ctCxMA3LmAgIpKk3SjuARdYkB4DItgEy2v39IZqIcWO/ujrMG/hEgZaXHG/tbaHA
HuCS+KAy3nWRGE9YPQLmHn5I/cQRUY26+dhjztkoB4mfEKron4qpcTCKQvhlb1P7
8nISxu+/ZRhE2mGDEAx8R7lnq16JvJ8oxgcFOwympOA56+DMWlX6dd1Rt4+jc4cz
XmfSw9Cfh5yINVkqgn8+9k86IBbCJ+XO+bsjLAAYgcBB8T5Q1HINpRGSPnOzHWyQ
2q2/3CV6mEKiugpqWQL4daS+v3Eq8hHZfNfXcQUml7VEFXREG/FZ6UbIKGzSH1lR
AxvyFx/n9HTrcFz6b8jd+ozCwvNa+YZZtZ3gPa00tuiXx+k/swKkoL88R+nVCLwf
iQUl5IUKI8F6uxoqXYzwKAjPE7a10QPNvQAaTA3kHK6oCW9f3XI3QykJmnIgCCD+
akSP/tLuuCdJHJvk8sXhBNkl8B5MUwpd2MvYDSwJrG0AwLlpKqMSk2FRzBKJG9sa
S6I0iti/Nv3bEYW5dTbko8Gf8ndh1TSbqe8c1B7O884NSAivBCqmIPixQn9qlmyW
qM7vd1LNXGgVh6pTZEvkBIAsuA4UgDJal/YImwJeqHZblC4g52VcHYOfaMQ5sg/k
SLEKkzBOoIc0WeCcsJejySVpPH2fy9lYFtl2VRk/BrxKKVaLw7qzbQSKZJuVbOxS
llQCfg5oOGPjZ8vpYBEYr8Fq8oM7Tx2eaPVbh5xQbWelcb3VGqn49tjOuEHzNFBS
ZhoAm4Aj6v1Nn7IPaW7r6JLg+Q3ENLlB7Kekrp+L/nARKVZjxy+r92obCp+PLowd
UdAWPuvqZe9jxzKAQLBdCkofSTDzawHZcjyL4b4BZvENtfZKEwpRZJYcp/w7lJEZ
JGwUe/cGgilj7o/qbYm7xILdWAEQjWZZH47/1glkyFgsZRYy4RGZgk4r/WNplHoi
8yjy4I05qOVIw+D7rj1MekLP6l6YYkCG3SDGeTSg1J5VJPNZ+E+Jgt16nUqf/FL6
UcESp9RjOtCNAMhtW9S/LX/eAGU+Uw7auK2M0TKSk37HDGVZuMAjVnvv7zDVrY21
CoqGbmOzIOOt4CQ00m1wJdVYuTq3xNQaDORZmvqfazeYjGcCMjjcBTSFBY+TYuzh
MMvLbNnR5WjA/bKFkxh+4m06gVibYxqGgK8eWF/tCynO/WH/3pUtHasd0z5wRWRc
DTfvhAd0C0J1vmaDjejCpbKIjGuhq67iVpXdK7PoM3RyBSqi5Bp+kUFWShQx8iD5
xUy0mblA1Chgl9EV6k/KEzxXlJkkC/yLXIQHS3QpHPtFXFl39jty5tsDDods383V
cuQ3m5Ml3Kl6ao2bgkTGP8uRrkXFQ/8tdtG3aNOT/07C0Ugpoos8c0E4KdV5svcy
UpymbX83P4ctvSa5vwCgXwFIE73reDlCiZK65jEhOg29V2L4vbw97ZTrHVPCo+bN
wnRTYICliWNINWnIFv/lgWTVEQLNPwdAYCS143ez2nFTTB1gPEw1u88dwAZ1kuSr
DxH2k5sf1yACLDZW8m/m2Bkyu0hYHeaTEPMg/NZGYI8wfikcg1D0qIAu8Xy/5O8v
Gs8AebiNRms9jlw3s+kAwi9UK8SryHOYBapM4ZaYArrMwdxIIPT+zRx9LXje3RWf
B1NjZthILP1Sy0nXLsrVlG6g2gjautSWqwQHRjg7zyBNHg9XbuissmWFmhvuJzhq
ds6d73AvLEvZeQMu23eemWpDpGTF2kYrmaAwOnR3KAq6L1kkZH0sihZEU8M61nVO
wkGj1Bon1i06eNeKK6uiN3cgVGTRQmXA0ZaUla/FezRJZEKnt648kILXDGgmG26o
DPDXg6+Req8ZLuNZO7U/PB95nPYYfNEgbtdXHb0CbmgjHVEwOwAXJiQ+Foie9rFh
56ClKq2yijsJ6WhGNYqE6FjAtCTH+KHL0HSQExlqLW1M+d48bMjM+AO+Udv55cRS
r5evrjhXnP9sqPVEvEVpUwPQyGirv+dwwgdQPGJecswuh9sbxo0scxWrBbTxxHUJ
/7QCD9O+jxIAFNtmWLvPYUYe8zAXnv00BtNkypKzD9Z4WhqX//uD6dL6o2sGUukF
e5n7/OZgHhkZgN9SE4DXSW2K65WqQQhEd3KYedty0jr2iAV3807N6MKtVUH8W11d
rFhGCK3jRG7ZhFId7JQ54AXtHnFIScG7L2LSksY+mG9a7jx708wItjhneDbUyEzc
aOmrSQ4TDGS52rlEmxdPR0x5pfTOIfmOe2gPU3CnCOKWsi4jzkf5gNVQcOZpt/Gl
4bO8YsD0gPeko+MPWDYXhKskjz5De6kPswbn66Qb1B30K7/tnrfQSFNhXu/0/2mO
xTuectxzaCGK1xm0jcfkSq8ohpsMK7ep9yXx6AOK1QGtqgbp/4AHLROOnM9PRhgw
3U1MjyhGSnMmZO1ys7gfXNKimVrBQRNctvQJQOeSn2kF0ez6aCjRsuNFktwSmLav
7hQLd6oBp5FCBHbNn7jg4tapddNnWv1sa6MXaFgJqD8xeKdpHjxXtbk4udrxlFAq
/OqXz5ZZKshFvoyv2FQwl3gI59WSROpZYCRM1D6FMWqnHzcyAxyFZKbbeXEVyQOE
PTyBe0frtodC0A6Yh+GL3LEyl/HlpTNX0VUaY/CBpYIQfzKQ6oPec/lu7trZysXN
DfuE1rZIxI7nZAeR4eH+S9NIThNXgZg6yzmWlAn1ob3wPkWrqxin6jj3aGQTIf6j
mV4qM2XDs6FVGsxNNUk8SlWX2/hcRBHOR1g2n76w1/HUw/SNo5rPcUod3NQxj6kQ
5ki9Z7mQXtqEgjmMep52RAgKgc0wnVVgq/fJuYqyUAyRM9i2Newo3Y6gzuO+dmES
aJ9XqXxVmGr868ZyrRDYi6MKYdfiHSXdJHJ7uGnX268NYAV92id1NRLPTNBxjCSe
2n+3ZU6oUZ45wjIpFoPkWLb52RkIoHvY/JsOZUtfF0JuCyPySc9M84wzho6ByPGa
1ZU/Bvlo/g60uPzUcoRhmaVziUXKHo4kB0Nu9/Thx9JCnLt3+hawIRFvYjc1up7f
Dyg7rtpFENFp7g/BftJaKsUHtRG40k+8QWvcCmA+nOSQttohfBsDtfCYhGtoP5AT
+dlWpClvpkmfyToJ4qqujS9KmMiQXQ0m86Tuu2Rs0iYyZFgoVycLmOWKFgopxyfp
bEYHbYaOIfG0tM7xYptXuCFiq1eQENQJE/M1Jry18wdkVYWj7wQpt2EezDR8a90j
ciT/PnXKbd5Rn5yddbJDNKvivAmGTdxZ6Mji/kCP1ztm5e58zmmYt/woVib/KGXp
P6qn63ZbQc07FoXacSUsqHOl8aWqR2TI0b7b8cnTPBCgkZ7UJpFMuBSLFb/Jmqnd
adQ0lZ69JCzH2SC6xxxDopvKXoTTzYVuxBc8Dk25zFrAHQu8ED3ez9XJGe+w9CCQ
H5WUNaS9KmmLtmbE0TS9fTLgIl2IeA7+k4x4dDxphJDhYAYaeXtkiRqh7fp/Nt85
Vfun+xq8sGafm+my5g4fHo6mdvodPTP9NvKW/LqCN5KL7o8R7D4ZcsLzBWG2q2ao
cuFm5XVgYfq/FNKexhpsTcNmYYuT7ZfChSze4Rt6qpd/mXOmzGpoQXkE+VxA/U2B
DT2nQvmvVGMawCiX8DtGlMSloKwJuMBoj5B7/yNFZVqqs1A6Kv95XJzivxkwjg2h
S7Itq026GKRx5TTSGWM1wcFeO1tUxPVSar9/xbA1KmwOsiJRbS0KbnvXRDjVdWV1
AwO9zmX5wkw7EhfpVl9jJYHincWGxqwMCOP+qy8gI67sO4rctWCwyV2ePQhfkQh0
J+eY1R2G28mzsQt4/Up8KOZSm9ksdzysXqHIaUnoJyQ3gA4Jfm/Jc9oB6wSSeIkn
n3xon/J/cTdcWnd0UDt4QlOi0ieOGFvmEFkWHWEgvnJNRvZE7qXae6oyiQGdfp+u
KvskEs4P7wQaZpc/zyzCKxMnf6uqP8mkbOBKDSVUktoUT5B/rx+AsB1FIdy8WW/Z
M4L8EuuZ38DaZPOvyGXmwCSMYUdNn1PzhmQuH4LrB0a2Tm4uHYdHv9ZCk+n+YBD5
3KNWiPoLfHPlIGxTHm1Xps/jPxYHL8xLtGbPGDuj57uvnJzFOkbXhjTSkXB+mfU3
i50mXR8vizifY49aYF6b3iI5OSwTLvgDr65pWXEgr+GOVBJ/5yp3kCzXtb4N5jl+
o2x8lgAHCBVDTzj4YzQOvyaYZ7QUgXbrD/xLTd37xxZf26esZsRPZOz9AeLpNfaH
xTV+p9QfoFgH4rtmHoZ21H2NPayg13UH2/+H+YIkXg3wAWgBxRBkZxJZbBoBmNT/
zMOYHHHFPx/eogulUGYE99ZjpgHPQMRqzH80EOHz3Yz7wsTZgCmbAl3mQwwomkqa
7X4aY7+yqrnuKMZczuoNBtffCFVAsBIu+OIfaZWxsEwRVcQWyca6BWD+GtXA+4oA
br2aAAFrJH72D7LO3yBegNn5TBGhQyaFxa9jaoe3dkJb5mZMMcjQZLiTr2yQEEV2
u/A77ZyYwCQs/9enVNaW2ou+X90ROi+LNBdkcwrN++6EIGlG10oNoXcXtHd7MKVe
vGa9Zl/UMpe6yWzxq8eJQRhkrpgh0T/uySEudAe8YVkU5fwlKL/W3EtX+LRRykVR
3D+GQYJBEyChe8LU3BVsZ1h5ZA9zd6xXAhnlreEvSKTGstcuq06bUSiziysm2nEp
MNVoTEvHrRGLsyDAWBVnaLDaZX/U0biJ9AUJxiCb4gO6aP/362rKq6iJC31/b613
f/A8oK7MkTdljz+2lCfsJxfZQbMO3GDI5Wz5iWkmGT0+DYp4uiNvs642zXkgUHqL
686F3eRU7TL7x96RGUL7o4GdGjdgoKmfJidLPaWa3y8PsHLi4oH2FMIerEUxfol6
9aQePNkVFm9s6MawAAlsJzvK3hfZanw8NHTI/tfeCVohV5qLHBGfTRPalDoB7zf7
nM9aVVYkR6cTHHpV1gEUWEp1ny4FlQe6h/WOVe4egtGIUuk3FjaNfGudB/qroNt6
JJPAyYEsB9MB4xLhwVuSIkjd0+vrRJU1VHKtQAi3RU0Oew+pKS1jshb74vQOwSiD
WacsCZ/bAdksRkWCnKXY9l5QdBrnuLiSjWGbshaOItxHdbRjDaWFxy3IjQkO+ByN
yj8w+/GbKRCK9tXcPXZY5z0qoSc4fjOnZl6nZ/8bcRkalFlrL0PWDkjwujPvTHcn
GOD5d7YjVaN6Rf/X1Ab9Bt3WrD40bQCyv2ibUO6ldhBD9iMzNj7NkHXddVlX2oRh
L9ZdV1l8CfjO+wUKsm9CC/8HZQmqeLh99JAMYcL/Qd0eSWN78t5pkExua0eYx1AY
alRGPL5cPgPPlRgLsNkw2oBIu5KkBb0GA+VfRqDad7Gx6HsSZv4xLpXgfHsKVWkv
/UIsogL5TcQLqUrAfv5PiOTrXmJBihjApRuYaLHB+2UatLhSisTqNdXEIpAflydi
6dE+kBsNW3/qvUWh2MQvdWxKfodyoB7woDNv1Rj0nFMiuT9cDVx1P/uvkYZhXwa3
g8VbLRBnJGyFWwHdLwdmQOO5+yYxnBXANvG/eV8sjIYhxGGFgN9EssQOY6WXHYQV
Hb5O4k+RKZ5fSGb9RKGT51bIupiahUWbVkEcSW0EB7ZaS+JHG7LpQddBFP+ufCW+
8OkcFKMZ5yL8tsiVpYf98N0KLFUs+OFRteHWWEUk3pLxrwN6f0peKOyepjNSrc6U
wvlOwQ/15cwB2lbnzW6azcEG+xVG/rD4/9NbGPtZkGb02TycbqtNF7RoX4XQS6MH
0vLJFmgCVBMqMTgKJpFA1/oxWbM6XveNX1Wm4ONKCnDCrUiBw3zgu1RvVo6BVEdc
WhxUhoPAoIKHTrsv0r6eO8fSG+/MU3W3+ekK1crHIiuSnZUPC7QKAXsbYq1Stp7+
btM7dKGAS8ri9oRCJXg1RCYiCjuPhE8OTHmX/v/H12/PPH9jk9Ztz7Px+bzAnfdE
vBNwJbHWL0jIi6vJcGiWWMP7RUNlqhHgRxFYedvxdc1Biuzkb8GqSZ3adDzWmnZ/
xnJ4noHTBRKbwJeHUcjcyw==
`pragma protect end_protected
