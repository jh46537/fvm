��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�y�Sy�;��>��&�MA�)Cʌtg���e�8~�����=H�9����.k������U��U�Xe���M�b�(	
'�m��_�S,(
>ɢ&T^5�[Kم~�WA��Mb�c#�<˃#:}��6͕��F��O�j�7���'AF�9��'�ƹrq�9�p�
o�'�w=��v��("�|��ӏ�I�\.�V�����)���cB�չ6�t3sꀚ u?�({��_x�W������!�`�e�H�H���|�-�YY�
ꆞ �Ӟ냨��e���S�kFd�v�e����y�*D���G�>����+�ᩜu�f�x�I���*��/1\1����r�2�*M_�4j�t�'{)ȳ:�A��!���ש��6�D`��Js�[�a�O[�G�O.�����}�9�����E���;I҄0"}̙�������@pi?%D;�4*/�asnq�k�o��Ѡ��+�tZ�h��EŌ�����A������$�5a��k&H�w�'ș1xB��&{X.�_�%��mƑ��),���ñ�����.�����%�"���B��]F4��Wn^ɍ@YC��C�Bﭸz��#�VyMn�3\�E?T2�;a�����ר�bͤ?e��������Y�Q'�Vx2�>F�����Y�4r? �����P���6`b��s2�s�z���;��^�fz߼�S�T-��}=�[.�G��M�e��P��Ɔ�j����������3��ͳ�{?�i�`�
��&�6��*��<�������ǜ�,�<�4��&���A���C��J��/;Ȫ�,�y�l�q�.R���렖��$(%���X<�x{:��9q�Cg*n�جQ.�Th�I�c��jI�����7�0��]��rMQ��Ē���A׍{�����Iu�������)��޿��ާ5Qt
Md:r�_X�<'t��@6�P���&6��2����3k-�|Ӑ:�p����L���N[����K�>ɵ�q���A��8`��R�k�{#Oq��CU�RHj��EӜ���i��E�Lvd�R�ʯ�N%S��*%wu�O��#����(�:,M�^:�� ��H	�c�y"��>��*����:q��nb}�3�zV�p����ʾ[�Ml3�t�� ���a�78p���� ���I"Mhx衉�S-���H�Q�R�h/�E	�e�k��s��-E��C����:�����	*���M��֙i|�)�%�*jƯ��4v��M���aj!�&�惤Rf��e�9J��D������<;�Y��b�,_�}K��d�}5�v��Z���Aq*�P碓j�@r��g0��\��(ٯE��X5~���4���eB���v�����.m���1i�0U{��}�h$[�Ф�1�tc����l�^yw�ٷo1�\28:/bc�Cѝ@2��^��>'���D9�BB�|���{&��<�ڽ�itT�ex�����@�W��3��U��b��F��ьM���УN�Z�t�q 4_�ؽ:Ft!�eJ��x�/�ni�b�7��%,�phZ	\dS�w��MٛFi����[y6�o����v�	�KN���)P��^3��NN�/��;!}�(��C���M��3�y��5[Yԃ���*�
P�6��5�#,o��>I��!�n�c�:��,��2w�]�A�������;�Ш�Y������S�0{i�Ҫ�wm}��]����4��Y�����)��4��_����|�N�����[�d�%xK��D�b�n�%H������H"��*�.iG�=�;�[�ܫ߹K���ϡL!�f̥F��_4N:+B(�蜸ȃ��?�����A��A,�Ij��\�3i�uKeٿ�
�CF�Ðt�o��Q�8f��@���7����@�	�r`{/�HLf?�R�t����
���\*�	��}�����ko,�
aH,xD>�J�}�Q�K�m���%J�k�8_c[d�J��J
oU���v�FJ��x]K�PMU��p����q�eZ����Hd��<��])ӏ�+2
{ه��Ж�O�� �<!�/ni��W0I�K�6��NQ����/�E���.`���,2�bfXP�E%��N�b�[8�!y�+�[�@d�3x�nKSҳ5_n�73 By6ym؟��O�Q�)�5A�Pbl��٧�
e�����n|�Y���J-�5侇D�������ո�|�)Z���R���?�y�ꌉj�#l^b�X�t����k�F�p�����_�yvs�*��0������k��81�֑Ԩ5����p�n0;>T&� ��!�o�hx�k�c��d�ˁ�:���?��H%7�]��Mm%$z���-k�Q$��7��O��E�3�����2��ab_�bb�C�H��˩����Ȗ��!��&|�/�����}��r�U�3{����xM4���c��k��w�f� � ���B7C��Fy��L����(]p�å��}�_$@�òw���(�մ;PD�Ro�˪ ̸1c��n��5�D+J{�!���@�@�	��_��1�փF6���rPv��-ɗ�=\2�_=�j�A�f* ��K��p���չ��U��@�@�V@��k)E�iG\w㵼�Ľ�����&m���X�Ǎ��Z�}�b�'��!�Y�o�h$����U��.��)�}��MC�kv�)�hjs4�3�NR��K1�__6y�2���n�mT�$�MusH�7�%\�J��Շ���̿O�������H��
�,N�x�mg���M�|9l���Z�� ;(1�	������r!�j���G� ��^�C�A(�i��0��1g�>]꣕SƼ��Y��d�W/A�UK��yE��!VN����p��BL\��|�|S'����5'����DO�֯�)1�-��#�T0��9�h�R�A��/��@,�xx�X%�Ql�o�(�׾b���@2{V�@�w/�n_ق��d��+9��:<��Zc��)*�y�yO� Ҋ*��W�SO\��Ļ����#nEp ��K-�Iu�m/u����`��!9`���x�=���Ь_��t��j]�_��~���=~��~�1�k���	z+���v��%�Xwm�"D���q~I�.�6+
 �a�Q��<��M��۱p���(.��;�&�����{����O͠���w�+�ͼ^^�"�w���A�X�@U�Q4ԧ��s���R��(�����$�λϷ��H��+dX�{=tW�����B��䄝��������j�g����q.x�ӏ�u5���@�θ_��Q����P�q>�Wo���5�~���`6��D%R_��/h���5m8F0q�C 0��`�@�=��n��a��� k�������|m�	R1��_��;���ī���Fn��o�gM4���.u�A%�1�d��+ӅP��ek�ڴp�/��8^����	E�zA&�L۵}��k��4!��w���)�F�D��5���9��TS[0�8�������"v��mZ���,H����#�R���C��ddC���%�.�.�^���i�u`�� P��'>6.�pyK@`=-���esX`����Z�bg���ϯ�H�a�p���j��kw̟��r]��	|w�Ȏ&B%T�x�0ʸ7ɭ��>���?P�cɕ�n��Þ-���!�cv���
�q��Z��L�G.�U��J�]m��z�
�j�@o|�kK�[�!���.�$;�'!�ۉ�#�,�H����ws�g�@��"�$�k�¬�V���e�e�r�kBZ.<���X����=�l��P�ƘY����=���l���R�����]�SB��=�q�Pɤ�����+9|˜�c7r�Fq��G{i���s�|4PU��z���'t�C���)'�a'ab�,��WΏ&9�N���ӕ���� ̉�\�vz �o��񨈬;?��n���[i�/���
u�%ðz�k�oT����F�cCE:h&�4�i桪��F�%��N匀�{��H�(��`2�!vD�N��N��ү0A���-5Lz��!�����W�ͤ�K��^&��5���:�"����]z��d�9���xi�w���5!�h���vfn��~ӹc_�r>+	��W^��pf�]�	��z���8�ў�xv/*��ގ����Z��yӿ�bK�Ύ���pz�����YT�x���0��c4����81m�`l���Ү|�VF���#5W�sEx�q�d��	C�c�U�xb[��(>���|Uՙ�(�{Y���7�C�����n�N����ƭ��<U���������R����h���X�E�<R9OK��P.C�t��x'V�4]��� _�+M��A&�m��5tg�]`Rߒ�ϓ<���@y�����6v�i��2Ѓ�t(���Rrw]�"tGa*�q.��R�(Cu2�@�r�V0���z3�2���`�ɩp��̈b�Q�ϑ�Ke�Ϝm��+�#��&p�"$���壄;�R#RA�:,J]&-�<�R�a������UO��@j7C�|��/�HE�]����n�	�d�p�i���EK�uG������v'�Z�����
64�D�:�'�@~ю%�)�(IQ �a#mo�"Mvmf��ӥNc\"u�wWŪ�p�<�`�I���T)�Ө�nM�]��lޙgyɡ��Y�.Z)��Z�n�e\���K����@/Q�a��T�R�PI��5)%�Gԓ���[v7�s�������yU#�`���ħ���W�X�=m�
��x���/L��ڳ�qZ���#�+Pi�)sS�	��>Bo�����xI;!��Wq�y��|gGᷕ�@t��tݓx�"-��j�������R,ݟ�2-�_g�I:������u��$�1��d�h����7JFB��f�ǂ
Ľ��tJl�'�׹�%���y~$�#Y��-p��-^�X)�s4CQ��jR�Zc�m�ᬅ`�}��?�?%���*����Y���� `�΢�`��)R�d�Evf.Ju�:�?��ް疃�/�����ᦄ&��x�6��n�2�kp��Ao?N���?Qh�,��(�0�L��c�yf�/�Hl�8B=��F4��tk�������e��C���&ﲕxv\ʵc�1��v���A�.rsf�5��J�t �_�NԤa�Ӱ��!
���\��
ȞZh��*mprPo�N�SS`c����UM���^s�ɍ1��~��+�I2��h��t6J�4��_��x!�wU�$b����먯Gk	twĶ�Tv�^b��)�u�S���pj"S�N\@���}����Cm����+�i����O��)�����Oq�/Uӓ����������{
��.�~�4���4�\��%��Ϙloa�`c��$!1�%9B�wdy���[�(F�C6A�4�b�|��gK������g�rR��Ae�x���}|S��:��*��ʏ����f���YD�H���P8BЮw7������Z����~Cx��ː����g��z#
sHX�*����z���qԬ=A����nL��e�����c�+Z��@P�I�C�8a��g���#,��� �<�Q~����22�G]�c=��9�wC�bn��e�AS���=
D:5�8���]Y�_���N҂� (E&�JGxg�$���>i��PìP� �|;q�ڝ��������fP\Ӝ [h>nX`��/�~�O�:!���ϔ
��`�>�v��1�<beP�f��ͬ%�%�v{ղA�I��(gc�|��1𔵞KUeR��#F&FLG��/N���:4l�3�>D�j��-8�7��۩u`-HA��U-7�������2}��#�o��[(D�Rl%������g5ӓ��g5�Y�R*�fY^��ͥA�U����wirP�[-.�/����
���������Ũ�U��I.OS'Jw���>�G�e=��܉4Sݗ�wߴ�r�`+��RWa2Dd�-�IeW�gڔ|��a�ad�9Rj�"���aU��ȗ�OQ�E�{�����;L��+�\�^���
�F6w�K��;lF3��ht� (H����\�3iި���t���_����9�6�T�c�P><
4Ӡ0�(y��6 K0K3�؜�I��'o~ֶל%s�}�2R�+]kM���}+�nE
ij����{�_�ɏ�8 2�^��q��ֶx���<)��ֈ�vY8�_�sW]�c�XG�����ʳl�Q�C�쫱�y���o(bS���'j׀���~�	�;���{7�.R���m��}��I�C��*1�Q�>9����nF��]@5�^$B���^��>�,����1Y-y�Yi������[�O�Ȟ�B?_�?e�Z�R�D�˧|���xgS4��d,YB3�/�=P����8�?3W��)�o'$)�]�)d ��+��<�jN�	B�9_%FǢ�o�����tMn@����VIo�BÍE}a.B�haZ)cgk��?���b���t�@^x$]�c��1~���!�:ko�w��7=�H&�X���pe�����"G�xG?L�Q4\��J�N��ޱ5�����TY��!\܅:��L�T����p�`��������{�1y���s?���h�O�b[�y�j�'ZE ˁ�!�����v����ooZ?��e�K퇍8�ݩ�tM���҆�$�f�CT!���h�����<��&�h6N��EZ�{��!^�}��IX�J�A��%��ž�Z��7�},�7�������������v)#�O�f��D
򮷿� wYI�+���.�g��U}(3����~^�ɧ�^8R����4��M���i��lV�L��ە�=� Ό d1�s�א�� �LG9x��ś�s�kc�"I�-m5�V	D����8�I>D[V�t���.[=H�G_��'�K��k&p����!K$%ř_���:�� ;0�1"�e��=0���3"�NH�8�~�b&�3�w��FΞ2Y6�hc�R�%�{�K{�4&��M>H+Ik���%.�V0ͺ]xQ�L��`���
k#�+��?yPj_5i���&T�">2�Sn����Ԧ*��)[�,�58��G�;;�S��ת�_9�{}`�����Lƃ���kª{:�6��o���D�ř��u��쫣�]ɵ7Ug���u�-r7�ENJ�D�L>�� ��}x|������<,���������A���^��ڙ���:%kP�
K)�G������n���Aؘ~#6�0����=��I��� �AI1�! �_���������߿���f�D�)�WԞc7����ݚju���Ws�Bi�G V!������1-��B�#\V��KCS��D�|y}�Xr,�+��S�!���I5��(m��'v�r���� .׻.%DڲC�2 ��eclԥC����orZ�<p�=��T���:��D=y! �U̔��p��h/{�(���Nh��X+��E���"�pw��1ߍ�4��4\��60,����Z-{'�H��m�݋E�K�2�{�T��UX�!�m���[�zd����5��	���L��>o��v��z߶sO	g�����e9b���l�h��ջ��  3��,У���Ҁ�T
"EF#�����O�^Y��mQ݅���bo�bt%/��K��ᕩ)��"΄&ZV4���'�%qcB+���>��G��r�c�a�t���]L/��"��8��=�˸>b��_+h� ��y��%���v�~�'��6Ǫm��$�RP�+�P{-Ij�VO�F��Hqm'L"��K�eܯXF�)���r����
�]o5=��&Ӱ$�o��^4�;I�h�^�RLu�.؉n�b�����Y��P�!0�m�R
�	z0"k�1�vړ�]�����d�W�)���'9ugE�SxfpTJ�˫����1��5 �hm)Y,<�(���\�:9-������!2B&X{��N����)0g:�:�Y�j����P��J�+?�������t��W��^H��} ԫ`�B��Çfi�0����e���I�a6U��?4N�|�ލ�̘�E���x�,�	���>}�ټܑ�csI��H(�C����yR��-SiuZ�Q��h���5�Jg��s{O.� ��n������NW�zOu-�Vj�f
r99�O�p~��͠�+�C]j��G���Z�Ҫ�*����
� ��r�c���@(�)���xgy���?� ��E�@�k���8����B�{vh���s��kq�C��v�o�!�b� X�S�<��wY�e�Hu�t-mZbl.#?�9�����R�I1���Mb�� aaSR�C�Mm�	����=0��v2m���괪�}�A�%����O�^�~�:su�]����4T�r��h��5%?dcmdB��I���"����t��ǹ���dA8�/���Z�\U��l���F%�P2�dj���Ǭ��>\�Oǿ(�]�� ݓ��xs�t/x�9})IR��ŷ�u�!����d��;N�c ��"M(�D1��yJA����5|�cE�oS~�O�7|�v� Θ��,]Di5�����s6:c�db�A/�C��ȍ}���V��/(���#��7Ջ����=��^w�B�a�ʅD.c���D�78�\�v��˙�j�����
P�p���7ʐ��??E;n������<��{iK�p�f���	BU�,�	<����e)�0��������XV���NM�{&�#J�c$o�ޯ���[�q]��
+���Mj�(��}j��7/D����j���Y	��xɈ�.��~����}�^�;	�a���H������ڙ���˸��~/8=�8�� p0&�2���Ta�Z�뮴��i}���-A[�򏠘V.��x�h��ȵ����	�~���F	��p�j��+bWB� ө���D�Na�C�hq��]�]O��:��v���뚔1FD�=�G�ߊ��*jG*$�F�4�XH��ל*�D�&TFOV� 8u�*���G��(78K������ٸ��8+�G�u�K�xG���>��:��	jk-�G��Ƹq��G'��4P_M���c�[�2�&��\f�]�{��2��e
k�^��3���F�c(�5��+�ӚHc�QXN�� ���>C�Z�4�M�_R25�%�q�k�A����zC�7�Be���	֕���'ȶ�ȇ(�WuS��O:���)�=���/���CRD��d}w>���2��C߬�t�Bq�c��=R|!`)����}�����@��b
u&�ZְA+�vRW|ڲ_��G�� ��M9Uj�'�v�'&S�*����L���׎�5	Z��֊�E
��q��j�J����.�����ro���t{7P��D��Y��-V��I�Q$`����s-F�?�y�J!��_x"�+w EJ�]i�u	�����od������X�c�lХ�=*`�L�7�~��C`0���J9`�(�ؤ���q)i�]�g��N7"�?lH��si7�C�DXuj7�g���$���a��Q����=��T�G���K�_�+�;`#jK#��8)m�B��!�Mo1��pK
?��Enj]������בRY��p)u|�Dp�]�^>DU���\nh*�ro@�v�R�|�~����@	�����蕪�5���͙[�i|aI�����_��8ӏ�+��H����?|�zLœ��ԯ�`���&,�=ُ>��N9���O�鈴�  ��S���C5��j��/t��U,tW�r%������,D��Ò�aa�>��o��w�&ȿ�.��` Jc��r�m}0��M��Z�8Dm����{��k������O���˂k�c�A�;��=��V�7�����������L������"��%���6�~\R@��b�0.Yzm���]��)����^�y��,#����Ų;�̉G�d22V��x�t�|m��ap��ZyTmi7������e�[.A��%��x���A�qAm�8� �p�}�`���|d�vt�Ð�6v��&�Ƶ����`;�ZZ��'�e���f��c�}#��#x]$��&~Үhs(q��$"l�c��=W�cϾ���K�}��M��zH,6�Q"�e-�	.#������e�d3�ھ�Pc'T4KuQN�i�B��Ф̵)�	�靊�����/���j�l�����try�!M��op�)�Dӣ �e	�ae	ʄ������'#O��J'�<�QK��ډ+%Bg�u��F��A�Ԓ�'����R�nL�z�to�hQ�4:�W�m�jڃ
���P5�wQVm�2c��?H�]w=�.S@{hó�o�P�.J�9R��+��~�m����<X�bF˺�1��:ڏz���N��Qͱ��.2�˦I��_ضC�0E�����L����m`|Qs��L����ɸ����<��S�U����'��z�p1�L�҆�xK�/��P3�nU?(�xq�\B�
f"kg��Q�s3��G��y�W��h�|��˘Dv��Q�Ƚ��@��ұx)�h3���RםK��i����a���@��P�B	�g���pl�t)v���x"[�wа8�q"������s�`�˿F%� Wb<������N��oN�����(KH�i�����E����fB��������/��eb��<ۜm_ �$捥vҺ���)�C�d�.ءyt>	�'(X|<�����f�CCa������L�	�9��d[}��/(��;�]h&Z��h{�tV�b0�+��@)Xc��r@g����Z���M�p��WXR43��Ă�"�/��ɹ�>���@���A�g���������2�m��Q?����nh����%7��ٸ��e>��a�}�K��9#��>�Ye���ȫ��B��n�D����3gJ����
s"����X^iF_�e�ZhTyY�L��RTy�쌝'��G]�S�8�ۓ)�9X�m�aG ��	�-��!�H�~GK� )��_=ܻv����Q��!z<�+n�毣Ѿ�F̕�c�;x�@^�xb= ��f��H�]�/��\Ӄ�} �C�?�o}��7T�{fJ͗��QO
�a���̳�4���Ջo+I�Mg:�90p=!����� ����-)Ȓ3��-]	A�uKS�́��,O?����OK�F�Ely����%dx��	r��Ϟ��)f&��Q�푝-��� ��'Z��;���j��e������9��".>"�!v,a���}�/HO����&O�e�;�!�Q��e{�I�� ����H�����U;M�ł�y��w}W���ͷ|������b&Agy6��zT�6#��>�7j�s���ы
�]����
��^�İ��N�ǅ�6��<�O�bO����!���]��d�L
TGT]w4.��]w�i%��L���ֻ!���P#2�lK���f�C��o
���{��l7l��6�Q_�c�)�л��qނ��:0\� {���+�ҳ��a�&�<!���7��AF��Z�dG�@��w=���l�墟����G;��������BȀ��}jr1{�d��)s��,�J-��σo�C����_6��;sg�1����,g������/X����;ʛ��=!3@�P������NH��*�~,*�;�`t:� ��x�|�L��Μ8i
X�	l�8y��J����񊒁4Lyz�#��Sˌ��ި6w� �1}n�kD��j?7��jŞ����uօ����n��Z$F;���Y[��� �g}��9K�����s�zao�嚦DP��2�PĬZ��S�8���&����o�ӣ�-��yU\Cנ���0(s�E����ܰ�g�߼Ex���3��c����&%���x���q�����1�G����>�+�gX��=�Q��[ a�J3��}k���	j}E"�߰cz@mpS�:��D�r�EGɮu�GI�W���P"!Q<Rt���q�T��;:je�y$�T>uV��{�լ�~ ��ˤD\����n�XA�HS`�b21XD�K0���Cԅ��ɀ7��B��W�%.1@#O:�v[�.�o�3������8��)Y��,�W�����IL���b:q�٨5�|KG#W�����iZ�P$�?����C�}�;k�+
�P��N=�s l��}�Ǿ� �f��r�uN�U=�"�d}r�U2����c�c4���tت,������)��|�o\�'������T4�k�D��\����T�&@��h� ��.]���?�����!��_��o�#�g���	��N��R]L�G-�k�GB/�V$�:J6��kU���dRv����S�(@�wVO#�	���G��t:Oő 0P�6�;��O1��s���y,��:�jz9'XM}w��@��!6��O��~��*R�m���q(V�uD/�i'��;��W�ϳ1Q�g�y�v�"��@c�4t�{Yt��q�����
`\�e�������R�f킉���X��-Y:�b�N����|�yf,Mq��كy�dЌ�q��cl�Ks> �uu4�蔴�H`p�x��\�N��~���q��Y$��G��h��A�䏻����/i�\q,��{`�~���+���S��h��b<8B#��E��C��M�Ia������]k�����/J���S�������w�R�/�`Ы���$���Q~8�.��^o"�Sf�z@���D?��9c��-9��4�@B�4{%0��'���'�b�R=t��{64i ٙ�X�ۼH9��"`+Q��S�Xh��(qm;�U�9rn��Q����H�3�f��w<��v����[.�?}(-�>��m�I�^�[r\4�#w�EiI�Ml�.���/��cP�qB���9�*:(�׮���wHB^����чN��f�u A�,�	��14f({�1Θ5,�e���<%$�d�K(�m~��TZ�s�=��$�<�q�K��������L�46L
��K�K
���v��)�Zv|�L����	����5|�1W+zrB5!��[O�@�e6�.��!s���5#C�}�����u�skQ3�i�%K�lA-�|�-�2e|� &t[$�G�� �|�+�P<��[�pG$YF���Q�r���q����7EJ�rJ��Ʃ��1����yG��� ���lC���g����ʭE���\���(X���O�' �:��4L;�<rMqs�s�42=��m�@���+�[>�%���k�
}���A�@(p�'ޣ[�Bb&CM���,-�b]�sv��ZǛ�m>�2uq�F����L�2~�w�R�W!"����:6�����y��(l��ȝhŷ���L�G�����h��	j~�+��+.��=T�aj��gO	��K��{��>ʫ���ni�޵�;HQY<�I��2X~ ��F�o� �3�K������x	lG���R(R<�И@4'���.����%��O����!.�6�Ԫ�֭�4n�{"<Oa�ML9AVT�[#:p'�t8�����bn�0��dmq�����?��ߛwD����Y�K�6�S�[<G����q��SxĹ5�z����I+G�
��>P�r���Жׄ��5h�O���ҍ�>h��}��&�\�] ���͕�؃�~�N�Q��J�%��7_&�Ǯ�)C_K��z�p�W,�J}̖��OF?�N�n+�e:����[�ت��H�x�-���I>��i���۞ׂy\$�'Bt�7-{�Rm�9i��B��ƽf���{�
��	�ep:=���H�(����"�>�h]�s���Ta�ue�=edJ����ց��p�>�G���ǥ��D\ZD �a�:�����Nk��~W.�_��kvA���y�kfCŘ�{���A�[�.��o%U�<F��Q��g:���{�*�<�9����)8�C1�sv�P�2�������a���3�K��>���E�˓�����Z2.(Q!!f�<���*o��B�Jk;b�N�ïΓ\G�ଧ�4 ���%���7
�e���M���ȝ
���.��e��8�b�!8����ec�#�~��g�=C��m��X��?�蓉�!g�����ru:�2�}��Sbߒ�J��VQ�\$,!2<���n���`{қ$$�Ķ��t�L���MsMܭS=�(>�3,E�B�
�0�1-�)UX����;�!�O����Z�fi�mL��@Sb�=���jPoi@�x�6�H�9o��ﳁ���aqbu�׸@�|�Le� C�bE� j���X��a}��x9\g|���Vj�!+��M�"�.�۽ �c�mؙ�C�Y���b�e,ַ����&�!^)d�gJ�9�<�^^��nG5Q��cLFq1#@�R�F��� @n��KY>]D����'SS�6�]4ˌg9�:��3l?�>����Z���u�"�ׁUn��|_G���a�1�~)g�x�D�BW�t���I�욞�e�Q����ʧT������F˺�S�]��D6/x���4�6�4������x-�4|!�QZn2��b�����uO�Ir�J6��)��	z���?�!�yUpJ�IW I�u�=9�᠀�M������Ut[��@�0��$��|�ń�ɇ�E��d|Ԫ�� 8/����B��[Rz��BX�ǵ����`ߝ���-�؃MZ�\W��CeG��Md�O]�-�2'�S��t�k~)G]��E�F�� 7���I�3�ե����?)�١�Ѩ�3���W"�������q� �]^�Ŀ�3��<Dlf�v�\��zClf�X�A0�@l����f4��{ҝ�?��I�]ob�TA�����J��ٗ,%�s+1f�ʡ��d*0)Ҝ�b��)T����K}�?�����7e;W��E�&�;�6yJ�fa��5�ms�����;E�[AN�2�`zwbh�<p��Kـ�}���=��)�E�R84�^�G���V�%��;ɑq�[R�Ia�1�*��cy�B���n�|��6�?�����i�I*�Q|��-��N�Ɲ7�N`�E�H��6�?�n#�D턮
MT���Ķ�[\�
�������LrG�l $5#�教	*2����o�t��ٿ�)�8�)ؖ� �z:%���H���Ʃ�:Y�:[wƨ�Qj��
&���Y��H@VD&gu����v�C�ǔ��U6p6y,��<A�a�r�A�ϋZ���e�A�ɗ�rL_�&NfV�2td"V�1X�� M����-�ۅ�#��F�
�ōU�tnsӋ��7��u�����v����c������a�i'v�^h��x�PD�m�9%�>O���r�qU�kz�3<����Ȋ�vLĥ42p��r�}��F�u�����F�W�#�˱��	��#����O���β��*�J��ga,&�}	�|6�_PoQ3:�PR����)1@fE��M#��dG��eV7�w�q	�o��NA&�r�q���چ�P� ",�.)��ȁu:��.��
�՞/�i�"=OzcՃ�1I�J~��D�D�  Y�lg:�-�*VDkU�W���[�:;��rV]`�-.�t�#ok�r��`�S*I��O*���@昦-~b�]Kh&���,ӯ!S����Ӿ4!%���k��̷��Uܔ>�U�����.���S���<B�:nra���� ���T(�xX��� J[�C!�q��DZ{<�-1����-�0�t�y�z0�)dKTT��v)p�X��������q�㘯+���|�0z���\���j.q�@����+���5l�c?O�s�na'g��2�R[a�u��Y����A��m#��o9/��N��ti��ݯ�,�q���+���u�R�;�5b�x��,��t%���m�=���ə�?�衵���Z���@`)^�.Y�eN�Ux�bOa�C�Ş�#ӈ����U�g�^�6��&� ���{����*@�WK��p���OE+�(j�e��3���HEj%�24�	��)Ƴ�9?���睩.j8~�]�և"R��vÞ��}Jۢ$��m6�ï�_�|W�>�1��29���M�-1��Շ�󄫔��#���oC���}��KbkIxmu
�\lz�|�DG�%'|'���3�ʻ�}<�_��$�D�E�	ֲ^�jki��,�5�7A[�QZ������[L�T	ɗ"� ��-�R�gN ]I�� #����_0��;B��-2�Y�<�#W��H^%k��|��aUF��@�lr�kdе�F���}���B�c%i�g�����Yx�5#��/� �2.'�]�O��N��O�t��FqWpd@�-p�GIOw�`kR�r����*�<��m^r�Mp1�F\�;�r~bh��|Q��swaC��`�i�pu#HK��v�����4Z)�<YZ��xg��p��+f�����R���^f�t�����XG��[cY�����~&���y�IFotJ�v����|ձM�z\�=��.g����(w\6������9��J���Q>�Y
i �����^����1�i���ǑyF�)A�f%�/ݝ�a9��"�Q{X�#�Hq'�$ҥ칀~e��(m.�q{�<�$,3	\�F�e�m>z*���'R�8͑��n��U,[Y�H�9djs-}@U@���;e�wR{-ic�dѶ.�����|{�{���D�U�i�W�* �r#:�J�9������,����|�M�~%n��X��u���k��^��"�%�s�"�*�dR�R�o���	�PBSf�4Nׂ7�R��C&�o�
 x�� ����-1�d&�E"T����jCi�5�6������AB�6V�WR�F�b_uc#���a�r�oWh<������mhΞ���_�Q��1���v��X����l��)QQG�d������[����h_�	�"C&v����Ί�zԨ҆�uoT���Y#H���\yӿ��AW�rBc�=�	E�h�s�!��c;� �~y}��vPm�&s�rC֔D8�o����������C���IK�ģ�{ufSٝuR
N�]����4��X5��<d���qG�#��j|p��Bo�=�r�5� ��lܧ�S�A��G��O�����X}�&Rw����焴��������v�܋�c��S X�"��Fxe�m�r�3rxb��^2�_�2��\ك��K�-�:�����#���yWK%Ƃ�Cv�=]F�+�,�1k��9�+�r���Zg G�V��6� ��
X`R;�Tkf���
S$.� ���fw0�Ђ^�$%����G��,WI�xsm�B�{�Ι�Z1���%h��M�;��EO2~�.��Cl�u����K��O�/�����0�K��6B�-k����n��^����[�����}Y.p;��ͽm�c!��S5]�¨w�(�.ΌK�9�����a�u�*ߔJo���rڿvj��U>6`�̶g�	d�)�D�?�ᓉ���h"�J��Q@����cꇍ�ȷ��� ������r4}g���C0- �'�����6��p�kS���9��b�Bk	4��Qɶїz���L%0���N� ��I��`��3 �u�h�IE�CD�e��;c�����w�E�K������)`�r5�%�7D�N�DYnY!�s&���"M�������&K��O4j�s
s*����ǡ�"騨T=
g��Z6]��f{:i�Z_��THt|2<�/� >'�obx�@2d|�/AP���) �4��!�R��1��F�ڢ���/SȌ�&���X���Ca2�x���ew��>�7��}���Ҽ�g?�o�yg��t�%�H��`�y�P����dM�k0�3+s�����s��L�by��D;؍Y�I:gQ�GɘS��͉g�DW��H?��HL#�^U����E�P��x���T���S�Q�͵��*��r���W҇�ϡ+��/���V	��`A'2��LO�m�W0X����bO����iԤ��Šj*W%�?uUb=�H?��!	8��z]���O��A^|;�B�&�6��8M��0���>�z<o��#XlP�������UЧ7���N�+���-���1��iu��h��dLv�f	��RE#�o���n˗��~�s����=b}hX*N6I�=NOlA.����0c�N�~� ÷�Pt��s i��y�G�'�MO���q��V��^��=$�P�uef-tM|�}q{�S���NFY�0�d�x�x{~��B��M�[,sz7�p9n�0���ڲ�_P����ץ����;�0�e[u��{��^��L#�H�A2~C~[lH�ӟFץ�nE@ín\��(�۱?��
��Q�ѱ`��@ j?�M��j�ȍ�i۵(�a<Ԅ�x,��Ae2�R����\.&	���R�H��qYY���<�D��0�����TՌf�i+.��gO<�h��'sW��*��>�7�)_��i���4@K�~�{�������`�5�/��(� ��4Ya���'�Ը��fC��)�$̨x���-�a�(,�o靎^2�:�Q��C�m��xj$&���_D�C/�� ���W�aul��J���v�+҇��_� ���A=5r�X*���g���!�K��ْ��Ǫ�g��bȗ ҚY�����Sɧ�N�B(F���R;��[c>�-]���Z
����{�[SS�r3F�sa� ����iʓ���n��W�?�A�^���
]^ͨ��ך��<D��)*^Y��-4~�*�M{�?���/����`ƔI���e��w�9��[!�B�$|���)�s�x����l�Hu�ŗ�q�����e�N=+���7���It]�G�t��F��r<�[�|z�	G��D@���H��{R*���i����C!��2R�/�����	�ed�5\F&c�>�vKT��w���FI�-��!�Z��ϕ��%����ߎ�8�v	�x����G��L�����G����qD�/�*ŏ�70:_o.��Z�{����X�����G@�V�F��-�}� aFp]�1�$p������ȗ����M�F�m7>������#b�`��N3�PP(G{�n:�@���k�$���R3b��i)85�o)�N]�фe�U,���WO�!)�{u#W3s���.���8�!]K^�焮'a\��d��$��+b�S��D��N��B"��é�&�AH�`������R��	�y/�- �Piԙ����IBw�Gq��͒@�e�l2f��m����[�NoHc���IX��S��:.�
����1#R��Ds��
Q[�H�Å�<��>"��|��<�Bgr�>�Cd�N�)�WQUw��-o��%���s�`�i�Y�D�m+�e�}.��*�g?f�1��!MI:��D]2�L��s��
��%iB!��sDkބ�y�
�5�^N��	`u��1B�ݽGp���-�٘f�ي�L(���tc�+*O-p��4	@�HÀI�8��}?@�5�8�4 �7��x�r���CV���)��EY(*Bk����̝�4U���9\y��U˘�`1����)�@V��Y=i��q(�ȓ�l���Q�X�6ɯ^pL7V�q�U���4��Ӳr'i�'`|��V���f�B�A��0�_C|6Nu�HZ��(�������;�`$@����=�\lG5w�h��.�'157\M�}bҍ��{a�Vu�]8��vwL��X��=vp ѱ:[W6)E�@�Qf���i�'�Re��q�����9#Z�*r�����Cf��x���%�d*̖ zh�����G�h�j�K�^��栎G�U>�꨼^�;��J9�8�U��騬<�/�*�ɾ��c���`���q�b�� p��0Q��tܻ�,��=�p�����PHk����6�{,�dQ)0/̢$��I�r3^K����gӹ�'�������xi��x:o�@�����Þ@q�Y�6��̜�" �Q>\'������X����9Ƕ�}ۿ�/�%	���s1Ь�VP�>0i�:��"�|V�>;�<)ۛ�K,ݰ��Y�ۅ�t�u�9�.���PG
J�b�]�w�zA�{gR��ac˴�RFa�p�Ԯš�����c$���}��ݢ%�LB"܎� ��Y��	��J�ƶ�<���I�t���H�a����`���#{.׎�5/=3����t8⨂T���}[DT�����s�����ͻs����k�G#��,�ϋ.؏=�0(����P�ّ����N������´�R�E�� f؟�AN��Xo{�V|�����7g�tdY/Gf�m�(<�L��!��G1(ߗe�C\}�yO����=��V�M��Wk���)9)�iL6�Ѻ,�;�[��R��������qL�W]�rF�ł�	R��)����c/��Nlv�s�R�b�J�P������.�
����Tl
(�n0�9-�Pu�(X+�wJ��V����3�A��aU���=�ij�d*ud:m�w)��Ӷ���f���6�|�uz#;��y�
�Iy�B�e�+��Sp��N��N��S`p��<�n��'N&'�63�"����:�ne�psZ�y��_6����rt���R�KZ��h��<�F��~�I�����̍�`�ƾ�����
�VI-!���7za[���W�񄡷X�����L2%�K`�ؙ���R��H�҇�A��j�Q�H`'�Y�I@^�7GP(Vc��@�1f��a���+�>��Kϥ��A�Ie
�K�ӝ��/2��4���ӡ�P���=�ޥ��	�B%��E�:���2��C[vc�R�# ��Q��!eWhWc���VKd�9Rs��E☧}�l��q�9�^�!� 3��,<A����=�?z)TM`4��q�˅ZJ��U~�PA `ny1 q�2�j�	�00��t���~_�A��;Dn��J�0b92SӨ�ss��G�ơH2,Z3����ļ��_��9tK�����\9�j���L��5��&,�@K�2-MO�BE6k�
ū��3����f����������nH�A����$�
��:�����u[W6%��}��.�L���@�}�Q���qQ��kD�s�����OJ>3�r�Kb�T*���������~t4£42
�:��1��K"�ٖ�ͣ{0�G9Uc�/Ѣl�0A)��z��Sڳ��h~�������~l&E��maeN�S�m'ԄR{!����w���(�<�Y�l�Q��CP&���Ӓ��)v�m˔q)�1pa�(\.}���Krt?B�ս�E����]��r�M[Gx�5ϩ�qh����R�yh@�������ٛ������m��4\�ĺ�T�����a�R�����g��hA�R���!���ѺXԊ:�O���G�_L�{�HT�=Ԛ��<�3	J���gGwI=V�HVR6�ĸ �HS#��hBt�WҞPpq��`��-�Vm���+6�}u��$���A(�h�͙�����g�S�R��ZT^���ѦO�)��R��C���O������*�±;��01>��%aZ���f�[�Iuʿ�'(1��U�6n�S�imE��%BO�X���)�G�tW�<%�1�N���"R{<��6g?L�w�d��(q@r�@�0�q 1gZrHW�Ͷ����`[G�&#!�!DT�D��n)V1\���{�,)�("n�� X�kcf-��˽%��,�G)�E���|8��hcjYh�.�h:{1�؂�ق��-�B�_d�o�a<2I:CY�������W���nITᗝ"ď���s��&#�2��۫rV�S �S����K�����K��CL���tN�xES��ZP-�L|x���8�Y!,(�itˡ@�7pt��[?nA�`��*t�O(CU��(7�g㤌0�� �6�D�zk=ҟ	��Ɛ�NpV�����as ������4�U�v$v-I����}�L=v���m}$��5��߬���C��
$�b�r�rޙ	�ぼС)<��٣�LKVL��g|��K{��dN�e ����C	���^n�Dm$�7�ky�׹A�!������������	�0ZG��^�����I�X�kݼi'�8Ś.������>��!m:w��[Qq7�iΦMh�R�G����B�W`nd����Lm
�Z+��Gp��Zq0_D�0#��`���﷌&F$�Ԋ��-�Rsu	�W�:x��^�="L�h* �ٞi����.\�����T.��7��c���`�7C�9lLRJdN���S�DB�HE�NՖ��K4�IJRj�$�g�m�m{�u�����2�LQ�5�T{�+_'��M&��S.26�z�d��c�
�^��DS�քK��7O
��f�nի3xv��1��{Q�ɺX�!�)&W��k�����'�U�р��Կ��MY8vB�2u������wJ�(:5�XH�$��kͻ��/l`��.��B?}K�/�aZ��רq��yߧVߴ�k2
�be[`�������iE`�,�ڷ.��B�1���'Y�.�e��j���Lvh`�?�����Z"���}��Mt��L��'�T�%���?;p�_3,����������*P1��V���}�#2�M��>kףE�~EO)k��y�u���9���/E�L�o�tG��H��D?����@U��h���=Qkt���� ԕD�G
=8��
��/���U�.�'�Oy��>ԕ�r�	�{�Ĭ��+(�s��˼T	|�h�N��hv/J���x���������p&C��Wk1i1Y���Ո��]���5"�D�B^N1Fh���\z��PF5
O7���	?;�L�	���s��my�j"K���q/E3���6�&��ç͞2	O����	�fB��+�K=s����ST\$�V�n۵��t�ߵ͠-�s�bܑ�