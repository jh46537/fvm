��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�=���,1�jӛXT�d݂��]S*WL�Lnt��V��)�ѽ�nː����2��m�D���#�o�֊#���!~�z�|��^3����qť��q�AM�:�5=l�+��(&`f����4�`TIC�����JO�8G%Q,9Ɏ�8���6=/^� Pfz�2!Z�����P���:#�
x�W�F��m�ƚXyH>e�����t�q��o����Du��a:�}���(�oc���(?͑�mi^�Ssxm�����l��w�����n�m���P�Q�.fԂ��dql�b>y�KF���
,	%�����ʗ�_�Ս� `��Vod�ȝa#K������S�^bs�0�Y9��w��+�ՔMt��@?���ԑ�|I��&�z9s��-�V&���ñ��/��ߜ�cQ�ژ�W�|Tybg��q��-u���w�~z�U�5�a톶`��.�� ���J���a��p v"\y�P��@A��Sy�_����:D>�~�! ĸ��q#�猡fW�q;א�/,�i��m����Lݩ"	Q���m�yB31\�m�(C�U�ѕ~'D��^�� ���6�_��Q|�;� ����������8f� 0�̀3���>�'E�I��#�q�zؓWd<�B�ȸ�G�>�x<��K*,O=��[�	,X����p����h�KT;�� S���#R|"5+�՗���g����4�.�]�3�C��ɴ/���&�|��(��քw�CL-��Nj�N����3�̐F��� d��D�(���Z��6�Y~JJ�|�X�9�Q�b�A�뽂�>LU���ڧ�擨����߽
�`+�F
/������ڹ�aԙ�Ғ�9���F4��/�gY��W9d�W��W�� ��B���+J��<�C�g!e}43B��P$�䴍d��rXUª�|����ENT@�g��rC	>:�!)�\W���� Հ����9:"�������S�H�!z��)Q������A������\�(�G�v�m� �Z��5V�#l�c�vb�cRUֱ�&]-�A�ZD�cG^~�mj��'"����G�e���CD�1MN�j���3�?���cH�h�H$�N���%q��<��50��~D�=.���CI�6
����/Ժ*f/�ǥN�-��Q'�a����D�-{�h�C�V���[� ϧ��B�W �5�ěNn���pn���w����^�n-�I/�ހ���blFa]㗠o�*j���i3*�I�tj;b���׭��LƐ���!�}��֢Bg�|W"�㓨)� �GG�^��H��da\�
�0��0��N�eUl����aρ�D^�Z�yM���qF���k�f�Fs	Z8E7�UIE1p$i1�	 �� ��=����D�ϸ��t�)!2O��t���<V�;$��Д��F����
@ ��r|���&���qu�Ȱ���㘵\���*��1�)`E:�s*����o�%��7a�d��QqЪ�!�v��dKC��z�Mqze���"J���,�&(���^=6E�5���N�����D�lo^��[���|���ϟ-�Ni��	�/;{.a����t�K6W���3��*�M���w`��Hĭ��S?%F�O#����A���W�
$eG����q�MEa���Όؽ�l��eɠK[�v�ھ����_����A��Y�w�b|b;���R/bct�&�6�h�b�)$�y:�ܪ+_H@�Y<CR� ���Q�����Q~J8�9}�l�Sә�7ZQ�?�T�8�p�@�P���4d�GmB �#�cH�������"�%�q<r�d�9�}q�Oo�C�
��<�:`���a2iHaN^`�dc���#�U����U��1O��p���C��
�\{6�/��Z�b��m����ҍMdU��3�H$�r�*�GçX'�^��D�N ӝq�"��iQ�Ӣ̒��gx7�6Y�^4�¥�|�S�h���U�)G]��!��K��uQ��|�.�oW��	��+�{r���jQ���ɈA���z��MK@�mKr�]ۄ�E5ޫ։r�-@!n5�{>?4q�1	̭�	!4B!� h�ׁfy)7g�7z�C�X��~/c�;T�r���S��<��l<�[���!^<��G���%�c4/�)�2|?���^Q�b7�lg$�Ѡ�A�A�W./�_�ۊŰ�p�g�I&�uP�f%y���Ig�`�1��ۂ�.��.{�$Fe/*b���r~D�Y�$N��nc�67��*MyH]֧�Jҟ�4���aL�)b�g㶿�5�R��VȦ����WZx4��6&h:X��7��u�	�y��!/]����`'����=N��,&��st`a��ɖ�L�{)��o�!˱l�h�yW�9���@�l˃b��8i�&��`C���WT&��@�#Y��X�A9\��`1��F5��a��o�U	P���b�d��O-I���[FBp���[�ʢ�/D�:�ׂiBJ<:���P�\9%��8��zY]�U����#d��Ħ�7'����6�-8d��ҿ�f���a!���[��0=�[@eͱ����W���h��B�����V�et�d�ܑmV� ���|#�a��S�X�Ku\�J�k�< �'r��_z��?����"n��1��t9'K�n�!D��8D��b����ڛ�Kω�A̭��ڿ#�k��	s����tڛmh߰jVGw6 T����Ky�Xd�ۋn���S��V�PU�4���yPܹO���d�� �B7	�^��v\�i������pG�1��xkO����0�o��6���CV�o���`���Gg�)gj�y���{���T�g%s ZC��u���:�����ɘD����I�p�D�C�µ$�_,T}�jC7)ՒUmfښ�;�I����GvM�E�Ơ���]�3���J�a���9s"���z�Ďv՞Jν��E�[�FE�]�Ta��`@���Ȍ5�.��X�E�rC]��W��P��[��+,��KY	�-�l ��h��R��e�ǌ�a\;�(��7��ɦT�w����̂�Lc�;�YSc,1͂�����q�#$1P!����l���V:�.������`�}B8=��cgܣК�����g�F�R (qv"�<%�<Ðk~ �oJ�>;�ё�l�P�;�x������j�R𘯡�=���؜�3
>�Z?��n
o^-�vEj]B�[Q��K��Fل@���6"a����nU�[SH��2ꖐ�ĝFw]j�Vu�T�K�ݖ�����h�1q��P둾.��%�L�֢�C���]\�6��j�~2?J�M��P�/tqDf6I2BW�e�	8�Cp4����f{=^��J�W��>;��|�q<s���C5��'6ҕ���1I�5�j�Uh�	"��G}��Bh\iB* ��&����ϔ_V�;5^�)Q�:/�u-3�Q1���y!id����t4wi�@�ܝ��5�ń��w8	+�´xdm����;�>�^�y��@����V�. ]h���.�0cd��y��
���]�X/�y�*l�ǟ���+_ +�Q�´���t�U�~Ϊ�'�x3#�X�\i+�0����C�'�ܰ�	)؀����"'�/Ę�qdhpw@��;t�)wb����6f�#���i��M00}1Th|i�~����d�B������f]��:@>V��=�8�s�>tnBL��-��b�?	�e� /�s�TA��`ƿ{u��#�|q���c$�:�/6lD�X�p�
���j���"ֵ%��sʣ����f5�SÝo{%��yd�9s�����I�FF���v)D�s=�3
� "�를�H5mB<m.�Z�nh8��4P%��/i#�I�`��V���e�Q���.#�$���&cd���I���sƺ�4�P�\�d�:�0)"�󅳰��k�^�ݬ����F.�<�M��L��H�߅�����r�&��j�NH���^�����y{�C�$Bc���z��!J2�jZ8������3ho�Sɬ�Dej��y��,XT��E��h����Kb �7�x�g�C6��ի���S-X7)�)�%q�_���>*�Jϣ(���ڦpX��(q�F�sU�jt��%�k�Aŧ]���D�/���g0
�J�������f��^!c��������VZh�ht��e8�`f�n�����iY�)(��a]��ཟ�w��M�(��V�<�ef}�ET�74OpY�$Á���_�^�Z�.������q|Ex�l�e	)|QX�Ra�Ӷ�f�*|����}�3�r�a��ZnS~9jմ�妺���V@'�3(~Br3P�j�q�ؔ'����^u��@��/�9�E�T��{: �n83��2��
y���,��m~vK�������>M�����͚��Mhmvm��b"�HcA�b��M ���I~��6�&=sL����F��\H�s�¨?�k����*ڟ��4���i# Um�C���}k"z50F���b�4C�M�k���y�ZJT�FӇ3�-h�Je����v�?��	*������<.��d����x��a�7�&�9u�h����r��y�쫓ݐ�%����Ыc�Ϝ��\�q�`_ғg���RC�@_JT�x ��"�K�a�s��OA������-��ƕ��a�����9l�]=��#�v�ɀ약�M��&`yTG�� chU�=*��@T_{Z�/ֺh"^�S4��ϕ
jC��N�E	����+�f������ �J2��*�[J��32W�T�3`��£�)H}�����]=��=���Y�Ыq�f�+�ǧ�B5�����!�|(Z<�W�[��_�#�/��?{X
��s�N7�2vI��i)���E���)��x�̓��������F��mJ�%�J�Ck5�]^��i�rc*8)Q���T����(S��P�3cY��k�K�_pYB��-�cU���?�;�t���RΩv��"ۧ�{�{g\�^�����Y��]$'}�H'%�02���P>z�"�Ca�k�U��s�&�EX;Eᬐ��M�Ϻ�m:�`��n���d�'�����^�kW�����W�KZش�a������#��Xt�%��Q�Q7f���q�W�k��ݘ.X�g��*�n�O���+&!Z�啍7�kitx�e�ѧ�c�*��˄���)'�!}FO1�{H��\j+g���r.�ر��9�LX�d���Ƞ����a1�S9���nSn%a ���O����@~������=���B�M�"{Y����J�%�B[M��D
�u�D"v�� !�gw�9P��n���)Ƈ`�W���s�rg�+�T�+������������=E]W[����K�^���FK�5lc}��g��F%kv�^��O����/:�eB@9����R5�YU�N����2BGuEq���	T����\��,;��!�/d_L�v�vB�����ALt(>$?�n���m��FX3�V�Nd�0]�����9����V�b�wm��Kw=Г!�������o�;G���y�N2m��k�{沧!�!��+�Hh0b_��B�A��!R��0��2Ɍ�C�����T�C��Z��g�÷MT�*��$���ی�~�.����r|� ��Ҋ��+H{��	3��T�Ht	b��s+2��Ӷ����x���8