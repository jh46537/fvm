��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9������t�qp/�{?I�0W�
�1S��^U��1=��Ѯ�.�ҵ"�\m�R���P���,��Ԉt�*��(H�K5�|�6���DA.�O8:�Pb��	 Z�B�Б&m�Q���ž Tp<�hB�7��pT�!NG�~`�/S�Y�_�B�o�ߒ
E��8w�&�����O����Pn�ZܦNeoR,��tZ{�	��*�&��m�P���z�B+����I���`zD~8N��	���d>c���%�]Z�ﵪ�7�O�J����Rv�2�T+���	�.�GCet�䂈ip�Z��%���㈳����g�H���m#+��2fL�Ի��fǴ��9Q�����
����>9�l,��'�'V�΢��~=�˾�,h�	d�Bհp�ӻ1D�Y7WJ�������:����w���	&=�fႯ�gO����=���5�^���䓭�yǋ92͋���i�����{�Z�p�ke	�]�DT��Y��=AJ3����:�xE��?���]�����N�&4߆R�k,Q)9*	�Z��72|�}��	$5eg�a(��C��\^Q�/~��A�c�ѥ���5|F"��M�떪�v ��d�N���-^�{%񧇲�]��֘�8%��t�nS����6S���-����2
���p�g7&n	�h���[�P�Ӆ�:+?��ݲ�I`��6H���d*ؽ[�
��@ȟ �K��e|�� �_��AT����1����DHج�B�l��ܤ8䣽�jl<1�Xܼo�����iw���_�3ڪ餲�3�P�?�~Y]�1���L��?�`��|��"U3���z�Y�S�13m�i�h"���Q���s��x�x�]-=�K��:�U2����Nb<e-�e�<ė\�>Є����Q8�\鰆�{/&M쁭��s����'Ϋw��ی�=�O�E��9�Zz�����R�"ݛ=D;�P뺠ǵ�Nc)�Qf���	�4aqt��q�ʟ�y��)�5�(C�QS>��3緢4�$�~���@����$��|}��G�(،&>I��K!�i�</�j�&
�l2Ӟ��I�?("0���F''�VŮIC/&su��k���y��A��3^��4�?f4�33�2*,�T�&�=.����S벜�d�8�rL�!�jQ�c(��E&��L`��j/%�#>������ ך�_H�@З����,���D���\�X�R��2�5\�'bڳ�F�d�#�5��E�J ���-nx]H��OǨ�g����C!y�U��w�ݬߴ���J�����3��n~��0ȼ�
�2�`�N���~.�9��"��,S����]�<-��5j)�⾒�J�����y��W�Pf����N��Qٮ� ���S �w��zR{�ݗ�݂�as\�Vr�����D�4�+��?j����w(�'/��z:^�Ċ�>��1&�1�:zb�I8:�50�����d��ݹ��M)�(V���TK�d�\?h%�����X�3n"Nš����О�	~`�^��Ս��D��?J�6`V��1~z�ˇ1��/hY�IU��K`�g����[�V�ƙ ����耤�9��x��9JȞU�S$��9������n =���1�9��
��a��D��>���J�\��� �P�\��ʏw/+�M���l��������4O��U8P�����^�\pVqd�=�>"��j&d�S���M� 9�pa����~ڝ�Dw0d�-��k�3	�U����� �{�����I~����;�Oo,�Xkg�w�Ǡ�J�|s�q�Q���1mZ�
­�id�
�8�h��oc���Zj$�̕-T��Y�,�&)�G����&��*�>K�}=|�_-�yX�Q��c�K��b�;�D'�������}���t�b�5�P��u���r����깞%���9r�{F�8ᲜH33�6����=܏�B�W#�Fđ�4�~���F����j�b��"#��?�;�O���H���ojÔ��"P������=�����|�A�4�,�3찲��o��1�7��83�����
$ǽ�G�n�~D��M�sx�a��~gq�v�W���U�������)�(Js7�s�B�l"�U��)kG�F�=!�`݋y���