��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�@V����B?:S���/���F�U��1w	%*:�X{a�6��rE�ʅ�.����� �jcP�麬�Q��s�L����z=	��z�]:�U�P��4`'����	v}2�R��4��i+�\�@���=�=E�](:��&ӑ���*���"�ɣ4��m�W�4��;b����Ĵ�^�Sy�������z�����@8������V���jٛ1��`i�b����"���},ԘsrgZƍB��9J�-lB�	�P&�������W�R��7R�d.M��'k�[h%�,�)���l)��Vy�T���?������ܱ���L�@g"�$兗=P��&�̒"�m%{�{�ټ�@5U]��M�����sU�*��� a4�@��g*������Zs�0^H�U%�U�S�ҵ4����^��=��!�]����-���2_��9Fc����yD�.f i�>�@������1�����vI�xv��Bj�� �����L�g���L�&æ��p�=.ܩm{��mg8��ԗ���X�"�=AW�O��l�?��N19�MM���i��>(W)An@����I�[��8�����M�W.��[]���	�:�d���1�[�{jxv{Q�3�k2�7�k�!�/�ٸ˥�db��$�;�)��Q%l	7������<�(����^��iΪ�u�tc� ������6l�A�s~���#�����X�NA�a�̃�Z|���l3+����v�z�}��u�����
���� �jj�����}�u[Ѣ'@tP�)A�#�lP���y�c��6�'fբ9�qD�0|w�@�Rq��=)V�+�>��I|7�3�z+�p6��%з��F��SJS�J�S����4�
�E��P1�Fg��5t�guaX�&kG���b��*�\{����YqZ�3-#01�Ms� �S��U�%%�8�ɳ'����
�����"�5�mr�$�����}���ɣ��cL�P��=�6��J-'귔fj�/�JHg����2���\0]4�a��-����Ù,�>�7@����}��-gZ�~�:MTy'9N��7'��!���,��L���Ӣ��w5�u�� �Kq����rt� �ʾ6�ͨ�?ߣ�5?��+?��5�����y]���zְq��Da��u����~�'kۊ3T�*%T�/�+2��v��s>�2��y�� v�!����mWT���z@�(�G� �{L|��A�Y�\�ci�Պ��]�MYr��\bj }nJ9ƪ&���#������I�s%i��D�2�e��:�1a�:��B�Żp�&tZ�w:^�@_�j�
������ ��ٶ~�:���rȏ�u�[xm�e/� e�ǈ9[��T���-f�~E�bM��liG� ��_8����63Һ~C�]c�P鱘
)�2�G	��6��\L�ݨ3���on1����CG� �s���z��J̪�QL�JP��ׇw���)�W�sY�\'脄l�3��]���i!��EL��t%�������`��j	�w�����p:[rrC���M'�u����4&���[�?���
wGԒ��*�T/�=��H����7��m����q!�"m�H~��Q	(�5����>�uv��l��"w/����ߩ�I�b�$<=l>1���E�2s���Ա���4���Z�	o}�ZM���ͥz�`b�z�xJ��ut�u�}�-��]S����}��/alSٵ/Μv�ޟ� ��0��x��!p�}���Hz?Qv�h<)�y���ذXT$��v��3����b��xP���^�5���-�����-�~��n�_�{������a�֭�U��?��Ў�c�||1f/��@�
��W:�C���F��Om{��@�N^I��q`�߶�kr@/\�����x3B�\ҩ7ȹ@�J�S���~�e��I�3B�p-�d�;]�׉C����M5�`:ԝt>!�]q�����s��tEJ�5Ce�{�� � ��8$;�~{m�ݝ<h�s��)����Ȫ��s��E������zi���ۡ�0��Rlz�@%P��0��
�4n��Fwy��*'�Z$��d@�9���L�9]�<�#��#�@ itN`-��**d�Dq~�U�I�#ud���s�`f�I���|���Л����#^��uYի�"ېS�+�ި�9�����ʅʝ�M�MƓ�-�y�_�?�I��{x�7�KP��}D:~��u���ݟj�x�Z#N̛���y+�d��Wd̔}��艚m�]L���Z�fg>5��t��!�!���N�Vu>"u�t��f��Z(g4�s�E�XN����MŢ�Ed��� �-b� ��x
MI��n�ލF܁�����";��IK�ן�§��t��8�P*qt�����|�Ĉ���c�q�YE`���(�u��`�v�yD��Ս	.c��s%ve��w-�@b�Ұ��4���KC�O!��܁��:�E���S� �^�ݪ%]1eZME�Rӂ���Z�nπ|�+șDЊJCI����xj��[�R��v�Fq<~��ҿ��V���f혹uj ƭ�>e[��|�)2Q{5��M����Ҁ�>z �s������͡Z.)C_���P��H�{9�j�\��o-��{�l�h��CՕ08)G�ً��ǧ�W�2�sN!���9	' ��F'	��"����*�!iRy���w�*o �H4�y"�� @��5JL&��;�#@Ut�|��\}�Z�����z��v$H��ɗ����m<�~,���Gx�j�$��CIR�g�")��
�s��]�	I��g+��kE]67{%�xbfE��EJ��[�id��Qz3����-�>hp�.������d.�����A�ټ6t{��`G2�`�"F��� �Qx�y�T�҆��������������D.W��:�'�5�9�~��[:�h�ƽ�%�H��|Uӑ�&m�:����L������ֺ��G5�]'��,A��0D�Th얔���n���䏯�j��X�e����?��-����{'�S�!�6y�*����5LC�o<���h��ɓ`s���K�����ǕW�8�gc�5���Z@!Z�b��[��w>+��kƛ��Ľ�P�p�(�y����n&V(,�O���������/|"���S�xީ�e�Dh����, Tu���h;�� �l"�SmL#{M9D�������m-q�*xa%6��������IuX���%�o^��h����,]���sU�f�f���Wr�'f�Vr��<n�A��<����6*�t迏��ӫ/�9�����j�����8��Oӛ�v�7��	ECkr)�j'Xe{yP�8X.B�����e��[��/�z��ݒwʂ�Ir��ڵ��H�z�1��購��M�^�B��<k�X���	��i��R`
���#)=�u;��7l���-@�����j�W&֕�F���"cD��u�S�)
�9L+�BN]�WU�Z��%�+�^)xVɸ���F�Y�o~���� ��,?.{d}�R�ɳ��ז���w��DQfL�d/d ��F��o�
@x��S�����k21eM�N��V��z̃���8�:�M��7��+�2y}q��+RҎG0	�����%��:l�dbGC�Nǐ��Y��F�}]��#9�7
��.�(�Z���U��Ϟ�����lP"���/MN悤���/4	�o������W��AͿ$�o� ����Au���&��&��e0#�	�AƔ�A��k��>Z���r�Dݨ�L��z*;۔ [h������)2�Z
{�	|."�x=���Fp�Ie�a���I�i}��t�ZCz?aaB�������򠠝�U��ǜ��'h��]{&��QYQd�s2YSJ&\;SZy����.GB17��2��]5<���0�C9qҼ�����u�-�{r�.����ە($���FCM:z�i���~.o��њ)��&�陂q��O�F��?B5Kwyg��tI�b��$s�bE�����)V�<T"�3�����p_� �r��_I�ÿ�g>�����=W��a�r����_�O����������ڃ�7��H�-���EϬ�M>��Pi�ݙ�S�D�B�<��߭�b0$8��>�c!��-o�z��q��P9\�'7�0�mD �R��1w+: k��cpH�y�p��5Z���t�+��������&X �|ힳc�9���ÈT��+ʃKX8 t��j�f@H�%}���X�k�4�h��Q{8}=��U�1����]a8���7�z���̃�*`s�I=L ����8?��WW������ST�S3?�J1���å(:�REõ�q�����T�ോ��������(�(���f��P�/�<v����ӆJ�V!!F�#�r�M�o������5�-�ޝ� ��ƿ�h�����L8ƨ�!X��6
Y���G p�O"!.:�4�*%Ӿ��
����Y��>��c����v��$��n?����)k5��^͡��f���Zh1�~�<�����r)-j�����6�6]��KvTC���xY��jq(=�H��UF�����<��EǌJ�3ʼ��I?A��o����I`�k�>�z6�t;�=���f �)�i�
��S%��,3 ��I.F<���%{���RU���CidO�Q�������]� ����`Nzȑ���e�M���+���<ÂFq�ޒ��3d{�tp��!�I��Q$8`��lh�y�K���Ƨ(�;�[J,��[ڌ��!LT���Jr��⬳��(r�ͤVRP��=��Q�n8!��K*���o���>��w~���6H�;OG����b��6��W�� �#Ͻ��}� ��8-J��
2 �<��"���$	�����&B_["#-�b�!v�g=˒@@B\�)PN����iUcG�;�m��_	r�ب?��W���G8ZS�`���[>�g�`�5.��z�P�)K;7�K�\I���L�<�	�)������i��,��