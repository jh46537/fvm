// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bZZ2w1FtoWvSkHc/7A9uonpcOY5568EDeWfOlDjnpp31E776FL2ja8AFPevr5KOV
6ufIbJyxFjwcohCOt/k2LY31BF6uba2rqGj7inAu6HqJqxTGWCme0ARMPyQYuyNV
SrH0IzBwMmPb8uaaftZ7Nz4CTkpMvgnwxgZcK/KL958=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 183696)
qD4MklhlFOGtun2astJ9oEnsgk9mG0MxTbGoi+Kwwh9VxHGUw4V1r3nNKqyhRqdX
sI3R/X4iV66JnfUMDJ2Y4RTWXXkBlPq1bxqDsOTTFnGFXfZvTJdFM52q2oQ8HYxD
nqlZaJ8oO84swvdKbRDCWuaLMsYDHur1GMJsjoYjz5a6pSTXJ3Q7A+qNLQ9HtcJJ
72J6D34C6yaAD26JvHzlXcUNREXRpg4TPXwRlAim/3psdoNMdTXpfWz6wLv3jnCu
ap6Ae6MqCms9ZNIHW9ZacW4f5gUXHW8k9R7ddDrlxzsZiFr8NdS3mDQHu/AI/8Ac
64BE3RgH5+ayq6TCoD9HMAWoaAKBShwH9EqjPUO107ssKS6kjfiPtyalE8w95WL1
R8lKZnTkl6KOZClQ6Qo1A6YMXjeAKI1Evu42uLCZVS/fOWiQ4stjQWqInQF9e/cM
qZcYp8RtoebXuR2h8ZCXoiJKewFdmJwgvwBYkSnW2BWA2uEnrDSUgLXPau1JhlZp
pD0hbUv2x46hXTb+n2N72JqfGR2AvU/HJk1O0aXWjPH2e0nEdTacTIsRRykQocfP
WIgNgbb/SrjDrzBzDKosfXZVATu8F8IhSf9YVMTLcLP5GMCLK0F862qc7Bugzilp
IyWQECFZ45ENlK2sopiVOfuKO1k1ifbZw9Xu2ZXqRnZPphK0Cnk6xFLAvYz+O8h+
ga4eYQTlf3QH+LNW5r2HZGmM7GnS8ZFJ2QKOz5C/R4L9oqCMF/2oaYiz9607NWd0
iSgbGhGYuYi1bwCWOE9ZeUd0gq880gkzS4oA252rRepndXW+bX5iqJHjXkfdczfx
RgQbh1VJL+AKkGFkQ2zh86iQ59/ATO3ze2ZBcldabHplCPfvUYEfxiivytIhNli6
5nz5c5Av7VPoUtqzjguxwLtKbHKFyHyX9PJLmmUIX9TAC8Ki4BeojAOn6/T5DlFi
UJJEOLSUF4NbOSAe04YMIrGVzalsyT12h2nCiWgeI8ArDtkEdvPTKf9jxCIoGhfE
0bsB1yZiF+iaC3PfLGxW4kGDWG/KB1kgWy90z7VIZ8RSmfaMlTTOAeMNZm0C84bF
AqT87JiZchDsYIcQZcv4mOcKiw6uofMaH2/6/tlIPoPY4kUvlRFeiz7IuQRLGSjc
O3JFqrUaxeeYP//+Zuf9/SSenqRBDxBMZ5Rg5Q3b1V4Do5XYtkfMUtfIiADvGjdc
j+HnWsTfxm96/K6dnGXIcIT08bYl17TpQXpp6Ptymkthqy+hSHRFwwmHxY08CPJP
enwMln6e3DYPCZhAnTW7pyi+OEhydfUkm+wKRvEdw3nsWOzIDh23CDz5zn7iPpwS
MRq0Q/E1YIGOY7NJkkNrXn0d81SG//lwYj7nL/f6vXZngo0xrrfFKV0CMZWm4SEB
hXfSG+jB0hmpTgfXcckaWW3zh5jfCAskf21m1bmFd1nDooMBv1O/RC2TQvliYOYQ
b6XHnF+yF/x7M0BdvapiOYgib2c5ImIci0lPBmGHsBAcjo+ES1Y9awiKNA18g3e7
hWWmBw36LteRzm9i+DJ6NXYyKQh5NhwYtXAnkaYPdrlT9CNNI7ZAut7uk3HzSM8/
MtEb2hpg4RMBTN5qQ0rqVhA5RVvfRk7qUSgJ0ess0PuFecLVgIEip1Xj18+a4zcU
TwyGCBYbo4Q0syzE6LEQWcQ9YDjcFC3OjxtF3SSTfCAhyN4EvoSSigLIv4UvPQJr
j+oOLFyn3oeBXPelsK/MreE3RYHnT1KbYa51LXrXJbStQiDAUziMot6Kmb7RxbL5
IsbSP7PIdxXxAf5p1tcpgEOXkRKjF+2v/KflUku5orVds1SALY99teI9UYF9QEmz
bQ0yPsyojOHjGYrUAfzbrRIkq9A86GDJ7/5FEzOxXjTCdEoxw5b88dP4v6iDkPWr
unEGksr4SlnTkLlJhcB6WWiYmg+JYnmjDrERRvzg/OTHPgU1avTtfK20yi39kdvT
DdsvADBj9RoYOGqlHgMcK3v7TXV3R0OTTqdzVC5bDqehtAY+mIaMyB2irz4af31X
+a6tFUTeDeIw4V3NMtokb8XtZJiEmxDRIo26eYkiDJi5633XlDW49iIb8ttJYfcU
wlwYefk3dnbC8REr0Q0XlYmuSeHmGyv8FpBYKo/CQuRXgADGFLMZKxcajpCXe29T
rrK9kt8dFhgMBElGOW9qNWXqz+/IPRTAyruU2aeLt//vVFITDqu4oLIil11H/Qrt
Ysnf41Pr4zHvNWm35gAzymGvjOdLByVQzOaTXemEgYc+qIwjrcmF9V2OLNFgTjD/
gitd6q1a02QQ3u/uQhcSifVjD0+CPOJapEc7s+fFVj6rG4Ia+0BiSOwdyTAorx2J
nMrtj2pO3v2u2jpWaT0hhlFoduN6Sbb53nqx/xYzXRJt+G1iTCr8rXPIIT09m7HH
FGDv1cbmN7N17uTs205etCPHA7rL+11i3cBeCaRKyPqfe8KPUbnEC9vMGka20kcA
kFsY17CuZNy3ILBE/UsjtlkgQ1KQEJn2a4Croi2tlptaAqHz3Ldb7T8ObnKP2dkD
pNjKkTLNGxeRqcRWy5+yxlVhHNJN1o4gBr1nBt/Wg3Uh1jyRi0HLeK6lcfaajJV5
O1aEoIePvYMCr7aVKD8UTSSQijWMQDJmHfTF4chgujaa8MBKi/dl20gX5y7NlmVQ
3uADC+Uk4eflg+qcNLyPirdFZ4qqlucTLTNsmfGHNon8pRYB2KDKjq+V67ktkGzo
7eUX0wQCm6ndR5j6daykSbT9ecNpPIpy99a8n3rpW5vy4L2IjXBieiSoq52KG9h0
TtE17f50bhkojLi+fLJrc425QJLUbj2oh63CUrxr65yXimrHnl+PdzKpFsZUUGVo
2y2bLyALGezpFlnt7X//4JHUAhXnF7/e6ILKgNX1tLkKAAOYZpIxtQrrIqH8F+mO
PDs7rBwrkx4UK3nbfHsrn/LYJv/UJzJ4QPThv6u+9n1gjzZVqsuA+atRyPu3A/Po
tquf/t3ul3YEl/KNffTWRvNRxjalNJyh+qhU5lfgRSYmD/fKGAV4bOSsPhurszhH
GeXtscM1ncq8QwVmBKURpxX1o3AgntKq+ekA0SA9O8Nwrz+9f57HZtrZ4ZijjgDf
D1mF1s5+ZKfedZbX+2d8T48Y50S5eis4SROvtP083+Dp8VEV/vAXMma4NVLL6wxt
YVX48DOConktbruWKIymh7YUarnGnkX+Y26NQLBv7O3z3OBTpRNPl+Ji1JbnTYJX
C9/ZyE8Yqjy8AvZckBZrtqqt273oJfnY0B4v7SK1d6pIm0jvw/h8A0SqIeb1lU8B
SH5Atd4vjYs1WF2tmeg7eNYINbAyYuieEQAvvSOKSIcfueKdF/sKUa1Pwwa0ytYg
8m6Bgu/KNIljeJW7mZdSN5qgmB5f4aXmKFSJR5IGWFil/YeY2ciBW1kj5qyh0dtE
PCAQGCuT5oy1Zf8/dtG0CbQtxwtEkjbePcNh1NLiP/zxvfxkXNaLClVskFV1/isp
XCCoJtOf4tkUhtis4Sq5BDkQ2ftMT6fV6HegiER+/DZwQ2bqdmIXL7HCiZ5OtdTC
j6X6XXdrVjdMgSdAaFCEgvPFz8bE/MKBmrjydcxQKldo64OzFXeh6ey5+3t3q2aw
WdPrJx9emxaeUmMAAxHMrJniyZI3qXjzSNmetxyPDQKEDcRTGzEYN13sW7dxRqhM
ZaA2ZczvFgzZXZILRzmIbUqJRElc914Yu43vp9SrKXPABQV1KC87a63ZoU9FQhcx
fVldGLqsSAhXyBYj2XuWQkCO7NbZ5+RRBXZALLWOA30eML9jGLb/c5zMqx/j5eVD
fauDIUiUBtOWCnQhlq5DbPk6cD1kb7GB4AAm5a+SZCTv6CEv5HZsJXyDYLluHkYV
H1XNRXSFA2tnQw4JwfXWGkvYZ7lBhVbL2KN80wItQMFKAuYGOPJ5oHX0Y6drFNUk
2TaFdWwuQ2H0pxNWAdgGmv3iEK64je31x5bfHVoMIaTJxX2tUN2RvHbuUqghLl7K
26siJ3vNSPV6Jq2EIRYbXnyB1Rd2hGQswxRTik3p8xWSeXkwN7mcs7yx8LlrepcW
OLl2ML9xg/RU6Dv6PxBpuWIKZrGsKuTu9ix4yotIqD0RdFOLU8BajXirbeOaf0eS
N0fiIAPsASUu3uTji9aLOVSZkFzrO+IYx6E8x87VF3gzLoV31m1zhYnrzGef7a7E
fHfDK6QF5x8daf0DonNrXbKNx9iOwUCLb5RYdWVJVAOByKgmTQRwsC8sOaql0eo8
9wH4v8Yix9S4UjuVOOP1V7WYU/B/lSHsXzw9Sy3syCt+uQtFdiJT48n2HdI/cO0F
0H3Q4sz7uHvCSPXP90O4AX7gBhzMGdkVkHWeEJrM645G9o7rZfRNpmOJUeBdxpcz
jqmE42gHALEgARHeJVAdbB2QnkzLjMctCMkGMw/ehQmda639dq+U2RDiU1e3vLVi
bMrr+Q1LcJC1OZj7fN/UFBxM8xTgfBiFx7otKvlLfWUIUMHGuzqWwMRhmVy2jeGz
kY6t87YMRKJhTEjMVw1ulNY6Cc3DSJqvgRsgQjKGkakb/HV3UQlHcAWw6P0E0J+J
QzOJvWaKZ22zV+wXc66sIiJIlY9kCKAfZgsdGHPCK9PpOMZ+Ku2vuwJgy3OqLbM9
L2CQV/01bIxzTd32luG8QyC3HLtfVK63Z9xxU5S7JR2zeoLmq7QqgevCzani5WTv
sWQy3yBgOLbsaQZZfv/j/D5shffkeOkk7kMHGpoTaw9TdRswAt1Flw2CbB3E23Jx
n6dtAytFjhNLOxyHTCNTec+RDAW7oT6JNwAnGJhzlrYy++mIB9EL46l3SDX6rwIg
WKohTFdCoiLTPQbPExie7PQpRfeZrTCmrv3Z0rIPvClzFWkE2gJpuSuKm+GcGegs
6xjKxFQE0hE/pHz8gO3Z4GWL1+XACD33TRxRIfjRaREMJcIDFaclxnBJogBCoQFU
5mShVKSrG718ad2FSvJ3hxloudb8e5mPZ5qqaKYCEhcYQCDqpHv9wSCsEkgZSmJW
14hYlYuZ/qWJTpUizdGBXk2kcrtoGs0mKYaKw9KabjuByeGHoyOJURZPLgA1liSt
TZBKiXEHSUyy0PUfmQkK8aSw59umXE6RwD6T5jssPs47T2bt9ANvYIokkJ8pnXSq
gQAoIQ0vbr75rvPwSOuytIdrOoc8UtXB6E47c7L2mNhH8bfEk4GO2nmESDZje+9K
gszN5f2FKXwoZYtBqOxc7khxcwwM9DZ8O2Didy/15XuckZC9mAZjfiSV4rWeTykT
eHFHgZ1SoxM8QYye+e/u1hYkBOA8ZTf/lePccjNdxeRqRYMih52vnBeDkaYbEzJ7
JdRkGAoGMGIlyLOGvNUIg55wT7NBE4pZ6CSv0LCRIfuPxO0eFNHMHaP/TSztJvzH
GIu7TbbGA2P6Q/Li7zzScH/cgMexxJtLXUsfRMEkbYO73jVhHofmOGFkFhfq370s
dA5VgMD9tWOsQoTIScqQnj38ZDoIujg7o3WI4pbXk1DeSBROItd/nCPZMRuDUGpk
L5IWSVW1LzkVrpXuI2tqdwQkYK35Ky7BFxtfrgiOpg/byMBhT+SLSY7/hh2iOyuH
r/QpF4/yyHts+eloRzzRAd7CqyBmLj5swukRMsxXB+s66KmuflTQ9BWT2C0+PBs2
m1VcIIeUfqjrXoTF1bWLku5lZLHTOf8MvP3ks1w35MvU/4DTJDgaDvHUypOL6UZK
JV4hCzxpYdVik17XKz4shevOQaYgC8TleUbPRSDFEaRZx/6hH7VZct81/SjUYLct
xI0r8ogtSh+KhkWHAtHQdESZ3XBjBM6d/UFFC53b/DL1LqzlrUUTpwMwS+4h45gW
NJ68Ghql4DnZb0yupDh9cBR5wALWkXpm+Scjv5bk/Wj3mkOuGEAMAPcK3DrWHHCz
9oF4qslho362CxY6zFVP0+fA034nvWCqvQmQhe8/yYbeDagRZ+fC+NkgTyqN1hUG
GMn8X5NYY7W/+c0iz1Cj4+3hwbgdavPc6FMbH/6LN4JZJ/e+USozv6pF9FzrwvVz
cXqxrYeCexoOv82t4MQ7g/QMF+b3IkUApZL0nMtFzlciELbeakZaA1D5T8LMxSHg
ymbfjFtXp4T3u2scT3c7w7953gATqsef2QdGz895JLWx+FMGfJ0oyOBof+SsLMZ6
PHfGzZTKC4vguPJ1mD4els4ioUoGbp7ZvBvdxQRlGacnRI3NV4TLV5XYB9DUzVH5
KzaUbBm/NxIJJERWBgUYhegbu07EdTvz9d5dNEZMHVQZjFuniGUFA13GCyqCXKJe
v1EKke09MV+gdGvg6IhimE6Ttw+aJZij+oc+qPQD65DaUynYvMqQDOcO3pQxVrnT
PNg4qEIDkHZnQnSpRDc8CrHbbKi0Z1FtU9SwwELyQiqzAgWG6knONc1XHV+Fz3H4
BlCtfzpEVDCLv+rI5+zlrWQwpQ3nPMCAPOmhwhZXkXFuoRYNIjCKwPip4DvjsLBN
R+/HRUBtY2mKdSMowdlU3ORtpvf68qjJ/GGu5wqyY5Bss8pVBOtkQiDxjlWTL4f3
fh8B/Fvfb4+9adASBMK/ZVdHe9CRuxRWBRoou5kOK1OLzVjSQ4I0h80K5W9pPQEw
v4eba37YYME3GUnc9D02OlGjOerUrF9TkevDPwdzAyhu4efl9NOuXA3jHYDPU8dT
eQdh0orZR/GGu3cWCLhp87+IXhE9FtJoEaEPx/K5pLTJ4LNtspP/90SNa0oWrt3e
fj3SuV2x8yjvZfMeTOy5tTT5OTIkGNzpaQpG5PH0IZefVDvRNsJhrKrEJ2Ik7f3Y
fwd7+8K4JYU3JyLb3U1TsAauVmm155hYp3fOGVT/YwWSWd7ivUiXVRYNMx6cV3Gq
9Ufvc4KCCzs6WKuDbyuetTwSPYhs5D/8mTwwJDjlaEEWtF7GdHi0egZq/o1n2qzf
U9P38MsMuydhegrvf0MfEYgff1MaM3SbD7XJNtPVmYa+awHKVirfrrEQbpPIhEyV
PyGJ7JZnz4N8Qxky0EwFAgsg4fjp2GF0X8qvXw2tnGLp8WygFep6MD1tJ1NLTiYc
IuiJaMGNIcLqDYcPpvFOcU7IGM0kuIMOULTaXg9O8OnmCRYRFbPKLhJSlNiKkhnc
x1JoeTHwFe8L62XwpBQmZCWE0miebQmLqZud1OiJ0rNEU8/9v4NUtUxrN0iRc/n8
ku3O86Rc8JgQIuqkp3XCPphdkycbStnbekvvrxOLd9/1dFugmPzfIo5baGxyUSWB
uich1p+bT4C5uwgYpS0SQE1ynSRV1++zqdBRVPkeBTmYVayyz076QlI+e56um7vK
tynRFdHIZ3rySIzqthNDRNFO6UNFFu+XGFHxvGQGnLqwP8CP8YfhJCT8DsNNoNVi
0P3YlzJ9CF4KFD9YxAi4LIZnqYZK9sxdOsmHewg4e9AbgqMtH7ayvyJwddeouMew
+H4xylPDt/h8VKduZhPN+cIiyJVzdSdV+hiHr8V5j6QWtV/PPDcGiLL3r8wuxRvm
hy2IOcCvGL7ErKzTMITcDXHs8BRugwP/K5SEtZNcuYII7uXvbF2E1O6qltNMEU4S
5TQxEsEOWtnawVCiaTPyuBEH8ErrTnTKUCZ1eOZjnDviCCLtGZXl9iiwnmWlvd2b
V/CMrejrpLCWP+vLz/+NFzsHS8SconQ0PTBkjRtTZo4FanIh07FGwqoQHuVJ7VIz
tLrYRcy2UeARQn0hvTUzTKEjNOZcLng9Q4kDawc+EFpWHeeaoo3LxQ9fG+QM5yPK
+etTWZx+Db8a/piUQxtcM+dfSJlRAbd4wlHzWAC/TVe3vH+uhkH/vQj1pGS1+bNT
ynmsgswPEqxX/pWyoUSdVH+m08QHU1Al/wNUAUUrR7J4yBZXqN/MQ+uAjLfM3YKg
RMRO4UJbyQm8vgTPmlEj4gkO8Vjr5Cm9rJvOyXH13IsbVH9MtyeXUaqet/zPY5DN
ZgAe04Bp0+PKvl8HznG7sam655wEgFRFK27ZF5RMRp1vtdwbnGJLBPRVwMQnuzF7
FrB47jv2FXBq429Kc5gJXbObzd9FbMAQVAQmQy7stWqLGNAtBqnkNENfhBSxfy5q
ZoA2OzQfTa62P/pnnyz9amuTB30bJBCHwE73WrhfEq+m5zsK+6fpk7MTF+FZpsuW
cZ9jKkJrz0s2M4bt823vN6Au4G6CNHcbcf6OO5mwSKzFBSpnUFg7RXfFNjbalY+e
NUrbMrugFp7e9u8z+ZlYfmk3yv2/dk1UKN5zAs80otWaDXVve1e96w7Q3DV5JhJh
CGrItu585W0OubHUNShUTs647vLQtNhAV+tny5vg1fzOYuK3L49tLjtm2aBHrBFA
Eu2saotQ1AQssRgSkHTD5HFfBf0TmB4tUQ1I/2tyWoGpj1C2j5LMoJUds8wE2YCv
XN3xmJ8JYPkeVtqLDDOU2aFRDYitRx2vEmEawkD10UVePKIXwB5V7XJxNESUvzPW
y5YhhKpNIpl32DD7D69nU0kLtbhp3fI9J6qcYSvi1Fa2HL14Fwg2h6RbfdUSQPzG
A/sqe2DcvphD/MuDsk8ccJUBPGGvVBdf9jop4A69Mm8sYxIkoeYiAOMzDayJXHaZ
apajyVd8ptOj8qxtm1h7gxMJ7ERLd6ZaoZ84u6X8nuFEqRlVrqqvthl+7ANrIDBo
FBhNf5GjZE0aOEk7DT3XUjnresmbPGjJGyJLUYYgmMDwBUgJwqUBzIxM/PzHhGAN
n/jyVER5DhD0dps1myO44G5dc8W2AofoQonGKXyDEjCgFgTKpHZPuURglYO3ak7U
AfFq4RSli1448RzitGBndhgeRciY1a7mVPArRx2iDdznjuAl0L1/PXDNcjjDcPOZ
Pyv7vPTSeGZYS1XGPfvbqGPKSgjK3aY51gxXaJzAq9YhAgoh1md1zaZqV+Jjf3bw
mTipARjFpcVOaufqB0v2ypg+6VE3mfZNtSXStg6uaF9ZfMsvKaM6xs9rCk9Diiks
+sgmUjbY0daAuu/rs2bGZss5HmQsQNDQJ3UZRDRJCOYp5nSwafeMpQgv3LFhRALd
SiyyId/lnltC8nPaoqXD39feCoDF+4BcFsISstC0214kGxl1sg4b/XQ8KaUW9zAg
SXXSr09KrKz7agzzROowMLbxunwRJMrtptIZZ1cOZQqZW6WmufMihkvSIlWQvMhR
M0ygiuQNmcfQs+AgJFcKXHj3Rpr5nQhpzxP3e41STfkBD3DqAu9xGKp2SsUDtK4B
6lRak76MdLvdkGcxmd8Dln3OJ1T0sxBbUXbjOKfWpUFPeJRiQ1PK2f/8zluR/16H
htQHhbut80C6Equ6oEQTVS6wzaK4ReUqwsguMwLKTLzk6cF0LhYo3whlzbBx+0Qj
R4wHZ8ip3zqOKgQVdYi2ZU3pq8D2V1p/zjBhZGUCC7IT/vLNh+YZfVMlTgICsbM3
Ml4Y5FY4gZenlZTdEyn8k8gfntzJGa9Y+Lp2JW9g7IrlPh19EX0ko6vuG2wc3W/N
2SYK70U0rw49lJwvVNokQ26Ddnfd5JyTZNSTVtS9kHruwXwaIhk5e6/Y8frbvBYX
LPQLooT10hMcYaxgtGSJTyj/+2AkVxnQl0xj+7MYhN8Mi5qt3ZAa4ZKjDbLJNWim
2HpG4m+vctZnmnKF+LMI/94un+nDXkS/88h2OXPxmWSjb3lq5LMlfirZpqKGbzPR
6fh3aAk99lzOLtX3Kd+vsUSUVIQyZdBiqz2zf9yDzy/EHjbOq7avp2OwxubNht86
97gBRy+rqkZDMKkvNB/Sfa463dSv4ltuz6677c5A2X++l8xpPwB8WrQ51/SLpURY
Jw+ylAP7NzTEyjRJtEH0e39PvUEGiFQv8WWuDHE48rxg/IbLAN5rQoGJK9Q0V3Wd
tX8YatGntQoeUlu7qbKcOZG/Qi9ZHvPof6mr/8pIQSG284a0SKPimE4yt4RoYLUI
vmw0LNL6+suUyB7F8NScVFgLDbsipNDqg9Nz5v48mAzPc4ZWjXC//1n5gVlUi5oi
8Kg/cesm/qqRjKhiw30tjqaqsRLrYVNPKu7MiOr709NZe7isKCHgB877KX3n9aEs
k2p7wHN7NBW2YdGPNzaC0RSzivsPAOrLb12p1wCPE8hHj3x7TqZ5bIILNSdDcGYY
OS9lmEyNadF5YFK3MQCrJK6UOR3iA2Lk0q3/IWcmA31Yi93ovvHB+2jAuQv+L+/v
zNW9kw/7kflZ4PXome1vJi57t3P7IMLTpeHmUP2lPl3AgZbnLuAZnJZsFWkHCJvj
fIqD8xrwoy2ARTx0LbrRzXteaJYL45BiPzoxOOqRb+cRtd3wSbe5Mqr1MdOWdt9c
3LFAyp+WPkUrJGDrNW10ipFdT7yrUD6cOP/2QByS/F9QYqFmojf+akZaGtQVRKBF
W41QW65IOG2sgXX3kpvIpMAmZB1OkpD+YOusUIc4TaF9hKraL8jMk6RGW1LfosMj
CXfC/3NUk6nGVyLeCrihcXGmiXeZ4UiEFj/dXZvFaVe+S0ylgtOID+VQmOELy7OX
Mv0U0rP6bJpL2o0rYdptSNykoYhiTkvjF2IClKWAWGDTjtkFR5Klpdsm12FV1Qhh
SsI5h16SBzUaSW1azToDijiBiBH+hmvVWhD8QyvgnN22O2l5/T51vZ4LZs4q8vPm
lSTzqLvHUu7502WLvi2vojF464FLDBGnkRsOI0pIfk1Styd2acapTKL5SKqNTNzp
om+tis/t6KQl5IS+aba4hDvUL7IXj9e0c0cWMyoywLxFPpJENPMN0HmXnQgxM5Dd
CDk0/5DvsxnhcBdy1Zqp3XlPBumN4ApARCcJKa4TiZ7roUbMeO2O71soMI8uh9TD
M2CEfi7GmJr0/c+CL8oRuUV50gKomdVa6qmFJuQU7O5XYF1CICfVg09UDuuMQGUA
9se5M35/e9V0TBzgXiPLwMlzI6uHX4Rgw9zlqDYWJeLhq0NigwS+Rs2flam0hH6j
hxpS1Zqpd1FFIAvOlb0sMXoSljUC1JBQVWuPveb1VbLl34b/i9YG0bWBa8OITIUH
ypl8q72f7qZVTUT6LBz+xHziiPq84JfKWy6Fvg89pThzta2G3pEQhbkQgJBujZEI
njWvTs8jQwTXVgs4fqasY9PTldo19qEwa2G1GDLQflX7ZyCrxEy9RKQ2IRvzTOsl
WaK9xpqLjc9YwilRoxHBRYD1QqAwH04nK5djJwTgRICKtVX2bYvEJj0KJ4BrwkwD
q0SaMjglKq95RVBiwTWWAAxrCZEfPHS3FY4H5fI9ic6sDhgZ9aaGFVc4urw6/r2h
5Z0UvWond999Fv6xCdT0tFKrfvi5xxFQWZZ5Krvqr9goIc+xC0DrTNctg5OtCHoP
xDun+MJQZJnj19m9HyOSdM1jwQggTSBVSPvs9MsjAb0PLaS0K94ff+l2FtWy496D
qi/vpP0HtpQmdQj0A1cuYwnhFg/WjJBQvY7zfZKqsMpdFT/pWL+8RTXq1gLyz+Vl
JS3FqunCX6oKSwmGsL+UCchC6LuxQcifiHhqf9s05wsLe6qakt2SQWprv1T4TAuJ
T/gA44LevbRSzabe87A4W0hF53VaQS8r9vpWrDhUYybIluO7CuqoHvvHLLzBim+X
dE4tXQ6EspZ0CI/MmoH+JX1Hzu23NDRe0cohDBguxVwHzLEI8JsJ45OG+fAdGdeC
Rsk4BKJi37TmiRF6yzFeqjzmegjtRthGzr24s5dzo61HeyKaFmZsTX/6za9l5xHN
aTCtqNC3EmmVtUWraV7Czg/+NlN0NjPg7XYuh9BG3rNksoKVsd8bKe5JqDVfgHW9
SAkcCzgDav0CnXSi+F2nympRX+2VTC7s09wao63GlLsL0CZeS+9I6TpilhmETpYS
mOAJFe97tZ1D9720JWM/9XVsFd3BRO6imRVo2t0apxZ8/baZKn1JZR0Ekn5p9P3b
6n/lBOv9Jt1I1W7GT/K8rOHml73cX6I8nVwwQvuEvpMehZXdHYHBq+vU6TGWgo+5
DB1/B8QHkcOB4g3pwjQC+/iXK8Y6JuGHadXMeTPz/AklFN1+iPrYLLBASnQDWD63
8NtpRC3jwssymIDkEL97wBWjkTfIlv+XzfIQYRjDKW6VgZaPoMHPFJCZJCHZjzT7
I5na8jMoqzAEZo4QqLUaFKhbWTrJgIdy9mVA5gTlEFNCbdMKDR/kqSFUKU0ZniBG
jNqvkyG0DTNvFEr+P2v8j9/+TXNbID3RFk3svypjdrIg8+cDql2aS/HZr4K9nVSX
sA3JHz4+Wt7wTi+2gpoJceR87Jh61glW+FrRqM+p+VVdV9wxLqDzgt4jUYsRPZuI
Cpd32pMhYpd6p9C59gJprQHZB7BMhStYtuLwvhFZeUPxu7dm3pjlevZbLQ1RyjpH
3zKyX5hG160O1fy3OndJS7/i9vsy/Urj84/iqWbs2K7QlnB23xEei8DFidE+r+at
6EPSq4XCfaHjS8DeKGk7yaQSDgtGPNp6QSKpogmm/Ar3MwKAiHSwKmQv+vNdp2td
6aboXaMneJp9YZ3T6eatphYHhX88M5o7CXyc7BwBLeM7mkmWvuXLBycvhUfvSDTp
kqOcDp55fkSuAPaMqNvb6DuP2ie3wx1Vnh3p2BmvAK0dGkJzNXrBhWzVXWartXPO
K3qcci4tnbflqCN05lBUmLRXS96m63dFKeiBs+AnU86YFWPNTrYyKf5x3QsmI8tv
hmcibG4h20htOON1JqVf9hnyj/qh5wVl0RpLzFzRFPT4KoCizzxGiQgOmGcTwa4P
ZWkaOjq9q2rj5rXFZINxRrECc2nDCY821pCdsZAmKKjGnCzmvMN1Sd3rixF7GI8l
E23LBY3ggwNLYACTmmK1PyDPiIX+cAvkKtx5XEynEnoA3BWgoBuoEEbjASudgCdh
+P/SiU8ox/H5ViAkk+gXoDrZXqsdx+1/xwW2kJz+bAUcTQBH4JaVX5AmjXDgIYZl
blJpZa6EsJJTjnSsUzsvUtFMFS8s4F+LDGtiMa9pV7wfKIBHnoinuNbfNM56Xi3x
DUgiNCDextx3G/8FRwNAwk2dNnkg9Awx3sf4YVyveYtZJu0H3/yaG90zKD7lRy42
XijV757kiihcH/6lC7tlG/aBBMh6AKt2lHm9lEhbAngPisLySSgcunLRY5P76loY
6iiRtNh3rWpqKnz/exDj3hsInWuJgCilPyGE+xwm6GV+N2y2mVVz+1kO069Lbow5
8Vmh6fLSX5jayvbQCEH0Y9u7yCuSvhci75PnmvRBI9M02gj+wqpT6Lyo4Yn5Fu9+
kOssscWXx/X2V6dP8fg1wwfVT0KByi/UZl/5avYrbeLfSUUmXb3IKYOvZFz7LVaM
yZMBdGBjjj6VQbn6AHJL+krY3Pf+0qNj3Ne2p5+MYozeKaDGQpt46A/hNc3FN7as
Qe+cwluKkz5Gt3bHFApJ1NixC8gg2goX1FFiP6AM40mYsBgDPtRm0BzjNhkBDLBZ
HZFFz7ON/DdpKDRr1pYa//VuvmAKgPp9IMqQLJkcAuTMamPRHc1ZI3e5mSV8oxJt
CGzOs1MHrlMhujW6rNXWVCC9ho5oXTqLaM+6Q3BnIrLpSpa4ZvL4UWamDTJhsL5b
EuRl/w4+G3Ew1W+lWNTs9mYUH7A5n3IzTMNBzyDPvBEbSoM9z9Vh9Fs5rdh3pOdv
GD/7oES604LMbSn+q4IQgkUMQK4xspeEAX1Ikw9wwqpkbVJ6wqJ5qsXLUEBp8z9J
4y6pyfQi05ci5gjXUQJ5Pjfi0Z78i8lPb5onR56uL7nqcmkT+MX5+TXnkHGSFqSV
1K5zOycgGMUsIM7rGY/KvUzRggEu1GNFgumh39zbeX1W7v56AQfgv50+iJA9YFIU
0ymu7WD2TgilxhWNsuBrzwKw0RaXd9FFI9Le48cOPAO28p+xufrZJd2OkeQqUbnz
0XN9TgGhQJlIRoDjX/cFJ6NS2QHda2HX/NjiXS++BKqooL9sD3WLRrm4y7tbZL4D
gtLyxFDZ38nWx3x7ZO4qv5elHz0d9KtRz7wvdR2fA+0zUu32ga17uwhLhwb44b2/
5cq8nA48GQLjfElkZafkGbtpqtTRD64egdhcPKzcsJMOq0E4IJN7gRV30/4ASBeW
Qmp7LlYNz/HIenZuieOw0Vei4GTqAhe16t48V1Dp0ES0t0QU4dSN8FJ8BQlJIZFb
vGuUogoVIxL5CfDJQtZLbiLhwnBGV/X/kwY0y8gtOKGMhiNevEGfeVstdzAzMAAE
dyuL7fWrZ+G1khNIiMGmbuePqPOAGaPY/lmRQ28uXtko14Pfe4DRIYGAJC6okOVQ
9BZcAe7K4z+sZewVjKE5nB4gmSL1YLb1lG2KCwlGChlWciLzZgPrbFIEYfX4am+y
v4fUDorAGw6YDi1RWxnAj00C/QQuMBuF5BqJxSeeTCjq6VPn+ynk1Q/PluUYmGKU
2L0KHsqiSHyvrV+/PrNDq8wN/fGCRr/vc6QKKiKUdaE+niCo6SJpLk9oKgSHHl35
8JX7JVw5yjRjDWiXRSMGJG+rnMaG1rz+2nDKo4iYwyn6r4q3nAd17/Fs6cSEaCDT
NleXN/mn+YhCXpb4Ig4oLEvA5htx4KWHMY1rGzzT6k0G66HptU8nOLcdmrzrAd92
y59sAjRhjBN06sbzQXnQSnnwLokm56VZyjBrq3rXoih9tl1iQOzmJ1fUkFgLQubu
rUoPougK7RiDSYLZvJK1fa0UTA8LGW+N4t53BVwjMgEotAOkylbKN1t8FfjaIv1D
QxFxyNYtzKyjN/OreailDET6d/CnOtHf0wVkh0ZeIeGdlWUi6DelPxQTmOGPnqlG
8TH8cszQiGjr3sdP2aF0qUExh/eYSuIA19BlMQ1JJMRlGeR4vcA4KbyB2GY69FT9
ab8i89s8KHFu80ITAivB/VZR1frtRnuGoSqRZGrVYzTtxyLQ5I7GEZ3bWadNJfBW
PAgOgvyd+8j8Az+UxNRG7HysR95uT0t469aYxyBYJ3xdUxMI8IJwTaoL6JArB2Lm
mFh8Ik2P79UNRgwJIpIVuzPLoz+8NFG8bC0NLxjbSHnJc68h9cDqVSlhlrcDqXPa
yWyOabpIjGz/FYi97vcc5lorVorP/yDMEUyb9kAESWRtOZ6vHV1+6Sf3geTvkf8l
I8UBQzK5s1HbG3FUCU0tiK8z6lstQ61ddaFLRosERQ8jBpLSvRMDdfKqlOQ4rA10
NMv0YTUp9sOfxj5ByohpgXM2dpfm7YXrA82tdyMD4jufyjHcu/c4Nh5Y4aQRzmK2
mVjztCeIOhWowzZq7XvUlfIrZ6VJPjB2SFS4UC/ESackshPDrCBfOVgJVi4oKohy
hik4B9pIc9RKbbUrPYGxUck/Nx9L76u0ubRoCi38Q7wxgtQMg+MDTWWklggwwSSq
N31+MSBiNpYR6MU/evOHDLYkFXeTHfr6DwuA3c23osP2XktWmTq0DLHOonDYGUJv
jgVaRmQLmEfSM4TmxTerTiFjIUvTb1Ezd6qQe5+sZgDdep0L989Rd8AYj2tw3SyC
DZk0r6GSt1J0oTT+KnZcUdKMSc8J0FirH4Fs1rRmfksco4lCbEHfxTaGnnp+oh6h
531F0yaiUkylP+ZvoOwIaI735wVFZkx580E7QQEXn4A665Jv4v915gLqyLyMLo7C
dTP7MmShNv6WaIxmOzf24cwXJVz3JfymCrr45kESn+uJCvRpFF3ghGgtcSSvorQb
/Z/OQOG3t/x3MmsR5fbHEGA/PcERaa5+yGgIt5vgpXGIHH2xBihq81yz7DD8Ch0J
fyGQXC4hoXG6WaO6f/TSKPS+Z5ZkTdyUV9xUUA3gfGd6trg6RtKOkeuyO+LXu3wD
Ra6yIJXVf27GfbLze/2Qu7v62Iub+aN/31f+dEANDFxQNEf/CXWlCeNr1fhHGA6r
tlrhQmvWzvbiI6v7XV0R53uxnURrC7ZCkrLXJ1sIxXtLZwI22dxvkxD6UpmhdYA2
2Q1SyjEmyhc9qVBfCiY/DgQB3tQPTCYqo6k+JYpwJHoWYeiSsi/3yBRWOg7M+dv7
ODi2siBNxOvu72WKigx+byAlUPELEat0RGSrBeOkxWKhcp9kU5XsEZqVvXsImPdN
qzABgu6VXbCXIR6Xfg7J+9GxhjzsclXbOYjulQdET3qjWaNUZ3lvQwAIhbDqaXtq
4gMfE0q6h7m1pW21+5c3xGaHotgvouyGaRbuH0aB0Msd03m40KXHjD0VbpIU2YcL
7LJvUBNB/aZiJqGVvpVe2J2BxzDuRKMnKPpY2Ja44+v4t/ohfiRf43CGFcI7IZWg
pWByxTbmOtTkC5BvMO7nMSOTQmUwxyaU5e+q9aDq7S6wXl9Sbb1DpYUhbn67FY+D
VX7yWeHrObYkhZyn7QD87Wp76iSRHNX8/RRST51cqygvfhMZpRyifHDA8fqNkwoN
mRcqDyaBRoVYXQeY2Z2vdC34FJsOTQeGWinhd7NAzk9SCRXl5l0KI206jqgzymTM
rC2nzmrYghyXD3yBFz94GxeNvWu6hj1lLm0ws9KsPNNqwK0FzoavsCatSYgNZspl
99ErR5UcBfR5GthVHmrX2tNX8JUVra/zY1b6fLB2EzcnaDdvPXB5o6VNqug+1ypf
+6Xls5e2PaXvLtAuiHm0gczGr/cu5iqE5KRue6uZ7EBRQzI3omdSczeI9PXweNND
ri0LyTMg6vvRCOXYyvq3MxCjbU7xCU7FFOF1bMDiaAxn/37/MieXp0170GKBswLE
FzdxNeqyV7HeytHlqHB3yoABPxWxkNIosvbIM5W84QNMk+ewpT85sLmqsDJs8M8G
o5tfhBiy0PGBFijDD1V7k2EfdfZdNvm4egFZD+usYj3JW/fbJJ6gsYm9fdN3w8hh
SAglInO/ABWQydRk2DOZBuM5m/2tWo71ezRjy88h33iCTm34UdmIPTRUPPHrlWiY
/q9K35srzqQzPp0T66urUsAyW1Mv8o8Lm6WvsTSuFm/00CtfR+vRAdHnko5RHgCS
w5Q9eVufbogyzYthVD66ffGW7nlEnvPvkGRDFyDXr5NRvUhUgm6j/AxosXYFC+20
PZ5nty5flTmHpy0KjkxxDLZFbgq8vaHsxl6j3gkU+S0z0YVPqnXbrR25kZFEX7bu
sdpgqoVq6UN237XmzHpnd/rmPXh9meZ0QvQotUTJ+31og3eWDzTjlyRGyqYCpBcg
3FjD7QBNsl0kDr4o+0HBwgnITZhNOwjIbSGHwEwbccRB1xnXjeuIi0nkGHPWqgnl
eA65rY31ToaRpGHjAFcZKQzRTbGN9NYoSuDCf8MBXN+DA2+5NmBgWJ+qv2XeTNeG
kDRqCCrNVFUW2VLhVIO70zYlRIco+peMoMlZi9/4lGvvMZdyZpl0n3xm85mIH2oP
rOXDeOZjZaB9bul0ewx66e7Fh4eaB+c286qZSydYksmFpsSOOQO3m0Uamk5tYsFa
6pg3bd4cosXb9qN+y4HNkykl3Br36TBq38Ti/qWcIKSjnEM3+jV7KH8y14Hu3uev
KRH4RUWX/6GA1q+7mg/vRATjZ8hcQJyzn5NcEEJ9KH6/FK5jHBp+y/cykno4yqNe
4TCqgL3Dw6v4gHGBODsE5gMGLfRWBhtYS6Uj2gGo4VFJViBCxE4GGH1g4WGus9yu
n0KI4zqz1wLdISv5tnBD3ahdo3s8ysEVJDaODYyx84Q8z3ZhOZUYdQDCoj9mn4+S
MNVaN0jELzv52hAc0/QgFCgF/WhYR7mMheMzgCAaJevHW6l5mGf4FwFFDErFq+Fd
9LFUYgZKXw8AOJ4mGK+husH9vPVqAGnHNLntrmLGwoUYXRQtOtIAYEJLzeShOtoT
a8tX8LwqhEKPrWrKjnL9A02i8kbQS2m7tjGhLS5SkewcXVyaj6CqNSOvCV4SIDu4
ZgzmVb87607OQDPhg6fPnrv33wfxk5ApR4al0+kjrgtpT1Ielk0lAB+JuokkRCwD
o3P2aEYhS2zCIpVB6DlB2C1/eJnVHVCMqiSEd43B//VsDv4BLIgdtHWtxWdpTKNk
i5OVDLb22TmxAlVylp2b2jc7XoqbuwvQYMrU9bB5B4NoTMGr+Dd67JbTtQWqKMwx
Im6egnGaOFqWUjSYNxYLWyYn3DS+9BXb/aTei8ZahK4Adx1rOpn3fhWaWrDpio+D
WGoz9JQ4+c94Rw2Ic6FTN8i2GQMtYiPt1Hcl+FkG9mEVR1EboAIQPSrVorgdKULK
H6V90HxuhZvnXaHVM0TNTUV7RUhwgNqL5J/hBhhpdLsbM9osW3/2okoNNrgTLGRB
rkx/j2iZ1isz9zARVZm0GwQJOlaMeedTqjmoS+f3DebaOY1Aqyb0D4KJ/LdkjxBo
C/zrGlrGSVFwOGBXx19fuUuHijF+jkxm2dxQXzb204y7GsXj1faHjEylIEUy34kZ
KEdUnc1lulb5FW0cglYpb/81PIcZU7SsIu2tuYynz36a2UIYoNWmQH4aKb3yRAIw
DTvqPoi353a9bRFQRNVne2NO7VvI3OXo11ugYSKo0YU0S74oqYEAEkwyGNnYkf3A
bUhX1v2mWIiiNVkg/ljtfTo/tDkL9wYp+v3ZnJl2FJXpIiyLO/h7mR0uwqAE93b6
BPdXHZ3oaenl3Y47rwOtVFCCQ8qS1hCaGqHMsxgpSZ1H86L1Dhx7OdDiJiM6EP+y
L/CxXTAe/QS6NuRDj/xir02JVjb5WiQUC+RjN8qAj/HJ63Iids92ncOyssVZ1Y68
QheqL3D5k/Bl3Yw/eEfOvB+gLXMeR2QYpi2BCx177YHlqS8SOcXf3cV++pvHABbj
VkzeR7wsszKgoN972CtUvGJURQnSgZ304PflAuCFiQ6I4cbDrjB1hefr+L1n/XzS
fcUoLVqQAhu/e/d8BHKodT6a3OWGw53L/fPea0wys54dnzXzoOR0r/WUCvEkdXaR
rFLh564JCBfIqzeEDtP6nqikbZfW6/+x3XUqGt4t1FblhyTCTNwp1MOYvmP2a1nH
NoOCg4Ps0sqUQyUX6SNwrO8dQsjpWLAYf5hNZMGIoDEsq/DBqUQTXvSsWE+TVOp3
oAn4pP+lG7OJE8Jez0u5ZCDiQJrC13BCtmCfC1eY8Kn7+W0xfzOcigNdVzJgl7xr
Nrtdl7ymFPa7Bd01669SjfiQ50WxNSudKV9EEJvidwVELv91KIESjxj7la9frxaX
WF7n3K1XPhpXrwbO4K3o6iu6kXV3uUs2ogEpHfiJnI5BQecKw3Ozx7kUVIsx6ZUP
WITYuaMjvvIlXw9ytInk6C6TR8ij99t+t/PskPxXyix3V/Exik6Gq7IKd28HbC/0
sIM99XaEkWnaGaPe3ScEwUNWDriIg/p7wZtoVIZce7fy28m99E1UGJthJf2wSdg1
1+Qv6NDNSh3yasaHE/RC+kZuMjDILb0GEEuAiTFpWjzp5zkgAihDRQrRG3mpazH4
NLyCftAEy7Lol8xvtpkIkjRmW1GGL+MQCpH7x6Pf7ekIBHl8fe9H5lAVaXz8gaTk
dVF2/afQomoPHhm0Bmh716bY61vnhwBp+52sHiDrFgpAG8y4PKN5iiuOsnf9Blu2
m1LiHKu0eKHDoXX+YMQ5uQsLVF+bvlrcFkse6kiCwH6r6i4rBAJ8HNjbFq5Rzd/L
itN3nVPDYkyBiXFpj7DvB4h2nHpesH2LoLdSCDBu/XfCbMFNF4RlB6DqtmQGfxfK
oBY5ca0/l5v31Q79aAQ+n+XHNSHfU06GoV8OWG0s6hiW+EzgA7Pz8K7+ijkQWO2E
iP4p3boCgb31H1gbQZUUxZ5AvE6tYabRxKzDJ3SvOnzTsTXfte/O92wdnqjIueeo
uUGOmVoVQMrxEnxM9v6Y1OIrO/8zsDWyrqs35ObODg8dMHSBwt9YikTpqZIN1Kj/
vM/8G6cLprYab3SMM/HJjt2ozeUzoaTIMDOf/gdF6ehv1OtXbzvlGVVXHkW1WxsW
TJsDqqEcilIoXQ6n1KpYJeYwhCpzzW2858ClhSzIEmR8UIb+eHgxiQpH3RzQkgOw
VsCkeRkYfllbvmhiDw4vB6MuRB4vKeaQl4CfRKsP7WXzWwDq1hJkI2kmIzcb9yzq
QoMRvf/4yzwqv+6kWzlRGo8zFLbY9u0cS88MhG2kYVAEOVuFjC038/1VS+gJ/bP0
n+E4T1aoAqEo3J4KEwhpO/6yC/kVSUnlYgzdpscuB9OMgS9vPZj1yRc3ceN+OFQD
sRYXV2p2WjZI3TuYP9OhqH086sa6dR9CwF7/mL4l3w+E3Je1hilvWSm+l7SF0dyG
TN9JVQ4ZxvZvgdr73aVrV0nbIiuld9/xrI7B6IbR07j7iw3qKHf91FzCed71wtOC
uE4uXbdIR7H9QLbhjFupXJjM+K+7IEa+xEvFEYso+coWrje4E5d32A6VU4Z6BNc+
U/f2/ZRnbps1/33RA4qe5LcckisbGDu4OC2JnihMYR6mdIY03nRuAtLBtR8Zq/a5
oifJTEhG269BdjAtydS0X8YN34BDYNrNqNCq8GG9F7YHHwCHOGNa7pM+5+5CAn/K
aDXbpSEDCVAKHpUxffS/kEIqE/nvK6K+m1vTW8/zO5mDve9u+WobpLNyda+yaLFC
avEnEPA1wiRey+ZHfgL8auJUrfJFuQc/7K34JlXbQ215iOhOt7Ujs2v1oNtlZVIH
A6Tys2Am7N/jxR4M8znFHADVr0J9lO+KonPtoOhGdo17okh65lAZ1Bkakna9+9IW
GfWGndlUUe9vVAnVc6OSHe11xUsj/tzzGHQdPBijOttaavmXvbgsLkSNSrAEAGXz
NuC2JlwGx2FMfJB/qJK0ZtVlSh5vOM+1sbsTXgx3m4bkphHX0y51aXXN/E4tFj3i
g0IKA968UIdUCE4BYcUW/90E/LpOiFHDRmbZ8z8tO040BFZ74NEU/fygntxphUIc
yE5MikyJLrC2Irgoh5bC1VoSAPomvk2EbDSXR11FFwsuHyP2yewRzjY7y84kAx1C
DCSfT6Fog1gTTsa8NWxY7nC1Ov1uQU8ICz5xcY5Isem5L0DuVRIr0chGb0ukrb12
fd/wOtTGXJIoF2W344RQQu77dfbX1fISM9jVcyVONqv3xB7kxa+ov/DcZLytEvkW
hUuJCqTBatraCEo6dibt19dMw8OMdla5m1OzDySbZuUtf7EqHpc8zyiBEBKDWbI2
CLc+rKZhK3iBLrveZmPw0uhO6vDXdW3Dk2fD8N0ng88KwcgeWzUlHqlNGE/AYdTB
TS1aR5KfsNRgsLdo+TQ1Bvh9Qye17EwpjbNb/uOIzDdQeK6VgtD9SYDXikcGpZq9
1hIo06DaE5cjOc/TCElK18fx+px9h3jGDwbwa1CkxnHVl5rTkfNnhZVq/qV/hWZS
4PRZTp5etTqB7awtODum7bHxl5/jXvaJML6Ir++ImL3HZs1yHrRoRy9F542V2d0p
eKim0VDVM1jtOat7UmQeMeuPcI6c1EJXCVtqFvAQmajU/XrTGAYt1opQ7zpWrQWr
Kyhv1JWdKD2slxHZA+tuIHuZXijxkzukWDzh23hFQCLeKvSM8yh2GZmZUehT4RV8
lM0loh3Ekqv1NvjgvrhXLWiyBmE9nGzy6sc76aar/1vfBKHx3feMAUqD6N/n1ScR
VGPlo/cDH7A9HMjtHh6Jo8U2PD8Qw77so1XoNplXqJ9oO1jH5fkuviXBsZx4fw1r
5lLD1t00uxeWrMMmJ8mKO89RhjQZNL9Por4yfKG5rTSXNaNQKQ5+viD+t+uXU9iZ
XxWApu+oPMW6shfxZcJ17mA0dgzWpZkLlYp7mbl97kKPfwd6gn4HaCZ7FZf21Uli
KjJThqqwJz4ZXTT8Nv62j8Fozn38PUrFliI0glOVcMC9czAX+JBv5Y50hLBxC96q
0oWWgd65ogW/2Qo+f8XdJaWvup80OVU9ibgfzyTHnZ5m18lO+BdblNL3TvQ2Ck5C
WptxReXOGJAnhGjQKBpSEESjIPeJCm1vCiFoPF1aCr9GRc3BxJxX1ZN8qJS0xnhB
Y96lGvdVD3fVpXn26NfHSfotUBQgr0+Ffttw3KusrWJ2kL6jDzXjHwdqsDHn7+7s
o3sPBhhPB9SGNgSq0l5SlX7klCy9NdZA5N6gd8uOmpGNK+tcPg1kblwz403oLFtM
27GW2OqGL7mkaxaYQzcu6HHFJSHZUCut/cMZYbNMUiHCp+MebMWlqngc9NCKMx9F
plUU0I3bGM6pJfoD5+XmhhHNHXIvKxtW5cKfmB4lITJnH3YI1rNJM+NdoMpKQy9Y
Ob1BvhRq7lgtLHmdzUlsb0/kfB5BeHVSjdfPjPzyhTA79O/WbarJTFdBJmfcV0QV
Jn4JzquLAfeJq54rWnQrv3Ia865NPnrzFhRcA4Bbd2UO6w+Hz+6co0RKFSGo41T6
6T6KFM09uLDh0V7aakm6w1EqAfl/NlkLa8Ei0+sYBgNFFhwoqMI1IQmIw16YlP8v
+BN1UqV2oZW1dBO5+cRHK5Ex/eBVX1R4vn3igTaBubLGKhHoWe1XjmKyv8ehG4lq
iXJNorgzQfYbyfXphErHnMiCDLshztGXX4yqouBhSTZie5HcpWhaYw3q/YWTaIVK
/7p+VNAF+7C1yxVS0XmycpftPlJl9l8+8ZiOJksZIyLwFAnQR9wrgIkyq0dGCw9n
UcfmfuC5AZJHlUR1M5js1v1lXr/eWwXptCXzwormpIUvup4hElp9W1JGrjHdLau0
dFgVZ2eDISnyrzKGwsNP/Wkn+3py7qHVgNNNF1IaR4/bjQDI6rTBGjJFMQirmg+6
gewPjOwflu/selbMow3hEHarZvWZLGCQ/uGL/4SO8AUn9WJs9smoYOhxuDSfkE2/
Iq44kYqpLeymL2BY0Sat5vsDdOv6I65ajQOv2EIktCc//JvluppPg3UHy5TLxDm3
YU/habtUd6frPS1I9u4AdApwzmZCrMDI5bFlPDXHxHOERq/8tMcCAsplyPYkzY5X
3/fcCz4YR37hJngH/r2w99/9cbC7cbuzJUBE7ZvviSpmBxjO9i132kpBu9LK4E0B
bTAgpqCpCRI5Uo4CCYSeMu9P6QBcbVOmrqQCGHflcPYLza6GgIWykqSdEDLxJMyt
KX+OfzRViHCIEJDXF33WThi3ws6hM4vJd6hIuZGpQz6O5m44TziSfirXrBzzxFmu
+gF4NrHodyfAU5Ejk6KTNMhDU67vi+x5Z+UUGEWCQlkkqlFOiG6gKNCz34g9RnAr
syNNDIzYvBNutYiStE1hhHFXVv86HpbjEgthKEMrDyYIbPfuFfl+2lfBhrYzLIMY
FzJ2FBzQVwoaqIg+qvBByXbg3U0ZU+fXATUnum8V482pfMdDqPG4hYDFGuKPJU0D
VoBG+2Pq57aZ29hS1h30pg1DW/yL1M6TbMKvDoDEcKISOvTsc8J46xdciDTse6aQ
rPxM6oUEeN5Cazd2/FqjLSumDZ8/zypuh1EKO3PL8n4FBIunyXghPAK+zFcvmfhc
NJPly+9kNj4aGmveURq9A4XsGPfzHpmE42hWN/eoyTN5YBP0PjH4JAtVZyYRsqD5
o3c2UFFcsLz2Ke2Y/zIga82qO8X3UMFL9QamZjgKTG69RJEtZhhxZ2TH5oureQL3
WTS6xyhWgLTjli2V1kDMy2tyMET0NdfSZdPzevWrGH4tQPGi3uysVu5iIJCWSRMl
EET/OSZPrFcgNimi6czU1rDaypqMCk+IQ6+VZ138DPtL6wlV9tzgdoUQSuOFCTgv
4zZea7LOgtzbMkeL54VoI9NG6pAvz3yH3BHIkYeolpoNYF8Sz6q3emHKbXQsdPCU
SfKJnaCyfpkNOfqnUFNX1E51l4gYOaRcfHawFo/gnvs7UoPHyVm8RIVsFpPPHZ6B
hNY5+F7kzTVVH5NkuFuY+OEcDo8geYINiJIx4JrK/3XDYDY/ZvG9xemce2AaLt3M
x5D5pAY5J/VtzXDWxygFdUWaCbT/dQiALu5ax+6RvwmzHyUIDck9k8k2qSqbvlFu
5k4DkwZEli7/afkfY52q05qFjZFAyb75ED6jbU0ikaWMkBwtSLZt982DPHZv2MSA
DGd/kphtyVIcwLIMG2xmhwQbiOfN1A2byCSLFge4CtonLx/ER33xU2fciknnWyDw
9Injrb3gKd7U8DMaDQ1+sId/RaZpD3znoLyVrSS90iyUlQk2Daz+2D+BwL0m7cAI
IRCutzboS5qrkWTCYADRFNBYO1PhU4X2sUBxRGwko74dTAyhF0eC17E4NWc48hqL
dFDJFHsiupq7vjDRgb+8XzqKsAIVlLnsoIQwMak4yOcpSkef/i6t1yRgEJlyq8mG
OWbkqTIhsapFm6c/5vWF6N8t1njGiJ/1bLV1/n6kSsgAq5kIZ05jxYWaKECETo0V
WRNzI+g35ukvZxBF8kLUG+7IXYGOUPs5PpXhwoQJhP3PB8WBwqzzOqfdmxzfk28V
HlQOPBUgVa8Nmxiz27JVfUOe9O+bkUMK8Pi7/qvo9pbtKTMxu3Yqv2JQxsAbm2pk
zHEaf2tyTsVM6pJYQdhR/+kJGXQyTCtoNK70rKh4txS5Ns7onBi0BpUJlUsmselb
LqSRMQcVdbbyH9N3kNG2xthpEI6O73YiPk62bybbia9XjuyJUgs+8i6Ym8Bto79l
GNRGE4u+Sgvj1r+VfAaxHPXp5bYO1j178QkWGhNAwxmOys1XP3kX+h9TaAJRjSVj
OJTmgxS8bk3fA3zdHOiX2JYuPRrtOfQxw6IYqAv9Z+/gB0+aCpWX9182ALl2KM0x
sAfnweiTftwBSwekdaF6H6L+HoCzG17H7eooJTxO4Vhl3gojHlqiFnlf6vwLH642
W//Fne73ZbzTLevCJOefx1fuVdsAU3DT5ZMjQZ4BBvVdjW8X8eCuU6vUrO+D80Z9
NOMzpf+Eo+6lMcVfdyEjSJkQHtbA4/mdO57KGVkIfHQ0+PoZgjeRf+a3ctPk2x1n
6KhieGwFXB5sixQnT9+R9FyTcU/X7WNcSo/NinpAJ40phkgY7uFzajkKhraTCEpG
qkhRchXFBMZ1UqvjOyZCPU0XOlzU8VDZ2rpiw2g4Ug5B0B5zXYVRoXkXZlKqGWvm
J03gRzhImAqEh3U7zLFplcjfkHDJHaXzpAcYbp1cCoa8KLqcPz31f5r/jyewRGko
x4H2HhIYQbJ3QhYiLaAYLEepwcIqKF+07fhR4ZuY9OwTAhzIBlTMvWDLz94EOlSj
oHjc4SnciXyIB1S2cuZ7d9eEcfPXjln2aYDZvkRUDjB6qq4HE4gskoQ86f5Mx2rG
Jd2ke8uudsmTaKmrHnDhOPgcCwCmbs2Bf5OAj8STLdlsHl5rPueG07aLwaBaxyXL
8sO/bsvaRJuH1lZRPrUtOVKkBRridPNfE3sYRI02Qb3I1Rc6AK4tW0W37DKyijb3
VWgwXpeb5rxyR440jb+Ku/6COfMf5Cj23Cyv42frOXQd7xu6fV5kPk9KcZuKETnE
haQr4smGFYb8xfsnLnKTrq35+JWK3p6iZD6WEPBWhUN3zQUvy+KGdeumcPmEOj8b
jQArT5/nGyrMGlxGqq5sX6Y9A8JLj74uJ5FI5TL6GvfswQxKbsurzUtMOoFB6GnH
U5BMyWbgsUtwJ/AdVQqJ/xPXj2N83Ca1Xj7mYUaWgTmgVQRrabvrxElyPkyUgzkj
OwmSi7Fzk9fkaKmSWmXo3kd4DPUYm2ACy7C6dbdJNE/mTgCfRpS6UpEDvIdZ6MzK
oKDT9DUrS2DLLKRUDO1EeYxmYF/xcjrKgeZ2nSU9hh2o9wBNoRwTEvEAG9myvaQo
q5mGPOa3cFOBVHifBIQxZwmAsti2RH7YWNrEPu6kpQsZUPUmiN+nXKPhCttXDLGK
Qf5XeKAw59wZbz+C5S0+gUfpglWqBbiyo4M+UwdMVNhY9MVmoM0NeXet6rXhOCew
NEDrcH/+m4KdifejUOsf3t35fhq6mZSNGfoAYYyeImg1uPwSucDysqubVOhxupWI
TqB0jyoXq5sIb2DHiXJ0dl6ffDGDa7qtaWWmuw9/VnOW7nrFXRvDESXY8LXYMkdu
eQrEy0gzTkIiVJuYtnSPanETeApwKnVzhdR4xD7ScvGlR1oU0LNhBIO3eALPQ68Q
MyLkI97Y2rpJUNSgtYxBqaD4FrKNykp+84VppZ6r5Y7zYqSBM7UnZcY2yUA08vim
Ob84XjWFRhnz1TLoaW8sbCRroexJJ3ebxPAfVKRaTONCq7L+aSRWH7qYoi8zZjIz
udWUF1wadCfIPO3z9bNlZRKdl5/lggKV89l+lPvPw3UUwnlGXruENU4MMCB8aiVF
Z9+snHO7j8f1/7c09ZhWI/pE9Q9ZbiqAZVyGMJTUQQdI6wVlu6hmrV/imv3d0Fvu
m/5ORLAYiFsjvz3Cc9aJGfISzy1Xc7aYHFzOJih9RKbWLXVOvNBPXd//X0cA+4aw
WaFc1ApXQ1dghCRZZYFHPSeZmEqvk1s5ZOwbYD/HzKJc0SAzx6SjBvCH2k1Dlinc
wJ1WJPbEqWOC3KXkyV+78L+FUDPs0LYJUM4MHA5sCuY38wiUXHh4AUI8v/DLOc3D
Mq0rgA3UgZlgmg7PaHsg8Oqfim53SZafFXRPgK0WfpD3Y3E7ZB27a8PVFwDWwl+Y
aSmiJvA8yUqcgLAXfuxJAMey5/zjYEsQflBQ2TMpjGrzcQ+jq/yB66GMKtzC7qw7
MwnSeoMrgmKpaKUxKSa1CRkYhLiH3HV3cPvVne1LUgYznuUzeKaIlRkojL9Og3UO
AQiK6ePiJdtlviY8yAQ+BhWUjhvOpLa6/O7qENI8V8zNrMFwCmJqf5/QehiT6ys7
c6wkoRTuBPrM5RS/WUNOF4OFmEl+GBDiPnrVga2GVfHBSe05k6kYih1DFRJWW8YS
kJxinRvUwPxSuB1jh5aVbV+aWRRpEWLK4NmruBiphQr7XNc9kAgkobNeC1QZ3Ong
RHRDHIdHwMzJ713KyNg4EXer2zrt/S5inOaR08gOJwNbeja9rW9GChK52Z7jOyoX
hgrv4TRKrXVdJVKIfIgTamUqFD78UhGxpxAR2BcToho0S8TkOkZLhdKTCFZRLF4y
migdTcMI+8YZ8+VisDDytbaEDkS7m0Go2Fcz9tk+RLfAKFIklTgE3fRQHb1v7gj9
83nmsxVhD0KM+W2pSjqNikOWj1SB2vSehy9Uo/pIvkWBjy08orvRlRwQmIPBjmMy
uzs+1y8XLYaYHEMJH5XPcIr+BGdUQWmVuPcsj2dyBPPnLzAmOlN5jtIt2CaZOYyU
cEUeDh4+osOcg1cG1p8k+yfVQP7qJsgm6w03vUvjXmcBp1R3HwhZ3H14KXwmmsc+
nZiF+Mld0Yo+l4CAuplLpGlx74sQQG+7k0XXsCZfoAnxv4LRVuWORtqAI6pOOLqB
OAQN7CBwm/lG0TuYWIn1nDu5cG6m4Sbb6L7gLlugI0/YEvhM7CcdADD77IRFahQf
PHT3IsgjBfELvL5r3reRSc1YLqhMC8GDoS+2iI00LIapOiNVF5kSYlNhOG45iYK6
EX5qv1ddXJgRt3svmZji61dg+m0ke7I2yah74gTfJU58B04I5JmsBDRkWhIOGUWR
YObUUJPgbcNaZ7PMjitNw+dIw1kOcOO6I0QGxpNEzjSrLmAdVZqsxw4ok0ETZPBd
mBFHml+UnoLTxrTAJIpJ1qMf/lC3AHiX6SmjiZIM36mg6KNHV9GF4aBSzq6jLqX/
7U6tMuHaM+egY2dqCcukt1NVqmBSGYdpZkioHc3q7HZfC4ggwWsOtkn3ooRh8vlb
Y2OGDt4LRo5CDPZVAR3F7569IZW7GeKP4bYtx30MVGmH+ClgO28qBkH/icOhxEmq
LguxPhBULP+zK2ISojYaQ1f/CTJvkrWQ8SjHmV1TfKL8kmZB0aDMJr6J3I64uPUp
UJoS0KYL3Lh8BWk/X9BZdgsxTZeDLHwM6LtRO6Wk6YCwD7I3As2OzO9tD/wDHqqr
b+woCITr60iyv725NSPN6ATc1N3/Ddvbj9ZyroNdntiXLmCVjplNHvnDIYpPQFuP
JCxqI7+9d+rs6yJGgLXopDh4+U+qXrqh1CnUV7ZBwhoiHCLK8oy9tV4K5qRks3hm
/okqOZCq67stmFkMeEk2Hm1n0k/hIwMjoRwT4EvsJS4Y+4KoPgRAWa6QljDdDxhD
nht9JXOjDybLO5sqn8VqjH+9Yqfb+SzSpUE8ybzQJAVMj5B7dHewuVY9ciFYM/hg
zB9N9GSwPQ19bkvwjhl6LivGS9EkkM2Ghcx2nlVK6AmquR/0qZVd4y73lfSss331
xhgFKKVZ2hFNErYoBkB4VY6jjufIIcah5Ve3gyYrS6EokPqq9jcFXSsvfwdi51Dg
COiuSImCFNJConCWjbX4x8+h86n9CrP7jlGILhibEfqMRLj6wkULeCMishnf5A7Y
AeuegxV1gxZLetciGQcXnScz3W/6JS9AaCV9ihOBo9kKuKM/mAEw+s2jspK/j/zp
azRybOxtry6cJbCh7agu1NOCuVnFaeKxrvv6uK7n+vVaetJuCD8qogCKhAuO/XZW
9p3T5h9xbN0EptpsmQ+EesIyy2nwoIkIHZPTJ/yaA9+EiSrqTlF078ob4yFizrah
9j5m8mve0+s0yl+eSSaJizYcpanRiLmnMHnR3A+OjuanTEs8ZTYqPTTj2VwZuZfH
oIUatzPd7G0TQxmifd74cBtOVuuVKTtyFu4UjoeqexVAeaGl0lfVK7XMOtp9HLpY
JcmExjUIfSgny78qpq/2/LqacgUIYPrhJhqdWhR6p0WLiB59d9OMqFXDo2Uov9Tj
E2OalK711IYHRM3Mi80HTstUi/lrw0fHy2jEz2irvwfboV+T4vBJY5Y+n/n/wbdg
2sB4ICHEQM18XR05nFNjeLrng2I8He5dTqS2aBQLeR8M9BWaCDsLjHTWHVj77U6m
uQf+e4YbXxo5a52yenO/6ENTCUHxEgyk2Ih/dYDaxyAcGfKey0VVai6JZumErI/B
16gBfffRLr8CPREe2qGQURrRKjgWkW6F0ZwDH56ecTKMNKQFYIsXkDN0ZGjuFoSb
Pv3C0rW92UiqElOOnHoTohFYC1qMp5r1iL4MmjEikN3A9/7/YbZfplD+98Bst1n2
c0Lm3ebbbOchIGb3maoPOpUaioEOnvtjmM9PlrHYCmLDk9npT6LMNLCHUs/vvFkp
uRRQJeTBgZQTgwJWR29sKP5cb2QyDxjGKnx0Wnf5CRp8hqwgMznZbi80btfsFY51
tHHN4m3ZpOlCLBN1sJwEQVAfdF+ZhnZrjHNAUOho90RfcLbo84HwZBWl2RjxuiSQ
nLqHYPp0msy15+VC60SOwcb8mRabcZoIi4zI2lnxbldCvtqpLKDMwzqpwjQOFre+
2wjgn5EGaQIAXCyJ5k/22OaHl1jqGHnbHDFAWSTQ553fZU+A6c51OMfVkVMtKQ2G
E+Rpm5Qmjv+x2nTVUkn5XnAYlFp678c2HS194/HUwBsg0seYMrXkUgEpN5z+Tyvp
/iPBlMzDSKmn0kbkqhEsaHHgpDPbRzJSau5HtVSmswC55Rjc99VSX2hC1l1gWkxF
F2Soqkw3SmIbYzPmyXAMGTPF5pQtQN186JEfZi/zMNNWdJEgNaEEwTKsquvKWl72
Ci10JsYNuqW+DhvOrCvSU+VKyUxX+ZfvZGjv6H0f0iF008itkTGDk38zA7T2Lylf
JMPtS5hskQbJFHnDaimGerx8LaExIEbp1drayLWj/UA6jTKxO/qkG7LaOSFXp0j8
zygGXRa/EG7ladrVFEUdBN8TOtCNY01Jkvl59tLLjcgTqFPI0yO5ZslSXhHtId7h
oInCuaWZ5mlCt42VOuH3phc85sspzv4mQF9lkqj6uu6YnlvP/NtMb84ELlZ5SmMQ
Ya6mF255GHa+AHKXWWvmKNzYVcyxqQF8Vot1660hP4KD9HaWCusTUx41v6JpHz2f
8QVcyMthqy0rOdgZn5iloWZ0fOA4fs8jZ34R2ibEREEgYkHk8irFGC/tpXRPFmEE
T2DSGPgrDv6iJqhJzA6vVlva2TN1P2d0cepSdDrnNl4VO6nAiosJvSnyk5KPhFCr
zYKNGXm/h2IgXWeMJ+ieVkhdmlJNiE/rFuS89OZyXZhV6W78C2RYTHy9zQdruWBn
w/JnwElqA75mKhFfYLrd9gFdn1/TLJUbhMU0e3YkHSmChWu9Afpc00ioyXNyd3YM
hND6+yhba66JvWTj+k9FcXKMa62mjOHrP431W/Nvy7fGt5TI5uOz8oGHPBwaBIJ1
eRctOaEseqvhD7yJEtue4X/VIBY8cgXDBHj6rjcsGsOUeqE42piDDtYhmP1UAA4j
ksbCHdp6NpcwPVHLpCmGBhRPU4a4693cvHChnqIAbmhwh/jGQhB2jG9h4xiDF+Z6
Ktbg/dKC2fF0KVDPvpzdEGG6xINS4A/ljoNMQyzUo4OYsQ6JkP/qsY+7tPmUxIRk
JtdZKN3Jx4e1ybWViGQp6cqf3Ike41coXX9qwgEOzo62kiABK6sBN+x/UvtxtgXY
x7X8A41E0sOfRdyw3TFqBQfdnyZHMjy90wTAA+UDd2wC6ox7FJ9IhHxORPjIKcJr
UjQucKDjcErYm/9CEQpZiJ4sfc/eQguukSXEqt9oLEO0KDiuTvPPaTwtKmPTbD11
NDkrcVu0D0kwxV3q2tL3AS01B99tInd+Lrg+rmeCfgCeHnSuSeyOcjEv8NOG3hBB
nA/O0eGsV8wqYdxMOqXoOITCb09bcH/kMdtsQnaFO5KjM4GLUaap29kgO7mZmqpJ
lDtegkOAXp9ywlPbcGUGtvRUbJoxVbOkg6VnWgdnnKuP27mTJcocA9W+OzUZ9c8t
kCVd/98LRR3f3+V6rMVHGashfbPMX0Y3TgArM2ndzWQLUwse+1Oo9BQyZ2I1NsWv
6FvVcPTqPn5KclGSSupaDFeSqkFUMZtvwzDBw4XebLypkqjwEdyoutX+RkLyuC4H
bhHxNNfw5m2J1sI4g3wPZG30Ok4PLB+d81RyfEKvclEKlVubDUMdZ/ZNpSRa6tpn
U7pf80Z9ZAyDXHLQ4cNcGlN/otR32563UVdM12c4bHF0XTjLel9O15apGbUT4McN
O/zAE3S7Pm2FQH7Ar1w4LKyBBeDLyd/8A4cHKHAmHb6z6I5hh79g/VL9v+REqqyO
44CdRh2XfHxmElLk2B/0qpZg2rxd8l+qA6MRLX8B0ieEOOeWQYdKu4VC1nWJT5XN
4vo8QDjuNAziTz9+vM/lswndejrvgs+mRLBDmGTamSvUB7Vcg14ZoOrPHTf6mn6W
BrciZr9sn8ZoM1rs55OjI9o6VFcLabEHHgLnfGQ6EG9pdUV5F1C4tzIHtgM8HFJb
F3UcVYlvFuVqIsOzuLiLzJCLoVHNgxxCmPmFW8G0AXB2eLfOBkH4unL9AYv6JYsI
ewUfcogWbA2v7zKSQjJirAVREpRc9QGFIgJTS4hl2xjZb/JCa/maPwioWXzOZtcf
8n6lYpCAD0NF8wOfMfiqlH1u5OMUAXF7xou7hJ7w+vK5Fw/f3n+W8MoLWe7s3ap2
3RLlkr5Gkl00cWTw7iKbFr8RLKPPUjxIBcYofzHWaZKQAO3BNlLayheEOiT1Nm/M
GAqbgSBI7XOi/c+RIf5gphXrAqQFkoTaOgA4hTl1c/14Pwveb3wXdHuCNVgP5zK0
OjwUxSdkJNyFFyPuxKUWzDTWuRAhkwYXjw6eJaNg/RgwsLec4lpyxNSHOLBnlGCG
+4wRWwD1TL50QbJX7RUW71HrUJiKBsOVCPo+H/0iTgWvIOevxGLM/7YGgznIsuOJ
CsV0gz4e89RtgBDH3/E3iLsGzGnAqgeGMF53vhmqEbXNpDc/4U/M62bkAOxeTHQJ
B3KhPoKPn+PvFwbBjH+VP+F5qTynaOfMEZNCWFuQrjcBKz4JXHvU+7RDOF+qETVb
VID+nCKdZWPmnc53xnj9qlxn52BZwj5vACBjMTVVrPoWJW2lzkowqrh1HsHWdjuC
51c7z/CImWWGk3TnNyX52qaw2ci/HwssDI8WVd7aBURNjYy6HL3WUS25moB9AqCX
u28CwZ6dvmZ2bW82WUOkP/sN+zpzfnue0ASe9UAOw1+y6OUbsvmvYj4/Z0AV4ewh
IgEBdXo3uHTCF+6crZPiNQ2SWqOnkZLh+tKLFyMuqOmImFfIwZ/W+iQTCVy+Gr+c
NRTYDHolcl+8ERfrSvTEBdbZmMxv7TZLgbMBO/hmTMdxiFpyTCKdtCNuHfBLDzYl
wHK5MWuy98DglIHlB6iVJwJS2GOQ0ArGnNdkKRpGa1suxmBXLo/w4Ow1999CIlK7
6HU3d4QOkRGlTZt6VkijP00YBs4FXaNcHj8tQuOrhuJ8RReU2NF2snIjq3tzRg8M
VEbDa9M3bWepSdUIUHU39M6ca/nlS8KwmURTGZTdiwBcEDjYgRj5eQxRoP6ncWcR
SMkwgkzs/+WK63kiusjNNEvwLOwXvO3TFINfaXIVfnFwDiw2+ND+uFW/cGDqqvzD
MEpvgtcAZ7DVGxJAEEu49toYBW3Ma1zc0kPkrEwY71vWtXM93q2Ku+t65vp3uquS
BuhGBqlfUZ2uIhyQiCzrnd4SPHfeH22kd2aUxY24ezM8u1OxwBd31tG7XLoAnjuc
U1xaEaZ1f3nAcq7szvKg+SM2hWsJlAseb4ZW7f8XqtYac+V5ga9knn30Vaepbv3a
/v1wUcKNhYXzb3zm5iCI4MKzTvJ8tHF1P3jNcxHKU5rATZWBcYnStL6pm6tWcwKr
KH5RFmviTeiFvZibbu9BuiABHZNN6kxMDCsS4XeaUCOLIREvWUkf5W5js+Y+TtmV
H55L7hnzhDIjYj1wlly37/tqvTvu7qkNR/4Cxs45lb6hYK4QAUNHbU15Pd8nYHrZ
+6TwYn/qkDMsgdm817wxlOJCkGiVxgWWtzhvyuO7+dmE2OKyTSlCr7ZBo5i0ESmw
2JWMnBMBzD/e1Wl+97adNu8rKEe7jMFHweH9IO+j+DkrgyH6b5JqPmY567cH4ICI
CTe131FewNa2iPbWA3+6vCK3q32pfjFKcAfc22eFkmutkZudtynMSEQMQNUK/JFS
35hy0liQRTeKSL80exZyxQeEk+hgv1Rpefj/uRkPfsBB5zMWokT4jiYvAug77m1d
ptrp0QwJ/d8rEOMzcQuVvwq69kapIfce2NqLfeJabsG5ZSPr6jgapXH+5frrM7e6
5tZuzq3MRaxXZ6UjMwMnqXTbT+4rdxxZvMgjyf82vfO7CPPeu9yL3PkEGhgMwE+Z
esshLC3dh8D1JAbxA/ZB2pEyG0BnjxeZYegy19d6EIyRplMxDvVCwNdJyRWSxMGR
Zlp3clWwnAuKGXruKRhzkoOnjH1eBRDOBHlsB3pH0I78n1lkAgud97RM2JBIspkJ
jbhkpHeHWmbBNeg/skCpcHsr+FzC9uOlW/+Tkwdl9tiP/jYU134GiCCXGEd/Y6Zm
V6fkPVagRG2u2euapDC2QHyNno4OdQjblsneTcMhfjag82dAvPmdSlix8Y7s6wxi
/sS0n8yzbnG8Ttnmt1qhZGSH7OldDvNs/+OYoZRczPnsIq4KcYU59ET1hoaTVzlT
hGfG25GQsevR/BlYchQ8miLuzR3sCI/Ll7T4HAVSki2N6aLQwfQyhuZpqUwMc91W
HRe3zDrzPch1rNfqy3n/8d8ycXzkVpPigK+ldQ2TnJO02DLzC/4CexYDNmiRY2DB
3m273syQ4ux22J9QoaPEpEbIRqk7qEbWi0e7uRcxwYsx/g3BURkFsMQEzzs75vXH
B1KC+zaDMk8HEFfLF28scB/DihYeSDoFNqdXlA6nL326XfEOe9cAUcHXrPFXi8Ht
r302/qHJ7jquoZ0YHBI3YrOORRlFqIkxuEZxyN2HvK+KDNiHB7umGkh0S3F3b5lB
KS3TtWLp0XYLEHd+xF+pTvdeK53bzDX5foYRRH9x0Fag7IjPVHCnrdNboZoSQWx6
CX836K/Vtrfjrkxx4Sb8tmKZGu2Qm9UZFcqFNhDDS1N6hfj6SIqv0x+uNnLSPR49
aFDuoLzSLoiw8MMQqnftxiyqeND/4XQqqQz+5qJIqGMxluFEjciY/mfQbPhQcXNr
7mkm3ZUWnwi06og84djzT8FzW8fvl/KkzcjwisR2CnSo9k/jSo1tXoBaYVbHCkmm
6I+04f45JclD0mIRRaJ2Sc32zHNM1cikQ4dR2vOsjCIxrzcClKtH88MWoFo6MHbo
VWDm0Bo6SDzecPKQDjk2iCnY0Td03blO1OXec3+j5Vwtz3SjnAPi+9wzNyMCM1Px
C148lqcDVAIEhNTR0jvHD+Kn/cnol7OjURutAWgbwXK1HbsxOyQiFFkqGnD3D/BQ
JlIXtPKMk4gHHH5pWfWBezjIMpr5X+2fIHk2Cv9bym9+DJDZXMppXkWpVYFZBPOL
F6EzaxtaPDYJ+eQlouYBlkrtk0ht0rvwoXZwJqK1ChGEeles0GnY8XkQHqPAPEfr
1NmBbCkMX9o/+UF9pWUB7oLXpW+q3ZM5CxAEvcObpZkWoQslpArCu8iWGQNvXclf
zKTcXd7aONKUNmpVYlLem9XFc36/3UucbdYZ52WlrUYkIl+8qGZ4KXAjkhVNJ0aP
XNAEYvDCJkRa9BzKzYFuF+wvaWNot/hRYBbnQ2deGGS+5qEBtXmwchSbUmuLeCoH
/9CYNRO2dIXceRklt9IXwT8HBqz6zspjjgGisWLEAsvyDMXujTYsAZyTrcCE0RDz
TLRE9B1wbAjcN/GtMb6x4W/joiuVhPvbKpmSP6HUYKvw8q75rmckNlPewhhnuTKG
lBCcYblBBYruS8uWXvyjdtvvbPuw7P0fwfFEwgFJE8yok3hivo2MqdVVv59frRhy
izRdr+XByhUWgXAuqbRMhlesUCcb1M73AG0c6CFq0rkHYtazOXvvO6dxxKzVFCYS
jTZRSSyje3ZWf151FPMdz4605hetsNLXYV0HPBcUBqYs9JxxqOCkdlWhJwSbyzuh
agljsHyufCjQukFycps0ijU8Opl8ZTMDHGeH0KdWPMbmk/oQuzJYDkjK1Fk4CegZ
bx2vT5Q63LqNG0M1M7kWhokEY37g4u6Ka04vr8mwNQxbFILNSG0fk+VztCwNi265
p7Rty2kiMtXbKc7oYqR7OL4ASQQtieSv5s8u2BD6OZsioavGP8Swki/V+VxQ8wSh
LBBZ5XQXwT6icGj4rMQ7oAH1FVXJVvha02mmm0YOp9TfSOPyAljpkDXplnIi3lqp
wSYR5+JUY4qqYrRw9ng97LXmRizZxwCCmQ2f/5O0vzTUX2CBOslvhc2kL+4Dcoqd
YUjsEgo29HvMU7ciNFmdUCQ2nbFLUDthJgXACcNkaE7GQTA0DMn/xr/ihp+LwpuR
XGNAD8wDZ9QJ4zDtOBJ2C1iuBfDsawIDE8kOvUeRhVglikC4CCwteFaefb+RH0RO
VMw/Ke9bcz6mItDVNG5agh06Gi+ze36t9Ju1ijXxGvvBbCunr4jRIs6RaxfJ2FWQ
/ACWmzvDYTkb7vWivolS8XqBGJegyNgBw9FM8tRiZgwjOMD2+tFom1xUS89btEf/
jnJZvENYEYPBAydRjpo+zgHpNs6esB6g6IB3iOB9YCv9XY1gGQPx9AzPUB1a3rna
lXWpJJcBn61csDdErZ0zMPzWpkQuuZ8KeiE6QYlZs3JwHQmbP96kqgZ48SLJFTav
o6LR6rFU/beygfLbzCFAxvd6i/4vnhMn5znWTEzSNfI7nMN4VD/lU0Lq9aNPZlo7
sEs4muDEH/PdnColcBRMzBsSS/YVoq3FfITsPDR+BqepqoDxQ9FgGMmJ3S50g2nZ
+4Saeml8SevcTbgj14SXXNbk4KkUKxeAgXzCbGXUlWIydeuEB2aDRG2fOk98ua7i
oMUsvlcmVAtixpVvadAQTGLMlpjN8Z4O0wTluEudQUQFkquVH6fbX+mM5JcfOkRj
CtHfUtUqc6QDauHPh8jVndR3ZTwZI8QphuVG5fwIsh6sM/rrMtBCVU9J7rW/hHl9
mfZZzHJ8ulQSS13jKp+/qvbtA3ZNNaaKaRq1+L42beS2UJOJdS1rycql5uSfW/2O
gJVxjcfGDZghXMwhXjrMqjZTi3yxcIDEiE6Guc91GAucN8KBsew857ODS62xU9NM
RY65S9ojzBLwGRl9YUSfqyRXNJYX1Q1a1jgXnXnB9A25nADtk3cGdm/VhhGj6ijB
Czfs2nYvoxNrNY3VH91jFD2NhBjTSLm9v4Sac8hZTLW9PlWGfmD7WsJ0+Y0iMO0H
FkidgEUH5/xZEwRCGDBmEXPlT6fcGrOmbxSnvZmcNC28qZE6qypLNnqU+YINkpvI
NCK+qUf9q9JvUdcW9FSK4eynFGEKeBcbXd0tN7LAaDVFNS25e/H17B4Ty8vmU2he
4/ehRPiQ395c/JM5QIZObxzyMYPHzO4tXiAa4f2M+WeHCbzk+ZArarNuyejdbBaw
SQfTGRQxbs4zS8UZ4fQYgWFuFcC8F1kt9aQVqLBn9h0IqJkNsYUeHaobveJqzYV4
5tpAAQbzLHhd3DefsYOlRnMUpw6mIQeOFv7YJa51DvEOvOnteeORjihV2YFal0Lv
NBd5cyTURXrVzLnfnaLbhpM7HOwfcE5W0FY1nCbaYERzgddQK5X3fcDmPMgRjP8c
szIOSkcSuoVCoURpZbmFQYc2XwjyIsxNa2HkCfOljmirq/rjR3iNsGxomwaKe+tb
7Wnp5lkmdxMeRjfn8tcEY/ykd7d7KhyFWGVDjqUkmGCQVtb5iVF0BJbOjdSPV+ty
zksJGDJMQTzUQLhyqQ/pW2NT6M5MOo0OtRCVwMOYnZETYjRQmj8Cd0sOuMi2J4Qk
ZTPIzCj9QflYCzdnsZQcUKAYrr1RJy2fZvRKz7zaZyEpT1jOannUbs5e/q0BqjYA
QziodamTT6UuJ5BR/e9hgisTtQ5qnbA70lYzBVl7XWVt3NoB2uQxPDNnNnOYosU7
s2lzBwErdkDu2zDjYTFW+Nt7HTQPAm+cqjrrzGIhVtr82ONcNoQvTg2jkBKH7t6Y
V4uxg0ymvgII44OdmTDoPXCoXA/9WJybvmDxSiNaRghj/UrbARpmzXHs+veRdL1K
tBrpFWa5+pCM/YZKRPy1PYjG+kA0I5r/FQEVr58umYOpbU9perPOx5znW5oi/U0/
V6Ge5GWBCKrwNbgKYUJikpBCpEi3xluolOuTJqzgI2kp4px2cZ5Dyf49beXmMP1i
k8N7Kkf89trzpTORww9tSdfkqDZ8WkAiwOslxDclPPDx7vHDfsOpkAYSH3Dq26GV
EPjzaoP4SjLV3a2Osf1mxUCtKBXTjUAfNUMavaQLwU8LbP2NIRD/l+SPceo2z+NR
angAQqfEA84xiYzvnPbo15yh4+qap9aYi+Q9eplJYHpMMFk4W2U01XAyvnFaKZiA
znwUJSG4tFzSSzZZgIaM8Cdh/e28ws9Ike+VduIjCYazp/VA+na71toEjk+3u1lU
h7V+XQwxYTk0cR9xkPxneFeTD8wnY+qDgChyMyyBwul+UOEkw25sivOQZCx9r90J
Kn/yblj3sggoRuHSvViPZpIVgsbLpjEnkWeNqPPVn34v2FedbBVy0cjLD22Mt/aU
VJQNJlenBAF/mCUCJgWzv7ANyWEUHu77JQwuPuQH5Y9DWGMxF6sT60qlntJMaSB5
ZBsWIbTZ+ZCZ/Nas7jo9yHmrL7pDToptRUBhv3hT62PpFlrEQzGkMps8+foHYjOG
ol/goykuCqrhIe3HJvGv9wGAawKe7EUXLYd/XrVvfcwbrzrpWKbd3xTGvWlZcJEa
73doQLFfUtGPDZ1Hd5hyK3Lt6OCO5xQCX/uaCY7IKO0lBLfm9B0Ha1YbSMPTGncj
aMaw1ww3NL6iB92plKBHNjdEwgRO4w8x+HtpN/LKTY1CJ76+N8SCPoY45OhsYHgG
Pa4N7wFmZjlzho0KNeAhR6UhKXGmZzvcjGTjweBjHbhs0XysCdxYKUzr/i+5EVe4
5t0frRAOTN3MfkZvS08oErvSGIvyGAGDU70fltgkaDN53eaKWo3zvfFOo74BgsiA
60Dt8XCGwXpm14YkRyyS9TTDNO34Ht3NSBGXT+e8mbeMgbcDEEsB7ClsOCS2VIXe
3ragtdFLun5vflBMv69ayze5WvepmNHCjqUv3chMZkkJ5ymGDVX8n6xYRowryCWF
yoHG/LR12MIxAK/hDoolmywIP/uSGRwhzHw8wKdnTLEJCND6sDEpmfq0DHoMw70s
qQToo6pzgTSzCojJ5mydSMGTndrM5rSHd0B3cbn8OOAuyJu8dWwOVPNigi74ht8C
2nLJnw0W1vyzIYE14iitq6MDUrq7go7dE9w6az4rHy4c8olhgVCOcwdIs1ZJ8RO7
dRS6JS1Zy6P03TqgHTXAAd5k5tKjHZ4rQR+Cp4m9nmklsx+NXNImN18+mzJalWEZ
/A7W0qA2WvNicSbBfALUow996HyXP6pwoYRB9apu/9o3lADOosaqzsluAfZK0mTI
/bbk/TjrI3JUTHciGxLX2yyPaLOlEcMvSkRbUEdzRSDyY58M3+TSa9iQxcEvkTEA
Kv0rEqWsQpGg3mWFvgGQhrjupirMCfc73IeSyeLjidmOOhBqyjAVYlkygnrO8CUL
GAgG9IAqy5iaIdkFBaNJifCw8lgtHPTN5cpNmJgjS4LjFdndOhWVIRh2Rg7jHGpe
f4V/m/plGWES1O/wzelQ06AMEntUyMNvxKY7zJRsj9sKPDqFzEbA6+zB0ZgTkjrK
MOckW1xWTDM/x0uhp7wiYRo6vQMdBdbNzZBrcJ8uLk6g4ubU1ka0wYXfurg5DJYE
CByXJzXzoq7D/NLq/BifY/XD6V1elTdVu4GyprwVBeSgb/04Bd857riYr7ALgGoh
DA1sE4QkTwgx+wixEpen6Ir2PKDZ4USrqEB7OdDsVyl/qUeH+ODavEwDPxPLU6Ou
/7+FPiYfpfhrKgbXlxS6o9xSIVFZpVM0N5T5x1tuMTbCjAlG1kINydp6P0Rc5Sgh
Km7+HRih7pX1dkU3U23KMIiFUgM83eQjudPt6JvGm1FAAv4J6C9lGs6oUah5ll8m
ToZKJ9SLKm5Z7WLQGiOhfhcD1unK2iwItsU+Mmpe7sxXj+jBOdeIClUR6QljdH9g
vfn3TflAQU2g1dLEjQqnZ7WWRAZRDkOfjnt+4JWyKqdTPVltqLpAvLGMAHcVh1K6
bFigwkf2I4lyQ4dutOEGFifxgiy6TDgqNvZ6NGlgdAbVXBsQj2Y879xF1rvz8X8I
WtWMlTKhOxoasewoxMweLoCtLdv2WkJmYYETBoUEz23PTMRyYAIHiFwgea33VsvF
90Tcj6TaGVfsdbLQwdPhcu0Ey5z0pH/k18YdFxlqq7O4uYR8nGkxYbwrrl1wbwbb
kKmER5xUlqEyN/1eRSFB7O/w1aZFyIJEWPOYrfCFoY9BUctUYPWhQXpHsD93dtb9
mtP0UWg1ENctcuLrBRfL5f1+7nB+HwtoZySZg+F+2oH5ye4nnK2S8QFdLXftEsqZ
KMrQLcBSYkSS7IrFBhJopLBZoelJO9oYhxsiLrClYLLPRIoNe7CqgI5f6G9EAqMs
xv/sEDhL3Ic4APL8n8qEc/GpdJfcejtmpvAJQL+Tjrsoym6uw4HsGPsiyJBzps6a
Zvz9K0zpWPnuwH9UJXGc1Mv68/UJLGLn9HlpmcPgDCXjKh6/ZPU1/2+w9mxUqk5b
vYn2IUugSOSjoSxyY2zxB9D5V67WnFY8HAMk9WBLhTChLDRjvDm0XTuRbB+DM/5r
IkWpjh9Urd/qCE4L/0VUIAqQPlt2VE+JLsBJ/79O0+26zeiwVEAJ+XhDFhc4Z6+S
lFuqaoI+T6QJzhPrdi5MGW9LvsUXQ2Ixq2QXuhU8BFJRVsloyEAcvyQPVB2p9gw1
7lxQLwWjl7NTigchgQMCds2N9F75d0INzkYz9SurkPg7TagMjBLAfzkYuamAYoA3
Iqb0jEG+wVhx6M1DlyCogfR7sUuV+1Ie06TgO5ozgMgT/UaQVYKSp/bik3l+cfJp
yN7MWNG2ccclkRr3Ceu6EsDIq1AIgOE7jSOJbCA6COn3kj85v67OGWSNe5rgyy39
CAntxZWMpSy23hOkWy0DMYN1XEs5L+73k85xj5avPv6YjtqHBtcKMM2PbgSvqB+s
K8ViIWN6wO6OZIE5WkvqyramiXI9DItJyjoR7L2Zn/j4Wj52iTLo+DYflKLLLXLz
eo8kot2AXRDkvQy0AgXTvryJbh5wawJFEoLBZ72+6ZzOpCmEEgCKNGArLK6olFpl
fj9tUSY57ig8zutSIJ1og+P43drf0qB5lw5tcvnIjGYV5M7XAjuwuH8YSBJhDDaZ
5fiLwYP35SJiX1lQwCxyegsw2brrpX7m0+g3mbugnDTGSXXFhqpMTuo4zvFK9nFY
TuPtZWk4lT65WyVQZtMHxf87s2eTnmcMXY65AU5DbCjaMF97NJynw7Z6HcSV7Bth
QsIn8ZVKPk90INdIdqQ+Vu/nqEOQbJ2dhJX/+xSLxLYll0aij7/t9w4jAPufMB3G
bqVzwJnxE96DTeqj4451wZhVhkRpgnb8YtjMRRwf9XF0c0nP/h3jZbNxilH5TGWR
5PFSwP3t6tDtjNG0kCGBIXUzOnMAmzALWOfc9T1hpTTbBQkVZlTWv1gBTHo3Cgmn
GsMecO40eEtEeU6c1WE4ws+RD7YR8SOD03aD0rtMRhP+3kcTL7oZBZbxqbplo9bZ
lCU5rgCL4GIxfuGqUCuaR5Q1gJek/ROMFSt4bKCfpMGw5q+ugFAvEZDYifWpOKPo
DNlJN2jJt0oP+pDdhj9Sxtf2ysXKpcGG6kvjL7Odcy2mSDofcQSddcTWr+zghPCv
b3vVfCxYB5Us8PZxC2zoEqj2taG+aKASiANoNmYy90Vw0P413zKKuGL6kr7faHKN
42ArLHVXQhZSPfcBB5Yn+5z1lFU+gUCd0O1OjORIxEXxj65muzm3GBSVVMhLFbyo
LQBgLxsD6rWIqI7x/Nj7lGARFJXuBYcI8XgR5/xop2JRej83WNe4Bl0oj/i4kDUG
4coF11oIv/fPxTdqL/pgUlKeH5HhkzPJwgCiYsesSP8sohFmD+55ToI2FnMM63zN
hx5lKca8qW8Xu3ZPvfVXZC9bOafgGtmkXSjMoSQ0klfj0BKPm/KVhW56kTDuL6MZ
RlZ36OMhNw63py8b91JRaT/WnEVTKA7xQOUHiElk6ZnTs8IoDlMLgV5bn5h5besL
OamfiECCYlPn5O4ERfjrfXuvrujJnbtq2qRVQmwC6hMfEsul5xlPfiBhyEzFW11/
EbhU9LoK17/0/+RVVLjeBREQjS4JACSgq8E97271v/jz/UWuk5B1pAuIvNCcEVQA
IphydbqpI8ruPaA6z9u2YUILNNmyJ18LL4hxCK7gbp9G+G0S1H3XffQe3wcAajr7
yMuJjz8pXcoin8i+Spkgu28kCYNMV6Fy4tJjq/lnU7IqTGM1v3xixmSWiX5mbrHL
z+/0YWMzA7Q8jpcHsj9/6xpuiMB6nQT2o1OHiqAvYquFU37CZwWg2dhDDB/AyVNd
Bn1V+flHXwRKh0PfvhKYlzZo8L3fu+XBW6iK6iB1pTgmlqpnR/pqWww/QZqWr17m
CMBvJlKv27L1lxa+ypivUZ7zkW11OgBzCb1yvBobMOFoAo1jlPNVfj2LbxTWIRtX
i68+oPeVEzsnEMRcLwaFoxrlubc0wGf0kILXTNQNEqcXHuixpBwMtq1hvEbmdWl1
toD/4gCBIqfIQ+bnar929zdJ3mSS1TJNdZxBOVqEr4N3hvTlsy81VfD8Taz6mF9I
s0wr6AkYOcSCUOBGRp8rQbsVqn2CU5ITk1EKVF/T/xtgVR+/LXyUkub0jz52dMu4
Ym6SXLCazO2yyGkedU4ndi2Zz3VgMLohKgdcmgLvxsHRHtC7KP4UW9hdoWHVhyY3
clIGJm5c1YLJ00dPCZnbr9Q1KgbDOP2ZmRuG+3DHzVlv9Iq2C/H/F0sN8+IGdNrE
NgqLk+UbsDkexL4zoaBuXU/o6J6s+QtLozxzqOaBkf+SKq45iUtv2jocaZR4V6jT
OvJ7X+pwIYgbVSDbhdorSDYhGeuamf10T5QkthYrduJ76Vd4h5X4n4WWuRThYDE0
KIte6ubNSXjJ4LolJd751jtdvizZQfo8Z2R8Dhbx9RgZyzKjD5FDEeWE51bIkO7Z
xzumBNaTmkdn4PAtp55hiBXwtlEg4qL2qaZ+9eJjsDzIkaiK9D+O2EbLBJX41Fli
jDPBC5Du6cpjU+tKyBXn1aBWO+e+HXupgn14hu/NpkNfQXEjH1m/WHrou4ZUqsnN
IAmIwv6835m5lzq+OYsrLxYgcdlq1Hp28pt5zOWkkpjFdQaFW0ZTK70ZlCYtenmA
3IAAQ24KZGwrfwQwZTSP97vGiKpmzw/ASmm74Xe9bYL6BWYMbrNpWWBJ/gXkTPLe
S2Fz2h54MjWEnZadg3tW7tGmUd3gzTPJKxCk4KrIhS32p5kcrgXdaw9C6sbRRdtf
uMHmLUNd9Cn+snan9EjnJugiidsownJGcLirL0B+b6vrlJOKylnwi+xdI3cUnXlE
Jl7r0Tgot9gBUJyN/1Xf3X9n3DDdfyS4ZbP1OGSoP09vD/d01eiJiBhMupYbtbFV
ckuxRtL8T8GmZwtJ2+JaS9lNxW6MvJzgtpEKK1WBCGuCrMphTVMQ/VrrmE1MIVtd
X7dj7kM1aBwg7DvSDWb7PsLG4UGK/74UVMEGDDkQNRbf/bSKUhLreG8WdnItfBIh
EGP9QzLaiIS1f6MNJDfliAfutMcU0eQQCXpGNN8jSIBDyzVksLvPXPuUEAgfBoT7
48FAFvdD8hQoOnj3IEss6iIF2dydHJCYlJ4pf8QtYxFJKIA/Ac7EWuN7KcLib4+Z
oUb/AnyD8zXyWQYiY2BUJd+ldp5s6WMlzMW5M0rLzU63EhKHfcA+sH8JhXeLnCRM
6Zox1KtHG3ejXK+PrS6j8IM554YTQ+3oMdfJ5Cs69Z2sauiYuUuRTTgLaOhB+1yo
e9XLPEyCFoT/CYzq02werYtvtzdA6VbT+8fkJt57JfpVuNpQpqJyP8GirI4Qb3n3
MRxVb6CFy71fS53dnXwgoCUIZHRDikiCg/ILgszpQw/g5kXpj1L3LdTR1s4Qcpri
liWt8kl+ySGHECjPBhVnn1DT0Fd28hhPOzdHsJHr54QJL1gO3Drq/ib2vbSSoBxs
kar1bM0awzrf5kn5OQJKrgdeYzlPqfvvyoIQpbUxPYO/5TwbhoM4dG53vm66vQo5
hbRe+y9ymJVJV8fQDn3tnhKNhlsKEgxQhxbouDnlEGFEHyREO/1QRR45Dhk/ExQ/
WOEoOZlNtalEJTC3U2P+gFtZSKB6Mbk0IdLgCnq3wDJX0HVQYoOw+ZFPLnWAH3Pg
Fx4hSEirsbE4KzlzkgO+3xvqX5X/33UrFDL1P3W0c8BNGc188YsBHaySedYsq65s
DgGtZJrz8dbC2dJU6knI9zUYUQ8A9Hc8VlZg1+hZeFRFPJmMy1ncvdlMeM/cPjCR
yY6zpQf1fJE0g4dCs5+SX9IqINnznzkQPZ2WTWBlf0yE58RHWwRoGviwITWVc8GR
E8fCdKYRwGOPpdaI4OO+e7h4tFwfrMpdzSrJKn3T7jkeXX4I+BYuCqw6t2n/r2Dy
O27zxrhBBXclbGZrdBvjlFuOEyBjwXwn9rVSaTzS/YiKs0XX1GG3p1OxQWQ6fkNP
ARAF46hPC1w7/honlHQDYI7VB2diw85GOQdqfVrap6PYPDh0bPWnX5Up6GIHMOyn
yeo5hBheXgYrpszdYlwpl7qr5t/tVY2h52i9q2x0/hPBXHc3j8UJHbZuKn95gdpF
9CwlvyvATcFE69Yw5fi6pk5hv6OjuJO1Nr77fxtaiqsdq6xcjt8xI0YGuKVKY2Sm
c5ug1bxAt2AO5XxH2JAAhqqcTWa25EIRk0ynYJ0ltHALip0OVvYfd78LOQBinf7M
HH9LL4evsMiHlKaaQQinaC6ZPLBQ1gMCpDLP+CntC6UCQim3jKRtafPxaEHYNwEd
ta8s4hoM011vxaoCiUQr+WOWqVPDAA+b9Zqr5w41ROJivix3UR/wXqhmaNlNWawO
UIOwlWbHiD9kz9ERnz7s9AQYYhWPw8kvybO7xwi7cWVf4J2esHsqMNGaAORBj/EJ
QGPLWFN9gesQSN2yuyuA6NisDytj2/ipmp3ZqNT/5uL0LLdZw9KRe72Ce3mWAuTw
p4rsxH6hm77M2dluVsCmJvGC3gEH/DDUxkggr829+avPR+fIXc06cvI16slZWJeO
Hu4t+VcUTxojcHS1ZYLmuYIG2RiX4wVzaZwoBIQ3tKCDrg3VB4ERWGsGDKRtqkKE
/wYyLNEgCkpZZDEOFStZfnobe9yxnqq8u/R7cDhrlmh+yb3w7fL6sujG4YhpsQ0E
Ax2X0sOpyZUoD7MIUssEO7JnO8vidT91FmDXZiT+QKs1eQlnBPWkRND5MgEegUx8
GLeTn+yvcB+mmrilGDAqkAf9uxHG2xwnjGYFnormZN4rWPRzef3Y9FdjWTG7cTmA
k/pvT0P+bVQXvjYBf1MkUyAu11f43wh00ardEhRKkmw5bdR47PW+qpg9NjVyhpnp
fSaTYKyU/nlluMvlsuz7+nKHausbf6tQUTti83rLNpjYOAfrob/5KqUIBjNid0Ye
H0Ca/hCQfxLHc6SUu2FxBLu6pQhLhJBrf8srph7GwdfyiXzhKcTzv+DFyhB+cIfx
PlUdCjjSVlo9bNob3TfBnSSq4EQ6sfqkZfFeoH2CVxEi7KtiODJENHBc8mQLIQ99
KfP6mwY+QRWYZSzxu8e2AEHHo940y+GmILLvKUl01DA9XH3JhmfXwfiGAu8VbAl6
a169ggnGQ66Jljup4l368Lzcj18Yhp9j7VN8Um5aNekrS3Ixon8Jibcb6UPuriUM
PpIjPqKAXvG3IZd8+6hNU/BPMcsJy4+WUDoj9SMt8OW+1/A7BXAZwbitAvaOoZJJ
Rd5ZPHk92DUGv680dyDXwf51kinVuwF3r9RNElJdOrGg4RMAmJf6cG6KNIMVVchQ
J7ILuaqbA12ESqlgp/nm0/ddtOuuknetWLdGIjQ/6xdzoLD/cn3gQyhZyIYcbrDk
v4E3S/TP+upIG8aXqNrEFq3OnMyJoaq9SI/4djxFQA83AsB9pvNfmcQS8LPNjVVa
rWJafiODLtmCIwvERaSHFZqt+3IRClFhSCj6kFZlKkrrotrYeY4xvMgO4a/TJNEy
7dvYAxg6JVmwF7mHHexqNxRE/evQB/hDFWtZDe4oMLk8QbbiR/gjrmEBm180pI4r
L0IJzu17I/IRybRjmB3JbAjL5CKjYhG7D3hXFQFkk0mmthB7eR7ZSE4uOdt07/li
KEMgDGebj4lSRiqIcnPKtSGyIbuEFMznrR7qqtdxhRayzWvKKNGh0KBJV3XyhGgV
xCqfJAhl8jEX1VLh/KGWgefCoyLx+VjFhsB2wROxdIHmWVG4fdTI0G33MY8qV+EU
C+g1KENbenbE+xKrJiJn9j71L5NaQaUwzGx7MJLhLWAB4gy3R05J4eRHTVg1q9GA
mP58VFUgG1UFI82yAIWseh2QeWeQsk6cnBlTPPOubrm3qJ8WAZcU2BDfIrgN8ci7
kDFU6jXz5UN0fIiGORwyXcZSMTmI/a7NCtOe4cj0MeOt3ja12mPjvidQWqPg/TOP
0Tmx5au3M3HfefXk0NRt8k0yAvSIQYHp8AkEBZs/uiXUhi/l3YApv8eap6oPLpZA
Xx/ofAX6XReZFId3t+g7uBzPG5tXY3qWsOMlhv6vSE+WoqTV8ja2xG4epWh/3iMx
uyLzbCfaerK6QXT8s5hVBB9XpfEO8RA0duXSiyuMNRoljxGuUzqFiSxTHEbTRVE3
aJF+FKAm5mzB3YDVflf2l2Kijehc+QO1a2KzF2dLwBAVf1hm0wItEkp7TafaJfHI
2lVVCKOYDDSUufHmWBokYLp90wrq0BJqrVxSsewZepC8rU/UkqZ3aMkZnnX1DOgu
/Q0D9S27RgtR7svqlc81ETdMENaCitn667V76XUW9uHQb7Tlt77uK6D0Ou4H/zim
ucK6w2G5GlUV0nTBNoRV0lakj/kjpOMMQUBV5tREbzRrbwekVjpedl68cMD7Vedm
gujNDIs27/VVDKCqtVgKOP3zlIcvmTAYi+iAjq8p1K96r+x+IchqL+l1wgm3MsjP
+YN1V7h3IF0u4SngdLjjDIhcQntODB4mSWmhayFrq0IGdfZ0EoUrrGzT3HR8XceC
Yct/GJtJN94jsd72P7kTUJbolCH/i86BOmoSOVB3DXWz0GotUU3vf4c6ZW7ZDw6P
aDjDE11jhQe7Nf5tTYMwwzzm80M2Cl4xL4qa2sQuGW5dRph/8jNXn62SwM6HrcKv
+PK9L/JVrgnSsID/Y1jo6K6vKPZGjz2c3zyRYqiv28smaIOTysmbqZV3yIdSjunq
sq53+t/Ow6g7nUvtSVsOW2Pig/RMRc23iIe9j0UGHogbSVB4ypNWYFFbnzo538CH
DSKTrPoRRA4uy/pGLZ46YX979aMmjpCDqtcnQiJrshZuP/91xjqSyaWJN2w5CmrE
MkDiWB+ya4cGgMK+XRMUfbAbMnzGFMvc8bhdHQyEGPj7fCz/la9mLd1uVkc9PZZF
0fwYy8nA7k4cfkO3nX3HIqajgRo+Q8fmRiOZjxNQ79cD8PDBRJ4r8a2NVDxcwKI8
hGLquYwgCCVC1W2ITitD0pGs9kgn85t5YEau+JOctqNoetmMBhvxahfHSVwyTuOc
SEXeB1uFF8j0waxG41PvdCCPrygf5hWr3Vlqi9jBSYMpEMgf8ucOFtbZ9eMNjqJT
gm4VSer2fKMjF74NaNXpDXk7xqgGeaNhd7jjmCoIZvQavH3+PS3I0LK/bBKRVgIa
putp6MgQ+6Oje51kTzJedNB07XvtvsOckItizOrICdq2YD9On78qtzO5xWhgmKmF
doR50vA1V1ovOVoin5y6jzOv7q4MFkrNi2l1M7eGOJSmAGHKdPVRGNrlPrqGW+oT
s3UplPfXIDZcv+43YkD2E3DtUCWN8rTq5qiovwVZ7UizpgrjEa0C7CdFoBwf/p1+
238Y7xt09wf2Xx+cql7OTfLdKBqVUgNAKPIcanuSx4DLYkFEeQCmmTdiaQYxibL9
HYcghNpGatL7jzlAZwQWKlSKKSIJZo95kTmPRy35CBo3qatK/JKQAf+nZls7k0on
Fp/lqms5uno0BO8LrGRM7CutXpOMosvcTSY7vnBit5qS2WfvOBWamgBrEaqsE0TU
t/YEEcmr9pM3gjs+RHQwaZuLAQxXtA1ate/ET9yKY4gJBOQeaOBZLCwGK0+KnO7n
LL9olqWvB2uHhW3xmCi/U9HrVuEI1X+yoeXObsw7YWyFZ94yE+VlUNXuHQRddtk8
ok5f9Wh24STo8ESPi0FkTMFZ9yaGybe5ZjygXC6NiW/8pDxoSvEiP5vBYjDT7vtR
2GuDoNOFDYHhruxyAEzCX57jSEoN5zdlRm5Pvt0U6FP5SkGy7Tnypma2wzkMbTLt
ntBLbv/Ugn9O4nsVoww7bBcPWRM2ea7Bn0Iz9tHbICpvFXMRsFJ8ajMB8HgsMF0M
EVs+KbxMBwUZCi83c2wh1WQZIkQq2h+id6ulchcN6ehNpo+xO3LBVv9X0A+neIQw
6kc0oQD8Tx+agb3KTJntAj4P4rOnIgu96sHKNyX0urqeEj7PvJzySFTvuo9KrXOe
+EwKUTALODt+WggpSNPWS64/BeAcN1KUHZVa0Lt2S1Nn0HJLGd0Hgitihk04Ahn+
NpIbFAjj9R8bdV5T7yJ0rsFfWoz7uLBqsHxGp/OkUnZK3l+y8BvjHk9h7EE1myUP
viKMYnMhRZAre7cByFh8/oBTx6ENd8EMLY143Ymb3ndYQLgfPRFK8HgFnldb0fhS
j/uqvPSIuy+wNLMDxCdrCBxcUK64addWfkMJvtbU6MQ1HcnwrIlqFgcQGNqMjTFi
86qWMDtS8gsfu2Debqevc9P2WnEBBfdLnbRM7lt4AodGgQoL2T1KXZd2U77X8wB2
Rn2dS0hlc85LpX2g2tXclL0verXKaeUGIIGFKAycAEHwAmk/uE/yxemmORYdIeJ6
KqBZJ4gh/oHfbxQFIVkKEJjTTcY6hIB9/7WeJqc8FpMQ6MQzEEoQp4/ai+hG2MLa
uVfZjytEBtTgt6SssGuuDlTqUxW1p79jnOJSOBL/O9mSeIZJ2krxhTv1bfn9k54y
8PuudJ3/Py5X5sMfQvA775W+Xh40aDpdaVCIEkgxGRzQmm/buIWqhIvBuGdLHk08
/6SuZludMrKjWh6j9Rk4jx9ZG1eM1FxHtkKO5aUhtQWLZGPIm7c2Y2VfBNNeklTw
0rzZNNAXVu+BXSqXSBpLnfIv9Sq5CzjvE8a/CDGkawFnc8xCL+/nULGvEQnAxNs2
Mw5Vv3KRYtAIZeE5sb6U6kbyr0tvKyKTTCamLU75jH3iJQxsKNbCMde7YCAFpzkO
RH9EJZQA8NuOQ5d/WTrHMyJh4h3jsSq8sXQDM9qr9LFY3NCkGWRfTt5Mm4p6qG6h
sYb6B9psbv6si/VHGyBRsimpyBUbNYo/47yO/TqBf35ymzJXoZvEu9bCI8h5jPFD
5O9tXwcy3xOrF+qsvb8RZzrbxGGdXPZVluZI8Br3O9ZTxoo8Ho4jT3Dp3A4z9c0/
qfdiGv2AqEW7UJ/H7oRfrPm2a7GWtkVd2v5yXf4KhZPZwBE6zdnnr1dDmmo8Yg3w
wLrMVO61ddS5RCJfhNca7VkfZPqgCkqEkoNwk9fIQX0lAvc8m4Kbeb2EHJozJ2R/
k2gNYDYE2fCWBLkcFSN61+BAaR+YZfBXTxpGGytaZTdeULUxFGv0Dq+ot1A178BB
MY8QvNvc44UG+cArWHR5eM5vav2S0Uw7gw+4PcOOfbuEj6WU5q9gmm6zzqERGtQV
xQgjfj9wHWLyv7K321zbHoPxKWXvCAlU8lp/I5t6+8/bfKcrnrgyzsLDev/G7CXK
22K91mhLk0ZF9JeEzH+sKBIUnBcNeynS+W+7iZpIAMKOYrLnbC3R+3ZW4NkVd6v9
dq61bsXGwc3i/5aEJL46LXdGy9bmoAwFZDO+Dz1epeIdFjKq9yPUzKEBLsUtdib7
7BwgdzGh14REY7AJ2JT59OXTAqQZSeDdOc7lj7koz3Ufb/88maZQ2aMvpCa9XVwl
KLsd1iKEAZTGVUuDSOzez3yd28nYsD4oJV8jBIoM43hdSszeEKSn0DAPCoGCuGbS
DCZm8Owf20LgTy4O44/jfsIGfWfqjMSGMN2Hkv3c4sESevrRhYRAoTp2ltZBhD57
gZ5mYx4lUKXZrUst49GjwlHOih4ye7a1CNFWXSv3K9OOiUgG/G278gitJTUxa0SY
OfHO9sH5qMjERqUjcARnsresr4ZlvTaPU6JNLe9Fu6WgzpMsrTsJYfnjWuAOUDwj
PgskNv4UaLxKvGkGzESEN70xpGBzcM6rhJytQztb6pgjzE44f4CbVn1P+OXcUrp3
SvJoD4eZZZPDMDyk46ge3ys+B8nFtpiclyM8px383d/9yfPTx7Eh2WaK7djZHJ7G
16QAHJSEoFFJy3QuLYVmD/R9M72EyWqhZ6Cdr0cQRxQ3ROpNJji1q/8wJpanXBlf
HEX3fTdT8YAnbsoAl+A5UDYTmguXs/Mogok0Ic5OMGz2/rQi9tg6M46kYkI1wfKo
ewuiT2oUijbDTOWDt3t1D53Oz7+4ok8VhUXRJM9q/FbZZkFdtjnt1e+xcYe88dcC
2VN+FKRmR0ZmTn3J6zcP0ww+4XkTOrFbWAbkmh57mlTi1WCSwDGv2pxL7rJz/fOy
EmqkIm6FC/eC6UJskdU21FU5GK/Qn4LFDAW8SqahIADPGmEjUWFg3DpWWjB9PpwI
xPwYSAGHouv6mYsCEJoOES4m7exNoy3Ig3JbCKbYElN1OT6rNWjCeTy/BniotH+q
RS6NKgNSITCCzW4j6AstK0HCeoZvlmnOJEd5Z0VIXWvvxg3Hs8UUluXvPShfBzUv
DoFzoKe5WZ0VAEdRBi6j/X/71xGOr31TtttUWEftpRp1Fo4CZPBfVZ0VySb5RtDX
pYBkPV+51vqdUaW1zEz/MvQx0nDeteZ6H3JIDoQ7lf/0bI5UI1kVcRm7AQnugQx3
u70wh1R+38mcrnjlivBx+I3Ce+oyFHmho8r5icm+wCvqZxcAY/VwBeqD1e2YgJzO
F9K91Ayk7eEheu8UBFf8NRJQMC9+qlcZoAaZfYVQq83tkoeiUM2YjN8oZ/S60xy7
dWk+KnUTxk7lLceqh41KWxwRefvIMxE/02ZsLOmJzDGQwVjKwOV1sRudbVSGLZJI
CYrM5uX9pJ6KdFItW3o9eY0RB5cIyiDZ7BiRgy/qTwyWJmiBk4wGdrNZG/tlI3jQ
qkxMQgnwZklLQSdfKH5RR5aMXKbQySlC05jLTfl/Ec15SYcV/0LSlbi56AXiANSf
Rxaf1ay7zW0nbkas7jJDHmJI/aiMHWooiKBC55ItzbZeC7pjXFQH/Ec7bvtj6H/+
6NdihmnW337+XLzSh6Sbcea0BwBVScuvyp+SpJ0Zj7XZL1AqwIWlISzbpbWlone7
DAjdp0lN/ZFVXthsb7xXUOYTnUJASIwUmN4ycudhTrcbn3zzGat6EcesEU/A4aq0
k1d4HkRPWjQSQ4Dc89WiMxtI8MBEp0/fdf9TAXYsFVMnL3ujLUIQSJ6zKyWPSOaI
owhBAJn5+FYeVepqPQqPPSrD4NBF++GhEHbBCszVxC4PD02YES104do/Bi4mhx++
CBwoijRKAg7Kj0QRNoVRj5e5y6IziVfHoJpiiVv5ohSji5lnPmU700AEhyf5Q3wg
NwjAHAn5pkiuOBBuRQbo5XJ5Ysy94VprbOvfnjHzQbyw46ldzK7AJdVkpVVYdiee
xbFQRpaSXKU8JSClFr0dknjWw508Qgrc8ic+Q2pvfnG4Y38pR+weZ1SXRHl6HH+m
u1r7uxpwzMus0Cs6b1afCiv9sJzrZpC4vuZh7f6Qj6t6HEA9PFiUxU11LONebGRr
VOssAs6dCYAYzOft3MfTHMVy/ToDEpfunZnq8TCmUMahI5lBiuEPmRyRXZzpKBAL
ONN8FTt1G7J35yVUycvyGBl2VKjF3OVYxJNxYVZZUA1GL+E7l0jqNCA2BdcLDuB8
YU2m8EKg6hXQf6TRghgQyzaUbCLwPDzG1y3sm20cX/ee7hcuL1AxZ8g/jk0ZXphk
ISRgJO1CDin2Ci/VVnhnLcUCgk/qJDziRPOPR4w6G9kMT4UGhSL/bZxIQg79H9Rd
IIsoRQgtzK3Zm4y/62WChMPR1ykxrfg2ToOugLXBvk0KFR9MKJzar25UU39VEaVj
fd+F5KabB6w6H2U1odYj9GUDpO4rtiCNNiJRXtgGcpcHffJ21zZ2j4mPUgoeCtVF
8uaA8RrB++2qXe8OS4NsmqKovJxtu9pt0uB/jlewEP1frJQr1WNWFP9iS7WvIzXP
54kzk/jY+uKpX+iwiXqv122IXqNHD65TUs0/zSZntwX2bR5t7wPq8eGRMgrLNRl7
Xcrj25Wj6OjJZlne/bEhSEWvVhUezRYtpa1f9LttuJcY3DFyu8Timyfsp6TGJiGz
nKJ02hCm1VjiWmQzwjmWOIiq3No9XiQOWq81LLyZUeOR6g+T+mEVgnjd4xLse2B0
PvVAgfz7e72qadONFGgoG4uj2oqYImzTdwj1NpUi/TkW/43gV1j4u+hpBti1of5T
4DFHzA8Nf8ZwTQwRMz3ZiwxpNKZGCnFtI/y8XKvsvUrjnGf3pQcQP2hoShzoUdRA
4SJEwzTNDxATeIsjbf6UzXxG/BrqOqluRS5gL658gL3+YWns5hpxp/xFZmNqrJpb
DN26NfJowfaYfdWCgj+6yxYONKw3BKEvfxu0uOAAYv2gWf32dzVHSlbJESWtv8im
5/zR5utYohUAioecwN36pGKvnvO4snClJiOZ4y9VdGu9RYR6xoQl2JElbgxKCZGn
UnRHrJn5SqKwnYz8tNQUw7pGRtO2I74QP7m2FDCBzVyDhJQ3SlOO+ygk/bRLk8ns
X0q7Tyh1c0r/dsTdmCQh8qGEqr8GtSP+LQ8YpXK0xbl9/zJzKVw7K+diPr6X3oNI
3z0XJGgozYoFy9DzOKMItRWCTcg/sblS3rsKVGUqV/zDApB0rPQ61aNxDEjP46BP
T4pd6Ru2CMj2jaP8aK5DDSFVCXhueQy2Kfugn4/DXxfzwSqMOJYtYCZ3HZXHmoET
N2UkMRN54cnzXiQQZC46p52BTK8eLUHOLK3wYx70Z5Qabo/6I/JzeZn9tAkBMbx0
lHFfs/kSGCfjtvw/L3p3e1pfJLiTEDk5dUDM1umeTEwtA/oF/yyW1NBqJ6hf+GJI
VE9bvxX8Tga9KpDHICb9sujn/vQYAGAPijoR9qD1gjrRV4lWuUDVYwQTElRJ2mx5
JLJsqpt6onS6b/iwx0sA7de1jdAwhETth8M4d7ezKsYriaRF702+FywMr2lgRzKD
L3757wVHraRtsCiSIxUcr92na8yCAOvRmNr8qrm/LkdmvGY6uo3c69WqOiHvo/YF
nVYwHJwSbWXWsn6ho0/UNyC2JE+XIxqfCWkWzLxLbrmnUMgtqIgQCxBsfM/c7ENX
5VGMeOpLuIUyU2ENfGK6IstFIJi2lly7pPs1cqDwVfZYa1omTwSAlc+asSAql1ez
QNrEgnhqfpg1o4vCL4vPPkAVX51jsmQ4TnaKG1iw4CcZswTT9ptHStE3CsjQrMMM
ZBE1gUezeQRpfpfjz/vDD1nyV9PU6V/A91RgvoIh/GaWq754aLVQPhlsSPOvD4eM
GP1qCri8G8Z9j60UYtl4rwVAzzLFlVA4Dh0fApamUelEM9icSUORJON3at2lHBJt
IT2/WHqOKu0ctFrbkds4uFtdihztXsnlTg69Ev+CwPkcAwD6GtEmIS3dMAyrdY69
MjFfZja+w11mYdtSe7yDBYXgJpbjo1VxD1cLN+qyh9+xTQwLuWmDt9DLoRFKiKFV
bb8McuZKhti3EJMCytIoDLYoyIeh7QlZ1v9LtBzVX2zN7MtDtvcg0ca83O/UEC+O
t1C5y/+dN41HH05HOjHT6EWW43iuYmtyRoLz4TEGa4jTfyowPV95K4dLBwQMpp8+
G6KwCrVMwSj3nDoyiyRXSa0H6BKc5V8C5gIKx/qHTsGrzuKTAo0xQhrDapJOGwwP
tvBojE6K2z2EAK7iL5j7qxtsAm1uFy6CWedqEg8IR2QALZ+iasLdCGDShRKgxt5u
PztNuwCzpZ0bmol2V11KXiJqasfH8Uy400/F8e9kgbWlY3nYp+sCbwR1yM8IIpXK
8mAWmD2f+M+F4Po8XkfvmDW8E1X3rVwyvrHRpc/u7o8Rc5gUnWzKWRlKNmbFhhUw
Aufu0o9URJdfQMDAtdWW/GWo5KgKLtVFq9JpT5ovPpL76LNTXqHyUTCSnbZ+HJxV
Rg8tNoc1YBNu8pFcIiKoxwb8ONiN5pvESbn0AjnBdSgFvTQA4HEk5vNqtkBMnkdi
GfWEQu0qf7HyGXk/s6KNezmySFaWEd++ER66SwoxhXShX9tiBDr7ImSvU7uvtbAO
lwOHBOOOGci19nZVDZQqGXowLsvuEXdfC+9xf6jdUtfX3+vgu69hGa59Q7EenZL3
hNYtutBeeIgO5DmM5sLtGpfyrS8/G0TxQeoZZmSot8H1kqOu32Lk4qkhnjLtRaWI
pAr6N8znzZs4ARx44BcIW8EkrHsgLl5gh1QIpn13gxumECy+SSliUpZv0lccU8xe
ZxhuxslnM4nW9thzDmXfxhaMqljQZwf7Xw+CG85E+rEdAmFiw03MQESmq6OjI57k
8pl+6QdjhBtg5fVM9xw8fKACmyC6h1tSDEipeBvNT+Wt2YIHNJw0w9XlpCg2jv5n
T+QMPDmnL/6th8oJNEDN0l/M7/1dKva+GE70UhvbNQQCUAvYXe4ow20FTAnbqG1a
GMtpFpy186w7dljboyjc7jSV0gbW5M6ISxaXpr5nbu9w+waFy/cqjQnEstWuwNaq
eYSi9az3vGMAP++6ko3OS/tB00T7pV+ZjexxLsAusUwzd9cHzLIlbzn9f47r5Cpg
wiUBfh18ebWnpuQRBeLT0/sg/WLMFX2R/rJXBJsouZffGNZjG1N0wfQk3y+/w/wo
M/lgJPF4Vdft1xrQ/npHomjbqb/UKMZQkWaR1VqZ14vsXFZSTdw4L4fHITcvGsku
O3twfCwj8AJXRKCSioVOmGAMhIoRf/CTDHZQxynXm6AS064v9pxy0QLh7jpTffnf
JKCJjXI8TQBXJ7k5/15xQwSUgU+FdRpKE2OlYqR0oL5N1sI6zL39HhkktjfSoc6U
6v6p53gxD5s2eo+Yq5FdRlRgE3x0d4jZbuYtTdZgrU9gpcbwtcHow3KhiJfBy7wE
nQyL6n8k2H2lEDfhkg6ryw/MwolViBxLoEUPt1kJrn5Lm40C2pUcxZIBdMky3J9X
e6QVu4hxD0Mbmfl23Japzu6nM8B+XLNa16pRBID119fxykAtvIR9QPYVK8CZaH3r
IlcM6vIiD5Mko905vjP/0uKnTHmjl3BaiDzH+kwrU22JEfD6d370BL1JllVLPvpB
izR7Z1Gwgpm5Z/ftB/26ikrP+8KDx8ngjuIn83fKkL7puu1JsTP0q2rtD4OUpqUM
m8Vq0yU07VNprITAEt3LCqnKjvXTqLGtKDau60KQzPG2JqsaFw6EfK1yczW+qUQY
BncIomEpuTk357dv1Am9gUMnvLbvy5106CXYCioyuZkX2jtvTU9oMGKprggOixOg
5KNR8gdEH1zppnM9STK/EB4mQ+pC9NsLJaxhT7RrrmyxpYyYnKfZnI/FceqiKvU6
QTIJYxTnUMAsCgtn28PhObKO0Bo2U5uKR8AaccP28QmkgE/blIWs8hX8167YlrTh
2NEWjJaWpITIPmbStuto9YGvGD2mt3fxnOTD1311mqVl3gvEHtAFOFzwPRZnU43z
YmXlCvva0DOu78TYYu0uBYVZMD0lklg+GNnRJzXGA0aJ3ZU31cZRNSBCcRYMRiGj
ztk5dKfZysjptdzT8WG1Es/J5fiq5EOeSlLU2ecnKNmm1AVY3hN9HXwL7RX2hkhG
QDKKr8HrrozvpQkKJ8EJpJPIvi3gjFTPbiFqHvBekqNG2TTVv4EfX6Dsb0UPQsQZ
fEp9lKasopPZbewqt/SScSQ3Avf7m/QQPGGVtbYYhqweaHMVRK/SLPvY5yzy7Up0
2XBKouTC9W4CYLjGPbQFsYmN+Z1YT6ocGMWkT1flfdcBI2KG1/VHQdpIK6EVVPzt
ATpNVI6AviZu7d2BC8OPPqRfkLZiT5tOZOchkKFiZ5XPp0XHARe+n0hsHBcpMCWm
SHGg3ghkZN0l3usIbk6EoSvs9q8sL8F4jNBXISdd768p+XoMGuI2PJsp2vgL+WD3
Lc2lZ8/JtJyTxDz0mDITR9ZdnFVUspmq2X959v8c+R3yL8k4PypiHjewj03sseo+
tAuiHLzWDkAOMG71L+Pe7UdnmbVgU+qmDHMm3juB036mpb/oKoAAF7wKxOwNp0Q7
4ZBPVA0UrfnHou8eazFdO94C4gq8nBbldNdE1yQm5HKEdZJCFh/X14VCAKgiikQ5
o+5dM3d1XjjraSlp7UewCa+foG3qltsrxegWugVNTZQ0t8AzESXffyYXe8TB+/5B
mzIcEmHqy8nayjAm4r/AObJ5uv6tG8FF2AMa8gZzgNRfb3t/aGqjk+SJXI3HQrja
4kNsIIpv5fmrWhRFUKHmuC8x5MIvH8pSxXIoMTRNwC1dllaH/XC5UUIvwydHXJS1
7LwtNXCM6BETdZceXnlQo9mKf3/LgiAnSj8sNpkGam76df4FwUuWCjo+3y9nmQ/n
x1J3eTELyMAxAY/kTz6aFNezakNBivmfaj542V9Z/bdUtFhHALy1qsPEUQkMOQ1a
2eoJ4T1VS3HXxch2alYoCrakLZ3TN1cWywm88eC3Mrd6d5LVL37ReuxbBLWOMO49
pFMsh61L1e5UoQoi9Yg7tTotDL7POPrDN/3fvR+QpWRvPEpW5vd5KAU499PLAFow
6NWtHcYjPVboGilYVu1+mAcZlYygRgT9EMjjdFhFGc43dcp3ZOmAA05Up43hsHx5
LWd0bnJ0Qd3IDotUktqY+48J+ri30XKseekt9LmfN3gnmE+PrzMkfYHGdnzlBHdZ
Tbp2d+MacmvY1iEIFId3d9NIVAqI4GaMbDQOk/FvLdyGB9inDWSMRTyS918vfZpV
c8DVS4p6ZQt4bO8R1wVkwLmpgTPu24dMffvfhqovQ1XiD3Xq4vbsOfTDaFd/ucnE
o1lghRDdQ856KJalHZyYxYMPxomV61ZBpZ4ZcVNA2soHhNIpOWxJPn398Zki4cWK
+4t5XE/HaJYdIU6uQmDdxom94NFBKDchueXludU0y+/3q+sFXWLSQyOMXgM96q4+
B2GDdoQsksCCHh6m7bFSyDEipGsfgryVreDyL1ti1RSuWFbY5T/39wy/iFHQUaoW
4RaxGcVRT1z7pfK15WxKCAQOqgRG1oZMwUn7kpmj2VqQc4KFSg6WkVMRbp7l/NTU
j9vx1eeTtOwRBkbvJr6imLrjTnrewu7m6woJyoTUgXelSz9i3CcTe1XEzbb6LDgB
4UvKvbSN0N3GU1isMBO47JjLORw+ViE+RPWGdkwZBXuWlSKNZNe42g80SBSBKaHX
khS2WM2YqyPmT/tg6l8iMOQnVeR+R/Fvc5f0yi/qwXGw9yk/+qP0UpgOPr1Sy0nK
YTahHzIV9lcUBytmqMh9aFAZ1C+soEG6AToOk+oDxdlOWl8eUXHqxgcjh+DOq6Ii
wNUfur0gyCBw1uqrB34pX2S9BFceCWwIBKPTLI+DUPhpsE1yQ8QOQEOGSZQszAHJ
NAy1EsWKwa77famcHS123NSQ4MmGKNx9bRKUO14EmmdJ07ySP3XNGXoIASk1cko6
KqIBkO3HxtvcjzlLpAbX26sm+3cgD21YtQ0WKR6BUf4xY5l/thKkUSZKu2+Ov/g0
nQLFgxK+SLv4HiPgCiMQU7IOHZs9GqFROsEyu515Anu7uUXN45h6S7W8gTdk1Jhr
SiwrrxfgFknoe3wBK+vTiVcm220IzMrtA9wGcVERdTOyeUnvPrHbOG1cdPZKFYEn
UL9wkY6EF7egOyH9o25+e9MzqK9APNl25sc4LsozNejeqK8Hhksak4+THcbpEveO
Lj/s1zY0lVdH1ZSGNpobYbQGY7dN+ZIdsEu0oD9gutiwtn1+oVsr1qnyhVQjA0KX
LiSpek2FqORbV9b2299OySxUGKEgkjLzDxaDw6oi8T+VHJDo0Ura5heMtoeGdy6w
4SlqwE4KAQ6XtGPKQAUiPDLsnadKWe7doUURhPzdTO8b6Tr3hd4oanOpBIJPYYny
RSLZCnrkAHjrjR2JXF9sQb2MeY6YF1z0qBl8moa3Vp4z2dQmKIZalm7HiRU+TCUB
e/KgKrXhljsEmCm7ZS2dkHHULISCBw7u/lzlWtUsKMt4yO5U/5fGAnNh5VAqoC5k
321xYECJa4iiESiB+OtjQXs/rOtUp4fpYKYAViaTO0JHfRwKy5TXrpmMhxBJvfbt
o6d5XIlBb8/vhkKjrnPJVqRL+8wPUG14WdZ8WL4L7jh3ZRBaTuhAQXT2r8ip0H1c
vPLe9PRZD0lwrF2bhye1uXXK8eFbh4VZlj/Ax/b1wnOTVO/hUzgCRw967UGQSJIi
u4hiZ3ARxgUzTVRm05qW5uMNtGhB3RC/jotytSZzvswypZAeO4ld20zpn88Y8DnV
9G3fvucEzoscQhBWn2vVe2zJsApCb+w2qd6L7krRHFuFg6itzUES1Ly0lfTL9ccT
hNwFn+o8KZFAwaXg49QGFAEOdMBWovDbedudKrsIkbdNvhEhd7GyakbMV9FJPVw8
TKd15skvEnJdDU6uVcbFO2w9gN81Byra3K3tP7geiOW4G8wLxGVbVZJAs5sb2hNT
eaVFY3O7Pv1LgnJey1J0iYQJHEfbWKlnjwj0ajUmxivLcc0SDXUQuRjARvpw9Qgx
+cjipYh13/zs510j3vqJaXQ+wrGIxGmu6xW2LwBITvL2HLPXczImcgW+zFNRH+RK
YKEhuAO7TXfZGteUJFao9Rr8RghBnRQdfUzHAsFK0muinJifISbvxvRbYa3kXJKw
tO7Fu6tuLRkoqWA78dmLZG18HsjoKPH43aEBMF0t/QHcCDcomsWAWMU6tRd/YcEy
NfR1wtckU1oOzhUoCSFCCvYEot0JjO/l8BYr/UaANDfPgk3AW539K6TnaLYW/cpS
ek5wJTUuJoSaZGcN48EHqTnBv1l8aOWmNlZyod3rDecauRC4tXNW1ntrnHjjLjA6
l1uiu+R7RFT8u7g6QeenRxYxGMKJ5is0tJ4N6aSRnEhALW1n6QpqcYAr2eXR6RvZ
R3KtcuON9XgQNEWus0ut7rTdCgdDGc/uhNeDZUflo+ICR5L1ckPPLPwG0ioKp2fi
Ns2/YWSZ1pPsXYjcT3eS2hM7I3M1zwW7nBPNvOiolVXbZSGU9iIsDuhob2XJo18X
2LFzvsNySqlLkGCmXICPQfnejHt+vh3T7UL07PzYG5c/IXvjcIF0ltqLoKudS4TI
Bx7pyvkCp9bJjsIjCDtfy+hyQsxYCMEz8+bU+uvd+YaFZCHWYD24ihq3G0uW7LKJ
E8s0O5yVbq38RgkYbJu4pbBMbuyDOhWOfZvkGGxhUgjsZkGI864aInYRJ5vSxNZC
gRXZT/NyM+IvlaIrxhcIVmgQLCMuk+/VbHu2XuGOEopd5SsMo5rRcY64LvIYdSWN
mJPl1zWXAxeoIkVkoXjrXd2iG1yAzY9lSWoW+4gw+HBlvYGYpEzkKbOOrpUIu/ZL
UHEs3c+7C8ZGptrwp3imwZzfa5D7POK1IWSkyl4TwEDuiuo/UmNbJF2fslO12ti+
M+Z5co0EB4R9YgT1cbeluHM4Si32296Pz9PvMCGu2TgA5d2ofJfy/Bv18rEiYu+w
wTfx8HYhu8KjYEI3YMzKV7a1qqSpeZK5VhWb9ezSn5C44YAQbabYjV4Wi4MuEUPZ
y09E2hMVmsiXE3XSPiJfsGqXbdmQQDWUMx258M8SnvtjJ7BaBa/pjvjUJyWhN5Bz
AK5qjKk2FVggS+sh3+cRzvFb2ze/0EBNI5HFD/adIWgd3FP+l8QmH35J/YgU3njQ
WPcEPARorE5oSty+IawYj4dwqAYFqLNadRpvqdeAM2tpAw1rb7pHYUw0C2TP8/eF
W5LwWtzkTWLzSl0MAmplv/ZSeFiqEvTmTmruMQoKewyXWbQXWovJeZZotXohdOPl
/Rom/52y9qXuMCopD0kLO6Qi+pOeB5bQsIE8vZXNL00nMPX+p6txBybKGRadL4Vj
DkOIYrfsHSj60nElUGMNtMVq9EJroubCri1wvn6VTYx8qsppq6ubQiYYhvoJqzUH
CjGbmIMgSQX2+hY+iZNwHBvEvX4k+kFm4WqUEZla8IE6M0DV+Nm5K/yD2tFFt3ux
nrGeTqdLCqzEMSFnNW1fakwbq7sloxFvMvfvzDf5bQQ/CGaflf53tNT3GUadOPJt
IuJcfXYWswKIK66B8AcNUEpBF+pxOO7PrmNRiXwnFEH66SgvtjR+0bHVbSin9LQO
MBFiOhAmXHqgF9D1GiKAXLys7XV442T3xornyoy08CUpsomEG0BzE8MkOjTKoQ5U
56JMziV0dBx5zPirPYr0rS5Nd6lo/lzv1WRPBA1aHTKCUqb3fGolM7VSY1F6iqWJ
dRIV+M8zqJVPs5/bieQlMvcSy1ONmbaEUVg2+VhvAcYLM6L0ZnBO7Y/lo45LGcZT
ZXbcmdKQlTdBMQlwnbmVAar2Gq7oRXzU9KdhgEnCmQTqGqk9/NFcKJlbbFWlMrro
TXcfuJs1uSfRaJ5npOjLVN5T606y8aS+EEkfPk43Ev1dHvAQgSHJYlDcCXqjl3Kn
K0Okh39zXDVNnxHq7Q1V8vUYGuePIrYXBFDV4nssBJHzViBRtwMic1Zck1V3EAIM
LYKC7Yjfr8r/JTHpeWCCl0dTmd2VJW7dkGQdytUhp2txttSKK+ICxZj9yJnOA5uV
y8FzZXuDngjzIkkyLxVniYfnPL4N/YS8ZXTA3Z+bBzk5PrNxPzvebPM6M52hdHQ0
h8TEQ2G/Y6yI+ysP8cX0EH0BcwVwUyCWHY6noOuwW9TuxXeLtgE2d0bsW4prcTFN
ncos95rtBolMZLZBkdsZ3wvvigcKU37BDUY9wDuxdDtI+ivYl2kHgQfv7fgZkxe6
b04PjizE2933/1PYL1sShOy5kUVDo0IztoGyvTAFRxsvuRX+FFbGCyXVUUUHmWpL
/12dj6EsrCoQioaH/9XGNDCdwp7Mzaw22m3vjx3a+PNM9z+HhrAuke6Kk8E3YgM0
BLzrPr335hsNRrUQkylhS7DPcfy87krEwI8V60u4R1qiF1XDHvulk1wJlEhwd/QV
J22wzipPe/XbMT5zj8XZHzS3lYtc0u67uJg8PnkrgG9xINbXxF1L8NVSo+eA1YbU
HtSVUXmphntx+5WKt1D15iyVUxPMAK2r5wNVDVhCRsdTBH8Ji36g4RFNLH2+sms+
iEXelVIfBvjyDJkx0+WxxGvel3ulC8Mm2GfKz6xq8e5xKYKAgR1eTyv4E5xtQ/1V
xy8G7ew8FoMNRYSUFRUzJ/BgE8KspvXUuVUyUfXZWwy1ZPvZL8/5EchxTsd/vaMo
FxHXEalHGjmpalpBrs79Nck04Sl8BnBo2RcQxjZ/FB6qMoNynCbZwmBekzVicXbN
nMDucHu7Oo9xEOyuL2tecBDO4348InEgDjVNPj9ENeTAhPyVp6c0wl5X/Zh1X0+M
o9C2/t4R5UMsHunJ6XaxkaDFEtHIeN2jINVnXMcomnkn4fevCEZOF7jnjCstvNH9
p5DaJfA84HOH43MYkkOyORLHVMOMvuUE4Z/dU5/oxvQjG4UiBBrJiWlaeOwNBsN0
qQeT6SWt/JqQgCvi60fPJgrN3QL0aUvhXnrcMcz8cnUwEdf6UWWF8BExzBSJCx2I
Wl0wc5zoxnToTdwc9tpL4kKq1tJ71sJpJEsQObdc7b4hcyiFTnhE8A2SO43vn+Js
ipU+awqDHDzg8wiH0wU6xo9abjrSrADMu2lQb1hFvnryO5xOsADkqgxKnSdvbNRq
hbpFwn27pNBVNiK/BSwPgbG+cFvakGRvaBdNEP7ISPhtArb3j6SKbQYLRn+STN7z
Vq3GKGraVNbW+T8zbUh6gWKBawX3XOa3JUgZpSpVW9IHQWpPKGFmTPYOh+hT+jSJ
vsw8WEGfi4xeaHU1Lm2VaOSJoviGm1sKVVzSjnLvCbe1DS48xnGxbCbBxeT5O17d
t43DaQL6J4W038K8+pYJWDP3fwuHexT/9+VbUzf3ezgJeiPIxcEy6h0wQzlG43bP
BVWXpa61ozKbuDnCpiyLlqfQMoHVYZnuGNXMOcmX3Q60aSngTjQi5JhF/tK+oISx
Ce68HpBIUtCRyDfOZBtHN1oKAHfZdfFGK2ledDOBOyQeC+c9fw818SRiB44XeZKH
XNmjcFck2tOfGmGOpT4qSzXOY4zbBhglxSNODjR2gle4ZIiVuxj0FJjCAdrGkQoC
ATqYQOvtmS/PV/MCHeTqP4Lhfs4YFDVFoteDIdR5TYCMuRowe47mecIuM0pO73bb
x1tLowtuXeWlq+stLa5xCmM1vvlD5/qUn+eYKIj5wiJtvTfqc0ZEjkqZ1eo+Gxom
TA+Kay8lbM6rxIUPD9vSli+XNIljvXQL2sUnrNv++7He0Er2cQdKYSJVttuLMQGc
sc2SEQacHdQRASwS7EqnZDs6pI4B6LDjkjpZ85ornYz78N/uoLzMx6R1mjkW0rRy
t+N68czkmkJM2HHxzkFuM82KYMIih4Ccemo4pfZErbe6ovGbMtQDdZZWJcgqL3tB
fNZyhrFNJXWEcD5Ac8ILMrS98A7faMxcMqd6oNEHqdbtvN8vAqWCzxXzPeJos/qI
DDWo8fxZGLzQAvEU4to8VvLSnNNWHEwcwIZLFU5DnkMHie8TGeESM6rjXVySaShJ
Q1+Xu3zc/ZydlH0jzz/5q4seRNN14ReTk5v9O0L0EkKrqqOeqQlGKShZ3fri02VK
5BFYvhMgWNgyiXwhe+7WLmzc3UDhlPRA+Q5ZotFGbA6TJbxBv5iwV8AsIBDPD/jj
IAqgAnh/F4yrsND4KckeNEZDmwRkFw9H3Q2Xwp/r0oajJ8rY1knp7yg2lKB4ECtr
s/tOL4FaG17c3ijqM6q0S1aKw8W/ShXzwQ4A6DubOuzk5YixouSPppI1/xpE9tdI
cEdlSw5ycS4fJkmWYFRgnF0N8YaMfBE82rZI4C2bbQq8qPmQYek36DI7LtwLEBMb
TW4oVLgAP+OTtOr+r+nUbKtZgyCND5NxKQNl/sqqu7nHuUfdFZFbgtONAb2XLjpz
FUmvekbHVhuobRO7HLcTgybKWpWFo+e5LW8odrtHOTZdwDMMELW979IUlGelpY7w
BzKmNpZaW+qt0lWK9KoroRDp9HUZSnRBaVJHgbIu7Szp1IXS9DR7+w5QB+wxug7O
x//8ChZfZAZ1sViVSjdNHWAjJAQQYQCqmZYjX9XEtN3Nws50V60cYUwlZ6i6U/01
SHmPUa5wFQ87uKSrg7QydPzUvmWrICqJhDvh6nFAuSj67c/XrvOzuA7XkQeWu/TR
R2Q7Yzchh8bLDRlHdw7iWth89PkPm7armVfjWKnD4+9rUWveQZb060p9VujD36O+
bBJ+bJyHh1jpkuw0EHPRkCG7BN2vKGcOsqpzpwQSuz1UWtjNT599RjHNL9+sxdmz
euX9KZz0IvmytSrB8YjmdM3KMurzI1cLAWlKX5ruPqK4OvkkHw45exmWppaQeNB6
2VtSahksrSd6ljxwRfrI330HoWoj0/WrPuH/FNbE+9SHkQgrcZmdKmy/MeGQubBN
Ru0yPHDCqJcb/evs1xbITPttV8y47m6b/92nzl1xlK1guZMFC1YJuE0msm7Bs2Z3
y85w4EqE5l5esN+qQt2JJAdFnxBvA8JPnoUnNUCwisuHjn1dnpAznifCh+IYsEgp
Tv489SYPJKBjm32FijcOGmLL7LdLOveGgd1dx7dUmcKXdQt3021n4YROh5IkZbOt
H4jYnAVdq/c4R+GaQo12qy1u9K2aKQEMol1L9FPyvwRq9Y1s5P+hwJ/JIxWSeirS
sUsfMEIHxsrRorCgGM5duUh+JoKH045nLK2dgRzS1yD799xFJX6mafRfIAcXnGHk
6m+V0xj32OIk1ZVzs+kkZndnSXIZCAT+Nn3i2Y2br/PNQF6HcESLl/ZExinsT8wX
HILQG00xPX6RrVSsQ9Z4HZyj2EbUdK7XV0w0CWzcpSQVIuhuxxKkPLN4zeWwj4Fr
9+1/7r41PfjcVFPTWfM+To+X01lKQFOnPyUOL0oM0G7e+KwUrNhsuVWE0o3FgySm
9Y7ZwwY6CxyzK7Y97dK0Es7p9Y65K52u/ReLTtyuj7txEnB1KMEZmMXr8gxnTirp
CCIMAwwl4+kKSUy9BpI4t9UmyClhIiRfIismc9IGvxaD8nV1aeYyqfKLVf4euQBc
pNn4jpl6fbE73xjtY5Xd7SgL6YX72VakL0sD/IdL9HRm2fRm2bslWHxQGW4W2TUC
vBUR/vXFH9xLllB/WqkuGLDeMN+5ETDYEJcxUXK9eHRkaT83y2HbLFCYMNyicHAd
aHsREigd9iKiITU/MkZo/9bo96gnZ7Qo1Yvv/KK7ISSdEcvcC/KIz7stfV7wDofy
JHoGMMCj8jumDV0hupyNubIjk88XR4Trf5MNN3X4JRS9J/I7RcnJww8bn78DWP/N
qsFPelLQ0m28SVFSHAO9kGprcULcguBp37MAs6T2sBGMoFWHWqTFFW+pVLnvUXOp
fEaCA8qfEsAlQbvUV4dfmRRnCNWSI/Xy4b1b5uNTHbtCuIWS72xVhqaApxkjyCX6
AcaGPlLbV5YwywcvQ3uoeyE+dI6O2hjGWWIJclCGNDueMVIi+Z+tpHnruku8fj/M
Z6jl0bsbipS3PQGolijAOfpJRUhXYeS+2JUBSp0NR20o7YGddksR9Iun2CCoa48o
KWq4nEhJ2ddPwN6IL4oWVb9/J829tyl4caU0mVmL31fRI8lIQf6ZAJwUZvHsZpCO
LXXPtfftnRf1t/Seg/oYdvMc2Q566UaLfJOpJpz+Nhf/P532nyEXxiVF/WXEb+Hx
a+7TrceEulFyfYFOsHruXWArCrGp6mt7xKkIn8+icUvPLxebSKnuBMbt6IV3yC23
Uo4m+/aDLneDqeS55/DfJSjRowAd6rrP74ssoDfY+FirwBPOygOjeHhPu1T90ng9
vi2vyRFfOqVF+jWUpKMICno3oy8Yj2mRSldmu8f+j5NHtyD1Ep/ZISQw2jDxnvOD
Xws7w6JePvuRqmd6Poih2boJg1WN2fHLFRXPmz27BcYjQdfnvZvfp/6PyipcbiNw
ZWsNjrNsawD6HK4axZJ2gGbCk9YLinq3n5uhrCkpVjAUU+5cEGW4P21rgs4Nw33k
xJJ1p6weT1sRhAVRJ03WCe69m2TNO/IN/xgKVsXn0KouigBpYG9d8OVOikcWZJ58
+L9NScmxsIPM9vfNpQZub3969KrsLRHctEEESio4sfXvDpOqhFykt2wyklmJH0bJ
sbxvrbUnj/KPIWtNlaOcBkFAKPmWETK1I3ifhWIMA+1h0EyWyyte8n3AtkPvfJ3E
u4xz2CM2bnHm1kir12vdUJEgxKnq1kDcHMoZLmqZdvMuzTvgc7Pio/9bjx95PdIu
RIB+TUGMPH8cxVuGFSW0KLkTINa2SY6uKFqz8ExaMXZ8G49CcjSsbJg1CbPWCgDi
0GxTKq22ET5O/8NhNGz10wxtG+NaxADSXoZ8t2FZVlYZvm25GQtNGvXqeYW1UiHE
SVvRyARk1uwwMk3WWycA1gtac5/h0XQOu3UEPo10RosZTQQ7im35dtQUThL38NDf
poHBWxU2c0jjP6a3QH/xNnvr3T3uOEzREpNK5XFRjpiCID45D4A4SJ51HZ3SeLBD
/NBWtay2JEAYwE5sO5HMCpucuV0b8/587lpI7HC65whN4Zbi0QCgXtuxtJY8sFlf
UPWaLYa3UEFevs8Yjdy3FM4QB6YoJSqwur+iXc1KYE7OF1iSBRdOMhYAe8RxSDqZ
M3bfWzFUd0lezGDaKCJf9YhED0m5ge3j6HZ82egxqMRyb6kq2HlmPrldfbsO/icP
zNaztTLaiUEzPc4ImwfGJSAw07iHjLZedkjmEHxFchmp9V5+KgIWTprKChuFKyi7
rN0QvTQu+yUMdXPbxCCSnUjY/Yg/yJ7a9eULDYzlGFeInTd6LDJKGfSMcsTpjb4f
zsMhgX8SCGmg8FpIz3ObA/nUxplCcH8j0KU/0VDlvKW4ISnnMuZoLXD+NJFyx7b3
9YQp138NDV4dyYNKLFB1fFA2GlPxBENjGvuZCbIodcfh9XkEPYYj/UTNKiLOfJxE
ev9mhADktTGQZokOvpcgKpy1yOHZdT2cD5qe7sbXTEBozQCM+iYVyuQNnJVeQ/CY
r0UBRoK/ARrP/bUnayulMEPEoUTyqUZ+5DE16syskO6NQoBQMe4KKZm3i2el96r7
xeNbG4qA01/Sx5zJygQDcX5Eo7U/PApz7heyignBT0p3FpZ/2qzzDsCBPy+yHCUn
sFw8a8N31O+akDlhFCd4VaOeIFGD3fxLI60Fq1wJpgc3Ncu7AfrgBY5C7J0bd9FP
PjaDet6FmdpOGfEriDnQmTMXmNLLKuH76mhbmHbKEgwO6YUpFhO0T3DhtCGHya69
CV923+75du5zjxXFWpEzA2o0z4H4GYQda/HEOxEjdrLRXVBsEFMkLY0SVssge6QI
x4jr1Q8jIpZhhT+8FHJuvkbzhOiZ/q3Ofu21B9bNkm5cL3vKH/nHqNMBdeF6evQk
6ztneTlpIlss3jVtzpxvpcmf9Cr+6vSi8z9slYQcoklqOp2EOpetaVxx0PSOPPVI
mCgXAdZvPiIxhgPqmlptzUxdz8tFVdyOei5MjuotvhomtTzYDKWK6Ur7I1ymKhAg
y6smZ2kAXI2VER13ih4PM4owe09QgC9fTaav3UxhYwgeJual+Lugk4y+qWn137UE
E++WPIDJZuD7+NDG72QTsC7mUwTDHTn+Ydq2GD6K1zt2ZwVU6RJazqPsUrAavWsd
PYwbTG6S3IUqrrstfomJkMzHCnpcQHX9YXTxVP2neg4GkLPM1jo26ffoxsGab8fB
Xys79mfvSLOvtUFBSF58+NhwhgyxtkGn9PLajgL+reYAq20UiRyIFGD0iB4T3ref
LUoAVWKU0j3nmgddfiEVPc7PADm7S+BkbMrVxgnMhcE+EqeTC8gl/hRDqLEQTF2A
NTzcVZgNZjoE5AAxKGZK0YxhSR4YpNDyZH0FrYrmEThgpWl34+U9VV6Jt5VdG48d
N6rVhiMY0CpN1dr2NyJ9TF3K6I8z6XLf+nEPrRKBYy9XP0LF6fzhMKcrkyt7M5BQ
vEZ+PTE5Tg1vzyDGCeyj6jJpTf52IuiDmWqtxjtVP1awPWcEBsvhk0TYF9Xm5EUa
/mXXruRldDxOw/bQK43mZcQp8yJ7euyN2eYfIhUexfqycMFFAuhWiV5/cUkUQp0D
1RzIKQea/BsFIYaVl0YxB2D2uzmV4XzGDAQHTYkgY2+JvbcAG1epSdrl+mDBEgUD
LGADuT/9TWgnmUZUqVhgPDuLLy/XU9uNfDgH6VnvGs6r0ehm322CHnFqBEHb38S4
rCbeVp4XnzZ4z4DfRJIVkLgRjc/O/0yO60MLVfx1hATXFR8Djv339WzG6wWcUxTc
Ox1isbARbDliX/AC+Isc8uwwuajZIjPLrwPfndeeEaUEUOlJq8UXyW3dP9axu48G
Tx1jF7Jqplom/Z/Roa2ozBPcaoULm0muPqAFeL4IzDhlimLPAM9DatcqMuAS2ahO
5A/dMSgIiN1jhholt8JCq4X6aPPb7Nbj0VOZWI/MQLsa7sxrVyDEuephSsALOIav
BYUkOywgiXFC3l2oZ+NLgcWMMkmTrajAi1KkFUvNr2na30BzckRTgGGUwdF7ftEm
/xUhtdTYilg+OAbL1bTpNMa/WZsqO+AvBlLmxRU/b66fZ03hW72c4HbsEbooFIYh
fURYUThHgkoNwPmILzI3xa/RE9ZK67CE0xWsuP7SENOIHcn0c4vEPyUapfvIcEjb
32z+tKLjd9bNR47/SFY6P/L8MtcD3h8G5fyyTdSQGXUq/6rFp+kN+XuG1dcJ8I5I
bXbeq4uJhz6lR63azgQCuY/eu3jNv4ofyILxMWUUf/ZW2mkyWqbWAvwZ3DcN2Juk
EXzt8F0DaTSNCPQdfztUmI7QnsL5W9N5mK3DzDQ69Mp9ryt0ZLVPXdSVJE07EyI4
zz+euioC347Z0qKTxPjit8e6L8gphFzlq/qIWcGFHAS5JPQleTEfmgB0ivbepFtQ
sY+IyEpypxK89P8cWmW9jDgm/rnCOaKb3AxKSe2RwhFVPfFnr8afrezrsTHDB/FE
hHP1HX3kehFu4+vm0LS00ADS9NziAWkGOCR9VoKH5DiRex+DUqQbRVTRG8oxSvSi
0KTLzEydiWiUT8QJAH7jt7Fju4NAecSS/bHTqj4XP8c3DcVIEp6shunptbgjjA9Y
TJ+694koRc1K6WrABV/dCqVP7GMpS4rV5u62bzQnSPW9qUvTI9w4wK+gCa1kOp9L
S5MAbQegbkaJoFcjqVYeWyK7fLYNRAKF5j9w6pUdaUf23cpXy0YyLmwYCZdeJXTi
xZdC4eWZXmn22pGi91m1UsCV7nxR/S8/I/HJJyZRkKahU0ePi7SuITGMerpFXA0B
HuHYN3mADwoe9nAQBJy/Wi8+NQ5M0HTthY28hC2Hza8pFLtufhtl12s4LrQfL78O
kQMy/7DB5b4MxkKlMzRMDoPoaLa7iUJ10qhB5r9aY5NzZYs4qgNC7s7xH5a/MRR1
xbuJenE7mjQ3nHp/vTUXhXtydaZA/ruoLPrlGTk6urVN+kgVQBh89OMPUGmUHOul
BkoXhNktNWcSmyycZaYTuQOUgTK0tPk8q0dImCETIMOKIgVVk0OjoQD2NLPgPtm6
TK9JK8qtqBN0gkik0+EQBXBs+8hx9631mOy+KZDQOdsP6OaaEYc9y1VNDFtsHF/X
ztjzmbFdJnrmE5Zjrh8JVnA4vdE+8732KttVl7KJNmJxaX8dctwV2ZyG04OmjsTj
4h2M25EX1dEjCQfh9SUNLkWPCkMDrbgUkrguNBrikHqrF27xZ2gzdz/nUYYzjell
x9jfRGGhe4o+Q54n4AOqtEIONYv7oRM7OD3QjzI90aryNJE07wcLNBUxc7J6MNhy
2jt3y1PmY6xbkUUyIiaMg60jccoD35Vfdr8w5jBrkWDGE7isldcbY0r9tI8R9/8S
7BMZtDNcShGD03MTlDgWKwm4gJ5vU5H1bj22YSrv/CxGz97y4+aBYk920fckp8cw
n4qf5uzB70c/rvXqViavscI1wbqFb1tOipBxdfXtANT2KX4Xyk+T4xRB1rdFP37n
07ihAlEatMrkrj/duhymsb8dJpnqtx5X+/XReRmAvnV7vfwaFRKtLpbFSxAnFQ37
29N37TLTvWmCnJtF0uuHvFP2wEgqV8lKTScdMbZKzCm7uEK3kPMXP0SPghV2dh+m
PxYAcMk7g/ptgd/r0zSRuWWN4MpalcjHb4BwuaJqSWFmVvZMRwz71FDGtV6awYHb
4g0NYWTMbA+tSKoPGMbH9MQlaav9U2/54UnWBtUWxPcz6DzPlmCoLym03teShz8E
7idbL+T5fBRfSpIR29BvibQ6yBSalQ9RS7huUUASNmmZ5X83GQGeTDUWS3CyBRP0
kJM4et07t4/2aW+dxCLO/yzrmbN21eju6W0iW1X/vNkTV3U87tyLL0fwR0fVeP4b
merWicovgZa1N4YF+JqOX24sdZDswNUE+Ho7W5J8S3OKXgdWRBvcrq8o9AlKsrag
ZF835w+BegJqAwJUrgYy5Ff+B8DYb5xQJP1XukHX8krZxM8TAXNoV2We3N61s6r9
vWRhPgXHGMabegh2ds5L38qStUb1hpgi70pzU6QajAgCTYOvVUhfjhkI3rSNmjTr
ZTidul0CRlXK72OZKjpcUgSmrKsL+g6RcZLO8EbXJZBhg/BzjK0gBumMEhckJq4o
LgXqXphCKNRRN7stiCKSqDoF13WpdlVA7toYp2cW6Y3hO77LTcCLuKDx//qPAByF
Qu15BIRTl9x75rkeyHN4WMUXxxziV3UDNpYZHnZgzM7/gNVBLc0w+UB5EVbmo/Zt
LvPTT2TU/1d0Qi8WuMH17WM8def/yNZWak7yMuZMBXt3H9ZRRpgRkN6kjCNtyGAa
kcyFxV3qVf/voLcokospdwA9oNGGPAndd0uwrABT/75AzwsU1GgKJ/QoPNUIbA+U
F5grQAGSxXhU7tobUZrw1uHxe3hATtK1EW5jezzeO8eivQq4LKjgeEzOfwe070TP
sqUOCCheXbR/wuf/jDWoYfmPtyUl2deMGT6VmlfbBc0T9sFDHrFzS+Nx7/Pc6yA0
UFMuhNCEl/6uBeZeSl92zQO8BnU3OyKBBXIBLcnVsm63lfOHbkSMoce431aXcSAF
9RljbbDHyxWkE6nsdfQlI6W4gOyHi76mVfoz2l0hohvq+GGHYe95AHL5/iTIyNOD
0jRq4m3Ytcte+tn3UssV6TGE4bS4nlALopDj4MGyWJIVvMWGdjVO5WAkCqukRFld
pOWYgXrgIcSgNYrVqS1sIDugNYG0SfFR4XIDR3gJMXwkZAterYy7Fx3QjuX7jW6i
XKUBWnHwtM0k/9afie4IaHd0CDNcZIhCITKJeh9CM6yP18eUZQBkzBVkvxHqXFbu
92K4nac5b79Hs7Of05O3XT+jhA2orJ+3tKlSAX1x1CAsgff4hVcSIoRqx1TkvMXi
wJSvyLlpoOgVLKdivCA1/ZC3+3o9LxaGr/doS/bFc9DknKj2Kc5xAFo8oMmODG3K
CHqo7OeDuJMVGw62YSgiCFyZOD1IoR0J5O+e9BMjPooeDo2xOOjIG0iNVw8l4zbq
Nf7sJ+jHbrbUsVFHdLc+nOLZJWp8qXAIcrvJu4FpcnHh17Dmbp2YYTK+U1yivQpc
490mY8bTHd526DrI4qPy0hPe//Jr6OQluHpA/SCqpYPbmJY9lKCr+CRJfdZxe7O5
84HAWt4iL3Uc5GklYXD6z+9iBxn92Mra/fcCwHe28I90+bNuSkdlkf/k14ZphJuU
kPeYLPE1qUmeXKI+YU+WHlblaUFPZ9+atHYaBDCoL4pIz9idYZgWSqQ4/UEJfYrq
0/Y5EPUPLk4wfjE9jUkxZrBRFqm0+FAqGancgGtPHMwG8lbpMz0+8yQBgeldofEw
HJS/QB8/NMCfaJ8gYtIKxHoauJmD3L904tj+GYorLLNzHC2g84BZFFngIkwpLSbY
p86IAZN8+QclkFD3ADXDNHlhPNaNJ+DiQjYL3KLJ0DtBc/F5bCzVQ6E+hWnjpcX6
2klLymrIgC9LimyaQUL7I5VsdlV/Dw1w6uTNrI3WU2NlAqpWxRJC5BCgdS6k+fma
jckZaAVuxC569wzPQn4GSym+GuRTPWlYVzI1U3WeMh+Nx0in1eHrV4bzU2CT1mZd
FWfXKODozl/BzI1CTNMBqt7dSE2aFniVVPSSCirQBXw1hVJzoEfMC0fIyTSWxVyE
nYXQ+slaTXZrqvmQRhG7GJNAVNSF6pbGVxGj2AyYmeeWQtVE5UWd2fFL2LVwxAkC
AQ9ai/m8JDFDxQuAibMWU/Bcs3uxyFkTi9rMVLe4eFemA74YQx9BKBetc3He+whZ
7oeqQ1iB8ldN43M0LAj2WtTLZ3bPK5WcKf6IUmqLp1qHXYHjVoiEft1O/aIQYwud
DSqeS9YzRXBlVw8QxOS/5ZLKyiuxlP2ue7lMObC61OoZWbZqmnGq4Y2+rSP9cKF+
GdPPksZgty0gAzN71d3iruw/td5F9O6Llh9dbaicqdviWmSNqbPADKMRg1qn2OWs
Wto//zdWF9gU18My5dLydzfylCCUKZttduXDI/611FRXX+LKEFBc5KTdPF67BldO
8pnXl/GDOzkqC1pny5xRdAXzMDKBxPOM2AFu7VvHXZ3PLOjWvlJzP4GyjL/8choh
bDJxHSOoO6jfztGfy+A/sx9oZmTWkUBJQAUNp+JhMtSqbsn8BKlXIXlsv/KVFK0c
4NkY2hGOMi9JZAyLA0EvkCa2MDJztyk+hCyMVE08xivOgGMwWG2dDfg9jnX905ji
EYmpSXHWP2VUJ6ie3fY51BrE5xV8hX7xfdoVfSsTVIwxneRBykyMinHNlOUfoNaa
HVTKl/IOkN20fojHbUouT6iK87v2b9gXsbqgSR1B3eUwkSC+n9Rky13Q5qNDZQRs
KI1v1WWCt4lrVzOtE2AXzo/XPsIXn6ucZNE/QgiayYHTlkjx9S56WkCVU86rNM2y
BNCktITAabdKrnbWuef2KYwKSv9EfVVBZue+SQJ3d7aEjkRTl0/dM7SMU70m4x79
6qGyA6tTCo6EcF4FdblbMhpBAvDrz2EYOKNmNomWOvXOCNCT1u5mAMDq2Kt+Jb0i
8dw8Ekxpq5yPLEFzTkJ0WQzFeFUExHL5htsQuDPIgQ/bS0wzyVVsSAXlp3ilFyP8
JCuecyZrwsPJustlecyTaz0eO4QhUbffTkKS+br0Cq4dkJUG3t284oDuSIreTlXR
XUrzBZGGzAq7j05m/MHE4p2NU6MxXbqGz+6AlEhBUyWPwpVqu/x7tfti5NaKNGK6
4fJ7LzGs8BBDHPyzHXcjcXdlmdGjRRMNOtAj/mU4g2JLCbb3BxAmr0/QURKyutvL
MmNsrNKTtNXfh5D3GHfFKRSD+OcAlOR+rz26R+qEVLiqNdN1RE2mQiszj1+D2F7u
eIHED75RoH+/C88YQaVwwpD+9E0B63z6uF8UsFolFkydAUi9ATcwo7kKgHVwobJZ
oVYk9jJNPJk4guc4WqqOW6D4J61TqwGi09PDqqNSyuN5rDWEQyXktS3kZsqEnZ6/
yEvZGdqU2Kaq93F41WaqBo6YLfbCEdyHj+tsCcbYBqkYsvkL6g0t/ebsSC0bpLva
4U3rJAgw8CF//5eeZfRPyM85VjKg5U5Lbu1q/a6ZUSSMbe2wzDCVlqhpC7+M/v26
FYV6XqT+JJdc6GNxGV0niYdZ3FGCm08EI19txfsSKIGtOMitO081Mf2/yRVxEusr
y6OJ79ipo/XAg8lCjwh1E8FgkQL7VLWiHd4j55XUhTevEHb94WqS/TtcJkNsyY3U
ZEAYd5QzjZ6qe+Syw5GBFXzsKgYiAxsoZZcqxm0TQGYaXezL0F1mjYxEZGsyhI4t
UpC21C1SfNyLQZc4qUITqbMqSIYxmEnhK8RMNBtZl0FnXULihrhSRb1FxBq86a6M
fda+T512nOIrocDJrS6ICDRFyJKPiM52bnVjw0XghF0TRMAIOfh6RJn7bFyvOWTQ
Df3vrgIsufKo4USg00rBuiuBH5J2G7TZAcxy7hR9J+QqJzYptH7vF7crBQa2M595
gUdyaT5W56kixk1k4u1RcUtbF8lNy8VuMB1ljFeH2eFCgcjW1czoiGCCsrcI1OAC
qViWkZek5dZ8K05zMMTotMS4gQ2+R4xjX4TgInwRVq3gkmSnKvKqfAYKzMKcHv+A
QSL105rYQiMOqecQqSnsEPGKZ+gXg5HrANQukH5AvWcosEe/xtO5wU56umxVzEI4
/oUiiZCLS8Cin/OA6ZzI/QJFaKZJ1M/dZpUFYKg5sQ8o+HIApT872uzYVgKrEN4g
O7fqIKcv5p6cIYrXU3ua6Ux/isxSaVPpMQNbo3JhFDCJaK3qY4u3BCuzjk6DNKXu
9GoTILoPfknAWOWa723GMyAGKKlrx4zp0nbwMGxHck4AznpwdbbMb/QHBfAoe3DN
dWB62r+JOnKuyM2bLtdjvAAFE2NOwHNN4FTaoiAYhN9o4uutpisblu8VWuxTPRR9
qkkxevDAQR2t9fTO7WVz7AYwIX153gm+9e7QjOZb2iXhBkP+7m2EJqb2FUHLbKQR
ghpn+LqMzCYEE3VAYvId2AQaqnqXYtY1gTTW7HC/Hq0rnZyIjlRv86wGyMXfWsvD
ebReAH1iNjGeMKU11AG5rIhXniFRGVYltj2t2rhZWw1FrZwjNPanrRB+yUqE4a+B
YepPNiBEalfbDuDpf5rBjlgzm6BZe0GbFIVLra+HCX8fRF6rPm3RwK8V6U2EsUnO
Urm/CDcHI6PEwnUh4CwMcoixD+3tOdm3MIMQmh5acJIBVYPdjv7EZVd+a6yyyEmJ
dvh0ZGs2rhhG74TP7kEeJE/LuVcG3imrthAaeiioHPwhVny9S57MaW8EOLMmsIHt
IP10OWGEVwUxZWw7CNnOBsVS6zCvjtsPGsRO9IGtG2AfwTBsOZ9ZRlRXSI4XZUJg
Cx4Mqcvmruio3nG/yRFb0FiKCQPjkfBStBO8a+L0RKfrcxM1SGsBRgk0IdAhYVJD
3XhzKRvRpi1YOC9k+mzyZbIJFwqpzMOGjW7V+7PxWfy/pixh3byA8h4GFiABZpo0
uGrVf94AJ2zm7ecW8ZrzGs3Hq61fdOHrhCAPvhsq1MTxGDYRwNA6r2rjKpzksEo9
N5l2YxnyDI8opbBszhj6a/IZcqEQtaLdUg90KpolTSvHDk9Wk3bVIcYm7R8Jmfrp
nxObgTAeMtRJGB6ufziyx2FawzFXoCIW0n1/b9bbkKw5mUD70z2INO7Dq4XeUXPM
I97BBiydxDzWHw3vW30qZ8BLB9Q/dn32k9tUSxvGnhjh9tfy91vqv6+Qhu52yBvK
taW30zH9Cgy3kYnBt1+D36BG2OyzMHkZqJNCuauHZBEzZ5O1GaIPGAlqIPGAkQCN
fgeMJkm2aVRXS7k3Q625YzXNUkv1cU//IxjxSta3iWerGqMSHrMBlFQe53mip91+
CXtrqCeRqF5oargOh99IgBTuuX55wLSHXvFy07tyIx7PXmQNa/w7Nl0V8HKpleJ/
WazWtGJKilXx17Zy/paYLe9hFbfJiw7yG+oulwM+VXrgNjI3c3q9Dwe9fCixcdcc
D88QuGWrffH7sr9lyi63x7zJ1wJEItGk+qOCQ+dWihn9JBJL8D1qz2RVHiwF4wxv
eCu3iyC7V8A2RiCiKMT9If6c3hIp/cHI7P2ggZZaWdX7peUFj75INyVtSPKFG+H9
TTbrVnjFt5ceuJlb731QV6vozNpd50v0qgHbFScFY+N+OrK41/HRHo3d8LQoD7Sb
w6aAVnGiHWA9zB8oLrsrODYxFxX4VojUxnjPiOj1vkpktL2k/6YHRYZw4E61+eI3
2yXD14sI+ZIrc5c3Ms9n2MYHN7CuUGAZfBUJKMXeg/CbN0925SvR7fsnyaqtTwu7
TuU535TGUWg6wel0w50GKBTbt9eLhupK5Jitqkv/RXV7RZsVi3C15ZnDuxLyULnf
fp0u6vlOSkIym9bq1WVz/QIlQ/ohvGA4pcnv+rwFblrdxAHXPJxNwKyU4ckm8BbS
1Z53/pk3KNgi7TLNWkq3jGiJhoDC5jJhSiBK9o1M9OVUYDjD/6vGE9LZLrB73GC0
kKNTUMG7FqGGyPvz3zTVXU2327MIffh+qTKAwwmqU4zBTDUV4kkAzSkHEQLr9YWH
FqRqdz9x4GLS+/1LOt7w79z0w3rRz2jDWCSDxawdc2sdZ6nQOxNTv5AQ+EGsfUUg
s8gCxXcJm/4YJumnOpYxk0vzy8sKOFaTve7M5x2oyZd88x2PyZofsxv2PuYlp0bq
oUP3em8P3Ukwxp1xrKm8ao51wWIzG5rn7HlkkD7CTHao6sD2r4gEmIXb9rlq8/uL
w2BEnjKkAfnnygVRtWleZ3/nO1AmIWYiqSAxS3pQf2V7jaiILvxX/PyhnnI/8pS7
IV/J0MNdfngrqjFpKy+NGS7GOi991xnJ4p8Du7zMhD0PP8v5u13QFSZtG5wSD2HQ
mvJuV7rxRUZokP8jpCGuzwWhgONgludn+ditZ+J8rFADOGVBgDJQP3bG4QsQjYK1
unE0IQrE9KJ2EEWvfKBCnctijStC4goMspPEdSDs6qLa6gWry2vZzqM0/oqmq52K
64RRZLQc8SCw2HMDfWZmc6RtppB88eO79mru9Nc/xiBzlLb39zFk8UUI2v60dRDH
B/z3CjvXyToOeBovqbBz8rYO+kZP8K+MiVOG7iYlNCZycZTZ+Qei8UPSCbzqh0A7
zLcO+XAKbLnzxfGk+5aBX6Guiock6OthzNyDVFW0Jvy68mTAlj68WOZtkVH4q6iF
QYmeXqdlVh5ah3qe+edaIgGCxRhgYoeW/wEkt5uqHeuryWmNtVDoeb2LHvOKK42J
DKl/qFVMKL8JW1uK86we4v5BPhW9gXhE7yHw4VK5SPUGQJfLz+W2rSiHKnPNSCJL
l3R2pUrkVtOidfiCa9P8JK7pbgSqaXGXNWhjqnq97+zdvcT6ooyrXS5tvkSTTFkJ
SQC4goDDO2LEEt5Pw4JoQwrEiNE8/EYvEUPoaLUwsfyWzArRmJkf7Um2Zajt4fEm
m9d3tOLzcUpxUNkcP25e5ojfRt6IXjKiu4Kwla/PR0riiNAjIz2xyV9Dr56bNKEQ
QNJ2NH43I452BOLFX8rO5ReMetEt4YBR5O365hciM9dx8xpSbEaCCD1tOVqT8KlZ
xivB5AdiLZQFGgzrhPvSbCaBrFGxWUfO2fbw8Li9ngxPFQZG7BxjG6VHsGQDMlCh
JVMzCyqnOrqs6sPM1FDI/MwpvWl1nBCOQ949CS33p9fbSAX13fpD78JO6RHhUp9j
nOJAQWl4AnSfs3/A/WWvy2fngrARuS2Rfe0UVxjZ/9T6OjNW4P7RxSTVn4ejbOOd
wOBKOKcBZc+v9qhhf/qLCJX9tW4pglxn+4+r3SBBlBElAmnk/p+/kB4Fb//LG88L
jlP9mCTFeZm6SEoOUYbQ27HeYFDpQN1n/gNHyVjtb6hJ4lvKuGesJGqDeUL7XmdO
ChfnIYLJmtzUEQzrP8wnUPXmFbsM135S5LQ+Clr1PX+TAy9Q/IS1FYL94FaQGcqt
JDBlqd6dLyvScCx7Vg4lq4gcIQnnoEwjnN/G9AO5/iegcjq+QfqjclQ9+Gl/GyJV
GvQYOCsyClHT71EYHAYPL1+02Bm305X/nR5XOTSez2HtmJDSljmu/p1n9hngsWqs
Js2B9EpnMCQO4vaJhgZ06+mR9EmhktqheGMcGhTxIk9TOJlsT98B2ZDxPNbFjYCN
LCaykViJSU3AVgCj1GhintfautDGgAlnaEMKDMmrNd3rEfWWk6PwbLt4kApGY6za
CS/daRQVzk70mbtOssFPE/cuBG9YNj1iMVXGtZUPTMXrJxJYbgap3+QxumeWUUqc
ZezQte0k433Jw9M9q/GcHDQV9hdKMnWNNyfgchdUAO1ALYBt+ySBErbytUQaaY6K
dVoxaS1b6h4Owkh8m3ipZlbEzBtLf4hYHiXbeJGZuzXVQecvIhGhuQ0GUPRgVQs7
DdIRykvUKa5HR67VBIJWRTtHlliuPqUSebgYaeqosOPLyKLTxFe65F7Ip0zqes38
gGNts5O66dEB8GVj59CeH4fxMdZpvhlTz9tYaOlwtYvxc+zi2pF8TnIWlgYI5n3K
60qWG8oZQzV8A5w3bSGb6hkGYJEu0A0JuaBLLHbEiRxpZDn1wmQkxj7/yRif5o8A
uihLoRLmE3tk3nf2Aa+CLQyFmb7L2zNeMxgtbwfTSZe0bJYJMKEPoiHzqBs/pIoR
hctYhvKdp0Z4NYByn5eZZ9t+aeni00EEmweZR04KT9vEwOYdA27SsuMGHyUAm1mA
cuaATCk5II556y88bFYzdZxAR+eatmU/VNEXmGSTKU3pfzSl9ulTdU3uak4E6MnB
Jk9bLOUfbm6f6tK5UsI4oRl7k2ASKDHGEg8hgXm511OuE040LHHnVwPr43D7FE3/
92goU8XVBs7v7QnS5CjtVVzZJlFp+x91kaSJAvFX4wnCL/SgfUznrtoaXH4JU1Bd
QMNnvPUQLQyG6vsYCw1C5pca0Rz3uul7B5OMnhRdVS4n64Qlq2t2kwkI0IkSfCdR
pA87CEGUIjZp9OfhzQ1Z1JmRNbpO8DvBodWCm+IkaMVzYYYBJ6owjhBLv/pIdk0D
fqGR04JqRDo40ZKyjsjzTjXskzKzFfILCLXyrBVsQyPMWXvEFkQt0exzZi2Jqa+B
ApaK0PyFDiFvnpGMAgQabilOkn5BsDuIVgDlnxPtCs1UTf+Wop0fdU730EBfBPQA
hoaemm76DDoKVQ91BrCap9eAss7Ye673QQufhjUPEdkXfA1AkkB1+GBeFmXB7cJQ
+4ZMnCw5bNeeAJ+W6E/Qga6Zllm15TeOw2DSRKXowRj1ivUzEMOcsU+FLBxms51x
tBDSnTGegzJIlZsYNs49T+2SNK7APtFzweVo2D7r/eHGnJSG+ymhEgJ3QcKS9P6Y
j7VDjEUKWgunBzDs2oNsAWr97MTsMQxwjZC6Nu5ZjrOrZO/7aDlN09+sl2mh2gX2
U5jxiCTpALPuQ+/R9+372cYn2jrzrnmxBNiVatlnLaSEM18bJEL336iKVJ9AgKWl
T9RzMWBGQVQUPQaFSaZj2Y6W5nNUzwsMObsve2D4214npyy3cSzT2xgCmyyoPpjs
Xr5OiBoWXuxqf270BA0aCN5q9NLyF2QtSbQfCxDc790ATuj0QAdwhKJbrZkurWN1
TqQ8m0xJ/IFapG1RzQzGsZ6OG4cAETXE7FodJ9HQVVPupgMpnU4QvE2LPsSUxhxB
YXoJV8AmMx6EE6QMx6tOL5wTqq2eehICpTwrmfKQMgG8oK5XiTwz5yEiTFHtzMFJ
hm+WC/CMMN6DnaK9YeFYR4Wx8Jc1fQq3w8PzL4ZyVzUw+ssKk6G+cj4Ed1V4zDDD
elFUawEtUHK/PHmSK0QkNnsqj1qErelLr/z5lrwa+yyO3uwc33Xp5/7IgbeEeyen
GYMNoSWluKv3hIqdAtMgvCkWzei4+Nh3RS3e9mkCpINM05DVMD8TwNZ0XqWXIA1C
Bx7T4k8Akox+b0CON2vEppsCybFS7J3rL5qlBH1gyzCBswwcR6zZlWk2WDYxNNxX
vn+TswBRCW/BHRi0FM5GOnYztGonq1WYeL6OuKCcjDhJEaHe0h8pnbLdag0n6YJN
8uOM1lqWUsc0dacQF+KRilU8KaFag/PJPdPnF8jh/+JP85I2vHF81MElsBa5aDbk
e1TyacvmKSifm0hERsFzW3gM/2h7mvfM2AXIUXyMZNKglE6V5xHsTvIE6jY/NVyd
VPkKYbUwoI2VVcgsO7jW+cJmp8yO7H9enPU6pb+Ej78mNdHWG53dtj5OtSoOmust
073Cc3q36NjZkOV7mL/zYDthAGPvrsP3k3SJ4t+fLUI9BW21kYFj1ll2xzzPixPv
OVfWe66yXgxbAUE7KUNiGS6XxT8HJHYDnw/9V/RS3Z3UEppwV/WbF+/QWn/fnTjk
PJQVTCLfSQTkXGSozs2hIsi0wMBcOnqEtH7uHZMInHCPXROINzurtyUbZy5UJ0m3
HjNXaa+0QyMlGxiGXwv3625uDBe4rSPB+gaGJiG6xcYeX3/74ByjD6TW3QVrSIvo
VLUV0Smaq+TTSIFaGZdogwtneu/BzmNhCoOryFPpGJ24bvQ7hOHHlzAL50ssJ0iE
4Y8cBg6RRcdUh/s5K/yMzd3IrhLRt1/miVcgZ6T6g2OqQ9yKJFQTUlG3YXeJu5HF
KrPd0GdqWqgLdmCaWQf9PIJ501J34eR/EF+Bnx1H3ISxjsAFaCey2Gqug1+pHlZa
yBVsQEYTVZtc8lftRx30JAJlHVhsbnWuLJqvyKuRyWiUgRahsf9dYjY1Pv/sZU7Z
OipYjcwzNYhKcuedGeMk4t/hYfMKYIEARnqRpvG65z3v0bWfPSN34v8W26EiTjcg
2CRUkJeY4ODboawm6yGuDA+aX3PjicBYup/IF8ZEABVs97dQhKCKSshpAzxOuSBX
Vhz2P3jpQ8PhwrytzGq8/WDCs/e+ob4d5FVvgwgNe3oPijAiZreCSFt7KtyYsIgQ
0lK3BnZUSQ+FrFQH7KYp1gbmdo3C8ac5t84TX/Mf5npQEXn1Vap62mJyBQbvrWHq
8E2a+mR56UkpKP7Couo1u7k9lup4kEQ4g3ylsYaHvULw0jzOPt/q5n2agbUDIPWg
OjGZL1R7QZazfGFggwaRpKIIqJ705dLoGG8NiieKlr83Hf502MwO9Nj/QU2U7Epf
XEptxNVc8G6+J4e/iVbHB1RzaPwwpcZKKkXsPfdARvoQIW1/KXlxktb2aU7+Y6eq
pfKFqx18Jo/IXcDWL2RXpEQsBI+ywLeknUl7H6bk0TBAvnxxjitZVPkojpgnl6hG
tyBeIuZ5PU4+rKno+u43kscQC3GHjfngGHImA1exhO1txJy5GmE1cyEifgHb07hf
jXhIeR3cDSpmc+UIACyyDEKuAFHkg32UG+FUfpFDNDUp8yfzcpX5F40QveOag1CJ
6Q5afS4RMPCPiOMgJSLokNK/Ys99mh15B0xi00zH23ZrCw0yweYm5y5/L6zaAnZG
04PKKvH1C/XToeUGc45Cl0KXjKjzPX2rWiLpGGDn+/HJHWWFvUHC2gdT4l072Fam
Z9fK/BDJ1LRYywHVSEitLrmXkNcWdAnvjku9/b05H0fxROvaVh5vLdlIQV0gx1+E
1hs+6OdWLy5Jme2AiWNnmTKa3hJYEoNt8c0meaiSTvWUW+TEyIsN/tiCpxMnCXc/
v6fSEGQUzZmjHv7TVmwROOXH9cgw4Fa5k0SMp4vUnZe2nGKLPY7pcVxMdSVuFWYK
6PpmlRx5cy2h1IiWlIbu0kKOkxZvdlRnDP67VUQ7UH2cmcdSJ9BFkXbWTFDhA0WW
qbWsjz7i2ohO63+H8N1izj3iMTb8b0O4plYdRYbEKnh4+GtbIdu0jynOIqR9xeU2
prTqinN95iuEfcKZDZmCtfGJoK2fuJXJ4+uje3KG3wnkT8VOopIzAQrX2Oijl52+
prodJ4vec5vxTxiWrWWPmgMNibzPd+sKXWXgnQG11MQn7REHHrrTMuCUj/QA3HAE
vYojFdjsDsi3wWcBMDi+lqwiB3EO0n2ogWyRTMswFctkzdzqN6acySwNdsuJjbmj
KfpJNFpxOYyU/0a7Ufnu+YBB6uINsQmkrX1BKlUqBcsXp0RjHSXakxaEHfRD5OLt
gHY+nA4nSZitcEQ/Ar8ei4c/QZE7FU18iAcZQdM1SmaFruGYGgOa7QrEY1tsgvfQ
qdtNtWrw/9ZHHxWXGavj+InXIfxPpyHtt6qSTsJWWLc82IboCiwGUiFTRE9i0QZi
aTEfYY8bM626ZtsZ4h0NuGD5tdQFGwDo7BeYrJ83cyAbOIG1xZhJDBow+F7dI1Ve
N5quIC2asHg3CjlYhUeTEmhOTCCuYd9PsI7p41vDcIwjFvZIodwQUvMhHCsw06rK
DJ/xl3/wMMHIAzia/v728itVuPcUpsqC4qJTQqxKSwnLfL5yJEvD0CIIFkvhz11o
F5zCJHt7cTIEiSV3qGRDXW0SaAeylu174tU61YxM7cBrqKEh6QAd3poclna9/NuD
Cc7OtiNo/2Av/ZekXY79nOirQ7LmDV7NT5thIiADhFoGv2TitjHu4JV1ZVJf0bBf
IZMWkv3U1/eGy7/keGzy6QAj0DmUc/Q2wu186ddjYXRTh+nphDTm4tVbpKD1w6nW
lcnJLDuaH7kwPFzbNUt67XuverRFqMvEiAlZJ1l+rNXqD5iVDO8pAX26NbjHmc34
woAgbsBagQ5JluxFVzHboSFRg7m2alBLUkLbjnqTn9dZOJRw0xTSVw5YI8CvGs7u
xxygVTQVQPc0x5Kxx65Aj2htfpeypg/MqXdD4SMXRYnOzqj8QtO3Bj+r6DC5ctSC
LUyatQggFlPqs0gBIdm59/V55cezqzCNxEqEJEvudeqGWg3wgW+cIS4w3c6thIFI
YCyf+lLZ0BuiLG7SMRRK7PeMnWsmGWTYOmY+wD7bJ51raz6tkc98wETiCKBLdBmc
ai+CeFnTDatv1SIqFI5eAMkdQqVwikITDd8ajL29NoQDIYl5E+L+bQqi0bYnZRlI
2PJqdTsf6VRt+vTvgyLDp3Qhch2J/fQLNPk8zVsC6KTB6I/iuUklNnDbF6OhehwU
nJE2pgPRFiCo2E4Hux+SaIHY2aKGLgobpMRyhZ/aAxT8vYMkLxbn+WKrCnd3IbyP
HZa92ND38yOP1+hE7Zonxd7kZyYDlbuPKca5k4TSAYST8TmXJegXCyoIW7vYZPVg
n+w3YgGH0CoSOFvTjXBgcZEQdbHJHzlG6c2ZlfokTF57FtHmTe1Thi8EoJ4/kYZQ
RQVjB5XQgI4Q0y2nlnqVRyJfCe2mGp6FEGP5yqNdwPFBqQOOnXibPQXHWxIse4wF
qKBvsKzCJvjK5PUmO8mnJlAbtw4P6FG3fSialVVHccVoWd6cj7NBPg79Fp+qHiCt
IyoL2jsgHSVY7NYg4RV/h4f04zpQS3wgHEEJ5HLvmlTZd9ClaJjHCnuqlPNjRiWx
oFc625M6JT8n+4g32vmz8YqcktLFCIxo9nQ8ztqahAis1zfWYVyLs3QFQN6W+mnf
095g8gMu7vYEO9XtnHMc/jsxS4w0KmgWa/gCoKoRS0rXttDm4LeOtxz6+aKeIgtt
TtII6I5sRIuta+OoRiaeENpXQVAIwAhA7/BiWCM7yGu+znq1hByMEV1K8mu0RbkS
K6CEBP5CKxn8StEy9Z0k1mgqaPpcmXpuV72i0ZGbBf22JKRZ8WcNmcf6EOn+7HT9
YzD4o2efUrBmoq3XTyZB9Fzdr1wajdSLF8Ny8SebCmI01Fw7r3CE0IbmnuPscCGR
5P7TVFH6Q8RYyJuJuyHqhzEKzHd3h/96jdF9FtWkjG7IwLy8AgKLdyLvfq+bIQyq
Ww0ckkltlYNh8+d5InSiLxH6DKYk4vmZdYwbU/xU5+TjJM8gh7Tp4+/7RhuaQBPK
tj/PaeGy8qZendjCzFppWaU9CnOG2xzi1M7VcIn2EVR5WWOitBKG3gZlOTtw3cqq
ft7upAXtTL4kwi8Hbikyy8/ET4eEf7QHYeB7jwi1M1uvuwGP/ui0zzwA8Clo1kGJ
eAIEiq72qJ8Vy9+EgLM1AUUrhOyxqKs43Ok0hd1HG81W21A725oIhmJW90kR38i4
iQbh9MSeoSZQMZA+J7UGZr12VeoUZrGUZlJYHwO+7hD2kUYrRXsEh0wsgOP2T+SR
+0gTJ5B3nfuMPLOE61p2Rc1O6XD6n/ZpU6tcNcHi2mwi1oHSdyu86dGuoAeZezar
UI79J6M82yok94LN+oRSoEBvfXCucXdSQaM7nzmGLolvDMDy0SRk//7eAM3Z/3ml
2o3VLj41CgWltN2uCkxWo6Sy0W9SfI4+Fz7eWidZYZ13bilzMRQqZDta7C/qZniR
VA5SFiOA5D7fPjI2NugdgcEe2tyj7OPrPwO0fDcoGRIOdtC4ArZkPDx7f9P5TLJh
HSpgMrykTIb8W/UJCcFmxTVwlVGZ9KildVBaTOd4KEIgXlK5xg3iULjgF3CLW93f
fhCcOW0joVtD2urcrV8vGvb1QeOW/ozljeN47MwEnJHV+Fkj7IJ4x4Zy58+WFl4A
16ojS7H9TtBVIwIoO9pAGBbmGJCf6y6OZOKM4ScmODYHaFlPGJ2AB37s9mngb2ak
vJibAnQtg5o/ntJa1rV3M1nwx567EvAQrHQ8jiXQPPx8Odjg6vn6Prx1gix9wTrG
HGpEroRDi4O9Py0B1SGfA0Y/aQUU5PDBlAxi25FkXH9gmjnKwIxsj3BO+qMUCcxE
VJZGX++IqV4y5tZ8JwbmCCELlIhRRLeTYqg/3+PQt2LAnOo6vYOeUuvnn5r4vS7p
jnjNro+0lC6OlTAnsaCO24Z69Z5XkjR3KzVm3Vaavz9RY7eFjCqU9fcooHffLbob
+0yZR6ifEu2CvZHQKK/W5zVorvWkMxcHx0ql+XLa4whMPk2xPdQ6rIXNqGs2GLJ3
7h5unI8kyP9iF9W9UBuySSin0mH9KUJAB4TL/Al55fJ3tdbaTF86BMK3CmEyZeQO
YGIffnQx10KK7kD701Swk/cxCA9eIPetM2mL2r0FfcU4umY9K/gm+ictr5fL8Jc/
CNTvNnXP7ZD+3R+tbsve3y8O2CybYCVOb7itUXX8u+NhqiabfJFSszgVS1YhPsnv
IxdH4S8a2mP+7r9gHf3daWHd8szybr5MJ/gCBLUY2Rfzr26+nkJWX/R8GLGffmcC
92jMZ46OPWztMuezq5ooadhCIAhz2z6Ta6JE8XE3RjtxuiZs6/8q7USGdIRIEWuf
UU19ZkBKVMrwd1y5H0/kAXq9t4RZ58WT5AZGXAFyGCnQ+tItzay7YAocMFAiRzpc
tvldGlOnLBF4qRatG/+FfcYTHTT8FOR5O5IesgXq96lGjJkLDo03J/c66mo7feJC
A1e19wEH/+nphPEamumw/JLXWMAcqTtsBf2rl6bxAszqqxKdXpCSjw+jktO/ELni
eH3CrCeMxhSw569Q9wQPXqYmUxsAO20T5hk0gXY0Zb6r6/yt5cveakTN0U8XjtCt
jSISy7xQO6pXbcjnj47MSjtnMLT6p1IGAq0OxjPesaIwgnlFUm4Vz6ZuoKfBu/gk
HxVVzbFqZoeeFvjxG1ISxVIgxvMp7KzDCnP7EkSLitYc8F7uRmUyM9Ma2nv43vLm
mWxba14RkCRJLLLpEni4Gql0hKYhV0THClICTL1mLqS9L8DDfz7lonJ+YdHSvhI5
IvYAZsjqBOCV0yp3khnQ6hr7CWq71K0t/x5H6NO9AL8dp8fy0ptKhdQtlqdnG3Mi
HYQrMRQquFHnchUUK8rbDJ1CQmpRMYjDCov1qskOhm+8SWIOniTLxj8WXB2zYowF
GavoROpCxMqVKdiGxbKdVwBunu+S1iKZEHUQYDv83AmA597mRNbAt2XliwcQciT/
/4Iui6+CLQRCxcAOfLEyBUHOy3O5q/8z2REE0NGgaucJiLvYMC4OiL4ljb9Fe7MC
vti1+z1DIA4mhXii4/WT7J7PWntQQ7BLnCf0n/O63pbxO42lcCzgANe29aC8wMeu
Y9vsaewOlsawsMt+bHL49+40JnX49nDFNIht6l0bnn09hrQoEgmdjN+yQhmHhyyq
RBwmBxthZbuLi/Izwdevd3QftO0F4N6spl2tYb57bzOcKmqb5Hk2+7t7A0Wqqtbk
ieGs08BWPjbsecjYxHwut4O8bpWqX1gMnvPQrL5ykXh+Q9wYtKvR7K2d4E1dxTZg
WhjvS0uOUCSeH4ymVnFCIakVzG41GQkNsaXbxYNr0Nr0YIkKvdMK/Cd5XJ0sL/Bd
JdT5nSa83hmkAuTI+Q/Zupe1UFyLKKIh5s6+e6rAOwZEaVDY4bkQ7Sa+fqYzApSt
qR9ILxQIOp9OmGpc+SJQ1F9c+P0L+A6xphoz7tKhsz2VcnyCugtu16h4BQqMZEdV
GPJ9qYyR5noJ196lS5Yl4JSMh7Yc/PUWPbc+6Ru2raaKhvKdv+1MEC3frt5ypGBm
+7HlGsQBxvtZBl/r3HiAcVLTsZX0YLAkROEUhaqS65ISe1sRBEbYQ9YB8qFl46vg
vPfaJRWoZMKWBggNqnuclNmU0YG65tJuqE6SD70Qr8Mg8mGi9B3hnOsVFrsPlGqd
R0VG4glvAc020rFxdR9TZWCcv+FmvNq6vc5UulVVw6gmi4ILl1DenF6sh7BA2xPU
yAlDAN21LHkx/ydxQ6vSCDRt2wF49ifeDipB9AlDR8m2HisPR+HlXMlpE4s4putn
RfXjgwi+LbYWw0WMfdSLP4XYrqxNMDuH8F0Gj4bj5XqbHfInCNkvKu3TCtxRp31g
kxwFP7/8gcbDppI2jFNN/TxK3CiDzpojHnnrzaqksN60Fkoy40UdEl5QP69Xl0pv
6sfKnmrcYWE2RopUcTdMQM+D9puIomJJV+Go95N3nNl571WR5MnRy6vkn5msYoa3
VMTAiWPOsEMB7Y1P2jth3K01T3rADyg/1H9QEnOj5K0/oKQC07DCF39TGTAEeJ03
2iImoGev/LLT0n4PaXdbvvksLwo6E7XKoevHoUdNGk3OyB3/I1Hk+AjoHcVduR34
p0oSiMfuoSDzEx6Ohrkn9nQUWELiD9w52GlzpP07R0TLK8qMJT/UBNw1gMtDaPr7
Gyzb8A8XCa8yS/xPZws+Au/DMEDMWkihO6cWImHl4Orw7GBVveT6N1eO/XBHHACV
6ovAhlLqjmiAuLrMj9dZp0GYUN8iqY2t+GNCutLnCJggfMzYPe3UH+tsIkmoeGMt
0nqqHMQo2s4xff/vRl7UU43wc3c/m3Ckw0Gi8j+AkfAM10zogAsbqvZY+KPfwgpd
+YHaWwQgIQopQ8xheVdJRcK0B7HBvpe5DGmQirSq4ybqh9mWOXTTXZSllpfwga/I
Mr9BDU9rbNyzd+KCkUUvqGU5u3rO55wx5eoNeeE26PHG38HeFjjTXewHzClxZO9c
NvLwrwndPX7ZX9JBB494LmEjOBfVrtNGSxwfJ8WAv0+SltrDQN3cAprlz3QRxvGV
VnFMqyubqQSHUwszPAtGvkKxXMOw8/I/D/PWz1H0Y3pZ+nMywhX0ZJ9/fYN64ELs
IQaNWPWsTunSoUHRhkoZHEo96aY9KMW7l0LBbTFDX8gH1w+oralohxdwGFaMV9/n
DQvyUYodO/OoS+IAbYXx446Z1ZzoaR8KJkNCRPbgE+UyUr3ylY/CtIp1sQOBNe8f
glylvT5SHMfuiQyeeeYv0pBfiLd1rUi2G6p79+O3otyDhb8tGSEWBHIPvZNl6Svo
HcN5NvFsLX757fC1CJHspu+r5hh1MTVNosAEbw1uIPR6k45JkWyjQCpxe/OmK1j4
kyIl14FqHv75QS1BKVdgs68ODJnAmdcUndiPihFNeGc+G7EYF3wCIHICNgW4wfBw
f2rc/ZJsYbRg/ENIXat49QDV0XMskjNNOA2q12DYw4y0PbB5+Ed/5gNJngMT04LS
Xr1cDOJVALEJDI+JwkRoyJN1Fw4G2XU5tHLlG9nM/Hq8PlLB0Vgp0d0tuU67Kj1K
9NFlM1qIJQcHG1CKEuVdw7r58GkOojoJ/+OBU/KB1PLu1wCizwXD59EOIq1uk8GA
/AtlujxaAK4NX5Ny8kmq7iN4rglb6sLoumtAfmlbHljJ8a5/8PXcRd1T3wMWS+g6
UueRWy8SoKl6hlePu+2dcQqfs1AyPT41Een7ZPgJt+zu6jg5gZueHNzAiZw5Eiif
+Ws1WbwafEXBOcGrgCjRLTSzaOWJzfCOTOtN9N1GfLxedtFyvsWOs5Z04NegepX/
yrMJhCRjXPj2o01mDrvOoyhEODbTY01jpfM/E4nLJxTQdbIpqmKRqp/e4CFGsRK1
gTa2p6mkNrO2in2VqDDwzrwyK+uMvHrrVlXmjWke6QQ+ScWukIaU57Dad0PHMyYm
ETArVCI6ibma0OKVAeiMdbRJgQc1Y9miJnIO5mC+m3KWttY3KrUgt2oUaHZm+CXO
zkKCDG0NWKA1q5pyDw7oMPFmxAYR/JZPDf89gLsvqrmqdPpZoqMbxVn4TPpoExd1
4l1oNH7RcHmtF2O6SEDMF0spT2ou+pdOlpcGLA7w29Z/OrsG1WzQWt9sUonNj+rW
qt2gT7gfFDRX4eyUg6Os7gQGCQ5V9oU1kv4fEcSMiZmOagxN7wJ3U6UfZZdeReti
IG83K6DLbE9/aDnfnS7MKdsu9L6D2a1H9aHziQE6Z0bJbDyMovcXM9yHiIcdr9pM
Ea1t7z4CRLSqli5/zz9+/wsj01MTfQnAhAEKrZAT8S1Flr8qi/pV6cifO0vMliEU
8IwF+N7lNRXUfGViEujcpmwDykSYraKN4LfTsRZAPLxi/hiGGpJv7fFSgwRJUR9N
goK/0apbo1iqxP6O/CTBpX3/SVuBe0BLGPcCEY+suZAPfO56XoBKdYowpi13AMGz
HpW5lN0gwhHlf9ir6qR3EtMksvD21EcLzfllAtEKSoRXk8pbQK4OvF5JFC25BkZn
eqo4JM2KbJ5g4gOES2CY6IzTwLoYmpon1mkhwqupACbp6wD48BGIg69euv3x3E01
YRPCJNqqmBkLhIv8ox85AgI5cD8oMzAK5bDZUEiJzMkP0Dr93MsEWGvepXLP+1dL
waTZGXa+sVzM5tfWW+LARZqc0L9mI1HbUxGlbkfda0WkO9jdzIDno2lQN6CJS9/C
Z+UFE5kmBGFw28KVOOIic8dMVEGpGjvRfKgCrFUbhS5LaZme6WQBevriCpon8orj
vzEBjt32qyvg9De0AIG0pRXa7sZRbjYXn1VYi/wI5UrBFsMgjDSke2kEkERHw0yR
pBvruN58RY6MiK3Mx/Rd6odGskLyBMmiAR/kKtwxuEv1kj9dJHiXgVBiYX77h5sT
nZ7gpRjCupI1XykhUiPhLsSxWK30zMt+WHyJAYVbhc/JPFQXONQyrZT2h052Z1Tg
62+ozhuq9L5wvniyH/zvrSwwTys0StSZ78o7VgwgC0KfORqifVqnFQEwL3V+yhrQ
nbSoBxxfKSUZDIe9s4kfV6bP1dGxJxxueMn8d9FGn3KhlagWMfL6/WI6aMqICFaI
e6eGX5LAAxOIKHWS58x7IXmmYQXG7/Pv6lj8V/OdF/jHuz8UM7hAfEqkryjpHmx7
W+K8b3q6dQbqWzm8mEEti6aWs6oifsw/DoQkbZmvptZhf/VT0l14iwcKLT1Yixx1
x0nMXg5wgkpGE8XDpSoa40uXbWpNAkWU4REX+IbI4DsFIL8fJUPGXcdmp6P/0FOK
kq94ITetpUdUyK01hrwhobc5Qbx1pqiOhJzBdJaE4kZ8JHYtbPDVFtzQ8eVvtmFv
N6U8J4dNW5hUP+VU2oeF6zaxg/NJHqpBUBHFhbYwv+lINWAByGMJ3v3YEsyQTjOG
3IiEeUpm9eKc8X/rYL7kgyj9F4iC6djKsTKYvham1h7t3hY97sCxs7AV0/ltvX0r
p9jC5eX6CzOJSmOo4W67R42zS0oGrLUi8HkAvSMf4hIm54S8gDPYVmMBGqh7p9M6
nQ0OjxS7+Dq88/5AyDe4krO4Mx/TaLECz1z/KRZEIaT0KVcwIjGESssM84aFasIP
DbHIIc3E2AuS95a82HJSQWb9YqtEMHAZEZVIrP4NDjw8Gt5vRmLbFob0x5ODKdrO
4b6uIA95Vh3xPFlZmDTlvYAvSWVBDXpAc+djuMD7DrqNxkD0PFfmYQizeMHwDH5d
Mt9y6acNsNP1BZuRrDoT9ZEMVYysDMBxG0D7/EG2M/gg4pgIg8HomvUURt6s2cxN
bANWw5kJFRCd1gPOHmNKPQFdf5bYGrVmZG9Bmimpxu83FhuUe1GbpTKhJV2S61eC
wwym1TxrD+lDpg3pHZYE9E2oulqYaHC0PTGS/lRX21LMxHfueXigSPwXpxhAByf0
9JaX/F0cpwBYi2UV9u4OF+FjZEskR6DMIliMvnmgHaTqWFOmKnidEFfI5IY0oN4r
Xi03ZZof0UTlJFugYx2ve+UhC/lsCt0o1oYMaGZKxB++UEL5/JnwbJjRQCSVdEND
hKBK8uoAKQnS7gpBCV7yhNCJJ2XoBWDr79bBfF2gykNbFHcBrJOEkNx9Rk7CSHLN
iTp8ElolxYmvuX8azWZM5IaBPqfzz1MsSQcXB2Y0Y59XmWB8pn945U0XhvmTTnWi
cqFjqrtl1H5ca57VZS6GzRlS+JNRds8Iu0kuQdOP87ItFYo2wvsxOZQ7hchggqEV
zb48dEZq5hf3Gvu/y+J+2diOk3dtVAp4/IbeQWXy6XmJ3lN5ds26eokKuk+/5Sme
wNL0DV0ADzvtFhNBncyMoPOSCGkHkwGqRl3ji6Y5q5HEYw4Fl4x3SsIu1RMV7pLm
plj/ldM5LUw46C0OjNHSX8Po4cmx5IfpnY/ZOGJnWp3lIcR9BOpFScnpD5o7+Kte
46BRpw2BoDYHjz2uF6aY0eSmPEo1OQkOl+iZHkJehhUidAFTaD62D1AGf8G1gvIc
4yl777jvWctrMnlykJh0J0oeihUekqnUEwYqAr+qOe43vxS13EMIq3PUOj0FiNmU
SyeXSdhbqAh8Ce76ODCTyqrkcfvvgyHDMuIy4RCtD2vKpBIMefl43nYes2kF/3UP
K2EAdPgM09/EHaDzvOJK3xC+/4+NKty3YdfVjEuNNuOKQYWUxABTSi1IBoPmXgHv
FHHkeGzGvkO01ylzGImHZBJ02u8MvavH1qZgmjTGFmCbl6eom6d4Z3w5UAplulPi
lvdnTOT/b2T7581/JvsX5ougG2126nsckhE71yE63XSHPnsdqWPj7pSgXMq+65qr
3ehPxal+6l1sQjkZODR5zy1QB3n5S76emEUXmLiWF6pV/N7fIy21l4MjVW07CMmn
BVafAxiMLM7kjYTu7BvQgbuas+aFYk6gzuFkLuildQwH3ieFplGq1huH6dXI+2ub
OQpXPitQco/ChNz5foPmvljjTPhcl98IYl6hFl+huGnZtrgdAHYaQMWM0Kik1w6/
Pfb8sdSZfRwAcRgVdfNaZ95RLgzKIHKvnjUnDkKZwAyoBPuNGCd3C6SNoi7nCfgO
O0xEzXVJKeh+o4ygfwgFF8ULmXXcIeUi8doMslsvMtSILJzRdAsdDsaKbAGQkQaJ
FeA6RiuEltQCIMAAwsGCTNEKZN9Lc/svDkHS83PACDT06W5+I0edyyDIm862ljYV
7o0Sq7j9KpH8lRfsuXin3HkxKzy2DUZm59GnPZP+YzBujcclC0wyp9jMWg6oetN/
PcY779zCCJ8Tg6O5m6pwb6MTk9sI167dNIfTvRGa55gv4jsGq4egpvQukJZCvv/k
w/hjz0fDdUftoji4E1cTPo9zdZinDiBeWpapnrvPvrOp8mgf9aA46Cryl3a4Ng62
lyd4qW9w388DVjNEKQVD3rOyvwa+PAUaLH/kKU9/5LPzGK4BFTsDmazpGIq/ew16
Qn4mKCm0MPtuF43B3wPd+uEcKakd+0GnSTc2nE+2pH78qqZpBf1/KQqKdsEDViwo
1clPasmf1EnXdCmXbfTWCImFl3raXdh3lJFTfy4hOF7HH8FMrz36uf+J8l2BTSzF
njfwM23wAIS9Mjl5aAu13Dq5C5K7IEm4HKr2LgCsqM7GoBtD1F9bHkfWhbzfhais
LPtyfXQAE6NK2BPxoHLNJDtqg2yKaQp5iHZFaVUDbBadU44GQqqAob7W2ODKgC1i
tdBAKZos2qQheYC1dkwN5/glIS5yJ4MQ/zzDHlWanYYOwL7BVIjAHWsiEm7ei2wi
VrBYJHRZyLF01wfeFi9t0Z0wz91lBpICqje3xL8WnKeGP9IFH+0fEgmOz1ID20UI
G5K3gl+9HYuVuoJFSdc18Lh6MFWRSnTpwRqya4Vo57wAw6y2/+QTL6+8afPU0lzY
3HJPb/+7bAykP1hs4spAzTt10iycxbRR3Jbt/z6PmLykrB0nR55yXFbUX5MS+d+p
tWg3Btq2HI12LB63zM2oUJ1A83ETwRjqnEOg/mBjvDlStNzgdBYY30PQ7EhRtaWb
X11Lyg2G7R14ivcaar7VvFlQKO5BYoiF+AFxNawamVUlDvovH/whyqPRUYkI4WtG
Bl+WAIksw8v+cTMG7v7Fn+nqtSjGSGTxiGP1VjtPqQYKZ3949nexYcHt8JeObySk
uU6IcMMXb2s3JMoqQiI3fa2wTb8oJb4afuvmBEWlmA2MAa4o4uuqUxCPoSDB9Fw6
frhRnvahxDlZMtSanD9aIacVtjTupV0q5RqKmL7eIfCXQizXDTtX0jWWziahQitF
Lgp5mA7OtiFVK2QQcFLHuKuopDfnKeUAzG0T4I4qCFqJLuMhuYUpk8XNHOqkz3bL
O8nbpDUrL9QnIP/4FM9hTHUfVR+U1tEkLw0djh55kCITdVqNKGawEBKFlNEpa4sY
zM9lcLb6cNmdLFF9l3GjOm8+1Oaz/LOGSmRHBSclz8uf/WMwXPuYS1daRp+0OAjQ
3qFX78gZbxFYGLSJqVbj1x2eSu7UJYYE7R4L7QZFgjj63Ot7W8LM7ZjUNHOCBuza
hXxiTAP6gv2igYE7VKXBtwj4xzA/hH6SNLpO24XBfIDN1DkH+ZjxDKkqjgVbyZPy
UWHk7LlsnpuJn0duSEZfK15HkXvZj7wINnzPoKk87cI7Ka0xP9s8GtEHCHqh8Gas
q6sE7UGTzvnVzYW6TYnc29A27CuT9DkitZ/D039Qyno16kyLKHdJfgOMb3fDNhiG
hr4XIlBtjr+86c1ie0puwifEhJgrWwZzu62IMZr0EdMx1Y/iGTMpDxpivf/2nYD6
2EtyAD/EbmLv6o8yCOSXg+Kp19qPGjCKz9vAqVkIPyRvVPBrOSAj8hlB7Lkrcs5Y
4yFD8kgVmC3vEQl1hl6X7FbzFwf8sOrjS+STRNQxPKgLWS4aV7N+n7N5RSTQcnJv
vOPGVQn6TYHmjMlc4bCPV0zM6fc+3r/5MzytCY4APPt4r9mazbjKtldMEitIffpf
FcRCeDCVxnYDywzZjfT3CH9fjuP5qzOXz8TaQz3Dr6fImbVrlu6Nw4V9Ow1rEYNG
/4Bp8SimbeeUfaJdTOMxGw8aK5rrsSuyZttQ53NJNXFMxs/1M9dm+MAzjwZptvgO
6aRDnTwkdhJCNEWJTphrYHUPk9C1/hkf6spuqDgRSg7rilAknciLsaPKjjea+rLA
hRKy7gtgwuRR17LfQ/JlwAb7ER+FN4AES4PTwMZCi6ABTslEBS5PvFpLOS0mEC58
nzrJoM5E8g490qFZSbY9/sRNJjD6Uci6s6iW6ILQH3XRhED+0opsUiLViNx1ESK9
WMwlRupldhKITAwPijxu1p7tjHO7Q+RbZ7Q5y60c2e03cA5izCd/6xUy7grxHZ0R
i2lqmW451z4ex0ysmJx94cfpO/u8S19PLwL3DYIKlKFuzLlzBvwFkP8VXKE8s9DL
xCZQTFzosHunZWUu9RvSgs4eQwJgi+XUijUFZdQa00dDWY0l6f9Ppp68rDxI0IFU
l6ufKzmOJNs8pC8CgscZ8+5hcVXykdLPwUxj/lkX/JM+dbfqnIxHu5PN+ZKTeAn/
xeTn5ONmK5+d76GTPv8URxx1xx5DJtkOzGal2nk9NjlErxeva8T0Z8J55Ar/82+t
CU3N0DZDecyqPUZYLTu7Nx4g/Eqf/uvqrx6askkLECeT5pgDvylrqjc0ybN3F/OS
LItpxoXgjJZJ/jfaeNgXhMfe3RN9coghTilZWRXLSbCnvbXU7qVE/GaynfcPmdCC
FFYAtBmubJ1X9io7UIkRTiJr1+wjoqjaYlGP1vkotEyIVqifXbKUv2rhu1M96X6L
og/4RO+ZtEONEAwprBaS6hDVyNRj7lkDYELz0f/hJDEcqSzyQxtmpp1pyUkz4Jnm
sidHSZLKTRXV/c//kY5pJsWWx7hGvJHhfZcpp3juLH/VN23LR8m192iPExjQ8RAf
wFkzL+D8H2FAHdFVT9nPpbPPJo2kEpXcGIhTC3vDwzRkBNJdeik4MDZBks6OsGv+
w3TggTw4WzGudfBQVSHhaICasxPFrjU6GvtvXiZaVUbis+2fg2FD3YlG92AhPvk6
9+QLQHkPxUjaKnlItBuFoWGuvekNY2khehYSUZyqbO2//u8gqpQjwAHAH+22Vm8Z
tDgz2NWxRTKWjIFkQhWdsYRKj8TouaUf1Efhr7GsfY7wmtxzO5/HHPCx0Wicbakh
3QsQklZuZeuC+QGVCkcxDeoNShfTHLk9guWS7xhfYFFMQTIGv4uT9cOpbGBgdlap
C3niXkIQ3LszSfQrB6gexDSss8E5i441a6nGNCq/c1KWb3Q+pL9329klUgJ6D0Zm
4wNTUSRdFTPmV/8TovV7tDEMjywUjE/zDMJtVFGZsupY0Cht6DMm/WNnTOp15ho8
Xj4KMniZja6BgY6YQBam7pbZAWULfZrxLEkeV/H/uyylLVxVeC+hyoD+4Eom4UdX
WARX4oohyBFWjKeaz4GZb1sxXFgbX3B9CIUYIeNWjH/gcQPu8HwgDNJsAY1cKy0+
mm2+fJ0Ut/Gl4D5sr2W9Du4YMfclFAMF/m3VckqNzBVxcimuUCrLp4ay0TQkd6jo
iOW1XzXuVSssn3hmvEiKV5KkwZ13vO3TEMXBxNjiou2ZHMv4XKdFU6Uvpe0v2O9l
ybjDbCK5dAxVblGz6WUxPJE6o4licKJDFrz16CQTfhtHWbBraYsqK5CPgzB4dST5
mRjjnXX/AFtrS7Hn3l5GRMdhRtzj97VKSb3j5TvqR7fw560LU/p2clrb7ZdBTUEO
3W5sjrb1FTMQfccu4kPKSsK5s5zZW/FKAl66QJRCNInl5vChaMIbsBdeVNYq57Kh
SQGosN0Lv0h8XKiAV1fZ+ALxMc3BDPPyhF9GRlSOvu2oh5CuKkft4hxDKZO4xiUQ
yPpQbZSX7RaI7PZANlUwpsP8PCQslNBQxv0UTTyCxwBU/VmDURBR6y5MPMk1HF5P
YZeFNwa6iIJi39u6EbpcIXAWhSdZKBD6Ex3lgPF/D/f/DS2JjkouGa+pJ/5JePhD
wsB3Amt+eiLJM6bGv5XOqJ/xS06m1iisLOi8+ayFCioCQJkB0cEeRUiMnASJuZ5g
xvqZBz7Dm/bz+V5b2OeBUphGoErYspX844/b4mmyawqMJKgA+SOFa/QD6xRMpaKX
106WHg6lG38k1IGHpgm3EAhe1J4xyAN3fXY07cl3WTdDBGAPTXNk/SdTDGfqScme
28ztrva2rC+0jHN/OhcEi41w5tTsIVOxBKHQGqwnC8UpBaosLE23ek0futdnzC2B
Ezy+oK+rkRUv/uAUA/vV7FMPzh+4PVyhw0GLsKgEHyRJR/S22z4wXItTjr0zP20T
+ouZ+X0brljp8dPCmN8p8WtEOHsJ5IWe7o09n+k6On0lyXmt2pXzyEUsUkBA5Txv
2NDXk+s9t2JQpSdYuH1ft5r0SgbMPrV5YxAifVTdkeI37a8N1fRHE5WGRfCnQHsy
tCSWPJ+wbAX4ybJPLxyaA6bJsHvTchwj9fFbKKdN/hrdUoyGVvnjxjsOoOWEBH9g
qsamLWQJ2NSzKRiU4TAk/L1FNRas1pumsuM2bYkAxLvs/pOr/f/Ciujl2l/sYRpZ
cnwjOLe9rODDkAxr/tyWZmc8lWzSD0jHkI+KReLomZKcu6/5E27AVp8msqC4TnXS
iGRJUtJu0o3nktNedGR4ESI7DS8Fy5BHb2F4WfQ1mUdDNvosXohA+LxDzfVfO3Cl
OVeN+MuhkBd/W3jVCOaVGf2ib4d4TNfrELvU5QkjslURNECQzpFS2au4E6Lj1D6o
0h0Oyi+fUW0WvzmzTPj48YCupU7F9BU9z9FHGt3mVrp1jKi1YC41dp8bzycSnM7F
mZxEQ3PLtkP0Pj+pWKx5NW0zYOJl6MN2iNnFHjtwIQ+TWINwkRlyxCxKE6QUJWiH
fH/xBrIjLpfr1vv/Fzsrdfjb3BYoOydN9rQ3W8PzJGJDXfWsuOh6H73okxEk9Co8
chqmWjhMGBL1QR8+1fO3XQSz7DxF0j0iHB9+yMPerwkiJFMx933SDFhw6xNU/vJM
Zc9gkAu7neRwaGw3rclFkB+sg6nznpQrDjnH70CVXULAn1pQPusHNUJ1vFkMbfy5
0I6eBq8A6UUk/fdTquynXHv/vlzhetGSuIMeQ0gIcBFw4EpgMMepEDaMMcuejc5h
fkTLrQy3cPmGfMqFe0BSTvHWEn36j+GI0OCmikErLdt2Se3ZtgYYdjKZ3XghNPea
r9rFHjFEgWYyYyjsic8THM1Zm8Z26s1hKxq3Pa2UJhHeOo4VGqoiadbG81MBHxNo
giARzE3x/b864udhGnqgvgnaXD+lDQ1Qxge2AkKKv43UyhM9LLEkDpRMuEQG5GJD
icvsXM1iyalO3acSeG2XthZKShra5Pjh/hcIcqvEkG+vYYUDQk7F1K8cYQtP8ayY
gl5psK5gqCQyxhnoGZvgMht+eN2ADS4hTRwdT6/zbF78O3LemFMY6s4t7IepoMz4
HgOUzAD1zAkJA2j2REsegPiscHMVeWwmhsNF4I9J/23IpVaqKDBpz7e7m0PaGr3n
Jx9DRu+XM5rxYgXUrh6MbZEMh7kbix3CBeQC+VAEYpH4QIioJVR+8dR5N4t/UhS/
Q1BmyG3OHx+tFHEHzY39H/+YXsuQwZ+7taaIbNMP8fRWuzpi+CtDHrHGv15CLBe5
VAIFbe9vXJw9xTnZmoeZqtqzqEQF72dwoGpqtOJ3Fw6Afx47/aIeWAiMRiGKxN+h
jECcd8Q9heqSrGHLrYVCodJMcWlZOTJ0vwP0McjikGaZGo1LpXk1KJB1dSkB4Pd6
cv2XLsaKjLvB+iXSCIrOL524KtRHG5Qk7RKTiiYngYOydHNfnxHvjZF4KzP4LGmz
BpFJjXOyN1p1b97wRg4w9ZrbNWdyjyRL1dMuS31/VTBznat2TGJsGsZaKI7/fH00
x1Yb7zT6X/ruzjGP7ojdsJvDwMfR9EGxfYXWeRBKeHVPayshP15QgULykO1wDiAr
67jYVZ7pu6pboCThpNm41mXJ0nlDs3hwbDXlS6J/8LB7KDtTSEc8UBVvMj47A9YR
fuSmKkwVdNtokugr5lGLU8B7Gi/W6TcuMcGSUw9xRWcGgFjcxebShVtOIjr3c/+B
ohQmAgrGrqe8JnGUgqQ/h8rs3nhqhGMVzJG3kMV96HgOxUpP0MIznTSz/VaJgyOT
XcTX+8EKF8CEt0zeqP0X4PrcrfrN3v/3ezjL/JN01YpiJ7pYUqHEShzcqwAqXYbt
cKoKTIoHGeOEHM1hQGT1j/Ea0bWoQU0aHsAVJ0eELrwvd4aGR1CCf7Hu0v3KFT1H
JIkVx3LtU3ZJwSSEFVAhsn7bacniG20wCWX24sazs4Ze2TZCYG55OxulQtpW5asF
qDXRdzAB/caZlUgDCZAUPmiBzUpX7T+tpM/HixXCJc7KE2mMsM5APvSZ+12Ogdwy
0T6ISjSp7mjqRScg1feeyIgc2Ucw0AizvzfFs+LI0DaDfvJF4qUJwr47BD1VloPH
CENiw7UN+1jCan81ufX1ym9gsrdDxaThDM3ftuHDeOmmVReHz/RMSc1lg459h5Lo
idFx8lD+O7JLk9uy7bFAlyDFbJI9i7bJcfcsKDAy7Sk1sK7ocoXFt1eOCnGiKCnB
vCZeXEUS6r3odaqDM69diqNC1jzvSGqXf4cvfrE0PjjEHVpnpuAVC2wvNiB5zk7e
rHAWyVkAiep6xxDLYejRNkZrv6nrc7xzmnBm1mKAd5eO7k/wVxwVyyRSLq68k6Jw
ohpnJxAHHPn3FTTbx9Xi9SfJDZdQGUnnF32+jGv0AIPdliKGYsfOQ43FFyElNXpw
qH+OpfXtyFbiPf+L0b2HM4ymSBMim7aFF/Cyf9B/R7Y9mzmNXLTK9tTew1PJG0SL
62fGtBmHo7NWwUOuCV3qiCxHrPNd8fBg43U93XnMDzIF2DohA9BsaswM9OwCeeBq
bQGCwdO7qQwZS7RRdb3VmoqCuLDedAKja64WwwfMe4zyHOVRkoRUTDrHUS38Ucv2
6N+2chR06j359X/p5Rr/BNn5dWkcsigVwL2vcNEdrzRSQznxJ8stHGTmCtONsHNY
AxBR47B7vudx2bpNQfWc4lD/W6ENens3HDH8roU0I/XgR8muwbKGapYauYFBaZaS
SwxF3US0c02/ThMmlfgQ67AJIEscU5Lbd9ZUkvwwSEopVijQ1wDYG52vq8YRkxdb
d+AJUkolNlK8hLa8bOHvckCoKxZ8h3IhQzDIBWCAB65IZkfMt9xM4YDthOViTmlm
oPLjyOuMqoFOSi5iWZ3fsrzu2NmJ4VLQEAee9YqENI4AqEIdUcFwrQa7LL40C9fe
EsonRWB0g8KE7ME7zkZnvBIZnWIrDe6YX66mtA+RVHgew/A08vYlm0vbRtr5vzFT
l7GJGxXhYr08cG43JQfUoo0K0MF3NjkW24sw5YoiB3+CGBK0FN7FdatkMTEBJjwg
6oSR3u7xCG1iu5elo1ECwUu4AVE/lFeUT2lbMH6eiansQzM+e6O9rauGny+mY6et
Cw+l65Hi5pPb5WiZhcUMzm+pziOK3U+Uu52Xrm0blXVM7GHaK3oD9HhzOyliGcBs
ZzG90DajRS5GxZfnPXE/vGyLWiT1wSeBuMa0FDzOs8ZMp+W+nQZbCt05aXjZLzi/
4oH+Uxev75uKuvZFaDITjklQWA1tGbOZ/Cz5zwMmZBI7lAKLIBphNBnEZZXZrCqW
GQdUlwoggfBHth+oP86o8umfX46Rv5TRYhjz4cJi74tuG1ufu0huLl3Gp0V874xJ
0QiOAwjP6/ofwJBoJOHHVlyeB7ueUgRqKCuv+89A+Ba1PxZk7fGRDQSiRtycmH0r
HtwLFfAZUujFGPOJQ6E7vED/nHxIXJI55WYg/CSHE3k5nCHElCytDk7zZFIf038S
knCBIbdijKG5VLfh9iyWvZJ2Ocxc1B50FTaZaBWuEC8v1m6yUTUDBRit2Dn/1hD6
cLQrFzGgwZC0hOgh1CKDqZIzU1nnrSZx+X/LxKNMAjf8fScFOZ7ZxuMbyAvRcbsb
jJRzS6MvZzMWxz2je9Qf6B5mw37Q4GhH5bpgCsufhGZeH68iIdTmUIedjBY14nPs
UNMDo6HgrWicPwVjnTNlNpelnOBFTTGolFRZ6/DB9d5c+8liQdkFiVBXiDcB3t7r
oazSU8GY8qH9UylMM1qB65lcOI8xq2eqe52FjFgCRygLJ9H8VCHcoqhXIHnTPiMS
wvMkvp6Tr6IK/7JCyvWwP1sJQxu0OWmlLk8BoHd/0xMc+z5kuYrpLqYNogjN3p7e
48ZRu2V5Ykp226yWlyoPyjEF0ppXTUTX9B3mVk/4gkJhEM4ZtWI11wmYid0tM25v
Fx44+74b6vz8KqimPm2ZKlCxC9xqWLfvtvPUbUZMYA8/HqL+BbS+yQcVLmZCe70I
lzTJ76KC5AZD3nRIn20Zqvwip/TKpkd/6SUWfF8/u5ivbm0yv0xWaTrqJd7pi6kB
X49UKEIgZxVdJWaBieaLU/kCfH+TJ8/BYwp9ljxnL8BB+PMPN+Pd71CB5aPxorx9
N0Re1rUcIIT7ecC9KNlrf3UVFaHGWToM1dhAXrkw1j+L/56lPqImCNY3dYYQdj3C
v/Wdziaxf7njY4UvJNJwa4pX4fOHdAARM1gu1PT5WVMtVbPlcKEFZAIXz/bvYz0s
e8skmVvHeP7Oj4r6DZZk7wh+Darvu81Frby/6qP4UTsSO4vDDD2n+LxSCIZChvoD
vn2MrxzD7Ho4aDfHY2tkugAw0DtJBe9ZimB6FRi/xe7vsIx/azTH6jN/kpPKJBVy
ng2u7PwCsVv/MXq8YkpEbL3Vn6l2V9GLW4Nygk136t5ppoHM15D6NtTYskvv6m+r
R9QdJvAiN07BKI0W1WyEOyeffWQhNYjjkmGM/wY81B1uKty+lveuO1LvcsEp1Hlv
zXAwCUhav7rU+VOqgcG9SNZcROEKXRfVPH9LgA8RtX2jnYjPKQbgiJ9k5uQLCSDg
ViKPg71xDDt64SWGL06AmgUytCVZyAVXBSE+x2ZEZ8NiHVn66awwQ5VpHqK/dkIo
iyUd1624/lwudcIIXQ0topIRfi5T48mMQxqptVMng0qfIwcYyjwN9UAP3ICwiJ+2
gfwE4b0MuwKeEzc1lb1IOwdX90y30oulpvIpQc0oGXATwSAlFsO4NLgeBAqFQbsA
FtoKildpvhQv+BVfWngTFz4b/lqI512RP7diNlp8QKweAIBt00rcgkXu0oNlLaMO
qJVgXP4acxCf6nwgfRYeeqUgtIClEWFYA69MvR260YsJBK3MlS4pKW8xoS6FTF2P
MO2+WtQI931D1MFzmhYQDuycpY+64HzBt7HwcrXL45yluZm4+9JGzC7HLsS6GW7x
yHpqASg+hZF9zVi4jKch1UJN6WMHsGebqzk2GZfkN5tRamxnMoFTiUlh+rHQjAyy
gWtgq8zAO7Fd33DsF5VXgVONbYxAr4wSyzqHNMzYpmIyzXdHQwLJe+vPi9TIvSu0
G62Os66z3BolikIsPt7e2nWH3jjO4CFuJhavXo7i1aQRwwcUwYJvPY/OeF8fnp7Y
jLruyJUnhdX0no5Wi5nBn86N6F9ZlvEApWWbhQa+GR6Sr2GWTk2cDtBJtxM+3U4B
NBTuTE10j1ITSS3J/zvBZlZ4mjYpRVR7FxRhi0qqTRmgx+fdS/WrwzqVSBEuvKsn
oj0Mt1vcIPjKlzKzB8T9ppon93fhZbyiMG7+O7J23E2QgfGaJ26tvQ416fOlthSK
IQhnYDUTyLerTtfu4oWW0ZPSsJWJdpN/44RtRMVSThYW+XsKVcdKf8SA/FVcgpGz
RD4qrTCaB9F0QdAvLUcOkL2JrxoL6FdT5Dc21i/k3POVRAaNoce3Rp5xLgBb2WHe
ofyrxIyciCPcnpDmwoCKRnlJcZj45lkJ8ZtApJxQAyTvnKxyD1b/SnYiRVrprZ95
El/UZ7Bl/7/cyvtH5uVxrV2++GcSIeXVobafj263lhz1sOW8o8VyxA8LPFsSz0B+
mXMvTiZxhEQG394vWOxfLNvGDm2+35dTeWtJ71Y0XSva+mhhLIXkVq7ir2CQSoqo
+vyYmRoQ4Vke/Ps9oheMSc2RvekR/OvaU54rmOz8F7chvPe/SR2DX07I+9YGsmtU
v0VQa3ft/OpABT/2xODTE115TTluaWhBrJWh0V4h3Rt46RUmNUrPm3iEAWwe3HxI
JDNqDliG20iPmXNxHEZ5i2FLRDXbl5oeH7cZNBY+i1FlXeUf5zWmaDrWSvYDpUTu
iQPE1pwx63dpB3TrORjx51JfS2yznAtDgnsBytnm6S7o5Dkaf27lsNvSWnxR/gbJ
ItHW1UXJqRohjyRgk/H9U+I+2lXW2T9DohemCw3Gx1LQ5mtKMG/Y9yWXK2INPn/O
O1JBdtWLp8UAX2WzGkWK3xoFG+jkhn1cA85kiLXFRK7XGCrP0ck1o9t3qJMpqp7k
jMReyxrd+BeD1rPu9Tp0kHA8KpRy2PSkVyD2UCRSD6lMDOZqTowioRqnNOiq/KGS
XFLA7GlrxtG83f1F4yMxiw1I1a/1y09cJ2jLhmJwnH51p3s2cQz8K3ISJv26WbVB
1IyTkrHnr8P9IX4PatDWJm2TQye70j8Uh2JFi9SbTAlk8hC+kk/135QuRQ8lUuUF
S7iZaggUSterVep3pijoqwyOGshJPC+yzVmJQHmovyZfTxOJKCIjy8FAEFI+C6TG
JxrtGrBnQIeWLzL/EVb1Vby6b7Lc1MwnhMTffYFhPWIvVp0KFO17oX1sOEmXEE5Q
wyHC+QbdyDc7Xh99vx0kJXM5+NYuObbqmc231+urU5lV16ugtGSCeSkQNYdGqykU
Zem8yjz5HrM6/T8kTh3gb3ArVpX4PwHcDt6HUQvmj0Yi6Ca5kQeFa2VMtip3lUDz
U+zav5ic4aSTJ2kDS/g9TlmOr+EEZSJ2CqRmilGn55GMcNGDjDfsfdNOGNITmqdw
xRvXZbCXZi+9hs9gmIhEfD/A4B1KXj+dR4Xil7fSDPjKZEukaVCE7oalOk/Il50o
yJAEsQjWRhadhvqytwkd5heYXxp5tx3wpBrVMlPNBKoYzFnKAtlWaJ9cVMIXf5Fo
QJimy8IpnGYxqzNIb2zcs1myD3Lvb+O6FVhN4oCZ4dBItdcDNsI/boZw+t8AnguK
Y7dIxym24chgGqhqh64QJIbEkQrOjQwRxcx887HWHcKH80KckPDQXj2wgiHqvKQc
iLgY29VGUP9c+g/TrugWOtVhFQVltl76SwJm4MOAF0tAhxryEyyPgHdKFQrJALk/
czWTEdY/UNRO+aiMoMFASAasqwB3HPBgR+oTyqxdu4+QZdYdhvauJb+ZbnuM2zvV
Lb3A+15dYHPImN0WrfCIm3hv3xMFL6UAvZ8kcWwvfUjVRacSErkxVidrcDl8Bwcp
Hqujwy9UJXIPCwK6f+3AnFNgAXw50kRpFpk//fVNDIUdo0ggqoX9BdE7A7CyC5fi
p7/uM/xhl1teJO8pS3ZacmPCD7MLmUF07qTV5Pz7Db8kWq0rKG8PNt7y/OflxJPl
FyV0yPmLHuhTkvddkEgRi11wLSCZQhGMnBstKSQILX4KX3sSSGzuJDPPeqALP40i
N0nKmZyqB7+UL/KiqRuZqv7xdU0CAVvZFftlZVoPk9B/OPDcFCP2QmcXNvoIv0WI
ell/PqISUgEJXwYqY39oPCy0fCpbl28oyZvzlseZgp9/ldo2+E9tw/ZHZ/MIMg1J
2NRRPJ0YeoKZQ2VmZpMMgi1ys/wlGzYJ9PzK9qL9EW5i86fQJSQtqH1vYQ3SThm0
PiVKzFKtFCCLB9hYlKcZWFZxQ7rpZjaOVlg1wpuuMNs0Prl48ayKoa1M+SXi5etp
rbno9dl2e6qBDaDTpqgyvNiqS/+beXvD7LCNAWyv61AKm6wgvOMjwDcyRpz4ssfT
wQ3mXgLaBSLL6n6Q/Ezz3Ab9gLILTZGOn9vY/n/ZhreAlm2PMwxT1jsMCtmg3afe
b9DVFN0JCvG7OQlCvimFM7tCZCwT3NcMJZihaz3Hj+BzMNXEcafb2bHjB0bp83+I
/l0cQVFGsZNEwa7TXcx1GXsTfRgmv9xuMm8YDPKSnDtyc3ceNbeJGpD5cVqo3fW3
c4JnzV2DUD+SJeO05TIH8+r1pUbQiHBIwnagUZYXB0qrtTX+Y6SHja7+AZAR+z3+
5OXRBWyNZCdVMvk2kKy3t+L/9q0BjzO18KyhDSDF/Aex/woc2TGga9yRQW/DTNkP
De9MhH2kyjPgx+tub1KaP1IPDlKiv9DvNWQkjMt+Hc6JnoCD8hl6Sd5kETx0HBAa
DimGjnw+Wy7HIT8WZ7+SaHO5sTPW7lA03H9lvQl/351aYDezwzqPjiYdR5d0OYTl
e89wc9hvZWeTc/YbkI+Nw/8Z01BjGCJrFbC2w3M5QR8rn9nnYBVr4TBKZ8+bF2MZ
vIcC3Xtqc9v7UaqUgWvYpAx7lQHH5kD0Ih6+kYqqoren/D86VvxusfFq9VHLx6Tq
oeV+k6k4eqehQEwbJSpPDvTFNJvmaKXmS3XrcKcZ3i3P6h/SycuHa+6ydAysqcZz
XOd7mFGXFHzI0nQw9nLxE8qB2HBuExeSIOyo+e4ufsr07zWiqtbSu67WeAt2+0yy
8pvgjDRRJhXUwSWNpUdukzGyDb5rj9P4kLHPwt1cHKesRAqmexXf/UU7vhe0MEU6
aPd69cZ2gJUOmKqhXS0BpenKXZkBdaAp8Sf+9LJMwFbtUWe50RaNGs0xAodejOpR
X/h1fo5vGkOmQTpB+ZD0X/v7gCllxAng/WdQBzOGfriDSqsBlmFFBGJggLRQiVPx
UMcMT6fAExSJUPRPItpZR/D5p2w84aLeSC64myXPRoJdBaz1bMEMRrFJrQaod+r/
j8oqMbBYH1UG4WdukKn/wG2FWiGK4rRaFBkqHA4kRPp/K6VtZhuyFYmpe1DMOZgi
xNeN2UySS9wkRdaoB82QPikyWDllR2ptj45RexFUuS+W30L8synoPsw7vgROlLm2
HMoc6hCV9NvTWA/jF2U4l6S0UVXDmj+HaUeafLGl0UDB61HRoXnAi/nB/EjYdWDH
P6kxAVYKTX0ELdIQt5b84t57BT10K2zLZveZd/fVWDgFjfo25WVJuQEr0HXFrk+l
SDMb2uTZDs/hUxTXHSx0/CUfGNo9Q3OpazRy9Tm617DT1Pgj77moB4uD4BhPDdtu
hyXWRkq/2SoZs24qvyhRpuUxP8vbaSZBuZFWRWPr4AlGGWndKtaDFeWuMYVCmFzQ
/4N7Ruzftg/kV5NTUnBoueIIdiPk3HdzVXTPzgGF0fe914FpW3V6AHNiadJBLpE6
rvIuUL2brHpPjz/xXH6aL4AagWZz0UB7wQi1nSKF2C3vVipxLDavX4oD5e3qkkrx
Jk8sy8pqec5aekvCp3bYzXdqnFtlazUFHND/BcwKzcvfYF1Ule7RGcYbA+vFoVFU
iNhGwdDN4m8KYR+WHHquTSaIDbK122HzmWF3C3mBpMcX5XbOkXn8w3RyLjSWED6p
/vRCbhcCIn50RNYZ+SrbvLJlJZ54/4mPRFzHZBtgxugmsUFJYSQHgBgBBkBA7dYT
7qPGQ2JbjMFfdeJLJOvwiBLo2ZKabJCSYaGLD+tTha3jt1Ud0YD0pvNZzwoAxKRr
o8LZ8hk3W1qNEwGordHd8IqIU8B/mnxglzGtE/DWPjVCQnw/+XtDZ7Jz/aRJ750/
GKC2QJl+JLcePjfa17wpWNVJTN2Xshi/9XOTWro6uaEN2qvKABeuR0AlHtaDVclu
6I2jbPe4pD6dOo39LIvX9PhN/L8yDzAQFpG1zEq0+ysOzsWeL+QkNsMQgzt0gx1g
c1+lHVR1UMKKJIJCkVMp38N0uIdeH+r9+RkSD6vwrpLTI7TpDvx+RpSuavXxjA/q
fn+rLvMqu17l3p4vEjFSdOehGFhrNP8RupNj+C2uF8XbW/Trro+tzF1zHIJ2Dh8h
TUXkdB2REUFevWsWIJZHAqN/luNH1qhMIQWyOvyV5DvQBfGC8pexNI64zK2SFFDx
I+Jy5vlXSGv14Xyj/r0QtJxoWIVpNOTK2gv+i3fMtrxAP7CE7hJUebH1tyE5VgkY
son4ZKE+PIltuXUYCIwHMX7l6oLFbZkCKJi6K3rHPQQfZ9E086BFZ2D5jRF7EAI3
xYglgqWOzusH8tP5zvglpWIVj4RmtRg61SVXYQ75XYtifOWfNxhwiSXZK/z1AgTR
1O8hELxGjqUuZL8QcKkbzjK4EfWuWMjWO3vt66/zwxBip4pI+hXsObA3Wiqkn6bf
kF3jOXwL9AHbBKPfDbkq2l9A49xdpUNKeZ8m+1aGaJQVyjVH3YHxAtFJx5RaQeyO
OHrKhYxz/Zlq505w7bcRbYPnfeXSVneVCh5RiV2w4qfWI2W2F6GeKw/A/g34E1+A
+b6a3bWZUmTBU7Stt23ZaxUpu+5haq+SVXyiJgR2js2wT23aQ/yAdVeKEY5WyIQE
uKDs+scaMNu/ogWRT+x4lmZiCNgI4WmxfbaG+ZzYc2rS8GzVDoTEE6INxCtz6xiC
pnf6QRGAdjOsoWRNppLzQFSHGSgf69+wTae+Z/VaDM6v9FMbLagBCO/ZAbqYe+kP
rxM4p0QChRhCO4gNolV7RO64wo7qQuIF68TxQ6ezFuJNomyXmkPy6l1sug/GelyP
fYQtdc5eD/jyUtoFpFPSUMqDrmiHr8IJOj3RvD2z1nQiXQAGHKBvPFEgM0Kpleet
GWHSO/B1Xh++/d+uyxC1/0XPYUwHUk23+uHuhBvqPu1JXAZDEiOGNIx+eJwfVrM4
jt3pnqBJ6v8QW8FMn9szXNtNx7MfuQMqeLo1Zs5Rmc9dAdvgZbLdyY6b0PsgbX+W
eRA90TBlcaBVIrmWqJRuFhyJsmciZpHokj5NUhsnZ1/QBgFmOQa+OoA3bTytEVDy
HVk9/8QP3WKRSZYs2zViQNoSov8TUUtmADXM7c/BcBsla5GfnKmjS33msWRRoSO+
7fgbEHoFypp57LbY3XIDQ52s+jULZSkJgu8/MzvJvKyh6lTNsb72L/kkgtLZtV20
jyk0JJRyvxkJC5dgNKKVp60UjThQCZfeQTI0RrbPifyDZQQdhNT/MGyfjV9vVP6Y
itT4WKD1aynnLrni8L/LR3zJhukIFMrvavSNIXrLMhJX79UH4FlytKf0YbRMW58R
SAhzOEigfrjhqP+9VGntAN3Nnaaz99HmL8O7EEa0xkxKXzwJF1+k8/Fyu2s8Wrjs
TMNRHASpz9eFPs7uZS6Dg4csq4VYWxpKBlKfNbb4I66jb4zI/xZuLhseoF7i5Nzx
8bHN++ULL2/VmvJKCbvMfCla5Iz3OQRwq7YEFYUK/sj6agVAKkJiewqEq0GJ7SbX
qw5p6YwrkoY6gPVtfMyX67RimcYfPHBjtBR5rAvRn7cWEI5JCAYZwqtRSXrnnUHN
OxlVZG5rTxyEEiVLSHPgYvTM6EmXo29rdU15+oDDA3qEm53k6wT+OhEmj4HDkKU0
VtyvZbn919aslLX+hTS15yofkhGyskAK54cBqrJl+av/Z477GCLuk9kgHrQicKRK
+phGPWSLcf6Ff9sl1saeaIF8QZ7FC1RSvMaOzb13XQjAVCnfs3/CCUTOYqcHv7BJ
kO9bp7hhYZqGoawulTf9zxbWj+wszf9Udu+o2isXklsaxdlUp00d/WUjQmh3nE46
7Be4rYi+YH6DnBja+qdDf8c9sbeDTq9/dQ3EbNDDFtOL6E03p4tiEMJHhLV3CjUs
idOp4lLvFKUIIxRBaeMBtfarFO2mJoyqmBbb4ycnpgzhYku1YLriikpum2YfoyUu
uyvIrlUpdJ1lD1yzOWGAOllgGjDDW6/6ABLgbA0elRwy8fdPx4c165GHaz46hV3b
ma3yL7p6/CTdhLtWRLvEGXoK83ZKT4V+n1ZgdHOGXxyrl0oxtrR4DRYUjluj43Ru
PFHy+a8qlAiGUYzgHf9WY18lRkZrdBCQaTbG6WKqAus3dYesa+nRyUtwmS9K01B1
Sf4vKGDan+WJ74qaoz/IjpXL6cdwJ958ATFLEzgdjQUOBM/zcI1j9wJhfTKGPZOQ
5wwdqrEJEDcOHkVczQIQHpn3jlN8n5teyH9LQ0EpPO9TdgEifNOJ/hn3T918+tw/
swJ5Sf5xmPaqT5A2t6Jw0XdCIkUxLkCITia7Cmi4DTIGT21o4F50zzk6Ce/WUorr
vzhcXmZLvelWo9o68ZBMk4e/g/tQA1nYqgb+caZ3fUiknUvkPi9SwBOmYaZbYhEs
96TTK+YaPHfxmZMksjGs84N8NbOl/7j91LLdBxfMvqXFTFoOgsrWcfsxMpHn9rrK
wue6yGsgp99C+jhGIBqCq1c3tIFrXbwbJlIdQTNRgoATj3q7B0wjsym+LSmI72QP
sVvx99Oy5MOPMdsIjfiobTyoXrAZpwa+Sl8/jZq1mjobGTpI22mtH5Jlu+XujxF6
H60uayWBjyUM5tXjlCk2+3tE6FrI5lvVGBfWR96Be72Bxcykww9N+DrxCsEdLH/V
bDaO5ipIIjaarSOvrarUJpfGW09kOk8LkX2MuDYS7D1F8lnOk8S+2FhHqc2DbUtU
rF5bCz1GrlcZ9pPuGzNkdlIsYZ0y7E2UpQJFssOAG8E7u342DIbjY7CbPTJdIJ78
/qVVcFqc9fZ7JBkdKGSfHEqPwDV2qa5vE38FM/J8NqkFW2b3goMRJ7CaF5mOpg3o
uOdkwECFYeseK1P4wIdJTno4TwHG0UT1QDCfYV/g6rzb9ygexE5mqrR0U/SzAKTX
asgVTVwA57Bm+srxjlSmSSFIuPBn/an8ob76N9UG1slz2SVukKJcBtpLYmm2DBCx
HiUYXXfMmzj2L2afujr4i5CkPuTG2nOUXdObrtKmALvq1vuCsN6vT+kU4+xZMTfV
JSvA0lNFiYvFkix0VYi26sPkUjSCw6NBwsY3WdBRszfkyT5MZ4ALf0XWdg3QzRuY
VgcteKJl331YZ74fsOttwiBLcgMp/r248O7pJvu1uv+kn9NM6bYgV19n4SYeA722
jmr4cNWwzftAAr3OkaCpgdyvz0yNkK41ttPgDLCDWSjZ7ez+U04XqwnortJRQVx4
zZXRuhf/Q8xeaF4MrCWOuc2sBMT2T0dSCi8LVr0wS39LkSSdF3msAnO7fynvdMro
l2KiNFhd+h2wUwAGPPdQBW/R0MbQMKs1pP6vhy0FOfX1yOT7YTPV2sDW5r2qhrZV
holgiFM3wgVdU7cdAecIQSnBGA6O4iKtHAtA2MbtCAdmTOpGsPFWCO7E+P+ul6j5
Ucs60AltUYCbimjvrgXDzDOZCOooNhcyGRXDcr8ccH4XkQEPAt2++sH94UvPuzsP
Qeqv/AAATMGPtcV0X9ESRUbdBr6LHmYiVGKwNrHy5jTmN81Qj+I6XXLJtyhO5uWY
E7BTW7VIddkW/Tmq1Zm0XoXU9uEnNwM9iLlGunbr+2moXFVMngmqAEmGVKjn7wfj
TWGWkh4Is03tHSEyFxts+DFx+b/eMpDwM3ovW/3qPqB78NPjIqcRrZ6zxJ2OdB+1
s5Pfx2kdw9diUHUH1iFpNeZfBVcE409kBC9gknZUslw3Zw2Jnqq/kRo+uYCo4xLh
ypspOxA+E4m2JFQj0PVXRiIKhxhOCRX4MLDpIrKQ1mBc6DKemRkYqNbcaNmCLiy+
84+n+tLwRXUMaZuvJaUQn9YLmwUMU/NWGAWJ5BJGB5XSRScAVzTI+kRGaZk8EtP3
nhaREWvn6Q0rAl6Vx9IH19ENqTO6LWQ+cAs0UncYlesnChsqEAMkak43wiKfDIdS
6NbxK1NBE9Rgti7vASW9y4Nns3G1vmI1Z3qfXfAtgtLNohQjBP8663jZljJhrNTH
1OiNvOCFMZqsEeP9os2wvBHmazTdbBOQJU+29sxzmgnIKlIT8GKZ06gjJMTl6WfA
5oKgE1ODtoNITZJAXQ5/0l7KUFy8wokDWv6O/9mASYFxmvll5Bgvj78oebKLH3Ns
bWNXdxpCdV6YY9SIwz88T+4FSZqm6w/XWIcKPnhHQQ30qp1yDncOo23tYys4mZOA
ySV+D6yMYxZyDmQ+KhEg619aidXoak97ury0amS+nqTQNtWROCwc8lVVaUf2X/yt
Ml9iZ2MfFrSkKkPxOJHZMtIufxRwXl985kH+LccEY8SgoMiY1cUP8l2nmRJ0iXxS
I0wmmtlugZCR9cHlt+UYpUwbp1wGBxb/P/8ecy061owdWMSQ6GoGGyXvaWfuZCPS
8Rqx4cu2JIb0pfm2LteyUDUw1vD7ejeWd3QppUNFifWLRz/JfaPpr//b8MDqh2Ga
jAxcEKWXauObO2+D3YGyiqB1JSIMX1aWnHxtdHcceGs0OZIG1B2Sfma/L+bQB5p1
wnxGmbl8SVw06FbyPbFI3M1G3cGhV2iXOf8MKTg2hkp6Z4YmEUPwSV5bVATswYDv
+lhpXLxgooX7xs8arojjD7siLh4+qIfSEPH3YfFGum8I+5GIXMNKU+DpG0lwpl4I
bOjqVsS0nNv9ScnBsHTMvfcbtOH8sGvpDM0K+WN9aeNQknyzjwzKj9YfprGo38xq
iWPC78paYYCpuGm86A0091tYwFPs94tGlNPDbAnELEvxplzFLowvBIo9ZzfnK+O5
mwGl8395YWq3PgXtPYlOLxPNkOI+qG5LUy7ATImLuHkRExOogjuLLm6TGAzhAokx
WYxt0UH/0m44r+gB9NXqVMVKZdbetE//cWAbWpcpWSZW8Dcq6kdTdA6XBswT6zm4
iHbta60YG05LhmmCg50sAkK2mNthcWHioZZ3xdgC76GuL2K/sD6s3EhxD2S6yv40
NYozoc7vKncOjhYryeVIlXyVONRSL2F1jRVfGEdTyV1zclacNJ999lvfnBI2PABZ
WLzclF71n7HTeofR3ynYdaSAWj9ZUwJJi11LDvyEAWrgXJF3dgLDSUmbbrrP4Vle
Au2x1u8DZvUDGzmVs4uyI9Jp64rlxb+PXvodz3wXyG1xes+L7Cr8MVTE4VPNN6kb
T/qObBa1fXNd4tmgl/oBWvgF5mBkKoB2NTi3q965r09AuBV9BgkcOEdfRzz3aniR
6FRU+VmqdfP4Zb028DHKRJ2UyHt8WgwRTzHHw+mrUuMHVcoMEbSU13jO/GhDx5fc
ScZP96V6cNP9cEr8mUv4n6c0yIs1QYZC6jyr0ERHSGOMitnls0BtqsUgNX/jTCyw
lAWk7PRbq0ZS6huGE6Xw1IKpD9Qzn0s3ANwqlchpuE7RWAnu0+wE46aHiJ/hVcjW
PfS8nM3afH4Dr3vt/uuXCMZ40wCM9LflYhrmSdg8ScxXOM05k5jkHUO0IWS1vS5Q
9yJxsAWNIJgK4XODxH329GmpQKqndmDoFFOMdYbICTNWXa44NKzNLnvTochDTDKR
OMfTScxIsjM8n8MlNRf4VSX4cJq6IsDXVL7pKUTAgnhvimV6OVhwrdoWZiMRR1rd
5ASGmKCqmM38uuS7V29fvFeVTgiPZ6XODgKEFL2LnNPkwpLoO5q3MNiIvRUl/Uwp
dtzaN6YTN9wv+zIwbTgCG+sWe3XmQYBAazyUPA62fLNpBn+7mZW/rWU8tGALJehU
QJIpwgLoQxm/n4GeMduVFK5RjcuGLYH9FIb0Xz/V5C8l08POLhbSpW2pqybtGVp5
eYe0u6s90PfvkJwllgJxS3Vxr7DOBQ+YxH9Joqxl3QS1KO6x0XC4heHRZG5egRBR
QjAn2FgvLR39THXI0r/E0MSL+v5/RRTVWWmupLeg34RnmFbIuGEXaiFExwB4oxYH
ca4vPqnenIhMevhX419AB8nshyzpc6F7wTNqNErx2q7fuyCUeJLIqnx6lxgfvWWQ
aIPVJiFqugxLvYl5LgE8uBHZ13MuPuUzhmeav64TNi4r2hLEzY5cm8qsfPalqR3B
9vKN0JxsDyiHSJqbOsSbGo/cIRSUpKS384JU9Kl5fC9Nf3aKgBGp0FOTZ0FPBj2z
w+bLPeW3+Az28nXQ5P4EwIKOgMjbbIVZf3NE6cfG719S1vDkgIur2iKePMVbMZGa
5KAJ4TLfj6zw69hchW8/n18rmJnnby0M7xc73gHl6DCoCD3LywWaNWXP9X6dg4QG
dtfYkTRIHKTJWUf63GeIisU8uJv6+yADjZRGhjpK+Q7qkifwQIB3SoYOQgWDppEy
pIgdHmermbpulR2UQJTy7O9TM1+ONd9rMfZcQHd2yIuA0a2zzJjwJPx5zcAgd0dE
kYqWdRcEITxykr0ao5yS4IQ3sRASgIysXIihGL5tv8VcfiN7D+qLZJYiFSSsdgKD
QfxYJ1qtcAepWQboTx6qDjXnqviuotj0R4bkp0LUiNYD5x8cV1fALKHmysJ7sYAZ
cw7V0ZYkP+PY2pnrCNo3blOuMEkD5e4vpybHc1fiRBA22OFo4q9gfSiXXkWKGKT+
SGSGjOERS2bcb7bsCRSOvnJZafvM/idp/wpIOclCr8X4fzc0Ug9ooS1Aqt1gJ0JB
dot3eWSAAW2ZI34Mz0tnjZKYcOagrgbVz39JuLF60O7Wz8y8efXV5LWwi00Ol2XP
TCgpNAS6q8KQA/Hv3Gw+Nm6o/DAMKdm7835YTqdymeVbkuoasdNpRmlqxF52WvAy
Llnf5dVuWiHlluucbX4/7iHCGMJlT7OcLYf0SHYAwaPphVfO1GNfjJFAXEEHD0XU
R2HB3aicfr7Uktp82wYZnFaS5zeML+5xfymvJUHYbGDXELFeMZJb+qgop68oydUL
YhMBOCjd+Vh8t4GxV+sM9sDelY8Bw/BBqqjG7/rp+ApSsD3+XtywGOXRS4a3K5Rs
PLl2ziO9AU7/42mxZFf1HpQkOzMoxYxj8nowzeJ2KOqMLlX0N393EN9LB4BUSi11
JIuvW5lw9W1W99R0GmMWkSRZpARDU+3ATJlzyxYX11huWjA1Q5haSgYVEPI2elw0
heN0dMPO4B8/XrNBf61OB9W6v1mSrBMS3uX/DVSIpzvmrSh5QksPyc+I0uRleGqb
Ht4NOf2OOgfaLiD8RdF+hna2ZjPSrZFdQ0aezNZLOshIZHGix9RDARkNFESAjUEE
qs6EENZHVJp42TdNT6RI+dIlee/8WiidYwKJoG7Zof8YqvpHe4Gk2IC2HKcUUzNY
lqpsrG/Y1W37pDcMjk4w/ZdscSpDPUwiMM0vrUd1/FqW/lxZUhwz6Eyj3FLPZ2xF
hIBkgQxAezvq05IbTmuho/g4VqgASNuIp5tTIZmcFczHBBW/bgs43SV9Np9v77db
FXI0poQS4D18OGurD0Ho5pV0OI21XHxR92j3/6ESpjkeRAfEAC/cjrNYEohECJzb
cLGO+CSSZYBffIRAcvu5EMSJVt/rV+71ubac905cxEbaInD3P2cN5IJjXEoR3JOe
toPDQ2m1sKk/UOYIzOwezcjPvU/bEDS459J6KGT0og7e29h5B8jD/6rBYZkmV+JF
Gmqk6v4nsPEqDBq805fjGEzNzIj1/IaUA1d2qb0r9sKxKZJ+fuioZi4Rat8aBD9j
dLmMebA9Y5rMu8BA/zR65G+gDA0V25dMLKkUW1RQs+DUrS91gmZaGh8R078MpQ06
tvWjuo03S4IaCV6mdWXXJ+Aam3Zk4luAXtS0zWbycH8SEIV5HXslNriGGKoR7i7c
QdpAkwwG7nHbhJxcD4qhU5rIT1pJvLHwrd6ljBe0t85j8/OI01JpTDbqKos11ITc
UlopedaaJk6FR5di0HH32HE1+H98c5+qg22Ye0DsfWiBsxIm0FJIxnrbzrVMyHnI
UJwOkqUZ7np3ZynkkAJAFJGDx0vUSkAnXreFvjGpv3i6CXa3sBa8ZuF1WJYASZ0P
zEfRLo5+1FETKXWw4qUHJFvyOgiSUCxVKram6io2o9sj9kWnjpULmYT+lAdIslqW
Y5gK5hY1rr7Fn3Dbxe41D94vkLuAnHEfNyWuB/wD/VIrHgMHtpGB8qYE0cP017h+
jjy01TcTzJZSPzdoouF4HoX+NX4SVUcQsk4UwHCBCD/C4v4MRre008NZrVuz5oJA
3X27Zxq6CfLFlUvIbtz3uuXDS6DNNbSX3cbYworgnlPui4RsL2VCk4NhIhfIHD6J
4Ld8yjvkwnlJ6w3vIAsKuGSKFq0LZ7CYsncvinDOlnS/cMdZZK1/NQnjAvUFjuwU
WRnd9J2+4W+eM3OGaJcSTMpNckSwAb/CITfvslrfDPHbq7NZe3chI8fPf6UqLQdi
s4MbjrnhVliUUJcZawCQjbu7kywiKuEmVn1wxuC542oFA7QDRLjCaeHaiUHd+sXJ
Fzitjq3qgKf5t4StY5qosEkNdN5q6XkEIxz8kq/2dAp3mDAPhcxRzzhCZBGSIicn
r7Y1Z1rv9VmJ4q3xMxP6Ujuo3PinsxH50tR22KUzAp4TU2D4g5tanZP0Sg996xVg
ldF5fCQbsZdkpXp65RZ4g5h2gn5Bio433ZuM62MLJQKOi9cQSOhZRVQavrL8WeX1
fNz035CZW041CDQ/9rCNW6X/k1SqSWnT5TZ+GT2HRAY9LgmX6u/EyNlR6kzHMl+n
K8moqSd7iQOwbNE4DQ21xUuw8UMEpqaMGMDbKzhGtzblW95h2ADFSY/g43G+Balb
Hm/IGKvDEYDwO2bbFV4USBCPJfAMneFVZwCbzf/AKUTnxXbcTpuE5gxeMZFLcx2G
qhdRoIczwAwY+zzCoDY528ntiHRoZLEwIW1CXk5oTVIuhJXRSxDYy1B35DUS/bFs
TOo2BxlIpoE/KhmYLoAiPF6zwCJjqAqayFe0bqfJK1LKi+XDnENHy5ilaHiMur8R
e88db3en7DjR4nIkIGPqT2MpLRx8j5dyIe0GdxpYqu1S90kak4thuJYg02hvez7q
5e8al9HtDpTz2/nlDkFqwbzp5438rR/u8T71MaXCX789O4HCvaqfQCzSltmVUE5+
RmcIpGWqngDRnOrAh24aFfaDXZ84vttP6a6LqGzWVOdUTnwKFXwsPZzUnhPC/y8m
C4FTqu7WEDcB2aUnSpUDVQgkZUYdaPbRkxqIa8l9/JwWWQ6tv5Ql/+Ey32upDm2o
4cFC3WVadIbSux6VY2qdtfaqalG5BWJwYb5Urj9L/oJpAdp5DV1Aggy2qeaLg1vQ
GLpgNU95zL2xZUguGw+JfD29SEam10MrhMLl1qdFszq/qV9j3hEBnlzY5ju3vFKD
knK1UliomZm8ijGJJyoEeccX/fSe4Khz78ivJcfkWkLulx6ICs/YERZeU8fS7Geb
SDlxMejT0QE0T9+yTRyE72DI66GgQBpzhxHUlIoxxn9T8kK8h/R7tlHurZUz/vhF
A+j4OYEnFGdObqoFcrWtF8ia8cSm3oqzGKrDkmEBpbCytCqs4f6vnr6gpEaVQ/a6
vYE0yEKdknmBAK0xI7PoCCkSbLx1V0g8xnH82OmloUmh7vEDAvn0/4iKEyZawntq
bWDhqYRX5VFJD8OUnGadhhDtgtU8p8bajA3zlg+/f85vK0XknzFQBCvBZ+GpH1By
tjvxKgSnaQRV7nUIFDpvGXRPvbGqgwThy55KT4wd9FCmetIevrN3BycJMaQOZPPD
k98CJqu1x7S3qAowwf5CRZMQMnFqk+A416PRH8Ant9kc/po5o9pnvJ5NpTjvk5GU
HglbYiXe/Ihi1LovWTgfYQcHmt1sUrIervOAO4w+OKmB5mjFhUcYSwxKamk2yQTd
RYlix/+Pnxn+4I0S1tDITxRhekkPbbA7BsAJKDbFn3cHzsw3opEv9OBygmZYMjf8
uKRpuU4CkYVJdoEBlKqamIdMFcnxnMoINkIivPVhRu9fdJ9hcS46DAtAPL/HXtV4
XoK8+oOPC7H/woYqOsQ5jvsyYOzkH+EUo5lABWxtnk0wqUpCu1XVkIb+1o+RrqRG
nAnlDXquaWv8I8ZqoDSuCui/FgUMjx57+Fo7fHIpa/y4TAlnd6wd3liCYkipxWaX
kxAHhAu2Sl4vRzmqtcKvYnKo+R8t9vkd9kAfAVxe+XkvLPzPPiTXjtI7qZxfwZa7
LDx63u5vCqXqsvPAxWDR7mDxRmExKFxubpU0wUZzpBB/HEQhDXI2s9lsW8n/aBsR
iRgjTzGneIzlGa0E7DpzBe1m6mljBH/7ptvqEoDp28ueMN8MLyxSFhe8hSc1ckeb
H7Ga1wZuNnzN1zCC512nI+WpS/qT7M5NxvQLi3OAE02xrZlqLJQy9LWTZ1vC4oqM
vyxEK+jP8GTPEPNhxjkj/c/bH/wKoWZTpXlzvU0pbppYOFy89l6xyKMxj3ywLW74
gQNV+WMuX6kEwT3DMT0gB/5NQ0prGJZsh4oHXJugOCxJr5lIdzeddcbrGkcM2Y2C
/7R6MuZFRkSjgclJspS1uWyst3XKELyOJ1rXFotkORxltBk558zY0F/ukR8oF/fH
UZEr1IWv5DvdZVMQGjueMhLTK0Dkp0tKzY20q5Upj9eFao1sMSUAb2WIi3xbOCOC
TATuMd6jbRyjXLA+i2SzvsN4EP62e4PRltYvytGeoEy6WDHe9cwFimfMLnYIbn7A
jfAdOo1+t5wMqWWFZPyJVpH8FNo+zYYbXrQy7o+aSeaGZdeguTajcsRlKVBwRmxH
/oNsF4v/KZQ4Vfsd744tQwYMQWo06cQ0AKXqtIYhEOvGGWZBwfPD6RYOAJrhF72c
O8s6rAFO1ZvFpWNnBaYrdqZtXEP/GY5wGQjj4JAI7YBGCmtUREeGnez/6g5BAfCx
9K306H4hqUxnTMmRPqJWumtJo9ShLYTBUz18QQzjBRUWGA/tW7bI2jRXwwwlOWK7
/Xm9zIE86E9uAs8tXMLK/VtZWqojNPrLAJOscNLQLJ7T2cEEsLfOtLr0ytkrhg/k
wYpTz9HeepK1jaCipS7OJMILb3j6I3TPCdqwy/NYbZjHeEaYPz8/QHTq2ESCwkAO
S7ozrgkn+wSUkyQltZom1AnS1G+6miQ7uwb0jCAvIyL2RnaOuTvoCKBzUYeCdQuV
2mRn1ZnT41Fjzx4WTnZI+Oy6d9gGjyiapfIh9G5wFZQLCRBgfH3prhXNSUvypA39
KNEHKAmf52A5Smdhjcx0rhpEyRGe3kkHAx4+NvQjN0VQRgCQLFFoRZVrbtZ5sZ9X
iNCXH2/jUFa36V6O7LUC1lRDd0+R6Fy25bRta0DdDva8At7EzFXH3UsVaL5/fUPL
gIC3C4CroOgAmgC2L9Rfw3ZYIF4YFOysTv8yMYBAw6WG8D+SkajFwd+kZFZI9Rba
hkFM7eBTwBs1mGoRXGAiqiYbKYrwwaB7CvU2ZzeRyXcCA5JGAqiTLmmGeBEjLcnl
US4pY1RVLts9MY9MaEJLE6Aodeq4kt7KFgrgwrVg/zVgA2rdU/EpJlUO8fjSe2mv
hFSDtEiP2jvNvdyGMeKwEeR82fWokuDTySc+66qV7OoK1nOUH01ilBt4ChRlTV31
uvhVD0RfvDTf/z8ifr35DaiCduCdpF2ks2KPPGqDvyCQ0r1NErnTUDElncBx+Fw5
ucaO+/RTMeKJ/t/IESde7WZGCkn6HoCr8wNlT6fHcxotKvxzvdDRV2GvHqZAbOva
kNC3ZD9JvhStG+edlWJ+lEvWJnqU5T/ctG0H7oxVQ64vTlYiqXRzzrR6RcdSpXdr
FxOVkw18NjPFVBnE5dw27gfFJ25EZT6+4bq00SdUWnCyPTWUttzlDxls+8OrkXXy
n80h0xus8Af3SvF4QTNV09+2c8RR6Yb4toLdp5YRYCiPbfGO4rfyzr8Pku5jdaDh
FM2CXEP+ItF2+g3F7ae++8SAsBHeJdwhBZMINuaBYldDphb9cLgD3l0zVJKL9FKU
767f3BACizG2irmyjXAEOD7IdnjSLk/us0vAQq4aqemYciJznPZqTupvSbWfUt6D
Azo7KBPl5wrXre/K5Q+WSLOwa6jT0q2/YANbK5m60KRXE21MyY/kTVDICs9svAG6
KRuyXsY/g8XizSBA1o4hz5+F4LJv4X3JHt3XHW0Iam5Z+ZBcapEDHI+alJVPlTbC
4HZpus0Ld1KRMDtsD2e6koK5SseNInMla10yjtrBILqqQLuDW+fpLrnRhR8/wT9Q
56TwUUeNXCnKC7oyUjVWB1Sffb5fn7WL/S16QG1ShxVZc6+nQ0FDRAZ7w34I88P3
g3QaeMQZSbP++MasJ0/hraBcAKL5xcnp4ZGvD1n1pK8+52C3bKZE6yq2nEuuhDxP
BHY6UgkWSj0S9hVri4uVR7dZHpUmzGgaaTD24NaQaQIOqmbIDNKS4eNy7VCd0Nn1
wCAl9qQ4j1T9DD5okbaIHtkGRTIKlr/Wup1NFZEedGWiUO32cADS+D8fwY0AtA0S
nZIHBbq6B2rdAyYOpHT1VH2CO83+1j2ury9T4ZMvdb033atK7+Lp48USvU3U8ZqU
dIih7uFTmO2Q/GUMCBaLcOqcdJBd7KgJNmxL7zOyKcynPsg4PQTWbh/l2f6LcFHl
HDjbmPF5y2hd+BgzPplH+uXtYUdj9iaEJ1wWoruo7F+VXKHKdTGaBrNHl8yfwFDP
JkNfeQ1Hkw9K/trEP5gBhjFy3voSmR04MCTupf42zOEQjIrgJ5rxj/1ZRF6gCJNV
7NfVIvoAaESlLBPRpZjqIFcvmKWft02sMoC/28gnktc1Ap2uMSssroIid424kHWX
0HQYzTSurd84tZvSILQFDtbSLWYAAnB0jUK2ctR3cCodErBXtGeKNwyVslGeArn1
4Bs+r0VnDp99s5GEhJP+4FH7Yc9V8+pGqCotUBiEZo+42tFi9Tdfr8n9tuomPZ0B
m/4loASGLs8h3HKRnlTZaF2OZ52eAx2MbS2pwT/mRdKXY1Jt7oF2BWD8045MFzEz
KxMvzN4pPfGbH4TsZRWuFmup+jIsuVuJ13dW6xMvmWNpjuxqV7ww02d/Nk2nbkNk
Bs9bUKgMhzbFdBeRGldcLAjCeAwDzrOGbxhVC0j4WVmm3ElTBzRt9BDhtgp63uow
wO43IeJWOKQfdOEMtZRbuITikaLh/0XayJxH88pkDYm9I9L1TqqkrQd/rqQdlHnl
RvIys3Mxb3vn5ma0vd5ITGK8IZzOyq5JLV66MPt1fiG7nWaPB7osVjB4FesYFzFy
lg3vENTNbrm8A/AkMfzo/WCsDc4IEmA8bgXtkGKtV06d82HUnU21LE11Vh9WFw1o
KNfDx6AILPqt3G+AR74f1zIgia0eeagI8Bh/PMVjOu4vgUZZPK6+FVRVW4kgW13a
4RVceZNy5SAvOpGO8hsjLOIqmc8Xbbm0jMm1HRzKTaK+sUAg6yl3vrP31VgVHHt2
yqC32jLbT8UUTbrIePMws43Y7rFDiWZDvRiTl5/ukes7FvhQEmvAZbNnhD3uXqqI
+CrxOgJTVBcUCwpWa3BDke5fruge36JLz7+YhBNMfEE1nYBU4DoODMw7O+UJhQWk
tEHUhcJc2aYKLyCdd0Nfgkay4Xqcxkb+b7DAx5HHgjN4pe4QP1HVaQCfjBbBfBxS
NNKMAZwV1LbyHefEGcbpWLSDuMeaYrC8I1bRrzJyJWINs9qRr4+4edwmxg8tlNIk
XOcUUID7fAceL1SLHCllRdDsc0YsackTNoSUTfGPdcwCb3SxnSkUxVu3N3b1jHsY
cghFFj3XtU5ev2VDRlXqH9bQvGmJVfg4j8QrfmD0kPvtyPai3pzoWE6ntkdiLYdQ
gfNLJrXxdV+bEg7uGQG9UHCWkZ5NkH42Ap+W8ZyPX3MP9pVrh3n+Wxzuy2lcYZud
uJHSuWXQXfmgK7ybTgcj5QUcFR7ZpGopMGIdx32/7iNmjzolmb+2GU1+M297zrf2
IbFsBA2mv6k5RjhoQUnLdxLdWTY4VSGV6yAq69gp2mcBcdkmb7mpoO4b0bPIxhFF
jpd0wXZmJnc0TyBbQLz9IaeFsyUd1yHMGtaxzBE0a/RX7vF4T1rORxxqqW4ivX5G
z3G02M+SKk4l27sc2jBmyj37OvSFRCgHs5dEWjxkFqPTsz6BTODAX8MbWTDuMQuR
8s70OcpWniC8Zy+lvcd2+qYpXtmc6RfMoSH06sRLzgRjHFpG0cRMD0bHT1uf5H3h
ckUafL8//wR30zv3veb8QN6l+uAWzXZQnisQMYvYvlW/sXGbIWLDgtAq1rDuA+Ov
yk7DDyjcjMdr1SmCq6TYYxFEpRDT4CDhbgqlgNnHWH5eGEHyFwxtKDPQDrc3qAuD
om75MoOXux6iZI6eaKayq1hcDqE0DsUHJ1g2t1Xr2xGF3QDFumYjbdpVviKl3mO8
kqsmY1jY2gSW9aOHI6I883KrR+Hy0X8Bf116LcVmEj65YCjoW5Xp17Edw8FK4HNm
rdvggO+yVj9s62oufjjTItC8CwAUFYaoTrqAKm4GXHxxRpss4Howz8AK7NvtvLQg
lsWyqYxCljxijycYwZ2JDT/GEzZfVkUBwLNkOFGUeTaAnLEa2mghMvhpTPsYhLwU
qK19Rv0+muCiZEp5Kp1RvTV1ZHqOYx8MzCEfcyPkRlitT7mY+Ti/FAFnzxELghro
eEFhMzf2GLm/dqThkMBcWJFm/Uj3jXKkKIt8muUsoclILIWk8pRQnXyyetOjgovQ
RZaN+HZJsXK4hL3zNUccHm/6MyapU6UaBdi/qWGZ/gI8/hEnerjMrVdztuA4sUbT
03vR5tkGHA1ff7BAUK20cCy0aEx8Mun4O04LtxWzfTShSEsH/b7TI1xu9K1HJfKH
xJz79lQWVWuXuf91d/faU7qH9x5X+H4CBSYX1/L8QtJl0Mb48Q+MV3lKAqqHLROV
H1TZcB0g6Wjk8CeGJ4YBC6/jv/eNMECi3d3YNGYkLyLiLIAhu4yaWo+Q2coTD691
uF2261inCr9/DSUZQkVxn5BDNyE6v1AfRXXV/P9d2ctdwEfYjYKps+Y0yJQdx2ui
k5TF1IsrLLVynQm4NrMZlCnESBjsScp+7INB7zejew04HQ4ZIvUfwvElB+oOCQg9
SEp0y+0nn1rUhTfRCBtOiQeGZPThGvNYajeFYyYKz1EMZIuzv2/5jtoSfwICrzz2
jnfpalXeGDLfx63AigL4ueSe5TvHjVKGyeoZOiThxMvLbWKazukbBioPxDnmFDPK
ZmrgNSdE2VduRE3gPg504XEV4HyTAHDY1xx4+3+wGj/Hbj/Awhn4XlO6K6Gmw4+X
eNGTAMvbqLMfTd/OZjsoD2sAL5gzx1fz2pxoNyUgfmSTlQWiOkU3kkiyI4K/m+vO
AzKyZMk0x4Zw1cqNVS3cuO9KokpjCnfNtb0yuTN6aj5jF0YtXizwPoDzPjI3CIGk
MZjW4Hj8fUaZTLqsLioWNaGcM3m0WKX2ivFB4oeHp8r9w+lPBpRH4oNc7ZdUmSfG
JJ2WE5ITx1q4YeyWEanRHqf79QOpzewnY9HIOv8K/FYshoY75mANahGQOyt3D3Lm
So+x3jXspO+SRJcmLiZJWOT0dLEV8haIqYSIIn66fhQz0MWlI2YpZhRIsUaupQX+
olR+5jsmG93fq0YqYLwKb3ySenkhnL+clzaeW1O7obxq7H8ttJdV3vl5lYb301Lz
ll8CSKRcQwu7LktgZNZUo0uxy8vUPzG7DQFWvfGBlroVdYSnBQdGTvCTeD/JmN4L
+AsJdfmixr2dR5pxrlttyBDrOOli+GHNMwI0kLupOLg5U3owYhwQODEm0KRUKpFy
kr5Vp96SoCg7qfW+5FPLd8Ja/iunSDurr5+tsCKl2jmDts51yCJA4Vd86vuIQF14
ecy4ZRisMJeKdNLBzSbD1dswBrN/1pbo46QB/urzd493yzBq+S3hmYtr/hjaazHT
ghBfp4zp78SxJNlHRck60o4KgDl5Zhywt+L/6kY75GUClgxwsb9zxWUVi1BH2H0i
5qQiVWNzwOFSAbcaFG5mojB8K5+QIHV+uenoXknm8VmOSJ+ZqD/Zr4LlBx+ytdI9
0F8MWCYsAmsCZl5YszfO8WMYJettdFyODr3SHBbNrtVnDNyOkrKD/mjC6z5V4Eq2
pmFreWFT6Pf5S3D+Qm1a8BAjaf3jF6wRc1u3ayTlbb/xdV3Ze6U4uH9kgx1SLpzV
q1Y8iGS05JDuowK363GtDBNp2XQcKcEKuedgaQPQQCAC8RoVlojmjeYIVHAVVnij
cwGQOn6m0kucwQyDh50/zHqjfBEvRGXP/NvgaD2xSHElmuDJideU6cLPUlMIiuqY
YI7OLxU8vtgz9i3aVCudul/fTG2u0syn83wmaDaGYYgy3qcwBxyL+PkH51PK5/oo
sadBx8PmLrLuwm1q1fpqQZUmXOPoRkUmEQb9yr7d0jGDUICCr07Gj3HM1DJoJ+8x
luQfW8BSNmsb5IeXpc6CsN07BmVHpt6QErTPRvzKUR8GH0CcNzro7+1gemQNjRy1
UtOdsQgjlxCPfyxr4BFNPtKJAx92xY9Fvmp354v61+CV63qUsgzH7W1CCa+nX4A4
8TKQF8B9c25I4ThkVFm7qj7zmCP8WBMAyYCN1D0ei6LglgiGJ5ywSEf2t8brqyJW
d0DHgSI1MJgmOWLy+NZJf8KhucKqgAPXh5heioV9VAy5dreDKY8oxVr4odblQ6E6
F+angcmkrGgzPOMjWeXIoALy3M0Ao+JNP7Z/hR5LqCwvH2m+VMbbDraM794cBqUW
P6aTPcc70Jk45Q3C5q+zEmUDxmy3H0w4KyvSSmeeRAU9kWKaFRLIG6Hr3JPcdsa9
EumJmkrr/HXlKWitdnPQr3x+um5IHbNgLWx44ix+Si1S3fr3m12uz8uS1mLab/ts
I6yscG9Xfzkj0pQIvskS4yJKQBPthuBxx1YvY2VUIufq0D+3whLoIpT/Qy9hRKC3
vf+x4qJFSgfOF7+jsRI7ktuk4Rgdr5Fmj+L1RrPsTaZngqNO215i9kO4/7A/IlMz
JTW3ENrdju6440k9bgh1Ft9pc5ABzPdszc10p8ue+59F/pTQqtK/YPLIP5eITtpx
GStWoK8Qs7AzqchlH+vvnzwcy+cdnTPZQm0aV1m1l1Bule50No/E54f7M0QK6fbV
AfNwY1UaBwVu75NkgB+V359EVSvAkVG8g9WGScRUTfmHi6l6SWHRv9T7TewpW/BD
+Z74wQ+1vhZwmD9JxgQE5gGQ4YNFIUZoqeGzcJtjy0E1lTbDiOzd77E6Igv85Plt
9/ZjNSdDYh1H28pJ5ha4pdWoN4aA59KKF/3jWm5SxwVkpvENnx/uxjAtRS0zQR4f
txNAlGQGtPu9Z0OK0y/3/7kMbNjViWZjkGFN9MWUT1IejNCULOhSp5VtxYpMQz8b
/nnMq2l5AGyz5qRvkwYpXvpcgSyvkg5JrOVr4Gy+TVSGX1lVOC8Iw9kTAeb91rDW
kUAby2gN6ufxo5xXAWct8ePne2ddD3eS6FRF6qm0M5G517kgbg3vkWoznJwsI+mC
jo+0Y0myhxftMIsDMVdVTIMdyzbPBAJl4W95tnuGKzblt+zNzNJougdAPT5to+GK
2tSAUzFuyjAsO9ebitNd/KaSTs7Y9dRtWH82eMxmdNgDBy0m2qy/AmfwbGg/hUuH
KPbeqInz/r+uakGn14s0ZnPHa6Id3ZZ5+aHs0MJ06Dp0SCBc9Ge3aS6fPlIGUg4X
JEp3l51TvV1XSYNleRfplFrZkb7AQorJm9OIlsjKr3egkDhNpNzRGo9FJaUQ7bSN
1++aUyRXeS21bV3pG9yvARyqHXv0Pa7uib4Uq3OBHXFOTkClSaH47bDFWN+mGwRp
2gD2Op35M+7DC0BM9h2W4HKOR/98c0X5+NN9uhrccJLis6IjXiB1iyUetjM+zMMx
OoMwNn7C/SdAifPzqcQtci7atZDA8RuQGWr3nxauaV/XcOs5BHgZAe2Nc3oPJ6+H
GF1bYw5zMHYdRD9yeA0MppCVZS/IQqy3HdpiKlVI7pQm/gOOgeIIfKq9LKw/lMAO
oSkx9OKpJf5TApQwZAc7/4N0sz82dhYCxhD8HM195xxDre8r1fHRHTV6TbxVSId/
FDj8ye3xqZHeLJI8/fify7P4BYGxZDbmp7edQthK0LE5YbfJD7RdTuR3/Ayv7WP1
q34PtFkevp5AmjOpBOAtvM9VQcj8nth9fgMoLyvty9HZNSiQOTKMF0vt44/2rdrP
cVgAlSistCysD1p+1E/l3EVx12GuQkZvZQSu2aA8hqzJXzAxhBPI4DbEi+se9KFK
zJAwhPcBbW4NJeKhgchjmGamFqZVZfVc8yTBzm3mLfwIpO6/ZPqPz8M+r5SywrQr
jI7OTAmpXK7+h/oQpX04+U3Ud52oZ6D2JUvQj6BXIfWENqOkqpkSSw/uEGlmsi3+
gP012IE/XAugZvv7OLGoABPs3NzVk++LI/OM8RYUPpxTd9KrVCqXZQBjYDZ/5N/B
Yi/VtNPkzxQ2MX4OOJ7x4ip1XQB9NO58iVuUfl3elgqammqQxO/IYEcxwSlnVtGj
Zjl5euIgFVeuBiiyJRf1FXLH2EYUg+9UATg9aiTbfvTGdtNZXJXGjuHzY34HAZ8D
cNqeLGOXh04p2McTZ00QPCiuiLTqAe0zDNV+MYkHSyYnUeb27ts0eIhRGtvgLuJm
a3ejuZZmUUlmb5LYNQSDwqVrLXuT0xu6IZT30Vqio03Zr9e1y5Yi/FuQt10ltHAh
t75nL2hMexzNf9lFCc/YQAI/DFt5PKqwSM8fbWvkBE0iV0kyuHTCEswjbyyULFVf
dEJAgvHYt0c4eis3OLhjbgEJAxsVAjZdyrlpAIGbJOP0u/62Ou7ddNBGIxB2rmQA
1B7LO9CXbmzkc8HQx0oH5WPmpXxsQ2i8fv+ELeMpLlOKoEFWSHCYDtZbvnnDi9u8
iVRFIP4MtAoHhRa2dU0SV9t9ewmeDSXx5exPMjlvY7UvUygGygmBctpPprDtig/T
fqh06Lb0MQXDOZlPTaUIo/vL0f9Aofnqu99C4jiY0fq37xsZ6Yc2CW8VL1HKy01f
UiY9nJ1O8pOtHmx6HrZf0omh0mjFBlbPICpoVFJ+oQLtWOIvv/mcS8EnttbMpgXx
QgDbmlGj/vQlsAC4p1Sj+7GBvJB+d+g1OcOaz5nP+1oQCwaQYImbpIrkRLf9aK2e
FLTzCt6kmFrpxYalAMqpNwhPxh1p/vcaz5kH05M7YgTgw96Pumz3splqSVuDvMXw
ik6fuG9vqqcsbWwDf3fHh2949hE7/O5G/MGoAW1TTGz1iXEDmHrw+IKUId3Hu3TN
K64kzym2SIfHSQYpriSCGkbjv09DFeNMBuas2XF4B/H6aJ/Eq2jtZUk6bt2NX3zw
nk1oMHtQPDKQPk953nJsH3Pe37m4RGXs4eAxGHfk4Wzf7EJ6as1v/mZCcojl7PhW
4Rars5vo+jfaUeFqLZZJcmai2KHqaLKbDcscLnpFDRRtwYt4oXN71Qn00qLToMPV
CtG2LObqa1t0XpOlRyxl5/2GVwoPG19ckPnry6d5dSgY7KRogfTqj5sdPjqCo07f
Mfm05gacK2kY8vuVPBHBThA0FOPFJ9lTS2JExe4HxHTuouo2GeM46xp/X1UOwmvy
rAKwROWs4/5yQmV2wR39o7sT2lq9GegRLpA05CqTqSK8KR43yp1WIlruwtAHg8kS
I1Mgyr05nS9nnp4Kt2Y52hVENPNL1FOOIxLcuh7tbJ1HdQ080ePPhmB0UWdSMBh/
PmKhAwpyudh7j0mXJ7K7qnRz+hx+G3VeX+Oib1ZLjt25O4Qpki1D9e4M3Sxd8gMq
ZKCRFJUHec2NohlJRF8iQhkWcCyyk+sdqKsh0QUfjlTRKmKfgFeKlC3omFE+cL8n
cqCYqDQsDvWpdxuaur0XWGGAL7EGkpBY+tZwPTvnKiYjpQoD91je54Oob1HIKVfs
+U8Bv2gT+ke22FrVFuI6skRlUgb9M8eK9gFRJqhAzGvevIppfzanW/mhTmouP4hr
puVqk7+Eu5sZixAIo7VwBa3vUCM7A659EcOD/Rsu2BJdaLoPaH3Jtgcp21OQhrFm
TcXPJ6ZgYa04CHF5wQ7PhH3H8X95TvckZoU5jbINbpgKCKrfVZM330IPYJEq0r3s
ZHtW8IkAbGTwfOwrtBeuxTlvpA/3fAC59ItoF2hfmVKDsGXGQL/TcrRF1hB1YC4S
iV4zVIcNTdPa2Gb7Vr1WSaudxvVjGFfFYWzN6Zr6mh3U2hjc7dS/8g531IFPIng9
xA6b3MR8ybXp7fF2ztZ/92QrziugWxEV8KoJQ9IY5VyZcwbMzBLdJ1SiEqMV8eP/
jZsXzXOgNsuL+AoWld26E6JiPPaTreZPHoVePhJfhHbXMzi1anfrpXJNB5Nk6ybd
8/W8Vww9710VJOARfRGh6yvG9h6Gbmd3yQmqy5pNj4gd7v7kZabGh+kWt8JGOSEl
WgLMxcsiknTkh70yKEkPb52OHSK7D3NVy6Rim3h6f3j7rhoAUFf+MO/in6HVdCQf
qERkDPZ2tBDRFgO31tr3I+KQ7q++AchG/mASr+mIqDDnexwtaVMg6z2gDZHmXxZ+
jU5jt6dU/guzfafIfSspVpFBNcAoK1vqmnFLI50qWVZfRC7pg2KF0W/3su6ulQVy
b70SyrKUuG964lmJJatWRBHmMH441NYbzEHPJQaYp1w5SkZBPG3Kcx6vi1v9yF/9
L1aXmjnzZ33rbar3DAlV9tF12hyc/IqmvLJLv1ChKtxZR9/4aEh9kveMjxJ5GI8m
qHYL+4ibhZl1FGvlNJLoA4m+MQv0wXYDrjlmmfolZ8S9hXkpN9nE/WQNfLQV4oIY
yvHMFYI9bXEzhzscDenzlMDOQJNnrS0z/FUwzZjlOgejtqqvDgPAOXaXU9L2a4sL
gKPr1abD82qE9rgyczQLCebwx5hKiV0zNvxCo8cYSgglUHmtXFsFeeYFEROXeCEE
jdle07gVnXXibTRlDRFuFIaeZISGbnL7Bk3fPqPMrOIKucPZ2AKc3wuZWmtvsj7s
ZycBNpo1GZM2tBWu6pJagkwmegEqmdeZDXz25P5MaHa6fKbo3379Al2SqVNUkLKH
6UVATNprgbOvHOKDJwNHWLuYUH1SOo3WGmmHUQKOenvRyqYQgt06ekKXQmX1xvNC
CSgMHtswlmKPtU51AafRChrW68YK54OQwKrsT7kUUWIIvqXUvOUTbO5QuwjSomg0
VE9zO+7w2bxgjxHdlhpskfteNYWfxFW0qS4I9+6LhuPpEkWf1Y3waQ+dpx8FT5bg
+xTdY/pHGPZYNSpMws4S8oPRLCcU4ViGJJ+LTrLhTeVhPQAwU9pYTp+gpUmFRLsK
FqhfvRP1F4Z53jcG9CokRmLxcW3bTNxVwb6nAJaLxC1jtXNlTa1RqCz9F1zGnXWR
u+Nu+2opqjRbX+WoEmx9vZC7RHg6ByCw8FbRZeeKmpVJ0wLWszUYyQt0UxKuAk70
amdq044D7YKZTMjkrlVm7dNbUrnF0gCdtZK+OAUAgZq0P9u4ppzd0ClPnchM6XwN
7KoRbF4Zasr6FzSnFoJCC5hceYKQYbOgRrPsggJnGti0hABlGc9bBja02J/UwEAx
P+pSkmt2BmiUUs2eO7NO4F8EciY8wXb+F96gt7XXfmvNrXD5iFbuKheLCrJTdlCa
0LMnSKDA9tpPqlBaWRXmi430JDgNRy+lG6KYVzLi4sbtSiOLyxqQlqmSSQp25xnh
sod2vot33uF4LQ2Qey2axj3pK6L/D/CtBf31K6E4AYRg+JnvRIoPzwQG7joyh22l
AD7rrXrB9L2+L9AgAUwjkxliFodIWUViC6VTDGxm6uDzwarN6e7BX1jNzU/kzjds
OIuIJt4nDq5RL3p+kF/nQ3w6B3GutkrzpjUU7kNAjmW4Zpha6RL8MluVrxSoDTtI
pboS4R4ybvq0KDVwnc3VUWZK9pZO2aAlCdDGAJfpzZdKxsSBwKCbpBhUTFmdIlnQ
o2zoQmZkM8b2Cx7jf8xj/CtRqb4iSIpIp4Pohwbz0m7RTOiAzhFKdhp2QAs9CiSR
4gnjAcW6twCqxoI1twTYB7JL+vH7MvMigiE7rHxCEe8l8u7600aOVH4A2mE+BUab
liilkbO/bosdutx497bd8y8EqumCjXjIX9FCpU76LZ4MdQGwrh50T227OJKQ33rE
7CXfYMzlIu+/c4ALMfMzDBTOzbbqwUV58HxXBq1pn1ur3Gd5Nvsn3/YmozRWrAHv
iN71SS4yRMDTgcAzpk5wohZEM41kN+qSu0rGAve2IbTC7Ohs486SANSo/X5IjrmJ
z4zYBOFYqN5+GyFObvg6T//6Cbx+YtdBc5r10NrWkw3qCjqf0szY73pKxqzroMI0
IIxCkHPoNJH9ZTncVsVdXHPfNhMHejh55N7URvZKDHyGiO1CXHQAImyhIq4m619y
qHsZ4L/X6+SbQk6wHDS5aCFDFLInMHuchvel1mv0jvVN95Ei5CS+JHWFiwUDFgm2
KEJBWGRKlgLO82iQakNDlLZEEWuqMAUw/aYblwBnM6SZQ5n9sOB7p+irqVL1A774
NhEx+RPu3SAT95ZqP9Naa344mvIg2I4ED3wadNHAX2VlWdsl9feUaB4Jozt33nPG
Cul0mJ5iAnRcmHWfRHMvDg7k/h32DG9/xp7gZiveRs7E2HiB+Nl6G3f9JdTAztrD
50P9cTkpp+vQs/Ovnl93twKppkJ5tlj1CERF4sztp08RuvzjmIw2EtdOfNV7O5v8
RZwWZ0GXoXFNHkmrbI9/RxlaqynYKGUZ/PEwWfSYprP9OJe59LQFH1HBgaIhq0EG
FjQuDYwZkQoNQcQx2pYTOactStSyw8nWX9NYgJcyuOKGV3fI3OQtitTj5wh/pNzy
uo931JTHq3SMFN4EHmxkgGDedB99m5urkVzXDtvTvvY3+v192+FaKfXUu+22WpSS
0vRCSweojOY/jJJGLfBQxAek02TSpmxj8uzyAq08Sa7BeYUFIc3TmbMQ+Lr+7XcJ
aZMVZ6ZyhKhX57dix426o5ITL6ZQVTJigojeO6TqmtW/ss1yBB2gdUDcX67PaM7o
nSo19mvkPbpXkgzEuqwcpEgXxoP0uttagyGmtrLtbYTxMSMfh8Jo6r9TMJ/gmeyB
j6zSCoRyA4SZtWoVdnNgv6Kc4AbFxukA2wUufHlAd9mZBzY8gjsWhCpxt7yNgGPM
YJMxOucvk9T7CWiLivSeOWf2UjUGQ4/TiWLf2TftK/v7BijPpTLwUqo034dvF8TD
0Bue8l7EC5NH1SAwOgtm3QF6dzUgbpVpbhe1+wHY9qVLcyFrAjyabEUPCvxVQ0Iy
Ds0cRlvNltWhYnsCO3YvqgM6hu+mZ+V9C3tg+oVoR64rLG6YzN9YupSVNR/JSuUk
N5eBGRMBtG5Tg21CiqkeH+23JuhCRbfIqau7r3zAslVU6hl7Eb798dnSvM7HX3ma
SrgC/QMPqe9Cb5Kqy6F/9Fl23rClmePQ36Jk48owSookO8w38DB4k3mopt204Zbn
hdcTIJZi3VweVRn+5ubZa9rum2XrP/pNRW/8cLJ/Yt2vdtWKHyhCgIQYHkTVIJof
t09ndlucy/qCAJ/op1WBrC0szRzi9NlBWb3pLwU6GzXR0v/FKP+1W7OYXwbsCzQz
youQ3xWF5/7itFfTVE8fDSIDFb6coEFBE0yIQl1+5rp8cvs+nQqyV8fCgKP8wEy5
GvLJZvREVkLi+egZR02J4U37G4Bkx9ne/KhPVdadj3CwlUFX8F7YGfyOCO6YHDXC
KhevgX8uK2Fu1/ProAxXvo4FMaf2ZQ53UPScpEl3HygJumuFWCp7EK8cnd+Qxhu+
HTKy0Z1g01+QAXNxRgWwk5hbFzUy0o/tSnyO4lz5C5m9+OJvfoIF9PuA0A4++0rQ
vApq3LxCWeXGxdpS0cg7NUlUVUEnW66umFzLrHF15KCK2a3EPdvOgn/YTqS6heGG
riWMjw1Fh+m/AjROvl4Gptc6PXUjt5njyJbZXPkZMGHfYbfjDG/hVL2IjyGDztj6
iQen96BnU9WnNoTb5zlcPsCd9sRAogQ7EgQWWH52SGCCZVJ1jeOzkTWeZFirFVRY
gfvjtb8W6eABblNZihekC5Y6nVysyg2n0jtr4R90gHZvaYVBtYxOE8I67MLIchLY
IGHVXkfav/de1orZ9+YTpfByTQuJUBSvvQ+QYZYCdqkTo3tDb0jXkeTC99BDGN1a
36+AysXWk/TxIWr/neDrBvxnBlw72Z0XQHsXv1d2AwA3APGkF3kDvEyy1Bu405if
zv5DsB4bmAjQP7dQZapE8nX9OMVlXEULPN9Q5B2SoTHnlzSzMYJU2l+LFMYwQILd
g2Yv8MYWVlliI1ndyR323mtonAw9qqhXyDu3bEz1SA8LSLJMzDDWpaa3H7mUuOrp
l2Fz+5zBQqezL3h5Kiq4H+dJtbCWrJFvq1UNiZ6ZLWCuNVL+/E+ByLXavGpRRATV
+qPqWe/+Hl1ZSfmPNzyuOipEnlqiGXGjUAiQOYQqkOvdzeeaOGS+rq0Kwl9Ij2He
X7roe1HIMEiTfZfRBJ//KzoEOydJxTHXOFo8iXAYAlcS3I/u0D6FVf8iU32dCg6N
0tjRHWJaE0/HJE0LkX2rAdy8+tAxuHG2EORHAHNBbn7mi0GXhW37pXFMME9XRej8
fJFF7I7UMzMljkrhiSWFhPJPBq39DVTtP7XQakD6TaG3gCz2pfqF1WZ9mtTYDOh3
Ytz7FWxME0XSDDK3MkUutsgZlGAAkO8w3rtf0g3fmLYV/WRB/q74NRpfiYRTUpKP
pxLECV5lyk5spmT6JboahXUU+VUsS24LYwELBrgZlJGjr/oqfHNbXHwAUny1kedb
v9zCWxZuqvMsjl8lM+ZzDgxOLvlE/RDTqnB3FMSvblKzRZubmvfQ9B+ir/h7Avon
D7l6hcgmX2clnbhOOmNoECCb3J+eJtRUSgMtKead0mbvOUSr10frgCKv4R4xXVxf
8mZsuctPM+NClmZNbqViSoWYLF7mMaKjvnAaNSDzErSmJHRfT96GyunIUPfxWFdU
uqWGFcX8VzWVy2m5hwHcrCvoMXBODvmno1/S+4n4RXNfvk6KQWHaEfPvofgP0yIs
3GVTyx02FkSlYJNXyVXzoGKhrpqD7vP4UhrXlFAdWkJKWij6cFnzcQ95tX9i7Tpj
jIZ+b6/vFfmG0pbgwWDWb04XklpUJ99vxqwMVKcapOxic4zkP2wMXaY+owAYUuGW
G81d6UQ0qavPtqzcFS8OUGVCOtuz175z6XfkfuDWpKbzD/KhxRTZMPPzTc7WhIdi
hBHHsZj35rl69WbEoA/zFdmpSHPAPRYXdbLibkXyRNGTmzpRGbViJDbqBe+JkXCm
PctSPk1J5KT14kc0a6VA2FlluKcK7m6H4c5NRhPluK4luTYTZE4OtVhcVXRIRiR0
wmhmn6egz9atbIDJcWUIKEd71mC2QaUUXVp9s7n9PHB9rgo2htKrA8F6+9E8fd5o
5uGxeS0yUtgRLqDSzzWc8Umv8jgKW3MeKDdi0e4RimFnrqUXzJQ8s89BU8uDeKrf
syPErBSzv2QG1fNupjA71LHUdJsCQpbpAi1f8A2eQtmXFum/un++/Y7blz9uG9UU
kb+5egRepfH2D0EHmxxNc0Xb144KOVsojNohounS2qKGwvd8P+jIbPpCjCwjq9P0
acUdVWz/NXOtdDUB3W9AesbkuCWERsINHYLtdhwJ+3ki8dWE7gA26+1XwBh0yf4W
6opyO1dPkoIlYVr2UNK9veCXK2r+w+IZ0WFlfz8+nhvLHVvEAi+g9bdsReSQIMij
umPL0abh1ju/7RYuRfioHnGwF1OvN/Nb1BzsMZ7oUEwOEK5hxNOhjH4eWQpVX38R
sj7P4I57gAo+d0HJhkoqjqEs0dmxFNwExvblhYte064K38ae0YTQPfPd/9MEhU8/
JgjMDeRmIUDvV+BHTMvkORdTe40QIstuyikMwskMVI/I14pii8Pnpp/UD1VywqM+
Ivg/0/MYJeBYgI6zaR6Log5FPXzYNGGGnpzr7I5npfHAi6DLqqibEzT1xQMnpXff
ovYs6YrqBMwxLRJIUlEWJ9CLOUOEwOJQmMZPEeba1mLHq/8W3kKcr42T+v4BEGMv
Kyx0c+t7XZSQod8Wa6Oh5SuC+TvjAWzDvKzgcwB/Yt3t1USnkrxr5/caNF3rEm1z
n4RNniud/fv9gE9zybXeSZRZUv6zO3Lt9Sflk5RqyMhJl/3hGIuUF/vbXnIZ1Mrf
lYl5ewDgd4bqt9Y/A/D73Wn75NFAG90/PdgJhpEtgQno8dJx0VYNU7AHXoeEp13W
kEdnRPcd7uUYKMs6ytGP/VEvfBlmrOPTXnUA2t2c/WKpb2bBxPJ/yaW1Kp5uvOEg
NZilPnSVwjuPFl78QOA8alYnO6JPs9Emvlz31+auKZywS+VlfmiI4MbMoIfrs+KG
2TfX4I3waBTTUcbz67YfCEnQH+cnHn2OSAjHGF2iF4iTLDlRyQTSPHqHBEdzrQoy
V2NbMjFu2TnnCm8xMsUUs7Aa1FwEIEne4Wi3r46IRt5HAtAuhlGWSG8gr2PaM2OT
eQOKIFoVHHoO7sZ+Btes5Xo7B4YL5Z9ux41OesSR3ASDSxFWa4RwbwXJktnGYMDu
rUAAVdbHOkPOeO/hiZshqXO9wp86dJH/HJBvk9+N/gp/b/IgDLpuWT0XSX7PJEhG
L2xKoydbQI24T9Bco/rdzS0TXurnfKU3wxZf5SMpZ0GR7hfqVci3VjzULF5kjuve
lxhr1lXjM4nLkszUpVypzsAm9Pv4ZfC6y0OZaRkDsKXkLVFV8oOOHbVz44eu3sUh
vvLQNir96pKY24xqrboXFP3Xqyg6C8BAIq27cRo6DPGcebZvae3jmZVEhHYDvVN2
MIL10vUFeikFNNQeuvjUgcGeIqXFwayISwdrMJZX5/9cBXEh6gHcCihjNOeQXA8I
Bg8ocfHFtMydnAJ2wh/e+CRA+Rejn817SGgJ6YBOQsZnK5iFXbKSbfgj9yWhTneK
Ta7DsLPhqD8cbZ67VvHN/O7xd3dCegnQ4zhEWsco0TEbaiggmhZDZLTC+rsGUngd
thNIaHnBpnrApRLnLWUJ5cGYwWJP5jjPgOsXhY0eUMdKIYM/0b6vnlZzE9rEOf6f
KezCQcVmmnVX4RFtpMfOGZD3K7MCK6nQtIwO85KuH+rfkgwZtsh0NXlqvIr6I8zm
OTE1IKrszF9r8Yk3EQABVUPSlBstUrplcvJEM3aOMFe0tYzzuhuYyPp5pDOgiyID
8Kyp1/QO+QR2ufkglOGpLtYUSbjchTuENh/z6ZmNGILgb6qHQp6htYiBflITY4yp
oUmk00tR6p2+jPXYcO+5zcTHeiqsGC69w/Aiujhn8PsqkUOBz5AMWH4hAP3NaGpk
e5bn1l3I0oXHy0juVKCQ/L79RlB9ZnwEeRKeVzQhHagIgqaV+7n3xvVtnvRWIIyw
lN5OpsNZN/AeVb2qvbvW0w9ZU+C1I2vtv1VfGE0LxVVq6uaaCJxwWzE+Ns289bwo
+RkSOTJ0Ory/l3jp+O/E233jCyC2E9wI+NArSTzOwC2G96hNNGJvMc4srLgw+uxS
hti330bYo9M2aiBcAK2J1X+52Mf6bhriOLxDVfM4ofiKYYQB6UivCuDSNZpaqMgs
iHAT52FElMQVZfe7J9vT1rvPeyyrU9ujm5ApLzOwv1UG6FTnwbMeZlZMc4LzQTCc
lRz5SKia8Oty2PkyekwYTihv8K7H2AOt378xUtdGybETCvuH0beGYyAzUkmz4YbF
iZ80A1memrqyD6KCDW8y2QNtlNRiVEPruSjmsP44phVolgP+5IbsCWAWPqI639ZS
A1ZsFLvUjp59uJ16cLJ8z3nmgql7qcg3nNA8L3yKr8PQ50fXVFRQs3R9vz5Mkna9
hDqe/YUVVc9S3OixGPWTYQ2zMFsoSs7KcPAXAmXelA4s0UyauvFhuB4MrtSfJjmt
LhOLrvqsAEBkAJvegj36YlAAYLPSZrVZjqVJpfurqu8XD+EP9QCUyW//3ISdxeet
Ieej7l2Hi3ERi2T49ndYOGi9aG8Z5mqepW6SRVyT1Y7a0Vemlz3eTT0YFO3M90x/
KgrU5PCIr8zl1ef/r9DDPwsuQqfRhcVVf7+R8uAEggL93VP7gUUXcLpRNO9waaFW
EI1FhdGpmHX0SfHyy5j8ZOlZRjb4y35QvaztYP+4DAWfYd1jnr94uSLa9MPNwpCq
T/mjNbU2Z/pkH6Zex8T7QVxbMfPhTu15A9y2CyzxUaAGHCKSiWaDeGMvTVmt38Hz
Q56Sp2y/Lh98CylsdesY/id/3F4E1rPRcvEPMAgxNwCVlCAxTnaG4IrDvci9sOVy
WXbJa2rHFh6wOGqIzS7JPjyhVqiENblXol9kSHEzSmq3ivQ/i892mYg9odWSEJ0C
aOhH+T8/VDAe6iqSehgdrD1RgqH1cSoToKCR6djegei0BwxAY4rtEmXT/NbPhYZC
zf0kH0nitpvv2iggoxH4/aYSFCTbVDskzv8ekk8EbAP+3DrVS23hiqaxsUH465sH
avi6E4jbKHPM4/Mn3R7rADIt96xmiSnE5tbUU91u40duoQ/tNkVSxOBFkdNqJIU+
E/vzXIYALtEqqwzz7ahqfxRZUPFhhEDCShnct5hH9Nlt8VBEF24HLZhz4k+X7DLv
0NbmDBk7TiNFK/dirKpc+SwFGVg5T23kpkAEDSK8vOmTCTG51UOGcNxhxH2+U73L
iX04UcseqgsKoQGYy1HBochg4XgsAXh8vrJRrPN/Qz2zna5blAYtTAHPcT4tUEFo
KCQ0l9PqueqDwDVic+orre2KBilQUqUj1CeA0B4N4e5tf3Rff/XQjDoGpLF5Xo8R
mpz1GkTVQx7g5SWNALUP4rOosttsa8e5NmDUYyXaYZdu99h/PYkXKo8wimiep1ft
OnAba+cZJo+swOAgvrps+gAXwWcc6sicv0HtXBBqHyOX9w1gV3Zw+9LOTiGWOM7x
QcZmXFvV1Li/d/3FP9buLFAJtgm4kR19tUMBvASvsv/Tt2B6HVxsj8cei0l+45Wd
zCCJP1+4osbGU26Fa56Nl3dnaw7TitO1rod7986W2TX0iAMIxHLDKECcuqnhRCpu
JtJCpyJD3/yJUoVyj1/y4PuYyl+WQNdTpPO9PJBZWg/D4RsPPUZZxsvGxqSK0U72
UcY8wNsX+UWqk1rVGCh3Rvb5sBfLTfysHPuFTkdJXUfHwhl+6YZJe8y5b4Nuxpf9
tL6ScjZCRAoYMOug9AcEmS6lBLFdohHJMwC6Fs0r4tAvs8jfnF1pLH4iO9Jern07
8F7JGz8spCtH5Si9g1c0Fo6h8xXQTATDZQkcOTp/PD9HJL6zIrUNiov114BImC2N
hkc7sVLTt/YwPvyPQygNK2zxtYGlWKDJ3To3rAMK7RuY2oUpeSGCi27XtECR707g
RB3x6BE8hu1SlyvtVado4BhzEQ34ZIkOeFetLKsD1PisTsL9Ab0BFxgofGceJngi
Ort9MuLI+PxOrlvJjalfVx27mLuv6NZ7vA7N+TbIfnXynsaWO7RSv9hUnsfSLHf7
5WKqgCZmzY8kUTFPwgZEODfjjBOTE4evn0DCs4QL3NqzHEroAOFNP/UiTjx9bQ8S
cJgNzPqTEGWSCojx3zqYdkBNwLU283+D246GkM8wE0PEWH/uPprMCAvKaLOyu8ZU
IwmthGJ8O9KCzhTprstJEB0SbkPfd3kyf7/pgE+mw4h0WCrX9tZh4d+xFoqnKlqF
8HTW4aJ9piAL2d0ZZ59S4utIHKXwK+occ/cqRcsLDuYi37Ww/naC4qjYyvrTg1X6
zxys4wLh//hj8NCsbgzCvf9mhBYmyD/uLrchcEwNNCuCuGkFMYCAIKEZOczdHtdm
VrXBv6fZn4ZCmmFqv1YLWlIsflumYS4Nyy/tS+X2vSSNLDexmV32IYKQqRLrzBdz
Ix7edljRbQ2SFX7XUL9pAcE90y517xzl9E/p+04xMuZmFfwzxmB6RZEarxahSl/Q
pWEh0yBzOSBreconVjgmZRgAYN0k7NUDyE2vi+m1kB0PDNf7ijaCDOTBjAz7hwJT
FuuT2eUO1VdYEfB/bbfi0B2TZ+xrBAmCtbRYtddbD36j/cbmYqzMACGtSAp+3jD8
7uhAC+fmFuxXDcetDBiqRGp6xOkiTbcIHTo6kFaZ7VQuUZiE5G/T62XCz50UWVeL
fZi9dcfdImPaEjMSmdDk8TLGNNQcqv4QpxMSBQK5fIizwhhIupJ/lqIXuEUyPpMR
4z8YjrowOHYFmESP+5vhSFWfxpPB6vTw6rQkFuTsj+D+AI8SL41/pUt32UoaYYax
vO7DdKa9OW+fbJ6QOH2wQxEmOsSUYYptYi6qO24ef62E7gcAB5FFhXD6KXQAwIUZ
gdvZhvDp/60r+C0wQZcjw7hkvkavDqvCP1gS0cvPuz0DB7++KUpu0lQ/CxJU6Thc
3YCdNIAeTNTfxQT4vpSTTmYy3rZ7cxdb+Ts5qsNOXd0LtvHb4bLsHHPoNAqToVPT
GlfJhnneZtvzgaVDuiAKce3afG/1Adfdiwo6m/p670ZOyFF3vj2r8KXhqrxkjQ+A
7Xs4ZdKRGpkiaQOMjH1U0uMGTSNfrWoeKUp1Pf5/ObMnxBZZc+EYIy10E1BtO45Y
z+kljN/BoOzOf8Y60AkHnO5Y+guCaYLdDLbkCojWmfqZ7KD2ndPCtdcR4G3wUlGe
H5qkvBDfxMqgGBO89nRivNM6N7bEzYLeoFahFRgYrdogKRG92P8bBT20AWznVjwC
QeRpbGjgyQZYjJh1bbJEGu62kkywPsnzeRV3b8J0mK70zCgi9mtF8EKQGStzPBEb
y08DrOIstZL46MCSEELIlf8QEebAHX/Mv4fgoTvJupApHmE3bqJ/DN2kFx9SIIl7
JJyXpu6x7oCXYeBBUNWxhvd91o94uR8i5Zu22QoVnx0lOYOyJMrLKMBqkKnnQYV4
dHkygMYH5kINb163asUkNwUwmDnM2YuNzMa/fYfB5TEo6vSs1QvT/tPzU15reQoN
Lr08EMaq6y47EIkAEAp/UAJVkGK9F5XKljDibGs2kT0AXjQLlWvEtEX69YPPo50t
X5v2GkzXpNHacRWa6ZwJpsI/fVxB7z7GDZr+zG86wb9r2nObpYXzlTHbFwSTt/ly
GIjcccKaDyZvUJKxwkFB4Dw0rh8O5UReAq5Nnf/gxKVzDjutiV2zzbPKrI4ZZTZT
AobfONunivgrWo+fTlwRnZUUT2OoU0LtOzCDy2OthAQZJqiD8350SfOSwHxkYkBD
NMCNAuWWrfZ/ve45wdIk1AL8suVnZeFVtSFl2hYcmWv1pVoKlxu90MqMoPODgf60
5C2ldS9XOzn2WyXVtdQNB2bJHhHjhos/4lBQZC+O6srOnBpHSNiTPz+ArmgurJWk
3u4+vBis/TjQvuRi0uRpetmboS21KdkG9TJ5maKSnC2VwiLCDaRTBhkO+HFWjSDu
f7fa8vCQd+ig2muma1C4EiFgsY+r4QeOz4/NHgc2BygAQg2Ta4o3PUMquw5Gux0F
kSF8CIoqdm/hiNdV5Uel4NwBeP79WxIPSXB4UOuMbB8BO4g1DhqJ3lqag31yM6mR
8IPPl1xwbdyBK1cM+Z6CVlQADfQb6MdtdHHjrCI2NIpxv7iF2jj8v9597zc6ikbj
SgY0ET8KYZt4B3m1lCi8JO6XTTPbmoKRk0OpKE2aZbcXe+ayqMzslZBFIjylnSqx
kl/l+OREKBskYqj9mffvM/tcazonsUX74eMJZqgbJw00xsJwwIH2wCgteQnHOMb7
7gHD3NstpXCRY34btMMW+GNclrI4206F9p0JaMFJFn6WxsaOuIS1R9DFMrQ9MUxp
fP/3anYBrUcD4P2dQvUvQ3CHzYXKILVEIem8mUJ1WyZm329zLbwv7AwnomTXgEaF
jq9cD75bCV1CGSbywxiTqEDzmJseqeVyv9QMDVC+HixmHGRl5jThXPFtmFEP/c9H
yY++FQ3Fa7QCd4KWqiGxS4LS1f4ZsO2cjBCUCahMIhqqTEH5AnVWukmvNPb7HGT+
8IlupTqLIymQleLmKjY/tn7Dqc3EzOVSNqIsGHf059dJY5GaT4rQTTw751bLKNgC
Ay7shqsZ4qpWqPTCvoxEO1ZiaNhxOL0E8ynSw4PtTML4K6vS1QvQJtR/mw6jGxIh
TSvwq9HprdWREXo5bZzC9HEa3ryUGqeSlkijX51riqpaH1BHwGqEFTxYxso5uGUE
ATh9gTMgKI+pxduFClM0t/FNmBjKatwDC5WOfsaYix0DXgbinv20JNo6GtPbNz4c
SEFBlQqOxjRqObsbJbvHVrGmftHn+JVYE1v4DhXrJArKflZVUdDI2UKpr0B0QP82
tGRguKFZJst1Q9X8NTLTubCA0S7W81NkoXmiaVYZZj91fpOfdd79plf3GT4sGAri
bHVe/Btwk98LgE/GCPC1HNjYdywSnSFZAkld1Ms+yXZ6pzB8oPq3J2yqwMIQT6lC
Qe/CcAbQbfgsL59BPjCyqZmAovYyeNrSijqEdPd42Tt+ZPOOU+JbDepPwFafGuZV
9/2tiBULplBLJf94xClpqeIvy7X20w9cPSU/9AwnWyh1BDS3EJwAgkLaOr99Fjse
7qMYFIM6Vhtx6Ob2GVpaptvHimLBlVEAJUDpDJZsDBT8LGOWwply6/HLa4GJLCat
NE7l187N0Ng65tWq2uec1stZAVLrXPTD88FMMCsEhK20CtIttRPu9ZXKpYvD8iuN
WnmgGu9/f4b7Rlk+zUsvUwWfA+UVGYnBEN/429aCkcIHxD2Oax6AcuA9zXq5UFyh
nPeMgC5ZQBKlabg7jlo0cZETnh0p/Huke14hQv+T7mMXrFALrpr0JxcfGiWyS0pG
X+dhso3iZkP8oeJ+GWwMrnL1BEt2ROiPXPkwVlgdsGJ+ULgIkRlWnce0fkCMeEuK
cbaVfoGG1eSt+yEpfXdgJrAuwRMa3DuNnyqrzhwW/1NaJogcK8Rqtksx7dBU7uDD
iDUY8hwTI8Lg750GpeftGTKHKGAVaOFISRf2RF3662O9qYm2iMYwguEcNHJQ/SYa
J/KYkZ8lC7e0shFAc/yuF85GdlJqr256ZsP5URSegFCzk9h6G8cjp/oQ6VmQdx9v
WI1BSIS2OP6lEKBgrjAWDzeAbW3RmNpubWCQrPR58no99+mpdSkdIqNRQq5TVknY
g50a1K4Ak1cmjEK7b0iMP/zcjgP2NQlsf5/0T818N78MZ1lCh7KJIhmqApotMCYR
z4SbPunScP6YUDYbwGfOPpb/e0n8MJTRpzQ9vrJTyRN/q342D0OYyp6Ajs/HcbNH
IyElNRDwNS/T0xye8ZYnHyn51DcrQ8dIj8zsgTHH55YeYbFu4ZWHq9Qt+kkyNByf
3BbsukzbC4mkj+PfgLVPNb0/ScD57kMOQoE33MwENAK1xDkKSv5gpDL0pXB1hKYF
13S/9rjGYcAQwLpCuloqTX+PO+xAupygKIVZ6bKDuM3wQny7tQo0HeI1keIC2z/u
VW2Uc2uTJgd617JuCRvO6lYxbV2idDG16wJeHcW76UcAugsZqtxwrgqjzu06BT4H
Lvr/JmC9YVavldq5WAT0E1i0LaVUJNaDvL2R6sb0Lpjb0Z8rHDsmK3y4CoUXGRt0
NXcQ/sMPPylN1cOvtWQHHDjzJoCmq7CGoer0t1iCgW5PkRUmjQdZiunhrMs5j0jj
2gt39Hu9q8wwWGspsZnHkclsHDMozi6G/dhRb+SdlOeyqJ+oZ1ApDUfzawY95LjV
ecaBcPrrZhd6tfzYlmyMKlTj8kQ1xRd21pUPlCa9uUEb0QeCmK5GFBtAeig+Xow/
+g1iTr4T3RRcrelz8DU2KywEXs4H5BGH5QpB5Xsbm61syCqqR5zYFlwKsk8sLbS0
Z4rI7Xki5mofG56GxRLnNvuj3LHhDBgftUfAdTGpTZCSzGi7VAha0ylTBjb5/v22
FXKyIQdh404U98M7heRHXL5eIDipcgs4N+lgWkkb3iH4lDjKdwBvsG7jlltCLf9y
LwXjuy3O+mZMCpqywLV3nkJmeNavErKTIBmWrgEPLB0uxnfvfvKKoFzhlkIvX4EZ
AJ7890yZzETBJ+HGmAjDh3qf7sZIfDVtWZLTkD0OdSOpyFygTtYACEy56ngKsJOF
apQSPCQkEYhOvOXHhIaonsuoYDlEpIM5tXLFbcQC0MIvUlPW25rhL0nlHa0RAUnO
nCYZoTWM1wgk3YL/OuJbXdrGCeNMlVhPtwo5MJGQNRMt31VtkYcVPzmESbkEYFoO
vHikb0JRCYaurcrNvqlvSfBW1w3ndnh8ab1l3EJdklf3Gkr7AnvyIL3vpbmtz6mJ
bFEmb92YHVxpVRIKtuiVQpmNnbhR1XevdzdDIpFxJOKQZGo5fBUHRwJGL79/70cE
BkBZTe0sI4JRc+PjcqmpBfjYpCGe0BzFAa7rR4UeEZiNxWSce7e3fme8Y4P8oJip
VT9pJR3otm5AE8LwvXRB+AaQ3IaO61Fy/XxtTtcenII/MztvRMiTKOfYdGNI1/JN
dTVs3AKINwNoNKdoP5e2LC2aTXXkYMk0Hfy1wfnVT6YHk0pc8mLNzYowzsUbROpO
yO+YKC/QtQ9rbx6BtoYqmOVciUJDsHD5jUXc7JWggToVjj0wnLG1K5PAdumH9anJ
i0ChDbpMgMCAnW9d/ax8s4dZ2a4sykqi6gd9EKU9jSDQTlLVdElexAYxmGlWeLzj
fIq6VzhBI9LzKqUdby6YPGt263iuOS9RXLMDJCcHnOd9125Y+lhylOZR+yPNMUz/
G5Qf8VmVeS/YgTl7w808XgcpPwvvs55RnPWIVnTa4ybXHZ2J5UodfUlnhIMvWhwV
ClYGzsAmgn+VhIz3dkuNpVDRbuoj5Ng9esfaZvbB9WujY+PW5sRbRIJ9oUmqu6Qn
1KhSkOSVyGeC5wiKMxkG1qDUBWfDN9XzNA+sciN9GbEy8Ble1RCWzQcm/GuiY175
tvt/7840rzogBjodzd7sq92SJlOdd1h1PB6ns0JLXWww0P4IdVcZ4S/gkyY1DRJM
Kg9PGlo6CkWBr9OcbhL2VNEtVqDfskmhrOlHQoxCMFGcy3OfBQM66J6LvJ8ChpzD
jglzGRmvLyBrB3q2go4Eo12nN3O/KWsIo0ihXVVkR4A8mFrM8YymdO7JHnztrUVB
X/7viOkd37wWDyBb4NL/3kKpy+5236jBEAH+NJ3D8uohkEP8V6e6Jm7VgtZ/t0wl
c4ttLTTJt2a42m9SiMpk0uJtkj+swMry6VRXASu1CqZXLIADNQ1er8jYDb/Oy/HT
bevBmeT+y8zO6gkrEDGA6SbuyTazX9zWJtyYC29PMnQRKwPvaChvft0YF/CAB1Cg
N2Zb+eMHWu1WBuqgz9W6qkcWrABpZT/VxkYoi94ambyeqG2eHIQGqSnetePlSuJj
zUcP5pp9L+yBaiaI7DLiks73zlW/djq1JA7bRuxsRxQnnQ4u5hnrOCX7VQm2oEM7
U3rI0JFHSvyjHYOJJkG061bkfNbgKQvcstE5Ls2xuUbjHYAQfP5dM2DymtGxWEKO
3hGJ5eUBS+NDgUraGoucZSTsE01DNsKfeEoyNmKJ8E6N1eL4L9teYiv2f+o7RWJu
9eaLxzksA6syy1VBJz1ZasOwZu5bZiGhOcI2GU4Pm+IkNc7wvsovuOBj7OyxkDpo
MW/caguiYG7QJTpkot9ms/xbkJYvzTNu+tTPjTAFkNHLHn6VxHOCCCuA9rvdt1eH
RA0RWJWUTEBPDg8g2oGKPL+hkCS/y85dL2+rnSbK4GANA+nW0F27FmBbYXHngdyC
Z06ZouURjDg0FZzZaXPICsZE89jGJp0ZFc8jQA6zSR71RcfLeslBes/lwcA2s5dx
wB7wVGw1gxrCvYrWvB6jcQpZsQYDZfQ6PmjdG22HxFwB/3TlRp6dqi8cN7BGShPy
FRpLjOVMz6OKXHN9520nnFq9ljGcFvueAjMmdnC1UYbLdOaEww/R0+Ckq6Y1uOL1
FlVuFvuxvcLgiZLLJ/ZAnFOPxHUTaVv5cE4lnLbqebHT1w97XKMfrb2CXzF1nLMU
95YaBoFnZZKxEwZ/cMFiBwMa5ZoyB+vA1cqLY6xjNW9X1hNaotNIO9O4wsLuLJui
i2kcKaVLN1PD3hBwCMRRqyVAGaBJHLQlCtA9NSYAsUOybO5NFSYfoOPfGgvTCKC8
y/fnXU82a3iFf9SCJ54o8QnRDZNpYKYTU0BLSK85v07vbSv/Uw/i4o/S6maLO94k
+filR3IQ2Iiqe9mZPTzn+X/s+kzAXlt+CcP8cRLfpBRlnH/0kBmyrqQRvKCAfeui
PwDcLRgqOtPkUJokDJFMhjeaFfzCrMrb9c1Roynlgf8lFmteVkl8xEgB1zIKxBZ+
27GYzItjEiJbexmICGRL65t6Da5zQw+TbdXCb2gFL62KLZtZCxYd0MmJYJVprYC/
sz3T6iOvh3HkqyBgC8KusKNSiP7Qd7uI7n6y7dBo0+53I9l085N5bZkMu5XbG0RY
bkI8KhxEl6G/jphG9zH++a3G91CK+TAGP6k2DMdbmOu6IA3kFXC3IllFbPC6dZYw
axzqshS/e7pHk5aE1cKAXnH5sPTqBXyOrq0FoJWncwNBOodUupbeHWYv32evvVKc
eKo0u/paF/yCTc7rZss9Rf4QQjO2oKMj4xKOPjHp5OGAm0y7oYOpmUHm51yt3GyY
s+10z5si+xeCHvOyF0BjwUY5yXsKVHBNTenBW3iaOyBLG3P4E/IRcrCNUgAfBHL+
NGURQioeTv+5Iqp7/+8PXb/EhM+kpsyyQP8Fs7HGISh4wJgV3aSkk2XnrhJBMZw4
P/T2rjf3YgwmjACxYpWtgBYKQa8lsWSDEzmtwHXQV3OdzX9TiONAMeF1nzpaNmQf
D1Uhz1igC07T/ch+S+yb4Nof84vQCcCrdzi97xXiN/yqJg7jZi7xJaJtouh23Y+9
Oqad/p4kQMCMvnqETDlpSxIwJ92mpBKj/712DG6tYacL0KHq5WZBQbstNeD4lIL9
LeY44P2d6TGh1u4XbaXOMnPLyCF6C4N6704Nh8ThykN/Zui4lBc+DC379aprcPfa
9WAqTlk3RNwoacOQewXfw9Z9SxPZMirLz8UW9+DPKy+fFmXlCNRfwMHIorWNpGYU
EuzZ5glNbalxRDT43Uo/klHl2unfXLO+5N0+bCqI2nulnJn3KKCFOnZiOTKuzTuw
aPbRFK6ZyBZ9Q4l1Tn0s4o6w6ztfuzTMiU6QMu56u72ndvKypMCL1J7ydL9tK5mj
a3VVS+5nUFIOHpnFUKZbzLxkdh9TdaLGs79a5jApp3WlwVxhm6p0Dy4XKTT1UPqx
9QW0OJhkiAtIzz8Kh3/dGb5RHUXcFpDMoGcZkKKj864HoReROv2RVInnpb6zG2Md
qYFVbQa4NTAYRvsii0qGQLq+jcz6RhxPpP0qF/HWnSTAWwiv2U6kkS0RgYickNo3
R7lEGvhQBXaYo+OBMbpxOJaQbrUSYFhcfNZqHdnwfkgLMqeIsbOJvNh3Wjr0YmxD
OQfuk8i6f4KOhLphsYcTnrPPeeTrAFi1PUNq0qAapgzR89S0VzotEZmLHl3CNDjo
bp4ILdvL30aoccqKDmjCwi2pYCBujfI8MqVlxKM/l3cMRGvPKrjmci6wOQhrdJ9F
8wssVw4LSy1CVvGM826UbKe1P3VpKUu4GZ+JHK/u2PM9wy895AXzypfw+NTmk9Y5
t5r1N7frCVdmY7eB6csoJ4Tmunm/mi9aFqZm8D6dnklzdCPNAg+7dtpTzEyIlGWX
FX7SruhdAo34pTT77ff1lXoAzphad85LnpiCqGBSwgVwqyIO0PGNAiqxUBx8PEAo
Mo1WmQIAZS1M3NPDupzHHoiY/wSQ0BC+Ip3tg1PMmakTPHPXTpqm2NaVcKah6RSc
/E3IcB9m8VSY7/4bHfBTTNwnUNQQtc/K/s2055L3mlAb3ub4cePSgyXZKdKgnSBD
zjfFSvTdQKpIS7jyhSHqSa4rFq8l1EUkATngo9Fr4o5r+wB6SI+/Igpl18jDwbKW
CsR+NUngLBcZPAIaT2WVKyXsrJbbRggOq64tF+5LfBDEuUbGA4r8JGj28/U4wJYU
w7wugiTyanNRj9WzXqb7B29oPVSNE+45Yn6ZcTSVx7YA87Tqn9K8KFpoYIjaCpyR
z2VF6vbKbcrE/oPVVd2uZ4w4V2FxRNSiCetsj2+lQt9zeRargukh3Ipswq4Nb0Jf
UnINxNKN4kwN5c3gj+qUixGw33/wahA5HrZ7LjFPgUZSEFkmnPIdBrfZC3aZ9X/v
/3nsnXvesFC4/lRxlbW62Iy8Kzi7xxxrPDTwH9GVs64ccNEm1D8ibwnVU8iDKP5s
iMd1nsB8KIGospqZKc0ouMH/QdWFSoaAFnSfgcmXjQgNRIgFzoAwYFs+SlNuaLnJ
SbUSb0rf9OhIAjf04/eXLbrvBsAJeh6ASnYlhEoEXIZ8qGta+cC+z4ZXkGoFCAeL
rDFucWCPokO9U+lMlebyPEoagV1Lix53pPT8c682VcvVRCgwKCZrod7en//IvnVg
CNq1Oaay5IvCrvEmBgkBoD23i0q7tnTvCw9e+UsKM11T9Y4ivfyFVsjC6RkMthxF
dOm4Bsr2bvtDdbkGC73oGrNBMscV3vEsuIJEZJRHcVmH1/sev9GJcrc6Ld+6i9cb
iKx3QxnfcExoGIlq0BXR79Tr5PsC9obf2f6Myr634tZVHRZO/xukg1XnSJEbCRdr
rAzguhgC59iVXpC7U4CSpf7U61RxrrQrezJZkL+7VEIbmWMsoLpXlhiHIX5Jb5te
tZis+dKEcznqn2zYMryEJmsOUil7emb3dJm/dwxbpfSQ5j6dfOlWy32EEDwDY0fM
/vEK5ycXIUNbVznQh2ADOUUdYj+yomvn2sR82czMfvYUCCxlZsDcm0lY30FC/V3f
cuhBhuC+ZMSGbUKKxM0EG6TDOw0jfodyeHi01Z4Iv8Sbhms7B4NeeZv7dcDSu3g3
80QwCGFYiOv1XNvdQKrR5/wM9x8haqFkVFxkKpMb31GZd7M6S9mRpPgptFKZh0+V
dHcGddAvusasMqcVYz8BaMk8JtBsjdmQsCD9c6Cf29wkzhPvSFM9le57Xuz0bP1u
xc1qNkpJN9zMSUlJRiTqO/u0cuapakqFbZ8AGhmuP+NUAiYR/kuoFHtoy6aRyCSs
i3/IhbaqQW6qWvZ9tOg8z5DjLYBIunwEIvEmCjrUwvcp2vg59o0X2TBRo4kTfrTz
A8qPhdFGA2m7RnKwE0mn2/qnOMmJDoL0BLrwEgm3ZyW+cCUPAMA2KpWtBxQ7Eu/5
jW1Ri5FGaqVTX9lk6CJuJxXZmmc1Y2aFIy25niQUuI+QKemNP8BP1xaWGqt+dB6Y
r47BbWuyhcUSu18tER+G4xqki1Zh0cQ39nx2qFHbbJ1BkL9LNHAf5r+rkeyRhqix
g8wJB8Uxjat3xEacvFNSEL5DzqIbnYf9WhXOtnecDykh6gMAokTqynjANieQIjHD
1WKHxfCRZ0rZqELuRWHxcayLmxqPqohvQdBMSEq1rFCq/IJwxfKQNlHeKMN/IYEG
OT099whWMhzqQESNJHcgBM4xB0EorHUzM8IUyknsAjYN9GaUXr1tmEqAzzcJ95lb
RkxkC8YczYMHSt57bSprHjE0Pn8vzvR1OkGkA+RpBdfxP5Zn0AL/vz1hCeBiirBn
yhyl/o1NVXsGWcq9rZx+5txozZIS88fWsfaJW7HSmiSeqQkwUYuJuuR4H069RnNn
zJwjHm/vbcMW5qWOOjrix22Uy1LoW+qEtUbiBufnimUrKpeVxhmOROb/NvkskJ0j
h+xa7zEpIaCQQd1XGQK3I2tIiha2WkpBF3aR6T+7GXvh8jtjWDqqK57ODYasYjTr
QZaiw9qF5GGNRU6JyFwpydppD/HfS00cEeuoNobJ8A8SJa6u5HrbjIftGVqEtaFf
x8Fci8ZdGISGaKsTBV0yHvjGhfvwHml0+IZCMVgUZ1IyYC/pTwlWyWFvFckJXigw
hixyd8hAiZFLATSrtAXV1r81oPFdZ08AJxob1mMuNdJdbfvyfWr36GIzKndS4pGj
RF9bZfW38lGXGiHFYeImx7TVx8OsSoPljvqF9OlYUlcXWuVK+EDDNetdeqh4tC33
8zdcs53TLrVn7AVYmKHkTS0gYK3FleYGyRllaZ8EiYWmH7SQd6AMVgE5AGKwL7UX
HPoo/G6CKJVCb/i/ZrWLEDHcN2TUc4lShD+3bhyawHloCfav+TnHQzxb5VS/pLIK
GRB8BBTWOLI6WDYqK3Q1+TNbsisNKTCHoKGDu+YfARcwQTYgzDQCcnXy0Bq4zcXw
wder8AB/0cIccVQpi+zBXDEWAcOecWqvimGGtZVsXXdbDGYMl27NKNjZGrPZzju6
Tz5dfHbj6s10RTea0Je7KxyBUsXWMtsazsDrFUEA8Mt5CNeHYDGmKKiYhd43WId2
s6acFcTQjq8jB3EQhxxBdJXjwQVI5vqeH9VUYdc9A8bw7V3RJvDunAzSL/RveBr3
jU428oLDZKOChbp9la60YAHbAIf5PCMh0ROeSLr36c8tQW19qcOgNZaROJ5rgiUG
dC6BFS7WXfUt5BasfjlKl0WX4b9cHW9GLT+SsJwiq8xL5/GfPkI05p91+FG8vCS/
i7pYmgshAnTsybJwJ69wkKCAQmhmCJwtFkIqQFD03IluxqU9Mk0kp7EGNdLEzIPI
qUVGQUedZEq4BAs8LffRxF/dlLQQLlpRXVu9uzzOHQkiL68I8CcqOfc2JpEfffPn
0IjUpmZYmbbkVo6be2ztPbag+P/NtrcQrcUESQtG4zXPT9a3UE6oxbk9xYbRTPdd
b0BUil67OnUcBlMZNnTL2S7y6eu0w8CZe3VxNANOqdv+ooh9Q7mc1Lw3Zq5Z6ZVz
UlTFK9/H8ehMePdK1pcu2E1sXM46UEL1ND2aKkpSezRTe6vCrkHCc8CxJGp4uUKi
i3YEMI4Dig0Yd8LZkyMCmzHQ22eBGRckdKxf7UGtPVQNIgYn3AqxnrhFJPeGHUE2
1s9Xc98obdPN6q5FsZmI9Z8OrVViYSFkKdA40WvQpaOMYgzx0ZpsFy8aeJnS1WeS
ZnsVqQKOYZLpHr26RfStmt+uN0ntkHOzcmhKsheNt0Ah6snefamFugH4xmMRO8Hl
fM51BIG8dZiQC3zBagqegfV5L9NGQ/oNRIi4TXkGJpaCJsIo3+cU9RoPzREvjigd
742IsK2Cye2f6Utz99/o+tzawrK8V4jguD0TooGr7DVlat5RXaoz1e526D2OhxbX
5HjA4Z2g1A3AqTzrD3U9ezv0DBt4hy7qQXeda5AfMDMZoXkXwx29XwLZgzbQxpMR
AtTz7Lagj3oC+VhqUdnkMv5nog65O0eTI4nLf3bqfe0sIZMClcxEvYSkxDzQqlf/
QQXt/JaHa/j22Qj1UqV/AZXbchb8FN3nRH+CnH7SROoWzsL0WC1yXYQLWtOa+ZLL
MaWPCiari16abpaYIFHci/CawEuKq8Oi5+Yp9LArMv/5sBFMEhyqsdRklKTN4Vnb
B/6eTO1RkRuKPcF3K+ifxePfRZJeZPOVl7yYwneVUPExKW4Dcf7sTlNuu1Bwsfuq
UIznQbRLKJ56BH0IO/nqbRcABKiRuQdeBtkhNLJbcHP3ge3G8QjGswb5ZMMpJ8Re
FPcfKgFiyIxJ4xYOUYNwiiDDRbUNuZZPirzfvSqRKcn0Vlq70A8lo5EEB4KPtJlT
w9YCZOSuR5PY6KzWHuSifrZlRFkakF+Z5cqFdESCKthkXq6RWqy59vmYxg5Go2Z1
smLR+y05BtodisoBObtcgpJ9gWeZt5gZ8MUVXky5k3CQb29+tBBXolu7KsTRJAPr
4Gn+D4f41KFNuOWKe9lrz/I5OXBSgEUk5SL2c1HprfK6p76TmyD6WklN1wRh0BDf
zQy9V2D8vZ/lfNPclQz4/WbsxjOYKf1C3aMYGTmYRGbHiZ8Jsb5BmKdPWJ9o1wt/
eMqdgD6rNkT/H7JHsAPNBzeCDTlEq/OouXJ1rB1y5Qadn/xMd//tTWl04OWc3VIk
jVhqn+KKWX9ZHB83YkqD+obRmAyPz3TwICpCLfBicX0qCAnMEpWA0JPsTGCloU1W
GpHKquOXvoCMzrtsoL50vlVEvOKIJwYNX/aVFloxzkmSPwvkdNOQozXXXtTRuc8L
4yye0EdtZU020HOninROsCVTsk3RRsR/8mnBfqS7MPPvHGEUE5vlV17rHvp4biYA
JsrvctEGQrwrgJqF+qfeNuRGHcmyUj3ESQLER7ZqnYBMMRqohkSeDg0m+L/rrvUM
b+IBT7y3MSKf9qmvT2qtgWQneflam4Cd6csJFd3aiMO8uPCt7YNnx5VCz/BfyHzB
5FN40FpMY4FRKjqL7C0ANntn2C8EtMMTmymK/Fyd0TTXhB68nsBumU8+SkYePIU2
t5U3iwskVFMlLc60KsUD3FI65/4K7MI9Lf4bvux/SqrKVraEJ5Fbo0lvEHZ6tCHW
QIGqK9kWR28nkjiKzEon0JyOoL3cJsLpr23fIGHYSHGcAj3vdlQPjbAJ4hQ8IyhW
c9FYAIkSnZRlhO8b392svFvTrbS3HOGs0zu+fUnpqq4Yfjx81OFWgM3lUwCKiT/Z
LLG6a79bcmvLr/HQfDgDl/vdIYLo/ayWJO/artU7txPFNF8/wr5cf1XVOpx8Or7a
uxzGSww1QkhOmd2Ee3EV5ZRTcPeHpFPJKbUyQEf0LF0vgvFaIkaxJ72UULEcp3ji
mU1rPdsQ1DzUmwC4acKxGUX1fy1licyYJ/aDKibDj017rS0DC9ppCmVL3QFBsQMY
UFgZgEeTogmxML5rrpIka8B0BzdLjowfUc4D1hRqDHKhx8t8fwgl0O5byOruIvnH
2iLmxAT8Ly/mzpkDkMQc5QQsJzmTwAIetgfj+f8BKV811eIz/0UYclmYnH6GO7QF
F+AyT15OO7zMGjHYcdEtlKnKzi5awiOOhKad761gQ8iM9wsIWyPQgh/6eTs5dpDv
D2u9ucetewJKHfJ5oIEJ1/LuKVqyAdv35RktepubVw8hKodfxo1aMRvTAwAG577Q
WDVAj/mzihxuZ2ZhioElkvxni5z/mcoRK5SysN8mcRjkaPimjTs9Uc0qqWftqxiw
raRH62ySFEbxQsMjdh5bdelvD3Vug6ImK3Pe0LYn87jn4cODmIBqgQJm1siK7sGE
CKlFbOmy2hrFe+lt+6NAYL0DJqW62qLx49k3li7w8mi+zVeRUVoicTWxoGJbyxWG
CksJdqZH57rMdjld+JfP7EDL9WvC76XGgF+NHKVFPV8e/QnkP/d1/BIBlMgX7RQy
kx/d03tGLdqSJ1hh5NsLdswtuj4hvyBVoa0ee2JYrYbnQPWoeY1ne32MesTaMpcG
TmSMDVd1M5P0IVK294h0CIaWoD7twjNHswRgTIwfufvQTPUcLgrsRjMrUDHluwm9
9UcsAbExtAWvAUMsiEC+JbKInANfWMvXcDEiHxS2r0DpNcJvcLEuAbZQqvwEi06M
JejfBceRFqPKsJzDhLprZKZwGonX0Fiwz7dyXeiCvVyNArb6e+60B8WgzXsFm/fz
1O3wf12qEXd7TpLP2C3j6gs5Lu4ljemMr7oE0IaqNSRHzy2JYGVHNLF/PPnXdp42
5yAFHyJ25koj77ltu5e93skEpUbZtgxUPZI9LSsarGMcJVD9CVPo0NjrVo2mIM6f
QY5Dbwepr3xL7Q3Z7ZqhX89WElxEH91Hv379E0e/15/+T9g5LNYhpDQJ/LUoqb3R
e8dOYUlNkIPSh6ll4SgTnluaKZsClHxinr2dmOS25CwrFnurPAA/IDDj60oCXnXz
MbZxJ9RAsZ4ms2eCsebmZLHfktZx7FkyJfiyodJLIqi8JK7JmwNuBaWDEAl2oq7z
oygNB5toQAl18jn2ZorTZ+GhnwY5wGp8Uz7+hgiJXb3ecY7L858p/TwybLeyHQqc
wTFuDAfmmrDgADij7RB9w49xBIt1wGEd+RBpr57N3ZdwhSNTU6V1Mai5bbAfsr6o
MfVx/YwGAkSwAVfTg3BQWBKYXHvTA3dv9ZzWt/aW67B+5lFxxVc3wxCM7YEccjNY
TkNLosRTB2RilCH/EJJ8zcQGem/Xg2gDCQ4AYOc3Og2n11zCUDnzv7QyCMK5nl8I
nJPDA9Ji91RWVYnz6/Rht490QftuB9xCeEKTJJ30BUpZjoipmnaYJSr/LT63t9/t
N3OkvoHkamHBOHNn0vi6I3P/Nyiytbe+iBIsbnIGAoENtvYOXeTr+h9fSAf6mvCN
n4jHg2gvVtfnfDPw4QUeQYxwiYrEaq8ptRwhlaVv+zCD5dI8ofV7wAuSmMUgKb6Q
Oz3nBp3qyeV2QZEkxWCLxqOr5HYehgBGoMepPomvQDaJPbu0C6hJ+UtdlhLRP9I8
lDGeKzMiohIwg2N1WaUGwDTCybT+Ii9mz9BHkhejbtBGv1H6ZEA+1c1pQjcgoewk
OFR7Xe7AXVd2xrTKdNwE0cwRg6oMlubjXbxknnHadkRVx4kd/NhkH/zyI3zgV6kj
To5OtNkOUO49uKTf7eDTjMoN1cm2CqzVW1zVKJHq23yH+L7yv+TkJzhhXehxzxEc
nCWwlHHxQIzYY+qDv5XYBG3kSwQsNk2Y3jVqJ0CztmPwBd58T9oRCJaCsKlmTW4/
IxbC4IeXhmws863ZAOR2I2XEsw5G9R4VXBXco+2tF/lJcxOO5uue79rWjkhDk0Br
o1cgMbujkUOpR5EUjWYBTHUR7Fu+faf2qdSH4oe7FwpaWvu9RqWVd7PlHMzMCBS7
u/wrK5o3YYbjZrLLRKY8hHh1MssCKbnVmhzelrgFBh3RoSm9QJ1PS+Zprx3ssVVN
XWFOQjxkVUaRjKBzVi7S+yyyebYTOLWtBq7F0yVEEaApxaCEcwbPRnqJmySTWIbf
fGNQyeS0G7w3rA6ort5+co60RpL24KNYJdTKmw8MRkHODjbGrZV6xAx6AW7OdMlE
DFMRlQ1zcddtOdVk7dnN2EC4/qodCmBZepjeAad2RDRL5+wG42YFuFniUyiRS9UA
tiULFvSAlPc8P+ANWAbeWKtpIDFT6EfQrSfQ1E15csGm6Fdk2ezk3nRmKAvmAkH6
CrOeal89LuMULVFWEzZuj62XEXELiT035ugECYFgg0YRPlw7k9a/g3vDJ2nM/fOr
XRvJ3vFEo9I2fImwp8YkI23RdCdoKSsMfkaz7oDtsvyITX3lYvwCxp75pJirHUMf
l7oj9gE5mKD/Jik9fXcgvsrGa14a4toNPB/od7LSgKEJy9ugshNEnQO++Bh3cO3o
AVtF5XShu+peCCkmKLIXziXKnJm6K0p2J8EI1/18O6Ee/Mimn+dNLYUgUK6thikq
V4YpmlZFpkixfLhS5zNUOc3ZfeBQVWEuqpgVFmu8RuZwy0w0u68Q/yJn/vtHgKwN
nCLu/4r/hzGWrPoATQgtwZK5NwnbFVcIxG01Q+uceveBQcWVnvIyGz+xjj+hyUcC
NgodfhR5jbIXGdPGOwhvXXGZEeM3oHxGKqsySSSd6cQ3tAXZG1C3f7lbH7eqP/U5
jKCJ5RBYgsqSbj5+Dn+T7xELEOhcvrRWGqLMNsZEfrjS9IOe5KwhC7jroBLh9VEO
urNUmAQcOu8P7yr3BtjGg7pHoy0GW/7WduRfnaWLRn3c//e1yozr8VtYhkojPirC
mIOZHOLS4Dzt/cbt/SN/XcQK1YUj83NuQ7/ncaEw8wcFDi5zFI2vtwV+I9N93t3J
hn1zAvNXpZV5DL16THdfPjY0AUE7akjlzpXULezZDY5Z7bdcX0INVr6chw9QfBuK
GnrNP7x/B7BcODbXue3KU47NQV/h2qW7ddGkhlySUswzTvugKYrXqMc0ozKPxdcg
B9XrD3ShTdI4t1+kKoyG+EtRIUBjbNoH6Xel/gT/WTY43Q9FRZN6KqcR+FfjgYt+
N+TQxIdvr85s3lPZbZlR+xg5EqevbPfIxfbonVB5+pkEHsv/ctGMoihm2uKaK0hj
dSd0Wvob1ouYwheomg5xwvA4YvLfRsZUSy3mBUq0h9zVzV48huZT+7f5bgatH2ex
TejHO+AfhYVfz2ceW10kVPLy0lstPfS8AAEL79hJki/jZN7MQzy2CWVAvTo3ZqPB
tiTFAtuo8m/SBR7M8isLbaDvUM2UE6cToQSOlyc48/I/ETNXM8QkLW4azM7ydizq
R6n65hdkCu92r473h798K0ZXC9jb0GasmMdnrbaOufb3Gmj43oslfAyaIRFmcmxq
ZogWt+dXvPJi2KPpa8f6DXazuYpSz/pd/M/PJOMNKx4GjhQ07Z867ehPwfoBvk8s
ozoVCL1L8bSDfEaRLnLyo+FHYSSOS7sEWbYcpIMdGdWoMyZm0ync3irB79279nBD
gKXopXx6pX06WsNWBwA9WF+B07UkmPvd9i3dbdKCeb1Tou6iyTElf11H0mx1Ov7Q
BBG4THPYs6UBTPPTLDW+3hy99XBHFIeo48hKIRrtTyD92fTJmATusa5cKj+lcGCP
w1UTUnmdsdH5Sc5vJK32wcUV6goxd2tipEfeMzsdbZQQCL3rGisTOA0MG4wdNA/8
z6T8a3xxbbDEKsOQ1OXNAnSh4Em4cn9ySJGg16+3LLcUebsGrGjcS1/S8eOPFKC3
b2k21rrthQ1SWdr0Y3pqTXP+4HBD7tOlIU98G12Azqq9Mux8ceqox+9QsPL5eHRB
uvtJhnoJ590FseLlS36A6mAQwyXnEfwE5O17Ih5Wqs86NkkR/kvClDAS81aHB/ZA
bpDmdL9L3QErOoeUIg8Diy1J4Fj1OnflacDF1zjO3r0d+tBLzSj/PWb9S9NFKd/k
JMWBtFFuOYCh4x2KjLxKWcWmVcTIcIIEb8loef6kKcKzQTpz/U2YVMLP8LgPkm80
cofRNPR2fr/hQu+XkmYvMOfYD3PcJqobSTMp6g/Vg5Li/rG0mg4rO+UROGdq9pmp
WIH8vfTU/F+hHn3ADHPK1CIsuZ8DN8Lr649ohROpJswsrhKQCtLgLUe+g7JLgYM0
yVQa4Qg7ozIMAJn4gl9i7mgTq71bnkrPs3rTfj7GDFZ1Q6yMjQX7dJzecGCGXifh
1iS3cPqjI4/jRzGr2uBF2cyltDMoClG+T0x+fVbIR/1LasmeDzT4TdzXq4vyZuct
T23Aus0YYuWm9jhQxi/pkDJLtGg2a8uMKWFSQAqCCmBzcs3SRdEurT7F4l++7RG5
/0ChPI95xShD6JIWtiSh0FN037zu99KvvwC0Z/jJw5nXarGKOo+k4dgyLJlG0Q3v
dNqs1MCnJgtk0zL3luMBA5OJBZDs2pMfjhVlAi5gLf2cYMvaW2n2AO4+eJReAYTL
/1phGKi//KE/KglGTDfQ1SeByeIx+dbJkXkYJQnWUNt/qtU8b2hBBlN04mu7qLAI
Xj1v6u8VcU03Lfx7cJwyb0TXcynYdOrCiRufcaHolo+Fa13d7wMLaC2NkjWJ+XOf
1jck+8lgnmqpT8TK+Oyn8BikS6O/tc47B+h4qXiu+pcg64kBZu+Ru9ipOU44S1iQ
dMIoDPIs/+Y7rapFBX6dHjv+s894N13lRCtJTOGW6hGBkptrf73E3XKFGpi3elyz
rGpqqp/+nGfQi05z8mrk3xrzy8aC7PrhV+CE5WGsP4TeaYSxYlum8SV+pxkOVSnI
SxRoABbejQf5r9vNZOy2Q2ZS40ZfEBqUm8vZYOL6cr/RSLJvmCmXy/1vICxo2Ssh
3Ogtc05CKCht6HxYymgmGAkcvlZR6DV/nFZOzK47DrO+bm7x2hSgF0wH0oNAhoFx
3VKHsR1Xu/zSO3odclwpV9Ay1ob0/jKN91oukyd6L8Ep4XbHhKV6XZFkTk1QPvYD
eTvdSGo4xPdjPftt9t0QNP8MVo8/kq/pQXM8oh2k5Y1wJ57Av+ya9h+fFQ18kJ+P
qYyNSvyVyk1MMmAO8uFEHKdCRyNNoXwTbZ11CJblrzkQripMI2yLAwmVQLwI361d
FORxA9kJLYSROjnD1KPdgLwo3GF0TDMy+XDyow9E1ZCuidg9o9gYZNmlwQhE8KFe
9IorZF0fC5IUeJxKHtX0RJo8me5/z4mCINaZZMdRH0gUxh1pQlWr2PpGwQchDq67
/QAEMG1RP2z3u1KeXz6+zqTBnHOSUYz+YFJFtGQl0fv2Zm21MuYoETuXexaVlDOn
I9AU7yPWSxq6ZEHoIrGiDbo+7r0Li7OA3oj+671W06kCQbzM+Q//PDTfBUk2LR85
Ge76S7vimxn+tvmWigqZN2//84O9Lhcm6UssNYwy1ZjmjF9qeoxd8OP/HjvNKJgM
jKdP316I8OYvkMLwjPR5WYDVEV5k15cH9Zbs68nzWIzva2NGDckWOEKmQtHkwhSR
YvgMNXOl/qKYaRvAGk0tIZUaIEEW0ViMv/ugq38aw7PICTJlav6WI4G8yHfwp2Hc
xUt3a2251/9+YcJhVVG0rywqdY8FTJxVPrXbfFCY60pBHyaHLGsUe5HAa8Hr542K
IbdQbU/VuJMnVSRmLYy2hZ+x1OMAcGQgTwrhVeZLnbYggNGfk9Cj+f8KOrJKzlCi
imHOmvRhJ6C3ieOdgThbNOB0+Jw2ovArS3fiyXvyfs0Rx0OwHagB0KP2wI/cOYCl
Tz63BmaDgNnQplinCCObrawxjSqqyem7GJQ2K9ZrdumoHWgbtzP3UBMGiiUvSooO
Y+gSBw8JKauCH6Xs99UEyWCVZlDQ/QbeOLKPfzSib/M9SsAHgV1JUW07EhQ2hqBp
JRwsb94DAHMKIDYkXwrKE3Y+VEkpLbFA3CBtis8/G+dpVdoc//XEveIn+OqVK/5e
ZcQsbDUd/YokpnhgBS621oSBliSo4i5l4obciniEQK9Ej1BiYcs+zzoUHV2GpT3K
Mlny8OYZ+a0lqFPUjPyPO7EzR/xSL4lv1fk6jBsmTx+5EOPRlp1UjycmV1XAHkT7
iRdOVHGyr0FgxVuglklFOnGqBEzOjQ3IRf6r7snwudh08I+6nLQOrzAxZvru75C2
o3m4uGFtx7caMO9KMvE5if4IhRtEN3thxm4uWtsKorDh+aTjFx1IIGRfvfnWv13K
UffyU4YzSZJisAp+E61x8t/Q+xG3EzAoOTAcCO1ygweLHqiNWeYlW4wgylsG2JLP
driNV+d+6DUm7GNVpmpTKLwQFFvQ1zQVibyjHFhL9d2Lxn5iXMI2Aw4hf5a7UkjY
dytHDt8TqBe37I3pmvE4mgTKUIeQkpvL37VTqdY7hmrUvAY9KPMXPItVWB6OdGDv
HGGxFZTahmcqmyIiobnMo+sn+AWbLzWBAmVXur7OZyy8cyNDn9gDv6IKxsQInWjz
hEye0saMP4XgHtxYIpAsex4wvNIQl1/ORQ31Gk1sp4UrN2D6c70xfx0X03J1nUtZ
pK222gkypoFJHR3WTXE9NoOHXbBynYkvYmfQPxOalOis+utVqzGeocuQeQbfeROs
bqsCrNF4V4mVzqibi4RVEE8RaTz4HutP2uJz56+/btrw6IYdDdxAJ0WFygzy9lL5
2nk1LeWl+ccFDOQ4TxQ3DhYWylrvvZ07fxF176DaPw4nnsK1neKa+pXPmqSDJsBQ
J/gsD4ZVePuUX3S72WpbvcjjlTyTNCIBZj3qRQmnA+mMfvU+u3ApB0KM3CWd/9+N
ifhgD3q6DZjHBlOT/UBQpcKesL0/s2CjZQFOe67QFHxP8b60uGuCyxyDCfGiKNFL
q3PbXq1s9m0mAkNKWsMGxhwSJMUD0uTDCWrD2Xt9qiGAo8TbspD29cFHvWm0kVYQ
pL4marAnuu5a47rTtx5u81DQ/lyutD0XSyexnZZ9Ng3P6cjYCFDmFAgqdf1LjQKF
zMWR7oFIXeiQV67MP1awaGsKyBjCs5ThhDn0jBcevA7LytOU1cGbaSEfntDyHSN1
vvuZmeuy7tkFiI+FwiMSL7mw0INzNuEwOwgLbkdWlJy0JoJoKfuudefDohJzbMTz
pRcoBJfxXxyQoMUX9985YMhDwgewc5Msd3kxZkg5xphpMZWVyVjrJJpSVhx4mGen
nU3Alb469DWDJNzPDyIx63lzzqIRdR2nGo98ZCl5jgDGq9dqQ7JKHa1M4RDw+1BA
82WQnQOq7Gmf0JczCknRe18g1S8YywpsgnJ1K7g0xjS5pURXubxxgwYsfNXrSSEQ
9UBBm4Sj5S16OjgDTEbsoWXrgOl0XVPa7w1UZFGpkhHpULdVeWY6fadJOsJpnea1
xjvqFW8Cpifpc+ljVnsKG8RkmjGb9J9cMhhZZ94TK90Ctf929PpdUuVISfl5Axvm
o/FgSNEkqUQiP9GFzYvi8HOV7EmNLwUAbfLm/eF5nWSMTu0a8myAskffERAA6bu6
ZjcsK6ao1h8HVnhunt3HPJTFJzR1q2HhQNmRBpQQce3AXmyuqbBRrh1v+PcDLs78
HvaqJMZp387HRWAp1di8l29hVZQOhn+ZrwYBtMxHAiEjO5zAjoQvaZw/cqBbPb39
RjC++yJ3EnVwAm9BiL/14SNNOqjBzBJMHlBKsdYAKl3zdFyjf61ElsWDsGNlMiDO
N2ApJ9SHwRAJtSlBA+sTwK01vFWDk7eklASkeoQYrP2hyR2R0NzM4AlFpQaiEe87
iQTQbBQxnAhqBB6FyfbOJGsF5MyxdzL2M4LlTVypO9OSnC3IIytwyk8hv//KUycV
e9algbBpMCsoH685etYAEq9rROQ5z8iA1LTBjZuLO98gRONX+ujQhJwtkC0YeyJb
lNfsV91SKA3BcbkvYH0/7HDb1JeQrOSPzDF1J1r3hnZlX9KoZFe2Nzx/KBrIqzJ1
BzFYAYltaJx/2kDO3hnliF75FGpA1cNy12ivEdxb+/u8Yz3sSqhQWVuhRuuSV46i
L2rvvYx0ngxBvxm9+DaIj+bGc8u1jjQOiGNNlkdPKWCbIESrdtM22ov/blxfn60f
kMhq7PjHWAPy3J0Rv4qSTXQEw1SJScI9i3btDWGxZghug3puMG7a1s1V45oADb8Q
LsAhPKWxX9QwVNhQ6BUnx6+Ss9DYJjIQ/kxX+frz+zaD4ejZS9MoJ1oU1jAwvo83
nTzuR+LI4r1NbEOt7DzVOHJPBtFYNF3TUAgccwfAS2WWtnqzJ99l/n+km/IvBOoR
l5TclBiebC8qkGuKTw7+izHA3NuPt6zgIYQ04ThuQ2FGpUMkPLMbGZ163P8Vl35c
dDNrj259c2FnxSOIVd78CWfJ3GeSASO80Gfz+gRKN1qZihHR0vwLV1JLIkldnpFY
zoD3tLINoIpDogUV7MCaXn74NqUwnlFWBXGB7GH0hB62rtYwDPhKVzeac/70j2gD
WdkQwFAy43NXPTZ86ioOpmMiWDUYBYbAuYCUIfCmOoCya9yXHiruy5ceBxwqxLmE
Ct8ZXCtm9oqQz9HafzDv/wKKxDkOb4hsVBc7KLEYK+PUI1O+J91MgNtTiW7TH+Hj
dVtEU/fDy/BgC7UsnOdtx0ldQ/0F/Sf2yXiKEg+7AguzlRlFgJPQl1qGIsVuXYR+
NFJHSUaygL14C7dYODeCHhWpR4UGbVn/3ZIqRBgmU/waMQZSQoQEkLycxsBZMCE4
0rga7KJLxSZ5A9jUX4iE8JCYfsWYyyt1zK3KJNexDxW7LLX4/1abWJNPQy9EA7dP
e/8no7mamEdgZANkI7zysUO7pj2jo2yQgKR+7ayUJK+iIRNbrVpy6v4yqFRVV8pU
GPG672HnHiMN7b54zcPrqdGFUlbMPpYKrrtp4dTRvsP1sVBpM/+VZbWRDL768p5o
EgdhlZLD1LidlMRG6AqiOuc2RT2pwBbVpnSFgs0X18jOQet+zRnIaLiwYKhunDBL
m0SO0jSzhg4tATU2aor2IRY7C4Xmhuhm38W0Vcrt1WH3EcphPqZyfJzc5ogow+Qj
oefeE24EzOPDvClleALx8JH1PbWhFEPfD9oOa5z9je8qILbgpRkJcVn3EV5c/JOs
VuJ+95WrvaIhf4m0VbvJC2TzEQhE/0pmmJRrVvZYWOvO0tX+L4elJd3Et/cVDEvZ
Det6cUZmZludinkALgrTbD9wvyTnvLORLerhsdUGtlZktcbSqAj6dasXnuWclJ1F
5bnpvm+Sfna+c+U0RJxQNc2Xj9zrXVY6VxoKM7OxZyzpBqYtTsvkweQmMz5WAkn3
9yimgCZypqZM6aniWLz+C7CP/pFXurcieCQcvIAnQu4qqco4qvRY1T6+ZIsLfuou
6fyr2N1b6mgAAND4HlJelQcXB9ViBYj7jAN2gj/KVM/OPWbm7hz56OYvoxBwQBWY
mt5naGS8qfpqpfOZ+vTx4O+QLg9cBdTK0fXu6pkFpICt5ogAB8dNxg5Bf6wRwCZr
aOIXLGcb7EDIoLA8dWtoHYeIXjCTzN7yau0VVYzCRKsFYX9RqGxTnlS00xk1A7IH
N73kbUUbk9oY0fd+JraWejE20CShacQXM4OuwhVD8bOO9IEqc1WO6Xst/PZ+4fke
+mODodjuIIv2bM4cYR2DoDTWCI/wiMm9Gn7sdmGf8PLotG+JQSacE6jAvrKeA3nJ
D8yTsmcg4B5QXsUq/E5oWuNc0f4ORdu7WwIyzZpnRG3i0qlGOs7rtCewf5Xa6npu
XintgLZ7Vetk4Zwm7pGjpyx1VlGAyGFzvdXPa5hMyvejWrmQhlVLx8Hb9DJwjPmB
kdQxEYRchbeAOnHTjG10w4pqcEp1H4OO7qMJPfzxrPdUNaH5i+jvUQdbwkziNxwK
CZA7zMpva4YlIz193tPCWexBfIlRj4B1JjigurGIOK9ZvK+9J/6SZAko/fUH6Ag0
0BYyJ1TGyudDsU5fYTdnxU1cyFIBOKdjkdCg7Cmb0Ebx/zCQk8nmsPPUKiqrTi3b
R+eRwrdcuDO3Hr+1YpfSyzXLOPuyOchbXtH3+C2jHERcf7WCwlqQYYM7kqb3Hr8l
vFUgoZydyIgeu+d/gE+J3dkWFcx3g5ZmVfLQ7P2fc+qTzmFx4C9EUPziK/yK9prP
H77l3U6ynR7mx1RQmxa01ujWQb04RNaniBzoShs8qSYbHN6SCWuM7yXZ4UIBysxt
sCpTPYR/7ubYFTslGcm/s4JNlJSbpz6RPKYoZmKzC+UNRkT59KfxtwJlioHDmNUX
tYpd1lRZxhoFKg7IhJBr0H3PgRrNHVBpDWcgsjCeb2Smnr9Sco5dM/TaoOVDK4Ys
VuZifx8sXwGqOufaDZzn3LuFE2auSTjfpTePE1Nj/tWJ9k1tXZr6kr5zL3ibkrNI
rVoLyl0PzBHJdSBSrJWPfWD95JYxqxHxbSQpgWmptZDuDzcGaOavEnjZFZdyEEzu
qfWOUNvHPNSRhxhDSx6qEu4dqC/M9ZfrguDgDhNvc2S72ZwR6DBEOnXr+MPQb6Fh
AOsjY7ti3dyZU0sPLoR7gsBU3BvhaMD0HeFSPgOU+cG4rSuvgR14ZnmQDr+bkgZ+
wPVXi1MFxA4bRZrO1CcsVI9QQ9WyfPhfgKy2qnPCc2vzmdOHZBHmqeALp3Jnd8BN
vKmFRMtYlhZy22odbCxyB1ydRQwb564AK9Vnoguxpbx3mddfZ+L2Mhvzsw/AOyBe
zqPHVADROYpe9XelTJbSwkb53pqzptAwxQ+BOmnmNIqBBiSS3YttjJkhvrXw3uXA
CoejyjBSJaZMMrAdf3tAo6RvSorh3Tq/ZVjcU6kA2RYHHdhq1CSc8uEW9yxBmc++
cuj/3xNIi3/xp2izNKT2E+GrYoTMqmKQneXXZAWiOXFJbYqRvwiDABGC7dvtR1se
lJzT7lQpiEzY60BybtKW2XCrOSsGYH/bV0nvO8fPESoJ4yGcQNp+YD+5JL8wS5Uf
k6uzAf3l4IKx5JM/klHDvQi+zc7MfC/fryuXxWEqgtiN+DWZoJ6+mDVSyKH7hJCM
5W7Wj/w+bdprVdzir5jqxVVPxQ414PiBUoZWhA+pzaV0zQh7wLLNRO5H/hzH5CC0
jRFeH8yA9Z2Bcu4FNx7s6njuick6VvomHs2aYt9VIyAtCQ/SPizGYTGb7Q2PnQc+
8/x6z9JCz4Djm13rSdL3BbQommpRIV6zO1rLJluRoY4mtb+EDSJPIYXLBQI9stRt
q/SV+zNesS3BCI8eKSBPKtAxzg4xIq6s7PSH8APvhdRj9dZm3PyWaMMfXLIW8C1J
EQK4mcmiykKZnzq347sNWO+d9Ds6vgAYQIe5MBIa2JotatowTg6TGTq4YlBjJfTK
TAwRIkzizv3P+xfu94bKRON6kkOCPALjEXvb7yXMQWjoGJX/UGNR4g/evwhUo2+B
9zW++wtMky9WtEu7H1rDyy54C+UAmqmVPmleiYKdKwXRXsv6arOoMCBdDlSo8gTS
AoYxe8oc0RrNZ+tRWwNstbc2t7kagZepsyDcldDfJAm1qpBzo6nupWA6Ls4njpP0
FnjLtt35yLiBH1zlahu9t0uKtvi+3O7dESUS+1gLwHe8RPe+Dr46kCxsLMmfoqQX
oHclBO+fBHgsHl5QTOTbCKb2+OIX1oXiLYIhsH5rI7zOiH6uFgBCtTwBy3xK0RJF
s9SrKsLMp7OwAwQ08YDX75E/w1seLhh0aLTU2lSCjnLmBtTB95lDxdUczoGV1XBI
J3vh/GPR3zKvkVoa7eJndtwFMOricvXjqDkwDN4//X+QhJFMZo0p0nnPWukEYGbw
3MBiwjpEb8cy8o/E3H1b4S8emfH7M0lEWZ5xIj9lY+wRmwOAWd7jeLwoLI+v/NVk
lkWGhXVMDxga8XqSCJrtArJ128xbwCmJrXSOMh6Ihs9AHNSrU3sMffru+CvPRF4N
FVMKbeZzSPYZHxtbofzL6H6DKWau9jH4eLlllR6V+7uEbyweVZxrVHOTQjTSj9sO
G4jVDunnphtsYHyvXBSAj0FMtNKkj2N3RVQdpIUIBSWSXuaPQaoYoSDgtvMixbov
w+43WWKqHd6hikUjSCIi5AeZ2t6CTORkPwL4JTWct7ZOeQhm95Pj/bTC905ulr+V
aWb5l4nAly3vnT96NNXtsFcso+SRqK1Q10Y2gfFAch5DXQYfp841gD0jT4V4J8f/
aTPSYG8oqp9Bu5Sc9JlgMiYCuGdJjG5HIdFdxg8BuaZxWAj9y558rSc8XwbyYdtP
hyTT3qw8qy7UjEOmeqrw8xq+9yxrHM5IGCng4W8R25j3UgjjuXA7D/Y0wZa0ABCR
SRZtsLeeTfjBKkZL2Lh9R3Qo298AjgXGPJfqXM+8QV7s0nJCWCL3RSVQCBCU/oHu
m/nLngFKK5gRxADo3LDU8z102gpD19FKCPQ3ONJk0ULV/3KokmrN3yHx3wYMVk1M
85++/RpW6Xc1sUMYZOH89CjA7xzveqfdOm2BHG6+rvvC03PKJ6xvwqlfSZBoBPgN
oPMv41hMF1nLlFDWwgo3qa41iIYCb5VJ18NUo9Q/AEtA7680F24l0gYxKDtSoP45
vkRKRDGAxx8SvlSswkLL98Ycd3DzCrR9X80qSxXHnF5wAYHXFV5BIhLzzzDoHbWW
bi9lc3B/f3LGvcvakwT3UMhr6oXtCf3tpc8b6t2bhTuUD92oncE6p+FBuDkmbGUP
/7M8bg7k2NaiOu9s3qSeMF0bnPo+EyH+aROs5Qdy+D7fbP/uREYAGSD33HWhrtGH
l5tLoc1mLiL+Ssaw8dlX0jffgd31nnyiDSPTnAwYpjnpcCUOv2NK599g3R1gnLhV
UVLP1D16XgOeuMCiQIeQHNLAaponxzuvlBw8snNZyqarfn5u9vmy1uKdRtWIVzYD
t+kVVPiCIu8B4oku1SNihbzrZnQx9/Rk2dKXYhaFOwckCnOrAJgeUqHbn8md9lfh
xzZxsJNDOc0yzgu+Bv69NeVTn/Mf2Y33mOt8OlwKCqxrYZM/PNprb8KO2XGk/dj/
WTeN2Bsj5TjL2Ja2PFjX6gG8dOlNIgigMw0xHyVfTBiTnZZ/imCFPQBfrS69HBQT
rwSwOG9h8sQ5BsXmjH+MjC5+J4Hs+hIMJ1W0lQ7buU+55B5vAu4+aClofM1yqvFm
opM/cEwQ60Ccx7IwQTHuOTSKS/nlOtHCJw3bzR3/3739WjpiW04bHZZTCAoXHcl1
zzQwpV9gvSjip6wcF5jZzxZTN1Xih2wI5z8jR7HBh5DEAhvQqnHPXKVpVXJRFrKE
re4nQZDxVdUtJcJNm4ODsBD3REnp5KW9Gth8gqhN6+0RiK5oFjGCQKN7p70ClTxZ
7U1k8fiGAMjO1H6ovBqJA7yUEHrxLW5kW1M97KHBag6p1RvraUzWMdpg+u4Qzir8
5fQIqb2g8jCvavqSgx9eUYhqHL3XPGlbEQAayJZVWbRBsOUhvkSOZvW5zH1PEvnP
bgI55JU2JoNPrpyg7DY85NVPIJVkliysVrPV5w29l66M0MQsO0x7yzDNyAAmycDW
6ob0Uazt3D5tyRyT8kvaFE5Ldla9/EdU3AcMEG5+kaiJHUGkeU7DEuUhIz9QlGuk
EqfeR2UhR89JUA+FG52H/Yo1pXEmA4MR67cY3Zzog8/Kt7p+kV/bqq9/G0MUnSnC
ePlyCzZsEPdMpcVbPehvCGvPgsu3rhzd5HdjCmFXx4N8R+SHrdwgxvzekx2aqHN4
jHPwm47ZAwW0ACI+cAY00TMvtFVoS3fLtoEnf+BbCWz1tXbgWxVn0YF7xGicir4T
M2MC38AXP1yNZEaWl8dwjkGOlinz1ISFxwKjF5fTIO5FZ0s3tngnHBE5KSxvxEld
sWp3nWUnCv8tF5ES1MMpPemHB+3u9+ZaHZD0DX9aFKu5vA1vzdgti9B9ba6fyqkN
NzN27zzqYEbtXtpL7DLk+O/+sA57UgRba5utZ947oDJu/+do54SBeejYjAKMvtd6
jFso4PMZAwYJqTK+zIDB//m5adRtTOqe9ukzbXE8i+12BPMqhHnEeITB2ZS1eVEX
dwO+etj0pbZFurHYoW3mOk/bdRySpk0vkx2wpW0RLI5uMH98zvd9sPTAO0oJVs+n
XyVvQGmMlyy4tgy1R9DcXaLTR9DBnlaJeMOK+0ueB+WP5nPau5V3FOTt9D00ZLzk
8Xmz5dH+C/y70BoO2jnQsH+YPQoVobCwoCXAMb691mNI2WKHNccxNb0eKnByAra/
YXjLNSPCD8O5In9jQNyihasGg45g6wDSGsdBI8fAqigCYcVjj4RHRT7ey7PIEQBI
JrsS6Ya1DBdqBevCe8j46tS774AcAj2el4/HUdG8x177uQfYtHZsfpQD2jiw077o
frgm97NI2sSAK6cXDf/erdciy3/6qhAJQ3nh+Uh7soS9Bkb8T0l8dGK55Or5hbLs
Nq0iNOhhJJx4ymlM2HFpp5HsJAVDEbko+42BvqH06cDXFZrKmD3IwGhXOTtAbcb0
Ky99xo9CLvdUpct1HsTn3xkYkNsFIxz8C+5GHz9ZBQ2vFQYtrdOMGLappcIzdxQR
1kirBbAVaKvLqY4KoAJQg1OIM9jEVwr1Z7VBsC/20dS9J25UVcd4AAEW8rlCvpCV
4XCND2Thf3pqpzFIdxz5ZdICzNpBe2ZUmw6OtUZmgIuyQcfRSEsPuivBjBCdSExU
NtPN4fAVa0Zngc/qveaDg1hp6gMOVuLK92yLPFjSpnxBqwoDD8GhRSGOBX7quaQW
EbYz5xECM+mOBDV6CWKlOpL+LtBgeJuduk4d3QtqKhc3H/gWTGXgBLSwTleQyd9a
fhiIWnr7KCcrTBF0jHnSVSd0Edhd75ajw1LmVcISeKLQGjv/P7inBj2H1ES2rLnt
wDbM4uYW7lPZM0Ds2UO3Htirr516LPrS0DaMFgXnUQyszmPp2ugaMYm3Fuhxbw9s
gl2kuETC03Es2F25H/tJwmYgXH3XdcRMYsl+LVwsr+y+FTBh8zjpR+0HTtThBGUO
zHb6h9SDSLGYhXJe5AansSikyBoYbn5fyhnuS3P3058CYYf3CukyMxgbV/NmCdSS
Szod8XCv0UaFjffTEwm4G+RZN3Y2TVPEoi2DNC7BWjasXu9VSExK20u8vHb5euj5
WejIcQVTjsqMLpbJRY24LujABc0HRqYCZXByusURimCbrCpiMIsbcRTW9/u8cPdj
r2Pej0ycgyBHYhjDzjvL4jNdhCl9VDFiHb+H4R2fyu2cQJRY5C6EgbkJyq99LVx7
p+nVVv3AA/LGA6x69BWRbmbGBBaMbrEHjVn/8lb69EZzZq5449vM8c4lNXI0HpYK
a/k5tCRe+kWboMj+PNbbv6070s6xcD0H/22NqCy5yvSOgmM3sxfgk4xkyEp+URuP
DMVnu1/vKYhUW7BpnzTKjl9tOznwKIpy+ZhTjodIReGohH3o63xD6VZWSHdU3gf2
+p935V9KC6M8hLlRCuTi4HtsUw9hL1mAlPccxWHKtUg7vSgNtCrevx+W5yZsf/oQ
Wnu06ikbMNssHN6ddrfNI79+FR/9MYjsd+pJgyC67BEP2HC6hCBKZxE3NFiVIjW/
fLZUZ67wEqil0hqV3pBtXd0apBxywUPS0X6w4OtM9wPqLHBoLaWvmV4Q2kadzsCj
O8s9egdw4+EU7sd7m2wSMrb4uqe4RVjANZbSHznNfXXUqMm2wgrD5geqSf8s2vzf
mh3KzoNc7OhXn33HeWeHnWjwmMSpcTaIEvNSDOseUqoDP5jG9u5lxiHNhgxv2w9N
vDGVIUKkbJz0ND73Fb7HNu2dkT9/+MbkpQozngY8vz3SwkYI7awWeiBkSOaCVdp+
vzKvQNMItOb3qodr088ohoukwWiiWQtGap09RcipVoFi+MrB8A/ZPjiw1aKL2V9d
1iGO8I/1jn0rjcIpLBGjIzBv1Cc7dvnEI1kKbg0bkjHSOEsVifPmf+VrMnq4W1Hb
1LBUpJbuGQoNuzl9wdPeTBsbHcv5+elP5KgPcHxUNbFkH+apngDL16p81tp5s2tO
/7Dk7r8swM2LlOXiejOrKrcoYzsRUpi+sZMAWTXX/7ti4watQLjRM7sr1pefZk/j
LoqPEdD3eTUBQgHRKehmbGmnWqZKmepOd5UbNunLLME2AqxI9zER6EqAJ2U0BEqD
P5MfOEFY7b0BbF3Lfs4stu23JcOlJQr8CBTIpBS064rbUaMFLePrJ9Sktl0Ept/J
ilfVV5tvtx+MzqM5seGQTnFNfVOuEgAAwfD1Nit+VwlGotAmQ/wdTCtwy9m5mgV7
VIpXobbQxJNpEV4KYtF1cQA1WvNT/e+9NTIQ42N+d1HPkxCNW24Xsb0KiJnc7JVj
xzK8PX6aKyoj93Nb+KaTiRlQjfPMudwnv3fxK1ZUqMD8sZnIc7qgkdlQh26u7UvI
XhBG27veouDE8aBqv+4PS+Ihg5iG7lQvrjZkBusdPXoFEOajmIG/dKOkY/wGKH5c
I3Hi1hK0hTnHBIzJnpyaE/VWLoahbCA4O0l9JiIZG3CiHxQeQagJE4wXSbF603My
lKXVxyOcdMcN/COO0I0DQXum9QHjG1jkUj0WrsgIedhJFcBXC+qwLZsHRAHvj//L
nBv03oVJ8HTLgVqqjVbLNgMVdkSfA/WqKnp7ssnhHzVa1QX4Pmu2nqg/z+9PhNbE
cPzJ3KFP+mH6jCCClwPsfp0aoenn+/PAFqAEZ9VQ64XQNLxoWTx7UwcQt911zCps
Q9JOAu5RpjqHnKYETOnp1L7lqbhv9l5CsI/T+ApTS1wwE8+kpnP2x049F5V/h0xI
jVsV01SJDkKdWU5JELKE6+PpqqVE3TUt5fholBZNaqawvFYTeNi6/PEMCGTCL2Am
TF0YowzF64Gc2jGVhRzHbae4+opE3G41zszM5sYzeOfu2navDzeetacjnJ8LV6bm
seOXwyvTPMh+TKq5dJwKHoeNaQPL1BHY3IRwZCXXFlAuptO/5MeahQUB1rsX3CBu
kZOEc5lpqy1EaJbcmpDqyQgfnDVtHeap44l9W/LbvGkJlqQcZrpX98iWmfduHzG6
iIwo0owImpqLLrm+zFcgFW6sDVdPK2G7VzcOdeEPXJrfc9cfr0gx5WOfl/NnfTnF
mSCmicy9EJfcTIUCKaUHBdMjt806VP2EFKNGui5qX3gt5kj0qPA7U84Kky/wnHLa
Sv77zKG9F2bM4gy6eescZWpus975rbOgh2b9dho6k4MMmLXvXagDSKvVBtlSTO7D
2d1KZV7anEKEGuqtFC/G3dAtnryvCdfP7aihOV0Rt24BG7H/iMlKXd1AsxA/ALx6
NQnCfYwmVz2Z3DgUJWfyhpiMc0YbjIhN8wwkeate49ZhWecb9NjsYXzrJ4OhhthS
/R9eTNhy+VhZgaZrV41nP/fhJtAPuvxlmD6t9llDhXlUiXNQk51gN4TyUROwJ/EO
Zwj0Fv1WIwaLZ7Nx+E/5Pj8SGYwKgjeXoMaaR0uHb+xC8XwOFiuUm0yLud9nQkUy
n5duhFtk4ogbblu1Z0fGsWN4FaxwMeJ+D7gqZ6qj/9pGX3eAB8tG4TJoG6OOIPnc
En3AOnNeRvDbot0Qsfv98PsYORLLdPLwz8/cSof+IvQzqzqIy0CV3CG9hTHuZoCh
aSn0HLtqsYVCIYOFSkT5YqJmNPAbt1SqV5hSGMenHIf8GZUfJfLlVwCxr67g+Ggt
3aLoDYVdUEZ8PtppHg+BoegReTZsmpTy5A7AXamSUs5bBU0E1G0KBPP4/t+BtgrW
iIGjEGuv8H5EN0tQd1i1pudvyjpGKXpBTyGF3CPasIEoNapcMu6rMZdslt05z5Mx
C/lshiC4aLMIzZvKw/8hMVdp8Qg+CUoNm1WtXlT9mp9rg7abqVbOguxcAycuyzZw
qzDkfpvUEEa9b3Qdh9h4I1JH4+6ZN7I0soNvpDWnvJCWTI5OowFzFBr1mAFxpBqq
08t4FDboUcQM0WiBRQ1kzGavwe6SPZh4QdS+xO3XdfSa4r/1A9PKsP84kOaGxU8M
/6qhBTfmSnuAaVeDei2ZNIt4VYuTrwOlD+83IvPmIyLXCIJmQXiJ0R0AE7dq/wRK
IUYOjaYD+wefs32uihWMtdwdDXl7+uPXdEUqEUafbTvuHzWmaWzELL5ZcPHROk+P
8MI83YO/H5TMHJhYo+wns767zDrmYV+PomXZt4cWjTQeevNFvG4hxeYtklRh9Zxp
FgJXKM0NaG1JpotLmaw9CXCVGFYi9nsvfO3+P+oGrRx93OehdIgZSnKDxFDTB2ZC
lUGzj/i7JTAMeq1Xh8OuwVc0Bw4x/Iqmq+71KodhGF2w8wFQX+mvpKLFttLiLISO
zmso4LhL0sY/w+abMBq6wc9mR7Y8M8RHklmgXMJVQGBiKJcHAksMBZDFJC1jL6sr
NNtOW8e9mJYZ/K0S4CnwmlY6oKftHB5Edbaang9vh7kTO2gCAnWT9TP+cwbk9Z4+
HP1DC7xwSK+LXqxjDjxcINaU5r2/whzl5CKCmkcOXI/tNN7urOoKsk3LM7MNnyIK
pcKH2VMF+sabBblha5rYxTZnPw3brNucXgP2L4KjZy30lnez6rC/UvANZtFHV2Dp
kHfCeBr7TL6exQ4IcwWajj3vSHXndHOpiKV5tVvWoVce46m7/RhJXm60f5nIg+l6
23Ch7UxZxKpVxwCG+Nj4GqUtqeNDNGza/OkB4U1dBwkujl+QEhRwJMRsRPTAYMxf
NhPUnoNW3DtYcW2qypG5XwfNAqWdPn2tG/KAnip3Z0ZTBPeqtC79Ul9Z5qEea1NC
0FmFPAvMhA4YM1G2mCmRK0gB/CxGFSE9hzyLt1ZwvR4sbAdv26JShMILF16GsIT6
YOWCdZtCxKDxqMLRDnZ0D0GnVAKo6ItwwxW8lu9hKYrcZFXwIlqzafT4n9MH87HB
4eHS2k7HVEj1D10YyDhYZh5SfONchxqh+6xME8+nvBVeCicjAsPM1ETBApQputHF
kNFcHTvHI48AA36X10PdK+RPX3H0QVJ1QW0ffDFmejwCjW4Y08Jg1mMJHlE5Ua81
rb3DV825plmU7jc70E+YWNft4/XJCKXg6AratlYFMd3a5lgkjPqMeHTD8/+ChNo8
CKnyoqsr2u0uQDibKGdGSvdQndKKI2PjIZeqXbV71hPKGEuSYHhMOXx5N1DAnOIH
Q+V7FgeLl/pFGNfqCaGVSruTrA/7M+6E4kaqPFSebdznh23PZbpXh3coReBrNio8
50jZHztd+NXFTGSlU4K5KDGLXv4fdionsf4AODcg4mx9wiULnvMO4NnFMn/teVpE
SIIu+M248w0Rz//LZJ/Amkm0KzsZUJNJHjnPAIrxVxog2sABUK+xUDVRbtQu3hVf
a4Pm+bRl8Mgp9PVuoWdgf3ojWNjqJRWBF2JT1/c9XZZsUmh1PL+uba52/xWoqPcq
OnHEhuQNdMJrRQIgjdwgX2ug6C2QGw1hjNR7r4GYG4YOlP1G7aqPhK3YU25PXXIr
eWSPXS5UrK8zJZz7yH7MWYqXcQW9SSLWVpR8+2aZNnnav8qJm6S8WK03X5VtvczZ
QBSjNdQkx6hWvL3W1PjqgN/EfCjDQywX9LKucfzTG5xP7r743ToUszSpEscp6QNk
2pr+0B3Cy2nU2cekrJJMYdYSvJ1tclES7L5c+npEt9KHQRq3dQ8KZQGTyQGvwbg0
eltXSrL/fEXxxdD5VV2n0ZrKTo9CiAVW6jbBCIVaRzYgPTYGR8+b8vHkW8k+w0nT
ZtYTntKT6uHmQ7DlSt5Bd32cTYLRlH7wwZqBpFv2T8/UavGQ3iJNdOou6Gtatnv6
46oT8hSBbM9gDuy6rUj4121BkITdtro42Qd/0cjOWBEuC7v7WzjbQdm33RDuOC+9
AlwwdOnrCBX9IyuQYv+UOSGoQTunvHhrgL1t2ErU+H83gQ3HYEfvWZraZujQJH8Z
q7jf5CE/YRdah72QKTBhHHWpAS65ZkEBLEop8gprKdfMWqsGogP3+HOQEzy3XaDA
/739akas7G7frG/DhLJMk+ffY60TluLI5aWg67ZFpdqda4Zi54zzwnYnjulvquOl
5WL7B6H/pHm5YzIKrlq443xSNZQMNttu435tNPrnQSX8ty+G2a8Cf2eYJTMB0giD
FZUCCI7AVz5JCn4mixccQoG1ws4DM3thRxKA3GwX9TI1TsZnJ4qDGKihygB5Hzpv
MM2Y+rrylnlmZ5e0VS1Y5oKPK5xwZ0WCnpyZu9N/JDp2VzSbNu0mqB+OlGx53UnF
/NcUN0TgmYIf1JtAFFGtXdcq2SuZUaq2Mg2y4PEaPXp0+H0/2le8RjZqiwYzcwbP
8g7dxSqMmhEnQFeaM4jw0o0r8j0nxCByq1RznGUfCBLW2vs6yzph8h1rkp+q7md0
i1qsG1z0Q4k9GI3fMIn2Z25tZmZi3VyCS/hDgAQF0VkzguFb93bsF9oh2hcsTb5x
mbKXcsClKeMggplqB4PzcdTFeiZ+ulE6AAbIPsalrZzFf08nJK2PBk+n/WAW5hRa
8rjxFLhGffcBLc0B9bgTd5iInCbLQEQXpmFeB2zPZKEcNSaBqEWp8yzx1CV8teDs
3CH+2hJP4+E7fnSr+gVIYK8zj/GerHVI+4I2FuUkeZCiffIVcHN1KoQJo8F5X7go
ouJJ+A7pVoLGD0sdlUqLDOKcIa4C9N6VGsxJpm1EthN9IVDK/cZBS9eIg0waiG1C
VRsCRe4qfrdD6N8DZNyc7U1znDHD19y9sEhBvRSOAhO0gqAM9rKhMgGV8kY1uL9f
8Ap+P0wcWHZTBmSmLTQtt3zyYUXhqfHhQm2TNPd6CZZmsFt9wCJ4D1f04XoVVYS7
1GLvjxNnltMW0fnKLvk/Ij8FdvY2xWhJ7eM6Qn63dHVM/tYhUOogCksGK8Na1+k6
rpAzUdsApK5ZeAZOF40L+BPaPIjwM4a7smJxlnX7dd0bJNw5SOcaYtrosNj7D0q8
O0kr8SNFdV99wuyMpxsJtRMzosL+oACaaP3s4nN79m71xSN2tHrRMW76leYwJXDE
cFch2kf+mjoKGkTPS2oZ9YGyAOjK62RonAxDqG5XEshYQVALrduC2mYCXEqA2wfn
grPxCK2mQewJPpgRk+ZFT44sF7pTnrXmapBTnx9XhD4IXLGGaBql9rxeSkOrbTEO
P8pGmnVsv1Cp1HP3p25gKdoVK8r0gaxHAY2XbO7puy69383Xkks64JxB7OCBrh40
L9BstjcbbDnRLz8CGDfAwNGyNINGQFFmGLU5YejuRfc3t43dk0iHywXlUdxPkNQd
3FLfrYEw42NcSLJ7oDuzvcYikPsvzauxqRcJ971PKcyXinnAPwsOSd65rG73JWdX
qVNwe3dZkIpgyTAKjyaxoQA82PBbcBlQHqisaK3nXncm/KEjzYnS//USND2VnU4e
a+SVCvHkYVIp8MkzyRYRe3YUEXFTiS9QpTzgfHZHaOHSG2gj8n00NlH5hj6x3Jm/
1zdGHWZlvuhkPXwUi4DPQY3oT0/3uw0egMDys7HYMbwNORyq0UYmmfB9nO0vCQth
5xVbb8Z49BC4os3XPnhiw0sT8VE1kU1Pgb7yq9lzRNsfoxHf2QWfkwqs11hfRkbG
E6jmN9HRb3QobpDze+mu60hyZaSwS0WRUuMk3olIsQGs1lJ2LYHMnhfDI2QGvpwR
YYotMy8weNfiLz/WAPdTUvWA6MvVjz3vn0uB4DvRNA8gTjLKizKgpFHow69wMypf
mGcQjk6rBrfdslcYCRYJV4Dv61RjWIoniDgHV2d11qKz4Z2KRymuwA6A4mdGbHGg
PsxKjNdSnetpDghG2la8xgwuzbHa+0Gijoa0Jw7iWp3cgwy2eEXGrGl84XJtnlLd
HHvRBEStV7O5rFzV5o9H8vGkCuZup+eXPcOTIjU4vde3ZHIhn4po21+hkTmOZ/aG
kEGmq3r/hnyuxhW0EKW+zHsGHnTF/czXO95D4uA0esMmMxTjL3NGljI9MHzYCFhk
g3RU345aYC/vMizdUjPDZTYKuT2CpzxGqThJqHfMsNnWYLF0KaybQb2C5SvxhPlb
A7CUAoA6j8zzb4s7+NTgcfF3P5tIxsYy8/EsqYDd8YwG+iBqmJbn2uGH07pw1OVh
9NxmCSVMT8vDNURpWYYUmVtqklZMmHQO23E4suutv3dByiBSkfEDSO2ZJCUWmZlg
aSS+P2oR0UJYklL6TI3YLT9ijdQFnpC5ST5YFVGL2/EDYMvIsuCQdb+dLITSZDsU
9QGHFlTiadZYYQyGzuYLwz6zBz64edYmLLCst2ubDh417Jzcz5gvqXYCKGo+0Ehq
bZ2DC06X2PXebnZ2nCy7fO2cr+8VZ+tR0CIWB+rse0hH7iOQ3q1N74xPd9W25/Ls
fhu4sKQsx3pZCh9zec3vHHoZpVJe13PrAEa/Of4/UTZ5wWUt2+7SJfe1wlio9Sjn
Xl7rRAYRaMznqsLTBZ793NDsqAZSlsF3vHCKhNSsHFvhzO3kp5h3woePZnl0J7BS
kP8q4VN/GDgh6ugTOLUJIq5SuZZkXyge7iEXfK2EaU5eU7tJVCGU+XsGkH+4veXI
RA4FtW4gQke7oBbeui5Tj5scI1ovWtPdrfgxARRoj1Q2quFJ6aY6tkXJSYu5HGE8
smPO2RxkRCD9bPHRhpEncaHann8XiE6de53kyrUmY4WQCwo1z28wEufUwRTOJ/3A
xcXS2Z3CqWGcMir6X4CVC27mGlAT8O6SVq2CsVymU7x+HMKzR5KlUb00ZtHlCvcw
ZataM1NfO+Bzx8xnZnEYnp7PESCeO2VnG8WHlpyMPcKS7lZxn8siSUxjOOn3RdFG
oZ2IRyJ2y2VZSbrWFA75/N56NbQ6YuO5Htt7Osib9XUfgiA2nj5HMK+/gr20Ifn4
4RwBZtIt7HwmVe3InQJ8E4KJrgF9ENle69Yfw9b8jTdwFR5N7cX/8kC9elOtb9z/
pwU+G/AWX+v6oPgAYjXfkCt30AN/O7lq3Cyhb6/oTHXHCY7LyakrZ/NbQKZBS7Vw
F+5eVw+vFv8QpGDyT+6YzLvkY7Ptoi7dJo7A2d+DsIBRNFEQMLnLJr6tD4bM6TKZ
dH5F4qF5pevgGAmSCHDIqO9DnRSCWd1FI69UIflSOe9gM1/vZYdbPta4rZ0W1kHX
Jiy2KNslWIcV92pjPZ9vvfkOZEddfeVdPT2s/r/JqtAy/8wsHerNcHy/amxVnlP7
ri9l4djTPuekZd5LFl4KTsW/RHvFLkoNO9N5r6r/uIEl0tSFskUSVLyo8bVi7FY5
US3lDdL1YskWfKjxS01uN92WXrbeQF507yOC1eNKLa/if+kTwJ96H2ra1+s4NDYU
cSMMJIncwWozSLFg4VbMmS3YDa6QdRYHIAB6vywwIfJA9ekL84wZZisPYfDwq2g9
eQvntLLhtfsmkD1/E3tc4JI1+DYzOFZExTApJmyqnoi2/2pY0/juqUX1tx4pmZH5
lDAVY84XRSLsSVgZ+HGT88kXB+2c8Fy892XiIkxK4sUh+PiKxKwg5Kk5BsOJ8XV0
xYbPdSxa0qbhP9dh57SGVxU4YtDozB48xtifA14c1Q6OgrcktSvkS0Li85/NX8hc
145wsxajYFKx3UCjvmReetiMfcCQdcKY2zX+j4wG5Bt92Vsimaq8SYyWXjNxKWnQ
6zSLjQsool/ww4khz8/jl5IqIdu4M7TcXqkR9C26OwtGOEG6x11tfD8zXg5PqcoV
VR86bko5g2iStKhSb/MsL8r3rUwV4MJDpE9R1hsF5QFjV315+dMae3cupPumhQPa
Cyab7mcJuWZyRYwxn9cw0Ln2eO9/y+3dr+8c74aizcLbQpvktQ8ryt5/FHiP1xPS
/MrzXVi5bS3LPx9oncckv/caZp0f3FW0oBoxO70QNqD8P+EUVB0nBGvS4LvcsEmh
02Knsx3VNCio7tQKFYX+0YAfnqsZW3F2xLZUE6pMgEm5wssFNPSQSUCn6ERHq9av
tvkzU7B6JsXoW4YZRMyj3eLWeBV8ctn6/PznPyZ5Mjto62VhwEtap71fzEa8l2Ny
pa7I4SDKAPFXd5nte5kjsSwf6JAS1lyqsCTLnuAoGcEGfYm24XkROy0ary8KCIPP
WbFjMtSKqmP0VWbcIDGbEwa+Es7qJ3mfeMVgm3wnmlbewfuQ6MTP0Ad7vl/6Y4YA
SP9bVGeaZWn7JWDdNcQst01G5zOT3/ysLHwX30nEpOTMO1p7H7N3G/wxbGLgdO+S
tNUqoCCBcTW8w7OyPT5Dk86piCQO0ndTJSFCnj4SFrNUZa0PmDTc2lRDicKJEF3p
S3mKywjKx75bMZo3Cxbj0ESr1j6a92IaGRjrrf1WHlKlcNQl2M0v0p4MIgRsbnqU
Og2UA+AGaSRX0WgFVWGchO36VStgTUOf3xlcoHx8aBkdNB31hctfv8njbmKvOacM
p71+x3SgwBnZHQBMnaPOxY3U1TToxeiwLiJOKZa5Pu09uZYy0okkJOgcw7x5L+hB
g1fEvHlBD1oaQ2OzVDC0R7uLHni0X3l/Zl4fb9V53EE3/JVb38qjxvDA4C7sODsS
01GoJwLdxI2v+lMbezqQXDFha61iYSrpkGJvqfGBCtWPxf0C4buFRt4wcf4qd4+U
eStm8BpBTnQb4taxffM+ag6dad+IHe5hpTJnbN49cs5kjMFP9CNKOIXwCKQz1dU5
A+2v2jo+r/nciVuvyGGJLsctuSW80r5cLLNcweK30HDEzcVlMYcRuJRZndxKJDe3
u7OC4VD2Ri3l439HwhGW9+xzB32dOmSYyH0sBff5EzTz0w+/6XUusKj2WP+1n/4V
TxH+z3FGWHv39Hhi1V4sjKrJ04y9WzApeWMEzpPcVJkBVMyOKCMpFOns0iPgnLvk
NCeXOGUYrEJC07Wlq49+bHKxmV/hwk2EVMYuFLRijFAdGIVbUlkWcgVp0AbR7ZMx
msGd4upihuBJqU/qyPYBaR2xj8NAc3vgEjrU7KarSUjfPaJv5YX4b1pGYjIS+0o9
gbqXCpb3tQf7pOhVoUyVqnjFJaVpTn8eL7VRnPoUpGSH+sZZ7yU2AGlCRhjDlzrK
W7Qd5w0QVh1rHTw+LYHNb85T6rHebK7X85gNb7wZ6wZnrD2Dwrd9xwEKT6dlQS0U
9p7erY0tVqoepxzynl86g9xga1rcI11FIf93TJ39xQk0oa3jMhd4sX6C2U20F6zD
z98ORfpd77BFNylv8SiyNMKmUPsOJuf1ZVc7nLldtrKx0PtmQZ7dVTGsGkcNoxKh
9zmlNoE0vVp27GzoEnVtBDN1gZCRfasAIGoVYOqYhygfvm+uqZvabaN/Uci2bvbR
Tzi8yrwnDnIg60Sf9v2vwPab7ophzz2MuGfSv3j50H7wNWhA+oGI9J5ejk7mUMPJ
04ez7pj9+54QG8i+I3SDJZ1Mn1dGP+dfBQwxD1AzIYIPn8fz2u1DRsXigVM914SW
OeMYd5oqoZtUDdOOdtjtR4iPoD5HCgeTN/CuafCOrz2tcffXhn/CkF8qa3oIIWnK
BTkCTJYLXTO954h+Rpcl1VSvtC8VMGROd4g3GiFbIxBYEgRr+yPGY6944/+WG4ds
Srb6xfj5L2wICLF8w3UuBx/k2QKakJRvTu0Bo5ItWgzDUF3in8yN5TNQKmwZ3i/d
koPiHtCASwWyhJI8z7DDRY2gK37ModGJuRL0J7DqWj2PibTTEsgwlqEogMdqdvPp
lrV3SmI+yqwn2v2QnZjrswFuujzkq+/ME91PLAn8tw4QAe0ghMYj32+JRMyR/ou5
dNiR3PPY2IjhgAkPXtYZQk6Ko6X84obVuX2vE1YOkJfKeCpIh/0quO3nxorpJybP
t5kZJ6v8h2KrT4KnYpfvSciE8WUlt/YO8/6lBIcHqxHHZ2Yl2F1OIW7jkDeukBIS
A8LjxBCAQsKyuaurNAJyda7GrdD5/sWj73r+nNH1Y8E4T3r2eSQwoKZB/4D6UlXZ
qv5MiL85vidZZIsd8sca7rTeIUF8Orh9a9xnTxH3WF4LYdRRlCaIwB6SP5c9pwTC
h7SqTuAcsUUGeBRY4HbrOp0CBXc2bn7CNzzJA7xyTNTBlHkyZVQxsUnlyFnw24l6
wYbX2nXbpxrmwKO+jR8bnrvRUxPvcMntCI4RQHg4CjKGr8brMPSRNJ8ihoqFsp6k
iVNGNV92xYyLEO7sliEq6wmHgLp4qu34/HrDZO0sRJqaRJJYa98XhPVuGOEtKPV1
bqpYUoK1unBJWxWlhpDGyX7FU8EXn6aGMqMRakaqs6LqF/dmVtqOXeOuqISXddy0
KQRMEK85AIgkvoVMMxOfjrj2s3jl2J/gw56bDH25328KisLzPJX7RRynAmuPwM+Y
B+gci7p8m0yzUDo1ujeQeZMVuG2y5bLapXceTECGeIbLgWGNuvrvny5w66w/K2sG
l4w2u4g+6QGej4kFYGNiWCpzU1HDNNtWb+9GuiV1bAJQ4301BQXeYS5rMWy85Q31
RVOBPe+KUzOezAD9wqbj+32l5oMA/mBAJr8qFGEVbDlIWCEtjaZcOU+X6EVx8aXN
uQzDjpQlLSoAcM5hrbKNRSyiatn9uQL/pMeCwisvK1lzN/KxRPqZM/lYwGM0v1Yw
kWF7R5jAxlMmBzVjOMz6J9R2BXskEewniH0zoJCl5kW00CQsaOUZjF1jE+6edyAB
ww8vDuqjUpwioOhXmZxJonAHr4Sc03skqpQxowKhUEFcVoh6bBZ3HIgrCHjacPDX
ioIUUbQaDcGRXO/gft4pCvJUNhWHVVS7QLXVYt3Ad6xD/7UDKJ/GqKtSx7t06kyT
8SrVJnJs6TZ4wZJ9ToQx6cjFNPrc9xjVNSxLHDBQmGVZ43jsuAIzlAyjXfSFV261
yXBsubZOI27vXZdlQXYxHwHOAo7x6IvZMQ6Tj0O6IODp7ViJ9pjU/spPRFNqTU8f
k31lyRFUypr46DjMcitmHx9+VBmAaMc1MboG+su5WmX8ioCh2sTch5o9Ot6lMNyX
8GHKQbc23Zyxtutz/ytyEChHHaPR7QN16wCC5/EYSkeX6Bqucuyttl4mjWyyFs9g
1opu51LZH+dnpQCWMZeh02lBDD9OHU31QRf+af2XFyLQJSn1qpG2snHmr/CIMlOH
ztFdDbMQw7qNiDBynUNFFt5aRTt/SVKgWIHCelM5EonHTmQs/80FhEzdIEMb7dTl
UR8EqKHKP2aaY8U/CRds8ZfOf16LhlxN85l2MDGjGfz39r/cOu83VaKEq5HR1zi6
IwhHQea9nS0YJzpBYF3RbyQ5XQnwTznjEusbT0R1Xc2o1cwWAMOO8EwbGu9ROAt1
kcPzQUl1rP5RvDQ6544SPSM+LqmEzoAPYN2To9QXbBsf7/fPlPtklvevCn/nh41b
hdFms8aMml/3aMMkrZCxplyJem28XWm31hrfjgopqKtiddxz41MgeLbV8wD/uYA3
SsIJH3glYahPpfv8KTO9oA4jq0HZi9w403BTnxvHp7wgRbljNKcLXMUDe37lAgk+
P6aB+DPVsLRZ3oNWfaJtgseeaobjR7nKohZczNVR6mLi/L3VEVE/R9HZrKNsTW/J
pHIXjsS69r9+StmZ26vRHsUb4A6BnE+bTJA7yjsZgevjA8tOtqZSQpAGzf+ggTRf
aFu1HUM2MLfcMdtgAw7YWnLy8bd3u8T82JtofpvAPJGTZKDhv5oBQGkxY4utdNKa
Ip4ieftV9CmaA+8EYh+HRA4jenS9j8ZL8t6vBnqEVkIU0hBratXEIqOPIj/AVZc3
Wiy7ZVZJL8lPALeIsWm9pPY9kUZ+wfzGRnDcwMExBPXrmkkSudjFfuCsP4wZRVdT
47GOoQ1evRLEbVedLYHufKJnIOb4TkHdTHaE32lWT7J4gm0ceUEI8ZhCyEmbK5Jj
0ukjFvNkSr/pLVwSJSE+0GRBwFRvhJgC4CKmlypA6u8LssbsNVLSen9QwgqK/I3r
2fdQrBZbh4RFrdr7vkju7ojhomNPdmelkcfkfTSSLFTgdFzGV/XUkieZAvYa4pV7
w2MDokxztbc4C+HKd48qhc+H4xPDjH0RQe+FU9JPS7hIytIOjXyWg37/PS1aZIA/
EnxahzILUCsfkqLhCX5bfcgNZgbFVhlBJI0u9GeU5u2jCuSVtZG+5ZJJhJrUs/rm
Zk7Fejv0MZQqVWzoADj6NcyE6Dz+3rpqeXbo6vIYoMM5HNGiYFjr1rmfpzRxjWsn
fPv9xhfMvcxMm4tFdtFzlUm1TlijIbcs0jB49GM8kD7lj3rMy4G55JeODj4IJEdk
1fIUJeVO4+miyWhkCIHJ4yJ1wJDALl7GY3Q0W2LIzIOLWaZVW9Xgd7PL+N0kXeYK
KGrHvSAbXGFkwXZk+DrY1Xk5oTvAFxzT6pto/27dbs7DNMxYt23XJsvqD19s8hEE
O8GVRNk8TSrS2XXZXolNC0bcSOTLVau5koskQh/vqL26CiWRFLI9dUSECjYdqjx3
B5C5jHhw3S6bxLGOatFUguKIQB1LRoEWsEvT6Epa7FlYfo64p2kQlcJImaT37sL4
GzNUkeVT+vTHmZ1hPW3i9imEn70IgIH+SDIOuURWotsjBLFpiQffV/fsLadbVPNb
kuTM4hY11AvwQRVXqAzjadBlmjKojcMSDud1Ve1EzzCf8Gt+bWtnEFJtKRV55WkA
S5VgSguduc/RwDsS60AcbtfI9iOKBLeIG/LW1TeoH6KCOrz16xURcOHtJQyyHqzK
n2KmVXYPjoP2o4skn4F2bGZck6cXHDFTlZK+wEdl82gZCBGqtcCC2HFunKU9gF+M
t/ai93SI4YcdOBHUGcq992GDhtH6zu13LVtlH34uVG19LLwwway/5m4n10SwVCly
k2jxVD7krlkyk6aEXi57cjSKzZDL+zVicecR8DQkuuHZnySPS0FMKVatBJlutRl7
nKNH916QiTeb4nekVcTkR7ct69w8urNbQsHGhgT3yjcIhcd2oU5LMTFGI0QDhUoT
uuBgLSzm/RjEszwmhgl2A8UtTVXRqoJzav/ENbhf99HGErlQR1lGJnjOmxC4jcOj
1YMwzTpHXOduBk8h/fiX/yac1zoS7p1UCqUcfFJvGhFDy6KsTE7sMIzfMf3VDmmu
pwRkSU37Zhk45c9ZtckSM9Dmw67wKWBWRlTPNP5gLT+J9oTxNb61Z1ZlNhkTKvLh
sCeTzz3q78hGSu/D+V0Ux6Nr0pC5+C3igE2VKnp5cJF/P5LijqpxlvX/hyhFywLD
VSve7ZJrCXFhiP/zBOa62DVwVBzqXoluDh8MkOXVcmugcli/fkE9YlUsVNPRDvrZ
x8Ntd6lMs9VctiLQmyt+ffBS7fhvhhPCCdriFf/zCdC39Y4mDOCuRT8u4RGjL1dX
ogsRgJmcRmV2kZApJ28lpe4HkuaMnPwyAqSJBRiGVcdhaD/kMSr4Dm9vfeJWSnob
ZMH6rpMv0SLkQ+D9ORXE+dA4O/x5tc+SHa/7dCStrvGmVwRlnppWewfEEpfxxEIa
0Gq11s3JxoiRZ8Ea9HGXjoHG3NJUHl02dmqFfK1M5OPMQuZgfekn+J4YEoczUFJ9
tLCcMSQeHVheOs4koHzd4C1othC3NwroiPqL18BV7LldS8k+U2JFvQhmX1ktkDwX
8/PXQDsCBlvpzTuX29qVDHEN8EmC5V5VBbc8gXJNWpVuU1y/Vd5HguldL6SMX5Ig
KP9VvZwvxOW+riIKYiOvjcu1thNY7OS1slbuXN9ptJ+E1HvP+UKGk0oSE2No8+SI
CySrSZMFSm9hsIxKyCyOwpVLTG3X72VzEiHo9RHNU3Dqho3ar4NHPRzDocGBq9IR
CdRqhpu6sClOkjAoIJEGb7VjtA89k1M43o//wDqdGzeiin7ifKcjW+Y+P4pH2nKl
/AQHzRLxpiUT2H15J05s5j+26FHs4p1e65GaNoS+aLnzA3o1ptWOMcJgqK4bZVy8
ypAFF4ZmHPIsaucVZAwTWMZ7mbPMNlcsZlM0ZorvBJzn0uHtErSuBpCs27yemHpw
ZHf5jpicLCkeOULp1qKuwCnBWFPozP66T8+GurTdSIU7YqtIWprzGzqm6G803KN+
NkUmXSneRMPZfrJ3aaqG2hz+B2VqbiJaAd9GJKKR1idDMrqCpZgjNBH0PuL0C3Qb
fnKOzI5x05inexuZNsfBWRzLzPkLzVQSEGl7YngKovfU0x23iw/TYf9Yrsma9vis
YndZK6UBj+AWwYk9intcEZCS7Y+MpX43xXzbftgZWWGllqtCGBnUSqbIC4cuHtVI
zYAWr3XxL5jF2jly0YIAWC9pj1WvBRSXj8xzXravC+scyQZPCvRBWuFWFcZmo8Y0
ipFWnpJn/bHfd3L+CDz4f5NXJQ+Wx3vPH3OshoGr1cR9x5eKCcv36P8KjO15YDIX
YO3YOFf46px3tOooA5GP4mQmWA7lFg0anvPXpbg1FyIDvvyZ6o0aITw6y3UfV305
UF1Bs9ZJcUnN2n5UCWArEz+Er67kciUfFD/NphMPvVU85a6sqawhInxPWiBTsDDb
P5ekrzix8yJ4saXPmuywdl9UmGm7U12X1i46Db7n0wrfApazhI+ZVK8WTQxV3d7N
4YO9cQ3KIypHR0xVpNiVTjJXBSeVk3r4vDlEZhLYfXmuSOxtl/NiGnmGG3l/ro98
PHax8kmcmZKPZBEkq1BJze18IWHAGqggLEiPMsZUkWUx3fPGPGYoetQQpmJUYteJ
EThQuXzsUMWnZDHpW1UuGVhc15xW3Mp2ATdy+clf8v76MzlhUJyMQ2yJwLC120Vf
gXMMY0knJQ4vUr4KNC4Ma8Pk1t7aw3E9uBtl/GC9/J6qBPVX0PiWIlX2eSsgQjWI
P0TLe0DjmkoMg1jO1Cvb1dWloHyoquALAo/SjGdrZAoEJ9H16qYL/HXB7GwieTQy
PvuwcYIdMDsZabyE5atCHlGcqT9eyxibw6XQNOktB0fmbDMSVeZaZSPgi88Fxryu
CrAI66g67VaArVnRtAYFf45q3T/s35+ZcjhQ+VEumtVGnY8bTQ0YLiBNFLdtxMU8
R6qBQ2jzG8NYyfoD5u5VbojLZhnIOqOIZGEUkSdPgQZlO8jz83Kvbp//Lww04k/a
FA3ZRheScFL52F7ILy2PmzCbVfioi9QtoLrD3+xivAN9kCUeBzHlDlpJB0zEC1Yy
48zTXJ+mGpsoBtge9e5ZIzD+N+0WwkWhOZdlRCsS8KqqsKgOyOAE3NFbQWZxT4Ae
p2SVONgiNOJEWOt/kMQedX2Ik2rgGr5ea/REO+3wwZFtLri9cPSDXxeDSFXQldK9
3yCXRZnaRzFPkA4OPtdRI9uMwi62miVJGosggvzFLEtGfMZU9Xp50dW6WNVgaTi2
86BIyNJu12YzRttMacmVpqHuGZqoI2wCWFlDPLKTqtOIPZeO4BsD9caRsKi3/A2o
vf5jihXyxmACCQB59GNVN/VN7VBbLmvN2IylGlMy7pa3oVNH1h0fKDoy2cL+0Yb5
uxoftmYYkOOYPHkiwQiyKYqRal84OiYwpVUg2M4jKHwaXt/vpiLNGO6b1Toq0cIf
DJ3N/zwEftFUin9Se5W+XXAb5PF/zKISpFJM5KA8TgyixE8/i08C8r0UEr/YzoTa
ouVXMenbdMyskyW7Dnt5s9lmi8GfDPzh6FW2byfn7aCEsagXFtqC94KdOAOIKcRo
cfdGRHHuTQU3csUJ47dVJcqdsQYvFGXAOslWfO8hphCeib2Jg/cV0HO7OJvWCJ1j
eLKCVykqbtgSKX+ywIYPkAGVbvQCCi7qCqQB1DQfYdqtmUyUU2ARfHcJ15QIru95
GLlzquJ6JYZICAW4PFLFGrrvfHbhhDyM+Yhq42J0JVoPudSlQmPaxPr2UPUdULGe
IJ6PijLxDOKCp3jnExbE0yxmFxvraF9P+oxZRBt/3wXhLirai9tFC3wdcgGgLogR
uJjpV00E9K5X8Vd3Cu7jc4wfhDaUIhcuGAa6eVLc7CsWqJlYl3kpqQvBhVI9yrI3
I9125qjQjl2lPd9oghpYsRbUBJXYcjAUrZrQjAY1KmAramJRt/CQ7UVFxttkmrST
4x5gXeWXNnQzysDO6of9WzD4VXNQptWPkBV6VPxBjiSg0CUArp5DK9JV0Dkn0yAi
0z2h0zp9jmJayJnH7/WqNl0HjljA4IcKxsTqMBETeAcGp+tDjJBexL1NS0d9JTOH
qJrlx+CryPEJD8YHeo7JUKpVunxV5zFYrWwATbj+S9TVSE7XYdH/muUqJHxRYkeF
WUKBI4igjd8lmc34duH86XaIYXTm7mqqSTXnHSMAc8ICetz53oieSQHFvwbxSnNQ
6MXej4HG4iJWfec9GeO5i55nrjiaYaRJyKWZeL4Etk/xezCZsy0Xns1ZEfyCzmvJ
OhpzByddHWpqPhtVGbpkFlWXNdE2XcG/K+RzKZ+/dQMnbLN4Dyw8uV/XbwZw4dwr
qKfLsH98jrk9NN32SYFsoepbMVX0w15wT5NX64m5GuKfSQsKhRilo9ZBJH90MeOr
g/fcgWIqitAl1e2GIsLwmAhBytFtv6v7a1RNbkjv8HIZa13vl7e0RrIhGndfwoGP
eFumVj6EJWkzscgOqzJOgFReAsPfR0MHZkShbxJNXqEPjk8fZjv12Ogiod8i7/4x
YlPDgRlgi6aLFPFmoBebC2GzsuWOVuhGGgdnJWNxKj31BONQU7+vj52P2Xo8GRcm
uvsq5dGa+lNJqOZDFcTjnCyykAZVFMUPwlkEhgQQMdZSw9TnQhL/v5Dnkc1wueCs
AyqRIJLxcCicezUkA1/OuRER5+yR+hw5lKSaVNiYJNZOBHkzHZ3HB40vA4ovJ2k+
eYHq6pXZxBXcxkNaD5gfb+hzIoF/V5LQQFWolWcZggBGhP3FTftdcQWmw1CklQtw
VDqJ/CJ2YnwgsvhQlzadFUWxDHhPeOH5g0tbRdrezr2OXcnY0BOWgUpWiMZ+9oT8
J31J0YFCFZjW3VynWSEncJJreGKo8xc+H3OeqEE7gcawXO/kVsmLwWgnueFg6OmU
kizIiEdjVyZnD7Za4HokI3NgHdDtnwstZxVYOB1sYpzVanm41YYcCPod6JSRXtiP
f3qaoUJAru0nd1EZtQNUehiPpRRD0o5XcRTWmg0JW3q/W2cekr+nKPoLlxSsQyVH
Te3Kypx25w1RdInmerHuhMkNwFCUYR4f3WXMm76S0c12McjJozdX+1M7q5Raf5bV
umo8xxKKeClOKwPS9oU6nILRjjDcDKiix+IitBmoHYrKujihSmkaj0EHmTvSs3EF
9dCnzMk2fpOlH/fcz3rIlWtnT6GRi8rg0o0vQPQms/z6X9hGNJzHwDqBly/dfHNI
gQ/JC4TSfON9Pgjhi7uITpnPYa5sIt8Kp8F++/9SgCCklcj1+QQuuqCN1xBeaTOf
Y00mwhDlo7433WwAeJQ1RHFUkahYp45dhkXjPZNRT4jLHY2GeGAJq4ZBlCykvLxU
+annS/ASFGf882rPb6nBweq9XDJmm2dAO0vE12/KSXkmGFWl01+qO/tCrJ1wGimj
84UFXthYz3UcmRTv5oo95VX9OBEX2G2eotOlo6yCJ++LbHbVR2axMjbDKASVsYIj
S72/E7EobVdVTDOVPk1yiNkiRywY3A7gC5jN9V6ylz8KcIdCqBUSkrs+UZoIt+7l
E1PlCFBGPsUVjCMieFjk+aDMjJoDb3UlKFNXWm19tF8m7rY7XG2N8GnVAy0lgbve
Sjhe5r5uJ9WxQLEDKy0utE7KCfzXXKPRpvYECUnnjD9aLlV0k03QGmSSpOIi4XZu
euRiyeGFsNmNHA7E5COnNnsTNDvS3JpnAGSucKfXHqBJAJpGPXHXYFzf4lwA5bHL
WqlG3Wx11cS8uSvmyHeI2zWkHbXOqW04YKp82JzeHyPrBYYkZBff6+cfKJ4V3AfM
JDdkwkdk8ODzJkxB2JUEFQxuOBy7tS2cWfiO9HFf++HqyPy/k/K8FW8+fd1x4jQI
uUeHE8eec3k/kGEdUQv3XHpctm4ti93UUB4mPZu5iZ9JqVR3Ukhttx2DSJA4WTXq
Cn1fKDVqVdEZjo89MvvIlXjXuo859+T9dIjL1suSMMmLaH3QIwpEdp1ag2OmWdT+
DfjoJ9b7pbu5Z8SwTYXqjVbZgw6GgGSYuu8DtXvIolyPLssNDvWUCuYnnlAulm7M
qHmUkamufQFtyYu3d/eiJX6KxqRHr2e3vQOIfFN0xXlLqewuPImkqBKyVCPDLwbK
bEW0IXSXmRaPD1W22MQKy4bv6l1NIa7AM6eSTFgaAjh3udWcoasUAgaDcT5Px70Q
vI6lDHezXqUYqtbJLTs6HW6GoLH6d1zUZ9/g+1mwHFA5bKT1TYFWJ8WO7jfWbXsD
lG2tuyTyAsyLdTDrcMH4hxJxSApDbktCNyoR0RHRbLl6HQ0r0pjLb8ZRsGqqXCLx
YibwT5cLxXvaELK3XpO6EqkARBzk13IYbgmibQlfLIxs++a/ga5cBGFHvlrrdP0O
YGozJALIU+2jfl92FGwCl54YADshiUyH3hgmFaKkhx2iDALmKqxtqicDePdJ1i/t
jNmoWm3MkRwfFVnij0FVxaZ2X10vXNag1CqjO6Oh+OWHOpvTsQgcEebBszBmbPq5
j2cQVLe+arK+PYGY7wTZxpMHR4Km++GCIph+Rgpffki9F+AGBdCTeeGO8Db4Jj6J
1EdGFEDOKMskv5+LEzMM5KneHGfRRsDh7YK6yvbJnrx0cfo3syJArKz0XRHmmgan
EcK5sYES5Q/jmJnUoX2STjXtNspsj6UkJFFo6tzEZOKFWc50qptpCmqvAMUWK6xx
RTOXpu5qlSYjDKKEPiWenXx8ig0zml35QMcxFn9sJ4RlUTDT1EwyeZwIRicdKWL9
J6MeZdylUzViEZDEgnr+rY/eJcyCsA4ZK3C/5OwE+RY0wsXxPoVMWKLSM2BZVqR4
kZsQM8RfUd5vjEi3Kpan4L+LcOiJgcrcWFhp2RZyxKj6wcdSiMnvi9fXz+3reX/g
TuXlaEw2ZJzLQZGczJElb0AOMZGK7SfGpwVxtIq61lPFyy0eJWJ95RwoO4maUfNX
JHcRmM3iQOAizP7DFxzboGO78KbFnShH986iPxXMtEewMd839PJv0RQT8EQ0NoPL
ES1o9hFkwDjixioIAVQ9X5mbFn5THmW9/8PvRBXhKQxHpvW5Hqu7Ah2bt4OkRGna
U97uGijwjiKyNJ5O+SEyCMnOSUHzyCTG/3fgVeDolIODmNVOdMreWXrd6SO2twOJ
gKbjU5IP3MTFrDzPLAqoVIrkkGR5Kj36hL9MBvN/xJ6i7Zgr0D9jEKG+pnR7DyCl
RmqPdS3XpBwffW6KGpxphguXPG/VFx1uGZ88jys3MvcVo3tiTWu9lRzFwokZr21T
F9sKponRD9fx7RPWy9Jwth+VjwrxNekSkdbY4D/BcQud6kBdTrWpBu4RuidPILzI
lx6JzmiqVtFrxzJNVP898BNbiNRO2XHYSgHaS4HyOJZyHYME4snPTdqiDzlWtu8i
8RR6PJfRyD5fOBPllbQlr47iSUlVlqybzfhnDeL1KCqyjRMgl86zR5k6m7SUWfCD
gUCSxB1Ol2lMU0NIBh6Mkm40frIxIVqb2AAyE1IpwyLja8Q3euc9TzXvj4Ke11wR
x8LHVxIkxGySEtIvI4BfJrlUuuF8UnH3/3uLw5+470BiF5AumVjTouOH24xnf4BA
buCUldBK6KcWvDay1G0Iem7d24zoRlJ05TcA9P3VxqlekliAjPxfC2ooex4jYevs
WPvWbdWbLftCgQiuLUFJujhxyYtmOX7Pru/jd1EVAV5bWnG+bwzT5w7SZ6fSn6Yl
pYqT/hhHwpT9iX1g7V76jlxpXNubBxEKRlLp7RLF3oAwMH5y04o/mLY5mfOK8Ek5
T3zp8oLobpDoPWdbwyiopNXdQMWO2TdX0YSV9+qF6PupARSg4ODwbiWnEcIv64A9
u+pVNKecauRJW3gvrmaIxaTJTw7awWpjgXsuphyqxN9iwkzNKVornmLqY9Ic1i/M
aVo4NjoA4pmK4yMPIdr+KsU91K9I1tosckctfJh+QgzBlCUv/Or1ThYUJb+pxnmr
VcC1CYMkpRBB2arBUA/KO9j33200XLDzgLT04NtCQsB72eI7LylSucWI+NPktrRC
xYcquBZP256XvRP+auT8a+ftMClgDydqj/BM7n3SKucJ1DbtyPqIgrnlMS/7kmuS
446o5jaCBYGxD7eZsArTx8LYbfvesStG+hwgaVFnItjdO0GF9yKlwdBQiLxmZjD/
2EfzQNGx4v3QlQviANuI1GCECvl0THlX1XW82eCekW54MX/qvq/lieE+WEt1zuvX
T7Zzg9rV4mpIya2MhgYdfzTqr2DEHOl0/z5ZZBnR+tGvFMrsa9hQOd+61ju9xbka
chXTQYJYMTnYCijjo3ignq0rn1+W4TXtE6r5QRnJhTaaak862twUGw8ICJ3L1T0u
wZ12no88j1ZeOaJyjHeXCkJlIrMe4w49Y8Ed4OXkmf3Go6LhhzyNIkmdaw5R/d/I
6XgarFG/8vHwDcoO44AHPvGj6DlwgRdLG+eVzKyIqNf9xuIGE4W6hD5GuOp+toFR
Nv3N2mJEze+ewGoc91BUnIws5d7xKGhZ857m7mghaU2aciV0YzGJXbTM90EjFKxE
qogaEErYfhPmfHJ1MlZTxqvbBQPv6YLt94In9jlKqQHQRtt+ttblKPziBLr0yUJ3
2kOat89yiB6vGGutJHl8CcikqgFv/ftnrsjTeSh0v7IU+FxcVbLLiWDnHEvNzywZ
fIj4XQwZYqOx5VZQup+4vG2F6d50gFJbpcBFcY7SNL5NW09R9o3o8iGlg47mrJwY
7/fmGyt5MdHDrjag611UEf84oBFSXTlXiXgIabBJWOvf5YDhzR96t7BKa9QiYBsu
R+1LyP/q3KVfGI2PgGFyIS6wbAWNZYeVmoqaU5Z0L7ccDqRW1pw4ZicBanvpzyoJ
85u/ox59l5315VHdoO9L0MBUuXVGshjYD2e8S2QTr9kYB9OWqSoPEudHgWtZ3c1f
JEM4pW2zMFbfz7KqKph5smrS2r43yzo7UI2Mi3HnbmxFkOnTXrzu5iIztNxrlADc
G23mMFCANcSob4g0puqoN0gOCnH/LF4Mnf/yZGt1pfc+JRuN8fZ6m7Lz0DKbx9zr
jICgs74u/Vl282WerR5x+4RDZveS6K9KGHMQhX9RIfr508NXaqLtgO05fcpPFObP
UX4OXBd6q3b1M1e6VQorJUvpvW/uc3YUdWaY2CQt5Mo/qHT6pcMGJ0qEWWL2PhE3
A3D6LRVCkgwiqxmEMT+OGjScrRR8TgOrrCs735ptJPZM67jOpRkrtpc/RlNnkgel
MG1kwsO3pFrHsVFApRnv7pSrPZV96Q6NFEUJ9M+h6CfaPm/1CPcGXhuzByxH9h/I
0L/PICuSedNBM8aogdBRFwmGKHeCT6DvhOwdX03IT/RwzhZnfG0Ap6PLaBb8ow2E
aZnb1LIfxEYf/a/28QUgpzcnS2AYL6fye/5lCbHPCkHR3BdACTImFOxDwhvdZVOQ
MC+52i8LNG49AQoQmQD4Cip7c2ETYGFGMHhNe69LpxlpjR6Q5L+NxWMY9GfZ8g3e
g1JGpb5ezSMIW/h8qeBMPmQ5C7/ZympUMmsj2nv1CyV1FzwRhbwzvyTpbuYsll0M
P8o/W0YHW2yuwac3+WrIFZKydS/ScyrpluIGzZr2orWNQSplBHQsBGtChWz8IzlD
AgovnLxPewgyer6EHBiyaikNO02Ed1TOpVJ6uNHdlK3PF3sUkVnMPHtPE5W9aG+h
7tqRYmWRXdUl7JzTcw+NrwWwitW20gluGmS2Eygx3miYZdEadOh8XlK+ak2czPCf
cF2j7lLg+NToW/FkkyHZSBtfy1G1BZUEFIDspBES3OEq0hHYxX/2ZZlrC4hNRBoL
W2pZLZKcm72IPEIUVPePZ8yy4QBXDP/4Aosk/a4NtYoMYDVjKwNERaG8K8r9A7RD
CztvFr+fpU4zM2SmvpYON12GKmV4alTMI3f9mTuLNa0DVCrW86yAM9XauZ6Ghp0n
GjYp6n4lpvVbSCRZY4/lLGmR06jCSjMvFrH2KZ4KSneeFWI3VP+BeBsmirrfNAjS
WVgBF7HhiOyNFTaUf1huEf3psC/ylCFewANbWTjHvuMBCC4tFGeLUaKaTuxn7dkw
yKvvS1aa3+iqM6oNMaHpi3g2pEJNsv5ma6NWe9bfLIhKfD4Xf+rzvMYQpDBEvpOz
Ef7NgmK4nZ0yChXn3cF2vPVSy3BMxp+t6jm8e+aOzDhc0MNN/cr9u8UneOdHxkSD
N9UN6k+C8XWFZalebys0FyRKi+FkVTAwTNON+NLe2T7QuFlYgyzJKuJlotzGRq1j
3SK7eCc/aIunv1iujS5LP0NA3yMqf+VsukBrBt1eQTpVQwYRwAcXk4vXq/eOnCbl
mVTVItZ/GFgSiMdi1AiMdxgCjAH2yrSJKHjnHI5hFMYUiFsivRLERP9oabuEZfRw
lFWhyj2/x8Y3urkus3nyYYQR/K+ogK1Y3wIQr21MhMGW4SjSDXj7LMXJ/YbTr/bQ
GbBuITADS/a0fQrFSpqxBt000Dk7qOCv6vyYfQpwTXJWMsmmCm55oQSecyt0/uxu
x6OHzezc7c69WKG/eyY0YYj3jCzKjG7SGyav3asQ/lJVTMUbyuqz2W5oxbBGbr8g
hYVaOVkgRKiyLJfpvAlgKW+2r2HLmSbQ46fpWzSMokUf5Wg1/VfIfQGLbHz6Ajsh
ZL9yFBJ0RhP1EqPP0bqz5A9Tg/0iUQ57RgQqcggMs3WnrS1U2Fa4xx0xV3t/L2BP
ZQSRmhchp/iB6g4Wa8de54moK846N8ZUQK2T4TXN2UQOoJvSMZjkq5XrhQT7lVeJ
tBSFgGj+sUHQjqWJbNBKQ0p05du1RVumnSsr6dssXCilSkziUt1A3uq3e0pn0Uf8
w3E4NU16zC9jw7dX0DSRBfq1/Lj7RZZzKAkzldUdSpwK66/vSvLzSrswdA4Ebq6l
Vs6yppNFU5bOGJwx1CXxSiTrMILTpL98MR1DyCjZXEsPSULdhaAbGIpe5U+rp2pR
AmOtkLGzuhbbBU6Rx7pzKWFBL2hackwu0epq2NTpqMuBMSsj2AIMhq4mNuqpZcDW
g5O6Mhl4BXL5T1AQE5q+S+OXjE9aQB356bLlCrxZI9HUXadPMLxXOzTmuAzFjBeX
nuddJL007RyKJr7Qa+au6xEo4s7vhL8gz9hVKJkLYsoBEUiSQH2hLS8T5/rEAUDV
eld7+RsO74W04awze4araAqKUbZJLnlNInL4gSXterTq7wRcqdu2FYhYQ6u0QxBG
000iK91beXE/4jc5RMcbNsPLvSmUHMVLVFgb5K1qrUt2TFZsoL2GucRJmKgAYXiS
0TvxnBSVZ9hdAqPznQs1ftMDwIo4Ax9RGBtMk3LXhABVgir7c8Ozqc5p8bxVbC0n
S7O6TtE7aflWfCMLAypIiA8DnxI44v5aIS+at7Z3RnSGlJgquoh5OulwsCeNnQMD
Soo9UkU9b3BwRujK3Z12n47qzcBZuA0aDUzLEjVGnp8EidjuTGBQzx/dvbb3Nc3D
GoVtBZxE7Qx9aNMcpRa1U1yDeyPRRdAx7tUfWbmBWDOWvLTbK+UxawqZ4K2MnTtV
0TlN8X2w97FR9HCJKFw8vKrc23wKAyaJ1gaDAKgjcL9LwxaBe+ij/qmzhOstJf3y
Wp1SPIy3IXiwNvZKwUNZX6uAz6NEalxWoc3aOV5AGf+DWBsZHdXyKLOTv0kJAspH
zPXAKFAleMs9uN4B8qHKgZhf7icGB/Z/FBz3ag5MF1rMDLsRaikrdKt8Tb3g8mwh
3wLZkZOJeRTzOjkGvDjthmxQxMAFHGQcXepvNk4urZUWvSqYszTfQacQNQBKQW2A
1fURfmj99OIYkYXl92BZPR579wn7tC/OxaeCre6LSIGmFV92WEPcFvNjqXu5sYfh
rEeYr8ODV+H/tPQP76+Q4csa9kRBlj5LyBWFcGWFUyt1w0XT5wmQV5ocGquuFoC7
GS6h8C9NCVU8qW6p/0x/Y1RXnpr4ecL8wR3ZDchDz5PL9pnOCivBDf+TMWJ97fXy
jHDDSw9wnEQR75J2CVeZP9QLxSAGkIqQa/YzLVoqf31oGjZl0xkoF4Ef1iFfbybH
ePkMwb4kXBUvsfhoIs6OBQznL/zvCdhNk9kpvi0eVLTJ8w4KOigEIPq/k7rgunhG
IC7kB5wEqiqLgfdkou7wSVYch7YNz2z9ddjotk42Ms1Ra54vSB7HEi2hU9baHmYT
teRVucfc4lVN7oEykSbftat2TQEVXc4pi+gzpbhXV4T+BZLPqicruSt2xI6AbLEE
j8LUKSPCdvlygeLVeF9o/pyCgeYjkXhvBVm2h78L32ZodC+v3qHXmI0W0eOEaa7U
8m3xDbctrCUKiCOAsFgvKMVbrKYDLuE9yIWPZLohZvYf4xRv/W2gnjr5zf4y2r2x
JAFG/SidrM92zzaFFTq/VadYl228wJrZJjDy6/HuTYsuem61G66t2eEM/GfarvhL
6rGq2FFgOELA5I3Pq5NKhV7EOZS+THppy8MOCi/AqPX74h0+zVtZnWZY38p1HCUD
KwCIVRQkMI7R53BsPRkXa4Do6O0HKkZ1QhA4p8FFnIfWjl/x2SLI2FVctSJL/nPB
x9h0CwpqaozyzMvbEf1B++Pt+tOoywcyTeNf5FgQ70dgZgEzrCarNGmgPcZBeoo0
IpGc3bjeOLZ+gJu1HIPCbFppC0/NUWyZkZlx7ulAurZ0t5lIW+UcwaUZSUzBbQYs
wNg/a62byHS0mZiLDNygfPbxCtXFSD0yBiFqUj5LnZerqubY3GeqQeQ6HPYgktnj
XKkL8lCmgfO885wi5rgiY7zylPZbomBtGoYF4fCela59+w0Eg3jdIVaWaHStNSDG
JohhucGvcQ+ArRC0PMkKjPGAihVyiBOVsm3ByXYi0S0F7oOZarD8fRlQclR/KldC
gRW5LlEN6FDIW9/Jgb4aAAmDju4nuHz+H9lDfnLrp79WN1SaEkQU5uLbq/uUNmCd
ouhCbJNPrsXF3ajLMcs6kGJdeF8uztOHUU7QxAXZvbTom+UIaBtdl2g5qhXA1m3J
6e4hEXIAgUSldhv9eDmmQ7fFRNWt5Mo+8Eni6wAS0qcE0twIqGlMCo/fUnoiGd9u
ZUAmelZuUhFHSCjpO8kmcyY1tz+XE2TzzdodR3KG6njkO3Bu0fdZH8oFP34QYIek
acqIdxZs0RlTw4TTRve+559xqL4Cg0N/H740iQh7enDz4gSGXVK+3lSjnFstDDWo
1SWnvwKUAFeTUqxMDCM+oiFakXx0zyV6fD2bTEQziL3J3kUdOsszT6Q5H9VqfJkE
xJl8LHuitk4mEPQtm1ZGU2g5HmYIia9WqOiMAM9sDaU3avRDsmuyA7p0d1KuaFHO
Ymk2cJMFdsM/m4gniH8fx+ZaLE7m15jCPLIcFOiGa9FMr9I02va4lGrJKE7JKQMP
Ast2TTmZBYgQOdM8QoAbwtPzeb34zANubO4aZ2i8t6dnX8CQdFPRTs5Vxpbyyyk0
jaKAXyq8zP3hD3h/jPxNfc/6w5C+FSHEK2zl4x06n+lPGfQpf2d63H1n/V8TPrbF
2iQACMs8i8ekjt8jdG4zMTnA0vmR3Upf7degM5Z0WR5cv2gfQxlcQz8b8G+U7TGL
2ASUBF3/C6So/7LG10osjYOLGMFpnbpwf1XZNlShHtMH52ZTphwRjREs1BNJ8jyN
hS99o7gL1VJLDWZwhWEb4Rfxdg23gJwqyiNa001ESTf5mLvBsHogxedCu5iyZbY1
wJn59rA520clwiySRQ5+FDA6sossl0SLYxYVV4yHdaa3Jh54BjpUPLc4RdZHnldW
138BrNLCMP1GR07rBsquBMTrQBTnCuOuksX8E1t2JxBRCvqsUfJLgSPA7aV73TIl
YELz4+wyvTf4JrA5PbWBiY9UMfHJLUoICWJ9eD+iKDTeCH5FC0QyGfFvwGwfGJaY
Nr4iE+OhXV3TUkK27ZorLVa8guCFQ/+SI0TIqVfwDMVvnisE/xidzDdP42Y2o7uc
RtY+TTOoIq2YFS9bAVveJ1oj8Tvqc2X4wtpETghAhy1yQs8L5/YvbNFLs2EKX6qB
h8PDaIU+RhqVDJa/AthsUWBqr4HlgPXuajJLVl4/fTKBrG4SsSUg+4xxIfhvS3VA
jCWL5BCSbKoew5vo6YB+CDG6OwTmojClkkx6J7SazAA0SWC/JqVEoXp8onZ5gW6K
YMNE8NKDZ/Jai985fWoAMImhzFhK0BKmO2TtifR2qjNLhXbAzSImATyT0hlAxboP
vom7O7BCMd4UouylUgwrTQ/4sXYuK/I19WlsVYcBTH8VlwcE4RZ5XQHbhJ7Y24L4
bf4K0v2Ge5O6rJN3F5tG/z/tXO6GlI49isAdVlqfzyhFMjZp+AFtIniarm/AAcJ8
YafZEI0FzV4EdR89oHBJmPPnJNKeLcTEjG//HO8bSgc4ouQqGAqf9MhR1LEe5kHs
AMJJLHFhF3Ahns52VajLdTE7UNG5lEfa2m2zHpjkC8NwNnUegSqxkQOBvrMdT26j
GAdFVfslsV3vz+ol7qA+rlXhQf1Yf8J3skyHOF5WkrbASJU+S0eW9VWpSaw5t5ZV
W+ypGJFzqz22AeSYgwCqYM9XGeK3gwiOd6z1g7qyPUYiSOFsBz4/Jeek0AhKIPbo
30wKPz8K6av76MVPuVESVkHndyZLKspSSyM5H5n/0X8wIi0XtZccignTxmmpR4ql
9sg7Ly5FLfGpSBVN1N3C8aciQqP29mitVAzPpJ/aLcUCydYYf2rReb5QTsKdZk72
bDRDFW4ryw9Yg+nXiFUulIR9fJD1rSk0u+5HghnxfR9jYlu+nBpBuHXEv21b5p8L
Ibl+NGKrIelEEXIVOa059xam3dqY3zF+WzCd9NAVTVa+VXThHfqk8eLJN27dvALr
u3SudeToDXVEpKgnWU/CsS0YtCZQOGjKJKf9L8spjrQdWpDDbQMIRFSsHUL8Q/3j
viqtygS2ufSIfjQIshZL6N8HgQeexuCRvH9PEp8S5z0pcREGjxwq2zJ5GokpJxbv
Qmbd1dgEVh6BC8VQQmqEc4pk8w4ExbistvF9Rlaw5RIRDr8CaraCeNa9JJANknmP
QcQMlsn2K03gX4R4IaJHkJOMAJIsQ3S5Whg9TvLBSHsmZ6g85Y265/ecuKQ3yrvb
6fJET3d+Mwhmm3C61YYiEjqEEnxaTmTY2+6QhnlIsO0wI59K2JKfqytWnhh1taoj
0mijn1DGn3stpeotmhGHW0nAVODECrTMpk0N5J5l6k6Nud8SKcCOrdOHetLp0Fpe
Dit7+k/ROSh0QcsqoYMlC1AK+grP9bAy7r2miaMbumbohmA8f9cn9wbkADJQoSDV
KVim1PGDxK1XGdva8mBCWyo69QZXpHU4WgWwWL1++nJ5KYloxhN6KUZTXCQ4nYsS
36/NhaZV7LFiPwjBZpTlbcIAFsPMSSAyn2FawPfLmlnAcBkMM8thZrI1aw/Scx8C
P+zwDSs0Pzm4036NpjR9X+Kpyt5mJTMd+JwZFj4G2AZG2F1KwXeSW0ZpqAGmDgDw
HFYCxfLiBoOp1Q8Q9HO1QoaNH8iEp1QHiWGbVzCw7PWH7XsnU6V9mOqmr2Ddmpbt
beiZb9GJn21NIRB3kJF8NQeRJz5A3M27rnhQUv2yEoBZXfJiaEZQ+bwFyts8gAeW
K+47uUfAicoRC+bPoxuMlwCT6EgqUHcUTJzhoLVp9uU6qVyGZFrXe6Jsuf/P8ROF
9bwrMbO4WBxheg7F7QlKWcYctRz+8+Iph+JCe3ig/j7hLKP1//NkUG3ZNJUGZArK
ohD4rClrp2OKB1kBowAz62VUwylTdghLUM+pacrqUxQl7YBoaTlIRGv0ReXCfsE6
yQlzyjw4jpw/8RtnHVwtRgfZCbGIRf+dlWsG4Wk7ZK/DRaGgz+mB9uPdPn2TFLVc
r1aWlTZsDBzRWOhsQo5fDheU9gOy7oqmNwLYYbjiVGughb6H7JX0J3CrPiv3182z
KCbPLrcSAdtXMoi+qEyTdPNZTmYM9R+pUJYQgum43wQ8v5z6u80bkq2Ci+SxYzHI
sgjb8KKBqdMt8kwAgyentFrDwnxgF1QRVnqfWWmFyXK48uRPOTBxKGtP7Mns4y3J
uXux5CQQA+SUk/NzFmh2hjkk4xHMUPnrvlArS1+QFtx/OjUrYQIGAe2+SMbZcvVI
zVU8GCzKvpaGKkLwEcuScmX7qKyKkXMqhdU+2cUdiYsGVLyqlgfwaPV04xj7iGQr
gAFtzBc81TvIO9xStVxA0jHE28MZmzQWFI+Tj5jHm4U6JYmG76INOci6eQFiYpDq
+RbAD1g3NB1IivefJpG5qmVufRL2DADnCitWfsH1fptBxqGORViHWISOIV72K0JX
x7n6sA6s2jOvW9D7Ui+VcyXV3xHTp4Qai1tUTSn3iXwaONCkSISYozTUCC9EZjYs
/gUz8n9LKnFiwsA7BBtrKMG6ILFWRnKOVoOTff5oyW3N5D40HZk7c4c+LhFjamSq
IVkzXEYnu3qwgbTDO6p5quriR1uNJ6rcsMNX8sWKrDEhHZqn0hZdLb18jJVfBkDs
PG34bAeBS3bfYuWz9BiR6fzozttA7SMcFmcmAIZSeNJ1RBXHXCXYl6cbC/yydoKl
/21peIwYNLJgsDPzdnr9SeS6WNBmQ3ehyDewVfEXU6uPKi5CartqtXOh9uJO1ssn
W0Onuy/qk5ZRNA2Td8K64myOYGw07kY8ZNi3mVSjzY77xM/fJAkeRuxOm+KJGrAJ
+Yg/UbPImVBLC+ThnKl/1X6y1VpjzoPHbqga6//He+Totjr9Dc9NZjg5uoMzkMGK
sXCOYa9VzTRphqItvV+zOvP/8/2Cg2LCNXwKo6XlydpzcYTWxbZ1v8FocFDwUSlj
mG5WPqWxjWXfGA+QRkt9qQXKEtLzf5YZidzIV2+nSKhI/yK/8/ZBj5tSB4w6Ap6e
sdpvWPWNtV+rBuZAB5t9YHlG3CzVi2vgPDggkOI4PICW4rtV0TfpXvMfKH6grpR9
wevnkgp1REkJtoXEww9/k51NZeD8Q97lhynV9mOE81bWSFDUJyFxvwTjuKzsmXWV
yqMn4nYn8CfcZEiY6ybPd1ifIs1Rk7ejaZPTJQYVZaeSJYCxeiOzrFlV9fHrfKbU
kNqLfkWUNQlotSBhdfPbNNDmRzLzj7ae6VqmcfCamsUjJLcmxiQ2oZCg/5yeRdIO
j8yEyhjy7IlmUXorE34d7Q0DvkrULv5zA3oQ2RnAND6OduFNvKnLnWxrjdT0ytO2
LakMtZ9f71mH4uHyxgHOFYPcQA+onzevaG7yQrS+vTd7Pkcbi+d3vAVyX3B6Umrd
6JM1lUtv8GITGRM4tF8S3Go20juVL3KagdViAD0C9ny20KDWAVzTjT1CIW9a0Ats
ytJgO8ZOOLT0zpXab5ZTmHzUBM7tENvcDXNST0N8bILWGVFLi1uasEl13r6iD69L
Nj4BaIvvDsinFSOGf7NyggnxRdKzDnRINj6ZuizVmOjQnUAwshhYu5knaSLLGf+5
0nVqLTcAF5ERYPNlmPAWtGwnN5rknqEVAiqloNPfdEYqtzt525Ej0AIidoKBY+NE
mqrS7y2brJlxMHfLSf1C2U5P4znyJX8Z6I/x897x5TJePK39/tCDdbELFVddhui+
B8VR0P9odhEvND0tJPzhGUX9HkS9AEQNat6MXjdXl/UzbJ5puuPe90Wcu4P3pGRn
gpTmGmv/dspVqWhIh3hPCJ7V9Q+jgaSwQmV+mJsRhV6nGkuKkq2wPjXcDNp537OF
7JanHYQmiRJ+bfRHlfUtyaos073KduLr3tl8dN+M+BPYi1bhqamY+T0Zd+Kv6dQ9
L9Smd6l+dGy7Tpz+7/M97oEkYsNAYujPKfFh0aP9+Rw1IoSzTHvep2LjXdeyntl3
Vey+pqkNsDzd84oFmtIGHGJc0HrXWVDMoWuRxUJLNcectAeedgiuvHKw7/mhkITU
QtYc2/jeTiW2gLIHpyKGwMabf867QS1tsZvHH020j/68VzCFWWm8YHqPbOBcLo/W
9nBdTmpQmY7cLgXQ9wzVaiAVgKj8j4OHjre3F7rBSMEBnOKuHCxzvE7YC1AwFc5r
jhOi9/vcz+U23shId7vpQLrBAkCrLUa7Y0Jh4weR9bQ2VT+USpLox/h6uuREM8kf
l6NhBAMfAeNKBqwAzMWakcr/GxkJZMitcgfOo5wzDM5UydwJYTasMP42/l6dWvoy
BZioey+f0iDGupzGMT3i/aEsbJzS4ksh1V235kw0fIuVc9WwhPYu/YovFFimTffo
yYjfAIe7Br8IP5FR0ffHO5yud/WAnBxNWpTKVbkpa07D3GWSMKTRQvYCrMbdFEGW
ZXclf47nKXmaf0hMtZsxVNDTW5yJnYAMoQVY30JUqyBRIQvRF/LF9g6KNhzB2anD
aMMgaMYjkrtQn+ga9WyWydqs2FP9XFH6xrEm+A1Snyq9mKPfaMepMRmU2x014ifN
YeYFYRsC//Tonb5pOqfYifFqQ1KgFa7lb9bw2bb0fTe/WTt43lcnXwX3IpUwayza
jVUMCy4jvgY9wOm7NYxs3oyVy3pbp8Wi78uc5wcEimoPi8q1WSV/jqHI94NnrKzw
7DTzPBLRL31Zv/8wPnU+BCbowNHOfJMG+1MJN5ytz/NoG7e9Oolajj0UJv/SasLk
gF90WS8of9pPVHRWmJv8RokZqdG1KX0SAyxPe3TKNW7gdKeTpV6u0ABpJC8loAuK
HHbT4u94jI2OnnPXREvqgJo+P/CUgsrvrYqBp6SwOB4O0VF1NbQKgucQYyEmoHgV
+Ru1Y8j547KWvoWpeCliQRnUTRs8aaVeUOUQs6jqbe3EB0vbj1mnFQtjDFWvPqr0
kMlP0nbc8f9zDdNjRvjG75xg15VC2m+UjMCV6FW15a2uQndCindleowPPPL7jWN5
fdXRsfzeeWkxFU//UaD2Bd0shIYSy6/bX5NfOHCWOBA73P3SAAXoJyFm//AXnJfY
8c8VV6PhMIwfqSKOElprBte4JpAlI13AYJvnaZzuG3mcr4JRv8vt408Uj1oed+rr
p0iuPErFimbSeZM33UqrZHko7LvMy60fTVnUzhTr3BhBu54GexO4GosL7XdmaiyQ
XzNlJoBaSCyWAduPUfHu/XJX/JrHOAg1kBz1exrDfYmiOyXvqNmsCSQGlpNHeLsN
79VDA2qd9tyMSSXyFlH/JwNEfQ/WK8/RGaqf7j7lxyPTCJ9VmLbsvX1qP2ZVDFMp
+W8fXjERsBUuEt8xe8Iqxj+1y28pgkStEl5WasyulH3qZTJxsiniho7h4o50WXFF
a+K/XOqwm/nk6NwitBD4qanITmJf4iH7tz+Ui5u4or1czWz/Bk4gQRgUdoCJJ4iC
CBszIGGj39ansu9Km3OC62ifWWh3ih9PD+QSnJ7ek+xPolpcupE/fhpMgvtBEz5r
2ZD7n3LQogj/Nd6wvJ8CFM2EzEIuMLz+Rt6Ky44kWJlJx/BwQz8+k+MmRLaOwKyR
d1UcvmlsIp7iu+gQZwrV9lFlzl+Uj29CiyMAkZRhuykJ//L/fKaeY7RuSfUPeNb4
g/uenpBzORjRWvgrFdQMkpO0bwH2OQGEvTOzs6wpIRRr4mVlTn/fX+FT7sTnXWUC
vtOJ6S5Vv+Yh5oflMDMzLK0W8SNDvrCElBepLRv8/RQOj+jnLEWqcqEC2KcG0Lai
cEVl/mOzvVhd18DmrWfsZnpT10i3LIUOHRZGpXbsmbnFMUVCJm8GJz74X02BFsZ2
iCtFu5QwaYLpD9SqfgBaN1HB8OVQaC9AGGex5x7m0KV+2I0Xg0K0VgGuu8LfV2Cu
mEjorBcAVaxOSTMl5vyMM+IMPE22yZdJtMw10R+4OLL1fJgiPLhZ3dTtOgCXhSj3
16rFkkqeh44quy4e+UiiZ3X1jaAfMljuFsCMeaTFtjlyQ2fP9wfCm0Q0Ib2meLd6
XQ5OF8QmlaAP38rbBQrCf/P4P6yMw7FUuwTASkJh9XG2FWc9p/xuTT3YDFJz8tgo
kFanfcISBswUIyXdBO5wMx9bWlv2AV9POVGGIu3SUb3/7k+LW3T65uC8hG0zH3Jg
6YVTkeu7BoSLtfJctrcjCBVdCyV6M+rwm15Ah+ZiyGwWb2V5DU76qjiFgfI9uSjN
xXpfE4UdIw9+24uZ94ynZCSE8F0LLu2gD5HCtKjrAvM9QNPaxmHSS9mWzJ3UrLQO
cl1h5aeM5d44TPbvuWuDQghmcxa0ptJbK51V2Yc7YYsah6hxD/HYFdFEIe8Ya3VT
lsqv/MCbE3UEAC01fYkQHAvHDvJqGtuYFscPQgOx5eaUMa0XiohuT5zKL1+fHe+p
9CCp9VdFQeeVWhxQqajjcV0FB/4YOIWFjkjv9hbAajNZCzqmi3ckr9P5OQsTiGdM
ioORjPyThckZJf/SHlHKcEXsHuCCUL/qOTtElOfb/axa97bFwCI/K7Ukb34/HOLs
VOfII7kL9DCmoPyR/OrTUJA3BlH0kTx7GYxvDkRjyPmMr1im6un6KPdzM4oVFtsQ
wGhdulTFBPRAqePHp4ZVEsjGNCwRvi3XVbCeDeGDesopE421usvkn7DVPMWce7hE
ym3nNV+S4qFZ4OSJAXW/PbU+LVkREoPC8IT4MxCmJxOywb+KuYW6cpEstj0XN1Gr
pepUfBUUGlkeWVBRINqx4VVPK/E1zQFHLPVlEQM/BHj9AU0wf7PYnZM3qKYyO7jO
k78Hzk/kVRZtf82dblRbV1i52G7G9EtjAT4Cd3+mW88XQ3xXvfS0i7dEAqUPjbyO
oA+Dmy8fPAYmrEa9cn3/TPpYq1clGAoSeleEiNq/DDa3qNJV6MHjY7jwynSIkx7h
UjUxaNxsqk+aRkgk1hpM0C1piFqR1Mpf4JQltd2EiVrq3x9MH69Bp9+rusW9sigw
SvI5XGXdkhCNZkKDGO0KJBTGg34OUCeWgifU3a1ZXu5sVGtZYwvO86RxyTzH8ew6
ISBwjvinU9WI5e00JkJNY7xrLQ0addTqz3rrOxsPnubOXJz5AhT+jlVk2h0FiVRF
T2nE5zPQONxCVO6PQrzwy5Lrj5zFIiGcwFtcThcuX09SihS54GxuUQgrY4KpXu1/
THbdVuGNsgTdXlJblkeWX46teHgwEMPJMVhIeN+nzVALw1TdH4LOAmpaEh3OgJ1X
TDch4LGGcUqq5uplqfd48OdbcI3ZkywI99+ulEPg/4pQC73LvoRro3NbWJc3CCkV
cxNNrSgKhOHP4pS5agLXbztC3dUgFDf7NgjZHprJ04wziq40l60EtVPszvbbe0Sv
+Cr2UtAMat2mKitRzgWV5uRLBq10W/lY/myVXuHMpRIc2AZgx6U1AO/8N5/60O2u
16FyVQIDSjwWSm6TDxveHKgHIbZel6aH09HOQH+TYE8E7jwULoJu9mye8iKvcCZE
EiLXFSJnA9lsrr/nuBZzO84LQOykmUbqRnL+6qFPTgo1n2bixV7CmhLb2NbdZ0g+
fqQa3gQzQ9ImCI+6a6w43Vra87owemkpdmDjVBwFPDKgFEqUciMFvDxJuNX+d06U
A5eOyGqu35Vc/E8nWUaSTLBO7qq83JDxdhvDL2Tm/l7cpcJbeWcYmEz1WPFB2257
ebzFHPNJuRSC+zgTnbeIVICUs31xkJ9NlW7DvborLRE0dXi3jS0W9hfxgjYO19Um
6J3u3+NOgMYkmnBXVyug41V/V4c8Sg1zfEIGVGVxchfQnpEUBkOXOvWGOquD+Ieb
+pe9vt9BM/KGV1DxO2W0pub76kFvhgHMWpinzJrLluWG2pczgXe2fNgejhaODGVl
/fAJdHG/+6zj6S97YawMW5ZtU5t5Vs3oXpCRttW2XDEbTbMQfOTJhubesKjM+Jyg
Y+GhwZgWNfBUjvXzA6ZMHS7xN9uvpD88OKlnEHcwZHoUbwa58MFTnLolAvvoUD20
3km0+f5M4p0x7/gLeW9NfXCIxmjVBysA4qWPFzJKDmmbZUYumqalTg1S4bo+Q55D
69+dRJAqMffUrhnaB65RryWW7xzec+HfK5AHId01C2+h6bYasZnmoNebsHLibn1g
DkzfOPqAHyp1ytUXXSLRtxeDy4Ky0VwbkxH8vOqx7uv4yw6vk+6WcEt4ihENsjxP
fE/Q0azrT6A2o24lrUj+cQMGfAu5vP9gykv0hYNSUiZr/A3oJ+qgGUWLq3Lhrt+7
U3w12DMBhhvMZnbT7K9nOuQvw8ApXiVlsigvlgCsgsG9c78RC2IbJS/SKY+VfhIV
9WRACD4oAHzYZU8jSpfevojD/xK6KhePTJaQY8i2xeq9486R5z2OBPe/p6+jr0Uu
QCkatNTZmlyPpPcQcTFSrWKr/7zecQiCaieKfgdUo9IAtkPodJokg/fnZpiPd+Lf
KW2KfgzvSQlq18Ql1oTHvPiRz/2fvDL/6hd3X1SC1kkCV1EkWSD+gV1W4ibuQYIg
73D9rwOp8uFPOuH179od+pIwoj6QkHOWV+5B73sgPb0Zlta2NXWQEKFXuMHY+evj
z0EGDoKp5CO8wfVd6iDuGbdoNNDBYURezLyKcA519lzAZfQ/aJWZmJ5hMuNYVrPT
0Fb/9pDZfvOfjwj07bLeVVYU+OudGbVER6K/UZ2EqglcKOL0wWrCSqj4vGBL0wsf
JulXHqaUGJZsAmfecpx9NLJBzkjG0bUrLuR2NtOrVgNF7b8sD1kfi4PGFPOaiEGH
Yix0gRXJO57HvYofi+E+JWWZNFOMzxYcq1J8IVO3o0r/Mw4ZtsiEyJJ2+z4rsgfT
0MwuME2gXKahxrBk8XA/iaD4xRxVcE7kM9uLwfvrDlNdMC0vhbVRxuCQUPHagx18
UKZoqok+Ux9we62EXMdOtv/Mwbs1utBrzQpMvVFD6osUgJ7wfDEc/6bGXsLFLbl3
HhdG9+QfdUbRVCXFnRxPae4SJ4EV9Zg9CClK7gcIQTQeJWRWrdjwBoPOWO8JeX0g
cCyU1/RmxEc2RCyFUiqi1oTSSq6YOFJpg0vUg3idqh2V4YKUeaASROZLYfmnMMoB
nH9HdnF9NZ8+lO5WbWm7ikiKi3Myb6cc4K31MPmZZtlqVsaAYO12Z2vJQ7KdQfr0
FWainU/JexPmO+WEMkoCOnkQMZeHfUbaBByVUKFcCRG91XvtcYY0x0GgefkCRk+P
oKbTGdFfu0btRco8rcbYd+SMOmZ9zmEB77sT17wApnDmXr2ljnx74VBNZPMElzQL
FHgdfXjvbWKam750MuS8N9R6v3oEFr99+knPP0cLtQ8NOB1PnA71dI/XFualL8kP
ZIC6p7Khfzh6aMXbRltibTonxCLR53E4ICrcTW2lzPlO7cN5zL7w5QP4nWKFt+RZ
dSg1BOoVkyOTogODvruoRxkJCcPnsT+AS87lg1gvKrSwvod/tmtufcKCzyP7Clzn
tMl5dg4NsDqNhnDSC2l41qgn+cAVs8/jlSDkb4KRRCZDC5nQ9sVSB4xJuRL9RsLZ
Dx5XWQ2P2iRJvTI8UJ/EYw2Lz+X/8KhxgxF53kbqKPaSCEmzcVAwFAqjPNn5ZAcq
23XjmPyUTgxC25fTg/T3XuSEBb4tsgJdg3F6oxDpyLGCYnPsmaPMFDq5xQY/BOAq
9DLhmepS7u1fga0fewmwDkGfCjjx+bfgy3XC2/0sRUNPB3DEQF+NdxhiEv9mSNdP
6oXIxEmT4v0HGFRK7tNnR3ZfgAv8DFIkWXwTwSZzoiCtEAeCKt0ZUKx5wQeF8FHo
eG2arFQPyn6uR+xJVHgE+Vq3DyJIs8Dgc3k5r5kgSie4AWpZ56/jxvjz6ZX9BVtt
79QkA2PstzPavXuFNMWpPqsrOwB27gNLWhbm2XbslBWRTKLJ4RXUPBF7aM0+U02b
jFQ24Kki/GfcKfP2GuqCDYYzY/wLkJUsEIRyJwXNpIT5pmPPkZ1qDgMKfFoE351p
kgpJWbz5EKtYSSzl5IX1/MHC1XGU4oiGVc/NnXnXsF2fBNbeOod8zs4xWQXf1NlR
K55dCQFYNVy8d+H7YPqy65U6u4cEY0J+fYLcwHIZDrtpQ1U4MusFp4Xjr1EVuamJ
/5uiMxYLf6FfXAKzHzdczws+7YpjZIF5Qo2J8ZywcrlYtSc4I+4rVNRjZnG5cx/p
cIxGnhuIKJj7lf23vCbA4KpTCgWvCAEUkyelznCr74+SizIReRQDHzPikoFZRpAF
8ZvZMfDzsTXTcsfhhVvs3VkJy+WPARbSfTGdHMcTZyBAcUEvnB2DOCy8Iq8Y8L5l
b14p/w6Up56A99X4GqyerUAzkdjMCkG6zzGEjhHYxctQHmvCxcOqn6EG/zaR4RJD
ZWDXe3qrefJBSk8IJfi2ECbgc/1y/bWuCT96C920ATnuIOkgTyAnn7JoCW6tCkIC
ta1nN5JRAcjuL3tw/wJ0Uf47Yq3OiteNw8Pf8cdAehiOBoe/r4CDIIw2po47r6B7
f4eWdgOnUHgghYdxIMoycXK7pGqEXpFLdHCX2eUrc8mMKLPXTq96RK0RCSz3asOQ
huLD8DN2eaG4sKpO1OB8J2Bm67CwNFflSFB6puF52w46lxeBDONyChdFXowNOmMs
S6yS22xfOb4jhHKe/O0M33Tf6vrOLgz/Y9QNn1k9q0+H6rgTREPBqjgyKiIjNq+j
uqtpjn733s/k1x2ErB+/XoZX2kurvf+2kpglqQcyjyidXkEhJ2+FTD3MMkmsOnSU
BXS57H6QtlNNIA8NcN/T2G9cjffwefRn7pB5ELYCKCNx9BCz8UXUmXKwomw1tuD4
bUqfa7JAHYHbgj7PuCVi3HFv0du9H/CW9cDCOwmzoxmj8JsTbNzj8SEyxVdSXtWt
NyEfMGnwAuTUDlP0lC/+JH2MQIXeMnSmW0yVNt1uDK/rHj4vn8UEYIbI4q1WHACq
93eqDDQ67IAfo7cl/lDem2TTOWKbxhusyeonejSIH9MMZbyBwmz8nDMgtYM0D8iv
5t6VpEMZN35jY2q8dE+Mi8efgnGexw3ENwuuido45dTZ1dr8a98LNU5pLZdJorNC
j8cVjHXe3bGGgsmBTlBpBNqSfrU+wRt+1fkHaAbSv4bxJouwe6LeOC2rt85R8OdP
Qzc2/HsS5vKLdc/KuaULjj1YAcUaC3BwyF4+zT3HsJ8S5njj88SCmUzHnpCFhmkb
cBdUU1VGJ5r9/N0A4riX5k69riXC6bHofgGmkqWmySfFApqxz0lXFCqhSLK9hzQz
I+rkkDz2bVWBZcYo1qepV4B3dEq1YZyJEINRdlwbs1Pd2QQqXWsmKAXSXZE0Ezdy
eWoPgx/KBxBilDkuSnjzLc21SL4wEWG/h7YszirDUuU88GIqkazbpAF3G6rlcTVy
hllKeql2L620ui1+cpuqBEsBscMPidLBXFI/6nrGTCWfYqtA2Kf2vllV2Dk5nXV0
hYG+//PNja2r/Cd1Tf3mPkBwnqV4WcC4JKQteIsxA+8AQa1c7ZTHH88SOkhjKP0e
wF4eLl++RePKsa8FuRUMICJXvY9uIztALrEswCfr5A8Jnle4Xye6KnSEXVtK27cN
vBb8rfsAA/QsQC4GP306xjbL97InkEzcFWXvTnoAAPe79ks01MoTokNkcMbXX+2K
0oW459ICAtmySqPGqA3GwnU9TiwhNg3oYlIAF5lzQtgz1cfiPALP9vOKcCHa2ZjY
Ib3n2g39nlGqCUo3gmen4+JMj8P47gdgDMbpA1KmVXViHDoBp5sNOx2kFBBs5GSD
n8oLjp5Ye5qPBMXmCzFjZ5AhYoU19PYhiJHK107UIEOW954AlhjwG/osbLNOK8/T
4OW2wRj5yAp9GA5s6vodcqNtfMVpOFtfmxUmFHjlbczDXLSlS2djszeEvhJq3DHN
ehOgBzPYb12dks43nHBFQxPIu0cJdB1+nNhZAWm5TH+uAQhf2zdvpNmpQNPBXaDA
n6t98MWpUj34f8J4zDIbLpRigbLPy66xrsAb6WjJvu3VdS0ygSFwFiwneJgJ0BDd
52a0al+T1Gw2K8QQx3yXJLAvDf2LH9QqKdI/jHdQLmmhSpoGukZEVoqczq362nwg
Erj+43LFRMt2KxoOu262p+Y39jjvJ/543FBVO/VGeo6RdSWdHFIR+rTzYF7Iv9ih
Btk8uxkMQYXKA1wRq4FRgJsfQLbD0ect5Vi86uXbwz5VXltnRLzDZYFgM14tOmLa
qeT8dTH4RQj5azW+qNF0vZe15D5vUFVrbvj9vt9EEVWouN1Ov87NT3TmnIbNH12r
rVpgraMuY6gjr4urfzoUSYv1jAVQibPQJ6w+c/wSFuTNTx6P1U35ijlO2xoWVVUi
KzSn17LQfNEfX8r5BDaEKzE3et0c3YxMX9xpLHLgCchaCmqGkCNPyRC5tPUhu8Bd
yNbPNUupBk9+Li1o8qOb/ykvNSW4fa9YXztMbwiec2UdW+bFwGS2VndPpjtaCJwE
Saa/KLTSxIVB7tEWvQ2ZzCPV04TWsq8IHCmc3W12OdOeCmD0dwLzbSJlZ80KQ9Em
gSUoEJaxPf5P7YxuGxEbBrMo+s2N0AsGmq5pToukkilWKjSY87QNPdf+Wmqz8iLh
jP9LhHOyZgVE+Pggz7H7MVz6fdkUjFGsH7RihOCftfm0NTARwLKpbnOm6cGfXnYs
ktshlS2gLGYsIwks6wOD3hy4uLGgqmkp8CX2k1+aks8P9XpE1ac9a5mdwdE/gRZH
nybJVa1PZOXKbmmqf+s4b5PtAgwT+0LCucBi3aWxCgdCmYO3TiODO1W6JcPqyV9d
qjhp0XYQoIO5h+89HiClLwAZKqeGhOJ6cpb+mmT1S8mW7Adb9gp45tYjmHid0GPE
p0ebXbw6374wB0ZcPBVH5UxklU1r8haJG9ceGAz2uAZxasKNKG201hvTsJ4tSe2d
7Xhg/Jv5Ifih2QttMhUSBMkrteA7Iaa+X1z1dt4eOJiW3fLpdesmEWsEDKInabX4
hnKv3XsKM20Ocodgt9rwLhgtso7a0GyNGMGTesw89XoAQjTW+12/pc+QBekV3dSh
UXU+rQiniVIQ4aoD6vAtM+vK54fYakcCfOKx2r/8/p0iSuHPbuFVuEoBjn8OvJJv
xKW0sDun+p5IUhFHZTlOnI1ccDTqIt1hRG8TdxTuq9ySeLAhLTAI1mKYU8rI125W
AP1tFAGrDZU6F+3b158xHhh04UuCv0mc9Fb0gsKtGp/2frd6OapBdjSica97aIKp
xyXmkBztLH1VglcrY9DmKfCJTfmeGkwEohBR3+dxdvOZqo7WAjnSIswaTyLLt641
+tSrYPCFYE4ks52tjyR1VMuY5uVs0ChZgsv4+T80an9exOLqNaAn0fF5/YpZ57G1
ash3M5TYp3pyltMryFCZSM4Mjjw3j3Ij8Sw+sT3U0OR3y700RWTcl5km1fxah18p
AT7QqppQhbxzTRcurHN9AmBXnGLy+B97j6u9fuxW+eIdJqsPpO9XNgNK5pSobceL
m24GVTjSw1/ufL0hPh1psPHvHHjEn7+ElNPCixNRX51+uV1YCW0XdffiE2JPaGtu
5YYanA3qLgk4oTahc8QPLiKFdSQYMC6m+GaJUYIzs5v14aaCG0IOppo33makYCUa
pMWTDQwtBKslZfDHgcGtFoMK9jkDdC71qZyzJGbh/VK2Vlo0XfbKChjbKy2/kuPN
59F9bBGSAS+OEhm9f9N4A1lYV6PfePKiXyjR665qLxavuawZ/3QFqMD2HXuNda0K
xySlTpdZ6NWWKRq6YDLAJzJOySqavDAL4gpLoG3AZSmoWgyh/XNVg5fFbPSWxYjb
dKUQRpNFMmrGjyn8/2o1KxT4kkTfMMrZyndZi2yqRldbdRhDR6PbSLt/FgHXU/ma
rxwaippXeqXCMZgwOG+1nXjmQU8eDd/Fd177BHpD+0/MSnelS2kOvJObVpVxYama
6HDFyNxDJvdTx4ZhiU+US5mH/CPrdZW/UKl+ydQz6qzEvVrPn8ky0fCtlcErELdw
cDDYw81RNe/s1rmxQD4ihz5X71dQ3Y8gCTSu/iUiMlVTkjMnHs1txmh5ebU978nX
vF4v7ayP5TOC8d5RJHQ2URQyoANn+6wkxQp5tcEX23c40ZNZmLLyhHascFaQdjOq
jW0ps8yoB/RIjTh9U0jnHeOKMKfL0brUpbHdPFNQ8KxC2wTg/QphYEjA4EwSjJMt
wBKdZs4Ko3SLvIdAd74yo3EmSTRs7oz+1imMQETZ7Q/rcVFfbMnvq7UjTZCudjl8
QG2EVJxQ+PdFmbponFzVEsqoQNwEohq46HGXZm6OnK5BrOFOPgEz7PJbEy6gxHWY
H9wJKTXT77NxCDbw2vn7E/kAlJmcd5q5ej/5e7R/iyUFp997l+fHkjqOFNnsdPDo
pGvpaj4JbUUqlY7yKqj1W07rwh78+AVNEKuYlsR5oOrRCgipo2hMmm4xynz619jo
Qlg0vV6Iynj5L8u2EJ9IU8/gH3z6N0QB0tbJGybCs2SGiUkd3dOTnb/V+ZCsSUvz
zNEXQW7QGz1cEpj4CEHBqfkLFKuXYCHF7+0vSBJBy7g+x6yEV9k6EQZhzhwXsE6A
LOZ2I199HcTscmfociiWMjbDp2rK/Qu9N7gYQG1oqZbvhK7RrYP75bQU9uWJ/5PI
ek7q3/6tHB+6xnKGiTe2KnsBTBqgK+Lcnam3Ts+znrv2BxPNOGsABYirLEqe31LS
BrToZ4rzfs9L+a9E5fbGOMCnK3GSLWNC4rv6elpbavA9xeYbMxwBHWfky9KMhA+a
ZB177/1sunO4gvZI7UfRlEneRV+ybKKW8N28Jlj5MAbNT2CxEJW0//eUEV1cg2Fz
2WkEsrFL6cKpHbi4wF0GVvhJofna5tkIEZ1J7BGLJL3+WFOVx7KAi6aKbOa2KeQR
yQM1ZDvA5xnx8THlFloCMp5rdwzcQDH0PgjT6khhtIIyirOXwhijWU1G0q+BWMF2
81MPBT07sN6vbgLzZO7GusJNZ/GW9qk0ZhAp5ehttQ3iQYXTuMhrL3AQ8xYcOkSx
84n53GFS3tbnW7FzgmoEJT/SoS73LlBmVDIcs157ytYIFVDaYQtcUTGXgIcjlsnB
2jaIxOt6BEIO0RHR6ZMJ2p4ecF9mOzvnYTVdXXAjLKBMmAO6Ltnzu6AmFoBi8aR2
WqCXtRKAbWuvwhdmmtRsPKwz6EWyQeIjtJRPaGGEhxiZ5AilY+kfu1kGK3DCS0NX
tpL7BxEX2Y/l9qN6zUp63xDgfnlRZiLdIbnBDVL82XiTiokrFOqxbbPyCAlSYZ/p
xv1jhObA18HbLzwjJjCBrKdsvRpu72duiNc9AHpjyrXuGjDaclUYUAkIkTsEpTCD
IzI1Mibp37zm478HhY4sT6ku7rCWwnzrrW31TsOyEhvfP49qfrlEo+IGzJQyJB2/
xvuYgOVE/7wDgYSIcV/QdmqpjPp6RiHJA/UNuIZH+ZHKJcsjhWUJXZuEJaV7UKAv
GJMgNTU0O6mOHMNuLeDqrUWLgDbs5AV7S8qtTdbIq/rgi00mcjc6gBHuGD5xMbTK
0HL/oNJyYjlQclUzTQhtYiPk7Qx9ma9PsDeOW1YBrVSJ+0DQRqjWzYb8iRM+HLBD
wzS5GbJ0UG3I7LLNQnwnpOi1PPDLsVOB8Vh33qvSVX83Jdw3C//plxokvaBURnfo
m4h1AlY2WtspWlNKFKqcmq7Dp1isPg12j9A8oRtxXacmLxwztfMufjw4aT78olM7
LfxrObNAJDvjhiWoH/R92c30cw338KVg+RnC4+XQcwbkPl86XG8jDtpiemjzVi4j
TVOfREXSnE7JonpxWGcSKi5GJY5olaMF9GwQ7WN3BOyxLaBrUU8eyZQmsDWrg9EG
9gYYsHUy9OJPbsKutvtPb9R9CCwZajDSdsoDfS6FXGy3iZsw9IrQUNrA9OxK9OaJ
sT9iuHIHLyVkXtWHmN738reu3PyHf3BphXhAZcIiOioF6ysPzBhAGpJNcwaJL1lJ
V/4248/0Ve8sLcUqIV7KlXcEsqA/osLSYAXd1rCib2U2cjQR/uDhWhD0Bh/WRFkh
igHRLb0j/NdYMi5XTl9wHAPYg8p/D1e1OyyAUz1/kMU898PKzRPfmgqGM1h3xQTo
s6dw0Dgo08iFetzovvONK8V+RJCIUd0ygjs2g+EJOkVv0GCLVYdvJL8HUiQxa+ch
73Z7VqSCl8qw32IWQUcQjcJzIAo3nZVcJO9Zzn2SwVEa9OyB31+PZApet41qztjW
9+jW2OyteFc6tlIoi3hFrjaGj50xvWEOthMM/o5qzenUI+/Bdmh9oyHs/7hhiF7k
oaBfap+6CDVBeYH7zLzT418ocKO3d7Tss+9k5h4wbwdzULvhTeoUYymvPgBKjHKP
MZj7gY+rlZyjJOOyM/+S0okWpggRnK3cdC6HPcxfaqm/OggMW+oe06rU5LAgJXf7
fowKNTxnE1k/WUchuXcfM8TSldbAFGdN3qJswCx1MoCa0cDkBzPHmoXpMwcgkLOx
djw+o+1VPTI1XU5hiUNdrWF1PO5BVRtx6icr+L6d8QopEnW4xTYBckP+OHrScn0h
mMTrzxSIc2vAM6BFWicuCfxxAMx1QmDb7J0DvLCZtvbJ9el9yHrbKUo/YMr4HFno
niges+n6FuwhET7QqAOV9toQPY3mXFJC4qVA0NUrGx+4Q3uapLV2WkNKxP3KyME3
viCynJye0m4jyta/4q/b7STK6z988PlXWpIOopV2X5VF/3IZn7D31CbUFgoAx6fI
ZJByS4I1umaOf3RtiAFjAvAakpNEXHuToVOsSkUDHEWnEhGV9d5eyHfUmfxeZwMQ
AZ4gvyEowdQEMzHoO7mhXZXP3SowmyvbW4fiOC5BjBYTjuXzXfHpDXLASO0B/zAm
3DCkf6rDy2u/r7LtkSzAcsf4hPAZmKBKjCHp0Ki/MImpp5XJKqyeD4Hu74WiL+gB
d9+vCJx5urY64iGMxUTjR635UKUIAeYRwyTLB5o+rKwzbIJ75ep+xQZ0eR04KVNY
LCLs3DONKInt32FNPWBuBk6oBZ2OlXlmRrq8MYLofcWap7o1Cl9s8ZpOnN46M6VG
y2KDQJM4WKnpagAAztUhFJ3c65yCajK48xbWRQbGjWI1bUnWWJ3PsGmMCXhO8mlF
seVQxJtaywoDuTg0MRk85HrdoxheHVg9NQdZxA3RYescKg8g783QwQcsRayHPR5s
nBI+VvZ0SiYcf6P5GYa2lZj+/3Es46KvHzu7PoRaj4p7SJd2aipqWe5r0hu6wGB/
bRFxXN13zO8IpNkRxnzz5GSZzhkgQC2dGf3cMKhACNxa0jM3jcDTt2EHqBLJoG/x
Bzbw08uyfj4L6CCtkFMsdV8nbd501QhkxgdwTxDtsY8nV9lzdkEx1r5bVKin+aRN
6NIpUJgwB5G9lwRJC4LK5kP9SI2gXzga6estU3wisIhiJV9HOJPxTEcSPPT2nIOX
+9JVS0WwOLh6u/SV0tkXJNc9pTlHGs47IEGVkiAVeLRZDS/AGs922mrE+FP6uqlO
/neubnoZNCGE9uTIDbjR2YH6ogzWwPT3dqajKkJrNBa3JODWLbFs0gydQE6b8YRk
NeoMrfBEdrLEJo6peUS06ygqLoY5BslOyXF+PDzCH0rwgHdyhS7Ab8xYX0i9dg3J
pL02s/64bHv3PUHldT7eTrZOlCzfCI2SAiaL5WgIsJKKkIjf5LRUh/FASPu9hjL2
20i/eSUv8OjG09wVuGE2f5g38AWU+nqnbi5AKIWxgCXsfCcutlgK1AprzVJhEWqB
yj9QIu+zP5ySJVZOHvq+7WeArX0qRc7IwKpvji/b7+5CXVwv3YldO9px0zFTNpi+
n1tqrrklzUOwPFLSEAcAHAsa5vTPxj07xef/EwF9cgh9RpuA9mEptAUCx7lwId3f
dK6tEuQVZXy4mIU5vJJU4zOgsF1VTkhldxGaq353QMZi0FXYnet+6eqLDpkSia0k
lbaFhGbfaAcg8zMWf8RSIQH2LO5czzKOYQ89sNnhKUxGUfkwDPbY8RdvVtqRq7Ez
wWRS8N7w4jlnRFGed908RIS1XPOqrsnyD6OL3FfM+zeVsKBTGnXPu2QoPbPLl302
zyWqipqggXWJQJj0piSMW+Jb1roxAtc6fjcIGrdjWihp4dgQ0TShre841vU68ufF
8lQcLoXOZaOJKq4RYry374pE/tkcoBTUn+Igj8rWgISH7M0F8AXTUvWQZgGyMFb2
E6UYNqWqYe7sXYfL3AdQKwBvInHrFjh0Xf8kWKp8cnbsre7pfFVjSGmwktM+lycD
runGt0XKbXjSxTJghzL/8pqu4BsIPdClR3E2+DxdvlLtqM9ShS3/j4YutVN92/wJ
Qv0VnOMemP/jZZVS7QNz1xYqB0bfJvwSAlgQxtAyjDsjr/G1gWdeM5L8Qv/XpleV
OYAgX2MzkarlX0uePvWpXJ9xpDJr4rxYUriT2Sjkv/wZv9vk1hp/8FaAuRauLPe4
vkr5m00U2NgQANaXQcOAk8ISBFwP8eVwgCa9Xl/JmELEkVjPq8hdw3mKS+ZN0sWG
JPJEKUv343XRox1878zabJjbxF/tpyKlaL5BxQOpGefo2QCfuBeaQiw6JKYE8RLD
q9feZxZcLhIjinuzsAbAy4adtq1jFanI2YDeT0SeBmr49t5qrc+/6PBQ3l/Cgo/L
LaDWFtyVcFw3AmlYH/hd4TXQBuN3j9XgCsQQOEJJfoKo9GUJuRFkew7xkOfDkglg
/qxg7Wexu8USs4bS3+PzLKmtXfT5j12okIRCcqBc9yaffIAFLoeUyDunOHSYuRNo
aLkJYPG2+cKO/rKHUNc/PO375gsZSp+I1FFpmAixtY8cD9wieBiACrrHkL8KY//A
zB4FSSOXobVZHjQvFvX/6KUuTUiIpSVj5QhTGpCTlPVmAhq1qghpPXdHdIgm0krT
BWRj1U8Z1xZgmu9oUYnrfnF5I0cRdueAX8AaNDWvXYzJrQb0VEFE9sqCpK7KZdoq
OPAFWTK/+N4dJWIpQk7AuJOBonrs23HvIL5AioTvDHBkPUdCLFgcRj/y7MjAiV2o
ErfwV0QbdK/bDmpu6rMB9+IJtNxATvOF7Q0PEwOcglG0tWKBELJdTD2EYP7Yzotw
6+iy3EkW0GiWdjeFXJZI/x/nzs0/vcEXeLpa9YyNhIXqaGCDvuoC8vUPr9qBBwvg
kI2lLibbV8zkhue/F4Wd29guLdb/XYS1U9p3/9OQ5rcZTiQJTXxQuGucdAeVgkTb
OwI1Du1Q6q0PtFHlQCwcgOCClTWf+ly/nkfhEybYo9StaVr5ki8WqvUX8VRafKuy
KXS+2WKRGK6ciRIMTQR5ijJjExQmO8CJSHwAVzU44Dtz06/3363zFq1TGZMWLmoV
67H2pPjZxNh4bsSjoLWEINq8u68C4wzkcuzrDNMX2cer9WVJJ8WGIgnvQsOz2ibi
Xlqk4yb8BFce88JIsO4xqvXnqKtp47RDkWu5Y1Fd+mccnAuDhPaSKmI+67vxBeCb
Jqaridz77KJV/ivw3MFf3lxt43U3lJHFEstMhotwq0veQlcDJg7UqMQ9h6L1692C
3ZabiaCSYc7HMbtXFibiEoCqlCNrNiMrVjWaEFJGq3pZjsM9HrchkTmk7YJBB9ux
oYndv0jdVBLhXm6UClnkGdJJEWDUHo5QmzMS/wzhSq+tFnvRuoFvsKDzOYc1MoMM
WBb7LBd7xaeQMX//G0f03auBbhz27xBXi1RSyIhAL/+f1uurMZbOsqQIwZWJJX+n
VgSoKAy3WjwpVTjKA1EZBHOE2JfRVOetH5JxiwEdYvM+sfmyuXyGW/4H9wQmnqYU
NV7AX9AXJa3TZ+ex0Pai2gDqNl3Ydt1I5UA0FJT3ikWhFwmcuCO674IpMJx7R+io
wMf5pZcHznl7JJzXoWp2RjoNnzo4I5eeHazIIZDKpI/132y1mK3BCuDiib08Z0fj
h+OYZ4GP9/4WABY+ydbaHoFHuU9i+uruDfVBKsihdzUjb3gvqKSrb8w8uKIcRh2E
2Yh3cdFCFide8f6JrMjHamuVeGBBb8mS9a7aK4xkXMs1uPBrbks5OsQPCIMbJglY
i8EE3TMV5NIiCGRuLiEKGwrI5nPMGIoiZMbjHDMIjbNwtgZsk+t975LiwY2JVNbO
BMaDBHyRZjvYrzhTEBdUfkzbWYVYbQH3Y3vHSlwejOxRKU17yClk3qa1SFp9r5jy
UPJ8XHIBNTSGhn31XJe8vh+zG6IMbAo1kWmzKqjxlDVSvirdUzRMQohFndQi0o39
mir6QJuniKQjGyy0x4A3ycuNVu569m3gFJdPFF/LUASI0tlXnDm/HV6RKohpsDfF
W0Qmz6xNCqaO7WbNqTPYa3L4QyfhgD+jZA6FXEbIYIVcQShJjrMo04g+wa7ruddF
Pp8ob9/5WcdgPw5p72M1oVo6dVYQbEHT4EJQSg/FFKvxLhX0MKJzxQMb5k9apDPe
+Wt3TsBB3DLXKhSw/0AbijNyEKkEIVlwHb7qeaf1vWQYbgFrJH0G+dp22HbUmCWA
OuMZKTSKWgfPPBO3jz9lqLM0UsXCEZgjZZfXpDMzcUItgtrOle9wd4VYm/5y/1YA
M2GM5tXqfN4Mril5NxqphRG02T+EDA1JKry3BR9i/KrbUxgdFxCN0GLbhwv/z6Pr
TqsLGxMfOKGmKJenZyaOQVylSylvovWJPl0xdVYsMMXzN/nUvjGbuhqQWebwMYby
FkzunDwJT+4vlAemEPMozjUaZr2cjwlpN2gsZRCYyX0hsXuYK1UkJfq2fypd2ZYm
wcKfNgo8+Y7dsIOvUc7Jpe9RacWc0i12FkDD0NDKL6fz7g5M6/MjgLAsCUur1+QO
GLz/GUkSQiEt1fajqEJdSDhUVJtgcFp6OSaJeBgIjoJ3d/nY/BguXRPOPQKkO+oR
lAa8OCm93zuX6KUGxBOLjhePpciFK1E4Jb4foHBF47HO+3vhNaBI2FLtDAXQYcXM
MMzzTX1bxeQ7r2Dbf1MPbERsQDcqZy4nutITtoivXXWp+qzCJ6b/VgyWWLPNOYba
L/FKyQ8jrLEinb+rQ1xAZmVkH+6E9WlSXkSbCLg4J4tMnFIZX+vc5WYp6BcOLa+u
oAx5MtR+41Sw+mPsbPOm8K8QIJQezlzmkaY5Wh/1ThLGVMIGXOrPyKZFPRmZLfG5
pEosURgrSnNu+qJdgaTjnNK0dazI9VsKN1rsEV/uC93ZmWj+SQzhPgdXL2USBHoU
CEkoFcrO6CciwdPl+zZLXYnPPjHsufPxTXVXkpOeS18AK6TtmheVoOaZSuLJpNxq
Ve4HmdVzbE8W0Uq7ATd44PY+RICQTMldMPf6uuQ1sbOai4FlxgjpCaYKKOqz3E3m
Mutkscyd4kzyVvQBXrfKGl6vdnjKMaD3wt6FO6xp3aQn+PQ9221Vb9UPHooeG+4j
UZUHIyj58p2PbBIdGhTkYDm+7qjjVgKrnj+p7xvM23pjE2G3Ku1FTnXFW4iWrSEk
7VCdOLRiItgXwlqaqiJRFzb4ISpFyLmPUBEssdhPGGiTgnPZFOsBrVrmOnjKGcIC
/w+bz+wos1EC0ww3E0mzq2UOfC8tUhSTnCPOnJ/dhO3bpVgOEvT/53mhz1fQIDER
jPdneJ3TRF8ZXMPe8AohXap4FkQuxZXPflOEoET9w3HgO5HYoiPUTC1mRSv/o9uY
aCkc+vxjDEGXfuhKtCK7a/2uF6Foe6s41ge/leKXEWwMV+DbxPPNBDRxxVg1ntwS
bzGSoZkDPpXa3Tpf55t25QzVk96wGKkTfmwu2teZlfcRx+/yngyssP7v3IrDlYzm
mOM57iUizqaPKmPUBM8aNtVLLxg++OaEubanRwFdjJYo2mwyvZ3pNzuWil6j3YbU
+M+xrAqbQnsZyEGFxK1McG4jdrJ85aTBsUx7LmzwTn1cX401MyV8HE4lOD7uvCti
G0nfF0N6pPl5mRiXMrCdSpNE71aet+VDjW1cjtvBtmGyOzwOPxH4koJjyQ/OFP2F
+X+LluspEQIR039u2aSsz06mkZkBlXGQjn8lWTSG5NXES4kxJPGJRtZV0cf/d2EA
FLTamCizmmIRmHS19C0In5sIcqVXeXA7rV25BMf+hqTqGsZiNaiktUrbjAz4OvdO
m8eGB93cv9+ulnvFvOrdZLU34NvQhbHlIjWGqtYOKLMB9PRZVTIeCVxAnJzE8XCg
V8/cAx5TxLMgW4hfJ2biTrtcIAk5MCZsTcIeERRE214H5lDBxR+1nKYT8RlLN0Aq
59OZcMFM6SKi4hyB6lCg9RPiknFeEtCdDf/1pfU6P+FsoA2uasylfG9ac3eQtLQK
YLdAFOOGBB0QMspFbv4OZJszDVzOVS6TihEDQkxc5T/qZSfZ9KbuA6p1ISqFHoVZ
NyXiPOQYRGmoGyBJY5d0rai/WbuBbxhqWyiCXtLAgZaFrFibuklMZFudKsa+1XeK
oFCMHlTzIkX9rn3Rk1iR8RpB6yPx0427EAQ08UlsU7GHQGsd1CBT5oUSbXbKzhhz
i8nAmYrNQ07vXEtWwjU0t7mYX3pbAplvS2idkuaVx7EUROBFGd3+zVO7PuqyX6kT
0sW6FwNtcnovMjW6fanEazVsF5JAUiGlmV8LEBXfk/WJ0GE1JxEBSYAqWpqx+IdA
8f0XDQYPjqArCGwLTi1/1HXQPmOkl0hVhEQwV/3yi9dc8qoyqn7h/ujAJ+4ODO2s
jlEJFi+8iexi7d02cPV95zZOazaNU40ZmdQvZsd+eLTzWEGcZP+Cp2IOX1I+UZ+H
pUap/3OWn54Lbd0Fi+ERtHduSKJMcsmmWRp3UfFaKd9xke3jdUaGrM0gebEvej3u
finGo8czMEk9UBlkNhR90Zws1qgbPXck+IHf9LxmGL40Ezk3Ku7ryx0+oIYiBqZ2
CG4Js8upO7dxY7/2iokO1UFRk7C2sNKTbsUWfWcom0FmNwQ7hw7EvsEbmmgMBLxi
B3D4Aeu6urNiETn72lcrws+EZKFbp7SCbHi5bQ6skV0RDHYV3PvpqDzbLVEfx9g0
f+9FVME9HWWLZgLODTsatTsFL+8EK0YcIqxmI2g3bkjLdbnt4hWjvun1oVIsBH5A
+g2SWnlLq6Q0lM0d9p7uW4uF08UtfF03diQqRrB28DdmgRGdiWe/qyD35LihQRZZ
RGZvWXnFnlnt/uoHoKZ0d4kNx3ZASxLzS4mP6TG+oN6v2DaJDksyNCWg0XrkUmuR
szKdIFTlkGlDmoLuguN0FaqDiTksXN9sa8NtaeaZuN1rxTLGI/8sRyBKlPiXfUMI
6Neq7FpAf2vf9NFvwL0ffYTGEepz9mCZmZAQOZUK6FLENk3MZc/L41lF3jQyIsVk
5WftTpF7LBeJPUHu1lYnK16nUb9WGzuTTHXn8NrMMg19x+Kdrjza1U31iRDyk0dx
D3US/bX/TRY4k/4AKppRjQld62Uaxht7fTvtbFXqeehw6YaiIcIC+tclIGg9VaZj
zj+ysDc2x54usDULOfhNNHzSoD+2M5xD4IuJeedOHL3sVyKBHtlLjn+VFCIor2y4
Od0WVwmuxUb4yTzUzVIc55rQLvB5DphE/idFCGaKcLbBySBQBl9HxbXORNMv6AEF
GMQuuAdwMiHNLOTaczWs/wIcAIS6Owqtl6AIOVkz0p2KFrfreJTWT1+72NGevC1l
4+cSMD61/tVIvMf1if8aIPzAnmk9r1j6+xosNu+1q5aeqMqJ5+BJvFKOgwdmOGL0
G9opEtFDKUWi/jwQTdbDZMub+ZWWCuKbUHKfyedwuKCNhOKJb7y7ycduBGpWj9Kw
eV3Qqg+2Wb/Dh28J7vC/a15Y9SnfLBV5021Z5prDjCikO9DeOoo6RfZy1duZ2KsQ
M6wVqQ/AXvuuKQzCAnGTADxPo9O4y5l7bx7U8AfrVaVbkblGhiwEEx5NqRVSRb5Y
NFIADcqEybMd0XWQ/c9JAzsTbI/53pbUQOTOxdUj9Yt06t16ryzpEjHqtG6ryLXe
81EHZfS/fV+vgtDysskYpV6zUxOKBBwAlM9PZqG8vqq8spk8h43y26ZPo2eKzia9
mvxMGB1dsYXlaI9gkXlNA0gLJ+IhE5euM8SVVYyEB9GivLebSATTAsMDdH0x7eom
afSUW0flJxVcy2qrVew6sUEP8/6il1Fe0MI10tJSDVs89Dew5sH2NoQwOQqWKorO
m4kZb69v2LP1i31IYptRukVa16YAvu0XandgVFLAVIW5sK/kjZcgT3WBwqsHh+lD
WNoAIE/BoOKSKBNP4M+l+W7BDuHCINoTR2UI+8SxXCQnWFld7k8sATHL+mRfPMm1
WQW8RYk6QmjTAgd8Cdr6uEIDzsekROd+AlhvOnvdzDgOobRcaL32pscYbbEVSVMs
IEuv9vr2Yx992BWIZdDRP2K77b8panY9PqR0pEmAXHQw5ECznCxGdYZBkty9fSwf
PPiHLApwOTRjkkuq5+kE7E8+H/e4x/LQ2t7N1460kCXqoftrfake20fcvYMA8MRD
8uwqSn1bYfBzSw4mLvKupoK1Rw9DXwmRazpCsjpTZwaMkL6BxZVW6oKh8xnLLGgB
JsmkjeDaTgPAHrE1KxyT2Bunla3nrpOuKZT46/wob8bqHdT2uU6g+TKsGRH+SW5X
HO5MV1eIPZCLMXBsiutaeOkvFuioSF9EZtKvdMNrgcykRzaAx2uLmOpwjyo6kAxL
YuUlwTiPRd6JeEHxk0TozMWXLNf3PievZiT0XoBSjTNNke2B9iRoc6o2JPO3ZjbM
nmKlxiIwjY5LVgGXhiCahZbZ0xqZb1Fuhe4MaaTbYi3ALBRclLRcHEAnmIzrLPvi
hHwe2MHcLRdUitm7cfUkzfjiCr+9FK0Qp7hvrFvsXa+xX9kKifyktHI6AFiTPwuG
ECvi7xGIhI9OZALo2ZDZhdwwqfooGOigyYhs3M/qjkG60aFWkC6GeSZVq4JEGIfp
1Oyt17EBEOQZCqkhjx1OaFgcEMenagv5uAS5QdFkikJfuhJL0kCQuo6TJF5QzLrE
G+4WJ2L7271GyCusN8FJ1Ap2DebfcWp0ZGSums4MkbXkiC8GRXGXv8t4JpS4eq7o
0pnBHhtQPGmMEXTauik62G6gGR+zY9gS0D7M8oMJsBV5UYpM9jFIn2pnFzJE5lCp
nlbQo9wZebpoHgYAiHWI0F86/gCmHqhr5UTgLGa+3Lnv6pJPJeNM0rPpSt80huof
ywJtgyna3v6nNIGu+rn4RFUUtOin6fTzhzApyb9V30kZ1CpW5mtHCV8vQqhpK2bz
yDKI73XPM7/MMGbhrzxMFDhlgS5rC4Cg9fnfVSteb1IiEit3VKrHccIBEkBwE+CW
EZHAy3bFdYfqWASEExjV+ukDVLZfc9fup90BkkmTCTGRXf9xWSP1bQ1ST03yU+GX
Cn8hu9ZUji6RMSSnnNih/DzuAADKr/tPvEQIQ6L+72DBUZ8vbQ5YONLqSyQr5Bc0
gZkFRdbMdlDMy+H/lNmMEkrDKl9weSZ5uElQFdBCqlKp7rFy9Jl4pi267PObokhL
FbDdmC0TKqjcq4rdSa8EfVDANiidEkBQxbC8lgU+ovBj7UHqXsqlYjRDWZRmc1SD
PPs5qgB2WPvxK2CmIJ/hk8NVjJxL+oO9/nZH8+dfkUn7LEOr2sljvCTWBrfCTgEB
gFSNfDckqM/OTEx8/lTtXpXL3nx5khPrH37ztipHJzG8rv2OfHcy0Yx0rEFmqaBR
AlB8T0mKkAeeHtZ/+0GDRajDSAHqEKs4sptWlSMo3kp6FF3abBHlRpw/xDG+M5vB
RYVgZ0EQZQ79qjT7QisI0KF2EAXuQGUr92CXrZ8TfaEYycM9H2sqHKdhAVmMOaQD
u7dOa5vN6KFo1hF1quT1uyaQqXljYQ0xLMA2WXD7i92wNLqfFW5DYSpqsp2/AD1I
Y6XGJHnWR1LNM8sbhA1rW46F+pME4BM0UcIU5mlU6CqgAHtSVu8ccsSrsz29PJKx
K15mMdNWCjBdZ2Wtpl1h5Et3vYTyl2OIx+tBV10/+zp16L/1gdECAms3QsXmAZ0y
Mwnct3gGoJ87gleLFbhNy0jjOSyOUhFW/AzbEPgx645JrPOrXO/VWE6Ra6MhSzb6
JT0AbRBiV3R03bOve5hl6ukZj+UlFTa2Zeo4ltJSePJuzdXqUKlNOGhFHYVtn81Z
OqDVMVBXBqwwbSqnU7xhP1CHSKvGOA+6MY9AGVDowkfu+7l1AOutCSQR1h/QLph/
+VAM4M508RkcKAa9kthNYlsMAlIls073Uibl6F0j5nD5bc34BuCTkZf2GApArADE
yLkmRxz8nnQg66Gkrr2SuITtlI5mC5PYq0BGoaDRdkvsdfv7udFg8XnOa/cSdqTE
pmP5yiys1rVTbF8ggkv9YmBZoqseXUpqn5dwuaXbAGhMwkxNMwROfdb8q3jVLmPy
v3jUqKiQK3ioR2yBlDbzD8uRjlh/TJNYDLwYxhGF7eiDszKmkyZFizXLjSXAQfUk
GgiEeLLZXZ3JMJiCvmUhwzyfeUkjRlcoT+w578gLY6z2kmUclfP6KHv02JGl6sLP
Yl7ilVVNoC6aINtoxFtA8EIZDeceFYrLHz+U25mzN2zHvT0pHz79Dttj3l8Y2nAw
hLw6/adHg+rQUZahNJC1NQNTp0HG4M86Azx2zoTQFNuspPhS39XD2PAlZad7qUGi
z7Vf71MpUM1PwVG+jE0yLCVS/40QqkHitAWD8bpi1+rQBbr6+NP0objbIzfxYwOi
TLXB9fYwbKHetIZckOXfXnE3q8jsfAI3F21/XI7D7q4KzjE5g1Pumwr1naOycD6/
JEp+QBHe6P3JUJp5xr5b4kbSbVxnYCN6vMvRJT+a1xlp+7b8OQnxb/Cgt8viPGEL
O9DnZmhL4R/7e2+RU2U3VTooc9VFVws2zRpFiUNf+pNGbEnHYJraDqPnndVfMG/a
GT3Ox3Y7iR4Xn3r1WxRi5enimzoPt4kcT/SxkKIB8oO9RbpjCHY0tSauVxMsaLet
Pr+BKm8vZ8eBwcK63TdrLLxSBmb3H4gTp/XDnDSZ1kzTWz/KSfmBgoFBmC3OZlcV
S3x4QZ9ZKIc3GPuZic1iMi/bBNsPaVpG2DvNNVf0ysls3OR9qeGnoYAwCcIAhDEH
DVf6fm/Uh1Fy5gCxzUKiK9c29pPm8Uzqq2zoB7KQ3QdOW0KVoZgIEimzGyIS88Ej
Da9ueDsfxrxrXINGHwCHGNhzeIC8LCFmvAywz2p1+UzGqzV/6Pe/8Hpw2uQxJK+/
JnzlAttOVLd418ZnOWhME7hyOnu4kug1jlC13pFD9CUlEhFmyfcw96+4CitwGZOE
inbM99ka8oU6GCk/vfhqXICNjTX0MZhnOWZichrA33ga7IHuIeV6QkDNkMfZXsbo
F7H2nlJFg4zWHKHAZp0WsDb2Vx88n4aGxDUCNICmm8g5Ob+fLF7O+Xg9rOkl5ZPN
uhvo48ElxWe8GlA7WfCmj8DoUE69p3wU8ZCwaXQVZpGc1YGxvQgqIOWcf899Jzot
fJydQJpMrDCheRkawydoyjfjd1UpG/3f8wCFFkJY6wkyWHPyhZe8OqDH77pxdB/D
YUCE/1tO7eCkFeRxeRZY8hWCObDXryJXIf07kDbcC//uIIioc8/YFxFR+sMkuoEv
dchzZDnWUMgNkz2wrxU0UmQngyEnTbKLMnbw8nJg73r0jHiTu+RDQ28NlFXLXg89
dUGwr5qnIXehsKw+Up5R9FhPjLLgUE5E2mHw4rW7K+JBuHCctBqCFsDbj7bwGqJT
SFN620YLuow9Sw8xnxfg59PWgxtvSpTCROF7xCT+luE1ryoPIkdR/a2xOJEhJEjC
UWcL4M1Nv/aHNDX2/BqOpHw0QT06yOBBAuHEzI67WiJAYz4E9SvLX4v/1jASUoe5
ee2yOJ+JOc8C4MOoSv9SIdcTivPo1WhE1xL28oybgPNcgEVMmW+hOfUDbUsx1X2+
B0mBiG9uNh7E7O4ykbPbR9g/DOyC69++BOgNBuFAm0iqezvIsAd4sHuAD/I8QHjh
QGMUDB6Z1R/2bLVd9uWbwwFlTrLXpNZHn2giX7LEBHWjrQOLYO6JB0cwOeu1p7BE
pJAJM45hxQcW4xAKYWb6AjkpUt3h7eHJ+cfJ/Y5y2GV8OiCHus0K856x0qH5wkFg
x9u5cDgTnzzMpF51UYah3NcgliqTo9epGYcIiMxlXJ7Y0V6e9QkDyLQh40+G7S8r
ZURCEeM2GgpTEKwFhDRcG1OVO8A8IFDlw4rC+6Y58u1Z8O2U0jMhCOdgfBhQ68MF
jM2UQYjmjC+z+xCTnEvOrd2/H0ryBmwTXArx0R3KhuQ5S6iFwI2us55B4nhq4Kks
z/ohaimublHEAwwQXsYpKAnlp6wqR9GTeti/zX/I1Qy7+3FOnUztaNVflWvt/OaD
kKp2CmFKBHan/noqfTQmNRrrQ7mwTzpGY8b8XIwO2GrBDQCXPWsPGvF0SMiQj6sJ
dd4wpcPQeMfLRougmnGfapPBxeALckPEr/FKC8WPHy8IyjTN5taWw5M5eLyn88AE
FJ0xA3hv9OihzS7jKjiGvIJNWOfj8qLmN/tn22ba/gUH3ygkNQ+M0+Rhdz2zthTl
Ws9y0IKG/V1K9R2694KumX98mif0IQ/70QHOP/bW0PlktCr5lNmwpXh/GMAbws1W
1eF3z9RbveFHi3t/I+uzYY2/ND6mGskcNHfXgR4Oe8VLEZMiH6Q7sZ5uS5/7BwbP
BlwnmiZjtela/mrUlHCqGauGSWtDsjMvCAaDniXMFXeRxtqAhSiV8iUr+H1zA9TA
EdsfDexWTH3k+zvFQwWKgBdiu5+Ug7PAPxyqnS0W8cN7VVpWMs5l+68X2ZDdInKe
BKG5lphAk96G1oQB/eRawNYmv+nHyzVP8SWDV0zo1Y66AZ7Dt43/EzK5H/Pk4ycQ
Ar3h+QYY7oloVHyRX7Rzd7uS3AlzY7cWd9HhgxxVexnifYO911A4dmfV91AsEjPA
NUIgYMuj6c58w1uAMx87TyRCXKUbr04Ml1O/DZUSqhnNAzcm+K1lOKXYUfPuyOFH
0uQQZk8N9cpL77vE0a1eDq/d39Tbmd7gDt+WG61JZ93XLd+YgkugqfB47gM/yweI
0mwTf7h/Lq+Jko9RAkrRQ8NY253b9HaAOIvAmjeqOM6ngk7Q7frMLRFjZ35OWU5R
qzoAatwk9HJ/Q/n0EDQKOH5+ZfgXv0zCN6zJHbbFucdgO3lIun0+HrsnOKF5/FQf
n4dy57Siw789qeS/1EFXr7R9NPpN8JrYHRiQ4kG6s3kO5b3Fs9Mv252OVeT0NSRk
bEeI4AfLJ8T+PoUMXyDVE/qMZVsCroyjeDf2yibVtAk7ybExrghMu7fUyzhOifGp
0F1JDDQwyOaEaz7Rw+BjpcVjENyS8MFYJs8er3DXbZUWq2IaW3zp8NE5JWK18lA1
eteuoIbEL8Lv/b3y7mtT5GgloivNqdpsGa8+DAHpnS1AXQhMpCSjOHip723S/VXM
KtMqjmItSTLPoFbW/9Df9/fV7HJWOZB9bp8+IJSoIvhxsef408LsiJgQoxLQcnBH
+Cy0cBHrHlcjUPDuEuYyUO+QSo0lwiI7WJmYYKkgv+EAz7pfK0KfIFW0azrzzlXp
RJRDEQ/K04pv7DfshLPudR0Ul1aHWBPuYH9ed8fd0NRxDp9TF0yE4hk0Lk5jqXkq
OX+Nkw8kxqWEtMknuGeAPPMURF8CgP+n4z9FqdxBLsKPSo/xEDpCpmh8Inq0Rgco
i82HJr/9Oh7wtZrU2SOpnxuZvYT5Z1N3cM4422rOlo7NNB3OucAjXyfDRLaMuYua
4OzvZEksIBiZvy5OBTyJc3BJ1IMUr+D4hdBaVaxyk/w9DTwZ/VP9+I2NJYUNPBMy
QG5g7ovyCbqXp6wbI/1Gdc4Z+EsbzkSeHiDPilw2CmNFmotMt4l4t/e76b4eAhQx
QOw1w9pbx9IIiH/uigm1ucUg4SjZoZTQdfeDeZLrpUShYEORqJJPpS2i8E/ps8RS
QUat0EJxL/ZZaaDLMps/xcSfKz5TPY9zryYQ/S7n7TlxLTZFZIjOLIicTg8LminB
BsN1YGU4Q6fIUrcNLrpEpd0S0G7rh4BBshmkgKgTqBCGW/Aif/R1QvxwyVYZ58dd
0WXfnDPh8jCOSg/vQItD9midHedfnsxMFhFUFfNdBZZY54nelQBIdYM/SIwKrj4U
xLnvBPPnC+zRWwPwOkcc70hdCPtHmHobavTNZ6mq5VasBqOLs3GD08DnJajvnf7S
FRkNejyuoezt/0cbbnvQK+gx8nNcCXbE0/e5+lMj9WMThcsVqwdB0ceDl6u+AVvE
oKQ8KSHwj2JzBho4ggk7tvo/h4TWRi1HDTtCBtXjwl+UH+888Kc1DQTDZS57hl0R
v0RcJN0VjRjRYW+1tsOVq+/flDy+b09pTwmCMiAul0sjvyODhbGpxSmffjN+eAEJ
oucrqfYcr84nyeH+G9NVOhC/iJux6qmrL+QFCVEKEch4VJdKcnbV+LVBSRfIkJ7X
6dChVy2xjp4cYY7GW2vnhlALr8wX8OjeeRawRlHk2GF7lAgFqo0mvNoa5IfwMGSq
20N3tMFW3CihP5r5ifovKVdwKAhdEzzgqHcT+/tBOQM+J6d7MbcB16R3BFraQkOX
aAwKDVpDEB1RB0prrXdzwkdquZEU4s1rMT3XbIXm0hsdp8sBBtElPC9vaOhyhwlA
W0T0ANi4P0RTa3Gdr2HchB7kb0K9QHrlhwgFSF6MCCHZUdAfxRDf5yCEiJJ7QcMI
j5DsDjOzomVAT6wrY/ospsM/JqCpcDu0vvHyEil6Q8voNfL1R4cgsyhlMA02GDWV
9VvPBxOyOMyy1FbANHTiKBSq4B4VhLDKHdZyHOVm08/PFC3dnP8f3O2tu1/s/cOD
rZ1Tp90CpWH7zq4YKtL3IYEnAyupmfkb28oJ9HviqdGu/eGYNnkxGI8QJXLRmXEm
iJe4qz+URFg5cW4dgwJI5P7WQ5Nk+YECFbyNMIPOTKbT5tqUIXAAzfFDwMPk8yWb
6tHrxklsgwiEkNbJZs7G7AokeEgvgr2uqt0jCYzEDaa8dqjErNpT1mMV25LdH2nu
gX+vokNtxsZvGjhTw4rEZKf0rQpp45vDRlU94EMj2ZIXv5Ck4e5yKcTXQVclU/Q6
fKx8pej1ZWGDi0IC5PFKGgNZYDhmDIgcqhmligVRQjuVLqjt2ZBHlUXGxQOsVfU9
cWtbmBK0GjFinSn2UwgiTcMeZOYC/k9XeRNL1B2kjVuyCGRylFsUYgJWnlGfCntw
iaxm6sO1GHg3kmn6vJoPD06Ax52EtJn64N/+Y+/g0pQK7IaE5hOIfje25ojsxZ4F
asJ50N38ufsKdoWH3dKa5pvqn6sa/PoTj4pTsTQiLvlF/BSq37c3gFITT4l6t8LQ
uw6NRyI9DkxG9qZ7IwDIuCu7ugUHP+cThSNUFd2Zk3IuhSsFkcllx6dNXGTNOLYk
FuHf17GYVC531cyOZGUd9yV2zv2Wr4IxxmHtypXSh52GbMwr3rh07ATi1Vcp2bkp
STsN0JVrh7shgFHhfJNFwSpfusgAIA4RevEgQiivY0cezngCHWaQPPo7kTM6qy6a
2cwKdIGD/nr2E2cJrsx3lcNz4QxeqBeKshnLapXEpTkTI21sU0vQw3I+BNV3rKuB
q+CUtvIZvH8eoM5ECiQ062ArG5ZvHLnHzJ0Kow4TTRwz4ozJxEIiZnnY43hIixyb
8bzqZgkjRkfXeIHVIimheYMVfRKZQK3cOhbPHJwvEdRQHUz9uw4DbafjHsUUB7WM
+HU8OUkxyc4pH3Fqp+X2003nEttk79TOJkBrp3vWrHO8Mte54uLv+RgMA84XyyEB
/0hNzRW7jWfNTw8bo09lZeKBznOiPcWdCQ2GvFxANgIY0q8IAMGJ2Qjq2ga3cX9m
DM6NKMhwvOmFCepqtCFic+vdP/zXg3iDhL6KG9cchSxyYjVIZY7v2IUuAvtz9VLQ
lnFZk3rZjXIEa5SyAt5DtovbbbwYz6O0QBQCBc+ak1kPGFF/HpiDzsMTmPfwswfh
PKGdmwboCYu3RJsg6EF9eRQpyYFalFPDJIcGDEJMCNLHkLeTa1KjRdw51ONYtzFL
SjfzGeTRYNwWiqBzIvzmZjgl7EZw0oFK5RURNQt1D9czJ8MwGSxw31IHPxYNwo/q
XBivgjnyfVNuO0K5gl2/uftjJxd7liNWWK3jzqUDDV+ch+vWsmC8ouNaX2VFfIDj
GR4sIn48n+/u9LDmb6v9JT4s65fEmPIFkRf29qiCUwhyTr3U4AoccbKQvEZmxW3k
rNP/b9AYbZxU+viWo0uqwNtpRQeZWp04GHaEzwK9rGyUU7v0caVHKgw53O9bH09i
5kVGcys/5uEaH3aVBmy7Lm/xnRI5XZq625x5anXCjyKFvMgRdE5kqOWEjzwQvcFJ
Pc5Kh6k3gjrHV1FclAky+DVsJu/mJ6akVPM3kjezM+vqzROmYya0WEHNA/DxRAyS
mVWQh3B9Ktwad76liwPuENXxWvSJL3/633Pu3+LnDvqkS4iCMIbqMhLJrTt4WAum
hso125OSBLJ9gKPjt3INU7sf3RI1QDTIiMu05hxvcFvLbH6v1hoE9ZvGd2Pk5Ru+
ASG0U9muyJvajN8r7ti6vHMqOrxwrgIXynyMnHWhUE0ltqsvT7x6t9EBpyb71uOg
GgzvGpqh08kHpxJIdTidkCYuPzU4B55BbJ6oEzvNVdZD1ElipbqRBjae2NBzg8a+
nhHZ8N0tfGQMO3WDuatTB0jfgdiMNkbyrdIp1GOmgqImx/31ll0DC8ar22i/oICI
G9uN61KTZMnsLiMlfAvnVGhsU5rAEO8kgqei/AmBi+49ab4BOeI0obyKAQWg/Msp
Iqi51MflVTSfgdQCQcbooFbkuC5ygIMLPbTTdZ7i0dHNxCGicPkuvDs1GY0S7ZIg
YKX8Nu/lhAE17y0rY5yVx5tKMh79CK2TJEnPrBeerlIJUfwOaCenY4XxURj4vMnc
whPvH+H0XT8Zx0n7DQFL93VgS20Ki1jluRlKjlQrlUbfXekddMYhpKaOTRwsMf4j
T+74giC74kJgx5KycwaKSrzmt02IRdjxv0VbPb9UBcgU762TV9tqVRmbT8NsxK4X
lyJtHzn+2hZ+80ewCQwE9R0b5vAeUv1HdWHa68mGNyo0R69wmeIMMGeg56QNheTO
8ngxH1XmP5Hh14Xx9QlDkSNls+vhlWIca+McvFnqoeCzXlTo1QJESp50MSr42rrz
89zwAZba9nHksqEkWnpXkRG9QSKnSjzCPTKopj8z/5d4+/xRsNLqltyzGL0mqKDj
TO6DpFEh17iUJBxHetJkVnjxI3aMvBfvTvevRkDrfq0pTRNmgnX2bLMo6BfIRfjp
r9tR/iard9co1gha53pnX1Teo9lchxwihyGNDPaKFV/WoszOotsd3RAFGNlU2KxB
gxgPsfQwKdKtcRBqT5n+xTfEJ+O4XkHTMatQPT98smcVR2zT9g1eBVr5o4CbTwTB
zezWT6YEDdsXW+GG+U1JULl/78D1LZr03YWGbc94USHJYTiZIMEdbussruSn4d3W
w9Ein0TSaSpUWSVf3WjKT9GcnXUhyAXFUD+9Alng1oQPBXyowWQBeNHNuo5rcBah
G8xJgWtUMfmWKKLLpaAvr1Hjz8Rp6bVuO4VmO/JIO73f15ABJbrLaWK5psRJF4Il
ramgqssY/oHa1iyPCO4vEl1l78iQMmpEHQgiI6UJGdTHKPXu80AMznNYkwE2OvTu
CWebxywK54Uuhu0s6jNIqrRR8VSsZp9BFnahVoaM3GcXjJiDAmVPrNvHJGvgA+Ui
PBvfDwA1QgGB2EXsIxEifyUfGUttgbECZVf5QSo4ZfYyeTV0cTAsOXIbe1j52HK4
9DwWVh8+iY3n+dK9dxOkDiW6cJYXmGLT8mUJqhTafgZgLiIW7/2h7YwsIdSoS61w
aI324lDr/VcmXkm6bzQi+DkLhDX9x0gw2mpCT9ePKv7bM+ouowdmhhFRttAWs/d0
iF82nncNBMHIijYaFltgwcdAA0uQGctFgzUWpEgc2eQ1mtHMbrn5Mmh5VXEU3hV8
vP5qaSfts2k9ei05POoIGy7x9mthrKzZZqMvyRaTOAgfc9NkqfMxaXA4vyaoChDf
436xboUq+E7sqCpLMFFAZVgI2f/t9AvlRwd6UkhVH/rf2OjTqVQfRTadhIacYWqx
Nyyxnrzg5C13KZtt2QZgdPua+fm30MMwcav3cRiFuFsZhkuY0tPos1dKOyBDbHrs
r4ew+plUZdXtwyjbnZeGJoMS15eOERfXGQb45qe0y3OvlI9OPZLkJ2wWSnCjutUb
tDDJgFVmqPHh+CmRyWYo1LAo9qG15w/8NesNW+DIGiTCKQh95fDj5cZ0fzTGlpm1
V/g97F9q3E8abUvsOhLwE1OBz9xEh16aS0BknHXqx+ZMmsaSFjs9nsNMWOkm/0jH
0IixSJCNJZEe1Te/bUuiHF1yPYEXbnnvCAXh7dulk5310B8VYTcKuKLKjFquCeI0
uTfGZjKitpS0AviGwIEDNSXDYqllQgLUOpdul1gj1WWlkPJ9z28Nutyy7UtWOlqj
iz8amvAyw1BbUU4mJ5Y8AyvQEUG2cDeHjFr7214mQWS4J6CBFnbg0Up8fQHQ/jyE
fW9DhH1Qf1xGP9nJNMfZXcpBG7NZM7idoHM3lzKswsx0sR/IKxVAyBwya6c3Xzjc
bLQynjYCIpPdk5Khflx0yGn/yu/bYkWYcyR6ZGCovQpiPQOvM4hSk72bXhYVCOT6
Opv0t+8sduVEqlzG3AhXQO4Gj2DADis2f+iag5F7SVDpYxcnE6S2lJoNH4O38rvE
6gS79jLm/1uJjg5/UaBgSdcouvzYuJS3bo0XuSUwZUVQHNxB6SG2T1kCA12mq+EX
KdaIHklzNNECI9IpGBMyIlYEg1DzGRKamWUySib/PPvECPioUs1HvhuaWwGcbrxp
XnSke/4/qzXFGzHbRUIk8+AQeOy8gneGrVoA3BqCLRJ/+QvoZkXON9b68XiwfHY5
R/2Ns0M9YduOCxy8Nxc2gHRZwltJv3FYGDPt+Kh5YnPQqrBdlrR0fu9P4EazZrdA
MldNN0q8VJvCU3lANMuaK/iR5fLtrclE7tlHCc7Cim77luLeAGEjeXTlMbMPKHU7
GEgWXRhBTDJ/ufKgyn8d8rcupQCZRA18xinxtoxqRY/hd2dGD4TMSV13/1MElXBU
c2NZ3Hv3EJbOaxgSuxM43mL0YyXUi8mnytFIecTFe7rPtLb3qPsYHipw/szn9qcX
zTG7UXn2e0+GrCQBv/cfyVH5r17qASSbletDO0ZVuE/TbgGGRNKEjWb6fjPLdkN4
EaM1kpi0nQMCJYzDysyCm/tehYI5OzsvchgYS4THOOv7YArgJGz2MGJ3Ep4kYalq
caJhi7jjT+XZZfBbDLoW1BJVDWNVbut6u+omUPV/uBxc7dD5slj7F2acUXgkmyi/
2xdd3dQVXZfcAN+NdJQvdqy703VTPciYT1AE5rkzqm0uhqRutPquX5OmA/x3Rawa
WKaXUyjHRh3qlse/XWK4la7Kbqsjv0tRZ+Fbno2kn8AqD5YMOkHtCisz6NCMcFVc
cXwO+W5nG5gBH/NBgTpcp2OldPD+mDwYeGA1vV7PaE09caQE9PDoUfkWXERiI4d0
qWlsezKD31IITYMjF1x7T5z5IZ1gwuyV/l32Rob1iKP1KaCmSRqJBlqEHsZ3Qd6W
OKNlDxdIMmdE6rTnML9BOjgCrP71A/AI88i0wJDaO7TVDcZgEKDO5cV21SRWEXD5
8W2DEnJoxfQJSymXpd0NyYR9GSd3M3ivgfDMHLIz8049TtnSoUEzlLJTHIisSkSe
dRPfAJuUXLj6rExBq9LvMy3C0lLU3dK4KCQJuIiIqw3jvi8ub+YAuy1KWeEq+adg
wJPalvrntpbn1H2MFENq4eH59rk7tUHfb7sKRJkCbqBsXHIa+QCDkOmPc6ibNf1K
u7FYcIJZErrne5msuWth8n0TkWS4duFb1vVwtGCp0i64qr9NH1/b9hrnDZkR2sog
NOrdOzg/nR93WJ7wyi5Aj56/fYkQTfF5GfvLlAkEkAWzv9/vzkpfbT4ElchFjhPW
iyGZOqbYGBA/Z1LqJHvvf47tLzJquSm5IkFDF8yvCxKnFgEXIRtcBV9V6EcJpS6M
eG/wZjDihqN7FfJICSG57Tv23Uing7uf6vI7Eb3rGOGaI60ZG6eRAUFJ08Fx8Dz+
EAB/CEzTHnIqv2xhN5DLB23xv+GyJEOj0AgIGU20M8zUtZXPZt66djXvBgXKFh84
9QkN5045byz+1r1eEqj6oehZdvUbpXltkHxIW/N5WbxU0oNI9mnnt295m6zCUGGZ
6ZpLYo4AyZ7JnXLkJvKnvV97tDXwpsy433ywZJm4safdpoyZFXfmQZ70V61Z9Zwc
HzA0E46ClsVHvgdQLSGNxFsQwrfPDY1nBKrlNaodmRK427mXVgyu9V7Jno4RqMDa
KxLC3XUQIjwz7KoBzoCJ9OKfImQfsPMz423icmts3nZRnUX88NC6jcSKQ501kVre
jkmY5M/fk6PmLaCgBj0bWxubjDo4Pk8T/yLev086PWUAr4JjwvKNkvakydzhT4KU
jdB1JpA0W/cJIQQPn+8uufBWu262nmek0TCrFWjct0tVZQeXLEkbbkTOWMMYdkCn
EzrZ+67R6MEaHjQ99NXDTm7mqgIdtWsBpCBvoYsDj8yRdYRFNRLevZiP3abKU2ug
T4GZ0Mx79EKQagQ5lJVI2kOtYfWsqVi+oNqrhZFK7MDJr57kKFlALmU5KCqY37Ip
Mo/DJsY3Lg5IjGpTQIBWVV3HekgunqGzzuMu7qPIx4Jn8qgLW/YSDRiYZ1dTAyQe
dnCXmZfkWuclnf2dHfcmv85Foxr9+JqRGU30OJmm461fTYkblB866oYvO4EN+ezE
IyGLC973nJEiPH6g/KNzIHy6hlIGZbOuxlNyd35iim1GbFXrAXwsnIcwYgtLWrU9
nROo2fX91vrNII4luE1yGOT2Sr944rzATPZCyq8ZeH/RTSAMXYHQ2kz1XIj8e5RP
u80Vhxtchk6SKFnxI5EHLJ4/QBQ+Qxz6uY62onh/B4qZMZn1LDWk0Qe63GKF3ieN
7FbuJwTyJfiRVBoHn+LNjb6T1w/KQXuM5p9ZKItiY9QSrY5Ztkvfxbr8pXhIr+eT
y3o/cY2JmaoCEA9BTMUev8u4w+PLNsZBFaHXTB+ugr/pWflENJiUO2wyWAn3gQdA
yYZed/T+EHVr7oszzy5FSX1AQLAfQUcpEc44g10LikfxdcDCGn1uXBL3MpErq04x
SgDjxRv6MR2iqOn6O+eW5XgcJqbFFK7kg8lRBTZa4Kek9e8FWQYP5z+S87IC03yk
+O7j/f6eVjGLV4+esCqrPam0X/2HMZFmOkJC1VdbB7s/+ZE+w4uIoVJIIBGmQelt
aTzuufy2tTjyo8uQcP8oY1PgKPtZ0BW/2rJhqSZv5KPNosE4pchFe6dkdJayR8vA
GZwWld5yozxvW/gLBHZdOFIRdHX5ZCJv8savvj7oi8/WCBJp/8AHSnNlXCzgAAr0
lq5Tk9ZDrvi1JjKpev4SvVMSZgevWP1kj8MWTjsiyrHnLhXJnPkGHbZCGUyrHcMd
JU/Wdx6ATv/p0uNMQwJQiXldO2NQGc1NJTypoyJ4qGwxX+Pen0OEBoOLsIT5XsWG
X+7iy8YUM0+DAF9bAF0A7wBReYYZgbXkQBr+ZwyMqxp6QGZlQNglYPt1K5Y2OJCD
vvJP5o5M4tvRkehuwqMzvA9oxoDzX5oVvxcdupMQ2KWPKQ9UCRWdP3+lRlXgvVEd
1E5APXYqonhTR30Mmg5F5uni4MobvnVCaWIC3Kwx785eaxQHZUruANSri8dx4Czf
qAWidaDw4bfdeU30rw/S8oEHppQ4PhdzCtYUkOHp+hk2OGMZ8jtJdbLCHjHGrvLV
nw0NVmpON3KH0cEbKvJyJdSn1CcKnFsZw1QuUEC9PhwceDT9FnllrBCR7QGW3hsN
NxXEeB+PQnMknoBcgHXaqVFWFyujLQcg43D51wJ0IKcFiBJso9QTSZg9SqouQJZV
zGJWpwhdPTqIv/E9DBbvkqeXsHcoX3rtJQyaD0oxTcdD4gDUfVkLzY3sy1vr92IW
6VI9hTxh50hoqRfY/lW6AXhqaFdRlv/PH6zpgpEg5deQwOcA1bhvm51uJGT+z6FB
b3TCPxWIRJ8ru9kSQZqyeAF9f1iseSg1Q/d3EejH3PXutsKQOaBaZWdrFqKIaapo
Llg5HiGiim8/9doy3niogGfHEJIqrngtf9A/79cNfDwGmWMQjUJm0q4uGefMmVUu
kusoy5ICKcmWx/hYBrc7qAaOj23Sw0zzN3IRRU9BhA6kKMm12EGOBNG4z8JPGyhq
SgH17u4vP3SOcN1zJe8MKWuX/Lx7W/xzgwhOplW35XzMEodKoeceh9eM55xuxL6m
VpK7Y14/EgJavWa12ABBLC4IFe7PXaipDltBaVQKWEkxJ1Kjod7H8s0he3FpxNrn
4MSbBsJQBR8Khw4q5xRia6DF6ZIJpZ250mlrcQuIdBsjnBAfcIe67SzQeCtY+k8T
B5vlCQjrZI4z8+7q4Bfw4eBMq8P0wzy23MjyE49QRnDOlDWFqiU+is3ddfdxLpc3
gfthBMtncY8Nosl7A6KwJD4iOKA3Eae06BUnbiYq6tYNHIOSjiUUMcD0vReLf5ri
LKjueWWfV3DL+iT9sExrFarvlx4j7o/Rx4PlWNCj9AxcgNFHzAWeN0qszu4PiDW0
9P7nUP8F5xOFUl/uDDOb/1DR0iFfoe/cTNYu9ZtUFjKi0poNeDM2JBYt2mKogZux
VQQS5tzHBUgELEqJXkGLPt65W8v9NIRrCpX+giaL1xDtQpOfuYwjMCEL14X/Us3V
kd0+YE1EdXIih/X/s9YbQVse3sPoKSr7OUNZhoTRQjHLb3UZTDQ587odZ9+/zWwr
vrtsFIYJhnkcVlg6ulKh2ndNzZCUak+TLjWxU1o2qy+5Z1X2Jrvz4qF3q9p5lHgF
t/nfZSObSRha6HnDJSJl0ZdAWxSzOpvJxdP6vqXdDXJcCV0jJeFJFWdc9dpACp1B
YEl4wR3LP+17iN5hGV7QLyGY8ppntcZENBZ5p2lUj3hH17FQ6VCA5ppbnuDmtwt6
fcr52LFONbPN07hC+pASyUBuy8upeXJZ2nQKuTJBoV0xouHy6fnQjt/fbX6C7WII
gGSaMD5LuAvETnCRJLNL+dILS8yZwSUi8cc7xaceXoA/mPODHyQoJTfgC9bQcZ9N
xZJT3+0CRh78RKot6zWbh3BmxzJPVQGr32aArQqPbz+2R1bvS676LdDc809Db+df
0w7cJJSEYscJncBjhunm21isvTl0SJ+X0a2hUL3PlaDustR6iLJosctU12+5v6oD
BT1miq68CHt6kSdMXMRJBOfQ+B5AivGPL7Y0xEq+17zFTLBdrIWUSXswNoEIcktW
hV6CsNwGEmVBZlcMLT2NOzO1ivqm3knCrBkF3luThNuMA8siNSyVlfbXJzDY9mOs
FZHVxiFPGxjhxZCaEZQVOSQyndFyUfjF6lelEdmnjtTiFaiwGPO7JM4hD3g2IDAX
8iAWqSr+YrmeS2EsKRx0hw5+/AQ3tiFbHP9RwgSZUuy5hOxZ976ZZX0CtPOxu86c
hHgVT4WNmwF3ieW9Sq4beuinARfscjw7Ek8ULxMoB30bTFJoqgRfSMSpOO46jQIi
rROplmPM0/EJ9rghmfvLENUVpAqyHjvYR9OpGJbSOtAsh3lJBqYq5NbnZCZ+NE4G
SpEPdS1JDYWFpvo6CK5bvqr+NwdSQOswqxaoLRkFjqaRyCk2DnlywqUHD7M9/Il/
yBNS7M7ou/0yJaGNQStv44M/4octBPX/xh/9fTegpOKVH/URhaUAZnEuUzA21Z7X
mB19kSFlB5Afw//bQ394+LBDdIN344wnbsEUJh34pu9l1U5g+EUH0+RdJj9XXzYl
/gr2BZhEyadDxFUSkYZHsXeZXMdjM1Dkpw/pdfZ3RYPrR6Pwx2n/7WT+fULLhWE0
IUJq5V2VyfZ/7xQX4OKSPN8P6SPN4IQd7DI3dLGvQFWL+L/xcVZPZU3VpyTi0FLH
IxdfHjf12Maz0z6OLwj/tzojJJAstwka6euutsF1qtp17+UenXL27tyuunpHS+zp
rHDZX52LuCtDrBV+0ojdueoj/IEDM/rVnSsQW5Xer+yjVAoMCwBb/DnrVdMu4jfp
yGBqYSfqlAvIDV41Ckm383PCaoSI0qsEv0QaczvroUK4smOUAQ5dCrbm6nr1ZdT7
VsQkSMxkWeYzEA803S4Sqhk2dmlue8A1oUNVSYY926DkdffAafSq8HVW2c0zkrSi
Cn74AtuPms4hnJ9JG9w1yPQiY7djcge54UVl027b1IByDsdz0Wl4j4Xwf3mq2TSZ
zmmZ+XpsNThHfusTPpvNOdT3mFEVF8eWZR/7IfkrRoFjb2OfjCKvW7+uMcq36o+c
sy5FnXagT1T8E66A6O6tjd4fTdQmwLyOIAKlOh2KoC9oFD4pS+jwtzmCO7wNKtu7
Hjbu53YQROII9OoIcsSjCQ4tJIgMQLPGYxZUGo8PiVbWCuyT+ArT/jDEW5EDw+Hk
+ht3fbflvSABb/Yv5ylGo+tbOB93miEq8R5uAWl1i+IQlTwWeGk6BRHMuDs3SLlS
xIVof8XYaNyqGy/7iMUgIk7EFU0+NIiMQnHPiSySshUZcZXJtUSXcdmWxIpT7c0X
/qGytwnXP5zFY0tB6LX4NZLVE2ek1Frd54yXCi44SMM0MknGltQvW+w2s7rWff+C
mYoiVXt6AO8eK0gkh/o1W9psQm/+Cv6UX9eV9ZiairGTh5jPst01QSsBpaaWCqqt
HIowlgiuVTFgaMM617KmVeeFOCK2XZ4A3QJYqm3vPErZN1qB5ixRqY+rkrhPw7G8
B9/W+YJbNKQZ8FYS6BksBeagfNW4q2Rnt/XaxzjOYLbHS9VDIITCeuF68sRNr7vS
NZ6p2/SK5FtVbJbcjyjmemdiq3Ewd4hdaMbKHhOZXkbC/zzsHsrG7NsgGJyqdiQD
Ka+WOKPZ1RgxcTOBy+e1L15UqluCwfN/Gz9jtL5TFfOtPtf61OgsBKjJyvDqqJpd
SPxxepxKCLXljx1YakKxT5BEUreuwb2OYpnLai7OHIT22NwV4LBH+HR8gOH9eCZO
VPLCfcPn2xuwPmXi98uMxtf1DDeLFHyqJuNE3eI3gV+/3pGAVdRXHr81FTn14Kkw
u6dliyaCCwH+XNuYbxH6RFyO5NL2CmipooqquNUvz6ZYXuE6AbVDx4DyLu46PKnp
QJUgn+3JoypSRV18/MrdXB4k6NEIshsnuogTcd5U7SSq0CT1K0+vulBURaZoRZHa
Us+ib4nepAcXWyXqkxGQaOOJl8U65YITYoC0LEcmt/Zp+sDruttGl1ncykdGLlZd
jcrCo0xssUWhWmJVtM3r5koHTb0OzejYH/oVbfECukcw4VJZcEK/DIpWyyiiJCd1
orMy/r7f7JcGxLzbBEUEALDE7CHdNQWUqhw5GWx43ZmnvM08D/1CeF9jD/B/NqFv
B3/vWDfUNZqso/Zto2VhsMJSlc6oAdQ+ggW1zJvIh5YTDMmnzB2HsfyZhXSwGOTZ
jjBDkD/FlfyYy79/uZy1s8Sc6IrUbQSa1s3k3vqyjI7ATZSYrZxGDquxTxQKqHlU
yXMgK7gyh5Yx6Xa1e1Uk2T2Nhu5wczf1P6a7GDRORZzs/x7XnKtmN9iwPtDqrkEq
uXolBUSAASmn46HvjQgSBEeIe/yBQhgbx3SDkLtP6QGOvRDrSBJT0DnuRLfza2WW
ndp2oaND3ZBuogebpBhf/CoWtgrTRiesKX8l5dj5QpHFQ3KgSLVnEFl3gXfma36t
7EkZGTdD39HNa9hWDrBzsOJqDvJVx0Iv5WXQDfggGoK+aYBMqZmg84WY09af/h2k
XVtG7RTPLL3nWOfD7Vrj24DbwgXlFbEtDEArM08qH+4eWDJDBDZzIXZKm9sHhYnA
HIq0QoYmazuxkzKzzud0YDYnhaWko/6BxDTPVQAHkirXpF8ou9VKWl+hwFOw6tf3
vMpSwj0nXjUKkS6OS0dpXWmTzzGAIblNx+13A+KT5OZgGUnCwXIWDisP6s/D6I8f
6xaF4yGTK2kyf1E6Bxxt7TXokHCcYJFbM1CcONRJF+aXYYPksU7riOrkcuMFKsES
wMukBFQwPGbiLJFCQ6LLeqT33zE0CBkcfFf8SERJnjjXr1GNAPHoMxlcAQjyt6Hq
VU6M0tDLqwWzCNl9q0pspndpxVrp2N4PhoQQkf1UMBwrjANKCwAMU+OhXBW4zNRG
sybOEUuIXHMxYh76xJOIrpdb5UATqlA6AqhOHmGq9J4xNMezkrU2Kv/NRIm9+sYb
zv210PQdqcg50oqeLkDW0pMAKZcTIXGXFPoDGPTbytdClBZJ6MbbeHlXnakPEE7K
1lhGkTkd0IuJVuEG8e/yXkzRCdhbYHN0MnmZgX3evc6RbtFPZu4XEBL95aFEx5ug
W/m9k3QOjgTRiibHvu9d956uMHICwTso4FIysOBlhcr+e+r3vUhsRbM0u2ifXdWc
cTHSz01+1MsNkTykUkjfrgwYYdd3pAAMLFWayQjzIT47oWakt4R63YkG11qA4w+k
8e+WdPypGlHY/xhhrH5FgGfooBH6lknjAO43iqfMnpAH2IMx+PCAdmTv5nEligQC
O2FAUu+J2F6NrCAYQUb2pYVY8f9iQxghXkU0TWAxb0K5bmQBK5hMomPvLxBwy5Dd
Vqy3N430d6Uxl1qPl24oRr7iiq1zvez5EusCvA46tZJBPxF56mmUeDUpBwCsnRUO
Pd7K6prHi08KhYEcFusRTQh7FvDu+cYCPkuLtQcd/eqK4RXMExYPuNp4fw2/rwd8
P75L02q9PKXS/LgoecHLY3N693DZvDeAguOuCsLn1rMZlp1m+7BXfwwm104CaewP
ojYF5nDujFkFf0BYOqSrclgt4JrJTL2rOfg17UFKHoXJNqhJhbXPuuqTioPIEeZZ
3gentSd+qWK2CPmEqLgDRXkWPVgw79Tlgt/NRlzMAwXi0Gl9v3EXP2vzVc8Ja6CL
L99Da42iEUn2SLsYbH0s4/IDXML7mhcbAS1kffCacw9jHt0cv1eyrb3Xc0yfF3B5
dnXnMeJJdaqWTadZBP5EQgdQrRcEUqUmEYVzR7Gq2hBETJe0xIahtkuLHblH451a
GWi2ME7M140TNECtWEI1fQY02qq1wKnyV1r5/dtjUoIz76jA1u0uQSVdECFYSkFW
PASZe9V+J76InZpbmg3P+FS1holNwf2y3zTuqqkIG6PrEnQzVs0duL9UQ9zhvvb6
JH+aMmpp+fF1qHYRKuSldZJlWmHdT7+ZCFk96nJZaXp7gepEvouZTiu1r0DqdYdY
4rTF1EvL/QHT+Y+/t9Fgt94EV6GE3+bieWOQfpxw17+J2oeo+aSwYa4Yms7qRg59
aggWTFUZApYrHDrDyblseJQBXjeIn4tLIaAeTHiIML6rY2mlvw17l7rGAiZw0NwZ
7+9RimlHFOzwMCGzuu122/MCOHQ6sKSTctaTYBQH+jkWBcaZ0MyzjltZqaHkRk7b
01wxi3cHvbuHQpsOv4HFrMaPZZyAOCY20QwBoBQ/VEUwwStE2FaYteGgBvxLsIev
Bd98QVCCicrwFTkIb8vsxmrUjMzNF188ARk79qpRMS5jQjouzVfD7GB58OIVuW7F
uAPgqDyXgH/hPbn21LtQmhERKQVjsJWOoR0bRFwfP48uNTsWaWr3uhCgMGAiLiH3
Y3M2XC5FkXirKV3ByNdxOMuijGYV6Rv1jfjiHxQd3vkjG+4gBY5PAR2hhW4bhAta
wPUs4NIfWVyb55GXRtaCflVjyciJQO9AMOmwr5DbgV4+hlj8C/y3ad61RZ7TH28j
cMxY/rUV6M3eVLEMg9cH1JPOnoxOJVk1rlxaz0BhXAxy2ZlDmL0oC8VxTUsUHTXw
O1znCwZtyAFa3mKndXKFVPcoEp3HF6NqEXlEEeVSRWW/q0xN2kmCDKsYTlB4Ai4a
RN4WSmcViQc8SDcuyfkZeNeUTFcSkPh6Fii2sX7yboprbmSTQmJPREHJJkYbAAbk
inH7y2kJG0UP9UJQuZSRIefMcq0VURQ/472ZyLKT6R3UhUEQYHlxX3aALoR1spj5
L1s0XKuKkrRiXnrn3xTutyIXEPFiLIRWqlX92jbB9tyYU/F2yG4aS6CHZd+nActH
FYgtPHSd0iuNaH7RHGi5tQT1niVomuB8lgYyNpT22nNXnyfuEOOzqRc2nDYmPS3v
VpPx3vlTGvt1bEeko0lLYPbeSl/C+8ddSSGa2nmePTi8SKMVzH0EQ5ZWXqffDkow
QCHlXP50HJDpp2HzZFhdKBXiFui/Zu6zkTqxdA5HjzoG59zVkjDQxF+JFj+wLrNZ
8aN86UyzpOCIwgVfhO1AUvfdUlENZXL7YXJrpeo+QGU8OeDUY3mar3f7afTnWm+D
nUh+uTTuwDNCcyVLP1N3vOXYCh68DpGvSSbKfwTWSE8Y6KFO8ViJ7knw/HXAdQQP
XrP0OyTJ+96+IyMLEYtnPxHxeaJg438JIPkz/FAFGF4aUaWdPjM8+RUQK6AeqdSe
K2uy+sjnqHXjn0UqbD1aATTObOVp9IRU72eYxu1rwWWiQO53QwPc7BHiXcaWLxdw
JnPw0PLwa5B82U4NcnKx4hqOT5kQLe7La+/Jz+oeI052qlHqbUoUxSwDakdUx8TT
PQTuFX+8y/WbxfSCrbP227op/ivPywiEhhvgZEYMvwRjoc9vZsFRoS0u+jHC7orZ
3NWFhYgYGYB8Hfb7X1rRpkO5XMGGZSLV92/K3p2a54v0BTV1b3azoMQkbSafWX2e
ZXiuzq+U7pX22xxmZiGMZP87y6KQJyEzhR0TM6rZnO6CZ/XXTdHIp5msF8J1OeGv
koKyV+GL+Byb6Je15PddSsw7WLWMz3TcRFyRWYHscDd4WXsMblUpd72DH+rQwDZZ
i2Hbm3G4V2sSuncdxtQtE+bpjbPJ5s7rdXQPr/1mVi8p3Dd2EGAxR+rPrqnd63tw
L/DgEbzkBp6iFhfGvHCmemIsX6yuECHrL1TzBX2RyM0oCUgJAtaYp4sGWAhV1Uy6
ilkIUo0beORZoOtY3+ZbAKLZ0zgocUtDJz59LJxfZFTHHcZqk6pnuxvA4JJHS00H
v9nNvps/pQCWL9GZ9ViUBny1aABv7YQNiiwMKFFZsr7Ge536AdpjRpkY3rT4srwe
pKKOKWmeaI6W/5SDrQO8hRplif+eo78EgNbBD/dAz5INSQzZGTEaWBr5MKbypFax
e8ZPV/8gCdTcim2KfrdHO8Tw0ams1nN1NsL4M/8q9sMPVgo8rjCNXFzSRTrjPln0
Sftvz943a7Vz3/BqoTAIY7x5NY3idPwL1iN/wpWDWl8hSzSOVKmxQre+XthtJoK8
FYwuxyPi745BOsE9+zHZngVbWBDIx+Kds6v+1jgqt5nvzGK/YPO71P6WqhuMpjz9
uFg8rxBa6l7zrJ08IT2hP8YlZ7m9D+HA/ywoErwe9WZzlUHo+nGgh0UpGdxyOihQ
cawqV/vYfFyHZKaHiKj86vQcehQHKPqWjHiudGbum8Y5zgSi6XL6rWx1/LKkYB3h
JVlvgnNmwnSUp51axu2+YU/esqMOoXwQO+PN8s/MBuZltN4OlaCKUBRRjL+LURkz
K5S70WdSNqG85tiEge8n3ow7Ns+Y6iQ541B3ztj/QAazcu85z7SipzU2ehUImNqe
5apM/DTMtunpntoR5aWDJMLxQAR3cMfUT1LaSMaRmOtdxJWBalo25F3ofgYG2vmn
DKpa8eQaX0HXWKdS3kN+3Q55nc5u0n2hJ0h7tlTIO/psEmxMpe7hLO3uxxCR4EUp
2tZZoAunAP6AXyPG6IyLEQrWKVe/+SzFSi4lfAqFzT2P7feIVYRf5UCZk6qYYZTc
Ay1NDTUD8dv2Vq1C6SpEuZThQSpuvzVtn8t1W55tE+mpXCcIgrZos3fpsCnwsPBe
3wsXRjxPeYH+CDr6HPnlU6c/rTHKGIsiUDNALOVLJSmyYc27+lGDT5c13oe5VxRW
VXM401rLVXsnqDcSEmzxYyjuHOJrXSLYvdkC+MxQsgAoJFmNokD9V4t1eD8sqy3K
vCpP2jPS3RblElCmvdcsbcSBIsV2diaYWIJelgA6/Dq98E8P572m1QYBWKZTIvhi
2PW2nfzzqXzNQaK7jIkk1RDdzt9shzpG60xWuvDczlc/BchSIwlpD2q6XzL/rBHo
yaa3V3EwxgjCYZ9RijIWOvgiVWPos2hkKzINPvXdW0w4O7sZaG4M97m5O4yJMqG9
ohsoHuxYRt6Ug2jZ48o8x3UT7vxqzo6bKGbmK2MLhHjn5r2SDU3AYlo8aeoX945s
mDOJNKdEH3bAuEStP898VeDIGVyt7gU5tdgoPZkVQT89uvZZYulYODWNg0Tnj2oN
AfvELRNTg8VYehyvln0UA6SX7kqCG3+FUwGe2YaJho2W0+KNLI/zZFuyOmgbxXx/
yYaQFCAuQjxi9jzbV3EjT+fVi9aAJuVZlCaL6pK0pQZ/Yg0R2RMizu9xyhrWasyU
npXtlCxQIx1S48m6doVYSoLVAKcqUPKjF4q6Ci0sIkyRzjnZ1PS9CdxZG1Qxlrez
UBtctEtB2NVhbExNrIXsHqI/k/549vLv155vqwBfawX0MUtW3KPpyyuVCEiTk260
DQ17zOpcT/GuQMkxoOP1aJU+pBAD3JxeVP52SfL7+T+6Fk8h+B0v5/YPwKVnZrrP
wpVaB3y+VlcIGvbdOn2os43h/GxrPXc/Ry2pqY5nGnqVGahC+zyoDf1ziNFUEs6I
LuCqXJAlEw6vU1VR7/p2qAPJbpUF+Y0VPUWi4A4m9fgGHW2TUrKjsHDNcPoVcEZ+
OsY9a0SNrHC0NLExucxQKcFB4uSKoWJml+zYkOtV5dBgv5SZmfOzH7h+p+1ZDOg1
lx0ne6zLP4+bzAF+uKyX+J3Oim6wWCJq+gLbxC2XYKoS0reMZzqGTWOwIWSQbPRM
frrIAdgG+fhZgB0BmTDbgUw0e9b0ey7ys8Y1IX1WVPZcS92lKXlcnygVUchrB55c
W4p8ppZ9xCFzs18vtL35ORWcSVmIpj4WsWKTQbd/EOFJLDzFKx5JgkHB4HBcyHnU
r4hiFOfD1MEDoqvFHgJxi6h4R7e2ELNjxMgSYJA9UtbCjre7dK07AWiSVYZYGK/5
+L0YLwSc4Zvu2nJlCFtCTvBFs1ra0CPsM5/1coJhR1xFLomuXNWunIWW1P7WmJbp
J9szg2SVrJmfE3VpPbgfyr/mdO6zWeAKw/faFiOuKZ/XKRjMh4clSFfO5qVNsX5o
tkhdk3KZmYnzT/+9bDh5LZT/zGonETvj9ynKRUqMV6Jn6UqwrRqmer2bV/xJr84R
O91Vc3AnnGfZjAdgjOyTPReHhZDIik0O2C/FK5ZVGIgddGTwum8U/vVg8/Wb6WbP
loZjCvqsG634ppO6XDCR4SA3swPEh2keVLirCFYGkCyulrQp4TiJV1rxENFJFMXa
3gpb/wkq57ekNK1eSFu97fJNdPGVXCfPnyJieIJeg4ASLJ/fndmlUYc7WKvyaV7Q
ZJAvgmT0iPLF/+B5JkRaoJx15aJJX8J46jOJYIu8zu0E/uVI9MKO3SDTWrtwFIdj
2XKTN0++fODrhb2j7PgvSdHrS3bMvEgtVJRsZhexR5ptOOjj/JP81Z+xJk3B6nCO
MvO9vfjTAh2h+tNFCptq5ZCrDYET5WfQFO7RSovtzaubL3W8MbRr1UdW/3dbCvTK
RLjFwB/VYv/5y/8cD+9Bt3JaC8jHlsRVfNLXlJRUdxCGfHaCAbtlSl5pY8Y14zU6
FycBNdGb2XXrlrHGGHmARc7wbtnM4NPtEx2Uif2YZtkldeaFiE/IrVx8BUlnbmNz
m+OFuZodFXG6W1Bz/ZonzZwVmpRFWESDuzNuxhyWFC3d8z3ZkxEaUnHLlo50zCEP
5An+mwj7EXnZqmvJnz7wX0LytGpsruL2nygM3vTr+V3+1dKx99fL5sYPzK+HsdEz
RG2bkY0yEhAo7ry19RLHzNCzKytmY71Jwcv9BYE1z4BoZij9oxzhB/NCUgAJ7Gmw
noh0yr+kbs/eIF+qDUmM+LdZEpEMh+K2SSopmmuhIZNuRkYdVjnIR0jvyAyEkNrX
iLFFSqKanx3Gih9YzamUNDaWhtnuLGtCgu0iF8SIJegqfHCujlniYNrT5SfDt6am
VW50pZzdkAThpMjw90pMW70PatkYoCzoDTqPvyxfQ1Opy8L8X94Hg92GPtsHC78+
6iV1/YZHUUVjy7Ks/j1ArvG1F9b8cYrtN2Mfa+kA3ui75MLiDVvTDcdN1n+/OuiG
nw4NXuwixvMW/vPu+YWo3kCEEkQyLTbcX4FTytHKx1gtOgTLNMzrKNr9c/Ezszch
pap90ro8cD5TY8j2Wu4k7Qd2hV6B1Mh7xnvX2mP0YVgpEUrgykySmvaj592FeHFO
UesiyBS4Z6s6+eKserSnOTlxe6BUWAhZNX2N5tmUzyc5tNnlHVjbG1FbqqPEfqGR
5FX0mJJihmw2wnNeG3QUPlq9kzi42X9HwgV1Ig3Czef/fYWt25k4d0ifSvI4MyW/
OqGyaNsffa/UyBz93vJlxDsDCDSeCUmcs5E4xxtYAz4XUvpNTvdH1sYVTkfZPtZ7
bC18flXXJlPW5A7YJf6mqkd+Vo79KRag9/47dGv7gTizq9W8RnJTwNc0mqnxpGB3
6YFW91TuA+RAQPKlEAl2n2VlBQNnVYxPEjLNprUw7ESodAiykdIHOyf9vgzxMV2Y
jODaH6uc7cn/adVFdUprMiHt2U5LwyTezYFJv4A8JZa4BBREoPYrbXV/1QDygrT3
uURwhMwvgEfYk0WsDDrBcr4uRBdCLeraeicaxRHO55tgcb9eslw7q8BZp0jT1Wo2
kmg3CbGf/R7arU30iIvJS9p/wK1pXb2ZKRqJ3SoActlTLCne3HJf10yw0PFZhgXv
zn8OB4Z9wBK20PREdxliOLTN98ifszH9svhHuS0hG+j6M4ebgU5/p6d6SGX93NPo
jbb/m9XGVcgE13Mo+ROfhL+lBxw2vzArehUasUgasgz6hGCDbUyOA4SE5nYYSUFW
zh+jyKni3H045EZZ1FDcf89xzBf8k22Y9c0fb6bdZYBBYLtkMBWOS4tRlEoB72o2
i+ynSYyGizKJej2H8SVFTSMjKJ8/NoBkPLcXA1AB5PKaJTo2hJVL8LAHa6wmjIZV
DWthPJbAqimdPUVkbrzHt4OfQZ/iXV4X1bCctbPFQzM00h5eANwD9VNC/51Lm1bL
jKyesMoxhfJTlYAa0HbgWHQBnNjov5Y/2h1hMG9J7PAI/U+QMlFZdEZEmqI4QDhm
YCookZFrTIZRwGDdRHVJSLbNgLv4OldJGoiJJQ9I6wK/Bx9ylE2hsq7DIkUM92Nb
emhZbiA36FuIDQV4Eo0NSoJuENSTenjalbzKBXk2Lxh0bPMICWuj4aCWdXIGjLSl
cAQkevpX5vL2hb5BmasxKpbz0dy28V/Y28eMlhdJtaPMZ1Lfp0vAnS1czWABwZoN
rn7Lx8vDlRyiUPBcziXW9mbMcn9l2uPoIxnZTayL0sFInsPlrdCf6JhJyMMl9EWB
WXHg8fH1RbVwuh09YP5o2f9rVGmmUMVJn/zh3/cOm3Dk0QvgYLRTrHMJCTZIv2/P
MT4N6znve+Zrc2Kj8UUAD3Zx1Dt0gK1leeLWHgOUOSMlHbs7Vur3EF1p+0j4ZDSI
STvNjAQrCVTCGHhJ6+OicWIIFXBLEX8SCpzxsDqygqkn90KyPp50L1llndK+7WAG
+KQmqAzPsn48R5H/ioTF0MLr4r+z7omLsTGFqPL6TkoNbaqmJYCnAjRrPggN0ORl
arFUrq/JtA+TZBfXegNaQvxwR0MjJOvux3lLIKk6tsR7q20ku0xM24AoGzGPyLuv
ElK1RxrnSAAnmDMQOdw1+W89cDwg0+TNOEVM2eatLVS1InTWs4FrL/CdwM+CHW/7
28q/dtH8nv3aaA5Ru81O+3dniO5xrKaOybQhOxhAZTuGGzSo2fgJB96r97f74FPc
MQBZjkB5Zik7qcdJ6jRpHKcQ3mpQXXYpGVFd031EdKe3lKOURuDH1/FYKv1UU+0a
KM/3hGtxNnWQQTa15nmOA5MXoMoyJelnzVpQm52E/AdmbR4VI4l9W7sXDwJqhdAL
MjUJn4XXqNI/96Ngr7eAg0MvLI97a6YFMYblSrPp1dfAFz8SgpssnomGfY386tJl
vD0EbdYW+AsTLMoC/NNIn+rEsevTiF2Hq7O/I0DlXkfJ906bPQ8C9TSPDE0HpEkJ
7AnEQSpHrOxjIXp+VCh/vQ8ouZYUWy05Mbag9DGZyIqmq7tgmxp3W73jBz94pIwT
hesL/9Y3LNkYlVLqeAHEER8rgElyIZGvzXcnIKuIVdtBfRB6FDHRIerl+0G02Lbc
XGbhoye9q29ZSHTAI88/6nKJK/CtQs+13VRN7hndV3b+lCQYqsi7ITSAAGrBbMPG
JgcK9nMfn5RciSrFo+J4NIFer67l516sfxRNC/YNtkZpSOUmKfo+xYtIVwVpbs5O
4HYJDoq6xn/RHR40amXXRoAabDkqPCVrbWj5Z7agD/FRGQJQZRxAsDGaFpBcZ6Jl
mmAgIS6sXbaWafQTqObPJRFz2ai+49zq1Jfhwpw6NAn80hFf3mD3AM/6bSZaISvJ
7lDsEXdc5JiWSlKIxrXcV8lzGF3l8SB2MjQxkCoLCZ/nS0SPEZ/fdDCh+ARMY0TH
UFxaAEybdvKyN2VqYT4/CA+7+fikETIQUfLC7frB9wCOvT0si5f4wZ09CXh+m4Re
xgae6vSLAIhtLIA7Fh1cI0/GIcX72G6zLKge0MFHyScHNQPgiTdCtXFytC/GRIiK
Y1t3BU5oLjCzEHPluTVflJfC6rPTHKT0OjF1lDIOP25tlyutl49qxkAYx/u4rlVB
xi3RVnPyXRwz4WTkYfjpnC2Pmr9kk3HRANUnFbbk40IuuuViNBD22mr0vD2snAkk
c0SvXF1JmC5mojpxmRFNKK+FiBqONHoChjsG4NzGNmwTEd2smbaiCMswfOPl/AD/
81QvBf945G5SR5M6djLw9Q2ddwHo1Yw6PAOU3urChSbZbt2nMu3QuNPY+GghK5p1
HmkgYAclGmWmy4RcJ0wrKMvTx7phzG9mr46xkZ4y/Exh1Qkk79wtllJ+UaQ0wSSE
ZDRAQ3qxWq2CJcgcLjO+xUdTL+Hk+T9NbOvRAQR1wYtd9YOSRR3KO8NzKVh3saWA
dxURTkrPP4USwzbJmSiz888XlFBw+mUBc4NqIVVBNQrM1rKtl6LsF50mGp6OgHSy
5OQ2InzZXusBh2s+ZwOOmIJynCmDmdWEtaIlZn8FP4SJKM1pyS44YaaPEneH3Xth
8QA1Enz7wfasjSMtvLQJZ79cnMfHGxEkkc7t5sO4okPicP7nBgL5r7mrtQvdAez5
VxLlk7cOI0fM/leYDokfo3CyNpqNbXehu/suF1kR5YtNpWgaNaOD0pqjkD42n1lV
NknwxiENJm4U2ff4UlQTw7XC7z8aL+9NaQVWF/avjUghXfnIP9Z8OTbzlZwnhy1z
IFxDu4y/5WLVIccLuiAxEvoK9cXNp8I7FYh9a97i2m6brf8a4PcK5Mxyie1b+qKj
fqT7mC6jIKFfSJQe0gk5qwFDu+jZ2LbgGhtlXFe+CC5K5FCgaAJeHM0TmCZWQ/a3
OSWVWv7dRLVurAUndK0OBsvDQhwbo2QEFrWH0ghw0depFPYU67BMbGGH8I24tvWB
Htic+tReVJsfmSa8adzFue/p1Az11KYIL2yDt9WfSApmkMRi0K7V/VobKQC3SfTg
K6fs3HhHJAXkXskxaH/38VcGiwNxl4X7oxXBvUre75dfB3zSIErXt97Dkj2gr+Qy
eJCjZovMGEPClVe14K3kw2gzlfMVS8sloNsVm5+ZEPcF34nBhQKXL+EBdIlTzHiG
iXt71pDOUYxU8jGTmXE1X0KDw0Xrsq45KJJHnQFFLKRUY4Bvz9tn6ReX01BCsO9r
nTtGXF6iVQtMtWa9LiX64JokkokxxhFxT+OkGmUN0BP93akqEPmtWEXWShCnfPQG
l7MbkXCSFBApWs7sZSKgF0eE6NUqlecdziuqCug3SmsLMD+HvqXyhkCK6QFWK4RK
0zXkGKt1wjvNay81najMqmQmaao6gLdkUsC4Sr182AQnaCYvQKPS/AjAFewFCxMk
m38l9hBHdjq5s46ZyJDPmFITzZFJlbwDXn4vZWjt/DpQ5sF+g7ZZiZTBSbIwJXDr
M8aZ2juH6itoI4OLkII5AmfjCk7QLtt6O+Vq1FxovRmEczvv1NDomqIyvmcbTDY5
E0wWD84cYBt8EgTfkhrdxJtC/uvq6YR++b3gM/fxJgMVOo3z8PLO1btAihQZoTd4
fHdbLy4uHaYudyOmkTwb00I9PesSkFooGPJNdCZ7g+Wu4mCpQj4mKhXYnzdZlR+v
Mgerb8FpFyx01LhXy4ko+Koy2lBkDGa7WBTedGw89h+u7VPQ5x4mPqC4HTP1MFCP
aHHEzap2MfvVqMgSom/EkoEjgCLozoHqAwNCj1P5eg6X0Xo+A/S0J8OKAxIDCOhE
lipHN3+54GCgbByrrAILBydpAneRgGozvosA02v0bZxAVmOPZr58lEQLShzw1uNX
6hHGrVwhvVuf+D6ZPuCxD1WWTfHzXbgUTE92tKOSTs1gVRZoD4k4+KItv7Fgw/up
KdY9ay86nQtV2Q3hXNbylnAcXEI7s7u5IjvMD6aBs6tpR71lB0LwcDJy18rCelT2
wsmdiobXDA8NNYSJA6Zb8NLke3RcO92pGGVZz7Jo4OijaOiNbNVdQj6yyi+iLB1V
PoRBfuTRFphV/VLHL4K6+YSW46Q4qZB+bRjNcI0LOYzP/MA75pSYZLr6j4A47hCe
M5DFbc7kowFWjdT/6birChmuoXLYMEZ4cvM4Dd2EnlZ/2F23cadV6yLv9p6rKs2K
EG9fECjboTcjKGANIiFnaGNzbrU1Xo9D3Zoh3NPkIbqJdg+TXLh4quM2IDtmJTqO
ER2+E0kUzFW8oQOkOCgw0+0rXPnUdHDvtS17S2RmziPiTm4YhE03GR81zWmR5tUA
EZYe6Jlpg63yDhGiMLN+GWFsp5jmcGTaTKt5Wnqj+wXgmAMn5kpjPxSH4uC+v0aE
pKyR7z85QharmCK4Tgsc6chXL07h3+TE+UXDi2mHuNxBnTWXbCTlk+yp0y7ZDzhj
mqU0NoVqf9sNyWwBf7Dg3fOx9vjL5nUemjhg5+RH4mFGk5RgzZJmjE5I3ts4V2wM
0jrRr2T70wVSn6kVfj6t/7uLFHerVe4DoHQnlwXcYn+b/S5rrvWYXckQzpFYsjFf
QaBsEFuF7Tc9pvCc04p9QFrzqwiNW2RV/m/CEBIoAhiCE/mu+SBoyTRLamq3DYC1
/5/K+brtGNMO5BRGYsXZje9FNkxf+BMyz2I96aN7NN08FcAlvKqihzOXhHF4X/bV
MKpVK4GBErIAqB3C1aeoxPIyEFO8yN2LRYvr5tS9BdZV5NMUZcbXSVMMpGhlo0zt
YoLz440ARlqde7tDIudsduE3HYFvIOdBjcM1dtq2IoHqgd8zOrVadrg1yoI0pYhy
ha/CbW9eUvRtgcZFT6FcjYZCFrXCm/b23qPgbAdEkjjbtBXsgsZSQftKR7uTNRxx
6OpA+ISIxjw9gIdFIO1yqkJfz2/jJg4EaYANM/2XPcNaIajU7qMq9b0MQi24+5T/
TlYGK411PEraoxldrEAm3uNfOyIg1xNSv7mDq9QtLhhHXWGN5a2n/j9JGv0YDWoN
L4uuyKg6+jjjzPApU0ayyfGYvamBLjOAAF7xmApXry6RQSeq1Etvhq+Aov012lEW
xPNLj+V2qPzEP+7EA/+YR8iEvfXzMcXH02IQaL0+xWZ6OqAuToBNGouwh3V8/xm9
hU4nj7hI8cRkTDdDUcK8YWc5vNpppyvMe6QdJo0vfMXJsDeIQPyOnZ5DenVN5mAX
oqRnRCnVfaL4LvjHX4kgE616F5l3R4RSDQWYmCKHiyzcZSJda+Dcs1EQ4yyo41kj
RyY3R3RVpa/lis2HrZx5mLxx9NE+nuOMk/HQlTaWdXllZ8S1+9aZvH5t/UwYUlKG
KXNYDZuxEqn7xLt5c2SHY6CvF0gDlnaM3sQ4voPzzs5EUpxHbnZ8tQQfC5EnX5YT
x/9SZsOEq8XD834nHLNq16d6Gq0yKS6IGx9licXx6g9Y6DagxZ9Nq1CWNmPsNye8
nzMzpg9OerrwqDDUt3JYbQksn8Ee6ypfQXhm0YumzpL6gbzlT0ui3G0WwayVr8RP
Jlr8KlHAvC5rrbTX536qd2WEay4mwKgdxxuSjkZ6Z3NvGLPG9roCRLIsTW6LTTgZ
/1SJUR372YxjtkFiA3PVjT607tL1uNHWm8s7fv+q9hKDuwS8Z29Wx1+OkBkEhO5r
0ukIhWi9ifQBMtR58SQ91y1JyPVmVYmfydKNFgZ9iCoRgZglpcS3vi02XLErQfNi
vgD/PzC5w79zSjSgPJvJgyZ2j3n2RCfEfK6RWC/dNDb0jJ5Ft/3hkcqbXAk5CsKJ
IejAmAkAd4hKtd774EqJjq5Dt1zcmOubSFZJrGts9pjnXKWQBHVtnJb9vwvl1iug
I84LQYK7dKSQdJGbV3izCVxfWaxdrxwX7EpCa4Z7pGV2O0rleVRqgeVHnSjvO/2b
9UeoKonjPTl3OCLCffROWnjMb+uQRZuNos72iP0KiyV1Wb7PeOidTj16VHYiz8cZ
XV4LQS9tuGnQU9HV3dO2cAKYMknzNZt7IZrqgkRHqoJgyXFwsQQTUY9p5mQnjaMt
MElEuKwrwyEt90zm45ZRU71x2gSbZsLRldjk7ZTgfPt2Tf2kmYsl8mAqgIgu+fQm
iP7Xg09qQPVMABW/yM/qiVEd3aol0OqunMMBM2habVoXXGa13Wu0gFepEILAaTSs
2Am0mV5Hnw9IkJqB6KhSh6j63YgEBGuOAYw4yxiTQL7zzwuunWmqdUy4UmB57V/k
hueOkJibGaIxuo4w7wUlSHH0ICxqcaFibJ3/MR9zG39cQSnii1AG6c6TXVHRyf2S
R8LdGIwqi8hZrxGQz0YGXqIAq6BwXmA8mz6AsE814bOgk54EXHhGzLdVtnGCP7r5
iZ/FZ5RLjZcSdsNUJMuUnx9QAwyQZBsbG/oWbNL/6ba73EoDP9DgitI38axqqyBz
cWoqgZU6YViM8Ks53i7cASINRET8kU4tFIVnnqal9GfDbIDwGUPDtEol7bbNZfOV
3GbeG8+J7AhMqWtfPJRlTEM7a/H/LD/5N1tGfOuUjRqZdm5Y3XerrWVo/t4oEYSw
WKI9i7oG5o5X9+m54IAtlmrecpSZ/n0lZMSWllML6+P4HHjHYb+KFpxVxio1TI6U
41nv0ScbL1bnEDH5O8iNDK6Igx5Pq5unO2KG8NHdaz3ClGM6Aj2Gdi2qT+A+uWGO
DJ0XXPtU5rCqN6yjMUORVka/8Q48smcMUYEO2NenZIpZjYYErtGINR25OBTn0pwr
Oc5Ssqp8ZJZP/x/8Q7XkLTK/3Rwi3tSWd1SHd9BuZJi3LgLQWlYmtoH9Pa8IkIGt
MhKF+iGZx+dvopFsrF4i8yA9o41Qy2LKW4pj1h6mcIjQxxYGDtM5BqiU6vMbgox7
6uQf2RbfaADxF24wyQugz3aH4tmFW4xirAe5IqKvqdjeP6cgfCK4W6/ttmHOzWAk
pFjDeJ9wMMM7IbsYhvoDhrGjqU5YMRW6o1AIycWEMngJdTX40hEySIe6FQsROuZo
MFSstuTrkjyYcGqCUGozINQ6pkIEc89/lQJLmg2RADqbMixKVfjE3JJQWTguKqVk
i4/THghURjwgfPoS+JxDi3LUZMbhiG/6sOARckscjK6KEXYlOwWBGQk4uv13SNnQ
aG7WQgELXjYpQxgzXS1kjD1BVTFZQkJhI7bwng/mZpVzboadNqmfy1ng9+b2EZYw
vaP/8Gxr8mHFf8uem6m1+IlpfuKptPNWBqRjVfw9YkTwtsrxn14jIBqNV40OL1EE
`pragma protect end_protected
