��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^��,�~{�q�E��	YjpA������2o&�0���c�LڄX?�i��+�#��7J�n北�����J��kƧ�6���+{E�b��pڢ v�U��4��WL`d%�Zx�Һ�|�N2L�\����-�1s����#�+��l��"����1,h�'� ��a��I�k����^	w��G�Z��k(\H�9���# \����5AA�f��~o�ItMi������)Mn���e�4eӜ�^�����[)�F�0�?��~��w(-�f�sS��c��7����3��/��ֲm=o@=0�*QR��$�Ym*2�ծ>"�j��MZ�)є���8���'.��]����Ai��b$'�c�]7�a&���S���,�'1�O�U2�"�7�;@�医�.G��C^K�F]���_�3ϸsN���ј��`a3mWQ����UJ��|���9�~�4�<�>R����t�����wt޲�MV��D���z5}/�a���o`* ��ք�DSf0�z�y1z�d��Q�R&Z9����;��X)��׃ec���\�8S�XNP��.dʹ�R�p�t�X&�p�۝�M����W#aŧ�W����oG�+�ٵ '�.���G����z��A0���w������T��<����4XJ ��u��Z�ł0�f �i\~� t~A�C�XͲuBuӧg����s\��©q*YfJ�ϣ���r(��Ap)V�۲��jKMw��$*?^�|Ḃ�Z�%�]����ښj��p����+�h�ѵp�0��4OG-���3�Z���w�i�˚�+��z������wvҜ%.�������?$w�m���p^�3�Lv�@���<%��C����^��q"����U	l~]Q��z�\u�d���! ���Ϫ��I,����./E+�/���҆�k~�(W�k*l��ܤ�h͵;�w���[M���B'�<j^L��Baeo����t����RJ�;��R_�f�>`A�
h�0H�/1�_�S�����	@������Y�e�8�		b`���5�N^K"��Ub9�Ώ��@�� ��o�)AǣX�^6w�ԍ�[3l���KdG՝��o�<S[����?:-�V�Ӹ!ڛb��bּCY�$��ۋO
�Y�sL�TG �^sʨ���Q��D��i�9*l�\2 W>D��#V,.�+{'�<�(>��~ �t��e�A�y�6��9�pˊ�AM��9��ʚ��F�4�R�w���9���[q�� o�*D��n\M@'�4I��5}������~q��[�Ǒx�|��d�!�2��y�g���<��R�D��>F�Z�ٴ�I����o�Bt�/���R�c�#YN`��M΍'�Z���O��N���VԆ���q��>:�>��R�v�w+�l8:����8�)��^�
�N�vW���A<�˳c��$XU*��̅$�����8p�3ȭ�5$	��=T���9!�q����#����N��m������,�m�тG�}��豮,�r0�}T(@���c+k��Su(��W4��� :@�nJz|�w�	:>%;��n�}���)B�̆yR��A�!���Wz��*C%��� rZ��҂�!93��L�(ϸ��&o�;7�9jͶ�@�
�G��j	��$�e� H���ώz��"n��H�>��I&�hFLg�����C� ���~�5gZ����M\��&m�0��.T(�G	�㙀�yOD�~�c_���VŖ�Tcq�'۰�A%D2;�8�Y5� s�������Q�����)�xW&�%�JR��j�X��j����1"q���V3#�X���!��25&��8Z�φd�ͯq���ǜ�5�c�����Z��wwo��3]A�E�c�{C�+"����)	+��?@�w5��<-���G_����/4�o%%�����E(F�7H��>_���k��X�(sHiO!��'��8lS����턋�"t8�� ÞB+�u�}E�����y��H��*�d����0���n5��}YdT&��4������ڣ;,r�[iFw.�fJ�`��:4_�f��Y��T���~P]5����>�,��2�a���?��x����wI���:���e�z�]ff���;C��ֳ�����ϫ/M�!ܰH�ݤ�����h�g���+^:���[v��Ω�pl���\8}aD	����N&�����I�R!#�R[��� h:%v�_�qOo2w.�U
��RSZ�e%�N�G�G���|ǹB8MƋ�.؆�+Q�Vf)�n��=b�H��0��z)7(���+�\$��>@����<��齰�V5���'rnRZ�����?���\�� �[d&����[��J�xI�6��>v���/L��Jՙ���dT��L��!�K�	$���;��?,�P�T��?�-��7�m�rzD�P="[��@�#r��O���O  ]�NsB������U���̞�x����t;�zJI_R�@A��Rb��˝OO�Zk��w�\��e������S:�Sv4��A�w/u�8������WYz��B��Y����x3&���e�jn�e�`�%�"��ţO�o�h��ĥ�����[u��D�Y�!��A��ȫmY�q���^v�y�����o钉��Y
�~��Pt�a ������(
��c^�SV4��W�Ș�8<�T��m�W�_b���!��-P��?��{����m�r-�4�g�#_5-Iϛ_/&p��
����to�cN�Dq��'�d�QDb��	+n�Jn����ao�g�mZQ���iߦȏ��H,{����$��f�u�J��EY�rԒ��l�z\�(k�@�N�Z��sC�X������E-	��ə*{��Gd�'<RF
���_�$c������]MV��:Q`��җ�=慇M>5g�I<jٚ�V���tʺH�[���a��o^�8Q�%&���ڛm{~p�X#�)��T#m��σK^#G�����Oo����]�ф�C,�E��-�R���_�Q��iq��ۄ�>xٝ�Aq������F8g0|�������{�'l�9���������J���?�|s����J��>�t�c��D;K�c4�/��Ք�p�Le`eG$Q'R��0�X�Y����R��_�,٦髏�+Dj�A�I�^�t