// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:42 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mFb3mofvVeefrfW+0d+Tfg594nFreH3tTy6WJbpVSMPxVUHD55PCA+I62BxnkWq3
zucxt22Ct4iBNMlfDAYCFuH3qahERXW4CMsmbxbea/9isT3l+Ykk0AT53i9Sboq/
0Z5uUJ+xprr7Z1SnI5mgYAY+8GXw7/XWw2Du8YaDK+Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30272)
s44jVKi2xJxx3/IWmvItDZvpsdbU+rvErQmceAry/5yL4RvnempH5jVmDKQFPb8j
zU8ZIwgNYDVM3AZqycTgcv8epalmkwFDpmscr8Xh/zfa53n6yKBh//zhOKXzEkTZ
LbxspzxgP6mT1qQHO2HA0P2do5u1yZu6fd0kZQ4nTNE5pCfkzEg/HNOaEOmd7Bto
v9mfUHo7fkkwaNPJYOpJU5AwQ6QccyMTNREuuzg8a1sPvOxCHbqbEZxccClgdLB6
HsH1sph95wlKKC/Lqh33cOJ2yPycg3Bu41xj/FpRMzhFqV5eyCtbOrjRcAYnhnsH
eF5f89iDyzg0UxkOgZk6jt1ElGam2pz54MjrPSqH4/rGGC5R96uP4APhlWNtLw6i
av3CCRffJ69XevgoqODJLT8scPImxiLUT28Y/CsEhi/u7kWEHh33BJjZAmYFXrox
L43hNnaBaza1Krl9JM7BLtIvbigEsLJSNCIEhPvSdW+wd0MFkfarPTzyoL4jiTBY
+rE//GKMSuwOO/l6YP4jP9bBdRpDforUF6YtWKPm2s+7gyWw3IJWClnBgPM5s8ej
tgPA+T1eVVWSm/RWfJME2YlHOwUV572kvpLqaJcv45dwiDJsMKThyZzV0LnI6NmX
fKsrvFnILNXcI9dXweOXt1eW+fiMQT/lDv6Qnli+Sw8tInUS0mWqNVVxd4+iGVpM
7Clpt1EIvRgiRyMQHpayBcktna/S3Mh2ANKkVEY9alwNWCoiiW4kTmJa7adDhB3p
quNMyZFzKKEyloMRy1n/yxc6OClVqRyz1FkM9oM/WT+nkzJilRYBzshVGR2VFlG3
D6ih0mA9IW3LgoRZlbJqBu+xleH8dY9B9CSyuCmclN+HhfTsprx06J/GuMiVwGWC
DTgTnK4/oKsRtIZTzjfXjG+SCRUtZGGR3CdYh1jamVfxHEXE3HHrKmdvKQK/8vRS
nGdxhqaoKn/MWDXLS0DRCHZnhsTTJQCRyBirdSv0YcxhUhmxmrRHXTtfJnHWl4Fe
Wwn9vxPUPpApym1qi8f92EqTyV7aw+ey2acpBlcbYe005f0kOVk+8dNOLITzTVki
fBFh9nLH5ivPLxRYaHDlPolPOfrpMmML9ucZL+fjeNHduJfXswp4hn/KM6DoP+AM
1k8219wwStu84HLjH/b3cx1d5R3hWcQIH1JYA/NsFxtvP/IfepyuNQFwsumiT7hm
yAyKy+r7qvhc9DRC7ONXlX7LCvDe7L1Zhe22i9qJgzKk0kR+5PLyXitMAiTteTY+
uoAus7OnF7WQVTkU71lpgJ3+cC7GdaDhmOzo3cmrhjHuNOe4iHA0JLOxKmj0dcdd
0hG1Be5aZn5OYfUJJZhQ7xaupnnCEqdUZvNsLkCkI8POB5YjIRuu/DmREl8oRA98
mp29wlJmoK25/WM7ZpAXxDlAdv/hI7gLPUQ+Ge2gjLeelWPS7rK2EF+k1DuSvX2L
3KWe5+64dy59hRDz7bNNKCHzBFb6AGG57TdCLzFD8KB1xJ5rWskEg+sanmyI73cr
UmuF2kyZS20ezOXOdEXrgc/YCG36y4dmYIbtNipPJoyrSLpfRVOEguD0lyUCsEMg
FjE6bzWxjZJzqu3vm9RhdxViqOE9XhJxCO+CLS8sq04ud/Dxwe+wYI8Uwcb2Jzom
B8fZ0eF6RUYPhigjl6c8Z+I0/4ntKgeWQ+jlJw4ptiPQYW4y6SlWohSomDDc5Drj
zoB0gTeO97esQH4UeanwYCTTH81MVa7ZDauhntUn5SVxmWTw6zl3fldLqt1w56m5
39YsKCecyYJkrcbqj8IU8X/fijWM9LC9dcjqNJApLbj5frsguBVgpXvbBvWWlzDj
svfxhz7hDE08JFDK7Asp/+oLnrm+eLX4FEDfIJ4ecQ4hXnf5/7e7Yqyg58Y9Me77
oLDPynLhnVHekbsh5wiF2eii6ls+xDZtSFtVJ7dNVesLbnLsjiW8jaL3xikHkho+
Zg3A0ZWya0Tx/8+leSrOkqw/yyVpTbxyq9aVJmqQwFa+wrPixpZJlFa0FuMWDeDo
QgT3eGnhfAD5cceqXDdxCZZFoeC4ysKZL0Q92sw4EABB0azATYeie8VHvY4yq9JW
Pkpjwv+my7Fe79rGLQM/VkkQAWfYTRvrpq/0fUhrtBwMB8yOWnaVA954xAJ81Y/l
2vys14++BWU9hV2b86D3xUGtXrnr+UGvY9refmF9N8wPJfKCTvnnCy5wrB2+ZkhA
BtXb9/PuW2pV50lJHlyvxlvKr7x6eeszIM77X3Nag+2BJShWQDDyyb0UF2Hyxjta
El0iOLjqsaWTBJb8mgzrEa8U18r1nCueINTw4CDvoNx8I3Fko1hvuagoVeawTHiG
mk0ITHhfZOZQMzy+7Y/4LeL+REGpo0S4iL4kQTe20mnFmyeCmjsnYUT9Xp6sCpIA
caNZ/+5gLtLKbS5atoZvpblWqKZkyTaqh3RcjF+acSXtVQnXkFgjeHdwXGafUsIi
2QowwbZDa6kgbaBEMNSNWVId7Y0rCE7ZwFStApNcpGOgnRwyjDYx56RSFdQdOjTF
T0Lv8d0bDAMlEf/naWesi51QFLWIrx03yKuSnPHjk0+ppHxFC3+pd2fcgxkw+iKI
9u4dmUnBijACTbiesUzsWMVRo98Dxfd/Bt0t6MjV29GOnce8fuWEbAc+nsXBdEj4
O7L9JAHbaO34wIalaCSvvLaoDddfgUYBmN6LLGio1KVXShXtgKHK5y52gaISm7aZ
lZEo2Dz0GroS2AHOGpMBxoiCv+LFru9J7Zk5/w8tjuYGQO27tuot67XUkfgwsX20
Z4PYNDxDS4ijr77zt7GiRcbsJhRF07GRI8+RDYxYO4nTuaO2NJf9Fw4MSOxqcsSB
yqyxNFbIaRNUlsN0pYWXTnozWYe/aCUrnkMc71krrg79Rqz0AbI26/T0/uKfB7kt
wXgdbVINJT7UZN7FTibd6EmgnPM9AcBM8vruyNri3DeXTVSga2ONzwJkaEAuhqwX
7LJ3yMbv86J5eaqLAcZ9GloZRdzs7Y1xkdL9a+wPi4kMku1ajI61ek2Virag5K0K
Ta2O9ZatNtyCrg/DFqIQC+ME9a9NEfzElG2biUKbiX0H7ptnnVdJclwgUrv0yBe0
eLDffEdBnzCciiqFyQYi5mK3YRiSYMGhU1S4EPTGm5P4c6oJsVHMl2UVTDSZEPEU
x3XzjPF4hp4rSqrZx63A+WosXCoQgGDBB7NhRhl5xyy2Meg0jDNOxtGzrSFa7U9d
9xhAf6EAYqzFkUyTjFOzYbvwBB6wGJKtWUEmHpN0KClsio0wpiYgo7ASRlYbOllT
Zt1P210pKaAHLhIDxcXp9zPB5kVqG0Zm6uWRZqNGCLilzia6eh9YVTJ91cjfz4on
AsMpeX9TLEmDaC+HwQV43B4o37X2z2rrJJ9mcEAbmy/zl8w3aGgKz6m06LPe2set
Wq6JYJXnqk+mIZxVQm3OoLl+UTNWgUcHfN1UiIRAUP3Faho4HYIjQDONlWweI8pl
CgtxKuHJBQ8a2ASIvCnFM2HxQRbjTrz+qnnw1JKoXlP2ufQiYAJ6MMfeJ6uyfv4J
98DtzkZPza0Dn18/11Z068nIwftjzkVX1IIJNoqMCo2k+VO4kwU5JoDfk36DrLmL
re5tHsFPKTtX2/cAr67z+3LLfvC11jBrdvAfF88Y9F82zlDyZM1hZtsjvN8rJKjY
2RhmRr4a4kz98wJkGvs2JSIUn7BpUJaFxV28GGJpihB/wwvKfeA7kegkhW6cPsxd
QI50g7M5/DhD6ZUNDBpQwBiy61fEfSfWlaSEog6ejAPvX280rJq19v+VMqMFYnrT
l5c/2eh9L6Zun7vFVsfTF+A7gzO7Od28BhPfEdyiwuk3aJLdyT6Zx0r0mYc1dXL/
rP+BNF5P06lpJVcj3Mfnd5HcmhtjD8iKMk8bt8fmSRZVwHX1lHkYW4fnkBPrP9+3
dNz1lq4rtoTzjrbT8+2Vy1n63HgD7vgc2eBg9+CEmS6iUfxnZ1obA+bQbyZzJm5K
JtUg7n6cBNE1YLYgyp20tRkuS2c7Tzwl4L07cKU1MB3P8gM4M1BN6sUEsf12DA3T
O6M0DgMQKjD7cwH5AmjxBJ8qpsfAge5ciELCClzsehqNBCRS6TlUdP+HZdbD6Qs2
rxcHh2OjPMTWrpe5wHXeBABjQxmUqQDRom/gOgln61VhMcsrKYVk79VpU/ts0LD0
vIAFj6l48Y7CRzBCgtI+QElEE1lo1Ppo7Ro1Fk226Sa59wZla5dRcV4Ma9DE1HZO
YC88dcT0C5rekBhk6utP9lKW78L0WMTuupugDaOErBcRKeRUMulmNCxYRojcsZ28
om17SF2S+kM+zeaVpUt1QrV+jtFEAjc2sZFyl+WZcAHYHIcb+QGnx/IlD+tLJVK3
1KDefEbqjwHfNdaH47Rj+ITAmUr1/wRPcBLtK5Y1bSLfFvtolP0kZdqNWUAMwciy
OVdCPHOlpZ4WGKh7K+VHZR7fVOlTDJNnNCn+TJAfZ4C6ncjBMYlDHi3crpXpyABu
dnDMFjT1bfSiJv6jwZHTR73/aA9EsEz3V0krDyeWojmbk/Gc/bBbS9Bd8NY7jNsf
nrd9aUTMzgk9QF43CwSLZRdC7BROJ43SGgDi0RTEyROu8WUEUOJlFK2X9G0GhCey
2ZpEosQuXlPnZ3hz94DI9PFvOSd38P4LtU9TmqVXK8ulamatlYzPvyrS6+Vxze0u
iGzPA8fWWmbGdVwssBA/Z4xyAz0yClPmS0maQ+aO57InqlVsx8NNngW/I4PAQn4i
QPpx8ob34D6KNzL32OLhCL8cLgDo2y28KWoe7W8CCoNAsHkqhNr3Hcff9ovGDiPC
l6clkw3Mc/NncBRjfuBHaS14yllTNC6i+aOcDwVispe7QgGbZerjLRB4TWvdFWqD
3bNbPOKeixY5SSH6NUjebMZb5XVMt7kdZvGWB0f0o6QqtAZzC2Y4z4gmqD5faHtv
8yRbykvcGuJOKqXefwiNTB1+TkzMaPXzhPc4itDZrbvldYJQ6PttM9+tN+69Jk7T
0wL7RgAR2ZJc5JU0jGksDNfC9/kfb8px66PvZyLkOy0mMPRDrb6xbmafGNl8J/TK
iUYlTi7p5PhtzoA+mMeHUUfxKko1k2R5pEvcRJkusdb0pbdok/E/PZ/sGQDqojd8
ODY5gcKXmT4tX1ML+Fsinti7Daz5I4QAwqgl97QVAoEcT5XSkLoQ1KJRmz7C3iY0
Nwzv77hbaVguU0xCod73HePud635TxoRE97mataApHtKMubBlrv6Nj4vS/X+cwbu
1xJdAstqFuuzgUDsoqB4v4n0UK1LNve/SPRX6DCMBlGhnhm4kkuwdoOGwZyTzrmO
K1SYiRUx3UrXCw4ZXFqklL2TWdN5s0XixVmRv1bIWQ1roPCh9TQqlUNuC+oM2jSo
e0d4VDTkhciPC4/V7HRqO0MXZU+qqcGyCbES2KgXusE7ugK9YQJzE3QOIYD2ssUC
X25uz//OqFKMyzQ1GwrmLhaDWrNv3gbZBx29Q68I7wOHRDZ6Qc4wvcO/yE0omZbv
0uJxGkXBcf0ttZcAq1dYe/smaYH0fTBTNkUfi2iL/5PLnMqdf+5zcvZaKmA1XBA2
9q9X74lveZPMGtjvwXrVIzwv3QBFQZolJgLiVdjNkN/ehaJyE2cH8crxL0iIhtaU
/mxZUWR5kIaCcS4BVZ975Teq6bkYJMdnlgOiLIDrfvPIX2wbn8ibFcfD5gBonlgo
7rjSvZYvupR8baMe+i+S3CLRSjlnPHe0BqdLFT4wRdv4oyWmP5EMdHBU3d9CAuKu
7G6OdTECqyN/N49HtYXgTIwe8116fizSxhx9eb0CzekKmLTCLz7OutXrSe2JuQo9
nf+4uM3LWFdqyQ5WDsE9sAEODvBVF0iJR89dg5UmLMZlr4/IMw5Zn+BxFy+BfxMH
tHNfNhGW1uKATb04EQL9aPkUUyMSQiC5HOvDh8vzQnA6OCai6aRoQVsDRbvaH0Z6
rmZ6J7AdMTObbCQFKbgbUhSdPZR2q8N6fFVv29q4enJCgvx95HNYmvXD8Ncbwdpa
rQZd9P1MMlM1U6d6hzL0DJcvtQXz2QNIxtzJeJBZUYeUkgVIhirbVMSR6fVvO/FO
PUiidQPODp9D6t2UzTHkiMB361bWMKBkdFqxJJY5cCI4JNm0NWfe1CWrGoh2xxth
SkTVYmj7hZp6xDq2jiwgHla/8j0bE+4tbyGg7t+Drws9CBd5MyPMr0ppXEHrAn0m
WboifEme/otjgECCuMtC7muivDmzuE5YkJxPKWXFDvKR/89LQGsMS6SOs5arckJJ
UU4R8ogvfRjtOSpTjP22C5o4PIUIZ5CkcfLtUfqTjdbjlM95ehat5Mf9uJoAygFP
SbaXViDZTKUP4PTYDM6ZH958n/TtL4OqUo5Y08J5PvGhdF5rPHn+Z9T8zEY9f6fv
gsTu2expTX+oaWHO7gvjB16p6hlhz4T6heChRwPfXphQVl3pYwq0PWIlE3zsKfgw
w6969TFDH8IiojffXjMteJWXXKA846c6ifEK51yC0UH79II4pZOO/S9y/r0SS4u1
nuzkzAASKYMNlaihY44XyDqM8l60kiJMHbvs5icOsi0B+Q682dfcVICxbBgIwpvp
TuJR2F7lp7aa08mkPQqEx5u7jMlGgJ2Oi7p8zwDXbPV2Zr2LQs594BferSu7jFrr
SPjDCFRpkkT5R7qYAAU9WlUh5gI1ukE93kOrfeqG26j6sFtmuWWdfqHQzJoLmZXV
6P6IXypD4tO3QeIuNk1ahCynXfvcgXIp/fMxvttCZTvSCFYlX6oFMUn5evoRWTzt
vG7MTDiafu4Sd7thDi07GcD7TB8Z4cmJQDtPL6lcHjBQF4sO2fPCjZwTv9wUF9I7
OIzNcvsRgQLmJnoB3wt9rGQ7V0i6DYUObWMcsTl+91Vv0Cl32azjg6jnGV8e15NT
yiW+MGYn6oE379qHrcjhz/KvF/OivkV5OdNw9wy7ITXL0hI7l8RPlsC5D5haIU4q
ZYpLhHX+m2B3Z0U+cMiaV3Roc90/4fJQAo3k/8bPzH0NSbx/ju/qHbyTLxs+iqtj
qyyv3ZiH8lYIDPIqIFUL1wy9E3NEOT7LDIC2EA0cNKkZ/vk52eReQz7rL5CmtOou
xAarSsOJSc65QBuIcGE72V2y3fmyt2rA3vxEN9O9zzac0fR3D4UgJyG78mtuJRM9
X2eB1ZB18QDMlvu77C2ZSzcKgPbteppFEkYR4tsG6tv7wL6FQm4OKoTA1e2PVHLS
LyG7dd2BqxVKfnhAXBXYfECYriicXm2a9G6X3Tt8UixcbLYzeNfMl6M6cvyRF4+C
uT0BBq0wEstUk1DUMcPzGMNdrUE0FCSdg7PP/f4EgpUJJMSeKX4r6HjytcGfKh28
qd5h7oTVuPhfrMaHzEotnawJP/UK0yBnFq4Mf7xCETmaP7vntycVcWWTvsHFvtLr
tECZWP5Cibn2Mlgye2ziKkMkp0ZHu3wcz1WoAlceqzfPP4BaeL8V7RJ7dWb5J5lF
qxbVMlI1hq4mnvi3OH4aygQVYs0tbZyZN/1F2iOGY9Bk4x2RdWxhUsddBFYvGS/a
txyKB3NfIYrq5vAO8vQ07iw62tNfiFGraJuLmiPqcVrHyoNMEQaDpArwFHsh4G2H
bedPzkftgOybgSKkm1aGOLP4LEQeWErkk92YVxGTHxjAtPsXqx0OwNmfc9hfHtSa
dJHl23OHO1ELGWeeDr3FQzX2RB4DpR4brndr1UHDH+BHtMA+JJ4991G17morV64S
483VUTf3ihfnV4RH2mTrJj2WuAYjR7Z4Tv/LLFGVeNWcyr8qrpZh9xEmCtS2hMmu
XK2ZKO6zCb6NaSVX6sU6uBrYEB1TvPpBvcbWLjjxafbPXItFwSy8ZRpf7I9oW+nv
FBwj0QfOu23V9oN3bErXoWrBwzP60O1lkOCL8gfbfNw6NVgPirxpYnDp6STz629V
Ukti3Z87/4wRMVCHh5Cwg6NWCrX8gCGzg1xJlTbWPfTrAWPr7sBSxixHVZk11EXp
uFvDEg1+9sGf6MMPhdOADv0CbCVCXqc961VH6fY1T9XvNQMPyP4SLsh/DIM+amrV
/DfluX8m7/ny8xdnKrcK8bJss3gZSSfc2h7agjDAzNCAFSG3WSBudFrVXUK5w0bv
zGTlfbMbDbcaPBzPvlIKWSkVpzGTnNT87/Ry4imGrvjpRZEY/11gYn0KdkpGJESr
7P1vsLMKv7xoQxXfvI4vlClO1x7SOieFDD3pdsWp5s50a5jli21co606FNqAcnWn
3wQcXxBleeGZnZuPu/ezK1EFAsI0e9BtIMHI6rojyLYuAkpcVakqBHQF8gv2lR3c
q1NTspaYCd2h144LpG2fkfSNaDPgZxdb0VKXp12aY6nzJYguUrlolPQQw9Nv7wMw
tEnkpSClLDzu8YR2UZngrrwumpenL0ldpdCKveV/MBRvaiUyRriNJY/eSyXzejSV
bsQ+mWFIqkO3HfRkzsx6wbkMvBXh2GU8eMRKEirGsU9Pg2an7Tdr6CaO8cYYjFB0
n7gF6Cfb3KahIr8rhwcfUCX5wu6ix7Q5qIgOcMf4kpHtXoioofX6QvQ7TvbF2QWr
37OF7Xw7bdKju7ebQnTtsUFJgTqb+8IccEfZjBskbxw3z5X5VLsONAvk6uT1OBcX
019pZvBwG5WtA0psMMRpZcN5kG+ZDEaHr/Lzu1IDz12W5pbWJm4hBZSwY5HSwEvh
0iaiWTk2G8218kjX0OdYO+NMCJ6ZbpliN7sRVfGpoPqMDJxXKhA8i37/kXM7PV0e
aI00wtXa5taevfJgS9uF9MifA4laRfjZ4DPrKMg2PBnZXhSmoKcY+SnNa1St86pY
L7ylx9taKLCOOXOsWGPdVzkaqWCBE2RAgiIyGy318NtLmc5Hutm1XGpyUTrYY6j1
kdO8Ok/Noy4I/G2uIog5OoHeU9a68VTazhXj3Xs3uAw2Y7TuAbV3p0EVireozopt
gdNWRMAmNH39lTK/IbD6OczcnvHwcwHay9vWCCLTWHn+VLQHfbkZIiBUhsNv2W8D
5SDTv1qyP9tNduhLAVAF1Di4EPY8r/dSmIjkJav4To7kj68JHWjV0P6gXQVWDmuQ
xik1CF4DNjIg0aqT6JYI//ZHVgmerlA4KQdyDlVnb5WPIIzXNA9PHxuh3kIDVEF0
D10xZL3KEIQLVabtx1jamdnYb/UwgJkElnhUKzTTnPkrzLDrd98JLiYWSfCoA0rQ
dpMXIs9ve3GshNo2TK7YnN0YBGqUxoSIzJ1/5zao2ENvoeEgjRqP/0mkZ7D41w9O
9Nc2XkoX6CI8mDiB1Pe98IX7SUtPSbQSEJvhe04K/ggqE1OeGvTgG7iY671Zug3e
4ZuuJkMn9ipfSgUVJV5kmoT2+RzDi2EJT0uHNPBP+GmYnG4t8s0bxBGnvTmMOeY2
l4G6ADNRq78vxlA58JDqzgMX26xXRKfR2pAKCXqLeIFUYlhAm6XUuq2facPJgdPH
2r6IpZ5JcwhJbuPGTFoA6iwvK6Y3CHfDtXguSUlFLosIerYNhbMms/obHIOStjqm
u6VvHZNUWOYI5hKqPs33912lDbZW4uXzwQdG6qdwGzp3m7i33BUs7mIn84a5YcL9
X4FpoteNz2rEOEaU+si71vVv1FW/1NnAJxhYUgP1HP0q2szuDHjI6SryfvdMAlcS
/wHkZHcjKG7lYqD9D/zHGvyR4xG2J235vrhAXI2Tzd+9skHgrKV5wRffiJDtrO2X
ntXPfaa9K6mYrg1eATNYhFQc9HH0WblzTyyrGZnJ2Bez3Py/crAymyobcDwt2rJ2
hH6BWCg9wvijzwd1ceqIPETfLB3aYhbQT4rAeHRFdZHEN6zM/NQKInjBa5X+4hHb
3yUSNf8ghU5q5gqJoWKW9FyBme3faH5TxS6v5VCAquj42ZXAGzJWqZZSxVqviaqx
vNXrno6DOuSu7/qZa+ISkS3l+8IAVSrtSU88Gc48QdFJb4oBWtXEv0qgRTm4a6zY
YGuTVdOnaM1SFTlRIkb17+DWjWD6aIlPXOgacDlCYpIWbGU24SlHPYEpB+d0naIJ
fgTpfkU/4ivfnpFCO7K+JKSnZiSFQbKuXWfy97X9Isgxs9aGEHF+wrY+/wLXHsXb
RRQkrNOGqpSMLJJT5kTmb4cMSr9IYkd34SRPXRejmxQHPylYWoyJxMnY3+3eWGk5
2NQb3OTFt7zMur5iExOzG5tSyc8BHAv9RbJXS3LOq6OXZF9ylIt9ZL7ur/2VSDGH
p2wWq/x7pVUaoceRc6QxsaeJzHOOCk4UzTjECsXgejERfEds8gZyv585tD3PA5Ig
vuO9eFkP7aXgHyQNHRl1xnmTKgZECMlPKDEF+6hVE+AP9o/f5UkosSBMg840D2N+
G6dqXifftXORSNsAe20FdxKdEMVlyxJpdyffIf4eRd3CE8pe9cQ8vKGLGnOlOrtE
Hdy40d3c3L38rp9phTOdXpWi4SbZxf3qXv9kQ/R/3ZwoPXNAhB7hICS22s+Lo39h
jtx1CNjMunrlneXgYI7V8krlQVBvdjP/W4Nmu+OZBdTV8a3EuOYK030Ic1s4VcNE
wnRRYOkkBrO2e89dpSfZCiOsG2NxFaeNSpq8IrYjkjmr0FoMlrp12lk9IgjnoQI/
sFrQ4GEJXKJk7w3MK9vEXQj6MI4lO+JGfw9nQNBCy8gFdwumEIT5QcGBOOKfxSeo
SB92TRDVmc/EFj7GfVr2hFo4ITDGEkIQePqBoZl84fiDT46ieITfjMqx5vTz8qmy
A6BSZovPtygRiMMjxRHtUvQGv/KFI0GaiqBcBq0o9PG0r2tD/Y57mZ5Chws2tZjr
p3rFO67EA1V8Tq0avTYXcnTKKNe1JEBuooKJZnWEIVU6cFptmGtR4qmpc9e0Cvri
Ub9Ki0jv6MUUN/GJSqMepu77gOtcnplYEM5pg80rAD29CjwrXDDmexszBOByRMWN
jM3oGvHKffp9iHg8N/oDG3t5IfMGQr51QYUHPMgisg4+vvFjjLJhT17qjSyVk6f3
MTQcVc/PHiC2ZWlL9psmtmzH/kO43nLUPxN5czwBEtUtD+hcPdDTnXkY9SH9COWK
lvCG7cA5BijYrbGagUm9pGyPQfFUXg8cWxwY6DGg4I7tVH4mu3AtEL/8RzVRKRw2
zh9nKRtzJoibEq9o3eVqpcMaFc+PEwkMNo5ZejPB6KPZadBFojrRCzMwD5qPUOuV
aBHvI1teigZi5vDmAUVJSOoG5cNf7VcCSBJ7+bMG34HdGGX8Rqy18AEllL44LNkD
BhQ6uX0c2yY2/RUEm2uTmohjhHQtMdqF8Y1yx5m6DJLWgzZK7N5cp5ab9bFl+Wg1
rQ1BfSy1rOcqgO8bLcDzoLFpI1MFQTz09rzTjYQIEPWCieYhpWyQFTjm2Fpq7kcV
KAVcu40VNse+vXc1P9lPmhuYPJWTJbMU917T609K+iSspPZiUiEl0sX1dd3O/Geu
+IebV8VVZMpMcsCAlCjQxddJJDidedaMWw4S0asOw7lVx3SJyXSRN6H1RAMqU2Py
AzNBQVHFE+BJje7gUxxrqDXS+o0Og390BuGMAE6NEVR7W91GdKGKTKLYgA2re2g2
eUU5+bpp/Sa5qAVYA/KedA0dOh8Dwzjxm0OmUWrmE7/MWtWrlrp3NUPaqGQDwWhL
NViYiPrStmuKeN8FScbGy0fwWKPOUeEO9IbUSVa+uCx/lcEPN7L/zpwEMcT69ZzZ
I9WXVGVi+27UsqLBcnbSAfvEr+jrc1NYhRZ+Yc2EGKUnl/HV+L2oZ6fROhso9Px5
SW7MKWZ6D6joMPY/PtL8AHpEtVyJXB+66l+ZKQ54COB96ryg1JGLd+JNlvx3xgIE
Wf057kWu8AvuSftuStbdIEiK4d59atYjb2nG057MTAw/Xa3J1REHtAB0eosEUkzj
5lUPC1WNF1j4fVo3eZAq5+WtgF8bvoBP72WX9KUnZeJgTs5MjZhouGUMD/Z6wH0i
DcrMlTltGsdtkv2NqSq2CRw8toFLvAQItsU9DyOmgrTOb6dsLtn+nNic+RMxwwiU
b90borBv9FZ0Kb/JeSYLi9tOnxIUD8sSM6dlxNMjrctN0ECE2bknXmdbaIz0dL2v
pZDJftbHMDNS2HFOsIDPWqGp6sYa8BRh8GoryTGA3HFCJwQY0qHmAQbz5nQBg75Q
CRlrCMNB2sV2Zerj2nLMdZMOVlom/TE/3sKn+MC26Oiej22F2c7WSrUANubN/SAy
9YYq4KAoEy5weujchpSM4Z15nEBZTxz7MEahjx1LrXDypsAAFZu6CoJUYypUbITX
TugX+rJkFUU9mRa0VhCCBMKmUziMGO9fQIA8lm9r4Kn1RG05DVt8onufbAN2EXnJ
NRPAwSWn+kKcea1qN1rIk05yJZGZWO36acURZI2JTLnSijqgcF7EaEtCkVVeDkYO
waBvQXKuqrfulU9O/gVK1hq14sZ+s/QD8Qf1ERazK3D0i+UaqoEjgyhcWj/we8tN
6s4Y5Wxom8WPqtgspg4zmcZSM19WI7+fJEm9UOvcDPrEfaGowOkkwurn+SY+O92H
ppsCCzC7HagzUtrYmTxFtfKyFnvbuKBwGB4dOzD7qMAdsiQZlY4dx2bFhgihEHQz
TPoAhmv1BMv+og1qUlfxh1ya358o4BAVokR2dT9X0C83JOybq8BVq2Dn0mnhzpA7
tvi/C7HTUEyTGibjut1CAsWSKhxJLTwFhuaZ9kMo71bDMfnOPvPrO3TsaMX7BhFd
NFZNBpZoUPfyql5Mw8C4WUwcu5tiPCWIlzGlsygL1PIGrR2yY+Dw5CrvyqYMnih6
/2M6p2B3PsZwNskJ0fHtXbzmfUEW1DDHG5gm7cUxfT6Erx1sjjp3ZkHbGypZy0di
mZ2UwAvJEgJys63sgNm3BSr+AJyAvZiqTmcJAnfNlCtdpvW/qoNrwAEKh4QQSfei
MhCbWxdxEu0Np1DLvw+4MNrgE0C3d0L/uxGZf3m4sOqvCHzp8+DMUccBjL7b0T/E
fDrWtUt3j1HwCkeKhwQj2Xq6/rkPBuA9HHTx/E+vjZcs4AljFyDxQCTqwVc6gKKi
dMVMbIUQ3G3ygX3K0d5l6bRNr/o0xa7KSqLygMudwDBa2CTv1aPnGJMscAz2ADR1
XgBYyjkZwMl0fc01gTrUtIeZg5EhM5dnjOmf6Bu6N9CpG/I7jnAxYIET9C23+OF0
41Kh+QkmacVifm4ckGuPAqnM9iTU45NnUQZPnRB+gURS5KbdT4L4evgOg45Zh0mK
2tFMq0knFhO1ThkVFgmXvAuaP/Sl0x62861L+tIF5fUhJvK2S9mldHXvB2hukSxY
GrSpZ67CFAYBwSfDk9bACq0GBLofF2BSsvRlhhsUE/6Z3pQv2Lxgmz+4xc/Ca7CI
gTwaG1q4fnffLCMM74lyzHoq/kyODZlCuZM+wcZV3CG3WzjewL8+/3b1jERyXc6D
Io1TgeJoOeXMlWH/8GPZmZqtmMtrVFXlwt0awBHzyKOqWeowsoHaHIeUncrD92SP
dc/km9+KR9MMfBFy9pYrAC0FIygXDOV09h1Q5/BY7FkcIYsqhOOwYCAmjqEUHlSY
+rPh6KKttkTAqK8wKWwENvuKyEnCo5yct6gPPtaMACp7znFoVnWPC+PiZIhd+yAh
6xYlujQ2nnElHGiQ73H9eiEilWfMtusiwKHaRbozNeN+RazB/Nhf3A1bigRWGKc2
D7xshGFHLfhgmHpDt2RVEOPmuSYSISF0IoV2lhHmS9st1Dv/d6esRqCp0qkokpup
6Na2v7olytT0ff4Ivna56OkbhBgxqIxLhk5hTGQ57feeyaVqdIkwnfrsXIcEkFVF
6nGbKX+dyYQxcXoMZJHqK/M4zFOqLYz+ZCjjY/GIZOFlHvDC98x0QEIntLEUEsJT
OqZ84A4Qyyal7Jiw+Znl84UVpCYhkljjDkxL13epmvJtVqA9/8wno05p+rMQFtxu
4TuKpUwN1cFgnoG1TuaZI9WembtF1aCZ30Z6k3KMO77/5pL0Fr3aJZDr8N0jFKiH
FvAJ/xp7EBfG7w6BgSk7/8z/Q5B5fSaGfXAGbtjZ9+72Ym5vT+L31WSBF8eoAnWo
0ufl7Mry6eeWinwYk0fQOYQQ8yHKed0Hj6SFXi1Rmh9yxwCe3ZBti8goxsouOztv
aSuz3R5anoJCfOwnC0MX6MXywtHSt07Rl/osmyzb874uB5Z0RenrjHTMRlsFk7PA
RSt81PWirskx5TVgHMGSTZRpoBG/bZZeMeViGkowmJYMxllQMTygbv4G2utKFMw2
Mf3gNnm+5hiafASk5CAg/eYJ87M1WvUBtaZlaRr+czpfpt4+6KyfF/v9KncFy1jV
evl+eWKOZlEECq3l0BR6pNYk9/MB9HP8PdaBW7Kv3Js8ehXYZvG9lDUHt3jraTJd
NboS3iK6S1B03d9p1uREWQg2cUUlNO0qiaS03oVWXNVsQIsDuZUjAS38Hwe7QY74
VsMQf2f5Ebhf7KPKr8IHjlrE6dRC6w111ta3Eo5E/5Nwc+5vXQA3/j41JAsDS8D0
w0HLwU3kabuVENNxzaW8q5yPtKOwTTaaIM/wZ3W1ZjVU/E+l+V9i8tXZ0YkLezK7
DbxgGudw0lRBHhLBMW/f3ElYZlcGDrjPRvSkPwHPa6dnBJt2LJWaIe5Z3bAblGJa
WpHdn6aEpRCEEzE/yjjgaxg0u4ozd3+Re8bvhBpEhLju5igJ8qwrMqFLBkrKXGyY
kJp01jYa7k/9OcKNmdpVeVOaB2UKTWisO2Cu7WysI5ML7kQ3QzmIb2QlfH8jQi1h
mv7JkJYcIGmcFu9XPmUEuEzfqC/COdozN50ks9067JiijvlHYpaM6/T7nfz2Wyjc
7NT4Z4yunHk+jFlBDAVAwawKULZmg/6XU0ecLGEj/BeyWUge79dlubfVT5kwFl6b
rAWHcIBiqMiv/TAFAJUFpqWl1RPD7evD8Z9ItwJlaCE1P48L3wSNrJY1Ea9jfLXU
Stmv2RfSlSHklKrm+8ylk0g7/+p6rab1EKBrz6B2opVt/1stetcTKP0chLlH6kpU
5+we8NJ+x/C3RAPEOOwEULBu2fTU0UA9wdfNNUfLIFzinpJwJyeqt/epF2RSmDfF
5o+3eq5ViAGFkCFp83/c2gqzbZcf5+ru1Q6jqeNjtfqdT4NJgO/a39o7PmMDWzt4
VY80ch2K62/XwTDPWRJMBkfp1xQ08aAIXSb8sNieHgrZqa+bzGPx9Yu9wimmgNsC
uj1btwvPkdRe6+ZgQ3MQ8lrF6ynBwAyAWls2Sgi/6ATwC0AHV9eVrKYi+ZPAfbw7
+shyBOK4xfunND1Aa/IhVkx0RCDp/TDTKxyWbYoOBUU+aywjuLQ5swQtrw8ybStq
F0dwp7K5rlxijDMjwYeBJ4jOXIYbp4YvJ4NPTOWZdbzpvAzn4NXF3HPPXCRi7Wh7
le6HobYd2LWc0s849KnMMnlh2veILe17tiZk/Mx3dzurGKrK9tTn/fPycDgi6SrU
fZVDWTPPot/aHB8F12PamNNiJYEL2uUPgJSiC8cO4z8wPJgKLvrHgD2h82UFl0H8
W5YwzL5seA6BgxTiJWILH9KN0pJNL7sIt4iClF+lQDBBhXmrbMDe3JFh+2a5RKXs
vm2DrCVGVKbaUCtAgm8IvLft/Dj9+9DO8BwWhokUBDqmJac9FHHGdVVY4xK2cxF5
GtevQ+Q2PVjIXmFkwGWG7aWh2/qJ91CRP0XqVJQZUP9baWHy7cdf1ZaCf8Er4BSc
ygiVSO4T1pEv6YB/YjxlNqD2BssUVsCShRNEftredupktYNCRgvUF0SuntjkcrAt
ubqCOBhDxSBWjKTYFuUhvrJTBxR7NTlwoxDuQzcuYKm0FrCrtPwrstcoCkylAEHc
Xy7LlBafi3HFNbcLlT2Aj8s/LGIr1R9PfHUP7NAdknmGXlc4zWJY1JX5KKqR3Dwp
IBkfMwyF3OPyBOUtOzjBds8Pw0VLcjWMJJWS1UDI4rnXkj/U9S2+NpK7/W9nei4g
CBaz/FmfWhv5bJJqLktKW1H21Mf76WB13WnczqRng1e9xY0X13D4PerYf+faAVOV
yywZdR6aL9hCMj8YuJ/I0H+zjAoD2N4e3i2MEuNA/OHvGj8QEQ3qC7YvO45JmqAn
9tQ4jt2Iv9Bp3g0VCg3OLgpVpNN+hq/eGBV2ahEcVYIkrahBVB8kNS8DRT4hsh97
dT7ZA8gH8wuaNDN1ScYREaI4Q99b4QxBKsK854V1rP+zWQeIl7NKk81wmxOCiQsx
+U9V6IPoQMquhZFhK01OwuZED1SjIdQHXP4coEiBoSfKcx8/hYyasekpA0izYPrO
KmuKmUScr4kN5C2XAai/MWra6ZBe3ejFNx597ghEYXvVDcquKzK5zNHtfXv6TWWW
yWPoJEo91DlI2Da4WNKlgAKt9TsNcWqpjo4lE2K5Va/NuuAtvM1GXMSWo1FXqCQB
aNkT0TtNI0rCPnARqJLQhcrk0FhqY5KK5J4Zm8NlWkyxZDfq0IxNEZ4uUpSYfAxw
DcFsSrLqnDn2d5GNKeLOPfjdXaPeIDQ4C9I1fT4lP5PYKXAAZTlAJ1TmJe3y46K7
gpNM47p8gVPiXEE12ZsOROfySR+mTPrJrLjoBAXUbHHopKlpD7qmRgEWQ2FT1x3G
651QEwWWWxBVn7JcnsyIamQvH3+5aNMpg1+lxlxWAbOH7t2wrk/dHj3VXm9xIIlr
p6Pn5sdiuNnsGxVbZm+AQR45IFCgnMDdfOZWkKwfCmQTmSIZZImHmBfyHTQP8atd
Za17+z3+SdXLkE17vW5CVF6VZ+pt1lKt8os5XfCt/tmwO+SNWa2eTFqf/os1nu7m
E8xqdbM96+j4qA9OnmXwtWlkbXb2jGvigNwNS08USe7XoQm8QiRWnCPf6IuxefmX
sB99MLtXt3tVBBscdHqmEV/u6NTAczZMOPtvPc2HzV/LToS1t6l7lfUIpJNBMQm1
AsH6nhqnNZZXbJE+MrEpkxqXcNUriIn90pWq+xI+q9qbGB7lvabuHdafMhG71D7W
skWWcwh3aPe3cAqmfpM4HbH0wBUDQyjH8o+gLID6LzWxVvm3C5pm1p3uN9FMbVf9
yowJ4i7lPauCE2uEGcoKbELJ0CnkJ5NSWBDgzvXDwxuEHv/tB/AbtUKREbvfpmCP
mH8MWLYNfx6yprr+q3eG4GbQNXi94NodcbxZNLk6KjjECRB9dDQaWuFZMwB/gSnq
J5jUsZPLn038+dX8TX3QztfytNYh3fqLaAQfcblDF/9LiknsxKB4SlAgKJdbZY2X
ZJy+23x+qFZbqkkTadMWG8ovLI9T+rw6UsGFnWk2E39QpkuMNxOMs5BOX4mAV7wD
LHOFOvqV6IRe1HnVPIy2Ydh5YGo4+PXiE63LZVKgACqgGBmVqUwxomfNBeHENdPb
IhPjQlj5nmAjspqyBy3hrUKK0xm1Ks8bhN482evKQ68MXvXfq+9i4SzEzEfe7EoV
5Fg9WIZU0WOYd6zuKXZF/AUFRwvetW1dWTSIqlZpUB+Dv7mi62RhsIpU7BzQ7IgN
afgIHrEI6eyRFuT428ZjSWC1XnfM3Ew2v1eAQTUURvRUd4X6cZ0EtGPKnT+RpEOF
8Rdm48uwxo7ZmJmRoH2tkaypHGD3qoTHXMofSz3T898vu9l7CzsuE+8qekrAlt6G
MatmoO51g8je2y/9QovxX6ciqIqqyeFJgpMwmz18vc+dvVYXP4VmzOAzkxSTWeLV
8X3ILrUYwGLrStOSdD7xpe3u5OFBnIGP1dJ+j2LG0BGt38Yx9vWglE/dBxb3cJBW
izgNbqtduoRkZH2dL5swZGgfK2kKrv81ghe4okEGbVUwSOrkIOZRnk9FtmBqLKoQ
Gx3OMcvNsonfBx59wX7wAdyNpAPAj+MoeKdYSZ8E4HodOmdg8Wg5l2Jpv0ikl0ib
osF85h8W9gTEMjA+ZZO8YpSXOX77HCkn1p62Mu81d7+/GzBDsbR266dbr0lWGnEY
qmm1PAjQnlC3xzCSXHwTji5I/HUdnRY/sRWKsmgqPgGdlJ5KpB4YxZEOZS//Qorc
dVsBsrPNLUUkuRlOONEByKtZOGVm8OZMeLCaUJCUi7m5W/mEL3a6owljvwWo1c8j
A/FsJJEGMG+fx+s5NX5MkkNvYc05I4l9w/BB3pryITbvJBNZah6dsHnuwE7XHqRg
EKaU6Pp+JAqKD1REv3L3DxFYGMlD1DOn8ySjLBa4V1HwGfOrBzzMhKvx2ia3lmTt
aIOG3+eGE1+HnwozMM51KXqOW6cg7J94Zm8BWr/8hwJBr24SZC1SE3QlrreZ7I/a
Q0UR2qFJY0rUcGwhia3zlVWZMYdW9wgLCh8askcnhz3QPhKpZfPtYpYDaZm9Wv/r
CVIV73v3z86ey1PnxT6zd+PqQCMGNTxkhxMvy4zDaqZg3bmpyhbEA33aLusVaktS
tn1KZiHHyGEl1D2Y0ux5mCS9Bh59k0L9EgFco70yrTeQXVx5+h6cfF/89XyXgFOq
0XGE5lMUA63Lk1n5RefTrrQ44O1SAId7HOQJwT/Gx+Dgqq46I2R7/upX8iMJt6cV
yaj/GX4hfL+nXtxlC0lDw+yuTlRQapeRsKVjheVyy7jkDQi/rVp0eqnm65rEVsAV
4xyRLaRX4MOCDRdS2qwdoKWjY6Ya+ha9+VCIybsxk6TakZK0h3Zg3hBO8cYfZvnX
RAoKw5o/YyKUpmd809XAWaBP3kw0gxEUBJdx27eNan61Phbzpn9esn6LhkbkJLeT
qgxoT3y7FyMuGe7xHHicbZpLnhOItIHEqth+A82yBPLimycj8wcgHU5e6eqCuizS
tSaPA1CtEWaqgCvKwcPVoKW+RAt+72PP9m+f6BYngq+6Kol+ee/SA1O/qH+kRFVX
2ez2N1E/JFEBL/eMhxZBzxVmJPoeXBI14ydNRVHFwU7RVpLU8oJANUUri5Rg9IsB
2Oqbmp+Zne2pXQ+vgOLzUqXB6hhW9b2ewdsZdIEvxtK6WhZBd4iaCuaf6gLnsd8z
Ri9pJ5QBUcGs3qTOGAo9f/pAzP9YA22fjPBd6AW4Yg4YDqpp/7lLns0T0OyjU/U9
ofmAQIPCwW3TjCWsE4BftIJ4EQOxPczgyH7Qbt6NBB8/A/l2e1viTKWFugMHJPNr
wtJDVZNsCgqbt+ycR6dFd+cpvoTgWP24hcSFcmhapEVStKgP30T1+HD4oA1/hWhD
sQGj176AjC52Et6808D72WEwPvgEKeLM2yCQzpFxPUyZkvBTiRdQVzNKNmvUXe9f
KB+q2WWs1k8OllwKbm7jo58M7pYSYTgH0fKXkXq3Z8Y2drH4znQwvi/1YB8aApWx
0UCmHGirUm3UfFLDKcmxVOaeNa3nc8qR+MeVqsBpUW69c/S3dk/vR9JDrmpNurCr
vPJQnqwCdV5jWa4sEJDm2iDtbqRMVlbuPipCdySaokgCxPwsl82GebfhPAOLkrGV
CiU93S3SHa+4cqUZCmgWEv2ZW/Kf0T+9A1ybredxFKyuvilBsbMSrbhfZe99cx1y
vaLQWRK4BYkpj+Z3Clrc7CDDhSiVkQh9f2Aqdsc2cPtLaKAktH/yi9ZHnlMlVlul
5OUv5dsF51nc7FCe7NXv6L6QZcX2CTcZHpweEasnTu04VDto+eGdduvLBZieAa5Y
jKSpi7j4Nvf8sKZwWbAk8umjrabtUi7WSWkXCb5Ro3L6XzA92VgLdHBBur/9kfOt
+tBaJPazabjWSu0JByWJR4ixuUUUtNQ6i0mQJvyxIKSprWoM0eIKD7wFfPtw2i9o
uz7m0oUkdSPiHZc2SASVTstQ1kA8J0GYpO4v7J83fUATVsDbwLebSyqW2zbYD8JE
2boqaXQfbx42zqY1NcL1ul7sIBqt0o7wKsmad62B5u48KYNzYbNW1QnIgnQGqm0j
a9yx+65GF5ecUQ622g6qUxqg1qbq+XH6Zm1pq6GaywiFl5++I9njp3TSz233XLXZ
H0u85wyk/9kNJeYrjOpUUZtrJk4oolIqDMkUlIDXFsuxKc+5/Sblkp6ouM/T1PK2
535pDw6tL4XzBSBZMLAestZmpbwFqHIXDvPV5ZwFf5IKgqG74ueP+GuOzvof+CcI
Shp88xAXqof44cmX9ZWAO6uYXy2nO3k1Y+rwJv42UsL4OvmB3kGbhHJOqYoma/8p
GMug9JcoKfjSV5Eofb8OAr2cWjGX6RMccpA1ziST5FYwk4YPnZG9maKJayeXwFut
5LJfq6F1KI5VQmiMGnPes5mncIija0f4Pq8eorTwTv5g1Kp4IeRQ0xU+L83YJJw5
7yHvFZOJLsBybapHxA4rns4ydGOd7JzTQHAuZxw698zgnCA3b1et/KsTJIR/4pJh
qiR208gM4JYPUoq793a6+4NtOyyNOfbXxPIZCj/0L8YuAw/GYZFGbPp5J0Iymp3h
Hm0Z3z/3orkwy6kj3VhA4eS5fs8rD/K7ddkf1+6gnRruVewW0gjWD0oyh1liXxTD
sTBZjdOX2q62EtqsEYer3Z8f+kx3x0zg8s8Tn3/oJdtrvXHMsJTlssakXhMb9N+X
hbTBXz5Pe7QZWzJrlAbqa6ofTGxVFYg0DveG9kUP3O2NANTQk/fgVW2WjO5Tv+pO
KY/hhS8tFfnJu4wKAI5HeSjewjYfrrydefnnN427WsIHxXEr13y5cudTWjUfMG9s
SBgJyVoEol7GK9y9IZvldG0hxM5DC9ZKo1Qh2q7TQHE4KTj8aZYUGpJVBWATz0Gf
/qGR4CnPC0CE7q7YELHJ3KDpLkju+NSQs3sHiTQVKBKbGRQVNpQwrK6Zd8/qEnd0
NVO/f5U/KLV4/g7vifKw1Cs9bL6DNSwmOjMyNvL3zDKBK8F9QE79D0t3EhxFaK4M
9hatCY011AEx0d+9XLjcihJiJGYG4ZIOiDODjAef2Qb+Jod2H58c4UpBqgTsBvAo
tT7H6xuuKzivw6ABhy8R0QDFcgClj46N4sWmY3MHVMfXDZDODY+DlEVo3s5rJVCQ
keWy5nAQm0YLVJ9cMSLbLE179wl8ofw6JUNqdgJNE0kQL+A9m7CuRAW+T4v0qC7S
9oYb81xDVIC+X29Gu/cAbp5ycp8sU53TcgZe15WIhnDF1bRc7PSTnmgwzrKtvKGE
LJRQeiKnvqXs/MuW+41s6oiiVwZV3i7Hbcs9w3VabOBR60bRex5sd+9aLz6CKaCD
3V/qcG6VkdyVaujl+0Xay38JdQQ8O9CE2U4KG7qm+Nnps14X6lRAaRg/VGtxuAo0
1hAtLnp+skvLPM8PpjDQog5wLcOVdfaHFOra9+5KWC5ksSGhR9KAvAb/tqCAgIjk
8vhW0UzmhEC49BSMHX3CU4Y+YbSUKRCzGktLAqS5JmtNPVKhHzS4hNiR1Qz8wAzh
1TVgfKNvxjdQt4r5VDkKBCk6VMk13z5HZFHjMRzZ2Laoi/yS96SQeAgFFhBVzzWW
f92PFcbOsBIXsb/pl3tGXJ24E2cRNjO1JbyM38A8o50BT8pWZmOIT36kSTQpaGzr
LyGiGmiRV7qOMtv4XlTyy0Fwu/9L5/4bkgnJs1b0tPqiBjLNjrz1fDG64W932yb3
67Zemg8T9ULS582l4e/c0SidD8vpo0poHqcpiGPPFdLGf7IKZPQCT9BrNG7M3fpg
PIDE3AY46OIP2hDxZXlbNiS0UpPXTOdtZqKtTJ20WrZQ9eynmtWqr22oKDO52fKy
m5BXBUr2oIqe7LW8pQ726IYEg1g3DehNXSY9q8+pLJ2gNdnIc7SIp7S85Wbb0oQC
H0fUBJdZMhk59fxcYEgVpAS7feonLmilKNDW+1TkgzZKgXowZwmjfxSZ5CIT8FK9
DCXaMtoPUS/6gZVbcIMBL7yRu/e2/suupPMd1M2gpQoUgZfp/azZcWv9nN8d1Swj
iH5AHC0QKO+2THKhE7XXWXxNcG5KocF5kQ++2k/ZqpJNnEyXsDAixx771Y3R369K
eiPxEfYoTZfO8LV5jxYUbtfRn4MAsBOlrqt3ceqDVN0KPTJ2I84zmOebcgZTOYo/
YmrfDEeKV0a2/Dfova6HzWMzUUGa7sPztUHfzvk4NaUnYLqvVxBid5k0FWHzIjCp
WVQ3dEPnehRZwEAPoLS+cDULXRfxw6Mbysu9HncQqLuwYRqx9e5TkOALl4MgM7xB
KIylO2n5VBAeCoBH3kxJKVtN1LY5Wv3qFXk6+hLQXwiifDcV4yRKHQSh1BmM0Vtt
uMWVVXqX1N86VrBEgMfPUmFGIxwhHBHG/mS5Y+CedpIWOOtr6Hopc0a8DC1X7S+M
dAiGQ2f3xDwe7PBQ9xaXJOOQmP9C0QqP0tPoKxbJvrk0Bb5N6b+dRj+NeEOJB0sP
y4KcjeTB7hblS4UknKfEgMMg9RQiMMLfjtAXdZD5R3zKPqbz4MeDPMQcfiUku6Zw
quJzpSl/EFQjcMm7RJgWS4n4bDT4STtC+8FGaUHN59HcOuFKVb+Ubmdl87cfQeq7
ihK2UT9bzNFl+NGlU0g+Rnv3KnwKWjSBl5KUsCbGflUAW5Z/xnOM4+S5A5Xz76n4
DKKucXuWWDtaAiDUht/JrS/Oa3MJk5okH8eYAJdPDdFiFvIhMVdOdBr2KoR3ivmJ
WnyO5jordu2dhBtAhHHhyvKCvyR9uhUzAWSWnDjEH/WsFfvMn3th94TPeSI8TT8S
nUM3SR2IOE8Nbdtesic62AR00NWI5LqOghlUyoeVmOj8yBB+2xSE07bRgFmY9r/I
k7PA/E3Yh4qFuLeHbz3g/3FmHesJw//A4R7B9aqI5DGek0ZwcqNs9qPbuGp01bkG
YBF+xDjXkapBOyPqHsOZTDf+WcZK+8RNBu3aiMSz49dJlrChaB9qkJktULg+VsrQ
GjSw5l8rosLjk41rkIYZ331Z7yJpzc58L3w+6vIleqVu7CDlDsYtX/C+SuNz+Il4
2CU7cpJUauE4DKZGEYrXGs+3z09WHlKMxwgCxkNhj+bMxH7TzaASQC36jaeZjPIz
CMqEJEF/Afzi7MHvgH010Jpg5hDu2vo/lprlREQreBs5BUJ8uR/B6ewnhd+NkqXq
9WAdAgExW3Q0D/7wUWXo1L4OdYoA5jQCnJTmalJoB67+Y6EFfpyyULnSz+qD7BED
I0RV2u8dM6pkFwNLMDLhbXrEgheESrt933b3IrBrn9Zkr7VwzJreJTKP+u/r0YqT
ZaU5DUxGmGX1kwUTIMc8kkUUt/N24HKaessjky0U9k1ECjEJEjIPKE+9iy7HPeVP
0XuCLWPlCPUPRIHAE2kWJc03TAj4dkBN1yFOZ2e2elzvBWz3h4LgaaUbPffIrOYT
bzxIVF5tJ3uu01A09A3vPJnsbSKMCQnXVm7YsJ0j3rF7kOP/v+pyJzhq1iC24u7q
uHfZn0s5iFUNm7jNG7Dt8pjLV7i+R7tRp1dpiEwT7oxIKndajKHNK79mxm0sdg6k
P3eB/tiPauW0QvXxLSKvnqc9mIqI/n9TE6N4EzwKhxINKNF/DkNr0zB30TO+We+i
eNK4FvtsTHb+t3dSw3M3t067FehqVEvyN1n/zaYsgwp5l6Zuqe8QsdvF9nM5EplA
kZOqjQsfrDPYzGJLSA4Sd90p8GhnQ6EKJVUwqeCTaprSq+DRYc/Ihc3LooseLb2T
42tuidDTJP04voUfmwywg7X5UPfr68rf9381kRgl1YMZBHMJ24eiN9DTCs4AxDvl
kFwgl2gU5keFb4K221uRKskjCQgzFcTRu2dzYMZC7m2uz6ry2ONCXBdNfzFFgwqg
oloFUyZyUq4JgLHFqxtzoqbGPgm9BK1n/zsOE+v6plL92TLa3jIeOb0eqVtF7d0e
Yvp1LpchSFIE40ayZoV62bo9IERfwYIVm5VEG/PWWCQiOeYQGGthTFnyebFeRRLX
BLbUf+iwns5PTcQo4Q2QM3K+v4KsPzySHvxn/vpxB6mEXE/7b0dFJuCSSGVnEN8j
EY2CffOesPxLQSX3Mi04+CS8KjaYrTg8hREXdxrtciChhX2aRmFVRYU7prjdVdNU
WQKKqQwzLipyZw3bldrRFH1mdAG8HQiBe0AeCm8JMQAlcXAaVjNDOmLxQ3dbwpF8
RBli9ym7wEiFqmMPOFDo2XyUHB4Wv3jBoyaUw/H9Jxh5d/8eCAgF5HLWgSPthAiW
VCP4t7kBpqHclMenfbTXg9CAqR+q73wItkH/WV+XK2vzYLU2sA0kYbMx012DMFm5
7Q3zaSa+scP2lU6xhqZ83C+2nYElR4bZThF57pUxSzowLEZvLb3XCXjpLF1aEmBv
pR0AlNiUzQQGcdzbHkVMHXQLIfVHabOr/WsZsUj8ghYD7AM4bPDyyJLIpGeXZqs+
pYQEQMObu4NnHY/88i55m8rpOdB7g6Dce5RImnMZ0hhNK8pxgYbsz5f9DN8Hwz29
WfbDlRjbre4KYJiN51Dk1KtilhKmAnLtKGHtNTq+zVrK1eE+Zi2txDH3q+9ke4Dj
fMmH8G7nO01FbosOvi+XxtYXZA+3SKgv2HnB+AQmIrAvhDCi2WICsngbpsH24LGg
cu2kCrp2THB3GAIe+IydMiparIE50cbpJg/QNVpVAQvZxq9rc/QOlhSfD8VULGBt
BMvNj4zWBo1x8Z4wBbS7dHKPCT+hzksgOahR9KkluuiBPdEYCjWBY70DH8gTKEIw
CeKBRcrgfsXAOv0J4aVZKi/TS6eH8Gc+ci94bynfyawB8B9WjjjXrDklEiHlzlms
PHNGP4AU2z910O+fAD47O87/QChOMivTPd6vPCOW9cO0LmJxJEYYGQU4jifZUyPX
u6vcxIVI8PdjMXkkeeVgPX18Ge27joX91Imv4QD91r0mZnLMIi/xdvDy685ZOt+y
N3H/exEKA8QR8iMdd5uzzj52PgNjRDeAZC5W1pjizXt2IcUstGl7lXuj52wTVk0C
nHFoqqCJP8xOQxhuC15mNFqZZ5BxgoM7Bg6M8l/9sM8I8A5sZmnLPp0VVbsw8fuN
RP+oVNhGr3KqXdl0o9MvvepFipP/reSFyfi2vuduYoXUVaHR9/g8xqjEwtiBj+UZ
aZ3G1AjxuL4ubuYqnGZ8Ym7dwpVG0Hfk7BlgJBk4GrveExPu1RFqXRpNTMLIK8PC
CPfT42Dx5mPKhzWtPtXSY8GfSk1uoMRWjB+HEq8riA/4yluhuGUAm70NY3lm6jcN
6WwfTzaNvGvyc9gS77tLf5Ur6vKRXUDaqh3PF3enwKyUQlNKtZR6arfO46IwBRFK
tvNP+l9gm1FEVb6Y1VWmvp3bUb3xAz7rACxvQVI+xjdpHmN7iFGpowIOpg/+c++6
Jchux4H3KNWiI85w7zc7V8j/dXnQVFzPyxjnJeo8rKNsrtpv00h7SIzIK7YAPLdO
MUaH8bQdzpCeCW2qJvgoa3Y/97qi+HBGXw/e1FkzsaXKZghyG3X/oZAdDAavtPtE
20yBvDVsa2FEYwDvFVWthIygiU8t4KNB+FT0XWYstvso4Ew2wGwaeavjb2qM+XLq
9RjRYnZPsI4paZ8enTPgdb31XMOecPVpsCWbSqwa7I8tRd+V78nk6TeQN5gZzFvu
8F8XGNT9Pt22mT/iD6BkGIYcYhXXwIUy46SwTV+rqmsCLFsCu1BI7BfUJmz70GeW
7YfLXDhq+OWUJxbwpvS7YSMeh0XThJOKpbeDP54fQpeEMYJ+PnkZ2J1WkEmbiOox
/i0W9j4pgwcKN+j+XILUlXDZmFg1uqTeaguosijq5/FUU4IZ19Cz58CNqPRGOLhF
p1WaulAXY2Cc/JX5Mhgor75ge+WI7Mii6YIpRq+WOC/bmNmmP0owR3pmoyZ33S1c
5UcEV1OJE+ClRvi4yY10+TQkZWmXCLUs91RUhmd6TWf/WUSRpvenv6JsaPlvOMps
NIei1bENTCcsixFz2pa/RP7t/TlDZgNwaQhTbVI9dVezEui5UJ02eHz5QKJ3Kpgo
WXycCJSTZDWNXFQFzbzXmZv0v9OE25zFEyxkHU+nNEdwiB6fyr8DLaTWe/mhHFXj
6iBIukWrAmLWtP/yTU/dnIYiqzdsZFlljYLNs2Y5vHS+1Vv1K2TcD+f6T4WXT6qk
6kIcjTBVK8MvY/o2KmX3HG4rP2YxfMRseL2Ae8SeEtepFGduLW/mu2Ui/+Ay/4yU
udHa3rVy47cTcq889x6WKej86NkXmiTSf5jIrStYPZYlDRMIUygUSMth4jNi+ypv
0flHNWF2eULyd2djhBQn8at5gc8E4DmrAVDEimmIE/sGEC/3+weWRzYzRxn4eUb/
8Kbqe3gsRtnwHk1evEyMOzeK+87LNAGvIKpwsi5E71970m4nehdUy9kAqFV7/tbM
Vvu53nwJBGfqKkMkaHlhAOk9Ji6P/hNHap0WTXNF9kjKzwzZDWE8RN2UbQNSM3OE
izEC7LYJ8NzLPb8XL5cmpawHepOQX6qQbrMEkPDhBbk5vM8Ylq8HjiHkTkNqA7dQ
+Kx6Z+gG+xaYVJUxOuXCLrVJ85cQCg3MCIn8rTkleKze3USvmYGjAZzHe09o+TA3
KxRJMRwUpiwuM7hh3kQK0d49ooI9rh6mfJjDnlW5rhT8JvS/ahksL6EoTDp0M6hl
kY03YDiEA82mjTnp2S88LKTXSnzvi9vfMHawzn3QqLU2rKqOkLPg5zU6AAjmRqPD
TizZQk9jHbJvJdtvslyxnQoL/TnQ+MLaiBK/+medqAptxNhBTGWseqFte1UUU3Ax
TaR5pd2WT6bw9NFmiboD8rGMOYmdjX3p8FC7v/1cUnF/SzXQ3gclGET5+6B2Jnby
AD+WZCQutNpyoOlCiJvEKjBQXudmB1Mnda4tn6A2lhm8If874CiwBsk8u3BSefJJ
fgYbLiOb/zpk7dkxYMXJgbYMf/cAzyaXm3xeO7i5cDPn3x8LkAY3OG5mo21eGCFv
kx1vL02kFB5I/M5WvEo1AKywq8RPD4/Sct4DEIr+uIpwDAn/9wFR8xxQn3W1p69M
ZHGIFGZDz5W5jGkWclkd+7VEal05uq3XIveOte/4q0U107BFKlUVR79p4FE8cTGw
0bMPY/dkH5FkhS2mkVoj4zBsn3+25N5juY38djmNNpQWpHaljFWlwTaGY7jXDYdF
+q1yR1P0J+iz+thx7ApiRfY7pnkE+4yVJ7z4cEmF4q96wQAT1Zf6v0Z7j5wYpS41
4Om208dmVz6yc/SCwBt9pvjtKr5DK4eFNzmgI+usjTHWH9GUx8nD6LVjvam6RGXF
B3V6aXshj7JAm98ENtACmzpScvUM7XzfvEn7ACPSWOd+yhCll389husL+5BMpo3Z
4q05sxEBLTgH22+L5rL4HAhSORJm7zE7efe3B+x+M3t8GCM1Y8V6pZQuKcO6TgbM
YdJZBpc2pToIejKYt9eWUC1PLuDkpZdMB8+H+yo8O7Hu6BdAMBEGJUp2anQS7pzK
yFCgTS7Ed+O16rf+C+dZmvp6MYjH8Ty7Xc6y0FJkfBwJuVN9hj3J5eKne7bFCo4s
g7kQL6K5KL9pBNhPCiuSWyQxUe3J33GIfH+gmYFf+MSShdQUny66ertpiFMxvTu8
TNpMKRmkqIn4efRJx/dB0qxlyd0u0UD/18L3FbvJk+Cp9cgIBpTpQ+CkNGYNOpaU
v5Lia4OIj/yGc5ekuDn4WpghBOdabOJFuwaUt8zf8PZeFjF3u5X2BRFdxv0ik+h8
GQ2dfKzqDr3rVBsVYxuiXxd0AVpo0q6PwmWY/8mw3ebmGFoR4CPt5lyQ0h+HSMek
eB6u49riZGKNIPVgpWU01ynmwvze3x35ZvENzM+IgjdyAcZ09TWaWM3vKCB7KoG+
RnzpLqqy5kxHm1YdrZ1iJyzO+AEXTW7O/l6udEVPW9b7Ciuv6Ke2Z3Gqo/kvVkxp
yyVuNpLBuKjAOA14IedoiTAZzF9iM6BS+4YvrKrB+n8kp4uGXlA+1V2FlyvaFkdV
23A+fr0aqdaQIGwDrDssyNXJljtO8JRjbT8bGYVmkiTUKgK09xbYBZSOf+yQfBL/
9zdll7At6TCUg0r4vT3hQLNUj9l5Mv5MrudgvA8q6uGmxTd7qib3ju14V5o53BDm
nZSMpyQCPVlPlWb4neWcHQ+rVqt4U5IQkorcULpzr8OdLMrFiqJWb7m0n89lkfMq
itUIPwbCZAT7mAs4qffV0vCQNlrcnCo8aGrAE34hWqHu9qiWcgfO3YHoiE0IEdLj
h9Q16kMiqXtFA56atzgaC47fUUQl3za8bAiJk6Xdj5ZiVpfunUq+oNY96SF22oUt
uiE2mxmhjdvpzfQKnyqEfbWE9S4NN7KtyyMgX6m2AcAlYAQgCphB/p8EqXVaxHGK
uUjA9Y29yp/UlDQHHvJNs8JEg47FlOaOGNojZK1AL9rEekMZP7+RQmlbBZ6CR2KL
JW8xbOsVou0HMMGv7W8Lhuyi9pzAlmPjgFboOyIrHkG056ppGALdfxrmhMuX2F2I
jGCjZzHXCc04pcW6HOXzIt/8pobZ/A4l7JyED5bPNbw502xlHr1SVGlEy6VlS5AK
46phG2Y4GrBcQMDQTaKQytVNeqtAeRAhYe7w5aJKS3nV/t5pkAjF9kaTM930MWku
anjh1RxBQkLz7apGHfyxeZxa23OllkbVdmTr0sRXH3E44on8S9F0GZK4B/ckGDwl
XlwRMV9GP9eDFUKt80fweU6idxhlrq6eBOsm6oX6+ieCzuu8NTw2t2CPzkNIJQZ+
38nPrWxWDe0Dd+yK67cgoDffYENDhwTC/A810z4EbgM6HyfeycztOto6BJbj2e5Q
IUpr1hhPMTIzo+f6i/8AQTMV934TnWFRDkCdXlbBxdqlON5caAAI8YSQ7nVvzcg8
pXPmiE3fIgZBULv6DnP3sSXlDnk/afmCL9NAX1i50G62ISi1TD55HpGGbYu4jx5i
2TsSl2fsSiODKInkbW0nQNK3J+gIyS52jj3hOx/2KpXOakGdz8VtZm8K/vE7u0fT
i8s27wQfmWUZ7AYT3v4MIqc6THXlEKzI+ML6MYkhSf0iOSRUlBqu1L0YkbTDPwyB
PY7JMCGuVMpRXUG7I9EC2Gh/46lrsr6GdqsJv1MhoarZKqDV+B+kX203tRmB1BZo
72U2Iz3FI3niteja6++QnV72wfrC1N1WSzgwupmnYBpg1Xyt0T/zJ7gncAtc4ODi
INExNqf+0X2KNHqubn4xaGUVq0fu+yaL7KmCEc52DyCE1pzABJpt6LVvCJlCoEHV
OUVljTG+CnmK27Ka38ogUrfKvdopQpOXUwl0O0lCPvM+PvX2CzYeb7re9cWC23Uf
UGZW7DkrWK/cs+Z64DwzsIoayoYvFwFJEOXnfk5mX/U/7JcN0KwViPgT5jp+XlHO
+OYG46IO0fyEx6WFzL3lPmGSknLrYGSYBCokpkGh6xh9EoZe99Zc2X1bwTJUxGmz
CtJnYSupBdDEkAkVbTB8Epl6kORpVk4HysT4z4PGW6q+109DWlm/XtTJ2FID19pk
Cz1l7hn/v3iplJ7V6igWTtq06SxEi3LmPQh3oqcnfYxS10Xj667w+2YTGAm2OJhX
GwW1fCc9iFy1qtwtxnhjcX4Z5dVzlTFwKP6XHLAjaTkQBrLMTG+pJYtTGvOLMhE9
bnIWLj38IlKrJon04z/9ysdbm029FRgAMnk/ScCmGwctTxWTSyNJrERuZYM46v5v
Y3b6k/8a5UDqDDEyk7SyMGP4cHT6vS/Chzk3xjxd202lWtZbDiKUU7wWh9nVERqA
4rnxoSlPLb7ceH3wqkb0GxkQtUWfygpEtaDtmAj58Xma1Iaz5pjRPKCPXnx3UUzI
O2Rd+bStL3L+57BdazdoF8az8P3fBxokq0McDYdNu2iHUnMhIgGlApKeSsreuugU
j/0bXi1kc2UuVyKl2paEzmQTpYji3F0FBip8e2FvSDImMydk2zAzgyNo1zwkiRey
kHFoNaBxCbqh6TiKRDG5NAMuRjuI+H+QH4hQkx51TzC4YWBWt4+Rcpl4nf3Pxihc
3UXUcPnCXejyrHm3O/Od9cXKvx3NcfhrvwJ/NQwFZMKPD4t9zscUfsij7WmKYwtG
29cTSgSVbubYF4qmohddDKtkUEaTMm7c2cDT8xwOrI56g9ss+4CO2R3wmskXO83K
V4Njcn4AyugIFv8r8bJaSyZCBEHHrYsH22td3QhJgRoT4JLl4uYR5n+22dgzFchT
uEppQPX9uXEpr+O/9eFtVyvwzV47ffpnKEwZzymZPDnkDJro4hOM939e9WsOZOW5
4hNvjMLUEl8OWV4vaBkTG8NGQY8Qdr9NulSvpkcmMAGryiJ4CcV6G5KaUkX4tjFq
RY6vBVADZASvTyMAnbOuKFNncv2yNYkJ7UAoABcHsuiN2TjQM6xgQFWTjN43nn7A
kklEY+IOiRC5cwBS3fiqvCUbYZvYsVuP4uvDzr1hpCkw9BRNJZQq/7TAfQOB1t/C
h3dfiMpuDZ3dG2DTvE4Ez6JrBZGI7sK/OZlld29pkUfUslvPOzeW7hc7V8otWgGI
xvftTC3YoDgV4KFzpwv1P4f4YT0uhP0RkNQflNAXftwzvrq9AMZf6me9N7Pmd/cU
jG5knq5JyzsmGG73WifGSonfPtfZF4ycqU5riRQBdSyRfVijYogvQUTfeXBZ97MR
izHOntQ+N/zoVFxpaTX/5+kM1CbYy8VIprUNabMmEjt0jfOGccEUQoHb6VlanTnK
9AK8v3qJGCLNOl62zaCBid06UO5pGZGNaViNUTMiTURrIqr3g6xpTsVSfWxhMfhQ
0+bzMuzl68VFSd6uLgSTIzC6PeRyqqBOl37bSvbXRmlAd+GGCyC7+4vWaIc71fIb
HO1MtffqK9vAwI7n4RQRnvfI6RDQssl/kS0uD0xFL9ylqEyT9RukceSz2WoDqCpA
uxRgexCVKaj9barzZJv4BL/zbzQfXM8oX7rCu3/bRndEmAoyX8LJMrE4yiRpQ2jn
zLfEo3XcEM3GG4IswpGSDnh/IZTs0Hz4YmenqKOSPyXTF+7TUWTZCXHQtJ7B3qwB
FEN6PggHwIRBrgPgs3wM1B5XGTaDTHuwPFCtNG09voh/lhgzd6m5nwrq0tYnXpri
W+NnLO0qndMaoFb8qw1EIZNkxLOdrr67LWfh5OiuPK0KJe9Js+9fx83jbmHquYQG
VMsnUurPl8ZVbnpd1BASlNOsVeTnt0EUq+8QS1TV3P8d8khmiPh4EM9OUU18TGar
cgOShOZletiLb1hbZh9o67dpPe2HmyySTb2IKKABJpClV1DsmckJ9LLjrbx8Qkjq
wBM5HbE9w2b/H1JyEYUwQR+mt/HOP11ptgaEPyKEv/F68IlJQshWfJHjISZcfgHY
sMhjSz9z3Rb/Af37E96sSv/Ek/uSkeuDWLprfy+2ISnv9p+nm0qrzRfRRkvSMO+5
LwT9Cr2csWMOG8gTXrHv5twhGDh6C4qWwTDWPGMA26/+JsEODN7TTABz12CG7vHv
NSWxZ4OEYxebku2pFdnPDUp5aZ09IWEI5yQdG5Dzmj1aG6MZ2E1GvmngKSzPeFQu
6D7I/ABqhcUDWCkCcGJiXFek4nihTY+8Lz8v9Aod4C3wv7U/aNtIreEXe/j4gPN3
0EjpgZSE/KzQDAUUgFTfs82SiIQBj1xMiEUgla4sj4SLuzkM9gLHf20aXriUgcTO
RSxSankn6Q7d7M40o7vXGzSLHlUv+DTzISMbJdzBB3VxytxDh8d5XWhzA+CW2ovv
tcauSJQ7j179sdZhRPZXz4Kk6PsPs2MqrQzWskJxaC46Rx1Hw5fjkKptuosUqRtm
cYtz3zYSZYt8eabr9vyWXycUkezHnhdpWOaCKpqy2tg/xdIVUXD2+8LeYGruKSqi
IPwIwJiWZkBuNjPg9Hf0QqGtXsN6UCiCluqqLc1evk/NANwcn4jMkxeDMZPlmJuA
DXPK3ceMOAR+AYtNE4MkZ9xKTTXRTxyPOFRIaId9t4R5fFDthwiRS/lov7MKm+jj
jLgmKNlUEN5yoqReE8kdvkDneGw19DcNK+vXlKN6XJEofl+0CtTiabLCYXxVXKRh
ECj46ExYBLzwywUiAteK1pBVvEGuBT1808DA2hDhifyN+/keLVzRIYeQxbfx/Ux9
XzST4vbZvy9M+EHcZJNS8fG2EovWiX4zQ2/+SS0Op/UJaPKzPICtWhCOcTOF4bpi
b/bI5oB2PHkdCJgNMrJDW0TeccgLJfScyaZkvcaZGg2KuKZ/rTzORPQ22dNT8/7o
Xf98A0gQ/buBdodxJRamrMrcIEoaG+akU0H2j5E/UBTCI2zEs9o+WJxROpX1XbxI
85MHOp0u3DlMVZ/JXZCZVxU75gIqgt16Intb50buWAXilFC04NTEGtNzUYs50dpp
F1bQaOgaY+8UlMtg6ImMZU0hw7isC7XXyNul7Dg0P5n6e1v+ljY074JRY1Km7gFy
Yc/yxN6Yx3NYeP6clF9c9jVOO5vOL1q5J6OrcDxoFM/ClPGRWpxqmySafIHKXD7A
xjkyktKIOrtaKoESN+KxpVsAhJvdVUNln3DUFWfZlXFhZzaUhm4a93fASm/AxA2W
O4P80oB4J4Zg9xGnLQDPF+fCSdJAqtOubkOMvC8Tg+++r9mg2KG5Bvo1qFplXTkm
4PbRplBECAq+PFLFnIK3aWw+0KsW1CQV3ze2LYXpFHnN+DmRIrpR+F/wPaGCh/hM
R3EUeOpMmr8s30e7zOenW/KvpDMTUsF15GXBD66VyRL8iDtT+Grmv1U14C16b/k+
rktQ2bB1nULadACcGyRYVwidv/EtXR1ajmRSGVARgKbNWZMdOFA1+FZNfXE1ahCp
wsW8WCgP4NWlwu75749yEElagb5XYnkKdyXPTKm3/JtlluSoy5Mf5vEqr1uU4Kd+
JfkZZepnA3l8+VhDQjcwvXe2T6yRzVr4Ew/e71qGaXr2rdUQKlnOUG99INefOpdl
9TofjKnoKF2USfxZdkkRqZ7khZc5PdaRzJMEuqoqDbPH/3I06prstGIf5cajL8Q6
0YTC2rQRYlJXJqKWH7juPoG/Ona4Nm+01ZlsuAvUR25SVbB+hou4MOayUdcFn0Sc
RhG5bHhaBhhT8qeeoOcMJOK9VZJQ+iWaGjmG74vvG8rcrGPKbKn/aTbbV8hLp/RB
63WhtKiw21tZtaaN7bkXftUv2WGN3N+gfiHd9uLGK3GqdZfLglv9rqtg+pv231DK
zSTgDMc7IcCIzs4HScpBMknXc7to1Tb2iuHFtH+JMIfIfFMxU3YkXdtPQyHkVY3N
5vk4e3HzjoguJFDfgdntCbPdX8VvHAqTAY+FMaHlwqhWd6uQ49v8CnJk9FmHjc8q
9adxcFaNVhHbkMItCT7B2nTq49jwrEyrgFJ6NMSvrvBbd1PJufTiQyi9YxPL80je
AvS5Hkdgn+97mIsUA3MEJsml4xepY0q0XCu7wZ+Ermyaiy8u8LlCgz64FJy9oYt2
kh9Kyyhfs4EJXbCbK+Cgr6kERh3x/hZlxhKqW7j6Mt42WuTkvLf5JoqPVJnt6J82
jDXfcdCKcZk7wOUxdu4bIcBe54vjihjfhtDCA7u9zewpsJ9bTAkEO43XoZ08cbQN
z0V2PS9AjhRju67JLL9c40+JZwPXFa351vD/dkzy1wxRCrFyduXd50iHdYhTVGjX
jNeCHm114k6noKRu6N9qEZPaqOyDe/yctP1wgG5abHH1ZukOv3R/CrBULNEIHVE8
TIaZHJ7khm7mFMu/mnL3tH40yKZNlK6JqLxgMBkYsjxd9+q7MV3Xphh4DxHLkHnZ
8vWgfCeYCWFzblVX0hdT7y1gDrTxAm3p82Gshh3ujtf3ZGnoSHwFJiNaY0ma8KYM
+L6R2hNQWsshrMDEeh2K7+Gl5D0G83Kqj6mhYu83lwBiB8e2MsDV3UK9ihRr8pIF
XDAS8zZ9RdfpbCFw8GX5GUDdWIRM44kzHMV5GkL6wRqoAR4T/an9S3CveC9DiBB8
iBQB4bqwrJP2uxAmTCoFUqezC58w6elNleHNz39kKQYErXUmN5W8l24bkPG6VqaX
RgjTkO0fr9W3sAxtj5ca/v1xkqUlwPKVPFKmhc/zFsleq8w+VyHCZJdyqbanbkbR
fdmnHVMKNrzs1wpLkyj9ot8xYgf2uFde/5sLifuOXUzqMvzZhxue038Nt20fjaJt
z6W81kMdNdsSxqe33s2rd3G3iz4mKGWAggpGqZEW53jjHbIBXPBwYhE844OF/Lkb
Yg5WGgW8GLTFDgdXgxdAxEQbO2ocl4ueE/PecT2x1aOWnsKbzpovJjC/CSBUs5Az
s4UKGr28ox1wQpPm6fBY31WVnfe7h3yQ2UZEEh1FZQliMR8LwxWabjf2yQjCVwQm
3OICXVHEGLdtcXy2EWSdFxitV3S0YHFeDLQ8f9cAc+bqh61ibeKa0myfDAScax+t
q8Bh8du1tvoVk/4Gwm5ulNfkWrtYtbjxblgrGroieeCt3eczOZBqMKSodfLqOJNq
MOJOT3vUzVJZ6Ign2Ksel4EJmIf32w3msrMWbrsXGQhbXEfnfyNHjZQ1G+yhAiXL
uWqbdOFzPdLqfiuv4ibu2+QD0VkKTm76hDeJZJUDZlIBUTaB6yMzMhsupVicBkgm
9EZlgdIqEoDX6HyvMYCxC4wTIxF+bAP27Uq7lBqhyjCfAFFfS1QRPp0V1H02yEgt
JY6dx1F9uznUT4/TZR0tb9uJ3nIWXmrs6OTFlRpS+jP/pdf+8HDKnhdzJRYu1Es2
RNpT3rdwL9tWGoSoCfZ2ch69zmxTzZHxRlmVrHuoavWAK55b8S2bCS51up2IAVD4
OZLPhuz0wYRJjqdeNxK59jd72xLKuNfWqbOJpR+ylxK+TlV0Ss95S9ZKhUTHvjfZ
5HlA1Np7ToIRjmQJvvhfs8MfijmjEF3CBG+kTMDnFlN7IFV0pmv0GcT1bGmczBcG
HVp2alaWZPYHJl7QtCmQI7tCwYNnjkFV+BD6RTwJ3fuIkh7FYfcIXlD/lEbdo+/W
vEWeSeu+X7rux+QGNyR48Ywwx2ApYkgcVNfof3nBcGR8ImYUagvo4b4f5mhX4kl3
ATr1CrRvUK+HW2Kp2fdUxzT8DU8OpIHIo1Jt8u//I0Hok+Px9oa24c0eLL5xFnDf
TrWSHWXGrrw2uBznKWdNGcAIDz0tu63VhNEKJcsDBg6PiZdK3W4gKPHat7qVCEol
Zwo111q2c0PgFMwHBvhrvK6yrQhA4qm2W7SQSjRqR3oyPyCTTKeUJ5fD834sxvT2
sMvnG0H1SFOLcOfZiyl3Q103XIe4U5hYcxSQ+tvoxR6odciGTTT9RL3sqC71cR0d
kbz1Xnf1KQy8C5rl03h3Zp9BnMJ7qsPA2G6iLQkwzdcozy08/+YMbQ6d4Y9I1GYY
HhZDNEFF96dMdqEXu4m6JilQVyV2NZtzKpvwCnBBZ2GvVq9w1oaeBUw/5JmYwkRp
jnXz7h5aG0FNPO6S7mRa5aU8ISLkTJJn/1juo5/VB7CdX3T8Ke1lBfU0/Q7MZVeu
zB8ppXceYC08O0yX/DFMReScKulv0iEZdVpG9Oi6UPV6J9/SM2lHrqVaaavWZrQ0
vE2r+h3Ar8+UEM/nofbSbZrs2U4G+7EOOpXpBCm8pSrDS+fW9Jqb6SADczSmk8g3
jXIxIHt8POfv6f8GID1+bUoibOIPDmimkfyGLC9Q6smouK/z3PA1xmy9kjnhUrTo
5nK7bmpIGjwF2UgW9yepMHznW/XpeOyNGGSvpmj5fQVfN9YQV9nF0xEsB2RAPmds
xl/H+I+OA4WYIftfqkcZc5pPfVa7tcsunrTveg3lGbsmoJ69CvDK+QlRRB6APsa1
11xyLCWHzXjhQ1q27eBZTCl+3IAbpvvW6liXadQdqVBj3j4nyf/gz+Pxl9w55B7K
vBkR69rCQZhtNJ8MR3KhPDb6eakDiEkpazDxk4lEk8EsxoVTvvkqANlT2kk2bAiX
FstfKMQ6p+9J5sGcD8Vc9PxlPU/bkSn9j/TvWKWFKaE0oxI2upzeb9wY5s9PxEMZ
wBQLD0pCFevTxme5CIF66Wjw30epDRnhSFfsTu6sQChSx6glyxyBH2bIc6GKbKTp
P5Z6yDUJCwO47UXUsOPKd8IQv8xQP6WmvkwPt1fPvQeVBAldt+eKgkJIdWdsb2Y2
1fFAOeHegfnUzhWTxwmx6o45R0g5s9sJN2Kip5EVPmZZQ2Z/WGOtqOWzEb6afcza
ABYOMoqrfLfXdNOWp+j7E0dfPDl06P/HE7ZIxZYnJyywkG/UP7r6/fB4Ct0xNa3K
DbPWS+luu2Pg0lqkdYWzd6MMuuUjP1q8pdxD2wQpZPFdIReTVPlnagFvcn1Z7aYC
8Yyg01P33yT5Gm+P8c+y57Hqfcm8AwgG8fUzBnaSTodE0gTOQl9GaiETzhL/ICxj
FajkAZzEdXlOSq1vNIzJRLNnbumf5dhRl578aV/WX+4Gmw0N05JEVScmgqF078fZ
noHDp30oOVdxtQsgi7nsk9IAn65/VGU1cIBQBqyBdEHWh3XvG6WrtSU09h+IHP5d
nEWibJNWtHCoIZoYPihDNRQkphE3ZV19h/nyyBYYad+pU7r8d4+cE2wg7RUTD31y
fbmzFL64m/1SiHJsl71UeRWGosBIKCgeBgO5CWliwdcZeJIE5PexJl/4yHNIeb0j
dcsdWR5m/ik9E6KxtLMfNbY8fnB1Ons5beA7hMl4LyhL7bGNPNxxHybTIkJOFv4m
91insTjWIGX07cUTPmz/Vi3Ukqo+phf6Cj/qtWZ7wGGPyClFdBnMnipzLOjBRxbM
b+vE2QiE5YOpknMme0DlyuPDFlJwVt0Ds+zHcgEgzfnCoQw9ev4NMroDJ7cCWaPp
0Pwn2mcuSUqxgMX4xuw3qcyjVHNOWNs0FALjgAxEmh11n9kiISNdYiH3s99At4nE
470PMBx97viTtRwj2jpxEg/Vl1KESY8b/k+QmzKTvaId6TLhPyMFhMyH1dl0C/Q8
oyHoverAf+yxPxhJKEmJRWdvfiufrX3HUkVJWIawdTmZJj9pFL24OVnCIefI6UQC
ei6Inm/sRC4IRgEio0oFPTl/saft0ouZsTaUOl3ccuUStd4haFq6PIWBOqFrsT0U
fHeKbyc9QH+SOLMtoSqoofHeAWxw4BwdMbA4uOh5jhTxTGzVuIumE5oe48qvGWb8
f4LRp2PvW8iXdq9w567ZR8bBmL3QQkFOG90QA/+nxrdW+a/Pgdr1TAandmOMFkhg
SOvoN9Yi7H8BBgtSAOduRDA1E6GldjrW4c8Yl3PzFwj2utdN4+oQ22rXhLuAlCYy
LxHSctWaV7m8tRJhr4LS8EpeiaSnLeDG1npmSlhINvXXtCHuSTqJl/MjUeJXBvKE
kC2P0lhKFcCxwon13yHr2F5mLnfmETY0D07aHa20KK4K1Kt7C4oQKIcm3yUQqdTF
dex1aDSx3APX2bVcilt58F8JYdm/SdVd8cF68tmy6GCA7Im0fVs8fKC9cJz4NetM
NEX5SaKoqcppqSlQ1oNO152BnEQGl7gdRaRRFGeLxC9/aIZOHMXSkVaH58F8FIeh
hVBGhpHsHdK4tgXDDgQhFOH3G/KZ7yhr/NswDtHhFTYKPfeKfzngwgIL71Hi0Uu1
0Hw6NobJc4bwgKNm4jtuI2cCb69v9dH14p4DiqHtBuS/UA+bQvQKybmloQt7MflJ
qmpAIxI+fpm5pkvsjn6E2pogwI2cEBx6LzpT0/EJi/S6xcqxuSLhALBdCTvnX5Mx
reZDep8YWaM/lGqqHp+3B7eRUIp+Sqc3T1VducTUPypt9nBY8MC4TWtd4ZwsC1Ux
0d18NvNiVibHR4d1rOP+DSESeJiehAPWufB9KVtHTiD8TbWez7WBQTjmxJokmzQH
ezd3Rj6pWNy+UvzyoZmYFnYMyDSoW9gvXkBmtgUZNk93UGkVUR8i6ypD7CPIfIFW
LLY5E+4keLD2yXQ7DTSy4gVDWybWPea+EPdAKukNU0+/3e4GyuVw/zn9zVL77ejs
Zv34AI3UPuTITIjJZajpbjzSyTq8awwA+Rq1PRbpYO3MvGC6erciTrIp0HLFctyb
/ZHk3kHZBkdKBqnvE0EYcN6OG2E54zmF1sMBkUyENkywxVbbU1Y0yVCAR8+iUFHe
rsNLTo9y9qT1JVMJPchHulZLa4VMC/JNttQt6vvlSZIkFzC2pIXmKwFkvPR1Y/I4
CpQf7cjFUcwfXPc5xqHrPmf4CXzKngFLVSOsEZ+8kwnBQ4zPyP2Fp9bVo5LUTxek
A5RzZYv6AN4qVFV9V8/DZTevTxf+BhbSQXE+aJYFKIyzwJwli3Pfc4UtLMqPZ/9X
RwgKB8nkzAIULLrymd4+nnDRJIvzRIpXjp3UGRj5alk7Q2Xvxfz2gFe8kxKi4LvS
EETCm9Y9W83orxDsh+9kCcBONz+KMem30YrrkGFZpD35BEVln7lL8anPzQbopbbl
3nlgY00w/EdYCyRMDxvbwN2RFgAcIzHCeUEnt4FRmKc0yVrbzI+Wtjtx0Zf4C4MR
dJZeU4Gax5RcvqToWQw0VRi98uCPfeMlNvJJsjdqoQ/COOfxr/+/uK0KlHXMtiKf
PXRwok65oUaiMfdyLNjOozZwH/JXBGS2tTkbJtgS2W4HAuZLhxhaKenx3eefGx2T
vZOxfNlj3x96GyYKjKZZcGKefmnfw5iEy7MTE9ukPlekjgW3hZUDowzToowtgfNY
a1OwibrGGElNrMt8z0bBd/8q6NZwEfG/vSBldup08AJMbrJ6bUEhB8cQe8MOVcFE
jiPrfiDasUzxPkG2h00n6XkwUkCGvYH6tHkY84cOpnShFPoV2Pj/FC5MGjwHJTUr
FYV/S3IwFdBlT5RSftaZnWo/hW9+uT1m/RjOI6x1VuP24Kf+edxNxS9UKsLR9ROb
3DKBT3X64QHlGKImGV8eCmFV7uErIsMreQsIfa+sHBDXL+vSt0hYHvrXeqIBqfdT
HPKKesrkkyV+1t2VPsE61ZSUz3v+Klsqt9zzxcdt9OYnus8TpVXmcC2x/4tN5AKo
/GUCqttQtUOOV+Vif0J4/J2m7vD7G48ZdMOKQww2G87rXUtOpJ/MlSYyeVWLS1DA
DhV+WvAw4D674JhEuttX/1ScsH9EpdMlar01u2rcUcQY6EhubwUr1UsA3xzxT0RW
gg3RKs1453P4Ga6pD0/QE+WR02Xrs1AnatxfZT3Mp5pDahHvK+hOvcbF8GLkWW8h
ldVOat/KRNo7abw5OWHCltUTbSsZyjcTUZ/+B+3/kRECpuPPPaumXsXJ8rNGkwis
E6/05jE+KIWZ/QNnJWdDM2bIqtEtAM/co36Ao+pl4hfniZSpXn/5w+A/88Vj7q0S
YVicOJNcGTKbS2Iycjj4V/dxo9clsnxA2D/P65e4MUukCM5k7WBKv6O2cPosWKyb
xxTqnzLUjJ9V66V8djv9TXfcxrPTy2JV1eVwD+rYg8ixa9REPcgIlZmBNy3EaACs
7jetPshHkU8h977I17z+sCo5jUK5Bf0SxuiF15O1/gzgYSczytwvLrsdqgYdrtM1
yyCa20VvrTSChjm5LRhKu3bxdQI0PI61qFPrQ71T9Joe9W99o4NaCGPuVPiMr5d3
BQpXdbj1srxImMsX/wUFPKvkLLgWbBJwV3xKz+MWgGw4VsYHM/Wk3Gd5cxrc2ysn
svpxrfX/PMM25p4t5rbBI4C3LTS0p8X13I9//a9oyQH2U1lwpunT9NxjQD8bpoi4
t2A4lKO6m6L+uBoZ6XyhJQ7kOiLwnbs3f9JS0gu/AgYOxvUKE31KtTq2bXUXx2j6
GmOxdrj00MddfO7hgNGftlE8Fx/FLuz/q27LyXQ3NqYxxYqR7Rjr2aBzmDpmuAi2
lkcpxjP3i3I/DyyBkcTx7gCtOYA1MXUh+ZKC6u6xI4r0bFxWT9RLwqaddGf9qRwg
uGUZBp6DExQlNUCe7mwzqTgc5Wzalo0dzY9/7CY2c2hEV1SHZioM4RfS1wRUrzYG
Dfqg/rreK3kJXIGqgMbCNJ73zltlZoAsotxWV2xD/t9Y5rta8BUV3gGlsHjB4gdp
bo+wWIUReKeJ0k8Tqgxbo2wEqycyfPLVAMXVxzi4xC9IzVdzy7f05A4+Bq2kXncX
RKyHFeLvYFYCR9pDUpCn53AcV4rr1RYhh2KVCpNi17dZQK1sxR3rbxq+gJEhtvy4
dFfCFjGdy9u5WoUUk2MWzhto1BbsK2rtigr3KFHpnAUcu50g6dNxZ540eMea8eZx
yN1YiczgT1H2Iq2VDXcXqinOvzfsmCWWwHAOtP1r8SJXV4SvKvDCxxhGF/zVWqdq
Mx8FjivcZJp/bFmIf9nMaJFM2zMzy5ev6gcNZ7ggzBk=
`pragma protect end_protected
