��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,VI�0=�E����pbT6o�!�R���#�&��ډ��)R����ǁ�7����s6��3�o���
dk��2+;���ƭ(�;B��iUn������DX*AM�U���{��S�� ��Dd�F%�r���֍͍E�s��h�3�.��Oc�����g}h^9�d�c�#�iS�ϺD*�-���m��h&���Z|6��{4N�CN��ŕ\D�!X���e�L|~��*�1Hh��Е�[?j��&�ʩC�.���n�<�b�٣*�4�ފX�g����4.�e�;,FD��f���1r�f�	U$	�c$�~d�1�PV�넾���=(�>�?߹ �7Q�[W�|�c'�(�{Cm.�����E]:Q���U<��î��:���[
,ɐ���^��9Ǟ���+�Y�϶GH�O�ws+{=��?���|�����3�V��:�};�N�a�[?`9�9ϱ×Z�n�:@�94�ZP��ގg���k���V�t�52�V���m#CJ�fG�z��T?c��{-�<y�<�m���2��fi��K��n!!y��_��Y:���f[����7�o�_�≁+��!q�<�~��gÛwd��]�|4��6u(a�rO�tX|��b.���}>_PL�ɵ*TAX�K�5&�����'�B[�B-k2ٰ%ԂY�P��� ���:4QH���^���{��zD�0(u|����d���'�/�����1W�cq���$e���j�c��N���!\��M}�ދ�B5�'xX���b�@�D���|�I�4��e��2���U���o�0��S�eVU��^�q"�ݩB�CGH�X��3���٦��'�M�"dX�T�@r0�b�Aؖu��$�g�><m3v$� $c#�'�� {0�Ũ퀚.�CG�3�h%�("d'a~�M�\堹�QѮwonfĺ��baQi�\�l�n�'��:�a*��Y>3ױ�M��&i�av_B`{j��5��CXc��F��������������t%�+~��	'�5w/��|����m�������i`�,������?�	�y�HJq��xX�߀B!0���k�χ�<m���j,�&��K�O9��g�T���fV�Nϐ�?ً��<�a�u����}������
kHA�G��-��ʢ����󜳣)���Pѹfޥ�v(����Z.ѕ��{�ĝk<�]�NQ	�|� �4��AH��}
�NulӠ��`���aߩ�6�,b��-?�%�ʘ֝��5E�n���J^�0ʽj�GH8��Ѩ���'�+z�|�z���U(��t��a��Vs���(�p��"����'���#�����Ȯ�x��&j0�r��8�; �ۘ%V��%��3��h
yc��c�3�rQ�w{Tp����J�E}�\"�.I./��i6��r�݋��ªqvJ��1b�%=�`�K.�n����d�
�Z[�j �L�*k�i���7�N��U��u�E`m:��S	�3�ˌFp1W	�|Ǯ�d<��<�Ȼ�p�q���D�ʥ���DgQ�v�\yh7� _�k�v <&�i�IYh�s��_8?
�ecDX��=�R{�&J�7�2�I��W�\�ĉ7M�ω�����j�g���"�d��������0��X6y�������BVH]�;e�i�/z��Hl^*��A$Z��UP~�H��+�s���C*�[i�d�(��)cO>��5����]3��~��q�.�Ҟ��eN�݅W=� ��[��|�L�u��[�7�Mo�����5k��,�{bQ�_i����_�2z�h��Ny��pD�;�ڜ������ӷ�2��.҄N�rf��MW�����T�}�2v�a��k��f#�n��� ׃se<��f�9��k��u���e�V�.
B���%��iPdD�����