��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{�J	�'=����5I��gرX���|���UK�xT��5g�Ul{̉��� `�Ƿ�V���H#���;��as�������N��!9٨�`��l�����BJmt�l%��
��[���j��]B����ԡF{8�ȍ#4X�З����z�j��q7�I[�����^s�T�]q��7�Iq~e�������*X 5��$Z@a�6ր'�!pZD*e�@���D���@t"��=-�p��A�WM��t�d�F/���CQ�CH��-���FOӕ뼘�T�?Xf3v5-�l0o�5���υ�v:��Pp+�8%c�������3k���ǌ��=r��ձ���jJ�oMй��s	ǜ�B\��,�!�[V��_�gv�]f`�WE�����X]i?k���D>��P��ћ̣J�����������Nz�D��3�p�m�.p���YH^����g;|?	�ps^g�jݽ%<��s�=���H"8��Tw0?����>i��I_2q[Ys�1�V:=�(Bu}�㟷.���Wl��G:O�`���Ȳ��q�uFQ���ă�[<�B��`��VP�'���[~�^���<	��}�*}��0�Isb�n��{�|D��I�/�N���O ��5�,��&Y���K����8a�`^#<���>���_�G7L�-�]5޼�����q#Ns��z>>"a�q�MZ1�|�(�!�nޱ��e�_�DBAp+۵���
M�:�k������o��^���RY���N����8E���k���U���%3���0kx��Tw\���;m�Fd���-���6���	�ɳ���(W�\.�	mݛ�	ԯғ�d���-?cn
E��]��c'*#ҦP�U�0d��~�)������۶)S�:R�(����1��U�l;/Xa�0�M1��0�@f�i�A�-��7�J��T�k�S��_�{�J4X�+�%!KX�y�l� y�:�9��â����
N驮�� �ٙ�����؜�g[<o,/������3�A<�Z4q��~��i���Kk�֔n�}Y7���&�Q����΃,��jF��5��C���fQ��Z���^����#�_�t��8����-{q�
<@ 6�l�Ʋ'��J��/꯳��2U����rӷ���O���z;��.	R�b�	_|�".��Mk�fm��E9��.��t0'(���r�-�#���P�� �X :����[�5�|2���mw
<���	�b}!��JC�R�9.5�� �SI5�4��6��p�<�HOm�.w�h]5�yᒡ���;1��/s�Z��-�ՠ�nM��즴��1PM����]Rf�����l�uC?������,�Nw��}U����$�f�9�T�/���RP`�&�i*D5�)�>!�c��ُ�޵�ika�NK��&>ۉ�</nW,�	��ۆ#X'8� D��b�hd��UU}��U�NaI�N�LJLCu����-��7S�_��"ZP�f�*5�z�zZ]c<�nW_�ע��I�Z����S�=eN� ��8I�\*L�`c�����0{K@�ӵ�=�;�B���_��֛���BIR����i��l_�q��I?2��F@J]�* ;����0`0t۲���9C��^�CJ��*�48<�$dO�XI/5�Uq�b�G��\]��x]�S+�j..K�E�X)}��ҡ��(v}h��{� jB��6(�UN��s�Vta��������"L0�Y�g�w��]	}������dl��i7��2��E�>3�yV���-_��Om��Η������D� �B���yk��(I�w��pE���!�	�,+��u˨�#܋H�{�9&�s��~�FQ��&~;���_�Ph�|�9=i����Q+7�@I��j��7�D�e3��?�`��޵��+���ƕ���/�f��Ǧ�ځc���/M?L�c�7q+TY��R�J�^��v���w܀�b�YP �;�'�p��:���z����A��ێ�'nO(YՎŔڑ?6�q����Ld�*Km���5�[�vF!�Bm9�)(c�r5���#o�A���.�B������}V���%�*���Ś� �:�@wB��~�9��\A|��.0��1d>'R ���$�!���^q^駡C�0����i&k +֯�۲O��b�T�������-�6�D��TH�D������m�G	k�*�nAKv�F�%#�i�Ac���|��r����F�M�s�H��K�hDvb�HZ�������e���"��1�iن��i,���`�c���}q��In);p��;�/x��⼔�`���z�vq�܇X��|�,U�Oz�r�/6�ʧO��c�������HW��J3a��@��KF��A�����&�A���k(K cIJk[ľ������G,�Ԏ����D9BJ����t��b 1Z��y��W|@�~K@M���A�K�	��A����Bz�������{��.$�Ӡ.��y���@7�˯:q������{g�,%��GC�.��p�E����Hb��wН���J�@q��n��KW�~�E���1�������_�k1����ٕ��:�վ�śm������௻�J ,H��6����Չ�Ԭ�
�7+�$\��~ ��
�]yq���oY���`#��̸��6�l�"��Ki������4k�r�