��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�p3t`�Q�|.@��Y�������i��<b$�����)m��x�2�2g�<���w��c�`rlW�X��p�tG�iY�#�iW׸I�5]Ś�d�gDG���j�c�r��"�4�zj��iw�ݝ��:esK����a��GO4v���/��G��˔���d�������>��݂��C������0�G00����<}�#�k�=W��R���T�u���ǋ�1%�(0`��p��/&���� 9-��.Vu����̖fN���W3%C�宾m����+�5�M2a#b|�aD9�Gh_�q�J���o��%U�31%��C�J�Y�?o��2�X6�̙X��L�o���ej���+�����b�/Y����y�'�B���ğ�PU�RJ��ߕ@Bg!K��5.C�kPK��j���6��3�oVϯ�>7�dw�Y��y�m���`�B&Z�%�v[��^Y�^1	 ���V�=~�%K���O0(�{�#�z��`���9+E>0�����%���ѴH6/l�~>'��hUx6`���Ig"��}5JRT��O@��^?�V�Vy/�&��}���B�Ir��8�T�O0��אf?�n�8HyM"S�)��A����bu�C�R%Βyt;��᪨���a�(���������b�Q�HL�� ����Gy�G�a�2ZE����6���9��LC�M�j�6�e�����lJ=K��Y9Zecc��Ϻ;�Fj���8�~8�:�Y&F!�����=��b�r
��E��#)��m��cX�{1Ms���DW�K���k{��[����LD���N%/�@��)�MpרsS
��L��S�p���D�1�.a��J� �Or��|���[�z�#X�X��F��ڝ��C��^ω/��M��_F�C �l��(�t�q���%1\��9�]Q�~������Y�JH��f�M7���<!-�c�����S�`%��@�F����'A���2\�A�/Һ$ފg�bD�ק��m�*�<.�K�=�礻9��y�`*q;�)�97U��C���p	�^���t� ��Y�a���j��G%�Z���%s"�hqB����^��9�:��hk�T`��!���B G�4�-6&�����gwʝ�F5�6��� �Hl�U��uf���p�zWa��FW���b�`C\a�)BL�8����6�P�=�r���-<��4�4��m�����T4�Y�4+1�	�����\��'�����:���_�u��~(vV­*0�^��IA�Z1�k�&PA�5��g>/#�7��9I8��i�hg��4��@ͯܶ���مy�GȮF�R7��~J�Ii�ߓBR_P��Wa�c��oR![���6R��X�6^�Y���\2�Iށd*D�VP'a3�-5o�"V�ѓ���yl����/��UW�������ƽv�R���Ɋ�� ��t��� �x���6g�?zZ��=۱
i����}Ն?�'ǉ����t׸�c����f %�6j�Ve��CS0ŵ`�'D�5ю�c��Wx�`V��տ#��~�)n�`����G<(�*�:��GA-<�׈F��e�0Nğ%�s738�M\�oa�r�0j�a���S��1j���2A�P�=���$�Y"�$:�)�-�W�{��gf���)���
DX�4�0a֪(�@U�U[�Z��-I�J�ف�l�zl����:�~�^³YL`v��< �uk2�T����+7�H�85�+�S��u�W�Ya���a�[�]�#)2`L����R`u��/���"N�h�,��/r����6�_"R���x��!�T�_y�d�~�y-��JC%�S�u�V"��@F�v�
zj݀�[R�X�k���3���V���<H���E�J��hH5.���3#�Y-��"��G ����~3��|�}'PO�5��_���K��kdg'�Zz�.�	I%�c�?,�O�.���ΓvD�
ղ9�>�S���z��8����#M[ji��h�"����[
�bN����upg6�|d,4�-X!
�ޘ/!�=$
���L�7AD��I�:�Pa��k�����Ǒ��G�{��ʫW�&�$��@ʐ(b.��r8����L��0s�� S�ͷ�-��-��j��������@d�%�o��O��.�~5�A].o,�;��Yp�s����S�{[�9�ї��ܠe��\1��S�O��~56��$#�f�h���ACF�ܦ�I�c�2Cl��n��!F��b�Q���P)n����=��k�)zB�9��>�_r���~0���,�ņ6.P?�sVvZ��u�k�<G0�G~s �D�����D�c��/Jw�������F����d��k�>U���q�Rw�J��M�R���aYWT
1��ՠ~���&2��x�#H�nhr�D��|���ݧ����*�t{��"ڸ.�k�)�t.������@�����m6'����8PN�F+��}#�����J�B�=W�ieq�'��5�k]Hʐp���d22�~��@��x�R�d�VXPK�U<d;W��q�ȍk����h����'�+vF3�,�"�@��k�֢H���GZ����@ZE�?.��P�4�Tà1�%�E%��=/Xb(�!�iԲ6p�E5]J)�Z|4�jc,1�p�
ւd���
�_�I��Quñ�����_	��2 |)�HS*�gh{/\�j4v� ��U�}?��i1I�e�a����^��<no�6����F���#t�.����=�(������A��@��,�N�1g�Z�F�V& �'5[-f=
a����c�$�1�r�^��"���#�F[��=4C'�#��~J���({[4�jT���1�����H�O���)� ��<�}�;~N����g��YUk	!jUqv�9<{ϒlB$׹���덟I�(�1�䞬�L�mؘne��Ą<8�W'\���tv03b�,���tŵ�&ڻO����^�N�F�w
!�0E��'������^e�	꼸�|$�� �D���Kz�O��T�.���w��Zw��;A���u���嗍o4��\�㕚B[ެK�LA=gN�Dy���X�v2n��oŖl/��ۓU#�u����5˒g�>�����}g�i�U��\?��ô�K=mS��Ϝ�l�+��|U���^��72�H�=fc���⭧	u�P�%D���i���(��ఔS�LE�N�..�����������X�C�49G(�R�:�2��b� b�zX��
�O,��}G(��D$�J�13E֌<2�(�"g��͘G��Pw������X>��Ρ@���@}I�B������|��D�4�O�C0O&�F��Il����l��437��q�;
��) �Y�G�f'�sa�ޒ�XeM�8�䁳ӅQM���������q�����7rZ���?	�ٙ5�nr��j��y��*��֜�����������De�2��{���d
���X���l���4���@aX!eq�L��.K��Ȑ-�'$U >JTՀLVِ��gV8���y���5-TzN&�n�~4vM
��ϓ'R_��=c6z�H�u��OpPnV��k����w�ڒH`��B>(@���0"X���A�����R�3�3��U�
ҏ>�n�Z˕s�ʴ���m�%����	Ak��H�P�SH���뭎��gv\�5J��J�"�xX�˕��-@2;�Gÿ�2������joX$)}dvֽ�P�M�<!Iu�B��6���w��ŝ���K�X�-KX>�A[hCSk<9���J��B~���%o ^v�!w\���%�4��1V'/�`�Y,���#�Y��~F���tM�~y=��.����]OT+�>�_a&�Q�f�:���T��|J�D5z�t�I�If���Z���fY��z7�ybN�]=��Ӯ�n�i�Nď�e�Ś�ص?n�U���O*���o[?�{6�{���o(ID����+��|��a,ײ��H�ѐb��;A3
$�����W��QC����j��4x�W�YLHZ�:����r��y0�6����m~��E|�-��
�8��,�L�3+��Pi�|v��ػoV�(�[��9 rFx�������oE��F�{W�Ui`���� >it("�e�rN#Ѓ��]�Yf �V�ر��U\��|�џ�129�躪7V����$�Y%)��Κ��݈#�����{���'ޕ�؆�|ۚM��г�򐡥���,��d�4�6��U�ݰ�������.�
�}Z�ߨ:?ed/�Ŕ�G�Ǘ�+�\��8_z�'�	7~��}�yN�X�w�T��Ѩ q�sUW$��%�����=���S���`������]y2C��h��o�p�b4�L��#�C��Ax����J�g#�U�2JiK%˅,��}�4`��X���������2���>� em6|���i��eh�(���|����"n������	Lub��%4m�/�L�����Ь!b�����9�@�+�U�E�B�&�o�[��}c��<M/G�OG�ƩF�=��]3��Ӻҡ�!�+��;�
�qަq�^:�(x���ԁ%1�>c�pfqz�x�k��!���Fpt��f`�+q>��`l��=�+B	�����Ԅ'��
]���ã1�����(���O�N��jئ�_b����'����ϖ����������;�Q��CY�@4p�J�b�����m�n@f��8N��C�:�1��N`��j�6X���#���:�@r�T�/�sj��3'�T��oz%�Q�<�oDP�0��%-��$�ݫn�_{�ߴ�&�{& �!��3RN��ϩJ�����C�hAw�鞅�����/���}�k5��U�:S���8eM����	���Ђ�Ö�,i�0����y�cf��'���OCqU�%D`➂&;�Re�ZZ��~m�m�Y���GKRLE��=��jDvf����|?�VKʪ�Ћ񹵇,Oֆ�F�jt�l�,,2E�y�k�!y�m�y�\�Tu���:��1E��_�Z�+R���g7�apP���M;h5|2&�uT(�6�����t��k ��T5YKZ��-A��k�aW��a�?E��dww�Nl�QPA�bTq�tm��(b���lǳ!�c�HH��-<:1R-a��ǓӺ(~aC
5;L$���L)����4�}s��O!f�!��8��k]j��9��k������j{��FUИ�D2��� u�3L���&91��ԃZIB�����z���̷M>H!9i���|-4�O3��?�Z����'vF+����U����J�Ա��#,*���Y	\��#N&��߀"����e������p��J ��"��SJ��V��/��:��\�P��r�|&�j�5Ue��/i_�b�@K[��J�x�?+O�.�2�������{F�9i@`��U������C��Ut�������b��_��E&�a�ɣ�(�M�C~4*��eG�t@�p3TDr�4y��-���?!���~K����Nyν���}�<a �cM2�ػ�~r "$h7������N?��440P��l����'~��J���Z39�Pތ��d\4� +�N�{^�����G���t,�m{%ޫ�=��ܭ"=f�/�y����jZ�g�`�D�$��{P\H������W��@��"ٟ��Z{N!���k�)�S>L���j�lE0�S`zr*�
a���|j0��6bo4r8p>[���������	,��^��KW>V�IjY/�B_����ɍ�$]|�h�J��m���Whq�
}��Y�E��,=�I�l�QQn=��I��2�(t}��zN/Ex123�7��Sp]���@،���O���?&��\���V����#kҊq�W24*9������-�(s]�	�p���c��_����f*R0�g�Y���_�X�ZR�bp(��;N��,���B?��f0Z뚏���F���7-h���n����8heF.�FvmVu\�Y�}5&�d��7Zoq�`�/Z�`L%s홬&�q���Q��8O�*�w�����g��0��F<�d$�j�{�2��3ej��ڼ 'q��k�'�r��{醹K(��XM8c,"�:Dmg�J!D�K�^�PL�ur�H�W���'&U'࿡�Ҧ���0r����ԝx��G�E������h���&<|PH��b�Lm� *L�F:�
��g��v�{�cb .�ə�5��iu�����+��P˪��y痩�����h�؞hm�UE b��M?KL�#�b��C锒�� ?�:��i�)���J�������wG@���T_^��t��`���U9�jm���Pg��H�=��a&%[�@��\���^B�!\Goe����,s2��.�u~݊�,l�����_�*Q�`��.*Vf	-�����whM0T;K,��Q�A�A0W=B�O=PL@hv�),B��ʤ3µ�`%�I6wW���x�m���BE��8�c�.�_�R}� ����}Ō�<qg�o��B�8�>�������~$B$Ћ
���*��s0h��&P��Z�u�Ǡ"!�mQ����M#Y��o��0���=A����P>_n��C�L��06�)��T�G9�;R��9bP'��f(c4cvN�F5o����"Y��F�����.��_V�:B L�_�Scm����� V�iȼr@��7"ag����#�9m$`-*�������@'���S��f����eH��3�}	�J�Z��i�:�ZM�E���������D>lJ~�.�FS�y�6oE�aͦMM�~�X�w�j��Xڶ?E(r��[h�O|��G��/��ҐD���'��(=!ab���,`�_z��<��w���^F�	I$HN3�˱�_�0���	H'�}�k��i��*�.�N��Dh���Gc���ϑ ���Z��'�%�܌�`�����!��l��]���f���D����@n�i�_4QDȯ~�1ffb�:�W�{�?J���w/�4^1v#��*�V����_$�4p��^�͊^D�{��$e�6��]@襖�U�8�W;�F<�.᤟<*�[Q[�!��p���~:��E��愰����(��[P����`7��k-7�r���O��ON�����=�"��I����^\��<d�[p���sp�6�M�2��x|A����>�e)͘-gԀ4S/�i��g�u��Q�����pC����eC�m�5���1B&׀�X�K��������^���}�Y+L �����,�U�P��މ|>�>@m+g#rVz��]0'��k�P�����~c $;��Mι���I�l|ƹ`������B�����Y�KM�܇�&
�~7v���3�̺\HX8��D���@L$�'fF���j�.���EB;�=��m;>5
1/\Vi�L���|��:k�gv1��,���»��P̐~���~���Gq�cF>{���Y5�(q�K]���Wv��wy�GiZO�<jq�Q-��Y�����PE�Lu:��
��%�b� 
ԩ	\�p�F6��W>��r����6�Q���`��)��L(e�P��ϥn�Oe�� ������9�rl8��G/g�Ҹ�Jfe��Ţ�K'�����'�:���eRV���grk�P���C��>�g ,0�Hr��{w�cy��rty6�Y$iL��s��	��X�D�}���G�_�u 
Й������چ�u�%Q���+q��8�F��&�W"u�&)Ֆa'��F�ٞ�T-b"�N��Q*{� &2�E�v;�,������,����3c7x�����wA��jق9��d5��aM���w���!�$�M���H���0�X��fO~亃�٫|.�{��`�,8����O�.xZ��c%U��	]�@NMu��r�	#�>������{h1��o|��J�d{I�j;��NL�����v)N ��0��{�@��K�a�#�����?��vr�5���,��t��m��&�]UI=�oR�8�����F�;��]��y�yb�+^4��s�#��^5a7���C@����v��Wi�F� 㸨�SokMQ����l[q��̳#�P�����˙����} ���u�� (j�"ʾ��e�(q����2�;��Kޤ^��C�����X!���"���a��Z�U�8LSduu�!�$�		?�~0��C�~��i�v������H̋�\�w��[��ƪ;D���t�h�a7���)&�F$ēQ�dJ'���&JH��e_�_v|!�2�q��Ӷ@¨�Z��x!aS���������7)�=c֜���7 �\/����q]y{w'�'k~��Y
�\��;��S.�TћWtT�n;k5䱥�&M�4���uĶGfp:�#��(V����PoJ��W����Mj|�(���s��hv'q��V��ȧ�_1��e	�7�w���N�E��g���類U>ew�y7@�&q�34a�o�ֳ�P#�����_ؑN���i�cu��Lg��39V���{�a7=^s�<�� @?�ЫY n��sJ���;���n:A?���R�J�O���,"	eJ:���d4�ݜ��WlT7	3񔑔ұb� ��+:S�|} n����������(� �o� ,:A��\E:�������^V���<���}����3�b'C��&FF���Y�.uf+v���I�4��x>4����n�'��#��l����s��4)5Ͽ��a��T��hf�O�>>�C��^�'٠h �[���)ͫĥ�����%8��F�|��37�D%�㴱�֟e��f��߽"qHLטW��ط��Nߖt$_U��V�An���旝f!4�A`���.��\y�$#��4�q��hwM} C���}�����D`���5v\��ޏ��]V�P�r@=kr������8�� %-����۬��_��Ƭ���vUT�.D��؀��o�q��^��t;���fl�*��ȱ(�R�pte��h��q�� �8z[ �v)ۅ�(������q;��Z�&�#y�-珷d���Ō%�2�W�����羀	V�g�l���/j�'� lkz��{؋f��u-�Hߚ:`��z�Cduv�ܯ|�J%���3f�"�6�t���!�>�Nv��x���r�KmB�n�{kAR���dD)�n���a����[q�*n/�lX%}�J莛of���. |��ڌU�?�zjs,�+iȢ̛�{�����p m�ej����e�[����
�4��rª�{�ٝ�U���g�(�K�MG�j
�U�#��ܻ/�_S�_L|mfv�N�E;&>�ѢŠ;������9#*/Xuj��Bho��v��+%�m]'�{z�V�.��
�������	_4{��q^���We�3+����**�P��ř|"��1L'VS�����<бʷ�#R6�h��d��Kw	ݿZ�����R���!�X_��6�75�_ �4#3�/ฬ{�Ibl��e �a��O�ݾ��8���SjBge��}ʺ��'�Z�&=��s�c�vb��>?�*U���N�lRA���3��Xb��5�W���]�R� C��6ڑ I�
o�߼�2���N�)-���Ϩ�.�:S2&=^ ���2�Ýi�>�L�:��a\�S�J��po��ܷO_�#��o��+�����(�*N��0]�z��6h�ӆ!G���|�j��0�Yj7��Juz���hH4���ƘS�Gn��@˛<&ZA��Z���}�d5����e[�_T�=�ͿQ�a��R��1�0����*��x�\�����i�8��yD�	�O6�G�\
D�����$�YY����W��q�ǫ&�Z��EG?4��c �]J��{��3����pW�S��rc�v|���~�{�w`�~���C�`0�yp"a�n@�Xh�&����� ���y@)Cjz6��%�Uk�6e5�R��1}佾�eTӑ���RNQ��j#�<tawI�'���EN���wI�eE<�؏�mI�Rë�QV��!�_(T���E�s=�����wLyM�Q�Զ���X���db�U��P.Ơ�/��.c�&���G1����?/p(TDg�(m���Cć^��`�߰a�FυUV����K�պ?�ၨ{+2p���/�h�63@r�!M0)��)�^V �d��vt'�R��$��Ǿ7F�H7E����;�q֧:��h;�P��5��T��pl�v�� Q&��9O���̕s0��G$\61�>���M�m���ݾ3��Y�|�E&B����~z�J�&L�D��7y��=�/N���ёcʗf����̴���C��(�q^�	��$�������&��'�:%�j8H�n�3��J+��/ �/��H�a�qm�Q��)Ѕa�m�U5����V��5�(݉��"TnY����4e�7i�M@rf��#��	_`����?�(�B��1�i58+ȳ_u��]щ�4�c���( ���IM?*D���#�*"�JS�#�Y�'; � ����I����a.fϱ@HL:��	 )3����#�Ƃ2���S�*+�{�;^�]�f�� q���c0c|Av�t���?�7F���Y$��)-V5���!\##���n.}&)����Yʃ�
1P�&����d��{�`9��:�gۈ��ڛ��9��7�K�&�$�C!��jj�$�Y;%��B��3U��N�!j.��0�ځ�}�p�^S��c�p1���U }W��� ����e T�:U8��OvH��浍�Xf,��ݵ���z���ly�]r)K�"��>7r�s
�GQ:[IH�z	�24�0_[�-ӽ���׼� b��'}���>Щ�t�% +��%W��ZI����ДR5��ߩ1=�!Zr9�Zo"���Gk�Ѩk�O"�#��
���,�8�K7�8k�IH� {w�]�7J���d4����(C{�E�L.�l`���`��e��c7�Q-�v���� �:�Y=N^mU}� _��(����HI���fi�W�&7����<z��\/�*֩P�?�>�ա�772�󏕤��j>�G~(mcP��6>�C���è��H5�������C՘�׊�8QK�bW�}0��c=gi�_3�<��aym��5�;�*⺱D�q�j��[���:��rT̂P�n���7�%>��n�#�?��fk͸؃)�Ȇ�dW/�z��6�B�l>GO��;�||(Wi��%k�^���;~Iж"cW�P'��V�q�y���7���AHjQ�7J3�P���za�>��I�[��Z.sdG�(�bE&�_����jL=7�Y�����5�&5ث��q%O��^z�w\�'�.Z<��9�9$�K�tL ?���:z�"��wtC&:�MӤF�ɢ�52��&c�,ծ"��$˞. ��h
@�!P�{����ע0dmHp��w���d��f2����)c����L�ki��\�D_Qn�3��9_��aa*0OO�0�A��O�>o�Þ�g$K��9������agC���P[WX���I}v���'��]A�*y�R�':�ܾ���ৎ*3�U��h���b�|�`L���n+��뼾��lGZ�*d��x�6�
RٷN�R�h��e�y��	�P��B�-�G��:Y��h�eJ��]^��0U�X?yY��vB�r��^��I���vJxå�'0M*jl�z���= ZZ��Ѧj�5��������9Wct�TbLa�Ă�Z+J@�sB�ؙW�<���M{Ջ���	t�e+၊uk����yU�;���--�:zĔyv�/F�s�������k!�:ˊC(�׮ÿ��'���|�[%y8��z�%������2����� Ʈ?e_k{���xa���]nD��e�>���#�M*݉�KX��<��yBS��z_������	�qZ����GVs�̒<V�v�qT�h�(����ng��{~X	g1G&�1���x���BA�lz��g���Q�>���!�i�a��)�
�����'�5�m4���X5_(��>D0���ȑD?�T7j|]dF3�+p�4åS���K�Tm�kGk��3��f��g�4�{��p����<^pTϙ?$s����-��V	p�L&��[11�T/n�%�.��}��~g*��P �o̴�\��.�W�[E%)���l�;g�[TJ��X�&à�&����5ֿ��'���m�y!l�4�c����_39�w289/!᪃R ɋ�K��t]�17KЬ�����֖`q,҇�ծG��?������0:���f�6��>��\��Vn1[�q�@�#'>�zI�Sާ���[�Goy�8o'j; �e��*�a+�L��[ÿ�H�x�V�9��_�3O�Pez)��s`� �+{�^3�<ҨUO�Ho/J:���)�e��ޓ�UK"1��h31����\���v���ߟ�j�H����Ѳ����rdΙ���I8ۍ��'[S ͸��-w�`�G��s�t����c�u�z���b�?����u��h��J!�bvlcu͢�IUP]EP�,�K����� �{�X�k\a��dY���+[D��=m̫�,�����xJ�����%�����@$��}����O��I�����,�)���oyF>��Z���Xy�<A���U�
,yۅw�:�� �&ꑤ�f��B�UDy���8C'{��Le�`g�?���*����9z��;v��r6R�]�[e����MA���&�:���?��́\"z��Q%�����(�4k6�ك�V�r]�gK?o]�_���|PŘ��J��늚/��Ｈ�̽��GQ�(V�:�h�7۶�p��/����A�)s(�c�6��&��#�_?GyZ+�2��p�rS��|�A�&-֙␷���Hk(z�({I�����\OӍ����i�K���5��f���(w�
&64��Z(^Ë�m�ʌ�`PZ��$iZ"(DH��%$������I�<0<% � ��{��,U����"��V�؏M ��[�y�3�4� �!`��;�)"�1�'��|'a����2.{�W�j�O,E@4�W���M~H��6t�=��"g���!�?�bg��5��m�trɒ�M:�1�7w1*0��Rq����{Քt�0� �j�I˸�I&@:BC^����I���{uq �*w�����X�R���������p�4���0x�)Gv�4�����n��ﱨi���媰�x��W,4Eˁ#v�'j5�������@D}��kz�Z��8�})޹LB���:�fw��o���r���Y����y���K�yp�&�Z�ܶ�n�Fe��v��0��z��n�$n1�h�+������zj3��PT6���{�����i��qM�Rfs+�vټٜ���c��o--F(��",�A��g�k�9h0�^�c6���������x�<���G@�đ�ax6J�4��œ�LHd�Yu�H�(�A�zE �4��y�U������Z';�ɐ�N��P��?����cj�]ԃ98J3F�'��+����Ƅ� J)�D
���N�ܕGBu\OS�a9��-��+.o�^,?a���B��۝0�N�-���$ѫ��9nB��.��:~�<��/O�g�i�g�A�|�I�\����J5����������U�ʾ`k�c�H*"c�T<�lW/�-ʆ2�g5̐#��]������Z�׆-�Yc=n�O�J�d�����/[�y�����:J�W�)��Q7��4�m��i�Q�j�7�һ���_`�1R-}`���O�@���P�"�N�����` b��A���}�!��@kO�{�%�u�^����R#i�AG�E���R���qʔY���3�`m3�~��ϼ�j?f�E6�0ݪc<Y�V�I9%�ݟ��Г�(���?��w�df�Vh�iU��ɍ�߸��Ԙ���g=57��RL��i������7�:��Á`��m�̖����HE0Νj�)�(�¿�5�O�;W;�R�2���G9���6�BR{�U�����o��CW�X��|��� �Guٛ
�y7���H���?��F��s;�o�-& ���"���V����AtN�E���)�������f*�y̥�JX�A�{K")��L�|�GA��|B,q2��<8��ɥ����Wб��l��r� ���<���D�L^ncBX��YZal���[�=��=m�\iy�xM�w0��iT���k�wV���O`{����p���z�� �,рК������th��٘,U�ͼV��Ǎ���(�"�@�5Ü���
���R� 6|�")r�GS�~��`�ȋ2W S���&$�� 
�w�����g��32�`}TnR5���$�����X"��������C�{~�a���� lZv"fWl�
EV���C	���1N��Ԗ%���D��s֨�L��*˵3�i}[e���Y��\C�;�,AeuBr&!�N�X�	�2��ST����,���A+C�B�'���j�|%��Hw	�V�ķ��9#-��c��Ұ�#Ӧ�T$|LC�I��a�@3O�i���ư�G�� 7קv�N��	�m�_óI�.��fEl�q:k0��Q1��_7�[$��e��c��:�c�6097^�X�����m� Qȇ�!���Q[�PК�\��A͍�E$��%��x������0�4�x(�UI�}�[G��Y0[zL:�[� uީ�̵��F�7My�]1�����I��Wo#^:E��y�"��2�-�`���o#@m3�`�:�ߪ����ĩJ�b���n�%AH�.�A�7u�A`,�.6ez�Y3�`)>�de���m"�I{���W�����~�j�/���ơ ��0=�.�D|�ٱ��"����( X70����"�����8�u�mp������0��X���8	��W��f��4��v11�kNv�]�)g/���A7���GI�x�p�H��&�M���0��&Ͽ�b`+2�Z����X,�^��	�3޹�����]"G°�Z���T��#k��<�����m�NB�ii9�����J�N�`y�S��%�Tz\cWt�-+] 1yC��3Q�4ai��dJ[�v���|�OM��R����'ѱ�X���Ʊa}�nRgo��hST!,�5<>�F�҇��z
š���ԕ�� 9��I�IX��`�ϵ��as�2<s���'���@�c���Ny� �S��0СqC�o�@���i��cL�K}�=��='y3����b�e󠯀+u���0#�B�d� ���,�C/�?�gn�G��F<�D�0S���;O���Rd�� ��nk��@�Ar��tQ�)�p"hv(�ʌү
�Ʊ�]�餭Z �++Y����Q����H1�a%Xۣ��H�~���Ĉ<2>5��/��ݑF��ce"��I[y=1������~0<h��y�ZZ�m�f:y���*�r��\�̚F��,	`Sp8\@�1s囹���Ʒo�n��q���Z��>��#����*' �������a�Г�F�;,�.:i�!�!�-��\���􋺣�����Wƅ�r#�",LF1Ῑ���|��Ěh��W�Oar�*�� `���Wrn��Sd���q��Nk:�`W6w�1���Q����B\�ػ*z�?�z���@ʮēA�f!N����_f�+��>w�|�]	��騲c� �D?=*��*�yn�/R˯_�X�6�|���5�C`�Jpm&h��c2���ڱ����r(��?�k�a8�X����e�t���*{ �oV� ��/nh�O h��r�uLq� ��"a^��^&m��Y��e|AAY�v�~y͊h�L2ei#����?a��/��`�5�����w~=A]�$�s[.Sت�H0���ml���3�����8�K]+���z"�E�͇4Ҕ:��?���K�q�����ǅ����-�f���x�	��V2�D�ǰ��򙽉�QS^�d)Q�F� 	��aE ��V��9���f<�>_Rl���g�JNG��0�v.�l|�XU��upip���1q(u׈)M9r��M��)� � !�S<���:ٵM��=�R �|�%�&Ú��;pm�w��{��N���)�2�ל�夅��셯�ڙ~��B��[!
���r���y���w�K�Z��3}Ǫ!�s$g����Ʈ�j��Y�=�1vwLJmP���>�+���X��X�o��Ze�	�g��_�E��AdD�6���3(����UC:=��+|ߢM2����9���Iqh���W�K�(Dv'�����.�fX�F�j���l}.O͛-rP6 �� �d�%~�� ��%����
Kiw�`����i>O$N�HN�^!�͐���3�h���?`�f��$Ļ�/q.�ǤJ��9:� ����}3���m��jB��pxsH�N	���ߜ��5\��~�grj�F���B T������I/�)%#,�$�o6�u�"L�\H_��#��~���q�X��=��?�1
%��2��M� �*]4aG�t/V� $��O,N$~� �Y�/m0��O8�6��?dL�H��m��l���qUy�6;�����{���\�	c���#sL�4�3s2��.S��ӟ��	��!�B1UY�.U����F�'R��<m���h~W���a�š�P�3�g�a�㈌K�A	�&�"빛�Մy��8�em.����;����J6��>��H�UƲ/tH�2@�<� ��EI�g�r:�N���w<�]�w�������HDYq%㞺ג�q����ۧ�H�e�bʝ����NhR���&d0���<��g��T�d8Y�~38�(�}�����mV��R�J�떧��S�a��[8��Z7r{pf_�I�lYoWe�#OMKAeNǓ��
i�Yw�%���M$8l$���Y���@Ҝ�;�����K�2[=-����dKU쭢��Źn!��vY�Ð���d3V昷����$���Z�=3&ˤf��"FZ��l��{ ?��*� �IxH��M�6�zD�ra��m߷/�>>�*������c/ȥv��p�m���-��J������9�B�Vf�G(Ȟ������R䬢�)�x���YȦi���@m$9�#�l���B�^��P��j���!a�Q^ή��:A*)�?a�&��l|e{�Q�l������5Mhy���]��R�fNÌ����\U6�c�y��k��\��*��qTȹ3m_*��)֐j/��(��0�n�M*��j��.�J��򔼠侏jv���%hL���W΀)��rJ��1
 �m
kQ�!�{)�&s��Dυ��3���v�=[_|�n�F,]��o�<ߏZi�*@�-��1��}F���[,�����x[��T��� �+_���$�����k���BqJ/��[(�d��:6�|6��L~���Vmy�t��q�o�;�Q^R�!�Ã�ep#r}"\��f�;�ۛi��V����2�mӀ�d�W$�4&��Н3� ,Ԭļ\O�T(�,��IA���<Pʙb<3�dS$�Qz`Cn� �?��>ۥ������ۄG��$���@�7#D�_�u�;Z�$P��Z�+�����)�ޯ!�1�M��ɫt r��6��g{�.oS��ԭc'Y-ʐ�}��L�2I7�?c���W��:��A�����<:���/��[���^F#��r� b9o�W@OP�H|��������D�r?Sk^R�iU)�\V4^8��|O�#�����'��g���Xh�&��Uԑ�x�Ԁ0����f}��,a��L}�r��g�`i�g�4a��	�!�{VG3����	���<ׁ�"�%�/���[cox��$\������D�����z�e7��t�������۸e|�)`;�TB�h�=f�-�l��q���81�� A͑OL��E����S@ʵܓ���-,e����K��n���ӛ���s�M�����g��P�z �ͽ�o�X�>�q�(�ؘ��E�G�B[3�Z;ѳ����˅%�U�˺�b��#֕4�8��<�\�/���˨��?��-�@�T#rn�Ck��M����#r���VW�� �&i�I�mn�V���7�[��C�s���?�۟�H:�o ^�Z���HT(2�����FV�����p�+yPw��B�l(_���M|g�T�f +q�wwI@���`0��!O�K��_7��%�m���m w�[Ù�^h㙯����~LZps��E�h�22��;X��o}�X�Q���6Z�J�X	�xO��U�%*c�� 0����Ϟ��Z�)�z�y��O����b8r`�c��+}mF�W�&��2u�"�t���u'qC��{FB_� �茯l�E�����5�=�$��֞�0ޣ��؁ ��x_vD\�&�yO�+���_���A�K���h�����Iijٺ�� ��+4X�i�5��T��������L���VJo�G��EfXn�I���gj�$G~���k�(��g���i��O��s��G���?�G�_-g�����? ��Kn�H�O��[ի�>��WK�.+�v}S� ���E���
�IA�4G������;,�j�幢���?�k*���0��$�����j�z�h����:Vowh��"L��tH�sZk���I�&���Q�	a�NX��l�d�^]�$��e'SKh1�9F�Jf;�s�z�E�f�@�N��G1"��{Zr�eQ�p\�5J�L
��am��c|T���z�V��u�b�˨qq_>����cq`O`Z57�L .�����ё�}� r���F�+�H3�,��3�,��D�=+/�a���^
2����~:(�9��C�G�"�el_���h���V����H�|I�jMS{B��?[���H�<f��7]��6U�֎3>^��d��V�bi��W��i��e<4�?�?'�`y(�ҋ�ݽ��x�d�v�r'� �w�W�����d?���g�遲g���l{���)�����G��61Ֆ?u���Ig���Т7�~r2+{��V�A��$��U�o�`������&M��6 ��:&��.v��2c�˾�����g�����^�M�H�+\N�đ`ݙ�p?�2���q5��5r?����3jA�j}���7�����u[�{�b�i IP����ŸΘ��tq6�|@	U��Ẓ=��Z?U~�qW���r~�M`�^.0GƲc��Hl�TMM��|	���8����Ē�:����HC�(�f'�Q�:Yݍ�����{��\n