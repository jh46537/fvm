��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&Y�%�ddؐ}(l��+��S<�{��-Ǻ�&��)��6A������<��j$��"�w��	|��:�NK���Ac��JF�i?�I�J���*��4���.�˻,Wһ�@;�xu�j�i���`̒F�u�	MR�.�OLN��K�9T!c�&�2u�8���ʘ�ˑu�H.+k�d���(��.e(,R�b���]w�U�sf�D�y&��"iJId�l j��k@��DS��x�m?"��H�@b_�J��ep���b.S=��%\�����i�Ew^7y��?����XXN�rz��[/D��ӳQ�ߍr|q�GUw���"|�i4Z�5��
�ӟ۬0�Do�z�_�?=B�n�`�*�0W9�n�f�j�
�" ,�X�n���C�:@0�0N �Yy����
/8	��$#G�,]��]����%����R�{�ճ�M�BXr��;��h2���	�t�	���/]js�a8��� t�6��3.s����c���j��iU���$�B�p�6&��������LK/!3�S5h��،��1��a���Q��.�w��ܭ��"�t`L���H��f�]��S����B^~��e͸���6U���oB�L���Gxj<�̾��0z7�Б�9+��I�y�������Gu N�F�eI7߉O��/��������
�ߠ%es �4�'ymn���9�ཨ]t�f4r�^0u��w�%� �b�a�m,����*̯��T����Y:%S	��,�|l�°��G����͚���l�22��� �t���	$FCl�����{��r�:���Eݾ�אN��~�#1M�>a��r��.��9��3�$�����f�s`�D���z!���ӿŎ�����th!��8ҽ5&6a�/��!��1(�A�c��!��M�����0�'!4�:U��;Ic�O��]�H''�鞣�RbZt��UMG���#�L�Jt�B�O�f��N"o�����z�~{�9�k�X?ъA��G�s�y�����*N+��� L�h`�D�$5���ۻha���1Z��Qd{�����`��(.��ȽU�܇j|nr�R೤'�(j4g	�8|����6k��v�91�P�m�wVT�[����0�}ws�� ��r�)
��{�ף�97t�z���ā0d��;�|&�G�����4���K�����k�j o\��Ƒ��(-V���f\^����埮=Ss�����|�.�W�i�6v�-y��iS�C�ɂ�VkH2禆�L���SA:�O���G�OVz)�_+8���E��T]lG�zO�5ϋj����),=��'f�d��v��	���]'�_�c?Tqu�c�^7���A��8���-��~���p�ʪ>���o��^]#�����(뉞q��{�n�>�D��cz�L
�+dφp��`�D�]�n�S������l�QEB�l���O��D���� ���,l?E����)��I��@�i���>��.s���Dq�@���v/����m���Ҭ#���dN h����y0�Ԫ�$��������K�:j������\e��>(��Q?��i:��Js�陜�}!F0pyU"�~?vqo�>��Tx�X+���d� \Q-2h�Ac�#,4��Q@�ͲX�s��f����4���1�YMOW��x���<̭`�8��lx�JQ��Xbz k:�ʲ!5�	�Ϫ7��N&�ךھ�.� �~t'��(��|8�v�R�n�#>��S�Jse�dRv�Dj:�X}��zG���jL���� �!�K �X3��Z��8�RƢv��Z7C@Mp?��`Ou�7K�
'��o����x˚cLq��MP���]T��D�g��{``+��eV�׆}�=�T��d���e�ɩ�4'�����9P�iPO�8.p�6�IF�%g��⇯�Yx	�QN�<��`�,�!�h������҉*������ʨ¢e��������n�FWV���Gu�{AAؘ�jEs��_����e:��/��O7Щ��<�U�0x����D3rZ�z=��_��L�����Rp]&�|?�(0��m�k ~�"��"Fz���*�dr�W�hR�ݸ���M!WP�fES�O�z9G �'(�p��h53���%���Ͼ���D��{��=&|_Hd�t��k�$�A��V�Hָ�C6�2���%�I�߅5:���� R����������ɺ�g�UÅ�@1(JؐğG|�'7�E�3M-1� �2(�mD����
��iH?ֺa��3������� 8��7���"���&jx�[AZv���r��} O���#�'a���m7[$�=ޡ�	4��w�j*��T�aٗ��#���O��}-/�f��e�?D���ΙCɵ�Yh:�[=HVC�z5愼��ڙv��^��>drá�3��+�ɓ1��e�h���� i2m�h���J��II���A�{��Nu|7�-Z��jW�����w~) �R����[� '5�lLr�Th�'Z�^&9V��>SȄ�0�5=�!�9jnm]/�tq�z�����h��/}bT�'��e�W��,j���	g7�.��<��pޱ� ҅��ٹ�am���ٶS��9��\���;"�~�Gc=3*�A�?�2�/w+�Nt[2��F4�s�A�@`�R�Bq��G���x�P�k ����n�w�(�ų�̓����oT;�;�w\�*�����uy�s���c�|��xۯ#-�9����kɡP�X[��8��:�N~����0NO����#߭��b���Z��C_zi�]�ɹ�}��o\�P �c�u�e��5�V���)�:���n�)�T"�� o:a�i%s		��@nW�?���0�]zJ5�-�5�r���:���$�S���S���ak�U�gA�z��'x>�"S3��޷����Ou��ǀ5�A�;����b�j��G@�N�$�>�<�O�e璤j!�>�{Q���WS'U��nm��]O����"�,����|��S�\�aUG��4p�D�U�ЦkQNS��'yp�����9�~��G��6a���ʟ��1��3E�D���k���XYa�{�6<taX�R��@('�t�'ʖ���/���`��IP;RB2�b,�~�y>U8~鹚q�l�X�E�"7�l��ܫ��"~M�u4*�#l3l��ߣ�U-yu������o(�J9�CB�/J�p�l���CX��>}�bG�Lk��L���sL�%ʟ�ڿu+}�2"��$����C�Tc��:1Q�Q��`4�/N�#�_-�פP�N��Z*u�ۉV�ЮE��f��6��=	^�$:�~�������ι|1Q��Y X+�GNM%s� <%�]��A�͚G$a��ޠ<KE�W~��$ܨy)�q��%-�.U��A9�=�d$)�4i���K�=t����L��y��0�Z�!�(���B�*K��W2�`{֘\K�@Q�jZr	O�u�ʳ�B�d��,MN��}xΠCx
�P��_§^�f���hb��쭰��dQ�~O�L��y=<�9�� .%NϏy�=���Xw=QK�,��&�(%�%�$��t<q�*�#ȼ)?(%���Gh��s[����*TzI8���K�H;_�@�*��z=�k�7�bd��*4	x0t�%+'X*�����0�
;�復!W���Nw����ǒ^����B�n�-�RԚX4��#?[S���͡ ���t��
ԟ�=Q�B��j��A�+�I�)�B+��"Gb���K�����kԠ�i2�z�q77��k�xy�&����Uɒ0/	8�~��/d��J��������2N-`F�WوT-�v����m��{�)��t]%��|��09����P뇭����,��eD7#�k�ɼ7c�Ux@�ts�y�+C� hv_͛I�Xt.���	ˍz�q/����r�>�P<sA��cB�Mۼ#�$l#%��"o�f���v��6.�����P9)�R��z��*��Q��䡜Tɤ�Җ�����d�N���=|����	 G�ؖ@	l��	(�=�ԓ�BIJ��U�\Dq��W	�|���vr�r͊�cPC6@ug�(��T({.�Z���^��X�|�*m:u.G��2���u);�������,����|n��@F��Gi8*}���8�|ko�}�e��g^���s"8�r�w�\� |��d�1*ܹ�ܑ��}!4?��1t���b�G[�
�Ͼ~���c��g;�fI�1"�W"t،�%�}��;��9�}�? ;�5*��ԙ=:2��3��BV�rNp���+h���Q��t�l�����}m����҄@Jiñ6�9����6r|��
��2-��vEanU��Oi>��Yګ�8¬����~[W��*�̍ �V>��R���D�!]�$#���,5��A�w��u-e����KU'�3�.��`�M�&N+>�C��rP�:��(����\P�&�[��f��%1��(i����h �Q<����R���.��$oؓ����,T9�8����q���V����l���ϔ�R$�紮L���ȴފP�q��'�Gۆ��������ڻ�}�tCu�����`���^�M5

�/ͅ���F��V8%�~=�%"go��E����`:�+�*��#֥�=۵T��Z^�N�3����i���HzJW�z�f�QU5XS�����U��+U>�/���X��}�)��q�k��Pw����_y���?�:]+�E�'�b9��U��	H�~_�~�[D�a�D���-�!��S��N��zL�vOy���D����b�f�\F�Py�z�O� �L)��`�43�%�)�re_T2����5:@_i3L�n�?���'�����W��@|�F�Ӄl�U�k�ɂ�V*6�瑟!�¡j�c�G/N_YE�=^�E�6���6���ji��C��ol�4}�f�4�p�� �:z^�
�A�0����G� :;�+f �-H����Y�[����V�}�[����\AˢB��ފy��#ʪ��$\H�b^OY�����8q �[@^F7�����C޾E�7�(���ZE���[q��Dl\I&�!��T�l/�t��g'��=�� h�LZ���QV��)'��5O��dc�n_k~�3�EM2�����!��8��m��B�sw�@��'~�BO��(LJ劈C�x�S�־��������*�+$�$���P�u�F�f���QIH$$���દ!���֐cҬ.�A1C"�
�%c�|ݵ���$V�H� s$9���3Ɨ9�t���v�HQ<�������3,*t���բʬ�A��FĦ����k�S��s<��ݥ'�U����Gb��6P�5qP�;/A2Ya.��0%)���&�y
��&�>{�?<Z����mȎnJF��+��N�S<Yd�A�[8�$�]�`g�x�p o���j��_INT+���@�h�4������\�g�pZJek��!?�c%R[f�p�)\ʞa�*���5M�)�=�7���@W\kk�2���0�?Hj��,�X�h�� ,��\r7$��ywo�M�>�� �H �3�6���3i�#��(�e�"/F3utl�@2�h�W�]�_kz�GTJ��3�I8좠k�j!���ǱRYE�J���9��ܿ�Α�^nX�Ʋ9_��+���w8H��:�q�fɏ\A��D��!�:��*z�ǎ���k�zRU���X��l6�<f�X9)4M���+��au�kH[�,����������DiбԤ�z��Ƌ��&ǷW�Ch:ɾ)n�d��|�d��s�!oa��'��ہ�N749Y�Ѥ�mU�j�L�a�[�=%��l3X} ��Lyϰ�������}zR+!�$���AuN0��`��˟��d�mZxi�8�I1-�p�|��9�
�28�i�>yw¬$�n����"BiJ$, ���C`s���9Q+�����1�c>��(�Qq
�������;5�!&69_���'���ȩ�K5�����wމ�Xb���=oB6��Y5�7��إf5�������t�3a�17&��Pm!mh^���)pj�O�_8 �})�);;U�%�X�#Z[>VW�74�m[��N½R����F:��� �
�<��L�?s ��#�bDl-t~�"A��V��D���b���^[[����9;���8��ό���y�nw��*n�8 ��߿r���b�)5�O��<2��AM�2U��=a�������Y�t9� ���%v7����m�T��!�A��6�z��:�����Y��� ��j�Ԉ#��&�����7��\�ak�'T�I�_�&9`Y�r�}�u�We��B�z�L5if(�	�	��x��x�����%a
 ?���EdµÇF����(��)����?M���Pf�Y7��$ja��{�v�-�ao(^�2�GxO^4 r�Q�]��ڨ���b;�}�GrP~Z6i�?oE�H����	�87�ʿO��1,��ȡ���(����m�8-i(��6r~��I4�ӒI��iLkC�!�`0��<ϥ��짊�����~l��^�\�1%^]����CM����zΐE����2���/6��Dnef!yfx����k��$��&�fο��q��ԏBT�'��hO�0
���Y��ɢ�m��"O�4J�~���G=!3еT&�f�",MsAP��?�3�W�  �˗.�؞0R�:��>٣Oo�IRdf�����j �<:���;����]&�R"�6���H�����x�n��Ɛ�;������?���&:Ԣp6k�#��~_v(�\������,�+�k��J�.����>���~b$�a�ѝ����K7��ָ���V"�^��&Y�6}�~v�^�>��yF~�ր���6҉I@���y>{$��&hP`��r\�랓�P	 �$���7�\�p`Ƙ����ռ7#1�O�Zg5���'P��lR��[.7)��Dû[LQh�@.c+���T~��簘Fk���b��d��Y��0X5I*86���Q�gE]T�f�bbƁy�F�g�2vd1�h|jP�d�1%�[���3n��(w�{�$�4�^��P$
�.^�>��|r[e{��gtu��3,L�L��o�w�ј�Bݨ�{���&�Ul�>Xn