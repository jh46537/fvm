��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&���2r�"y��4�] �;u�F߾��Ye�hO�%ROx�<�G����$��Om��B8�fb�&B��{����vK����F\��Y���埾�}�#�njQs�i�ad_D� MN%�
�=}�-�/uEn�5��Ye��f�����OM�Jz����VW��N
�U)�07��c
�����&��Z���sȿ�7����(��.��l���-ھ�F�r٩�1"�*�閎3���L4��_�'(buGE��?���8���[d5�Q+.���m����/�߷Ҋd �h���2n96|��PǦ��:ЌyP���F�z��k��l�+	�/�(��� ΎVĔLSq`�s�zƺl�᰸�B�ۜs,n�/ޯ=F�ca夜�gx?�Y��剨Ӈ��JseK�G�R^�B.���_Wi4S�$�v-'�wѢ���x�I*I���v��4��+0����j|oic)��H�9�+j�!�F�tF�5[P�[�0]KEr��1��b�+寕�!+Zi.�N"ɽ)����aL��bH٣���ڴ��򀲙Zus�p���,����1�jҊ��Q���y� �հ�s�9�K.ㅇ�4����J����x���{�mu���n�"���;�Y5�a�jL���s���C3�Em��K�g=P�]�]R�QE���T�~m����b8|�݌�U���ԓ�=��fkW}ϺE�*�\�g*D�,Dn��WX֩��E=l�	]��L�إ�#.�	�����&>ۮ}Ӻ1%��DI)��=׏^����S��������a}	�3���hb���U�a�+�ma��N�o-���h���H{��-����Ա@x<�� _��!�dB��F�w��6�4	��QCТ���G��Yo:|�5G�jB5�k����7�Y�N���HIX*�RX������{���B��:��U��W��	<xr�@��v��`!�Y��}�G��	��2�I��o��� ��22���<�'�p1�9*rʱ2�w�ct#Ĥs����(�^���M��>Id$�;:?���_�&�D%�y�V�gK$�W���_���v�����^H[,s���v|�t D�7�wU�{��G�S���A����$��59��R ���y�hw�����{�>2�l�`��
�ݬa��Y��Ù�/��X�z:ht�3 /U�_(>�i2��d+p����:j&.���;]��m�o)�dF���>�(N �/�w(ٯ��W]�J×��`jg�G��@ ��\]bA�^Y:���嬻�A}c8K&!�n�#�������o�����]�ܶ<݅�ť����0���%G)��/��wc�Dū��d�U�+�Ti����E�f�G�(K�~Tv@E�*�-h<k���!�SN�ebW�K� �q
���fG�5	o�� ��N[,,N�ے�-pH-�܇��Fz��T�E���k����hhZvҾ�zP�2�^��3O�!�k:�q�܏��~��Wᑥ�躿$H�Y�+�̖��)$����a�&_��s)jU��q� �M��7T?��x+�ӛ��]%);�����Bh}��Z�8�,�b)%���`����� 7��mz� �� ��1������z?1#�Yv��>6����d9��l?�q��Pz2����èi"̿�I�4i�ᖮ([~�>�������.T%.:X*Fl#�JwԉB���*Ԋ�i��W��Ԩ��w��mH�������ڸ� �Խ��q_�ҫS%XY_�f��~
d��Gp{��N�vK����C�1�d+ �+��m�"�S�X�+Wq�$=Q$���[s��-h�Y���/�8gP�9B���(��Ԡ��s��1����
�.�Èx�;�S��E�
����HA��J1A��Rk[�jo��S٘iۅ�+x��ֶ�W�9�N�좀�Ay�f�:�J�P|	�Ok�H�_��1t�-�\Eq�R��N�HU�P���v�>�A�ct�Fʍ��UU�A0�|XW�p��J����-��Z���?d�%��u�u1zpqe��5�k[�e�xП0�1�����|Sz�.@�ۤۢ��v�k���ň�ģ辺��+��{Dօ`L띉�A"�ߣd�U�7p�kD�7x����72|oS"� X�'���A$���e_p?S��#�^�����w0��~��B���#raʶy]� ���R 
:]�A�>������oq�J����W�A�d�4���g������N:�R/��Pݬi���2F����T���+ `j��PZ���[�w�@F� ^�(�b#�w~z���#e�M��(��a���HAɒ���&Y@��j��h#��[��-kAD.b���_����m+捨+]-�A�T֐�_���|�G��5Ó�He�$�_�Ak�~�,�22(��9*�&�5�O�����E��@��t�2�������b�w�F�0ƷL�a�S���}�h�V6�]��uKx��5(Cτpw>ѿHs��X���Яp,L�A�m��/�r����}��Z
ڞ��!�W��s�Ԇ���l	p.^f��}ڷvf�� _½2w�Mk��5�+�qn�|"�6�>�,GΏ�b��ΟT��G�^��x�V�=ת�;�b�V���,8g�`�H)"�:��I���9G�:Q���	�?��iY��R�q�er�S�8�^5ty�e��ۘ�N6��}E��<1ا�X.JK���G�"v//r�`a�z~E�B5����[��+�9�+�� P�%���F�dꀸ)�d';~�0qn׌��8�43n��eǷdO�����"-	{�����p�lH�UU��T�`E��L�+yY՞*w(>*������6�Y��٘<h�Qǟ$�����C{H��OQ�,Ų5J5�}j�Kd��q(���H(��4���^Y��G"@^���rÒ*G�y�*Pj�f�f~���+�?f�k��n��A=Ć��G{���^��S²`�;`����﮵�yL|&&�Ȟ���6g�e0,�T_�/:�9����aI�)j��� �N�(�^;,$�Gy�W��sp*m��eU��I��a�/��Q�nL4��|�7��"e��9��o�ac�%�S�oA&nd)�}"��VdͥT_�DHb+IR�;2 �C/"%n���^���`�%)8e�%��W��,���55W�z�5��g�J�-����d�L2�ų߷<5�5������w�����!�O��wn}���9h��=�{����G=����3��d�6�M����p�w���;��h�rf�CVb���%��aF#����e�W�Ţ�5Y���^x8:ɗj�{�d/D��~]!�����|���օ�>>Z�:;ԗ-�e�G�;�!hݩ.~�􅶽&��3�r�0-T%j�6A���G����1h<�[�h˙Z�M�~�YV�qF����m+��7�>�e�#�"�)ǈ�����S>���b2v�^��,%��i*�U��Z�7��E�σ"vh���_kJ ��� �^��-��\��	�,��3��;�������.�lM��:�ls-v�d�8D��"��}3,�tN`$���l��f��e���r���JLE��$�k����^c4` D��٠�];'I^fQ�9n��'���z� �I:���+�"}�c�_�\��Gg>C(��8O1��F�<N��Ț���W�gL��.-�;�Q��X���8O� -"A��\�mXd��$Jt�*��ӏY名pϻ�Z��?�+����w�mWH8D'j`��A����[���û�*a���A�܄��<��2/�@��eL>B�B�9�,Ɍה�C~/;�Ѐ&�d�T�Ӆ�����0l�4�ޯ�������	�u��Æ�@1����f u���*�Y9(&S&-�/O��oD=DM�2���y5�qe�M.k@m�nտ4	w;��v_��C��o���eX��2~��b�q�b;�N�Xȹ���6���c@�����KA��҆��o@E�����}�(?~o�O ��z5;2��_'����|nحɘ�	�N�n3�8��t.�wa-$�9�oʥ�X��Ӊ:�\_���"��������xzjAσ�Tzib4f�&6?�a sʰ���.%��q�X�H-p��i�f�9Lo	��/3_�Ь.-�I|h�p睮YX�*M�hu��i�)>6=5RF�c�ӳU��V����,l@���e6�|�b���\��W5�-��P:�%�3��\]�� >N�|FKs(w����Y
�흣���eŢ� T�t��]m�\����ʄS�Ȇ�g\�9�G�w����wo�d5��?"�:S�j��k1z#<?�&eZ*�dK ct���� �?����>�ƺ��5�z���:4�m�w-;�6\�����]'�Ζ�"Hʋ�|H��J��A��F�Oģ9N��"я���	�y�֮ᄱ���D�@�pg[�����3�
6d��3����xT���0�pq���@��f���/�O�l��9�$�"ż��1��:�d�܅8l�S~߮tҘ���{��}_�5�7����S;�C�6c|�k�{��`��{J|L�O�ܪ�B������Uoz��/D��:F�H"� <���dYٞ����U��峉�\4P�uw�e��z��ۿ�1�j�{B0�:��0����dm�b����� q�N�M��3��^.�����X��hP�	����K/.�/�����R`�zT�Ģ�z��T���Rb&;��p��]?4�-�3��f5˘(�[������z󌭕x�;��RZ��z�S�{������׶<���_Cf��o�(��P������EZ;�S*L�K/+��j ����\�G�x�Wy(��q%E�Z3��P��n�f��U��N��������y�[ �M/4�
�eH^��m��;�)e��fz?U/vz䦧�9@o�܉L}�t�#�[9#�9Ua�o@LI�e���i���Z�;s�%���Z�Ȫi�)���� ��Nٲ���R�G�r
Ф��*��/$���2��X�f{��-N�'�1tBJ���_طw���) 9�b�?.�4�/���,�y�1S������!H�H�g IhpZ���3A�T�g`ɷ�*R2 �d��ݟ�}�"v��&�:���(Vk.��oK��c�Q-	�U�|�+�@�yIB�9��<���	�j�M�Q*�c�G��H3�Ю1�.<���q�[֩��4쯅|��ps�<���3�p����+�����|��N��#'����F<��8��B�&��؎�i7�_��{�g#�	����X�/j#���R��R���>t�1O�l��wD�z$L�;~m�Co���&TKE��w�X�f/����.xک���"#T�J��Vs� �xCL���?6�lvy��}=0	 �m�T����]�o�E��=��$>�K�Q���"	���Y���#�p���9~�M�0�
�k����R�b����|�{g������<�ISB�U�����u?�SMD:A��	�0�c5U�嚅��Y�tN��>O�'��y$�� Ԃ�z���J;�U���V�w�=��$���}g�k�5)�F�P%�ی.A���t,D��q�וA��!~�}�
(Ԥ�!��J�����H��7�~.O�CZ�G�QM�?c�k ��8����s]�1
eJ-�~�{�|�a��q�0���RI�_7U�,���U���W�9���wqq�ؽ'o���n �8K�w#՝p>{[9��f�j�F����E=o���f]�ZU
!]��tS@���_�Ut<NAe����6�Y�|�~�V:GS&w;q�aSaZ��BI����,�h�Y.����z�����*<��&=F�L�#V͜�;�2�P�gǢ{�#B�s��&ȩ]s�C�k3 r?��:�K��k� �g�jN�ܸ�3���Z�L$mp�!0��z�P֖�_a��nGRgơ�͍��QF��L~i���FZÁ��	�X����]�s�8Q������4�R��(*�_Beefo���N�(���\E��S�N1���ؤ���� ��Q̲)-ԯ{+Q�	v�IN�)���E�T���E�dy!=�)Y��6]g\ϲ��|j>��6]��V��#�g�EZ�y�P�gm�JLܒ'��O!��(3��0U��OS�g�j��w��r�d��ٴ����$�C�rD�Sz�>���A2ظ� [��_U���:�?Ws�ld:�
�m0�����	��*�*�Q� �b���qu%2�p�x��%>�g���`w�7r�6/�g���Ve��֊Qlx��q�C�D�^G�Ul���%���(s y��!����u��w��:6|�(��*��2���t^�tyB��"��@L�h%K�/�O?F �i��⡆+��ŗ�X�t����V�M�4�Y�rڗ �^���u�a�ƙ �I�϶ş%V&la`E�!�_�!�n����>���X����=�w<=�?���]������������75>��ڶ��&3�@!���-..CV���>��̗��.|�������ʺ��;�8��$hA%Q�{n���l༈�����H�Z�FGI�oHoC1��	 ]%��Z��M����;^dba_n[ �l���p3��]�� Y<�p���_�ۏ��Q"N�k��@���S�V�4|S�)�/:�C��B*�]��5HP�"����9�����kTH7����H9�\r0�����j��i������~��8�%(���"2LJ���e�����X�G釈������Nu*��_��1������H~���x��%N���5 V}����{�a�՝s�f
ЦUzy������	�܃~ͭ�}{���7O�D����b�w�D�oc�E^��s�S-�|C]u��0N����?Uh�5�e����D��!��!/�O�P0A_�l/΁)��=9��a�p��xL$xh[�\�ڈ3T�t}��7��oK!�CS5�W��-づ���G���*R���vۋ�ez*�O���*�	��=��ݏF̃��Ut螁춼"����.�hl�T�+8-�n����@w�y�Ne�����
t��- �[x��P&�o��MGT��B��Lq��A�PZ�*�N��$Г(�쁚���:G䃧0���b�٢&
�P��Y�@��9�nq��VΩuC�[���D����G0�����p&+{EL� ��ee�
��\_�Pv	�F��P�7I/RS������<؃��d�vNL8x�zP�!�J|��Asa$������)(��v$�[s���`� ~�]º�f@�(n��">(��'���<�ʀ���Λζ��w��A[��8��K�Y%5,�\q�h���C�֩J�v��1S��۔q1l�[�.�Ǭ�F��U���?"B��@��Z�A��x!������p$�.�<��l^��	�������D���Q�'��6(�v�O���eF�7]E��u>�&H���~��f��Z����_ߢ/7%�V�޳=4���͍T�Y��h8 B�Į�����J�ڼ��en�PxP6��76�v]~"C���v�����$�&���?ڣDE���B��^�#3���q��Qf8�M��v�&>��w]�G
_M�͒�{k^�$l|cN�n[BG��� ��X  ��3��R����j����2�l�3JB�I�G���;�����8bb�<�[-����:LS�c˒�:�����9�䩲�r��S|��]<W��p�)*�H�[�Y�ߗ�w�ǤG`�Ly9ȱ��C��
ނD���g]��J;
Ը����p5�����]{H�^\�7�6�^�Ӵ�ɰU=k���7��1"�/�e�K@����ɰ���"��h$%���9L�5�"���0�}q�G��O-���"�(2��}��,��]b�N���ٳA�A�Ԗ�2��g��/sBRu�at�n��/�8���ty�J�v8y#�H�K�	֛��6<�|\���!B���,S��?7���d�/+W1��T���b���=$��MI"BaA��۫����'ju �l~��h�SV*�~l�֠^�V?�%�h�P�uZiq~�豯�ђ�cXE��J>u�����`��G�7T1�r��;��@�gQ�o�@65��;%~$�����nqyӤ���|)�{9�q�"�7��.6�����t�LDs6�i�l]�S!�"�}H�ɳeb�['h�|��g��*�)�$XlƯ0d��+uϐ��Ə������4ϩ(�TЊӝWNO���\U~_,';7�`Y	՘��А��:�F�RF��l�G���:������ӯC���?M���1�y�_ӫ�����S���i�&~VF�Bn�'1�&`D2s��Q=�`�AY�ǌ�e�Z�F�\�q� �"A�HC�DĂ�� �ͫ���M���{�;OZ�9�V!*W���wpi�{���`A�X�h����᠌�V�|<��r�Q��>]���僈E���&坄0PB�ā��z�&��,	�\�"�ŷ��v/�\�����v���M����v�3D��Nx�#�������5�JO'����C��H��ޮc�L��C��\زu��ّ�ճ$J�t���@v��t�h��?����5��e��v�O���V��g�՚Z�_1���RR���a�ZchQ!�g�DNy=FX&l����!�G��g���հ?x��%&��.V6���A��y}'�������6�oߘλ��H7D6�f�w�$�"RǉD�����|Q��1"<�N�[�-1�+���c��[��bG�5CQ�B��b(I_
�ڛ�ov�L3��1�r����!����'&�e��4'�4u���n
�0]����*#�.�o��kcQ�;92t������2|��(�96��-Y�³���i;�%A}�� ���3#�p}{j�I��/|s�<a8̳Ȕ,Mo����SPZ�(��'[;�ꋞcÆ���γ�V���8���q�xO ��
*��uݡ�X#�}qN):*�-Y�A��G����[{tκ��a ���D��i�sB����Thv��HQ~X�),��t���A�!����l��@4����bP���Ҝ�%�(K�zgH�ÅG�o�n�IH��Ed�wM����[�IBj��2�|VA^L�NM�{�a���0qw�5蘛�~� b��)*#�ʺ���h_�V%I��Z��ClM��<�W`���Zʠ���l�U��fV����boA���v��W�W��rͨk����=�|β�(O�CT��+�~��t��j�!�qßC>�3�ʅ�sL�;�i_a�R�рq��Mk!$�� �0a��/�����!n�p���k��N�퀤b�!�����^�`}o�U���Xfĺ�t��g��[�V��e$���cTN�2u9�L�.����[apmf��W�i�g	@�~���	�-�N�����§����xU�g��'p�pX��*�^��_�8��F��x3�<��鰭R�����J���լ^��&�8���P*З;���B��?��Z!��V� P!�A`���)R0������y�G«>�� ��S=�jk��s�g#����L���[�����>Cq<g ߘ�;�G�E�� o�N�Z1��ؐ	���eSՏ��zV�tnN�ٛ�Q���ݩ���*)տ��iM��o��S� i�}���ʹ��Nc�[5��'2�q�!�wһ�4#]]�8U�����ʓaUj(Y���*ǅ@��,�^�ݷf�T�~�(���Ӓ�P���>:ï037���J�1�X�\�HY>t^��n|���z-��x��Ȭ���əW	�0jXt8Ҏ�,�}7��X�]����"AV2ӏ�o��z��_�,���D�\Jl�|��L��h�� �����)$���=��f���nr���}N�.&3�D'�D��lE�[�F�wq<���r��k� ��J٧�q�l^���~S��!8[(�E���s�f�l���E�dǘa�Y��K�9_+`����m��w������8;���cp0/ �8-�b�6�=`P]5�������t�c��гݱIT}�SdT;�(bIb�(��8��R���^�Ύߞs|Rރ�Ʌ>T��W�Q=���GC�a��#���3^�)C}�Ùu`�0��lӋ*~3�O]S3c�2��c�D�D.���B"��`P[��rR|p�����B{��TCՖU����8���7F{�@�d�u>32kk�%���i�5��h?�K��=)]��wĞ�s��j�-~�;�I������O�%'�'�8�?r�L3�S�55n��3�)�v���a�U���;tWI���hS<AC�ϥ~�S_��������Ǟl�7(E�q���8X�J�����`^��C�	w)@����J���U�5'��۔L���;KQ|��;%~Ư-�t�ٳ)��TQ�^	��N��t��ZOK;8�؄��O��=����g"���Ѥ����/g��9���S��ZU��5�!㈓�n�mjm#_����$cdpz3���م�!0�5�O.\Kb^�����pou�ܪ|z���Y�팼�T�����J(�2gr��5���`�>�W��r��:�i_9�SG����w�֙E{�Ѩ9 O޾�����0�7���%/+4L�ַ�X�M��)���q
�㖝}���W�F���5��e��>6���a�F���Y���nHKƠQ,���G]��\;�������%��?���5��ې�b'�8���wM7dV�h�IW�5�/a� }-��[�����̀w�v�@;<�z�/dz�\-��g�s�
�22�H��P�5`�|��W�'U�����m�*������*E,����a���#��	�)?������p`�������O�KP
�$�0�ʢ%>��9�_��}�ן�7�|{����V����g`b��{��ewӉ�F�BP�'���^�z~B��ӝ%�q!I��Ak��3��j�f�>k��~9v4}���L�Q��|@����I���o�t�M�����g"&� Ym��
T�+u��u����D=a�%�H�6���T�O�v�j5J�3z��>�*~.o4Ė͓@��@���>+���AD|�8OJ:1���{���Y���'���z�c6N�a��L'�/Ɉ�igo �a�}�����J�`������H���q �Z��N:�= �[�E�4���H'���i� �]�fiz��e=��9�*�"Ǩ�����]�~����&+0H�� ��v��H9�/���]�.�e��f��Rp1�l����Pc�����kj����.J�|�^��N7�j��Uɋ��V��Y��>]+�X�)�է�yY��̿
\=eіxPb���(���*{_���YL�`]�Ik��I���\�p�d���X5��)�n���x��t&!��kҰ]��%`�*�K�/�yɋ�óX��ϖ��n����d��B��<��Ia�D�q9E����j�t]׸3���"ze�9{� �����<�{�Jm�8L�&�] ��ku_
X�>�,I\���cIZ	�n6����@!�0�sT?�+A��dg�sY�U��/��?|]�0e)��r��3�wiU�G�5�B�/8 ;}���kݗ�*2(TN��-r�Ǚz��ȥ��z|�ȦӍ��݀rZ�,�&���6��-u-���E�ի����3m|i�"�@��t�C�vIp%��~p(55�E�P�ڣWk;ŀ�.Ѕ��(��|��������O�
�sr[�e�,�]��[�6E
H9�U���Jl+�\�`+n������3	Ȱ��s�.���R �k����� ��y�0+۴u��<ec��Y�ޙC�!|�_$����[[ ��r�;����Y��O�\?��S&z�O� �j&[��+Y4�0�S�����,:7(�VDgu��� B.��MF�xm�dc��)����'6&��G�z
H���UҠ
�lK#*rfC"�ܻ�lئf�"2Q�oKB��fq�$��d1$������h���3�O	/��]vN!�cn)�H�]&Q�3=7\H	�>��y�w��"*Z��~޸��|ƚ����Qp�>\J�̯F��a;�G�F�R:6{ogV�Q�D�ቭ�M����s1�P�%�W�5��c M�N�}*�q=����b`���mv��3;My���k��\���k�:_
�PH��=��z���i�q��j�[��0���TT
��u�0���VF`�tnd�&G8�����g?�wc	o�%�E/�K8vFX�7�>{U2�8�T��u�4���X%J�?��%�"�BRDT4j����ӌ�K<YbZ}�XBn�Y�L耿�,dڲU��F�: 4
z[P!ғV)�$��#��Q4ba��Թ ݊�:�ϭ�u��!�8@]��R"���C���`��Ga����U�z霹�:&b���ґq���=5ȓS�rw2v�e}��c���`�ƀ�S��뒤2�;}���?�B>�v�ņ8L��Ԅ\b�D�'�ƀ���]�D �t|�/)Rc[���DI�₠�z	�lT��w�i��V��2i\�%}py��7f͋���3d��f����Ʋ^���qxuՔQp��HgH���/���m?�Q�Js	G���8��.("g��e��I+#6���(�(|��WO��*�������bk�^���XN�x�� 3נ"F�^�g��PQj����~�ص�8}x�zya汆ّ��VP��P�ȝ୊<_4�x�~4X��G���*=Z�(Ɋ�]˼e=o<��h�y��he
�
[>?d1��dǴ^D��M�E,�&3���x�R�?Qb�8�2�ֱ�����㨠2-cD':ϑ��{�߀�3O�<�!\j��ۯ;J�V�� *�:6w�v3�X�LdU�ޟ+��]��o�� k[r*��\�/�U���,�+��(.H�dz�YF�ÕyPj��i��,�1ɸI��W~��"�iKR���>��1��Cw{VV��$��ޥArsY�����4��������.�p"Vڞ���6ĈcG�<b
�5=ը�>�(���:tiDb�N�����̓���v��J Y��"9�pD:�� r�K:Gf.�d �GF�!n�%�����5�:��F3D[�c�ƙovtr�RF��1A�ڜXaDZ{��:��</����ʚA>�j90�t� "�� ���
Ҵu`15��w� ���(�{��>��"w	S���e����#Ҩod� cn��ʫc����x��<��X@������t$T��+���~r�s��@FvVFj��BAm�A��R�&��SL0%
��[�@�Y�j�r����b�n�0�&��_�����#�(���n:�A�~�}��pG���Z;�0Õi�7���_�Y��[J�.�ր��>�O>3��}�.'�fRn�j0����I��S��ewP�@n ;����I;y�����8��޲ SW|oN�{㌲Q޵@�K�g:�LJ���Ph*`0���j��/���%�W�H�g�������r���D<����e�<ط�+5Y�A�l��uK{��Ш̖���
$Ar���h�9�w�60aI��ѽ�(�*�)��d�i�5y�j��N��"�m��h.o���&�� u^��`s_I��[�\A!^�1�x*�DO�^�0����ɃU� ����^�����v�v��d�N�������289�vɦZ,P�3}��sB�[/�Z����u.}�`��+P+��QBbqP+/�]ꡨV̰R\L9������2ߌBъˆ�#<pl�!�����͌g�;%�J{��;'�׳x��K�T�����B]m
���c �P�Z
X $J�FJX<���p�hR�䍯�t�yī�"��ba�Jv�D�w�2��(�ź��@�g��+�!S�pKR�WrI���E�y��bՉ h�a�P�g�IO�6��6՘ߖ���r?t�Q4���~��������KQst�G�0������ڃF>7$$�=2�MQ���61���������3s�;΂�Q#����V�\ɂ;�����E,��`���hh����"�Vh�a���/���Y+â �u��%w��<��M؝z��m!��dP`C�hm)��G=�b��T��3dð��� �D�<_�ҟ�����O6ɂ^��H����yۺ��c������")+�Ul��"���V���u��yK_y�Ļyt��?��X.�D5H��5������f���09G,D����l�V��V�3���g#j���Fv��"V��� D	�(!���l_��`��p����i���ܱ1�H�P:�9��/˱J%��}��b�Y�T)����õ�����
��\Q�<gm�9�cr5�m��o|�~���5����.`Z?�L8����i{�37�2{^����m�o"��w��҅����t��
�@����;T���jT��ɠ�����;M���fȇ_�~�I��x�fEG&�p
�^O���8�\��D#��=7�Qf��*wU���,�����,g�����H�k9%��Aq�I�cO��i9TY�\�Wi��˷f���v�s�眘�"Y@}UA%ƀ�UKD�Ȕm&҅OtJ��&�}˝�;��=Οf�b��ԚW��*m)϶N���~Y
W�K����$�>"x�?B��㾱E�GDG7�p���s�m�v�ct�}y�:�����ߓD��+�6zh��,ڇ�z�+h�7�$Ұ�B�V�%.�O����m]���&h0#آ��G�1�b�;y���!b;��g���8��zR��=K#$�8Kv�q#:n� ��:5�G���5$��J��4��t���8�QBN��;t�;���e������8�L%����-?Ɋ�b�w��r4ٴ}��
����{"�_�|6�K �	g.\� �d�c��/c��Q@~�r�Y��%�Ka�����N�������\��\�`ZNR3����դ��PL/@��z��tF�3;�w#��@�F��~��u��$�:�8c��^՛Z�Q�J��LDN\V� ������tc l��p[Дa (vnL#m��'�X.�B�H
��~�%���]�u��7��X�{����M|G����I>c���+�;���\Pm��u��-@̲��i)R�w����M�$������T;�OA V���C��K� �w��%t,�ࢳ�J`I�Oܔ�Gi�"�?<�1�ػ�p���K�,M������\����Һ2�)v�h�(yf���ʉzl��_����'+����N0+�H��U�+yw�"Su�����U]<1����;O�,i����X���v�F�u�.��`��FEE�s���