��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbơ&����/�
R�A��$Mf�s���/*�9����+�Iy	�E$!\���j���*�F�53�5{����z��3���h��B��XO����c"��r�v����q�Po��������:�-�DC�]Eam��q��ma"�������Ƙ�rW�[��r���⏸/7�'n����tG�����Ě���mo��Y��V��)��6׻\�p%i��NvjP��iC_����i)�}TZ��ҚӆmkvG�2۩�J�{iU�oI^�^��� ���A�f���a�k^o�*pz���tDT$;�̉Xg��<R��Rg}��g"�?�[}q��q�0��Sr����C)�C`�1�!2F��@T�=����B�<�,f��>K�9��ϥ�X�mr�7����6�I(�LVIRn[?�]���lC��m�Bàp���?o��(`��Pc��W24{V�P�$�%�9�)SQrQul_����J7���;ɞ����X$o�6h-�E�zl����])_��}"��K��)a0��	>rLG�&��k��k�����I���>Վ��`�$���	WK�m�F�����Z1�������ĥ<����".��Y��l^s��`�哪�S@��g'aᲙ�d��هM�X�Ǹݕ�iZ��lJ��V� E�Lio���`w��!�Y��c�y)8F9����sy%�����d2bX!���&{�
Y�%�	q[1��H�u%��n��GQ��Tn<?V���͗�XY�&�����us�l��3�E��]-�}� �C�٧��g�mXCr%�q��7w�!�>h����z����.듮����r�E�����D�_�i\)`\���oȈ��y�	L�K �'�r��gM�����ۼ	"��z�q��d��G�N,���2�S�hI(�a������-s�d$T���;�7&���N��S�Q�~�Q#9=�~<#C_߼[�f��;K����*�4�N��[|��
�8�7�;�-�i['���+~���A���wԛ��nͲE���
7��J�yZ����=o�F�gꑲ��$���B[�v�.U��#����y�ʗ�j,�2C�N�љ�t��S���6Q��1P���'� ,�{q/��+|����t�`(��\�Nd�!�Ш���0�v*|?t�{V�;g�?�g)r&��`�ɉ�̌�5%j�	�Y%���Z�A�(�d]���+�q������G�U��0qh�W�����C�?�X���~ ¦pڗCG#gB��aD_:K�)�g'y�5@�R��el⿨�gx�6�.eSx��0�@�r$3�s
b��_͵��Fh��_}���NQ��H�nO���縖�s���T�>��	�̀�RE�<;�����&�Ē
C�Q��ɒ,�J^Q�����d�PO�sez-\s^u���|��G�����V!�p��c1��8��Y���7�n�<꓈*��J��*�  Ȳ�oF���kv��Cf?bq9W�����`��.�>!�i��wA�����mo�h��L"��sд�b��̪^6��}�|H��%P4��8&oǱ��D��2ֺox)�$q�~f��%�_]��t�r"�S�<6�M����f(����@�`wAk�ŏ1�6���05�����y=ݏ��,4D�l����M	.��I���?_�ІT-7�d�7�r�%�T�&U7�� *������/ha�C�nyqlE��v\�Z��S����ۙdWK�h����V8j�0�b���ҞF��M�R�\.�.�]l�xhO��ط�.C{�"��K��/�-#�%6��"gG�E����@&��ٴ���#��ռ���S���vђ��>���W�˟��o����iB��N�����>a�K_�u�+�f�E��z��@T�Y���i�3�)����Y��V�n��4���Qb�jL{.�S�U�#�k�{����}�m)F6��,��k"m�ȕ꺔�<����@�I����sيx�S���1�GIā���_��ѩ7��������O	�=�d��vd �=hDJR�,��EC]P_?��DoH�	B�l�6��Y�9h(+�����?��l-z��-Q�+��g�.v�ņv^p�O�A��M�؋=m�g���Qz1�d��r����(�MƂ~ڡ��;O���y�7�VfnB��<F�6���������>w	WX9���)�v9F��1�]�I4h��:�{W�k���N#���G�q,���(N*�\kgjF7V>n�l���|�}:L����TP+kH�o{ �l!���!�ek]��"��� GB8���[[�'*��A�?�uy�CM��g� ������Z�,��&����)	�g:�Ƃ�E�}�ѻ���6bNy�6C+�T��]�_U8|>-��i��=ɨ�^A�UҖ@���g��a�p^�J�iԫ���OQ��P�.õ%,���B�*��$���L�yܐī��hֲ���yZ�zv�
nhV��TpN9U���fQ����߉���<ɺ��������c},~�_kk!�~,��('��������&�D� �wݐM#$��֩��B�D�NU��yj*i,��J��ր����1�X4���%�8|i4��k�^E�J&��S��{��\�s�ͯ��I3�d���Q�^zs��'���k!c�Jt	�zF�ԃ]�?6l�T��a}���
<��l��+�y��	�+�m)�A�D�qZ��K�}s�wS�[�j���(K_zW�R�T�j�/cRs���t8���i(�1�X�`��Gih@�;�t�,��q�k��F�ıu$+��'p@�����@��y�`��1�O<9�S]p=	c�������.کT���Q��c+?3-kMXDj�Ӯ/��')���t&�rМ�_�FP����_��JBw$�,��^B$W�����%jy�$�޼�e��k��G@w�}��Lf�k����q�����C8��Ŭ&
�v�&�8�7[��[5�#WeN��b��>���o�J���%� -0�Lw��{Y��?:+�mjy��9-��JW��M����F��o�^d_ۿy�ۅ�g/9V�3I���1��%�G���\�Ⱦ~�1J���R�ad��c_d����6�ym}=��I��B[qS�a�@�#��r[V�	8��N�U�d鹆ٻ��(�� ~e�ODq�ٞ���ʵ'7�<�pT�I��g+>Y��4���M�a��o�N���x��Rm�obY�,��:*�of��T�����B-�j+��X�����0�D/�s�uF{�@:`��4,W��ߥ�]Wqq0�]����}�"K��s������A�{��a§\3���.o?⧞`���!c�F\�<��vb�쳂���h�P=to�45Q�A=�s�K�и��X��lA'Kr����з&#ԶM�&���;���S��>�/R����*f�Ƣr��#��d��H����d;�^��mأ:n�zV�%%"Z���9���.XM� ����[C%xj�Qʴ9}�IeCwF�G9��7J׋85�oQb�H1x�/�>c7'��i�|SZ���]�@����o�GK�8(w�JFͣe��:����Ƿ��{�ɮ�	A�Q�rv:)���D��`C�cCp�>1�R	`����b|�0x&8��U���:U�R\��ϲL���l���~P��a��j��XCm�۪s�g�1��>c�!��		��]���i�)<�E�~F��j��0M���F'n�3^�3^ծ�a���$o4q�i�R�w8Tg�s@���ہ�����^8?\F����^$�χ��)�Et��n8�������u���8���9��D%�KZ�.#
"g��╒F�Pw�ճ�[�Ch��1S�8)7�p9�`�W�o"
�(�o��F̵�ax�D�g�����ms��Pg���>�߶����ǼE��?���L0��ϋ���oi�2���]���q�<D�,G>KGҍJ����&��= g^C-���Q��Y�! �ȉwBx5s��E����}ɾ���y�l.��:�vN@��e#�.�V�|g��X��~�� n3-��*��q�c�6#��g�� ��� ȤƑ�?���G��^{)ڈ�,nAl���[��貧"d�z(9�3�9��7&��?�),�ۺr�ݕ0����m�@����ݣ��(�-�iy��I6r�(�&�1���=pi��=j����c��(��ނjdBu�銫[q��/��kC�/���M��k��Mv4�Կ���l�AЖ����$�Kp�"�������Ƌ������Z��-
p�i���u�n-*<��9&�up��~%ou�U;�BkS[�u$}]/�Pwl<���ʯ���p��-v��YEG��{��$�|Nǯ�����<l�(V������_� %�0j]WRTx~�m��G��t"�(a-g��n��oP����>%-��Qu�NEXc����ZI���	B�.���
�� ǻ6���a����@^�����Ɓ�1a��i����0��"}�A����)���S�G���i�����=JrA�[d�7�D�Qe},��4���iP/@=��XHmw�1X�W��I2�m�m䨂F:�;������5��fE_!�R�!J�!��	0�(�V y�>ɰ��7���>Q2��K1��n�5m�����R7�hρ�,��X�-��(9��#/V��2�Ρo���������għ�	��v�|0=VL �.b�%z�� ����$�%����O'|�dp�'C�{)A~���b��٫�3e��P�Dܓ�/�%;�"���}�������B��ʃ��>t����F%E��o]���&��S�7~�_&A��62�/u|��ʤ<��f��A� �G�������S7�|$�v��5��v�c�Sh��y��T�q�S�z���+ɦC*�������. Z�xz!��:�Ǭo��p���	��EQ�6��K(A�&���WIn�{6��c�5-+�e�o�e��Q�~��J��Y�F��ۧ���C:[=qᦀT�-�|�]	B\��X⃧����a;�k�{i��T_������p�4q���Sqw+V�O"���~=�A퇡SA�r��cY��5���[����r�d}p\��@�V���(� m$u)��]�[|k,+2�弃�0#��|�o0�Z��o�EHZ}�oOdC�l��P����5�},�sKY�K�j4ƵZ&`�S�ȭ�Xn=�/o,�w$>XcS����N�|2�G$�[2���;e�5�p���N�y�q_���ȫ��O�����\9���M�;��K�* ʎ0tD�;�G�I�}�`tcyn`}r@�������צ^O/o�w�*+"<�%��!^�\���~�12yOP�e��'1�P6�;*�1�
����v�!�{o��p���:��h�u�M�6n��7����T<�K,�nڹH�r�Q7%@�Sض�,q@gJ3��i����%
�T����
��X%~�\�"�g�<�L���Do�ψ�\/<h�s��&��[!sd1�M}�؀Tݪ�7۬jq���a����KNc��!�7��.��H�����I���=l��4�hU�&�7�fD�?�?|�v��[Y��D��鏯|9�nI=�Ձ)CS�Z�Z-��� a����Xr����ɑ'�t:����gJ����5L�f�A�TI$�05�PB�����"��H"]�V+����я�V�|�/��2��@�ށqb�h%*DՂ^ P3z�ӏ
M�$�� ���9�Y�te�C�(H��FO�䳈���N3��ǃ�Ax����o��Z��A �v/ӕ7�r�jI{?��	�_��[�jPTݚ-���}J�T����7V:K*;e�6�}�}�� {�JC�X���_���_Wg�/��4�Wx�q�-Rr��T�l.�Eh!��ɂi�S��]e޶�B��_2�]יI�5B��G�b�V�����[����T͗��I^�9� 
j$H��6��60�e���v����{���r��%p<�mK�5I�w~�v��� �[��^XOޙ/��9|��E�o�]�@Aa��]�<j�U�KU)e���Z�l3�U���]�#+_�ɹK���'�����*��/���1d���->��}NKA,dy ��&w��j��۰<�^:Ș 0�&;��ĉe���ޱȉ2���i�f�O�սb���L���ө�0�߱>�hOsQ?��5r\'_s�M	����6�י,�R%~��B���"�ߔ�6��Fgw�ᄤ�	\����y�3`���X��JIAZO!GZ�t۞8��A��������F(^�Zh3���oZ�FG��2�/�P��A����N}ԛ۳��1ɂ�[����s ���,��j�ܢ���Ւ�Wi�<C�O��X��v��*�����&�l��k�^�r���[$�r�us?	�(�����4�*\�HN�P�m%���C��Os��m��h.
�#����O}�$����f�1����e�ׯ���1w�+%����b�rt�h��wA�C^��� L봘sf`LT.�M�X�h`������С���������0^?��G�*ƛ�H����P+����eqAP�����ω�<}ʧ�6��
&�e�K��oڒ.9���y>�I	R�a�"�� ;���+)w�6b=" ;��,���*��L3Y-��"�f� m�QKȟl��VK���Կ��e�Su���O���@%��Â Z�[e��}�G��uyRی������%bz��J��{[\��1,Se�m�f����B��3z����qg���)s�Q �?<�x�/[4�:´�Ϗ��"����O�/�v.��'A�SWG�r�".^�#.�]5��d~S�Tpp�I��M���t�8��4Q�n��1i<)�m&��q�[��v
��4X1�:9N�]CѢ��+�{��E�����D[�JIL
�ͲXQ�����-��"��F�(�耶���_�|��? �4���GO��I�I�Dε�OJ�h1�E�nϬl2JK�ΫP���$�
pe_J��ܨ.��(Bj�f��P��,�'��T���Iig �NY��V�ҞЙ_;R���7I9cT�����u�;�#�°�<dqi��8s�p�:�e�F����:+3^��}!�Đ�k�߆FQ������{��ɶ_��z� ć3^�)��Ǳl.�CYZ.@�gnA��� `��t)S\��p���� �|�L����e7&���H��cESԎЪ5�/�	���(�Il^9�|���{s�:�U���,ZY�#-�rދ���#x^���$��k	ƾ;�6�	��>�	�}��@�'����i�5�h7�)�ˤ_'�q��"}x�XU����PӘ��r�g!�7���Q�S<x��}�" ��:颰�9r,�u߰R��6+T��w��}S���ȡh�ҍ�cG�Qnp�XM��UN֣9F��:ep��vp�������{���)H8��!����n���`�lVQ�r�| ؊�k���ߜ�A=9dŇdER��y�I~�5�^�	�U�JxC-����P�2	ؽG�cG��^Dp��.-Ԑ���<����^ I��,T�M��l�0�A-`�Q�_IHn��Y��M~l)h%�t�ODTH<ft-jŎ���df�?�;�A�>v�a��0�)l 0
���uT��y�N7j|�u�O��G�f�R@d�� �2�4�\-�#�eo�f4�����
�[9S���c���nq��DwA�i�<��J�%M��N�6�(*�`�Į�׵@XA`r���-SQ��R����#�TH4�ר];�0��Tϐ�����@�9`{�\�.D�ʃ��BZ�e	Sv��L�I�d�l��]�<���0CU����b�� ��(�~�t2:ȮpMN�]�r��6a���!,|��	�/NA�x���YUI�#*Pμ�]TJ@�B �����������.���a���/֋�w
y���=����kB�T#���:%���m����t�����	���f��8�`��"�uE|�vA�r��s���n���SR�Lƫ|>2�
�_]�=:ӥ��@�@�X����Ʈz��j��>�e�����$(��OG6ӾWs�#��O%h#�w�[c�J��_�� �@}�uE�RQ��_R�-ߡ7B��y���
�>{ƛW�(��-��Y[����!���"���Q䶵��|����s2�@�Ĺ�݁L�2p��-Akj�ٸ�+z�nG«�*B&�'�р��$8�/��Y����M�oBr�r��	U�Z����S�����"d�ɋ#��'��9���М ����aO<�GYa42AE�zS#��sf%y���ES��i+�?����b���ğY	�i)�����L�e:�MH_-S�A���ߡj�P�����u]P_G}:hՌ ��"�ݚ�.,5�lo~P���0�/���_�����!��zɯ�fFoD��S��eǌ"��d9n�-�c�u�)K�u`��:�@��+�i�`�?�7D�W;��a8�7��'o|�x����o�V��^_��I>������KꉽAw���!�BPk78�[F��"~LY�����U��r�g���3	V�^0������4�T37*1v�5�����)-���H�|z/q�nUO�8����7�����z�3a�t��dϿ�23(�B��*���Ͳ˔c����p�n�B@��:y9���N�"��=��w�ZM�
�}T`��d�>�q\JY󹠿�頪X�W辶���cc5#M���~XVi���w�f��*��������; �J �C딻y <ĥh�^��t#QF��d���\�4HvU�����MfF�r�H֟�F9���9<&1  Y����7���	�o�|�űK(:�~��3�m�C��vQ��}�Y��h���+�� ?��.σ6m_b>b  ��h�	�0l�3�&����:.1૜���)�]R�XJf �~7w���#c�,����ɬf��ֹI���y�6�N<L�ە�g��1ٹ���>��I`~J�~ޮvl��`O�E��P�~ʚ���|�.u���HS������3ȱW�6��l�b!�J���"��!g�.ø^4��V/�L��Lw�G8����7������5n����
��Qb��Fhj~C�C=�~�?L:(%�+�d��,8l�)�
�D��Y�.��P@�~��/�H.����L�7`W*����7���D��]J�,lѼ0��Z��j5�%A�u����	�����{��^:��2{�5����ti�0@�酕j�B �k�p��	��׊�tJ�O	!)��m�|<�O_1�+���-�(�M����C�B���c��(2�0s�20�Z�*��)B�H�2�^��2�D���j��R~
���F5M���+�<wU�[FB/��ʠ���tg�*�p�Z�4�l�J��2��u���誨a��N�K��'k,i�$D�#w3�FyL܃�� fC�=�>^��
��x^�J�	ȢQ��PF>y%l!���޶�!4�`���v��#��m*زťt9I!84
���*r�J�>Pd��z�;�AW&�n������(�Yb`��zCԠ��/i��$~��A��,�i��i�	����|�d�S{��,q}�L� �p�ڧN͸��앻ܳce^n@e���J;��r�կ��3�S����wb��:�� ���Х&0��e�z_4��	���mnܠ9� 7��¢[��)�̓�i�V�l!_�\T��M��M�Ei+���M��|��m�/3�/�<�������ϑx��j�D�a�h�����`��ϝDd��,��X0�߇�}%����z��8Y�&�t��p8�E���+�6'ZD��87�(�p}Q��&fa��{��?h �ʏ:n�L���k��$�:��`l$C�����8�k��
�_c�yc�E_?#o�b`���b�~N}H�� �G}�%��Ks���a��s+���ʼ�����R�}���2����"�I�]R��Յ+���g	$z��Ot�-(&���Wn|C������U}֥�_t�F �b�aY�\�B�0M���Q�O	7�����gX�P�9���G Aь��&�.�ہ�� 5��Ĉ��uK�����o�*"��
���E�t�s���\|vgo��T(i�g5% �==%�VJ�R�]�M��I�qvT�>���NQ[,�2q���CN�=�;����#����_��g}Vd��r�7a1�p���*�Jx���yQ�%���ڈH���x������������S���Om{���&�����5�;�y���j�ڣ�U�t��&>e@�.Q�<;!Q��o�^F�����lغ�̅E<*^�E��ܴ#=��
���kϳu�����m
3�� `b_3���D߶���9�6�KnYB/*iư�ݢ�0���
aH��=>���*'c�5�0i�pmE�L�<NW����Z�O[/���ew����d�7{"X���]S�:�Ƭ�O���\��Rh��(�)v@�k�kCU,�֝4�F5��3!L4M��=�L([y���B�p6����$�l��a���!܎��L�%N�H�.�d|����骶/�=��2�DK���	��o��{���~Q�31�3�����Ԧh��̇�PĄMa
h��|%�~S���ת����0�p��fk�t�B����<6��[0#K䋉.E&��#=�8��^a�F_�Ӡa�7o�ѽ��>�T;/ i�� �hn��� m��u]��V���ڂN79�,T�!�&-�ʀ��/�+�m�
8�
�`?��ޗ7��;�n��n��J��t*�����S�V�l|�g~+�Rd��_3�~� eĉ���-n�p/׎�DP�x���>E���:���ͮ�R�O�h��u�4�E���4���S)�t�1���f�?\:� �5���}Cv��lV�F�H 
�.��*O�J�~��f)����Fz�U��K��$���8v�B�L��j=R�20�p���!�=�7J���K����0��_%����c� ��)���Y�Q�����
��y��m%���Ԏ��b��x2��߂���!��Yw �uo�L����t��4S�A=7��N�q�O�$rK���{U���Y뇞��U����&�-<Qt�XG�KZ|�"�����ÍE ��:5 �n	aX'!i9��]y�\~��K�Z&�.��(��.�uC�z�~ǘ��r�v�GͯcT��g���7(M�m1�gO$�c;~J�Z0�%'!P�3�DWWhpzVM0f�nG�o�0��z+����wX3�ͅ�7��+�	����͏������=�)�W�%PL��:�a�=,xEb:��~�m{�n�	�lHy}������oQ���Y96[|cLB�4<�z6�1��8$�ьY{�}X̄���L���<*HJ�R2�^Dh���|*�pT?:�ŉ�tjR�Z���wo0�h����	в���v��3&��p�a@���vY��[+��ϮM��c]����+�܉e�L��'*�Q�i�S�r��IY=�$W��V�����F����~�Rv������1����Z�A�����s�����A��`���2�/[Ms�ww�h�a���5$�g�@���td�	��[+d���0����e��A��E��D´y$��
�������GX����F-5pK�o4��p�$D�Ȇ�_u]^��n*��Q�+L<�h+ʮ�$@!�8���ʂU�S�Ln��@�����qZ�P�ھ�D�� �Pz7���N��X���ɺ��c*+�y���`�����|��]5��s�cŔ�	Gk��\<K,�pĶ��[�+G�[0�C!�.�lѢ�����Yp�V`���Q�$��fu�tHa����Bp�0Rb@�	޸�Z�s�p$��׾�7熅*�2��Z).3�M�sX�w(�ClO�g`R^��b�vц���J'����f��� ������v_��/\���/O��. ����.���lQMo闢�>`9�VZ�4]C�������
e�O���N䖀a������N^_-Z���ꪸj/�ɔ���[`�4ۡk,�g;pE�* ���&t[j'�G5��-�d�X�N�H���s7�ۇ@�Z�>o���D3j�C#E��$��W�˨��V�2��ʶ�'�wR��p����L���R����_*���`
�閖J+�Ʃ�jn�����g�O	M����;bg��-
��V������S�zW#���ѫ�2���ܥ�w��}�Y�����*ٛ�~��2�«��3@�M�E4ǣ�p�:�m�Zl�<�dL�@����Y����A���Q�r��Q�ƨJ�-k���3!e��-ae�T+�~��8v}��� _E��VoS4�nJ��-���QOn��AY�o���O��dVj�&�fv�(;�@g>� v������$}�*5���v�֖mdѶ  ��&	��u�\\L�^9s]��9;'{���?��O��Z�Iuv���R��N�/�-e�~Y�ƒMNI\	��PR�5�4̥h[Pe���:�c���8����j:|���ϔ�y�k�m��@0Xz�*A����p��%������GUN
{9��^����r�]�M�wx-wa#bA!��k���/� ��y����oY� ���agB�������e�_��*9v��#��ֺ�1v���B2��~1��%e9+)����b�K"�
�)�����o�KU[����p'A��xծ�U��.��_�����W��
vk��ܜh�%�a�ߛ�K�N#�q��͘$�/4�Y�fH�|���_.|�'�y�����k_�uFTBņ6��S殅�I=أ�- ��7a�"��o��$����O�h�u,�o�	kO���;W#};(P�r)��� &��ފ_A��T�Wg=;��C�\��<Q¿�*�9�Gp7e���q�H��,�ܗZ5�^���67_<�c��3~��f\���w=�])��	�~`��_=C���*�Ŝ��1޽ݜ����߰�Bֲx)F5��2��CA�����-9.�)t�Ĝ��h�΁ݧ$W�����L���j������,!������	.ӠHz�?��5��r�)e�2o�E�z�y�xny��^+"BR7�$���fClKY��w�o'$�?z�f�
R޳~�E�&`������+S8�{�Z��b�Ecr�~Ҩp5�b�i'l�DlSs\o�;r�X��o�`ʈp=�\h|Q��x���(����U������+���$�#&���H #݃����آs�](:*2�N#ׇ���R� \��x<��z�ҋ#�f�M�M�Aʠ��Ω��[ƚzvp�X��RJ�7����h����N2"QL��ۄ\TY��$�~bd9<��/;1���4����-[�iY�O�M���i�"�����7�`|1.� �w�s(J�(8N\��3�?�]�5w�)��L����,�b�S�F�K� ��^D{̓���T�ɂ:�2AMJ ��(�la�95�'��e��^�!Q��AQ/�g`<<!X�X==��������39������\�29}L/�ɋF�����~�\D:���Uj�����t<2�k_I�����'�6���=M����z�ױ� ^�ه�PN��AU�o�U88�bRj�1���A�
,(������+v�t��@>ܧ��#��g�{���		��`z�RI�^,÷%��-�lR~��]��z��:�A�*�A�X!o$���T�xW���.Z��i��f��7����r��0H�D�V��Z]sv�U 7�{�S����J�gwˀ�[���o~Wo��qnH�J��D��I�w��B%�zfh�X[m���Rf��G�Ɂ�'e
RSGON�]@�����9Jq�B�V_g8 ?~r�9s��?ҕd=��c�{�+hS���4 4���k"@���ː#���j�-��Y�n�G�����ѧ�>spЍ]!o!bjܢ��Å������c^m|8�U�e[�_1���@�}��>Ra��kG7�~�4���Z�y���Us�k.:�3��k������k���``����3v�-��BW�¤O��d�>t��r X�.�Qö������Y[Յ=i�9����jb���[.[�5�c��[��.���gR� B����j
d/�xԌpeAAr~�]_r�x�f���+��&��r��o��8���^ R12�r�y,�ճ��\�\�{@F�e\,�#E/n�%С��lD.��~	2A� Z�|^�匿��y[��h��&�C�����/lO�凓	"�>.�������8��?�a���c���y��A�A���C���V^�,{����*�4�q����!���;�#N�Լ���0����c�cX����lFy*��,.ŝ_���*�TEdÐ��[+e�^�PX9����|�v�����4�6�I�tWJ����9���1�kC��T�v�y�R�� ��W����U���	���EŚ�ۃ�(�I;���,�V����p�It����!�(!p ����lg3�V�E�_S��$�.�mS��e&P~�=l��$�>Į}�>�q��R����v��f��"4#`pW��$�N-u���͓(�iJ^�������G�;�C�H�����^���0c
ޝ�\&�J��l��]�+�^#_2��z�t9�P����������#-�������`͞���;G5ȕaҟ�XE1�)��6����0����.)W2�z���Ⱦ˾rLG^d^R]�	 �Տ��b1�6݂��
ǉ���~k���h�\�"?� 4 ��m�ݿ����r���O$��-�#��@-��h��\���OIC[~�r�y��#\S��������EE���n~�H��+�Ʀ8ދV��a�<��$�\mv�w�B�栎1���-��=�ǋk�D,���SU�ٵ6Z2Ba�D���
ցd
"��=�k:�]d�O�44HKc����Z�A�4Ə��b����`�Gs9���M���_q�5�1ـMa����3���h�`\�r�jط���~PE�~HO��6�'ϛ����Ľ���P���6̯I���l���ΰ\��u�<G�8A.��3�P��V��hDb(� ��@4�u���$4�9�k����4��U�ϹvI��;��V���5Ķ0~,�9�^�3Cٿ��3���(L�n*@�X���o<z�7�L3	t�lP_P©��a�M�I��>w�j.�@����?���
���3�xHutQ���.�xdu�hǦO��L"ː�k&=�~��f�)���ҷ)���t� }�Ly����J�!����m��ڢ�sD���f{ޜ9ۆ���d5��E�s k�x.�*��fp���-�c�����l��7�U�������k\�f~A�!�5w���4��.�/"�B94(�����Z��e�����k��5�w�Q� ���� ���h��j�K���:�(��rue�V8�_R(Br�ZOJ*�	�
K0ok��0 uw���*�en1	>��k��򠯧I{Ȋ a��GoԳ
��oڧ7����F�h�7lx�)���v�b�����)�����I*#�<Ƭ���o�Ȩ���8�W���o�B�Ʀ����0d�T�a�0D�s�֓)�c�*��uXm�Oΐ>�������L�m>��qT#O���ĥ�Y��ha��ˈ������h����$s�l��y�-���(^ʦ�#@�	����u|�H�Ej�����#��i�<l&�Pm���t�-�~#J�&3�w�����<-j�K�