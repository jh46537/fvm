��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c����}�����°ȣVhX��M�=?o���.@C|�Z�1��i��g��-�5S*#ƪv��8}�*l�>�	�D��xL�kkg5�K8�*�$����)8��(d�Y��j���	�}�d,뭭�.��0�q�����b演��{���Ѓ˧|:^�h.��pz�+5��$>s�P%�kf�f�f�g�@N��dU���HO�ʫA�:T�(cF���3�D{��k̈��S�~��6LΠo�->�u(2��ivW�b�q�*���,3�����y5��A��5�����Ǒ��$�߾�q8?�j��X�B�当Ɏ=.�a���� ��PU6�UyP�����Ɩ�(2 �F7*J#Ea<5F��� !ƷI�p��UG=��m�\)RF�Ņ֭z��f����H��:"�~_���;<��ѯ��y^���q��<u(?� ���9���\aB\m�#2������3�m�������e��P� ����k�b
i�����gL,�l�ސ���	ۀ�4d�+�ZKpV���S�dg�6T�r��})�3�ӑ���<�>�7Ӵ �I�}{������՞�����?6�) 4�
��=���(yڎ`4�0��URH�}�� ��*5�b�>���/M�	c�O@č5Y�]��W��r�ޤ��͑y3�(Qb�x�`Q!s1����ɽ��`�N�3������ln�r�������v;{ �����
toڶ�^��t���O��">�g����ݛ�lڦm�Jv7�k�_mx�{���c\�5o�)�Ȕ�fٽϮ�B�H7�i�����*��, ��̖�������P�0���Zx��S�UE�1�\�v��;�&���}��~=��UHBX�>&@�ǳ����^�ޘ���B6R(��	�Hj���]�&���b�1��<{�R� 8���^����b ��=�󙠺�m�эs��$�==�D�΋<��%C���jcsw�s��ٓ>w:�uF����C�F<8���h�X��,x{��9��P�"F*��H%A���A�����Rn\o�%Y8W�&se���BR4F��s��*�X^뉚��j9l���
�w�M��$F�5
s*z����
��L�`�*����uo|�f���M5jg8_��%�6�J.! �U�VL3�l7�rC��k��[���V_UȬo��b����5��Ҙa�Cԧ�UW۱{�>��˛Q�#4�H�,�ꀑfiyD
��~T�s	�%3�bN��24[,����T&��Z�g��?�o�2�(�68<�zh��6`���b}��h�����\�t"g�b� �%p"U�e6STJ<�vj#��F���
+�U�;3��Kq(���~���m��R#��zĖ~�14O5���3�p�p.�}��i��j�I��|Ex��zg�}K��|�=����p5a\g���R�\�׹@��V�|�:��Do��y����\��s����7�i��0$�Fr���'Imfb���&��륋q��.ƹ@�9��������"��J�-㟀0Y~GX
��]��.0�+�\|����ԑř������L���R^�M�	�E�����nD2x�����ix ��鶹��ܔ΄f��D)a�K����.ם��$Z�)������V��IQCT�g�����A��K̳_��(��FZyq����(�P䵿��
��eL�mU65�l�6�\���1�V�e�h����c,�;�` Ҫ�GCT&�&$<̝M��)��v~kYw/���Ep��S����
u���#_!jT�Q�����	D����$,�)q2��1�.uC^7x��K7kq"�}{�z��F��+�*J6B�lPn����Įa�15�C��۫xp1?������͔�܃�8�Bʪ�v�+,��]������R�4�j����B�}4}�I�(�-#����v�Tp ���9U���==ڏ靷E�h�C���냋D�S��EkHݍOk��_"{�gJw�������{!����E*?��)�<͕4t�x2w�}`ǻ��a#pKˉR�F��f��/2%�w���4��F��4��[M�P�ĬA����@�[BY�0���|�(�h�^v! ��(�0yu��� �D�+|CU��F��\�,��l��x6���Pgl�F�RxV+�TS�Y&08NZٳ����;;���8�S���;S�!�5�XŹ��.r���K�K�:��]��.*S��?���5��K l��P'�����TW���x�3S��_���M�v��|�LPc��KjC|���!:�č�)�uS�f�H�U���p�!�J���&7&k�^�� b����{� v.� #�꜄����z!�F#�C*�J���G����Wmp���x,̠�g�+w����ڻ��"��4��t12�n�����1���8pa��i�S_taJVȇog�-
���������T{7��_�l�4���_���'4\d�?$n~h@t�|c�ɂ(����ƨsv�c�oH�9�.H�ʐM40�a&ĭ�M��K�RF��w�s�������R�;(�J�r�$���,�qV�to�J�v��_�Ϧ#�9qT%���˩��ϻ@����C����{YI{OF��&/�Z9ȸ"���by�y<$)!�������]�B^/�����cϏ�֝F�f�O�>�'�@�C��~!T�k�i�x��`���9��w+����F���=��y?v�uJt0q�ۻ48^bQ�|g���5��#Sh/�������^��8Sg[�Z��'�P0�b��A����!n6��;|^��ۙ�T�@rTd�@50)��y\Q�rY3��u��]��%u��2�$5�zR�����2��Kr�0F��A�Ԏߚ30�QH%v�6�S�Q�U��׹O�H�$���P�C�2��~_��%@4AnK�އ�>�z銘�I���������/������/���.�E;�~�4�Q��]xQ2�9����Jq���lu�ԑ��F��Ǵ�<W�]I5��?�v��T�,�X�&v�_i���z)����k����7���"o�^J���y�p��4��!%4#ȼ���z�&u5��`���h��ġX���iTB�������b�rp]���{b���34u�R�ƴ���f�,s
�J_��^P?��9�eti\�-bS��`/���m3��7ÂEV�^Kt��N��X��|8L(K"oFU��0�_+��!������@���m��a�<�]��>������R�n��Kȯ����_͛�B�V���pb�]�V�F*ǁ�@�j���|��<4�k:��S�x��F�6��X'P��|�T-����ώJ�G�ז���4�ch+xH#�a�F�s%]�npUs�徼��T�3�vNG!�-�4@q��>�p�,1�����D��V�k�T�;��V�)��~j%J���^���+���ҷ>��o&���&�<ߐޑ��Nnv������[vH-b	�0��!��|��u,Ph'K<�>Y�5[�����a�*,���%��<O����es�n�~)8��y�X���GF�b���MT�u$W��f �+tϧ: �5����	�_�q�!�0@���!ϵ��i0.N����)�3�*����wd���с�YE_f�\�����U��%�Fm8�
��wPD�w#K�>��PAZh�[�Q"�.�^9=k)]o�����5����k9��ܛ�܈�p�޸�� ��N!t����T;��"��X�#k�!7'H/'1�r��_�����P��T�Xg�\���yc�@�]�uQ��
ɣ� $�+p�c�"���F�p�X�	T�u[ݧ�l�3I�]��a�i~/��v]&�P79٣#E2M�
V��㧎s%���%�ؿ�4�P��I8c��	��N���jʎ�?a�E�x6�.�^�"�n f,��I��:��褼 ��f�Y��\��`�kV�����(3�8�igXlK��=��I��$n���㫰���zUP�;�G��%�Ylb���Z-���r�tڀ+�_2�D;lF�$� �HB�kܼ[0� ��J���vEe�E}��擋U�����#(�����h����*j?�x����'
�o�bqpЋX�-�eJ��/���H !��Ƶ��I�^�A,ۮ!�t5'����Qf+��fw��j�#ˍ<3�$��h�b)�����g���a�:�s��`���5�4@�%��J֏��u��%!Q�,r��׻W����w���Eav�E��<R,5�b2Y��>xE�ګtJY���'�;H���K;h=/j��Ů�A�F�'c�1]��_^�z�Ҵi�g��e}N�Lt`/2B������'����E|������$��(h��p�I�
<�%���|Gt��s���Z_�j��J�*X,a�eo�36���Ă6:,ïTE�w���p���-9W���^X��z�k�jӵ�5\p��Q,��A���N$e����?X!���Z9�d���c���k|՝�?V�om��,�����˘�����8�:��Y��#�8���7���D_\~�"�ezjJBm
}-t�<�C]�.�e����Ά�������v�\�:����Mj���ED�?�*W�ɺ�D؎�o�<�Ŷ1'@�2����3T���Q��)ޗ�{���2:������$^��F�{�c����1�׉a�L��R�0fϜy�V޻<yC#�=6�VvOW��:�1���X��K�W��j���ܼ)f�jVX3�"�S�\�D`(��	)�XH�n��^-�"�`¥E���yѮdH4"˩`iH�tE3m��Q�
�W�!2�"�Y�9�ۈ_�8��L��+Yc�f�o�$.��G�޶�}#=N޸��%�E-.˵T� �v�W�҅]]�P�Ɵ[�;n�l��ES�h��8((?����f{�gD},�E��
��Bi ������u�r|=�ٗ�&�.|�G�OD�\̊�����ǮT\B������U��mHW��<õ��W�H?�V1��;�8�h�q��L7/����ͼnO��Ԫ�)դr4���=Y��uU������m��g���,�"�%���a�R������+<�,Cc^6&ӑ�z��漹�@@����e{�D��rʢu���~"�X}e4����6���b�|��t�/ ���VF��B�]��3��1�~�����k�@��VP(�'�E��{͖�p�_�x��d��ګ��� 7
�͂��[q�����⤞_��S�0c�#E�5u�%í*�K�猆��X��=-?����S��:a�[b��Iߥ��Q��<7��u�8&���9Rrn����S��޾��|G'p���E�K��=�~`Y�ӓ��\*�����kP���m��ӛL���}�y;yY"��C��]��߲#�X>�c?���+��/T(D�!G�?/