��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]G���B�X�x��x?ь�¿Y���5�1����1�y���E��AjsY�����|v��3Q4%{4��@���y��u��|W:P�ݯ��Qci���Q�z����-�?�a��ǖVxJV����.�����@{����M�G��:���mUjݥ�M�$ļ��%��G�?�jF�ָ���Cht�"������$o�n$���b��JD��.���;�t-�i����n��nn���=�~�|��ۮ���r��[����
��C2��yc�А��6,�ew�U^�����{�
������a��9X�'7\��3�I�rksE�Cf�"��t�8(�IA�'�2�%�}%;�$ xG�XD8�ڣԅ�#�W��+̅c�� ���W�=6���2zq��߲DY��>ho����%� J(rW1��� ��t}�L�4�BRP��<r�KRjV�hy������∑\x�����I�6р�b)~C�I}��Fcz�L(C<-%�W$wX��l{�R�PĔ�R+t���J�9wm��8����;#l&XܵV�uP���ƌ�#l�m�7� ��^�ڊ-?�S|3�S�ϑ�j<i.�r�y����c�@u�ք�ȯ��Llo���Y:".�����LA���o�;}��L��m?��Bx�+����;BM2$�m�j���L�`Q���	�c6����Z�_��9�,�@:��]v@�qj��^g{Ӗ� �62�o��@J��'�)E�!6J����Xmӈ���ƞ�؝��p�}�K�'K[}1xp1ï���6C�9��WÄQg�N%f��]?.�����������h��W�h0{�<2�$[6�
o�w���9�Ҿ�$&cU�\s&Җ!z.�İ��)S�?L�P{��*���Q�%v�j�p?&�X�G�����y�UKMZa�Sbc?�y����4BebZ`��OS��`�5�>�v���ǎV)�{w`�-��\�$��銑'�E�_�Y
�� �@�G�6�޼��	����b�0T���U;p2̅V�拉���r*?�^U�f���|���mNFPv .���`��ŋ�N^.a�*G@��N����ΟC��8OIX`�i���>�uo#��;ES�*\~.��4i����]Xy��wL)��0V-���1zO�����9�tv�����t�����*<q's���G���۴ĭ�LØ{.$vf�st�7�w�������e��Ȩ�:
B"8�$��G�����|�w�����- �G�b���h�Z���zhb��dӭ^:���9(U�W�U����D�{���1\=g�
�wD?�Dt�_�	�L��l&��TNs�OH�����>��/B��YӴ���۸n���>�n�!�\�{W\��}+dݳ�9>אVH{�L2 M�=��v�}/���9�I��'Pt~���D(������CUF�^��B�j#�BM/et�Y[�2C\��Q�b�&��N
{)!�j�q�=�HB�%�l�.X�R-�A�uQ�e%��m��py��6�'��-�P�Mf�V�贿�-Y`�>����۵����A�5)%���Δ��ۑi�ُ�z��T�M��w���B���G-�f,��2�7���಺qND�2�;:k���1��<��\�z^���\�)���q�:i��\k�^Za�R�$�oW�q��|TnTqu.ک���L��A���'Y���S	�w�PK7ey$��-x�OU�Q�sb��̑�7ThJ���Y�aZ���Z��`QLϽ��T>�J���zC���������&�ѣ��yj���ț��3H�A-ܯi�Jd^>���},*{.����A�D"�A��`R�����K lkv�ZY1�oaf����3���22�i�(�j	@*y�U�$8�'B�C*z�	Q�we���
�9���x+��,�
�

��:w��MФD�:_�������^��fo>'�1��l�=h��a�Jq��X{�|��mP���5�/�%N�/S�\ߚ{�^R����������Sp=	+�T�FY�?���n�O�ဪ N9P2v��G���'���h��X�"��֞`)3\&��re��� l���m`3�\KE@{�!�Iӻ�|8L��9Z�����DSr%�k{W���Gq�AHpc@\>�΃g�'*�CP�@\�D���P,��E��+�ﱂZ�����r��=�ް�ْ��s�/���ܹp�Fj�=S!�"�GuHM��)1�"#7z�F5��׫��½���uD���;uW��I�����n��sH�PN��%�	�ɽ��i�`������� 1ӆ��9��h�;��
��̿�\�D��_5�z��=�՚�9�?�����l�e�M���6�wIQ�ف�0�`Vz�a��(�r��I-�zͼ�zJޑ�[Kn ��b/���������ך�������	H����R�*Hnz�ig�n��G{"�戁�Uz��{N(��u�Σ��:�0*�N�s��}[83��^=V�&Q�W4�17���W����Q �4�I�`c�ʗJ�'�u�ѮD�e��*m4�����č��<��~���)��������Z�,��o�'���,�	Z[p��E�,M_��4���OTi-��G�v�G^M@A����9Zt��v@���9�OǀC���`��v��*s��B��&lǑ}�x"��4n/p�e�L.�?$�ı��i��k��[�aK�8Z�d�H6U�ݑ�dU4�V�CJ���cB��ha�lp9��NCٺ4-�&��^'YO|���!%|y]t��y�t�IAt�V`�1s:�j��%�(C�<2���z4Z@�(�ctń�Z@B�u#8e��s�,M�%M�1Cș}�(���lG��c@Q��j��70�_a���hJ�X�F������ �{��!�Y�p��_7 ��D���g���|J�a%�ũ��D�J�`W��e8�D�pGݎ������>() 脅d�XQ��.��ʁH�����ADT���zd��y���(���$!�G:^�L���	HQS�� �z�K]-����s�paŢ�)�F66^$p���A{�g0RG��N�{��=qc|#��E"|F�:�����Ab���@[@	@&��������$�2�"�_�J,��.�s����l+�(�$e��R�0u���3��:�a^a�
� ��zG�
��%�t�Q�AEv�#���|r�+��[�+#�a�W�K���疁���Ujٗ-��=K��|L¶t��H�5��:�b��.����,?7A��VLp!'�߁����\1�_rwג-�����ɺ�
Ɋ�m?O
�|ʀ�e[��CP2O��J�i)ƭ��d3���(c#��S�NH,� IV�.��~��W��-VU��h�%�����k/��KW�-��c �Fw��A��?峞�œ��$�~|��$b�"-N���$lZ�ĭR�n���ZnV֧KѪ�M�J9jxڌ}'���w$x���p�_�L�#τMf�Aۤa9�&��GnG���SEB�}lA�j��&��2�������Z؉l� l�a��`�p-�L��R�_�8�e�	��:-sl=���[{/Ih����T�=��*4\ V1N��tq���П�K�+PصT��PB�&� ze�yo��c\;��]�H,�{��|(P�P�ӣ�Vos}�;�p��O|�=���#E
F�cAֶ��q<�z OE]�~af}�kc��O�����-	cJ̙pɾ��Ӊ��h��8����d�'�$;ZyLQk'��&�pOz򅎤t�G����FJ�_��G?��ѡ �ܧok�Jcf�><�Iz1c����X�hTǝe���f&].��(!�0��ߋ-�
��Sg�8�; T��*Kk�_�VN���N��8����=���R�α�9���%C�Or�!Ng��hj�������#:8����k�����*��D�O=;.k�'<{W��!D��<ik�-
,�co���}�3�x��?1<W��B��h���)�ccxMs�zɎ��2Aү�H�E�Px&���X��b�-v���+]/�:��!�]��N�r��b2�%�R�muV/8�$�ET�KQ�}�Ŕ� ���}������� �P�	���a�I���̱���?�0s��d�;�I`�s���2��_ ����LQD�U���~�|ѥ�Џ�V�9�/S}g���~��a�;|�����I�	��Z�"��v�N3c�l���R7�?.c����1�+��'���8<�H��ڃ��˺43]^u���j�7��Q4j7e��\O"P�pD�^j�0�?�i���B��k2���p2����gFX�1�nf�㳍s?�E^q�8�ã��MG���۟��r3'O�kvBl �k[��)��%
�|t8��4����͍�9�"6�޽7�3PZQ �Ⱥ�D�ö[1x:�RY��z"a~I=��}���y�v6�ëe�]�(+9���6���\��N3�'y�d��ZM�3���ф���J�j
�&�ZNAR��T���������aL簩w,9표�1�W��4��ATn@ի�]��E����{�.F:�Z:+%�QD�Rg �Zp��^�_ug����`)�F��n���~B�O'�n���hĖ(+t� ����L�-�'&�� �4R�����`��Ke��_|�躂����<��r�`�d0�	�z\�F��4�4���X�
nB�v��'���rǃ:����E�Kg׉;���8a�6�|+�	F�6���
� ��P2����{�P�X�O��+9ᄦo����$��6#;(�E&YXLC�8��C�N[�,8���,M�JJ��u�<�;e9���}��L�{����ň@P�-�����%��C*�b'$�OΟѡۡ|��?^��j�E�e�X;Sq^(�-��+Eu}�_��a^IK�-����q��w �Q�6����A�p�y�A�:T�M��cg�����}��6��k�o+:;��f9w5�#ׅ �F�6.,X��d1IgX�w[�x�7�2�}�}��GQIތSlC�Qѐnn���+FO�Mr[���ˮ ��b|����AJNw+��`Z��%>�=T^s���Fع����x��UMV���Sp�̌�6�^�����qi�E0SEz�7d}����8c�t�[���WD��- �Q,���0��!�Q�@��	���o�Hb�J�c���r.Y?��6e��a�f ���u��u�� T�
H�;wN�Z�ib!���}:��^@�!�a�&y�ұ��CO�����ۗ���僓<CD0�e}�2(�o24�2��n�z56�������q�fMZ68U�		6�:���mw����ZɆ�8��)�� ������c�EhYl�l�XǏĬ�.������ҧ���R
�
��Hp_�8Z�@խcUOGy��=k��}��m�v��6�S.|������D��_�VREv1E<N��,3�s�c�8p����@�E�e��Pc��A2Jհtڌ��������H�|���ڠ���5����L�?�'�<�����,ȋ��ߜ��bKz檹�@K�G�s����dV��L4�<��R3��  5�$g|`