��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���Ⓞ,B�$t�{����c�,�-��� k�4�	��[%��B�?���4��\�@e-��� ���u����'᣸߬Hӣmy� q�`L�S�L��-|�,���Ξ�<j�����̨O��f��U�,ﭵ�h���voҭOu���[�)n�g*k�<l��p�l�O
?7�""I�r�<ɫ,�$���?��,�EL�8�	i� ��#�J�Dm?u9CVCI�ji��Ĵ��q��
l����*��%9aI��=we��d�Hn?��sU�����?�KDG�R>�>.�@m"�3 �Q�Z��L��n��kl�z�K��>S�cl����a���׈���NfW��#|T8A%I,���_܏ܩߕ�'�3���^�:WÛ1}R-��^u����
ӭ�cV�l���?�,��d}a�[������~lxTot-i�k�L����z��\V)LL�h:�<��l}�g�z�F������M��0tg��1�Jv����a�Ƥ�>e��m��^����ߞ��YF����@�0�
��^UZ��<���lV?��a�C��;Y�kO�p�#�h��UF�(tdM�W'��D��=���ĸd8_�N�h8�x����S%�k(�\f7�A�&�%�v:��<�}��ל��(�� 4y� ���	tQ���eH���Jv�m�@ɬ�����ؓ�������QP�F�2-ID��Շ.��3I�4t��}-�/�$1���W��/a�Ig�Ôh�q����!�d	FP�,k
�.�yU�'k�u�in\�.<J��0��WMD{�,f�L{Cfx�G�\ۉb%�lh�^�}�d��g��%���{��7E���/m��)#cRM�g�>c�:KO�<����q�� ;�ܯ�X��H��(N�T��2�Ui��p��o+��{�<����$��Q@�@`<���9+�k(��ME��gdl�zq߷S5o9s���
r ��a�>j�k�:L�|�����b�q�]}:o��PA�5椕������A�s�� �.lTH�نk!�5��̿�ʹe�4��Y�N�zG/�	�W�ְ�Xd�d4�4���Ԯ<R��sj�1�\�����t� J�r�|"��ѴƟ'��}q�\U;�Ʃw�9am�n�1����c�F��VG��C"q~���C�Dd���6!�v�A������&iLݪ�C|
I�����N��>|��6�\�8k��^�� $K�9�&aC�7Uڨ�����41 3y,�ճ/�<ֆ�D�&T���N�(<2�����s|"�,�Hǰ�k�F���J;�a8g�׊sr:�'���o�wR�y]V��p�ݙ��逤|8_,=���J0=33v<M�������Q&��ṡRzi�d�`W+�A�h�T���?Q�
�͢�z�GRz�e�@��� �,������v#��o��L�W8<��d�38`�.�\/��g�0Ѱ%c����H�U�0K��-��A!�j\��ؔ��;ll�n��5
�)9�p׼��&�����tS?���)JȰ�*�l*�	�15��7C�Og���t�$!_��MF���o�;?�P�vf,�d��������sY��K6���_�"�<��<��O���k��Ĭ�PJ�(���*΢����Mm�:7���L5�m���������D8�-�����Guwq{�� ��k���_�m��${�,��$!IhBE�2��⓫`���!(/>�!1��|(�:�~
aM��t|J�M��5q`e$�o��"�H�\���>�WJ[ҁg��R�&dFҡ8��@>��Q$:�P��Nq��$���6XUC�T��%���e "S�I�8�Ⓕ��Dͽ{�HT��3Ä�=�����Yt�f0��S�m��5o�a�۝B�EƱ�{��#��*@�Vi�<	i�&�T�@^j���y`�%A���y)�h�b�4t�7�LnN-�h�+>�g:{�v܎L���F�T(���ާ�G�-G�`u�Wf��3!ԇ1���m��	U3%��`4�8���Ooa��y����r�3�C0'����xⷍ>*���$.����J�!��4���TP�:�xDew�|�a����£LB�O	.a�=���I��`�VxQi��8(����S!y�!�n�5@z0g3ܥ8۠܈�;��h����FP*�]�to^��ӕ3n�J5,��NDϑ��I�M�Kf�+Y�dv.ܢ0K�9�w�/�٭9>�zj>x�Q%�H�ʮ������z�Ԇ���nK������evP�C���F����lϠDE��հu�t6��ad�{�� �TF��ݙ�ء��r��������o���irN��ɧ
Ѷ =�
���)>ݾ����6�� ��a.?I-Gt�Y��@c<s���җ� ��UDw���IRr��'fd�*r�,7X%�	�:�k����xq��qV�"�.c-۰:ٳ���Yw�{�n��I�4]�&qv��c�e\?]f�� 18C���6�[Ok��I�m/M���E�f�jt�v'���7���8�V�`~�%`i�J��b�1�y�}6�|��m��U����}�a1*���Z�����������6T0ϋ5�T1k�2"�d��$@/�Lk��ux���Z�/9Wa�(����y��h�DZ9�Qg�j�Z�Nd4��F9g?]�S'`tC�Xa�Y7�7��놢4�i�Լ&��+�F�����ֹ�l�X"��EܟM��7�ԛ��	�G�B_,�J�{1Ϋ*IG�9Ϗ�)���U�p>��!��y��k"I"܆��B�w�� t�ٶ�vݦ؇�$�v\VkQ<�&_X{�u�$P
�N8��cǔ�qno7�,\}̉�'�H�d��Eԝ�7�]S2A��r({��P>D�B���2$�0�w�0βjtt��������{m ��e�*�%��+g.�O����|��!q
�41D̷Äd� ��/�`���<�_q�vj��ln;�S@E_��#���6�s����t��LE���4��ZW~�#ݧiǺ��fR�]ki��Iy[�VI�\�١ɿ��tG���qU�O�s��o�a/��8���}���(H��m]\]k �1����!���<�sB��|�MG����m �4�yC����nc��F�b'�>.�$1�k4~k�M[@y|-SV��ɡ��YCO*��c@�����VZ�
s���@o���I��1`��%����w9R]+j�H��u�9?����.(`3F��Ժ��g\m Rza�}�\���+�wv��z��V��]��b�҄�c��$E�Y�L(Hr��#$��)RreT�������!��ż�B�����F��.��k�,V���������@�'��F`���
IH ��}�=��RM�8OM\�6���� �ct�X�?�_����r��c�Z{ 
�L�lt6�Q��1��G�OD%�U�R���Q#/�@��b��lVS��e�r�Z�rO>4��±�o����ٓ" �ܕ����/����w�W�M�sAْf3�Z��-Av�k�"�s�!^�6�n.���a�q�,0�-���I��A���7<R�w&�N��$��Sq��$�<�$d)[����JzO;'�l\I&�u�Y�,>p�`�%o���N���~�*]��{ �9��伩� ��9���#w��xf�:臎��o��E�f��9�5I����*���ɲU��mH}�؍��I"%n�L�=5n�{!�pj�ڌ��%۟��Wg�ǡ�̥����5�����ʐ��B�U\�{���xX�=4�+���@�i8N�4��Bq$Q1}8h�D p�۶6�t�',q�1��o+�^��ҷ�	^��}OӠ=��_���q�l
�5��N�ٌ��G��l���N]+D9�f��������V��f�H�K���u8��i�`�.`�sx,։L���ML�/����ԕ�80Z8ou��d��Z;�#/���4,�\l��6��,X����!�b�����I��'�D�IR��� ���H|b�H	�-"u|��U8H�&9/0��JU�1���C��V�z$�@=�%'|�
*�`����B-}�Ʉ�Y�ҍp��Q-�����m�g����Ce���d��Fɍiv�s^v�^gk��Us�w�ۀͨ��C*�YA|�}(Gu�h~�J�lQ�в��=Gk:yɌ�~mz⼟��+?���92��?Ì&������l�r�������=@�\���S�Y��5�5���=ɜ����Ii�.�&����fqJ��uB�C̨�(�w�Q��K�#}6�Z$Q�{q���s�f} �U7|�����5d�/W���~ӝ���\�z���4x����h��H��p�2hD�ų%;�1h�}�E�|h��V�l��"ʡN[�#��:�\}��<Ȟ�ឞ�z�;��h��%�"ĕt�f��PM�=�=�N7�����QȰJ����ѿ�Q�*��q�Qr���c��(�UC}��⪡�W0#M�Jt=��E�d���y�]-܉�7�OZ�swA�љ�;,%�|��e���Q��ti��[�O컟a������,(^}`:b�n��ځ���:s���q_���r:M����|c���²���&� 
������3%t>�QR�u�� �w�T�N�������SM:�����٘/¯u�z����{���!+�Zn����-��~a��i�6$��ف�h�5���jI5T����W��U6c9�0�d�¹b���qa,�/髽�b���SZ�1{���He���ch��}_����5^� �����cS�_~K���N>2�/����{Z����I���,P�]ߒ5�5tL(R"�/c�g\h��M(]��D�e�p�w�w0���l�D���	C�r���T�s'̅�aZ��~���`
i>�3GE�򺜯L`Y�C�vN�v�A)�FD��`�4�-~�zdͳ���5[ޫMrQ;����d{��jr�Ed�����U�t$��Z���|�ξNSrZR����
���3W�|L�9�f6��M�q=y����j�^Yx�Nl����[�>��>J�;�^�BA�1��,	.��=���X�����=���j��Y+��+��[��D$�{��#��)�����)S���3�n��-*��!����b�b���r��]B%�,�.;�"lL�Ͻ�/֘�'^VI��*��D����$[�m+��"���e\�ԙ�u��������%[��{�7��	�SH[������Jbܷu�Hg�[i�&F9�5�\�׌M�K<�R�(I����J+dT9�\8�h֡|G{�4�O�p���;��S1�abU~��eŃ�M[���f����tݻA�w�����e��á��5����`�n"־�Dy�}n)��Ȼ\i�|���`^ڻ���a�%�p�.pܕ���icnѰ����$�E@T!?c͹�����(��.dS6��l"lǯ����Ĳ&�o�R{��@0�f�#oXC#�݆k��I�������G(�+2��3��p*������*+v6xE�V�]j��[+����� ��y`MZFS��;���E�	M���o����3ʻ���OiS��� ��/�X�<{��.

8Qó4��\YZ_��2�����̷i�bF���*���o�f{���Y)lbr*E�$�=��i,g�.��8����թ��<8�K|H�j�r�N����	Ⱥ����  "�(\�%��:Ħj�N�6b���d<n�����̪y9���ȥ��헔q�j�e��$���QD;�����H�o9#�[�������=x���쁳���������'Z�pD1�K1BP0��rr������5�ԵQ��/�m�;A��۟O�M��фA���É�V���_��h���yd3o�v���ʆYﹿȜ����ɳo��"�.���AQ^aStO	 ����\62�(YJg?j�w���P�vٯύ���1����5��#w7)��?"�k$����C���@�����-�8���	��t$X�\�l�$Ҫ�А�s�S��".bQd��@�4Q/��	W�].��D�=��;�fHe�]jh,�1�I��gM�X�6L�a�`�|���EwpWu��N�yQm[O�����fh<��i�k��2�T�D]АB�����DZ]8�Tu�/�5���ƶ[�4t�1Ѵ$f����Q�e8�j̠)�������yO���@V���k҈�:(dy38!��H��.�k��C,s����_�q �`�'���}ٗ	�'C�.%l����⡩B[+8F'���YAom�臓	�w3��M�Q���TWN�:__���2/��f��ȉ�e�rD���[�'@
s�I/X��Mg�L~������{#�^m�B��]�5G���9|-�����V�S�=��L��c% s<m��^��f!��q��w��1[Vд-�fO���%�V�1ܩ�Hu9��e�'�Q��!��%S�]=-��3�<9�G�idZ	�>?��jћ!2��s�l�6�95¬�tEn�.x
�Z�
VtCl�f^��]a��W�;4, v�}�%�\����� �d�8�Ջ�V��D�ݖ�t�F�<+�4Y���n�mfK r=��Lf�\��mAFY��g��K]����a�I�c�J��P��h�7؛��g����)�#�ZC�b�����ސh9cw�uP4~d Xàb/[�6���/d!���^�:G��L'�\�*J�_���T"'g��P���!�����"s���S?ܤm9�8�����1� sn�� �PS��JӪ��t���$��}�
ryVَ(�M�:\g��v����y�vv�3��8�y�ʟ������K�֟���d����8�ĳQ#|(��]�}�IzW��ql�5�Jӑ���W�/��j�%����@�Q�n�"��AV�4)��O�J�l{|U�h'��[냴���Z�*�C}��R��(������.=Ă�ja�5����B���ߓo$M�����֧iEs�G���絉��S����j�$���b��$x������}�(�^��GZ�*�S�������ˇ �����N@��� ��	P��dA�4 �y&��/Lu8m�W"�ԛ���{eg����<?F�~���3�Un����i�O�b�e~q�Jd���8�6�[�Ù=��T�����7� �+�8h�4�c;�)g��5/�͓�#ι�a$:>&�q�P��w��B�s����� )c��;��� z���[T��A��u���qu����?������c�?$�C���A|���2����vS�G��C995E����c=��3dh�X��L��]O7(��U9k�^E[�i���̐�F ���=x2�V���W�l�f;XK&��`Ǥ�g��ѱ�obIv��fap��Z�p�ALuV`�<�����.@z/�x��"�_@�9���-}�
&�`n_r:X�u�9�ԇv��3ִݡ�'�U_�M�;z�_��f����?�K�{�ǜ߉`d8�cK��+"N�sY����A1���ݐ���R���mX~D�<!��ɼ�(�A�V���Q��e�3�:3��W0��Їȧe��V��y= �4�O�K}6��C���\s/�:�o��2�m�$���;�,\�8������!�L��IFrԭ�����p��,�Gu��LSiHA�v>³ ~���;���qf���'���X�s�xb�
�4Bn��y�p��T���p�L�ֆ��q̹���1���[�5XcÊ>'�� �Y�E�CxL`�%b�F�׸)4aǩA#�0^�[��: 9B���m��K��g0�?�I25L���Rj� v��2ñ@��JM��Rd���T�!]e�j�ܑ���+�C��ᬁ��G$�Mǘ�祖2q���aX<�rmuo��˩����a
��n���x�a���D
ָj�*�9U��F#)ێ�*��=O���½s��NV����RZa
��ԼY�q�m����m�"����-c؆�nW�]J��	�h�n��w�g+�Lz�>�L��i\�_��.OPaM2��i�y���r]��&�h�~�m����?Y����^z���Ww5:��K���!�2�� �p�R���R�[�XD\:����&ұ�]ȣ�K�Ƥ􁮻	]��{Q��f�s����m�����#���&���y�������ɶ�&�����5w���� ��:�
�	�Ɖ�jd��{�K�}ӀѪ���D������d�f.�=H�c(���^��!'&}2$�EO�%�sܟ��ϯhCQc�5;r y�m��� ܨr¤�>e
o����1:Pi���]`����z+C����b��y�)��&gR��u�|J�!��b%a�F�<�X\���F�gB��\&i�/rH�{��i���,�= �G?��r��G��alD�pOsЌ>J	�wu��:���$�GH0֣*W-���r����)/j�W�~�+`5�Zq����9ARS~�h�GI4�6�i`��B��}g� %ic:��B��ͩ�$�wT�ޠ=l��pbj�	��g��a:K� }��p��� �=,�h�"/���^1 ��0�`E��ы������q @��q��������?�������٤�-섲Udł�[ܯg'>�gU9@�@]`�����.),�qz2[n�P�k�?a��a�G�!*��{(+4ԬA]���Gd�J6v�`#�A�x�EcJ܌dr}��>6���<^#���T�3��[�*-FH~���'����
��PVp:{o`T�sTWN�^�q�{�ǅ��u�	���#�9�@\i�$H뀧�Q�X,��O��V�z���MZ~
+�O�6���e`�e�i�z1�	i�j��e]���>�js>������Ω8c�V��G<)�+'������)�vo.3��+:řj�*ZFܾ�\���G������_��R��7�y�ɩ�0)�_Oe�4���,��Y[��-s7Z�t<���E��FN��R7�>�]�{�F����8�%4t�z�k�HX�*�1e�_?���vܼ�	��00��R�Ղ��Mk6����C���>ɼC{���/�agl�)�(���qU�����ߌQ��:�f���׈��VS��4,�3����9G��%�����'�<��N��F��&XB"���[�ۘrW�(5�B;���$�`F�פ�b{��Yg��+$����������o;J�wC�B�Ԯ5RU����^��\�(�3lF��8�{'�Cj�1Z��)��:(mr�q��^� ��L�Yd�`�p�X@Ϊi����������� |���@���O9��}��9$���f^�j�B@=�G��o}~�9����r6������6U��*w��m�Ŷ��8���]�@�&� v�xj��朩�D|J����OB}m���_�WY����q{��Y>�~��C -�]~cٳ46cO�!d�w�'
/��.�
�NB����I�uۄbLm?���|7͒h�܂��xfeL�y�_���XX�z�.GXXͯ������'	`X:����Do��ʽ1�P��&Q�aDŃ'y���gI����U?lB2�я�A���^0�$�d2�l+#�B�kUpn3�O�T�?4sЊ�r��)�u�L�yXAN^��(�X����������a�:6q�q����o����:�?������2qn�2�əxI�Z/C�d��I`��9�m�V`?\��\G�˺����(RD8u�HhD
Z�z��v�*��wC>�)n�J���L&ʫ����5s{q �^n��q�C���xk�e��#�����s\�q7���
���ޤ���]I�bFoF���J����#ux����Ob@��çg���wL
;4f��b�����5�V�[�<u�/$�=�T�	��滚T?*�������N�j��2��>}�]�}��{��R�O�PY���HH�(ٟ���:k���l��:Sx `��j�z,.�S�^�6�a7�rR��>�È+�G~c)&cF3Q��,rr=z}�ʹ,����9�v��<Ya���]mSyS�뼃6���d�}1F<]�^�.s��k	�]�b
�������Y>!�kv�73��L��W�9C<��� �~�*2�_��p�W�Ɲ��X$�2^5��z+ ���狳���]X�/R��'~��䪒�n�/tB�~�H��!�a�M]�'�bܞ�'?�?�72�V��AH!3cS��I{�y�Xw��*vr#���EL�o�vX@[0ߠ���K���|���hk����YTR�Ɨ1�4q�B��֙�P5��a�\/�S\7�W��/�:��DRJ�ݻ_�r��o@=�y�|����ǌ�OQ��j��]4W`�Wȱ�DxI@CJw�MOG>��w_�)Q^��N�G��*��K����㨜V��:�Qχ��J2����ݟs�BT��d����D���� 1�����4n�����RD�����!r+����R���&����8m$d^_[��o�F�`>'O���:��1��}��I����c�<Eӣu��/j�~=��&U�k��IUX~Z�$M�k�H3;������$G�b"[s�^�\��V;���bx��m��p���yVV��6���ɮ���¾*��=2�{�0��9��m[z�@���H�� .[ԡ�guJ�5��p2���g�2���B�\8���'�Q�ŴY���e�A��v>�X���aJ
p������9�zf��F�q8ti��L��D�h ����G1-���wĩA�Y�P�X���
�Ga��q!aC��־�ڕS��0�C���<o�uZ%ݜ����_&a�[jm�]��
]C$͚/\��_B�Ϭx�k~�^ˠ`�U�V��tJ�]�M��ݶ%
;䱛KW|l�*�&�n�fh2��^rs�N�d?�0?R���ϻ&o�Jn�HbܪD���q��M��<�B�X�M|d�����j��'VZ#��Vy�+�\�MLK)r�xsw$�U��r��%�t���z�z-��L8�?�ԟ75j�B�;g��ּ*�+��O���C$#�
�w�:*�Hb3�_!�j��ۄy~�����nl�1/�?��!�f�T-���lޓXx��6�|�C|�XβxL|������T�W��7g�T3�5z�ìM��b/�$�`R�y1��i`�?�ё���'h�/ �M�G�S�#3�� 1��_���>8-��4��UfH���"X��ۛ���s����}T���ѡ��z��zRFF����i�zڗ�٨��6�*����_�8���1�R`}�	Rҍщ[�P��'g�2q��4&�h�V�N@15�J�s������)
�k��;\�+�����P@Ll���7�H����?*��"8^V#̋�\~�~?7�����è��>�#˴C���)���P��Ď��"�5��,ꐌ@�:w��p�ɠ��>�`Y���8U
d�'�AY}�}C� Oa�%ԅR� ��d �_���kf32�f�Hľ\��O׭���d�e}G��y̏�t���"�zv�����S��^zb�BM�P�@ޫs�,���g^l?s~�\��/�]9�����a�+o@.|f^�"��L⨗T�%�C����Fd����� �ˈ���_��T��?�9�>`��Jj����y`2��tr���9"�I��T�P*C��D��/ y��@��1�-0I�,g̃�)�{i�%���ӿ�r�R������j-���WwPH9v[��P�����B9�>��\K_��2�ER��;�z��f�k� ����--S���_�Z�ڼ�����t��q�A�.d僙cM^�N�X`�f9�M�D.�:y�xbܯ����%�	!�Җ������X.�hr�*p��`��0)���ʲ+�v{��%�I�������Ƣ�&T��[�(�t�����|a�.k
E��A�P�nP�Z@�glf�j�2�� �
p�7�H��Yh��/�������)}Z�o�1#8.�-���hd�(>E)���yd>����8��E:+�S������|��&N e�rJ`����%V�m��!��)�K��Cc�w�:!�u�ub��h
y�Xȟ�&���`�����X{�?b�8be�^A��Q�]��J"�Vp�1����^���[wUY�mѦ�Y)Q�61�|�?�>��0^��4�A�|��\�c�n*��d�i��D×�e��j4^eꗹ����7t�p�ŏ���>�,��"��^8BZ�bJn��X��P`p�w�e�EN���Z�FruG%];EV��<��,�[� �K򵙫V��p�|}p�Ƽ�2DD&*Ĉ�)���|���������;ա9�,ZW����V
��Ɇ��;E3�J�[ֹIˉX`$4HؼH|��x�2,L>�-^���&�`ݝs�R_J?�ӹ��)QYt_N����w0a���Ɲ��u���wz?2ʜ_zrq��1���E�INT�#�9R���3�1f�q/�{-��
��(�`uF��/�K�a�1����b�Hg��Z�0<��kg,�=)y���Ŏ�7}ӑV&Ɣ�p��Ub�DQ<�' 2�wp^�{_���Irۥ&]o��78��R0�E�2&5��&	e�Y�oY��V���*$xm�μA���C-���T�C��<���`0"c��E8��{�j�rw�v|]�k����c,y'{K���i�4�@�����t�ISY���i)a+�/ی���l�v�3��0��m���0N	�ܣ�#e�Pru�7v_����ީ����J�l�cHE�l���b-�\�������z���g��}F���/�uj��"5V'�r���-.L������y@@������2�Ϥ9MQ���J�MB �HP/�8->Lfq���2��D�7p�ՠ$a���p�9	�hn��X*+@�)ʎ0�~�+.�4@���o^cŖ�y���r�2�	&��	\X��P��h�l�lw�(w|�&��3�6��%��ѝ���l�$t7�_�)p GL���ֶ�%�3���<#cjZ�d6��6�r_g\K�C�ʮ��\�^\K�^"ߑ�OJ����?txe���D~��<���K��#5kn�5C���`7/S<��P{%j+`�3�31o5���̀��|V�G#AQhr��3���N���ޢ~�^��"9V��v�VX 8�֩@��	g�*�~eLߔ]k�R�&o��#�2pJ=R1�z������fn����W���K&��0�H���k���}�f�	4��.K�[G��'ۍ�N���I�;�	M�?ca�;C�yqnB��F&�ݐ�c�t=��Tqͪk�~ǭ��� �>�S�b����0��ʴF�?�l��Qy��>׵ܳ)NZɇ}��ʩ�<G��4�O����v�F?�9��b�D֩�uF�O.ژHP��2���F���`�A���ȥ�U���5������H�YJ��t�7e3�����$ވL.|y� �:���ts�y�� ����PBm+w�P�@���Ef�W��9��,�U�I��q ��0��^r�Sp�B�S�qҎ� �$�?£�Yf�>!p�~�z(��1lj��Ș�W���H�s��+{�47��a�y��208w��YqE�i?߉1t��z8-���2�y�"e�*�F�H�������V��I+)������+3����>w�ApZ��~�Ydd��F�Y#@?R%�� N����p�����f�'gZu�w��v	�ejx��6	z��@K�<>�y�C\����SSP���Gݣ�{��s�����5ӵ!��jR-^�P���.k�7np}�y�Ts�r˒�7� �=����[S��� Q��,�*�6��4tc\��f?EID�uRu���&�d"�zhJ83^S�_�.Mt��r��>D���`w IU�{5>HPD�����{�?�n�Ho����e�����8�Q��s��X� v�d���p�5>P�rZp�$g��3�C�	��DЊ���kW/l��k�#�GHk��O��f�}���TuE���(w��άpP�GN���];��f��hM ��1�+���>\��T���gB@�\G/IOs�	��M�7N����8�nu����w:��{s3���l���[��W����;����� !���hR�X5�qY��C���oh�BZ-�9no��j�&�#Эwf�}��=�g:a�"��#���ݧ���nRX��j�����U��W���l�H�}�a��ֶ��'�8�ORQ�hn����&M����=��,��х'�����е�֔-#���)(%�qŵ�`���AYi��V?F\�U��a%L�M��`�ZUE9�~�Wh�a��1:q���%��C,���"g`�H��8�P���Y�1^������6�A�ʌ�k{�CR	�g5���pA�аH[!���%�&|�5�r!�'%O��ň.EZ�|�)��w��m)a*L�k�Q��/���X^Nh^k���d�؋��a<|-/�	��LƉ��e�q4�����|]�qM;
P�>�,��:]� (rD�m6"�BH��"��˺V�D�X�4�z������Zˢ4 ��|�v������/�0��lg��2q��IS0"�a�vfg���/6��C_��L;
��S&XIkt�͇B���9y��l��v��Nl}W���*N����Hp����jt���}����եʬKRO���L�֔D��B3N�n)G�XΙ3X��}����ܪ��r*e��<Ư_Hey�Bs
��;/�!�Н���|��|�W�������`��.�B�����@ե��$o�;|S\i��?$v�)&
c���oy����Ȁ�bF�P�%@��jP���ͥ� ޔ��CD��y����>���8��Ԥ��;=����0E��,��6ƕm>���?��E6��-��W*~��,�Bi�����R*qW�����!۰;(L-}��Bx�U8Kl����B�w�Y�L�r�9$�t�~��Ԭ5�Zt���;�p���ݓ��\^N�&&��������4bPN|����G�aE2���G+tm�=j�R�G_�[b^���(r�`]
F�kf-�9�h���i�jmv��"�T��Tt.������Pj�ЬnK*�*}EZ�)K	?e�y���^&����%�����?��H��T�;��^�᠓�o�����T8���͞h��-�y��蛰T�*��$��P��]�̊�3�
n�'4m{�
��f?�}h�^$R?�l���x֊��]���!�0�6OCx�ݸ�u9W�c�)VU�X��*�jB����OLo�)?�n'�x0��K�^�W=����ٹ6�Y�����¦e�(��(͝T�D��Ց0�1�S��6����_[י���=�+|f���i�6P�s!9K�ۡH���G�\/�f�db�INC���_̻I�sx�34�04a�ѣ���r5s�ķr�"��8�
H���E�3b�t7^�L?S����H���kz$i���ٔ�K�IX1}�u<Иg�� �x'm���vlmmc��%����"�<�2��b�
�E`,����𷋠���G�/�:����-��`��)5bG���d�3��-����wBs�y��B�ð�UO�ʵ_*�\ӏ`)���|�ȏ*FE�F%���[.{�⨜��F��w�M�[A�qYBNJ��@���߀��h����>;b4z���u�p��������	3��Y��JNS-�Gm���f*&jI���z�8T������+�L�X$щ��[�R��_�ؔ,�'�ħ�s�I$�8�ԦZew��w�2�'�"/�%`����`�s�嶔U}���W|�޻����K�e�p�F�0~za�'|�C�t��
TE�>�
�CP�����"��q��J=|LD��`�}*���u����E��G�A����?ը^�	��5�[@l�7�05�u�뢸���^�p��yܺ�T��,J��-g
��݌�j�T_����ֺ�qc,fu��V������W���S�>����f�������{#w�۵Upyb4��#@g2����D٩�lU�����_���dD�<ݐP�N�����c�&Z 7\)���Rm��j���_R�J����� *��\�ÓZ�Z���L`9����x����bP2�$fZw��5�nO曤c�~�3aZx��Eq��'�/�(~J��Or�W��d0�ǑB��Z�K�>�pٗ��k;4܈��U��bÅ�$�MZ� 
 ��3�s�͋�F�yVa	�\�kԣ��hIh�z�U�~�>	!����Rh�"'�}��e��5���8\�80�H+XK�b-Q�bJ	��j��t`𻓨��GM��PoT�4�_t'鰋n�{ob3�0n�ڭ�t���cS\�ʡ������
�!� R	^B�$ϩ�)��ƈ>Ê�^d��膚=M#d�N��䲢#2�N��e�Σ�V��U~ŉ�T��i.���иN�cf�=�YQBTL���������*DT� �K 
��%L�[a�Q#b�t�OG�#}ËQI�ʳ��o�[�Jba���Qd���Ԣ������ �3ж�=�c�O�@�mum�J�im_�aٗ��X��w�y�gϠ��(�;&�|�w�u�Ӭ_�U,o������e9L�}���WC:7"0.�Zo�<�k�����\����wOW�0�-�oyQQU������cQ�<gn��3K��b����=��p7d��Rm~����(>���3��Nd >G��>lF�<=�~L��05����K��6�r���/����1�'|4htU�@��pBf_Y~�ϗP�ڴ�Tʽ�^ү�>#�0W��,ݸv�t�0ˊ"s���U��f9�ZD)�1�/g���!����pD"�P�ϏT�32z��%�L�òr��Y�r	�un�c�%��(ah p�kr��z�㈚s�d1,-����ԫ�b:c�y����tg��ct�$l��,/�d�g�w`E<�����6�P����x���� 5��J�:fZ���J0O?�Ɓ����� �Xn�N����5�g}�k0�@��$a*�P��l�,�Z��*��wa����Հg_x
�\k��"�'_���psh�j�h0��M���]���5a��7h'�t�(��D����|,L�ȡU��ם��GFP���b��ą�c�+Z�'�)��
l�J0��s��P�;��C��{�[ܚ	q�?����֘�&�k<��K�>t\��L���{�[�q��`0���d��s�ұv�*��%M=YH0�V��D��:G��-��tn%�V)��R�9C\O[:l,�9� ��0'O�q�
��v2RX��ֲdT�m�W�
�w�>,�a�>�`� $�j�U�\%�VV��8�AZ#c% U�R�J�*֏(k�-��H�� j�?�̲D<�����5d�³�j�f^�F \Yέz������U.a^%���cw����eB�<��,�����38�M�/4S�=km�5��w�1%�����*	�6Sܷމ��5+Ǚ,9w�V���و�Ň_?��m����]Ĵ'�e�I{����N��?�F�Fv ;i)��s�k�]B��J+S��4�6 M@P� ��=I~G��KPn7�XEY����/9C�p�[�'�$O��t��f��/q�;K
��5%�fn��b�Op*O^`'Z,�b�%<b<Rq���\��0T�Ô��4�I<�� ��(;�[�lq$x�z�	�:�Z��.L��"�@1�<yP)P��'D��\��o�Vڧ��"��ܬdQg`ڙx��V��<�9��e��#�J?|��H�V��\�Ǯ����XA�S�k$��H���*C���z�{����ŭ5�j�k���e=��J���5��Ì ;���@_�u�im�#V舎=��e��X��7��)u�������Y��,�Zu0�׷I�b�"�?�d�F����_��\`�ػ�i�J �䴏 ����t��(��g���E`�9G'����gaC�Tz�@ �׫�O#@�vRz� k�+���,ǧ�$J�����L�xsm��e�?-˯�R҇��*�#��`����;����09��wk�G�eT:"W�� l�w������OU�$�9��K�m,�V�0ք�4��ġ���V����
�dGk[��V/f�e��S �*XFA]za3���:��K��DI��r1~"��t�+����&a�(�P��|�ڱ��kVo���^�f��1p����sY�q(A��ʸ�J�N��ʞg��6�2�6��u>WQ���Yשft�q5v�N��x�h߇��#WT�g
�>������.�r�~Ѷ�6��?Aoݳ�!��\}[�3���؟ e�:��PW��A5�.��tP܏7>H�0��=9)x@�� ��@)��Qҵ���B���8`i�be�d�W�����-�� `��~�77�mG�϶Q���.O�󳴄�!��B`�j�٧fWӡ�x9���w��B*F�޵��iR{�T� �Z�7r���F�����i�1T�-������eY\�w��m��,6��ݽ��n����خ�\�lD�����mdV�qhɊ��z�xm�>�R(t=A�L��:+i�@&"�_~Ϥ?(�>�v$h���?���;����}X�~޹>��VP�i#T�=�#~�����{k���D#��bZ^bvx_J��(��
��p�bX�|�G��zB