// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:22 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jc6vv6X7dvD+9qNh33180LAumfNHuXeekfgGoyfenoU4cgFGEXYUTRYzIwgd6oIG
PVVUnEsKqDRji3866fhhWrkg4fitPpZwEQS903XXcNe6eQxsay2MhKUIxm+ah49w
wFyPYvk5uzZN0Y1U0LR+ZD9TwZSR6eYje9Inmm2AcHU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32160)
hLsd7+hVr7lQP7KH4eHWy5nMudesuqzlFGGCPV7BotFMJ0HOW6yIl8hXlGf57Mwf
zfv6+RWOrZcJ9inuEUWWno4NBRyb/Ys6plDc2BF0jiV2JYCd2aoAI0DR2Tdv7xlH
NPDTsMeBZVfyUVrWVoI+7A7lLfcevShGfFxYSLDydXMHkcKq4xw/MYjMuJnKKMok
jbqbWDAUafuvaktOBh5YvZnYLMshi66kYWPTLLTNn/cOZMqKhTUlYAiodKcuzskF
soUCidhNKT/B/rY+2V5+JvXDdVxavn9PPppJ/mU3301E7tplkT6fyhCpqoawpPVy
W2dJnrrFv9eVWOidVaguHj4+xdc4Zax4Rdr5LBU1PHFu8wtXW5tAUrP0DGDuwHO5
pYPech3yFRSe/FC9iulhikzMOKHGZi6WqhRGIjMqWDvRDxXmt1lJGH32P85Pw1s/
FQy0qijbK4F+QLttU0+/EMs+ydYuYaRXQ5RRj1RDBXP/Z8CmliY+Gm8l2ulatx6t
lyjEWcyrc7zkFZgzHo5HRDI+RyQQZn7iUbzdaID3gi1GbODeO/noEMujNk1F8JDr
DtrekSw3dKwlj99ahSTcWlWoTUUq03eq5vFf16fDpNFfYcrfYyOWYwz8Lv1Vj8n5
nzt6jkWrk0X9H/xs0Q/Ce0cDxhnw/9rFvYsCRxcJkCSJ2sA/sl3zL6i8IKX8anuW
IL0eyGD6Jedwn/ai2RzBddETIwIZIbdhkZgq0N+vJFhspKmbJgP//vkZnFISbvQi
bKUmGHyI+oY2JoGPpmnRUHswgyBsggpegYFDXTL1nKlyiGsy81nQl9niZDH6uFry
lz6A5IPpM2ZhnkAg/WoJHVVUDYaW9MCU6wdVFeZB9bhgqenIx5667At/B+jr1khe
9ysrV/ukmWTXlmAhYH/mntBrz7Q25oPx3vHl1yK1CSgu+yIa+fArRO+aWpk7VElj
nF1YvMX+1vnWXZcot6mzL+FrGMR823OxuuEQ0tYuiLObLqwUlrojQF+ZUXapNRlc
bn5Z0wdRESl+xPg/6uRZ0Ki8Yd64rzejZVWoX0FOZX/OG/RBFJP9crDUdi9flFJc
VSzcVhpwjroLlsLJcSogfTF/g/6D4Af49x0nqxiKhvRVZiRKtPGT4wyCnWt3qspZ
HEiEU1qJoKBYQOhKuJY9KcK0fuFwKeZdznaZpsbSxE3c+iffI8JghcqF83jeFf/z
QiwY+wNjKmp8dRS75t8+wz2qhgvhtjfMxdcwcOCSXEOWBg1mFU4HtlNFSiUl7ZS2
c//8TLRYDu/xv7EFUAgAnOIkuBd/2iRrRUf6YoEs+18nRPfnLS99fXVqjYqXaChE
Blhe9DJXdHj290n2LK0kx2NAfvrlWI1vw3df1RGYnv66EtZtC2BL+n7mrnQGRkQ8
uKWSskzgBBk/kni6cYogc2K4VD+Vp8qmb/l62xEkWMksURN9xNkW+WtoVr2zC+rB
pV8bNhylqTO0xEa9WqQyz5SWAQXr6SjD31IU+7j7PXUpqof+Ju+Cmq1B9tvmKEgB
wpKtW574ZfP9wr97BgpvWjE8ziGXO+fHSMm71aZlLiVa7ezh55sEyblBGWSTVfoK
wAnKHdTinkniontTG9jpbLM0kacTrmyEiv97kOHx0BvGAHRf7QKXjCwDy2xHSm/4
x/20g43DZi+5dQHBjAUjsBQcUhgvy7XalVuFUNK/OUQtXch4+k1XNhnZp6yELejH
8sJ611XhppfYPrv1n99sJE5Asj+SN9nqDbD02xrx1phxSGJQ5mXTzo0MIYZ9PfQp
LP+wh0/Poiq+Z6fj12Smmd+CIjrAQn08ObDEYeDJCqU5vh0gzhW+f596gvD/IBeT
k6dbB6YNFwxF1egOhss619/PXEsdE6ssaOB3NluVNheGFHo4jLcoeIGfn2iG2ZlR
cj9a9UDuVRpFqHUf1XFZpwgWeEFgXfQjlq0Y+gYQ1lOpMVSaP+/0s+aCsEzOQQ09
GmbAMCgVi9fbpaI/drScp9jm2SMuyHi656oNZ14wqtitiyr++/DzhU9G+9d2wTnj
kE7ayCoAiivwpNz0W6820dr03STfsXZe83JV28W4K3eIV+lLn4T0Gm2cfh7m0Vke
UOtheDUwpohI8mtaoZmp6jTFCR6f0mXzCy6vOkebrAE61sHvYmRt0TiDTMob5C/R
E20nDyk/xjpymjYmpXUcyX6Z6GpXEpci6JDPx6DucnYHP85PUGcOBCg9z9/TxEVE
uiD8fQ3PZwI0LWdV9mIn0iEzP+wuEmmnYcGJdfUlxJIZlwUaU8+iwTEg4pmhAwf4
KD29E81sEl7X/jWVQOEYZ9lvV1/ycu6B+qbgvOs4Bsvdc2ePtFUPBy5qW9M6xybD
Z30QhPYg7hoWPjC++btuZNfi3X6C6Trc2OtPiLCx5rTFjQ/q/fUehNPM4B3PqLxz
x7gYioSJS+8O1fmAdeTuYnlqDPQ4ngWxDJAJSmy2itM1Jlo2v1sL/WwmgKeCt+sc
S/h/mIpxbqZYVT4DrDaaO5DgcJzdWawQp9RCJgCCv9XVjHMrB+1qyXlQoXl89eRn
czJGHfFzSACNtFmCqv+IiiUpMQg/34R13Bi/WnWcCHoMTaUR/vHT5NC+zN9b5FgR
00p3k7PDBm7+1A6fGKqi3C8rURpe0B4KImKTgRC1iqTPc9HPJPbWFuU02w0RBQqv
jxPsV9xV9OZUHgboFzdEiJQjT4uIdoR7AcbL8vVzpOYk5+0M5FD9Qxdu38PAABW+
zu58H7TPXaGUzvr4eZKszelcLBi9sl3vvJCBG+EPNRtP8Lz1GUtqHuzxbKMbke/M
S3LdhYyu0WIU3wMtpluLU2OzF0SzUeqcrbiW6+CHJrueyjPVTpcCcqffWXtkFu0d
nz9OB4POcbsLqIlY4+GAlpbah6Bthi5MUjqHs2eFT2djUhgAF2Vg/dtwhEJwU0BC
NKDvQBNv1p96HqIUg5sIu7tZabE026ISM/GrYvLnltK2C8fd5npmQBabnmTKoPCJ
jDq6wUeygKnSSLqQ2ooLe9Q8fVqZYyeYes7Q5CecD82aiJHACuXRpVGshISv7E83
W81OUMlFybw8PsdlAlVw7Sx35gVUamScj1qWJ2dl4Yo6f4V4YL40qjxSBylr3Hxy
vRST9YOI2dHXfU/mSH8MVBtM0Ku5/R/HHwlLMGBjtwlYc6UL7OgV4x6RRJkrtkeL
4YeMF7Gv5+8AZn/HIACxol7rNq79TYi7oalgV37/xtYKpFQ7EO1VkEcUtKDbyGBz
hOWTspZ+g9APh/decFc7apX2UFiWIPSgRHETrZJjOo4svgECmaNWadULgac+G5Bv
+FiaNlnig0G/0XiBb7SUHH9I6WGz178PN1ClHhrBU/dynG4dOwaJt/kwzF3NHoSq
AHDbMivY/3xXJBXqwYER/8HjZgYr+gYacEEaOtBT4erk2MWJuAcBeMPQaLD54fl/
yJCunsr+9yF1bQw1qlbg1SOFGHAL4iWUSRb6GAaW6hgOlYpQTxM0W3zL+XEIpTW1
ZqQQ3/hN8wVXWmTSfdgeb84inWvmYFBk9S8vB05fGmWti8s4kxe80v+tzlOPebx9
9XXNNBZn6IGmhUOkxOXCMpxiBGCO16CIP8Wy+I4XB377RrQ2Jwg1TyudHbppKhM0
A696pj6B66A9rfJjCZihcCfxj7DgdfB4wgGR/LlR6/inoPwFvCgimIlJ7Kequ31V
1bZ22BL5W28G1Tvh4iUZ/hIxrVbiYYeCU9SRKQ0ckgK5yv8Oe1v9KGOzI5Lln1OD
2UNv9J8HhLAM03a131izuowgd3sPT5FmjJtOg3fU6Rft3M9pfBjtEstcNEMVdJUZ
MAXzZeFC5BkoUUz/Pi7q9Lznw99GYBDqAZwS5pJOnBUwqN4cuLNZtXCKbvfU0NUA
Zx9dv+Ygd3vUiW4alP6MeKFEce7Hgz93Ti0o9DixoWhiTCCFkAUhDEMZ41H0aZaR
1UVr9ra7FhtljIsgP4dALVRBIoJpVqK0BJ1RKv34EK84IlXWrde1K5tnjH0aWt4V
DanYgC6802dW6tkBa4s5ZPMKBy2GxfWAUd8Hn1t3iixy6sFmHWvxEsX7sBASNFjF
tMB+n6YzPprlvi6xbhMLUFvzSWcr0tUnMZXo8eXMTe63beh4ZDgf6vLl6h9Wy+Vx
o9ouZDELH3+qWSDxoprIVft6I3xi1YEw8VEAE6l2XPvVqRcWt4Ov6D4SzUXf+4qr
vuUUbhdsSPk7vGav5SVVT9bRj+90ceSSEYRHIZ7lPyGgn2c40aQYSe1vZCPxK1jD
CvcRxJk5I4JMsrFJDnWe0+aT064rutBRJvePArY7zFVqVqZ2wBFFbLdFaQh7MW8H
NFIsRLQMvXqE5vwbHNx1qhTw/h3euDyaZXE6FND6POveLz7UKETsWUGiltw974s2
ZSrUs/0dghjd2m+b3Skqux17ZsAIb3Nh7SURreYWwOHnQ+sVIkC3HMoxGgNJJOwP
kBAghTk2cY8xXiUCcJldiuVFkoNfcv/0PcQO0/iBf1naqlwpF3icF4xQpoO3XpAm
5AUyASRlpjEkxm2sEFw/yamAi6h/Ct1SfdPVaiBRjrIt03JRPzPO/YuaRCX3o4TD
836zLqhuSnqu/qthKTUARiWBK9BhoHXvNc+TZ5WhZ9WtRk6nyLJ4nn31+Cv7O2fl
JfhAA68ihbGozQdG7m08otH5I+zWr14yGTmuAfiHItBq7mu+O+oK4p725zT+aeHK
G6djHDP5NO3ElY92eVl1PXv0JwluatqHyBEpeGGtpGynk0JX3qOscZHRmPtTlLCx
nhBg4oNKRDxJH6cEqAiITpr5W63Hjms2pLE+RMUKe/TSPrsQ6EB6WpYKOVsZ7U8m
Gp4niMZqweGKJUgxBTvI8ZE9ROhiJSHcuWeZgObd1hQoAhNPpn7QgdW0FWBcEMnz
85pt4SqA22xIhBDoFB6XUXGt/Pan4hgXJCdOMfoph3/Gttv96y9YghQeLsHfRMim
9vkvTLolO0cvPron5CRPknNjIQ99gbdnWHVg1xLsfhCCTemL45rJ8/4DiKSdSg7n
dKLPHfk8NklKbAQhYG2PwWkGpJ8OgTMDpuNx94pWaFORkplu1Tg0g9K5NzkA/Pya
xUj+FuJE+avjZM5dI1qvsU65ltqJDn2zlaBNMF/x9WnvUXdaxkP8MmxvOFcueyPX
DU77oD0xVZMU1Zluqsi6Mj/I3tLQ/vy28y8cce4WY3e5ufrKrn9urZmRNyD0X1m0
IRf6E1oVwbUoJ1CKLReShQye9W47miH3r2Kr0zYTwcc3JP3oaQ1SJopUuajuTjs+
lj1vGk8HctTAoZmmqM2I4wj7CThqh2LuWoVY+IlNZPJ95Ux+6sXvJ0fIQTMQj/bn
/y809Gc3L6kUcFVY0e6VleLy3hJSD5furluelsVgZzGfJR6dzToLJv0DxrVewxox
S3QIqt3KY9BcJqR3Z4D197u/9VFNMO5Ss7/j/+BUbOKjbF4fR++WrMPIudW9Bmih
eU4Xa7TimQJcc1AAd9DQC7yLU4iR+hAWdzgM2ms/QjMvPMhg6nu8iwE2JTTaF4zj
otr1rjE+fDbqDzL5TsXoap64KxKHPa3a0SITb1ljwo7WyUJ9kCbspvls24seZwIV
1eePCx4o85QQBTsb5xzb96UVkfZyVRkSdauKqnhqMapS1dGaN4TI2G1AW7vLgfNe
5OxzvKTZVOtilVZdgb8t8B2d51WOAvVnxdiGt27Uxgn4wd0cvIQp/v4vi59Q+YF4
+Nxtx2VvUPoOrG3624F+HxVp+KlXFXL7ZVoiwfCaGTJl/VTF/XcLJ733EIjQyHUn
hFbT5h3DJp5ypOqF724d5O1rKEaYLuezx6ybzRjFvB0cPwBDUErIMafclCe4SNjK
V0ikw5gRKKs6aGN86WOp982wWbHjMIjsGhmig0irVtrJL8BwlARlTrEUi2n6VfMS
6Zb79YrdkzC/XqXMTZT0p57n1csxaXeXAey4V+cJLIxivpsM62MIcV+TzW0o+F/G
1HijcJA5qiGDgRgA/tojMd18rZmjVM63+fu+TffBgZZzIGI3HSJEf/zPCePmge6K
Ir7X0//RmnVcVW5Bw5ZLPWrkHKsvxWvV1xTyYMu8CTtVMt3q271im4x/hgLy1POw
YGR6k0naCVHjoyElEbqBS1KTWqv5q7Zdit8uvSB5/EZcXPxBR7w1FyA3C3LswL8F
ebEtKC+42UOXN8XHw37hv6dPzIK9mpq6RxTi/ptRMoB72jtHa177rCIPamfoqJJg
K5MKcyOjJ0E/BUTBWMXME1yuP/YZCX1aLM/OdkoQCNofe7TwWrWXugXQQQxV9vM1
RecyFJqyQLSLUP8t8FXvVjYrLD2njRCaBAmroPk80ND2LqkBP55nds+7tBuvF5F8
q8SpBtQJMvLiWL4v1wf5gfmOyIgcQB1WM5Sir5VHtvceXgigXNwKKfFN9b99cfY3
ycUQpXuWSz4xPlgcXYpS1Y6c+NgpeZmY7D0m9LaE48YtdkiUGyPQLFS2FsEAVWmu
Dk6aP/D2BVIsNFos39jx4dfyZ/JqRjQoPMVB1VGDXQ2c+We+Gz7rTpV4z+BU465W
oKIfV9gNImWy2HNY6w4j19/R9wARI/9V+oXSN5N4BC9lZYHFYG65pZKdOZrZIV0U
tE+xbswTk8GFrY/Rm+8vaGdk+pzTajIMpa4z/BdA+vRcnxpMeg1ULSLIezxwwmOn
VtUt6klZF3y3kHN8XtvK9IQv1ajoofSJ8cKeFCoEK1j1rN2v3+jyCQOGW6gHDEfq
HJTUvGVY3QznZCA5b20/JNCU0x8v1fpuqrFYizlQR57qda5BKsQ3gu9x+cBFuOip
TK4Eg1NQqwHE4iZxs0g+IZWNkKvgGyjY2jIPbsbXnampKgoABAsa7tZLSkvop7HN
ozbDLU3XDcGPsAp840jYVoJql240w88ETmOXrVFkHcG2pNZAh0pDnheIu/RSeXNI
J+hG7UMMIoxHNHk0Mpctw6MFxD00PaPPPYRQ9Oiv879TfcG1tgnkX0wEvwAiEODx
NomFnmtHrt3Ghq4WgRtVT2JgBYUnaFrsNjTYAoqyOk+Tg4MDmO/SxqorG8+8SJqV
vTKnPWdIiV3b7toH+Nuuda6PSsKqvgkSk4TgVqfSh/eDh2O7vYgU+npuIqyIOcXR
C1TOofQKkJUq7mPK/21MWa3iKZWu+U/IgPbsd9YsDyl2sj6U8vdjk8WrrNRT0iX3
+S55s/ioyeI/L50WXpGJgMMT9jf7jOxMfqdBhJ2L7Oapu5KzUu0zKm9nIbnajfzU
f6DWOoBh/cCP5VAeXya06HKEw0NtFZ1yk8wGhjo2oUyTu2oDcd0hdHLA5dQQjkbx
S8/sKiLM5nFK3lTyqyYPdwz9J0M+wR24bpuEzoc+m+WQhd7an9E/L5AeVuvzOnOo
0cDLxlW6wXKkwKcQnHILOQXaKHqPH6lhXd0uVwA9+AKleAykwPVNOUJPdiEFlmb0
FHqihuOeh/NaToc6Q9Sq4bxLibqDwOLU8cEtqxQJRg67+sEQSlCuE9Emte2dBDOm
4/8nrgGyNcxYdMQf3VEmMCD6pumO2WHVunwkgMbR+omDnQPeakCOOuLQP7c1Ep97
oA2ZE68vykGLhH+hBs2KV2FjIAPhQl6wpVMDesQyqbigZc1dvAWTwnhf8Lk6D+gv
QTsgM4RPzaaXXZfftgZBMtxrDLLgH7dkrono/mdLXujdRuiDRBIj8boC98OHqR0B
86E+X8lcRrrn5/M3pR3Ki4441xu6sflFbRniSYjdirlKO7hGQUseQlaWSzgxua5I
2tCJk9+aqIHaD2jQKnkv2p1FxmQUzclnMmVmQbUdeiKtrX1T4eDxbvN7v+XxaG/K
ssOZkqaOQ4hDSYtzXEEmEtM/TgKx8wzM5V4+KE5IcGNSQppJ4621axLW7CZhsH3B
qoHnmXDuA0xTZNeS2S/i3mWosIFS8tywrb6tdk9Br4wGi5NazYMjnHlNukhdl8CC
GuRLAxORW/HcAy9vI1tnIyt6+t4U/ocw+pB8ZKjxVmCeaKf67sW2d/bqxdcsPsYQ
oEnO53PEwfv8KWWSgYimGwC3UFy82Cn2OWNndflx1efdMhPNrV1Dl533bitXmK+9
86QgUIqKPHTo1msiiDRQebd/QhNwmw4pV2NVaVYSzsMaOoBJayVcU1p0XtWfpZLi
D8SUIUxv9hRG7r4WUI5p1RwTLCUwwLJoRezBPDDptBDWiNfltgfS7oRvJ5rB7FeJ
P/QjOsRDF18x8DvaKP1AHQK+iwfcWHVFHV9s6J+smsl1bowuwXHoYLZ+pyzGRDh4
pDjoVtqvU7JcksF01U0op7cv8cqWD6wb3rNo4tO57+2zH3XjXP3Tw3MXbz6wlEQS
tfMftM3KXA1fHGh5wIN6O5HjI4RTFeYvlHYKTsrMzjHA59IKcJAgdXQ1DkqwCMMM
V0sl0ZSVWjKW5R22oT1IVrw2lpy2XT7ppC4QS0vSmaZ3FCXCDNuVstdOI9cWBR9G
GXhip6qssHNxUFJ3tqdUfGcqUpJD9A4oM6mEnnnKv9P3Jxo5L9FChcslyVF2DFyA
ayLEWiza3of2YxrI1EQzxa8tWeC2mQKqtwxDNrMei/1qEFr+nvl1Y0ESksWX/vKM
RWKanO/Op8abJnIh5vk9IQbE7UsuF3PSe1TKxSn++nnn+3b/iiio/Aa+XNnfrdX3
XJmFdPq6loa+V8Kg4uclgRD0LVZPRwN+yMgRDxH3s40edwHijaXFJSUa+JHYzh0r
IBGzeQW67d3pGQFxrbqFT/cAzWHLcncV/zdT6lGVVFQcqeU9UiIHs1cZ4eQQqs5f
ynBcXmYYUCJ7EboWyauoXKgVO7oy/q7/nnceYZ6UJournKMbOycRbgtWUg3aRt+X
pOqgtsE3H5wmbwGyetEMfDYfohYw3g5AFSrgD5JLQskUX73gzfBH5WtWqLtvm+jg
V5XLRbFfuoDH03h4EeGN8Ggxrpg1JvroxpcQ1YxZJjv9xsehRtMpw9pOTttRQBoZ
tb0VDGO4ecCB/WHspEJj306GjkiQXwJ9wZROddYQUMuFlrgYLcQTeWiUr+zKHif4
2SVi60O3I1s1XO5qUd5zud/j4QWClCgQzBlahLhY04nCspdVpoU7pwIACnxdvDpQ
W2ifofrOSKP8hHRSdXxhIbHtMom2XlzvJoVAKDRTuMKK5cnqu1oLZzuIJgQO62St
Qus/JKIcbqMPITThZsPCwn4uhvdG4Q3QWiZ8kdbeP+e+2AI3RRDqeCR8utYWHL1Q
s2+yn91GhBOnpKTYTotwGwiPtU1AGJ7JHOmVvhPl5XhWmaBdzseSZ2TQ8csA+UzU
+JSCSLfW1ztNxd4+A4+fk8WTUknfo59UisesOXGjH+rbXsSLyinKxe2Kci7SzFzD
8xc7hj+Xe3YyQXPYPIuJ6ZlAj+GVEiZeyZGWMHhE3NBoj9zxH52w78tiEc170+v1
A6hAunxfRieMyIPigqSRfzpl0o/wJmE/CNqfaRpSsOky3YrKMtoN9VOo7kEOCh4I
3u2dHUoKUQWx42Oz898CUWIl+ffttw0JnNPkO2JBC6KtSUrjycWHGKY1xRBn0CSf
JM6y3NWd6IypNTpwMThabBAgzCwz6Tutt8Cwj6RfklBGZ2/zgRMAbd6/UbkzwUCt
utyKvN1Je2Lns3mBQ2XvynXtbc5FLJoacYUzDSw+BgdgKqFCS3UmbysOFcShpvwU
DeoDRkbeiqOeVMBGryNN6RLASf75C9ivWR0jL77khGGrCXS3GeI5+3umRnHfswGF
txK2SV427lckQ6QSHvRhPbnFmbsqRLpqQHm7cX4Tp92cxzFLHfkchsqk0U32vXkq
ctI646QONAXYYhTfN6Hev0Mi9gWxFCAi01lU7dPrkIAulu3Yf4XuyS5DSdsszYNK
GpL85aOLE6EWKPJ2zSM1EMe5zzlyQ/vDZJ8O63l0bWze/DNGsRH88u3mof52uE73
V6+nr1+kMV58NAPXnXes6hkg+BMfMX4gEYOIhoGMar3cSw/WGfYiQZ5ZgLOHTCAw
fCUE/Su6aP5zbQtZhivpd37NqdNohlrIFJBC0EBjrM3jRdwkoAE3tu247jwcJugQ
BY/sS7VALAAgkk5s7ZTuf7oc3Us8XD9Xqzv8aPxcM/cgqGq1xjePjMNwVK6JHIx0
c59/MUaX5jyw4SeT+XKaVXQlQgXTohlcbCwKEwKyNT5811gK6qwqk1SlgvVjhyll
bf737Ae4UklqPGPX14nz7sij4lGVxsc+JvUUm0hxIqqb6V8MFy9ksT3aK8H+huYV
hH1iSewpIdYPTGhVpdr2f/6aaIgl6fZSkMuC6T2g7/+ssC1L789q6Dm2aOJhaU4E
aiOw/dRweDjXdswDzZT+hggByrOs3zpyeFtpp9sT1SZ++ufQHGH+VZ4v9Atpuljj
8kGg+zntokYXQB9ni1nISQF5EmigZYgMbRuQIC11vK6H2kvjnvIT1TzEyXyYKDDF
F7jrS7AjCDa1ewets/D6xRmnEQbWYjQ052LzenoXE7HTliCcQ896yTgBLlMItwON
mxRmphOHbyuiFOzeiVl5ZUcLskytYUUE1wfhnSuNXNO0i6MfOHsIDeYjMN3Ld03l
tVjKKhC5cWNCrkob0DfOp2a3L4NBj9E+iHFEpnySFR3ozoVZYWsF3AHx6CQ5GG3b
d+1iJPqaD0KTOMVlBZCwZ+NzIgzekpTgM1xxnPRpAwqBwFNqyqak2o4WVaP4Hsn3
GtM7gdNBIx0T9Y3dwiJMcACmDjoKITW8mLr8X9VNGCH5/oNWYD8bm+cGIXX/xqQy
OGMW0v1nq2RPBkk3KI1lKZQ3Ip0vj7kR70sTFMaEgNaizoglRLBJhCNOxRbATVs5
prEh6tQMJW4OrwnCU9L+tmgbt+wn8NZcmUSDy+TNTlM+Nh2D1Ixt9iT3WOgRfJjc
xng+CZZNA2nI6n018lB0xQ/xfrSck4sqCV2nBzmurHd0qLX3aIZv1fJRaF4bM+Hx
Kf3ceSP0tB4Y8gmp56+lykyujIUOTlIKed9D2IclRiPantwr/oKtn1YYigwugYlq
gi6RQNzdabEudez81khyLVCRLYDmerb+NTY8xcTXgEv+ScLSN9022fslIMYA9Z2H
RjkW03mWIcD1tLD1sufW6Px8VdOLQPz/ECMYgfQ8doTIigPq56huQtYAGuxzsYls
EJt329wtfpfOcDE6jQ5oBa47LJMJ6naWdybTM2McFuIKG+ComKuJp1IzPdEB8BbH
81Fjgjac3ysJZ2MOprDo5I1TBtnx1cEY9+kJ4T91SZZ3kB5XvMTg6MD+GqYqFpId
l0AKQa6Rpp+OJXXl6VxTz8pBRv4S04WU6Sb2Eu36mfrtTr4w0UE0wdaSMqcAjieD
w5IDZbSBGgJk3dOW39emtSvdFtqRzU11JkW0fl8qN/Rb2fIfkdv4J5QNidoaT3aL
3obvO74+HizdckUjyJaCKemmo9PgHRuuWmXeJRP5Dqi7PAVfodjIaU0Osn1VZb7Q
jhplDEjktA8qnFkmwsNmQ7I2s+S9zRTfzPSj80dVMM4nChvGirQjo7e9JAkgagDu
zzwZSOPqWdDT4t+uqwi7QpSsj86N91sigFtjM1LNlmmb0d+1yhsvhtTfaWWXtLD8
ZBlAOFSLcaZcRIiBZP1UmK7cGFNV9c8nOVEEm1KrS4kmae3hNGVP17cfLKhNZhmx
Gukgyxqq1yn9kM0VgeqpQum1rTfqvTRnD1v7s8WEh2lFIZm0WmhCbMPS6usl4zjH
rL2C+f3Jj8k2S7qWXiT+hQ8D6tccd6KVwL1cxP/4F5V/4vsh7LVtZNK/9EizRbF7
y0ZtNFapaPLCQZreVKdDMn0AuBr+yHfYfj1gtksp8yQHoTgRdbzkb7fCcXWvoVAP
59X1NsZDH06/CVTZpV9KIvSuvMxor23+yHHFtOq9aABsBUjYa3mXWg2GoVcMeoFs
Ryp6qnWRbMkdfphnnOSbuiGKniF83JOqSSc+WlRxHYYAMiHRI9s5a45x8Ep1YRXV
rNrtzIjoaKYMLBgkHgI3kLnJX7mjdOEOG37zTlXXrOuitpdQwZ3mGyXhmvjGPuAR
nIxB0YpP7uU/CZSo1UjXTmeolDLJHWEPb78whO6bORbnthlPTv25zl25q3IduL6d
VkGCGmdBO11TtAL+eCnz402H23WA9OHGrsgSBZWwK8MmRdFSxxbSuh7/ESrlOMvE
EMHpgswdc2uokxFdOFbSIhZHPk2J2OfaZBawMGUqz7mpTO5IAJZ26aOnYNP4g/dH
o6VKuBDARA9fs3GUTkkCMdm3p0LzZ8SqS7XHxWY+Vc9EOGqEz4paqKQkFRErY+0a
SUvBm+Od9+v4a+o/VUgp8c+wIvZ0Ised6yzunAr283p8zuXKCQKmga8Tq/sl298A
/UJQBsV1x9JEOM3xF6Up5GOsqWlAIS1nBi/i863+yUi6zrvJn/sg0ydeP9JpLLe+
Z87H2XlnjZVZC9C6k4mPeeVclbCbmr2/FNiKPSbWjhiT12NjuWfeabB1q0/o2NJB
zBQdsBiJazDiouqbtnri1O2/zgRvyLwtTvDYi5pHcZsC7LZxbsRtN5IowXezc5n/
Sb4nwIZtiu+sO6iSfLZxRGQRJTuE+kba2UGKkUXSD6KvIqPgwLncutuCAjjbsjyV
4JdCUFqK8S4p75PM8boMk4Z7PVhD8Qlwi9T2mCjz60RoKmRWl/N6elQi0LMbZ2TF
Snhqyw1xQwyAGiDgnQ4W8sydlc2KyF9cTmMO3k9a7PWytMCSpa623mhS7N+jI2nB
5u2oPw7Cht46OavcCOQXEPE1whnFUgpUqwyPxVlTo4iJKfoUin9EGJYUTwUBpE0o
KvsmfxTk+lQhNxW5c11S0KbWOXJXRChm5ayCpjWYYW8GnQZ/MSKowjf309DUWLHw
YZS5dIumPO7E0SOWgptxsiEvLHsgXjeb07w0PYZaAkHkh5Gpte0SZUY/AIhhcIlc
WuDp9XFGX+BXI5XT/QLF0q4EbT+3JSHi0UqXy1juMmDASnLCuLHb+KiCdXBugLCP
DFLj+8ivzG4dhNWnWjXFXF2VkmukmX8dakxV9P3E5GFilKQL2SMNnhpa81ul0MQ7
iYLh39NxZCBn1Mv/bcGQA2ATwhwNUlSYNtrs8uhTMZpGit3RSdxKK5dqaqux8bQj
A1j+wVVQRBXE0QsuJVLOOkPHWGweqX+4rDCIfch6DhBwiaY1nub4jFZw6FJ9ROY3
2HTKubAjjneSfIx59nVu8jrqBEB5O3iYQagMQ4pkoM8vOUygfVoi2h+F7Lk6EZbM
HkepLvpLBKWkiBT/xSameec0rceQ384UHNmI75dwe2keKnJpVdqBeFRHYprLrkDV
JTpnolovJHvkX0soAaXa5AU7ZH95N3OM1pceC8DYNw4VW3z9i2Any+4iLqW6AwGF
eOnHJ2WNm/W6DZTrvQcmFj7nfYr/6CNFnZgJ/lJjM7IVYBohkFQvb7niNtdty0Fl
59KsBSQrAHPKzxHiBd+1pcni3LuI61RrgBLgiLv0LI2c21QfuxTFCrlFIhgM1gG7
2GRpvokdP0idd2ygLzJ78AC+S/lLmeGrV9hUAb7p3i3XDZUiVwsnoZBFM3/1Wn/c
xMtuRAsug+tG4G0KN2WtTKBnlMWjnC92KowBb5grETdnzfIw+kIZ3wDNZvjg7QcL
mgyUjiTsEbBAHh13Z3htQGMGVYF7UCzdZ7cKKCKNx2z+qYbE7R0lDOMCjvUg9uua
LZzNxhTEYlzlkd0FoHFaXUuyYzNI5dfuZv5X7TDvME8+l8ocLIPBsCfxz3h7yaK/
MOCFWKXBn7VvaOmcmhDeDSnXTqoJVg3EycqXGEIA5Lt7rhZRVYhQs1aJbJaL7Ccj
DhqXl5ch4MBBcgv/yQeSaiwM0ihFQsisFxWK2IXVTKVcQXcOfx33yKvF7tVkvkfD
m7PvNLYCZOxK2KZ9E4ABecFb8vZCucbjidqdJlTa0mSm/4xPjrN8DO8ncYF7AQR1
QJZLp7O95WZxj0NOVYwoab3roIPy7i8HNOl0AhMvlNVp+1BcNnzHY5DHyZv8H9Ay
ZW6IND1cgjUoApAfadbWd7rEaA21A6RdT3ecrKyZAoN6n+QKv/D7uEpf8/ayhLYg
qe/2T+S4xZ1RtSO0lgbM8crgsjOHSVtCVDIC0i6eTudbLFFFxf64NBH47ZtXtC5M
7qm8v98ACy+gZR1hfJ5wjvW2zaTtDR5kic86XDoS+8GzzumDWqSZsbw6Lsc/KV3Z
wmGJPM9Uv5mQbLISGfW+Rot7jf63cK67Dw7sUk/Ryh9G1V9RpxX1dGtv2I7NcFZ4
8YFNi4r1wQ4K0kbcVmJQl9XIeGGQfjfgnOhN3qeYbTPn8vRcyhwHHhLP2Yh+/LGe
oLKUsytKi+74ZGj9LoyMONrhO8V2r9uTCm71OZOv0rGTDiMY4VuR1mSzZB+xMpIh
TnjFsDfPVRbgUmUEbdGEDtYDyD6o1NsvV/inGgf8yGAYygiSMHwXW9Ku2ixqrbB9
fGvBH99kMZMXyTH0w4ZOond1quNDxXRtsDt6mkmDoDlfpjibp4Zpix9bJE0vNx92
PhnDfKK2f96ZTikvafNwvX9Xds2jFQoOzur74bRC6Mg4ASn5yKO5NxsTU4K85Ws7
OX1rvsGCy5ZPpzwECqhx/Nl7Ne7lnws6V0XUN6RuEIWAP5+z38HCgqifVqfo+hdS
pi6x3PgduKIzgC3L83GNF4Fm/m5cp01jGZ0uMoS1LLbPhzrPty84gJBng+vOIYM5
MKA9EiHi6HtjSp6DfD5MdhwEyPcVyrg4dVgTLZH8NWUxSb2NzbDZD4LybJPPPrAb
pcoH54J4U+VFwD9qySWR8YXfBXbypeUAkEF0T6hGturs5psPMJz4kBAcZt4R99uQ
4daYfeXnB8ncw+1iZ5SqdkeB1BDpR5f8RDYCAD8hcpZtlu1I7m4/DZtE00278g7c
0lhX1nnPpEPnQOIup/WVIqS4p2c3iKfVettnT9DYmO01rJZy/oBb5i7QGxsG1jfL
TmrxVjpQ39/YOkAycgOcqgkYwq2D50uyvBoTd75L4gOBcPXt52mYLIJScZVylZtD
UWry7QPKrPXadMn0Ef2w3Agch8iJu5dSrEupUE8AeHp2gPsZpM+QELtKIHgzovp2
nT+36yzQZV4bDIvLNVwrD4CiH5/6h1LS+tkt+u68rtdggAZOqmlrB7Z5RR6caPni
VIDdAYCy5OW8pWKnQ/GJn8IZPsBGw0NDtpt98DlDAwhCNLigck/On5DQoTKxSkoo
DOc7mSE1v9eKQwx8a+Jbs5fCvJe8j3pKD5RssblX0yqw9SggNU2EoMngSFry3blD
olxS7WXZNpOVY5WuYXfIVU7XNJ82IGLpiimgsryOu7Lte1QhmvsgqLbjBPcBuj9J
VKEpYEPrPqhKvMAS/IGYHz8LwDs1r3zwvTrJO/C2Q3u5+aQ5kPZhzrOmRB5+L6TH
8Lsaqs8NbZEOg+ZIXfb+wWR164g28xnuL0FqzcXZsPv0Ju2Y/BTZ+0ys8HNKawJe
1X9DxeZ3jrSOWubPLzcoSNgshc7rIZU6LnuGcZB8Pt4ZVoNntH/q106nSya1CBvI
u+XuqkS2OAXHEGphgnPT9clorg9FBAu2V4WnhPs92hOEHSKPB+cs6Jys6/s0Xtcm
JKwEnfxS6XBfchgWq034mPUC08qoaImj1E3QwweK63EsxoowtVhsIJOV0J3lwaBj
steJafkgXPkSLLJTXNyEy4XDMeyb8+H9C541eHjXdlTJfJylmfohoOvEjcO5rU5O
J3oq+4WfbPqHfYruj1Hw5c2znVcFbwIpHoMo/0l6sxio9XCxXSPpgRy6ZQ4dkVOL
h3ndUClB1Enmokp1W33qlE0gEI3kXgEAy6RUXnTT9wcNY2Ac7xQjCvFH1+TX8VlJ
qsCwaQ/d6P8pi3PHWtvfIhSCELbyx4FfpgeGDZpUJ7XfVXepH1t6sWY+2t/4eloy
W6T98d7VMpYqTVCOll51AriMnlwzg4ox07ZbEBKEZKYAncGCSUGwrvTgW58euth/
UmTQGeldggzE278/Av83AKarpNhTVi4V6iUrH/fOZyaVNOyzUWU0l+SdkYkXBF9Q
XHRrUCTfff0zQb0ODxqtiSEBzIobXFkgkHKdjum5n1MuJ8zBmz6guqMBeRD3W4ID
gejeisdFgm4D2RYJsFo6MmH8b7NuVHZycEWETEZ/LPDNoiyTISsU17FotvuuCtdi
ppYKpuMolfKUrZQnxcZI5gDarb3Hph7vz6KUKjP+9eWz12CM66h3DsFKeIqR/+SI
GkfHqa0vnCvVuWTnmSZiOWhQOP7bU9t+aTF2rqHYQEw4xZaXCtwYmvIpGEaP2UbO
pUCROiqOmfHvCeU1Sht0xCZerDZrTGM4vrIIvIkhCdIe63UqkQRUx3Wo0XhhL2Vu
2aWsq7jJUU9kkwa22H9hAkxUSt6JW4lAePhXeftiU6V7BVy7gXqWgxTEQkWO3hJw
bf24T0sjzOh5uMwYnUw64EGpckjg+T5QC3ZTAfq3Z+ePmVBK3rXLnd3JrG+tnuaZ
T7d+xEnPc7iyqLn3MZsNf16pcpJ3VaroRdcud1t0cnHpZ9AnSgrXBvRh/UL2f8WV
eK41i+/0VzBvaAlaLcHuK9cE2bxLvB8wqLQLVLzfB6r2/xx+RZNlBAzFOhVNHOUc
ZIfLasskcOFqK5Tveeg+8VVjTOvcw4Q+Ekx2YaGQPwV/Q1kHXQpSuibGH7JWsuNq
4UN2ZsmWV0BbUMc5FJaHoUW2JikxxGTJUzcLLX2LBVcj1VJRGFaCJPC5ZU4+Pmq5
mmH6iC1Wu1ZgDFSAHOHiH8TFj+gXaYK8b093hSO6qROzahZGUjXy/Uyh9JxmVeSa
/yu8XwsYPDSV/+pM3VADuRwJ5JB6YGf4jkwgHorYnlhH3mAUNm0GiRr30oIysoYo
+vIUazUji+085oekJ/M4Irfl5gn9TaVnKpeGj6Drifuj6/xes2oLJQk6Vv2WPAgm
aICY8dKbHqM29eNDWZ2qU93nhCy9fIs/VrLBHt6o5MBs2opUtMi+nMYp4z746JZs
bT8VHXlRqL6ey6Kx7qK9x4Y1N91x+qRdhzCZYBJcW0UV2Sh0OhUUvcPlU0sC/9O6
iS+YaiVIwWw+gniruivH0uCYoDToa782glYw2FzXzdQBDX9ByYtsFD3RwVkwdMyn
osb/xrbW2ykn0ZRhUrlwrK0E3PTwoCBT8DO1v7nn5oKwCURABMSxlnFTgzGO8SaE
pM/zD6yC67ahorTerUP8WUXPn3u5Jwmn6r+KQBAvggTypQsVY3VIHCsknfooO/sd
GS8HC/zthNggntt3e34CWuauohl5eb8t/hlG+1bU2UFeRyJZmo1CcPFkqfZVkH6x
e2phuqinfbotwkB4OIVzDdG4vvsn9sIcsKaqZ35M2ptDXCVKzZMWyErvK0xg0rS8
nxgMT1kZvcVF1PIlzU/zTfgB7mE4gyVRt0dbaAxA97blaUb7gIj2j8y7nLtwC/4l
6LwZ3PnScZUoa224HVqWyWbNzDzAqChy04eN5Gq6OwXzFlqKJ9yOwVIQ1EQQzfHn
81kKokwqq7ibfv/9zrAxK3QE/nP+FuBIkDjKCDFuZB5KA4ODRYKOXBNhUQxbbVr9
1yPoXTI6P/c6UuArHtbaCV9EXy498EtbiJzsHa4FYiCyLGa6OMEU3B/3u3SlsPoG
nJPGbZF6T3YYHzG2dNykz7fpq+XqDYGZZnWYG+ddMn1c7C8xTVuP84ByGoyAGhXo
RqcknR3XakgP+a8vmmQvJqeRVB0vSWDtzgYN1PK3FXpPaWfeQ35JzNOnGUh22CCA
sDAlQiZ7hQ59BI5DNFGMSzpg6SOh6II/5ygZm4/UcLIHjoUimmkqh9neBnUEzMdl
dKdjDlD0bvT8KV3Yl3owmEGtayTtHoMei5SbnHHXI+fB8bBif5Cuf85GhfKhi3V+
0CsQjJxWFK+YBoDu/6CJR/LIGbebMIrJAyEIIocmg1K7HJmIQbbJn4Utliduk9pi
0hlgOy4/lFSQZGlBlibuto0Cgjx0XprrxKgWSHaOHE4/8kmBUZtiQKVpfTdCHIAc
w9NJeN1xMy7xSq2jV056WMkT6t9v5OdagYaeFF9/2TbqbmKKuJF8KUmlwEzgVV1/
UAHUz9aF/NJ5Ju6cG0p3DwPKP6Ps+whG9oqB7nAo663JP50G9+IFUKwQIf198dv2
mAVaabEr+Qv2KA7OCdkSYoNnk2C6PhccRpaH1hsUygwSMOPWeoO61SfyIuj/cSQj
SmaMKJG3HwGFd24ASy4L8dJSF0Du/dekvkMc3JyfhLkX3XgmmiB1wYufGZ13GOfo
Tc8N7tpHepHZMFjFtb6NKStx/iP3Rqovb4AfVBctwv6UCcu8V0os2IVOxwWQixEJ
VpUHdLSlKGbP47y7fH+cYVsMZkhONNtMNotS9ZMhT4c0FrDwj4m8wqIG4FFaKr4X
UdZ+8RnjPtMad2Vpbe+V2KwLNpJBIBTiG9ifocR6nvl4h8TGjwTK1rh7Iux0Z4nE
489wjG6W9LsbdhfxuJbpF/rSoCSzWWYcGvyFdUAziB+SY5nhDozP8/OiFrEmoudX
oOHZU7lut0T7KmK3kSEsfoHBEeD94t7dO5D0LVAotjaFOsTL9r9+xPug1fJHFa6E
z/NX7D9g/p4bx0Omk9Ka8/utRKn8SRcdC8gAwSGrn/KXGBAP1gbLon6SQcK7K1RK
A749YYqmcgW1z9y8I3uSmH6YjvVoBCg+BdU8sjn5JHPr9Z/0f4o2QTD8gm9trp31
gTpNDHDAV/8oCPZk+v293wHi8PfVdeJbZc7gTYv5kruJaHxwMfB6AMS9WXUoLujn
3uUI8Ch6hIlhjzlnHs38/hkfHkLzRy/VvErZwftCBhKdkLYeyrHyOP+X6D0VwdbC
T8A+w8FZLFDMt4KY19sB1XKrk4+nWx+87It675dN8WVnJLKZ18KQQn9PbjG4HMzU
rzi6K2b1EQT5JEKbHdUP+tbU8Q2ojwrXv9Llsqo3Xa4EsN9vlj5fDiI8kWmaAwB0
4myTjf6saSjExWA5Kun9C5ImIMaeehgX1hbp/I9Jv/9v40EUCD4xX9vZGzvQPvWG
k/SyDn4067pzOG7WWAJGrZh/grQ4UF9Bff+WcIPQJV+XAvI1qzwOiFgUkYPf4SKt
iS8kuMXi1nRflicUjbUabPpepz8lpJH/owFhx0G0D7MopUomKvPBwaImnsLqbUQL
QNw3XDLu6cIH7gu4Zi4caaYSD1CMlUivSJKFqXUHsUZRPAB99JalpBxd8wEVvFmO
Gh7LMp/mhLY5AagaQkFOqGoaz17YgFI2XUzJK+oFEDV0dVdkZ2dZ12zmyhxQOxMU
tK8G1yObx9bSGOhO0j3zl7RiBMT8AbDJs+ssjlFzfdqML6u/U4xhWVTMC+LKK97S
XTYn5xD/m0qIFpBE6km1A0Gp2HhyKq7FYviAjtDCk0tnuewHmMlPGkUYgWVVBMDS
H2Wxu4Zd4Qmg5pwclaQQaXmtuuUgcq1ehVRxxd+ykmYpUKeRsc/ehRUjnzRlv71p
gnagqnU8eJfC9PDVVVpzMbAf6pRJVFNW37P+lAbetmGAHJiP+kHTukZeLhB36raZ
QWRwL7TZEpaRFkeY88JGHRL4w/U+y574fZDAeOiYqlLbmz2UzSwDKerVKKxdMjKI
Dsjf6qhAKUlH4FTozn2Pb4YwmlwymGe0rSuVFARL7xK7vwWaIXqgmL0WDJs6C3aC
cjO5rSpy/7eqs8nqreO+4MOtv8sFaIAsJG+6mtg9mBgcFLuy9LeMLJYRXuOSk4ih
khyGZWFQKqRh3R1CQPKdFo2VC4GRZQepXanCqjw/sFBQjDa1w5K12g89JiMCDk2p
cX87WLJJNo2cYO1HcqJkgMmypo0n0t5jiiBw1PEJdT/1KprSzwW9xXWVQu7mz6uS
WNPQF9+Vhk9qyv7pchYaUt7blDLr8c+TTNv8GJ2tTM80PnIlp5DI6UTwk2udhsTP
s8GQ2CY/I8r1BOt9rIBFV7QGtLcvnravUsHcdMLNM1xAsYg22OZ1TGBW9k30uvkO
BWP4iujP9UBm55q3Ny2rKOfomWfrG6XCR8hBevZMvBNHjkUosBF/juizs7/wjJ5C
3OFuwbR+2Yvw8uXF72cnqMqGPxG7T5e+u9RkeK5amuU3seJXI/Ih+FOhEsT374jW
+vLZBCJmIy+NqdEBNG9YH288LxgWJxCVJDaz7nF+r0VKxTKmU1+gGJa576mkXAbm
SvTmT87DfWfA+VXXB5uxHyIvtCGOxataj5ZlHgmRMT0vrE3ko9X7s699GlZKp8xO
Zdo+AvVX/4JQKOnxfex6K4fgR6fBzPFsoU8cajCOiEx1qEMlOejEXMs2kDGVFWZn
1U0YynyZtavfLiv7Yc+Of+4tGQmX5F3JC3r3ETTAlSecdO6DEBHwGoH38pmjbYRf
G1aAntmmuTNcFzK8RCG7YESt6vpHeKHVKKfSLAUPR152TyKUHbpYI70zeDzycNHu
EdhhhF3+LIz9amgM5Xf/7Qsr7/3/O67QBuFVW6PSBmVgY/xv7ruOCZnV/5crunDn
bS6ZDNpDAcWj06Dn3CjDbAO0LAX/eD2c+N1yzXMnVF6Zo4XgX8H4y0NExDliy0PF
+vbqeqVHhZ2kpzZ4z36ID5vrg8B2BAW500vwnxxP7AuJK+2OBXLHQhjo4p0u6ppr
UavW6IOQsFjaJ++J2hX8LYpdyZMlrHA5HIvryyg3cWCc//7t6pa4yxE2n3k2JICA
yTXqmaayYuk9oczDnENupd7iJEeZO36fCHEA6nlggKOYsg+SlTzIhOA5fIKKWhxc
rsPcc4FouF1lwOIh2H2XJBsiFrEIECykaGBOXRc2lg/FP3iEbbtAvXPXFqhwkj4r
mM/K7MH3gRNjUWnFLbb8yeFMO+FwnSbXyIREDesG9VKEn5JI5kRk4sP1+MQtScvE
/ks5USmN/4dzmt6UHyxx8wvE+I/++jjM/pWzzN6EkJcu8FNljJD9QvgV9f35Jd6l
JHNDRQi+tIGkAPs9flkSleKkA3PzvRBRSWYASkSBzwcIbgNKvn2zOBZXzMq8FBFo
gpqNAL+vem00Yy9liXRdD7LN6XmEY+TbDtawq9zrfhA9UB5iB0Trlm/rq9rs1ueR
UrRjtgdccOCNPFk89klqP3t+OygX6fWgK8iuzmC1+fbidUUstMn12ui60WS2DWVh
JnoFpSakKMkPUoUv3Ub/HLDRXtI0ecdgowsQvlZBnrgaRTqClF/XSIB24ieJ64Kt
LNKJaU+ZRy1uw2/geRek897lgwOjs497Jq4+RwpLg1ysNQYXwK91e/cSenJOESKt
2tbvGsc3Ip/prXhjSFnPBd60wYQZ+jTU/PFak/LB9dqmVkbMfimLm2Otu+17ywd6
lw6NP1xQ3l0BS8fvGldW/+jAkdeIygH8p4F5eZrA41XpkEIl5sJyGzRk8oVFUPWJ
hMlWL4CYbpwgI/lhGhEXEMfP2aJzadFqnGj6WmO37DGBAQOMjsFtOIKJRPn+0Fwe
L2Ne0oM+lIBrOWGVKoyovNR+Fg2B852HshxwstavLjEHTbf4AnxjDK02oRW2TPWE
Vx/01CaOT1/lPar+U6nAwkOafvj7Yk/1ojz6OWYSkeBfsrE2hlxhZ0CkXT/AxRzt
vtP0lFV9+QjBn9OeAUJ57Lt44Jt45b40kIuMTYxlIY5wL2f8MbWyEP+ZBD345iHQ
H8xkMpXf00CF27cQr7Exo7ekM7nQp/PlQIPJogq+7YBGyU7deNIwwqtXRIL9Dpqn
lHJEgE5cowBrUcCZum0v0x2hgwztmVdy3EZP5ghItT0nkHyQT9Nh24FlAIF6cvxy
FSBhekT60imiA1Ch+ewt+O9Jx9MD5difyXHGQo+VLzjZ2KH0LooINtfZdMpJx4kG
8a3uDwjZNbWqN1x6nIxlsAMVjRABzbdVxcVII0ocWBAP+3Vyf/LXy0bQzt0Ucd+k
IPwMC5eKyJjQB32Y8CpzSpHpM4qFUGWIzDjZX5+fRi0d8kDZKyb+EZFiFluQSYHX
6KwZlfH4yvd1hKDyBKfVTgm/FPODrRcmJgIesYIaUhK+dgf/by1fE6a1/TEVt4Ep
qTEt/u8dqdO2JrGUoDhCnF8DQ40nsYkU70jhsOllcEXPTD9a0XZgDzXnMzx2TWuQ
p6t/KTEXmJtpux2guextOHnl8iziwZtM5SkXUDvA8CimXGSFDjKiZLYI5QHRuGn6
mkPeLQh/bazGm3SEWUbQVvDp5A1tUVhaGBwdZrZHuEZ6/wn/klknYkQhpUofzDAz
eZ+WiWNvhpFKfgfC95BJyI1QTJRwZSECpBSsqkCce65PTWureGUyitMyXXiFLBYJ
b23X7KAB2thKSE6nm6N+CXb+27t15AGqlhOA+YoURxQcAgUaX+3HocxGDWkUtln1
/ymOH259TeakaDVy81t0BiagYZSbbIHcIX15vHnWmiDSovyJRy9mf83BinPXfNQZ
zAAZsJMu+sxzvf+zKws9ytR/5cwc5cVcWmxVSY0yQwAs60SSL6cmvkqGLxCSsJXv
dYyZfV4P09qftMu8nzzV1lsmxzfYN6Tb0mrNZnQMjOndRlM5Dhj9MibPSCTNRetO
jzJpj4F9xcKiyhc/2nMKAb8s5RnZCRcLUnxryYQPD8PwJEXeSDgg9ivU02rN8Vme
f6CwwIxM3/MdBXxpq0cSG4kiFIOo59Y6BBaAZfJWj+2QkI0k5SmKdD7NL8TnQDyA
YCkL3ZAL5t7JxkUg5IpjRzgEexotwT0cpLS3xm7xFuqNJvTWFVdc9fOdQ2CpAA+I
j6OB7vyS0K2mDmYvDYOce3P0CLhMtxr9lJ5h2f77ShtzoJ5cLJsIVr2qAwcil6wU
rdGyAJcqQHij9dQZtgjQHJygdGZ9ioxzIQM81yNkIi1DZb7mRuU4gqThYqr0eq7Q
qCUs/2JDyVld0GZpcF8TsPSabKLal2Ek6DdZhA7FsDZmWzRQC5OsgjERj520nGV5
Xui6n1bLZIaAr7xK/NbqrckVe/4lfOst9qfhlPXKHUe7EtfXKDjKKV1Xg/SVHzPj
axUidjg4p/ZEU6r8j8hn2xsnJmSMXAjcuL/UVlBz8sWEuKC0njlZqQ/vc22DJh6U
MMvMsn06XUPMgFic1uKXWW5sb6bbIBhRJL5gw/PviqcN8stytdW4nt6HlssPcrjE
NAxRwhr8avj/ixjpQJPP9o16iAojvea5UDuTF/Pdi6KO5K+EXezRVlNq+8HA85La
E6eDLEgTbx0k2sNiQpsk4sFI2c2+hZE2VcOvu5y7PxOyVkATUtPZew3bHpZuwX8/
GQsMxKDTlzT8374S1uMR678oaw3PjB6qt9EMOv3ywtHKwau+bIKIVT8dIMsjvqF8
P2OKz1AiBQAgsdO7CSg8jCtM0fCIMqR8B7X/OzdAwPj+DGDdEQTw3UGP4V+9NH3F
/YqQJFN7IsVKSPJ7KtN9xRc1qwBWdG67c0QM9Sw86z59mQc13j92JhG2AfwR1cF1
RX12D8LQyyF6C9UyGceC5hngjL4DcD9mblkESGG/xYMZiKdoq7Fd2E2LOymJttsx
Z3xvOdCRXOiqaI5LIOoK+T0hlEYU7mw+8Tm1/oh+RY6CSF11CiJ/CS8co5mnP2g2
9ph+fWffPTWLnrhTYWuZwu/ip4RTk3uum8YDUeXSIO/Arcxn7VrziKPxX87orBjx
Y8wzEalC/jCELS/DMbAEYff6yVmhHXmMFyHW0rvrYNFOUTbeH3qmRDAv4iUCOU20
tV/SPJXIPk0QDFDklJEi3SDiM6yPB470WneX18EEj6TYiIGD/l45r7CweK0EA/Gu
mojj4StJ8vuOGC0+XQZe3Z7UhvkLDiB/tN1xM2EVwmsggjbhqwUw2pB/MzJDl58h
NwEjqx/YeDhVwsekq5GVkjjS3sDUHsu9/2Y0K7U3QvtVyDMmgzgr8Z5UsOf74fjF
BJvMbWy2BuHMVJm3dCnFxY8G/obE4mFEJ/KxfOagtltt061v8SpR1to7zVvyHeif
txK+vt7PzAFTFLt3bglv00EesEOUfDVp2cACZ0m7mfAElckM+hLOPZrsmqlquhhg
yKF/2UrEuybIwHcljykRa4mAFXAGy70MadQhQhs9q5d1RLFoOv/1DN2q+J7mbuJD
8luNldDF15eEO2TRK8ryrp6IXZKEC/dniWEmM8Kc2iB8DuqzKnYYNTdwI1Vrsqdt
mkCSGr1ouz8FnqjH1sxwzD5F4KOwG6IIXkp7AHYV9NG1W4bTeidMEOE8xV8z3oTk
LD7FIT6KQE7xcYE7rRR+aw5u/vQZWHlmyVfQc27HDe67By5vzJLg9M5l2uSM/pgC
ddH+/GxKTGubEDtAGagJSRc+3xzNzVNsk3pZnW2FPwcndgO7F/AWZBnamQ/HSN5I
jYG4tGlWrPzDmUZIPGGFfCpLGY8yQ7FsYOBuitRQ3hx7TPNzqGWtSbjUtisZ0u3F
JyAfGJF++LeaoAcT1A9zqRin1yVJJwpOhwIQ8ISqXA9YvrIcTbHVo3bKTVpoDZGY
CtgpswrJBGQ60pkXSzLmQHalskqbEBpLLBDYmvQftxgXAn+XDqJTu/To06l/ib97
jdx3yDcnw53zeMMbO7J/p7pJosXXspYAc/ecOZu2+E4F4b0uUmdp5c2bz//AP1uY
Urz7nHl5eLqdLAFxR6AHegfzpLMIIrf+JVP7A8KH5y2nUtxMyCUFME1mU7zfqcCP
eCrcW2TfmPcXuzt/Pv5mLtS4SJWE4VTKhgRAwASl53zCBkkbGHnPX9NqxHHaONrj
ouD53EmHohA/oYyj61/XYwcPBqgtDlXYUDwvZjX8+KO1v2g4iJ6hMe24cg4TRVHG
wJY/XA/bA/mvfNq+CNGFTX5USLMv8XtGDjqh800/q+2jVMsznpoKwQPDewbOB6gl
rcjjquw4oiV7OvTojXU1T7RqaFLK/g04kiIl5dK96sa+ATKZJnMVk+abzKKw6ItJ
EV8cAAgu1KdMhG59vF4SZ/wCc/27Pf4I+3HFpXkTKOUTwWl4ZLBFHxJnImLbgmkG
SnjSofpnqp6FDztbSl+3+wMl9cNfEyG3XeGbhcBM8VszCjeqSdpoAnDojMG7ucCa
m+bAyHDJGtwZhOE9LnoZRvr1njg4R+i2tK2PnrRPe1M6aq5Px/IlsV/RvHUMgTYR
drXAnFGyVuVNWGPv0ifBfhq/ne+eKgZ4PFVoYJ/5kCihFmmdZRrz6IgPRU0BhS7b
XMM1CQukJbtfcttnxe/SwCuAA02ldgxBEpxFRqQ2AUoyXyqq0mFsUIluR/lIVy3M
f0jOuDWZZNSc7Q+lFc1WnSv8hTPDmUMM5glF5zVp5w9K9UjS49XWYjT+ZIGbmFBP
44yJ0pdY6aEkTSf1FrlwPuD4p3dLBUyTrrcDbdGEKP/+oaJRc8B2X1u0VQWXY1Hq
6T8OkZRO9n1QctF++oS/gJabkzwcLhzZkn68AinYWMZ9/tixSaLEuMk3MjhAUZLT
I0ZkJ6leF6eJCcKKmc5QaNmaRb+POhwLzQ3xTYuGm7oL7yXCLuSgqYT80aEwHWS8
SuBu/Lw/08gj6Jqn07FFIyrI6kEB9o3Xzr5Sdyil+MYzLSDnX6i2bO2wvQTDxraD
Dnri62j1waDwVrhdumr6XqWwEmAJnyFR/lTJtSSIxjy4q2qG4wpdoCOwkFlYxTfx
8oJzD2iZMMeN0EK/lE2hrQVpmO0HLA4ZyZyjfRvjhuqB4UmHp+XICCQqFX7XubZa
1CyTLGKKuCkMPZIw5n1dvtMMDiups/45nch0A7rQLoJeQ1mnTC0TzFxzATxURhl4
KMhCl8Wke/SEyN5RPxPWK/QB1AuqaRlcbd+uVw8VUkqRsX2vwzOgL/02IC2DlwtA
k4CyQ3JEKJDWjHgG+5n0Z1kc3TOpXOupBtaDPfpUuRpJlVEqXycZapZQJnrG3uc4
768t9MFnVW41CR+VXWakBfbFcKb3L/PHRRJQnJz72zB/Mj2zH7PaDmyvF8vRSdrP
OO9obCKWoFHeAnz47xTzVkd9Y0NTh0UOGYrEKvG1E8IGYsqB2am1h0nDVJ8l7dA7
d4BepCXFpLfv9JpC5yZwH/BKLV7vqlQOKOKHRwLbSIhNw7yOMzR80eTfayYXrpio
/gFE/hGSYlviET/jxIH5H6ZQns8PtYuHTSDsqlP6uHyjufotDo28aBQ5AX4JJaRD
PNF/JzCLPaoM3uLZJuJ4954Lg7VBbzzd/Uzf41grHshT2DuN1ZKfVfQSDk+M0+i3
0A+yegeAMxjE1lGqWeqhYi/dhFcpGyvUQLrMVwyIW3t08Hcnu+PhwRrcXb0zwdst
oqxp2zJ/t1XTqTIlMBfrQ9fbdwZbIMnELF2H0n+p/ihIOd8OUAzGIPwViPdiHJ9T
J/iR4WpJNbaY0P3nOYeIFkrwBhRvX02WzRp2ZnBGYND8hn1OWz6zZJ8dIkR/Wgh4
NJFFexqkanjqHEQK8iUCRmKDWB0m/WYBFD1XDMmfD8Df4wPjg6QjwCLip0bPa9lN
QLPa8QlVI1Kfxl73/FpNXZ+HzL0I8XU/W2GaDbY8SdnrbBaWoX5jcLsyeyhygVAQ
0SIKD9CRpcwLFVmL3ya9/IpGbExyw16TcxGHyyaGs8oXGGJ1munDDBHew6X4QtT+
Gw4OILfEKoPEXdkjZIVUKAS8cEfoNLEXsZL+iLvDNPabWNXo9SoDKLjdKOrDpwVy
wW1k0TEIX5lk7qkdtNHTNSlTyW4eGN+aXDe6qZagXiayrqQLDr4ApTCN5O0MagXO
oue7aBws4kMN7Z7rgfiDs/Wf+SnVdTKxxDRWtIf/E1jzt2vClOdNa8AhpCzKOGqK
l0KwUXtsx6Jmgg8s31/DWosjUu6whIOqXroOFnIAknvkBG8KqG/MxGPn66/YSIjx
Lsel7ZLOWrAWw0OzAedG8X4P9f1nfE4fyiza5dMubtnj0vt+qip2+6mF/0VVQ6X6
d3I7xEQ4fBllt9jL940C/vXlJ0WOpn7DMh6zOg3HXAVLtGq9ATyFbf+XK+P4fcRu
6+BntnNkksrlKSFtDIOgernMg5/eQtoqPwYPCYawNIirzL9+PK0zMxYjbxTcMbnI
Z76XRjyo/rQjDykx3hG6Zhl+VCpHdUPHhsEnQdP9VHybMkFrcxKR20d3rDWELxdQ
U1rwguXZ9DYL7eaV7HNLhdtnkfp9wMj5uKIURu4OcHon800RcTJrFuOFZfDPMJeD
xZ7nqdVrlH0QzG67fZ/vInRmZ51343G3zkCzCl2JJEvp46O7g4dyV+bNJDti09ZD
04OZtGvCef+mVQFb5BFTW7xqBse6bHQqCI+VXKLcLlIxW4NYjyD//S6do6giNo0G
AhEsUxA/utWVhPDHbIfl7v/FkZiXNHsDr3NoHgIqkXIVHSElOE/KDz0hh23ApmE8
GfDSSIm1+uLxCibIywUvVSy2g+DakJkKioskfQj3Rc6577rEiQh4BeCRCv4f/Nb3
xDTQBmgVsfOqmGcvdEzp0B6MQXDIc/txzFdl4JFYg3UwmhB8SGzEnBY/RfNx5aQJ
UA+rjQQJ9CtJe+TIIw3RTSzjA+CNgc0ttb0FuCEgAPIsNn1SHHB7f9R3F3vPRPQ6
6btVMFoU91W5uNiBEabrbpAgeqXxhbcw5gzva6FxZRple3GXUgdQQHNPc25hpdrl
Xv7bxjE9e49JM6UMQ5doUfMcNbx1TG51nRTTZ8CSf7+6un4HT4AT5i+Q59J9cDZl
EI/lFRDlq+ozxsHozs3AdLSx++vM0kJLZo0KgrgBPdo8/FtcWQGNByQvuI6F7lTR
S+SOA1jzmmHhzXmewkxIen8fvJufT4fvNrdRdf6xcwKkaH4A8uCln9+vD6EXmrMs
PTGEAPBi/wXcT4ksq6fHVdpk2G+PEosfhKCyqMkyDjfXktW6Na2ElyQJ+6WlnPsI
+IkkayDIfqfuGNGAOf/DXQGSGGK989TVrrm4S66F4amkiXkurdc5AT4qhumnCC17
uSXkiFgMy7kBkaZkqdRXFONYD8HVzOKbDqjjxz4EY7Vi+6PM+35Xs7rcOUXqOToN
4TdeY0KnigOuYBDbvoDndDuGOWkMi753MqzZU6LjPI+dEsEM52lzpMrpDG1WrCap
pvZ6zTyJ4waEvK4bh62pfOJK5fcQDDQBym1teQgPDA0S+GlQp0estYtIAFIwOQrd
MIg8bBQ4dvrBHd0pgP2qVVvwUbhxsmoI5fIz3uygv2c1wlSISTqQoH/XHj5LMADf
lJZbS5hs4mLGgW6jCUyHEaAI1oaBHaTe5Tp3AVU9weLog8kFOXGacdoWWS2xH7HG
zeQECheDWRoXkpn2IV2LTI1XyGuNCV5928n0MpyvzTw2SRBw3l1n9ZlonP448jYM
C9o0viDp1XRDh9BpADh8pq8YpngqE+bIsONdcmyjY+th0/DWVpVymrsjTm3gsri7
g6hMtMGrmw44xQZehrqeF+UYBg6JMDzyG8/ZAXxAY+Be5K+e/1uANibzDJ6lGMZK
17TPpTPsNcAM9YrjuT5r96qAF0zIm8oPUcFyF+C8yzbG8xQmZZ8EeSGvqmxTQaoh
v2HzQeRaZtGik3U+VrjeOjc/LegmMTDIQ6s3M+AGvuBbe2PWoa88E2+vd7VzL42W
ICdst6smbvh8UIm2dnWVYZeCzHh4VuMy1hNTzdgficqkDfK9+hZIPj/6UQtfi+8R
puexOYFtWtp1dGWSl5o+OrGL50IUw9LdwRkCfMv2/R/uyAupgSYuZdDalx59KzFr
bfdq9zo4BYAFhY/W6oHTJ1Djueh6OiW4yGkgWKkGEt5wq393ZGvh3F7KatkIDYrX
1mNxfGi+BsqYq76mzrPxKEkMFRaWrWQ4Ix8md6S/+EZw2gB1aduP3Qm7TCQFKS+2
24CdlnwsnkGeRpMTeg40lDakcCv8arKHlvgNOuolUn9Fg/EFkT2X4LuQoLkGPkmW
Y3umzbmavw99R1NY5rLLso4CbJbgg57VlZtYHSsSa5TCrgmtQtbOO88UyV8kyoq0
S+qf8Do5IuEphegG7t1z7V7PmEUPdgsamtX9QAYY3n+EyjMc2/qc22MFOCTL28j2
+yF79JVE/UlH4t9hLb78w2oqZtwN+octLuxNGNEI+kQBawOi2cJcg0n9mfuDzSpS
OgLUrSH9k6lz9EAKh659UdM6Hd2p/gUQNjwag/3lybhjshIyh+HfLX8mfSy8r/uB
GDhpXb8cegl2nChq2BPfGQYxZ+RANuSAURHQlzSPZtCuKQ3L6DEHZoWPX0iULbx8
FjlfdV+hattJQBSGuPpGvBcms3/0sA+bzUbtbf/TXfuf1OPZmjPHwM6OFPAMrsCl
fhm5MDEUDwPc+90VqOp3mPNxZ2E3QZ5U4LqAr8RKWOTS8XPC1zmfQjNESaU8T18v
AnY//0aY9xkN12yvnjUCJ38Eh/YtKsHph2DvyFiEvILKCZwDToTAkYKVy0DSwLYM
bmLn9SwhnVylib+2lGaLXeRXb5Xt+80LSilyHkA/2pNJ9VwD5uPo0XbAFRbLENGW
oJbczCcVJu2dFXmUSGcSae72gVvTqqsiU1diEbhngJFwlb/iOVYTTZylXqpPaxI9
ktelWZop3HSswokyj1EstrUmKyU2xz/NTicFFOtV88KeSMyghxrrW9PjGmpweQN2
wPUsFsYNwXQ2g3mouOAnIetWLAoT46pReuPjFMIdWWpUpej1X4CE8EOBCCV0gS0d
eDBGp8aNRrR2x+TwQayWFKeUh5XnMEN38bJpL6Kg3d2L3kkFvGJGlZ/sIOGITabp
KWiKivFNthvmUFvlbsETonwhtjDfd6bImz8/9tmnjj5IaV/I6jh7AiquInxRKFED
mxUVyJ/+rcU+eyfb312cWBHA1y/ewfY4ypqXed8JKSFhleBcVwWNQiSTD2rdEBI3
lVUklfohdLzSFapXaORbz9sdlQDlAt99M85CX06Zj0bvD00q0T4wr06VlU/89j3I
TfM45kSNDh7pqdgrtmRoP8Iuhv7pDkmmEKXXsoQmkMNGi5ULPYQ46dYSis22k+Rk
82cf8Do+0aAMPhkkRCSBtnSRR+A/AdlmdEEurnUQPGC/xSh7IpB9nvDlsZNQlwaE
Oyl90G2vLjjGNSIxL7ZXszSqCOKAM1qswiLoRfr9rFSGpszWDhiTdplKGQ7OMRtW
mEC16LwZj3748pYecT9IlIUz4Cw4kbI15MNQXSMt+mlS3c/8Fe2pFDQ8icDA5DUA
XYLqExmfyMYoCrYFeVhscwjPb7vOcF87qpJZioRGyZ8wMwPmDEHKAx7ONdF+hXAr
qah/jCTnFfFdxXZwvPtS5f7eAAoieyX2A/FdT8Cr+1JXdbWmXHJixf9yAL6bWW62
zuas9HJ04dXdeJHZgaN17Y/kAatD12sh+X7tKCEJaPgwoJQKOPo+/JhWj6i4M0yP
q0/7qHynX7hXxgeUd7iXB1AA92AZoasbETI8BkKuC7/+aX5/pNx2RbD1lgmKZJOG
EgmCoPhh+Vegppufy3tptuo7pFjnUSTDvDqeqjVwpJZR6MP1bTfY0uOfufzN+/n+
+cjjxcEench9lDGXJgpfYWeKHesZ1s86g5ND5MBFzhwAKoXfN3V8PR/cYjTbPcGW
EpGFL2Mg3m/zuVubhvq6E/g1tozV1DntgawfcmiQlqi5UFwA92Gv6DFgoXUla03u
+nWxT2D8i/fW6V9hXTh0bW89YtVO21+j7t3rQviouG6fQrXN82VxfW78mo5AFErn
0G9W+sQt1nnoF3fioD3G+FYCDKzKmfvtQuZpzdoLTVwnhcpkYpxJ/8w7dzFcExzT
ClXwD8tEsTJvxRGspOTRJbb5/VT+vvVtTGZIU7i1nWgTmWzF22XJlOo5SSdKIaNx
DmirPR9WUbTb1ouZmCh2KmDuJuKv/h1GUXvFEsZVemiDBaFBT73jQx55/0e9ZYGg
2BAmCEqNbrFguWY2HiMVQ5IdxtOYcQNeQEo/+ldFqOjCrmX879OU8J65tgSDyEpW
kakXgjEhuCO6EZ9nSA00BG/ghTIAMJUuqKX0GMW7tinM34vtOkQA2ZVaTtkukiGd
WjIjCUlbxG1o+I/2c5gGfgaGBrbjNvpBVfnXZ4Rr/H2uluD95trWEn/IX+pjLvej
zPFGLJgYd0n22ZtJ5g9xOClPis6VPYpYs3qrJN7YMZZCkTP8rKclEEpW7wH1A0VN
nKVGMaKfQQTrPORkppCXmIv0cvPDzist2try+z3VEyHcDkrQ9zvtaubHvlocYmPt
iiT2Goyf8utdS2bZIRREEbvd+X8A2nUXmIWGhW/piYOirkq/czgma9ATRhLqFZ/h
QOKrgyQik4mbKPdqwOHU6CEDtOh67H5z7b2Ecdj42jFbyZEYQvAEOXz1uN3JX6Kw
cA4c13TSbcu1C85SVsiGvN6NOHoje7UW/gmOYOnBdo+RLVXc9KDa0OhdxTdXn945
ibTlNW240EXKcIg+EKoRKEa+Kbk0Ku3h1D69Gid+i2sAWXSeUsRB16Bu1HBfOLje
ZRu82aFkT5vnkAhL3e4o2AHfQ4Rzor2Wclmvcykq0yuAa4LvMnH30eOPDe0THFJs
VF3WbNG3AorWSDrZr8PEpL3suevzd8UR8fzXPZtuYI/BFofWuy+II110YHg/ljYE
y25PGXABKApWhufFiTgoImhtiXrIfQOFFg93uO+twIWQvEas5IbGV6V9uW0bHUTf
haM2fkv7XtINfqb29eCGaHAO+sJ0gYgPKGeSFD7oTNWUTVuOuNB4OoAy+l9a/izP
QE9BM05NCbnV+cekczvFLRbhGVmNfIYf6OTt5GoPFYM9YL17QaEpADsjizybuo2j
Ls8ccxCDWk227AKt+KzqaAXMfkvm7fTzxweABYkT4jec7U+Ydj37zkYiKoLmtHKn
Y7h89Z4lQVMkLvXUlGeg1aGXOFvSfX88g6yAdtT1Uh54w7sOprlg2my7a7/hyMnt
1l8Xi/XETR9noIDhrNYCIpspFb8O8GT0MrEHEdgSn2S4Z91WmsoH7UhB+lAYCy3W
XaDmuFD7C3wgJAg1W7DMQRmuOprnLihxnGlCrAifmvjWUgX3Kd4D+JY0EBjnFRfd
xmzvC/8uHEhB5RfKHdcXBGaZ4YRkmjp6YiM9W6fHxEuNM+wvSPEIX/yJQIxBMgDd
jVLkY3boMzqcQqmq5v9XK0MMl8sQNJ5jQI8Tmn3I8Ub5gNNuva2BN/EhHjeKpO8s
ltVXank7Qvu13r/ep2xCrO6vedpyjnl0AyxWfpzIzWNGM0++WZJhUStFB30Vn2dm
pUT/9II0WpmKKOPrqYM83eZHHu4+3NUBXRbPuSxY8yE+zOpbNu/zFnM9rDSwBOAJ
DRNpjDNNGXNaeK/3DzTu48yvdccmtFCw7Fo6moqG7Z/jlxK5OVFQ4JSEhnVC8yqL
4/I0ijbG5upYov03nYwIa6gUg/9gW+/hHvo/R1J8K82zl/PSPwRdaJQcB5Ke3CfL
dCs3fPRSDjoa4jrNkcJC+Uv10shxKmH/mMHMNfrSa+Vxrh11Wky/Bt7XuWuunj4Y
IpkUaytMWi779wb00FogofDKhe/7OtJ/ruRdvXdu7bpDBFZD146EZaWFxLn5SSVG
skJ7os3osp8AulUAKgXMHsoMJ88pw+6hVdN66wxrJrhSiMFh3eveVaneMRQaVri7
umOQqHlnMO3yfo+2PI8gXkUoJ474I+38uFJhVC/bLi0IaBO8TyaOlKzlHS9OBTOw
4u5O7bLOdM+vd/aG51eyUN/WDRSdxijT5NtYAoesdsxyY+lpT4qxKw0P4FyIhHAc
bizp7f3LBqVVZlndj59T/kJjWw1Sauk1AGzy0cjMmN2zXqArISDKIJ7JWPdIS6va
EKpQFx6Das9So18mDYnnHTuQNdiTOIw9mdVjgjh+TXiZEdz0HdWB0F1h+tGlMxSq
uyDWFa+1zRmkT9hZq8NWWKaD5U+QVmDzW4+a+LJ/dpber7WFnpuJoRGNWfFUB71L
Li0/WL754ggRZOY0CgtqKlPaItiaUa/soXYz/uroXKWgSqL6mRhfSE1VFZ48SJ7/
GbMEecxozfhzz+ORKLGF/ClDZt9e4liHV97KyAp3De7exWLuw3QtwzfojNj7+KVT
heLudarO6dt5QCANvr5WagvnZuePIRMPlfC/Nf1f2ZzC1qwpK3PY4CnIUkfmdrU8
oGBrmHuy1EzcdQ5BSDOJUHmIh4ycokGIsTAc5xJZxx7abqmhZ4Inh/S4qELE8pmn
KPZLBs7xwBsG7bxp+9aRs9QEyHwuqbVI9AoL8NctOplcKZy5PncBiRafwofnLiCU
FJzDpwkVzD8WTV55ZktRzMBcwpydT2dz6PDR8DikJkhJ3c1vuxn/jYXQ13c+Je8a
ds5y2dXHOlp+mOU5R4k5Y2mkDGZFWSOj8WMwXWUFiZFs4VIMEtJnb3puZCFYXZiO
QfyppDKBbh3/4G+B4DAdJNKyvBVK0o0Mb1fcZVkDdaiLC0Damunq+Qp/Sb5pxQcH
Pb5am5ya2TwYRUpELfyWQJZZwqmJv+zU5cCcCo+Xr4vcyMfIeR+8rmt+EQAtdmoL
Ws2vSnfSQcqWYc1zCk3TPvKTJsFIDLs84GcyA/q1DLrZt1FgkLlOjV8/ThYLt4vk
NXkd6FfAWii/I39YunDkavLF2XL0erNAVZ7axfZ1qaUrUXblITD6PGp40ZbWYmR9
q6K2igUrI9kD0ZSCYpYnQnl9nHjPhKL43cyHgHrcJmftpoLL0g0aRhn0LY7dK74I
aq1Ke5a3kkgpPi1SE/criJFZLtna/CHgvdwNwucREiD8IsefHJ42v/2Lyvpchz6U
7DupWUs9Y3LMhfPX9mp6G43hpHr3jdAOvN3cSOhDtZMtb2c9zR8BvMEyeb/71lKJ
7RISLeQReqoQEblsA6w07ma5Jo0bZ+AMu1R4WtICl5Ijoi9vg9gtHrQqZiQ0K0Ls
pby2y/9bZzNtvS0FHEjZpPuD6fj0Zds5tsWZctGaebrkzgUvaXU++vccqV7ZrQqK
ZO1EZkOibhNmAZqinwmHz09HDeSO4QjngQFqagSpWWFxuIECCx8MhnnSfAZu3NSr
Id0zWJ0bntuIdAyumYAadOm/mO1FArklOLDfvQp1bHO7TQ9cNOb3rwTcFRqrBV10
V7/t5wVTg6K1DE/8QtHHMZWZ5/KNjxTnf6iXkGhrHaGZYuxFF5Y/YWs7mthj3B7p
WyJ3U2TVy7b2/TIUtJ8nzEg91IyUu5j+R1+Wf1vtejBO6fGLbL3jfsOzki0NmWGF
J8ppU+QaiNHcq6bacndkLp7sJxHi8AtxxatBeVukXx2LoxxxaPez4Xu123PpVAXT
K1XZ419y9U3JOKXeB1FqiNC+1sJpHR+xcH+gQ23HZYgtyp+oWfDLspxVE+WQJ0e6
DEfRNf0QusOrE6Rp5rd69BNZ54W+jZRzKUJecJnxVVULvOecAJXXZjaSiWKJdtTh
gKyeaG6mVmFyURUjjFSGGkh2EHOEK3x0TOFaGW55WFs1oqdM7F9707KqgTNkHdb9
6Ue5ykDxa09CF+/9iVL3j+qFMmk6TMc1E52q7LdzZPsNzowfJGSzIoRAE00lYf8o
v2cLzTutRk37H1GA6UNe9NyofIQ0N2IveEYkzwvWbMhlZkovPvI4fjnvVck43/I2
YYkEdvlXTMtfLjoLuJ50az7my8MszXo4Ls+GhUkVzy9ZF+WiGOzCY9N5uJV5cknR
TG7uVIFQji8Qch4G9udKugDXvpAqPtG5gJUHUFWSwK4eZS7XMn2JuJfpLthN+9v4
6MVY987lvC0lJKl5FZ1+MlKXND9QSnaWzD2oG4lsuNJWPA/0zPlSSafJEQh6V0sy
/uMJ7my/CPku5geHBpqdgNEFpUoDEss4fvBQJ7kdEEfZrSMpGCCy14J4zOi03UKd
q64ALTwBSrI5c5URCDauJu/m6HHxN5DK9bSV9D5MHF1TA10FfDaFWeAb25p4VyfP
zmWw1A8LcpO/Yy8nWMVZ40xyNDPVhm3++cesVHxxSsoDArMpDwSjmvtAmxhbvxgG
xVtP61QnZKuDH930vpoyCyDt3YHmd0eEGYxWncRK5eZGGF53HEK4nJWSx1abhyqt
Z9HQ5uMRDeztH37m2wLcGZgnvAmuRZJ2A54h4hLUjUFcGwjeQaorSx1mFkprw7rP
3aT5/ykRyxtfzoB5iYFK6JcQ6AgY37we8ak71gUHwS5O7z1dA5O1elAkGPnmf2jJ
0eyhaRpdvlB2fgRsY4VITP5CFrK0ArdD+0q+Sy4Cpto3nD4Gp8DZk1ixeWS/JY9o
bd09EpjL0zDJLBTvulrewadBWjnZIBjJ9D03FlmKDUxRBoJgv5DFugj6VgSOnDag
XbM6wr5hN5idzwzOdzTUIhjz4v3rQ39nHTx1gLEZRFFLuAIW4rUs6Xdxj6Fh8Oft
ml8UKhdQ5XyLYyh9/eSMk3SHkLQrhnNiJc/CX0RDk1917ldpzrlAQVUIq/YeWU+k
9hGYbZUjU1kWwgti8Yu8aO7lpQ1dAoJbDT2u9dMa9Fz0se+qHXyAhrog4A8z7OSW
e8B/M9jwLGUGHTbuBoTLIFKaDyRXXGuywuuVdXOt5himaqmX2qTisys0xid1298W
vhg1+ZzheUfFUIIRlf32uF9j/FwAoq3yhqN6XMgFF+WKQHXmYHJ9cdnhOo2emyIb
q8DLTnGXK1iqelPSRZDZKEUlXctVGiEcyFXGEmu1vE3PZlc314UWaGy4wh0hIO54
DapJTasOwx1tlawcQXOqRC64WVTxo4aoJTZjxx+nwNFFvIv9rdJkVJtRqzrvwnux
hlc0+KksW1fOEAUcibN3DupNPabPgsf5h6BDODU9Ls6C3J/J6+3ke3rIzXGVqGtD
i9H9jEQqjaomiAtMmvim7AVcm5ab77T9x7xuHPY4FDv4VwJcclh4Y6aI5D8d9t/K
MMCnrnoZR9/Fw6Sc9ajcVqwR5qfTaalJh7/nhbqaE1xysPf1d3ofjxyVwo565HBJ
TA8aoyt+0qjEKeH83sb+afwIwsbSHwDUuXIklrDqI/UtEP27wteG4MaveT9stBQK
9yljMRJFFcLt7ahrRR5TU4e+69b7zv28PyFhsbFqNvA6sSvpssFNQNLh3YtzDZw3
gigElPU0g6JZcl8sIzfYO+ajqU2nFJ9PzoMRJ+sDiIPSUv71hUD+c0IwNeT9DMAW
CSbq21Tkb6xEQNor2vm2tD6MlLBubGe6eyldU5cFEK+ZBFY63sdNOHkbGqNZozHd
X/Y5n9vcOmNLkM8Hgu+DjdXWaSJS6lh8dn6MHTo4+zQUq/cTICbiSvadlIqZWwno
qKPQ7kf9RixkqQdC9GZbybTj5KNslIPnJJiGBPAFeRqF/sDOuTmX9SN5Ed2mZBZE
ZV86yGouJ+ErMf/RrgJeZ4JH+VznlJzhN5gD1SuVwrgw3OO9AylhMlhdnnUbk9JS
Bl2oTig3sdtnTOPQsPiwjsTRjU/poOUR2woQwmdnPFgdIj+1z7owVvjW5KqSQszB
LqtcM/RMKhC1r/AC7AKel0FtaZS78Lwuj5LFwISuLvE2o/nycDwjVCBtl7A5oSWv
04eIRpqFqIOg2U82Q9ASdF4N2eu7fVF1B8AlzHyRgSZ1iZHogH72oJICrhRV+5uz
+vOIEQ66NT3hjDhhp8rZqAE3HjIUnUX/VmQHO2bHnIJNsaOSC0dBTIE+tTQZpO2E
eEvyE58lQycQKqJdoDaCHv5LAjLIb4VrbAvq6bG5qvZ7DQa4XuI63fn5aVw4j/Hm
6GIFyj3kQgHJJLbMR4HI9pXLVmwPIZ/Wzn3KgWHo6V6Ipcdz8+SI2bPsrLVdXj6E
R4smp73SAuRzlFCoN2gvpPdzPGBfvEjMY2AnyoWh0H9b4B4STo3HF7ptKj/LFFoK
JizLbRAyErb/UYIch3NDdf99AqrQaBRc7IjBa05aDHRL2c6ggtvr83MZxCjR0Z17
elMJIQMtHkLiAnDe4BBGVVJ3Ly21XdgymeI/JWLbDHfQin76SHCN+O7oD3DwCDzn
jbzz0rwWyRvFq01G8GEnMgK5/kXor5VvrD0dxziWBiVnK+Qa7GujcNcUEyEmfWQH
VDlRjjALksLB5wLihcvM/HHJ8lFcOLfMSY/noCPWrqw69cspuTBMCxkPyEk9wpV0
HYnLNz8L7PCPXhmgaaRZop/8ap/PU3wih/jnSJx/OdcWtyLAN+2/dbgjNbP7vuKd
SddYCNlYkG05+mydjzCbMqLGiQCBXQrMon2lwLSWE74XJiVHGim/CAmZeReCYltv
dig2PS3XUhKCaHgb+IJ9A4LEqhEqABYG1eVUUJbmTRtBG7/vm02uSJ/0b0tfcAKG
tyb5tWPD+V/fGrgL7LmO1HHDOnkOe9kbwCRz/Sjm8aClAwajX3kQZlmuw8j1Vhmx
um9mNkUPGmdUoBklKhWZBNbkkzKgWMY2NgsQQxxC3MDCUXyHT7BeVAXLPRvlnQ3H
iUmVyuA1t6A9TK86iOF9cqWkRs0VNnuPpHyFueByRQij8Ovq3wGuGbhBVHbjhm1a
BBxacxzHm7g6QAVckiBElGREvCqZ5QAKqJodTvDAuTRhHYbT5X/5zXfkuEkibNLL
6pM5C3FZIc99dRXc7pVWa6uxbPejMU6AcidzrB9FUt9Q9yv/8ujxux2Wm1vpxm/u
JJ3ZLL3jXuVUvHaKfWuZITlTzxrFGaiCCgmS9xFAijj7Gcv0+XfO8XksIAHr22ja
SI/0//Z7tk8LPE58VTZNdrBbfngErN0i0hotBywAIgtr6qoPy8VvuyGb7N99yJqB
CmLeVVVm/2z27jjh5HJszSDWfSvvQOJ/ikHM6o47DuR/vDwBpfHsgSO9iQ6rah9Z
L63zxpzFNQ3eivJmChaVmHHckh271D1GTb4OBFQ+fnZyeTUbYiSOWP5BZqK05vsw
ItzYa6IT7qsFHKvuY26AruWpMjTkZ3xFjsTmc0q+quCnHC0Dg2z15IXsl3Rlg44t
mCgDE+4K0ZeOXsYMWM+ggzfYONgYKCv8XMsQ+L3a9SK7NN3wDE7imtgwRngnV4h6
ljHVCXegr/gJ1p3kXYU6MWrfF0s3BR0I7LLUGSnXBmJvgEZjADxXnUrNGkuZzHvE
F7BmF1gFuzf0VD7p+9cn/NFFBFCf2F4yXbmpBK4LuhkiPCgXiIqXejHkcycacwGV
Y5iVq+pVsBCapYjyO0SrnCTmz57YMSOARpiZDMFX4VLmLp70SPpH0etjF2rryMLe
prfHal/NVA4cVPpvuvB9AXsmOrpOIpMohnKIvsLnisyZD7m3uxxRrSAbwrv/aTl5
AufcaRIQSporjVA0bPWzMr2y+RWKj4ZcP6vxau9VZUFnqXs6SyCnozF6sYf2HFos
lw2ygeitnRhvsHCR8cuKQ0NAqQUmQwhPaJcQF9j1VxvKqEWgstDut2tfuwCWJFTS
UsD6dhUw4fKkbzjkqXAM2oNtf7QBTipON5A6vRVPbV+lr1tH6ALzJ4TP2se5OaL5
Ug5h8Sna70NSybt2hGugZLcXYBIwggYbug3GlM5j7CagDrGZ9hfOFYOHYCnPTwkn
H72J0h0ou0LM8UKey00umTXdT9GaNdSFidFo6yqTZhNkY6tvQnr/EK38A23JlTzC
FNktau3ysf8sHEd1wR/4UlSCOcpJ4r2kMYGg3wBfb93CcPfWLgiF8dXGoWOMLgGs
d3FO6+loYREQw2tWt+cjAOE3e4oCAxphoIHziv6CwjaajyJFvfH8uePQuX+bkRbH
r5BUVla28Amjv4w+mZr5VWcCHB6boIiTw2UEARenHmyPcBGi0rvhOmdEtp+jieIT
sNgcl1loEZ7DNrohhzxmos6lLN9Yipo0S2UfDTes6OzEJErqY0Dz/0fFKnGFl0GV
UkjopGTAK37wz3JDFtcas0BM1v+Y53ESufZM/SHwcN8ahdCAJJgQvJM3do90nt+1
eZDVbJmqSbG3/r7bv7dhLnTvS3+0YnSa7YQ/yFdIoIVW3pmDhLTbGsN/pJSdS8kM
tOK8woMVzwWe5AuMsmQ9wCpX2aMYNZ2qtBuBOC9NsTEEdTXLxXHF8RUjb2VoB2yq
KFEjO9I7RFORkO6Xf1edo0U+3D45WlpkKbEFIOBFLqQ0EfVeCoocKP4eKq4feYGU
mUGgaE4polYIR0tA6V1kp3GZtWYofWVx48Y8tuWXaZ7H5kvBWcwfvAm6hLVlrXGR
uLjxnbX03IbSIoW3/g8aoYh4QXOgJVcgn+6NWvXE3GANvwnaIAlP6YDWbPJ7Yvy6
NiAqsg9kjKAGw++0Bru+mXjAFe53xcYp8zfl3z/6uvf+o7QHpKSPh8OY+P5/7Sou
Ajcg/HBcCPxwXzFU1LrpOwsoFazr8aRmd9ZZzwIPlSUogEECj7N6Of/nkYvwQjiq
WYsize83SGkmtYe4nksgMQSButYB5LkPUzrSLeeLLtqk0AVdQ5F9N5lIgi/OerdG
AdTPJXiUrco9Ig+VRlzKq8X2CredgX+58rwHzK9d2lFlP565pRFUYXVlWFQaWhiF
g8hWXQBkN7SQQjfHzs1FEanzQUtjKjgz/mFmYtJksTFzjPO23ViyIqjZsE2j8tdS
MpgluJcIo2wWsl8cVkyNScBDTonHmyaHnRDGng52utECCE7YdQYvURq45QuVZ+n8
RzmIHx6zX2nkdbH5aYx/uE5TbsxY1xofRiQoHlXW1qAbcFUnjwkfckZ1KixCqW7S
kB6m/s6Fetu4fsuBs/vbwphuJvW+/veItGva2tbwcjAUDyyKoXHzU8i//L2S4feA
88jhvqw/dQUWe2OmpK2dHH6rMEcA15QC8FR7PnMI2loqjNC7RH1ulV7la1f1Gh86
wJGiCRkztJ2zEwZN9W407rK8HsvBP0BAFe5Ijm86qnzIsBiB7FTXiAh9i4ClWCTH
+W4fIxuPW+5b5TRhvMS69VlcUl1nKeGnlGlsFCkaGoRj61Jj+00heQw0RLx5SMdk
qWwiYGitPtZaSlgewt1CRY9kHB3w2oiriSH36OLAVWn70/0CTccnzd56I06Ty8Hg
Jmc5pRZ+FdRBgOjvE0NkxqSnB4NSuj6SFFFOYYWMzidEVmbmMrsgoBXJfRTo2J26
u+lFveFfjrH8cXAbvTt06X8neg8z9ZQztwBQmfRjQB2W/gyeP9EzRXYd66Of/fEq
Hfj0Oou/nsyuITyI13h8AXvkgFz2TTABVC6zOI3eP9JVUgBcl07BQWNhCdt3fAPk
cakCymU4hwoI9MQNxeZZNQB1iWQ/kOctJ7Xy7lZr0d1MuFbSUrjDfNo0CZmWQ/jW
enUwFpdtSfriWiXVTRfqgoccjWI1kgNuThql0/Sm0NL0UZfntR0qj8XIrxDvYfwZ
AtrPrOYfHnpi7/s33zk1zcsNT/kHcgWINgmzvaIwoQHvAVSE/GUXr0wPEWHGl8hg
gyKv0g1J7Pql/h5WfaC2j+ePEac5cM3aoMpor1dl6EJIE0iaqxl2jnPqSddBqeZH
cNA+kUK7eFSwDZ67aZUaSsOGw5hdulXL0s2FBees8d6gfXdXOKjYq7Rw2hsRNWlj
h1suingt9713XKPjlMPJY7TbvTuGQ8RMQQFNho9jHsB9dEH5h97AV0F1Wngxxunm
SGqQJNA6toviAjtmPECyIL/VlIHc6K4joLRXB6sOydS5HsmPZwvxoYZdcFbetA0V
9PiynNWWNyuvQ8AniLIoYDR6exDIWWLrbaAlodJDyiGBeSHmBBSiik6WDrFW52Dl
npYUvUDtL2iy/GhqgJMI4KzWUTkZ7rnlHktpR8lv8TdBwtkgQEaMPKOzDeAPxXJb
3u0G2niimyEYM0ua2EhVERwk41GfgMVnd+o8fvVP7sMC4/d/zFI8Rw6dKbvbumD+
YVJxMVaJG0FJZfsENhxXMmEWkyva/vo1E0P6ZoIVDcuqX754wuSTW6HSgRCJ6MwH
ipBRmoQI9JMV9E3ZpuWe7vxZYh0y8qmUZFZ5QSkdu85TN6HAJ5vKpiNIMCB9n5jA
8Tg2gn4yi0CgC8ijKJIk+sB1PboHw5XUT9tG9cWuRr8puZM0Qa7gAPOnBN/i/hEp
0NdRz/wTa32SrbJDcCmsqbBn2ISFtxUvUNpNxF1LT7J6Zjai3VL5XlD9gHsLGd1M
DTthiXfmP2qiK8t13rZMACjK10n11HSyWGwmISniS08KCefij7dF9kZJ5um1LcJT
bye9anU1gDcrnUHtIkJE86+l1UtaORCCq512WN+erI5T2zr6/cTMf40FDhRpnPkn
fpP+QjSbXdu5Icls3pYtVpb3vqA2xLBCeFTU4Bo5e2996X1HJO22loc4ILCRKhvK
RLepUVil8i8blbnyls3ff5bcPkapWouX1VY/SF/9pIB3pdLMpRZLS962VSB5UcjS
2zmGKvkQILWNKMrmv39NQZbYcI5bgLCQqKlxT/S8yK4jNThUU/8CiqLdxrXBPLKr
r1lzYPLPqeELUjcjgFH9UUFMgCw00OBYzIii7WK0j3OZeR5Q9XWA6476XgTreApT
/m/qIgP9tUm9wQIYfvXaYRiP8W8Bu6fh1D9ihRjzTKk64EPmfPGQvXbDONapvw7d
zlFcInOdIdeLtlByoeqBwcKImb9hmH8S+xTqmTi3f/JYNlKCrfGOXDsPmTEibduB
uR6M4Eo7JLzLFieQiKGFFlZDloxVlm7NbcugPMjPBnymsgV0RmtfGQ+47l4Bmnqr
jcxMNb+QhzlyeLDsmTGkiYaTYMLr4sO6u/v6hfYVccVQpCoElkw/bk31gZes8eFl
j9aFyaFQ7sN2ruhRzlTVswc2G+aJQuUACbk5pPwjk4qIfGjAiVOi+TNzBefPufP/
Tkb0Eb7lhnkryInuzoNuAOzZKlpSTEm6QP93iKUi7iJ6K7c/M/jr5GqX4hKVekk0
SWwChdIgnaj7cQ09yxebrWm3e5AhVddmHRD02Q+QuJFod5N5yvG7+g6T5CBBdzNz
fLxi6YR1uywYM1YYMM2d1/b8kgsK9yjl5Iv3gqYIXmJG6z5QiSkY2CdWbXin84CL
P7GVpFDUy5B21Zg5HJcIr9MDc2g1vSWqcDo0eR7Dvz0L/zg4Lu1wvD30eBsKq0Os
p/8jycJP46EqeRFrI32rF9XmLmZiuNb4G/WiKa5OJQxgCGTdNi45fCNioAmnxZz6
w8ZDdsDn99E+7MNJ96zEQ6wCKRR+RAvUHOiQi9VnOAOxs37U3C8mhimASkoaA5mn
AW/0r5zNX78s84LBmqqlhwdEK2u68Ta9+4Zc6FdyrAp0UqRG3p1HtEaWYO6kQxsG
my01j1VT1/iOlcKt9gmLJYear55of5SQuePmm0U/J5zN067q02lwHaftNNZliIaB
3nRZI1/0aZqJhBfarxMqxEOLMp1ci4ZZEoahdZg+W1CZyOAqx6OnSU2Yy8e8ZTJR
UtTed6OcuQ/cU23UOaZOhW27P2XJOdDf93TQdwfYM3pareeING7g4TXKAcPb1ayi
ZLz7/Pc90gmbMGzGLq1TQt6iyLaKG7K1tICXWU4zfQyaNV2KEUJlX3JTsIBBo9hY
bRvoju1kZjw63MS5u2m4+emxdZ8iwMmkNWS6pVs6YEaXE1RwQbPu6hYxFZhiio83
OEaOs4eg5GNjRs9b4K7BLaY4oxYi17Hf7RQQgEePz0ThAZmKhxJbAHM6uuSi+hep
AwgmQsUKgt7I/8OVgtEapxWGiYiTWtjHPus2MKzW4qiRdPC0hDNHKcxOkRg1JlfY
r6tNeB4PjTYoeor8jrKrVaioHjl2NR+nOSu17kjdWdt686HhAFlEv095+kHIpeH4
UXD+i5Uw93AeVMPetxJfEPGq5Ja0ivD5YMApAppSGMpt0QUfcIFleIN409RfZQgN
`pragma protect end_protected
