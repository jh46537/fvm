��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��x� �u J䇰`#����������T�jCQ�g���uV%�+�@��m���v�V[����̍�HF��a�h%��PA�1(���J�ȍ֏��*��<��2m���\L��f�'e�B3���YrW+��oa������Pg'��CK"k�1��c��R���
��͇b�����k����l���h�|��6	�D=���]K\����u�q�v����IW�Θ-.�F��*\,����X�o{j�:e��ϖ�"�wb��x.~���~��@
��ꦱ�7$��x�4�EP�AO�~�Gn�,~�qv�w?��Dˁ��?�7�wer3���Vo\)m�L00�xmC�r`�� �J����a\>������ݣ`? ��hO6C�`Z�L��bɽ�$�H�r�cA�vt��:���I������ǶH�M�S9�&�qr�q��z ��0X��87n_�UL<���%z;"�����Y,1������\��-;b�^���������e|r�b�s��S�3b��5%q�o��;,Q�(�k!m%�:�o��N7�Vf1���� ���6��W����oc��$v-3�M>������s�b�X���)������=�Q�=;��b�-7$&�=9t�����s�O�/BAF�a���hw�E�j),҇����ӊ3�?ݖv�H���z�r�u�]��Z� �{]�H&�+���o�Y� V��VE�D�/��A�M�P	�|ɍ�Lޖ{��J�Z��B��h��1�#~�,8�6�<���R;B>�ً~��V��6����)1��I�W���6�S�\[��A����W)�>�� ^������|r<C�'�E��/T߈��α���I����J��v��.t@$<�5
�=�S�1c�.�`�ZT�h����J3�I��bv�Z4��[����.�,��s��	��}M��}j.������!��h���o�k^>
GsNPvn'�_
'd�\�Q�������Z ˍ��\=Ӕ��JhS�� ��̂��[�4�DM�G=/d��$�,%@]��đ��1/��NV-��8V,ī�F�y�� K��ζ�n�κ2{�)�j?D/�$�J&�7#I�iovC�EC�F\�j�D��j��PCR���9��F����'��!�p7������N:;@�*A�Y��L��_W�e�RPKC�b���|5���$���~ӎ��\K�r8р$"�Y�;��mF�C�z�)��ۍ�H����k�νR�(Жg�j�a��
�Ol�|��Pӊ����\n �h �B^IH�`��Φr��-���P�(��9\gc�z�R�t��A`���lHFn�4�d�1�~�njT�$fQ�>@�(����$Ș�S���R��x�^�~��C�i��3�F��p�ܯ�G��	��Ju��ܑ�r͑���k�R�j7A�^S(M�e�h������^���B�x������:�_m{�}�Sԣ��K��"�9E��Ǧ~pD�f�!�;�ru\�6 �KLMF��{7�T�Β�����:�zL���k��_E=��Q^y�����鸞!�\����UWk��UJ�P� ���4/�JEV[�>�a�O�ԨV�{fD4�<V�������폤���5�%}����V�:�t"Ǝ�h#����I@���j�K�D�~9}ڗ}Y��Ċ����S��-��!H��-R�%��7yQ��1�X�%�)���\�Jjꅭq�����`�D������)��wr���.�_� ~Z����ױ��J�@kF=�S�t����K�ڣ�{�}����U��֭���>CV�g�O�&�i��3�y֧��v�N	�փ���U��{��d}he�0D�3��%��;t�����Oy$<�[n�u��؍��NH哽H0m}�l"��8f��K%�#!�ka�h�v\�[�[��P�?s�f�d}�& ��4�p���2��Z�i#7�tYW�̙�\c��v���{��o/T�� ��-�p���{}�
��@{3h۔7 #����,��� 1/�z�ƅ0kߖ27�r���z5�0>�P�[�-V:?U��;�N3��f/�!�R�c�m��!�^!��dӺ���Z�1����f�����p�۪CL�kYD[�����(4�o-ڄr���ѱ|��m�n��|�e�����g��b�D�'J�������k+W�