��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�'�I����-���p��7��g.<���K�K"9t�@���l�m�]5v{a`�6��'Ґe� ��ƻ����Z��ՃZHۗ��z�Z�5��U,�=��n�1�?�'��B~��sh�4�,17�CԤC���!S�&M5�(5U�VS"��qZ0��������)(�X#~x��,�25��-����Y��||�󦱤#YjmK��k�=��p�xG��%��Lᷠ����\O��~&�פ� �V��
5�z�KP������7k'�ޔ�k{/Ѕl�B���=���F���l�0�y	ŀ�V���&� ��F7��﹌g��N��]�\�EC�ࡾ�`��8��\)cDL ���-.b���QH��{�=��h��;����F���>U�)��p�󩹲^ג�7��HtR!�#lv=4��<�昷����j'�Ɉ�S.8A�6A��(�����k�_zͫ*g~�Uk���.��<���KWp<����Q�b�Ƿ�`Q�E#/��
>3�ϖ���� �o��k(`�v�c��pp�2.A��Fs�\��8�s�Du(1� `�z�8hZ
@��D�d��?b�]��L��4����X����h;'����!^>�<~)ĥ���4�@]���?�H�������:%�*��F�:f]5�bF�3�f���NGrT	��6�I�{�'̬F�~0�}�������&Zc�K5`�W��/&�A%ʳԭkkd�2n�Qd=�Z��ť�w����"��/䔱�T�m�T�1����N��2s�q\}R	f�Q"A��C��YP���୳�J$*,Dc�V~�r���8M)Y���Y�g"���<9�ό���1�-�R'T��}���Q�2�AsldP������[�Φ�t)�G����Պ ��㟋h��R��\�ڛ�_l�4�.uG���B`��r����^�y���5�@Lz�޷�-T���"�ç8+��YV�����C�:9;n�E��|�@�y
N��^������7s�Ɖ�����?��H£�Q��q��%�hQ�����v���*J�U���Q�;tۊ\Ñ����nb���	B��
�;Vg6M�eGۈ	�l�F��xd)��RA�O�,��q�g�Sa��x��+uҖ�*c�҄�ykU�[Ґ��so��ܷE|�!��9O��֍��Ҵ|����p��Wu����������qag2��˩Z�U��}�{��;6.�s%��sM�%�#�t�iV���O�N��sLֆE�(�'��Ϣ&Un���͵=������~v'x"M��g*s�E@PN�o�W@��y�P$:�.A���^`#j]-�rtG��8�>���E���PVwC����DJ�cF����[�����N���)�''fy��vw�W���[!Ovо<��?�U���ðѿ�eb)y��&e�t�v�} �h����բ���ްX�[�dD���/FF$䟋)����1�A�*�F�)OH�hӶ�&ܙ�Bw��'b�+q+����g]gI�?>�G�Y(�B?���%��+,,��ԸF��)��-27�^������Fn��g��%��ڐp:��݇�'Xe0<�P� �w"e`��ع�G��(U�neL�ۛ%k�{�����S�`�I{���#p.1/�kǬ`C��Y�d'�J����ϑ�Ą)���^����&_�B�K�|����k�=d9�F���\����������8ֳ��]���_>�W�<#��Ha1	;��PT���� {�.�w�I*�P�ꏗ�t�j���45p��R��'��1w����f\��c�uJ���?�T�����*b�l�#t�����Z%�|��rQnKy$����	@p�f�h��~:�Ɣ,�0���e��rK>�˱���ʭv��84�ԁm=�� b������9�8wj��ʉ�j�oݧ"f�>�>���WWYJ:up/C9�Z/����݊��{1��w鼖�yMeI��`��q�� ��so��ǝ��7P�i��r%�TM��ʝ�j_���)���� 8(Y�F���/�TR��� Z��x���S�zu�L3�v�M.�ٮ6ts'�# ��!��D�\MM@.g��}�)�rZU~I(�/�"h g�����)7��8zӳ�i�xz[ ���5Z�͸����m�b7���7�wz��$����u��?�@�c�*e91���-��mO�QlAp�m0R|!�w�QR��^�Q�i� �L
�{���vQl�#x�`M�o<�j++W|@ݍ��i{=]�c2�{fGA�M�7�5�}�*�n�6�����D�)y��;l���Fb������M���0���'�\@]��|:��+�Ȇ4�����f��s��4�f��M�ѩ��$���tuCbY�𯨴����2�5j\)�ij���ĞAن��	����1>�`;e&��&fr����f�.�Ӷ82����/�Y��n��6� ����U��s�~B���3M�&�!<�L}������Sr�C8�C��'!V�cfP(���,1�>tZ܌
Z��-�ǽ�Qr|��L�^A8P��ݫX��R�o)�+���N^]b�v\ĕ������l\��S+��N@\�_���pڄ��r_}N���a���Z>X6c�b7��ϼ�H�1Ł�U���0.�,��=Ղѣ���|)�ݝ���oQ���{������L;��H/�Юgp2=
�L���P3d�x��ݍ�`�����3�\���-)P�n!��1�O�ɝ���ԳE������ډc�5�P�GۀO�!׏n��
qq\�2�n�%x�s���P�-�R*��6�Ȱl�l��P��Ц���PVk�:�!m_��u�-��u������G0T��+�P�9����R���6굗瘱X�#�D�JYY��ߊ�$�e�1;�^�0��n!��ev�j�R!�q����j��7dR'����+�}ԛ�3O�.��jAn(�{t�\:�&$s�g�KZ�]�6�Hy�X�\�޾�AaψΠiG2θᙪ|��}���x*C�Փ��uد)�i���S.��j�h��)-��;�`�D����Ԣ[�@��mu��f�A��z	`.i���3�f����q���i'g�R�ɷ��Z �= ��P�BcT��WEr�#bG�	�4����}��� �[���Qgb���z9��"�`��UIV���&x)�A"��M�U�L�U���v߷lRH��L<Ef%����[���,4 6�S�"X�)���.⌽�}o�#p"��-��i�n�,�q�w6A�К���q��ؒ1�sc�R�(���-��]���#���o����O���V���R�F�I����,��^�'��7f��?$��NR:�4��ɓ�~y�*��n�N�`N%��������U�+cB=N���!�'�U٦��t����ƪ������Z�#HԒ�4�Pp��6+�Jxk)����F9���T���D˵e�����26h(-�	�+�0L465���4�?
��ǍX8 �q��V���n>'C�0{�QN�kF��N�	��M[�@6e�4��N�z��6��Q�����Չ�s1�7ç�h��$}����<��/�n~ZMÎ<[Q布�$�=��U��#���;��6�RP��ߥ1ƽ�x��!���xPm�5� �i}�[������u���&f- !PUh�GgO2�'���O��B$��,m]�n�Cas,��O$��D�A\�sI$H�,�Q�f�4X�81�=���xR�R]�2m�@&}�"�����+\P�j��"���%&�Š{��h/�=EkIA�������x�a�(�S�(٩�jNҕ���]٥²{���H��`&N���;kh�����h�Y���ލ$�3�R�6�	v��a��f(禕�k�]3uc{&��gG[�����O��)�B��#�s+�WB2��F C(S\���l��}jGM@N�s�:ս�Q�Z3�X��y���B���������#�g���a��45�Z�r����6zwU�V�pk���F��Όʒ��
�آ\�H��/��+����Y6�rH���k��y�'�$�??�k���S/(1�Cཝ�_���뀓�H����!J�x%�i���B�Q�ke�OiП�<�)��yiIq�V�m��.Dl��2�[��$i9�k�����%������&�iW�W�;\��-��W*y::T#KP�jd�@�����	�
k=t&���m�GՏ�s��5mZu�?������k�D~B�_A̈́����U�i6���
�/m����h�����G��A|Ȟ��Ι'�x܃�8Do�m�(�)���MDټ	��m~��Nm2{S�P,�M��O��&��-~8�X!�#�|4��K��"�j�J�A��{襖c�(X�=RZi���i���M)_I���#]�MLx}U�
tU�_
y�9��M>֫��4��YQ�*eBk��jņ|��	j���Q;G�m��4e�k�)U�I��sۋ�|���K�4�%g��٢�%��(����F�p���#+*�����~�ߢEL��<�4k�f������w5_��m�� �j��z�C]]l[HM�Νϊ��&�aU�n�*'2�����w���r�G��c$z�����>��d<5�nOڢ��gY�~p�L��+�=�5Y4��e��8	(�3	�����y'��T�����ǅM	����yV^),�s���]p��7J=s^������gƁ|�����!���
@�Ռ����=	FHG�p�)��r��J�o��-��!��bML찶�)��hp��u+�?o����$������"WJB��B�|�����%P�L�05����H��3���1���?�(��[e[��B\�I��;�Tap?�4���0��x^�&�����:���u��C�(���?5 *���bqc���o�ÏT��a�י}���2�Ce�us0�@~��ai�^,l�j��^����n�
~�CB�G��˗۰B��45b��WS1aJ���-��ك�"�-�y��Z-ZCr��飛���G ��t�QB��uoϒY�U��d����N?�Έf�>"�Ȏ]�b$���<-ҵ��dc<���LM�g�!���ݶ��6�=y�Gb�7T�^�4d�-S-G9�n�z�d�����Y�k~����*�#e������W�J���ʜ��<�A�����C����@-M��b F���<xPk���pޒ2-I�ee�E��UI�`���8!���f�gRZ�F�2��T'�m���_�O�<x>���-����7҆�xG���@Fx��\��j�B]0Q��u�O1 �E��R�Gr!Ъ��5�At����_���@���Ic���Q�Z���<Ys��R/��P�g6sm9�J�� �Z^�cڇ�tO��N����ՑQj'Je�1�\�kigQ�O�nf@�b�\��ѫr}80M��ݩ�LU�Ĉ�*-@�� ^��(�|8|�^oQ�"��J�;t��}�ac9SC5Q.��/=4g%�d3y�N����]�,*L�8Hw3�*�r1jT%a=�W���1�zx�V�=[�K�7wH��7��gjD�� Y��8s����z�D���1��`b��vv�M�b� 8����B�&?Eb1�ɢ����ǣ�����"nsL'�M:�*w��v�9���}-����{>��4uߊ�J�_H�Ye?�}���d0�f�,7�`b���!���'ԫ�e�w��P�a�L&O&b�����Ӑ���иz��\���5����,��Y���,"���lVK�7�`�q�0,x��;y?�3X������Y�F�Y�7��BY�Q�����O��Zbܟr%�P6�0���i�ѝE7)�8�����j"7�ٲ'7��4��?������:����0[-�im
n��ȵ/�C�:�i
c�,�3D(nCs�̏��PZ	�����2ܱ0z=nS;��D��
x��I_�̟���~?q���F$����U���ku4UB��lO~l3��t��#K��7)-9�m����">��g��\E3��/�C+6'�/R�#�Ø��O��h7&�D���M���N�I��A�;����D2�Td&]KZ^$�y
��z1����խ��^g�bg�Y��~F-���V��.�"�Y{/a6���(�ؠ)d|dW,���Q�fQ�S��J1@��J�7�
c�ܲ�� "I���G�?
:��o�al����q��`d��TU+���kز:�lz��!�����	� �WW���4�E����2xXBAGE�go� ��A4LH?�d�#0RH��1-O��N��@UH�� ��9v��y%*����='�Z� h�Ø�-��_s1��!̓��n��B��c�}��t����ԠEH�b�T����{H��o�i�G��ز��>R�<�P���k����!
����	˹�-r��q�c8���]�T���c�\2����'��U?�̜Y>���\Ӛ��?چ���[3�
�8D�a��xЍԓ�>
�!/λt%ځ"�4�ϫ�jOh��3K�ؖ��v���vZ�ԩ��^�Yn�o"g�Ԭ�YfG��y�PeX�'��XKƗAE�߆ҋ>/&8�*e�����a�������n�q7���N*m���-���n�~�S�y���A]^CM�Ȧ����A�2�7|,�	�50��A �ѡk,%i��Y<�Jv��p��aL�����?;�	\&'��A�ƞk}q�먕b�D�n��]�Л	H����.)~�� m�`0�\�>`�Y{i�C5zL��{��sO=nEf$:���3c�H��'p�����N܊Sq����I�̭���w��,��y�������=m;�X�=�(����G_��m�9��*�|���e�r;�I5Pu�6�N��jd�b����\��\VݰE�z�
3�O>������e�7{B�cM�Y�����Q<Y/��pE���F�Z$r�3z]e*\�^�;��[>��ܨ��G���w��r���i�������2�fd�=��	�v�AR��s��V���M��5�[�!.S�+��kB����5�$#Na��ѝ�� ����휾�0�P:�Q+��)r�s�S��L���{��f�AC�ɽ镦���Y:I?��S/�A�c#	[.D�K���Qg�&J8酰�q
H�-�a^���W�Y�*�L�g/O�K�WH* ����Ye/sM��+ �7�ߣ/�<d;t��x9��I\�����&�����r�rN��"��g#��$�Y�'��)l2f���I ��0jo`��G�bǰyL����Gt�9��L�iY���2�!������|bSs��K=5-ej'q�n��r��0�,�O�[Uf	v�]�I� E�G�s���&�5&+��RY�2�����5��9�cɴY�	!��Q��̝��oU�K�t���6z�>�962ڋ�Ъ�wtA����^����S�`V���X���KE7�Kؓ�ع�K3��v�=U1v��V.�+�R�m0�C��V�4+8v~B������!����t��������'�m�t��[R� *C> .Z����Q��:75:��לI뽌1�6�)3<�)��^��g`��w$ϳ�'QWc���md�L����r(�-��8��x��Cy����)4�M*oh |[C�e��(���K�RU��+�2=5:%�A���d���q�){U�����P�|%�b��VK�1�B�?�*�'|8 ���	E5��<�g���`���\�2Fx-mG�����ؕ��r��bb5l�uS =�e��f+�@�XL@��K�����sp^^rS���h�N�J�7���x�'t�5�s������Qa��t0����5Q�Y4iXx��Sǿl0�{Y������!
�V�7[8��^�.ù�qa��7H��E{��V�u����)�R��JT�c��p�ʙ�6nN�]H��\-:A��4�<oZm���AA��Y��Wݳ�9�����=k��J��2D�nń��TT-�5�\�����#��yp�,�l�j�I�{*u��cf�2�g�8�	�&�<�.���g�8F���}N��
�m>F4���:�ݵ&2q��X�����WC����
��X\�!M����*B�����Rg�[<߶��fW>�h�+�d���d�)k@6�A���v���s�)T?�;�����[��ֻ���"X��V<nQ��T̪�u4�"Z�}���.�g}�k����='_Q��څv-��ӜXM�P����i^-s�U�Sx�⁢�%�a�,ӭ�D��6��y'�@JӃ��t��h
WY�YO�]��EW:M�L�n�y��u�Z�=|t� �\����V�݂�[*(���{��v�b�l�*���t���!�B��oִ�gb���`�O���`-U֦������ے�^WG�Bn�K���y��rC���Tk� ������#9=3�G4�~Y�٥� ��$�֒Ny�ڠ�.m�M�,��y'%lF�5Q&f������)l�t?_���:���w���4&'�x�*A� M��g����`�ը��)��D c���*�,F7h�!W�/
/\�s�,���A����М��娑4�5�}FkԜq����7��m�Q�4�+
�Q��{`����G�"i�v��};������kxS�q�ɀ*P7�4,ݘ�-��-���me5*�%����zg�R�G4��o�1���d2y�4kb���i�
�`\J�2�y�%Z�r	j�ZD95�Г_�Y*�|�c"K��¨�y�2`��f��5��+��4p:8�W�������d�$#F
��Y�PmE�K�aHa��7l� 	!�9�|��5�P��\tn|q�b�iWF���=o�3�*CC���n� a�JO��Ԉ����)V�ɱЂ���̻��dV������D'��f����aO)��υ�RA�}�c�
}��9�����<��+�1_�`s+`�L����F���/?��@\������?0��F}q�$l����x��E����� �W���-�{𧖟$��5$�N�?�ij3������8��H�ū����C����M0��b�9�i�2����k����<���}�s��d',���t<����HߖP��bT}�y�O気�To�~|;��*z��xၧ�[�P,1�?ҽ[4�/ "���N����L0�e�ѡ��LH�I�h,"�V_�X�v1d:o�/c��)�ܞ��<	
��Z˱�}�A�X�Ћ���^��W̬�O4æ��E*��	Q඼1%l��ʟ�/(���;\騎�5�,�#�%`���̠Ĩ7<��ODpp)A0���f�{�`�GPi��@�M�}�s�����q� cz�0�4L�{;���
 ��M�}����9�����O$V���.|ᕇa��Z5i�f���B?�����$�Y�=�.Ƒ ���:hй��j����l)�E(bz$w��r�X��d�w��r��cק@6=��J?��0�G�+(�&�+��1��N�Or#�"��MK��kR:f��luIB�Zu_!���1*��0�p�(9��2e@<9]�#J���XBcE�[m�
p;b*���S�C��$�4M��P�W*2<I���h������T���/
�
i
��\���G���{�>`�0�i�vh\�FP�Y�?[��*�/�1W��L��Y�d���)�����y��aLѧ^]2x�v$бi����5B���q<��}�M�ה	]?([=l��ɱ=���f.��9�>����v��
d6
�D6CK��7nM�y)m��$o�
S(�pCT�P�y@:�/IŅ<�D�.22u11���V-Mڪy&��U9�m�9��[K�Wm�x��|�	�!ڏ�ΩP���@d�V[�z���D�z"�l�J
��OR`�N��Pa�'���`2<I��׋C%[��m/t#�Ic]�Ǜb��l�j���O��ڒX�H#�}�s�Q��n�Zk/�,���T��`��é\ɚl��I�N���!�7�2^`&��Y��[�y�!��Ws[�"��'����hm�Yr��[e��ʋ�ݵ`�RѸ���I=�*�;����I(	)������zg�{F����R��V�||����6N 0$:�����Ю��B8+FM	3��1��A��K��d;�9��L��σ�O��:z���j�,%�V�?Cv ���A����3G��<�WP?c��yX�F
Zq�SJ������)A��.؀Kpð�$��O����z��1�P���3��f�K�t�>��}"U��Fx� �#j�f���Rf�sᡇ�y�̸������=?���w�]��e�$\U��_�k!��:D��ݽt�5�o�x�&�΋�4ɑlUQ�[<�����bc�~�}эѸ2��*mO��Rێӊi����G���q�~G�<�x���j4��g!� @>ȋ�,E\"]:q���ibü�̓������^c��pG��f^�*E[�LB�F�r]G|]uη��2�ɹ*:���JZ*���LAMgd�����*Y�W�H���G��Z�����" �l�U H��,����@��j7�%��#����[�t�?��D$�M��R��kZ�����r���S���{���H����vcbtE���m0����Q# �ز`��o�9�"�Lm��<n)��5�	*� ���ɩ�cz�f���z�[�a/�2�a�4A*���L� �|�F�39��`H��Xs����g��8ĞiWÔi|���?���R���S�j�.�JM���F��{wk5�VO��}aSS�I�o,_�z�B�U�%=����1�5��V�.��**L������vp���,���ZZ	(��ש�����dW�1(�(ͪ� ��@׀���z5����͏��36w��M��>A/C.>-JM	2(�|�D�O�b��[f�6/3=7�Y�Z�ދ;�(}5�pb�,���y ����#��Q�V|� Z�bN�������9~[���o�,>�d���<�%�	�B��h[!�D}�����z���a�DE����~U_q��Ѥ��V5�a��W:�&�L
 &C�o:�Ub�Rt-z���?������I��
�KiV�SdB�r #Ŗ�",�,�����P�,ei��.��z��fn29�|j��$���,$�نΜ-�c"����=���VR}�����pƒ�l��j�I��v~��M�y1���h��e�������{��h�έ������=G	.yR
��^ݍQ��-B�H���'�1��`Ҟ�QT�`���ky䦞�R�>r���Wb���'c�Gv��Q�Ѷz֎[�\��Ŷ��(&�2r���̴�27�������U�HU�WQ@������b�u's�b�S�O���c,��
����sq� ]����K�yY��}l�02M��+��������9�|%H��Pm�D v�MX`}T*ui�nI�(� ��f���F�Ξ������9���Z�rS�B�����A�\��Pi�j�'�Q��D��Jk#|	f	r�nJ��J��E"�|'��p�̹d����%�=���	��d�gI>"5Gh����X��]O"��d\Y-e/'-7v͙�+��㰲��S�j�7�����o)>��j\�|�
��Q�٦�7�aoBE!�U� �ڂx<�gy�f]��G�M���=8~��*���]��S$>XE���Zk|U�������ݡ��)`h�X�����|*���	#���%V�Pj�+��GS�����
��߽U����?��ڹbϺc��N��G�-�T]�h%Z�Cǌ1)��,{G���'�0��x˱?~���D���Q�|W�rRXЈ���quhM5�U�g�W|ݼN�3	�R]������lkJ�2�D���n�Ft�Y�����`�V5�s^�He�~(Q�꒷���,�V�dw��¤'N��:��t����ѩ��h'NC�3��s�%e��c���
���M� ��j�A���oi�������?*��L��(\y/i
߳���j�cYdǽshO���Ã�X���ʣrH��<*(��N�]w=�2�Z���;w�~h���hi���E5 ���/'م����w��b]�Y�ʧ���T�r�qg�H�s
�y��Q����dn�]��g��="-�������4.��Y�!��e�u q���%�`��	����Ezv����u��������a�1��po�@ڇU�(�Ok�6e��?A���r����]�f%i5]{�p�R��l�#��OM?�B�\�܈�x��=�J�o=��a��wE��f}�l��#�f�__x�`J�@{Y0����Lj[V��:a�Zᶌ,@�&P.hk�@�8Ì���ۓ&4�۸"���S���U����ꗜ
~_�8]`�SV��ءRR\��P=(12��	�EF�Oj����n�>��Hv����P������x8�1os����QE��
L��Z�ϡ{�^%�MM�eX�ܗi�����~@��7!H�mU�olv�"�|pr���~��[f�>��`[��6��+xt~/Q.�u�o�v�Wѹ� ɮ���Cf�}���\ҳ�1$�PEBhɏ��о�j^lťT�\����u��Tb����(y=&����
�4����N���ؐDэXG����a���2���Iz[�U�A>l����͐ ~M2��!]=@jCn��j����-�`cp��"	F���ko�F��
��G��sc�ॊ)f�LP 9$�7T�#��}���F�<$��0m�����0�$���Q_�g�.���$�V����J��Տ=^��՟�˳T�2��f�;�cW=��Q�'���^���	w:��]N��(�W[���9�S��	q1y�"�"��qZgQ=�@t2 ������Wmi<A�����|�S�M���<��2��}��Xp��S��\�p/�K3��UWZ�Y�acvG�ư�ш�W3�(��:ke��-\uRV��D#��R��o@��O��;�8�3*)\7�ܺ�^�� �Q0�,�p��7�Ŗ�[H5FI7
�����|�b�Pj��Ty2hxy�]���C>J��,�\�� ��m�ze����d�5��ω^��YhU$Ow���S�J�~Q}�����Ws˓����){��q���%�]���
gNm��ϲi�J֣0�;����ކ�d��׈h�Ş�45��z��5c�d��l�ES���K߷�&&��tn$�bMvD
�HA⓯�_f=���2�����6ʧE�O��8 ��>#���Xo��ꖓX��tW��x��� ��M��`��ӱ�v������,f�<2���ጚ H�4T���9��#�L�¥������ �����ڠݯ�2��M��'��y�ܿI��d�y��+�U���60q`K��T��.�$aC�l�����)�*���]���Y9�����ү���]��ΈB��X %�Uu�[�;rF�	��k�$�ڳ~{j��:[�6lf�Ju%�^%��Om�%���B���D�q�*��6�}=��xG�Cĺ���^O�%j��*���.��`�����!��2�Jdɤ�� Q��{�#�C�K(l��,b��)B�)%�G%��=q��R})A~{�ɱ�X��
j<������t0��अ��)$�,����������""�_��n�2ɬU��Wy�*�=c1ҕ��4k�WC	\�c^��B��p��RS1y%JJ��vI[�)5y�KB����,���hَ��=�;�L-"�`xpw�ŭ)G-���$ʢ�����U9�������>ܣ�r�v��-��|P���HL8��rh�t�?f!��b�-6�2��y��qLL;w�L��w�fe�"p�nȻ�C1�"�")�A�?$�/�9E|�ӕ k�O}�����4F��|���YK�߇�Ĩ������f鬾��!��XT�c
^z�,�u˸��t����	%��h��H�$$�6e���(u�V��C^:� \X�VJ܏�G�q�� ��IC)�X�ZxÓ���p��X�u4���d�׾t�+[6��\_Q�<�z�e2�Μ�z��ۃ9޼�Fi0j,M���7��웿��_�[��y�ţ�� ��"�%�Z�Y��\��Lhi|�\L�����Pa�{o�\����wB�$}�w�J�F��j�6X.�t�|oJ������B3u���3I�j�(+�|�W�@��_EX��$�U��$���M�1��P������?��K�Q��3�6�k���2b�T|t�95����ze��8k��e���/�.��1G�I�sb���d�M�c\���k�0�W����X��2�����C�^x�n\rgIOp�L`�.5��"�P8ꫲ��~�'e�&�p�|�_l]��@N�@У��s�>k�X@s�]H6O�NH�]��`Î���'s��cj�I��g��%\��J�q��'��:y ���������!rR�j��v�bP�[j�M��]b}y 鈈��A�M9.����Y���U�+ŰGV(wS�Ax�E�d�2��.ف��5�:�#˘�(��Ġ.�/�
o���Cb7�&����-�;�Uw����s;�#Q� ����=����[��ȢS��ۮe�V�#a�dI'OZ{J"@4�a23F�j�ZϠNaq�t�oȾ���<�����qu�;9�܃閎�ǋ��L��El��U�����6+D���˦>�6�e��F`%�1��}�M؝�E�����e�� �!����I�(!�fYPe=�pnIϤ�ĵ?A�i΁ ���"ʊ�3����Z��,�1ib�֯K
R�|����R4�#ކ����x��f+�E�u q����#vG��)��{���N�,��2��Q]0�)a�"JS3:����uV��?�/]�Z��@�[fl���z&�J�6��*u��gy+|�w�y���l��5���U��,_V4��q�y��C��k��ŉ��8��4��)�dЗ��b�i\l|�3Rd�I X��y� ��q�U��-�D��5oG�F��#8���z2�B��gY�x���7m��R�48�m�}�"�/���k%���A�s�7�8���)/�5��7�k<$w<J)�z
�����>�v'�2o��$e\B��4p�nm"%D?�4�L��(R�������1m�QMEV��B-�4���\�*��W:H 
jn(�8�U=`9�dC���Z1y�70�qywҭi8c	�Ia�x�C2%|0�@'"��9��n�>o�RT����RTf�Z6i���4�}� �=�ƝZ�	��fl$¢��P�ؐH�
6Y�`�N#��3���[��l�7�$4����Vjm���|��";U�[bI��s��AM)�A���۔�h��#%��)?J�uG��h�O�< *na���&r���`Q�Dc6.��ͥ�̧7�Q�)���?o��r:�� ���-8�|63��A\�g�O�����=-޴;^v�هiperl�
@�?��:5CP3�2�V{�y\�XR¶�R��Ky�u�H눥�/�U��AH�k��\`��*	����b���!8k'}�]�^�%����[n�S{����8{��̦�ο�|>?�q�V����Cx�1�1�g�-��D����(ȅ��C��+OD�IN�I���6$�06�.��SQk7#�z�A1����<�?��M$RQ�#��e���*�%�
�"<����f���Bfx/�P�p�uT"D�  �	y��!��:	^Iڧ�����!��TL`Ԣ�ۯTm��l�
(%�
��TW��e� ��h�5e����^�1Xp���>��P2�S%f�<��f|� ~\�Sl]p�
�]M��nz�"�2aQ�w���7����@&�߸��N�f�m3�1�5�=�mK@6�|�T���lzG;7.�f�M�C�wb�lLJb�# ���Q}�t�R`H���.C��b��W`b#�-"f�0�U���v�������s�+�u|��D�'���������5]ע�,��b�N�1�l�n��e\��0�w+8aʷ���P�FȂ�7�Px��ak��i�#WZ	��,�Rk���m��� [� �|��id�2���p�?bX^�I������T��Gn��Ͼ��x�{���i��H/�H�����}��)���r!�W��<zEY4�=��n���u'�^���JdQ�� 'u���Q�<�B��sW��l�Ღ8�_ V� �T�� �:xķ��.Ed~��=���=�遆A¬��!��ގ\w�J�g*bt�UN�@	�RS�w�%a^��	]�#=l"5����`���v+�՚�h�G���{
��Zຬ��� ��I�ԓ�w��{]iw�W[�xWmTG�i�38<V���+��|�Z&;���Z9�j�	��Lh�X���{j�!��Ff����0��%璭��)t3���H� �߮� =����C4?e���F&������1Vxxp���v�3k���p�f�/]%��f����m�\� A�L���s��Y[��ݢ��/T����ov��f~Q�X�0�m�U�r͚�ݗr���\z'\cO�?,����ց٤nJ�ɝ6���;��k�.��]:�y�b��|�u� ρ"B��d��]"�Zy�MR��1q늘��1�Rw�n۟�wҲV�\6u\��F]VT����M8��H��l|��ܿ^0tX�/�dD����4�,7姭�8��Q�|�<���1'�/��oV����nrB�F���{W�7��{��й����詷:7IF56��JC��� ���ռ�u>���֛M@3��^�r���KM �쀘#��0�|e�$��9�q�:�y�W���X���d�f���7ߧ�U ��o�������d)<�k��<~�N�!��ĶU��3����D2	�(*�׿
閡⫻�P�-7�X������SW��bI��A��)-��y�_5.�[a�W
`�3E��$��7f�"c�=!	��a��i������X8	ǰ��֕9#HQ�q��MPC�`��=�b���\r�d�� ^�z�	��azoX���2>�fM���]1~���*�Ċ�#���l9Y�m�0��͔��ΥQw�`�xL9�("�I6�%�:��^y��<���L7��ԗ���g!�fG<킅��78|ڏ���n��]!�J�)�,���-�]�S�<m��[�3�����8��5��*�qGo;*?������wf��'G��hs�j�n��'��c� (h�a��az��������1�=6\1[n<�],��B���C<)G+�BR��[i�7+5c�puS�p�ln`Y�n�ߑ�P�PX�T-��HC8�=���d~���‹Yn��{�&�J�Ƨ���k�ۿ"d�M���� �1
��6{��{5u���/����x�O�P��N@]*à�U�	����p����7%��!������[�QѶ!���L�%�T���4���Va�T�͘d�E�������jD��m�{e����j�����{�Ⰸ�2��LcǿꇰF�@wFW3��~\��8��u	�EL]��'��z��
�K5��v�.>�u?����K0e%Q�'��O�x~���4����:� j����6-E�r�1ÞL�`崀�E�5:��\k��{����?�1}�8�"�u6�[�'�f��R���`/q�O��p�{n��i�X����-�p����د(H �z�ʼ��C�f���\�Bd30�/LG��$`�Y�L�R/m@��J�q�h��VcE3a]-�����w�e>�q\�s�SAC$��.֕��c�is�[Ebt�B�<ag��3�]E��{��줴�E>���:��ѹǈ�l�x�FP��v> �#�WE����������,鏙��Y�T�w]�ܽ\nJ���		,�t�hBKq��)����U����4O���ޝ��DR^��U���7)�`��i�Mzī�8桪\x���ɪ������/Z�G����1�Zv�)%����닉���Q\��r�)��W�Gm�_ů[�����^2���g��J�V��2Ǫ�����S���.���b��v��h�ɴd�����D��uK�G�
�v�G��E����i
�3<����Z��?0Nۆbb�X�E^��Y�ƺ��+�{
�Q�$z�U��R�>�Ƅ�>�0��P�t�C]D�܆�f�߆槿��j
`bB'������G�1� Q�ح�*ٕ
1�܊�#M𙉷L��%T^�}>�f4�Z��D�;�Zj��c��n��_12!��D�R@�%�{���|���B{yʻH�Tx�pf�;?LO�|@kM�]��?>U|�&�Mؼ���n�y/���3�Q8(Z��h	�jެK����'�N<�e&F3�l�x<����alc�X��Bj0@������ �<�|����{K�����蟕pt�N.�k����q�x�L���1Pʑ��7dZ_��i�r@6j�̑f��\�)��7�C�P��^��o^Y�ݒ���W" F��^6�"��[�n���o����(�������l0�%�oX������y�k�]�bUF��R�pRi�u��)�^��~�<��f8U�"�k�;J�_�7�؏�ƜV8U6�!9 �VE=!�C7��d�
���V�)�FU��ؠ�bl�����4g	����}���ػ���>�
]s��u��X�,؁Yᏼ	�U���K�j�ߦ��x=,�:�?,��\du��r��g�������5ʑ��N�ʠ�L@�5��B�EQ@�M�QϫT��zP!#�EH"&��g�72�?�Y�y��
�¹��xiʣޯ�������v�c��eKӾ��T���5!�o|Q=��V=]>`I�b�f�ey���ܨ����}�Ha����b�6^���Z�F�2ةFfMg:8i6!3/�{ѹ�k��'6�~I3壗�|��UK���H�����Kk|�W�1�ᮀm"�rX	��MkM_[�|����P��pF��P*7
��ļCdGD� J��[V��ƕf�y��:R���>�n��ވ��y�S���H���:.㗹R̃;��%�|��*�#��P7+���}z�]SB��L�Ls)��'�K���B���?:=�
"�=��\U�d�"y��{e���V���U�rM���[Q�����%��)�����ߦp��������������5�ݰ�,�W�T��_Wm|Gq;����4������$��TE�ᢅZ:��T���T5UV��f����@�z���jo�%Io�-���0�f�O_#��k9���	C�j�Jr��
�T�F-��.`�4P�Z��P�xu���3
�9�
�/D�B�I7%$#��թ�V�TdA_]���[=�p��Q���?N��$׳a{�@?]a������,	غ��XV'�J�f��q�<|9�M��l��׵��@�[�����"˂���_%OprP�_�s�l���S�@��s�����;\2��)d������4���Hp%[���i%`D������BG�ɪ��@:��ob�#��w�	q �R^����aE7L���y�.��u�7�t1pWm�?���M!��g�5�_cR˶�1\��4'^%>�}�4s@*|i�zrdB�^�Tz� b./U��lӺ��F]CA٫�w��$3����9��� ���7�e �F�Rw�Z����T��[�&5w_s�ÿ�s*��Q̠��u-��BW]3&�vv���x�a:��7Ѵcz�hTY�sȐ1C���p3n�iW�w.�����	ll��Wm*H����qT�N̫.4F��j�A"�b{)"�M���, ~�L:���fz$ �D��J�����`���FT"s��@d�V�:}3Hui�s�@&��~0!�8�����#�j�l����LL�W~�5V����Qjr�-��Y�6���������R���r�.����#��DS��G�d�U�,ZV4�װ�wҦP�0��v.�Ghg�����4,u�
,,��! �-q�h&K���V�j���k����B6h\o0��/��G5!/�V��6��ͺ�ڭR��d�Ȍ�̃�s�p �izL%�a�6�yr��uP�V	��$2"f�n䌹T�JK� 3�ʿ./�u�ק������ �Fm�h�xdy9_;��B^^�{�E�X�8����/�]��^���/�"�c-
%U��LH�ԲA'��g��6��w3ǭj����̈́��>W2�l���+y���7J/'�#���L��%6E��ӱ,Q0,��P��	�C2!�k�(l�M�{`�5�:FqQ���*Λ�u���=�Z�A�K�}�G�F���E��iUv�R�����6�x���"��hR%r�i�-Q�޼�d��Z���[�\��%@7\�s��{Jn%f�Bw>S8%)�á- ��'3T��fxX���Շ5x�LZ<�����Y]�]p+]�� ;�6KJp*��Ō������48��h��cHV��K~9��@jw�0��F��c-�ԅ�Q�π��<�|�hMz@��yG�/���f'��8r�Du��-�}Dj������Ԑ|�<<p[��8f�F��e!�+M�5��[|���"�X��̃!C7�~�4���7�m�5��5��bӼ�!��+��*���It=����M����w��n1�?�D�ﭛ���koS�~"�HA�n�%�@���Oh��@�_�������;6Q��8��쒛�����9۹bIf�����=E���x{��K��p-��,��;4��'��g`�i��f��ǬC�RV�C`�����lѧ��u�َfl�
�����~���6O�\*���duW���7�V���a�jd�0f�3*���E��j#p^:X}q���:��A;���^���p�K�]H�H������9�	��28QTE��E�7��N趃��n�3�����yκL����]�$$�f�+_�}��s�,Qf�"A�O���_�����i�?�Y���A`����R!���5�K��KT��|�� `ܛ�����KK��W��3��՟�T��?9r ���Ô�E�.���FZ�9�OY����H�j�27�v��H�=�o@�,��O�D]���4�j�aê�ؤ���x��A��Z�Osn)+�'�D|ʜ��j�c��|?c���G!~��7�tK5V��){Uٸ�C�� �D2�]Zg(b�;��!���G{?v1ܔ����C��GL���z%���sҖ(ͳ���ϖ4T���!���d��z;C*�ƍ3�m�c#�(W�`ģ��9�P���d���<��'���ы�6��l-��3�v�(�E�7�.utՑ�@�a�I��-h'�GEaJ�9>�HE�2�}--��;�/}p�HI�2�AV�V�q������y���rm������	�-9	L�95�
��Dk���v�=�O�#��v�1˦�������V�W�V����0��)����KW)RhKk�W���C9���ŷ��}F�M7a2)�|w1�"�џjb�h�g��j�4��L4\�PpL���Y�������ز<���bu��� ]�&*����b�����j��y�D�nI#�z3�:�w�e"EP�S%����A���Rw~Ȍ*Q�S=�{%��I=k��fG�Az0�t��(6�D��[,3�/�yc�۴�-�sw�3�9��_)+{zӇӠF���
^~H����ﰊ���;���MS���
h�^d�0S,���\��(�<�E�@�zR?����ي^iSr§�;�\"��gXD�Sv�E4�rV���Z��نgsq*,%�Nر A;���X��t��Y�<h��d�j��!%����3	�.V��@�i~���P}F��Cw�;b�