��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�~��"yAfEi�)�����B
��۩C4JA?ϋ���n����g�ҕ8[���!�܅r(�=����UG�O((�K�`�0�t�s��hP�D)�w�xJ�[K_
�ԈYJ���LݷV�2�콷iF���}Kq�I�q��h���H�i���m�����-�bH1�)��Z�ٍ�jӰtr˥V�ڥ��L���|��qѷ�&GDq��ʻ<�����n �Ꝿ��d�T�\j.+�wH^E����C�]��b��`g���[~?Ӷ/�}3�oN��ѭc�2!	�PC������B�+q�z��*����� ��z^˥���ER�J��d �-+T��o�9��h�:V�%|�]�i�E�GJ��4�G�xn�XV�Gü�g�4�a�K����ѥZ5j#��T$3�"��!��K�jt�%�8��2�Rk�h�ﾃ�!�����h��4(_�YY�ꍪ��w���[�݋���\\VZq������'so^$���%��E�3s��N��9_0�����q�-�����B@�A�7pVbX6��з<d5��J%Mx�)6����L|������n̗���n[$��g4��|ٮuc:��vBu��Ko*
�0H��ŏ��ʡ���ݚ�z"P��%`~}<T�s�r}�
�C���m唜[5'p�j9UB�Y����l��m��Q%?��#C���*H�Ne&$�
 	i����G.P��k�R�8c��%Is��h�z�������Iƥ4�7hm?R��yC0�z<㿥�ϣP'�ߠg��>�������H��[}]\J��j��u��~�V�m�A��w��������L�3�ŭ82V�2l�9�DD��E��B�̀�XI������Qn=��dh3�3�k�"���uu�}2����$�ZۑF�-]����xW����;Wz�D�Ӷ�i�6_�c��>�<dw��I�!o���RuVG[���?`ѹw�B�'�ҫ�\4�}f��dϖ��4lk��X)WBQ�ŉ ��o����V֊s����Yp?�.6�8�y�։�Q:�,����ѫ`�~���x��Au��0���n���9�78�����K���e�<՚�!K¬����O��\�fW^A�K慷[�à�A��{[퇆M��Ҥ�,�`������1>}TT��V*�7q�it����Цt=yBK�&�Xg6S�������
�k*$J�
�,w����Q�#4x���T��E4%�:�����;������gĎ�B���A"p�A!{�� ��8���w<����b�Rc���!�	9F��b{�Y�p���*��N�>��(d�*7��\,4�l�Ф��y��<��Y$>�]������w7ڌvZ���`��x�EvX����P{��/����Q���9�f-<ӧ�����#ǚ����):�vrr����FJ6��=���2��j��:�T�jo �/Ԑ�4J�	Hd`�ߛp���s��8��4�k<�534<�������)�~���+�/���^�u���0�"ލ��~�'�[U�ۧW���MwK�����r��:}%����m[��0���нa�jQ��U#��א�M��@����+�����P��h���:0�vɼ�F;�O��>��ƒƹ���*U����;X7|d`��1%�I�N.�p��r�mIK]�K3�M�5�Jk��a����}"�2V�1��_N\CՒ�&���+��AP��˵I����b�I4BI�5��7���_T?����FCZ����f̹���0��z%�IPWsUػ�i���~����{2{_�/�G`�(�j��D���hx���{��1��HR{�6Ourz1� u!0�F�]m�*��TЕ��[�(ם�^4Y-vɺ�%����;��\�:2�`=�7ik_�U���0��ܢVo�PZ���!�:��ׅ�m����(_\J.�,��3�+m�}I�M)3k�o)d��kW>�u����ݴ�Z`�E�2F��T(�ܔԨ�2�F�x��������bP�i|LL�:��6H[k��~�f�_siL?�]�g�!'�]�[p9A��#:gu�Y6M*=�&B�ݦ���Ժ�c\؜�3!X[4e�=�{"9�>��^AhNB��Xx�S���2����F��[�nS�e�x�hRЅ���-R�g$�nw*����Q�Y���-�����7�3*r���Pwhӝ���N`+�`��At�!֑� g"�5V|�ĵk���)�љ�v-v	$m7�T��b���cT����C.�.��1�,��`��HFQ
]{����hg�~�o��j�7+V�8�R>oj�]!�*-�ef��.�ٟ�sSL#o�����L�<0�,w���-$r��D�E6�J���NV*�w�TAr�	�(j$D�!<��ճ2E��8��	᮵u�b/!�2?}��ew	Z����u'�3��ݪ	Ф���.��8C=�vS�8�Y��=랠�\nn�⛂,[��i�[�V���	��rǻ����dHo�CLU���k�P	$r%�����rݦD.�܍ɸP�Ŋ�8�x�kߜ˭�
x �*P:n�cV}�^�~���,�6�L�G���Cڬ���Ĝ�텥.�\Sc{�-���;���T
����??h;�.q�?��������2yk��r��_��*�Q{7���;��']��a3j�|�cJ�8��V�r�B569&6�@�}Гvk1���A��S���v�=�&��Z�0 �֋K�B&��ϒ ����L�u��T<�n#z���g��@�6hF���M~dm�K��g�B7�͔������^�!��B�?۲d닱�E$���ʪ���M]!˺8}���]�����p�0T�E�Zu��������Y����\)g��O�d.M�~�2�[���A��IuV��Ҙ�֯�O���Wl�R���X�B+�q�\����F`щ�L�0�D��L3����,��ɐB@d���h ��;�$�68eA}������q��S�7�s%��1L��,A9�Y���n(���C���=Wg���`����;'��j���#��J��u�~�B��	C�*�{L��2GxC��M%�ਿ�)�$�'(�jd%# �zq�TnE�S�8c�ڕ��@�Dٲn�
�A��JJ��_��
������H�4�?��V��D��O2��xN�mڋ
�ÈƆdb&� ��S����a/���h��Iֿjv#�K�H? (V�tѿhں#�zo���ċj@�e�@��\�KR[(����{�����:7m¥B[w�P���s(�K5�1B�,���4~+Ǽ�y��v=%�7:�䟬��m�uJ��+�9#������vW��O#{s�ߕZ�%�XH8�Z���-�B@�1k#�0�p�]��l��7�^��If��)x���j"�!����?���4^��f(\=�Zs��V�"�c�����	���G'�[L���C�ڪ���N��:�
QtQMԭ&�BgiA2K�+�'���L�ޱ ��
jg���C ̦�_Q>_�e"��)�}��������r��L�K�1�H#bs��Y���2���)�u&��$� �Q�������
;S��멱�M*�;"��E�L��a$ວ�`)���uB���@s{��g5���8tJ�F�~	dK������Ci��!�c֘���$̊v��"8�D����8g&���fs�NfT�]�V@�]IȠe)�a3C��"��q�j��0�Qw����/~�f�B�RKY���i�i�uċ��-��0�y����AC��k� _x�d)X:D��:kPw�P	P9����FCL�x�A:�k/��W�+g�I�/��;�r�G�r�A�y�Wn��Z�~X�:o�O6����t�x6������Tu[%KŰC	iց�� ���S�6 
��p��{ټyA����r1���
#*�mZڏ>U�F�䒷,��E�v�:��/� 9�iY�9�CM.rdn[L˹j�)��z�/a?�Q�NTV��.n�1П��P3�'��@�`K�Ӄ� ��C����$Vp%�r����36�_t��(�h���� ���'	���g��|�3s$� �2�tM��P)�>48���0~��-�he����raX="�4�y�����ʓ��C0J����[����F����V�`�7ai��1BX(3}�^�<)�B������<n�&��D�}𬜮�3�K��7���)�����1*��?�>�#����l5*m�!�����T~.q뵁�"��s�`��$ H��*���Y��i%�j����:�d1k�Dcn�:�>��]���՘�yք���3��6�>c@Ql���B�����z�F�'a��ݍ�I�7�ݞ�J�'��5ep��d^�{1 �dt�L3,�����ii�@��YY�Wٍ����U���e��ж�&[�xW�!���.`��v�K�p�5���+�;B�J{ŧ���٧5������h�*�	
�_�4 C%n��N�('p@�|T@���ʰ��W��F���t:�_��2�bS{�#�,)�m�n�fϪ�n��z3���4C�����G�a\��k�Q��d�ڐ�.��,_��So4跍�Y���{h�J �8f}n�U��*TJZ�GS!��������qXۊO�p
J��Bh��($��g�!�:�f��@��Su��kԇFb��?�<�b,�֤������u5Q�Y�+j�I��8		��5g?ג�^Ț�m��H�O$��sL@��7��uI�:B��V���:fX�`״[.�9e�P#f��5��+�Ӂ��;$G��� �I���΋�2-���/V��<l.�9�i��|��|D�x,j���{u�@��#��+A�y8�M���ZD�{�6���)��VT[?8:����eJI�z���; gU���")T�/��K�ʡk��V��qYF��mū]y��)|���!A!�l���K�VY7BT��ԀO��h�u�&�v�z)��hַ��Q?��Z�rT��G�����c�)�*���k-l�L�U��״�s��NT�v��2u a�g�:��B �Rh������y����6�ē�2Fz?����ʷzۗTO��@�s��c�j�;��{��q�$���W{�5xL��6 ~�ph�m���e-4�ش�n6��e��55����laS^ܠ�ܣ�Bԅff�|�hִ�h�By!u����[��k��^n��Rr��#��=i����'Tc�����.�pnA�/��s���w�Ir�}

��Z�U��Ci�q�~$�j��O�f����`��Ձ����<�k��o*�����]��k����Q��̦/7(il���ˍ�ʨL��?�Jb� �豜��>iy�%�VGF�cW7��f�ܛ���ch2-e��ϱ�WN�OӐ��N���ݚN¬l�z��ws��w�. 6	~4���=n�4���,}���5o�v����d}�s��i�u2�l�5ON� %)���T19�Qg�!�/�8��� -���g,k��aUh�6���V�}�����g�\KE��'��Q:~�����&J�Kl�(�����é�6FN/������3fTO�z>��g�`ϥ�;��j�
Ԟ�����M��xҀ��-���A���k�s3�U3K6��$�'���ՒL�p��)"2��b��ᩳ1�H�V}��wZ�<��(���a����G�����oY�Kܑ�ˠF
 ���ҩ��R�ֲS�Ɋ�Y�o�}�1��ƍzM��+���sT���ݲѝ���m)<~X�-U*`N�H���C7,4���3 =
�����l;�ZMÑ�����N�P�D�`�����nV�V6�KX�#�wd�r�"@XȜ)�D�uҺ)q��_�{�+���7�*�Հ� `��대��y�BV�����h04�R�>�c;Ԓ3�Ƕ����6�Y�Y#�_��]�(P�k�v��Ą��Mt�s��+��z <���H��Sx��(?��i�P���9���=��e��Z�劖��u���r"Tx�?�g�~Rv��|X���<+.�C�rY8a�n�fN���~U���dt�`l�r�o���S����®�>���um�~�cu�G� 4��-�3�#P�P->}��n��I�0ɚ�5��
B]�@�"�=����aW1�p�sF�e!P���g�C*��Pm:��>vp�v����1v��aP�P	3�)ɚ��@�ܩVHvr�\�J��Z�"喦?���S�� +��lP�@��ݕM�sSӳ0�t�Q9a���Õ@s�X��N�o_��ۍF��4�(�u��*��'�������ydI��� �@�ޭ{u�CM)�[˖����s)���X����W�_L/W8 jޞ{V����t�P���AN�����?Jeέ��E���S���+_�B���Gsӷ�6M�"��F�o�[Wq��ΚZa������0~���������v�?�:)�i�/�l�Y׬B�w"$}5��� ��,��k]���U,]�P���q�t'(�;�C��I��˙�X
!RУ5#ڏՉ�����'����$w$����U�D�ӡ�l�%��/T@�y�+KG*���� ݋K��=I���4 �"�+��x��A����rB�I�� ��2�[5��叆Sp�p�'��½��4Mj���F����}�).�p��B��ʒ�v�1���]�G7�a�hr�#�j�F���10�"Ҧ�#�	�j	�IX��]z�?fEQpNx���􋏽��8@/���ی�ա�3��A�Q0}��gK�ڒGLQ{&�T��H�#�8�Ux�O��C؀X����5����:�h�j� �F~��B�����~�T��"������e�3�(�u�=�>(���H@KWdxռ]`�",���^īU+fXU$��EŒU�-%�.-�)���~��R�>��t��>,*6:f�)��*��S�ӊu�A{��y�ۀ Q��U/dDf&>%l��;��4w2�R,�
���3���dlٸ/��rg�����`-�||�34��F:�*/x��m%�/-�f�'0�J��o"r�����΅���ý�_�����CWD�x�:�="�3R`�6>Y6akS;���"�`s��Ĕ&⿤Q�$΋_�����*yU����b�k��P K��`G�`2��U���
)r̙�������S�����#��A*r��17?m�&��T[�>2�W :�����(��O�����W>�-Ed�198&%�S�����Xu��)��SeᮖW�bϡ#'5�3�OM�N^��0�F��z�,����L�xQ�7�	ˉi9)�].�Sᚽ!��:��B���̨{ͳ7�l���SY��U���c6/��z3:X]����y�̻]�+YP�ŕ����KYo㇂"��P�8ߧB�~dg��9m�
�� �8hZ1��B�G�܉�)�L����/|�h��I���/6������9t�[�{ ��YD7�\�t�&�,WԿswF
�JWG����^�v�e��0�'Uor�x��8f�$������K��{�s��	t&>3t1)z�9�~�x�3�r�]!�;U��˖�g�hZ�+��B��%1Z�J��N�����g�\r��#ɂ�B��@�r2Tg�l�`�]�"��s��[8|d&<������믰�E�/�Zm�E@��0�]U�%���ĸ|�ۦ�Ic�F��v�
[
�F�_D�2�0��A� �d��TLV��z�A�9�x��K+c	�2�q���;��q`�X�#[�ܳCB�J�L�����ܘ4z{
&���ynO����Bd���tN��R׻�A���BPP�%!ͽ�f�+�*Enޠ"Z��x9����aP ��ݬ�E)�Q�/ƺ�d��T�2P�������!9��/�]hd��(�[��n�&(��1�Z��^+n�B�]�>*�:��(u|r%�g]��&�rl��7/sQ�0�i�k8����^~���Ԓ5�N�䵝����jqe���Rq_��ץ΀9�r��!�O,���0�FP����Q�L<E��7��@��S(���n�"nZ>1��	�T�SBM~Ju��p����T�����
\K��Bv6�t�sX"��)�#�?����DE�$-��W�(��뢲T95�y� v��>I�"8>���o��v �� Xd�1_*�$*�Q�y|.y�[�7���g�]�6�{=�nh��s��pv@R���婱@k}d�P����9��
��M���/�Ŝ���p��6�KR�Sh	K�R���x�ږ��k���ax���>�f�g����RFA�����3��s_�g۲�Vaj��c�Pw�o��@���.�z��@�^<G;��C�Ӷ'�!�����FQ������G�#0�fm�m0����$�)�ׅ���+����̚r��i�Ydl���;�-��z�?�Su�c�թ��(�p��T���P&�QQ4c�
�x$bCd�a�c��އ1��ŵ�9Ӏ�#�~.8?��SԨr�����ܤ���!Ą�O�dG|6��SG��j��k4��E��c�����j�T�<�L��n��8~�Q�n�A�բϓ����5-��?�֯�X�S4�K��R��y���7���]O���N� mK���dL��B)s��r<DD+�c#-3��#)��4ٯ���}��r�v���nnu9I��:��3�I�=���T��|�bx3��B�G�{
���#ڪƩ7�sw�y���[��7
���{�P��yD�f ��3��S��:��q���a7D��%���r�S*p&UNb�ɤ��!�t w�ye�a�n�TPe9��@�Fe�7�7^�`�(�hqN��_=�'�W�OFp�4H_���O���MN��	>�n�(��MRmy=�O.���m��^���k3]n���zꆭ �r������Gb���q+�����Ы��}A���X��@�gy�ܦu�<!#���m2�7ؼ�>�+�O)�%�,�r< ��$~W�.�,��>�+�	6�(W�5���2�.れ�Uy�d{t��w�bs��҂M��sF0⿛SR�tTw��"�6_���Ә4/Q@D�4�Jk�5 5��.�,-�e��Г�#)�>��5"�ݣG�9��c��<�g�e���2�f呮#���
Y���cW��1{�,�����Gv�?D&&ޤf�g��.z���$D19ſ��tR(I��V����%&���|�TQ�Wɛ�^����0�#t���t?I���G��b;ْ��:"��׆^dQ�I��S�J�ML㣌���l�fO�V5�o�Q�7�]~v"�@;�D��^l�y%�������&.�iG��r�ˎ|Ԧ&�)�dJ�4+Ӥc�i׌x��=�5Uh�����cU4{�ً��$}��� 0�A��+WJ7�]��T�M�O�<~��c�u	�+/6�|_Я}Z�h���CJ����ouL}0C�;۳��er���۪7Γ����q`f��]��rUNLzZ*�0��%��yRu|��%5�0As�7��΋���M��nY�g2���:��,]z���镚�JV'|42P��V���5EͨŸF�J{rv[�j���eޓD�C��ה��0���4j� ������
^ �V5Q��+9���-��?_y ���ë�^�AU�7e��D]�r�$زl,1Ck.��ڿwr���d��p]@��4���V��Md�A��
�r�}����b"3��_;ʃmњyH'ǀtz���;�.{(J�2r��䡝Qj�!c��d���W�{�:zw�Q8��������x��*)�劶�����n콛^�B����&8��Ec�:'��!������s�D�2Ki��3�S3+>���ӰÉ������{�E��Q�`*_����f��������x��9��Ru ��0�؈*��8͙�ׇ	����\u~"��C���L �P���~��⠕�O|�I��-ѭd-�#F��ՙ*�j�4�DQab�(9 P�O�������q�Ul�}�7�L��N�N�*mQ��t��F���,YNG�W�I\;����WĞ��9=)>^t�� ���򤎭j��[��d	{8�[	���&��&�Ȗ$�X�9�:�}��_������$��b �"|��H>�(�R	I���6����L�=Rk�duD/x�鋏�-�	�4����3�q<�����D׺d�Ä��҇����u�AHa���Y��4hc�>�r浫m�����M��rE�O^��_���Q�:�֧p��ܶ�c���-��Z]����MW�����0m��'�9@�;�����eh�u���c�)���i�6'���P���o��m�<c���m�)t�15�C��н{Il$�j��:U�;DO��5�2�P��p��w�6��zM�XS�vP���c]�%�'��d�) ��� `h^&�x�s���E�����{��}� �{��3��qk�T�����,7�!�� �7��i�&�@5m���m�'p:�i��(O��2��F��ײ�N�Ѧ�l��JK�z���m�j���4�)83Hy[�2!�/�~�i��l��Ct��bHZ:cؗ�FK�"C��W
2�+2	�A�Z�4*ր1�җU�]�O�?��P���>0�;!8�W(�
A�ub�ĝ��)s�_�%���{y�9�~�\u�F���ه;'5EH�\֜^����ɴ���:]�Iz2�V&�&��w]��NYn��{!E\Q���B���)B�,�Q�X��bXٴ�N���ŁO]��?Q�Y߂��������d�ܽ'�-*��O^��}2���Q���삵�I:lm��):@$^���#�q[�^b3�T҈4�K~b�Q鴜^�ô�B#�RCu{�_�� �Y�ҴƚM�K:�.����$��#�7{�=�/(�+%Z��Cc=�V���u�%1�����BA�����9�ІB�+�&w��cL���k��,TU͏�%`�ϗ�.c�$Ncd��d��q�(� -Or���zx([	2��{��`;~ʡ,��h��l�\%�~�� ���m�ȷ�@uW�Ꮦ᪶�.�`���Y]�O�D�N�u�	2(���7�F&ϝ��֤�,��W�[ҕͤ�1��ξmBU���;$�6��(Y��=�
Y�����fXg-��6ȇ��t^nc��z���F�0�A�s͎\U�>�PZ����bkR0t��1�6��w{+?ȡ����v��L`��C�۹S�Iu^��Hmv��8{��co�ø�2ҋ����jKȯ�^=/���w��\�X�����L���9��=翅 +<,����&�N�գ�:��v\V�Y`�~Nv6�i�����#-C�>adS2��WC�}��k�0���t���ھ"w�N x����-�B��
�!YS{�w���=nՎ�ʺ.M������G]�aF>@{]�����]8Z1i&�{�l��+�XOV���w`��I;[W#���P�{{��$�1�no(i������K�>]��穷�kG���)��;l�n-�_����q'����v.�qL�p�ɲ��m�%Z��I��rG��߹K���z�22��Y���ځ��~�k8�eD��;�(6�A�T�ϫ��q����~*�;x�c��w�X�tB�b�BS�	�ϟ�T�)Å�F0�:�%�G�>�0xSG��6Fj �� �6�rm�ڵ�k�-)�+��۲���m�}]���n��;�Z��B��]�Z;et��ٷ�3���@&e7,=|p��}ԚHE�<�¨��V� �z!�7@���wqu�^����>��U�苐
��W��V�&�W,Y���T$~�z��N��n<�c��oB4�zcL$��n�vάn	�K�N�-�}v\Y��|t���"��¨b-]���0�(���̟8���r3Q��6T|��5dE���?u�h���3��T�m1^v1�W�~��I�{�H���x���F�g���0�ԛ�J7��h�!a���#��s`��+���/f�4�;�Ew>���YN �����B)^��U�&��J�������v3F�v��9�d��o�|�4�U�f"	8t��x��z$P�o�~���q������<~�(�"X��U�:�S���F�}9��ӻ��#�����!�:�]\.���ݐ�`�-��ǔ^�x
��u	}i:�E�D�����4���̍���2���s�(�O�hS���_u,��_6�"L-�~���dI5�������A�Y��h�����%��l�h����)��Z�Bf07��M��2pз�לꞋ8wŕ�FY�Ѿԓ1������Bވ�$=$|��FSW���f�ɭR6W7�&�E��5��j��݅8��7mņGR�soc]�6h�?G��L���3���c�¸��>��c���VԤ:��p�eO�U������/����Y�.��l`��v���M7�j��	��,K���<��9����[�]�\b���'h�|H�@��PN/����W�s1Xpw��Yts&PSRT���n26G��u��F�o���U�n��Dޏ{	Β�n�j*3\,h�x��y���
�iY��UR�8_A�Z�
����]�+��5Ԓ��������2X�����E: �{����T,�M#�]\�Ԅ���j�̕ŤV�+F#���͸ZP�3�D�Y4ىbk+8�my��!�G�	�v�~z�h�V�V(���]��6���2�����u�)��M@��<OZdvb{���Vs��%(A�C��*��&���������g���>2�&{ZAEg������2 j����>�n�'��ʐ^��;�w٧h���L�|�A��%rw͋lΛ�-��?j���Ѫgp��4�p$UeW�v��������8���I�u5w���tqX���N)��]7�M�x�=�`G���ۦ���^p���*����c��'�h�Ƚ�iCD�oI��@(dT�/7'�l��i�|ۂ� T2.��o��3r��N6p�s��}4���A�5*�_�Bn� �a���%��!3�P�[yV�$��-����V��L�Vl)Gj�_�}_��ub�ٷTw ۽_"�Z�{C5�z}���XtG-����|��d�>\߀�&����W�֭�h�2�`�����ƈ��V�������]T�G����m�N?��+՘�@����y�:҂N'ӥ��Cy!c����{s�]�\G�M�7� 5���)�g�PF��S���T(${��\��Ni�O��.�P��i����4�a���fT� ��jv�7t��B���t���
�o|���\��h��R_O�Y%��% ��خlc���1�	Ո��UJR ��"\�t�)3U��OՅ�t�d�W<~�75{����I�Z�i�I3p�����oH�W�/�{�ZKP�&����s��}���T/^���(I�3�Pu�cRg_�My��߻#3):�]*��QN�jڨ��
��1PB?dpC]eE~�u��w$C��';t#+��s��J���9���z��x����Y�2��$0˱3�X��^�2E�ͯ'�wVEP��2����{�/�p����"�&�����%.�2�5�!�G"Y�5ʺ����ҔЕ=>�h}	Ml�e��!^�#�I�{��LW���A�Y7�]��	�N�)h�%��%m���_�n�ؖeϲ�˩9����0M��ʯqu!�bl�s0�p�aYU�H��x��]���n���8'��_����]�h+���_/�S�N�x��~:��p�@X�"��@��t���̭%h&��
�-_4�I����m�X|����GHw���?k3��=�4��~ �=�����6"��@�6���n�UA��& �������b]�&U긤ȡ83_ .�D�J�G$ƛ�Q�����zSM�V��W���}�d�����S.�4H]ʻS>&������-O8�T7;Z
0�U~��������g'����%X�d�x�e��Ă�.]+I���r� "TPq��f��n�(s��AqDJ�߾Cf0� |=��Z=���7��O4����I�}��XPb#����Bɡ�R����U+�	7�[8觫�Ys馱/������O���;l\h���iJa0�m[��� ~�]?���f?I�ח��t��]�W��n�ɥ^��%�A,C��[D��c�g#4�+�:rd��ιz ����p���2�#|�,�A;��#��J{�ы���\�Ӛ[���Ʋ$'�a��>�{DM�?Fu"�8���%�۝���?G�c=���n/���<tѦ I���P�\[��fkO�3FWXd{����:�5�y����*O�*�4�1��]�6��VfuXS��~T��r��u��*k��";�K��o���� �Lь`�4�yC�":+Y�h(�=L�\��ϯ���AöyOP�~�3�k[����_�J@,{��e�X�:E)� nA*��ՁJ�q�b��t�45���,�B�>7��|'�b"3wY�ӄ*R�� �������-f7-x�[���wS�[p�G��������*��?|�����%��W��uYj}�g9�J�W�Ԥz��^�A�1�"�ϐQ�SAC'�Z�9Ct�<�����&��X$,�+���\��Ԁ��w'��P�)�NI�(�[����	F��W��2�p^�>�S�b����i�K�����������>�seŨ�2>GCd.Kg֘���k?��+k�����u���M���P��ɜ�o�ډ�5pv�򩲭d��o�8�p&�7W�e�����~})m2�i�^��	S�|�O>W9�g󉈲��TCӌI�/z��L�M�Ɩ��ˋU~;�pA��J!��H�q�23��n������0���X�BG��H?�iv�=���� ;�=�V�����7ЃF_\��3��dD�����6�k��Q3��,����L�enM�쀘�qX�����#����B���
yo�w�P%8n+������4]R�����a����Nb�*����ǸD@v<a�-��ȰE��p�?`��o�@>?�x�/��"g��ƴ������ѭ+k{� [�o��77;e0:Z���3���B�h
���3���(KS��ӡ��Hw��|�,��~y�y�f�S/�↟�\"�56e?|�ekM�C��i���l4R�Q���퍉2v�#��gC�3y�\��3N�Y��O�5��U`V�+���dk���`&e��U����`�����n�)*�VS�A�`�s�q�(1o�br�1�'q����x�|�5��K��۶m����p��E[h"�6�I��b�q	*��)b�U���=A�zRT>T�h��g�P=�ݕ�iJ��`�'{������ (�;7CY��;3�����H�>�_�Qƚ�TX��9�9.��*ȁ!�����aY��M�ٯ;Ύ���C��k3��@.Y��tC��¾�>E7'�)&��9��Wؙ�p����O�"�6kHd~�$�S�k(`��/'������N�w��|Zc#'%֌`5�����!-�h�/����찢zMO��Z�+㏓$�u��������^F�,�*��7�_��������	�v�lH�<@�^p�!L���i9�@�k\��jD�=&�YlĀ���2G;�-�6�-��L�g��o�?�x����n�4P�8L�a/n�	�B��Mbz#��	��a��q2�Q�i�_Y?�n`�]�	H�6�<.������(ʔ����GJ`�&��D�N�x���ww��G�n���2�{�(��)�|C���&���(�ȅj�h�WT��?��vH��>��_�U6���-S�1
�<��U���1;HN8�iX�I������A��L+I&I!+�Q}?��i�≄bn���:�<�c����r������H��gc�UI�>�mS�T�G��L�@���:����H/���OT�ܮ���ጷM>�ǒ�^�<C]���v�0�P��O-b�ɪ�g��5j@omZ��m���^&=z�Zw���h�E�����ZXb�9a6��MHG[e�ր(]����k��x���!Q�O+�������걪uY����I%�֯��,��!�E)���ط!�����7�BP
Rk�Q�P���-�=z�GѦ�m�h���S=��N+4.*�hKiF�s��q�0J��B����,�O�� �}3wؼ�R�7HTE�y��Hd���g2�_N�%��O/C����{I���ޙR�l�p}(�ޢ_Ԑ����x��������?��u�06|k�������cx���xK+k7���(��vfd��^:򑤻����*�6�i��	�d�N��-����UDe��������E��(���s���QJKE	4S�Ӈ��Hf�y ��2*�D�����@(�8��:�î���.�f�n���Su4�I�
�:�Q�g]!��]Rd�S�T*x�����X$�"��Z�A5��!{�G-Rڈ��}̟���E�}�����k���U��$���)�g{�Y�<�����v�0���
��[��\����d�[$�/]�R\=p���/"�)l��h��{;j��;$r��9���7L����p�-y�*?O� \�H�O镯�u�X��a���������{B���	p���<%r�s�!,?��ը��;N��j��o9ގ4./���!=��R�����#Z�S%��J����C�]��5`�@>%�"���#��b+v)��eÝ!������k~�*�Ѻ����ԺGI�;nj��^�y�+�	F�h-��Һ�`}�Ƃݗ�5��D���I;��Xp�`���f\�q���_�6�`(Pv��a]�̓ߗᣨU)�S�b��W�^U���MC-o �)��7�yO/
ŬިȞ�8!�*������t���XS5-W���^26V2Go)$��6�A�q�j�=S,fX%gj�w������C[���޷�������aM*�߶dyo]g%�ݨ#��h�)&��'���G��<�D���^�*�O�����#�5��(f�lD��G���k���W���J���A��@T�������r�ٞ�Y�?<�k�m迆'�,dx��%L1��e�4������w�x�^r���׋#�Y;]�m�U�WiN?AH1E��8�+	ZSG{[��l��Ni1�� >Hg�n���t����D��f���k�[8a�:�t�{��Hs�7�~z��X�:�v�? 0���Ҩ�ͿY�7z�P��*�v��P��3�ʹ��(Kv��ٚ�֌W�dd�<�������g�>��U}%�� 4�)���R�k��O���j�o<�jAgo>MM ��K�x��S<�S���^ �I#��>r��X���1�g�a�7�U���+�Nm8a��`�05ґ?��:
�����T��[V��ݦ۾�**��c�54^�˾�d /����D��S�C���eI���i���x57p�P_��g�G�H2�0MҕN��l:b��k�O{E��=��UI,��c��<��Y��r�M��ps����L���~�?I�MdíLI�}Y�ꔮ����kT,E>���@c�[%��B�(����Wea��[�J��9��XKO�GO�b�n�ۮQ��gӽ�wE����Mx��@�1K�DDZ}�\�72s��e� 6���~3��s]Ω>�bڬ.�<㥻�Α6�q^��Ϸ{ap�2�� @S�7��B:�Q�<�v�����T`_�/�ABT��	�=+�Ͷ��$�L�*��q�=b�|Ú���q�������O%]�,E<���zi�h�'�b'�7��#m�k�=�(�<��v$Hޒ+-xy%��u�����)�Ģ�E��O�z�Fδ]���!1w ��5F�3ߺ��Y�>����a�����
"����bt��R�  ���c6��|m��z�]x��O��C/눈�=#ݔ�¬�'��;E��Pר�]l�\�;F>�9=I�B��]T����L{�\�&y��ԎKա���r���/�:2~�Y�R� ���^����R���W���Zҵ�p�����O�Sn��$޷�S(�E�����z,ǡiY�)1fB���*(Y����Av�;����>�谜�R���FP���X��u������Vۢ�=����h���G�O��6C� -xY��i�5����Ge*W����)Z]���
b�Z�`#R����-�P@���0dZW�ˁ&yO�p���g�-��-�cj�{��{��$����A��Y1I�?�|��`���[c���<�Y�*�dl�/����>hK���?�͚���k�B���w��y����N����$�L�!�g�J,i�}dl�Z��z;��~"�� �N��T�|����}�-$-4����)T�Xlj�z �?E	�!.J��B<7�>N�$`��%�|�/��=���V���>�7�f�Z�3�I�R�������*M��A����30-}��Tk��W��N�gˬ����G�?�AA�qS���v�LST�<��s�B�@�!Hy�(Zd��v�-������疵��1[E|����~����_se��{���#���$µ�@\|9;(;����ά���m�$����)���2C�;'���x�`���UYuaH1�SZ�p��Ȓ�3��!7�Iʹ	�bQ#�Ǫ#�fGd,Iı�Mj�b�O<k�W�g�PG�N�:F�R�|��P�iF��>.hPsy�prv�Epd-�����Η!���*B|*1���gn�e�(��+�k8���7�
� 4���/��K��VXS��6�.95��q��G-�,S9 �1�8�"#`-���O��"B��K�����|�rk߆={O�*T�!CD����\��'&bC�$�X�1"�b�>����G����hv2|�q)��Z���K�A�2?�d��_�"p�b���ҁ���Pt���ܸ�����7�h���=|��}�fgҸ����ZiIQ�,���m�>9� �)��.�aD��̈��w�K�ݲ�D��G��KH�~E88����f?�%%2��`�Y��Ԣ-�*�ݪ*m�������]�KSA3/;��dj�v��G�55���kg�qoM����ר��g]H|�xNQr()�~�>�3�)�	�*�,��j�jE}�y���gU�
/�G������ʞ\F��qJ�'��'��F���s_O�Ŭ��hϤ�*�c��G��:��0��/��Lv>����ݚ��2�a��]��ۗ�?л�gHj����W�R�P��2Uڼ��ӎ3����el��t�+i��F �T�6����q~���pY%�^J^èY$y˭L��6z�a�bcg*�{��Kn=Aװ�����Y�� 4�iT�F�����k��SP�˒��qpȞv]����I�,��PV�1��[�ȧ�\��^��A�h�*���X��1^����io�a.�7�(Z
�L�kGW6Σ�Пۃ�CRRk���P?*.^���U�ۄq#�.����G�C;6�De�}1����~�E�֑5q{["r��m��	�[�E�1B��.�1}��!n�G��/����߷I�С�߸�H]��t�Ϩ�ί�Hq�����&H�=f�^����ď9l��])��T�����Y��:$ �(�;�n�,���>�8�������TS�H��oe���2��?��髱�r���3��4X8e[D�4���f��<�y���7���u���HbvJ���b%�0m�-�i�%����]�G>r���m�����/�G
S�ܲ�V���̲Luv�}	��A���2g�O��S(���	�@^yER9�&��	��dn��'�'z.���%y��be�1����)�ׂd�֧S��jZK]��*��#�������"}d���Z��e^�@|��;4�1�I����%z�R��J���Cd?өWP�C���!T��d��Pb��ng5s�}*2��v:*��߇��P���42���M��\��I��������d��q�'��Yc򽽸��e�>���F!��=�4��US��w���:t�
�;(�L����}�r�G�~L*��$�`�17�:�=>����2�t\��@5��`p�nG��DS�4��ָ�0����"x�_�`7y�u2�-U���~S����rx꧇�>�~�к-��!�Xz�����ب�2jk���屯K,�bP�fqkg��c���'m0?IIe��>�X�{9���	����]��(�
^h���M̠Pu�'qϱ�#�s?]�{T@<<z��26j��eR�����RUT��;C'� �sܓ*�Y���7�mA���h8m���V#sz��v��������/��T��K̕4��{����<�]��;ޅ(G���3��8f?a�ٻ���q�,�f��
KV�A�m�����!�̼�%�d��Z��#���%�u�,CPUsVt��HQ-"AT��UI�z��9�[�?6�`��FE� I����0��D��ÖJ��Ά����d���Y�R��5����z�ژ°���I-�_jⶠf�a� �x�41�$�	޷0ydj�Hy4�%�3>����lO%6���B����7��7��jb��J���ӵkڢ:�y��<c<��5_�E�u��Ogx�Uv)1G�hݫRQ#��Q��k�ԫ�c�»����m�x��ʿ#�ˊgt��_xJ����4���T@�,B���!�;�X���,EáA����l����{G�"ǯ��0�m{��>1�}�s����/b���Hr��o^58��zl����;�b��.�q��d��_]߰E����I	���=eY	ڜ@�p�#*���O��A?m��{wL# _]�u��FS�EYnEV��1鏒<���7m����+�k#EC��rH{b�yЂ1�~N�N�����?��_[R�@��8e�`���,�DR�����q��U�63v߄�K7�k ��ս���e:�i��+�KV��z�<�G`SQ]:��@Mr#T�vh���{o���p�OY=B�j���A���Q� ���ٵCX0ۄ<1N%ͼb��X�
��t����&@�C0+���;� �FPNV����&�1J�T��(�Km_#��lx�@)�nפ�Z��į�|_φ���>=<[Ѵ�����H�_�f>��D Ҝ�O��mn�����1��f'�+κh�]
�Ӣ"����`��37�O��n����v���{:ӷ�����)��XlP�0�~�3��zA���C��r���9�U�q��>)�0�d��Hv�h	>bn��*��)jR��˔�����1�Qs%��Ԗ�O���R(gl���p���
�¨��b{۰X���s�?���,Ɵ�J�P�8A��m��B���p�6*;~=�W��N9'�u�T�.�'4Ͽ]	+�	�d4x���B�r��+�[���zB�^���ʉ���k��R����?o����'C�ny�g�M��`���-y��5V���U�R��kg}���-}�c����<ʶ��7�����O�i3�."~��`o��yi�(��@�$]��{l��H,"uȋ�1�LQ'� HE�{7qT[���T�2�%=~�Z2�3
�K��o���W����e��)�xq4��^�5�)\(�u�	���B��/)���r0��ψ��C�MF|O^3ݰ\���Um� J�|2���&���Ъ'[��Z��keF���5
�R��ܐ��t.�]�Ķ6��)�w���d�7y�J��b��.��z� /a=�o���N�8�����X[k��_��#J1�(��7�ID�8�AE���A�3:;�n��qX�z���a�c�>Y�.jGͧ�T�X��Q�ʿ��me�h_3��p�,t���<�z�z�
D�p�ul�T������R��� K@���hs�P�J9�Mx�?����6Z��MG1d�՚�d�6�uӅ:P��i���(���Wj�]VP�f�r�����X�N-K
���6j�2[!jу.�|-���,x%VW.!#!~\%n!m�+��Iˑ������C��y!� T��h�!�����N�*[��Z�O ���Y(	�b���w��C���euˤ�q�
ɢ�8������pٰd� @Iu�w�&��pWMm�)w}�\�7�T����@���^݁2�;i�g�w(�5��\9Q [`�I��Zd��%�z;�;j�	W������н�|��EWzF9��Xl��n�Q��r����:C`f���=w�}�γ/�L*ɩ1er�Ԕ�c����Z"���"�������ˢ�kNK%\Z}������	!����r�)�'������T,�&��ƅ72m�/!������Ng���P.��j4�����x`c_j��e� M#�k�c�'�ԋt��O` Z�O��.P�����Z��$	O� +���E�<�٥�?X��&�˴޻�"%��c�7o0���:�|��4���*�(��y���-B�TXJ�E��ε�|q���Z�F���1��r��+uD���.r��w��D�e��Ltي�|�$]����;�9cp69�9��\�:fF��^���bn�~�h8a��
�k"O�{Y��'�<��N�/���u�|�zp܆�uO
a㎄���^ˍ���c� 8���ue��Jx'�O��8��M���?�7��22f$�1p�
�Ъ�,f������t�)N��,��b�T�0k3۴�%�$J��T���!��fi�3��Oj]r��< �^��S\��Yn'ɳ�C�]ԋ�^`!譬M+{*��>������p�����I��#�c�9���k�����Ȧ�׌��U�7����Z��'�׽��l�c�}�ɟM�&�����`�fUUzfx/ �@x��P%�]�4-�Ey@<dtkbo�9�r �t��<�4��>D�͇Sԭ�ً馻 �ҷ	��؉bn�&�}L�P&�`���Y�� �;�n_ѷpùm�ܣ�ۂ�9�F(��_��=�|�@]�×���E��a��d��:e� �1�)�9u�e��`ؕ/�$�s����y��(X��7�7S�:$eh�"�8�1<��'W��q�}?���"�U�n3��[伧t��f��I���T� T�j��f#��PB�C��!���>��y���{��a���@���!!��pyE��Jө�V�����@��H=
��� �[��RVI�ꀙ��:��|�V� ՟X��h�s��v=P���V~��O�7=Ё��Xv�W@����_g�,����6T����}�-��	Z�-�4J^�a��a ��E!I����kT	/P�L��l�RQ;5����+��I��������A���k�^�Řļ-����Vg~YW������I÷��J��3��zϓe�L�*y�/5$�d%��i����]&�,��F��'uN�Ȗ�l�?�6�lj��?o~	oЀl��H�X@"Pg�^Z������<����1���m1}|�Z5J��+x[�	U�&=��S���К�oŤbXxdL����$yS@����D��NR��M�E%o�M�z�&tU�0���#���+u�-�Z�/��������<��� ����<CO�ɹ�����/���ItSwk �h�!SG�}b�`HQ�Q������W��s?`$�O$�*�
'�2�4��3l�0	��۹���wA�C����I����`��1���G	}�b �E!�O�eO� m�C��(��$��-�݋by�*���Ke�#��e�?�d�\O>�����eׇ,��;��	4��#$�-��YfhC���&觏ª��&V�:�3�.��8گ�;�wtW,n�@�c�!~
D�'}��q'4�59NdYʊ܎��B&C]��X��Q�<F��R�QEF��@���VҌs߾�+k��&Fh�a�������Zc�y���ݠ��:�	T���+e@�C.�-O�z�}�t#�����Z�y��N= :��D#�Le"�KKu�䯒y���en���6�n���{<� >���q8?Q���̏�����9+-U�)C��ǁ�L1��h��B:�ߢ=���M��a�%� 8�/�P��w\���c�_��aWN�����(�*"1|�`���p�M5P��,)��{'OMn?ĺ������f��$���v$Р��I>a�hR�>��q�!���~���c]%�'b�o��{H�� z�R������bχ�x�6���A��&t�� �z�vJA����[���: z(�qvA��t��p8��>ɏ�6�LsN5���ۚ�����86F���#Z�	(0�rM�k��$<���;$��!��R	�^������Ӛ�	E��j¦?/����r��E���N�@y�����pڵ���*۱����^{D`t��ge3d�7/\�����ٔ��f��s�R0hQ��[!<� R����Ts��&c�Ʀ[�M�O2=^C3�7Lw���͂�r�
	~������'�re���Tf�u��d��s$z,=�c�T&���F3hh��O%�d3x�Yc�į�%X��ʐ���O����A0l
��)����.ru���<�D~�,��,��7]�R6���<aT�,�Ӄ-AT~5oD�41}LV��1�_+�O!7GdyDKr˜}�O!�U��EF�?}�`Έ�OŃ�A�C��=��x�Э��չ�u�_��@V�-�Ox;�e��ě��d�^G�o6��-���"��\�O�C��.�J<�)���G�|mF^��*"��
tE�E~�߇̌��f�l����T��{���`p���4��#-�4Ķ��E�"��S��<s��I`{4�J<V��2p�O�8��#f!z���슝Cn�"%�}^5��;���/�;C�p���y�Z'ю����Lc�=۫�]0���(��v�3�}��'^1��(�����Dk��IfeJx�)S<d�)�>�η��EoV�^/FcLvD/�>9����O�]�2����θ�Z�N���1���Լ;�[�G�ꀘ��pT֗3&��L��%�r1Q��h3����K�/z��u�J�c�߀:�[�x��V�������zt�@�zo�-�׶|khb��=��y^+�>>�x�"����@�7z�!h	*��;(��~�����۠M�B%�>q;s\=�r�"����+FQ�=�6��B���ߖ�8`�`Qɇ2}7��v�D-/��&�� [L�卩V����{��R�k˾�˅�!�2M�����s�O��hw\R&��
���Ԑ��1B �IyV���L�]��l�>zϬ��C�M϶y9X�����HjA�/!�b�}!�]��%��2��:TY���čɋ�q�c64�a��	�)�5��u10�Vm�F
(�Au_�D:|uT��L�!��?�*�8�,�0X-$\7���20�O���h5mk]2,��6B\��1�����L��.�m�>����T�����x����cUGV]�Ғ�3�?������℩�"*���
ޯ1��!��hm߰;V���nV?v�� ���%^�AX�V����9�9䇑�]��j��%,���I����|yu������!P�9V<Ño�&����s\�G�	��b�O#�%�r�V�?�H��z6�@rͨ��41��ؔiF3��v�.�c�M�1���7�����01��]����m�����>�ޣ a�G�	7��H�_310�\\��$���ύ�EVf� �ԥß�~���j��i~�_[_�Ƌ�XK}���%�]����2��j�'۪���
e�|fQ��	���`��Du�, �u▖~��1�y�J�������L�}�{L�ؼm��6�RV^��/c-��v>7K-��V_M�}�ꛐ���D�op��Y�<�bش��Q7���Fω���@3�p�\��-ȵht`1s�lS�_6��f(af�Pw�姥O��G0�e+^��w�R�:�R��T����k)��;7��ա����p�9��~$�2��i�𓎶,��F�.�l����������u� 3�
�ݤ���-g�܋څ�F�?.)R�-�\���\�.�Z�GAxfk��(K������B�3I�2 �&�D?g�~i�q]�z<o��QN��l"��#�r���j�Pmg�(�sq�_�����0�ώ��̨��XS�p$�x��:?�&���:��z�%a����h�t��da*�`�D��܋\��$	��.֥*_٨#U�^_�]fȳ?�b4�&b����e���@��l��ʚ�nZ�K[���ӆ�M6,�n�|�嗱y;�h`����/�Ξ���eQ����]h������C.u!���q$�Y���Dm��/��� ,~��LհyRu%�SԌ��/�g~��So@
Y���Xkn���몗,{D��$��V&��G���#��_5hxB�ۼ{����1��B������;�jq�ITHH:��!2�B�WRu ��bb��Ӏ�\���`���L�~�#�C�c�����~h�|�nK�X��4!���8u�G�ߍ9�O��%s�?H�C�ש�db_*:�H��؊�\��O3"�-M�DT�e�������/��zU���?���/�m7Ó��E��H=�/8�N��V��w'!�+U��Mw�ӀZM�DЩ2=��ד��Sԫ�W˰��x~��a�M�O��/t�E�G���(�����2��PJ |ڰ2��H�R*2��C`�A �3��wjXkv��BM��c�g���H�Б��ĊX�-�*Ȗ�����l��@���]�Hz����J�m��F_�qSp�LR�O�σ�uP�t;	}~�gct�őS�"!ڂ�e�Lz�Ӹ�ӆ��npԫ�xDM��������VE'P��H��`W��3��6�9�S�l��t�����{��ؙ���$͵�G�uc�f��iC)�Q�π�a�[��<�7S~ӯG{c��p�\]����34�ͅ�5�WOOW;�HH�����H��Va���g�R?8��)�ţ��o7^�6x{��s�d�`�t��W8�ݩ{����v��:��i3��Q��y� �<f/�����]���q�����ǅA�{��F0��|AC��vQe�8���~�;��[[H���Be��fui8�h���-�B��\ZS~�噫�c�i��;�!��L�k��$_3q����L�3�mpAU F��3o��_���E:�6^�ܷދl�9������]��s��؛*u��dO�ˉ,��Gk.��A�Y���z �����G�1l
��TA����^`'6�x���.��bf)ގL�D�ƕk�=~�i7�C��
L�2�פ�W�[�4xn��f� �X{�����V���b=;�h�q�P�06<�W'x�����&z��v�v��UV� ���@���D�Zy�B��	y�9�`�z��qK��s�C���yG$�q�d(+K�/�4�ӿi�F�����4,-@��>5�R
b)��t`/�Ϝ'fr?�=%1��Fy}�m�]���
ʻ6�+(�1m���z`��|ܜf�.|��3�[p�G����Mx1�D�}��q�Zn�lN >�h�"�.�qSl�%��uf�k�je�E7����{Q�V�QQ����B�2���F�{�5ݬ2�U�������hQ"XO�,�lGΠ�y�����V0 �2��4+lk-��[���Y=k
3[�d{���ɓQs�1��q�G$Z�,�ߙ1t�9�[����j�Zg�}���x�%%��f���C��\����am������J��?�˰CT�c�[R�wNw(�>���wF.{�����5���'y��}��.sR$f;G��~�b�N�*
��H��Q (u�MH��S�whUN���_�sX��@ܜ�T�T�?jh��4�itW1��Gye{�����Y�_�����դ�lp�=�㩠'���,�J0�	����T�
G�R�~�i�ZK���A�Q�� 	����Nm�!�X8=U%)���^r��4�ao��"�+���TC��!i(=�������h�6��e�v��[ӌ p�����Z&~&��9Qw8�3��4XX�/��0N��jD��o[�1VB�xL��5r������"��5�vD�j��y��YV��}���tX=S��r錞
hPČ7���yo�m�BU�r�e/���?��۫Z�۔O񃼴�m��������( T�մL��ZQ ����j����y�z�H�B�ܺ*K^�*?6����@�W�}�T�Pd z+xT��a�����z��r�� ;e���8��)�ՏI�2�u��Y[��g]Rv�9��u�4��Fz0�� � �8�j7]��lH��v�fq���Q��i�hEfkG��j'Yk���L�ᕱ(r�J��Ɛ'�B\����]��?��ݫ��s8RW��٭��k��
P-�bC�xã���$�V�\�)���c"@�(WO1C"d��
�E5f��������V����1�~��
������ws��^�|S�_٢�q{��X��z8p�O�S�C�(V���>x*=(��-��N牉"��^A���	�aN1e���5�o���\YUu��>�#4��iŅS0R?a�� /+lZ����I�����7m,��������E���Wn�M���S�15�hB9�Z���!����	^Da�k�Bx��q�d0�qv�V��*a}�P,gzk�Ĩ�Td�ևҍ9R�^6�,��]�C]!������ ��P���^�.zE��
���D�}�)E�i� %-�h�|�3�^��9�m�����gQ�Oy1J9-�����qbiF�=�Nj>����b�y45��)M�Fd�zL���C���W�ಊ��U���E���q�l�{��|N}D���s�&�3�vW#������<0=��q�"�jg.q�Sӗ�ReR�����ZR�쪕�H/��9(q�5;]5}��ޅS�	��u����C)�Ͼ�/y�`W��GnC"��#�L@�� �����p��!'"Qj'�8i��㖟�>����?`�5��i��#\�_l�7��kW�7�|�Ͻ����0�lK��'�oc~L��"��R�o����yǟj��W��׊4���Zi���
���;H�Gs���Ev	66��	�H|`
�����@��kը�)�0MZ��|ww�e��Ȕ���KD <"������nY���������<�A`�.VP^w�4�K�1�w4����~6�4 ��=ޗ���K�F��~�6r��l�
���1Y��{�X.?��>�A��
2RԢ=�g��s����"����IA�)���c��]?�X9t�����p:�KF���<���Ҧ�GtK��Hi��V��y�a�0����>��j�4ąB��>A���Ԋ���B�5��Hq�{�U��%�Vw�tm�>&��� ���dekj!��2��69�C4*5s�@��;gy�o(�����+�����k�|FSx���ijt�R�	���^�q�|�d�0)�ǝܠ C휊��W�C8?��5��j�/t�ĭ8�,�� � {��7J�C�,dtG�LV���Y�s�ȏ�r��解k���v�i���ki���.Jh;��YO����D�W��y��!�}�5�E���j�ɨ�c�
P� ��a%wZ:-ê��&*]�-�E��KdJ�ߍt�E\C�>�0�����f�nu*�Y������V�h�4�"���6�3F�Q�]^'ʶ���H�:C��Z.߯�h'�^s�Iu{����;L�cp`�5�?Oִ�������f]A,c�!��Yᗪ��!" ��{�OX4����n&L5HD�U�c��<:ݱ�-(�2��*j�#*ܚ���q:$�5r���`[%_Ȯ�(�/ĺˑvZ�VL3�%�g+�/���ژ�kn&�<8xԅ���Q�*���ˆ��r�o�\Rc�=�-���GVn����P�n"䢜N�i*�����&�l����ԃ�ss��ޣ\���2 Up*��ξ�[,$��R���C
�d���h\�A,Y��m�&��%}[Mi�\n����͠�%�������� 3�G��9����A���f��#�-���h�[x����~��c��g��wU���E�-Ňsē��|��#V��>�cd|������w�ג��
q\ �<	U�A�_0�`��O�	����:OH������G,��m~�+z#ރ]�\[ϐ��S����A�P�X��%�bK/e80}:���R	�x�,&ᤋW��k`�B]��\m5�0]6]�>N��XZ���`ߴvCD����Ki�_Vص����wCB�$�)��r�iey<SJ��D�����G_�9_�8��e����.\����>/�QڝB�B)�zA>��G XWP2N��2��������{��"�2��!�삖l�����O}�*�;��f�5�x�Ӌ�4#=�Wܾ"�Yј��s!ddΒU&ʥ!ו���םo�-�Q,jm�5G�  _��
��+.��ȿ�o�)��r������Y���HY�O_���}/5Ai&:=>��\>6ho�`�RՋ��nq�(Hg��A�a�����V�R{�#�Oz6qh6l�f!�կ�  ���H��n6Q�'+)�8ЙQ�vD��`V'��^���ř@���iЎ�y��:�=r�n��l����YA�_�e5��(�������\r �P9!�k�8�h�4�%%�@H�f��
=;b[M_�U>�}r��n��P̼dh	�2���zy���puOȆ����W7w�_�D(���E������ߓ����[^�
 c�qT}��P1�h���c���WbV���]Ȯ��z�3j���̬�w�:�n"Q-�_
�>!���Oہ��Ul�?��i�K�"���4�n������.�u��\ pbr�.R�ӂG�D�y�����\b]e�#�?���R.�[�d�ي�x�5}h�/�6;�w�| ���㋾vݳJ�j��
dȄ��n���������P7"��Ӛ�k���W�L|�$���\��*���h8��uN�/_ac����R�H�Wb��A��D�u݃y����~�|���4��!�S3�b�Vj]�$��Qqvj5#�� �x5�6�\��]�JTG!�V���ڗ�'�.K��a�E�)������{��^4��)ۺ�Ţ�� �§�)��-W�ϯ��10N��UT�s�1�	��87���E�1����!�V��2���Ò�8V�`����Щ�]�?��3�1��t(�8�Wy� !g�	�mt�JğJ5�إ��3C��&��"P|���T��7�Q�}�֚ŮHЊ���5#����,p�:P$k�7`]ȳ.y� t�����H1D�>R�ҁ��ث�L�p��_q@�����,?����D�$��a��
+�d��;�ڌY$ǔ��|0��&J�Ch)��pAܴ�bx���Pg7R�s4��^q��3LF����/aX�(�{�"H�q�f0g�^��6W����3PX��>�����i�����pٍ)����1lb�+D}Ck��}~b��8�g8��;������
FY#�J9Eo�e�cĭ�Uq}��[��l�$_dwbw��u��ѕD�)HE>��ژ���?:��犃%�t @��?��?�'�<�n��G���6��6M����/��Bx"��=̦�J�Hn�����t�N��O]s7��.���g�Q��)ݿ8�+yJ�U��)?����\�|ǗK�2\�be��0����T	4ZBN鼡� +j��N��?��>}O�~�o��*1����9W�J�>)�q|����=��*��cP3�My����Ӑj�:C��5[���"u5���J[���W}?��`2��C�[X��ŲVIk������hg;)MQɺ��Tq�mM����^�c8���a�=݆4��q��c�9�!J~�1�GN �l��f/ 肤�˧�V�G��@�?"&eU�X���X�a�8��ĳ����,)cB�Q�W�P��+�40�'�m�nf�!U���&�pMe&R�� ��s��&g�ly���5�e��O�"��8ԇ�O�1���8�D�V��I\�}  U#͓l'�&`�����g���	�G�ҍ������c�Ս��&�^Οc�+����
�L�.l��$��S������T�w���d��wf:nJ�2zS��q�@&���B�>s��������M��SS�P���Ӊ����%e�4�(4:���1��V����q�!�It����|$,\!��ؐm��+�8杄��O�Ū`�Ģ���X���w�PӬ�:��g�R�RW:ǿ(Aw��d�ԓ��s�dv�"�����@G0Fژ>Nq� �7����V<��b����7���[�<4��h�k�7'�q�t%C�n��2����S�a�+x.���V��3<�[�H��"V�IOC�?Nc��3�iI�6�������v�� ��&SD���BرN���Fd�g�p�ZY���"��>�	Y۟����b��WK΋Mǧ �0��9dl��y*��,q� 3$�{b7�d���R���b�����R������?�4.� c�)g�֚����[^�
��(�!/C�����\��[���H4:I���Y�]�x�3��;�^�qX${j�~�&�:�Qp�;	)F�w�D���'����h�[=� ��:�p��a�����/�������|0�?$�B&Ɦ�������w�;3ؤ,��
�C�Vգܧ62�&���R�4������\��i5xf����⮄Ӆ�n��m;/���-�����IC��r�w��޳>�o.5� ������ݦ�7N��^ɰ�J)�l]EH+�i3'��~$c�O%��}��bL�${��:�ڼ��[<BD�L�<�ǡ��3i�\$��m ���+��w(��)F������ �FwI5�ᚺ� gA���:akmRи�O{}D�!��o����[#&t�7�a&hܬ��6�� �g�
m��Y���Wdq�<��L�_�"b��'�'�������`ye��G��������Z���
�����v�SC�� ���u4H!y2�ƃxLk�AZ� +Ca�v��4����U7ע�v�am�[���-Nb��F��9b��ž*Ӈ�F�_�ט��p���Z:�īErB�[�)�M���chQiP��@@JI��nB%x;i�32�W�+�JU= �S�F#��1)0� ���PK
UB��<p�&q���{lz�|���^>bn�*+��19�`��J��u�d��K���WO�B���Y�
���Jg/�p=f ��׼bj�IU�Y����L�
3�O���Ռ������\u?���ML�֝�V^X� �h�&��Ԩ�z����֞��F:����%N���31���"���KP����M!��0�ф �Ya��u��Qe �jf鵵LՆ��R��@��"����SRO7 "%�c2'4����7�-\�2���7�E��g���?���$��H񧽪��Yʶmn���QG��%��0��]�n�RjU��
Q4ڼ��`�'�:(|�O��4��1��|_���0c��W�L !ڡlhO�}s�(`�P�-���h���n�������g�4+\$D��2��H�96��A7�צ���|�͂qtu^9ȯ���SK�����F b�%��>�i���W�a��U�֓�U��r���8�(u��^ ՟ՑA�#���m�2c�WFK�`bٺ\șp�0>GZx���0�E���E`�+�!���A����ͷ�~_<��&iJͥ��5��H�*�ݱ��h�~�����`J!N��q7&Sz�0��YY5��h�(����R���W}��v��D��D96!T����嗰�△;�9���V8���� ��\4���.~�dv�S�#����lF`�O�����L�H�����YG�5���c�:���w����T��g�,\u׭n\�~�A�v���GL�T-&z{ZJ;Ҧ���eG����݃a��]ק&[0��K�6�'����p�~*��X3Bl\�hZy�X��}��)�Tɭm?k~S���KBY�꿼��ЃԶ��-��(��f��ٗ	rk��6C;n�ѫ:�;l�T��K��Ly�vs�oZ�6 F�qk��*�NY/����t��!���3�Kq�*	O,���w2܆�`e��%d7R�=�O,��2��9�5��	������Ik���Z����S�c$��F��FP�� N�I�Y=�_�τ3��mw��I�h�U��j�I;�0�l��W��&O�D�P��&��A��w�IB7� �,MlܫuS�Z�_9$���Ԏ�͛j��׀���%�) blb�er�8�S?�c�_�g���֧���%���_�/���6ˮ�-�E�ͮ���FV�R[/Q6�mHA��� �dvX�!�Ie�g��R��gR�O�\���$Z�|��z���;���8Tlnx���\��Xl�}�V'���d�����7R��o���h��v~r�	՘�lO<�Q�6�K'"_���	�a��U�Դ~beH�t'��r�c���w�R��	�vn_/r6v���y�'U0�s��s����`K^o�E�>;q{6_�ɌŦ&߻�5wK���e[�9\���%ϖ�YCۄ�qQ�o\_�0�g���Bbc(kV��+�ո���Dm����K�d�^�5�(�|���cv~��C/��oK��} _Ӛ�c6�1BqA\����~��7W�wD��i��<(��nC��Y�cT[���$5�7?%FX�׎��6�,I�n$3�_��ZU�A>`��N�w��r(CwN ��x�����u���N:e��w%�2RNCn%=�z���e�{�Jۨ�ط^�c�p7:�ޔێ�:�6�ܘ�HM��#�O)	��d�b����ڿ��&�Y	�HY�v���	:zP[�����o�D<��eS w������;��b��P
T3|�o{��kU�eag�^c̍*�Ѻ�%�i���v�ޡ
���k�骛g�\N��hSd�|��_kz�^P`��F���Q�3| j�1���zw��ZȻ���������pmr�^_�n�q~��PP��i�BT����LP:4�3A���J0�����1[�h��?oY�B	zXBT1>᳓ǁrƭ%xSwi���A�6�֫a�����/���wl����c*�;�|�pULWpđ��V�X0�6SxG�S.y�j�k^�E$W_Rl.�e�T?=��Q��,����d��K��{u�������V*�(���(Z�8]���q�����V��	H��|�o������5��h"�֘�*�9	��[��|W
������K�-=�XFO����Ԁ��M2�t�4J_���ղ�ܛ+��	'Sj!u��o�aW}s�]�O��Z�}Э<��m4��ܻxM�lXpJ�\E߬E�v~���i���=D�-�z���p�,_9co�?W#�=�0�Ϛb������AK<sI�h��������.��CnhY�xzh�R�KQ(�'ե㡍Y���~�6��#'4�9��'��CV����LT��h1*�ԓ%�[p��z�߉3ů�Vۅ
�0uV�����Z�Kǃ�^�_0�F#"��t1?S��Kgg�R��i	�X��6b�kOO�>*��`�t	*��Ç6� ߂�hȬ���Q�F-@����C�A���q�	�	#�7˯�Y}~P�D�ӵ�ǋq�3�5G�FY줿_>& 8��q������ ���ELſ������ k�� T������t��W�<\S�`?٣�[>W�M��m�ŝ�Y��C���..�)��n6��OgT�G�"כ����-=�iI '�Q�Ć�R��P�U�:�UTC�p��ݼ3�EG�Y!�#?:��QVʢ������O�Th�(�;��Ͷ~^ϺcS���<ᆷT֕���uM'��q�^�Wy��ʑ�g�m�O�9�B}Y�U��-�������sc��'����6�"�ה,���{ɖM{]Иt�8���g�5�>B�?{�*�����9�d��^�Fq; �_�;��w�S���r�����beq�Yٮ,	���:N2�v3�����6�R��y�:�W��J�]�55n��ra�R�(=ӏ��ܕt��k������멨�n�@�M�+_�'���z����P͈��:�:�-;$f~~���Ш�1�/]���� �G��Hd/0�sr�Z�k��m:�;��q��X��!��T�e�����w�#S�uY�褟ן�8�t���p�5�2�����i�à+��I���t��ɡ�z����=|m�塖����ޓ_�e�����7w�^̄U�*�P&)^�/�lJ����ߞ><���_�r(�*��9`��;	�?5R@ݙ����Qn(|'Zk�G�\�tA���N�T$ᴦ0z�:�un�5�����ovj͒!˜c�{
��B�L&���÷2�BRz;|�>��z�DK���,���ҕ�~�5��ߗ�'9t?wi���Y�a:䩗ƽ�o0ax����gk���k�w�*�zĻ��&�,:s�Ӝd���9�,�m7�(�
��*���Q�Qk�
N^����V�[y�hQ��=�@(^��6\�%���f\�P�L�7Ul�EF#%���`�:�t�^O�O
7v��/�<��=�|�.mJ9?��O���6,rUq�8��~,�.\�u�^�3d��>��u��6��?���r\�aS(��z�10����H,������$'Ea�������z�7�BK*x�m�������SN`�]�I��r�E;���uG_������Q��(8�4�[$�2�Ew~JCl9���})�_�+rou���&a~Ͽʸ��y<���!���)
9"�M8ǐ��6�w��A��L>��͂����m��c�x{�a����s���#��Z�-mr� ���oy�k�� �L,>~4��ڲLm�fдL���jc6E�9o@�9L\K��������D~p�����f���TǗ�[�l�(	���ed�Z��gR��Z\�<�3����"��u躮<�������)2VgT��Urh���Y�-Ch��a`qS��8G6]�5͹�*4ٿ��!�r�.d�j9��5H�j��Q�$����?3�`>_3�/͊a���D�q�@�γO���Q#�	 p(��ը�ۂT��R��j�c7������+�]������*�#���0�I�� Wr59�Q+�ikǇ��N�I1c-c+W�5z���rXDj1=��b��@��&�"���o�]aVw�y{��	ї���v_�Bd܁�#�����5
m�]͞�}�sr��%z��z`lNmX�`ͪ��}{L�#��E����8 V��KB���t�[����,H�ũ��\�s5�k�>!sbr^j����AW�a���o$5�_��3����.[K��͞�q�'����7�D�1B�s�Qi�M�ď�6��V	�37F���l����Vֺ�d�`PO��K�@��XA��z��QP��@Z��h����P��A��{��
�n)*�R%�Bi������!��ihm%~�^��ڞt:n#-�?�g~S��Dx���X���zʼlΓ����7���i4b��#�4�|����Fj������s�p�5��,Q�f��o��Qj%���X+k����)_�vg�� -�d5(�S��{�:��Kt��$%fA�7�#U�W�j�
��g���G!��H��Ӷz�P9F�Xd�,�Bm�Q	�F��� �?��t�8�5V�J�ނX�0�y��iF���:���}�3B�����~��� ��$�:�$�����DA�r��._�q,k(R�3��7ER���ݐʐ~
pq^���j�Y��=�g)�P�xE�%����MBǈ
Er�`�S�����ԍ�p)�9+��u�V�I!������u(Y��KS����t6ԏװm��C�LH��<��Sm2q�.(b=� �u�l��W[_�v��i�?�"4��Yrq� �ىM ISʸ��@4�	���$�} ����ֻjR�!��pASd����
�|`��v�$�i�2��1$��r��6ʹ�S��-s�Y�I����4��i'&��vm ���sB�K�?���bB~^�w�����:K��0��vf�vR5�f��Y���]�xT���:R�^Ә�a�L6��3lwOZ�
-��u\���ˊ�����3����N4:l8nK��oS�ۺ�� %Zp��<`�okf��[���
N������4y�.���l�w�qj�?�x�0l�����	A*���{���ة��1���i��5/����,8����Q1"�)�b+���{gT��H��H	#>f���J���	�t^ԯ	d��lE��o�$t�|�} �a\k$g/��e�J�p��x���#��kR��9�D��ze�	f���l0����
����L��rW��ar�%ݖ�\��3��1v�,|����M�pkW�֗�a�x�l�p ���+!
�>|����.zW�=z :� w?���!�[��Mę?�Ȑ佱
~w��ېi艇ن����U�5�	�lA��b�t<iYrn�9|��A��bF;���f\硝���,�'��X��(	�y�@��O5��s�N�.��'�kM�&S���D��H\����e"R��9c�������px���Xֈ;rM|�ָ��3�p� �n1�_<*�L�4V�gRc�S�6Vؖ�b�&��cP=��Zof;����wށ�$i��tk[I��j�U�������V�׵���T��h�ز����;8���FXh��B՞�H�&<���}:<_�#���;��ҕ�r~�/�*L$uq<��Moϵ+�Įك�jյ>��L$�H�Ъ��A� �hD�e	6�!�\�%sݵ��o]V$J��j>فDy���ԇڌZs|�l���x|7���Bq��r����q�d������f�NUhȻ(�����J)�('i�aI���aDQ|D#N�p��N����ގ�����g�	��mJA�+=py�e���㦻��:���`����F��d�����ev��5dR�����L��&�J�͢K����$���p�7�n�����4�Δa�>�� ����hH%(��}��e��Bjj������>z�gM$}
� ��q%�H'h3F��;�0Q�9���ڜ
fr����Vm����h�|	\#�4mD"Z��$�!���]�|�aJ�8kl�Л�a�1c[C�@|i7ϙ�A���l��Ž��c�mY�6����=p^fa0K��aJ�S:P�P���r�J����-`y>�[���Nn�7`����]�NGFR]�sRcf��?�s�A�^�M��ԣxr��K7���8���lӽ�P���e�V�P>�-���	�E��w�pꯗ�m�N�e7�ݫM��_+���::���|�oc�U��`O��r����v挷#9	�ñ���>x��[�9��~������`g�6����ﰝ�5? ��q�6̡�9Ύ�A |)�g���n�E�z}������#x�xl��'؍?�/wbE�����)�(_6�-��#�Ky|����|j��3�#n2 )�fcğ+�୲n�г�.:Cj $�V�;"�
K&2|͗�	s~�q	N߭e����ǿk������ʳ��r��Ս�D�&�`��v���e_Nҕ��Ǚ2�}z��ߨ{��2���Y�b���.wrԺ�o����B�h:��f��(Q�)�E�8"�_F-I֔/9 6�ҏ���tprJ��U, ZնKb�Ӧ�D]V�swش5	�6����o�O�.�2m�˅?mg$�9�!�Y?���L�<Á_3�S��_�	Q���K?	�6MQ����\�C��7�g�CC���ԁ����o*Z`��t�94MsQɽ,u!3���eEq",\V:1��<�֕9d+�N�}|$��#�5vi��S3����d�7|�C����yZ웒��=;���"���}�J!�AW0�0�#������������<����0���!Жڪ��4�"x�s�y2V�|��ͨ���������O�\���g�|b��S��B�9�����u8$'1BQ�..Ce{s+�-�0�W�F���J��L�Bb0���r�h��|�X�m?�`���.d�C��w��y����I��L�C�C�W��wl�fQ�~>��RF�t�}^β�_�9?�^ oS9��s6�,v,x�n�Ѿ'�Jy�]�h��c��.��1��E��0����zd��2�mͤ���Rb�ͨ��p�7���ښ:��)އ[ɏ��H�4�{����ȩ��݄8G�?h���R9��_��&
�UAG�4�
������k��?,�3�h0l�F�s1q&�����n-1����TXf>c�A"WOE�=v�`�g^�, ��"P�$�ȫ�l&x�H��@)�s�AZF9�u���M�8�9-���´SB~_>t�+N��p�PaZS�����A���� n;� К�nZ��[$� ��L�PR:
�s��KY,��vPl�d(M�k�l��ڰ��G�
9IS��m䓂����§s��=9,�r���,�/��L��}ķ����HﴚVt����� �I]���ķ��c0��B������%�ғ�6T|9j��&�r]�X����p� �`�2�f�ZZ���Z���g�?z�M�8�~�̲���� P�d��ͭ���ta��Ԩ2�XJ����������^p������s���f�Kz�w���xnǴ+T���;� ��i������{��/e50��s[��\X�P�L��So�����m>v������j|��FgA\0������D\(�X��k�[[�	t�R$�^1��g�x�Ǻ���)�w����"��5�<=�"��=��_�Lqb��d>X�d<n��12%���ĊvG�sP�&l6��6�8�r��?�t����cr(jby]ibJ��#(B�^������8�NPk�O��^��][�.3>�꼬��Id�2�&7������+E�h�t�~��6V��k{�I:�)j��@�x��6U������ ������6R+D���:����n�y%� ˝?��*hޢoc_ȟ�t�n�%��%v4w��@3��  ����R�SHns
5�����㼪@�-����^��YǍ��ت.j#�њɮ�0u�~� �#�طl����p#�s����5���6�l�bV��hRz�w���vm���H�ŨC�����l_�s�1I.�^fʮ;I������M��è����#�Z'�l�d_^H�M���3}�^�D�Td5ך�C�$I28O�猕y�̭z��I��l�o%-ݳ���6�>�ʨ��R��n�MGŜ~t��+���%�.�+�-����~*�(T��9����1�)�ՠ+��MuOr�IhQ+yI����Iz#�Ν	~?�� u����+
K¬P��%��faۑ�� J��E:/����^m2B����	��Yl���-�>r������#�<c��D�"��j#w�<#��41�3o�8D�lt�ƣ`l�>�" �QmL�9Z���ƴ_	Q G*&$;|��pX��쐤%�j�ԗ�nv����փ?�'~L���T� ����L$���%�*!b|��!*��E`o�3�x!x�	XNM7�>X�$M1���a����%�Lq�Wī~LɃ�$g��	s&���~��=���y$��+������Q��Wjꉔ6�������X��u�>LJ|U�˽Ҳh6顣u�G{��BJ���":<����)��7$�y#��[s���燮	�O�������/�;+�_���@Nq�ғza�>x,]����;�dg�� Y`���铦�	^��ߴ�/K_�Ry~�Kpj!�~�j ��"�23J��>?��xL�>�Ɔ'}y��]�V]�=��F��ެ�N�<�@s�
���r���^�^���w�i�Lj�,P�	��sB-/R`i�lI�[F������X��T�Ѹ!�@���S��B�x��/�V�
�>��� �69�Q�����xZɈE�(,������6~#S�ynC��AoɓMw��3�w�uj��5�aX=<
C�����/����4��t%'��!wK�W���ḅ$
�����W�O�u�x�=mh�"������-S$�l�����	2�_���GG"E�+!=����r�ŠV�.��f���ܕP���{"�����aX���F�Q�"@�0u��Qm���="x���^%,��HǄMЃ"}]�ħ�ւh���gU��b>��H?GE��t��f��� ��;!��6��(Vb�����u���5��޻t��NMn������X�L�t[�}���@X�/�N��ʎ������eD����2+��~
V0�)�:q��I(�,�H�\+��fZ��|dsB[�����yl ��͚�b�:I��+;/_ÀP���*��Y��L}-�0R�q�K�7��?m�pYF6�=x$����%�Ϩ�����jg��"0O.����}e ��F��NY���HnBVL�GVۀj
�:A����%�n|�������ۥ��X�b@��D4SLЄ�QUL��4wS�f*��X��D8-`L:��<oy��Dw�֕�M� �_O�a���`�������_������pq���L�&|��yyo8���E����E�m�.w��i4�b�����&�?���?j古��朰	�C?)Ggd��;�2����DX�ܶ��G6Q�$(�)jj���~��Oκ�n��vb���[b�iխn$��?���L.n-�#��S��-�$���#��PL���2s�����y��Q�f��_�iڲ���$2�a����2���up�ú��i�`���Յn:����Z@3_z�<�-<_��.�Ũ6G,���_�R���jn�	��JY�$4����A�5 �uv�+s��$�����>-���C�ո�#W�.q]W��2��������z;��hT��{��!�g���8\�U��I����4�ZN�l

��X8����v�l�J��tʼ 3�T�c�&n!0�mc�3ri&��s��m�15cq�)�D\����r��[��k�f�h��G3v<��'����e��#����q�
H6�~�C��:}J�f꬚��������,�ayI�'UMv���>F�|�JF��YB''0*
�R��+Ʃ��*J��U�;��d�F��O[�6'�Z���T�,9�C�����"]���`U�c��T�iCpF2���"��Vw9�6cmSȸj�絤�8�y\�E!awG�ip�ހ����D�H�v5g�K_������̔;�H|&U�&.�ޫh��18�[l��ƈ-� u���t��	r������X���W���
����[��-^���e�$g{���⠯R����h��U��KG��9��t>�ҥ���7�]��j��GF�Q�opv�rz��#P��M^o������e��LM�g1�d��P���R}��ߚҼ�R�ʗ��uAϊ�tc���ͺ�G����4�y'��EN�w*Q)J��� ��L��_�����vx���9�A�YN�N���8�����{s�
��GO��]U�at�gZ%%w�x� NX�`	�� ���N�N� S�0&�ԍy#�A�m5�ry��A���e�(f�$u��׸ܷ��k��C5<Md6uƐZ�J7u6|���X��;(���'(A����G��FG�] $e5�=9攬����9�� ��e<u
���Ju�~)*	h4k��U�{�d�v
C9g4F�y�`��(Fձ��d׹X�u�KӠ���^�-4���T���C��P�W��ĨovӚӦO�ѣr�z>l�c`��QdK����##�����.������N:�,�s@��9;�\�h(I�щ�M��m#'źrr�]j���2:�PpD۱{�'خͫ�>�yA�i'p�@Mb�d�L]�m��{o�n6Pu����[|�n��G�1�`�V�E��������y�ʃ[dSə�q%�6�w�,���z�W!x�����L2�9�^�0!��{����>�)C�o)��X�KPW�L�XD�������8*;�3	+��i"��I�Pҽ�����	Up0�kͿi�Od
{��t ������W(�-?(��&���A������[����7"g�DOVE�"�"�]����gh}�Z�/rZj:��:�Ĳ����V�cMx�Q+;{O�`�w�Y�Ref��(���so���+����S��?���[P��*cd��d��������t̪<?fg7l\����`�^ާ0��a���G���P�uvvp�[��`�qO����z�M.jә!T�d�>���}`�6���=&�FB��D4��&H��隌x��J��=�\�r}7�����
5F��X?��?i�����H��o��go%+p�s�hd�@#ۣH�?Ϥޏ�nV��e��6�p����}Tf��#�­�z���QE2��=�v�܌�un����,%n��k��R���8��
�����D
���U�����!�X~9�X]�\0K&�QR&'2�9��9:�h�l%��%��tӖ��y���
P�;֤
t0ӷl�N�M�bۉ�C�||$T�a�I۹��d/&�'u�F�f�n�on[KT��@ǌ�摊�wx�4�^/L<����}K�ueiu�0�A]r�̧dݝ�ӯ��j�[�"��1�j#�P���q �y�x	`��U����Q��r��1-�'$
Ng?�#'�\t�|sytY�Fe],�(�h�$X��(W�IL�i��~e\h�<׿�,Q�����F`��8D8H�`����h�$��FY��P�q�LW}����A\�͂�eɣ���|�kn;�#3�(���b�]����Q��`��D$��[��sS5�/%:���UDC�2���P�C�� 	տ���f˻����aZ�&"/
�̳S�U���Y����d9�	X����j��\�i�?O3�^�@<��k'�zN&�����3y�b�㘯�u�<�:m�E��>nb�f��]�b�������`!m{Nlcq��}��+�d��<�?N������W����5RѴ�V���g (q������U����"�	v@Z�g�JJ7�SKE�/+�8�*��V4�XL������c��E�E/t�=�F��cn�+?!�~��y!ˌ���J����b7�Q~\.�6@��~̭^p����Az�%���FB	�h��2=m(��?��$!�X1v��$%�
�Lv�ڋo:���5��d�2nS��&��a�1���i��KC��m��\A�zj�b\����g��h�����tz�� �8�x���8쿶O��@�{��Q���i�ϛ_��r*�+���0�΢��B���� ˄([!3�_1Y(waR흹F�m��>u����-:t�d�윻y,DK2I�#j�Dp�Pm<��){���� ���o��uZ3Q�$_0��ಚX*���7�Efz~����BMd�����Y��JݠF/i˼7��/��d��p��!l]���������`����s%�A�Sۙ��\^����}�1�i��_n�-{���9�g�����������q�[2�˱-�EBy�с�^ �7��0�&��#bUT:�_LA����
��P"r���)
Q�f�Ou�@1Q%p=$*��[<��?*�Q��όx�09dXI,��'M�"|�1(:�KE$�����(��b�ܦ���>�8�rŚ�61��?�f0�9�c��բҙ�6���:�����ۮ�R��;n[����ّ˭R�JVr�L;���m����w� �jwE��wHf�ZH^H^��V~��z_}�	S!���d���r��CVo5���7����#|(��Wy3ϏR��/���%���U6�Pe��ܚ��q��� E��i�R��׼_�B�I��L�W�[T��Zl��De���Xě0��>Q��g�QG�xu���]����"���5�S��S��1m�9�!�$3V�c�;L˯]>�d�~���"[�x�f-g3r�{����8QjQ��ۗ�.�B�,ד�̥�(���׏Ŝ���G4�r'��=���3��6nz�bا����- Z��.�?�Y	�%�ӥO����c��P���~(��.�E�"y�2�1�(�O�9Ե䤘�C�ʳP�N�lX_�`��Ah�5I2��l)f�g�i�Yo�8Q�A��!��*٫ �L��\�8�D.8���!�A�v���(	���ʈ�j����?d�����
ſJ(�W���O�D��jSU�o��D�ܚӎ�r$G����M\6�? �Ѧ��WB�u9m�ӈa0[��R2,��g��#Gwi�|�ܒ�o�k)�{��L��f]� d}rP���uא�,��@�2h�&�G� �������f�-��|3b�^���@���x�Qa-0�X��"<���Yv�=ς�,u��	զ����?���%��9B��&q�q�Cֳ� ��N��!7�T�_��X�l�'�vU� m��S݈Cp���b�n�G��W��r��3�p��`>������E:��&��sYN�X�\���L��t��n�aq>;}@~<�	�3Ewf�0ZW�ŉ�e�pc�|T\+V�7� !Nz�Ł�QkX��A<�G"O�f�{W	�?��)M���Mx&���<LM��@a��{*Uыy��1˧$q҇��#D���Y��'����Kz>,�Q��Zw]�&!��)F���*��-fG&n�3�m��=�u)LP��R�Z��]A@�'x>of1��vZ:מ$���^�;i�N����n�g�ᬯK�&޼U�%p@I���c�0��9m=�Q����Ɍ^n[#b��H�
'wm Ma>�f�߭6Y?�J���S5��Z:�
V2�)���WEok��b�ʴ.�P}^�h�LcQ���ЯpX�8��i-.7��r�
0��]f�P�!�)(�����9>�M�ĸ�S����N��{ �A��d}
�ћM��7͇�t��s����z5�s$���;~��l,�Q����L���D{�B+���qg�]��n�{s��oܹ�]ɀ�J����&a(֫�֕j��j��a�CVD��v:��m1}�6��P��$%��dsN�Ȉy���Å�Q@}Kd��l(�#g��i��霄��7�1@���gQ���,E6��=VY/��U�_?�c��ǖ5�n��~1��� g*��߇��ULB]���Yt����\� �0�J�ݾ�o��t�I���ˡ'|^�(���w�P�F��N`�>��C��"���^>�ʜn��crz$U;�K���9?��7ߥ�o�S��{���#C���F��+LVj����V1ɺj���`I���¯�,,2�&Uj�C�Uz3+�Pfq�q�����^�'�����`࿔�L�#�~?�t��r8��م$�@����6�hm�� ��g�:
�O	��8�CVg��0z�˺�wE po6,9,2Q@�x �^��)��H�7-�:��h�xD﹂c����vK͚v�C�Ⓝ�z3s�4��լ�Sӌ���H�Y8}����X�R�7�����Ɠ�\�+T�M	ֶl,���R�) �������
�Lܿm����x��A�� `�8����e{����\���CXx��'F�*��;,��v��/53d��x��J���qo�#���ӵ��Sbw��41��XΘ�F�i�D�7�!R7��tMo��I��>���������Rg�-t����1�PW̏����F=�H~��i$�������t�+c��������ڎ�n��x8G�s�`�X6�:�(7��Zo�$��U2�'qɟXR�H&�"���������U}d�L���&�rQ܊Ѹ4�M�	=���k�O&m�Z*���) �QOYE'.t�A����G�rǻ�z[������W��ᅲ�]�L}u倔�ܡ��,%��`IvD����ߝ�W���T��Cq]9���W�2��:t�@�y���Rş�����6U�4�y�r�D��p�������#�az*3YU��w~��Q��X^���"��+ۄ�9����yƵݐ$OӴ�_�7�]�6���f"	W��~Woӟ����e�9�o�{�X��t��Go��GZ	ΐ⑮%�(1�x"���o��	?�gH>���z���A�5}e�/�oq�A�ˎs�@�2!���3�۳���EDǎ�u��n�fv�@ծK��R��
3W|�� g��'Ƅ�_�\�?��9��]��L�5Ik��Q����d�}̛-/����?�������¹�zI��.���qd�u�5�� Y�r>�ø��)Ïj���yܐ�� �L?j���3���y���'��ÙGT�,��F���y�]�ȏ�=�i}��pR2���/R���ǚ0�J��{�*o �n�����\Oٷ��Ъ�gb�Ù���9٬v�8��}X�c�"9��;�6V��w��G��k���q	�-R�F5&�Y\�S�3 Ţ��<���;ѷb�Wm��0뷆��RU�!E��;LO�2��]Eh/��B�u@��Ⱦ[S�:��l��l���|����t�oJR�p�&1l���T`K��Q �3N��W�&B�G��X�l�g�g1������խ��q��>V��2���8"��}�fd
�,�
�qͦ�/�`����-ܹ�;��R�7\"�ԚA)���g�9�7-w�7���9/}AA42� In�ګ)P�4y�k��bc(��mlA@�̋���������؛X U%��[t=�.��h��oO�"���l���"M�:��;)pl�ͧ�Oo>�ݚe]���aկ|�/�v���"Q���� ��I7�߄i���`p<biR$!����\W	;�^9j���9_����wv����	�������Y��H-���5=�]�6Ԁ�X�����D�S�y�CG'��|���E�H��?��o(��sRR��38�ω^l8@�Hח|%�c �%xC2�+���T��~ �]�a��o5'��"H�5��d��j�W�Nt�y�'�h]n��Q��{ɳ��|v:n�6S�E!ɋC����`�VZ�m��4�.ь�	�����v��[ ��U����B1䃙������B��?����	yx^��!PdJp@C a��ѱ�
�7@S]&�D��h��|�OX�@�M t�h�v��0r ���2�p$TW>A��w1��ņ�������כ�͓*�oF�����q��4��j֚]�~�Y��U��r�P�ј"�o��>�2��$�J�;6n�]�ګ�_}��Z�,�@�٭�ԧ��>%��|@��j�?E!P�Sg[����^���46�߿:�4�L�w-*�Uvx�5��x�dզ7,uv��$M N��(���#�5���!ə��٢U�޲7��X��B����=�]Y��/-���'02x��&8��j�"(��IK.Y<�=�m3qn���{h{�f��L^�lX=�Q�Bi7�o2�	��/��Q:�l��I��Ό��q��3kg��Y�3�g����(��������E�}i�o�N�\���,t_Hf��w�|�a��]\�S'��mΤV�8}���-Y'@%��w�� ��0ǌi�N'�X� ��`�.%�XfE���D���B�=M)����)}�`#L�˂
�&>@��z�XV;�NK�w~��CͰ�҂v�F\h�5XOa������_�&f���>�[��{�6�F�m�4�8��9��H�Bi�������O��m��-��ؗ7z]ȸ��/���""��﷼]��[n�oԛm�Ȳ� c�f�����}ѥ�����0Ӌ� �Bڍ�&2�>sb��B��?n<�Ԯ�8�4�4���3 ��p}ѿ|
����'h2u?�s�yFa�o��;ͷ5�|j�YW_����$S8u`�����hY$=���N�nsף>�Pqq��/׭x{+�˟�:WROU�܏��%?4�%�ꐱ}Y�9��Ґ�����#��j��)(�,�k����G��6L-,��`8�U�_6-��9m���t���B��pL
_e(j�7 b}z��p	�1�J�_�38����u-S�Fw�k�/n���6<)m�%� ,��5Nv�6�=�'��v��Y�f���ap&x:�w9���'�у}|r���I�Z�;C�r������x$\�b݊'>�����W�"���5�ӆF���P���u�I�ax�<ə�|��/������˨��U��l�h=@ +>`�W�'L,��G��T^�Ơ�!�m������ ��h�?B2P�~�z+�tŔF_��oG(4b���"�-ϸY������VC�E��c.�.��*@?}f����{��}F���8�ɣqXd%�hX��@��o�P	�K����u�50o"�d7yX�2�\g���g���V/D�uPW�}��	��}e.�[�8j~Z���׿��}#����V��a~q)��RIA	`�z��L��6������ɇ�ͅd9Ɵ��>�X�'����煊|�/�0�9�j��t @_)�Ɂ�(�"��ָ�����x��,p���?�z[��jbom����N�y���8�z����~���G7��݄50��u
�Znr��Ģ���\/ĺ��:���!A�Ѐ�z����CJ���Y��|��-����6T�=W0J�*����b���S�p(e�N��E�7/���6�;�\���)9�$��q�$󍸋݈b�t��-3����������=,+�f���p%-��xk���z�,�+ݠ3�|�Ho�VG��bZՍ?���U��C�$�qM5�}I�}$I)���_�$A)}�0���1:�	��S͹���i|�'F����x&%�"��RNvwE*JT��EuJkJ��g�tF��]�B��9CfpQ�z���6��z�}u&qf~B�ٕPw�qR��#�axQ>y��?r���J-\�?��.*S|>4o�TkL=�.�w�^���&z���J]��Ԛ%��x���������RD���"X:Lt#~�P`v�+���I�O3G� �	������B^�N�/=���7ٚ��$�'4�k���^���H
s{�]G엠������K��<ׅU#ހ�r�#}"��`j���/�||�O��mJ%���t� x돑�A��	�J����P�2�HjD�	�>>�=�1��XU�f�����ڕ�z���,ce*9*�V�s�Ϝ�u�i:�����ZƇN��XS�I�C�ug�i�B˟{�� ��e3��=o��>����"6�_�Q��2wW5���t����Î�Ur���;��S�,��a���b�.d{��.4��>�R*�Σ��K��x���q���kvR�2Sk?���`�����8XŧWI��;���=��Q�'�0��QGǭ��x#���0�08J����(ް6�����ֳ���?V���,3����UeO3m�� a�_K ()h�{	���qE�1��:Ay�lob]~Lt���hB�L���$^���i^���0�2��S�D�ް�Dg��=UM�j�38� f��\�qd��%�a��x��V�ї�s� �I�*�hx ��5�]��ՕN����=x���Ʀ�����o����f���w_�"�bS}�I:0���x/c����:�D�'ą+�U���Ҽ���4�J_J�9<)��0ٿ��J;>We�љͪ֐*�k|�� a��w>�����+� �;��rú�υ�sŃ=�*�!�r�ʗŧr�)\�jZ%��"!o5���"T[�E�x9x�㡥,jz�)>�&�L�` }ΜF�J_P�f������A��Ĭ�����g�����.o��
��֫�B����4�c�1�{�V����x�ƮX#�yRޫw��B:V�I���w����0
[n˘�d,��y;��ܤ��o�jbD8и:��<E���J����)�/��q���_;Jw�C��߈B��{��4����9f�O�L�'Oq�0&�� &��!U�$���h;�w��p�&I�%7��V��jc�9�!�$UЗ�Mn�l*'�i*�x�n%����и�gi�M$?��N����� �j#��/��&���J-ܤ�CH��4���ω�q�Ų�1�+�'%��br����;��{]|��NI#�}�[
�&�oC�~��?}���oXͩ;n�I�������!�?��3����֙��5�zCK�1��$�Z��Մ�V��˂�R�`|٬JW��V��,���ܽ�_��>�4���Ta��o�� {��0L"�
��oMI��O���t�_"����SG��D��xI�+=�'~[a�>��h�}昅�>�����4S٠e��Q*����,.�!���&$�ֆ?j�mgrl�����dQ��;|'A-�d@��MM�r�%Ɛ

!��H\w�'�G	`Hׁ~O`��r���{ns��/\�Ȁړ3]������U�6.~���1隅�bZ4-a�6pv�Υ'��(	�#��?.�Џ�&�{�zǵ���pX�g���ϔ$����zH׶R~��[�v��$��{�[����ܑgY����P�HY۬�_��Xcd����8m4�s��6�����:/�v��ޏ��U���O.�*�N"�����G�u5| ���ԟ��Bbó1\	�Bo(/
C�I@�WP�v1w*z^���JO��C�`���ӗsu��)�^a�����
�O�՗ĬXx��!�$��k#��ٕd��$�c�43V�7����`�:.T TS� ����-��?G�5�aZ]����Q�v��
;P������(�ٜ�;��>��oj��!����t�)5%�^L�~@����f����{m�|��?�����
��|v������켋8��2@�If���-�5�y����ک&b�q�9����f����x�^�|���َlL�쭁w&y�n���O�H;�=�X���v�(���(�>0�kD�V����*�ST�&���9\�D]j�Tx�|��7��:�j�p�Y}91�>���v�z?���׶v<�|�D|�Xz����u�R�������Y�l`�w�u�ET#�
nzql�����j��+�L��@M(�g�n�r��t�ڌ��)���Д�Uv�ᄡ|ʤ_��O�l�8�뷑U�z��o��
jm×M�O���4�ʌ����"��>���#���1E/��}�@CϬcG%)<|���;�&y�f�� �}4����\_�
�/S���e�b�@�O4���c<�{ϐ\E��s��L �#��J'V(�v�b�6�^#TԟW4!bJ*mPWM�=�~�m16��4�̻^[g���JM[��_�b�d�R�Xv��L��0��-����G���1����c賷>�O����9�>!����	�&��E"�7b{*Nr��?)p�����٧��׬$�e���C�ǯ�a������?z�˥U���y^��<C��+M�05�8�v�?����M��� �['UMbj�\�	���ZT�ֳ��Y���.�ɽ�J��[��"'�W����?Ɔd�1���W�c��	k�qsdMt��t�+3�.�@��&��r�Df���I�t��8�R���VV���}H�a�j�����4�-n�m*����O[N����4��|��b�eu���!o7��he�|w����n�]���Ӵt$�R�"*�TeUc�c<U߻����!UPA��$~�A�������f���z4k�̀��
F�1�w>E5y��ϝ�� Q�VQ��J��V������Q&�$��7P��!&= H7��",��H�<��bD��
~�-[}JQ�6X��;mZڭ��T�������Y�z��9I{��MW�P^ޗJU��ڬ�fE��{����N���u��SB�xg�V��v�V���X}VrI���'����Q�-]A߆:��\ �+�Ŏ���ŧP�1e��JXT�3������A�z��0����;���r��K����7��q�[�t�,�&2�ÀXckX�4x��LP��F�jh�����Ȗ��4���H	���a�>walE�J	�RC)��dH�]鶤麄����7>��ŕ�9�N���`�֤JX��+y�i���I��6n,�u8D�8��Ğ��A���������AF�}�E����L���Ix��ç rvx#5�R�;<�Y�adh V���_�<�)g���d�g�˹�'�b��ܐ�md�K�#8B����wd4��2����w����*����^�l	U|�zx��Fb�����7�|å`�z��C]Po���D/�[�f�N�]؜��T+f���25�ɀ쟭����Ζ;g#��[����-�!�p �W���>��ǖ������ށ`�ǎ�����`С�bA�@Zj%�BJ� ����B��p?)g�-���t֜���Et����v�J��7()CK��X�NƄ��6��Wr�K�-��5���9"�*DXKJ_���P�,Ř��ӏ=�/+���򝲁�(��h����/K�0nb�P�b|vu�`"3s�u.���Ӻ�2�+4�ϕ��ܬx���#"�i��X����$,}�I!3�<<B�8��
n�"�	 o�44����j�a֠b��Q ��W:(�����Y��U0x낰�Bw)�sMl��������4MH�����c.�'��ƿ������o\���B$��T���B��Uq(����`˖b��߫��t_!ƖZ���#Hp�\S��bL��3���q3�n���@�\��mQn�g<P�B��ʳ:��0ih7����{'�c4�75��D:g}M.��4�����T/��r�/ p}�3���K~W�r�C��!�yf��L����Δ��%�}ev� �O�-��Œ������� X�r��뀁b?t��ن���xr��H�E.kA j2�\�۔�㮵}�Ԫ���M�����L��eU_�w��q�"�����G;�aF�s�4��zx�,�_��s?��:\�s|�K�P����:6��jK�UqrlY��0����^��؜Y��?V"��5�'���6�S*��lD�	�voA��z�v�~�ϗi�9�_��^��c���\�M�_��UYh ������^�C0v�	���9t���F��5�.=mҗ�d�9o�#B��C�]�c�L���S-j�c�.۔u�Z@u0�G����nf,Z/��cɑim�����X��G��o��T��x�T�^ܼCI�ߖ� >��ԥw�u�!�S�<��9<����}&BR�7ҨY�ȩ�8}C-�����AΕy��`�0*0ct[)��,���7��F�)�न�(_���/� D����^̱BE�v�e��d�h����	�T�$�>��ܓ�9��ٞ�zO�U�����x�XW?D!��F)SҶ���Ӷ<���pH��\p�X��׸��W�!�m�� It���pH�xG3?�V�<*OfH��!+��%Yg�0Y+��B��3���t�O���OI=T�0�ҽ�j��}d[���$���ӿ��"T0#���9��~/Qs7����������<�D�y�l��HM*�L�7ufƅ�O��U��E�!xs�F��)f�1����^��n�hz�I!U��T��Go�d]�Bk��q��f�l��A@�oZ������n6a�%A�E���u��~}����L=��ײ���Ӭ���}�D�Sdk̏Ѷk��Hʺ����ڃ�f�Ǌ��@��}m���^�b��6(��89��%p�\	傢���F��I��K��rh�#a������eˁ��kZ��,�-N�He�o�~�#��
��ihJرQ��L�z�ܷ��B��m=>� ����6]�'�-�$~��%��E�{��+��ZdE_�%Rͻ*$�6c:d�^�������27�|��V�u�����0��I�F�G�ƃ��l/VD���6���A�4T�Uס\O;�R��`�H1�Y��f6���-�TG� '��������i�sI�ޡT�{b`V���a{���ϋI�������P#�je�&�K���$G���_��bA����IU�ہ>��Z�U�2X��S�7L�2��D_�	��E� a�پ��ԗ���?���o�9�0��g�M�%�"gWYM�C�����3�FkZ9$ּ�&k���_v(n�J���
�?����q��|�!ϋ���[�Z�ݩ�CG�ר%�4��n�wV����]�}Y�48�9@��IVD��N��7��~>���'����j�W��h�.)�X�JQ�����o�nҞ</�:��v�"ŢQ��X�ׄ�N	M��R��<���G-B01,؃�
�'���d�O�khҎ.9���.L3��I2s��Zz��L������p��b����p�n����
��DW�� t�ᒒ�+ݿ(�o8﹕'�JM��~A��W�sE�^�B$@�р�w뚯����Ķ�LҰ$�!H� ���E�~�vAW��I��4�Sp=!�ا�6VL��3O������:��CR5c��[�w1�l"�A��w�(�
nbzI�������D��؄�����������
1�*�9�P����n�@cv�$;چ��A �b(�5搧�6�l��Q�eQ��cd������P�;�8\�P��)�e6zu�+��l�ywr�S斷�g�\�8/U-���M�0'p>�ѧ�����	jOpP]�G|�&�2�@E��s���o�˘`�<?��c~3�δ��rJ�˳ё�Lp}���9 ��Di��t�A�d�.�dm~@I�E�5�Y34����)��H��ĩ��R�	ֿ]@�/��My�n�{�{%|1-a�-���UNmG�̿"�-ء�Q���vO�k�Ț�O���v�K
u_t�k�hJ�]OcZ�-iw֮Z#��C�}*y85��S�[xw�Q�a�d�s��E�Ҥ���2)���Fv�ì����O���C�q�R��N|���V�i�dw"��9��ER�W���k�u�,c�~@�	Ln���뢅�z�G�Q�˄�&e\�e��u��d����	�`�U,�	yw��n�qeș�����{(��$>�ո(�]}��VΊ�f��5v���)���f����	��a��%���Z��ѥ/p�j�4�ǲ�3^Q�:u�5��M]�����y*��ui��M)�}��/���:��fO+[��[�t�a�b����ȿk`�~!=Ѯ9gJ$��a���C6�e�����F�����s��2��?7���y�2��N�$�����RL:�m����`�4A��!�P�9�N*��!w`3���9�/�W�p�����J'9-�L����<���g ��ǊOK�\��a㘖n�f֘�6�6|,��y�h������!y�<u+�~��ׂ$ﻇ0G|�Ί�!��UkR߀���߅�Ζw0��w ���|��$>8B�b�מ��z^��c̑TR��L�4��'o{��0��uij��UɘDW�+
=��Xy�9:��aKR�hZ����xqT�md7ߗB���"y�^[I;d�A�5H@�%�d��S0}n]�N�D8l�5�� �rO�$w!ab��k��8�����SK��g�*s���� �鐦�m�w�|==�6h�_b.�P����<~��5�)�Ɔ�3bu�&j�t|�~B�l%��0KLC��X��t��,�B--S톽���o/��TS"JA���6p|�k&�)��!�Jj����X�[Aז.I4<�"m�J`��'t/�03����\�����������o
�o�0��~S�`��Y���ݣt~p�OlH��g�48���~Q��
�**IU3XDUw��V���ZZ#�x������*�Cg��,�45v����Y���>�go4im�/]�Fs���N���W�u�CI(��t��� ںh�9oᾼ3����.��5�Yo6p&Y6FoQ�յh�()��4u�vkfpV�I"p��D��T�7@]�����|F�6q��9yb_`���PkDK�؇|�P�J9��v[>�u�g�:@u��t�����R�yRR��IY��ۄ����	-+�+O�<p�� YcP��_7b�[�*�ރֱ��|���_��MǐP#�RV�r/2����K�0�N����v5��|�vif4;��aaȄA���z"���RԴ�@�PY���d���R�$wƘz���2�$����OL���@�U`�_ꮏ����|#(����\���2@2�ya]�6\��M Au��|,�V�B9g1�Y'>@������ &�!��-�<吤ߖ��4��~^�:��̈���}�nϞ��Lw��wv��gY���^xJ��f9w=�{-C܈�s��dU���qaG������r�z+�"իa5�a\�.���?.X54+����za+����)�T"���$a�%[r粿��������1�I���l����ُS����v��b,�/B���\��Czj��z��M�tc7��M�]�mA�$�p%�R��+����A�Ê���{8h����7$xP���3��=���e���b�Q�3�Z��WU)
￵��|���-@�%G�*�{�y���M�So��f۞X�4�=�� jjI��F@]��I�۪����J����2��l�8�)բ���7q$ �� #�XE���*�|�� ��ӺD~V	�eW�RW��f�q�S@�З)�-�ۧ�P**b�ż:��5��8 ;�G, gh�jgl}L�Z��[(�]~����[����
H�2fz�|Q�`�0 �KB�̨�ke���H9)̈́�&F�4�"�o�6-�>Ju����c����1��g��65t�A���1$�������1�����&��ܸ��(�W-�f�:�