��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0�����(�_?V~��
�r�-��i�`�oD*Av�a��*��c��A֫~�K�l�R��U.l�ȫr&�|ހ�Ҳ�XI�yD�)�����aP,��'}�D��r6+u�5���C��H�zx�?�(�hr���$G��t.���t��O�"�j(L���7@P�D�ML�M��4�~�%S��C0v �
��:i4Q�K�Tҡ��`
�=�d�fs"���4�.0]U
W�yPwb�1ðt�ީ'�<�Z?���@3jeNF���K\�����P@,/�<"�3U1;M�@�	i� ?%�<^1JE���!a^�=Z�P�_�ݾ�L�yoH�iX�z��h�9��
��HT{����ģ��m�>YU@ߤ�����׎SZP Ψ�?KP� Nu�����{��N��s��R����:gO{X��ɷ_���e���Tv��5��V��u��kaK�����6;x�B�� �[�k�6e]Ķy��ӹ�4b�E\&T� �`#.�Ʀs�i�5���u��m�٫g���K�f�թ�U�G ��&���u&g��d
I}��D�Re7�I�F��C̲�tIA�s"��M�=z-���Ϥ��1+0��X}]�1�0��mx]���1����D�4^����b��^|gR$"�C�@����~�n�૴_EH۹9V��u��ҁ�%�q�tp"�fML�ā��B��
�tFZ�4ڎ����x# v�g�K�,53�5����f>��	y��G�N��T H�#�~�T��~�_9��`Ǜ*i�"8Й�5��1\pBQq
m5��&}B�=[O��P�DM��{�d�o�g�d'.C���WU% 0�iِ�	�~;�M�r���u-
X��⁯�/�p�5��Pp�t�?u|����2��g��MN���p�;+\��z��j��m�0��F��(�Y��ܷ� ܿ��D��`����.�&���F\׺Ƨ)\ �L`Ӱ�ŀ(���wvn��@�0kĶ�p1LV�0,bLFʗ<�����=��м���/\2���
�}���AuEfZUs�����)�F�t7o��n0P����:�$��@,��<Qn0>T崒��s#G:p��1����I=/�2\�^�]�C%aJ`v�3��9�#�'�d�/�ts={�6�W�g�b9��ͬ�d�}|f�!�)K\��Wox�p���je�捞t�>��.����W[�A{:�0�p'��&ҪJw4�Na���ݺAgb���U`,�aE��fRO#���) QE�f�c|�˙+��롥�N�1��9�y�<�n}mz*��ˌ���3w���@�����~�W�/H�T;�VR@\C��x�'�ن0Lc���VOL#�-�TW|\�~�S{�F;e'Y��i��0G�S,œ܏�ܑ�&f�t.f��A>xU
�`����Fg<dI�*���9(�=�L�ɭ�q6�(�u~�x���B��K��Trg̭�g��<������g�X�Y(������<zP�� �c�l�0jA��}�K�� C����J�x_��8�f�\V	B�2iQ��]�W��u	����F*;ُaO�={���]<���ػ�f�����(T�	�\󜲇nTm	����Ȋ1֊gaj�}��Ҟ�| �&�E�/t��<��LT���K�w��|-�	?�d�;�5�܎r}eҐ�Tm���R�W��q�������p�}��a�-|�<�4tŷ�"� �����I��/������S|��a���"�_��$��fG�m2a�;/�g�Ϩ�>/����o�X�r~@'�~Mp�5��̦I�"w"�6a�W�%�Ȏ�h��+�]�Y��h���=v�������3�����,8T�������3��ںF�����
��H�o���� e��ǒ+B�s��d�8�k�����P��B{g��0�ކZ?PՖ�h��x���NI�s��>���^O1A�L��M����>��b��:�J��*���1�I��Ax�|�;���Ktյ+J�$.��ڴ��f�v�l���:��B����L��JN�����XiD�g��ؕ����pZ�zc�������K�����~w������Ġ����K5t�?Ф���qv�;`������-�m!��H�������R��e�:��2�>f��/���xR�WQ��� ;D��U�sGò�cē��5�&�p5���A�-��i����D*g��{�Q�#<�	p@h�����o���5_%�Ί}����n���Wy��� BB(�M��"EE�+�T,���AQ����`M��Gl�Y��4W��dXӟ�#֛?�C�{t���[���<���e�+����6�}P�(�Y0���A�lؗ)u��yϦp}IS��� Ҷ&^C�ɮϏ1SW��է��@�����4K>lK�w���	ץ�B�D�M]#	���	X|%@�=I{�ْSk�MT��ҏ�5֏���KΐXL.�k)�j�b���4Gu�WZ�)h�U�� 8=���Y�=;m�@~!�˰!�y���a%T�w'q�u�������&��4E�wE�{"^�����9�.��J���C�~UYZ�d�-r~��V�#�dpf9Mwד�;(���T�)L��7����C�a{�ka~H�߽�L� T�Yx[t*�Ϡ��7�Ę~=u8����۶C�e���B�nE]���b�yK2��'4p��I��r��R��;Z�ɡ�Y�e0������l��!