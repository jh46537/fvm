��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\�#��t"�9���!��� �h�
���ɀZ�l��\�����o�P�V �(,�=�`�Ce�t=�b�؛Y���ft�^�VHͽ)� �<��9��q	J�$��r.q{.+��!q*�Y��u��bk"nܫR���� �p.V��&���:ǐ����r�'B���iE^6W�z �W��lj��-j�'�,g����ג��ٜ�����#��33y-~}�6-� T;}VۮdQS�"�wd��|�E��]���'�AGz�Cgh�����i����|I�?:S#����E�����˲�_a����"�X�8���_ke�RB5���c#����.1�odO�33������OK3UQ��G�?��ˍ
�a��_�����=��0�j�I���Ya��|��^�3��x!��tj���(R${���iXᨗ���KOP/�l\1���s�6��ula����e�9�ؙ4%��A핟�ЩC�?#S�ZXH6�e�U�����E9���~����F�b��H�/[E�P?Tc��1��j���#7m�y{'{ʯ^����?f����GV
S�
=�W���D[�H�q��=�Sw7-'�w*ur�Z�nn�Pό^.L8\H\'���� d�F1�v��T)C'�fh��ݙ�����N�V���[��-!-�E�4�aFY�i����oqӃ���?-\t���h�oLVv��[���?[��%�@~���Lћ�P�C�|oQ�$��������AX|p9�����Q ��[6AA!�SGJ�
\��#��b[|���Ԕn�B����nC1��z�{U�X	�8��Ɛޖ~�����\;����P���2Ț��x�,�����c������n%��b�঄�ч�*�ꊞ��xɾ��Iƍ����CP�x�1p��e=y�ҝY
���:Ñ�qK,<�p#�λx8�t�v�؄F5 6 ��)Ob�Bz��-MԋL��S	>8�'��G�_��<ė9��xNdoڞ�B����U������n�����T��w�s.�����p+��
��4q�c�|	�'���RW�9FTX���X�=���P6���!��+��*`N#��nvR���M�}l1	���Ӧ����]���9]����tL�,ư��??�G �R�Z&�%H
�>oxV�So��}v���c�$�M5��v�O��� �=���C�� <���D#�ҔJ+3��gMY��3��YĹc����}�w*�%��,FeÍ:�s|l�K��/�0>3�[�܎F�dM����E!|UlЋݎޜ�e���I;
�^�Y=<�_N��q֥��D��A.���f5*R��d��YWBP����>�1�bF�.{5!���Q6o�=��`�;T�Y݁铔����x?��@��S��H1��dz_���{��'��x԰�8\
*��LzD� w��|��:ُ��K��L�&�M�S�0����iZ��ّye��[
<�ޅ�d"�����z�V�0�L��Y����ܹeM��(�(�l=����͖i���L2d&p7�m�Z�K����H��z���} N_�^�R{�.��Txx�	7�t:���A�5���t|&�XZܩ�@z)n��1�vw��~���g��}׀�Ԅ�\ً��+�{��מ�I]�C�'E&��Up-֊[_��_t��u�v�*I�輥[6��������!��1���Cc�*���*�?�{dP����(�?i}MHf/�F˪m.�e�<���z�]m�]\�wX��?�� �Jn�f�^����&����#e?VE|I��݁�"�pN{TJj^cKGL��)�ʹ���A�wϳX�Л�
��H
�}i䅟��O}�7��vn�\"�k1���N̮���J�'�/�nQ�4B�r$�s�Lԕ�X(�;Ց0Ǭ�-���N����E
��-�E�#�m�w��:P� Q)���\����f�e�i�oA��VsJ�}�\�����"��&"Re��qH��zmT������x�#W
{g�܈5P�c�`��;O�(D\��\�c��u�ghbf?ߍ��t�N
���c����)��c��!��T9	;��:�+��-{�&�:�S���������M3d��h��ڧErT�䠦Qo�!$k�U�F�.�@Dd������ �{�����;��!34��K����ۊ��XH�q��W�Ui�λ��,�Hpf��������#>�㪜e>e8iR�Ӑ�P-�O|e1���p�7��k�(�Ч���a��\j
�0�H��M)��`Vf����c��U�����؇��<�gVE)��T����':����e sӋB�v��X.��L���\������4˓���i�=�1Q����F�mр�1��]���4P�*��9�K
`��]�SSE���%ࣷ?���*�?�Ƨx̻��mX�[���HXU�V����[*Z?p2h̅N@��,GXO��UF;�a����e�r	�z,SS[2�-��{��-Ň��_����WZ�jc��\���fƠl���9�,?P$ �	��6u���D�4��L݂�6FV׭g����x8�?��#�g�X�C�����(>��!Wj�[zK�����Mk ]�"a�є*��Ø}�SY���NCQ�
{[�x�:ܣ��U�f�woوnQ�)-L�������	�b8C�'8���+Uq]-KK� ��7].�U�j�&�J~<����$Ȯ/D��G�(��xLbK������C���b�?v	���yc*�h�ɶ�m߸�7Bx�F�7�%�lc����~>�X��H���U�Hb�Ǟs����zK��o���j��}��]���XI����ͅv\r�jzS�I���yհ(��i@�Y ��Fw�EӠ���.���2l�nHV߀j#0�i$ͼ�r|r_�J�r�MO4J+ ���Ɇ��YYM�5���H�ՑG<6Ȧ2�;C�f�iͥ:��I��`ܯ�g�#�z ����|O�-_F��ޑJ?|L�$���i<���g}3�x���E?W��p��者M2��J���i)C쫑[\v[>[b2�i�_��bA�z��p��P�nbc��:���xT\'��J��w�����S�:uo!a4���x)f��JЈ�	3S����$��M�'u�1�P��2����JH����@�_��#6ޱЬR��r2���'���ld��� ����U��;T�5tz1�^`Z��^��3�<�F�˛"n�E�C�����()62�>����-��o

 �A�<�X<�1H�p�^�6R�Th`���� ~�j���QԿO�X9"df��Z�Qf#y�D�qp.�+�N��g���Tү��C}AN��?������1Km��U��Bo*V�`�1R֒�[���w��%.�D6�� Y�ig���M5QP�֣�9�Ā�Z�H�2�6u鶏�
�].�K�{3b���`�f��o\�=�����F܉4:��7Q��S�	P?R��i�G!d��Ts�d��f�cf�ֿ���)�o�m����g��b`n�gZ����?���
��5�Quh܆N@�j��Q[�k����#�>�c�G���IA�/�=<��Y��?��?��*ߛr~SM7ÎG�@�}�
��o��צ�m��2�u�N��2�J�dYW�A�xaz�d�˂�P�28z4�:	�хI�%�7}l��Gޘר��ŗR��)����;�ܢ�b�\|T��z�S�ȉ[�(��Y�ޜhDe���[�0VGT�����jҺ�N6�R�����Gn���"����z?M
�52�]o�P����:��n1���.�GC�0=pUT�X��݂����5Fކ)�6M�&�W��!_A�$����@�2[�+�=��`�%��[G�Ou�J�9��o��L�x'>�w`	;�a���e�X��{1��
3#)sUXl*Ҷ1':������Zņ�=��]��&|�����)���h
3����u��A�
 �R^�� ,��
ĉ�gI�"�b� y3.����y	�[L�J�� n	-/!���������U����8����qp�Ŋ��`��2�X��aK)�=	�<���<������S:�-E��_���F�<\4��"	F�%{4������j�tɺauv����`Ht�Eڭ���|QHG�.�U���w2�n�4�9�v7g;d���}h�9#I��#��hX�ͮZ?�j��ʞ�V�㔊�S�u� �QL�*����ē/�%��"����N��� �H3r�;K�BCb"
�J�	��2��1�e��g����'�V�S��5Ixy��|2a�t�_���:��È�K�ʌG���j�W�Z��⎦�>���*�^[-O�|(������{�?י@�'�o����pI�J�_����v��9��.�~�-�i�Y�-�1Ѯ�v����:	�y��^L���1R�V��<�I$l0��;bL��� ��S�	�����{��G�d�1��V)�C��YU
��\:�W
��S�H����U~Nr���4���͢�Ԟ���s�a��^��dA��黖�ť��^�9ѫ�L�i���Ҟ��uH
+���R~)�c�S޻�2v0����>�}��o�Cwq��w��T��L�%B����,�~�������'�9ظ���Ҧ��������*T4��Koq-�;Hl��}�Ҭۄ��G�y�RE_�V���6�E�؃�g�9Z`����S�a�>F��J��	v�)��BN���9�!�����`^A���'��/sJ��;�D`��qg��MR˭9c��q��ך$m��s�.���|�U���PCz�#��@:��.4˧�Jq���|�[$phX�X����^ט�"�������C�
`��:���S�9�DT�,7.��> �D�ȧL[9�"�ֲ 0;��sՋ`\�"�X���:�,�F}�z4 �XGyV`64�[%�ĸ;b.7��̋�a�ؖ�e�F�5Ӈ�,��J��1�=Pܸ�c\+�,���Z�-����MY�/m� ��V��'����q��/�<���Nk��Ε�*��Q%�y��z�W�G�h��H�;1�ry&<ݫ�C7�U��=w�hV�hQA*�~��3p;�