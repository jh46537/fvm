��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&hs���τ1��E�"a�;�V�"��k#"U������P���\.4!pں�L$�u6�����90�G����w��-� K����Ί`���K�`����F$GkT����ͷ�����w�@?�x�)�F�MV�+�8��6}\e�_����$è�����=9�7$H�i+�Y��H�����x�Fw�M 1��Q���-���/n��#�����> �9d�m����C蘂�@ޑ���0�b|��мj�Pb�� jk�SaR�4�:���6a���1�*S�5Dh$��=#lЦ(����������A�t/+:v�5���d|��*�>����v]b��AI�r��,g0����)��BYe�
+=q�����Ӂ�
f=�e�0T��$�z��,q/����V_NH�RKPz��bi44H�H�E{�וS�hq��(D3�F�.=�K�_��9;C8�Sh�\���<�<���Ӎ��n��0�;���f ���B��C^�Uk,p��]8M�5&�'0z������Ui:��������{D�U�>@t�<��m����Id;&�g��r������x]Z�F�/��'#���b���<�����ի��&�������oV���vܘz�',�r�䔦eSh3��/v���2+v�5bz�=�1�����m7�,�6������:�!�þ>�:8P�	��Ծ6�Zo�X&��6)�p��88�|[�#��7ά<f"j��cR�b�6�6m��Z.�3mm���V'�ԩ$Q;��Z��c�&}^\ݞ3�2��~v��Q^@*j��HH���V��,]�4��H��\��d/e4���,�H3�g�RW�^��d��z,���r%Q��j��wF4f�6x&0�����AtDTro<�2�7��6(�tʺnE�LY���b`��%D1�� U����G�1�j�Z�Z��.�V�8U|���G<�j��@7ӵq�<�O௼c�2,�����:��w�x�Żr=��)!�����a�I�i8�༯BE<6Ȅ���ѡ��lBn6�3����W@QG���2,��߆{a��4>O|9��̅����,1\C�VY��q��o<H�:�|yD�O|f!��3���^��/8XW�gme�6���O>kٵݣ&�nbF)>MN%�4j�o������Ĉ?���$�(m�)��>���c���[�(9Є�Al._AHہ�^	�� �=�氶iK�uDZ���r)�e�NB�c4L�jIw}l����6"�h'�bm�Qm�*�$�B1:5|���=י�j��:ىM��p�IW�lzt�x����%�Y�����G.q�Tih@��<�'�PLی "�p���rv��3Y�/ﴝ�-�ʌ���!��T5�qL��3���Ȅ�y봵�h�|wdNO	�w�h����J���ǥ���ȼ2����Չk�'�J`'�ƈ��.z�M,�����Z��m{������LaNQ-f���ʿ�����3&or`�������t�8�q�޵���k����B	�,h�do�\��)��%aaL*NV���r�K�!�_(BwB����|;`鄕y�22e�Z���7����}�w��*⚣L��7�n�Y��SʈUcગ����-o}��2�|~��?��ߩv�B� d=�2��&0���hL$�T���J��1Кl���'��@2��3_�;�����u���u>�<C�M�}B�=��3���=gWi�s�����Q����; *����h>~�>�\0�����,>
�%$�c=k�_"�)�C�-E ��� h<��-ж��Y�0Xz�!��`,23�9Ġ��yH�T���'��I(����~Fr݃~��;�v��l�г�$�v�,����Q��.̡(W�N����7&�C��5�M��%s#a͡����v�_�Ey|0���'"e�a��r�P�~g6�g��/Y�x���	�� a$�9մH$F��l.�[��Q����B���u�6eNs�\��K-���y��E"�B+,�j@E�m��a���$��<_[�]?��u�8��SA����e����[EY�JC�Qr�P��w����W��y�
�{k�qh}W��>W��T��'ۯ���ٰ��nyql{�M�$ ?H��=\QYG�%�T����m��F�pwnO9[wՃhi9u������I��y�E6��d���%���?�R���qN��M��Z��^�\�r�z 52p��vRD��]�: '���P����s(	>P
{ۢ�ň.��J!����ufx.܅=�DT�3���	��I֍�^�b>��o�'�ڋ	F_���^!�|�Rf�i5�O@�yܠ��^�9Z����jHS�l���$��ϖ�����fp$gg=�+�R���C��݅CL�u}6����'<^���_��s��iƛ��8�C���zn��V��M|�JmSCd��U<kK\��,s�U�Oǐ����vv]�Xr!��
:���E��I�g�������7kf\x�߭o��]7���`dX��9N)�t~�6�6������!�[�&G�W�����r��sz��<`��b�I�"R���̀���*�-��RtA_f%>J��^PǜP����n��)ǅ�S	k����#F��9-��ٵ�(t��c����'_m{��-~����8ֈ-��D�扰}�B�v�K.��&+��5;��{"\�W�^ȡ�x���m���`�o��w�՟'"�iz6۔:�b�
�p�F�@��8-���2nt�� �D~��y܉㣵-���T����/#�r�F����x)}4�'0�y�P��\
yS��YI�zƏK}ց!�oZ�OZP�w�n�&T�Sm`~�ԋtN4��C��ԃ�f��!zǒ���[
���ǭ��bi���˥K��}�Ty�zr]�c�BA�~����b)*JX�4�$��㱏��̆H��"3M� �׶��7u�����.��ʜ~/�r���`�ȑX>W[�d&WP����S>�M�.�S	.��v��?>���rJ�؈�[���chk�ѐM����=ҁ?d>�8�]�Z�o��v9�֖3��H} �U����?T�fU��Y�w�;�ŉZ��-ک#�O�3UZ��\�/k/��˦x�t�yI|�=f�1C����!,����G˪9�p1U��~�G$�0�B�6��If�kl���q���Of&^�&mo��@�H�mGH0\B]_*�6�U��Ș�}���l;��4O��!���Ί�)��PM�}MVM���@�
�b���p�:�xI�t-�̳�R���/\K��d}�`<�~B��*#gO�_�#xy�jN�bX��*ǚ�_�,�D�#�g7���d_��<�?����+��h��cd0��{��Ў\�R�����Z.����{�p�+��Y�tC4�Ic�<�mQ�bn�v�����$�����Xu-�.�C�hf���u����i%*�K�n�0��_��D��Y�;%�4��ES�W�5�Rq�t�Jٶ��l�� ���l3�"u���^���Z��$	��@�뺳�E��K�w�Q)�Ua�o��1��3L�gS{��ʶ�9,'�q�ʵ��e>kNK���&��KڒAN^ tI�Og�\}��>( 7�a���S�>�h������/��6n#�v�p_�Ì�3���獪�|���+�������ϫ�|�؊_�fU4�T�`g#4ⶼs�fϻb���ؗ��Y��	�Vfv���>a�������A}"��NF� ����	3��� �_fkՌ~��8}p���'��-y�������7�6??���lxV'�φ
FK��3G�S@	�ΝA�,������ǜU]h�ʄ?8�I�xS�rG�ltb���=Q�G�����%3���&�7#`9�s��Y?:��D]�O��d�Ck��g r��hJ�~?�R���o����e^'��xpb�-������(+8��P�5w�z��q�k��L��^��R�y�7#��~8�:h[n�'�:���Q�����i�\�m��U�������ve��?��:���+�#��f��%(�;��;N!���!Ys4���-�M,c�	�g���a���2��<bv�A73{�	�'�a�VW��) Yd��:��Tx&�\c�=G���
˝|���k����1T��>�XR��1yUnY��v����MAfut����]�Oy�pWVQ�dhn���i�a�B�lJ00]T�U]�m��-�FX�ܡ)��Y�u�B��V�����P5��7J�T����)���>���¹��я/u6��_����ۡ�v>$�ȷ{�7l���[�c72��� �n]A8�����Mf��&�~TZ���*��e�C��@ ;��nH�\�\��W_�0�׶����F�n�.6x����j��Q=�T/��l���u��"P!݌�\	3Ec|�}�U����7�A�o�Hy]�#ǂ�%�q�����s_T��W��V�.��a�2}2 S�(�%�2��2+�� RgD�A?��������)́�k�Y�i���>F%A�(��F�|��E��t�,���@)]��_�X)�;�|0���؞�N���NXd�J4��z�����ol�x^��|�+�2.D���_�����F��p��/�1��
'����(u�
��T<Qx|Ù�-N�W���� 1����U�jr�Cd%׿6�A����ls��D�l�F�G�I�V���gz��89($�X�z"o4���/u�.
�Tv��Y�	|��L,B�E�O��FҨZ��欳��5�<��V�4%^6����M8����}v�BP.�L_S:{VcyY�PN�ۃ7��@\ ��#��q ��h
&S�eV�0^�>�t��k�ָ��J��Aa"8���}��{~�u7V_[�e��V�����9���`���0;���2-���2Y�:��?Χ?�i��T7�W]l�F��S0�P��1s��?��':O�v�A�����"bZ�}Fz
�=�y*ۍzC��T8���º�/jdL%y��5��^Qν2�+�c��<�*��-/�yH-g�/�g.��t�ձ{��|�i�l�5��.�N�0�a�<�\��4tXPvHh��X~͛&:���
	k�#�����P�c�p��>y!��Ź���"0����� ��I|{b��Ce?�J�Y��ϕ8nh�M1t*UOnV�<�#�g~f������¥ߙ��_յ��]j���JJ���;潠�-`y2���������s�#(s�+�[�(,���p��Z��=(#eՄ_�{�ҞwF�^ekE�5�.x����e[́C!1҈�P/{ 7��V�p̐��%J~D_h<Ӊ$_�"��^-P�g�<�JGRK,'�xw����T�kq>���d�F�Ƭ�U�'������3��*�{�[�&��;L�\Z�͔hWA�{�&c[��,�+}�4'�lv��>��xK�:G�����_�%���$��]*��Q��`��f��-94x�3�����QC�g���lN|��)+{�Q:Y�-SK8c���E��|r�i��gˉ��ј�A�{��	�< �*� tŔX�����5e���UN��x��+wV��=Ǣ�i=P��+/C���	�f�4]�.
�9�4����ڿ���o���ߔ�:����P��LdM[tM�G�ӸS�uZ�v��0�b��`�=3<��[��ȴdV��]����*�hwf
V�/��%G�Y�Jf�9KT���u�f��.�4\mqQ_`�*�Oi�.
�!{�Ĉr��Ս�҅��~1~��)���~�N������BD��|�x���C��ȗ��i7���3�Í��Y��o�|�;�<�r��+�T�=-��ڹ̈́��ܾ�{��D��d n�i\�<}b����\�a��:\>Hކ3�h#�N�\i�f5���opr����&6�s��6�K�~*��NH�/z���).��I���-�mǫ����Jh����	�Ab<AM���s�y1z���b)��<���Z��H�y��rz��♨�RO�	�ia2��&@�^�zʠՆE�:O����tv�f^&2��o��	����t�s�< C��t��H/�/����/HGz?Fg�X奖)a�2��l��k��ۜ�u����Â"������@^_�@��ԒH�'�)�Ҳ�^��s������1��:/p���KoJ��f����IϏ�1?�
����j�a�����v� >���?��k�擁����(Y�XJ,�.��sj�`"q�Q�A������*��� ��ّ�t��F?�d���kVDW���F ���TK g����hm��k����.�-��6��6���0�X��,���E���6gz����@? �{�\Ȭ{K'��mn���"&d���U��_���s��`��� 8�Ҝ ���7M0��)�8�X�$_�*8Z�u_�����b��V�Q!��f�߾ʭkCp;W�u���D����� +�ZY&��[�xH6����`�P�
��h%ǎ�9���C�>��X�Z�@�NG���Y�qW˳cL<߰��˽���k�y���t(_��W
R�o	L�ڡ�6�LO�]��p�i��w�X����''��~�
�b���i� nZ��!ǿ���8���U����M��q̣A&�#m��?��Z��՚�YϚs��%� �(����d�g��~�����C��oOE����H�FK�T*r�Yh��	�!��)Z�����D�d�P/�q]��ڢ��Z3H�x0�7=J�:��~�c��#�,��S<r�$��SXR?��̩i��U��-L��E;����E���n7N��kTΝD��DyV�; 3����!���H��{cMl���A�(Q�"�"^NU�N���/���@�tQD=�b�=t��t�ȿH� V6�X���!JA�H�k��\b�g��x�Ř�,l��ɴII��uc����]�:��|K�#��:�����9��u'�TLq���HI�`�ܫ[��2>��~�G�T�^��-��
�yAүM*;Θ�rF�����a(�J�a.n��!�wS��|�3g֌)8�S�6�j���Z�fhڥ�����t�
�ǐr�L������|�![�D���^�XM�b��@���|�5�+�9��%�s	��uvv;����7<y"���xv2�}��b:�V�G]k�k���+��x�X����T�\���	�����Uy6���I* 
b�Kp,�4(��o�)~$���q)��T�=�ǋ�?*��:�U���^� �V��n�P�
�?5�7�E<|w�4w�:�x*��D��u�ι��T�X2���Z���`�ָ��������y(�=ؚ�hC�n>�,y'�ۆ^�g�G=đ�TS鶮�UmӬDvn2K���ۄ��+$��3Y:�e!�ޥ��������%���ח��reu�>���;X-8Z���>��;��d�D�z�|8��ɕyaԹI�*E�>�3��no�5ἓ0�%���˨�2
}�g3Ӈ\���|S�u��l�;o���J1Kx���(�~�"��(E��J1$+sC=����_���\!h�_��İ��#�(e�_L�Ú;��3?'7��-��fE(����+wn Va7Zn��:�!�j�\�e�(ʙ���F}z��'�AA��`O���z��W]�%_�3⡗%(FŲR�Q�)�zx�'�����p�*�L���b��
f������+�bI�if��[QJCCk�!eߐv�,!=����x�'~�>����ː�"%^�Y(&��e��җ�Ȕ�r�B��/��"��_��>����P���Dm�2o�����i��-�1?g��
i�,܏��4	_�,)'��L.j�.�h��f"v�Asz�&bs���D��"���rUO�uI���@��.�m��?�)T@UD��K(�u���3�ɫcW����p+U����Mŋ9�YJ�*F���� W�:���/�A D
a ���9�jmY8pf�dbKu�`zO2��&�hT��DML�"j���#�$sf�7-Zz�a�����]�J�𽄒<|��/����%rБ��LHJfP���
���3�r�<��}{t��u�ٰQT[�����;����i+���dc��o��@�O���-
զ8d%^�Ǽ{+��[�a�Hf�	㹞f�wq���p�9Ys�IT���Uj͘q�f��w���r�~�_"�[����w�٤��F�X�AӾ���υ#����]W�FZ���U ��w���5xAW�)ۑ��Q�/����~2cFsk�`ۦ����7[�r�e��vA<1��0��d����=TL?����3�h����P�`;�l�|�EX��i�k�:2�	Ym���0ȬKҭ���&s@:�}�b���iQ�-âW�)�pt.�������DF]��,�������[��C��p$�������G����털��-�8���>Q�3�x������Z���g@�>gV�]�Mo����p~wl�Éy�Fu7N[s3�����97�Խ�y3�� !T?R��v�O��~LЯn�
y����[�L�k%{��.g�Q"R@k�1�y�2��������+-�},�境rҒ�OE|��sz��I��*t�}���Ci��Yꪸ6�<�k�"A�Ћ��U�rt�Y�����8v@P,���-Xv��{�ˢ{ɷ$�)�c�>x�A��#}q������#6vR�@�hR����ZaUsߡ���Oh�G���G�q����YyT�n�}�l�z�A��o���
�u�wg��F�e�o	6{�����"����w�x��Z+�u]�9�<U�����āW!�E�Ė_������$A���=tM��^��7J	�K ۰0b�[�Z����mo��i:�?�Y���P��R[��jr�\S*1V��g�3=}�e<�ñ|
OB��F��G�n�}�[Ӟʈ�'7��'��c�0"�M]�*���ڭ�)V.o;P��O����r�m�
�$J�)�E��Y�h����CK�aǪ�A[��
�9��8��Qh��Tu�	"�M�|��JH�����S��yt�N~i��MedD#(���|��ty�_!�X��������+Md�|���D��������]��9���O>�Yǧ=$�\��\�꩞#�;����� ?�K)�#��[���>�K�s���\�`�s�*��2,���wa,>��n�^������}�۱�A�:nu%�f��Aʭ)=��41 �?�CHn�PY���
��K�%��,jcE*)��Y�14�b����Q@�ۦ����C�R�D��4ﶄU��>�E��!���u\@��:98��Z�1tM�(<z��"�^�ݓ����LQ���3f��j!��+m����9�~?�~���Z��L�=9��˽��³Y�0�+1ŉh rޜ[c��c��Zb�`�YAꕰW0��p���4	��"d*��&.J-�7�+6=�$�����SӇ�vJh��+��"į����n��+zp����u���6:�&4�r���"�u��y�Ҵ��xt�"#�\^o�����2����Rno{C�ڰ�)�c���^�$*��>N���+rV��r��P���lok�)p|�:����w~_rc�����8�k�h~Cy<9�	vZ��57gם�=�Q-o�����oΏD!��J��z���g�C�l�̨z^�a�_)S���b��H9��*��Cj��O�n�	��%-����Ks$
t*�8���@�=B���=��Y%9��)�D��ZY��J��J�%0�K���b����_λ��Dص����Lz���{��
���e8�(,�G��j�oy�A��CZ�đ����r�a���·���Hr#zi��-W!z��R̵>�۰�F������qgt���5d!���Ľfp
%�HR���h�T�Lef�����U�y��F����5��}�Ūϧ��	^m'M�؜�H1}�(��p�I��%~�(Ư��{x��{>�h���I�w ����6D�q1�B㤌��i�z��s�b�S`V&.� g���Nď���,�N���\�s\�0g����q�7�oe����Dӗ-��@���È2�����]�"�4cw�?����6�Q˺N����̹��-�)�d:��6�N�_;���J��|g�ӫ=�t�o1���z��E�1Z�����+�e�ǹ�#�ԉw�H� 7�vل1J��'}�M��1F�i�>K/ @��ޚzy���ŭ_#bs�D������44PX��-�Y�s� �Ć��[�C�h�ɺ��ΪK��aO��"���_�$�T���6��Ҡ�X�}w���z��VZ L�w����u?iO;N�~�����N���|4�`K���{�U�% �N�z�)��f���`�F-���a��j��^An�1S��U��W�~~ޣ�YsVW�yl40~Ӓ.9����"��ҋA�,���1���F�GN���W?��6�Α��^R�T�A+(j4��������p�[tS˓H^��)��_���6\TKNCHEa�%t����0ԓͣ�p�z`˩]�������k3h�������)���4Xh�G����ze�a�LB�6�rثU�䁷Ԏ����-/:��nD�@�K��k��+nWg})��~���'�v]�8m��xJ�+�R���a��� vnm��ep��T�w�&����#�ͱ��y&����#$0W(��$!�R�1d��`��t-Ĺh7Yc�o�h�����4�}M"��h���W-y��Ԍ�Pǎww%��0������T�|������ȯ;k���_p�t� Z3ޒ�g����ŷ��4fi"���08��c=oQ�~Iҝ�mX����5n��F iATt��tչË
c���Y�ŵ�5T����;�e@�f�w����42��v�C��"0��D��u�a�~M�h�ޑ����2V�D��-*�!��K�ԁ
���������g�:�m䂻�i�yu�4��/8�,eq>�0+-L9v�1�C�$>^���I(NM�+�6�;6ּ�y��R���_��X6=�/	2�B#z�l�:5(��)ݏ�f߇l����߾j�$��,���63'k�T!��Çs�P$'�EӋR/��� ��������X2��J*��O�s���[$���"Y���|��P�.5�C�(떍3_:�6��$���c��p�"C��%�]��
_�OFzT�fи+{	\]�y*׍\	#�Q�����w4�zV��˨X�a�m���JC�^�<�,��7��k��qS��i�N�ɛ�Ք�/n#�Z ժ7`�d޼�������z_��lN�_������g*8�HÙDh�k�޺k��v`픍	���^��3Cm�?ۮ��A�8԰$�+ۮ�&Ԑ]�����Ud�+��9�%��.�%0�~�U���yL2F7e��;vB�F�}j��4��/�4�A<��h�ћ+dZ�&������@iޙ\o�<���aC�/�8e��&�����Qc�ne�TE}�H����hf3>^�P	��Ѯ�H��S�V5�u+b��yD�Zys�q��۫��՗J����;D�N�w9������
�g�t�'����=V//���Ȅ���G����𧽶�xm������{�?�lwAJ�)LtK���`t[U9���DjK'�hݑh���G���9�)=]@�3�ǰ]��Q}%�%�W6�8�"�J�a��{'���*��{"�s ��NV32�ĳ��bb������4A����V�+Fg>.� �"B��8�I�ZJ��D�j%m[z��G�KŠ�(�v�K�����n��a#���Pv�w� �٪�/�sDp���:��A�7?0����>��]���E+������_�V���Ջ�M���������I��8�rZBѭz'M�"�U�ͺ��I���]������?�.�V
$MF�X�:�Ώ�]g|3Z?_EV��� �$��}U$�=���黺`3YY����b�3˝��K� �n2���2�:B���kW������F[�c���z൵#?��ok$:#��יPw�-ݸ���x�t��F)��#��]�m��.��z3���"EG�p�v����ǖ�W�|E�}e�Tt�TY�����#G3�W���$�K�,I���v����f�ݮ�s�5Nv��,����'ڮ<�ѬҫdB%�8'���VT�I�A����!��d�J�uz�
!�2m�췄ƢS�P�L�y�a@-4���]�aRALD/���U}���6��k[~�>b`�XqY7oC9[�������b�����.�ZDH�ʞF>�$=���zo���x�㮇 �D����P�l(�?Aä�7�Tס�7�[l��~N���<�ʗJ�S�Xj8�na�UϬ���q�ܫ��c~���So%�Q��C0�a�"��b� �&y�A��9��r���i���'KE����B?|��.��_��D��깙��. ���)�݃o�i���FR�M�����d/+l)��[�ϊ�1�0D����V��g�	l�"[�r�u9ji\c!����,�긹o�2}�ʪ���,4����&��_����,Kĝ�-����3_�ӓt�팽@�.��m=$���m�I�U�g�_�k ��5ڙT�c֐�f�y����a0����@.;�$s�K6��m�"1#;	��$f�8�Q.0�Xy�b���ԷgɨY�C-��Hs�A��+��ld.-�b�k�ŭ �5[F�����f)�J�Vy�*l/���F`�!)�+k�'�ޫ5�O��+T�E��W@�'�����^6H�1IDC�s*�'�r�ۖ��I1���z��n��Q5��y��*�=��Pzj�y�����;�;@��!O:2���A�����W�F��$����_� 5(��g�o��~�m�lھ�p�
g\8l+&g�\�Rh�W�/��y�&,'Ax���d��X�=&x�{!��4�:~�o���l9X�!p\N$li�N[��7�n6 LZ�Afی�w�44�}���7\������P؊$D:p[#nLl/�i;3Y= |�D���&#ӥ�e�m����z�v�B�D��ڛ��Π����ޖ��gԫQ��q������ĦC�7����{��YE8#y68B��g���: ���:yS����	�4��:o(�<q]{��{�����,�Q��A��"�ZI�����]7�<�1�*��Qk���>��i,�N���E����ғ;�ցޤI۴�[eS�u��5p%r������wk�.pa�i�[�_��E�����W�t(���roP>�y�ڠ.�̫
�u�F.�__v��"}\��ل0�;�(,��o�4vn4�'
�|t2�c�w�Wt��&BK�ɽ ᨈ��0á��h����RªVl$��;%:��TO���������=���n��7��`"h�h$<�/
k��T���7������*�[D3gr�Hmavq�� "��lWQ�hY��М��%�x�!��⏾�\v6�}�O^���٣���4�KC��,I�(��'�&�Y�Ы�3�֒��s��Y�`u�D��*�8�U����C7o��[Ш��J"l���sF1�.�65��=8w�����"R=PR���&�=��m�GE���)�L�5Ãh��oh)����\h��[e��=�Q�ӈ]��b�g�y��]��*Av(F#���q��"L ҟ*G՘�����i�] ��1Z%���l�_�*ӽ`����g�@�sZY�	��7�jl5����Y�6;p�����	�:P�0o�� 5!R:q-�����]����I_��͐�h� jݕŋ����S-~-��GH��u�#e��,e!%a�x@ZI�RI��ՀJ�Cئ��� ��Ӂ�燠��=V������w~��4$7G(�شM�,��Q
��+��>X<�V�}�B:*�{�?Z�NԸ��S�B��`?��_�W�r ^���%�,byݚ�
�ִdg"��Q��s>��I`���W<2�9��6�N|����ht��>�҂�l���� ;4� �e '�+���-K,�,Ҷ�2UR�D��i`�f�����j��ݙ���Y����A����󊅞H�x�+<��i �W��#O��MeR�3���x��+Ѭ]��̀_c\�铝2�n��X0�]wn�W	�~,X����\7)�6��<��T�:<#�ApR7��m�C��y�㵗���)��L0
��ޠ�����q�߆$,�Jڻ�i��3�[����
�IT��״!+���hļc�t�f��l#'[�Z��.��9�#x�M&@4���|.	$j�U�<���C�%-aq��0��kg��DR��0��$G3��֢�̳%�rԏ2���r��$�vu��ڐ⚂���0G�e\~�lU�\�5�{<�����Y��T�}��s:����=ȵx��Z�U�pMv�Ҵ�8���w8���5}�,9�$d ���W
)�`��`r���-�g ��X�STX�mn�]����"cɿ>��s.I �k8���Y��?naa����K� ����cn'���9��=��ᱜ`����ӥ��+5�{9���dhLG��^���'��ʇ��ݚ�`|= ���������Pz�t�-~�G��߼S��,���8�����?���t3 �e�g���Y���&h��Ӂ�ۖ�)Pc�xz��Kh�K0��H��*x<�E���Nˈ6��q�)I��}|_�k����텍=wN v�7������})��Q����t���C�F�_�8ak�VT�pr�����ω��������1>��k2jHKTi�TOul`KB6����l'r�z��}�F���ެ����B�L8v����ٚ���(��O/G��a+�ij��_�jK��� ���w��� ���c�H��R���YsW��f�^���0a7B����}��@����9L/Ǫ0b4�d�݈=����5l^��������ω�q�E5A������t���=u��a�N5���vu�nK�y��Y