��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0�����(�_?V~��
�r�-�$�6e����<a-
d6����L�}���W�D�Ѝ/M���`^��5b�L���OB�M���3�
{�8�bvq�62b�u�<\.����U3��ZÃ�'�l�C���)��J��}Ѽ�ҪI���e�J\+�P�j�?[��CO��P���l��1DT�n��*�k�K��~kP^�θ�����Mz]�Epæ�ĉ��Q_�P��t���dh�s���bN`���F*�3��W��E6�;�*'xl	x*+�}d|1��')��*�w�W����}3���?It2��_YlLq{���eq�SP%z�]�s��E2Ţe��A�j4�G܈$඿��sЩ�BB�8���kK� ����J���dў��\�y��bTi�1�[7�0H}�4�K;Ț���y�^��Oc�B�IE�W����5�Gj�|�rN-HH�lH�ix��z�g�^�bР
�׹6�?xV;My�-�?Rp�tBKk��mǩ�>�A�%'>�j�6I�,R	������)��L>�Uߜ�{l�E��b�d,�mF�6�!��c�T��ȶ)�Z�,\Pdr&o2,�-P?�bK�12(Mӹ{!�dC��T:̫\�OS	����SE��%_G��-�k�P��lŮ$�/���u��y���fˍ��C���DH��3+
���Q��cY�X`�h�Wv�������ѯd���o��?u��Ƒ���1(�vuuL���q��sRSa���"4/�${��j^G�%Uk�+y���ߟ��=��\���Q6�5���K4MĮ�wSAIc^��RW]�6����!��h�13�#�+?��� ���|m�2���U��>�L��� ��G[O[#5z8J�α`���̰�1����f��rx)KU�:�U�.�.��O�EB��'�m"N�+i����?U��c���*h�}���7ׯ����H��w��8��H�p�á�$��{i��H>$r�s��qGH9���42=L1z/o�x��M}u[�r@���&��:���@5Bv3�g�\�h��o7�E��~E����?���4^$7�+#��� ͸�U`Ш�D�����ec&��)��|r|o��b�a�&2�L�ݏM��c`<{�=���$���9�׹��lQ�+W*L�&�^��Esx;�_#����l���Wx�/źϔ��84Z]��4.��*eV
]���E(�Њ#�M �猢K�4��4�|L�K������N��{�����������1;���M#��Xj���#�ۂ���oR�.П�D� �1��dx-Ǧ���hG��2Ϻ��v��+���S,��\C�%�Pt:��t�u�
[j#�SȰ`:��`�eR���2ցu׹Bi�g"�%��hؠo�0cd��Q0��X�M7�\A]ɵ�)�+.?�����C��.�Y̀�O�T�b��q�n%'W !CC���<�d�]}9Zj7>��6wQV�o��k�]}���^����3��?�l�
�>��y��jGy5'�&d:��	V��A�~�GP6����H3����<���2�R|�.(�*5��̈�H�-o6X�m)X����ʊj(��h��[�<;4�g
�Wأj��c��1Ft�[
s��Ý!É�+�C�杸��UIN�l���1�3gXӂ>�	�y�sV��
�~�>�"yYhVL�&��Ge?OKOӉ߁��W������l�5������ G\VN�����X`�F�ݎ���*j�<4�%e��]�oi��#�l�ް�x����酿����<|��Xn�~'�aY\F��Ǽm��H҂ ���d�,�����-j��^�7�����:�=r����&�i�M���@�5�1��]��R6�Y��۪UQ�� �uf�Y���,�!Z�k���ۛ��9#�x�2ڢM���h�4���j���ٙ�
W%���{ݸJ�l�k����r� .j��F�a��+���져W�����*L )�|���,=�q�pǔ7�'�g��(�z���"��t�_�G"S���
�
S 9dm� hڍjW��=�]��lyt���fga���C+5W%��(�`^١sr��4&����� S$�(f��Zi��.�祙ހ���Z�h�g(W�j[�}�����h