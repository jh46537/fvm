��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>����rhhm���%�ñ��\X}"y�GM8�,�eP��:h�Z�{|��L�~�t ,������DN�F�	�:j-��u*�zn���{�h^���C��zlC�Wg1MH����{[�rx&R�+0,@Q:/��ц�?yU��g_b��1���C��M����훅�[�>F�?X�	��ϟ�]w&A���E t��/y[�x�b���튟Y}
�]�w3cGTe�����F;;�A���|-�¤��^�{�w\e�+����"-�v�E�`iӆH��n1��Z���Z"9߸���֦�}Q^�t%��$w��=6�e�C�?'G;n�F� O�9�Y�,Q���X^��"�p�񔺖�3ЄQ���W*�'0J��kq���>|6d$j���V�+�{��Yf[�( ���_��qd�pY�o�4�8h� 
��ɴ884�|�?�d����R�T�2� 0���Z�@�ev���]�i4`_���񸝭�F���f�!
���:���C������VQ3�l�qǓE��	&W�00�E��UN�v��/�T׷��;S�O93fu�S3B�.� fM�3+�B�)�UW�Q��e��dCc���f^�n��j9�Qs]�8$z_�l�h����S��OA���7��{��L+ǭ���"�� ƴ�!���A�w~%4���k�\!X� �3?�ª�@��O���/����<O�7ۮ��cL�*%A�qA���
N��k�؀jj�@�8q��K� &/L݋�I��<�P�ȊU�LnI^I�Ͻ�~F��|�))���]j��=�L�Y��q���❢.!���Gqeg�5I��!Fڅ'F�]��(�a?곸���������^�W�����*����Ր�{,�i��2�T�|޸�/��`3��1o��V^��|L�dH�Ir��%5��+P}��
^�JZ碜C�.��Y^�����H�:b|�.ʤ��ț�n3��C����A��"�\�k���*'����ؒ�5g��ל�!��U|*����h�5�[�����Ᏹ��f�٩�i^�Z)�<�Dĥ��Y20�=�Í�g�BX���I�b3OY��~���۝���0�OY������Pd���#���'�Vq�2�W )�w��&D�q�o\eH'M�	�t�s����x,w;������*ޭ'��e�VJ0�?��;wn�^%�k"����M��a��u��G�w��>�V!���#�����Q�ܬ?�����"س�2�^�����҆
�+�$�i�\�/�,�yD���r�m $|�˄rc$��|�{���0 ���
�F�m��Ҫu^�D꣸����pX	�W�����%d��1�3S���j&�i�f_����!岾 6!�kJ�x�Xw��:8� ����F��f,�J��^"���.��Bb�CE�� |	Ky��k�z2�i[%��Be�M5v=յ�0? 5�1�d*�H��C���H͋dߌ��Nzd1n�5��A�6�n(�����B[<�>R��b��l����"Tř�üUT��O�,>�n���Â_�aX�,Ф�#?�Vx�5�� �7����5X������X}�T�b�y4c}9s��f�������թ
�e���vۤ��:�·��l_.�Bz"6����toD�����> ��VHM���%Mj�i�>���(�V��v��ב�)�ts$x<��-+k���MT�u�����p�{^��W \-JwN��1 #�#|!���s��[N?�9}	�@¬�eqb���@@ <�Y; N�݀$-��$�檵�c@Q�=�b�[���j��e���E��8_����YE�o���fk�{8,���j����q6�=:n������^*�qT�/^*��]Ǽn�p"�4Zq��<���Mwe�,fkO�7'�2H��-o�P��� ��+Bf�,�x�?���D<�"��&'�K*;����_oY!j�mW��~!�^9xC��Aή�%����\`�hgv&��\��)z��ا�[�H�F�Ѓ�q2t����gޝ%��^�%��Gϴ
'Ti.�60�ڞ��C� "k� ����������G."�\��=�����c��<+<i.N��� �&�tlt�-��i��<R�M7)؈��i6f��;3��e��/1x�D'�(�r�HG^�?��[�,NMD2X*��e���n��p�'^�t�yj�EV�Y_�ɧ�k�[t�:o�|��y�-�>H�<��w��c7.|�'�M��EQ6�r�3�v�peOץ��K��ڌ�SK*��t�xuGT�2,�[���,X��n�z#�Ѕ����.�̞��1��Z�X��1`��}��i����5�A�?�B�1r@���B��?
�¸m��ިU����X��̦�<Y�����j���SXH<?��!���[}6.�y��m��N+V|~SO �r�H���/C��Ʌ~��\�)U�C-��gR3$�Y�mKM���vu�3����*׷>)lv�' B��(=���3E�ʡB�b`���H�������O�8�'u��<����%������)�i�;�q��wn�9���I:m(�]xmqE!�c�Õ~4Y�k��7���GVڷN��-������@~J�b�@��)B/-r
�i�����ތ�g�9Wl��5YʦNt<�}��3��	<�d�%�	��~��M�J�S-n�Z[�Я)�".)[��2N��/M:���������VJ#�Ŗ���y�ƃ$�>���;�(M��x0�aP�Q>�P|;I���S� ����j�+�w���4�}Ut����>����׹�,Ǎ=��)m&�>��7�=2\�;�g9>�
�$Vx��kV���w\|bA��3+Q�&����%���Ы#7��gD��h�'���������eIG��ݼP�+��Nď��16:���Jߡ�Z��:V
r�_��P�>�x�p[�K�ڈy�~��+�Y7����0�Z�y��!�a�5�s�V��E]�ǔz��qM�VC���"�aG^�q��P�[����|������� �F�?]�e=ʋ��� �i�;��9��x3W�o_@��%ˋZ?��q��R֎"ĉ�z��"�����9��P�Htc����'�蟊*b}Em�;k�:#)��+�z|�Ks	�|�yl@ufǲ��:�Ƞ	K��6��H�3|�'h��B<�ݶ�u������\K�{��s�.�S�Pl�d���`V2�O{��S��C��YM�\ ����W�Dͱ��uW����6H^1u��bɓ������E�G+�A�-��It^�������(?)�=��{Y�v�uoD�z�4�d_'��l[B�G�?Jҽ�ܕ�T~�������5b7548�/�4��Ngn�8@�z�7�-�%�}��,�g��3�ߥPd����vC���U�O��������leU����h��������?��f�o�mL-S�Ϯ�e^y-|Rx�,�ϥS���#"T2�ze�&HOb�<5�'RƯ��V�f�U��.��ttU~hc���І�).�DX7��
��mu���ro+=&.M/;y�'��	��^�(��굎5A�lF������M�ݍ"��B;� 5�U���Ϡ9K�m�[�Z�4�%����������~&�Q7���?���FCɋ�p9�6H}��*���o�}��y�t�^�"ix���ό5e*��h'�z�[Ȣ���u]�vAw��3�l/or&�]�):��(T{[F��#��.����=b�)b��g��}���+�4�R��+����H���$�i�A�T�]3ѯޚ,ky���	�>�񩗋�(p\Kd"럗d�k��+�5{�'��3���~q�(�\�v�ƈ�̦c�0+b�Z3r(���%�6NG-��+�άq�'^�8���I���z��)���
��,`A=��'	��<�b���ٲ�� (�k����\?{|�s%4XZߍo�=����Ev},	�KyTo;S�t�����h
�Q�ҠNҺ���K���.kvMA������Z��'�[S���<��)ą�Z�!)j�����|��@�6(�o?�5Rc�[Z;�K���W _M���B��r؞��Kj�&oZ}�ged�=9$��;�"ch[�z��u���@4XRr��
�������(��)��\�j��|��u�o��,.��l��`r�;�4y���;��\��Ϋ��|��L--�ߺ��IS:Q�����~x���-��p�s�H@����̋H9���6�m�#l�,�����y����c��[�f��<�wؖ�	"nЙ`qh[F�yC�d*�@�V��[ԕ�%.G��D�Ap(t�N�L�h��r®i���uL{��^ �k5 ��~�9�Ƕ��G�ö�%��)<����^���t2��D��y�={�?�}�EY���<L��͝��X�*\m�u{@m���ȵH��ځnn@Az~^�&(uwھB�bU��\��K��[�Ϧl-#�z&�U�U��fO�x�숯�O���������x����-�B<z ����;�hS�q����J��j�.r�8����r�L<3��[