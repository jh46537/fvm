��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħP	�(<�%5,i v1`��Z��7#��e4��������UZ���������n@�������
�{�.�#8dGo���^gAT��d�܀����P ɫ#�l���Ӫ�w:�Irx�J�}�ō����@9I%�W�(X�vojL��WQfr*x�7Tiy�3`���c`�t-��z��&��<�ӡ�<��p{�� ?T
���#z|��u�hMfl������2����0�MI���oSNP�<���/��=*�����@4m�2��߮[��bf��$���[˙�
�
6����`�:ΆZ���y��n��◩�|�g�![�a�Lv+��!��w,����3�P�����u�$�e�؇�K�D��*���w��̺�c[��.i<���Ʋ!ݸ��'���]�X�fŻv�
���x�Ґg�)��\&�3�e�5a��ib�h��0�M�^֙��(��{������~M	;����=|g�k�
>g�!���WP�-m6��?�����_�1�"ˬ)�)�	o����L�ܔ6O�)�)?�'�  La��C�!�Jf��djz���5ψ�<h����lefH �]CI!����݋=-R j���vDѩ�=5�
��D@-XVű�����y����F���J����G9�sA"ѽ�VQy��J*��H^���~n�pFsl[�l,5�<��cSdḚ�i�5%�,[o,-���-r����x1&��g���9|���3Q�=7ł�l�½��^=�X33��s�4�	(̍�i7�[D�E��ʀA�ƫ�V����#�%rk�o�cl���\�Uϒ�[�e/b[Y��#�΃���'�R��f��-�7��u��||�` Ѡ��t��(���#�)�K�<b��îx�&o0��x%�IC����Ț�b;6ThIH�w��{K����ʕ�����c��Б��1����b�ŏ����7kK%��>'�6@����,yC� <m����Em��4�E/�/thZ��s�f�.侙7Xec��8ш�K|~g0�=�9�n���01����q�����Z%b����2c�%�^o�[Hf�d��*�W���gy��]{T+����f��w��g1�Kv�^�[���b��
�:�{J$��.뙄�SN1��ĳ=�
�d� ����_	Qg�Z�]��P���h	oS<l�e�z���"�Xص7f�w��:���v���\-��%pU��A��h_¦�y�zvj�H;l�9JO̝����79M�)m_p��������d�5;��f �|��gG]�z#��ah��8"r������Pp������x�vU�E�Ip�j�\�h��+�ZR��ޙ�Q�R�
�9�G��(����������e�=ש\_g�d=H�A��Zt���>��	*���c�6Rd@|�?I?����u=�'���ػ2ӡX�ws�����ߢ���G�o��4��	k��6�k*�\h��$�$p�?َg�5̲(���P�Ж���Τ���p�Etp*�D!6|��w荓�pT�����GJ�����ɂ��Ҥ�a�o��lo���
�'!��5��[���JX� :6�P�"��H�:[e�)]A�D{��X�7�O��C�!��iu��f��l\�t���.� �H���.y�w ?��E:�%�Y���O~���kH��"�SY���W*PSp�7@13��&���~�N�e2��?u���5�w��j���i4Y
�v)+�{���&,o�W�)h�1l>B/���ߪo2���(�=k�_��Vy\F9̰�4�a-��T�ayn��
�5[M����B®���:$IYp�J+���2�����m5�+��=Yǧu\��d9�_�A�6/�B��ޕ�7�7�r��t*=h����\W~D��dd�eº�fp%Tp����H��U��a�Ɓ�;�����1�UU���{p�N�s�@M�md�;��6n(�2�=,�0�rnJ4���-H/>$Q�ad��ܢ&=�'w�5�R���؍!8�7;)��'[�KT��	�wt����cR���I )&	n2��t>�l�$A�@���i�`��4v�g"x��j�/ ����9NvIu�M���1��r7����Z���+��q��a�#��: w��5=��5�F����R�#��ǇdЂv���o���}�&h�h_"�G#b&P�!�j1\Db��
��oUv��F�̰_(*��1EY�� ˿�1�N[ϳ|��lb#}�~8��06C_m/���o���*��y��5�&P ����K���z�3R}�P�KT�e��a��9ga�ӯ�����W�H�A�xx(����I����L���8&���3/�=��|�N��
8E�%�����Z���Ȳ=z��H��).�L_�mG��Bx�U))U�-�HP{R>&Xc��תz��H	7�^I�n���_ g!Mb让L���L��{;"�q ��3`�����D^��G��C��[�ޑM��"6R��hޮsUȴ�_�C;�r��4 q�q} V��FA��A��g͕H�QE�_�� ��
�տ�&���1�tA��s.I�+
i��WL|��SLϪ멍��49k1[���0P۳M���&���$�5�O�D�rf2L�A=��X=|��%K]��숡��?)��о����g`�;t���gME�7&��=��?P~Ɲ����v1Wc��8K� ���R2��i�U�/�����W^_ε/�i,ˏ��`	�"')Ф��SXd07Z��*VyI ���V
�:i&���)�)�۴�<5��t�¡�v�i���Ֆ�w��̼:wY�,d!��n9K2( �)��>�=���Eg�^+�:��w��f�K���(��>�~�xB�J�s􆞲�)N��Y߬-;Px�6����S����;�J���PvC�%��\��"*Zo��r?�U񣟓pw>�8�ӕۻ}���oQ�xv�4f��N�K֎�u4�iƍm���y�Ç*�'I	?�^�����^".T#�H+vj�O^$r)�,�̒Cpl�΄�v,����0b"�1��T=?޹i؝�n���f���❥/��|ن��I���4UG0���ƌ�>�j����T��~R�_)��,���r����@�,�JG��d�2��,F�>���)���d�&�P�O�D==U��3�;T�w@�d�=��3��=&;JI��[̉����ޜi��=�n�����3��+&�����Z$�?;j>��?|�V���4;���	p�-���ج�q0���#f����
���A�`	2�8.���PcDT�����=�L�!\d�f哤�8�R͓y) �|��so
ڠ�t�K*����,G�9�g��J�褬�m☆�Y>:�c��!_i�\��п�y 	��?����0o����I�O=-~/mY�8"�*��l�:\�C�eH��Xg c/v�x`�A�J%�w1�є�i.����/�oy�j����F�=�h,�Ņ���ԦҔ�p�+9|,�4�|��-��I��p��4����d��Ф�`���~��I�h�p�Y�}<��kB_��5|e����vu��x���F#�-�U\�v����Z���P��{	�r������j��lٚ�6�/����҂����F ����˕�K�D����r���=*Z܀mw�u�����q;k�����\qO�R���<�M����4V-;Hz��r����G_v�&��r:�h��V>����բDk�+���1<��X{c�

��5��g!F�b��� �Zjm���&3�Hu��S�(5c�� X� @q��j�RfŽT~6���.��-�S��8{�Y����S���x�I�		��[n���5=�30ތ�T����&ˈ���'-�*9��M[?5CC ��bׄ��k�г�N�W� +��i�b��My�~�0�/EgK�mЎ���d��C�ѥά���:�	���J����F6�������	�8�[�e����d>fy���nɳ�9��fs���םN[���� ��������[�>p����#oQwd\;�>�_a�N�} /��e9;k���%��O?��$�R_?�R�\>.H✪=ĸQ��v.��c6-���D	W�r4�Ͼb�P�F�`'p	imeB�i	��'_&��m�i��Y&�i[&Ԙ`��4!:�S��Y���5{4���m�kr���<��>U���]|���f@�)J�6�e�,h����m��eBlw�QO�d�#�����J��t�"&?��qԎ.�8%]�2���Õ���FE���ppJ52��c��,nk:����u�>s�>R=}�Z���t9s��9���|�;�8ÓnnM���9݇ax���<۞#i�*b������Tݠ��eT�z�W&e���B�B���T�𮯙������m�3>������z�M�Mtw�{���)��Iؓ �����sb_E����P�S{�iم4Mu{x�[a�'bz��Ț	��W�=�w[�§�����M-�m��<�]u�*	lJA��-� �VӰ�1X�������+wۏQ�X���Ֆ��Hw�\��c�l���\�&��}V*�~����T���L�{t��d�����-]�XVA�X�����}�^��R�9Gc�w}l�V}������f MVv��xľʭ����W8e0������'X�Y5�Y�H���S�F��R���	�t4{6䎵�7�|^w]���W�7�z&�Ph��,��ӽ�Y�-�)�A�.����T!�1�w8���e��� Xne��i����X�u���. Z��O$�W��̸�]�br�Uz�,.�ů�o��*7�������ɊՄ8��7¤QA�g�F5~5<�AQ��]����c�	D����f�yǡ+�\���j�T��a3��0]Kjp�^�N��4��Gԓ����@	< >�7�����ǖ# oʴ>
ٯyB�#��35d�<qyx�l��Q�u}ȡ���R>Տ䎶c��~���!���t�s���}��D˰-M�c1�]@�����n	E�%G���=�Ό¶�I��$%?+
R^bz�54�uӶo��`g��	;�@8�YeEI�?J�i�n����5��&�w��*HV�������/l>��K%��δ���g�f�qA��J�6K�R��޷���%𢦊�7�Yx	`�̱�����A�����	�|�t<����|(2Ѣ�����f�P�T��"t��� 1E2�rr���E�̏�wv���ގ�O���~����O��%�F�y�!_�W��6��]7ƂX�._?5F�S����a�`�P��)���ud��k���&����^b�g�:�<� �! �v�s�N)���2LQm��|��V���������߁CŤ��\5����{EL�Т�l��|I��B������g�[$2A��y*E�!|b
9�)9����y.�gH���~�rq�+�P����s�MV��o���)ˤa��&U��@(_g|��0[>�����o9$]s�K�:�3����!�Qñ�K�nò�[�|#��) �N�B�|�R�KZ�)���'�cb��G�Ri����@ip�w�L�[���?N�v����3���R&<^����O-�T�r��z���i�c�K��S���9������)�[Z�г��OS{�T��dYU�uZ����FF��Y� �7�S��ƺ���dGH�F��M�9�3j*��&�3w/3P���) 41-���z\D�6O(�GQ�����Tl�V��9t�5��D9#�ڲ�p<Y�(U�꽒�V���v���e� \�%Iv4�������u�8=ߔ@~����5т���I��W�\Z�N�\��t�`q\�-%�!B�\փ�?(!���A�dR��ܦ�����u��I���O�:��O5���UH�mOh�L��tz����'f�C�v<G�疸���|_^Vx��I��b��'�X!��8���:���^�ԝg������;�r�/v���5O�o땪������gByH�z��>»��s1汃_Bv��Z��eK
YM�*L��~�+C{�KJ@$=�.�.�E��~�\Y_�܉U����ܮ�`�\�~[��b�^
]��r�7'�5�Ս?� HV2�#Q����I� �f����T���aG�?�<���Gs;��|��|__���������:�'(�^V�VTqf��"��s�/�/.�s���"�	���s>e��xiW���Q���%��%�Rϻ�i��)�s4d�z���0��pi�3��s^u��L�e�q���Ъ�W��R��^;/�8���__���ޘg�b9h�6R��+�o�jx����6�z HjP����#����q�f2<��:�v(lh���uD?U2���3ܜ :i�m���[�F@Ο�*��c��ه��	~\C׀e�&�`�.E��� �~�����K&RD]×g�:��1�e�����b�"W��c�3�����}@;��%ezәG����!uK�7���CiE��:���p�W.��w����T��O�2K?uN�LJwJH
��׍b�#���E��{kmE�}'J�m\n�|��Ĉ���6���S�۴�e���wl��U V�G�x�՘�"������;`�����؝}�8�5+E/��J5R�`�#JN��AL�vp�D���s��\�/p� �ؚ��������� p�f��>�+�l
�h��MU�o����5�`�7��rV��\����0vt��3���'F�~�r���[���$|�����^_*�s���3�%;��SU�ӏ�;b�h��9պ3���IC;"L���X�|l�Y�N�7���t@�οm��v��Y�H�B�dȴLTnn�Հt�\��_�V�G��55��v.���������p#�5�]	�:Ԙl:[!ʃn��+���1�
>��	4BT��7�9FN��X����2����N��[/��-���3Z��`)��o?�w��� a����<9�EZ��W��/�5���\T����\"K9��rV�Ep�C@��|c�V�լE����O���$�{jOR�5�q�S5(�,wZ��c�<�gMu"��d��«��7'U��)�)�F�FI7�[��q�Fy�g�l	Ą�\�н��𕄥\V�o3%!��̯EG��?T鯇if��������>�7x��o���c���S�&w�P't�2��|B=UZ��G��s4��hC|4�Wˊ�Dt&�(S)��,%���g'ܖ���)yf!��'C�k�e����F�%q�vu�NE���j[�+� �m��������A3;�F�V_��?�YGP�b��#���R�;���)�J^?z�&����`M*Pnj�'�U��؎T��IQ8���y����`f��>g[��I�@(hR��W#-FlI����!w9u�}���d=�o�?�^�
�3�3ހ�0�@���&f>������u�����C��5��,�o�~E�jYT��7��^<�i���^{(�	��KS�(%��ό��s�X��^Pw�>�s�8e^.d>�߅&j�MΩp���}��')ڠ	;�����r��y��J5j3Oq���s�xw?�u��d���ք	�._V#&x��u/�К��hw�+��5��9��9e���F3��������9�*/��C97忹���O-i�6��X���h�.W�(,f��Y�L���J����7m4hX�w�;Q�U��8J�/���� 8�k��u���iU��&�6�5U	��u�!�\ʢ�/;������Ra�ˁ��w�7�/8	�n���a�k�ze��Qw&Q��SM���}CƲ���7�(J�a�6����z�Pպ���zX��0�s�},32P^'zv��.� �()��'*�f��LQq�̝Vnz��t�x��d�So9���,�_����c��w����1�{�9����
��@b$>dp\��W����ȡ�4�:�#zh�?
u!�7�8�6��P�-'L�EFT�q.Lg��O"8��>��C9##�(�����T���"�;��q����84%��=��GIOK� {��3���8v�b�-��7��r��O �wQ���u�C(�Z3��jJ��0��yeb�p]��%>�w���2�RR��O�.癴\���P;��n�0ɀ��A��MR�u��	��m�g�C����mP���F��C���f/���D=�զ���rw��`[�`��a��t�5?��������E�ONj}x����n�r�?=�H�?���I�kZb��*{������3)�������M\͡�4���*)�չώ�SxqqRa�E4���9��5̉O�E���`����@��L�_\�b	�uF�ۦ���L���LA���0
V����V2� M�V�&L���*OCz�v�AhX퇣^���p����\�����/Ub�n/�@�|c�P����J|��q�D�h��8̕���p�Ȅ���j;��^R��
��q������{�Ș�ͧg����+9�K�Ԛh��ZU&] ��I��_�~Ot����^��7}jI(o3�z�rX�q�i�Xy��&�>_7V��̀�62Rʱj�cw����s�׽2�������:.c �� �Rq�zg@�r����4��󌩚w�H�3hJ�l���A���3j�����`� D���8�w��
�u�(д48� Y #�t.	��#1��ȶ�(�E�B|�+^5�/��`4�Zr����)�U��ظ�S/�nϓa6G���	[��Pr(�b�\F��>a��!C���7}zr.�Xʎ" p@jޠ�
TY�k~2��m�S�A*{_̲"8d��l���]�_9��e-"��!���5Ǵ�Q�_}�GI-�g��c���w�;��͍�����*<ե�Z~�B�aV�v�!A��_3d<�|2�2&�Y:�������0�sZt�onQ_��+g9�#NP�d�r8m�+�A�����5SJ���<�q��1�ge���#�V�b��!T9��ڊI���Ӻ���k%C�[d'� ���T���Tɭ�0�Ǖ;Tk�S�oLY��pp�'Nݧ��*�� ����,�5ػ#�S��w�^«�K7�\�%Dt�u��ڢ�c��ӬW]���H,E���V��i�����38�2���S�yӼdDxK��:�OA��Ơ�FiA��?r"t�S�m��~��@L~+�39O�V璘�:bG�;Ժ=�b�$�&Q�̧vG~0OB �����<�Ly}E���p�΁n^���Mlݩ�o��[Y��	;��p%�D���x��"Y��6$~/����XS��Y#�J5i��ON�����K�'O/l7�����,��i���@��t��S�C�\&g���*�6���&@��0��������ْ��ٚO{dZ�a�'�����_�4ؒ7rD~��b��� �6]m�����)�O�Cή[�8ʅ�-Y������=�k���&���p��9s�!;������q��*�}�n���Z"2T'0��Gy�{�����	,m �a� FG:�nC;{H�=��ʶ|���֨�5�b�2����D>�ܹm5��-l1D�"/�p~��Q���S�u|WU�SO�N["����312=�������1��l����:2�ܓ���q��+[�-�$���J��C�#�V�f^� mm�~��9+��_1u��c)�aB���2�� �j�"��g�1���9��9̈́�Ŵ�#�%	�7>�Ph�BԲ6Dt�f���c1��i�Lm0+.Z�Fڎ-��.f�1)��z�Ϗޏ��K�%l��?얅e�Q��^����:͜<kStcVb�_��#zv�O��U�E$m�[	9�j4-���w�,1/��N��؆�k��|�iTq7��U��<�O���z�wA��,�c�2"�B�v�,��|�.�@��㎁�B�*�`ꬶ�.����2�t��6l�UK�nT1r<E���5�n����ܨC�-v("AW;��
n@r�ī$?�ތwR��c��4R3"�=�w6�w���l���D�$���ML=�̜Rm�O;+^��T?D�H��>��,1�P~���*�M�%-�Th�3M����;!�eZ���Wۼ��~`�q��RsA�%{<�Ҟ��/�m�L�����6�tUߵ��\H���J�~wYz�qZ8�w~���F1�D܏N�r8�WM��V%�Y!��%h8B��Z7Ա�X�b��%�����[J\5B���4C*���eim=K�Iˍ�NPx�W��i�L����_蠨�d����Z�� BW^7���,�d�����|sB�8�统�>�u�h��k��E�(�6]za���jO,b�K����e����c�;R1齚����.ɲ¬
�B�
��E,��T\�d�WJ��#9H!��R�`��r*"�Y��`��H�,a�.K��R�FӞ�J�r �3b{��R�0���B��vR�"nRL��6��/R,4������*�.�\6�yT,�M�9k�����e�3Ϙ]��1�(�I��j��f����k�"�����	w�3�����cRG��T�9�*,� ����4+/���:w�Ş�O��ɮ\0̤>� ��-ET��<��0Gڈ�WsF�1C��;��(�쪨ق��}�{�($�(L��5-���a�U���
X�	69��!�P�:�y�$��_k��/I� -���s4)�K"n�h�e���oP��HU�H���@�	@�=I��QF%�~�z�̨����B币Y23s��{K�:�J�r�yF���-���=0�c6(\��@�E<{x��t��s ��q%��Vw�����.��Hy�:�ܐ%�I�ď�/���TϯϿ=�QqӺ��կt'�=���� ��"*u����a��.����H$n��<�,�Ί���q�	;��ֲ�dq�/T�0��Y��_0M��Z�"Ĉ3�rX2�g��'p8)5a��$�M�� ��Ӡ3���Nש��O�0%f�ae��K��@��Ko�7����tX.�� `�>U�wwQ0C� ��#�I]^��w��GT�o�n�L����B�ډ��ީGL���>=��C��pG���=�E\��P���nV�Ӯu߇�V� bT���V����7��