��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9�c���]�uJ]�u����`�/�_.�~���8�l3
�����[�U��:����x���<}t!ĪRC����������j�}&JQ�8��6>(�Fz��L=j;����H-�&3:�V�a�y��`G�$����a���ż��P3�_���
��j�("�/�����T�6X�9���� ZV)֌{6��eܣ�d$z�g`��  ��(ړ8�	�4ءR]�����}���R���K���a����p��v9S2H>��Ԫ�$,��)����W���Ys)���O���x����]a@��>�n�~�5�����GK��
���Ф��4�$q�U4W@|��{î�`-������4��bdQ0Wޥ�7ɟ��פ�������vA�G���K0�Rj}��c�䷃F�$*Z�{ �ǉ'�춝�(6E�V��.Ti6�D�a?(��r��*�RL%)J/�Y/�dK-����C��&������o]�]��m��b2s^�Ȣ�/ �׀�(1�I-o��Ι���ҷ5K"G�� dӫGpThԌ�!�ǎ���Î�p��Ϟ���I�ROHp��Z�X� �΍Y	`Y-r�IV��Y��RJ�W�ܙ�:C����ډ�Ċ��z�MnJj��8�$#.N6�*^��l�z����݀T*G.�	��`�ag�7K��������Dh��j�^�����7u�U��f�EK������y���`8%�9����,P�	O�&!��;dz6��B��da]������p�e��0_J�1-)`��0����~�͞B5UQ�c�A��PfC�n��`Fc�ȓ�����)�0X�8�bR��:��h2��̂�����-ƫ�,I<�T���>��YBʶ�R�"H�_�ܘV�(cQ�`j��-�_S� ƭ�g����T�G�l�ؗ���o�7�&�_NSr�0O������b��x\��}���B�^�"����=kDpMw2�ߘh+�Q�q중�S)��z�ҳK���#��ˁ1�B!�hjc-<�xe�I����YBCM���DB�>��������b��Ә���(EG�I���oVym����9ę� �7��������-�����v�yan�r��'�q��,�(fo�Y�8���\�ҏ� ��gIi~L��Q52��ʘ7�
��U��y��̓}��Mö9ӈ��X�����k���%��#q� �o�g7��	�;���1sS��@ۗ>����m������cnm���e�j4�.~��~��vxj�wkZj���G� C�?�<NQU4���W'��;)�z�qD{~�±����Q���T�N&<�DZ3�л��|��%�3��n�"�0p%Pc�-��a����g�>~��+�	��sB�-����h���S�U�m�ڤ��
�3����±ũf
�>3Aʥ����4.�-<��Z�>��:�cO��}���%I���_��O�t3����;^o���=�fE�#�Y�4��t�&%�e�	�(!d�S�	��̹8�nl+�D�"P���^(]�,wo�&��*�Y��gC���P^܍ӝ���x#'-��uW��p~rWJ��;b�+�1��z)�g C���sf}X�*͡����� �����Ù9���6�:s��x�Db2a��DS�33-��b�m��`d�)3�_���}�i���,�9�ƣĪ������,^Lb�#Ž�<R�"e��R����\�{��Ъo0��R��< Y5Y`���=-�Z8��yz.�����iS�3h'<1W!ѿY]
n�ID�	�}�͈; ����9�I���0B��9FZ���k��T��5ju��tRC�3v�,���&�� � Jn�'�`#Obљ��||%��zD�����IJ�h=&���Wsd;}:<��h7C�x�X'zusf���,S�C�&5�X�1�OQ�g=�ǩ�!+�g'A�b���Z���G��*�,r������/�k���R���q9,�Tƅ"������S\rQ�!U��Š�F���Pd3]��2t�ԡSe!m\$��e!y���ڙY��t˓#<
`9[�ر�U̅�R�![
����6�Q�<)���T���\��Y@_v�8�O7cG����m�!�~{�2�v��(�7����x����T(P�/{�5 S�V~�=�AA����c+ۥ�-�#�EV���<�-��@�$ �#��A�U��?�Ƚ���$�6���})o��a�3�i5�T���-R�_��W��䨖�#����i��鬴d'���i ���h3\t��Er��K�ZpI�`���RfvD�!E2�����;Wt��]s�&�K8���ۼ<[At��Q�[R�Ă4)A0�va�F�-��1lJ[tVe�`)���;wJ�^���xca6[[�Yg��q�ө�KR�j^C��˽u�,(�w4?]��S����;����6]H5u�q��zۅ�F��:�V���?��qr8�.�B�iV��q�mN���s��uf�+G�*��*����Km��IR0��m8{���<a*�YY �v�l>o=�c^e<��Vs�5ERW���8�ubo����_8�5Z�NV��b�m��!qu`ϴ=� y�=���z���L��C�C�5=5�2k�2�BT���4��ӌaOԮ@o����f:��j�B>�S8�f>�� ������]��Pq/�$��e*F��HA<�/h*��cT��}��:��M��@Kn�i�\�SG�e�J�&d���4���ǗW���'���w���{>�F$8�