��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����G��l��"�Fe]=�/>�"�3Nع}EJ0���U4�q��q��i��[�3W9^�LU�3k<�ҋ�͙.$w{�d#?ŧ�.�&���\�FaAG��Ƚ6�o�� ~[Z���~s��c!��ء���]N;k����h ���ZAcd�q�4S3�*S���k�!�[�>�Gf����tZf�ث���Ta�z;TcP�.�Dz�Wt�'�KC���h�����D�����5G�j~7���w�q]M�����u��ɲ�9�#���ƈBt�L�Q1.q4���v{��і��гX��"K��8Z!żD T/�P��x^�அ�#�U8Kr�%��;��<F����Iv]ɾN7"��x�ܕ�R\�P�~`��WI>Ru���^�Z�W�h�1�p�|�P�T�J�����(�S<IH���sWO㶕��oЬ�!��ɍir4`�2�g'��6�$�U�z�µ���3��
<�o�C�k�Q;
(&��^ �R�p��p#y�̷K )!�����<��+�ϲ}�*����� �$?��F>P�O'�0!K���.���OL�^N�]��q��#лKj�s>+c(C�<�Ŭ�8@X���4@e q�^iJ3�r������2U8��im�b�O��`����.I�S��~g v�$B�9GK�����-;��}�b�ah]>	���h+'��`�A\>Ƕ���LO6��$3&rW�!CH������9=��~fu����L��`JN��a��E���n"mD��R?��I2��^�v�Q��Y�'@���k*EfV ��3���6�kC�$¢��|�=�md��]w���@��Vn�bB�ߛ�=Fg�3��27f|����Ya�poy�j�5�8[c���r��G�)G��Yi�Nt?l����w̉ާ�__�b�M5�
�p��*
�dqh���׬�ü�rA5Hgc	=���3��\_���?�K,�D��><���S�%4�9@X�$�Ƕ���>�Uy� �C�h����[��SXh�1��;��u	��}���H�E��7�����&�}���J<�G�E���]��fO;��[�1: