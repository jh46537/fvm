��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���c\�esR&{������o�T�e�Z�/��`%�����1�2��g\D"[ޏ�FH��O������XĻ
��(3�k���]&����.=��g��,�4 �Kz��%0�#x�S'aV�?ϳ:�7BX߬QqQ��SPw�>P:�Du�χ���1Ӻ�]���fޡ_֢�MEW�i���ܬ��UT��)id���Qq̧��^�k�>0���i�dn�#g�9���#V �,�)[�n,S0��	F9�A#T�:���"A&[���g�< 0���#�m���������A�G�&t�Q�����@n���^lp�"tPNWWQ��Vu	2��0��.(*Kk$��;�Iz�f�JX�H�#"���g��b�<ԧ�]
Y��GrY�� (�V���9�C�T�a�9ld�V�*:3��O�rH���!M�oi"��1�_�O 4˒�v3�	�4z�;.�s�b.s�S��,��D��?g]�$:�7�J���b'�5��i%�p�}��%��f}ISV#YŰO��*cK��XU����wi�Tv'�����J��K�89ă)��4����]N��^'�i��S9�r{3<� ..����|P���G��!j�<�8�&�U!�};���5(� nJ�}3L$�6Y�4����c��s�G�$!�@.u�W����zT�W�7썇��>7�1�a�j'�y"�MȾJT���+3�|eK�K�z��.l���AO����;b��+Q�m�{s1B6�hE�}*��T.ƍ��lz���E�ő��̼:���ůB_�\oh��F|�����J�Qm�źo4�eu�4v9��y��v�S�kn��(��"z��K)]�w��H7�{s��d��)��.��b�/^��e;�U6d�����}w���<��Pb��b�5�����fOƏ��ʓkH6�b:��3n�)[ݮ��ݟ�b�����R%�����}x[��Q��$lYܰ!� A)�/5E��G梋�^���N�S�G��O �ڙ!244���"9;p�m 00�7�E�FXL͹W7�H]~X*�����+����x�q���,�9���O�jTY"�$��<[8�[�hY��Z`�`NȃC������)m*Y'4�w�p�Y��'$���x�_Ю��|��Lf�8}���^+y��yţ�A���q���=���Eg���գ� ����CzI���=��,��(_��AK�r��D���_��s�څ6�ˉ���H���Y��͡d+�F��^�R�In�L*��m�Y��S�!O�0�?HU�ޱp�4��]��W�Yn�Յ^�0���^C��,�h���uZ^q��ы;e����f,֥�jQ��5Fl��Ď=�����60�/�F(mrZ�ľ���Z�U_ 
��mv�9f��*�SAL���[�}@|CS@������Iz��)�u���N��%���y �l�j��~=И�rF�<��60��9=�^�A �2zu����_���P=��O��E+�^�8�+�^�bj�<����Q��i�Lɦa-ۢ��ێ�ZjJ��(�p.�V�	���T�(a��_���L�2J�Ht�[�x�/k�t��Ѵ�nq�t���.>:�,"+�p�\E���r���#U	^��8�B%�#Еć�p%1�J�Zozi���!�wR�
��Wkƅ^I�e�cEM�=�4"Y����t�qX0��ٲ��1�_��Ğ���܀� ��]�@��OyㅋaJ����8/�r�o��J���+[XV1V���2�I�,�!�&5}0��?T09��FtK����[A�s�{7�����^|���ɫ{�[�b�j��,l<[}V�ñH̬AN��,��n����Idߚ����eW|��V>#�IP/�Zi�K(�Ё}�*xe��<�ľ�qŊ֬��>���l�8�>|��8�������UufY���%W����|�v�Sѧo�=i:*��̰������D �4*�cj�C�)Y>|�R<<��u���<A�枴���D�����=>̘!3z�u�9�k�NK�	���nS�?�:����2C9믃���E:�`��_:
D�i�X��U&XEZޣ#D�	��缔��.��/eT�K0�-�Z�ʮlCXQ0��(D�������i�t�t=]7�V��#Vv���^_�M}D `����A`v��u��^5�E�#��a4����ww�ɨ��d�W���z��\���L#��b���{���OO =�V4�b}�4���p�ylr���d)11kP ݫ���̩~����#&��0��`�Ki�O���${��	��vbO�p���
φA�����ZJ�q�4��N[��*��R�	!��E���qD?Ή���b �)\��S78R C�'ژT[3 ���L�=�|ϦuQѸ��&b�J� i�z}ؚ�h�gۢ%��#���[�qJ,��4/V�F��} �Y�V�
a:��&-�<�LA�:)�맸�T�͗{\��E���1�'��� 0br��!@}��[�Z�S��Ŀ����&_4��g��YQ���H��8n����-����M�"�h2nj�xK�Gy��E��+��x����"{�������v����l�x�F�|g�1���i�3ThOc�j�VkFu��Kχ:k��U�dEԼ`�\=�zL�P�\�X��s+��5�f��H�*�Ǘ	}?�[���4{���V� �~�����)�����o@�l�&Ǆ��0O����oƦNd���)ި�sTO9��MY=]����M��.:�U%��{b:2���I�Ǯ,6:fn;�!ف��M������-�XpY�T}dgL�1�^���R���`ƚ�/f��y�TlR����eH��
D'|�z�7������+���L�VR|]/UϠm��߂d}�3����L��A�|�t���H��{�_0���Z?�(�j�uK9���Ž�t��{):g$g�j���Y�k���j��g#Bi�oM�aX{�v���GNH(o�~5Ǐ�s���d�F]�.x%�i_�RK`
���fD(����k9ZЯ����:����J�c�z�Ə��WW� �T�Wnp%!�v�-�ٚʷ�Bb���9;�S����o5KcB�2�������Dh�<����n�٘1L����7�ͳ�o�_������`1B��
`솫�M�>��l��R�\���c�>�a1�v �@���ꞈ{��&�o	�H�]Y�������@W����<�>Wv%43�T�8����n���d�@�2�i�,���� �Mk��rsG{
%�@��az����2qӌB����q$ەQ�Lt	�%!�	�|�G�%5���-w~�V>�9k���2���%59u
��<��Ʌ�����/�[��;a��� �3v��=:ꥦ�\	"�fwfȝtu ��ZN�����;<e��=# ���A�S�)���,��V<��0l��*��>[(&ۂJ�O(Z������%�VfBD��=�^���f��w:v���|'�ʷ�����s����Z��G�_��}Ξ`�/>�+J��+�u:<}I��/f=����bɞC�  \x21�ze�,���Y����ɱ&>�.4��y�6)�r*��m$d5��x�-�5e�&�Ͷ�dh�7�y����f��"�A�?I�Y��Y,���U�<�Gu�;��?���O$�I֑B���r8r'U"P�F*npF*_��z|!��Lc�Z$ҝ�?�%�Q�)S���m�EXI|5�hA���\͒]��<CJG��MO ��ٺ=�Q2��f֭y�N���0?9E6!�gH&c�����ͧ	�>S���Z��6�.�'�a�yq��r���Vf]�veUF�,���Z��ďBe6�<��� 'v�#����:��Y���bu1"n�9	UOS4)H�p��g��
�!7��s�iv�Ol�[}Q�# ��c�Y+x:���k�8fzQQ���2�\�Oq��zb R�a�l��1e��
��$��=�� /5��(~�l3H��e]��T4���{���nu�2d�����:X�S��/��m���t����QB�8��[*,;���$젵��oo$km���-!�ZX ��u%D���[�-:�=E���h�:����:\������8 �T�{��s�+R��8vQ�UL77�_-��2lĻ�.�e]��V��ؙ<���U�U���9~��.e��!ݽN�*�Z_ˡ$��wCaO������Q��-_vU�T:;p��y	�7i.BWc�ZX���p��&$��3&�A���!n�ԟ��!�cF9Lվ�Z�
(V�S�����<��=�)�
�����g%�%0��`�17%6v�'��;1�Z	oR�Y���SB;�S�-�l�?���+AT��e�QiNHӤ��g����H�+Vզ$�4�����\*n%ʙp,f�J����,"�\-���J��u��y��?@�_����+��D)M�F?��7LD+BeE���=��m����N��Auu���S~#�Kn�@�*�Ղ%V��d�'9
]t���o E�O熜����.>��B�I۷�����+p����ĩ�P�n���G�\.v3�e'��Q��,o�y�uY �?:��l�~��:?)�Թ՜�r�F��Mye�"������[�>S���k�jGк2q�����Q0���%z�zQ�"lD�Mޝ�#�!յd�Nqɻ=�B�3��1 �C�Wr$Xl�;�Dy���3�q͘���P��n�nc���`��r�D�6*V��ӱ4�x�����8���n3��|'����+J�S@C����T6�>���l�$�t���bo�U-ܦlA3}�a�(&��T�؍"_p*.;u����%8���}:���5���d�o�r؜\�`�,��>��Kvzx�:D��֞>h� ���PE�#�]�ζ�~����5Ӝ?Jn��T��ź|�{�`a��L��Jo� ��j2�sC�0�X��غ��v��8o�ދ�Z�^�9`p�=��o'�gTlW����We=1`0�2:Ȏ�/��N�_��$��Q`rJ�0!D�����b��I��lHK#�٬�^7�i�q	R���#��>l]��(�rV�ρn@��#��^9��uڝt���f�E�~S=�v8���~в��b�M5���	�H�L���|K��<�C�((���reN^���ykO�p�]��=�z2�����OT��O���+��;,�b�@�����k�	�UGf�3̴��8���;��gH��]���kH[��&���8"
.6Q.І���q`��n(?aM�aL�ǧ�g	�`�vW���	G�b��U{��.�� ��nZ���|[��{�ݗ��?�t&Z�����Z��Ys������ˑ�bEWl-k���Àm� �S�=�xH���_�b�����_"_���C��	�j#���ɦ(1����W���Gl��:��g�x��������C�w�=-� �n|�:�mm�<�gq��.Pژ��h=V:��Fz�8-'���Y�eut\Y�Y#�>�	�`R��҆`"�������bǷ'O�	���gi�Hk���j�&,1 O�.��Ct���3����;��b��y�4�[XX��uΆ��o�y�����Օ�>��+$pN�n���$�dm�����?�:O���T�1�ީ���&Z,b��a p��g��R�m�ίk��x�z�����%�)�`�p� �����/�k�k���C9T�m`cLe��H�w� O�ژ��M�ѭ�>�����w�&-��=h��y����i�i�5�q�7���m�M� ��It���y�IC��Z�*g��[�m�2pZ�\e�3���[����4Wr��w�r���� Im��k�}�H�����Θ�����'�/A߇�?k8�_��8�s41�s}�u>T-#��y���ъt3�I�A�����!���M%	��}���9����~�	�.��")U��g�?���+é�]�E�i��%J(i�]7��: ��%�$= >{�?����OVz��o6�����U��_��� -�&�	L��=�!�sɃ�;"6�)�L0^"���D���~[��e3���u��e¥	�Ϣ�*��C�qAd�ǒ�He�+OlD��l�
z����@���$+�W?���?$�=(<�L��T��g�p^f�(�څ�U��������֋d�7�����Kp#�,���g�}B%�,�y��U54,8~`'���w8�F����ZG>0�~4A
���Zb�?[���ۯ)����q�34�u��'����՟3@c�U�d�/����qbğv�x�!˔;o�uc��,g�9eC�}�	~�����vˁ�눵�s�:����)��������)Yp�>]�����Wb.5���\��u+�e4�g�m���F �t2+��7���9>0��L�t`�ܭD��9��mF���T!��F��<����R,���P�x\,ҧv���$.*2͌(j���r����:'�j��%,=ܓ�b����;�����j����g_�[��^����$f���н�Ϧؿ��oo�s���b�)1��S���_���Ҧ�t�0#)v��g���>�eV!�*gJ`~�3��g�3��}�r�[���:K��:��u�F2�/�NWy&� l�k���搤��*E��V����Xwآ/��y
��ϮM��N�sv���HS�9�uS���Ƀ�,������°�t��?��	�^5���`=i`�c��
Q�u�����Z�mR�v|"�E��� %��(`�4���K�����ߣ�w�
y�~�M+��̤~���`����k����|�7�(�3?���� ����N(��%X��z|{i��F�S:-?z	#4vU+����ՙ��:�-���dA��aV���*T��6�eW�f��[7��x5��gE�\#)
,�
�����ӭN���á����� ��Dɼ҃��^*�	J�7Q��3�v���ڂ�1������ �涀ޱ8?�TaH�mQlS7:9��C��SD%����?3� öu>�7�>�,�@�)�2�!ĳG��ȝ@��v�u�ț$>�ȑ1�ٙ�Entq�7��EӲ�ř��b%xsd#-���2�X8t�,γ���z;^%vo�@F�
����K�L�{?r���_�i-N�$�����Θ�L�M�*rQ�AT���Q��u_��;���}[�o������Zs���7�@֟o[v>�n� z^���&�@◵ ���n�K��$�bLrѣN�����w��/Ё�M�~��w�nQ��=��f�{W�9�^�����QG�oN_n���NU%�!"u󑔠s���v�ƫ��DH7��8��I���I���g ��*6��yD��ƅD���)v��Πn�r`d���ў�+�JE=0n�Iu5>�H��?��q�-쇑�0y7�p�<�{��WS��s*wN��m0:���3�{4v�E��i7�-�yW������e�#u��A���X_�q��b�u���X��}?x.�;kUB�N���=�L�%���?���pʠ4�rG)�ʗ�����F��:���L�54���-Dȡ�L^�M$�c�s��{^j��
�2�U�eq4���L�_��l�a������p}�l"�&c�ݠ��{�ԇl3:�� �����h�- e>��4
N����0QJn#��v�'���t�<°䃐�P�a�>?BYwݨ���2��:���$�w�V�m=A�H�܍������<)�[^Űim(t�&7;�C9��H�k�s�\X�	� ˡ����^�=d�$�Vq����7�����^k�_-�v�S�*�x�hK@�:P�Q��|�{��;����������]o��4����s��Ic�V���:Z|I�	�����l:���Xj`ݣƂ������|�o�㏝h��k������^����`�}���%��q�`RA��"�R���^Qw}LKk��d�DOs�sG�;0�W����Bk��j5/��&���;ێ��z!z��$�)[���5ӽc�M��Ə2 �MȄ��i��Nb�R]Y	�����V�Xk#��m���ukwC�����vo2�c�F���w��}c���s4__N�"W%�"|���~��濲�0,�$�j{L��$�@���5|�j�C7���V a���%W�?L�܌�Ձ�3����n�J�V�n��&�1JDo�Q�qC�nv
\K͘��X(N�ƕ6����o�rD����iI����fmw��J� �/b���f�l�$~�&�o��=�cٸ�:�Y��rU�}s��^{�1��<
�Q���<MA|��s3RVF���y�e� [���aل�k�؆��`Ûd�+���!ꊚL+�����u�����>�X��~G�F�5��@�&:w��f��� �1�?�̴K+)&���3\��3�AX@'T���L�������;�i��B��{�5���T��3�ҹ7��q���h2D��7	��CI�H��n�ݪ���/��Y�!�nnSK�� �cxQ���ÿ��}��q��q;-G&ag��+?�#���S�>�ꑉ�V��f����s!C7m5����{ @�4m���t�v� �@��e��'�{S�U�7�}�0b�^���M�)��aڜ��6��+��fϭ.�
+-�n=A��C��ȉ@ � ���3/�I��D�SeI���9�a���j�R�~��/�=���p)ch7W��{bb������ʬ�!;;J�2�w���h�/�]x�v%�H�k�;0�
)��N��0��R�����x�Fy��G��m��MXRQ�e���wӏ�0v���� �8�"�R�y�`��#o	_�	���Q�#�m�L�f���K�{�s������ь,���ӬR��h+Kɲ�ؓ `n�Z7wH�����y �y���W,W�$+z3� ��3���N����5�
�jٌ/Y���V���J8&���c>�<
�>n�LW�!ɀBDAe{u&Vα 1M`�Æ�c�/[\������7�F*��\��iqܩ��{��Մ���s?{�;�ƻ�,O��Z���,�����੢'���F�i�t�t���k�@��ҫ��S2��;c;�dOª�LJX;���&\@�����X�L���io8|>�'r?q��B-a��J&���<`��'�jO��Ŕ|$Y�m�bJD��?y��$�q�G�m��-|�v�,�ܿ�\����bWz�;�s�!Y͑�W��v��y!��\&�OŃW\�GM��j��r�k�-c=B������+5��lA��7y5��+%��X�K3@ý�(���
���ⓙ��-��:�\�'��n"�k�z���f�O��' 2yoz3y�I6�b��%����i�o�Ȅ�-ċ�6S�Zz���_]��է���P,�η��{�:�Z'Hʣ�W�c�`�{<���0OSk����1�����_i!������5ז)t�rZ�ꩢt$�m��� n	�a!:H����DL`�4�Ͽnңਕta�$�Xe�Y�|�^_�@=�����R���s��p�|۬�{��u$y����@'�~s��Ǳ���%gB{���8��UhE�ZrW�-��,��_��@�U2����a�z��a��,���C�W�.X瓫��V6>�..2���<W��m<�ƥ��T+��l����$��̪{���~�
�ߊ`�gvS��!Y����s�*����P�������(U�\3�o�A�W?ٛ77q *r[Gi2�p�h��� ZO�,}��d3jI�H �Q����ɟy���MR���$��_�ڂ��=��.YOVwZ�˞2�L��GU,�M��pi
�Gx�	�/.(V�Đ)��7t �;�TXxߌ���?�ڹ,�讠Sz��T�(����Q�p��Hx!V�%�&H�ܧH9�K���Z��Eш҇g��.)�� AyÈ�(����4e�hb�*C���?�`��:l����N�i1�ϵf'&�R� ���b���N���3�S�$7����H���Ts^������Q�߸�{@d��n(�-%4��2� ���W]�2��iӉ��7i�!�]���ȼF��) uu�
�Ć�����,Ax�'(Eij��*�ڽ&F⥺/Q��ܡ��-c��:��[��\%nZ
rӸ7!�J�)Q�8Ԅs�#�+=��<]�B��^L����F$|0FI�bW���+�3z��l����6�����_Z$>�ad��">���²z�� ݬ|���K� �L7�<��G|�|I��x�2HO߳4;L�4��s����a;n��K-|7�����X�vl����dS�40�_�%b��26�9�#B�J{ޫ�H�~����S����.v+�l ��<j�畸�^�mv���,,\��Z<ؾa�u'���Y���ǎ]�ky!���M����>����9}���T"u�qIϹ}��y�I�w�r��yFz�fUʊ���j̇o����e�Q4e�*�1H��7��41C�sKN1g�Ňp3�&�|Jj?�W�������v�	5�+k-֔|�f�������TV�2�U��݈�����*���/��+t�4xcP�+7�b�`4O