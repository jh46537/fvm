��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�GG�mV),AeV�İU"�؉ٲ���B �mH(\��2��2*�CM�D�|��j���7v-7��a{8j��,���U���ϹJ����Ӓg�1���^$�0P�S+�S�*����dz���7&�h�V q���k_�N���֛?(���l�r�<Q�2�� �utL˱a�@R��NH�@�:���ǠyZ�|��-V3��������*'Ca:��2��#,�㉴'���2L�՗U*�1mU��BI�l��h���o�ot����h%�6`e�-(���D�й0�sf+����z�[���������1�[p�[���B�<R$�2k�����4_BɊ�܆��=��6��j:�U���?F5�obzv�ȍ���|�?�{��SI\�6�h~��HiR�mH��&[�p��G����5��\2`h�9q|�Eg�7�_T۞�4��e�Y�A"ntL�=��q�Ɓ�������*�7�jGZi+��n|Խ\
\X��'����M�`��#UO ���;�~��]L�k��`m
C��j�N�C{��c��86'd��b��-�W
j\ϫ1|����ƒ~�-��ĵ��.)����&U��M��e�_ q_G��ď��E��*(���̼Z�n�x+�𥤲"6���6S(ɶ6��c��wd�r5��^�s
�m�v�J���q�Ĵ�֮�:�Y	�M�E���@~��Ԏ���E��ݹ���Qc��ۡItF�Ӧ�D������7��̤^ti�v��zl�Kij��NҍZ�ό�=���&5���T":rB�3wD�e[pXr3��e�ˈ�9�J �,T�\���ǈy����"�_}����36��Kg)���"���@|p$1� f����,�Lk<�x^z���L?֨*ǌZy��7m�7e@B����<����k>$bH�K'{���\��Q��ܔ^�o�(򚜇���pw����Ahɰ��<Dh����B�w���NE�1�	K�C&�7��G�ZSd���սn��҈�s%�r��2��Y+��Z)
�{�E����}VU(���Z�c(��[>�Uv/�|c��-o~�f�De���\d�E�����A��0�A�:0-O��m��a�	���Bu��y�8p5�
{�3��4H��J;/B
o��5�B�"����;����i2�i�)���l�LV�'3 lK�W�I�e�!A���P�����W.�
܃97�ڱ7RH;���UWI�;��6T�To��ܤšj�}>q�n^sW�����(�v�ѹ�o�P��WR����Ip�L}�H��Q	Ma��P����m"֒S	K��q-�,�}�E� �ʯXl(���#���&�k'h����fq/��n�����L\��,Y�!��)�����23���hfR���x
F�I����Ҁw�zk@n���hW�V.y稿̿�s��$�NڙJk�lgr�=��8an
2�p�x���G�gԇ-Y$t�\2Ɛ�|m���5�^���Ӛ���Fc_|u���^)�Q��k�����Z`���Z��,I�n)��>���)U@u<LE�_�<�e�� ]����W��]�\��f�@���KI������y���`!�4^�,ݿ���>]f���q�I|��2���!p�Au�5�f�>K�{��Ir�&g}��uL��dZYq��l�q��Djq�P����`�:޵�xeÛx�Q,XZ�3_�X*�2�c�n	�Mo1������_I�>�Qa�!���8�=�����e��TɹW�Xc�.�E�Y�AUٕӛdpbȂ+�Jb
*�*O���yUY���Zki��vz}�:�����/vKKפ��3S���ݩ�Җ>��N�ü3�7ܳ��������Ol9}��4aĠ��zQ�r�Lgzo֯�/�cd�'
�E��1��[JS��3�f�ߘ`cйYV�>V�S��a��C��� 
�B�������cJ�]n}=�'��}��]gI�h1,3�Ј�	�\�R/k`˥�hxn&�P��)�D�5��v�Wܠ�sݟm�ɥ�P���n��D�G�_��)"��=a�Ejs�n�e�uRF���0G^h�ܿ�j��_|?g1��Yo����F��ׂ�cĐ"�[]�"6����	��&J�7��f�qU*9�����H����;��G{`bq�����-��h1��K'�8�# Iz�,	�t�R�-m�� �v�GоV�a�W�e �p5���{�,�=o�1w��bk������c������n9ơ��>��h����q�G�GA�a��gf�Y�� �I����#`���͚<��6unh��d$���NT��nq,�G)�҄��~�Ov� X����2[�Z��
'w!~��x4���U%E�����e�
	���s9��=<�TjNfѼ�����C��Q<�IX'zڽ��T^�dF��p�I������3������xف<3�x�F�����q�W���۵��2�E�FV��W9k���L}���(�C����T޸$U���턇Ik�S�-ѝ IƗ�L�o2���CK�Ր��#G*��R��*|7��w�j��(�:����M�l¢m��T����V�7����r,�A�.����nj��kk8N�z\×���u��J�4�t��Di���WB���=��0�D�E�j
hRJ�P�>��o>7r��wDKd�U5��]�~��P6�	��Q��p���P�ᬓ?�W��U���~��$�m����3-R���r9"�� �4ЛJ!�<�\��aO�W�>���P�f𯮯���27����j�C��l�+o�l�°-�'Q��Fx���ن%�ө���${N�Cx�����#��������Q\<<'<嚧4^��g��Qj��X��ep���7��6�6��~��:e@�&�?��k�Iˤ2�0��ط�P���7��� �G�K����[�b��M�?�Q�W�D��=�Wŉ5�{#�'DP^(�Ŕ���ƽL3d}}���1�,�}m�
�}c��ٚ��[����S����hfr���q� 8����Ʒ�a�>�M���;^ O{c!8�_Ú1������a���]C��$ FwD��,��m��@���/�W�S��h���4��< �[��G��!�ϊ��v{����! A���%��^��>�k�A�p�Ru�2�w�Z�D�Rv�vB�(���E��	����9�_C��O�+�r<��.{Oj-/WX�d�1�Q/������R*��K	�{uV�z����Ow~fB	�T���1gSN���	�x'�1����������l��\�N�R/��"<ͯp��u��Im!�X��#h�)���� ����K�C�R���0��M��cfLJ��U�o�H�2�˔�_y�w""T�S���=��vs�v�8��	Тa�
�L��O�?��h��h���^s^l�w�m�������J$j�.N$�-�$����X傪
7ۙ��_�oz�4��Zg�4R�@`�[���k�<��R*�{X����G��<��V���f~�h��r��H]�9�b�9Q��o��>]^Q�(#E=���!��a��ݤ��@�V� �l|Ib����m�z`�ٯ�8[�Εj��Gj��.$A�|�W���f���X�Ec����zd%1<N�G��#�[��<�W���lJj�ޕ��֭�KO�>�}K�p��Ϫ^�"������[�3��	RY�g�RK:�kW'�������!	��@���'by����6�b��Tޟ���:x�A�)��t��0C�T��0�_a���1O42��\����@j+Y��3۵�#��Z�Hxe�yM��Lt�R�7�%p�.���VBb�ֿEF8:G17�2h~ƺ�&\CkfnL"b��&I�,��P=S@�o�{?�5ˊ��rW���m�؜B��"]�4�;��W|=����z�xy>vn�he:���cznb)�:¤�kJ�c�n���7�B�qT�b����s�r=�u=��2��Cr{F���d�$̹�z;Bf�i��M��/�MN�#{b-̻Eޡ�����3�^g��N�3��dFYN�.f���=�e"X> Ku39ɔ���4�g��u��%��>�|��/	��j�˕���΀x�G�d�j�R��cR:v
8��W}��߰B-%��n�T���P,3R��eݎ����޵Q�d��/wA����:��V<�@u��}������3w���'�¦H��;p�2���fKj��0b�'ƣBĎ��R�\�6����ov6C�H�)�i�ᅶ;2\�z����E�����-�#a�Z��7�p�N�j��U��}|��'dh�`-��<�˻@ʒ�x�1Fܶ���c�gr��9s��<!��L�,��+�F��FK��?~(����0MR�<��8�cO�5�H�gp�6��ۘ#�����nB8��!��J�͊8�H�߽��+�J�H����Ev��DyX��T�P�	�ON��#�����/�4+�+8?��_��P6|�]��X-�&��-�v	&�ڨH>�럋�F���u���ar(Qf���]�hlA�g�l�نf�A���i|8�B��_�*f)�߱��=�v�+�Y V�O#vh������ȴQ��%`	�^��-� Fe�Ub��d�N��\`l3�m�(ƛ�8���l+��3o��zo�x�c!(	�,p���=��fve���	�w������t�X�	/�,��l�!����yV�y� 	C� ��D�����}�}V������x��� �����9��֜�����hg�.=�;)'�U`S���\afe��u�s@��@�3��"_�������k�c�������a�����
���K�f,FQG}���t5�+T��q������,Y���~��Y<<�҉R)ً}˞ס��]�rah�����ѭTK��BȂVϳZ��)��������+N��Wߎk`�������(E�K� �3��(��N̓K8K�Uu�&��S5�-6E|��\��*V�,�������.�؆�������;Mf�Z��F��2f��y��y�詪"ϣ6��Ӱ�V��6Tj?Ý|C'��u^o�KLV��|:"x#����,,�F$���c���"�k�LW��g�H�*��$b�s;�(=w`�Կ�+'�qH�����������v�3>�#�e	�/9����8�L�մ�ɂչ.s�0�ꙑ��1Jr��`��e^fs���<]�(m�c"�Oo)ą&�$��23)���\��ZD����T�]�[;�-�@dϤ���e��q��=_�N�3��R�:%ȳ�h,���v�y!��P+
. �-qMD��`si��K#��M5�n!�=��yeC�d�����:�\ G�9QT��%�v��-�dkҿ�t@�ץT>.-��,�����Q}�?��{��t�ުN�R0�L���8�����[cG7s!ko%->A}i�`XR��RD��O��~�5��J���U�ZYŁg �T)g;�A����2�sMcza)��l�#�t�s���uLkˀ�ʨX��ʕ����4�c��3KZ�DKM�W�d��<_P�(��L�
�����SO���0;�|Z,�Ɩ��щ�5�fV�q/�o�B��-���?�q�}x���p�֓��D�M���Q����?p�h�m
��8!�怞0A��u�� �53OV��x�I�-�u���֖��P�lee]�7�@E���$]Ei��Y.)�_��ާ�v���ȱ�;4r������_�ѿ�mM{c�z���+�+.,S4&l<��QN\Bт���1��p r ���#� @�r��*=��E�T4�c �o�N��o����`���Jb�𬔷�����)���8YWlT�=���h�n�.���%5�Dv �(zK�N�C�=�Ҫ���}�Ί��/B�U?4N*�icK��,-����Xa�A�J�r�k0N��;$��=�S���g�A����Wo�>���m'&��	��i^�j���ᐒ/�𧼴���� ���a!�a�!�W_�[�tT�|qx��6�mZ,�Y�BJ$�*�A�"h�(<��<����p����b=��ݗjYx�7���� �Jy��ryy_������sxāZ���	�*
D.�N�?�l$3�5
�"<P\�`��U�ߩ�ec@���Մ����9�a� �c���Ϟ<'�v�P9�/0s���HS&��.։�~��Y)�B�l_�X�W��6c+�CRK���_${�0R��7��N*E�����l�iȚ�ZQ�7x���He"�Qb�cDhg��~�%���W�`��|qQ��ø��)7��ys[6�TY1��6�x��?�~d���hԙ����>�N�)�3L��:���G�_��϶��)�����\^��<#�Tb�y���tx�P��l��o*Or��ii�r����~������΁�M������:�6h���ϫ�0Ӭ[A+�Uko�}��1ґ��\���
���P�<���R��.��� ]���J?Et���]Ւ T��r�׳�	�k�h�V�� b*HH��uo�-~�#6�y<�I]3��Hj�]y;8��Z�zC�'�3?�^���j�P��%�ſ�I8k��1���U$�`�r·]�8���1r�%~����j��n!`M��K��P��ӊ�"�{��W�Y�$�w���\��|�9�J]��P���~Ӳ�u`ݚ8�{BܢcI���$��~���y�Ş��Jj4,��%d��(_M��eZ6I@�f��Կ�:] �I��x�<�����G�!�"��H��,��+L_��+��/��Pq�����rd*�9�Jp荲-�7��Dy�\����#��y�zt�L=�f�)�Ƌ��Q��⺝�)��2�i��Iީg�� ��6j�  ��M�8	=�ѯ�*yv���J?UA�ARD)��&m��_쎬�}^:������׾�!�d����;8.���灢�2�]�Nb�S^�� ���#� �AXK��8���i#��Ǔ^��	eI?1W��Օ����o�^�{���J��0��뤮bX����-/��J<NS�k�o6ŋg�hv�Gy�	�����^9s�=����?c�Z��J��OF������
I�#��������)�S@x���!j0���.�a�`5J���j]ᲀ�����{��S�3��/��K�Z%f>�rX�#��sf0���"8��h�>���G�*dY�=�49�{��1���P \���Hs�*�m7�^��9��_#���k������~;�"Q�l���Q��h����2 �;�0?�L��8	:��-٤�+Fĥu�\=�fk
�Ւ���!ߢ.��P֦n�,`p���>���4_8�C���}��1u[³[��\��=n�����R���w�.H �&���Z�h�ۭd.r��G{ ۂ����/����h���L:��C���Ys�@��I�D{G�Q6p���+
���q��D�^�/A�ZN2��&$s��iv����}TF_h ˓�]�(�ElD!W|j`��9U��V��td��$�J_9E�U9��N�Ӏ����? `���q� �ސ�}��ٱ�(�mt;�eM�D{kcrt��R
7}��o��Q �b�Y�/�n3m��L��y�'.O�����M}����-�c��%_rQ}9�����l��o�VV7�D6��3d{%051:�_4�j������!�h��ڒ\:�z���x�l����}��['=S�6X��h���h�mo7���"k���e��FU�_Z��q�s�� gx�ٔ�s���V:��w�Ԉ��;��K�^�1����eл��9h<L�, dB��j�K���"H��h�~����e"1A�=��4�'��W�n4�/��zLCF��6���X#["�^�8��]a�x��p��g	��3�q��o�tO����J�K`�O;�m���v�r<{*Of1�oR�� 0�+��0��Ί��h��$��G�i��-�C7��Bm%�΍u{�>���-d�a+mǾ!��d��'-wqG!��t	����4��j~I'�[ְ:c��q�J�o��/ψ��"'������v���R�Q�Ȗ���{@���1�n'���U����7��E_��u�&7�i����!�(���y����R����7���Н��0ӤZ�\E����8ne�b�F��D�r�e���΃;��{��z�b�oj^��f�T��S���R6��p�@>�_���Pw�g!u��~�ϫ��P��1����{+�|zVMd17HIy@H�yh��#��(�~���4�u�?U�f@-�3!�P~��ZYAV�Jǐ�/��ͻz��+wpC����b$I)�}�ᙁ�[�a}��	����K���
0�:ۡ�}%϶
"/������ߩ#��r�Tܽ&*Ǻ���� ���{���]�/?L��+�\�\%�>��c}����ʳ�D,�)c��Ƙc/$X"�Ewc$�Y�VK@	���cMY��B�W��xy�o�jj����h"�p0������Kh��9����� �ju�}�aS����{]��E�* �g�e�X���ׂ=I��1 �E��og%*���_�w�b�[�}A��\P�"yAGtn�dO�PK��_���d�y���:��v�c(��W�9`B!)��u2�,3
�F�*���L�ٮr��z.����%eA������Y��n�����kk��w�͓�󻒶͞?'U����bN�����?Q��2�^-Y�p�e��0�<�y�L�<m��Yiס�m&��I�3������.�;�n�{�)�f�[�d�Gګ�F��F/�������X,����H�%��U���TW:�����ߞ	��� ��m������No�Ё	��eL,�@���:��ߧ��s]���a�u��w62=�ИD� �&�?l�-�0���GQ�S/x=I���1�q���='�+l�6��}��7�{��i�W��_���LI-���;Q����pG�|4��87���,	������q��
�A:�fyd*9�kJ�`^/1�yNY�S��^�����yhgl��6��N��	:B�H����Seb+X�4���A���T�]C�o�٭��v�ǯ��T��� '����P �)���%����=���XE�$����ZW*�K��gO��Z�a]H�Ri�뇿rC�+��]U>��oL0};��+�E�H����[�s ϡOv�w�h21"8d�^?�S呲��$�Aĺ'7WNY$V��I��]�Ql: