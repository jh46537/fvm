��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�0�w׍��SΪ]�����E��>��顗���="�Ct�QJW�����j��I�����1��5\W�(�V����������<l��ٗg��h /4Bܟ�G��Ls�_��q5\�;N����|��A>���X��/���d��x_�{ɧ��������q����5���2�a��(���RgvZ9{�����m;֚�h�&�L+#.T����?��M��AYmOoNvG��$�b�&sZ��K<�E=FQ���[sM�0�Dߖ&u����s�*��!c�R,���:�-<M��:N��ʃ(���6:{����,|�����8��.�}���t�J���?�)8���B9#�8\vVKbo�������&^}:\��+#O���T��!���-`6��e��T9��ų'f��(!s�^Y�#��$2;����I[#���N�o���+�~��{Uv���Ii!�H@�Q�~��J���G�~��m
eOCm�C���
�S���r�'��`Ԧ���� �	/Y�M���)��F���$e@u����"��R}f�,.���(�d�i�n���ݴ\�Ϲ�
��@Y6G̗��T��������ѥ[Kp~���~�+�`$P�{=>p���ڇ�4��q�����V����ҁ��ꋑh�uo�������Į���Y�ń���_B�/c(r�&@"�+�� ��B�߳��q9�ηϏ��,�� ��;ƭ_q�h>줹̇��΃(�KÞ�W��8):8��1�k�)�Q�S9��*7po1� �..���N��)e��
�h�fb��v���ΣmkF�n��"�F�E^dt�ı�8�`,��ͱ�n�Dǫ�0e�=\����<CB�[7� ��r|���B�q3-���]����F��h3˖��br��H�����f��(�Ԭ��<�[*'����A�a�~U�}_�u�4�coh�=�<�������f�I<�g�`����CϧB!���`��.���K�w�-�Թ�Uo�ʆ1�c�%Y<G�>\[���<縴E����Z�,XH�;��-�,��G�
_Ko8����@��+�.�Qݚ���7��5�4Р���!����հ�ϗ�]eI4�[�j�EﱦW��㪓��(�=�)����C�C��M�!����0T���0���4�0AY��4�I��������E����6ZW�=����j4%+�N]o�/���SMV��+��Kb�X;�s[��>�l�Ag��tqc�~(Yck��MWŵ[iT}K���z��`ĵ#]�N�n�9�
��f�Βg��./�xt�����ϰ��n���۟_�b�.	�[	����$"g�ȹ�!���ϔ)-��O��y+��+.��y�O�WH?�3e�*(J��
����/rq�l�&�;�s3GT1[^.�|�5���{C�`_J�!{�����E�Z�F�	��������j.��Ȃ��]���[�sc8V���ټ������������Q~��[&&�i�kOx�h(�4}��%��d3]-���X����m]���1����3�1�&bGa0�9�c��l�[���]��q޳`F%�:`��H�}�ң��j~����+ٷ�q��k��$Ox��V&v�mT��C�ގJ�r����~x�-�/TT�=ϙ��]���@��C�"@C-y�9�85���x�)�@^x�f�b��Y@��_���~�]�3�P�u	*��!��k,��y5�6>5�Y�ܯ��uc����2�ϓ�_nl�f�^Đ8#6��7�H� ������nu�r]�U6�5ա���R�&�uص�6lp 3�rb�t6�~X/L��
X�f��4�䳐܄�I��$|k!OAKu��R
�۟�Gk~m$6`纑����`�7��|'���l��Q�=@`#��u�_���W�m��PB{� ��4qQY���,��c���s?��I
!��P���w�0����8iE����0J%snv%��X�����y�H09y�A�$a�t��YZ�Y�#��xu1��E|Fy��#"���yP09��3�3T�'�y���E�2
�#���3d��Ҋ?��^K=෋�Vj�����ώ�&�F�vC%��2JW��ԑd��)8��K �jE���EFc�*���49ť�	8��Y���D��}H�K@2�-���2�J\1E����z�s�5�T9
����h/ە�>W�+���9���\���֕%���҂l�;��GF.~#�����pY�'��~���TZ�p�2U6�q/ 1P��A$��HJ�kM�V�fA҈sc�?;2�j��*����w�[���\��=d�?ѳ�O�dY��Ag�S#���X#�γ���-?��"hj�,'�ލ.�ɍo3�P��N��(&�a�R�A;F�J]6��1��H@��!����n�F���<��bh�Rd%����%����"���@{��Z\�+^:y.�i ���ݹq�_XYY�����T@!F��?�+��%G��I�Ş�H�K;,�����`��1��<���8/�z*��O�A���9��o�� ��# P�qq��Eplrw��ʍ�5)��[|x���b@-y���L���=I[�U�j!6���h��q����B����������"u�~�e�C�0�jw�Za�O��?_����a��p�x�wW_�p�g}n�v�p�&�&�=��+��~����1� ��<b6�@��<��VG0�zB�����܇2'P����q�U��+���K���w�ڣH�k8���\T�aj�Ƹ}<�m�� [+�s)�h�\^�J#���*s1ի�ݎ[c\%�( OQ�Qg z���(l�4�p�����nOP��OBA�?�[��Y��Vj���P�➋*d�&<�R��yU ��('�/�N;x1OƆ��#D��4��r�L����A�#˶Ϻ�5Qr�\��78���Cpr�a�.b0,�5%=w��/�w=v��%�CZ�q:���S�,�,vՌ��b�#�ʈ�b���Sڟ������R}e̟����=)Y�%��v�]=4��V�ǰ`/��E��6�M�,myk�M������.�(�� ��T_y[`Ex�S�C6z����9�tVv|�L[H�Vp��j����:�������@i����P�"�q���.ؔU��/*�ʁ�
	٬���������ER����G�a��20���)���<ܷ�N3�ŚV�P����ՓtS�Fc�q�T�ժ�n:�g��Z��qN>&��¼!�A�i<�O���t
��NP,բ_��G�_����d���DG��cRepF�!���f�T�m�2y��J��Q�ב��H< Z2����{~G	OR��}�r��yUuN�O��=4c�~�2���}�H%i���Ȅ<���Q��S�9f��z�5�/����E�f�]T旡l:r�H�(��Y��z���8�d�G9�D��M�k�
���%K)���	mݟG6\���r�:?hҲҒg`+��i�!!��^����Oo���!�n�
�>x��&,��c��T��9�\o�$fei��>v�j�Ϙ�����v������r���˷{{�YΥ�TFP�YU.8����N�&��A�U��8-�����m�F>����P��m�/I����-af0��¨cp�f�>�P��ד��	�/�v���9��酂�%����PA�,j&�T����;��oԒvI*��G�m*����K��k�S�M��?�:Iu�5?k T����%������
qt�r��x���W��TJ����N�@�d;00����+H�}S��)��a��3�U���U셚'�Be 9LѾ&�Q�ӌwE2�0��}��aO�@�t�h*�S��?���&��0���V8�@Ny���BBߴ�5���T5B����A��T��B.�o�0������`6�t6��P�}`8�� ;���{���(���c���,�-q^�&Z&#�Z���ؑ�mN���Pmk��#��1���ג�E�Ӕ/cf��Ar���ϳ�JEr�yU�-��͓v�`�(+`�g�t�ܮ��}�M04��"㽿ueI[jG�0��·�4���D�����*����d9�����`�1y��e�D`�,8�Eb���3C��c��v��%S����IR�o��*ġ�{�h�x�� ;~.�8����N����_0�����4�vU�꩟��4LE��E�
��%\�0@9�lH"D�~d"�wG
6��G��ٗX[q������!�]?C����]E��l���A�����BQ�%�n����/v���H����¯ITB�(�==$0z�*}��.�bG��`P8-��C'�4���}$0�H�Ɖ~tqL�/g��$/�n��	�x�7��T��M�̫�*��l�}>��vD���Zb ~�IS
\è��!��+�t��Ξv.�	�:b�3B_I��;�]�ߟ��d�LL������c3x��(�o_���)�j������?*�Z�#vo(��`1��^��a�F`�,��q��#��#���]��B���Nj~��:�K���uoD�fgaH����8��#���zk�L_8 �\;��([N�B�r����;��O ��8�h�X�L�1E����t��,������f�_�����$[,�ܵ�t��)NV�+T3��[�,;�|G@��':�rN�{c�9᪔W�?޴�-h)��}������'(K_r%�8�]�#�Q�/9!J��M��(�b�+N�\U��Y��Й?{3S]�u�K��1k �� ����ԩ�%�$�$otB}EZ.0v�� g5B���ʄ1�BMI��b��7G�ϋ�Lu���ƱV+d�7M<C���&l�t��QTʝ�Fy�[�hxsew0��v�B9�#�=�)� "I���)W�/��N�	��w�=!�f�|�jŏ8��R�L�<r��֭�4��/��E+S,_��8�߸�j���O�nze���p�`X鶗�����L���uViH�6�*�T"B*�=���i�Gc���ajѵ�^���4�*���4�/|̯'�Lqm5�~�� ޳j�����z?�~	���4Q�>����?�m�՟e6�RzV�(�@[v�d�	ĻN_0��^�2y���Ҩ���n'_�1�G���)��c�mp�
Ӵ�j��һ�b<�Z5{��\�)����h��]T� u����dvd����@�a����u�19�qC�D붵����k�H�x�&����^�it�R��&��1�-2�t5��>�Ƣ�qR<e	^i<��i1Cv^��%�Ei��eΥ��3�4؃�G�6��Tw�Ĳ3cT�$�>�_ ���ݭ&KL�ϯv>0��^튢�?Z�ɋO��9���aN�z`�����X��b��|2�;pq�aHj�������,�'�~k+Bv���B�=��4�9�n�{����R\��0��)�˾VK�=#�:���Q}R��^��=�<�v�o�i11�I2�\����(,p��_��L#��7#� t"�R�ğ��.�-�.Lx���;���Q��oҩ��<(���A�8�:���h������\���nHZ�Y�����j���.�ǨLE��(���������E��?�E!%�v�A�H��Q�*��S5��4sm�b�L�
����)|�j���� �E��bȰ��� �����J�pKk-Mܑ���r��}*$� � �9<�bp��$�<��OF�w]�UiJ����iqO������ #���JHCs��xE#����{m�.���\L?߅�ڿ�8`��/�
���%�cg�O�_�l�UsI��Ekq�2Ae��s4��-���\���Fr B�hZox�.�� en��>8���ݱ��-u23����Vq`[z��ƽ(ipT��Vo�u��:���+��j�?�1R�����Z��;�W��۔�\��˯���Z�L�+�"�k�h���o�tLYD�^�[f=�N`.T����=_�n/�%c���2-�ǯ�
�Ӕ嗭�z8��f�p�(&��߰�g��R�\�*f�:2p(�/ˋ7'p�k����!���1VR�ԟ�<�>��]���V�*�� o��Դ��wQ�\&��"l����p����[�BdK�P;h�dʘa�eH���C��d�y��/�f!E�nz�s��ȼ��_�'EI͆��{��f��sqn,ԟGXd�����(z�>|�&��*��V2-V7��E�e�)��QF�4��7m��LZSZN�&����c��#T4K� �%>6���^��\o���o1*��_:�
���2��ċ��������ߦ���S�h,Q�j�ɋ�$�&K�� 3�wU\�e��=�ԓ�R$�p�&уJ��?.8�ެ�Y;rtVw�L!ubֹl�����J bJ5cˇ� NcC<�;�U<A�v�8����;l�	��'�[�q�6`/����9(��FA�ҽ8g���9$G ����}Ƣ�+a?��L/�;z?ria�(,�㍂��敟�%[X�RŖ�ؚ1p���k�����Du��=��	�A��Ȓ۬[����ⷊ���ב�|㺵�/��52�/��]����s]T{ ��S�<m����^+U�0Y �P��@�����Zzέ�V����X>'��}�S�l.^W��$ē� .}T�]%n�	>���9��^f��u��g� E*�6�T�eHBY7���`��0�;tp3�778#
���U-�d>�gA;����S��Ք��u3$?��	2�Md=<g��a��,���\ 8R���K�{�Cuԟs���(eS8�2\`!�LH�  >Q�q�	�N�#����#�S!Hg���޹Y2�A�M��ӡ�X�l�7��A[ K�;#��`"��ņ[�ǔ�=Q�?��i@ú�Y�F6ho1��M%����-�5�wsUv���9��;Q��qa���s��Է�+���,�1*���Un	͟-�a3�e��,%�;�)�f��+��'��aG��Kn4%Ѡ���7����a���Kʹ��Ie>��e�w�ek��1s��~A̕Ġ�>��������@����6:Kt�!��Q�F�����#>b����ꩧ���������'>1�?�R(�n!ď;L���S���R�%1�Igӽ�S�R�4��܊ZM����qp	��T��4��VNu��P�1Jl��m*0>D�Lf|/�����KU�t^�p�Ac���AD�_n�~ݧ(�A+`2)�}��8����$��}'"6u����4���:8�g�&&w�E*�m�,9R�~]S"/�n1�`�#(��w��A+��>����%��c/���3�3L_;�c��V�.��7�ÂN��΀QF�>��,�C���x��7-i���e�LQn�*2�$0N#'�b��2�ͽ���Ӎ���w�E�L��ԭ|�=�7*r�@Ϛ2�D�g1O���D����[�D=������>1�3�zC7�J(/9/�%�b��'��gA],�>Z�b�;�}[PD��t������ȃ��J4�V����0r��l�����H�m��I������L1������@�O�Ӯ$�tu�u{I�!�DcEV�>�0�i�o�5i����N.5�8̡_���9%���4��z�(� !S����//��������؄\l%��x/l�bEqz�}`�6�e�!I��C����b٩ځ(7Q5V�3����#�y}�h��KzDT���Ճg3� %۱D����<r`=}4q�P[>���r��y���D�0�) ��ګȐq�ѥ\����W�uOl���Q_�W7�|�K��s���X��˞^0MQ�8)Ⱦ���p�D:\���	���H���n�#�ǹ��Ѓ�G_E�����l��Q��~vxb+=t|��f�^쾩)'Iy8�^mUt7'u�����Se^t.���U��sMb_�AR[��(ȯ��ItX�E��5.���"� ��d�R���Jsb�*��VM��]�k�"P���?��0H����3����{?�V�>u��M��~��#p�*Z�ȭ0�'�g�H�#{өQ��-��C���j�m;�|��:\A�	̝E�=���ٵ��F��4VY��\|w�*�!V�܉�3
kR��w v����n"�4Iˮ��/� ��*�hX���ڟ<����	`e�7֜�nj2������t����C�^nJ `T���p6�7��,w�?���O�?%E���{��͒56�[����C�^�������]�ߞ�W�YB�|m�������,�h�B�g�������=�R��O����?P�|��3/��0"J��S$bDS�HӼ��OX�����f;�W:C^}k%�B�'ș������)��m���i�ρ)h�����]^nf���)������kD�<�K��9�<�rI���HL~U-�5�w�(~���`�k�.�VN��ջ��|Ü�A\�8U�K���U�fC�'�ed�Y�(���9I�	�n9�l� ��݈�p��jys�M�A��Aʚ�ܻ�Wx�Nӆ�����-jĉk����/�W�nͦك���Q	��-��Յ���ap'J�Cc�&P�J���ć���e���1�$�5�X���|{�0�o��Ydw�×��-8��6��7�៖�����Ol�Df +�������/4
��"���y/���$���v�Y���:7�H^e'0j]F?�tE��1+-n��Y��:�u�[�8���! O#�G���%��{g�)�Z�݈�3�z[�D:� �*�d��V#�a���£����t�m֋��°�
�����q�ݣ��u�ʽ��hR��!��С�.��f��j=g�B(!���Q��B��k��2�Uиq�d�Oݦ���_2ʆ*�I��FL�K��Yn6�-=���F-Ǐ�#���ur�e:r�I>�h�����Q�K_��@��N�Ɇ��Jh⠸Jer��)%�$su��Ї?m"�v-1����:Ω�=��PŌB@��	�p�މ���a�a�D#$2]��,�'�Ә_hÄ�i�(��O��$�� ^!N!�%h�c<a/����R�E�n�!s���+�/�Eဇ�ћSZp������@e��
7�A.��;�Ě8M6K���h��Q7�\K�����B3O��r����0����iwɹLS6_�J1d/J_p"�^b�#���2 ���O6�w!'L�b�A���=�4�2�-� �a߷�ɂ\t�eK�qB,k`C���'�׍�ZF�Z������-�ș�#%��P��%/^=(F�I��R�T]
�/`�9"*�ѳZ	���R�z�2RDZ����Ѽ�0�a��zT~�%�𥣽Q��Q��,��D�v�I���lyob�D���P��~��b�WpY���h[��/� Q�j��E�Eݧ�ܢ&����5<)��d��Ԥ�m�4�5���%\�5�yvBJ�c�+ۊ8����X�6P4Q���4�GI�˥�N���L��q��&-��h����3Œ��P�D�U�Ny�x��p�����l<t�uڑ�O�I]��Mz�<9�(s�#tU`I������[�Ҁ���ʧ�6�B#�*�1I<����� r�y�1m��;Y����s�ۯpſӜ7��m��5�����S���l{�/&}p��	E!ܪ����X$i_�8\Cp=�/i����n��B{<�}�Ǳ��&N&#�Ջ�w{u��v���Ă���va}t��4��c�;S��]"����Zb�
&��d��p;h�T�U�$�Ԑ0S{�;�R�M�!���(JBJ-p�`,���P�`�����OJ=>a`ϳ��"�X�"܇B)	d�ģ���V�*/���u�Sͫ����TC�N�������|s1���9�.�6�b�)�k�X0ʺ����1p|S��yp�0�r��>�|�l"��Y(Ĵ�&C�Wj�B�tl̓�.����hT9�=��F�x��@�ϮNѪ�1R��+�8C��"��ɑ�`�Q-�47_dשpa����0��[Ab��Ei=�N��M<��,�I�;i�x�!3nXa�Yz���� ��,1s'���}6���� ��~[_*���'��\�R��,XKroI���i�4_��C#P�ױ_xv9c�=է��p���P���߽�ܕċ�%���ŨJ�-[�PIb���sY*�(LDEI����L!x�=۪%��v�&k>�����Jֶ�~&>ퟖ���(�����rD���Uי�����Jװa�C���+���I}�G�JR��N��)+��O�R���6�Nc�;S/�޻䥳�i�����H�~�b��N;j�zƖh��|;��ল�X�M��T�B=�s��XS�%�wG�2���T��'j�=�;}�!OWWk9Ǔg�_QsX1�>b��e(�k̆�4�Jsz���б�r5X�����h��l��i��hE0�5�� � �{X�!���A	Y"<|�d���&�z���k��H�5�yqgi�Q<�7s�е��76�����g��5�D�w�}���R�cQc��p�7qggm�s�[$�x�N���Ml��5��>=�o�U&�]F��Ia��O�F�����XX�y��ƴ���vIL'ʫq�L�p��_�=Ҙ�Gr���7Q��03LH�4@a2&5�]�ؗY+\!�a�R�8D�Fǖ	*Z�3�0���֥G�c���?C-^�ڥ�@X.z-B$�:�׉�4�Q�H-18�^@�#+M�ߖ�q"1h�\��زa]B�/���DЊ��2���o���p~̐� Y����S��������a�ה"��^�l�^���D���6���/N�w���K-.r�xB�q�[Ĩ#���z!���A�1Vz?HG7u�O��a����G�"����i�@�@�G�c�G�G����ٽ��Q�)�*����(&Ѓ�K�dzEE�ei,��#ښ7ad?���}Zr�_�J����M�`��)��3�/��N���`���c8��,i�>,a��}C�O�����=vS� �J��^rOU����rT����t�N���*Om� ���'�;b�������;_���}��_�u�(��}��f�aɼ1)��bĎ��to��B�^����.}��r��S��.���c@��Ni|�L{�}캱9�T�j1�Rsͪ�!���!����/����q��J]�D���՞.Yj�~o���pO�@�w��y.��޽ї�����$��s�}�����m�6��[�5z��*��y6=Ѫ�.��
�����×�A�Mm��8��#�S)�b[��1o�G�,J{\'#*c�hY���i�R	`q����xb��r��@/�
����ɞD��g�|ꄥ���5GU��¦���D�1FS�]�A��e�M���WH`$�0�s�禤�0��D$X�F=�c|��e���Ԧ��s��%�,a�s�,��퀑�x��dB��L��S�mu8��SKg>�H�E�3ʄ	p�>���o��iIctp�\�M^�ğQ7!S-�Yd~;�B���D�xg���4
���9a��=k�7� 7�O���$�顩4Ys����ᘂ��Ua�
:f3�/��ڤ�ut�(n/����놁)���:���zEBpw�����m<i��(��*�4�wf���<4c�����ӳ>��6��������>!����|�) �cE��k����}ƫ�U�҆y�Y�����D���!��@��ԭ��W�QZ����Ck��+:���`Gh���o���P�CBZ�^C�Q�ՔA��g-G�[]�Sq`QO��f�9=��~s�i_J&j#����"7bNFg˓�s:z�Ʀ����������~nDҬ�[Rk�,u��%�=;�?�x/3�=�Z$`6"Dask���X�Vƌw�'�޹�k�K��Nꟿ�3�6��]�O?Y)�N@��N-X��!��9�S3��+�ܱ�z�]1�>��>�b6I� ����nZ��W0�[.�����؎�s�,�Z���WV�nG#�$��p~_xHay�$����3���v�����j���@x�^��\�Q����ˡ:E@yH��h& �D�.0ja<9� }<�cZud����,�=��4����lR�@xGq�	�mH��}�l�ru�ɣQm���_��)	#b�_2 �VP���;�PS���tml����a������\iJ�1j;��_���%☝�sJ]֛����V)��թPL�%4�ችO���qN�]����y�_�%�����!s�q��k�B������6 ���HL|�鬦Ew�n�8� �i��G��)����.w���]��0j���-X|Xq��Qx���*cP��$s���� ���u�����|���[�mڴ:jS��Nʮv:���[ 
��
�H����Jڭ؞p�N]���US�5�B��c�]^��iA��CO����ʉ��ܪ-'�a۞�b�`<�C���%9]��_p��aTZwi��@�fkj��]����؏�_ ~��c��gXUy��~K�L)�t��)���ٹ&�`�&l4<�����)�^��C��_��b;�0�Ш����*c௎ή-� i�z51�g<����&~���.n�(�|��v�'�TٗU9̋�����n��5�q�c'%s�՞�;�q��˫�.�'~��C�%v-�iG ��Nw�<Ö�n��3]i���0=f���^TZ�o>%�>u*����\8��h)3_��ϱ�f��%Q�J/��ř��?r�U�^?�����yMY��ݖH:���aPt��nj��Jj\h�=�K6���ξ�Y�+��L����F
E��TfJ[�	Uv!���FJ*#
&\���&Gv(��o�������BK�,�j�Z]a{��$��}r�F�O qÏ|�q��*eudAsmuF��Q��Ӎ=�^��#���4o��鷽f�����ih�A�X�ϭ�*�����om�	�f���/�n�>	�����qO��5�bT69�B�q�9������|�	�_]z���������\���MA$��S�`g�/TҢx��c��%n�peI���� S���7��M���O#'��t��h6�Er�3L[��*2o�.  H���;��+�K<��nU�i[Y%�Y����xWN0mNiD$�Sy���
|������@3�������P�}�i��������(a���<�ڋM�iL�Zz�����"���Z��������`ո�ol��΃�D?3fC�1(KUf�	0�_+c�^ {Z='GD���Ʈ�}�>B�JOМ"�:C6%��7��.I�Ҍ��myh�jk_��L��s=e�ħ�;��u�_}�`�E!�g@<e5 �o2(���UϪ$�h�\�J:9���ҵ�����I ���(IY	j�>���xO7+�md�FP�����H`r$�m�ۏ�!T"���"�ҳ���&$�c���=����5��E��Y$X� ��'s���Fi�	�E�+�Z~m��:����ʧ9�? >-���]���i���+��AI�T-��F�M��Taob �9p�Hj�l$^��B<��x����ц�&=P�������;�dۤ�y�rq�$#_-������D�&�G�}�-���Ȁ�|f�7�ߟ����3_(���볷�i�R3��Q��s��4jV���ARu��� �f���>p��}1���6j;�-�.�ˍ0�Vl�/m��[��{d��ڛ��_%#6H�-6j���3���8�8U,#8M��^7�a����M��F	�n{g�	l;.n�!i��-�[��-FPGFa�W���t�Ώ��������y�|�Y���{Fe���_Ky��v\��B&��jQ�%���Gr���DG<�[0�AY�����I�	&�m�� |[e���Nf��s�A�=`���:��j��y��� F�@��;�X�y���������$;��Vj)7�7�<װ��6�DR�3�/[����;�ʶ�U���b�w�qI���mB��1FK��*B�i��'dQ�5�q+�a�5��G.��d���J/O���v|N�o;Յ��	�H�k l�,�u����8(!�fr+���6>���e���g����mH?V������.7� ���R��rܬEFZYN��c���}��}�c�֊�mJ��e��Fq?��2 lȂXL��xg�@�HųJ@���6��^'���j�H��A����M�TDP�4eh�f-�`�����G�0W���E���Ķ��"�<,~�viA���'��5��s�Af0p�r*:YS�&�=�`�?$�v����`
��G�e�#^q!�q�Oе�Χ{j��L�I�
���H��7g�����/��%�Őy�5�A��-�R���O���T|�0�1���3a�0��"[�\I�, tS)���3gŧ����	��
���x�n�n�MP���H�o�"���pf����~��q��|;�Z� pu��z�����_a�I�ۗu�R'�R���6<�
��?TU��m4��%"��Ө�W6q^�-�i�`>��\��;�����K����X���1�����' BR4�NhPG�e�	�x%e���=k6>KIp�p�c�M+6�݌�'�فBf
��G�9|�rV6��޿�j����Q\�p�L�\/4��w�:Iv�LF.�E?IIó�����!k��rG�����\�DJ���p��WM�j��v�H@|�\��&}	B"��f�5!6�F��-�@�v� ��y&�7	Vlх�	nV����yK���=I�{SEh{�h��8nW��b���{O<�/������e⟸��p��lɲ��d�QpԈl�TZ�S�n���J,�Q;���5[���НViSA�w��|zA؇�c�6��*E&�Ϡ��8�8HX�,Ŏ�7)Y����7�K�[	H�����6��(��P�)�u�E0z��E�y �U�eb%��i����GLp���_ƴ�B�����'�cJ���q��w�lw!��[F�+PZ�[��GŚ�j�gB�����9�L�Ҋ\$��թ=��`���l���D;�8E�gw��ܭ@4nʍ��&��T?8'az��ۢ����0�W�M܉�֑��a�T����Y��>��N�ج4�O`��$������k�0a�z���
�uh� �Fh�:�W��z{�T�ῄ�r�]k��P�YUǽ�p0����op{����B�L��7.� ��!B�sLj�����3��;'r!��L���-�N,k�3�#�o�:�F3k(0W��t0W�b:��o�:R�&�E��M`|�� ➼P��U�D�@z�j4�����5&�r!\���&r�1\��3�BW��׭����@���#����(q�FA�l�i�̌���{wA71�Y��4T��5<z>7�43��PƲ��Q�C&E[�M�NT�BJ���<��UϠqS{L�҄� �$ �'e��cb4��>��49#��d��џP�w酏Cf� H�~#��oumo),r��tY=f/�*�y`
���I��~̮��!>���>��<H�LO�������0ߘ�*yF�S��Y7�S��{
���f�+#	.<.~m�Z�r�����b�3����e0�����υ˩�u���n���8F �t8( ����� .8��M���.�AX����*ő*_�4�f^؁R>2�^*�=JL��j�sAݳ>r(SF �41�]C*+�e.^8����M���oU�#��cr�R��J�Q�e�@��_�O���B�q����Y6�;Ĕ��i9,�2�O\o@7��]T)�A��_��F�&E�'¤��߭�����`Wׂ��(�n�{tp@�Aw�O�����G���N���e_nA� s������n��!ri��1�J�0_��M�]������y23h�Ӕ�Ƞ��}��7d`�/� ��w�~�Ӧ��$�1j����}�t���Ծ��}fH;DZ��~�Y�>���Z���0Z���B���2�6�Q��y��kU;V��'-��YW��m�C���L���#6�֤|�t��'��B�Kg��X5 *�D�����G�͢��[�ʧ��c�Y�+tT��?��LD�;�s��K��i��]��.ɲ�=����"?���z����gp�n*�ѿ#1�&�eSi6 ;τ��>�{4��P���u9�`�=�ܢ���ͧ�&^y#u����_N�WO@'%B��p���F��,���I��~�쮞4fb+�ׯ)6�5��\n�5C���ʗh*$0�FQ�(�+����kT���M��,�&z�6�ء�h�;~w6���(`g��Z���.�ZX��v� I=u����qv�q�
�"~�4���4-�.�O��b>S%�ؗ蝱���*��\��R���2bb=M=�d�u
Va��f��=R_ߪz	z�	�S�ed���W��K(E^��m��c�0���i���k}K?�\���G�)x�\v�uЦ�d�������_�_��k�!�����5m+�_2���Q��-�.Aí���%�5J�����f;��d��M�&I�Gi����u��p���icZω9�c}�l�}����:ﻉ�V��:�����C���KO�9�44�wT�ʣ<�V|}]�N�k&�"*���;V�����ϖ�
:RD���b�C���L�˘[?�9*`nΏ+���4��g���u��L.�lp�d��xڏ�]�xT�:kFG��@��I~H�}��R��舙>^�KKj-i@���lP�������>6������L�
��e�2��Co��z͟DѶ�
::�ZQ&���Ă?��T_5S�����^$*8Qf�� ONu��O)Dw+"�