��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7]�s��^T��N݃a�O�BL�z�᫛�䣄^oK(r��*��'��!N�I�f�M^.i��Z� ��g��G��>zQ��G�n&��� P��z�� ��Q�/���}��nЂ�;'oM��^7<vx�V�A$�U����<vR[p����$����%7���ϝ���4L �Vb�	�l���#8���
k���*]���
���C<ď��\�zm�e���o��b�kdAK���n�\���ɷѯDF�ĳ�U�Ũy�VM�Bi�:� 9e���B���G�>�%���(j�e
a�|,�۽�����a:��{J��l�������z�t�&�q�p�	��$v]�m#|�j�=�b�ç��W�����|Zc�,5�C��@�}	|N��
\�f�!4?��~2E����G[���*o&�m3�7.��S%�VƼc���ʝ�a9��%u��J#�n�a�/n�2u���Zsǣ(�ba=��u�Uy���b(��{b�.,�X]�9�=�G��c�M6	7��+����7T@T���Wc^;/��А��v�q�V�e����5��*2��nn$~�41J V� g�K`]��	���o��4�I8#m���R9<d6�_oGj2��9e�(�mN�ĉ\��?��E&�_
��[��9t�%����?y:�Y��z� "
� m�7�R�pQ��*�j�[;M>�
<�'c^��#h��8�x��>�F(�[ZݱtE�^�
��VA�^4����k�;c�Ɔ���,�.Z��Z�61L1�C���O:0����<sUI/�'tI6���L���I������i�K�������3]D�58 8�*��V���ͭ�,�wm
�����wK�5_U�<fb�Պ�t�� xg��`��U���|b�\*��H`�+�Mk���{����۱�v�;5�|� ��fd�YQ3�.]ǫ�?þ���eW0�������VkϷS Q�b��d.t�d����,��E��O�wϒ��ח&isT����m���+�}В�M^�����u�6ٚ��nm*3̋��$KMy+b|�9�o��\<A�%�Q���!+��ÈO��9��86��&8���l5J�%i���#&�&�h=~V��w�q�[.^�?A�l�,��c�@��lQ��QC�g'C5W�v,����\T�É��{S����_� ΅�.�� ]|?p[�d%���?|�|�8Jp��3�)�;٘�yj�w��M�E}j��ɦ�@}��~�FQ��{C�Hf���Ɠ|쌀G�f.����)��	����σ$ђ�=蝑g��@j��+5�/��j	>��E���K�'wQ�ʴ 0^N�o�Hq�S��D�|9�*����������Eun�m�3�|?H�ȫ.J2��%���	��(N��L��w޽���X#��!��c���{:�ƚt\�M���@<�#ux(��6&��s�C�1q����n�ˍ[V*aH�>���0���[�LqV�h�(MM Do�TF���y�0f ���+��
�b��X��mZ�'}Z�8��(�C�ߙ��Ϯ��V�߆��O�(,�&0)3��������ꑢv{�,U�Ikm}��ַ��ck��+ӆ@��p��icY�cPP��oF�,����R{�8�L��¨Y�SO�j�%�p�o�i��~�����%�%([��<nB:z]�g�;ǌ�ԉ���n�j{�UU\��>D3y"B��Z�z�����B�5�ut!(m��<q�j��NIf'Ms��0��u��Y5�֍F�ub��L8=��M��;���� +?���Gb���¼���`t!�ijlOf]���{ژ�U�����a�-;,�>��:�ܹK���;���J�n�d(��9���ĈA���3p�����D��S!t����/���ۜeq�� [�arj�Ĕ�����>-1�j��j�W�Ӑ���B���g���j&��/���O����қ	�SR��{����|z��M��?��c�B'
g0�"�IJO��P��V��L�-�S���~L��cٖ�3�F�^��34��x�Q��|��ր�ʯM��&o�N���B'gt�faќ��>��l�;���!�Mv�U�:���'���	(4�	�{�j�]��)̐��A�8)��*�̖u��&J����%K����l�ekG��s�r�B��9`�>��ޞ�{�%�d9���+m�H��C���l�C'�,��]���M����t���:�,�ʕZ#g�6�<65'ݾ-/�=K3eVw 6�1:?�#�́�vh
�́w8	��ϱ6�c
څM�g�F3c��D�f�d���]��iv�S�$��{������+��! ���	������pHD�U�Tܿú%�$�L�! ���џc�f�Ҧsfz��mؗ�fB�HE���
�}��2a���Kl��/�>q� ���e��SN���`=��`d��j1�*(X���\�A�p!�L#D?�'�(<�N%����P}��1�&1�SR�/��.������� �K�v�&�
M��w����Cb5m���9�2z�8�,.z�O��v01���0��>c�>�Oc��ױ,��E���	ĝ�f1 kϰ���y�����{@����gj��ǅ�̍��;�����Q��L0��3k�����g�)c�m��U���4RD������{��IǐNg�pc�b1���e��,�,���{K���%z�P7!�ngd�ԵH���n����Ɂ"=r��Q�$�V�b'�F��� )fĵТ�C�Y�Z�ؙ�p��b7��Qbb/>�����Z$
L��M�r8��79?�A�&��ȅj�A$�l�_�8�7S/�T��E��$��f{�z��p�`������_)�:��@e�HSH�@��	�q�����4h���@0������raa]. ��h�\��?wU`v-����d����=rx�C��u4ni��#��H��r��c}�@S��iet)�X6���W�.��ǽ����[�i{�%���i-(Q������V��?� ΰZLy�A�ă���q�Y[i��J"���h�Y�wh���_J!�2�al�*�D���t�ze}b Q��Q
�����,1��~�tC�$��J��d���h��V�D2]n�p��b�����G>����I7��"�'lwKk4+�Ox~&���M���(6�IS|�m4���V���T��prwH^9�������W2��vǿ��2��Ece0�bs4�|ݜ�H�/�7�!��m܃���0�<w��>����og��;�:�/�~`�0��H{�T���!l��[ ��匂�����kj�yESy�nw�b���{��%�V��2\f�b��tf�ͨt)�Md��5�ȝo�U�]UZ0����L��‸?u*9���V���[�g�w�J�SJ��ϸ�vSy�Rc�����ļ}�/W;������8-�a��)�/�h�=�}䤄���,>��؍��=Y�\�O|q1��H��d�"i�j��Ԍ�@��jh���n� ��7�W����^���bxiyx�>�y��Ä��3��~�d���Nz��>��j��˂�ݵ�@x�Kl�U`ݜ�m��Ƶ{Z�E���'��������RN�M���
��x%/X��!CFg%$j*	�-GK��$�O0[�[Є�̷~���n��gq���%�?����O��:�/)ɤ���!;(,e}��;�0�k$�C��|�,�~آ�h���\ +!\���|��K��"��t��J�ѣ�(��M]y�.�V��{%M�Օ���$k4�̾��2�i><���gE׏���Ǥ� 9��X� �s����y���E���1�H�ֲܵHF�k�<R�j�+�Ns�B��߫���w	����k;$,<p>�����G.0�W4v~����B�9~i#�ߺ��tWf�a���������gg�����I��6���K �am�y�٪3��
o�����H[�)(������U5��K���Z�E��cy�m�f��m����a�خs�X���7~+�֜E��n�ߔ��������d�5�7!�b�c�np��
��w)�1��������0AR��z7�V�BU�<V$;��A�!,]|�_.�<0��M�ep���76�H�W�ƭC�F�����̨`&;Hq3�O[�U��G�8��
Q�#��N�|�ä
r^���&~0ߔH^6
\G�@`t])�VEpF�/� ����t�S�N�"Pz�v�t�k��-)�'v�8�W���� ����=��Z<� ������+�[lL F����~�:�Lؙvb8�vƻp�4m��Y��3
��-��\�nA���n辅�j�bɎ�^��F�U���ׄZ���Q��#�1��ӭN��y�v��N����'͑�칷�O�G�;��z�)yu�b{��`[G�:9�+.��%�h�{�#�+�����.�v��d�Q/�.J�+�uc��o%� '�V�.����ǖV�,���t���Áu�9L����H�H-Q�� g�Sٚ�,�>}Nդ�8�8�M5�Iu��� ��9�L���p[�EX�#�=�'( ��T��pCM!���|P_YE�Y���e��	*�ͭ�J~��
��ͦ_EC�B	�4����������0�����%L� �Hy�������f��R���8�q��"��#v��B9�NyzHL��>AD���987���Nj�jnY��Tυ��:�1�,�c){-E��Z27n�s����BO�ɔ�Ta$!)�n3"4�|R�.m%������/��"�/T���� �����Y�#5ZAh	4��Ṱ�҅���Ld�*{wG`�ka;�4��ow;�1`���&���&bޭ��%lG�k�e�X�����>v��#fZ�L�Q�ޤ��[��Q�@�� }2�8ƹ{�N�cA�H��K{8���b?��El^�*��񅓎�,�+ ��%��?6]s �e�%�