��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^�.GJ��-��?f�b��(��ҥ��Y�����!���نϊp��=׈�kS(�?D� Y�S���#��f�����V8?�_���Mg�\��gѵ����s=�B_M�E�B%z1�����U����\�����ZI^C'���d�_ ��-[b�DU�Vյ��*�0��/�^�]ݚ�Z���r �Ї-�l�h� n��ࣁLR�5���e��G\"�JZ�z�!���0�.f ^w ϴ� I�L�J�ȷP>���ө�,5�%%�bK���>�͇_|'xƈ�&8�.�7�ԯ[����!�X��fŷsIE�~O�l�d�O!*�W,��H�����;}"���9��k�CD`Y���r|��# 媑6�x��31�_y����ъMd����<y �߱o��)a˘Q7���{;L��:�:�6�w�K<�&W�u��wK�M���b�[���h��������HC�δ�;ի'�(�����Ӥ�@��$ �V]z	u���#���ځ��2G�#�B	�}x��G��߳~��Yi�y+�����(r��ꕛߥOy?���B���W�uuB�d@�Z�ܩv��x= �ap��X��(O�vNleJӣZy�D�o��/�?t ��0��犢�?�T�*0��Z��}N�YE�1`>�	r�D*�>���NqxVJd� S�3459��]n��H�Dﻅ"��7w�a�t^|�p�v�5U->���^� �}�c��@T2��)6V豓�"S����Uf9�g�$j��j����{?��S�X_�H�_\��ݞ�D��.V�H��BF©�;)B�6ƨ��J��� [�uK�0�=��D�v!����S��Nn'
j�z �x9������#�1Wl�v�ScѦ�$���+殗�#�l�#2� c������h�D�2��ݦ���)��؉T�E��:�X��LO�l�OǞ����j��~Ƈ�LD���2�H�"龺Y�����!.7�hU����j̺�������IE���qx�;J��w�V&�����\�Iҥ�2��\z�<w?�\\	DD=L��j{m�φ�J�s�ު�c8{�w�e�!�obu<v���`�Eʏ��Ju�����-˹�l��¯���Soe1�O���L\�T�Bgzk4���C�K�t��"��m݌-S��2�Z{��.F5T���u� ׹J�02�:�,�S|uUD(���`26�N�PF����?'x�-��!��/��Y�s�<ZV6+����}����g����J ñSkm���g�owa`f]RC���=u��I<�۲g[���Q��E��!��C-8�|�r��Zo�!��@�g��'s�t��ŵ�.̩���d�7�B�;�8�r;���cl~�q�b9`������m{�[�U���OMU@�V��׈���aJ�4�����I��O�����_�q�Y ����V������E]AܒZ�p[	���M~�[�-�q	�@r�	6O��{ɧW�Gp/�Q��[%�)��	̚J���a?^�?G�>��vW T���m�󾇉�5$�)�K,�٪�N�|�le��c��D��ܰx���撄ʤ�E�O�V㬈��z�ˏE��k�����ҟ�_<1+ٳ���ت�4����1�˗o���a�Ą�	�Y�&==�2]P6��
��@���V>���P2q"�y�@W|�J�V+�h$/��
�=}$��3���bݸ·������F���U��o[�L�X�7�i<f+�h!􂓡��J�#��VB�(a���'���f+�z��᭼{k�t}^�-v<&:jc��`��/ݩ�j�i^�r�]	��a��w�igKSG"�B��jj�(nB��y�*�}��+��
�IGe|n�����)���-
��,Q���oaP�U��6�!]nс��P.��H���J	�N����C�׏��O��1����̶"L���S�L �`�v� g���c�[-�� R��s���a:���3���"5�lp���|��v���`X���8ѭ�x��*w{�<��^8*�R˧ޡ�C�&bU��>�d��U��s�h���e6�7qI���C������dX�BD���V/��)5��K���J�i���AO��e(�0�g�Z)�e~�j"9�N$���K��
��w�,O����a�i{mjo3�p3�T_�U�?���D���A`�F�v��S}��
D��H�c��&3Ts�M�����b5�V �0���E��|�I'��8ǹ_�&�_���������gO	�x�t��>���8s�������繡�D��ST�m+'�kw�]KmM��a�i��RTƇ��J���o���R)崃��x��R�C����-K���[�U:�bRE`7�� <rA�J"�峅ʒ�S'��@���S��F���o���y�I9��e>6��	�0�}q�0S�B��fLx��=S�юt$y^�%��gX"8�i|X�����{�Η�j����W֩�G`�;���p�L�l&�@��2��~G�l0�l��8&R\e��qj��M�|�,��@��eˏ<@��6h$=L*���;H��̨�0�z�[ر'��C��2�K�Ȑ�jq��Z�E�����Œx,}Ӫ�����A`]l�7�Iz���c45��[e�=�9Y��񹮞��::ޠ-�$�Ӑ<a�J�=�ә4q�t_��
���"IxW���U��NB��,�R�AtO����kq��ŭ�@��5k碌>S#�}36)�L�,�K1����;R�$U�M� tʟ�Z�aڤUΔ����k���Jk��k�3�2\��e�-�����S��rop���eDk��#>�����y�Y��\���tܗ��^D�+�Lџ6P�B0�:b���܁[XQ
*/S��J�xIL���k�wy�%��������HUfp���<B�S�����JOe-��	�Cd�E;��0U:�6�<�ğ^PndvQ��{(�'ٟ��H�_w������w��W��U�9x��qw_���W:>�T��澕y\_.~k���V�3b�Э��ǻE5,4�xEB.>'U>��Q6X{B�՜��Ky�7[&܊����A�� ��҇�c�����@o#���t��睰��uV1VX`LVy�d��`uǃ;�u��5�s"Z�}a{���,U�� K�?��g���$�H��dg\���28b��U;�pL�/�ӰX�V�8�pzAߘ�{wl������3A8�}�u�Ծp�"��$�'��<�o����	����9C�$[�����F�◶d�����kI�WkjGj��X[T`�B,*Vb�����a@Ӯ4�ǭ��v�wxT�iMe��#8�_߃�ob�5l=���h�/���)��c0�h�U��(<��}s&�JL�
(��ʟ�͜���G{e�6��Rcui�r��έv����V�AՊ?������� ���
����瑸حߐ��I���d���<S��`*-I���ݢ
Fu��bn���n�-Vw����NY�V�Y�й�i�QN���2Br_qPD9gIR���~$���S�� �C�M����J�O�K~5g>�ܙ:�j�ޅ���酧�7D�!���0~Z��uG�*x�s�,�����I8�b�śWu�j[,���Pd;����B���~x��٭�5r�%��7sh��J��$�"U�Amy�2�������Tϵo[���5�魫c��64�#�y�[¥��c0d�9������eӇH퐵�dK����&����PX�ޣS��}�T_|�81��54sw�^������a�M�&�����~����H�%RK���qs^�SS�>�I�j��ͼ�D֞!evv�7��p��є�w/m�E�᳈��_��q�}4/GL#7Z��DQ�Ƈ&��]'��=2�S��3�h�3F�v�j��cBY@��աe��P�lA$�@Q+f��	�2ֽ`:���jy�UP��q-HL�o��|
��7�3f����aY���;��0�Qb6ۊ�6CyS����w���B�Y��J��QٿT���7��Vi�Qۢ�-o�G���*�� t�WU:��7-���kYmC>�#�KͪcL$�K�\Q�E$v+�D��-��T�mO��a+0����%��ˬT�y���*2�U~�'U��[�!E��5�:�� �>�[�#͹z������^��Wk�w��J�j`%c�1l���B���Y~���ߺ��>Ae�%L<BQz�5��^�sת�&���+�Q���h]�3�!J�OK4!h|�
'# �9�~��c���3���+�ؔ���Է}�M���*:\A�[�8�7��D��П�
 脎��݈��m�d`�DX�J�"�ڄ�*1�Z����.f{˜� �
�a���Y�`#�ŉe���S��=�kؼ.;p`O��÷�(�����a{3�城���t�p<�*m�ʖ��ȯ��L�P��V�x��a�����3�G��!-
B���6�pA�Le�?:�\�L�2�܊�����1�i�����HOE�k��0�mm��MBߟvu�)�ds��ɩZ�ynŊ�2��J�+C}P�j1��T#��CE~�J�$�:%b��-�i�=����̸j�k>��!���O���3g��?p��_iq�5�u+��O�v�Xw��g� �L,'~���^\��M��;�*N��3S��+�Pa�2��AZa^��D%1�I'��Wxp�U�_��\(�qak��W�捕m���=�j�K�ٽ�G8ƃ�k���-��Pb�Ze�q���Ǜ��]�8��[��t�����e�-#"p;��NDx
�����p[*�d�3�]*]﵎�
y� �^���b��r��G�kHz����7/f�G�_�Q�n+�J�tK"��f�ȷ��8�G��x�T�fŁg����">�m�j����^]G�J2h�5ٓ��Uo���K�YR�b�Ē�h�1<�W��'	�%?d%~��4=)J�z�H��i�d��%L�jQ�>��%�.w/���pI�wObkYc�@�t��0s��-<����?[=�n��x���8��kU� �$�V����e"�M��F\Gq_q�T���w�:k�׾np�(nQ�^z�X��
IN��8N���:xk	���WW���0�2��=c���@����ß4r�s�z��Egnׅ4
 �@Ѹm�����4� �rC��e��@F$��M�'8�8�2)�40�}��b�M��/P�v��KU+�!T��00PȌ��k�B��a��5HC�-�/�z~7��Ou�|���f��1+�� (��x Q�9�����I�Z�8pM��?>�<�9Dl��z�o���~���z�W�џ2�H-'>�j[��� ���#��z�5M�O3���[�y/)��N��<vJ֚n�]�a��rW.#���I,���3^e�#Q����� !^z&����1�*m��v�r�[ep�Տ	J�G��Žw,t�z�]������DT��ܖC13r{躹#&#ol�V��޼���q�RB�׫sߦ���mEo��y]�cs�`-�e�J��SK�[��)t<�+Y����z�Y{DT�6�r�ɗ2�F3ql��b������e�_�D9���7�x����ŭ��8��A��4��cG���C�/F@#^��E#ԓ`�����R�����K0�������ma�w+Y��+�8y]�a0�)���9�BCwt�j��-�����jU~ݭ�Y�� ;�n�вgXU���뗀�yLP���P��Uj�5!.[�F�=������98���R�����΄����"8�֚-Μ���鍊'�����KV!���ٴ��cC<���\�(ԙ��ze��?\�|���eC���;��#$����o�E��׋�����P��/WrڅX(�aۡ��.�zn6	i�����,L�A����������46��"S`0?�QIԾ ��5;ֳFm�B㜫�u�����Nl ��G���4	:N�>���5�O���8�\\�~�w���k\�PM�s�N�<���|^��I¸�W���?F������_���G2+5�s�ݗ���Wz>�ApLiv!�S+�f����{���ο�!� -@����v@��7eT�]oT��7�j$j�L(�#(d�����:s�D^Q���<	+i�bI���礊��&*�/����7	/���/aLG���[]�<���@5Ѭf�&�R�2O%ڦ_1�n����)FS�⾨Z�$N�Z�ٺ�&�_r˫����o9�L?�«����~q��	5f

T�`R���ǝ��{�$���t'�{��y]~H����=��Ї�G�t������K$d���*Y�yK���0�߶P�u�k(b��)I���T�j-�Ѻl����s���1�(q����yyc,�8���V�\���D �o�7��dM��2�I���<:�ZF�}4s��7�� D$wp	��J�/�1�b�Y�3,N�W��m��92�d�l:Y�3/׿�B������z�r�X��ݻU�L���F�j�|�5����	����8?��H��;�%�*�#}�7|�u��g�P��2\�A~9BP^��|Er�Ϝ�\c|� ����uG�J?�!�<l��2*O5�q�ZQ[�`C&�%�G��9�(��O�_�"��e:.v�S����qbY����BSbk؂�CR Y�E&,wC�%��>�H`�܁�GMԎ�&��3��f]�Y�ko����2�.49���p�#�:���7���1�R��ʳ ��wt���6^Y���\��<�����"�3����Q;B�%�c�C)�P���h>f+*~�4r���{+�yJ����!i�ޣ{���eBWj�:/Շ���I�i����4|[x�}�dg{�;��k���w�N|�Tj�X(�)#