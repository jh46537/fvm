��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]ǂ��O��˰�	JL	B i��M����@���>��y��ƈ��	@'����N��U�z0�dw��`�I���臏p蒎K����>�+L�����Џs���a� �qķ���q��۹����
�2+���d�}D��dMP1՜�+M�Sc�����ɡ���7���,{��k;����u��UU�[�uvO`!��M��B��e��<�,�Pz��v�[1�*�7�0��-�G����_��2����N&f��]�z�l���v��	f�e9������Ժv6~��n1�D&װҦ�����2'�*{����C`�0_b��WL��u�lŵ���I'�g����߱}�k�2����\[>a%�)_Լ��(�bd��.�m|����1d���2�]���0j4�M�YTY���ߥ:�j�ر[��w`��k��`e��"�^��4�3�|-)\ߑ�Rao��