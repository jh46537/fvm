��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(|����	t!&�
��7u�"�@�G�!�>��q����7>����d�E�vs8�Z��3�!�i|��L�����0��	#���4�0dY;i���������a �c����G�h�
�s~���J;��`Jʨjжzfŏ� �ې-"jPb����x+T�W��ZE8����'P��ܕ�IE.v:NA��5�!��
]��횠Λ
,�7���8i��sD�> *N�bTq�tp23l\g���4+�&�17�ᇳ�6�^}��35��$w<yZ���)3������^���){��d�m�Abd3#����-���1�h��u���åB���9��%�oOb3t�u9/����}��eG�Q�v���&�E��Ѡcn�x���9�7�RĜƄ.a��j��c�Ý]&;�H5$��.�ۤ��v�Y�o��t���I�e�1�q�qf���T�f�	s.�Ve��*�v9�l�Q�$�~��'���`�����S����%��k���11S��W�9����~犷�������NZU=FY0IBh�L�"P�O	o�S��E��o�kd�-�\����)1�,H%U��vU��g�PK���21�q��M�(4�1�	���	��Eo4�gK"]wS�]N���"��̜�{)/^�^�oO�1&*������X�n9܇�� 1�}+�0뎓�-.̚ca����pz˪ITAfA2�ҁ���EP��v��I9nQL휩ihbJ���&�M��!���*�_���Cg*�>.�:�9��һ>�!��O�6+�aU�.��~�<	�$�:�l�bh\o⢈��)!�	i1�% �Ɖn�814p�w���,��	��6QP�sR�rV��;͌�.O�S�|6�4o@6B�N��(D�﯌7��̲a������QOe*�᪹n>F2�q��ͧW�\�֟�#�L�T�KVv�.���1�U�1Gy�'o7z����I�Ƹ�����y/�0�� ��?"xiVP�TW̾C9�)\��/8�߮)����IĊ@�J�wwwYDg&
�m��K���̻,�5�p��2ڪl�gh�3 n��_�w��כF\5�TI��g���`�=ʀ�9�N���)��1;H�,/
)�H>o�=x�Q6��Ag��`֚غ�A�|)�}ه�Q
%ܜ�)�n�j�MjT�Ι�/�DW&�\�ʌ}փ�A7pW��f���T0*����Y�Ʃ�1��t:�n���L��@����˞!L��6 �xF9�A�hM�>L��2�.a��)Hڈ'�#��\���S��6�y��f��@C�39� :������Z$�g4��-�|��q0!����M���-��U�8-����N1Ҵ�I�gX�$�2���㛀�U�C���"��#N%q��K<���yӽ� ���k�d���4��tw����Z�,����&�I�M� #r��� u�.�Dì�_�2�w6:qҤ���<\}�'��#"O�9b2��|o��֐<���%�R�aj��A���}[u}�uҞ���`��Z9���%jjA�B��Am��e�n_|���$,�0,0�Y6X`���,j)ו�C�(<Lc����"b]��v(��B�]-�X/��g���]]Qp���
�΋)�R+NQ��x��6��[D^#�+id�6p6G6�*�ˑ�ABy)֫Ae�-��ˋ�;�d��|߃2Sq�J��ތ��P۶[����ގ��별�� �@����V5u�2�gm�/χ΂`oݽ�:5=����m'�{�|cF��m�=��.J�[0��f�Tv�Qd/�ց��+�xh�Ro��OY�疖��I����=��� \(����s�����O�����-��f�'i�.��z [��Z���;�⣄�=�����5��Ɔ�/!����bZ?��m�'F��Y���wڂ'b!7f�����n~d���<��^Bۦ*S���5�	Po��[��X6��Y1���J5M����q��`�x_Є�B_J@{���Ș%=ٲ/�~�h:Tc��9L�Ɏ�F��m��f̡ZB�<�*ԡOR���E��	�u�����Ǣj��x���[���Z�ɦ2|�d�Ut���H�2G��lĝǙ�[Ī�G9ܯ@h��S0�2O��>��z��D�>f�"6���$�������r��%��# �Lz�~�i=�n7�kβ�I�Sp]!���y�n�x=�+C����G�h���-�:pOł���/�x�S���([��ӛ�i��d��\_�9�`Y���=��t����_"[�)zB��E����D�9j������-�q�0��x/Ί�;�ѪbPm�hL�?����&��gaOy\���W��͗ԗL�Q.^ϡ���I�h�E8�ӄS'�����/�(�\G0͚��{[�<l+7]��r5=�8J�U���Ü����de&R��/7ly�-��8U)>� ��]uTf�^��n7�'�by$�d�k��S���/�u���R)��l��Ԅ̊A�}|��4c���:���ʮ�6��1� �������8������/��AYq���}��N���&�3Y�[����3�V���XZ��'�.�2��Ǝ�~���y�@�"2�r�D�\Eę#�0�p�k
`�>��yC��,�����#�{A@�}S��p;]��vuMỸ�9���T��ШP�%��`L?\�lA����o�����ܹ�����t���J�m�,���{�i�r��+}�����8F�� N��V��Wz�����=�m�:l��9Q�%� Dn�M��_���|�9L�%}���z�d.����,����p�5�����Տ(Ŝ��t�I=��#�L�OȷTĹsFz�g�f�Y���VQi�\��@8 ��"2|RBy�#;�j�G� ��N~�3�io�No�!|"� �����i��H��P��p:� 
��ՠ~c����K<P|�M9���4,���&�U�z�9 !d���3⧹��Z��x���@�L�_4�U[�5�Rݑ���#+���T��)T�������g)��>ī����b^{�c�m+�����&M<gm����U :�?��)��aV2�ołJ>nC��5k�I��/�v��<��}=$
w���S���:����,E��������8�)���o�:%������?�p����J�z�Q�W��1a���+�;�y��9N������	'�3W
v�oSG�����ar�w|��]i�f�����{5��:qpi��Qv�l*|
��*7��7u�Y�>T��ӿ��Y#�RV���t�Z���G�I��h���Sr�hֱ��85�IQ��P_���=挍�v5�q9����fHW��q��n-�C[I�Wb���)�_�O��
��C��"b��W�|��]�/,������:,��"LF��`~�{u�w�g�ک�(�o�;i��@�����C�~�&�bV��;^ ��ّ�h�ƿ�+��#���>@�:#���b�ɜɁ�U��q	�џTK�7�)iW,@W��z�O�e����"Q��$_�A�3ǘy�=�|��=���œg3���BX�_5�U���{�8sq�]��ͨz��yX���B�ڙ�P� *^�_��s�k{Vj�)t�������"^m�`p�/A%_��q��ӰZ�,�Q�`���ܻ��|�}vz9�=E�����=�\Uŝ�Ҳ�����[q`�o�����>�}���ӛ����A�:�Lkn<��|�x�j�_ub�.^�~ݴ*��X~�)3k���cR��3���DM�t�6i���w�5��~��3��)M�Ɉ�z���Zy����+��E�E�`X�w/jYi�����;ƥR`�ݼÂ9�Q�|K`HL��8��?������|eߗ�Ψ�yx���>��J_��w=��I���.j��@Yyj�ί#�'2@�c@�km*6f��wӰ'�r��ߧ�IchL�a`�� ��`ۇs�
#P����m����|,I7�<G�x�U3B��nyn�8;����@5��v�����E	#c�mz�����y[A�����FD�z��p�������V����~��A���{W:"PY�O�L~d��g���H]ќ�AzXm�F��+�c9�������6��ڜ��y��D�t� ������[�x���)XNA)��(�L���8��"��,�`P�-ő��s|���hM)8~�ș^ޓ��.���3�?�3ɖm4� ��vM�\�x\����t�?��nC>1�	jr|,���S?Ba�f��D��z�w�~M�_|(�;X��n��>Y��l/���e�CǙ8�tf����{�g�����a�����
#'[�tg��F���
J���
�~*�~[`2�b?��
L~c�O��0j�{�4�iju��>�����:lo�f����v�dd3�q<B��k1*ʽS����.
8^D�M:S=*#}�>Wx"_���u���7ܺV�i�T���L��u�}(wT�OmV�)��}�%D�^–�I�-��
�¸�����vH7"-F��p�[�93o���l ����却��ZzL�����.f����� E�N<�
��<��׼Efʀb�e�Cmv[~��}��������d��t ��
-D�"�����&��hḼ*g}޷~4��w!�D�F��L�nm�bmT9=�0�}�g����	�qAg��SqD)	�[%�%�ֱ���l:�]�}\��D�\ il�-���K#���{�F�2-ʰ�Ĕx���o��5;����)����	3֑X�O!NU�x�~W�#{