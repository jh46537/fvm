��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���q��՛������@�oa�R��Iz1A�#`�ԀP��Iqh�3��F�`�ҥ����c�
K4#����ge��T5��G�z�4��R��\3jU�;Ѫ.Xq��d���D��nmac��V�ܕ�;�)=�(?0�י+�k�襮=�%�YO������鏷w��>�s]��6�t�u�;]��4���!����q��
1�xF!b������.����\�2�X���`���~���4�k2Y�a�w�7=�E�u��#��_f�g�:�S|.�� �֞/^���J���,\*��p�#�0k�|
]c(��7��ȩ�'�Q�	�kR-`~���Zk8�$'��x��A1����Ko�� _'-l_���\��
+*�q�k�����V�LZ\?rŮ5�xwpP�V�22m��w�j�{!��;�Fs����]U�ӂt0���Έ'1�j��	8m���}��%!9���X?O|�GKހbL?ҵ�S���Z{���Z�6
��N��6���]��w�5���$7̙�����B���Ho�ɩ����.G��gX~��y���RnWN���'q����G'V���Bu?�Cr�ݏ\�r�Z�;]4�@���D���輀{s�`0�λ�m��$�(�E���u�O��'D\���sl��Td����h&~��|�l����C�M�',�}ÿ4f��H��i�����$؍�<`���=�3�L�P��&\: ��v3�VJ�E�C]�$����vQ#�6��~���D
��=K
|��"�$��T�^gǊ;���{��$�JW����Z�>�Q�a?���5팷LP����V6Q�?&8!�r	72H2��\�fPc�2%� ã���[�ԏDS{r�`p��rf�JV�q��'�OZ7�;���WI��8�+R�[TrH(-��&mL���L��2��?��f{Hrň�E�mC}B��=�S�k�����mk�ۚ:�y���\s�=T:�(�4LY���=s�O��a�� ���Za��˒7jҼ�
d����ILt*}�_+/��/�nR�\��d�T�2�F���8����vzQ,n��2�o3V�������k��L̵6j�}���6����G��#=��~K�l�ax����F%NR����J�w��=��"�y��b��`�0��!�p񶹵8;���/L��C+>l�n;�B�'V���9c���7��pT�~7��X�.(�֨nU�A��"��1+�jv�k1R���q�D��:���V����Ghmz�噵�T`%�K�S�w����+KI���'��+�yj�ȿ����.B�0GS.��J�t��S�>Ls��G�9c�� P�j�Y��(*#91=ΡFi+8o>AhN3;���:;3.+�[�pz�T�f,1�cL3;,��LMHىUs�%z�~~�V�i�p�"�	F@I�c����f��Շ���Ph#JɕR� ?!��M���״�A_�8z����PsE�O��׎n��[	���8Smȗ&�S"|73#���Py
Ow���|�RU9e�c���G���q���E�*\�~��ڛ�!\��������W:�z��A�:SlL���b&��i�#��~�BT�%ω0q��K��Rq7�IL�Y�~RV5�KWO���sk~{4%��Lg9�W�j�m���R/9�u�������mO:)�̾��u�V�X�P	91˅�x����4��'�����;� ��:V�Y#���\4��f'!_�$�@���y�
��z��'�`YUbn��:���q"�*��v[_��y��59����_�F��w#�ҽ�g�>�i{g�A~��x���y��ZT��30"��Ag�3T��g��Cʍ�<V�n}�@MD�����Yd1�2rBeՔ�r���{���Ό?�cV���sxV��K�~���?���M�>
��9�`LCUD�%�s1���4}�	6:�i�hZB��&��O�1�az���v���@�f	u@ �*�6WR!�no�͒�[���)�$Z4��+�q�AM?��x��de����}⧼
�RDًY�GG@���5$� ��w�%@e�,���> �iݰ�(E�s��s�;S�bΫ�x��UU���i�4L�����.@�.�6�]�,������(L:Dnߓ��QP���ْ���F�%��Ld>[b9�� 0��b�b@����8S%4�>��H=�&^kWD�Z^�����	g�e��F,��|RRg#��Γ���(*0~��ȮV���^=!gv��<8�$qZ�ʭ��P,qC�E0Ԯ��b��B8�'|ސ7�˿2�����/��`�T��<�~�q���BA_#*:���
��'�����rc�p�TR�is�2�[X���n���=��ʟP��~���D������Uӱ~3�-�}�6N5ciA*Ϛ΢�:�rv��8�OUJ�2�3��uNs�`|1��*c��c�������VaK��"�rw����o����H�����SQ�muO	M�ڣE�t���ӱ�-#��k���0o�^!4T-����!痫��~�_����w�-�	��7FЙ
�P��<����}|�E%u�\�&
�5���)��:�
^�q�@��O��=C	��W�M�az!׷k���G@���Q~��A1ݘ:��Z����V�W�W7 K5E{2~�`e.UyS]d�'a|¦�Q�.�筆"��
�e��F������_�Rh4�*�Zڲ=�('�ߩ����r@�k�ؤ����x�:ا���@��n��=�'EW�X��(�$_`J���c�of�R��?��!3V�RfT:�V�������t��ܢ�4���AxW,I19�v��#���k.�
S�抋h �F�x����4�\���0^��w�����K%��f�
�������j�=w�P��b�n����KɄ��hպ�w��H#H��c��%��N��Nr+�忱�
�p.���4��`�=�H�>}F&[�[�r�{�h�~��E67������z��V�5��L6WG����n@_��"!�Rj�I�����:b�
W��n�^iq���d��rMBV>�R/�1T�����/?��\�v�+f��8,��#�zs�̳�[n	ͭ��Z�_� ͂-��S��f�*�4�{�8�^�w���~�������i��I�:���Y^��5W$�J�"���)4D�A���-B�A�|��r"̅aI�5��{P�1�"�s_<�I�J|�G���+y�O�,>Y`����$�)�M��*����S��l��n��~}�i�z���6d$���o_�~V��y�(Kp]͋}��K�����_FT����3Õ��]��Ёi$W/W;�&������N��Vx�|����v�=�65a���[bz"�dEap��~�Պ��_���1��H{������#5���r�x�0W�F��O7��	Xw=�o��4�g�e�[t�d�H�@^u��OBY2�����d$�7���	_�	W��j�u��P7��܎�F�K�\Y	�����> �p@.WEc,J(duP��x@�h�8��@��G)r��J}�;�j�^/�kBUrq�^����H�%�d/_����7�^a��
���lF�1�I\v����֭�^��-�\�K�|c�5��c3��Z����h��"+̉�*��V�i1��I�ד�e���¦ImN6h����һU&��#7ި�}r'zk��g�VRm ��µ8Ù�v�����lXƐ:�̳ �J;����-vw=��T =�U�t�.�����ey�"�7��}<{�<�D=3v����35p4�Ӟ�Nf�Jf���D\W.Sz����S#X������������,�y��X��8��j���*\��F���Zhd�[R�׫_{eP�6��R�1��{����r���cL��������Qs��!|���oq�?�]I��7�!�.%�����Ӏ,�\����������"��X�h6��@0QS�$��� ��e_�!��=�n���Jc���S��jZ>mi	Ž����pC_5M)g��;t,�Ԁ÷{+��{�>��G3V�G��+(�������PQ2!<ZbF�s��\��2�)��>�v���.J#wl���%�Tt��ԑ��vb��,B���b���؁�@N�Mm�]�á����oK @���(p��d3�wύe��)0�߂A�4����?/��ǥb��Zّ�	/�%F��,�?�v_�U�+<?�\%yu� �Uk��/�4��?$)#J7$)�X�7���=u��)^Ԗ��b��C��v�*Z�4�c��\��S>�H�;DЄ�����Q�P�7��l�4E{��;��������t�������<BN�m���n�@a,��;��1��bخ�谼�s|(��Wlbr!���s:s�>pB�ӝʻ� O�d�tR�[�y��ʠ�ArB��y���[�X�������o8���B˗��by6j�u��H�%��r׹��nQ�[�wq�?����P/'_��@��!�M��������� �%��C4�����k�|�Li���x��@|{&)v��ޝ큅�q�嵠�[�^S�a�f�싺��;m�,p�m-T2Yd��EL�O yiU�}A��Q�t�0tM��ù�3;�A��j��Sa�:�� /j](�7��7Kh�"�;\'�䂵<`t��"�����kkpfK
E�6(wd��q/99�N;��͏�+:�M"�ы�U���g��H�ji4q�j��R#����X�go;jZ��?0����L�k�����dgp@�|��o�UP4{�9pTv&��a��Ӈ��г<���������̕�ιT���z1�8��ۤp�hx��=��$��d�f����L���F��:��5:ŵ�k���ts 0ݢ���Rm�K%��=���tR>���!`7���t/90�uaH{�'��p5����{+{�@A�����M9��a<E�L�{�"7��u�m�Qd�6���]��xo?�<ӓ�U���sLK"gV�Kˤ�T�t����MOo�I��TH��R���Y�f��V�UK��?
��b�^�r�֢��fY�p�@P��w�-�� ?��D�y3(/�^�x���B�-�S���@6Z�#�/��+�qH��=U��J���c�/.�$�Q"��l�ʏ��/FIjY�:��S��\���fap�����	=-���Ţ���.�B-2�G�Ґ��2Ŭk�z��wX}�2��{�1�Y����d	��m�'w���U'2��`Pp5�G��Z��9��MQ�|`HGl
"l����@��FC�����w�O��iN��Dx�1�B"�X��JƂܺ�f����YX��1�T�8k��KK��K�6?�~9F�j��T�@�%^'��f^3@Z��l@������'p��Z�$V�4�(k�����Mz5<GsG�3e��p�ȁ�.��,���"�䍪�[ts�uy�Ǟ�5�/*�A�&�����^��~�g�u5�m���04n.Wڲ��z���LdX������D
�*���|�����3Q���Oh�Vf�Zȼ�I�,��zp��+| xp��S�_�ߺ@~]�t�+{ ��C�����C�ŧ-�D1w)i�Yt:?߄��v`�jo0���D�W�w�H��Y�+�́�&J
I���nh�8��e����(G����դ�xu�����&�J������	۩�ۛ0Ê)ݎT�O�%�G�;08j�E���@����(F"D%�&2�_�D�X��z�.29��mF�y��OϞ�