// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Dq7EL/AvLsgJ63vyIW0tWDgPPv10FREFPLfASXjSM/dvolEBMnIisAnHFrDFohu0
tjUnFBzJPcoaLfGu65KTyFFbX0upX6gO1XnPdDxmDDEWPAhez2RypGQ96xBqBrQ7
2oEal308DFPfdztfZshNd4NsNKZIgtkj36CSTdu/O1M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11392)
PpXW2hoHa3ruN+Ft6QI4Zp5pl9GC5sOSmjTiSJaIBfZgB6D5GVj5Q/gZTjDQfQat
9LNxXdRp8lLb5FSxntfeCFkmnkhnm3Bpb4mhDKXrJKXtjzfdTQTJY9Edukuaybr8
HFIuyIqPkBI39pLGpKhZe9Q/ofIZrlf5tLiK+GunKnS/Zw3S2yRG0M4l2ozAsrbv
HD/J8svpakjpxo/O21I28nLhfa/YtY+bQQdydeMXAnIaE6rNfy71flWRZ6wgc4xw
yod76rFhjg47P6xkpLBxWCqb69wuQTycCKHPRR2UXFPn5CuMhfdKe7hG29cz17hK
pS5WoNQIlq8YuJv875NgLcRYW/9xGD3veWdwJMhKwlksLS1QsJFVeGvkiKs+tqf7
jXLAzWW/LxhgD6OYUaK+h7DmGV12GuaF3XRV4CpAYg7XNnzHKmiddU5W7mfa6Sfh
wU3OGulTKKuAHH8TRAc83mW/PMBJFCQ8cucj79L9xxXVAhWudFkZCULqpXev1WXR
UVUg7/Pp0Dhw3k2++bJqER+iuR4+ajdrso1u+yJhMtkUnryYKkaMJweLd7IH7pUN
friAxNhhzjwVypz1vvHOwqz+DNUZXjzDyEmiOG/a1Cq9eNSCBrMlpwKagKHNx1YV
pxYcspL0xx0Uj6mZF02o/y1lznBl3raxLIrgJoXtd9zNQyLPdew784nBoJCcMCMN
z6BZyFX64WmEa3pqE3H2GNaTBTMTe+kWI4nj46S0iR1NlQimKLKrXCgInQGIqT0K
V1Gj1AsxAtYezL0LMQ6JObK2eWybGsSiSnQsuyCjxwJ47Sclzs9zTVhOc4wYvevf
OPTfB7HMKObLgVP8zaM6qRjb2Otk/OvokgJ/9+PSBHEs6qrPMUwB6f1do21nd9Nf
mBUtvZplmk1O5MgTDdQ4wbVVfgSDf20ukYUb9EnM7dXkOQZWYvbY1iHSpH8go0AY
F8+vg+jHXnsFrFSAht5XU7Hi9fL7Hevhr5ZaJAY1YCypcszn2R87SRdtduWjRAoN
L1cW4Mps0FglIde7dalF3l1XsAxpyHQCdKR3G2otOrgLLLAgVG4Pc0x0yoIoNFzB
6/F0hN7HjyB2GkptaI2hcxO9n/gLfXUk6IABPsaDBR1DF8teqGAijgkznqRCgUTX
sHR//yFIOCCGiMruBDC3vEwWhvlALIdBITl9iN48aY9OpXSmcNRI/ymfRiTKmH0k
5TZYNSLg5txpDe8i+sJlZilIepWvkqKfUVyzJ6tp1BO/C4BR+YY9liSkufFi5sR9
zcRFDl/CvTI6aTj1v3K2IPpKDVybhQk/5acgyT0R9+fEvNxvoXJX6hS6u3gFQqyu
kK0lcZuylQQNuZ0qXtauK4K2D7cPl3VDTF9plj254yVRK69SZWNoISPfdg2FiJze
PJybLeNPvRZQqz1HgK7h0xbKJpNr0cwg2i6Bl5rGaSe11wCrhHRPM77NYRMGVnfs
R28u2EAUZTBY6aZY8iltidPQxlspGQd4XLGUf4qbXeI8CNa4SjSfGnMkd+H5tofG
GSLuArb02X9vB2PuM7OWsrvmcEM17bWzf9EZeWkDkatUadIBO47cBQgZxcoA+4Lz
Xu96UyBL5grl9S2FyGQLEpfnu9rksk97Z0SvgDaDZ9YJ1k0bn3Ks9UkPpk2YAKx7
OJWi0Gy24LjqapLJzWlQOcNdBkz6NlX44k1hYBh2UorYnZxqgo7ysOfbUMj3qH4q
f5BIXo0kuiBe69mAnKfBcgINFcxbl0f473l7kLFU63J5Uqr2jkpSDZSZRmJ/YQLP
ezZOa5PiH/OjUQtEVC44405fTB1ULxZIJQ+vzMr79Ba1ZyrHyQlYdd6djcKSGs0i
r9atTtnTAjMfI2+3026DCc0gnmVP6I9SwIrNaOlDnfkDanOv5d6XsH82SYdRJThC
IqmAd0WT2kKGbRy0McCjljA/zKu3BFC/CxAwCb09nxmhTGRhIfP845DhBCGOurQP
4LNhTuBH2r5VlWzwVIeZc6lVE9dKxVXfCPY+vm91mtFKX3i90LBHFryFGtKlL9fW
Uvo23lvbni/+vIYWp64twEusVoaopa2zl5JbqY6S8GoP7P2DM6zWKt0PwN9oSc2y
fWcx7f3z2xJlj25KeMEMPCZDF1gWVTL0h2uCULwzoXWcDkPGhnqR1TCRCqeTfdzF
wrRLjcreq8UlFa8cf/+0a0+OhoYVobOQa+ovfg5wdyUCRGFDhLDorDeQbBkfBXIR
3tRzfHdNH+nfUjzE5jzQMvqILRsD8ct2mUryS5ttfGvu4n+n24sGnEMSaf60BH9V
ZyLO8QZu+sdusaHs2Sd7ALdeHMhnmVHRsGUd5bKvj5pseYpaF0XQs1GqLbEnGGbI
BpuYNPuOimg3Okpz5SX5fkrDMIcs84nJUr4DOI/xjH+wvaP/718/7wbp9UnhXOZ1
6FnBnYun1bpJrXsJ0zWC0FuCEO2q4HPR3WdhUWd21XHziWuZIW+ejOuF/7LnKDF5
BrNUAfaAYvSpKdwxJls1+EQFPeny+53rZ2Oj0F4Q+Gjz3NhPWz5AbbrJCzXSdmpL
bS5FzhlRLXqniqL8zy2sqX16l1RKyiXkse0dYsaFQgQexpGPN3JzDSFC8L1ZLQux
YgiXZLJ8vat6xHPUi19dcZAn4eqRuwX/z+SrJfryBfQ89sEDM4UZ0c3env+9vHX3
Gtksm3ceGwoBlGdYs+Z1UgDfriYlbf9fD9KyoyVANml8lYe1FCDGr5+r/5V7L0ay
Y6vPUqF1p19NCZZb1Gyk2LNxnsH5pKClOr/GNc+/po5Ll4nmgbrWNRIN0uLtf6Rm
2cpF+Y1kmK7u6zwyQqQMb8PBBffq6TXFR9acmWhvrjxjWBQJNyFN2iQqdrrTvmfh
UVT0e4/KvUbJHaHcAl4A77pvvHPREbgzFEcoVCyZeiIDt/+u1nXoR3vS/uY/GrdP
haZUSRWBDwU7qIT8gn3umAVkZ7hIfQBZPXBEby7x54OzDNf9EKciLyUdlX5nS+o2
yQDfiFf8uhz8Jyfu4AFA2Intzs2da9ZkdjpCIvTwivrHCrWIcHHp/QeZQubLXZo1
D7mLG2+c/bho3QK68yqnaCqUbXdCRBQfE8G0ZSDcPSzEi6QizRrrEIoOItMLFq7u
8pnakq7kTZ5oJDb93UbWkPE2Dg3WrVViOEwmN7tLVuFE0Ieop5WH32zRXpexWtu1
Wv4Mlx4/nX9y3pYg68jDL8fH0yPc4pbq+pu97AvyHwOPKyMnBdaZV/wBIRidJLyq
BeUTxGJB+Q6FvYhGhUDnu16/O8lKwvXY5WgTofyxSw80xzFtIT6DNSH70rVp0pzW
BbjrzB98o54Kcx+mACaDiBKBHYO7+xGnHQd5vxArP13UKuz7HLrT4vsE9T1jfHE/
1EESHxwbSiwZe4GrSwdpyRBxIlGUqU6gTf6lYWWicrnkLJladQ57NcvNFDpP7Ajb
X9yz7UHgYwiR+Sdur1Ad+jbP/LTnA7MsnjSkyP66obwn4qNa8Y1WRa/wOpDKwA4r
ntmbeXnuH/ZF93uYgQh1pR3PeG8ajjJJWjJWo7rjQZ/f6/9icRf7YPKaj93Yj4X/
W8Svo3wrNuE8pc6F7Eiu0dr27LtQ9hMo5B4OqPxuP0BKqMFnKwVkLN+b/6/uDlhp
u5KiL+Ue7LYdGe5xBLOr/dgobZ7sAAV3BbmtQGmSmKvyyWxX573zi17a2WgWcSSh
ATQGujZEsrwblc6R8mewKd1xmNyc7bCHyFk5mv2mgK7xwH/t0EtgdifFoI5D4/H1
kzQWUl6ltlQNPO0oIEhWUSFEhUEjMBruQN+YkGdSDbVrhrtdthf2rgWgUuAgJoFN
SpL1mAYs/eSb357noh4H4VhDJmDfUuAAb0X4ZFpvw7PdAB11Go/6v04q62idQpSd
oDXKn3vBfyIUdH+saRwTIuQC5W+l0o3sRSwY8eL8NEjr1lAU2Q5xLNpJDNMCDh6P
eN/ca4Vjm/VFkEomvqI0yRbj912GxTPH9yP81jmuGR0We5qw1cNFWGWpbFtplRtX
m928AwFMO5PHSdgzwq7u0Xl7XX/hCv7vaBgrhp5UYbG1XBtqcnrEagMNurPjVHL0
Dl7URQrpJBTtVyjeFd4wlNNSvTwJcy7rNNXxLpcpJQD0mMGqtq1VcKBLQK1kI/HS
4THxiYDZCRgazIkqbW45+w5Gv2OuqVvsTfhRwdPBO0Kwn7/OhMVZmnLZa3sLgNuV
/rv7Ot7XKZPSj6QKIjzO2Ee3DJB/QVcWCdlFvOh74cHbwNSkpLUAi79FvxjO6Qod
XkwZNjLGJNY9N2t/2/TiYZcCf+Es8UCIPTwXVmKmn+V+IxHq0zLtV8m3vrGltF1k
BpeZRePst62EE4It/zY5CSSlJ+vXT9UD+hjefy2FSM4B3WppXacsJY9Sh4Mdq1lE
iLV4J1+jYRkQ7qvcL6USGgcRDymo70NpxGJsQOwIsDef6oASAjknFukc8tYkwloS
L94tyuy/pDN7XgFP/vLjikcKAHqVTOtn4Fcr+3b8E+hoQZprQGCgoao3DP4yj78b
/2Zymowl4b0St8B8WlH8yva5GBwNMP7/xpwFA5ZbzjgtEHtI0NYva6q6dmeYjAD3
L8MPe+hnnhXhGDWPq6SqEfdN4AUIQw8YC1Yo5RsbW+x9CDBL+8/ZozveJydU+1Az
jjhyDCLaTjvWCmYulMBU/r2ZpUdmbytvOmRAAoDYe2GrB04Ew9i/qtdc/vi5c42e
Wy5jZc9b68pYZm+IEMiX1Hgba7JyQAQ402wxbNTpO8+MFkqAJr4CQ7Tg4LLBjAuK
jXRcZX0fpT7B7Jo1nGEnfbSiNnpuskEZdBechoU6VLi/JOf33B4WL4Zdv6vgsWoL
xYiNOt6vXZPtPiwAWdEzW8zbj/QrgtwXK6dhQHE+uSEjyDILUgxNF+ovNIK6CWjA
RO1h9rymcjgVSuHnFuRi8uGVrwAK8Nj6n0xZDBm0wSBA/tGawQqZrANJPZt/OowZ
QA0NO3RHphPJC22LqYH9Nw5iLdjOEyRnBevpKnYA/YtLQghlzaYpIefhvVTegJcN
L/nZi/GyN40dRpUfo+7D+QQF14pT0PHv+0MV6lCCOZes8iNY29fVv05shyfWcoNt
C9MCkLhPzHxR/8oI3r+LoG3m7bywvskXSaROaqWQWp9DGG2DLvKOVcZlk5Rng5UG
YffgJJhc5z2NGhEIepMG6u+P0ZgUUcbdtB8vtKeM5zQWR+GsERRTA6MnBpbqnu9z
Ygx9/NFhV/1liq6bh4wg52JtXueXti590L2g2f/AUQKeWxhK13+dSlK29LZWZ47z
UUvAFdoXMpUN54Ynv8Scq6gU/Io68+NdTjFlxRrr5HwqLTUJh4rqZafOmEzQsZ4/
TExwOdV5+DXlojKDr6sZM/I3tGbezCLvkR1/fsoGxZRES95FK9olAl3391ayi+TG
zeXx0B6RANe9Tmk57T6P8FH19rDOtWNGFnLTlDyOssH59fnb8cBTDFmNwFqUK3lq
4MbXzphH2y+QDOJkSMKorE+gJW5B2Vsd5EiNQVqm7ii4OZ0oyW4i6qZVOu6pATxx
j8Uw/GCrshVZCSn9YVGm8Hpbhm8Pib7iYA0vMvvUINmWwQXG4zEj6HL7Ad0598Cz
xbQFY3NWnMsT40PEAtirJpJjw/nryTxUNTcLmdeg46rw4DB48/G46dQevJ1hL3F9
RBNGZgCnLjZFQaejsw7E+odAQF16FWOWn1/viQe9JRIoWdfRvMqTA6s7RWKQhOyT
A6a5hYdx/kTEU9SMY9OcfpaXe7WpgZMWfH4vwFvbQaYWfpV5dOzYrlS/cizdADyj
GN/NVLkTFevHJN/AYA+XwoQG92tDtek9emuJeU+2YharyFO1TqOPSPsgwnMTSPtd
NtdgpPw4oDkkLKb9ghCqu6eGeJMb18ZA/OEnPHKJWfyHbqT+mNe8j3SIAKNE/1Wh
m9e7UQLlf6DrAI7cFGniNAJxayvQGwDHyGNJspHeahg2DPobP8K/kKXdYEKDz6dm
geH1DN56SmKYI4/twWGTUrMs5GGkj9gp4FqNhhQJdNV6p6/rOkgqnIq/9QeJqi21
1zbtmjmVyYlG/HYi+oj3cPN5eVXWPd6Nr2zMNBn4iyPXYd6pdXGj+GE9m5i/hzLE
PURaEnDvq99MlJaDrp6hyqzHdHgAQzAsWQaFju7yili4+K81NEruCMncx5OqR2zA
Bf/a/1mwUCHVwbEL6uiRpkef5iI0DcZrptXpPvpOjp3WObtJzYHN2d8f+y2naj1B
WlQypZCp3sL8pwU4APVlNJRmpZhOmtROGW6kr+XMQ4OQ5kDmxtK71swpzldHJcdo
Nombj8VyF1vU4ub/hSYMxpIOkaz3Vi6XGk/QYqqd9Ynb74Dl5cS4hyuebtvrHYea
UbmNZ/X03OJWMg+RlpogzCMYMILb6o7aiGUSfI795yt/TbUACYPRInMPKR0kdUuJ
xfwyRkO24YfO5vG3l8ZW3u68WvU3wGH/r8EPSQ04ar+D8a35jdzhPp+2aYiLyE3Z
E1HBg273Qcr35r38Sack7GHakxNW1Yxc71XLC+8llKvs2mscbZeUsnrxcgrwoSOl
XbE70hQWzLsxX7UTN4iaKtl8YR1zLHaRaofe9RP/6kRGEgKZiekp3p8MLxEY9+8z
zR4wdbsG7ORQqed9lVAHKUEXLRwIr4jzpCWrKwydhNiixQgBOSEe5fyF+AQot4YH
dvPmM/6+0V+DQt4280x0mEPJEd/GwHd0fzctwcXwaqXCL8gHqd41nR11aEQf37PB
1am2rdaLRhOtFxJ6OrwLer6RXUtlQ6YcbwshjGR8GWvWsG2BLQEg6K2QQXQWN5jG
lBTcpEcvnT9H9z8yiaIg544UBZcGH1rC8Rj9VwjTvDt+A+Trd0RVYsIjYoqDWJlL
EnLbkqrPq7NPIBRCZ8ESrTXG+hlzSqVpSTcMm63WvwkWP7bT8bYqefAek5kcb58+
YPGnsqUGzXOajMgwA2KGiQNblRBpxuR6W+tWs+eU5cv23Xl6iPOhgMrmpfd/5KRj
Hm0YoP2voephg23QSlJ/jB9aWpZGDmd5jgZ3OPw8vzwlcMC2w7VQ46O8pWwZUR7v
4ZWocENhjlDOd7XE1RRDz2HQX1mTdTXyAwDGnMWHmP60y2Hta0tJIKwYxyWxdark
4mUm6RUflcR6Gwi1OjWJoHcrPTGZcHlAs7U0BKm5BXzzwvA+/+b4TtOLTeqpH6YU
QjeDZJ/PBk7TE/2G9nLAefbkUTcYyknM2Q4GGcvU+J0KsD6fFAT4wzEA1rC022Q3
O+2aOECXoAigUeYp7NUHPo/Ep5i2fujyBXGYB6mtVDPB3ws1R5f7vtgANNRauWMj
V/aCtjgW4a8054UAWUkmb2tEEuuJ9A8mYBNlHbzHODaKf2Tg6StSPNgbujtJM+62
QVk1RlceShZba8NhDk1B7jAoXLZ162G1oc3bTeE72yvcn+etch4eoPQhTqERzJAA
5vKCn9UxMpSxv1qC2wHgDRRcFhnQ6GIAzgilcUdHdrrRwGgv7n7nycFAZnOJB/j5
UYyOhsBa35RvVJnZQju9jXsLqsCTOcexGPg6KEPC8T8mdTC2hbJhR6qd3l/1j0p0
IUL9it4q/LGsRpn9C2pokCbJA12HoaOn01nH4m/3JYW6MQtPzFg8voEcs1qGAB6m
iCwYhCFqjg2nQ0MI9tmMBDl1NRIl45Z/b9WuNjbZogXi0fYFURjrkrylKmT+1Fhy
PWuWpK/r8Fe9T2ML9Hi2saG0V1ZDikl8HWWbPUx48fMf4KzPJFwzgHrFOMDsVBjw
sU3kueUR2APT/eWubgMnF7Vp9MtwV9FOqBhMd49FJ98jwde9BInc4ZukX2YZS8lL
2sV9/DNcuu6f8fhA1liHuS6LXXTIwFO8GSTiplu/iLgrDEfzquKdVGd25bQMNvPC
4SVjUZtqMrbb0D+vwra2u4X+yXW+tBRKJ1CXdwJrGGngSvENDMAJ3mIUElxkyls6
22hVuhPPZ/tNPW6dGBUXz+8oOQ0LYEBAVGObH5ZW5a9cQAi1fHfhL4iCB8OMY0uY
Bq3ScYgd+AMOSicIbRfC4Dxd918cVFbuAHebV3pgFS5MtwMC3qbTq5XMVQDs6nf0
XN627aPQSIQli+LfTuC9BqVUlzfS3lC+l7/chmUny6reBxtEzwp/lh6NmNhoN7Y/
LS2DTscFiMWy2rthsBwTAGon//fNdV3wBO6N/6yCRi94HNmW2b+Lkf90GuHltrwx
PkYE9KRWEVX+CVT145IifvBLcLna3Ak5igKPPBIMv1Oa5RwrvE9qs7BGlFbMdaKA
Zl0P0dxiw2kIn5PK/pSZGraHDV2aIVEgoYZfUf327lY2kLXxF8VqoBAgWeFto24Y
O3VlHllcJ5MZw9747ca+hUepP+FrvpOqhyD+PqAmg9SBC2ntognmJ6DESsFQClCD
r+UymmsfHPAU3G0xr6p+osu8+425ealSwCDboAzpjgmnzN/mmm2ijeewDt1Hs3yJ
LOGWEzJcQ51t4Cjz2SM4zKrYPZAv6F1afp8b679G2EarxVdo6XJ3f8AKHGmd7c6I
vi8xQWkkpQA45vg9ay4DIj2s5qlj/D11WkF2GB4vB08cd2SzI6z3BHn49Z96ECGg
wYwepRnYEJVGvIqAhByGwRD7qr3woEKvh6IX38F1nTNoRvTBvDCvL+1ylGXjLS7A
J2nSmrVeu3hc+WGFFFv1gqAnUnLSrLyk/T3wnOPnRw2nZLx2ACTNO/FipaancFV5
hCMTkY3ai1C8GIwoZYL40wXIpTY5h4vKDF51KrNsmhUnc+yvOAV3OCns3urIFfhK
GndFqjW68BfIaX8rgMg2dMkmlKD/Am8DXQIKTnI3fsCEC5tCm5yABXXEWMjVo/qf
bqODLj+V4SeVNmufiDh0YUyQWEKXixOWTGrggYv7n0UwtOIoLdCvWsjiVqk3r9nL
8JtfGK7skEHyxQWJ757G3zD1ciohSt2m2r1wYS7mvSxHl2LEO3HqRY+o+n1y36OF
UbH/tpNFbhlAXcGRkUY1ynQWpmyKCeoz8BRZHqFtcfvN/noo+OMBJO2J4Flx2mwb
d7ECpc7OzeAZIn/uhzk2dPTzdl4FjzZdn+Y2pYLiQuHjBUmU9TCULTg4fSLle/DG
0tW4+03Lm9lf4eFnXs47zHBooSC42n1Ggb1NT79z2PnKlTKIP206ROeTTqNQ1h1B
SqfSp1myh3MvhBpg5HfaimcAm95U+nmIZbVeg6t8ODF5GgNg8QSErJzs/R1f/rNJ
H0XBa0tIlJ+EyIOL0InFbnm+9blHZgrQ3vHz5mSm5PZKAHZfxjn8PN1PIGLJYZZj
43Gtomt5Bt2qupiYXLM2eSLf7Faw77+BgOrS70rVpvOUODvlzGsrTQ8CiE5bPvKG
LShcIvob1QFpSdzIotae/fmuqyKcyfBFPE9dLlVFkDW/JaxvUKNoqVk8ozJK1jHJ
43vG5XgBoUtCksqH9ZPzl21C/5TDMQ3KPsaMBMWy/j+Q8zLxowpfCKOZ0t3ZyuT/
sOAX2DVeOXzCXwPScCAfy/d3GT39Qn38z55T8oi3V2nceMm3Ds2Zr2NkjIXBj7e6
DHwX7xjlphArgFlsQ+0avvKTQjJ9SW4hLL39CEOo9+p/nQH/3Z+J2UQQwMOvUc+p
N457fIER5rtAxMc40fs51j1tu7j6hwp3xsVS+TSKcBkEUcqRvlWsC3o79pchCYcn
IJtGlXCTA2qhRQPI/z8KsrPsyk8t2an2in+Kk7EcV/awM2BO2sRODGFE3StJ77FO
YTViB7Qtx1yQLJG4F+DqZlhi3n+/tT7/+ahD/Lwzg34N9KCFCyi+ckL3YfketLHk
cIiSGm0Ch27x5DSuOB7hUJ+bKMImnVMn9kh+Fdk9d7tzhsUIQP3jDmmKzf+AZ7jc
ndNHZzT//0OUqfhw4iPLYQzOYG5bz55XMMRuwutXjGlpamyxVm/FJtE1XLxAi/ZL
r3nH6oR6hKNSghchD4yhEUt5wDVDQ98GliE6QsFIAWRraKP2mnyxfdSgas6n5+cR
BE35LSTYHcvyvqSDrts0oRSqvSd+GlZa2FRaAvfrLHGmJc2R85UOsTFHv1qbz1pR
cWs4lCS32g9oz9WtpAlgCLEwX8foVpsh7oa+s47G9VgoKOoMPHPHs7kEK2DiJRfH
QOS+6UetQ1zWmjP4Yv6W5LXi9Zrwqs1w32bbEDAPQvrOZT4u+3/sCC0O7XzdimqQ
fLVAfRRjAC7uYfzg9kluCSp6Mb8/TiltFhFqn3hBQ7lVPc7CGBKgGMA9FHItc0u4
mnzxKsd1MboPipBzvymIKdALRlxyoQYA+YkczkIqCSqeMHZ847X9wTXtbElUzhiU
fR4KruHmEAxQd0899uptfM+8AhZZ16Vhu2I1L2vUDPg/iaG7QxbDxPjArKuWxAYf
QwgG0fYTYBUzwqOU1x099pqPffxZ30EsLjJyIkkWk0qvNyO4LeuZr/Ldc6nXVd8k
5SW7gRa2u6DMqUzlSxXKRUw7AVe3J4iSXoE1Vr+VROGbWaEB82I65XB7BuiWxrEX
7VBXZZBDTPUtU47zwQ0/HpXJpVN3bE1oYIs+cOxfow8xpVuKx0o4Sf4IgH/Cbt7B
EsUD6F9q8Lx8g5lnzTebozIEUWsJrAt2wjxv6Q3R/vibmWKGrxgo+74TrZDWFc8v
NXjGejgk2kERPRo1sWSOoLgeGgRHzFcyvEeFvmW6c3cYHu/7XMpblfjEEJzAXxCB
uOZZUWLyC/AL+0jeuslcd5R+9t7BujPJoe8AhfpOpynXbQ2KFrGAVlmXsC9ANXXe
MpECurMNHHGCD59SXMJU3jvd1oOsNE/a6HN9FYT99c99TC1u8/vzBOVhvUn8eJa6
Q2eGVhU5zj3gl+bRlg7fhz8JBl/pCy3L+bXNbQ76Nl7KNEc8cjaUl+OnfpZbd873
aErXShse45i2r1/hLVz3OZaNnbhGBOrjBZ5TDvFzRjFM5CvdiU8mfmxJVceYuxHM
loFkeoL0UXZG047EkwQKQruUp0RkBPk/r3TgaW2GDgc1FjOTBhW3Z2hD/vGErPyj
lUw8GggiobzLNRaghOczGc/U/PEYPZ4iZC/v9RQNThVR5gec+ly8rv5mObu/950+
A3BnDdL8rLOCkbtFvm6EpkZ59FB6unZ5/Oi1JYnzRvvKnzv3CXxSeWuyhCe/NjLs
8X8WJEfkIbdfRVArdGG5YRSpILzeitizRTK4UKqO/azfQ7HgL2ssMGdk++6kFAzj
gWpLNSYLQr0D/ofULkAW4q1f6MUm/VdInHJSop597swlcAf4jpYZlL+NWpDGGUu3
mBlR8Bjr0jgWh4Q1nJgHGKS1IlG3ND2TT113uJ1MDa+hZTflC7CwqkzzZMRkqqO9
VOc+kt07SdsPQKd0kfskIkGctvD9vhsAB8pYqYmSV6uOJcBQ6kp4kCyySnFfyRB2
9GbhSh/IuC8GEehcQnz7+rTYijLYW9zbMtbuHOVGCviVGsm4Yg8kGKb2z2J67Lmw
sWMwTAw0nYg73sY4jD2b1y+z1UpQ/S4fTdTajdjzObH6nex7ThrwAbNuU5toGBTz
KvNVTdUF7h4wofi8PPGiundO37jd/dnGNFEKy6nhq1c0JeIYwwHC1cxNc2tc0smj
4R2MWyRg3ivltZNSfmSe8rSxMTyvkKhoCl6GHGgBXCcr5kDy9+zyQyjvlvcxYiGP
bLuRh8gtCBFCHBzKR509OGtqqcx4ZSji1rBCIE9kOv84Jkonrp8N5EU/4vYfqJRS
S6wDq14qo6s1WmIqnoKSWTeiLsoAR8O0HHAFS7QT9Qzx71pFwETeUK3xue+pi2XO
H4HPl0bHbqu+XtkAKkOWZBzjDJOqUuCeJDVRRqqfJbekB/d/PAYGdw2ZQgtxEjK2
BeBE+aFjSHzg774jU6Qg0Md56qbkRlvC3UP0gGWDA+hZrpOwsbCpwbJXLIE0E72p
YUh7IuYJHNzKB/34JgeRreOnQu8qWKP06wl9esLBbf4Zr846bAgufte/Ms1yGfZ/
Ee5JJlDtI1PHFUaLPt7gIAaiq5tCkqSaK73X8q5ywpngpZhDYEj5FBbfj7CsOkXi
5p9wW0IzKONkhzNSozKa6gwywgJ6kzpOWyrank/QRwUxevoDPzSdnbruHyuHJIvX
H75cQYDGJSzjrHf//ogsPsfSbmgTx9MZpAS1nUxwKdNY3x1IWaSYlGzoCRyL2mqH
eDTc3vPpJeY9H6rtV0WiOKTtonWHv0mz7o/1c0EB6y7m0i7hSYVjKxU0y3Go04zn
qvF+aeKYY7ByPsWoVwPHt+huU3xC1phg6fE7/fDKCBqzSzUwMKPERWmbQkcINWfV
voQevQt8RidTVCdycDGn12TZbJCb+JWK3PgcHMut3tjBqHHpGKwdr6OXe96Qgm1u
YNQNwvPF3MJ5DGvE9Tet3j6jZ+/NRTkAjFW3HggsRzOcqkK5PGtM85ITHhqEtYVp
8frqlXRMIDLTtXY0tgrW/KMFuARhSAPF4+emYA89g3EhMt04tL6ziJC3DP/2SzOi
e4XKYFD9qfcd1ph5wnHCDevEwKXin6q4q91OQq5cdy/AEEDdSeNfEuKHWd9YYD5J
1jAkO4w+Qauj2lPm4q9iNk/F8JqPcVLFuOTjtlgpnx1CPhANeFzjFS4w+fuptNgF
lcQBvzsak0iwErC6vpOviaZWyetfauhazf/kOW3uTORVQAj1M3dKk24ZJdMq5I1o
jlFd7jDDCTLn7dHdcORI4CdLbsRSAY2LTjXfaUQr+DRAVctiw1uf7JWuL/4qK70u
6HNWdZuzvcWS8MI8Hmt2NzKNuisExnSIapHvAm5V4FKUpouesv7/l8gvKVVMnIiF
H6dSwwzIkA5AHRfTJkSpACAf1nvmVUfoOg4cmnnDr2a4M7xKtBe3etJ19fvnSUKn
XWOBI41IzzeoKUAksHw/xFNV1awc2UPyj88+ZYdRMz/sP+xD1gSseahzoigseKNr
Ip/WmlOW3atdXId36Y4mNEdOc/LgSOsaHZT3SAeCuUeZxisnFZZzp2w1kaC35Ct6
NGz1YPkzJp0GHLk6YHxMsPuXOxYMO0c2ptqEPeMpBElbo2kuzyp+i24EKU+XeH/h
gRKY8QOrHpOl2AeCDZT0wRAogwH0gA+1PWrwGxUbtSUeiS+4rvJ4/c5z0pYlriD9
Vrj6DC1bBi0d/pPJ2AbHiSzMka0Dy+ahiHxVBinnHuODDY8tK7pHyoHky/mNj7TD
eU3UeFfpNnTrefxNCF/dtaxvK9K6m5vHlZRymTKSY/zEQgsI3I/JNMOsm8EGqTDq
9NlnVAz3Cdl5VYLMNz8mKQg5+eK0tSYwEomJZf9Tzc8GaZUpTvpruabWrR2BMTNU
Ga2iG34xicd7g8Owb8PpmN6l+vV5yhevvO4nOicZwv+rtWuH+30QswK6IrmFwd43
OBd/MJuCP0ksXjIuPRoa3wkbCcQvDEH/qRM497dTBYHgSjpPhYG5D6Ssv4AiSeHa
D4T7hNfiqwUReA1W6Whl1aoMEY5AA8ZGsFvbT0N9fINiMj+FbD8HMFkDPFncZkD7
Uli041Pozn3tYFw6lrWqcvBUS7sqB/LWzZNpOVrvzSBAGeUWe7q2RxNf/5GYcpW3
OjttJw51pl6L4GbP9zapzNdPN0vMYpwEuy3Mbxkc0iJvJvtWC/OEXwp94BzBqSwH
pv0tq0crAR4KvSgI8t62lC2Iow0m0HEzPNo1ep7Zuk80DjJhERhkWXtBF7vAfpTp
gAWQZYYfJb5L/ZS/f57ksI5mQP7EoxNRhBdZlnp3OojYoRuePfY64wYdYKyC+FsQ
k56600QKrsVC6nblUlRm6CVT+Cj8mtbgKd0mmW3vEPOzZr29hkKeHI5NnMdHBrmt
ko1HUxl/QVG51cB+UI4tJPkogVzYrKqyRpScyE3Vtk/tRWtHbuZqRlr1ITSldUWU
sIlRdWQ9OgKjRfDtPyH0goYVdY2aib1FtWm3hslbBfbIvyX7i8+5M51+H+qrqJd6
Dn0hhnBik3+PmpE5zL1H60oiakvx2Iar6I7T7XhSeGsyJ8DvbosACHNvhbBJbNl5
Xup1syLR/uUIU6fO4S+gTMcW3VNyReUGZLvU8sVtp6DidzqFeIUmdNVSOmzmZJrX
x1EJebv9BH29gYpEn+XoAlrWSSkD6ZmEWeYEGRdj25vwJq8PCWQNuA2524M7NZlJ
enRk1Bc74IShnICJ1CGgyIeY887tQtZci13JQDOQZb13wqefjWuhhcSHvZYIsVuZ
0bJkOv/Fwo1+j3ojrRlmFeMDTQq7aGR3t72RdHXBJT7SgWEV+wUENLllDQ9FOuBF
iUYoVRaaHZmHgSM/zlKhS7u8O8oFzDuR9Su/xfo6hRCc/lYEkPwwI+ezHmUuU3Ks
DW1urxcwI02mfz5fO+UDM7QQjfc6Azpx2Nu/CQLatTh8UL3+r+qJF+0c1AaZG8HP
6tmZrKYavpRc/kvyBsVh2KxKWytfqwltw9to2Xb72T4JoyyC5ttmRzFoPfrFgvqe
yTaVut2xkGXL/ycfS0uuk0N1X0mn+6ZKIg+PQzNItG6WVVQWo+vR0r+902XrHJyS
v4oikmlED9CGz5kPLWh5jbH8q/NbHNUgj/peSChPghQGm0AJbu6hlNPaoq6ERUqO
JHlcrcqzGjgiSJIoNditxVPwq+9n+MwlxvL0yNDgYFxLss4FaonxPiE4b2ioH5HB
Wfj8txn6QXfbcZuE2DIPKdknTpWahMG8fS0t6g3Mv3Tbvuti0JN6SNvLRQTzgy/e
W0LBZ3geJSQmI4gWCRuYVEe5j6+ODRAEQ5xvoCqkNU3UMOxjBjVQhl1jWmbFI+vh
tH3nqOpNpYYmaUJfDkvqaqx6JF4afNC03BkkSmrYiTn6fhTq+E4mLOHEDHaHxYyR
EclA3GwTjbEkQRbXA6uguGHaxeKfvMRigd5p2hW+Q0RDcBwS3NxtlnHEA0eUpWYI
h00iK6YUz06G8JuaHBa3OQc1hszejXpW6ISnMq0z671pAoEOopWL9NHM0v11yA/F
ZGIXxqRar8fQt2IO4GLzplhlQLqeMvAYU3g/xfkb5N1xXOtS1ONTQSoDbVTvBawk
0f1o89MyXJiI81MnvAU4DcT3MWO3aeuUSlRvIj79KBdupvKsWCmJbvlc3FyfVZLk
rvUKrV6LZ85icuC4VKs3UA==
`pragma protect end_protected
