��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbж��ъ��~���=	�2�:fg\V?nJ��á�_+���q��jz��^|�|~�bX��2�[���|i�c��B!;�j�״�1�r�c�<���Px\ƣ,�t�I�q�*x�"���i��3�JH�b�͙��񳞛Y�UQ���iL��'�.2��Ā�e��,�Eo b��ۅ�i���_O��bn�%F����\G��~�%*P�3J9�����(��N�YNH�ж�\p[E����(4�8�4;���u61*�������F�ؓ��*�mI�C�Y��j���Z !\IZ�T��9s�-���-	��v1�J�E+?��g���0u�u�'io�W�v��H�gFo/���I�Eg��&��R�s���Ǜ38��C6��2W�Eґ&����P)�v'��lM���08>,��o)P�z4HN�R����N�Ꮚ�_�����غ9*���\(�Ô�$.�Ы�]���2d�8�t�|��}W�O�O����4���\%d�)�C/"���1n���a��~���m
���]�pӾ7G�������θ�[$�9"�3C�'�dvK�.�|�ZT�c��nxEm�0�?<�(e���!�#k������)w^�\�W�}s��E\V�XG����9+�S��Ƶ
��וB�F1��[������G�s)����}��ƽ�a��Wy#��VNlp�3�;�,����`7�ٽ-i�r���ԗ08�x�c�%��z78!��6�ύO�]�^ �-x�zQŇe�˛5͔��B%hO��		�z�6����T�)����\ռ ��=�5NzPdr�04�7=���=������fu��ɨ�rAp�X�j�^�'��Q�z�F \L����Z��M	3f��Ψ�Ռ�(��,�YN�t���p���ӎk����4��c@�,/�@�Z!��*�KOD�QR\�Rv�m�$���F���V����jg�zjьV.b���J����7��F�~}h� aß����m�\�eg��Ѳ]̃��n*F�Hqq�`��0��4���F������EF?`/�ճvF�Vf5F��Q"��"�v�N��(�﯈F[
��YV>��:�<�btu��M"�%�F����W������ܗ/<ɰ;�;پk��hjg�Y�q�vD�%����h#/�Dj|R�s�6.�k�Ni��9�C7Q�-�J�w���:�1�]4��.�!W#/��@�w<E ɻq!֤���I��Ȋ�Pcx�؀/l�0��WE�f�������	��s�T|#���s�D��v����;��4������By�l�&ӥ�/6���W<K�(pT|������&�����$-z*���\�zQ�]��`
/Me��:
Ԯ������X̜���V��Ǹ���o�**�Bk���y��t�ý���%U$�ܬ�o��Ѩ0m�Q��ިk����o��)D]��Wl1�.zv�L�L�U~ϵ?ښ�_��[�A|V��i���bxBX2�ʣg��ѯ�l`K�]ŹY9�䭙%j<�7�>)T��� sn~��j>�Zᱲ��x�S���z_����c��i!�|����[���ީ3���N�B�P�븯A��9�*�Fj5����-2(���M2dS?�<u��jM���'V�a��fr�>��E`�������k�P��-��e��9^�5Y�Z���0n5i#�J�����u܎a���<�0�ȇ��Z�g��$�d/����e�V]���j]al���R���Q]���\���Y��9�mA��VT���n�W�泶r�B��qbMn}�=e�y�/�6V��5>\o?A�G���� ���r����XW�^��*E�c����*'π&j6�ӭ�~x=��E�	�:����� (-D���ɸt�BN���B��ÿ'�ep^����1�����*�4[��2C��t�L���1���z���띙d1�,��/%z�ޭP93�����#0��-1?�G�������U�[��+o�^���_���`70���+9���3Guq�A���?�q�U��`�
�ٹ��7'D���/b_��k��ՐX����A�����&ߣ�������	� ��8q��Q�vd�J�KP,��5JY��,������R�ة��
WuH�����H������I˂����,�F��n�Q��V��ʞ��&��R������Ƃ7����%�����صT���iA���NіIȜ�x��_p;T܅��PV�ug�`~BU*>�Q�_�;�����0�Įy����Hb�b�2on�@g�4�2���O��X,��Yd��s��	����� C��n��诇�V���C2 柎��Z�=b])���z+���㯆N��wәLJU;y o+}-��5�4���,�Ѭ�N�� ]����e���l�VP^��5��k�OCz0=|'(�X�fBm�סU�?"6�0��h�p(D옖nM�^p�Iip\�ֶ�
.m����Z�p���A�0ԥ�3�uu�� e	�8�s/&1�L�޿�c�f1��������5�{͙�v��Ō�G�= kD�Ff�9�����*������{C�5�7��~DI��2D�dJdZ�>ʘm�w�"g��v��9�T��Ro[�&���Q���ۿ�C"�=� �=Z��(&�!��j�_�,�R���fNoZ��8���Y�� �Ia*=���#c�2N=��6�IX�c8损&�z����]t���B{��W�D #�L�Xa�n\굤�uA����7?�,�u�7��j��ޣ������.��|��-��������6�W��{>y����݃�����}�����N2��3�6�;�8�i���Če/���7�bg_p[&4��qW��S���ga�c����K��$�#P�ɥ���X�Yh�1)7�c���f�C,��b��	4r����$���X=�-`�-��dn�r��?8�^���4!�{�4'�1El�S���(��eeh*��)3��ΤuU6R��<���$�9��d�ԯm�uku ������v�F��-�z�8 ��#}\������(1X�s�ܕ?�^��DZ��P�(;NK�Hu�����K׵����n�f��@�%�kd� �ܮv� ���`	598�@�&$g�~��L|��6��e�**��pl�T
�U0���2$�ҳ�}筶��(��+H$�{���dBF-X�X/�ޑ��� c<�����A����{Q��p'�����5;o�'/4�<Kk���_��b�ø5�d��s��#�2"9C8\���>w�+9�
T�χ {N+"K^@z��T�Q~�g��vJ��{C�����'O���ژo��c�Ԓ6��TQbLr�R���YGch�w}
��s�A3!������W���?X�)"ȫ�f"�v�����a�ɚq��Ă�#�������Z8�9��p�7V%�WO;E�T8o�Y����"7Lb�+-��}I��0,�
��:^�a��` ���}���l>ϱ�11����S��t���`��z;6Kw��a���5�00֟�p��;7hөH����m�qY�,�2�	iRU�!�(=�w����p�T�5˚�YE
��ڀA�/����/�mz�& u/��rp(�?L��m�@�g*K�Q���铨[Y�:�#i�h/�K�+��0L� Ja�$��|]���Z_�8v�裈Y�k�HёL<Ϣ&h�#
7��yP֖�hi�4�R��<_l�u�Z�t���x�o;$�'��jN��ҍ���k8l ��a�Il������3q���5b��F�\1����5�01#�I6k��){��4�F)5Ϡ�_\{���/iW;�1_*D���IE�F\�<(#�.�E�O�A�DB��|�O��t��+�<;CS���&�C17�w��#qqb�~��h�ՈM�n@�Q�g|���ɹ�;b��n�w�����Q_"u��B���J��5c�I��5*Ʈ4���PecN�쇫��"����y�ߜ6 :�a��
���f���7[j6��J��R"����}��K�GD�����2��C��5� W��*F�k{���ܚD*�4����r_T.��U�q܏�<��}t���xQI�i\5VzZ�:��.�m#1(�ϊ�ɣ�^�Sg|��J;Q�
�H��E�k�H#���e��:V0�ɴͤ���,��ϔ�&�.��T��ZP#~V�B�kTs��7�=o�m�E�!'��(s�9�zj����!�J��d L�>&�$�Z������X���Ԛ�ń��� OX��U����"�@�޲K\��������/��#M�}Zm�$�{џ���Վ՜%$\'wa��{��[���b�ϯ^�Wp��0|C��Vs$k���&릐�8����Dq�,���'�A%Q"��K5�D靯0��=�1���s�x)��b$ȏ��3
���c׉�W��ga����uy���n�䄵����+|Ζ�D����v��P6X��-ҡls[Pd1Ә����!���2�>)�]���A1�5]s7�ђ��9*@�o-40x�����xI�g�����/�Ú5����-�A+��G�^��/U+I��B�(p�*�xq��� �BcD�3;���{�/T��K�����n��Xbrx
�30�c�Ѵ4w����Y��R��