��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xMMh0n��f���X�h�ʨ���H�P�e�Iܷ �>Z{�hT����r1�;iM���ٓP�d���U;Y=i�q��1��);��I�'>�8�9������6eH�۷���Y�����.������N�X��Үd�_h�<݈ޏ��EN\Th�p��P�C�>{�=۹�g�Q����4�1�VMu�K�� ��q�sM��n��C�ϝ��j����`�W�_�ʆ;E���6t�� H1�mczZ���.hyX*͠���T(��Z�7!/����6;�6��ң��P�[��N5RZ�le{�'����_5N7�IrG��o��7T}��W��Fxҙ^Lui��<(lqd/`)��<<��S�����X:s�"t$�><�$%���4 \����Y�v$:�kZ�'��}���0���]����̟0���L��Tl�6�ZD<��	��>j�@��9�\�
& 9W��t����y��A8����q��e8�n?�@��`��#L���pS
l
�k��5�wa�<��[�V�=�M���s
�!��i����]��Xnu3�@OB�;-4�8[g��?�n !��� �kHD<�=��șmp
^�W���`�3�waB=����b�h���d���;���j7�d�T�B��9�1����h���[�5;���n�&g e�QQY��K�t��~�a�a���,��bd��Lҍ{L�<�Z��W[K�f���ܧXE�U�� �"�M�!rC�G�<Y����3pl���t���ç�je���5qL�B`�a)���mKyWz��N{%��FNn�f�:����T��6W�m��$h��AvL1���0���Z�t{��sk{s��Y�l6��5~X���?S�����U��%�{Ϫ;���x�5^l�:u������e�_�k�î��Jث��7��R;AD��q􆅡:O-�e&+���΋s�c��fs�8Ѩ�A��>��{]hU~L܆&���p�}���*�o�R� H��m�籜�
6�CiV�X۞�x)G�8$6g����8�����7e����/�eW�fô�ț3G���*=E�cW�`>�p:5��?4�ͩc\䵑��_%��\�����U��f��m�t|�n���	��#��|��፤!E�%�3h��z�	���}%�[tov�v����,U�ߧ`�2c��� ����HG��/�Ge��(��L??W����y��$.�@Mv�2��<J���m��cڃЕ`�v�Û���wi`AZ�d�2��n�=�qY~��Т~&s���L����MP���B�>��+%�x��������?�}�Z�ZZe𹏪*`Cv!�\s�π>�4
i� �h���'
4���)����IY^
�������V7�'��ER�bu�E��|+09>V$Z�Ã�-���]�|�Z�v\�����iC�/E�����/Ɋe�{1�$5����5� 5�i<�A�U�a���e:(�b�N3R�`9�?-��cF�1P������<P��wD,�آ�HMٳlh�l���۶�=����^�[��O�\\���� �����b��-5�S�0 �7'�E�+zlԠq�w�1��z�r�Ƅ��	�������4������S���%;��Y#��(��L��{	���MZ]ʮ�꡹�Uk#Uv�]�mA��؛�s