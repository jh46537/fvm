��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,����t(��3�<���W_� �_t����:(͸�����*���9�%0b+Ϝ1�/�O{���u���my�~u�~�6�x���Ώ�	R�2�g���cJ A�s����d��~��{"�,Ny flW�ӚȦ�<��i+����(Kw�3�8Ի+�'�p�u7(��`�5A�% w�7��P@ۻ�j�l��_?�}�ɯ-�1	�1��|*��Û�li\*W�P��%��xҔ�0��oL��&3��Q��9�iV�ω�j��%i�s���b�qRT���
�z뾹	F`�v��B��}Q�01�,���=y���.���ەW�u��������v�3Z��:�t����i��߉�
߹f��Ss���"���[kó�-(�����$��*�Y��P���'@H*��j�<��ϒ��Y�Xõ�=��m$�Hl�l��˕�e�x謬�&`�d�@�ˊt��t�|�?&5	6����:�M�����K��L<D��^eMl��4�w�ӆB�y��L�Zwl���]o�1?E��Ms�M����P��� �>QKщ7*�<ܡ���	SO4$`$�aꮧ�QjR�D��t�B�+9U�N7�B�,e�=��r���J��c�uf2��}n��_1y���h��mR�9�-�:�s��f��bٯ���Z~4	h���-��=ϳ��_�Lh�=,�T�*z��Zc��O��3<�{G��9�=��C�O����S�Z�v�����Qa�ˀ5�E/l��>!Ba_��?|_*��B��i�֔�5�Zo��}K��4C#t$�[7�b���5"���2�-ˮ���Zu��s�J�*�qng��CM����ˏ�kd�o(pb����@����F�7�`X�x�){����BZ�G���q#��ͪ~���#
[Qx�!:�Il����ߤX�=�3"Xծ<���~J�cG���� g������qO첀�o`�G�Yew�6���.�@�pmGASO;_D������ط�WN��G�������L%��G�`cT<s�t��,GSؤL�L��G6WO���*�Z��@��b��^�
gx�M��iXBUʣ��$��I�X��(���bA�fYq��j��P�w�qI�����ҝ
M�!nl˘eP4��7߁�qRԁ5�f��E�1���}��=���A,�<�K�Dz���J	�<���K��N�e���~�dT�|�.�C�����0���?U�����@-\���V�#�L���Q�c��=='(�e"�K�(�g���O�� �`{m�x�-k�+���m$�+#�x��C��� NP��ͯݽ�a��$`d��d�BɄ�~��>�O��.l�k�Q�����G�zA�$C�/e����{��P^:gvUQ��u�����dcy��t7W�Sn�;9�!w�} DPx㲞��z�Lt��x��|4��un�n�_)��^��[�&牢�I���Ol_�,�����K\ܺ:�����	50Ά��~t'Uz�z�os��E�5J�/����w�<��(j���i���Z��`�%�[��s�z�J�ʝ!���x��i�����e��_�L�\��bHp�n���[�
����k:�,��� ��GHhE����>�-���v�k� �4֌v@�X����#�����%p��s��YG�)�Ay�91�@��k���N1���6[.dȬ:���<t�+�8�S�G��e�����_Ǐ����֍�'�M��G�F��B;��|�t����D��
T#��X�i�!p	`���8�B���2�M�7e$�� E��5��.��T��m�$�oT�ϡa�ca07�^�l$%�}�EK��1Ӡ1K�\g���V�LL���i���LF��"*��k����xc�O�>�t
$ʺ�"k��N�>� ��ҷ���qs�-���@K��6��I���z���R��:5ã�� �q����>2�K:u�Ţ�(m�(��5��.�.��',cݿ8(�?��AJ�w�,���a	�ggܩ�s+�$U�Aksa�څ^��`�1�ģ|hF,�IS�<��lя�F\I{�U�Ֆ���F
40�Z�v(,x�5vu�����f6̯2�L ��9$��%Ȇ���Y��%!ӏ#s�QXNKy>�3���D�V�&)29��5չ�� �!�Zj@�oȈ���>�=1�,P����@w�{6xj�/+e.Z�����Ibi�����1�`y:���9�k�zy���^�Vl��D�:���x�ldkR�=���B2����=�~����Q�.�)�IJ��������xh8 s��a�����=�/� `�(��#�u,.)��KTL�ZI�E��^gB�u�E��A����-U}�&z�2s3/kNG��M�K���3��b?�� />�=��A�ThD���0� �V���V��c�I�	�+�&���.����i�PE&���27l�=2	
ĄNq�{:�_�@'ε#���&P�A�V\<��n��|r����)΀��Ǘt�"����N���C�1�fɆ��s�i���M&hBD�Ƌ߯�Ln�zJ�m���-	fv)0�@�~0�a$=�Xڛ�K�S�ш�lR���u���PXv�wͰ�]���WǑ3����SaT
܇C�FHNM|;Y�
>�;��6o�Y�"������MX\�~OI�xԸ�"�p�P���R-3�h�}��?��:���e�Z�Z�u��o[�asR�M^?Ɵ'�=��|,���;0K�c_I���ӁHf�b�.�o\?�;�@3�,d�|��*Y_�T��i�Kq����\��['��1Zγ��
������|�����lN����/�8������ht���+��Đ֪��xi|R�)��N-�E=���}�B����T��%K�Ïs���-���I���4�{��j��y��~م�F�r6�|X6���%�V����2h::*��g�HX��Y�m���������"���X�������<�֩8<oD0��S��4�xEέ�G6�$����U���S���ҝEԼ$��������������|��2�4�y�M˕��I'b,���9��w�=I~��Wo�B�����R���	G��$s�1nW[� �u�JO���s�T���+�;}���4І��a`�_��T/��ź���=�D�����s��P|ۧ�`LZ����$��G�߂nGy�H���rty��+P��Lw�>��'�3a�KaC�.�j*����k
씯dkb�.���8k�٬�`X��D- ��W�&��Ncgq�j��^�C@SO���A�:�|�Vi_gČ'D���
�p�Ҟ!R��(��+��M$����d���