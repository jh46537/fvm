��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�k���W!�`�����lgX�5U� �!:ŗ�	R+�Iq��lYI���J�_��+�\��� |^���c��K���� ��ݧ�9G���=��*��\-n����Zҹ���3��Z�2U���ױ��U'��G��ľ%���&��D�gB�ɇ)���sH�V��.��a�qtޭ��U���-�8�]�R�������z7�p�m�xS����t��4�	����oŕT�f9p̱(��y"��%4�xf��ΰ(u"'׈o�B��H�\���Rk������bQ��ɤ9#Btjت{�uh}t�����F�CSr����~���b���oT��LG�AwuU��2��a�ߐI:�? q��)2�MF��J(eZb`M5�Ҹ =zC�9��Df�0���ZfT��<p*S����<ZJm��孤Aጢ��p����f��8�����
fd����eC
�	L:s��!"vy��.Y�mG�42��u����T�H?�`DQ��pbS��T,��&�=
��%��uqat�h����.���ck�\睞c�SF�輑69a=��B�*Xg4�������8����4�;��̋�Զ�(_�� c �f�ll>X�X4�v�f��
���r:>1 'b+�AKh���E�����]���&���E;<�uPS�4����@�~*���c)�6`���W��3���b7�v��*N)����������c��? ���||j���k'�<��
G<�0^�Իs�9O+>� ��_���Cڊ�\?��u+�i�`����z����5�Xu��k*ᷙ�D�F�+O6����I�ΫIEr��Pq1}(v�2���]��=m�@n�c����#���-��u_
u��i�d���#�����wv��BGK9���{1�H�Ü^���_��^P�E4��FڋH{hZbRs��(�jpi�Jѭ�K��Ma� {)D2���K��.����dk�9�
�]lpp1.E8n�d
��{?�c�����Qr�	�ςyI��&T�Հ^�P@�����a�44�?l;i�Z2�k���&�B�6�ΞXkMz��[�O��2;tZ�@<��O��̩��E�J�h-��Q�}W|�]&�V�O&AaЍ)��ۆ�@k�@��#B��͈nǨ��줿de\��
W� z,�T�/��m�'`�_����[�4���垼�|�Zf^��6���G���馹~��f�v�6��@�#k���N~��]�����
�:q����������e�/j�K��\ӓe��:�#-���*�jq.|G�N����#Ԃ~�<��j�����	��sz�Rg��G-�z��ģ�0�v
���©����7ء���wM�^����m%�z�X�f�jz*$�k�C@��[ҏ��{����Z�2�c����B*[/O}�w2�����p(�?%_=�ţ9�8��Os���2��#kt�9fh�v.1��FvŹ�^6�=w�,������������Б��~&��,��k��ֿ������D��V�H�Jx>
�ʊ�=?�ɛ�p���d�N).(��/SW�W#ZT�R^ZV�#��gMfIT ���G�H>�։��Q�Uk�O��@��Bߎ�d�v9��:�� �x�2�>�2dq]�+œ��SK�D�"PtBrH�;/�����U�І�+��"��- �Hk٣�ּ;�O��R�܌`_�Ol�Z���
�[���5\�Q�q>��ާ��&Q%�x��N$d��B҄z��w���H��H�ulX��$�D��`���v=y���X�����Z�����qp"w[߇����	GX�%(�Zɐ�@EP� l���AY������^����2HE.����{�sKV[Lk3��� �WO��>�b����-l��Y#��3�&�|�����ܧ��s�|�����gbO0�Th:G�1O�AN�R�Ү�u��9&HEC���-^����p��7��Y��y�*g��b�%%�����;���@���-��j!�%o/�ܸB\-�s�k�ϔ9�q�9?�.3=3 U�͛BK)Ӹ�x ��Z�Ay�LbE�/��y��g�[z@��,�
�֩���%Cf��%�Řh��05����	�n�:���D
�v��8��D��ĕ��Tgm�]/QE�_����TXу<9kp}�v�%<Ӹ�mdh���.Eԡ���Oh��V�&.0WZ�o�l������!x�T��] j��Wې��*`v+1�/JCGtMG�A-�紘���b�[(�@�ث�2���Ť����h�2�%O^d�6H��ͷ=n��f�p���Q܍8æ׍��G=5��dc�U�@{p���3��y�S|f5�N�*�Q�І�u�v��t���ϾY�$��Ǿ>��=�'�������N�Wn�K��O�c��4�)ǡ���%.@�s['z6�w��S�x|�r;�v��4�{^��a)�����HVu	x��G8Ѧl�50�)��A>l�k�Y햫���[M"J��f�23+���k�6U��