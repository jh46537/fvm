��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>����p�0�F���)�ã~d�:����f=�n����l�@>O�Њ�۸"�#~����f����S��UT���������בJ���\/��2����r�X����`Ir�K_�x6YV����(�/�~�k�q}����;)���3~�=�FgBBKO.��}�@��z���̥x�6;���X<�����~2�M�2��$)�sFaa��4����9Q@���e:TWrt���z6c)�<�~q\M6�'����/ q	-��# � � ?!3�m���{�D@� �+P>�e�<>��]zF0�P}��N�в\� �Jy�Ǚ�j�qAw�IX�Q�2�6�o7�O�7w<S��H���y7
W��w�Ӯ�T��Qg�"D��^�U�L��u~I=�5U�$��n5p�V����B�E"i��z�MPBo�,{�օ9����Ka��s\�^�d�hw��*��V8l�!��KSG��O͹��=��_^	��5��|����	g��R�I,3��q�,2��bA@
�C�)�*݆f��,SY��_t�F�}��u��eD0��U���b��C��F���n�a�5��������h|	bM��d����h�t<=�%�kJ�M�B<��᝶��=�N�)$��o��eZ���ڭ�'g�-�A�m,b/��.��,������ꝳ��n*����#8�B������1��~m���Pgj��-0L�6�ks >��~_�Kg�:�s݉�cs<��=��1�Z��Ry�2��Fs����MdIi`,(Bn��d�z�w�SKZ���M�{� s�$�=��^kaP2�Cu��a��%�� r Cǀʎ�	ǹI�y�07��$��G�>�N�R� {�Kvՙڋ���r��I�z��眄I��JJ)B�v�7��~&	�q!�
k�!���k*��ZA܀�L���H�^�ωk<�Y�	��$k� ���^8�R%�#�J������A�>��s�đz@;9L�X�4j��p���/�:����T�����;�'�F|� 5�{��]G�a��[A��Z?j��Uΰ��fp���'�b؛�ۿd�W+��i����}�������5��c	s�Lo �� R�|�������yZ�&>��rK/�eN��U ��'᫷㙙��Gm/C�z5q��+/>�=�0 ~�w��a���ڋh��p���B�;ń���g{�2Y*`ǮԾI58���7�CCnR�g©���$���bM�K����K��
�r~��"B��Z��2K*����A���9�[�Z��c,�2�)��7�E�v��yR��ϨWc+��X �hȫ�76w� g�6F9������MsH�N��f4�3ʘچ�4���� ��1My���#�A ��ʄ��~+�ް�$���] ȩ�R��ʪܑ�uO혔_vd�-�c�K]M��A�v��v����������
���X��YE��K��s���3t�շAX?ƢK�R�� y��^�}I'Bu���w)Rf ��������0�1��`_�u�i3�''��NA��%Yˑ.zl& *p�#�RW�邞~�����²X6KPU��SV�٦�ʀ��f�	f��F�z4U����W"egA�
���"r~"!���x�����UUe��Y+�3vǿ�0�2�P�@�b�]�a}���2�ˋiX�����&��k����A�"������̹��'�nK�^�a�z�^�(����e�����i������H�~�A�w�f��_���2.�	Z������9���V��/�{�J�}�
/��\fC�� XZ��J�c�_���ۚɏ�|m,��+��»a�q�u�i��
�Ǚ��������I��6����Q��z�%�-V�!V��?\����[1w���Ի;�]��C��l�^����ޯ¡���a���Z��ոBM$L%lf�յ0u�<*��LN!�����%�'����o禑�M z�e�w} �
�$fl����!8�B/�����K�p�8��A��KU¡�~����U{��pY.SC�3��p��}�����~����U�N=X祱�M� C[WtM�/J�í뇙��K��N�Fë�K:.�#��eOif��)Nj�A$�=�=BMq�dq��߿N�.��גc�/�1W���/5}q��p��^�7]��z%�K�"Y�F��#�a�JLn��NJx[H�am)���r}�(9:���wjcؒ�м���V%��(&Y�ܝ�) ?�tz;ցE#¢���K,�$=�������&n-e=�;T���f\O}����e{�yi�ћ1�&�sQ�,����Cp�R|��Jm���[K9���$��^C�9�ӧ��)׌�8��v�ik��qR��/M%����w�!�-༮9g�^.��{:����ʒ�B��D�[�4��2�\�h9T��2���r�Yk�z���4�j�Nҗ�n����d2��@�>�=?�)�Q��qEFe��^/)�pq���ÀE"j�z�����L��&�s]뚴����1��*�V���Q���|)~�8����-z�*V�eC#tTL�y�Х{]x8=\}�U�۩����/[A]��]��b���g[�B󖡚j0$�
˭j0=K��4��vA�r�I�����
@D�	���;���f%^�<)GO.C�h�G@f�7GJ�[i��J��r��t�Q������"�������X���X�L�Y3~�o�+�E3׷���v���$
�O����E#.��B~�bX��޴��	]�����47pً����7��XE���[��>�ZG��b[�7)?�ތTΡ:1�!6��2.]�Xl��'�dXpy~���n[�^��3@��ܚ�r����#��a���:��Sa�D����4��хn�����4�f7��%�DXt��K���/H�Nm�*zܮN��v9���D|�B`�N��)�[�o����T;}��@Y�t�Y>�FN.Yg��"�S�	'���"���A-~f�A�t��Y�4�l��wb�]���#a
]:�Tɨ�����M�·Y�%�1y���bX��ξ����Y'~��A����L�YN�w��a�v� h��`p�L����@^7�-�S�9W{td?��
��W�b���~���(J�/�K�ƱgP$5��d��Z���'�g�vvǰ��bN�˃��W��w��#-ne&U���ͅm����k툍ezX�ߕ^�^�sQyH=jA��Z���;?���@9|"�NA�	�>��G�sA�b�]6e{x��Q
�$s_�R�̨�7�-6�Ahl�"Q��S;�.�u׽|��c�B��,�g�t� VR�.h���0�[�����s��_��OA7���J�A��9��c5v���S�ׁ�x��y�#9a�SH^�6`�x���g�jx�K̙��S.Ȣb{{�A�$��id,�.�#㐑�p2���2
v��vb�~��i��KW3�<3Lw�j^8���Iy;&��ʜ�s?$�޷��N�h�7�G�A�x��:�%���5�I|J��>oѥt�� �lrm��ئi{�/�BQ3���d��i�����$3�Ж�򴶐_۞���D"����3� �J���{�V#U��GX`��kk鼚��4+���J{�Ձ�񭱵{ܸrJ\O�\n'����S#ɵv��s��t��JBX�u7-ަ�Lk�+S��]�cMx��[r��x�XX�Bcƶ5�Vy�h�애1S��+e����Y���ޜ�6%4����b��q�e
2�[Z���\J�P��������F���+D4@ܖ��F�V���b�W��z�7���2�MVYP_p?P��$�v�����[b{�3���]���yFSN�E��*��I)ih���]�&�,�d��%��~��E ���������s����Μ%���9���G�2&��CA���j��$�Q�J�_����!+�#3�����U�@R���s5�4k6��C�@��Ϯ����7Uo3�f�YK}'���*����
���*&Tӛ�;��1�I�n�R�0.2��N��ť-���i�%y�������d��0F�&���ÎJa�.��㭣���/����+4��+p��h2��\��I-�((���~�#Z�DUU6rV��h�|GV�e�>N�-�c=�� ��T�+�W�9�	�\-l�5Ca���|vu��E�/jR�J �j�q�ÆڲSs��Jw��@?���́l�.@a��\!OD�L&�2��O�A!)\�:�� !Vi�W�lK\�]!���E�ዌ��%�pymZW�B���~�)�?�����^c}~p�X	�CW8�ю`t%�i��j|�i��*����!�
�\?��'��"�e"=z��%��V_����.���������u7���t��^t�8�*�_:~�T��ks��7���aF��	�(�d��$6��>es�9�X�B�U�M�w �C�
c��SC��[�!�᎚YH�r�%�t�mw�#(�\�`=��U�Gҕ$�y�9u]�<�������Bh3�o�nMǓ��J��H���v��$����u�+����&�n���^�R��]3P��}���#��_Pz��z�f�3ߤD��W���q�֢�=���K�y&T�6���Yx'�P��^G�9���H#^�A:�!��'-ք�V���~�\�ʜY�g�(�@�uΏc����`vd��DRT>�R�S=�d{���)���)>�d�63U��U�,���h���4��!dG���bӾĭ(9�ȿ���sڜ�y�Ų �ђ��F,��0YPٴ���kA���R�[Yn ��Z�L��f>�GYώ�#���Qw1	�
)�������~�({$���L��@r�[8v/c{!�w��\L��A�]��ou��7��;��S��GbT��	�TǍ��΃#���G-�˟R4��G�ÈЂ9�_V(8��'(K��t+ P�R,�E/A�pf\�~9.'4�J�,��~�el����y�[hU�j\A��G��%�B/��l�sW��lb������%[��K��6#~��	�aa=�.��1�jo�mI�P�t����;�[����~']?G�[@S��
)1�z7	~��^e��	�i�]�uq]iGf{�7wr�ʪ���?��9��'���f�bl�6-����>��|��Ja���o�	bε�hG�P��͢����H�0r|>��Rxu�����܀���Л�9Z��f�q@I�ZP�c�T됱8���$�b0����|�|�"�9�R��g�7�|P��G@�X�k�ى�2�V�RRl�\�7-�	��@���<��Ԇk��*6~��q��+����#�
��N%P�����g���xnoN'�b�G8o��B6z�����0���e<�U��U�9R:��W�U�U�b���K�1N�+��w{A��쀿�GRs��Y}�kd @-ȷo�2��tՠi�}q9��G_�-*ߤ��H�5�Q���(�|��M|��7�5��z�03�ب9?�Z�<�dd��[���l�5��}�^��;��DZ�W)T��C�r�?6&\W��7�l��&fu�`����e�(�c��Z{��PSC�E|9j>�8Q��2/�"GvuŅ,��G�σ �AF(���K��IB�q���X�z�uEd��S��*PU[�x�1WRQv����c��t�pB�I*�eHa�"�i|�'��ir�����n��KF��K�����ʆa��eB	 m�]| o��S�{���k��G�*]�V�1�ed�?w,���M�j{I��;��z_�DF�K�7�(�a�J!�)Y�wePD ��v1�����0�r.��}d5��K$���P���S�O�@b������*�sC�7��2Fɒ��xRz��m�'
��m[C��_];����6��8�b;K۴��XM�؆����hC�c�(���dJ�4ڐ��!\����/��&N�"Sc�n�+�[Ya����~*���2I�'��l���,�0��<��I㭬����S%O�r��Aݹ z�:~-bh�����{�`�le �AȻ1�U��϶�|��wB�n�Q.}ח4��0�Cѭ^��6��FU�%��J\�_#�vdg���2�;�7~��ES!����R?i]=�W_}�����=�m�%�<�OR�b�+Sf}�>�ƃG��Vw*�D=̿�J�O�c��T{��疎Ou�ˣ��y��h}TrHHb��Ɓ]	V�������������nΎ���R��bϽ6��������w��r��f���m���&�I����0��tż�{@��� �/�,��S!�G?nJ[<��D��ɚ�A��q�J�-	*stγ�͋M������yB���(6��S����jF8g�K%�~��Z�$] b덾崪�	d�f��C�ޗ�_���(� �D��o��/Cݴs�>]k�o�g��/�~�X�#P��	�NL��َ�h�V3κ�VDC{���Ao!���!���a�59e?MK<��WK��f�Ǧ�/>�����w�ilh����M�7\����(=��r�b� \k�磦�����G���4,t �g�y(�=Z�^�B�F��"��Zi�)���*��p@�3L���`{
\�S��ߕ ���S5jɪW��]��`����"�ۅ9R���]�v�a��^��f������ΚWt/�D�lH�-�")��ƥ��UB3+-#}���ִ�J��E1���3��v��4�ϕ��I,�������Zh&E|0J��ܖ�_J�&̻/��ܫLG����L��a��=AK9���-��N��S�R��Pe6�B.x�w����V�_s���Gz�E8b`�"���N��~lϫV��
�z:/ ���l����B���C�w1�*D�>(Ĺ�|QZ�j࣌�ą��a{��OR'�VCӤ7��ۺY:�5�s\4t��+iQvv�W�y�k��t���h��V��%JD�q�2'�ɤ$)~^ط�����&K&"�Ş_��{��0d8�E�O�;q=�9�/�Y��%�`�Bj2�����t��
p}�����or�E�Y@�L�f�v^�{*̄,���[m=���R����$'����> }܇��BHs�}���Wt�5�8 �9/z4�?�)V��jb�����:s`]x�U�ΜM�kEL���7��������?�#ֻs�.q17Mm9R_	����7��c'�#$�3>���IN>?1'�㍱n���8�/��Т�+ � �6^�}=��J2èr*p��挖��2�͂J�v����Cd����-Y9b��Cc����	5s�����G��;��� �3�^�� �M��@3�",eD	��ិR���A�eAJ�JSM�dQ~ಹ{�&y�;���'�a�^����"[�X�&s��G���_U�f�-�-�q�����"O������� �|:����N����P�}�|���X?�1�d� h�#Z~b;�����%$��G�B�;u*A�� 49z��l��
��*�͐ac���W�L�Ґ)��@+��O�bn՟�r�wZ��l�p�6�D��heܘ0�o�θ�7�����l{�1���?r��1�\��a`%,�@ϸ����T�'�aǞ�}������n��М�a��u2[���I(���1g��`��Db��ל�ma 	uzT;˷�dc��k��܏]���CY�@R}�=��,S�{,�	&灧�[�����1��u����j�g��ч��cu����P�ߵ��G���PO�#QjH+�2HW>,f��pE�%�=ׁEr�T����n��Be'<h��ѡ���[�)F�s]VBg^-�h���Y�W��"��W��2�Z������oiaS������]�?�#�J\7#�ڕ�I�8n�KX�?���y ��9�q�U�|�?>���?�t�:�MI���f���.*A���ga7�i[k\�x�:�A�I g)�-�(枛�p+�j�!ʦ"�L;�9��=\	1Iq8�'�E-8��Ϻh���_���m�l�|I)�0�n�զ�ĝ���Sb���3lzh	�T�2֋�va��E��g��}�34�c�� ����� y���;R X�N��Y0ޔ���)���ʢ�'�x�/�{P��+��\�A�@�6�J������|�U���*�˹��)󗯦�"�����{U���*�b���[���%���j��_�� O��I�1X�ܣ�׌��]�Q���j��]���E�RV��8���C�wYK������-�������X���v?�À#s��R1ۤJb�%���9{��VX�Nͭ�Y|�6v2���R�yni�I^៭%6DBG���M�gi��߉��u!O;�%	�.�i`)���TL�6Q��ޑ3z���D�nC�Hݮ�"a�@�� u��/O�X�e'��o�Tc��/˖oP�2���4.�����ܱ�1Hk�2�p��6Q����G��>#����1|����b��L;dbT��*A�t�p:�ų�;��A���ژ�!�dg���[u���^	x�&LYt��v�`��L$ĸX���#_E�����KD�=lDh}۵�rBoy�������a��1�%@�c��/v�膝�t0W��Z
S��$�%�qU�N���T��1l,�i9F6�+Y�|��ZT0����?� mp�G��ƛ	��s6!_�K]�u���aXsힷ����,�1\����8��[մG	/�ۗ�G����S>h���)}[�� ��V�1�C�7!Fy�J��S��b�G�D��)���72�Kk�6��~��-?	}JRmg��y+�̕�ƀ�|?I+�^h�B��񠊫���s����sk#�W8X�0䜜�΅���o�j�d�hSQ$�@�$�S� t�U?M��|����������%��
�����.e01�§U;8�Nɽ��?BI���'�&_�m�����q�5�?��n���^�vP��������^!�Z���?Ի�AK�:sWfT��4���K�ui����
�%W�>>$�A��*���`δ��p�������r۵fZe�*���Wήk��2�,�018�	��N�D�"J)�Iͭ9��;��)"9������J��P;�5���w�Z�lj�_\�a�Ă����C�?��v{-��Q��<&YM���F��\�CX`��z�.�ը*\��gx�+]Q_d�sN,Br��Qfi���I��pٙ�q��nW�M��d�?��I:#:K�b�1��e���ê<�+|1�h��I��� >}��@*m�[n^�p��� ��`�Ф��g��x�Ɵق�2��>�e�x��KX������bU����K)
�60��J�X�,��a��9N7�kdڢ��ǭ���I��/��[$)��)8�<�S���8Tp)K���/���*��3a�6�`�^@g�ZIM�'88�-�{A���3I� ��a��b1�RDƤ� ?E,xg��{�ZK�1��PG�T��A��^�j��D����?���FW6�� �Pk�S<�o��<[��tv	JQ�5t'���&�ϭ������T�ŧE�=7 �h#��X	�1�8ݞl�m�]M�f|�h������'���'�7�l|Y���-��u]	a�؆D��Vc���'y'��N����(�8#oI.�$������6��E@����{y�u�?Rb�CBM�����:C���U������Eϋ�%�0���>��W���1Q�(�q���۞_�-ŏ"ݫ3%*6�b�@�Gw[G�R<��(BN#��6���pEj��|A�.N�9�C�r�^�3Cq��uh>���+R4%1����?UA���3�u���sam��*o�� ��_��lè�˥-�r�k1��׌y���:g8���/�ȍ�i�zS��u�`o�Q�-�<��H�N��z?��p!$�^��d�@�R�[T�p,���J��*��Ms��M:=�����O����,h�8>�[���%	�� /6V��n]x�Z�mֺ��J�+��YMާ���,��1�t���s<p�yam���ff�x$y0�;]cSE'�N�l��0O�\�ߘ{�`5 !��mf+=�����?}�]�o�EO�f�����)}¶��q�)�P���Oͷ��?$s�� �R��6��1�y��=�qr�	��[�1k��'G�v 9����~�W��cY�$}t\4x+�T���f=z�%�����Ss�2��0M���'��d�N������,�X�^��X>�"�Q������64�����Zr�����Z\�߲������G�SˢRX�$�QUG���W#��������׸�87l�`��;�x!%`�I)�}���n��Y.Æ���mJ|����u�X�7�j�ُ��8�yřtw���T��}:P���K �-t|���uƢO��
�b�0+k�l�=�h�����A__|��A��H�1n��2����{H8E����I�8ن�?���%�����'I=�������m��\=s�K=���ƛ�`�1�z�-��"N��T�	 ^��Mє��گ]�|�����0N�0��}������o�΄>A��FW�-~���M+�����q-×�bvE=\�P�������,Gͻ�P�ϦD�� Ə��޳g9o�o�:��̪��������:S�TŻ>�r��T,�����S���}�ܞ����vQ�{@ذ�{b�r@�.�6o�.�0��^�/���F���Bid"���I��jݚh%Y�^���MB� �oS#8ӭ(�M�-����Z�)�Z��Z-���N�9d!�WTΉe�WwJ�o�YD���=��vv�<2y�o�F4��H ���p�Q�s�K����M����V{�R���$�1�E�Zp���f:}���� ��[ŭ����ջP��Z)��m���骿��ݷ��cŕ��ß
D��<��5�{�Y6��Y�b^Lt��)H�:�7l x�2�䋰1dyG�2�?����̵��H�r���1\�3�x�k�K���hEE�34 }��6a]\��9ٚHU�(���Q��\�2�e�L�>!��Aˋ�Y�e���#���Р.����堶S꒷D��}����a7���9�UW=�Ӑ���:͜/��.��t	�FNN�*g-�y�p�d���<�Њx�=���f#	��<o
8���wz$��x��^}����˘&��DT*Ȑ�ܿd)sBp��W�"&E�W�ьhŤ�x�Wm~�
]�}u-&�\���������_\cS���Ia_8�!�����J��Y�3@SS��?|���I�E�6݆��H�zР*����4�|Ġ���DY���*4�⊛g �7���PwNÉ�=ևtؑ_<p��JL�M월�9K���"	��Ԉ����$���j�㘘�WV��,	� ��s�)'���:=�����5ъ8��x%��At�r�N�f����?єA��д���џc ��VD�%v�1ܡ����C��I���h	L#�O?{:�T�,/�]�9|�Sl9��E�-���|"nnk��]��(�z6# P��]D"%<8��qn<$MX���!���
�Ƞ�D�5�ܢ�����{�拣� �q�M��qbUW6T���� ��iF.�?P�{�o�$q+�������:�k"��I�eh$�C�%Ӏ�W�+�sw����ӑ������jU$*cn���j6Doe��ǜXi�f�pӟ�!��Ϩ[h�1��Ԡ��\5Mi:�(T�H�7�'�R��;�cb�xZ�ލ3Q%�)��a_ /�I��1�9|/�A�1�H��������:��	A�۱�>�^��0��Dg)c.���Ae�$��|�dj�������tM���/g[2�r����G��eɛ�O�G�G�B;�}����`�|��Ye����r�	Xh��{	u�~�ȟ�<��}P�"��P��9����L�ht�y˨��U�*l{�7|��D�Bpl�Z^Zw�_��FC��*t�s󃈅����~@#�h�����֬.���\����z��;��
!����}^��^s[�ϑ2"��s��F����R�h�Y�n�^�&%��� ��%����p��<�t��F�#W��L�]�.�U������ �k�(�WnE�`��R���6_�'s'4�=��g������ۇ�����L\tj@����4
�EBYI���>2M�h(�	$���sL����x����;9]FY��/��|?22���+�&ؽA@��r�û��qj:�i�즷�R�A�]���l-Dd{l�=��]�jb"3�̵�4B`HL� �����׿�{�V��{I��O�j�g����PW���Tg}hq��" ���i��$�5�pp0��e,ko����%�M��ī8~�s��4������H�z'6R�K��v"�~���wg���9~k8���$��=~>lF��Dy��Y���]�$l� ]���K����vɭ��g����:�[�j�նrȧ�d�����$�v�ɏΑ���J�x@Y��x�*�S�Y&�4N��BYf��a\��I�qvh0��i� $���"ʈ[�
Wc1-Mi�✾G;`}ފ�R�d��*Vz>�� �R���W�U�C::է'�[w�`t�����[@�#um���Y��M�"�ZBĻ�&9��h��(lD�@�%�{��"I�rJ�������ʒ���1R�"�rE����}�0�L�FGd*��.�����:�U�(���R!&S��pj��+3��譭��L��.�t7P�����N���c3y� kg�t�י%�g+G����1���M�N�ݍ p�
���'���e�ܺ$'�ҟ���~�=3	�?"*���Oo�S��=�muS[1x!��W9���+pf��q�.
�����0�5�>��Z�5vʅ��>o����c��y�����ZBd瘰�QN��14�)�"�BO��
wW�9Ķ���BX,��_��jm����8��'��*l�ړ8$e�ο�O��v���n#}ac� ���Uu�%r�f8�VXF�U��(b�V���{���o(�eg%zw��i��9������2�'�}�XQ��N���d6�K�����ә�5�����O7�½i�[R��sh�+.U��t��i��k����ή�HX[�������[�ؚ�N$ 9'�H�����~�R���\�_���L�gӐ�e���\癛�	�,��x� ��Ƽ��O�i��y�S4��v5�x�wF�1W���m�^��u[���dݚ�BXn>�*هa�s����V�.�@<�����vs�s~���(��E��b��
H����L�"����Nt�� D[�m�� 4��	B<����s�����Z���y�1��\�!^ؖCJ��%�������!�b�:C�����}�v��N��o��D��	3��8�b����E�e*2�������2��!��@�h�Hƴ�����e��*}ug8�ߖ_�ۗe�G� 
����`��6�X�(}� �
5B�!�HX��-��4��mE���ء$IG�2A\ՠTl�sJ�"�a{Yg
z�v�����i���(�NQ��j������A,~���0)�n��9�,+�-Z�������+�#䶻��a��Db�6Vw���]8�u��������C��n��}O��ri)���U���~�v�Xrj�cg�cj]������37k����M�����@�s�˛&
���݈~��q�^�á�B�������[��9\� tt�#��$�Y�nsa"���j�{���o��ޅ�p=��Cڛ��b�-Y䘲g�����g;��B�M��*�cJyP�9�2������5����I����Dtuv�No,� \� BR]��N�њ*�޷��=Ժ~��ᨄM��_#�L`�K�~���o�Q�wҒG���R���H�v����������B0����v{��e3�Q�ι6f�q�����P4I�r=6�M�$%��^����Z�>=GTNp�vs/]�T�����I��/*f�ԋ<�u�S}�\d&�3O&�"nN����]��X�{�+jt���Ƈe}0��f�i�
.���DV�Ub��Z��/M*�*�LR�@�E��00���G	^_�fx��4��~�D�|P��Kx��,�7\w_o��i������L=�9�>�p%s��m@W�][?K�K�3�S_��J�aօ�ÇG� $�d��B�҃�)�E,�I�����iJ@�� �H���Og)���ׇ��ՠ��IW�;:������2�T�v���Nx� D�� ��[��ت]"�F��([Hr�FO�l�WlLަD����1r{9"$�E������t���\]d��M�Mmp�=I��@�0�F��ZU*w�>/U6@d3�My�3<3�B�xhU�i����m�2��ޚ�
���'q2������L��C.DO��
]�����x%؃�͒Fa�*vK%H��!����g���ߝ�4�l2�]>�ygU�g�G0�+��h{r�x٦�f�9FE��=l��dUoi��]!%����ʅ�f�GC0�|3^6�!��
��Q����%gѮ��>9�ny��=:�,@ZxߜO�a�JP?T;&�۠�.���v3b�Ny�7�-�+.T��>G}Z�Qm#.d�ާk�4@o��(�f3�������
'���>m�d�}/�����:��/~\޹f؀��n��6��?�����F��+���C����֌,��{�vM�WhZ��m3UA�t��oFN:Z�ݨ�t��@z��^�JBG
��3�2(�B�F=���j��A������G;Œ͓�b���۫z��%��=0���bܗ`�ZE�����H�#��I
��ļ��I=b����ŽbA��:�=A<R>����w��,� �jf �2�X
�ꎪtM(kU�^
��Z�K#�dĴtڌ*�J�,[�0���ذ���5�px�>����c.�Z_��Ѯ�V��|yO���0 ۦ:f�R\�Rk����?��`�/�0�1�/��n�_��`���H���X��4\����p�i�u*X!m�1@F)I���K�ۨ��=pj�pR:,�t��프@�{Mv1�Rm-c��'3"��a�I�k&���V�8S 1E��ܮ��:}D���zh��ޙH������\�����<�X�(/��A�6w�Sޥ�s��7qb�Ũw�Q5��V�*9~�M��+.y�CgA
c��mMcë������b C}
������J����N}���$�V+�� ��$+��!�h�8	��V�+��������M�il�ف9Oz	d�1a����A��n�P����LчŁR��\�� .��?��<��z��
�y�~cE��t9���1m�r]����q�(j~��aDWK������oQ�
z��{�/8���p���W}>��L+0G�������0��J�+��2��t�1��g֮�.��`,;�S�f�my�ʾ)��~틨��������΀��p|��3��C?2�r;�9p"%4�a���^���!�ߢ��Il�������F��:��8aܑa�0*�����ܮPKr��%"�O_�yH[��4ڍ�Ȟ�c9N�rq<��JkL���{��\����
�|*L)Z����kp����Z�7w��g�J?<�i�gNJ�p�yZ�S���A���4x77fj�CV]��5t������1�%����I���Lh�Pu�"�C]Ӏ��'g��zq��E[}dΖ�+��?���� G�]eP�w.F�?10$U�[@�[5ޖFb�s������#����	!�V�B��J�����
v���ϰ-p�r{Fi���n
�Y�������bܝZ�x��$T?Cr�:A�K
	Q��ڭL)04�FR�GO<��ĩ��+ `���B�rv�Ϟ��ߕ^c(ȾS�����7ϤZg�j��iT%��kq�n�����P���D�?���i%fǔa��(n��lL�n�5�mc���~I�����)�st�ڠkih�}�-���}��竃���+�Rp��^���"1����̬b*OYvӛ{�%��,����ף����L��UΒ�6��nKu���?����ٶ�/�U�߹�5����ώ[[;2}B	���}�i����E�],@NT�A`t��4)����LT�V��Tut�ar�hkΎ\U'�KVGn5@Ӌw�Ї��\8���}�+�Q�')_?E(���x��'�}+E���|
8�|�U�x��od8��]�i���qeM)[�vw��6�k�f}��o�>w��7!�	o���-J�/EyPbt�>��e����]�fb���^�κ{S%e��UgD������ �$�=W����"��`���'��0��U�^���u�8K���k�h.��h�Y�6V���A�
�cbH�K�VZ����x cP��^�V��oW�W�[f���f��5!K&ĺ�s�_}��T�P-�!T�*#�`SY��Y���t�q^�q���c&5�}�#K������8��xPCʟ�}*�W(�I�v:�8C	W{34��)�����$�G)�����`���6������Iu�ռ�>>(��H���x�����c<� �_(i߀��
3-Ę}�@!΀J��,�j~
�r��Ad�iY��:0t�jn��%�D#\��5���o�v����h+]�]R�E� HiT�����է��5>���y!<oŭ��}=����/�V���mR�9d�ǁWz4�E<k��z��ت	+��*�Yh:�Dａ�t(��S�Y��/�y���AJ���Ʋ"Ѐ���SAq}޿F.��J�O���ġ!�u=C &_�МF2=��~��>&���:���Y:l����-�˔��K.��sQ�}��_N�uK���mTQ>S�8Y1��;��u��Z]c
��$��+��8��#�yG��U6�@�p�n;�Ws��������^f.�AR��9z�!i0e[��jhm��
BD��ݡ�'��Cƣ�N��X�ǜ��:�*�ح�v8������lD��y�����_�P��6��fg�0��1��@�n{
��O@Ϯi���E�(�Ti��h9j*�<��
��t^�X�a9:Oo#uy�5R������k������F��8���ժ����#�'@��.
]��{fA��<	���~�2��}��|��f^����0�9�̵���-e�_[ē�O�`�����v���>�X��&�ĩ	�Y;%���ib�o�mF$;�ˎT.�1+������@�6h�N�7bV����LA��Og����"]���{����$�z尽 IJ?{c�t��p�m��{�M��$����g��|��~Q|����ir��#�1������� �
�ʞF�6�Ň�"��'��1��*t)cU
�ӺL�fM���W"�-�5�!om�R\M���~;0����F�q�'E��Qx��24dˮ��՗��ѝ��ۦ��c�~�6h_�|���N#l�}�\A�M��m�1������9.�Y�M�ߓsx�҃'�װ����(ဪ�[�M�kx��m��^ොOvpС�!7�産��0H�$������nO��u��ѴOt�����J���f�b�ǁ��~e3���!�!�9��]��:�a��(��Jo�P��7RI���68��?��T���T�`5�.��?�H���J�I��M�+���D�	���*���<E���;�T嚐t������2J�,|rOw�8<��={N-������ЎD�iq��a��*�ۗ���%ha���`������夾�[P{ /7�Ťma	�E�0��_�E,0$	ET"C��r5�b�FX��3Y,1����?��Ţ:�GO����|R]j��,�+ �����8��>_�?�p�FX(���1ྲs/�HE�ixm#��$�T73����c�����_B�Vx���p�ر��b7:�0}�7�2��֗Q�c^�
 L)3�I�����'Wp���_��X�,騮J�ғ&�7_��R>f����rZ�����bG+���~�)�*��_0�Aw��9�Gm����e����|1��=�&��dX+I)�gs��^)i��H(P�Lp_�c������G����P>qbm��zlwy#�]�&%��OW~�Ҕ�a�YRoܲ� b�
 \V�7���f�~���G���ւ�� �+z�cT�@�S�b�7�������|=.׼8��^���8*�\w�*�ƶ|������wߙ��..8*6�X���1Y8���z!��[�v�O�t2���Eu&���Sz�BM�� ��?~��9U�5.���9��G:������g�Dq��8�Pl�I�^�L�ք����Z�?/\!<#Ŀ�H�a��+e�LD�F�i$��xL8#q��+��DC!7�%�4g�����}QdX���utN�ԭ�lq�q�ޅx*1(� �9�
O��Ef�S�sZKnn�I����/�}?��A�����G�T�&��K�0���'��s�O�e���*Zr�+d����������m�Q���C$���}�X�7m�/f5��Ԭ0UA>�ؿ��65�oLr+�C�g˦W�D�M�����3}Q�=ՔQ�����Mt�J�s��@�f^j�0��w���#t�d�;��S��7�KS��\�������n��4p(�0X�d?���w/�.�����-h�H��,�L��[��P�h!����(0�u�c۱�ub���E?���F+��
�-#b�+�'���h���<��Պfd�ȟ辍�T{J�{"E���Z4:�_��{�蟫�GI%�ȡK_�����XH���1j{@24RJ�b��Q}�׉"�$��$2B�7j�c�h(�0��J��s����� [�j&�w6Ș�3H�;�5x���+��N�F��]��B��� �I8�N��8��]A��i�����P�efGlr)�6+�vAb����^�=��9�'�7�B�1lٛ��#ީ��X��j���Q�������̳�mS&+D2�(s�Lԥcd&sRN� 1��\}�zE)L�X(!r38,ha���]��$��(���3��pѰ��B̏2�Z��.�7[�$y��Ó���f�����=�rk�=�<E���o�h��t�Mh῟g)YV0k��o�_T�صvK��+�	@����KT=�J�π�� �_�<���w]*����j)�������T��-nθ�pkDV�fK?,6n�U(_�N��N���ʅ�
���g�W����&�\习�̒陟M�����F
�ybM�MB�hKS�����`
�\-��e�!}���5�n�YܯC�9�dk�[�x�|�z$b�O4Q����?��WW�7�4�(%`�?�QQ��2E �My��?���xxЦ�h�d�H>Ek�y�?���/`��kgA�yZ69̥���QD�=�L�+i
����q�2f̑��,ވ�K$m��7s�cq�8<��_P--&-+�-�UB�j6IB4K� �W�Oo��Q��gJ�n?U/L���X��ͬ3�=���`�:5�.����y�Ri�^�$�ғp�KL��k$͋L�Du� =�$���a �:��2%�,�*��4+���g%_(B"��P�y�i��R���'��|�1��&Z_%|d��Gk�\G���B�ך��L�~�͡`%;�A��e�g�]�@��b��ڂ��WP��B���U�������xL�]��[�y[�Kܲ�>�'F�z�R�Q��)��+�H�e�� :e��L:`�(&�L���"��*	H�����NƝ8�.M�w���Ay�zh*j�<�fU�I��vη���ό����K��JGM=>_����U�Pw�\|~D�f�JW����'j˵��>�`���w�4�L��/�i�A�h�mgvF]�P�����l2�Ȍ���d�ُtJY��GjWKD��RVDa��%�]O�&��~������������"S��ѵ4��vOV���iJ���h=���Q���ud��Wܸ��`�NM��!��<��j)k�Zٸ|�uC�d
�n#�>��"���;� �����>���W^�2�������V��Q�P� J|�1|*i����@B�V��@|I'`��J4���^���f�"b��q�e�=Y�3�jb����v�@�#��s�t��R���3�/�5b�+�����Y�� @�O.N׎Lnc`!(�a�r��y��̾շ HX�ga��R��E��{˘�dLy��Wb���{k)�rk�'�-�B F<��hJQ�NKb҉f��3Wj$8�O��[r���!V�TwpO��\ �կ�ɱ"����p�"<�on�z,x&�-c٫m�[T���?�a�@EI/ռ`�8�|���֏�(�,��y�)�,D�`��㎜�e��)�[7Ƽ�z
"2^k���n��/|(�-~���܃��p�}k����o�{~���(��VIw����<ŵ
ya�Ҧ��ga�E;_G�c*E,H��?��'&���yD_�"Q��	�:�pPB�!��ݟ���#�Φ�-�����Sw��?����;D�d纋��4�w�k�����w�M�.Z7~c�,8�sˌ_��rbEC�0h�2�z�t�:��F"���כ���2����s��<�_r�9��	��P&�JۏS���ף��'���矧LK�n��#�j�������l#�l@�*!�ZF���^P�V�Yq���7E��ȍ�F]{컥\��ZҖ�O=h_�� ���g��Z|T��`g�5�o�Ii8q�K�k,Ey&$��"&n����׌�)ɃP6fY�5�q�ν-��B��u���ϳ�o��$,6E�,�UH@�ؤ#�(nžs�!f#����Bן+Y���f�[E�
��A}�1�@��]�M>ֵ{#M����h�E���Q��\��З�t7�T�~��� �PF6�N�"��;��NM����M��x�u5q9��L����j$�eMTū#��qi���yh�G�#�Ɯ��(3q$K��8�J�T�Iۊ)5��~I�W���b[�%��ޘ���A�`�i��m'��~ER�L^�jr��tBf�X���`��	���A�y`���쟶�f۬��~{=��C|�f�ϼ����R���Y!>ӗՈ�L��b�Z�l���m'�/�����1�q�O	�ۂدJ��Y6�>�u6Y��>!l��_QՀ�.2������U��FHӔG�c�#���bҀC�?����t��5P�btHo>�o5w	�tN&^#F@+?#GY���pR����x�8�|�O��)Ub�|�YZ>PP��7�-M��Z����p4�	�#>�"�N��NE~�rP�k]�U�N`�x3Pjbz�$�0u`4!��3
�n� j+�Zy�<Ova��%�{N�'�Q��N����A&�j�&3a�۳�gJ0w'\��穒�@|D���\��%�[.qL�����8�e��Z�,b�1��F)���ظ:m�^��<�^l(�7���I�'Jb��^-'�ݷ�j���P�J�M�Ŀ��jk�ʀ��`��E��>�]u|��M�~<�3_���Cu����A s��5�|�
�A�]��i��`��$X��5�z���a�!��D3m/�<h[<��"��Is�x���N�%W;�vf�A,窚��0�ې���)`���O���iN�`�(^x�fl:n�6�5?�M@���'��z{?�N� <�)��r�;N��
k/+��]8 �
�ơ���K`��J���t qiX�Ť;�%D��ЖW+;йs6���0e���416$�DO��̈�g����[�B�sT���=sy���_���*j��w �x�_$Ts[�XVU~�*��F�f��r�R�ޏ�U�w���8븙��� |�y�֦ϖ�j�{{��m�ۿ��T�qU�A��0�8�}��02�1�K*�-�8��f[�/��sR@��}�x;�[����!�<OpX}h�{�!���ߣwaQ4ˡ�Q��Z<YxuC���:ٽ�o���Y�f	ͥ�O�us#?ZJN��T�a.{�W[���.�� �aE멧�#i�@�!�ߢ&��(� ��x��WM]�*:El��J���@�]sv������y<�����Q�5�������(����,#('��AHOk��5I����?�������Vv�����=���_S�oi�ĤFϫsh�$�$�!�v�թ%��|�Ǚf�{.O,])��]��nc��h�O�8Sl�!a�'uxf9Ry�I|���y�ED�X�׎~`=���nN9����x��.B�`�
��idg+z��8bT��� \Ԣ�<�� Hg���<��{ t�u�@�*��b.��x�6��[�$0�)�jK��5�G���LNp�hɶ��r{�s�`v.������A]�"dJ�7@9 }��zǣ�����z!J3K�+ �(�L���}�z�#c���������g����;��o���ٞ����O��nSo��ʼ���b%;k���5�,8�cNy6Ԙ������#�"B�)b.�Ylke���{�L�|G�]�c�d+%:\gңޯ3U���݁1q�
�%��8�U�.��zHj�p�É�`j���?���= �Oh��>�TJ��ePA�nş�р�딪�=m�4çG�>zY��G�;�;���/�v~� ���/UVھM����]L�C��P٨�����+R��djOli�Et�>

vu��,"��� 3<�4�IxQ�h�Q>�~�߀��O.���|}��?�l�G5��[?t�c�O�ҸV���1W������!����V�b| �jB�2x��8�^B�a2)��#�#��PË���Y�ݒO�_(��麼��`��j;��Cz�=�S k��t�X��-Y۬d�1��n8����B˗g]0�í�.����4˾�N��� ��r3�-z�:�*�C!˓�p�{(�J%!t��,%[�p5q��?����<�\�=�X e2ݙ#euJ��!`�:����,Q�*4�f�P�t��Y�{�+�B1M�HV��dzz~������¹J_ge��][G�Y�<+�-�y��*por�S&g���̐A�Qͧ[{r�����&;�pW��]�1�-�U�U��EpF[�Q�H�T��R�"�:�B�N�ǉ�M�-����M���1\�N�k�����$�
�\��GD�eK�����T��s[���������NS�%`!'�Ԃ)��(gV �-�\n�&O���q4�jYmklî*%Y�p?m��5h>ǂ�_Y�	����q"B��*T�� ��"u���4B�,����*�8Hy�j0������ur	����3D([�O�+L��.����6�=W,�A4��S��a��8X�o�UѸ��_Ĳ���n#~��"&[R/��4D�z~�䶪�Tj��־��������
s�X�]�%�W� �������"<(��;��Q�g�늦<��M�@ʭ���	�����w���!�*�qm�4P�x[�	���ƁA�J���ʶ�9!��Ϥ�3��h�������P�N��L��P���:�Z}���iQe�^���p���i�Q�SC�v�'b�$0��y`uS��X��J��3v�j�u"'~"'�A��"2k�)qIm];�u��gB�C��Թ2 ���~��zyX��۰�@4�|�݂�����J�6�`<Q���B���;�;��|�%܋w�mf>;QM�^)�W�(,�l�P<�K�A
˄���U+C��}pR�n�N�2�(�6�x�p���呫�І�Yߝۯ˞mp��<�uV��l��I=�X�2�?+i݁d�g�fC�>/�}��|\�����f5�fm^�B,'���*�����&��dR�d�wޯ�{�"�g.ۑ[j9p*�L����zk�z[.�p�=�g� gu�u��e��Z���n7�R�Zc*��Ȭ���	c���1�A�}mT�f�i�"/��S+�LҰ��Eؓ���v�N�+$2�֦�&�4���{�"+uB�����s��.��u����+9j$%;����&pt���](�Y�*��S�����t�gt���e���ZMB�r��7`��\�D2K D��,6k�Z��5�α|G� >i-��cwj����؜�)�w=��@�-�:���t #�˧nO�%&��m��� �5�>�ѡm���Y���L��I��#iF
Qv�H��� �B�>U��;4V�̺�Wp�gX/|:��2r�U�@�ѰJj���ĖK�Mw�X����Ȕ_�*��vb�RnĂ�llLi�i)�����)�P��n�iR��h�r��/i2�D��RŊN284���m�°I�_�G/H{E�J�'IJk�	��k�S������T�o#3���*�P�45
{A��X�Bf��v�>������x�A�f���6��@^��Y.C\9�6�FN��H���L���3C;_��_D's�tb��X=%�>�h�r0���h};�ڕ`��t�H����r�:�#K�֬a�	E�_m�0J7�5�����C��T�/4�^#VX�:{ž�J���)���<{R���ih�-r��jTO�ё1;|�5�AO�>�+�P­�Trӊ�s_��e(��|O�+_����+�[R�Q-ŀ����o�&i)��ӘWJ7G:� �l#��7��rbM{ zg�*\�Q�������5]w���p�܉RD��~%�������$j=UfŠT�&��Z������{�W�Qrx��
�<?��_Y��m5�'ђ&�Fk���p�g�T�L6QI$9�� ������"��m�x�Ŝl{���̻D�v�qA/L�hDo+Z���>y�{>Y���46�F$T-t�>�S����X��*���j2�16�*�j^4�?�.aYC��=֗����[��5
(ϩ_YJ����re�حF��P�o��"/�����﷕Ý��ݢ%���׋
�(]T_%$�h�m�`���k����>O"�9]>ö��!�� 0���w7���yZ����{@m[��m��7S��<8����E��\��ļ��E� ���0�15�	&�ٛg�+��_�Q"r%�����ɼI�o�֭�R��`���[j,��)n6ɂ��	f�����c�1�D/� �� ���WeL�
 �����@|v?EEP�9��/����n����m�La�XY6��@�f]G�T?�L��~7�J�!X��Jp��m|�P8A�A�s�ą�CK�T�R���곦m:��g�Q9>�;m������?�i?�\�MtN�+��Y��]"#�g*bh���)�Y)��&b��t�ʉ:�X��x+�;ʹ�{������[�j!&A�:�&������A�%�<fl��wC�04>J 1�p�*����J(�����"�=p��n��ù�S�E��CG���Ł�`�pX�:�����K��~ CA�^�pA�y�{K�	� ��61�}����bk���*���`_�X��J�n�n/U��f����!T8�7��?r\C��'bi^'�3������ٲ
Ϭbyf�ń�u#��#�t�i`g!*F�忭|��\�����i&=!�x�C3a��'mY��nMl�}&�;�� ];]�r�R�����C��h|��"���&�k/�f-�u�}�Ӹ%@MW(Bk?Dx�F�]� U��Z�d�B-Q�bl�����ò��`��.�"���iʫ����� 4	�gn��-I�� y�,f���
iU�B$=_�+͋W=�|���-��[����F�xƲ��Yށ1RJ��Kq��_a�k���:x���#T#�����7G)�(��C0�S�F��Ͷ8���5R�;�������Nj�R�v&]�E�["[�画u6PG;ӎ΢?Jż8(vE8r�I+�hQ�^}2���&se*Q�2�r�4�����T�����sG�ȃݮ`���Emny_]&���)�P�i�����ys|_AQ�hg��v��}���P�Oi�,��m�m�F#SC��o@�+��-��g�B���vfd�q�dSd$�< p�ܓiI��hY#&�d��4�՜�h~>�,;L�|.��������0�!��������~�xڿLKa8��� t��q�w&LZ��v!�YUfo�.,T
��A�Y4T�5�%� j�&z@P�S?Fw��ў�K�t���|���,�ݤSX�f�!�u���m띸���]I��ox�9�~`�1�ۉ8ё*e�~�Q"5ﴤr�M�����޷�	��>4��1�V�Ӷ��E�7ɬ�2DG�Z�(��1�i�O��Z�5\�1���ҥu�cj��"2|������t�Zr�"_�SuU7[]l�׊��[K8�#
��-~�c��$���N�|�x�F8��7��V���>8j�Z���&p�}�N�����%А�b�r�2��^)Z:)͠�i��b�ଝ3���b#{����v���@�bV�j�:T7��O�:<5r����M�S�&��K{�Z�=Xf҅��Xv��\B�W����t�c�7�g+ ��J1�2KV�զ�g���&7���t`�_�k�O�a��Y.�D�\έ ?<�d.ƹ�令SN�CB�v�u�i	�%)�p��	S�0>ˊ-	;�/���$�Y�@�=q�^�Kj!]�e8<�f��� ���e�>���D#׆#݁6X8rdL@_�5e�H��5�!���vP�x[�yi7�A供���Z�ߥ�9�_�	f�@_w�G
Alc��Oޏ�N���_'�9_:��_G��z���6�$���{��x|����>��*����� �N�)��'���*�~*���S������wyI��-�sM� `@j�e	�Y���!��R@��@�8���4�}�J.��1&�C�	� �c"P�<J"mLv~���������~��0QKb����ّ�{p����q�(�J��Is9?!��qJ������֡-�-�2R/eË�����Fٺa�m�I)�%�d�T�F����L��I�5��h�!�����'���w��s�fB����\��	�����#(�|B������;�S�q�տ-�7r2�h��&=���n�I��8N��c�Ea�I��2�$�u��o����X��ha/�2E�y�7m�>آ�:Ɋ,e�e,�[\��6�������-G�(@W�߰.w���D���I܅�g�*6�Omg�L���6B�|k7�x,����9Z.4���@ ��\MǠ�㢂sL1����~&�Ch?�s��h'� oX��x��!�l�*s�x�����a�L�/����/w�]?��G������uٿ�� '����R�x�*�_�?�!�M0�9T�Yä��u'�c���X�k���=�k[Ye��ƪqa𮻨��`qO���	o�W,�m��
ȯ&��W|��1���y��y�� ��S绀�=N6BxD8a� v
�	 �ׁQPه
8h����v��x�X ��w���������s0�R��	���am@�@�N ��á,52��U%L�^����U���b@5�k�?�l/w<�Du�z�I�O��&��5�P�8Y�)~��fW@����� ��>�ņ�8�}��ٮ�
�G�鎤�E��Z�67i1[[Rqjq2��bp��!<�`�u�=�s�-�L�(,Z=;�����'��<!���@���1!ަ(`�۾�5��%2r��4�8�cWj<O�>��CD�}U�D6�r�)�}����M~�D!,&1�5Z�D5!�*Z�Ae��5��z2vT�ӂ�jp��+�ZN��gy ���Q"G��j��7ߙ_)��	���-i��Twc�]gowhЈY�ۧ$jf����:G��]�!���Q���z��4F��f��%��u<��!��2��n�}�{cEq]��Wr�ʮdUXe�+uv�%�i9y����C��Kk��� ��z;ڽ�E�]|׏�����+�\�9B�έ�X =�1��U�����Y��$���iZ�g�6�@]�h?���_~�9��]���%z���CQ��b櫳	F�k3��n��ˊ�n�a�?�����<{���5�͑�DT6y�'�������q/:ߡ�[�����0�����C��sG`�����K%�O.)��5�yN3�;o>�%��t���;�u��-.n�q�͏on��+OQW�M�i����)2�ɳą��4ɯ�/��FEI�a��7�h��Ϩ 3d��:��l���Y�ˏ5���"��/'"�Ċ~_L2���#�<Όb2�|�ex�a��|�$��pj^���/�X�6���N��^\f�O�d֙h��''(zq�T���ޭQ�6�bKy�fy��t�ي���(,�s"�beҤ��=�b���i��s~�h�ڛ?�D�j��O�L�*Wb*P�E�ҝGpr��i�Co�c�Σ����;�a�N�vA[��fu?m}�P)81���;�3�.޴|���j�����M�nPP&�����Y���G�&�N1v��wٲN�K��Ә�Y�ݯںcAI"�#�����Q��Z��(��o��a&�}�?9Z Z3��b�h�H�Ru��,Kp�Z��Ivll�җ���'@}BYypxMv����"h	
�l�jX��k�, �QE{��{��.���q��}�My��F���j��"��U�y{?�o��B�q&�pE����Lf�kz�#�bU
�b�ݣ���գB�VN��/2�&�i"AT�,5�����k���t��[�rn'ۯX!`�J9���T��!���z1S�f�V��������6�A��b���&L�U�A�-6B��/�Q��y�lm�*Q�wޱ?����s3�0{G����b���w@�F�>#��<RUG�,џ�7P1�k�`�Dk%�w6=�w̲��u����#r�-�~�q�����QB����҂b��:+(j[���R��Zz�Q��p{aڟA�<�x<����/�Pч��kpgx�
��U�e���538ćh��X3g�4!� ��6� �ZDI�]�?)�L%xN�*�Ib`7��ݭ ��,���1�����`�͠��-�0ȵ���8��ݑ�ᩇEUX�)}�P�:9���c�}'�x��c�5D)XQ_���ZR6p-n���k������t�3m�������V�Ν��J��s��,��[��no���r�θ�v�[���N��$�(��S�G�ܬ:�&��������0�=�P�$~�34	���)�Q����\�&)�@�S��o(��(��Dc����_��U7͉� P��]'�O��G��]%o����`��r����k�D�N׺���ч3NH�&A"�D%U��D`A�{H�zs"�6ai����=�"�L�U���1UN�0�E%Ma'W���{@�iQ�
�U�5=K5[�C8��{S,{%�jj�N�2��� �y�+�bb���~
y�/Lei���0WI�܌���4T���#�Eq�H�fYU	!����Wcٽ9���{�a����=���r�O/1��p,8yS��V���J����@ݍ8��mi��)�����Yb��"���!��{��(>���o�x�dd$�f�*�j���xM4�;�6�Hm��d_�u�?[	���QU@����i��ܟ���_4�j�
��"���'�3���ں��� �i��yi��ȡ�#���G?�0��ְM���0�Yt��e��c�6㙥�����QG��&�]�֔�T�et�Z����o��x\cA �,jF�z0˓�J�)�ǰ�};�J��f8��$����(�7����,WP��R��6�lq�����Y�0�$ZXXlr��v��+��g�L�_��JdU ��M-�g#ɑ�� �����j��O$P�r���+R�9���S��9ע���/�*�#�/6�$�|uF��,�g�F���-~l�=e���4�~�s� Ԕ%.�:����e�^g�C�D{W§s��������(���Ϯ�ʸ֬i?�I��a��b�Af-��xn��k� 1�p�������(gՑ�Q2	���C>ߵ�^.w�z� �hpL�t�'~��P�mq��R�7��V�iɅV���FƜQm2��a�5i��R*���-v$L�-��pS�c̡�VN\����1�#)ɐGо[2�.0Hx���l���<�|����[]��LƷ�iו,X(jУ�6۲|]��ف�X��6��Cf�s�d�P˃�P��m*��M���.W�>>��VH������4��KǪ�>ꢓ����_��Ͻi��:P��n@���ʏg$�����_#�;���&@�2�	u���7�;}��s8zxI3�*`��8�X��D��K��)��{6$�6���̠�#�>��wܦ��` �)Y��ͮJ�����sq�Sx4���u�\���;��P��zy��x9�j�YH�G��3?.]��~�L�1�Dʮ��+S نh�_\К��P��o_H~ounyDPq��(@��B�)Q~z�ʘXOo`fr���y���+��^n|�)<}=���#9���m�z+
Y߯��')�y����^y�/_�S�BYl9#�]�Ά+\
������d9S�cQ%�quȧY��K�<.8Ip�!���o6�Nc��T�I�s�_���G�T�{V��+�;:np����ڸu?�V(�a�ڼ��� ��ˑ�u&c�(����i;��
��	#F�)�P1��Q��6�I:K�bx�$�1��6/��f<T�Vq N������X9;ޢ�Wl��d/����pL,_�=��=f�������
M��[�W\��s.�����#������
��̦�$���I�ӳ�J�'�U�p;�����&��D�v�I��`&pHSζ3?�K��V��vV�����Y{63����(n�Z(�?��?8
0f_��n��
bA���PJ�;�r�oً:�Yy7\y��@�ýXݣ�1��?C�R�&#r� �ә��M�~�>��ڸ�,���8@DG\U#�K��2���?yN�;��TQ��Z��H������1�/n]���
�W�rЩ��lh�*N\���3Z,Д=_�
�_���|�f���N�C,�¬q�-���\'6#1�6Ȥ`�����]K�B?��\�͡o1���u��P�MM=�4c{�r����nC
E�X��u�:�2���"�5�٨|��� ���v�v{����w�����Wyp�~�������nQ1�j$����h������C��I����m��Zw���=z�<M��C�/\(N��V�_�|ժ�{T�*օ�e�+"�Ֆ-k�}ٕ�U��$�"�ʦ�dW˱eZ
���nZ�������]{~�DX�j8U�M։�9���ZP⸲EQ��J:sfā��4��*�,��w�ݴ��ZDO�}��?���\�����5rƞl�l鞅@ ��)Q�VF�y0�$
��ߵEw��?N6ڑ���s�¿�x��
{�V��v� �gE��f�x�{��'���s�(a]��	���L;n��^m�2��P՝��G���	Z�g�y,w{�{��C�r�����L"�~���V��p_�A��1�%�Z������sAq���� ����!�qslYM�u�b��I�v�GW08y<;c�f-lH��֐+7��I���4|�0aJ��mY�p�
�����X�J�p�~q����*Hld8��p�36�a�L��B��՛־���ۼ���X�����m��%T$���T��
���Mh5c�����G�H��{Of�˿������+l���t�ճ�|/�Ζ�I�7!�y���Z���kR�T�"V���y�5�+�_�D��o���O��:�e�5��̩����������1/�\�i���q���+(�����/���A���9	>�OGD�YS��R}/�^���̉�3�`/��e1B@�jC;���6g��w�@w�S*�M[˛.����%MYv��{�eNBm'��)�G�xx���Tuc�������:�P����dm�p��N��I���;w��G��1��%p�M>�N�k2Eo�����/��pgH'�|�ء�-U����	Do�[L?������2��x��~V��+dX�O�Ѷ�B�C�_ۮE�9�Z�* ��=d?L�z\P7�l���`Y������]�r��]�(���9�ƚ2�ſt�d�oDktVA�/��}\#]�&/�NR�^��ֵ���hI*u��3��=��G"�T+;FX�^�]rD�hB߬��E.��o�� ��z�t��h�s��x�N�p�O��[������5�`e@��`b$N���Q.3��8v�Bi8�_X�@U��ê��{#�#�1��*Xj�>F�N_IU|��EX�|6Ӈ��S������'�D����#E���/t��F��l���{��0F���XyP��b��#籯��fj����f-�ʆ���x�$nojN��w� :H��J~�wT$�Q�Tz3��C������3u��U&R<y��p�E�5\��]�6Q/�oq__�8+Lv�G��~�P�7��l"���S[|����pX���T���ꐥ�%:~R{��Bͫu�
��|W����RJ���*�E D��׀B�%��Wevj\�! Z�o��n2;Q˞I%�O[ţ�9e����C�ň�gѭ+�g���[[{��jR����&�c������z>�{ȅ*��5u��ʨ!/pw��2l�4��P�������V�K)�6�՛����n��P�
��@h;�sQh?%����Ӵ��G�U�>cs����m�yǝUvp�̙< ��K�j������
 �J����u����h�n���"��i�ú��p6'j6|��c8�%/�q�[Z����Eo�0,U�7e��;^/�W:�ք�t�'�{�'��#>�aӑy�*��5��jv�G�f��k�����q������R�▉/,�}ʅ�i�v{�yo���f��0�{<��Mq�56D��@��=n����`{r��;
b���nX�x����u�{���������SH�ƻ��:�j� ����=hW[3��.�rH�c�`G[oxb*If��*ř�数�3)ܐ��U'- ^x�1���)�U�q(��%re!��_[��E��*�ݰ�qV�n_c��5�(�>J�.�[�ώ�Mv���]��`0A���B�;x��JZiy~�#�c�U����.���K �^���w�i�4�&ڭvT.TA���
±��/?���$�%S���.�'5�t�.2�v�Nh����N�%�(����l;�du�d�xp#����#.��S���C��m8A���*��j��"}VD6fjk�K%��SԈ�����b�&�,ѵ3����O&���o�G�G%�����Tm�$�׊i}�/���ܦ'2}���Ѱ�?��c���f�4���9�$]r�r	e�*2��F%@��~�ܭY�� �r|�v8a� 8.C@%0g'���;R̨Q�n�0���	vT"i��®��C�]����" � �y��G����ֱ�!ۛ��/�ે;��͒�Б�mμ)��f&l�m���v�}If*�Mh�,�pt�� O�k����j��]�(-;��UI�z�v+sk���r�k�Ë>TEU}%�)G�r��x�.���(�@ΛP��$�ce$�arӠڐ��������4ۤ�p��u�}�tg���إ�f�����`��lq����?�iI���JiS��g��: ��zP;��)��!��Z�_z4,�$"g���$WH<��)�~5핃IWa�RqKr�����EY���N���$�G��v�/�``݄F�Wj�,Ŭ�E�ȭ�Ma�žcM8�� #�cg�tɥ�����C�U�ۺ��lp�S����h$���-~w�B�{�7dyJs`5�?Z�E>[�q�>O���OP�; ��Ñ�� oӉe3��Ҏt1�x�҄��}VU����o�cZ����<~�W�_�ٲ4��%6�Vf������K+d�m�����Z�	V�
?K�ݩ7o�u�ysh��C�g�]�T�Q�g�$��=�=+F\be���'�0wՇ��ý"���1��{R6�f�w>�sP}�	8D����b�#$y�"�5�5:���ȶ�_zu��Wfom�����EKp1:d�z�E�V	�d���l�SlO�]����W�7-�`����M3S�����	�+}k���D� �%y,a��v����=
L�� B"���?���?M������z������}�b$��J�r��,�o�haHz�G��RcH�ُc6�n��j'�f j�>�<e)�,���+��Mΐ�������Iq�ʦg5�:�ƴ��5�hO�`w������-�cu�'=Ʉ��o)�x�O�9o��o��o�f���b��j�����$$6����c�n�r���XG5 �&�+���+4)���`K�B�+ j������rϭyvV �ӆ����F�qd��L�B�c:?̹���F�˷�0�=uwh�� @:Hf���1������+��w,�t���ц�C�V 'ߵ`�m� ���-�gjHe���E�%���S��(�*N�'��������������%�#���o�x�:�y�C�N�[�C�F��P( �,�DĴ��U��]iw=C^��?��:Oj�i���9�Q\%���fۼy1�B��n��p����Aq%�T���e�pPz���}6"�Ȥ�,�qP`�D����{󕇩��"���'d3�Խ{����:��cY����C�p����f�ڗ��x�,����ڋ��mC�PY�Cha���d�����������٪E�������/�����#�3��]�������C���ss�\�OE�9ǙF�< �g���x=Hf@�O�L�,��s�J�q���fv��� T�1����G��X�� �0��$���?3D<���N����/nv
�B/���,`�Q���ԝ�˶
*Y�K)�����V���[ݻ<VH�S |F��3�T����|��Z!����h�c;O���N�)Z�&�����N�{T���6�o��m
���ty���5����*z�JW�)��ZM�&%Њ取��pY���JF�3C����O�]!�D�b0���s�x|������#�����pt�c��(�ھ�W�������C��0v��"	�dV�h�=߲�8<l=�*�^���t!فkw�����IZd[��d�?bׇ	.�?�0�l�n�Qx^3��҇�S�S�-�\����_��Q���J�&q��<�g����`��R$��ړ��&o��@�UMꭀ0�v�%8��;���^o�/7�C�����@L�6A{�|:7I��®��v�)l�B��@O��~q*н�
�>.�)���ÄQ`��]	����H�˾eˤ�>#�M�Ep��)*��-\�_7{� "�͒ũ��I,E pnRX{Zi�d1bYd�&3N[s^!1(�l+� �-�v܂���U�V+GRicw0��g�G:+���l� �wvr<������>uY��|�eVa�I�4���㲘�t ������颥ƹ"���7��������KiL��p�P��s\�*���=0� bj]��A"'>у�P�3o��`�R����!�o$�_�N��੟��{�U��o��`%�k���Q1�.G�"�P�U��i�῀9��I��Ϲ�颇�r�<惤"�B�ف����fk�����sЁ�&����%~�,ղFG`iZ�p�-o2�;��s�A����B�|�l�>���-J����������Y�����f�P��H�5�����O�Y���,�[��7]�CX4@��s����S��Nc�z����|�Ku|�l�eʡt���K ��9�9�x�.i�A7fk<B�O3Sfn�=��d?sևO6�4>+	%#I��o�q�g3�G����oK�����O��^���� �`����p5
qa����i��H����3I�*p�L �|cn�<�{�d7�h��E�qV_h�݈&Y�X+�gQ���]����(27��,K�pt�`���V�< ��
���,�G�y�{�K`�Fޞ٘B2J���_e�َ��=�7��aʂ��G�ӊS(�E��~����Y�
T���f�gNq@nY���37�$1B�eɑew]ܖ9)���� D��*�I�e�Ԃ|\��/t�-rR���[z�Z4�I�}5>�L42�N��`���/>��)�������
E��{C5�V0��L��F��)�|�L�{O��p����XҒ����\��D�y�0���+�/ǡ���� ���|;�#�.E�b+I�i����=Ww��S�ƣ�|ky(@�`��T�?�JZ
���]y	���q�դ�Ou�]�ǲT��eY篢g��ܽ�z���w|"~O��v�W��s��4x�,�J�� T�i3��r�R���;R��:�0�p>�� �L������)�	3��$�$�-_�u��I���f��@�y�����E�����a���GzfA��|_ޟ�!$�6��gʂ��̫
�Ţ$��F���vM�H\��B�֦�������G�=�-wAI������)��b��䙾���t�C���tM}?��L�G���3��t�YM}R*���^QՑn$�DH%�rBx/�S��ˊ�l�q��-<c׭*�v�Ql���^�ʆ���L�)�A�,��@? -�D�8��8^
�ɾn�Ѳ��C������$%�9QM�Vs��
�fn��j�(�)�o�����0�P @c�	�bt��Qr���
۝s��9�N�JWᘾ�#?0���-Cd��\^y1��m��rV�jGW`�N�B���b X�	���}��������W{�A-ZC=�kn�ن�"��0��g��co�G4�$7�:�&�z��~_�k���j��c���`��C����5�5��R�Oe�:4�'	�r��s6�.�􏳜�ív{�}[V�*k�Q����g�l�0��h�4?�kN�'�D�t�D5��G4b�ʽW@yt�'�8z`�����C�'!�ҙH+yZj�H|��t��جųj�1E�S�1����t�x�R�`� r�I)�;f�o�L�)aWT��+�/;g� � d\�$�M�P�i(ͫ����xP�?���;�c{�h�Ó׆e���By�ez,c6�{��6x;*�z%)̾�V��S$�fl�C��S�� �A;b-?}�.?>��$_Γ�����l�R����w�%N������w#�ga���+�o�*��97�#&A*�+	�c�'�Ӊ٪�yZ"@������ߥ}��s����l�M�_ݬu�@(��V��y�X=���S�"���]u�%C�a	j�V|������#��=y�r ?&�0���=?BUC�4�è�ֵ���,�M1����u���;JZ��Sd�=��䝛�;�rn-:˰��J��y�V?�C��ee'���tEL8��C�4�䂺����hmͿ=Q:��r}z1w�f�!��
ηt;�x�Y��G����4�O$��0n�$`�u)���a49��Σ�uI\1�?�4���jc����e����,��&�	6&K�@�|�v�eFXgxi�$*t�����Y!`�RMݝ��`�훭�!��!��krr`l(��+v{}aL�����Z�oH�����9�ʠ'u;i�u�V�{�S��gu�@��${DH��&Y�P��*2�U���G`��N�h����D��.[Q+�$J��&�ṡ=*����`L�+�)h��5e��/+>y�Q�&C��٘]z1���;RBO��uv�<}�&#�Z~�g�Ķ9Wь�)2��=	�8t���*���?Ǜ�MC|��0-4�M��K����qJ�rU?�-d��or���?��V��ǉ`����Y@�_�&�rjv#	�%c��Xn�x�8'W)�H�7�)�w9�śđ�heqxr�1�.�����G���əd�i�^9ȅ����6����6��q����ΨnF!��b��~���i�EN(��q�}?hݞ"���IM�@��R��뀩�	zT�P�3��S�!�|�o���5�;�ra�B6m��J�p��w�@�,w8@�k��G�"�ikjΌ�v������-�ɲ����;�Բ$�?tΦ��b��z�����۩�4ͪ=R���
�4m]��KB-��D�U���"�i�T ¢Ŏ�������'���S��5���q$���T��A_6ԯC4���xeM۪Ǭ��,\u �j�o��U�Or���✚��]�@�b8��u�צ���oOJ]�W]I��O�~�Uu���wl)����DpJ���Y� �%d{vq����{Wi��p�i�{���H]�]T+�3�����m��:'c&��
�+�'����tuG3	~�t�Mԣ���x�<�#Z	�;S��2��um����J�7�^
YM��5�D9�x��$�Y��:��׈���A�������O���!��Y=����&��e%��X�ʅe(��� ���q�֨�a�_�D�N��N��+\��0ͅ����p�->����_�2����k�8.���D��RL����F��õ�����&CΏ	qJXB�w�@��N��tAU�]F�QC�݂|��*�#��9\٣X��w��2�+6��э�CC<@�q���� ��Q�i�P|������U���&�u�ycr������ߨB����T@���1���tC���X�vI���F�]W���F���=����t8�x�,�5��L��A������a�Zw;�X�>���㏙>�'o�C��|�S!�:��I�+�����}�-�衦��b[���Nˢ^W$�cɵ�Fv��M�}����'J>J�>n��nK�XYa�����s�ٌ
E��'=�S���#(����8@ڐ�N��]����0��.�-c��siAbT�i�7�s�r��;�_�9�/�n��8ӹ�6�G{*,$�H���@�ws+�S��c�� ���+>��|��ޑ#E���͎�a;�pd8'�@���
���nr�;�k9��aѳ3�r�*_�uB�=
"���w� �&�ո�� �LV��%o%�0�l<�╤�aN�Wt������G�Ʊ��dRf~�Vu�U�Oi��<>_M�󕻀6G�ǰ�~��6a"W�V�г�|��dpǝ/�l�u��ѫ�Lu�y�u���S>Q�2��%�-/���#^vLVF���?�`DT�/��Í�0G�N��F%���@����������m����g1*[�mWy>29x�#�|�F�x^⑬�ѡ)�밵TH�J]�	�}� ����Po,������8�[+����d�"Dq=�v�ZsQg������.�A� 5�C�.�*��"�[x�l�H�cS�����*#y�<-,mF��4���0�d�6��-aP�yզ�f�}oh�Gc��!?��~0���h�h�1'�d���b�M����Vm z:A�N��Ƽ8X�!�[2�Q�Bc�����sĎ�"��%��0@����%k���G�Hj-UU�6}b'1��+)���\_jυK.fu�Z�"�MLZQ� �YG�z*�*�۳�_ĕƱ�!�ԫŪNKU�UzA�f*�+�է��<�;��	>r�pE]�h�w����'�q�uH3�S�O1�\�%�l��|�c���%��!�\iaZ�H��w�E5QWtV ��-�I�My�g���!�MD՛�itJѿ���s�uq�.�Ǜ��A��l ��)��~j�)�F�ȔPy��;��u��f%�O�"��y^|��r��^`��p�+P�P�iif` 	�ac\*>�6�X�e���o�L�*��xp�*��+�2F_EZ�Pb��%;�n�Ig#�Z��+��O�ٙE�g@�n&N�a�FH� Ce�����X�g�s�"(��o(�>QM��� Z���⅔#v3�������$O��V/[���j�%m*���ًhP��z˞z��V��fbU�ٝJ�Hqv u�?o7&�Q���=N6q�Z��Źcy�^>�I�h��� �:�,��s ����A�Lh��vƉ���D�Ջ��z����"�$�Kɒ��E�ɇ���.�^��xۍ_�q���;���6
�e���f3�$O+�LEK�I䢔��j��Rbj1�?�3+d����n�����ѽS��2C/����n��������}-�¶��9r�!���1a����o�G"�D؍EM���<C�'r�H�,���S���FL�uV�t�weh��`�x��ɮ�Wv5�M����q J��u4}
EG���'��o��F�J��F�Q�@�������>#,�ʳ��P:���Jn��G;^�?U�t�_�D�K��^�HVau��F��ͤ
��ezA)�>���|G����n����Mh���B��������o�-D��XE�N46�*�0�I��T?�ߗ�YD��}n O�y9��D��<�n�|���F�:�����PC���i��<��9~�UÇ0[WA�� ̤l1�x쎫���rx�-^�J�2k���4��m&��.�&&Fu�i|���b;I9��F���<������]�ǿ��fa��=0�Hf��s*ew"�gOeŃ�>�5�x>. 4�$(��˂K��!7�?�n'e��4�@���1�7�?��oզ,����I�k`g�!�"$^Lus<�c$���{�ﲀ;��z��CQW��1��-����9m1>���A��J�{�qQ��;}[��c�<RJJ��� ���кH�`I����D*��O�ʊ�]��4@@�&�M�7���Zs�CX+03R#bK3ZTTH ��y���%��=`��+���V����\L3"���^��S�
���Kc�}*�Mz����V���&g�H�T|�eۻ�7��B���$q7�a���=K�Ƒ��sC���y8��#��	 ��e�5ؗ��Q,H߈ғ�%
��-8�|�L�	:�0�0�/���р�1�\���=%�u����܃69�ya�'Eo?u�ا��K��`<qM� �`����KX���M�������WS����-�bԂ츲$w5!���⏘����َ#���4�3<;�X�Z&�6�5&����B��UZ)a9y��vݽ���`������>��֮��a`�@j#�5y��
�<�H�BcUx5!���2ګ�#c��������0�)V!'΍d��L�͞�3��\b6!���i� w)�d4���d���>JR�M(5g[�r
Bī�7�(��	��R�tM�K��s���ϸ���i���k��{�С�K�4�lwZ|�?z=A�a��W|�i��|����	����/A�ז�K���>p���X�N2�w��U��5lz3��������_�t)h��	�֝S�m$��������JqD_d���$߮Eh�nI�zK�r㋕Rp͝R������)t��V̔4yx"��<��2��w���m�%F_�_�܎s&0�G�~GC�Ut���ł��4Œ���)U��0P��*S���b������]�a���ǫ%Αq$��������
ā=��U�=��:��h�ߺńFw�7�,p���O�Y>
M���&��n�k�`���^��F�|�M�ʜ��N'ܿq%O�l�
ٶ��ZPe��`��;�_+���Q��A�t"�Z��� �5�c<�,%=�"�N��PPlb�F�g|kT�(��\~ɫ\�"��E�$/�~�V�l3��q�Ր0�Id�'�£xu������ri��������4��o�pJn9%�&��V�!��QJ��X�+��u#�)����R�ZO.����R�����,..�4�_�`<j�#kK����c���g��� M��Z�Ӊ��B&y�g3E���v���qM�W����t�|I�>�0i����+�܀�2��{Ay)��|�g�2Բ���/'��PԘ`����1sBq+Z��\���S�\6B	��3�UՒ�X� j���؇s���8��?���z�m�U
�\���ld�bƇ����ŀ�@a�\��%"^Z:�!����X�EVw3y�c1Z�U�<���DVL*�M�vTG��$t=W�'�BWֺZ�^^�P/��:��#�Gպ�/sR�gQ�9��Z�7��׉ph��u3s�u���޸�1	�t5��S�IEq�8�߷9�3E�v�:ȏ=x��52�gh�3�^�w�½o{�s���m��tL Ǝ�x�Q�Nw�#�����N�xɓr���p,���Wܲ�-�P�or[�F�����r����@}L-5�x�x�0���و�>|[�"�/�A<E�Lľ�Ѻn�+��h��R�g'!޶�(����vl�^��tH��z�t��hv%X�`v�ݦB�"��f��wg]:����(=Im j:�c��;~ډ��c���ə2����@�S �b��6>A:*5���*�5��wh���t�D����E��U�p��t�T�H�m~�`�)T��	����&kǸ���-�*
��������(���T�J����D�]	GrX#��m.*u&2ޯ�<`S�lp�ɻ�k ʽK$뿯0��=~���[Qz���d��J�K���JOW'X���P�d��f
�b!�M��F�����]G�B�R@��RY�踅�ѡݻ+�ˍ���%�.5eod�ݧ���p����>S�KK��8�a��+>���7�-����eܳ�EqʍC
B��"�.�
E/�+�Д̚�&,	��&���z�T��c���~��Q"�a��К��萙�� d���&�Ņ89�TDZ�^���8eU�+1�OZ{6���rd��Uz�ٻ;��z��p[�xy�O�ӓ!�zm6)����9}�T�M<JRL�@`/�[PMz���Wy�c