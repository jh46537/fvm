��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbж��ъ��/�S��۬니]�~��8�?<iq�:N�?�@�V���}��¸����n4�U(�ѿ)���R+bw�T�- ������t�HC�iT��	x⫂�K@lʭ5�����ƅ��ё�j��%q�[M��d�D�j�<a�'߱�~�.T�@��?K ���l�_&$Q)`��jR_c�K�l��-X����n<�9���v$2'
Fp!.�n�<l�����qt�C������;?�󊢓*J�#D,4��w~����L�>�n�|`Kڊ+��4��&��^RD�����&����aA� �@�A<+jt ���fH����'ܹaU�p܅��~+"�L"Z���V�tF����}��	 ����l�]�X�ڗzm�mX�w\�I+n6fꞁc��S�S��B�L?@���;�9�\y��x�J�ǖ���Q�#G�2����2�#`ݣ5��A�h!��O�����U���8�Җ�?�h��'?ġ9!/)��<�F>���|]�Y��C_J\�dGfk�f�p���v����fĂoHC$ I���IGUEi*1B��f��{�O��uJ��T��Y��{����F�����\��P���0��z�/[��l�v?΂g��3�����0��%w�`Xm���ey�&{� `�9��&&�1�#HE:n�)�r=u]�@X͋Wa�4y�7�	��í���x�0�w5���s%-��!Ԏ)�e��D]`�U1���w~7��ħ}I{��]
d����̓~0�'.Y.p��1E��_0�4��E>@��'׶�)b�P�� '������7�zW>]-��K㾒�k��?��H��d�L��p6Ѝ��$�+:ahI�\tlҷI=.1-���8f0 �ˍ|*���O�*��U;��ҡ�/e|�'kQ(x�g����ri1a�d�(���JX}ǘZNZ�z=�{���2��F�m�>��>��ɰ��v�¬������C�R�;�]��i$�F[���ȿٌ�d<�ip[>f��qF����j����֬��x��! ����<�ڞ��M��8����rD�kÎ�є(��w�sp�[��t�z�@�n��9֬�x��#��d��K�H�D��D�Q6 �H�]<}����M/��y{�`��"���a���zb��͠Dg{!w_�L,��k��7�t��&�Y�Ҳ7�D��#t��	��rA�&&�g
�%	��y`f�|� ��pt`
uzB;�C᪳]:�4��_qs/���3�C��>��hiͯ��Y���"��nӲ�㷛�"͍�sӈ�zZ�,����#,�9�C�iJ�W��y*��+�q)� �n��V��j��P�Ώ�"��0���pZ����Ě
�����9�_��'�a��p��󓭘�����z�p����]�.�|�)7X �IB�:��r'�"д�ׄSX��鰖[p������v��[��5p���z�YN�@��k�<6�qo��M�K�@��!��2��B" cϐ���B�xM���to�5��u�4l�����b�,�x�8 ]4!���Ș�]`���颶]:�Q��]�Z��:׾���]O�'�o�䝷��>�����=�K��
��'w��q�^f;>��$�KЉν�����(�c5�qm$�rź
�$&N�&�-�F��:=�W��S��V��*�R9`��."�l����\�S��L]O�])��R��ҁy��FPbnm�Z��D�n��|)�Z�R�X8,U��y}9�g(.^H^�UԂ1�� V6��_�e��ڗ#z�4Q®��������K�M��)�7�����e�,cr��=_É#�j&�d<�(���B$� |�~Xt9��b|�7�J���٢�"Ē�\��5���$x| �N��([ 6��pc?R�e>bҀ�����΢�w6y1����D�����L��p����$c �$�˨�c#�X3��6P3T��5��Y������1�帙�>���GIv�:�,�O��ʂEj���\s�O�s��ۺL�g|�?���,S��h��W��zh͕�J�����h%BC�=�˾�PDI�Q�a4tn���}.�Ub�.vVvK���������WV5�Oz����O`Xo]���Q�.'Z(�@��A��������K�|۔���=a���}#���?����@�RmRZO)�>�տb*�嚆27�s�Bf"��+�Wf��6W�x֧z�wK|�G+��w�W��߅�:n��2����=a��1n'8~ W�z��������ܞ��H�^҉���r��r��.^��TK�L�y0�`ב۵�uz�{��r�"��ky��v��?�{z[���tE�N6�u2�{�ejPW<+�V�Mwk�ٿ³LP]ء�w�ܸ�[�=�+䤮	���y${H��mⅶzc1Z/��^�*Y<WP�鶁��
y�FW<X{q&"�GC�5HC��>e�-��L�c�������ٮ>�1|~sk���l�p0A�_�g�qY �'��,�	�;( 	��p�@&=�@{ۨ_����R�b�D�0E�x���޵��d�@(�y���9�t����d5|3�8����^�cZNAY �����.��Ñ�S��T�*�b0�0�7��KA��}cE;Й3.�Et��w�:�^~3�A�m��CIF��5H{��o�����5��M�d����x����Ry��X7��ع
�gS�����W�U��������N_�H��5��;oou4{��V.u�q���Ǆ�m��NbZ��c@|g;Y� �+HL<�#�l�jۃ�5��|��W�ş�1���f����]`���z'k�����<w/B֭��l���}��Z�&;���0tX���r��z�������V��OJK�Q����c'g�N�����	|k����׶ӑ�0��(�z�_�?�o�%��W�&n��f�O�K欢��1�31}�=�I���/Fy]���t��_�I�Q!q��9;d�ڴ#�c
��F�l}
^�Z��I��q��6J�(*iד4%��2�t��3��S�VA��΀��N���@�p&����M�+�2��M%{u˧�����gL��v�E_E���p0A�^�/���s�������pp�o:<�We���
�x1
��{W��>'����Cs�Ġ�7T
��F��a���>�'S�f��Ȝ蜿l�U7+8ަ���t�<�����ٔٱ�BCQ�{�)��F��l����� ��/`Rr�Bs��>��S�Bϸ�T�X�biz�M�wg��y����e\� �L�8QHG�(�;�⩷٧�����	���pJr�w��]|�w�U��K��ꙍ��w��"W�Dڐ:lR]i�fPߝ:b`n�&taˠ����� $Dď�Og�[`	#�^}�f�����	��A�'e"�����J"�^��/����wv����(T�F�"�]��긞���XF������i��]�+��w����N��~4����?%�~����?)L_�Ο�X$G��m?�B���Fu1�Gm�D�p�۟v1�Ԡn��H�c	��mi˲P$��/�Hsia��2a-+�N&֕��0�O�ƵJ�VB
)�)�4� \�l��p�Xr���n�"Z���?��CT��Ƣ��z`���ES��Y~��?k����U��*ll,0�� PM9r�P ��x}�raU��&W�u��B�#>9q���%)U�S�;��:��okqjKLHx�N�px��~#��|2��4�O�bAL���ZߍLMV+A�)r>��=i|�r����3�^+��#����I"<v��n�ËY��Y�i�b8�/ �F��cv�pb�P������ y���CҾW�WMV����,Ń�L)P~E�K���E���m{"c����j;�r����M�����GCtW�W�����>vZ.�OVPz$Q5]W�����ɶ�q�� �]�gj�
)mk�ᡤ��D�~���