��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�I�X��a22}�<�����kb/�1�������K?�v��]�j����Z�3�ܧ�ћ�����q꛻�Eqo]��E<8�s<n!����(}.�)-#��S�Ry[��N,��If��{P+�#n�R�=~�3&��I�6:,Q�����9�ts�2���m n��,-H���
%���k�3��@��\�����d^�ΆVb����͛`��1��?Æ_xxY	�̊���(�zr��*�_��q�]Ұ+g��Tځ�D��:��������r� �:�e���\���m@q-�	1�m)L$lf$�% �;��br;�S��IR6�IpMzGD�/�![�9�5@����l$�2D�-�'�[������X{c��#_�a�h���yͦ)�4�x^=:Y�S��n֤e��D�JYU_c����Ы	)�4�(
��bK�%
�(�g���Zɘ�P�(.چ����Njg�6�lhϋuO�m���l��/���iǪ�؈����a/cqy�-=ɶ���ME�=�)��r��ɰ�D@eHS)�$�D)f)-_����J�u����6?/���U�k��BI�������S� �U�����ni]�^��h���h#r�A"5��;3e��Bb��2��ƦF�f��U���&�E�qqJ�s��x�m$h5��Z��f4[}���~A��^��^��{��k����g��V�W��$ۓ�N��I"���Sl��P�}M��拝�S��5�$�8��j�:@]>�z�:]�6�U���	s���+q�3���F���/�'��'�˃���M���1/C$�ixIu4l�`B[{�Cx�ظ��3��=V(�/�<8��;-����k��]�[��X4��'m.�������V�|�t�p�〛"���_@��������.�{�1/���=��[s�^V���;�@a�0�Ć+�:E@�|w�<�آM�#i��6!��4X�� `k{hL�VW�����=v�4e#eD���"i4�uw��p�WM	�5�iJ��AA����?�I?k���k1L��<��a�Ҹ�Н�C��U��#���8�j�M��s�ȕ���O���"hD�cF.�S�aH;�����c\�6�e/��Lwsҗ|��bz�]HE�/i�\S��1���ί�L5�Tp��Z��`�RhuՍ�1sY.J��1����
�ژbc��ު��UY�6y�wI�l���o�y�D��f
��*�����?)��q�z{�}�(��>��: Gf�":�f%�!65}��~�[�Em�f��-{�;�JvR.Id��vo~��9O� �b����>t��r��n[�3S@���ip��Ԓ�>1��r�� lfl���RfE��*��K�P�������]�$]P�fw��<}��f@���=9��f,/n�'J���݉0�n8(�LM��?�'���E��oA��=;�`�1,�3���ȂsTy�����%�ش�3�6����ӄ����h��ۤ�*^#T�vx���c����LgD��ē�v`P�p,�����Vn�v3_�h�Ǐ`���M�kM����"5Dџ������}aw��E��rdQ�IXmk9�p�
��N"�N��QozUk�5	Ӻ��9��P'�@h�N��ݙ�jq��[\{�DEؽ-I��op�p�`u�6k�����uںX�c)t[����h�6k��-���N�z��`�n��T@'�³�L�i�bǏ� �6.�"��?���Lil�B��s[4rc�1������X[,7�+�T�6z�wND6d���'���Y{��g���g�%�0eb}��i��H.��^)�;Y��88JZ!�S�v;<7��1E7�V
I�E&炄�}3��75:M�u��'�i��%��YY�e�M�jumU��5�Z|�vD�#�<�H	��/W�G���~��ݗM�b�10pEc����V��2�hi�d#i+��╵�&%h0+f�ؑ�b�v��Q��ox�7)m�
��qJ�[���_�h<�,�V-5�����	3��+�0�Y�S���Q�.QU�܌��[U�m��'츪��P����#/��K���"G2�'�l�~1��j��w]和Y�9��c���>��3e�G�$2l>*�]-�k9��4������[K�z
��{�L����zQ<(�2^�{`�QSu_�F�ʢ��4\Mխ��������)�g���b3?U5A�_�������ٜ`%v�ҟ�'��	�h�&j	�4ơb��*�7�u���7�����(U'�.e?(] gΠ)j�}�\�"m�Z�^7D�h�3����qw��洜ޟ5���go�'S{�b�*���/�����e@���֘���V����S�}6�e�v�^4���yW�-ߥ���o�K�����=چq��{@B���]��;�j�qY��6?xs[8}/Zi.ނ��<�)K��%��5���b�D�R�mB1������@Xt�G��g�}�:����WȰ)a���`x��s��L�(�R�h b�nP�lq;��/�M���b=b���4��D���|Ykĸ^s2���@B��L�1(�p/o�z0�]42jkOE��V�,�s�X�I�]�8��
ҋŻoV�����.j"\����C&��Ӣ�k�ᒲe	=�6y/�	�~+,y�r�d��q��Wc�/�m����=R����(0�,T�N.�a.��3��:�ǯ�b��E�!�i1v��E[�?Fz�?�6��r����b�[�����'��峇��u�{�B�]?+�1ha�&ʀ�<g�
���3U������Uu��I��I�U�:���A�D�Jr�|`�������:�4p<O��S�E��
�-���x����Q3����� �%�?|����hb��1�M�����V*n��DzHuE��Bq+��=e� ���itImV�k��|{���i��W��-����~�|5�Q�k����
crf����Y��l(�T#�ڏn��D�'2��,�t���.�^is�[��@�Q��=B��@Ty��!aN�,��Z�}�q,�)V���kπ�j�A)��a��j�#�.%'!}����-wF?ә佂@u�w �7��pZb:��`���c��ll���I/@�[��Ǐh�+%��bF��~�5���I�������
�.���Z]�����K�Рh��2t�X��&�j���
�����Uʭ�"�S�}��S��Ǌ���!�Vq�M�yF�>�l����SOT�ʸo���*���XŌ:�م���mP;<��$���>�8ˊ-�̫�
+p����0�Z�Z+��uB��p��QG�������������f��X��R�L��֕��v��Á��0��B��^6���I��=:$�}�W;�fo������/�����*3�i��Ȋ8L�%&��s��/�yNd��ըq�#j�-�$�y|hAu����)JǬ�$�5����b���^�����ji��JI/n;���<�U��m i+h/ǲ�CC�ShF���t!���%�V���L���ȓ��"B�W � ���|�4��@?<9݇�7�����5�d�<e�TF'{����j��%'����$u�9��HkA�;�h�+�PZ�Ad�9خ���b�y��b����򌜆�eE��RB�vM6t��<� ��J��|����5X�o��>��r���/|��,\?�1�
p����������`>=w��%R�����M������6(���C�?��}�Z*��t ���`��%�`�lTs����l���~dwXtV%��-�eJ�+tq����W�W�=�`�4[���'�z �9.�P�c����bk���W��z`�n�w��(��V�#���j�P�iZd&\�����Gb׋c�Aw�p�"Wί�0���� �>���g��Sj�j��:�4����i��$�Ϫ\�-�
��.Y9�'U��1��U��?T7%`a��= ��C�Ї�\�����@��Ϳ�m{麂���e�tI�`����ٕ�*?{ه|���ؔ���*��N�~uj�qV��֏@7�V2����?�!X�!Ω날 ���a�p5���L�Q����#[�h �QE��J9��~��~�}��1�n?�Cʆ^��K� 1�D��ӣ��ґ�I��/ۇT�7��S�b�B2�Ͷa�J�����c���ǮD�YUw�y�����r��+�95Z�l�׽�L���0N���g��U���'4�_���H�^�B�o?T�F=�%՜�R��g�kT���MK��P�o�i׊�3��
:��}�����I$�sv8 3e�/IU��s��QW�t�3D��QLh����?�n�ϗI�� ̿��u-�+�1u�.�����Ҙ�׊����p�!� +s��A��W�u���l9s��&�k���EN:�C�]�>R\=�c�O�JB�9����@���`�0WM-��<�WX�rr�	#���}2�y��kl8������;��e(���*h����2���i�7�a��&�'��{��� -���$ (���x/�$��X��Z%���!�o&vVAw傳�gih�GS|��� ������
�/�Vg&ֿb}�t�HdBb��PhU7(t��ABT�`IW�3��Jc�`ͮ�q��F�"�2�#�����'OKݵu. ����T�C��|#LTs"ae�[:�bB��x��9䰭_FV%�&���o�C����e�Vx�ϧc$�A�=^)'�����n�؟��ʚ�Ԙ��1K��H��d�ۃ;^�@f"��	��h{�T�`��������xpjh���<�� �d��;�)v�-�+�J&�%�m3}�7�u� �49��f���ɝ��,cZ��R���D��&b� �U����˞>�$ś���mC�k�'6_�	?H�;���ī!v�핦r8���2��Yzı�s���h����6��y?�ktM�QҞ� ?ݽ���8�h�����Ƶ��Ҏ,��3���2��J]xb5oL�x�� ]����"����ĖX�t����F���qE�`�ƛ�{����(d�!η@B'��o��<|@�����o�K�}˒GS��C<�sQ��D����x���`�"i�5j�bѶ�_쮄%q�D'�W��y�ƥ�Ⱦ-���|�,X��?sЀ;���!BS��U����c@̄�