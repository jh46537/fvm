// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:29 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
m4Z6o5ouDE041ArnycI8sl9d+wkXXr5n/d375ETwPTmDmStVF3M/7Ex1a+b0SnJW
LKDfGHloqcvubHAwf6dVccVWByqNNNuWgZj9AqRygqdLGHWb3yUROcsptxxSIvPb
pcx1Hhu5eHdJ1gyCAUr6JTQz/mer5F8jjjTN6SuNUhM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8480)
32ihXXsPEGGZOdvNvbUk85H2z5j1b2BgaOBJFAAtJvax1LXRJ+9FaFyWtPzSkbtR
SVu4bQSPTSae3VSjeH0CfWdgE+0STT/EKLy3XWA6cFUXV1IVMkeQBY+nN0ftuBm6
4fkHQyuiUh0/ygfw9hu3pjdDZEJUggfWhcEcT1O39aP33UCQ/OIm9PNbj8Vyh5GW
535eeBdWHfdhOqpRoGTlpctvzIbM3uiK7cq6aW9LInOMm0QSKpEgJEMzpFJYWy9T
s7qhK+pQU0htRdnoliKcXVADJJxEc83cfY2NNdUGrAsYq6w3XYj/H++lFfOOAn1V
qWhh3VuQJO2fdP6t4X+WUdD+ksoO209HQLJpzjoQ5b+s94IXrmbfAhUZT30oVpY2
+gw6SiqTjK/w0237H2wIqW0qLp3d82sKJjQon6ZvplrK/qWMH8BO79luDGbiovWz
c4pxFYkhEjqBHQXwbGrG98brstIeVF+wV+By4Hj5WdGzKygB1VTRG0nPg0bhkaz2
npkv0C5Ud93rKZw0rt58Klap8+zb+WAqRUPSWXqZHiNZ3LSMmICg+OzRtlkPhgZ7
5QlBAuKz3S9Wq9xhPU/op1Dg65d21xAgxNsCNhIHlJY5ckJZNyh1mY+zkYnQrCoT
n8XaDa1F4rQ1lEq83im+4UN0f36r6CuXpEA8TuPSD5On4E4G8a6EculRW0Q2OF45
FeaY862K4PI2qL4kTZ7G2lLiItitxn1SyaVt5TbHk4i9kEheTsdbZEbsLuYHqNLS
njd+JaYSfRbsaekoHPG/VM3og2aMbCTfDKP39IxBCGCzDlkelfoCURvy0047OoiT
MSNOyLlVAl+DGu0II53+qqbyLVsSzsGcTYz48juAcnxE3+StAyOwYi2nAvqRPqqy
H34RilKo0k1YHO2RPTDNuv4MBtM6xebcETBUWoQFIC/o/0FyesqLSgGtw/y5Wzny
QAIQL+7+04/RTcLr1UxhKfMTwZIQyqX8IF483DsS0yuXtRxoleWDZlZYE07GMAjY
xi/3LsYIkBrQzJb32hKjFS4S3F8DyOFYUF2a4m5+O77T1cz/5CpmzI3BmPrV63oT
mgPUV1vIJLH4TqZeEonogIcdt55aNoX/wPJMSNm3bV5TyAQuS1OKOpSGp4YRZiiE
X9K9YJXDyLKYJcP28cE9aHCq4Ogw32MHnTaeEszqGGGM9QRj8oZ3YUidqJghTXUb
R0NORw0BZsvlQSDHnnBzXYPYiQ3CQS1lBwUqnlsWE0EIDyHCGmyBveq533/3baXl
kWVgcBYmaC4Vbs3CcTPVPq+zYoYGzmwhRQytF5/rxTJ94GbFu0AjIWKEm3k7wsgK
eruj4SjYU3qNAV2QgTmsjpbTna2fcKm2PnJx5rfTxmTDiye6uJhDJ1zYUZtsWGd3
IhbfIiamZDmWG24/88bczKc9bDxGk4g8dooKs+1TPoMG+DNZ+yeVbSCd5CdyZjG2
g2errAGE2YEiTyovL6C81nHowU3DxEZBOclx6+uwPTaLzXziH43/9kZeGb8KwgO8
tigGnLePBBoOvWXxGgXiTf9VKZWpMbqd7dtAb72rQ4nRssZKFsgRHM9Iv9xQDE/N
0z+4TbKR9tPzlcpJh8CJv77moYhLWJxCUEYcP9/QvNH3zLnlsX2pizi07y14s4Qr
hdj8jsx/Buzrg/vBcLpbLnwxOZ7K5a73qfvP5jgpD9tJkqLL9BGCbhlUIxmY4SxK
H88BR3ycikFRn+UEz++aMr8FSHOT573KpMjgbeFIXgEU2DGCX3TaWhvdFcn5TVcB
JE809FObIcOkvh0I9bOQBIVAbwh0pOUOCoBKuhnv2nN5e9MPN9U/EVJJc31MCebl
Nc0hvGsCozD1/cbxbQDs4KTw7iJPDH5LFyHspjisKRSXaV2io0Z0H+uNQvD8/z/j
LY6HINeu+a0vEzlw1hVJOaTrvSVArbYt9Lb8BlXtgO4I6aT4ryn6vFg7kR1xOdVi
LIZcb7qmth8f1IiWyEFXIYkGJdogsdFcZrHYgA3/Xb/67evEUj+ycq79vrQ7EY0X
/V+s+wZW69ZfSyDkwQuHm7te7ymBl/VT8uuH9q0rlK5bQTCbmXkzjKfUCuyBc3/J
NA4tx27I1kBGm3nr1t5SJ8NJjDcalkH7fMFl82j69sRNte68KawaoK1n9/1eJElG
pkhmqhjAl0C7wFJCI4w8FB6uOUTYMbhlQ6cZs+6/ZPG0Y164JaSY+wY/MK4JVX2l
GNbCkr3bd2LiKhDKiQgOle9jNu1Fvf3zpYHz9pVF/O/4MCEcJLc/iOIkXSIOgAfd
E4cu9HxMPM1jsyuhZF8DwNbBypXofagkQlRo22UekGYgK5qcB9v90bvoXjj/SUqk
L3rQ7v4VH3s+MPtgYbXukgA4D50GcPS8EJ4tKEkPcPPJ71ac/WS7Ejc2fnpUXymU
maf9YhH4gQir55mLsg02B0z7z/upHaNmf5gDkAnLuvydzoL+/N+egBLHfeebXRBV
c7MHGQ3/GUtVKs0jdkqDsV30DK2PNyMgv1AuNcvuKAxarqpArid8beCjrMt9lDxC
SxGrnRvPDFI+WbjOqAgZR9tuIi8YPu5oK3YxgVFzadtY/qFM1e1ig+an64ul7Q8c
nLzOkDtDJrcoVX1hnmx/L9zxTuzRHoK8s5OFDMIYHooQkKh0Z78eOezSEUT79yC7
46ld9T19UdjAEO0+Cfmh5Xq0YZQisgP8DYhOGgVhbPTd1Ku2zn624N6AzFh0a8HR
JtfVq4eRlJRn6RQXJf6UAut3gF7Y9PYXAf5aZNaGknLA0iQYFvZtNPiK0FSu2Qmj
tv+pHybtd/WmYPmispXyAqgik85fwbAWSxO8rpl2UkmKZxuykXYAf2y7iZW2Ecaf
gzqiKg6lrwK9L1cxSEJqJsZfAsQIxLt9PKRQiQRgdZy3WstRvc4DpS+yCKkZjAsz
Pp0JlRHik9YHYbiyTGGGKVvjk8Zkb1qulVgP0qlV7HRysKdj08ym6FyfiXwXITP2
Bv0fGJj5mOZba2a/afwaBYzLe6jSaK2OgrQPyDeGMLof3Q84qK2RB8VAYn7JmcwJ
gW3vJc8KsnTFPXhqt8LevLAYb6QFVa1XMfxbdE5iAEakZimyWoCbyzWTwqMRG9KV
SxmbYsm3lzNbJf+45XXqrKmDqHodVqTRAiSOliVmQukR7F0rLmo1NeVjV4okaIam
NzgxCy+/bZRcHManbDw+yL6Qym57nZ5nrqYq7ilrlsdZIJGoRZctiZhDEiPcbvNm
9UMrUb1tWKpeXuKoRpWS35wmKBHDEO5ZW/W/i6XPa5tKPemteL0puu7KFLQQ761Z
3bjsesXs7UCXWgWCtho9vlajeALh+67I5/Sm1sfjSqZV+YU9jJl8jtaPgRy1Rlck
tSvbQUw287WD4yOvSl77LgfYYDaDoaK5RjMlWcvGw2UOpi8glwk2RS6YIfLedu8y
RJgC3K7ktqaHULSDXVQxpIRphqXxzPYTECtZSVg32Ctng2Gt1Jaiu3x10cYWlIIs
XjtsZRQZS5MU/mmOqihLJOF3kpWaxl4BP4MPC/qKkHYeILu062pZluyZyL9TlUAY
rCqviGhwLgBtAz6EYI4p95lo4N05CMaNCx9Td7u5oETPwHg1lAgzY2HlYpfWx0hM
GHRYCnj733nzbM33O3XCr+aI0PkQ8v1nlWXqOepo5cIgrDOtYLzCtHqQi01Au3vj
HFszdZx35HQEdiU5rT0r74ghz8htN/bIKF7msw7mHdh+1TFN7S0RZlTrqywMH7BB
MDadyzvR2u1U0467YoH7xveW42HlziesEfI5yJwSBaNWvc3fKl7QDDc7pgI8wuGe
Popr3FleMJwFQKjAKaNWxwKGEZoVnY5mkBdrNijDWLqqJQpOsO8LGB2sD85pdL9P
TGYloo2nWwQIY4v8qLJoFv19EztMDOp2djVl3NTyWyQMC16WfFHfw0dSkBvQ8I7f
ACLBcTk0gltcUlPscVzEP3j5wxi3pNeyPP0tzf16byFCG58/oY3GbgYVTIqsHYOT
sf/fCYMTIFWRalS9tgzNr6XtoZSlyg3yQq3/JTmwoQlReBLN89UlnKxpbyupEkrp
Jq9/kpiywgRlnikMRPqPN4PZmfscs0VBPfrxJ/SVmTzle83fJ8kQ7DSN5PYjK9ur
rku2VpTSi+a/2ZsRGU6EsBTHKxtwXiXKPVObKiTsTQZpTZcCT0PMi3hpn7Po+xYi
FN0qTdfh/HQT/pZKocRiZOZC6cKE7XtQxtFNvYK8Uo1KvavpH9PQznKIVI+vCaTC
zLJcxh/qLIPrno2LSVU91q2wvBnZoYEoV1vsIfi8O1yERgZRyFlLUtWxRDp6+Qy8
gnblDqnM0Ll3Ov9iBZXJgNENDYSr0ybhgZKC3D7OiBm/vbfLNa8ZoOxim9aNRG4/
QUD2gw8pRQhXatPZ42TvlxgQ1NWh1RYj4hGpbG5Ua80UJjwLb0WulRMIwpVuFuka
nFMdWY7DXKk9nzubBD4rOTAooAmmjqQdMt4hDlI4ncJEpJqUAD10Eyxmky8PC/BI
Lemy4vI29V4bKDtCQBpq0qsxKUaRplQpqWNxUGmGvuMOx4kdyA5lpagK+r3b1yx4
WgPUk6OeZcVoZ+xoU0xl4BAR3dAU6ML7tYqYeBxLiqvdNLiIW1BiHn2sunxbgMbY
tW7or/U29W8wsEr79ZsbRpsACvehO0dOlkQJetzBlFkjVDF5mXpk1ONJJl6iM3KY
aUFU7R16DWHOrKP3p7dxcu+j5MXQlWFb2yXYVK4VyWbYZXm1BAOo4xINNdF+9Kix
BIRpTtOHSmGpAlC/6BuCmEbpU7yIlbt4+NhyGxYx1La/f6tcjbpCT7jwvT79sT59
4nNXhOfWrBC7H2prEe8qLk+sxUNtWKKsI0WuI31LcYZQUBFRjRKadnyOvbCYECbD
Dp9qf7io6vpc+Y36XPnxUSxjf1imYYoXk9h6NtQuowXb7WnW6j1fGUzToP74UPoO
O/N4hu3VxYtYAodG1PTXIOJXYlNLxH2VQE9FC+6SLxNScl+6w6xVKW6jE6ThnlRG
r1wC5fWO1zb6xELbiBu3bTxzVGNC6A1Y6fjac61wPzSKDL9FtbZOtrzips2j124A
FUYtsjNEACS8HKZlKlbixMti0EyPnbRC5M9IDoIZVG++E7db7hiPu5lWVZSn1v9z
YoQMkCnei8es8c1sqW0IQ0KUTx6Hakbpes9zwfqyOG1ymh4oVghCoubbyFOAjoTS
AgDzHAqwkoOXk0b39/E1oFEgGlwSaC+YV8bP05G7j22b9+xSgRPb7YBdHvrOVgkt
s5WRJub8YHEMaUPp2SJsC2t1iFRWy8UZD34lywOzNUpSNtLHaVI1cv14xBEPOz9t
AFwdf4C+7siUcc8SPonvPMU5KB7KA/1H/3R9MCw2wPh0Gr484rXspi5CbLDWlh0y
7GsyP/CboZ3/f/Mdp8fMEisF8uk9sBJU9AY4TdBoXVI23CAjs20TkgD07ohIPmFr
TmH+Ay7dhP+7rYUC1EIlla9LGws0X65DXyIuv2DpnV+5nTBaLOggstavIfNy2VBJ
2NJ/nG40XukGcOA/+dgDpBn394LQ/7zpT2n4m940ULVHoCMZZ7lT+ODzW45TlmUA
MW7JuNt7WummwdHjxAjBtE10TruZxKsd5L9cKrzHPcwLNnl94NnbYUeGwIk2Ui64
6Wid5dpw7pNCfDImPnbW/h08WXnaIpfUNyXldk9FhNt0V1+hI9oX24Pxk2XDJbn3
ezuzd2mYY2TeS1z6pMB/uTS19xw+5T7Dm/z/mRq8bRPhXzqfWARo8jvda+011g5Q
jRQBLXiWBBaA4RS+vWBoxLeDHG6iA55NEafwkq02p06Gy5w97sCtWTACIss27Phw
0/LOZefpLRFM6Gp4A7kWW71PdKzKKlWV77PR2wxVYiJmRcKuwYj+/00dZBoNrjru
TkvDDJeAi0BZqj0zIQNTAJNnakcv16hVmPniUqE0d1u6yBYGHVY+3fPvKbpueP6o
EvRXS8wL2iMjM2mQTOQXVa48AyJrcnRaCFg0gdTl8ScXd5hbCa5d8Vl6uHInrEot
lkBNlQS0DOgCQoOE7c4hk3LzlHTDEz7bNtfy7wHLMK2CWNN/UdHA0TxQuw0iO/TF
H+6OPAQmCBvM56KhtRHQKUmZbAnuEBTbUB44xUQ0zoPLBqa1SbjwijCRCQOm/Sbx
dXIZYm9efOIMoM4mGq81KoAOucWh8L60TDoyuMF/mQrvFzxIuGpsEFvbbz0tk0AQ
u/nXSc6wwYB5Xw1JibzzKOXBhTePic4U2tmfOcgqAiqeP7JqPt+/euVpUt6vK7JJ
s4fUeQF9bCrwaAKf6XkghC0MXPq1qZ1cqcnayeEOMIcaE3reXXOfd0TPw3ul15ay
oVpAPZLUNqN12ym8ipEwvw0vJGYCJJiETE18AmVv7ubYblPkj2qbvrE2fV4F5k9m
/7qavcCXv2xPojbkC1TG6RD2Y3LOSTRIR0UKTs4Yxbc9QvxHtOpSUrCKXVxtTJRY
XwMJPTzMbSHdG79ZyfNbGNUVIEI467PFWuBgl9E3dP83IyD0OsyEvb9yq/JbO+J3
PUbo+CkX9RYsyA99Cl2QL8Gck5q3iB7c8ftMXuPfyxmAc/AZloo/wnGpFXvDw1Jp
KO+t/c046XtdQcoipxQifqlU6u/Q9YVYbYNaPehiACYnSoDF9e1ATQffDFuBlQ9y
T4BBwPSRLT2S/CwNjK+NWjvvRk+VLQ9nb/mbTi/GemofCpv4G0Pm3uTkZy3pRrDY
xPw+qpabc5hfIQFHRIuGTw0VFRaMoZXZuRT+npPFwJF4Kd6SfmV7ABe76fx4vo7o
SP7lyNX4uW2qdYE+f4vxmoFfmDHH3oWtCIm/WjSHLLuD4dSy58FwxNooOv3fzSEd
hF3RuMSfgwchDYzZRB3tdV/GTF1uNhS2vp+HKA9U4aTJLAeHnhMBxcYPkTniv5UM
8HoZcglb5DT297LAlT+YLYXOGvtjrSjHk6gqQd/6ktIkq4SpO9y6ikGaBI75PmR9
Y3fVbUs/jHoQ++slrJZvSbR+37GizLju/aMJzv4RwjjsUQ7xqqcHaWb5vv/ha/xV
ovy/gbEGJnzrQTl94lQ3doNmbjw5n6QEm6dkJ4OzDXtOO8iVIc0Kjq7EJv38uJhH
QWfwe5aSw9X2FT0ATguG96a1N1R/5y1wLw5txqrKUStnrivyNmC1VV0J/4aEDR0s
HD2nvvDyC2RXBRM0D/85+FCni/dRWc5R+IfLYjzu/a+ACEgQjTdF5HMdPkb8uFdk
cxbluqxCry9Ulk/bvmjc1R/zhfcc3cpOAHp3BEbTN54t9/JTpjR28++TnyBWD9Ir
XALUoMfr2QBqLSFoct09UE6yTLvLsii72eLUEZLRSJp1ZzpJKuMsCO2bl0M5DEqc
MOoVOwZ++TddOTVLZWCb72ms8D4/pr5sO9rvuuf10kzK7ne2qdEv3ODw+9/lkRzC
ZYi5jx6RXmV4lNPEz3qx50ZcLGY+3iOo6TBo4jeAiJ6dHggMy2hF10lQmFOZWzZt
n0d1p9x3Ov41+0Ob4RwI8uOJe4SKxBmcQXXBM4H8OoYNFKbeQBtslvUQoSjA/sKA
wnob6qg9PxJw+iCu4rD07H2dwbpWPIklMwN5zk9j/gFBTflvQrdQwmVkpxY3y9Lf
wS6nyhol98/fr75Ew4eZCQ6E4c9q5vgKAGnW8z0Z9qOOtPbHtachOjGqUzq8o/JN
rb3G14LwybNIn5/Ko5Uff16oY0xp9gaKYEyslxvIadbvyTaad2S1uD8g9iVpOnfr
foi9qobmA2CizKNNwf01WNpG0l4kJoLcZSnN/hTvOEsyy7nEx6XqjPWlwDSSX2gf
OxIt9SRY7bKO/WUiOxQvGR55Dq7wSxn/DVxDJeyxNIzbTDl0FUMv/d6mkN0N15Pu
plHZr+VHb2Zc+Uj1JnUHaEpdDBezeb3oc5d9cJoTRJMExGdWm4ykHUbBjMtCxUHi
CJymXAQ6pWiZqGXyBC+4qdONeUe+z4bRbY3OAkLa6TTtyqTJlMc/EobaCjTDk3Nx
qWnyhUeQu9msveX5PGCYYaQ5ARW47pGZbUAtQisV1SKt3PcolqR05GWzqHJPc0gF
TRnwmdgAM5aCvvkKLEHCa7wMyYXqLO8jmuY4EJ9VLJXDBFCL9t0JIcgbjGO/Hu/M
/nlettp/7GtAWjVJ366o2Z7Ke2RTzLU+PXgUqh6Aj8MAK+7ON6wyRPhXpbzQFxyH
2W7wZJNmD72WWla1sfOOnhXaEFRxxrtVB3ZDCjSXF87lJwhWd6T57Vbk1ZpEhARi
xE3XwnsAdxZHhfE1yc+5KJJ7xOTQag0kbUIWKLhDw880DO2NtYXrCX3fMfTwS1Hf
c2C1WVYNGS/aHQFjNjl+XEegoOSCOtXnwMjDmxLmPyDubSZD5AN9rgxHodifTc5S
fyx/K29Mzm6+TsG63vSM9+XQrIqleCc0XNg2hZkVoBEHiuR12LAUNBLsRuJr7wVq
BFktxZayXW81FEG3egbzuF1n3tm3iDtH0y3rMj4qGQ77Iv8SMlBzjEvI9baNmW1W
iQojInCUUXlZUb98Wk4kocvuwo4UBnmbGulmn03xPrBfJRTUKFt6eF6OVS/Xn89s
0T87kEdJOrXvuKaHGae15bZylHQ/qpKc8Y9krVQdURqCHqZ3LWtRh5vsCQmPVOj3
dDDQTq88/lijpZhkbhrNgkTRezf7YrM8BaJlGApjlC7FKImRdrG1SqISQf2hzrs2
nzT81LCgFkkcmFDm65NoeEU12wqykv7qtzhMhUNX0XZ2Oz3n1ifF0GLgh0IQeVHa
7p/b8AzIjByP0LTN+n+7tVirlSMdl8ZEEUGOL+rd1F3DnZt5c5Z+NZ/+61kwSILX
zFWYUTPx6JX27icV/zgiYM2jkwsWJXSBo72dLoV6TJCKpsFV/SVuJ8Z/IFvEAHTB
ZPAnz07nf2bK5p8tKCKKxj8dXIDjj9Qssgxh6EC199sUs5rtLGzTqrPwIWycB2DC
FO2Ebn46RSCynAIj7J5x1Hrw3EV047KQd2ZFzPgRl5C6SCVSpLMo55gJ85tfBqWZ
U9ALb5+4qT+HO+QrOrBXgkI90itPUUoGuUGxK07sN004Eh+jfOMrWA49wG+AqHuM
qkSDUHSsUYZYJtpqZuwic6gDvczmBgejhEYscHJ7X+f96PLUWmSnDuTBrwKYwdGV
1IrCDIMUd7jLpS56FeyVEYFJg7gU/UbesDOxwv+yI7OXpBwa+30x2nhdMbaOyFZ9
zK0dq06ZR/MH9fVaqn2ocG2LsFFS24/5WVU4oqYS3WfNQHmCRVc0kLkOSFvzK7Gw
VzDefAA6YUmEGEG+bw4DZX7p8274Ie+W0t6FNDTPJCRM66Yu18Z0pOpn7RqucSKk
LZPYJZhB6DSsCSWrGAXwG3IbPPTjZTvHuJq6ms/53qUDZnbBdYyZDHJ9qWLiC4+w
fBDhiXdreJyufCicrzj1lfRK2a/Qg0oGKX3OcVdB7OOvkzvtBIz/3LZT3RbAN4gC
STN3XeNEoCQRn9iJnesgGGiITrO8OK4UYBi3ki5aqN2bvvyKY5lPnXK043Thb/cy
vGWBA8AMLKb3n/CaeHNMOPYogjw9+w52bYmLq+GVTwtghHq+QjpJwnC5qREx+dDo
gOS1VrzTA/Z+gvmZFGwKgQyuBkQ6aUCP54Zs+ZQTDklX40e5fIw/Mot96MSs9IB6
/7bKOp4Bq4/mjApIcW8NZpVQG+FIGmIqjMvU3eFXu8QM4VFLaXBbasb9ovmNH2qp
DVAUflnWxqebt+GkH7iy+zncP9ew87XEC7g+yxZPeczR8nuFijmOaYbtZA7F7z2H
jOFHdsCiDKY5xR4JJXCA5cSRlUf9ZrVMImidb+rKy/Sog8zXDKcLHDW/9iFaylZw
b1tnLpV3BB40aylE7Qu7fTSPsbbRgiOiVEnIb71NZJ0tzswmwld8DZTfzmt5sGO+
csPyOxhsQR8T8sUI2VFUn3XVa7AtGWNLBRM1UhprnY6lxtAvRPpU0D9FBco8odsx
9gy0WY8URNs36ZWLVIp9kHhwJGXUB5nhyeOHrSj3W8l8xNBouuBBQyn4BY++Mc3i
F15V7yZaHRe6XMAldshqFRd1Xwl/BTyX0d4txBvGSDrMFJDrDn0LwFiOr4tntdJB
iPAY1licI0ECcoT7+90DTt4QrV/ULFc7GqUeRow0PYowmghs7rwLzfw5nbHVnQF3
z6VYrgXZfirESMsoEFuii1WGDysBNN13k/+kJFsfGz2joq/onUqJzOMzYBlzOhTV
+zhzFYQv8If2URED2yJHpnObJYMQKfOazAZpcZkgpaOUoCXnN8bwTTMUhYpVYiN5
38rn5vuYRUY2qafeA3ciRt8AIp7n8qyupJYkN2o2K/T+HWrqBU1GBYrrujSEcNAN
ykizws/1WD9NBXHCajQp7lXQS9KG0lyboTW3wb/G0nden+7V8ik1+oOHBqDJzkEQ
IgA4OgXP49a7PYuXEtamrGO89PRu9EwuPcIVj4wy9TaTy8gElckNiWUtNZHUH3b4
uc9qPhrgbDND+SqCsH2RWLwoRp0K287UkEHpYyKwZOBF0EBP0AV1lO2u10PX2EIK
NquRm8CbxAQbyYfk8B5YnhvM4/z1/HpnOPW1kxtGxrqONsvnItKrZXXz9XRa56O1
T91SCCm0lgn/WSj3KDp9bsHVVFM8gWZOq2AoNwmoEBTGTrMpyqzbSEfsO4IAVcFB
Nia/Td4sQMXhmT8Stxv6Xa9gVcmcNoT85tY1sffbQ8RFlhwvcVgKCGzcb+9gZ5LJ
64Mpdt1kC6mWrbWL/h7CtZRuXmYktjbr6/vwgDIo94eW4NFOIwy/c5WCabfYQaEY
/DMYr4lMnWJNPnnijcLVRnLQ6GZ802Z+TfPO0drEn08/2/26rLLOwWe9iuXazqRV
P3x4k7MNBbM1p9ke5t3CHg3n9VwiWXxwJC6x9oKu2EZu+81ZKgryWRBmoVvRmd83
BbPGb23TVUJywo64hf1VNUXEMi2PY/BbGpYJv7MZkAztsOsXw51N2uF54oLZ5p9r
sHJhTKFrBArK2ZpD1ot+Kbsh0qUEmQ/gMRb2w4oJ5VMMd7nARNvrL7NXE/3Xq4eH
Eki3vXqlaKrDwz6L/tgzxaov4/zbtPaEUXuVYQSN30s06dIeNfYN21u9gQlwiGV0
tjjWIgVnh99E4U1jeDvNqk7cKbv5X0qoyaolJAptl9HJWTyVBfrr6CeM4kzWNwC8
M0XxNW3soKLGfRohm2PqKTTpqw50NTHbwZOE161usRo=
`pragma protect end_protected
