��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-�1�M��[�
fL��l��ߛL4��v����Se������;\�$�u�I�z'<�%�'N�$��� <�a]��֨7I�������7�͕-EӱZY����:іg9�{0D,��u�.j�-{����
W#�8Gs�1(`U��2	�����E����1u3�:�nBk�������A�3lf�0����giPC��z�P{ov�Q������U>�O^�-?���*3W$�����k������fG��T�`xrJ.��Gl��[u�|+t���z2�3�*![���8i��?����@}���F���H ����J&�����e�	F�����yR����O�@\�(f^HR�zTo5jT�N<�T~�{ؽ���15�4�k𬅘��c� ZH�Ny|�	�N�����>�o�q�gح)$xFٚՓ�+9��v����:?W�O��;�G���Y>�-�m�7�9Y�hԡZ�$�����oP�.&7���✖۫�9�a翫�f��b���r
Q���8T�$XK�W-^�IQّ���_c?���3?-	�toꇕ.��P���˚�3J��啝���L�6�L�0�d"�����cj�2��ƪ�*� �cI~�����&|���$<��,���m"݉�AA2�
���ҧL�4c��X���)�#�j�w&�S<Bz���#ȓ��1k��q�Euo�o�����	0�9��)O�|��j.�����3~�]�qN�6kH�f;n`([�mdZZN��J��ޟH]�x�S��O!���9�T����L+���=�EPd�+&�`]�i8V��s��������#���R<o�� |as��Ш 5��/}� .��>�A���B��%�����χ�m��te��L*�Y���	�|f'��^I���S8��F��OoZ~��.Y7�] {�/v�d+N����}���P���
0�FGĳ��5�7����Z# �k��9��&'����_��PZ	���h�9H�g���C�]�+x�� �I5C9P���[�wU5�eՎ�	���B4��F�Il����f|�yYY^�� 37����$�n�l���*%�8��w�R+��y��z��PI�!Uď�W'��˫�]JW�]�x9R	Kc��p�3n�T��2PQ�_��_û�|��T��Y���}~���󮉫��
.�nF���&ǭ�`�+&����4Q5Qz�n]��<Ǿ����ba��TՔ��S���F�3�]����U��Y�r9�-�55%�{�6D`ˠ����m`5G����7�u�dWe���(cǦ�䉙Y�C<kE-X���8������=�^��(rPҗz%�Y(s���$]G٢�D�d�8��WO&�zP8��WV����m�3��h�ge�sJ�w��B5�*TrR<���-K>��_�׀��/2�d��p�c��=J�a�:�c:r��X)N�㹝5פ�&Ӂ�t� ��5!��*�LF��IڹX����0*�>�9�O2��YDh��vlѓ��� O#i���U��|��/�� +O�Q��(U��˔�o~��B���	�,��_Uq��s@X����Z��T�{�FqZZ��_�z����&�9~~�Y�x�(>5"%z_�zv=�n|�!?Z��吮_R���o�b� �
¨ڻ2,����?�M0�Iތ��xGJ��E�;��]�%�b����WS�SJ6]�B���,-;l��#=�ŏ��|�X/���р�>,Ī,4��t
ƞ�[1и��@��#%�3���pC��!f�v�;�~�5��_G� Nۥ��ћ�������L��o@��(�>�dd�EDV��1��MK��� ���&P��k�+ �2PL)h�o�+Bu�7E/�^4w��xV���%��L����乪��BY􄻴�� �2d��L��d2�s۵��ak��#+�v�e�QI--Yx�İV��N�~��㕆M���*�~��·9�:vY2cj��2�;%���{ӯ ,<ߌ�RT9��%V��~#m)>����ۯf�����gc�>Dس�%JlN�M�в����
?f���F Lʈ�rw�K�r�����"E�g%���Es(��3�_s�د�;8E2�((�v�z�$6�};��$FQ� �n�5��Q��|֚��3R�{�U�7���u�\*����������8��z'P1��E�n^Z$�{jd	w1����j81�o61K?�-�K�ņ��?�C��Q��L2��7"��)<c���2ql7y)�����/R�`�>%v+��KrI��H�#It4�'ԁ]�Fb9ϱLMz��#P��)	��/ q^��="���P>�:���]��q�	�.r3���^�Gq��*YL�G0,�0T����J&Xw�����m�8��XUE�(|��'�>�M	�s����]���!.6��)Jt
��c��ﵟ4y��~��� �(���e��r����(�:�q�0�_~���t��yY���= �+3���w�F�"[��%��Y5̒�s��"�nՎ�vC��jdi�Lq��,qiQ�q��׉�.�� �?(��m�Pi��w<��w�`atr���Ƒ,��r�hh�w�����$�����b��^`zw�Hu=��LA]���q %�Bx�i�bv��[�������Y���V��g��n� "
+o��؟����v���ϲ����^-��yH�.��?ߗ)�w]��<Z�ǒw��w]x.�>��/�l� ԭ��J) o؆�_�5�&��I��ہJƂ�ސ>N;	�1��
a�d4CA$���$�Lrg6
�& ��
�O�8��0���� F��H���$�63���nS����t�U	���G)��E�Dkf4�o``p[�bR�TZ
*��H�����U"���/�x����!r��x�ma��������O7���n@�QO�ŵ����?b�ciq�� m�ܧ���S]��V�4Nl���@Fܰ�[��M���M\l�x��p6j�#\ET�v"�l�[%.�L� Z� ��D���5�����b�5hK����L䫼�SQ�B�#�	��^�r ̌�Q}ˊR2xʚ.�<d�����B���p�G���E�K���m:�>����t
�y``�+�`Jj�
��[4�D]����(� n�p�j8�>޾���p�]Q���YJ��S\��5�^v�i��n�_�l�	�#d�(3RF�]�UIyq���ɮN�Դ84��,��$�!ʺ \;�J����.gz�$�6qZ~�ؠ�� C�D��ݬ�*h��H!���f�3a��t?�_h���Pْ�Lvo�徦N=���L���$���:=��NE+ńt�:��|�i��?�O�hlK�s*��!X�GU�k;�Է�/P���+�vM�C�� ��q�d�����]�������ǎ�a�j��B��`z���;y����'�{O���!�$�N3���S��h�P�Ou>�`��,w��4$�#Tdꍶa�ˑ��,�m���eo׏�с!�ߊ;�Ds� �r{�`&�'�+MR6�e	r��� ���~�tTm�v���t��h�h�ז��-��`� ��3��������������c>g���AW�SS�%I��ֹ�thq�S�3U��e��b�	~�u-o���C�s��+(��\{��|ڀ�?��ӥ�t�nP���Ⓐ��ˣ��|�^������������>��rD�F,W��}@-J���.ܳH�ΎK�5�}^�R:�2re�������=�
#�YU���Үf�������T�<�*'=��]���P8>�!:�y��9�]J�����(e��_�r����͑��b��=�����fI��LYka2Ƶo$��[
��}wQ-�{�1�x��0�����!@Ν�� �G�*�gd]���m D}mS�S�O�XeM/�_�f[�����r1����M�µ玬@� �!
�;=b�n�AC	��$�����-�t�#p���<3F6�\�֗dR~��Po��[�� �F������Ǉ4��������G����H���E����7�����(9���@��`�#d�
�g&�&�6ߢ�/I�o�����=�F�چ�ȥ�0·��ʋ�*aq�k��y[�9�x�Z���!
Fl��GrGl�,����_`}"Hĥ��Aw�ykXTF��y�+�k t2�4٭��q���1�c-8��Q F+��j���Qt`�~���{���`vk1�$Ԁ�z�yuϰ�o�