��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cqL �$��).y5�´Ik����o�2|�0棷l_�������.���|U8[�j��r8AJb�A	;�q�$t�ٷ8�j��R$%�jυO��(G�q'Pvgˉ".�!|����=)��
�po�7�j�"��a�X__|��+k��s��Cuג��ِ���V����ǲ�-
�#�ե�1[f��gR��(�{^L�WPhwF��pِ_��&X�DXFL}I�?2�n��v�C�8��4~D�	ì�8	 �m�WT�h:�}O`��v���ֵ(���n�Q���v�����ws�����yv�fv=N���&���w���*�`1^RX:��a��b=kC�����a����h��dj�^������W��n��=���E���|�ab �9;[��Ǌ'���s�e��+*����?�l�b�3QK6�k�pޚ��#��;���5�Tb:ǻ�ɔ	ݺH�q�~��/}��U�#�\Fb��C�^�T���N��������M��m���cX^*`ˀ�Vv�����/yE��s���*������F��1K�f��|D��^H���*YJ�N)���$�bq!�Ga<��=��7�[(W�zQ�G)��`e�Tu�2�mR�������:������1�J������8�Aϓt�غU�����>l���#Պ��v'O%#Y��n.�����L9�=������ ��5�F�� #Xl�;�T���w2��PY�'��w������\'����r��%"�5H�7��޸N��g~�Ij����˨�l3�_�V\F����u�˿5>w͝_�j���MiM���q��<<L�wd0<b7Ľ�)� 
�zbY�w�_F�p���!X�(���9�����ޣ��PQ+2��9��ح��*G�i�m&���ֈ-5Jں1kC�4��u'�M	J�F�kUS�)i�JȈ$��B�z-����^�X�@~�S�R��O��Xc�{V�����R7�u����|�������)4`O7�b`ʮ�k�w��g^2r�^��U�O�.�
�K��H��d7�6T��
톥�����A��_�}|���Z3�]A7�h�-�r��w��t��^4�+�x3�?G��&��xު��%���4OL�v��$0\�KAۯ!�a7�p�+�q�d(�M��j����WV���[}���!�"o4��O�]�v4�S�MF�vj�������H���5��}�������թ>?fv��'��}}����9pq�r���r1W�g+N���ԑO :<'�<�� >c�9���%W�j�'4������mv!ްs�Ӱ��nX�C���4l�BO�Z�b�^p��~�.�08�T���"��?��#�R����r4�K%=$gc�&1��M����~��ł��w�8�BU�d�C��+S����=�zs~��8�2���H�{h�4=���97����
N�9�<��;�?��䃧��5N�~���X-zLn�����$B���]�F����D�:)t�#��R`�_�F�m�E)'}��;��nY�Y:{�����j���h����jt*F^s�%=��{dPa�-���f�P?�(�i�bިY�d�g�@"�j�k����N�q$���E#Ecy ���}B)u@�?,mIۗ��<6�U����(�ú���7G�b\ʁ*Ss��{�9X�qE�g�0�1�8E�U�7�x�!";A	�Q[�5UT��� �jT��y��YR�w����"�+_�p� ��򣢙��E���8�����Qlq�6Qo���O֘�����(�l��#NI.,�����'f��@=�#J��.�����u�\���R0	��j���w͑�b3�����@�z�C����^Z�Z��xh���H��k��.�[Yn��ƌ>��U�X�.��.AoF�d2�3��K�Б�6l<L�s�pE Ԅ�����8�ur�*m{.6����/���=����6��:#vkUl7Ur;܁��t����3���W�i��l�_�0��p}�W[N1Uh�|���I1Dd�;����9�"E4���69���O����!'s>����.��+3�D��S�^t��IK��o`�&" {2���
;�oD#b�f3�8�z_O��� ���1nSm�#Q@�A]�-�<*�իI��s��P��9�#��.�_#�MyƸ	S���+���O*�G.<�tUqN �QI�|���?]��.�Ѭ�ۊ�e]��Lf���jشÑ�ޝ8^������#�×�ץ�0nqzC�Sr��l�	�X�����R�9v��3 ,t��j���)-;��$�A˧��p��w�ą	xj\�튍1#OAE�X�)����0���4��1!V'�1`�:d;��9�̩�DV/=u��R�~�=��o䝲fڨ���L�wy�	���G��J%�]�b=���h��I^�O��6#_[q�~�ť	c�qwꨧ@F�\>��?I�+&�;��^c�T����n$A��g�!���)��ֲz����aˡ�4��(�R$@և��y�MOp�|{�f*R7�pw�MwΪȮ31h>%+�i�����F�n� L�H��1A��W,�D�s�kPT�Q�+i�։Sv�&[�{��>���uCS�N������ǌ�L�M�E���m��L�Y4���vj���������M��%���
���}�FL�,{��+��,C��t2��i>�����~���8�}nx0pġH�l��?o +us�*�mxf��'� �'���坆��v�0�[����C�Sm �(Hq2q��z����_�z4]�Dr`��TK~�9���]��Ѻ
��9��C���LQ�@����4�0����:H4u�9Y�a�)m^����u�ViE,_!Kݗ�'��DZ�Md���{�:'���5'�i���j����|��G��7��]�ΗA~Dg�X�V~���0$��4N��������<�.mk$lR���l囀^d�1��ؓE~�*h�����L���=����ta���NZ�/08�r/�Dc��S::��5$NJ(#�PqgRǋ�~Fx:��p�h��,;ű0�#5m�_=����d�zK�gމ�TVDm����E�tu'Ԥ�'U���~��0���=7���p�!�605hێ����ZC��/Y��,��؅g�!-C��C�Z�Ǒ-x����w<�|s뚣��[fTP����t���H�˘�=���вbN�zqN2^@�L�f���Zd���!q�75K����3"�Ǵ}���'�G��7t)��>cq��2�\ɳ��C-�V���>����ڗb���5Ԝx�oK���Wr��|�\���_&��@���m}#gYc�`!��gY&�/�{[�iw��'m#ӿ~Gl"L��ȝ�� ��W/TY;{'|G�	�����+sTo��3Bf��n@����`��f���([
n6��
�J�J�P��Ҿ$eec^�/�hu_�[l�|��h�x��\C)�n�T`�M���{�(���f���D2���U���� ��D�T��������7mYMR2*��<�ᦘ���������� <ǣBnz���:��VT�;�%���Mۑ%�Fu&��W3�-��~��>��*�����<�E�ob@F����_>�������J�>��Vq�`�i��,>��ʼ��~�g���p��d��C�~ȢS�֣�CS����=2�k��N��	�0 Ã�ȌxEH؞�����3?���� KL�)F���ɖ�M�JW�A��Wҙ~��[V�.LW�X%?��@�c.Ͱ=@���5�R[��l��ܻ~� ���\q���;���Hj�ڿ�� M��������5�ވhb�j�����Q���G��/>0蒁}<���4���GXL�uܴ����8�Z�2 X���=pi�KRn�4��Ce�2���d,��H�-��97��ѯI*����kҽp�͵޴���&Nf�|)Lm)����%9˷���E
k9����Q�A����1}�6�BK+{ntM��db)��ߙX�:�\H���%�	�Z�H���A����֚�{EH�4c�nG�kl�5����Uc�]Q4g�(c�b���]���؛����Շ,�������s�̫����F�O���+�i��V5e>2�b�ϵ��Oܱ#\ZY}l����� V�F�N7�Q�����߀*�TQ�fu?�q����J�?���{A�rF_A��33�}�!��׷��Bx�.�$�f�<q�m󭙑Z�N������x�Ƌ9Z��dD �GaD�1w��;{�(�й.�?w��g���7C�M��N��%��"p�`ßm%�VM	��y�"���u9av��Ƙ�˹�<T�j���Zܠ��`d��R�<�����/B�wz8�c���=��VU�����`ҟ��S
U�d�

���`�J�;$�#]�w�/�h�����?�&�]���fB�c�A��� ����W�g�Ʀ�w#��sKâ�
�y�*`�����шȪ�ة�hS�e5k�,�����Y�4t�`�+_ی���U�eK-���e���zs	V��9?��b���͆^�8�M��H��S�����O��a�Xѯ�����u����7&a���-�����e���O���2yN�-�7�����O���h�\]_�aW����~��>vSg&S��07�}���@�5�R歕[/൑Ǎ3�qV���mq�7�i@���2�Cl9(!�D���0���%�5{O�Uf��m��sWb/����Q����T-�A�v㓨1�VO��]a9��DZ�Co^:�ouE�Ɩl?��0(|��-Š�~�E��)&�1y��je�	P`�^ ��g�K�h�r�=+��n/~�P��酏�'_K�5����$��} ���ܹ��/��������϶�43n�0�a�`^���qe��R#��h*;=��v�3��(xE���xP_�D���F�b��H{��C[U�WqZ��3\ۏ�����^ �#���k
�/"8v���?$��M�z$����`e���k!�<S�LZ��3�D
��0+I���*4I�ū�LNg�Z$	��_�!��(B�( ���g&��z? ��]ު�:��O