��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���q��՛������@�oa�R��Iz1A�#`�ԀP��Iqh�3��F�`�ҥ����c�
K4#����ge��T5��G�z�4��R��\3jU�;Ѫ.Xq��d���D��nmac��V�ܕ�;�)=�(?0�י+�k�襮=�%�YO������鏷w��>�s]��6�t�u�;]��4���!����q��
1�xF!b������.����\�2�X���`���~���4�k2Y�a�w�7=�E�u��#��_f�g�:�S|.�� �֞/^���J���,\*��p�#�0k�|
]c(��7��ȩ�'�Q�	�kR-`~���Zk8�$'��x��A1����Ko�� _'-l_���\��
+*�q�k�����V�LZ\?rŮ5�xwpP�V�22m��w�j�{!��;�Fs����]U�ӂt0���΃w旫�u�)�ު�z��_�s���w%���0����҉
2�W�e	�u��9�P��-���
��m��ȈR��?N��Ir@2!��1N.���Ф�����_"v3h�K��-f���X��w;�N�-K��S��0�ΧY�[5��V�g�����ֶ!0��(��x�����)�^��ٟ0\V�x �u?�@8d %#���6�o�B��A =3�i�jT7��!9Ig@�?t��C�5إ��	�c�����m�C�+�>%"�W�j�J$��w)e�YjeR���½��xJÈ����蒐r5�Z���C�c5�	�-!)�S&k#H��GwEdOuuwF���E61������~��N���G���m�g� �V�]��:c��!=� 8��-4i��B@j��u�3�� <%V'�|��k��2��y��-l�l{�P��=�9�_���Ǵ�J�m�M1m��;�!{RaDb��m��Ԟ��p��n��A�{�7�\jߑ~~.��y*�YGBҼ '�W��5�y@���M�&�͜�Y�S��]䀩m6͜�6���?u5��
�����G��k=�!C	�`�$JL�e��ӑ�V늰��Y�xo���;D�л�2����1|6�ь��K$
���
��ꒉ�o��z�a���Lj��� �OF��ŀ`#s����j�L��H]�����G�C�E�/}P�Փ�t[�>��Ĳ�[Od�i�i�~���3�:7nK���:�����'�}zs�|�|��כ��y�c !��x�OT�dj�t"���=T�9:%�����V]
��[W�:`<�����S[Pyb�:���?Gm�w�&ې����ܢ�D��Ñ���;y�Ȑ#��d+4u�����L��K�ss��,7�L��GU0�?Kzݣ���
傆]�+YO���I@�����Zjq ��f?� 9�2vJX]oaN,�����Y�����������xz�u&�-��2)Ǧ��,��Jv�>��,L�X�5���Y& =w$(�u�g7�F�S���8C��\[����U��Q��S��y�������*$��R��	-�����&ɰj,th��N-[�b�$˭f�F}U����3��{e:�%F�����R�<`5��3��+�^�c:˔����qD#++�)U0&���'h�|pt$|I#��ad-sV��-o�ƅ�Ŀ�Լ]����
L݃GD�Ao��5H��1XqR�P���Q�L��pCI���L!�E!'��x��L��8Q0���U�q	d�9��ώ`eǢ�%�j�h�]��ɟfK����(�h%>��8|W���jV��Jqb�97,ǣ���� :w�YrCo,��J�X���֑/�؁�}���À�stV]�aL�G�ڱ����Dq2W���҆�S������-(\ʈ�zrՒ2ՙ�+t��;�|���52o��Յ%g�e����!�G�4R:u9w����2qS���3� ��9��k�!������m�e$�э��n�-nlE�۱��gI�>���=�&����|,��Y��k��;;�������"ɭS�v�W��w[����l�}��R]���S6a�߅u.f
�����`�#��JL=f�t����Iς�b�*C �D�Z�|�a�	R<02��G�j������/��tUp7S5�d����������!� m�ȴ�O�ne�g[h]`ɳ	�_���OH6!�E�|W�j-�ф�a%�i��p��-sJ�B�;�+$��x�]��+����9�E.}����OT�,Z�Y(��������r@������(j�sƤMqۥ��cQ��!6�mS;߫��B����%�h)���4���㣍����1�����ס��X0u�k2�lr�obX^�i�"������55�ƙ�D|��}��9S�bn��N.�Z�]�$k}���-������ONb@]i�EíM7�"�h��߀��*�)�Y��t?���<���vK�I���W�D�ޜ i&�j��>s�Y6�R����Y��߲��x�V�
+�:?=FMw�n]q�g�a�JJ(�����0�	�]�V�'�
��YXU��i��>��W��=o��(���=-�y4�9��A�'hT��H	���1Yw���¬p$�F�5���|ߜ�� �����S�?����Mxv���
%x�V���MnS�p���5�]�y\�6�Ti��PzfB0���w�C���*��>��IKA����I��~�0�O�;f~�ٲ��Z�Ô"'�k�{�-�6ިKRE����Z3�$�:����܍�vɫ� �Kc>-z�Kv1�;�YnH�
��<�����<�(�z���$h����Q$]7��"rP��j�H�Mn�U���������R�R�߉� ل���##A8W`�c��
y,�#����&r��)?�{�`�>���~�a�O������X�����ӑS�CI�z�x!�i���΃J��i�a�����N���湃!��ԊG��w��䣸��N䬵�z]�5ҹ��pu��iz
q.�	D�@��<|� ��6�X➆���=C-�"�=���w�h������^�cBn��	��]-��M�Cr�*�xb�D|�Á6�w��Y<E���N*��	���A�K�騟>X���w����+Y}z�('>�b�����j�ObAԑ��4�y6�\�פX�*\�`m|�:؏�a$���TF��}���\�����tp��+�
&ۓ_H��K7�\T�~��+��(�S�(3�S5���4ys��j:�;��R��Cթ��fF����t�	������C����w�����ш�Z��X�d�8�����f�?��؉�~L��̰�X��o�jX��ۓ�'����.[ �ҏ�����U�:����j��y��1�s�
?L�e[
��^;��}aY�JW�e��j66+P�V�z8	�
}!h�bY���CA�����3��@�Ҳ'Q�*f�_����*Z]��G�����`��<�?���I��������\Ϻ��U�)Z&��k�dt���^ >x�2��W �� u����Cā�F�!k���OT�\Hݡ�p�a�R�IZ���o��;�ۙ�q:�B�
����w��L!|��ב<3�����7a4���d�׃�̈cd�L?���S��r��2D��L�^EO����o70r��G~���{i�\k�c����K�-�$����P�jػܩdWjv�)io,&�����䊯��T\�q՝�6��C�����񰔰C�5��?�u����.�m3�^^�^*��t!;��HV��#�!Z��N� ;�ڥ8h��كӋ8�V����[?��M�r|���gߐ����v�߽����6A9´��6WZV���S��l��;�1����~<����8���(E*�2����n�\'�b�wN�\���EZ��A�6��$#m*��ĶA��	P����j��<�	��%b�o{\�H�����Ƶ��G1������Ud�M=��{%C�8�����( �Z��>Ę�S*^��Р% ��K�ao֊�JP.��
l4)��B?�l�܃�.��e��_c��CX����0��Ķ�P��1>*5_�$���H�LM6[}�����=m������\��
��E��nx�,��"�3L�)�P~&tj�ӨU��Se;U��wj�$ۯ	����.j2 �E���T��cOU����z���(X����L��
����-��p�ňN`����"�y�xW�kY"_l}����<����~kS��*;$�|���[Ѩ��"5�W�3���ț��X[V�l��f�d��E�=����#��x�Z┮��$2Kj�� ���aF��Ы-��%Rtjιq���^�D�G�X�X6�[�H����T�=sO�._r��M�h�����}T{�S�B�2�Td)�j�u�t��e���Ws,|�ݚ����D����i|jg������Z��%�-�0ܽ�4��qɑ�'��*l��Ofj��#��^+���p�'�n.`������"��]gC'[��PHvp U�A�"9�N�c�T<!�ܐ` ��rM1��-�e�=�p@��@g�ore#���+<==�f��*^��c3�}�1��g$��|<�Y�����[Ġ��d��hq�u��3EP}����Or
���$ׁ,���c~�Neg}�6�c�%���ON�2�m(%�~��` ^뒓%t����C>i���U9���|�(�_$S��.h�ZǑ�;�t�C{�t��/C�YQ��F��=eP��j�,9�H�Ӟ��_�$bS�G ó֨�oD��/�} I2���P�����H���sZ�|���k^��)�g!x���L�p���Ǚ(_ɡ�#�V�h�A��u=���*H+�(��#��4T����Þ F�"�?{��(��ĭQ:m-�c����%_�_Iy�x�_��*��+�ʙTH,���A�3��+j�&m��}��ݦ8$�7�I&�2���T>Ԓ"�a�k�ޜ��y���+eBv�L�V�,����i������ yN�|�<��-�2���P��,�Dֆ{M(��R���"߿c�6k���X��p����"�G�X��7��$Yϳ}�v��z��`���fD������%���0E8K��|���?O�Y�d('4X~:^�pA�7%G��H�#}7=_�_R�C�&�a�8Z�C@�ÿ���v$T�NnǷP��K¢�>C{��)��P�����E ���Ca,<c�N���^Q��1�H��<�`��Y�����h5��a�\�t��M�#�i1�H$[�Y�mP��"�N؂->�#��аa<;��-��3�6�#!�n`�8Kn��a]T\+YPv���?k,{ƴ�Ss�K�Ψz�O{�2N�z�w�[�XgrqU��gA|O�,��L��2���ln;)�4�$J��ŕ�����)~n�wPc���,$����'�5�c$n��65*�*S��0;NG�$�E�n�	|�aj�6�i���
)J�_\+�Z[�7����5D��[]�N��oa��Z�Tv5����M���0��LcߩT6���m�ГW�~(���ʄ=��i����܍���C4AT*�]tq&�f@�x�����\\������d<G?����A�t��]͌æ<�5Q.bf��M�;�X�|��+��8@���&�R�������-����`���	�!6�!�7�X����N�+L�.Ӻ�Gw�,�C��Iw�g�P+�?���Fa{�C|R8���[���ǜ3�U@t}��/��puƮ��L��X#���6�}:C�`s����e�v�	h�J��3�5Ѧ��Ʈ�+ns�c�a�H+�s�[Ћ�Ô��!=.���A5�:(���P`�n��2E?'�ϼ���UФ=Q��ht��?I���E5C~��Ś�k��;|(NT�qI�5L�;À6&J�����tL�y1`�X����s��E��Wz&���Q��%�δ ��C�}����7|��0S�݌�ñsq��z�]b�W�U3�b���-���ʷE����3�GKb@{�vq����!�������S�A�T��>�4m�vۧ�.�YZn)cK�?�:�w�ݡ
�����m�K�k�����.���XzJ�S|C����'��8�*i�0Ŗg|�&c�=iڈ����
��->����|�A����4��*|#�B������#�u9�D�.����F3el�1O���o7���S|v��TYy�#�(���*���ݪ��u�Y��W.R4������%j����;7?�%6��l8����I:�A����C�����+���2�������@��*�5yk�}�`��)����+� �*�D[t�M	Ќ"��ݣ*�(���n���x����8�A�?��N�_�?o>�Ǣ@��®��`g;��X��q#�lOt_���뀨�<�8��ú�ݓ���o��$ᨄ��_׿z� (����x\���K���n�Pij��}�dF�@�R�iO��}z�0��A�r� m��0�E2_�
�M��Z�e��#���9%B>W��Sกuv�����r�e��
n�_�����`4�e���Y�,�Y��Z�@�� �dK��I�n�v�/4��m|YG�����P��XPx��5|�����$��DL�zQ`H��������,�n
͉y@�VT�1�T�3�]��62:�/��p��Į�5{Gu�b]Ay�}��Y�ы��?$ ��M���>���E ��"�®��8r��u��ʣV���Z��`0O� �ܭuV��{M�"m=�+k����v]�Q{�X��+ԯ\�/�h�Ce;���~5C�6��8HOZ���g'���0dEF�0֫=}y��39;j淝��`*0ʡ�����c���2�EŜ���p.�i7����N�Q��!�.Y��>�m�rŽ�Ö�W������-xP6�my�!g0�Bb �ks,u;����7�ؖ҈�� �x���y�b�1�ȝI�JR�� 'm���(Ǜ�x8<9�L,��j6�=%�E��/8��u�"8���N5�ݧ�BO\{DŽVG�q�S��p�x���`���g(�<BoJ]�	� G�K�2_airߓd���(v�|�5��]8�f;oym¨�O�)�B��J�Y'�l�QQ�k�|8z���=V1�q�b ����B��}�9�
�Q*v�$��"���(Q�D�G0��.ȕ��P� �(�"���9؊�~����h���]���e�d`��Y�	��铄ox���0Õ�x�~ @A��Mx�7�x�
�|�d���]5kRtLC0���)�Ĳa��ߝ-��D$�R+J�o��.5ĕ:���\s�_�^���CD6R���B�1ʲ�4��N�}d�{�C)��9�R�����:"�� ���O���<M��a�F�����D���v"��ސ�=��9��ߢ"�M���\˖"�^��湂�d]{f�Q�;m��a�V�$0 G+���:)���<�2T��ND���g�o. ����a:�pV�G�,O!6j/�E��-
��²J,�r����zc���D_5faF��BX��坁JB���}V�Ԍ���>�cЇ2��*�Z˞�^.���)3�`�h/bH�x�J��(R�W@��	���JO/�C���#t��ir]��}�y >eh	�I:�c��J:[��^�#&�����E����s����o���Oa�oZ�����M��8$�ź�yH뿲�
:�)��1��r�ڵ7H�u���:7?�Xk��o��F��]{�ВYNܦќ���K�\4,��?�F���qr�}�e��W��o����O_�����
<%!/0B�.�.V�/!}��L���2Ȃ�I���&���)<��5a��!~��=��|����L'���0���wrV�!*�c�|#�'���% mJ���cc�tG�Iô:��oMb�R�!�d�4U]����#��wa:܋r�tv�v&h������ "i�wf��6�=�pn�M��l�1�@�dA."Ny��8��7VV�9B�
��b��J�}	�z�@ws���¼�ز\+n�2�1.[@i$]C;`FhZ���F��1\��M�(.᱙��>�����s��E:���ŻV���~&�睜2<:�zʁ�����\�����q�{��R�T� �7�wo��D�Z$�i�7��}�f����W[fUSi�w�F�����G?C�:�5W`;o����75��!+U�o<�0G/%e}�+��}�
��h�^�q�K*/��O�ڿ�x�|�?GE�|���r��.�`��t#���^�ת)̔�mh��z`��K�a���{�ӵ�Њ�u��Ͽ=)�.[���>8�'���)]�������·_,"�����{�VFW��̍��