��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���<+�qlb?p�ӟp����K��>�Vc��e�Sd��n�NmnX��J�#��A"�'��`����N�,�_���j44;��z�fTi�Y!���FP��v��G$Z��$���o~�?`O�,4��C�m�^-+��yUG�T��D�g��1�"��:t���*�&qd����$��ܯl�dX&��׎;"�$0{}EN���hgA���6b�(�M�Og��z��wt>�{����M|t��s#��r�-�4E8�:�܏�%���G��A����Ͼ���O��Ss�k��������M� ���=���hfP�`�}��ζö�&�`����Gn��SMF��7���R��Kޫ�e*-n�R�߿9!d��+-�|��1Mς��K��f��Jv��M�\��\��#̞��{Ϯ{{M �{�n+���6p�hn'��f���>���xk3��x��ۦ;�� �G�{�r����9�*�1��%{Р��ܳ��v
��Y�͛�r�(zT��廞�	�1��(�K��1W (Ej��i9�
��]A��������va��j�~Pi�wv��ܠkL�7G������R�K{a9NC�q��x����$�%[��>����[`�i�D��H��q2���r�����tL������e��=�Cͩ7�)i���R�)���� �zq!}C8M�/�Tw�ϟfHj���9�^�(�|C�<D��o�/2��W���L��q�i��@��7��`���AQ[{'f�68}�>\xP�UY��`�a�-���)K,%�r$��bo*���&j��1Ń^)����Z�R��x��u/��r��SV)^8��}�ֽ��x�:�O�J��s{�������4����-Ė���2�V �r��p6Y�ǼH}c�>�z�[,��*�E<Wy3�F�{�6mD*R"��XΙ�3���Kfs:s;�Ѕ�������ӳ'��߳�+�T뇼���GA��=�'Z�m�N�O����(q��}qX��PYDC�F0�i��MΤ�_Xߝ_�j��㩧-�68U�����) �CaD����(���;ˢ�YG�lC�>�М�*��BS^�R��4Z��sȴ���1[�O���i�dn���M��#<�� E�F$�EM�'���!e��s�%�"=$ַ�Q����!Y�I�*bD�a���?�j���W�n+��h �Y��3n/-2jJz�P�ɰ+����H�D��,=���V#-����=qp�
�s<�Z.b�Y'�Y>m���ү�mO������:1���W����������'[g�s�\{*�3_����lvս�q4�?�ᷚ=�|�[�A�]dom8rPm�+8�1��nRn�R���ע(JP��{�C��L�/��>��!��@�jA�к5���[�"�� ���9������؅ʨ�H�*JD����1��f;��P�9.����x�${��dc�آ޲�7zvl_(�rK��'��������FD�V�QY�#�1��i��;;��21��֔��Y&1��-\S��#�/ �.��C�XZ	�9��W;/��j����>&|7�
���nL�n�=��Y�l$T��0N�A%%϶P���ʤ���_Z^��&��U���Q���w���)q3t�:۟k�$@"��{�7"�����u�m�c�ͨ��;�ظ�$L�m�����L�H�r��3�bSR"}��_��Nt�[��g����a�?����߷�W���L<�}�avm��$�>s��6�P��C��I��a)R$Cf3���VL��	�"�3�D��	��/�!��fF#�(�5���^��^�N\fb�(�F!Xb,��;f?[��4-P����
�vU�=���Y���=�ׅ�w6�I������L1949���&2��o,^䍐���!����$C'6'�
�YT�lr�nh}li/�V�#,��n�u|r�[UL��ER8��ćSz	(�խ���#<_E+!X�����	�.�O�6��d��3�3��W�G����nI��C�$z�P:�/�|��vz�X���`s�F�����H`F�bf���\�=�Pڪ��A�^X�rѾD�9�;}xbh>q��F�k���K��{D�X��x�	<���cz��6a���:(Gĳ�Z5�ć�� Y?v&X�M�!9�v�G�����Y_�v̔a;#+��W�%�ڱ�����&�zu+Z-�ib倱�����"���U�
x�y��b��:DA���Ȥ��f"�a��V�My�����S�v���v��%W����)�U=x�(�M�����hQk���%�C`}xiI��#��LЉ��'�!��sE�[L=�c�)�'�'y#t��~x3��[�%~��b.�w9)l����bi&8��z��w7�_QPp	�/�ZƷ@�+���M�ܙ�i鵆E�j����W�<px=��3�!ܧ��lY��Ԣa,Haѽ���uہ����g���>�0� �^{��0:����<l�>\���B����3���|($�Pd��ϻ����i�u��9�I)���~�F�3.8ڛ�[��&�4T�6��0ϓ�p~�f���	I<VN8r��{�/؍&6��TDt�I~�ז�t��B��S�x�]l��9��%,V	yP6��=�9�x4�5^e��:� ���
���2a��7�&S��A� 3�����-�������!�y�����c���N~i��5��E��B���h��b��T�*��N]+�K,�g�ߴ{׻�@y�*0�o!ы/F ���F�R8vƛ�F����i����z���n�\䑈j���U���0�I��dJ&5�8Ƥ2L��F��#��hG����/zǯQ���?�ܥ�BhGD�gwXh�)�c̵�q���4g�cK�U�������\��K�V+� ΰ���'g)��/�L�s��7q��U <np}�9�NB������	9�����C��qL�ᑐ���Q/�'���6������ ��7)�3i��:i�I~8����&�r�/��nǉ���� &q�WU���;�їǚ�o͠�|f���l�l��r���������W+�s�Z�7l�3�g�ݨJ����9�.�W@QS':1�3|�qj�&;�78�/Lat���|��\���%w㣵EK���V�%�8�Z^�����ُi�Ȳ
��><���R.�0 ց���o8j/��ͼ�m��7��a���fa��M �*u���o�}]���� 2�'��9��@�2�������F���#L�Do?f�A$�(���+u�r�����R2���y5Ѧ#@̔�b�S��dg�Qz�]�<�HW�#:ٮ���~�:l@L���!�����}%p�O������ &�3~7�X:̔?��5�H�׸X��*�� ��A���t��C�X�-��?tV��:��٢�P�U0�?:R�R*ZOuf([�_���c�WT����WJY
��j��)'�,�F؟M��V���/T��#�Yf�x�V�b��Ș52�������p�G����,"�b�qY$������ؘ�d�gd�DTϔ�Ҵmʣ��ܲ)RD5� ڟ��'�>�ٺ�m����(��M_���kw���m-����[�Վ�'�`�K�l���]hm\E&a$�.j<�w�@7��eH//��-a�ĳ��ݟ�/Y��GV�)jo�@1��"�mk�~`Z6&T3Ė�Ui@�<5a�~�L���,k<��r����R��6~[;����#"�^8�����8rd7'���H��������ze�V-���\I�q�{b�+�rčM+��F�t�~h�L)9VO�@���������j���W��0�	Bұ.dG���uC��c�[�(�S)G6�n����	��&湒z��U�i�d�������P*��K����Jϙ�nrV��j�q9
^��PQ���:�*�'�n�5�P��%�r:��Ʋ�UM��W{qڂ	ioHb=r��~=3�{��j�@��E�������r��l�A��.Z��Pȃ���������!&F��INq�.r�u��+[ŭ���X�Dz�!���
��$� ��"�#[��.➄���4~��&g5FJ~Z~u������Goh2�P�Qb�ܾ����8'�b%����HA
sz������"�jl��:@��ⰻ��^C@��G C�<��Tȯ�x���ħ�m��nH����dJ�m����y�z�a�˛pl�A����V_��= ����t5 ԙ�5�Z8��RѾ�4 �D���*�C�5#/�nP�2����	Ot��)����p& &@�C�3�F+z��%��Q*���*�׎��_����. ���#{8��;j�NY�?v���;u���;N;�Nc���~��;!|!?nm��b�v=��Xoh�7E�GSF�/~D/
���q�u��'0<HQ��쩖��1c��t�3;�"�~�U�3�u����<��$ɓ𤏣����K���
���� �J:��2����J�R�L{���Ĕ3�E1H��(=i������L&�ѬV�k�ҖE��O^��ȕBx�eSb��wx��x��A��
6P�΋��Ձ�G�.po�U#�I��rm��z��f�}�vo�ߤ
_E���8�����'�qЃC`�6�~�k�=T/��:.`]�N���� �z@�і��>߾��f�@�81#/���l��n���!S��O��mX�Xς�<��F%�zۖ��H�x6tOP��PJfم$I�~}��������H�<o�zW�������L�_K�X��U�b�0$��"�G��s�u�#�&7ǣbiyͅy���(?������s�<,l-EyV��/�����*��H��Q��Y��)���3I�<�Y��Z ���w��;1H��W�6���D�,C[¢�k�L:!L��?��g���T����}j]fO}Ku�LK
��ΐc��<������(�g�:�誔�*�w|^���\�B����K��
AƑ�Պ��#��3����,�x�M���o��M��g�S��~�Η����ҵ	��VN
�ò4C�R��jR�b�,�s�'�*5*Q�L��)����B]f<rF2��XZ��yD�]��ݓ���?�m�!��2��8�=*�Q�����8}U3�λ�������3L�%�~R�v��ĕsIrJ��Х!yϏ0V2 �a�6N&�{�T]��!c���x)�w��F�5�ɢ{�J�#j|���H0HL��C�blN#}�����HM�W��(����`�o��ج*��V�}e���
���Eg��uD���:�U0	�Wc3��m[�`�L���m�A�KS=}���q!�������H��r�4G%�f-�M��H+]]�?>e횆��	�4�N���Z�ˤʫ5j�5o�#8~.��z�Ԃ>��<�8�?E��$���2X�.E/Z��F$2MO��S��Ո�q�Fԍ@�d3R���"�ӣmD�q�rl7�[�O�8U}`�I��R�Nт�������xOo��k��˖�?�t���U�r��G�ܬ^�T�I��O��'�n��y�)�Lj��=�>n���%��a��0�x��Rê�]D�I���
����k�:�`�i��8��$��`�Hv[���(#�P����UgQ���6������5m!f��,R��:���,���GB��U�ݛq��J�X�m1p���aD[�-ӂW #L`Bk����VU]���y2���ϴT����
��:�Nm�m�)4��!D��e��b
.S�A���H���՟��^���j~��p�@�"!�@T�<�k���L�ihiȯ�]�`�D֦R �cW"�]�����+�.�{�<�B[�`�w�>�H�V��,���4���1�La`J���xs�vVn(ZX �=�v\�4�5�-|צk)��9r���P[<1ӾR�1Ѷ�>���B��B7n�cc���z\����p{�d^�XsܝpV������v>܄Ѳ���L��"�P��<�B�h�Vz�{��mw�Q/���g�{'I�ޚE�ݏ�õܫ~F���I�qq�X^����`N�Z��S`S`�q��1��E2޶,�^-������j�h��&įJ�6;ib���r ��۾>���9O[�Aqe��b�J�v~�A�Vځ�g�bŅ���X��H��8��
�0��-��u»t�(��e�H�_0���`M܂�ߙ��_��c[ %ά��&��%2'�譞)���Gה�;�{xEs�z�P
xn9�rp'%�}� ��x*4��O��7�\���D��=�D8���NWL�G2'����	Ӓ��MW?�%�a�����L���%����6�׉�y��aOx�U����5�_]~�{]��tp�����r�Qf���|����)�n�+��0	 ����˶߰����&r�>���t6�(�^��}����)���$A���sZd;�.8��h���Tc�m%����4Rdu������=�D���>sd�)�P�oץd�i��ޣo��WJEY�b֐¾1������1.�n���܁Ћ��㞱d��5k��t�=[��
W�=sg�^S�`ét�  �oU��1̈́'���}�ۍ�`?τ	C��1ts�!��M�hZ:�'s/A���WϣÚf���׭-�(��+�h��[���V��6�O�~8$��{g�2��'�|�ޞ�RSŧ���3�37]�4�|����#���l�����pVwhMB��iZ�k��ΓE:h�p�?�[WW:��O�:u���C�G��2�EJa=b�D�h?���1�����ʹD�ּ�l����hG��k}����������4m����O{��i1SNj�{�*CNK�_�Q�G��,O$3�eM�=�h�,� k����=�����Əa�un��V��m<4�(�'��x}�;ʻb�uj��4�(%�QE+�{+�����df�)�Fo�d^�x�Bh�x��	xH��&������M !Ks	��r�&1�W^�_>XS�N����sQ�{�!�~���쑜�U]��ڊ8<J���(԰��;�a�Nk�u_��$��]4�$�š�F������ò��Ii ݠ���O}_�����R�*�^p2��Ճ<*2��+X5�K�F!��|l�;��>���zg@���ȉq5 �.��w���n��|u�_uҷ~|ǹ�>g�8��~���Z�?R�����D=`�b%3�<3Pf����*�������bnyt��`B��4�-��N����(�w�Eq]e��Cq���ew�!@���{�X>�s�R-(�<�WQ�/&K�0��[���33`o�� ���p&V��o+Ю:%�;-��2݋�0>�ͦ����	����?��~g��5�yK��|�i�3A)�y)s�N�l�ޏ"$�xWM}-�"�[���K�)�[Aͫ�DGV?����"d�r�m��ˋ���,L8.�ݿ*M'��)�ӡKc�f�Gl���c�KO���`�&��I��o��ǅ�8l_I(]��b[LF
�
���v���"͢��������}��➹h<t�ll��d\���Z �}�Y#�9Bp��.1�c~�3ݶ���������C��������D��	J�?�|�7Wx��������3&��q���� ��`��&�8���m��}��6I%�c����X��5`u�%[�<~2Z<|}�q� ~�X۪���)R��ؕO���k�gu�4YT��u\Sd�
�l��VIO�e�����`���9ӤU��(�b%�)��a)��dE�;���2�\�S"��T�0��7����V5qb��x$��5:��d������w4���q/B�������ye�|�1|:s2m�`���.ב����;�ʥ�L���62���j�w��,����]-����}A��Dt���H1���ث����3�5�a�4!�����祭x���� ��T�yLs̯���DH�h���Nn��W��)Ѷ3�K8-i4�im*�o�72��L�"ݦU����W�ɢ4!?7U�ox��� 0zq��G.��/�GC�8SQ�W�3u�PX��^��/u�J���e��I��P�w�;Z~����D� �/���`)S�����X����S����7dw�n�0��u� ���c\�ZT9�f3<5�O��͢�Ί`���\ �]N�4���������bZQ.j��!�[#V�,�`�M^Q�N9��#����?��FO���T�p�6D=6�m[N�c�Č47:��z4�{���������j�Nh�%V(�v���T�[�n�V)����Ǿ��!����ǆ��T��؊nI�Vc:�	��
�7�'X4hؠ�bx��zՅ0	/����<+���s���_H�k�gf��+�F �o^�0���y��
]_}f�yǙJ2�_]@�|�@��B���T�tN�����NQ �=�`t.S����{���գҸءquZ|/�'��1}��~2�g��QM������PRzuSb�����Q�7�8�ߤoi	{��Ey��;�s�~7��Xk�@�ƈ����c��lٿ:ȥtMX�>ًo��	v莶)��� }��:VK��b�M2v��^¼k�p��E�H��Nt�#�S��eNpj����c�A�$���]�ջ4���
���*�r�N�k�K��Jt�.�h��i��?(�K(�J'!�1䁑���������0�Sv*��^�����?�~v�?���u��Q�M&	e�g�L�'fb�"y��.gDk�l��l#{������}�0���рj�g�lJ-v�(��˅�oy.HsX���{��/��cj���(�g}����M�����.�%e!Ä���\�2,�<o�g6�H�d1�����k���(Y�t�u������c�)'�M	�շz�����ˢ� )��B��8��k�	S������z��$�Fx
��I�glm<N>��{��g�gt���J�C�j-̶��v�m��vp+l�����K͎:4qz�"q��*�W�f�	#�i(�*�TB4�z����v�����ezlR�+$�x����#vw�Af3�a�ՠZ���V�1m��l=PfY��0�p���V����f!�Xs+���XdD�� ݗ* �'
ﴄ��6o�t��(�P&}�{��k��=��Z����ЖR�N�����13bt��'��)��_����+��C�n�Î{�寓׫����՜�v�4?u#��VI4$��%���w�#H�b�t1�Fk� c�g��gm�z�	k"�z��-�d�<�d���mf)Vף�E*��k�V������?�E8^R�˩v�����l�T	�PRT���zՌb-�Bi�A���:Ӷ�����#�4�ؾ�38x��!���aq�����r#)�K�:���6�2�8gq r}�x+����D���56�Q!Y{��׊r	ҏ�g�>c{�X�B��ܙ8	���s�*N�c!��j')���U0�1���Zi�B���'QW�%ȑιi3�,4JB�_~�o��m��f1^cG�Rt�5�iv�s��hBdcO�����'s��Dw��4ƐsϪ��Ќ�����%KA���C��%x�&/-�L( j@ܽU�L�z�b�
�
p=�}}��J�7�a�If*�O�19����[�4Q��/��l�v%i�p�kV^pƊ�bS���1�s���2�vsΕ�VT�5�9�5�V�#t��ߖo䕻 z��{��p�R�_[�S����2a݆m����3;$�66�F�K��Kg\6@���ڮxi�4��q|W���P�"]n����>#Ճ �r��ktϙC�>���m����7��h������?���?7�'���Vp>YPi;����U�A�+��fb�ܮԆ�ە���1�4A��q{H����.�G��$�l>Zo�Kމ�i�|�a��>�%�BS+���H�Gk�uQ��ܵ4���ņ���{���w�����j"��[5;$����.��U�:q��;�]���vyt^�1�f����XٙF�|	� P�Jm��BRBz��ր���ݽ�/���Woo������N�j;a�	c��{l�gZ�$��C���VdY�����\���z,a�*�k�m�ӧ4�T�d[�CJ9��C����9�Z���8���$>_�`�<9��E�!ȳK)�]t�����H�=m�� �2:�����[@�uJN�>kZ�Ī�<y�{��Y�
��W#�4u�RWB���)YdvHAv@�Il��,��/�#D\p�D�is��E��f�D��I�}��"���8�nd�b	^I<��[�rQ�%<9��O4����W2�K�������a�t���Q�Q�)iVN	�f���J}�A[����\�(�n
��r��v���tT�/�JG�����ӌc�)��h<�7Z�4UoM?��po��\��/���6����f�?V�=������_��L��>a�5�j�k�h�>K�+��<}�|y�5�Jvo�7SO��i��
v��k��D��vP4��Go�@����[n�f�c��]�b8�Q��/�wc�����6P����pdǛBu��.'yR��2�f�)i�]����Jwh�cE��
z�2K�rJ®�U���_�.�㢅�f'��*��p ���O�hȶN�Y�h����jY	�|"������=�ۤ=�>n0����i�C��I���-k�}`��Y
.d�5�֮o�v��.9]�)G�	���o᪲Ac��znk�g[�ґ��@�h�J���[s�i�W2�����y���y뻕@׮T�5Ԋ���-Br��(�v��UY�68��EhUr�-X�c�o�	D�!FK�XH;�A���\C[�0��&3�[�!{K�\OOUW-�k��Lj�� T�N��c􎁝���G"6��t�f. z�W>����<J�/��˛R^�+`�z{|�˿�A~��qk�\������6{�����\!�,�gIR��"�?�x�ڱ�썔���6S$�ITV��7�RR�xePb��4�&�'�����+#E�y-�$��(�6%F��а�?��D���^���@j�t�������ט��������YՁ����3��d�'���t�� �>����T߬�0��W�(T &٤M�\�:yj���20�d.��r�l��hO���XZv�h�1-kpb<�Z,0�z�9C��f��Mw2tU�+ZY��7���r6j 9c�5>-H��lM�uͫ�Tfq�1�� Sz�U�@����0�~M�R�� �;��^�t���^K�����g�h��CڢV��-5���c�3���Q�]�؎��n�_���z���{ߘ%�����O���T�rZ�N�{��C�̷p�-��j���Y�����:�d�6B���b>��f�Q3�CwO��\?���6��:�z�%E����