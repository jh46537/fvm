��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^�.GJ��-��?f�b��(��ҥ��Y�����!���نϊp��=׈�kS(�?D� Y�S���#��f�����V8?�_���Mg�\��gѵ����s=�B_M�E�B%z1�����U����\�����ZI^C'���d�_ ��-[b�DU�Vյ��*�0��/�^�]ݚ�Z���r �Ї-�l�h� n��ࣁLR�5���e��G\"�JZ�z�!���0�.f ^w ϴ� I�L�J�ȷP>���ө�,5�%%�bK���>�͇_|'xƈ�&8�.�7�ԯ[����!�X��fŷsIE�~O�l�d�O!*�W,��H�����;}"���9��k�CD`Y���r|��# 媑6�x��31�_y����ъMd����<y �߱o��)a˘Q7���{;L��:�:�6�w�K<�&W�u��wK�M���b�[���h��������HC�δ�;ի'�(�����Ӥ�@��$ �V]z	u���#���ځ��2G�#�B	�}x��G��߳~��Yi�y+�����(r��ꕛߥOy?���B���W�uuB�d@�Z�ܩv��x= �ap��X��(O�vNleJӣZy�D�o��/�?t ��0��犢�?�T�*0��Z��}N�YE�1`>�	r�D*�>���NqxVJd� S�3459��]n��H�Dﻅ"��7w�a�t^|�p�v�5U->���^� �}�c��@T2��)6V豓�"S����Uf9�g�$j��j����{?��S�X_�H�_\��ݞ�D��.V�H��BF©�;)B�6ƨ��J?����(��-���4V@/!V�c��\���>]Vm��#R3Y�;
#��h'
){����Wc�U��B�"�	qB���L!�v����܈u�hh�l���-eQ����IP�����^�O2yؓ�Gz��H�A��~U�g�T�
ΰ��g`�J�'�dd�	���(�����w�� ��/yk=*[׳��n������%{��@v����-�?ţ�n���M�I�X��	Nf�d��T}n�Ph�Lh��{���?KUiuf��i���nq�`���F�d��2b|���M,<�R,aIx+���74���Ԭ,������J�Nn��Jѯ���3 *�Y���VjJwz�O�=�C���M܈o.�����k���T��r*<�c��p1i&�~M�3�a<v#�?_��)�ܻ���Y̺�eU�&�r�]$�^��oYxό��R(Z���Ų��<Zʛ �E�TY�.�� p�A���vhD=jɻN�pW-ꔞ�^�G�b|b=��<L��7�[Ф|��%l��+�_�~��M��I�%%���xk�T�:)L>�,o$��_Р�� �4>*��#�mY�{�R۴�F�I̸�F�]�=�E%�\�馔�ɾF�*=�T(6H8�50(u��=tC����M<����щ�`����K1%ر�҉'{��(��b>��^Dؑqzo��z�����K~��q�ы������'S�gzi~�u	 ���ox�\e|K�)l�F�rg�^5��rf@$�;p1�(b0�ƌ�+V��_�z<����*������

X�?t�o9�����a&3�z:�E��(4�꛻J����m��c�2ێ�=�Ĥ��]���l���b����x !A��~������q�4f��r��3���=Jc*G����g^��7��r���6�M ^�b"���WeV�	��/�����iq7��E^����B�ڤ"]dh�[Ң�s�3!�=G85i�{�*w�|Ń��?�G�B#���!p��r��E�Z6!ȭ^�r�wKE��c��SC$v��tb�7�������0H�u�zC@�z^��o��T��� \����S{�%UM��v��wM����9
䇙�}���h����-�R�����1�o0/�o���H�(un=�ſ��A�R��HW�/d8�%�>e_��וcx �"K��*��ت��	-*��M�K;�ח��C[B�|G��4�b��>V87�f{��?��f_�g<���,�H�����pd��8�����_j�Y�<w!&�AjOtkR�ue���:w8w�X�i�{�����X�N��c�C"��.�5un ~�d���rۄ��*�3�\?��?�8���U���B��m�-D�2 ��ς�sC��Ơ���#���������J��;��t�X�L�Ϧ&D���rq)"J�0ܸ�h�ZR0�+@�˛h�e�p�sq�����ȋ*��"��~��G�_��j�0T�_�{W<7���6oϘ�}��S��`�`d�TW2�^rq,A�&����/�����?�����9���|�k��2�����M�F��o�#�b~�Q3�b�4����'�e<:\����b(�5G��f���A�w�*t{�R9��xV�H�'�Z��0/}��a㎔,0��i�g�I�d|<��w��sd^��mt���c�dKAJ��4� ;'�I���VT:,GE����7��D	�Wo|�^�H�Ka�^�vk��m�#-zʷ����j���C��GA$W�X�R�䵦ǔ;��6�]�^���:��z	�仐�GO��{�n7y�=��r'�*��m
������Xb]V��>wд�rD�\ՅR��*��~q���g(����^F3�,v��;�m��ᣊM�I;P l�C�.>˧���T�DQ��<%J�OS/��at�ߝ�Z&�-���&�fM��7ci��T����?�/zs�oKoc��%*�<ĵʌ�f��_����*v�(��s��
͋Q?��[{�Z��[ߌ8�)P��2�e��u7�[��h�%�h�f�\c�&��Sw�Uٰ1K����ɻxv��W�����N�6�G��#����dF���Y��r)ٱ�C�)K��m͛u+.�����og��:�˚�=�X�u��b[a돃��0��cֻAx�o/��b�/������N�?Ï����\��.A7c5�џ���~�m0�&�H�,4i<OopE�iм�Uv�zT�$�6�Pr|���b�1���2q�EyW^J��l�ķtE�mo���U�([VQ���`�`�%d+L�:	�cR7@O̯��EFfrw�MHG��3'L��Ϯ��2¥�xM�[�J/�ێ��E�����=֍��ǯ��ة�n%]��!XH�����+و9�?ǀCJ�	?��Ʉ1��<J������9h�ھ_�a֧&qA_ٙ���z�6����/���ID�O:;��p�ל˶�xٳu�H A�^�˒��Ό�.߅yY�,v3��m�f`��9�s��"��0>��љ�41��0VD�Y�IE��1��	��%v�i��Kٝÿ�8��iċ@�Є�㈌gS��0��@f�6��,��'Rv5$H�UP�p��8�ե�j��(�w����v���"���Dƿ�rW��s���]7x�"S]��p���i��Xq(��.,��a��k!P��dm���u��k��y��n2��e�=�2�Y�9�^���n�ſ���y�⏸�&�T3���j<�;'	�K�'�Q[0(����J������\��э���l�>�_��i�<��%�.�|Z��-��[	6�~��<O���4�E�_ Q��Y�b�t8�0�a�"L~�����`N�-5Ȗۻ�!(���\,���	��1v���4�;��������QuWem�w`@x]�&�ٻ� KcS���?o"�8>��L7<>��~�Qߢ?m��\�'��w�@b2p)	.TF�+̱{f��!�`£��u�G���*�{Y섳W"��	�T>�&Y�AP/.(۵����\3�0"�փ����vj??iy�ɸp�^�=h�!U�j71��oW��>�MFԚd2r6!DhfR��T9<]��:*�S, E���cĂ��b�����i�%�
$+�}� �aH����ɶ��[��y�PG=������>G=4�N7\��Su��:�r!�hH��볆Ie���H�wlJM��.
�NNL�S�i˞Q!F��Z@���N�
C<�hZ?��Y����H�B���~B[d��A�qй�FPr��[�Ѯ%��|�X$�����(��7q��I5�߃9�5N��	h?O�����U�|��Ҡ�R��D�!e�~�>G���n9���N7a�}ZY9��
h����1��]��P��ݟc��`�>� �X����[H�3ա6�E9� r���J���V����.��N�'A�b��$@�s'�
d��=�S���\#���~v�h�[�㗩���f�'���S]v����W����Sȓ�Y|gg�3-�Q"�>6�����2���?�O�F�E���h���%-G0C�̥`�N�􊞙`�$"L�P���U�6����TH�<`�l�!&�@�	�V�M���l)�"����h �8sM� }q�C@���)ԁˊ;Q�jṇ���w�r~!`[F��A�
�k�ض��|�8�^�6 �aws<���؋�ʫ�5���҅�N��>�g<٩�|���cklO��^8�Tw+2i�t� ���I+��Q�x�ܥ-�qk.�I��\}%�M�Gŀb���
��u�sbp���kA�b������q�9�@�?P"���^�LT°��eP��������`Dg�[������d�v�Hj68�k	���;^nL���|��p�׀���Z;m�k�Èx��]0waP��^�h����R�`����`>��v)����r�b2,��0U�2�H��W�W��S��_������uu`$���G���2����@{J$����~�gd��V�V[3k��q�{Wt���O4�,�s���8Z�o�=}��֗��߶eי�e�(/� 0]�-�B����bh�Q$K|� խ�X�����H:�Kߟ��<�w=m��#xɾ��_b,�]�/�,�5ד�H2;D�T���1�F[�a���ℨ���̗Hmkq��Yj͙�NG��	��J�9�TJ��h���V��I3���B�u��[��+��k���]�#�� C��x�`&C�9�}��mQ���78�H`�d;� �/�{݈����+�G�]�G�s��)������s��!<I�����������	�
n�h
����k(Ѹ�{�S��q��Uļ��Z��o�+
mSP�������#���A�f�� ���B���F��F�-�n��%*�P����lY�۾��gU�q_�l��]f	�ӏ�Z��v�>E�f�yh��f�v��N�r_[֔G�w#�ʼ�vQ��C_�E#M�3	�k�
$ L��o�\5�� ����-���}�y�[4A1��+P�Njhr5�˲!�E�b!+jk�{B4�k!^
��m0�$�ź�?T~cew��NFw�f�Q;?
4��	S��HS4m�ت�'Un �C6�R/�ý���Z�]�&s�s�?T�!Ss�LU�j��G}Z%zjНl}�F���Cc+:�LV�u�m{#[�`?�:�'�w�]��EyY���)R"��� ����QҴL1�O�_���L�Um-�L��"_�Y��f�,��n�����޺�ʭ����.;�����G������Ԅ��^8�M����(��f�8�s��1��H��I�糛���Ǻ'4�*�7��k~���=| ���Nm�r�e�=��eu�"{�i��A��U�=M���v�\��$�U�H����ǒR�"Y�l�S����˝�g%�;��������lSҪ����Z�z�ń�Ԝ��
���1(�h	l����m��-{<�}QN� G��u7���8C�Ɨ��kC�� n����|l�F�1Xr�-A[a�n[HA�apk`瓼l]�IO�W2�86� ��6�;�� 9l�Ǫ���*��w&��0���]��9� �ޜ���&��px<[N�L>"�s4�������O���L�9eZ�e�����
��1�'���#7�&�5����Y Vɚ��}o/�/�^4�]3��U:��V�� �-y@��Y�G�R�k+:�lڠk��e�c���U�6��Mn/�ԕ))Ư�����������HqQZҎmt���jO=�T�9�ѫ�� ~]v��P@U��p���;�=�:+p���{��� ��-]Z��Jz����a8u��D�7�AjN��	�)IAbdf7}��O�F�����D�L.� X� �ŕ�Ǟʪ�o>��.��z[v�u�$��e_��FP1$�4Ȕv]��%4Ѱ�U:+�T3W�Ǭe(D�9mBt����	�\�߶��BJj�
9#�ߒ�#D���(���{��R`�Q��ް� �۪%hB5�JB_�V�`��=`\q%D5�,;�B>I�4b�P��>Ύ����0Q�f����mc��g]��\��>�g��#�Ae�->���0PnY,˝�E:���q� �]���9}�6I�%��:�U��j�~*5�j��3̯���ȏ!9i����/@mælw4|@��vV�+��ں��-��s��΃��^?x����b���\:��B�Q�]����7�ɰ�͝��/�^^�Vf�EL����{�yd��}�)�)9�k��W���t,�4���-���w����]$�n8O#��FO�n}�u�/S_��[~H��=��B�C�/�䣑���h��6_o�٪@"�[����&�T;Y-Be�!�Ч���\dw�d��{��En"�JJ�b�Fc��8-��K���:�����拂,�y#L�\a�2M鶣�Q�?  �V��
��яWL�d�'(s}�g�U۶l�eaS��Hq�#e�������?��y�����؝]�������D�d۞��L��c.��^��.�<�n�*��ّ�Bah��'�¾��jǿ�Ӓၼ��+7��U�"�e��R���N^4��s����Dz��9��6XU� ��lTZ4�!2֝@�T�4�N��U���� -Z�K�Fj�ih��0�6� ��o)��o*�#��>�w�O��?Cv�ڟB��?J�)�C	�`)ɷuKVr^HO����p�`?CF��F�RO�&�Ϡ3Ήf�TE`�{e���E�et �$�c��E:�p�;߲@8�ŹO���>V��	/an�PxB��
ȝ��L��)�~i`�Z�@v��Tw�$�pC�{!eG�s;館of�GG�����Z[���&݃ig�~e�2� +��J�"�k�\g�]�A� s8��n�YYD;�[�I���}1�Y�f6w��~�3�9���ؗzE�(w���ͅۉ��M����,���[ъ�
-rUPG���wJ(į�E#�]��M	�L��5q&l�
ū{�P�B���a�XS4|.�F����K�L�Q���xWuo��ء�'���(\�R�X�8�ZǍ�f�[�2�w�S��h�����䣋x�a���ɪ��^��PY�S��T_�'���J�O �u����;�
��;�`4�B}5L&�w�Im�H�������EBRe4���2Ԃ����.��~O�Qo蝀6����P�^�1{v~�sz[���sY�D^�P�Z��"��F<ѿ#8ME�G��7oN:�����f��9�:zŏ�<vp��$0��1�nY�o��1�Z�Q��D��t�ı�L3���\$M�M����ɛ#��Y��^>�
��ָ3���L]iUԅ�$��Ƭ�Q��$Q���A��g���N|s�o�\�!#��M�t���̫�kc���:*��1�%6�a�7�2,\1�����S_J�����s��B�8�m�WhM�d�!�Af��E��R%|�czJ� 1�f�_����Fg��*�Q��7I:1� 75(��z�J��v�����L:ߧ��,q�+v'ٞ8��*�-��f��!�d/eFЙQ��_�;ѫL���Ȍ8���:fj���L�����z�p����iuU�@���m����́tW���T�5����H�ǽ��'���m��3L�*_#ˢW~��Y�=��L�#Xa��J/2\��6(��0��w0�x�ksd���߿�~�!�OU ��W���%邤_ٞW�{��#�Cv}}��D�"DA{�".L������Z���-���(>����}��^@�BN�N���N�[ �2.�N�)S�p�I��οö_ǂI���E^Ӭ�'�Q��^JR
9���������FZ��q��00���u��b��
/���~��]�R���PT*�r�g����ք�8��%���R!��?̵����x�����9���zQ���E�
��]o#hA.;��i�򿒄��Y�]�DE[��8WG�z*�ؙG�u��8��{�pRE���W~���u7��KJk�����N.� �x��d�H!F��FN_`����W,���R_�~�2q"�ih��ÙO`�^�0
zB�{�("yJ��xK�Ao����t
ڨ�b#���� mE�)��[e\����Q�}
����gN#w� �<�H�ILQ��������J�4��%X\�������'(���N �����rBu1el/2��xU�A>�6�V�����<8������@TOxr�|Ѝ���ړ�:�/R� N+��+N�W�$�G�2՟�HTC��P�������K�K5�_�x�ʠ;� EIF�n��~ۢ\ā�����\��/Z�+�D� �-)��=��"��S�y��\���G�=�R|���������(s���p�}C�1ϣ5��g9�bB��%�+|���#yFY���,�#*q�|w�:���j����z��`�]�Ӆ�z�qݛ��s��&�O)�TQjT�=��jT�0�*�[�
j}})E��xd�Z�,�&'���3�9=��-O��x����M�ژ�%>v���%v���_�V�a��{�Z^�F�[o�_�^��h�"�s���@'*���@�� N�揜53�Y��<�my�Zh�84Y�D6UC�Yd��Lq�;*H����<��,���������"-o|r��)͵3�1~�7�p�5���*�z�L�O0�CQF+u͙�C+]��*����}��wD�|r�
��x�v���m�Cے'Mtt𬥵Y�-N{�æ��d/����x���èà�(�O0�\��[�q���0����<��V�:�YICFzz.��g�h|��+�Ҫ�g�n-[Hj�I¯�1_�c��<���EW�r���4N���Dkn�g���&��6���At�ځ���}�6d��z��j� ���Z˿�5����i|�}��I��o���G�F<�w}R*�HEM����Nh�jj'B���F�5�9�Y��iNv�j�1���x�*�F8�0A�e-V�~u��"J>c�4re�P���*�� Y���^��"����&dv#o������j������6~�	��@�D�úg�t���ÿ��$��}B����O�f�a!?,u;C��A�����-;vw��||�)�,�O
\����ʇ�
u� z\t��Ia���u7���cKY1�Ņ�rN��3Z���\7����-��N.�Vi�斣�=4��V �Br�	�]��m!\���_�^l_'��~�7\:l�0�Zv��fBQ�q�n%�C�T�	�J��?���]x���~&�n�����3�x�EY�C��)���LoEQ	�u��H_H�x��qy@�]��$��ph��[E������T>�h�iǤ��<ҡB�i��1q]��r�һ�F螤4!�]��ѕ�A���/��2;v�P�)k3�`Ą�)���Eֆ(ww�&VtJ��g�#&����̂��-�H����z!L<���u�����A
�g��QJ:���P�ׁt��̎���'�wI��or>�G!��U�9�֕@��&�ϋ�yYV�j|R_y'�9>4Mev��ӗZˑ��r��6�m_�昰�pv���� Ë,��P�65t�[Ǻ{w���p��v�5V�s(��쇅��@�o� ��c=���Z{LfʚCpL��)��..�͛��3uE���%�T�t�;p����E=���3�P�<�砵,/F=���z5j�h�����m�J)�+ً����@����E����R2�j+}�!���,AP�&L��[�(�8ai�P��g>����O.����^gRM�=۬��*� �x��ctZ�d����9=��-��,�Ϝ/�1-�^��8H�����L�h�P�א�-'>�b�b[]�w٫2��tOu�ő7e{3��!�Y���-FL�t�H�Б��!�˟������D$:Jt��f@��@����<��!^D�M
2�&�m8��@�[!�N��8�M`�R�	��F���f�3�ǽ��ҭ@��G
a,@���D�[f�}eLO;{����~tg;��|/0廚�ͯ���#���ã�@l�Lt׌'Mط(o4!���QLI�4�ab��7rWۛ���`N����O���m:��>�%l�q��!�[+���;m#]�g���9HfҞ�fܣ��Q�z�}�+!�W����)��gQ�Z�����WN�B~Ih��>�[Ͳ�.=�͈�,�Ց�v�Z��m22��vU��rRƴ΄њ�;�b���I�i�����j*����[�U��s�Ȣ�N7Ғ�OJ!y�G���Tw���p.q�2�RKZ(J;�m��sxDB���>X�gei�u�!1�S��i-�e��PH��Hl���)�[��E�o�2m����6�%�xc=��P
��M�k���l؂�n,�@;\~��c/��pR4��Ҏ�.Mu��*s���I� ���Q�H�R�\���?(֭��Q���^�0ޱ�G�����
	���;� -O3K�[�|i啀	5@Wdj�my,p�h�R��\��~	� �4_4��&�)�(eA���[�1�-���B��IS��6���J�#�W�?��߲f6�����	dn��T ,<=�= (�����T+;���m�(<���k���aZ�.��m�%:��K#�������nu�K �Xz�L�R�:ܭ�&�4]5B��z9�Qi@����~���ҝ\��w}���$p9���%PUD�= {��̰�1S��r(�)Y�x�.9O�<�ȟcTh��=�Ɓ�.�N�y�ə\��R��t������LŒ��>��eߕ����<n�5_2�]t��O0�H4�Y%}6��y��5{jX$q��>�y�[��[�mM�G~}���ld��r9k$�J�N�o�oN�w����u��k�]�^(_����X����DS��e����f�˝pd_�n��=���v�ڑQ�l0��9����,_��9�q�������\#r���%ħ�I�E����5��h	aԫh�����y��a`�c"�J�x����Xj�`�C�8�����T��U��Z��3{W��*qSB��[_n��4� M�t�?��1� �S�+�\Mz3@��x���\7����Jb}W�TƦe���bzA�t@�$�����7���/��h���!��0qE0_]�w��>�'�{{O��E'����z ,-՘z�o������)��n������cULXX�:	ޔ��ܬ�z�ۅvиB�B�3)�l�B� �2X А�G�p��q�]���Ch����(��s��ژ����s_�S����Z��c��^�J��q5�̻mr���p�z�L��a�Qf�ze��3����g��o�V�	�R�ȴ�� ��9�nY�t�Hīy���[��ԇ���X�����/d_�WPx��ٯ�ht�`�"Q���,�(=_��P��~�O�0�3�4�bq��x�aT7Ë���:i;H��� 鳋���ن�|6[QPW5�v
�TX'9[��̗�W��*�7�w�#�~#{�k�ۓ���1-�K��&��~p.]	��3*����Iga_h������~L$��Yq��mD��υ�﬎ڳ�ZB.'��rJ�PU1��`��R�vc�w�Y[tfV�䯬�)�m�+6�b���6�7���$AHQ�@ڞ��u�^�D���ɖ�p��d&�C��,%�V�:	։l$�D	�M8T����䒊����to&{��C<2@W��X}��q�
^��n�f�ԙ}������Ê
D˹��w��e���o�*�kǀ嘩�%�K�T,_4���!�����pd��H�@�>��{�@��L�%�$Dg�I^��5Pd��'���|:�f���)�igr}m�A}~��=.��������������b��̈́��[�ˮ3��Yk�<B �k� ſ`�vaR�=���O�rC��$?b؃XD�j��o)�ŢI~���>J�e�V�����O0�����C4��X��X(c�-LB�L��[_g�e����W����Gĵ�>	L�3��Ex��nF��>j�W���VH��ȃDs(Y�1c�< z��bk�\�ʥ)&d���OzVb)�ۃ}�ؑ�|١�;��G=�|w.��'�~�\,(l^��qB�_� EJǖ���[�B�ߛ��4�G�xd�
b��\�
�^%��LĄ��w'�%� %������A����zn\�$��AAc������~iVh򿙊�_�O^I@�^FD�.O�U�5�Ee������:�lW��;�С�0.0�o���,^[b�>n'�����|���`R���"�����Z�����R7d��ЕLu���%A?�>�M,f���F�gFrG]��������o@ݾ���ƶWppr6�Y�H+6�\�o�J��ɸ�k��1�M%�2��1�>ܛ��Ԟ��K��b�<:�ģ�Q�9���m�0z!k1�:Ҍ:01-RE%Hx-m�{=�<w/w�sB�r�Nkػ�9��	�r|(��nS���+c)��c�S$P������XF��[`����Uu	[`0@{�t���[��	��X���a�� �����e	��W�tRjz��0���B�P�~�ѕ���/���Qi=z�X�Df��xEr�V ��Oh�h����S��B+(��\8�Х?�9_f��������iIh2�s��q>��Ͻ�A��E�8�dJzF�O`�qW�Sp�uw���5\��]�������;ͧ�*�,[cU���Nr��_��Oq+�!�8�����o�5 U��d�NY5��~��p����?a�r��!Y�4��W:�o�7Hl5��۶�����:�L,D�������\�Y��S5@��2���>RC2���mea0.Wh/~�X��o�>���
���M^��#��j��d�w�G�h�'o~L����Q�b��q�is������� ����~t�}on�� ��O��v!Fh�埿W�^�XA1>&��'�)�f��f�K-=C��,������v�{W'����*��9�z%�Q�Q|��dѣ?�v����.��J�|��<lAK�
����A�l�n"~��(�
�����ގB]ٝ��5�݀pr �2�%�h��i�"Gg��Z(U��{�-������*���煪�V͵JrI|fJ#�q����ď���"�g��Y���J� �N����[t}��G��݀�}�{vx��fG��`΍�3P�
�68č�Mess�W���e���ys��/��`�8G��s֯�?�u�x-z���dD�(.y���GlP�3C��N]�ĥQ������D�2�.���vɯ5�"������"U��c����l��;t�x�/)���0�Ӌjq,�