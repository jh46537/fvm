��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�؆���o��9_��ʵ�Fꙣ>��IG��ɖN"�(Kcf�Gޚ�cm��ո^L�
���H]�FǊ�F��ak-W�e/��fJ�|���ia�o`���:�D-e̫�/4�a�0��v��  �L�ꩉ�h�{ͦ�P�6�9	��9
�]����(�H�����UC���|���c5�#D���D��˭�s��U�w��2��0���s�\]�kV��)�Iz݆�Ґ�����qֶ��%d����-S|����7Ì;2(f8� P��`�l�-i�r���)��m]Ӱ�H�r�mM�z�9t'"J���=��0�Ͷe�W��sh������`J�i�K���Ŋ�Ѡ�O�V++�6R�v����$�W�Y�^���՞j\��>�p#1I��e����D�M&�l���B����� �5��O՚�ڇ�O"�J�Ī��V)����|*��G��;i�g�$�j���W�&��2��Ƌ�'3+d_��Bq4o۾^��o<V M~v���9S����GF�ړx�������6{�E��e�Y#��I��O$��X5�	���ø�||�o��o��j���a`�@��H��P9`%å�/.p�v��K	�S���D��C��g������<n{e %���P�VHc�����pZ�.�������Z��kuN�^p3�J�ٖ �>�[����^�]	J4*\���U����}
�-A����	���:gOR�E%ٷ53��-�4���G�T�|��ޣM�.	Y�Ĭ�5|�����z[�W����l�ݛS���h��s�6�P��T>/p.J[ ��dt��������H��23�J�����>f�i� םֺ;_����|( ��}��q�>4�y������2�&v��c8��1��\��6�m��#�?�߉?�kv���Z����m�0P�6H�}a�訩ڙ���G�*��pO�]·�N��{��5��޽59��Μ59"(�`{�Vˣ��̈3��U���q�c�?������, H�g>�7 �Sd�ǀ��;�䆬�����u*���"��5���>��A�d�h6��c��@K��]��º*�\4��؁eI-[�Z�OF`�bb�1��}��R5+�	�8*"��&�����zr��ys|'Q[ =�z�
�)��e��O�[�������P��=л��8,��i.���s��6rzgc�G%�D�ߘ6>f����`1ĩC��6���PU)���I��XA���E�����g>+]�)@~��O���ѧ"����h�ˉVo#�gR[�xԁ��2��D�z�w�&?x���	s��R�a���� dz��z��%%�'��3v��=L�����W����:��(�z^�soG (��}*�0	�c�PŠ��y�����e�p �lu����Xu���!	H��.1j� p(�����:.K���ժ�<����̋Ţ&��iGs4(��.���f��+u��~`o0e�z3������wo!����%&�
�Hɠ�v��w=ՙ���ʈ�w|��|��B�ޗ�g�R��녛�;�?ks�� r/����*]!`SNQTU�WL^���D��pf��m�O2�u�|�2�7{�E�s�>�S�au[�|������9����_)�J�BԎ��_�|ck	P,�=Y�r�v���+[����I����6�C�K��K��m6�JVFۑ�irw�^��v=˦�����M�+��E�9wV��%�er2m����:��Yo��o����E0�t��i��aI��#@6|�
�C��-r(�p],�Bď8���x��<2eМ�#�u�����*OiS�`������������|��������,O��@��X#�T��2�DI"'2H��MI�V(T'CW\�����&D�7Ma����G���T�h�i�rO��ݗN]�`f��'�`ʈs�G�F�b��k�l�4v��U,��:^��d-����{K�漠�z"n!�f�d��� َ�V�C��
�# `�B� }~[��l��(��=������/�ǅ���6�>�]� ���yN�s�x ����]�%5�r�?��6�S�$�O�󿺵�MZG�Z���Ct�X�����?j��_Z�y�!�q�k3cJ�� ���IH���_S�.�u��-�ވ8uWz|�A� �"�~P�h��7.A��!L3H,�7�F��[s��.&�SqRV�Q��JR���"�+�;&����9B)�r�{݉��O��Ђ�,:[*�δ��36RF�)oq*'�CV�w-2"�pI���
�޷y�i������~�
P�pqv�g����i�%���(N��f�E�?��JʹQ�����R���,�l��g�M��O��K�QDM�e��?"�(�)�B亂j������Gy憥��]�z��}��nȀ��2��K�.kԣ���Mވľ�_�����u�G~��p���c���c>�L��3�
s+�;jv�eu��л;�ش9�uh��a\c���}�sB��c�Y��	:���G�7k=��*@�TҎ�y�}ԫx��'�X1z(o��~i�͘���V@Zy Hd@	���K��6n�i� �|2�K��;���.��hU�+�Oi���G��kn�C:�G�<	kBk�$4j���c���X�\d�m�ȇ�3x?�[������i�JS�d B	�-�3�*s�5�����h�g��9j]��	˺]��h�B���6�<li�2�=��F��f�'%����\�P����͇"-�a�+RnD�������?��
��r���d>5$WS
�����P��I8�;��EH9<���f�ց�A륃�l����|��a���c�U@û�c�AT �-AD"�ұF �Kw�\�o���z*;{���i���;�'�o�@d�͗|ήH#	�Uj6�j�x�!�)ŕ/�_���*�[F%ֲ6�J��dXW�̷-̒��$��Y���@5D���������ұ�#�&���Lt���-0u�v��[���ţ}\;P��0�R8�3l���{�E�=�S�U�<���T��zA��8C�b!��fzl"J����E�)�2=����Ȕd������&f[խ��g*'f�fa2�ͦ;��̋l�����<�͎oe:��ڸG�k:P���G�˄���	$*q�,����3:@��L�ʡX|S��<,�!>�c��j���ց��xP�qV�Mo�M�J�~��[��K�b��!����� ]쏊�>�֧*�Z��C��!�S����%0�\Y��>�vX܍`AꡬvQ��#q+ѩ\>B˽�>�?op���.0=���-՝��v���s@�;�v�U�8<'.��ߎ�.���.��Jg�,r�V��Hxs8�JC�&����Y˛�����ݵ����9⣲��l�'��uf�fR��i�^KN�Lnq �7��&����	!_e� C$�\��A��<)�s~�)}���c�$v�1�]';�)�;��0���΢$���n�0��m?��~}$��W�nQ��CQZa�A/��-@,��:�
�]2�c%�ùp�ե���7'����|U�6���H���)FA�?�e-р��%�k��X�F�Ja�&�R="x��&_�٭Ĭ������F2� �[��e�P��j�TQ⽾�3}��i	f:G��T�B�+���r��t�B� -l%X8#��ʡ�PqInN�*�>4z�;v��$���v���YLp(ڻ":���C#m۳����+����6����]� �C����~|9��f�p㛚�IGtg�&��^���/�!��7A���-��d��^�ǚ�k;����k���|�ލ�I�Pvm���[��Ф����K6m@�G6�(��&�R)ܯ�㏊�g+�e�!rE��P� NV���9�|ɣ�@ߗ���[h,ѲT(ο�byC�ղ�b�c��,k�3ߜ��2S�'�"/Y{Uq���;-�5{��1�?��G��1\!N2���ZL/��b���P~��Ĵ:��D~�0N��J�`��YZմF.՗�`�ȍ=B<A%������Zնǻ9v��T����y�虬�@�����u�7�)��K�N��f-:����Gp�3 u�^��������E<�k#B���E:]&������~�O�`/�����m�+��+�Z����%P��>ּ�S�]~�*����
/=���bn�ˉS�K9��X��@xX�n��L�y�m2e	�(�M3N�������朻j�cV������T���-�aQ���Y�w6kTX����=1w���Pn!ꀼ��}������[�c1�w#��XuGdeГE�������U���[sɨ��B;�)er*�k)E1m�����1 ���KG��W�Z �����7��Z~]Y�W�Sa
��g�B��G�v]%67wz΍��A��C75힯�Y������`	'��AD��_{��7y���*p��I�Zi�6��Vj�kȌ�X�{O����I�n��b�V^�E���t��N(�}�qz-��4�}0�q._��(Ӄ�ۘ����r��ɼN�"u��1��b綰A��t2t�'7���`0�m!)���sZ��vU$E.C�ぶF-�ѣ��
�U����C���(Aj3�6(��J_����丢�P�R�) �峗�L|TWn�UΉa�!Kpo9�\`Gvü7��m��3s��O�~3��_<����fnRMx�ो�n��I�*M!�z:nN���b���,�a�G�'�)"D��$��55"��������,�_�������2_�(*4��s�)Gc�J@��+	�pm!��"���|IX|�X�'%۶�1.�m\���k�6��[+{�|"E�- t�ffҦ	��|����؀n����{/���F��Y�T���x��9���Ω�ʖ�&#Y<>A��iu�:�;ċP�0�bu{n�*_ٚ��}t��� ��\�u.��fT�2���:����p���e>���<:�;�W���Py�6C�&+��.�Zԋ�C���