��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"�� $WժAi�.����^�r˹��<�G���u�!Vy@f�=��n���y����v�r)�z[��v��L��^p�N�%�yï��PB�<���8ܮg;���r�f��B���ǳ0�bA�$������!O���d\���_�N伈L��|����u�e}�
���ec��d#��d�j7��5]�e���w�G>E`0|qp}b�c;�2)b=��XN$�J�s'�rZ��}��)/T��|	��o}�h2:�զ����Sȿvd���8v:���;��cn���1��$��~;1Nř"���X�����q�B��cE	[ğ�JJiΖu���O��Kn?D	�l�7��g���O~>��4��^Y(��9�ꭀM�Ȯ�놙���4b� � �����3��R�O��^��Aa1ݢ�6�j��,<C@��S���0%[X5�g���1b�i�O@+[vl_IǋR���: ����������o��px��朑fQ-���J_����u�o��C�B�4IG�t�C�IVu�L�ѿ����m������
�i�'���
�Ob�r2�<!m=�H�[���uЏ��9�U"A��P��2Zy�)��L��x ���.q��ԘH��9V2$UW�I��K��4�^�d5�gxM 2��U�lH�����-�"�F��Jc�ѽ.TX��~7���8a�Z##NR�}9�:W�T~�D"t02F��c�M�>���L��N7�0�:9���6��r������a��Oa��l$?�
	��5hC���(F���z1/���^j���>�N����[nu�3p���P�0�2����1�K����NU����� 魱dv���,���a���)?�E����VRv�A�j,�ѱ�y\��A�B��f�ֻԒ�N?�%��89�hv �`��T��Y���J`�\�}w�A���%�}�Y'�象�\S0�'j̜ �#ȡ�|�Ȍ.&��@����*�=sdɀY�w�cem���h���{)����d�>��!���^w)n�%۰r_K���!�;���9��^�yU��,W�������~��Ia$=�Bp�_�`��w�/$���8k�5����^"ϰDq��G��4�<>�l١sէ�v��*� ��7��V%�#���D� `Ю'�RIl��̗FЉ��E�y��t*���?l�-����8���5>�c��dK�q�r��J��(C1A�EՄ����֚�P��%G}��x^SR
���:���t��Xe������!a�3��=��k`�@�,:]���]����o,����P�Ld����I��v(�g�M��/�}5�C���ޔ5��׆��%�����'�M+��_�y��w`##�Zq������̃������I�ݍl���p��Ƕ��g�lswe�n��B�Yyo���SB��'�������L#�V�ۚ����3��c>���5���D���.�y��������f\����K�Q~�:��V;� N��YOt���4A�	v���� 6�㨎�[-��^���G7*E
�Q��o 선�n�@ǑK�