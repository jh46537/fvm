��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)��4��S�C'���Az�V���g�hN�6���~�w��(�,곗�%F�Q鲩+^���t}
$
�o�3r��a�<���j�������+��'� ��w��W(�m#�Ķ@IwK�F��� 2�=�V�;"0�K+j\lb8�F7ZL[1�sY����|gl�Z�Hy�b�uv�m;>�-�=����T�wȜ���������ɤ!��*i�bt�����0���o!����ksF�H~�I�^�"������ƹ.q�d�w2�9�K�r��	aTw�'�m�;��\>����"7��WL#�{b�V�|[p�i�@6�.�mA'+G�>^Eg�. 4���o>b��	
c7a)uA���\�=_�M���a�ԶxB6�S�kJ���uW�0������|��R�c�$c<ʠ�	I;h�{z��k {�ޜ�5|����N�//{!�>zԉ�%8���:�:��Ƞ�B��۩״���DYE@_dL��Q�r٤g����O�. ��F�a����w��d��%!���/o#�����P�YV�X��kr|�ӹ������6�L]V;��ģ������W/�(�����oJ��,1��?=��M�>M]��I����[��3��u�nSug�b�Z�#.�=�\�GB��Y,bgۂd{�h�@���vUu�	�\�:-�\tz�;��:X7��}k���|p�eo&y�_ɖ5��-��w�+��-��9��AK�
������d�73 �1�����;��y*�ۂ�x�$�.�5�����[ku�*����`L�O���~�0�.��80wH���K���~R�0'��:��\�~H3'�/�$�v���N2��Y�jx��[����IT?t�W�R�c�W,`��#�h*���Iwt{|�#����im%�l�h�6�vU�!�^`���`��Q�f\r���84!! W�n\����!�t�NÉ6��@��G���5�{�\p�m��ݽ������n'���Չ.���~ԉ|e!��t������Ǫ�A_�A��j�x*�����6���KTє��T�͍��]��9,4�gC��##C|	�b��xQG]�X�����+_��6�}�KG��@���J���O}��&G7��+��>:wB�j�}�:� 
���w;�-8M���E[,�I���������'�.8�:�W)<�x�?'h@n0#A��N�p��?�����Ӂ�Õ!j]ec��VXu� �	6Zg�6�m��ߌ�@R��J�m]�]o��A�-�&,�[�xLfhtX@�����CTk؃XNux�w�o�`0h���
�)#�l�'q1��%	}H�U�V���Yֆ_�vxT��	Ǘ��V ��Ϋ��jO*���t:�7��j������Z�ͯ&����NK6i<��(oA��%�S�!�m�[<�� �5 ��-�H2��t� ��ӳ��mq���P��A!pz�цha,�ԣ2����|���xj���d�)�MZ�Xȫ�����G�	p�Hq� v	�`�c�q�B���81������<|y�Hd�ղ���%�u���0��ٛb�j�7��N�RD�a���LQ˗�9+�W�۱���Ww��+K_H6,ۃɝ��=�� f�O2}���Ĝ��(����u�T�J�|��� �cF���@^�\SO�46� �7���{�ʷNB|� '9@#	x�T���8�47��:��u���}���L5�z���e.8��h�/�y�nϮ�ۢ��붦�PL��>҆;�אx�����i�NP����%Bw�\Y1�U-��Bqk���W����睨l���F�g�{�v,ٸUdSt��!�,��x��Na���kx�����b������c(�s|�v�-w�j��UA5j�Z�C��B�%k��=�F=��N���z��o��wR-d�a�5v�����s]q�<)����Š��������7_I;a����P���B@�j�UwUP��v�xo
�6N���ܺ�$�d���q�
�F��J���x�<��&jDHӸ�KOe�E��.�Kj;��c����{(��\g��w�^�1��6��H����Ld�D+2�n��_+�}��H��-E_��c#��d�k�!?/���W��Fw���6H&_�s�g�Ko\�;�)U�1
�3Ӌ�����O47�n�	P9��!�����_��38�Rj"9N�@5
���@��p�����C��)�K
��4%ԣ�$ �1��,�@|V�Ѿ�V�g�w�[����������r��(���S�B�u��;�Zb�{�+��˜w����K��)�71h/̏z�4��� �m2.~;���-������t��J����� \�����+�N�]v��j9~���E�O��i=���Vӵ ��IF���[�=��+6��x�
{CB	�]0�c�7��%d6��tB89�G3�����p�rى���BC����9e9��i���@�;zք4S�N����C���@�V
Ů����{�r��^	w[6�v�f҆���$�1vf� }c�[х]J�g�`���J�q���8~�ZT�>���)|_�;i1U&W��q3�Ў������SQ85������Y+�9/�rx��� @����Q+�r'�D��)bSȬ������ܰ�Y�� ^z�aҭ��^�.#�<�Z>��0�.tɮ'��w��su-Q��8��7���#ṡ��54P&l�,L�c�H��]gN�y2b,Aq�P��(ž�_湹��(VxE�c9��[-7������dA��|@v��C�e�x�35U����梀b����e8�&�l1��=Ҡ�/���Q2�ŻT�sL7�9�&mZ37q,���6�3��>t�]��vy��� ?��4n��`�=)�##-\aw!�n �|�7s�-p����Z;�_K�!+�$�d�W��]�:��������:c�V"�<�Ώ����[x����Pq�ti�dd!��[w@�=�T�����;����}��h��w�场5�h�&`e�й�?�К��%6[�R=��7Ϧ��A��:k���z��r�^4polx���p:q�*��ˬ�R���ę���n|�Ж��x���}�e�����K�d�zi���,q��!I�#Z�4l��n��D�&�)�B�1ƛI���\~A�#����	2$�i7GEi �QT�����.u�5T�}�׶&EQ�ޥL�|�dSǫ���67jCL"�KK��w����t�뀸�u�|ږo����ΤhY/��4�� c���m�?O�>r�Qo��rl������_4�q�P����:�J(ɖVCP�o�j#���l��,?��K�2�`���p�D�o�x����7��r��Cu�(�QB3O8ڋ�:�����x��8����W|BXQ"�`���&�G�}WO6�.\䆯���m䶔�W���m���oK@�qӷ�5�`s�����0������9D�R*������eD��J4]*H<ܔ0sv�n{y�;�����L� ��,��y�s���I�f@0C��	6lb/�z�w�܈ӵ�R�6�Y�+;B�*���ڗ�-0s:t�>2=�m:i��Rי���;UȀ��������D�$6��/��0�G���w)U����g���3��6��e�3��y]M����[�����	�e���U�֝�3�����9 (����@���m������;��vR:p��9P�31S�h���!*��5��M�
���`6��ϼ6WCn�i�yY�v�cj�:�����.~њv�t0N��S�#��-yz�ޡ��t!�x'G5 �֠v	��״�T�u�1�^u�e3g,��:���ԖR���:n#�]��*�����]ۻ�Xizd��#�E��&�j�h��Z�2D��/j���v9��O������|�鈡�f�jݞ5~'�?��]����ͫ�_�@H¬�x�;��垵�W�_s6��,!�d�s��+��쵊v��V���$�Q��1�gk e�@=(��~5ڷ$�2K?J��̇�2#�>+}�4�ќw9�g\��w[d��~�=
	9���	U����}��^�KlE��v�)�>�?����o��F�O0?R'{*��N
JC���l�r|�f7(�t{Y��J�oELSۘ����匤#�>(� 	�]珜`�#m�K�r�|��x����F�q��sZ%[�Ϣշ�
 ���~�ʅs]�G�@ƒ�MQ���$����f\Q��G��y(B�>�7���_��"̊�s��t���8)�G��h�O�
P�H!+�^w.��8C�-8�ZMG"�k�Tރ,��~}l�X����WZQ��]ψ�S42�.+���S6���t(31|����J���3��hSV%\�*R���i�mO×�66�m�([� ���T	o-�D���`�M 1'e�0�U�Cb��O����WW��A(�f���=���y�"��~��#ܰ��y��0 <3�-m��8�YM�}$�m��\�Ai����f
��ݍhl���p��˞g�+x	~4{KZۢ���R�*S�~]�������%u��w��+����{����O�?�<[V�	�	�48y�M�ū�EyH�ׁa�������"��c.5s���`� ?��v�����g������<��\��'~S�!�`�k�5C~�;��*�����[��x�&j�N�2/�����KX�s�]�� ���5�
�}���t��,�x��u��yw�5>}d9M�R.�Ej'��+�W���)`�,�(3��
I<59�5K�h��V�����d����==.0V-��A�~�{Do������yڼ�D�F�W�)p�Wo���GN��*L��@��?���0�L�]�nW}��N�����Sz@��i��f��+On�'����	-�kr+,0�vB�&�^4kLO���r�$�K��	���f�U+�w�e%�O�X"/*{x/T_��-���<�5���&x�9�Q]���g긶��a��t;���t�B��E�F���(_��� {����%&h`<0�n1��-�k�g֒���т��k��}�����B�Z`�L1}$i����?��-ڊ����2�+I�GT������Ϧ��vS���9ob�R���*�pa��pL{T�Y8u��"4$�@�P� �5�Ue5������X���/7�.��!��V�;1�I�3���"���Ho"^n�4�>Xͧ4�]�ns�5thiK�s��j��W�{c�E�����$��'���@�u�q�v���������/h	�<E��%
��4v�������l�w`- �+�-8̆��}:i�Mf!wU�OM1�cv��f{��@*0&L�-��GĨ�5��2���&Y�L�u�zZ?H}��D���7�Q�a�c�#=�#A��:����Z�ǒђ+8��r��h(�h�wH�� v���
��Cb78��M�J&��f��8��(�[�/Q�ǀ�`���Վ�af L�._����R[7[݀�l��'��� �%#�+F���� �̿�\h�4kS�)Z3��6��o���;�if�͉��َ��9��&�5Oy��χIk����cr
@]�H��(J���O!r��OD���|n���8Ѩih��%ũsmX�IWB�P�ǅ�/�ҭ>����{����W}�ȓ�;pp��5����P�g`hoe�>P��X��Kك+�"/jS*ZO\� #�*�eis�'�K�J��*��qS��:Z��}�� ��/X@+�n��M��>�qD]�v��(��EW����;�z���%� ��[���ؿ�A;*W�=#Ku�7'M5�����L5����EU%���i�ر0,�[�|er�`��`�^�HjX�]���K"Q��CM���H�$�d���QD=yxϐr������@z��Z�?Xo5<�Bs
�)���E)�Σ��r��+wp�s|3�t�T�X`�9���/�d�=�Q6��3�`M7�j��k��^(���c�~-7��t�9x����9[��������E��pF����V���{���!�9��bWX�-	62k�;D�Vf�~�8��ti8"\�K1�d�$�xy"�i�H�_	��~(���-�Q�;�0��y�1 ����G�:y1k�LʊK3��Es�Ɓ7���X���/�B �Ҽ����2������+�o[�Θ���샗���p�ؗ[B�t)� NZt���J5L�,z�RM���F �o�}�:�|q|=���Q�gii-֯��U�2��|��.>�Cʪ���DWJ��S����A�Ħ��%�%J��5M2չ�k�rV���iq���-�����Nv�=� 
M�:@$b�!��ա�c�Ǿu����Q��&$���r�@Z����c#�͋0=2�;�~�ZG��d��ԭ�|�@)����s�ɸ�K8�A��V�Co��9�,M��tJ1��$��Q���#�f�V�L��4��Ë͌����8-(�f�f6���W�Q�y�W/�V�]z�6��@���5Չ�����2�7YN=�y��4�[���-
{�R�&=Vd<�ك�#�cp6�PuM��,��yT�T\m�۟�vX%"m�@h&�ri/�7m�,�3��ዚ:N��<ē���-�mȇf�w�i}�t��/��F�vh\�7,�������r��(Q i�kIR�c}f͆�.*L���=�c��_�_Ep��y!�"����/�/}�����
f'��F���fP�d��sa����G�6p�g�[s�.������>��������/W�,�������cs���r&	qM�����-.ֻ�E��r��Ԭ�=1�v�xr����Q*��`�A3p-�ƛ�Y��\u1 ����$��d�N��t }܄�T�>�qB�z��@��s><ԫJ�g)|����T�e �� 0:��3>��jl5�.#f��A�����S�����Шm�
B�{T��H������%��S��c&�//M���lf�����!��h����+(^ܻ�8Y,`tK0/HәTK���:�K3,*��L|p��=Y���퇊X7�\Kj�`���[��1�T��(��o��c�6�7Cy�4�ѡ2�N�݀~��H�H눖���}������˛����7�?���vI�N�S:,8!5C�i���J�ҽ0����N1�4i�Q�lu�-T�2�������t��I�?�.ؕ��(�j?q�*��f�D�Ð@��_�|�L��z(���F-�٦*��j���J���<˦:�s���"~��?���:wPǃ	~S��Ј�ܙ�?�^��2`�ˎS:Z߶F�k�p���`��>jL��Q���ۓ�vfxF�=};��@�q����b��6���]=|h�{�4��֥���{u'ux����K7V㷢;v����	`�:-H��ދ��ȧ���5|��3 �C^�ۮ3}>���2	��p���'Fi<\aL�zs ILQu_C�/��Ϝ�{B�[��p"�:3�QY��r��po�W|���i�2q��:��w-�[���'=�p�|o��h`�#0��Q�[�L(�v8����Ǳ#{'�m��8�C(�5�����(Cq��&T�\i������&��^&H}�wa���(x̼��*z��@��M_v�c �Ε]�r$C\p����@"�*��p��-}�4_��K5P�e��@��O�)U�ʎ{W���j^_��o�
�_Ix�G��qZ�nSّ�`A�Ƌ��]g��GmG�|��2d�k,�[�	��.��O��F�X��ȿĿ�Rj��VK�ezS��Y!���]SoЂ=�)�����C�vW��j"� 
�G��<-��ʃO��\��DU��%�Y�@�����>�����7~���t�Q��J�����]� ���"ՓR�d�x-F�u���W�H�1�]a0B�xG�����@QK=��k˔�_"xC4�b�?n��2�����xPAò�=lBJd��w�P�[���Tm|PL�u�)�h������ͫ�T�v��u���A��_Q
7T�섙��[#���8�`=y�͸:}�}<���<���_�;sw��k��T��	�S����Z2��煬E)e����pז�Y{�ϾL%�mP��2��_h�a����`@4���U�沾X��ōH����ĝ;�QM�~J6���y\�L�+���޿$}|܏����W1�����E��-q�]�:�٢���W�s8)(������J��� POp0�>��	���Zf����aj�_�3�r�e����IAL���mRC�9�aV悫cJû� �Q�����B�l��b 3uh�,4����h,%��(�8<n{};FwS0�q�^h䈞A�K񻲦=����nH!57���H�4�Z���6�-�a����(�Xq�4��M�
����[���3=�3S���ێ7�қ2k(A���m>Ƥ���o�w��4�����*�Ӷ��p3O��+���R�V�������.a�hX�l^ׇi�
���YEΓ������t,sCq���i?NnS_��� ��SQ�(�� |D=i$���j}h����9����6�ܗ�d��J!��z��C�L&Ae��T!����?���
�w�vrs�&����+��$����<�D�m�[�P�P�Z��w�3�on#(�J���Q�bˉ�/�8�Y�v��ȸ�eW$	嚅�?�ᩑo%���FJ��n���}g������Q�+�G_�=�ј��?�2��XÊ�
��wfH�ɜ����~�%ƅ"
[xb�+��D�7�p�ձ��g�^Du�(��@�0�2�+^�26S@:�������Vh����V���&�[lN���_ ,؈�V�	r�H�%�b#g��=�,-��̄@8'��n`T��Cz�+U��ҏct&�v[|����^ٜ�tE��a��E�_w��G�]���:\�& �A�:t���F���!O�`ΔQ'=}��1#N[�ќzCJ��o���ݴ"�������'�� Tl	 �M1Ê�������T ���#��ꥐ�G}j����I��&]K�Kζ�?^�<߸Zs<��+�#�6��e̍�"���v�9�iG��6W�<o����c��kZO/DG6ݳ��\�}6E��g5���6��ӏõ��k��*���D7p���z�������T�H�?y��t��h3[���$Q��夹��j���~�,�lC4���ay�^Ԍ�S{l=�O#\��+O>M`���N�ʷf���*Yx&	� 6I(B�������%�gj�����n���cQ5��
f5n;B�N��ׄ��H>�5��
�KǙK#��
a��g �a�`��0B/(/�S�?[�]#�S�`g�:Z � �����>�7�~�˛'t��(z���>�iԕ�t�����$�r���(��-�/7v1�om���x]���"�G�:��z�)��'�O]���U"�{�#'�� ��F�=����j�D?���o��^���bx����[5Z�[f[����P�s��%!�uύ��No,�^���^~+�����y4bU�����k��M��˚�>�A�"��z#ZOJ�]-���^B��h��Q��FQ��IO*b�4���Ƕ�Y�r�Z}�gs!����$�5YP���/@�:�_N��.����q�A����K\!�l�J�b�!���L3Z�:�Hũ>���{y|��M��OZT4��������-LL?G*Nf:Ԅ����\������]A�1/�9
�i,k�R������^h֓�g�}C,���չ+L��S��;�x�ri��b@�:'�8��>���0Љ���4|T;^P���.��n����d�^�wP����1��)l=�zE\�9*jֻ�|����e��͕s�=�cKߖ�,��^Aa)ӫ � ��#�'�����Ӌ
�$�?1�#��L���:}��׆��F��o��VsX�G���?c,/��4ęR"�B��
��r���d�T�f�E��f�r��8F�d���(fQڳO[z�O�s'�ҌA wzl��J���ٿ������k9��.�\�"
l�t����	�_Gw&���K}쮵����4����</�uc�uY�'�48k�Į1��)��aeR��w���R��/߾�Vo4����#t�P��D���<�Bģ���'dx��.��cּ�GoɫI���U��R�87�yl�mH��O��:�}If�丂���s1���Kp@�����_�ɺ�B��6{9�#<%/��~z��}4���!Q!��u��"�d��6�a@*���ۖ���6)�pY��l���p)�$��]H3�����`f>��l���m��*ϒ�a��Y�vW�Z�#��=��7}^��I�,��Y���|����(�H��Yp�5�뭝�ٔ	�;)��B���`�3%�V	��v�]?L�����rr��ǒ��,8.�AiΧ�6��H�H���x��:�q�Ku��b*l�m�N��ޕ�E���]\l��ŵ�x�v����0q'f_�C�+�x;�x�ڮ��/�2s��F��Ȁ���K����N����usN7�oXlFh��@��c@��]�?��T�V�B�#*�!��z�� �[��J�	E�&�!U߀#hK�C���t�s�7�_���%�G�$���|�X�|�@���r:	��:n�y*x��zƿ%a-`���k j�{�ٖPfZf����J��|�Ԕ���J���vݢ�j"�(��v�+��$��ǳϔ1���G���q�@�1¼GO�4�g��[����d�X/��
W��:ȹ��뚖���䜴WFV?�9q��������iH0T�ķ��ű�y�������pŬ�׳L�8ڎCL#����矏�5Pة2����jآ�ˠ�_�����b���a�8�̗�%�!������KCJ��&}��쌼��V�5R����|�~�Hf��TDK��cm�T1#�`�,r��}� o|��D4H�/�1��C*PI���5���IC#�$��j�G��0}�LpY�]�R��=\v}����qʪ�zw���]C���5زf���K�����vsKƹ�@�<�n�
���K�WP������`�	�~$��o�1g@���n:�~׶7��IW#�2q]Î��*h��]ĺ2�e���ם/ll$!s�<N��Ά�\�������a-��sd����H"��m����ҭg���*0#��L�)l="�Kz�`B����M
��`唺��K���$�f�V�l_r��?����hg�fb"����i��o��>L��	���Н���J���fæ�E�$�	>�[AT ��*�}<댵�VpNV}'"ժ
�&��*x�v��?&����a���9�;B�\H�efgw��w\��E��rOT�^8�I!3͜�qZ)y\'CV��wlZ����ڨ^3�wفt!�a]�,��k�䙧8�5�xm����� �7��������}N&����b{s.�yJp�Xnxu�ގ�u'���� �&�'xtNI}5�ܣ�?E4Gn��-ڛ���t�>�	���cRV�5�z��>��ƣ?~hc�9WT���5�nr���1"�ܧ��<� �<{�9uǕ6�_��׭D�H����S����T�H��s��-'8�\C�'����D�{��%Gah%~JWn��%/YO����k�<s��%��r(s�-kx��Jm�!��A�u�������/k?����\1��V��[�����۾�ۦ~�^ O6�}�it���,�(6���`@`r��s\��~緖&5I���9.L��8#?�.�Rm_��������H�T�P;ƌث�W��v<%?��䓰�,N��ߜ� �p�������֢d'�J�L#�CaJk��L.�zk�b����Oj[n/n��P�:�Gpѭ�0sa&Y�%z�?�� lj��Ɩ�k�w{?<�l1���-*�Յ��+=�c3�Tj�_i�] ٲ�y��5���e���$�m����f�pW���� ǧ 57����;�.l��A�
:\� H/��P���U�����W�-��T���\��5�na(۫@��ZnY�4kM�G�m�����G�k���sO�~�f��y]�y�m�q����=a-�|5I��� ��I������b��>y4�9B��-cؕr��Q�� �����|�A�7�,1l��ҏᜉ(��ae%�|���"�{�$�k8�^��uo`3S�]�\�V�8�V{UȾ����HT华ǅ�ݹ�������t���0"�h��͢t흐zD|q��Qɻ���h�?�B�N��a%@�cw|⹢.�S���Ш����9���O%��p�[Q���9��J�Y5�+y��C쳇0/td�J����:Z�*l�n݂����CӬk��W@u.�S�tC�3qX��l�2(���Q6��.�ɜ�`��y~TQ��\�ƞ��Z1!�R������u�Ԃ���7��B m[��	G!��d�gx���ܴ�$��d�(6C�/�����E�'A��ziG�b�Zjn�4�[U�c����i���9�ų�H�C�(�u.!���,�f�G뵳v�f�qoGX�b�7J\t���E�Q���ї�u���韏r]�z����.��.X���Ý0Y{����6�_�qO�=��W�f��Ϭ��-����;�P}��.�G?\I���ap�z�Sڎg��!о-�'�.yW �V�Թ��p��Sʳ����u��G{�P��>ϊo�c!@��ń:G�wk �Դ�ʭd��Pdj�a�R�����e�C�q�~_
lP�>�@2�L@]-h~�>�_A
esx���(���ZL���&���p��%�	�!�S
��<���
���5�]�*����j�E������9�ƋE�h�wq4�!��J �I=���pHAϑ���֑�f��t�c�y'׺.�d�&�j�o��[�EH�	�I�D��n}���%S�#p�N��QT>��]��h䓌QV�I����!��P��?oV��S!�r�i�)���9��"ּ?b:ϐ����l̪;�=������5LkB9qD�?�z�//O9	���A%��㦛��:�,��R�f O����Ĉ��%F��/R���%�	�T����*W�_[/���GumZ����?�׏�k��D���r�$��TS96.�6EM�L�<���H�cVU�l��FQ� �L�l�5f ���^_2�я&B�fJ�5}�:�.V�8��/��5���HO�� ��2�hT����/Z.��.ł�O�f$8���VD�,Ax����(nq��4fݔͽ~hZ�I�2t�!3����z׌Ϡ�������F�
��z�J�I��r�]\��i���0*����F��K5׺V����P���l������r������;oˤ��Cq������a��d��xr��+%93�J���أL�����HZ�JbuI�Fb-b���7�u�����Ǭ> ���	nEe��J��h �g*��+��,=�|2m��#*Q@k���j1������M�SN\k��:Ѥ�?i�$HĢ���cV�s�\�x���Arj��Y3p��07�j|r5��g��a1�,�=Q�����C�H��S'��`e�_����F+y�B���a���_��ϔ���`�{���m��{�7��y3�p~�� ��	c��{ϭ���r\���3�6°<�fPF�����#�l�t�J0V��EGt_5$[>GF�_Lsc��*ŗ��}֔י	,�����(ӝb �f����G')=[J�/���·���~Py� V�\4�[��Ao�VY`l�$_�r������,���/956/�� ���Q��I/L������3*_F�6Ea�O����R���'ӳ�:�}���.8v��%Q�������?��r�癿����x�jp�;l+8��!�3s�ō�N�	u�k9� �>p��������^yY��e%O�Οu��ʕE�p�*~.t�����dL��e<��,_K�5�9^�f�
��a;v,�r+;nQy O��A�C=�Jڇ�G��o���lP���s�W�8�[�z�]w���܃HG��i�əW� ]��hM������P�L���@k�̊�q�uٝ�b5�_�F䆷��w%�+G;�
�c�{UhU�J�4�_�<��7hCĦ՛M�ϴ/"�Ter�j cWTp4��%���G�9�!gh�@����� �3~��qI�� S��\���2�B��v�3s6���:��H�Nˋ��H��U�^��jA#s�d�/����Vy�B���,���_ �L�p��9Nۖ;��y�#U�u���p	l�^U��W����$^�5Z�����&���=��P?= ?�{�w�qi�U��t&����r]�*Rk�D3�XO˲`Q����ޜ�����*(��o�a�k�Q�lj���ڤ�9�0�a���~�)��憎�Ui���r��%�x��­��v�*�n�W ��K)/5�}|�ȭ���g�ӞƲ�u��r�z�ng�.P��ŉaovY�,4ןZ�}���7	f�=���iaD?�\Ι��eC�Lr��ޢ¦����e��⢟�11w���i8K�1�TrN�����x��~?K�9��8�8�yavH�D;���
�B*�4EI�^_�cT�0;?X�t��� ��E�LK�=?7Wȿ�
�b����wS��%Ckr[d�kP��'�{3�WDϓ�}ePA��f��|c�{���o��O�e
y:e3E�l�W߫���>Wxx����/�S����ea�)�d��dޓ��c>��>�<���0�^����4��3H���g�X�h��>Eմ��Dm?�5}k�/�uUx�ǯ���RXx:�K%��0��끶��N��
��I�������n�ǖmߤ���&�,o
�|o�����[� ��]T�܄�v0�d%rK�F#�v�v��K%X��n�Ȼ��Ҋ�����A��a��JW�\��h�:pZM�ه�1�%G�H�2&%R����g���;����6A�c�К�?���0���w<}?�nNWS��t����!�ew!�ݎ����,��փy�(6��=�)���26�Bi�k6r3�T�� >���h��i��O���J)����^�p<x
�4���Ks�KS��p�V~���J�¶�a��B⒀Ր&�,������o*7l����T����q��MO��F,��,@��sp*����626�z"x�h�D����7������!�����,�F(L�Ɨ�u�XcI��$�ƭ�5��&��R���c���I\�n^���\�	��0�Ao���y`�䂀�,�p+��W[!7��Ik޻���;��EJ[��������Sڐ�A�n��/�ߢ�^���q�~1p�-�����VR}��#,q�<J�E�*�>��������e~��+��aኚ�ĶeE��0)ٌ�ِ��JI�O�)���FBF���~��Y��1�뵚3�ǋǇ��鶕ߥ]S�@>k�{�gk<5_3�}�j6�g��欋�
�.����NP���9����N~�A��Sm�<��*(KO�/�Y��+�
��!�̯���{�V���#p�
�~�fV�yR�Z��K���:�&�RkW��pL�뎧9��b�	ŦX��TOP�xRkG2asm��cd�2�N��66{�CM�������'�\��nwWi�6��=����s�ɫ�&�|�s��m ߷�.oU��{����J�u'I�g�/3�X(z`?皩f�(����o��"0�-]��.On�' �ϲ�����K柍-)��^>f��9j�H�]��u3�D��KՍ���j.��!�j"���#M����i��Z�nzh�
�����~՘l�$����|�L��v�ּJzד�#����0�vwy(~yx�V�ap�?����6��!zՆVN�KA�>}��T��*1XA�R��,���,�M�dadT2��8����9F:��
gҳ�ӡ`��W��*��u!?�39W�dc��_}�X����_lZ�飧7�t�L���.K{w�w�� y�z6�Y��]��Hfpe6 f`v%	���I�Sh5*��ʷ��S/����u_j-5#J7�����|�-�N��)�:n��!���%�kȚ��2�+P ؆��� އ�/ޢx�\�	�r�0��N��`~l�0�i��rc1Ɛ�A)�V�G��C-��x����v�y�l>��1m�tC�q,���&�eJ�IH2�h�S��1�x4�jՄ}'����m
b@#�5�:#����8HR�%D���`�J��A�L�)�����O�[M;�`�ߨ�x����5x���Ud��K<aJ���u!d��4V*�pcv����?�E֜&����w�-���;�}�&�h����{��(�,�Gc�<~δs�<f!C3�ʼ�x.2rc^�ǟ�c��Xq����p�������y���x�}p����}����I�
�2h���o򚧦�H�*�B�0)���� ��!�2�4��??��c\�v6�o�S@��־��gjF�!3�[S&R�n��ڸL��h����j��3�����0@3����S���&�ǧJ���x����mح��i�}j�p���pe���W��i0o�"���LA�z*����<%�U݂ey=������6x��nP��?|��_��|wcd���y�?�_���I�#�^."dpc�%#�����P�f��(��+Yj��T��4��� �a�l
���&���qt�:�'9���M��R�N��$�$"
�����%XӘ��|�̅ Z��P�ߧ��v(�XT2s���k���l�d������J!���h�Z�|�*��Ķ�C�s�/��A*�oՊ�W��ᎩS�=٭��֜�/�r|eڈk��,
�OM����u��I�gɈ��Mzp�O9<ǫ��ۑ�<I!	S28�;���{ܔ�r�%�6S��4�R���	-^��f�
�Q�߅ ���ŏ)��=N���Sa\S?-2z���k��9Ǹ��>�*�(J��Y���*�[xޑ{���7P��A�5@S�i��^�����CD��%��:D�o]���7v��vӦ�}.fЋ���&�09PA"Ȳ�a^_X`�o'ߗ�f��،"]MU��ʡ�1�g����ؓc����/q�L�_����m�{�;c�KY�{��=���ʉ��%�F3�!�W� j��刏ס`n�g���QT2�c(�N�\�=�~R�ٮ�j!_$����3XA�l��8�`a�[�y��+y��0�|=�P8���R,��&&��/��j�<dKT��e��ۅ���
�L�V�oǐhu��^�)��)�����E(�IM!0�P����M.�w[��Qô-�h�oƩ�Z���=7�\�GDlر�`p��Q���CXGr��8�עٽ]�F�M�����9�N1��U%��$�d�=2@d����B9̗F�*�
�{k)�Z�	US�2!�% 551�Q��7}�� *�K����`��g0�Ԑ��[���h�������G�Qa�W��oV>�9&@Qі_�胈���Q"s��P% ���&+R�"�<���; ���Q)e�/�[]��:�+_��*�����:0 �4=�Qw_!�4sJ q?A8e
.�3������o��@�g�_�U'����3�(>���
\*ʨ��f�,����F�Y����Y����|��.Uyлd��,��j ڦߨh��g���Ϊ�ǝNWi�o`��j h�*���x��S��)��w�N0����=�l�1(�LPI#��K�9y8;�j(�$��\��ù��ϛ�E��9��L��tv;y��i'uG��u��yߴ�#H_��J_L��m��"+�5S��{jr9�{T�P�������W'���C��T#�)Q����kd��`tX�.b&���!:����p���VznI�xl�����d��hϝͰ��CJЭ�wjjNu���� 78zF����E����M��@E��f��s�+�$�:�QM�v�{����=�(��4^�0���,�b�R�p������o0v�Q�V���!�
-'��F�'ދf�����1pTNC�a�?��0�l�{$-��,�_1#�2�yVj���t�~3��x�#T��Pb��e�p�"�K[�xu8A�?s��IMc���`�Z��籴�T��_���Y���#��f�׃��I3����̾�'ZSNAƓ2��ܬ��C�;��(i9Qb`�Z�H �<p���"��GyT������f��Q��Mt�EJ��v���+9ǈ����Y�����J��̚�k�=�МYҀ�-�G�o)��&V��vt�49q���[]��1P�������X�H�~�����l>��]~� Jh��4�\e�G(�z5��<��*������E��,{�};sƃ��C��l�!���+c���Qo���q�4J�dޖ�['�R+��t��F�/�ы�'q���aQ�Mj/لH�#�	 5G;(�5�eY��
܂ e���61�3:%�o���4��s1~J�r��<ȏ4b��&V^q��� �=�_��a�������㳖Q����w�xb�5�����əA�X��c�.����WP�@X��'��N���- ��|'�hw��߱�Ү�듕��@�H-��⫷(�H�$G�_�*u�~H�!�Z�b�XW(/�C;\�¨�z�娝Gޝ�����ks��u��q�7���$�)<ʬ��A�/R�ɥf�nT��}VU>�j�~Sn:nZ�u����Q��n�yR�>F?-pv6[��f��xyW�0�VD���gz���zm������ў�R�p��.���Nz���q�X^��!�N�����}H�ڮ�A�a��U��f�v�^��u�/ֲF<\n�Ϙ�5�?'��J׈�:���gg:O�f�OaE�E�'�)�6Xp�c��f5��K��հ�����=u�v����$�.����*����E0�:�*�Iqّ[9�����^R_ǲl+khX�,'[X��6\��Vw��B�ԉ�(D��gg���pɆ�J�w��4~3�-׌�km'�=�[-2ET$�����������Sk@T��]�jB���me��諂�d�Gw�ά�:/+L�C`;�6�F@�0�� ������%r��g�>�j�P�makd?Р'/e�NmP��gnh\_�R4�H�����%U�ս�k�߂��p����u�*�R�x2�-?�g�VS5\�>p�
��_q�1��r�q���	'ڍ�H�N����u81@��G;�OBP��Ղŭ��I<�
��p�b�e6��V��8s2�9+	����O�8�G/��B< �r=�"�ԷI����Ѣ��z����
���[��}�oB����(2}��>>
 :Wo!�n�#r3� h�h��p�/�:���Ƕ�n])�?�qȲ{V�z��Cj�[�yY��L�%��^Kvl���%v�u�n�3M�����^�YJ�O;k�~�&�p�A	S�9*�z���	[�Jgc����/#�ɼA=�$9m�x��b���CK�<�e� �%�.ᰩ�	�s?�?�VN�3���s������KS�4�*�/���z�H[�-3q�״��g���E��M8�����K�����~�_W���?@�o�~��F�G��xmЫ5 ;��@D=D"�X�5�L>�� ���c
s^�'�����,v�k��.���i�ct�%�6�N_4��>o'�𤚂���=����0��djO�'w(��++�M�23b�`��p�O�����mF��c.���4Ӽ��C׃[�;ZK��_���`5|-������f
�/9����q¯��M��:���ա��S���^����ښ΂��᠏ˁ_T�з��>7�fhh�yY�ݼ�z�s���AC��7F�S��d0S~�g�9l�\ĥ����#������rd?˶Gy���퓄�/��jB;7J�4j�w�4��;�*�N�hG��Fu�P�{�zǩ;��H�DC�`j����h��"�-�Y&�(g�X�$�P�>]�25o'��f���{i��9!��z�β:|jh�N�
�:�Φ.���Ʈ{��c�f�˖�����`�WM�ر�:b w\P��eN��)z�(m$;�ч_���N~)$�,a���dK'������VnGHj�mi�ѾV̓������%���T��+���57,�v1³��&\���,���ٳ�f�9ɓ_�I�4�����*�ǑnE����	��;�o��m�b/����&T����>q���������M�R�[U=���j��o�2����{Ҷ��c��rT)�zY-�]�W��[��r빌�&�gz��Opcn[�rB���	X@��hh�[�c���3�>X�f%&�\���O4DpG�ei D�]�m��jB��%
rc��Ujz�!E��T�NO�b?�jB����[+k��=�޹�ݓ�*�,���k�>�e�9�g��`��P\P7���#R-�W�(�S����0Y�
���j�I"8;m#aE�r~.*BSƑ�7��%xY�h��-=g�ɑ���Tj{Ҹ;�4�%>zt{M4\�~+�`P�%��4�#L�4���6HV�w^�#��D�+�a�cQAʝ&���_'�a[�R��¥m7�f����R�����Uj�����,��ỹ���+c�D89=�JZ��*�L`�s�1e�
c��i����C>I����.�k�{L�7�`jW���X�f�����2#�� ܝ.ú�*6��q�8c��99n�/����+�*g�G`�@��9Cnp��V���c�v��W�֓�h�_51�s�B�߸zEx��Eo'��c�[���藷��Ga� �X1�b� ���f�.9�{5?e0�zLg�����s�Ӑf���<� *�:��1SDdw����"�QĮ�`��D7��!G�gs����"4���)N�Ԉ�ó6W����w�;Q��~���"W!
"��-\�q�ch�ِ�=�#	������E����g��� �����]�l�;���I5XVi߉2svmO�Q�v�/�Y��Û��Jp���S�<�XOmP�!�/㶍�B�[u��2vC�mq�����=�w�L�� 3�<��$���=��{O��ȧ蚵b�mb�?q�.0|�:o��3Do���HN粎�%�v�Ωa�\|%�34��0��d{R��$FUC�q�MM����F��
�T�|Xͪ���!H������YBe�����r3�3K��1��δ�-����Q� Չ/�������8YW��*�4�Nz���MH��+���S���s_�b�2�a�W�ӮL�ˑ���h��Q��)�����0�VI���8�NI���j[���}|�^�b4��粐'�_]����YP��#EO=�}~�m;�O�+�FB����#�*=:��A����x>bE��3i����Tz�y�G��2�Ɂ���Z�Td���U���+��&�9��^���b�ٰ�µ�1���K���n�r"Av��9Dwbع�QnRj��?/�$z�= $�_�o�q�R��QJ�t���"KȤ�S)���Z�����v�X�i�/�K�y|��X�!H�	��#���D���i����)�X�(s�����1�*սn-OU�s�� ��~"�y'��������xii:Eo%�ޗ1g���T�N(f�JY�N���P���D�$�#ؘ4���<Y�V>���b��v(��/T'����s�eF]�t7��!}hR �u����yH�z5ZΧ�C
�N��`�A"4��@������o�L>W��j�w�G��.� &P�R���p�G��"����7V;�a��.��~>$��bc�p�F���pG�_�}a�r9ǂ;55�;ǯ+�;�rҋm�y��oM{�|D_F�\�z����>�@�ѕ��(�P܋�g}o&`vK��.�'��?McU���L�ڭ
��L�z��"��N<!lڑS��ʬ	����H����m�:����cm/�ѧ�����ne���;J���:&h�Ն����Y�)�4��^����G+���=�[����4�1��5�-�4��r�3LBv��M���]v�֠%���++�u�Vwp�f8���Q�!`��0��cǤ��*l�Й�h�g�����+��hvP��i�z�b�����
�g����*]�h�1:s�,�घ~���k�4���8Ef����HUM��T���T�<*�gO������!t��
0:!��kA��12����C;��ޔ�D��]���ap���w
*�g����8)��g�f曅ݯJ��� 	n3�U��)�D�2�s�ca�ŕ�y�hw��9�m�ݫ��J)��6B�N�i�Ɠ���}�56��i��
�ނ�)���^��杷X��b�W�fև��LXNq F.�r�	�����ΤP�e�̤�_ƞGDU��C�6˄Uģ��Ն�}���|ʑ!g��5� Z�朄B��3��.-��ss��Sg�uT��6փ`&������� ��W�9�o&?qQ�rARGh5G�Fai��v3�Z��͐7u�����F#A�ݫ�K�U%�x��H�G�"�T�7��a��E�%_�C�E?�2���+�%�
�L�T���,��]/G�oq��)N5�mȁI�Z7(^��=��
W�m�K�{C <)µO��#DM��,���Կ��/��β����i �&���"TS�-Y��.?04I(�M�[V�탋�%��C��j(ˀ�M��H�"�t�^�
��H�2��$��J9�r�q�JA��hE1 �&�;N�
���g�2H��VM���Yj7��m�9J�-��?7N0G�B
��6t�oN�e�f�GO7��4O��l�ޑ��!L˜W�+�67N��ƣ�	@��"M�k{P�L�aJ�=�֟g��jjz��������!��e��Q�Ǆ����,�� њ6&���2����2|=O��Ӂ�n\���k�r`��d˗a  :_���_G���L����DO��lj�G9gПr~4TvZz���]!`&Đ�t.��[��$��7=у��e�����p�c�5���Ȟ��r��"S"������y�	�R�S��/�jr��s�IGhG�0�p=�8�9u7U��瞲k<����:�l�#N'�.O��c���D��׃(�m�"�
�[�
��ڐ�k��"(����'�|�@�D�_p��2�'������^܊f�t�As��rO�l�`8@c��%�:enew�η58POA����RYp������ew28�y����q8� �R�e�M�����[V�0*�
�#�4�w�1Wܲuw��5�4JQ*m\e�6�H9>�/Ml��|��s�:;R�j�kD�ˤ�p��M��4����R�f��7�Ng!��Co�8�\),hC���'���ģ���X�KW����Ⱥܨ�W��&9��A3�P��m������9@Q�>ߍ�F���;}	��t	 9N��<��Q&u�L����-Lq��?T�'�M����RiV����uO=� �BR|��:Au"�5΄����.�ü�td��c�&ڮ��Y�N���֭\����������t6���HP��a"��?e�7T��	ʏ��-�^�NI0�"�M���ӄ��E���S;ȫz��?{m�hֹ���պ���
|l�g/�1'�������h�Z���?��v&0�B�0�sj7����yv�B�]�=<~%�g(�/�F]#����%�Y%�)�[����.�ҜA��'A$se�z�%��t[�V~�x�������w;JŬdC���Ok\��A��a��ՓU=v�7��G�l$y��f=� ��s&B&g�u�ϳl��{��0���p�C�1a4X��X����N�R8��\D0�Q��&���c>�|�P�8��)˱����X�?O,��ʡZO��/S�QQ�f��_%�4p�K@I~E6㾳V�b���$��HK4�Q	���B��ȵ*M�
�M4'��K������"z-|q��0%� sp��H�ⴡt�`m}<-�$�t���!l0V�̱O�
�"��j�V��=�J�5K(��]�6
r%�k?�%�Թ�CМ�4O2	�_h�,��u/�]H�AW#j�G�T����ޯ��@	��grGwW;�v�u�n|�&����w8������
�	Cg&�E�,���f�rD�%i��|� 뱀��g���=���0�;:o�Ah�k7��A����IQw̘�$���v����y�i�����>�/)�QUb�y�Jҍ=[嗼�w4�'��k[z���v[�1�o]ZǠ���`
J�U��`��+<�PZFB�y�V�0�4
fܝ>Xr�x��oz�����m����)�*S4Տ��>K�'L�QG���4��o�a��-$�~��H�m�Xd�g�^���a�*����!����G�������3�+l����M7C���h<����+�E/6�=����0��h���>jG&�}Y���+�;�#F���Z�Ͳ�|*!�Q+	6��t%�V<z�U�Y�!���Y9'7y q��
q�s�>j<&��yO���~#�hr�5u��[Y�k��э�nBRb��N~�J;|<����p�ե4���G/���گdEg�4ɛV+q�h�P�h�]�?Q���S�E��y� �s<s�a��L�� �`�d���	�-�ڑ��<�&����2����=Gz�٢�=����;�eIQ��Ax"?+*ǍP_L[O�'������` �7\.����EMj�����- �;1�r��b~Q�CZGhj�6Q�iQA��mKa���ɍ�ښ̫�N����7���f<J��0�Û\�o};� �Ze��]U(x��`�J����b�2�}�������H���X�.��rt�Z���jW��m�R|ZY�D�g�p��j���:������\��^:�H�|�c����U�ɡeZ]��(��s�9��:@��2/�7?!#"o��u�4����]j�?e�[�n���1�WLׅ"���yR�R]#y#bR�	/���8]��V�j��n��w5��ſP�� �+Ch(]�\��P��K���'2(��O�0OXQk��s��})���ăi����V皯�fh�+�}?��x8��=�hH`�:���tJ}�+�o��V�T:���C�鱘�+�5x��mcxx�%(� �E�N�t�Ti�h�2���a�CӸŠ��0"C�C�P��!TT �ƣ��I���9.jU��D��\W��	�C���🽮�3y�V����t��\�i;�s�K89z>=��KO���Q<�amF�48�H��h�N�W����kڵA+H-Z���T}���q��8,_:"ΥF�'��!�*�e�^�x�MT@��|�� �$~����xӦ��1K�$8�9��<=%�E��	$�,C��#6�{'�����<!��F��Ƥ�Ǔ�cR����C��-Q�[fNּ�b���-�rۊ��z��u;pZ�I�+/P(SL-�D�K��:CKȗd�O��u��c�tW�w�5g�Uo���i����Z��:]���,��FIQ3f�ѷ��>���Įa0���c���_��{���F�#�y���?�}� �f��pdۻ����ɖ����6���1^C����PX���^�;M;ړ���bٍ��t,|�Te�y~��� ����lM?�ܙ����q�ҝlƐe�K:������_ȗ��_��z�bHPO�M^6��%}nQ�s��*�\_���"̋��7�+�����=�g�Zc��-Ơ(��J�Z�.��.p7MD�Z����Ma�����I���;!S���0k6�Kk������BIA>���Ϥ` ��G@���'�n�Ns%ř�����r��t��爀U|��P)��Q��R��+��`͓���<:�V�Hnl��k�yO�%@�"]�Aq-)͍*�h�@�P����C�?�ˣA4
 !��vJq��rI�o� g����ls��,Z(������}yD�#w*�-��W'�F�U�z��fv��І�i|������Z&�I5�嬃~5t�rk�pXQ]i��s�-�-�����-hVK�̳�	�Y)�n�U ��z�	1��S�=N ��2JXFj%�#�lh�;�x��"�ᆟ��?��pZ�f� gm������>RO�#u��󫣅�%FL�j�&Z��[���v����J+0E n�v��H�;#_�J$�C,yf�@���QU��A�?��r�eQ���E�{� w�*lb�����9��LA�=X��`���[?��mp ~a`�wv��s���)��Lp�� �89����{�ey�>��@�r�zRp�b�� T��(7?i�YU�~�J�C&�����˷]=5R�U��`N�	�����R�s�ںȇ��|"��?T'x��=JN�]g�ed���������6�L
|pZv�n_�ն��F��[p�s���(��E9�s��E��n��C����������,yx|��`;#�l��Τ|�&�:���S�q�5vH_��9�����������FuI��떒��/�b��=�V���b[W7��{�w��LYd��PQ�d96��WE���e&-4�Aͅ�����x� }gd����L\<��]�����}��s��9��H|�ѵ�YP�����W�{�aX~2���6�;���QV� �qk�V���c	����Α> ~ުM�x�d�t�Ƞ{�ͮ���^���6����=�ͱ}�mpW0�4")$5�����T�"�ֶ���;Q���z�l̏�ҀPw��W��JD]Z\�r��fR�Pe�r����U�װ3������OSy��Z�	�zsI�ӅL	E��.D����p��X�?�gL�}%��`����4�F��"_t�������뢋N�ۢ����l�JXl�n��|Z�H���ە���Z��~�0Kf��T~�7����ze�.w�jO��k\�oc�<��6��=c*��B�{�/+RN��C�Eh�z�c��������Ԩ�s����|:A.ԓ/#�a��&�}� \���nv#��o�5z��xNذn7A���8苹�.�ȗH����'��������nk���Q�A�\�UaI�G�0�>�>F-Ox#�k}�i��{���R1�1~��՝�70�2� �M!��FGk>�A�jE�u�<��Y�P�����0Z�C��[YH4�ļ��ޏk?/�4�'��~�aξD�Z�'�-���T��hl(ڠR�6|N�hEp�U$�{��~�m˭�҇*=ܓ���?&�1��ϣ�����%@�M�a�)�Y�:a��ڻ�X~P���I�soj��*���('��R�O;�,"Kж�xjd M�fm�3�蠃���|�GxbT{�D���`�6�	L:���*6�� ���8�SD&(NS�$�%��p�zV~ٞ)� �bVh�i��fG�@�UC|S�R�[���X	~èN�]�Eh\ky˄��|N�#E[M��6J�1���K�b7�
�yL�<����Է�i�b�&�F�|��˾���mŉ��׹�~��F��H�S�����s��f�D�7�W����)܊B��*]��P���i&��;�	w��{4�^tpUT��l�)� �"�.%#��5r�����{M8n��-�j,0�ozvo�h����Z��8�%_8���M	��Bق����)p���.�K:���_@�4%7�JH̊I�}<C8�{O�=�CǺ���_y�k�R7ݮ+�A��^�J"��8?y�m���.%�q��c'=E�@�wv��K����K=�6'M�B$��Z�,����t��m��'
�>�s�;q�`���ǣb{�ׯ��B�44��v���Q��� �X({OD�Sz
�Q���ěd��a�53SL�g�zwe#A<V�N��$Lm���ID��afw��sE��Jz�I�.�`� E��DK� ;����c$��e;�ݗS)W��TYKY�⽴����جn�<&�J�H�jK�NQ*�
�4B	..����z�
�-t)��n�i���FK���-�W:�[�7��QS_<E_W�mnU�*��d�S"��W�,L݁o��E����uQp^h�|��2����ʀ�$W�R�(,<�I�foL��Ԁ�G��9QF���l��b�nM,"T>���=��a�d+�o�H)�P�|-�4-�R���
ʌ�s��M�XM�J-|��X�U�g��X������MR�`�3r�7�36��5�Ξ�}�Q�q�3%�R�0���������W�"����r۷~ްD����n�
݌�g�t�ؤ��"L=l�(��v!�����	��f,��_�|��;�1��.W��3O����si��H��P� q�����/�F

zA�{J�����F�K��+����}�Z%����p&L���#�Y1E�S�N���f]5���-�3�|Wz��w�,��v���� ����R�;tg����]��'c-Iϝ��� �0ͥ��}m�Mk�,Ń�G���SǛ+K8�U|tK7#���q���9��1"/��/�!e���kÜak��� 1b<Fw�4wVT����I�/�c��lL5���U���{%h����Ra]}5Rʚ��*d=���u,��P�#fw�nI�cZ�%<D�4ʯ���y�@��z�u���C����\F��9��uϦ����)��S��Z�Â42)��op��e9�����ΠJ�Eb�Ӯ��l��N}�By*y	|�8<��,̇���v�#zh�%����5�:��S�i@P���*5A	�ĵK�>]�_�sn�������S�D��7NG�ѿP�x����.%|-��f��E��*+1����ed�8f/���o��]��_���N��xF�ΜoDs���Ћ�s�J+A�ݽ�u�-S���oQ���s�e<=��d�"�����ƿx%5� ك-�?��Wٚ���<��?���r3�S����񢺪PM�A~}�`m��Vą�����py*5��8-��+�nj�K�b�������-��Ҕ�S��*�?�B5�o�[�>ǶU�WC�fg
��_��<�:��4F��� [i^/� �H�S�QGݨCҍc��Ռ���v���W����%���6h,V�8ǉ�H6��#�6IOr<\��X^��kKl�
u7Y��Wtw6�抽`cTo����� ���A�cM�Ů�kQrJ��ߗ} ����Q5��u�T� YeZ�-�!�eE���d���A�M����TY�~Ү�Ԅ0��׏U�r� �wE�
u�̪�]8� ���?���h��m�ʆ���]�]��?���Rg�l���s�(� ���4_t�/o�Ѷ����!�tY�bZ�lQ	̝vPPm,(�����h5@�B�ֵ�F�#�&@�@)�߄A������0�\�kB���պ��w-�<ψ�*V�d����{Йq��Ybg�:�\L����?�
���R�������oC\}�w�U�\$�4�]IC��Ҥ��6�O�F+#��ҋ	���)2���MN�~��ĩ&������!տ���)!<��/=l�;������&�>� F�Y>�m/�x~�/t��ڋ��p�g��q�KL>%<'������7�Db����4������'
c�u�	�����dǨW��ݕ,Gګ��C(�������ovN����J���!��=F�`�1��|��̎ii(b爛�d	%����t�r����'��dӌ�z{_��3�����d������ ��P/}�[}��L'�y�������kI���סP�O�4�!�7���S�$���? V*�9ڝ���.�Ǐv0��`��1���uw��[�@��4Zؕx�6�Od��P�O�ui-Ge =��➃�O�kY�0NFf;`����]�ӷ�q_\��ˮG}}bً}p�W,�6����.�Mg'�ݘ:s�q��C�D��$�5xAU���d�HZcC�H�CY�+&'R�[��8�7�;��)���&���\��>J�LM��~�6�_8�%�$�'��cn�]��
����L�+9��f%���
��8��1� �$R�L_��Ήl���ɧDe�R5W���]4�{B��4�fP9���=j��A��S�}	vl�e�X�)U%�FA�Q��gv���L4���a�C��`vҗo�n�Q�C��9?TP^�v;���Lg-V�������q�A�Y8j��L��ɣ�H��MA�>zl� O�Ny�����kJ�@�ʚ�,�p�!�̯��='=�D�u�G��i"��Qr���h��ɜ��O�>��짵�囖�h�����1W�WZqhʂ&����)�T�p�Cq<�� �g/�3hA��Ȉ�-g�F,�#Ҳ3$���=z��%  oSr|C���B���%���Q0���i\�o�Nf��9��'�ِ�X*��a�}��w�Ԧo�G�qw��h cp���h��y���;���~�eS�K75�����&�L�n�/2�����%7�4�Qp���Lmf7�g������\\���ۣg�{��&$�xJ�����͈a��6��{0?h��kVjAP�Yr��ʰ	e:�՘�Ë�����W�Ƞ|���m�;��������w�D�9��P�C)�;`[&�������ܱ
�"�o�2�ؤ]�����Y�֢��*����qص�if�{�cwM��ʼI��h��9�*���m�Ԓ�ɜJ�8�
�X��W'(���FQw�1��2O~���r�A\�<��
œ�����.�W� ���ˬ����ˊ��Q �M�a)<�9Zpơ/�mL�'q��e��ȗUf��?���"��j��>�y��E�8;�P�� +=s^�i=�.���w:��:�s��G���9�oϲqK��W���^�� A�jL�;_6ۿ�mB�sb8E����
�� �p�s �
2�u���^;�tk���$'��+�/�,���v%���J�c����XP@5	1��q���>9z���u����9��u5�W�}�uR�|U��~��"u��+���9Z��q�E�`�wu~�~I�i�E�TF���Pc�'}��Dˑ)����q�^��iߠU\Ay�a"�peG��i�(Y�BaTC\%�a4oex�G��.�]��Qm�3��U<��V��Q`Z���b�w�P-�
 �$�Q��Ì�Dz�Q%8�k_�G�f;�����6��Lk�X"]w]t�,d8�ۏY9��!�ԓ��N�M����)HL)F�٧�<�%`�mrl�-�:W,'O�=��E��#�
ohoe�޸�W���?�qM�ӎ�>:�H�	/�Ϲ(���qi�=��{�-faZ����n]IRx���ZU��ܺ\	B�
~&�S��n�.w2,��R�;�y�s~�����yPn�5��2F���´�ن��r!�@{����Tw��_~wGt��;���Kn�%��� �g�λP�jz2o���o?[��Ł�9c,~��t �Z (�]6�>�h�K�Pv��77C1I��_�z`�w�ݣK
`�)>1�L:�QZ�����D`M5�I�0 �ʒ��Э�4�/GV�^ϸ�55�[�/�t_ƃ6R���~����ϰ�-;���Z���&����~�3�b<]��\#S���0#�a��5h+�G����p�.�㢀+h�gcVI`�bjoz�}5(�'� �����7��~�Q�r�Ҡ�F
fT,��e}8�+M��5�Y��
� �7�]ԿpU��(^;S`�swM��B�X/�����-�I��#����/�<�������bE�֢��Ψn�d��+��K���8�t��Xw��5�k$$d���8\�~(�'Cu�!ʜ�]�?Z�!�.�1Uh)z��F��kp�{(�=��w�K�$D2J�؄w�{�S�7D<��9GK�	�y��]=d�q����4�= �{��-E^�܇��ۆ�i�u1ܿ3��e�D�;ה׏�L0%��b�|�Y½�٬��"g>����l�C����"���|�'׶T7[������Oa�+��0Z�gh��\��K��*Xg�'�5�����l�^���,�4$ �,̖�i j�Oߤ���8),3��Ut#����"> ��(K�)ǯ,�5A�
K�6-[��$~�.@����l0�A~�Ҷ��f�Ğ�i��.ZEz�KS�]�5|pz�ݪu���٦��ƴ0�k���*��c���=��u���oh�Y�֨��*��uQV,*&�� ��Hg j�+ ��᜿y\Z��>>�x�^g���Ƥ��Q5;��&4Y�|��YDD�@}qr�1:������ڒ4���nx�����������i-�,(�>h�9m&���턇r�ʖ�k|�'�/���b��r瀲�+���p�|C�k=Ix�uT+oB^=Yӓ�n�H�V�~�h��x{�T�r�5�2�Ɗ��7��i�L,g&�X�����%��|c��:mY�`
��
�1�~ň%Vg��5a��Vb+8	�w��U[r�
^<��mX��op�� �G�nC2�'�(��a1�2��b��w�I��[pg�/e�ʐ��7C��!�o1�&�)���˨�y�������h�X����;�e1��xv�f$��g��%�����wv47���o��GD$3#�/�y�"��اV�$��gq~�$BH���W;�Gx�O��7v!M������o`�7#{���y��������8��.S����	�UD��9�/���02���>�?ݏ_�
�<@���	wU��Q@N'ۦ߂����3+�0�!�td9���kѱ/�m!�g
w��]9X�n�Xr�Ze" ��~�Uc��9&��m�����_!K5��G�����9���4�7��2q"�;�`�̚OM���f���kN��XUm~P�Fa�¿1g����=�* y�����ܪ�U9=��z)�^s#GjMۈcf;�)Xj�}�\�3VU�4?ǀ��ĳ��#tLo��`������8��.���N0�2OL����c�|�(d
N(�6!,b6	-�+�$���T��e�L����cLN/T�.�C��f�ym̗9{Q�RR*��g�}��*��_�n�,�۳K+֗�E���
���gN�~)��[M�h\�͝J�t�$���;�r͂\+?!
~q���I|�%��ܭ�S�����f��:�X:�~%�yk�c�ۋ�%�b�n���=� ��ʱD�k��I�8B+('�l`���v�G���\H�weӟٱs|� ձ!���k�����_�(��Ɏ���5���6�&b��Օph��P�i�Q\"���Z��&��S��?Qv:K�J�oN[bu]���r����]�!i?+<�.���I0�B�y�3��/�&xc����m�')YH��`Q�+��]��^�d܂��d<�3�F����/L���%7?���߅�i�C��:: 'r������M�̌�?���Қ���Y��`��Y�@��DN�0·����d���H%ϸb�
v"��m�:�U>��(�L��N������cѰ������v�97L��8c�%�Hn�Z(�bcā.8��Jv�#HE��I(�W��6/W݆*~��_K��K97?_(�)ߢ��7W��<��}|Ot3mp���-�屈�~�7?[�S�Q���_VX]鴢6CF���&9S
*�?�0ʢӤ3�:���.���y��1{�=.!�������ރW�ʾy�#���!y�b�B�i?�#��˱���۟��79�^�~>a�po�����tk0�-��^�n�0GH�w�z�!;N鞗�O��?��L���Y������Ƌ��{(_m	�f������l��K	3>Z�C��1��žL����
i���_��qA�����iv���+��)o�֦0�Ha+�u����?���*+͙6pq���A���KMq�����>Ћ$�K��7f�;=M���.�}�w�y�p�V�J�ڻ�C\H�?x�V_�S�s�A��1�2{/�f�vxLs;Th��8��[�7���pz'�c��s�ڍyը�/�� 6�~������6P�ީ�jL�}^a�U��I�%.�tg�rMOe�?_��^nEl�G>�����M���%6�6g��u�^Zah�K�`�e.^�4J0�2�0:�q��-���=|��t3��"��Ŏ�@����d*�(~z�.�{��M��z0S�v�䡛np�iS �Xr-`I�h3d��mLX
03NƎ� 5㍀G���(���u𼇠��y8_'�G+"��Dy#�t}��8/�}I� ��Tc:��hݚ)"�t�*�&�ң���bTy�"s�̳&����]��V�ul�2^h��R��F���s����Z���/�1������-!�iHQ�96>*]<� Gr�~N�&����t�<�����"�����FL��<,�Vb��*�`N�*�	��@� ���\�#�����M���Qn
w���tk5x��|�xE�!��^��w�PաB\ ��n�������a�QkTܢP8^�Z~��~e�K%���y�Hy���ݧ|��#�>�q#�^��h׸_<!m��-^CB���8���U^�;�H�����H�૵A��o��2��\��(5=���/E���~MMy���-}��¥�u�BЅ��Busg�"�����'t�( ��H��z~xQ�",uZ3>�Гq�.���EZn";����q_�$��A#� r=��4����r�?-�a�Z�$�qy4���H8ң�"�9�s|���Q�`��999�lȆ�~5�NP�Ҕύ�gj_�T-Yy�}@Irq�I��g�XrfK���K��#�@P�a���A|��p^M��	^Y��y<�@+�bK�jR��4�`C�\��iKT��'��}��	�ˈPd8��2����	[AN��Di"���)[H(<jfo�`�T��,��D�9�F�1�G��ZY��NE~�e *Acăo�t�1]`&;A�/{"�N�0�|Ti.�K�j��}�����D�UG9�@@���d�����x��eKۓ�.�nϸ�$akQ��>
�b���5�#�.�,�������U����8-���Hљ�
J�]��^�i�02���ji*Sd^O�'��o�C���KҸ=Ϧ�1����PI�քm޴yуo���Iŀj�"�|���u3;d������ϽU�C��z����4�$�"���X�gş�T����2?��eA׋��[[Δ�Zבo�i�et���p��M���u�L�V<Jyb��'�,�0�=c/��i⽁��
<z?n̰��׺pv���?����㎫��a/�F������쌍���P>�ZJ��I���?��� �YT�mz1��+��K��No�ݸ�=��-�-lh��6�# ��l�J� A�6����J|��
A��2nc��l��Md��l&ڤ6�����!�#�ү��~�e�{�b��� �d�D|X��RρO��J�C</@�x�I��y�W�W�*�Zc�TP Bߟ� �c�_�`���E)��v��SE��⧁"��,�>��[��b����#�6}�!����fK�#��}𬁃�+��ϕ�^Q`̳xO��Xq�7!|�%pRN�֩V�Kn��4r�dXN���S�.���&�LV�4G�H՗���5�@J� ���䀹.if��e��=i}�x5\��8�������0�Lr+Su�@���ШH��b��)CA����KNX?qND	`|Ю���{��a�uV;A]����2ȉ�˼)Dq�֗ߘ�Za�4�p�gBl�����������9��tMr' �Z����}����ω����IJ�ڗ�i^w4�`�SG�]��mN\��ʌ��zw���-�t#���#t���g��x��uIC�(���� ��c;#-=�\�ڽJ0es��3� ���I���z�152��ϴ=�1ܢ0�{��BK\Q���fHge���<G�ͭ0KR�aZ-������%<�&�f+6Y6���u��C�'���gc�0Թ�HFp�ޜ��5)���dr��W����i����a��&D��!+$#�Yg%�d�� ��i�5H���"s��3�瓧07Ƕ?�Ʊe�欉eS�?ht�,���r���!�4h��j�~����V�	[P�]c�%�U�N�݄3��P`���o�`v��j�=�c�m��Ͽ�}�(Ʈ��Tݼ���$���4��,��~�u�d٬��3sD$r =Lo��$���BZ6�ˤ��,{���%��|:[�|�ŏ�8�z�q�S衙�sSڌ��7�k{���K%���b���NA5pw2��?V7��t�}'���r�J%^���$��KE!�l8p��CQ�Tt�z�ƨm���;j��GL��S������+���I�(�[��jd04�� s��l;���1�ځb��'���z���V�\�svf����kLu֒CטQ��9p����#���FKHO.�#�6n�FL��;ʽ2�ǝ(�S�`
�a���5���+��+۪�����ePTl�dʬ�����rbW3+�-�P T^'�u�F�	��P�=Z���S�� m��E0�4�����Y�̌�H��^�r}�#�:GZWh�*7�x��M�"�����x���TAzR�A�4 �l�ڳ��Rͻ���0"�6��|�6ZV�j�W���
�7�K)~Uh�K�C>Z�=��H�A��\�Kb^��29r������t�A�F���k�N,\[��R����R�]y%��5����9�d�5��*�8R�?S�%<WD�Q�{�~f6#r��qG%�q�/j�������g��p�2]���B�C�f,��[#���>	������������9�gt����V���H6s�����%���֜G:�C*W!�� t�`�]ChejX ��7L3q������m`I=M�`��w�dË�2���T��S$%�:_碎��%��omcB?�O�Ǉ�;>m*��@��Q�˹��o�?�,u���M7 �Z��i��j3|jj`)ײY@��j0p�!/�Zuvg�Q��U|����ث%��rMb��ZQ1�%��n���B��\���+�%�=h>���D��J�P_fH)��k
+��.A�B`Ţ��i|َ����4HkҢ�5�,ڝ�8�5���2Loe����y���RgK$�h�q�n b��T���#�b;��
ۥ����Q}IP�h��+?����-n I���"5���#�^6��`�v�=)�����3z�ybn�S]�=}�ǈ��xpW�E�5����y� ��T�q�1�q<v-�����,1��]>���N+���vC�S���*� @3Ú�Fx�7,�({���i���PB�Js{���{,��WA��9��r�hW��Sr`+2�[�����˦�5��^�<{��#I�:'����򼱖6Ю�m:@�w0���ËzG���es��>�͊W�R�P�5�CBX>�`��Jn,uІ^�3�&��j����(�*&�y*��3.��Q.�=���au��EVe֒DR��g��v6�Q��щ�P;�%x�-&���f�Q�GA�X"x� �ǻ<�Ѵ�V�A�� ,�n$����v=8߿���-U� Yn�-X��W�q��K���ⱫnɌlf�Fh�@��-�-/�<�@�r�&H��pm�t��8x�"6��7���&@�<40I�ǡ�\W����u&��:,��HD�ū�"h[o~��և����={�4@�}�c�$���|RkO�t�,L0�ѝfō��/C���U\�5����p�<[���=�c*&��!�m�����b ��9ɩ��A�+���g���uZ���6�
�i��	G	�g�O�x~=/:�N��Ɵ?`��	N��5`�9F����?��\� ���W���xr��P6mf�^V��SQ+���\ �@&�Q��?u	�R�� ���Q��� 6!t+jqA#����W�8ܹ�x��ߞ}$�p
{l�ܷA�7&�qŐGxr��nC}p��RZ�}�]݋��NKؗ�mX�9��yV�X�=��_�Ʈ�i{1���=����]m�f�m�OH	��Ɨb[Bw׷.D; ���7�3��20�T��v��g���X��m&�w|`�D�w�9�_kJ�o]��j�so����̭]@�꾜XU�Wt���C\���6_���ɀ-�U��Acvm�)�;/�-�F��v�6�3��n�����y���9m�;	l�f*�{I�7����c���%�x����B�l�S`���'�!����Mr�81��}����"G��qL8���ԨMőmM�$��UFԎ���9o�<�nt�hէ�)���P���ݑ��� �l`R�,\迪�� _�L�߲�`{OV��Q���4���~���_-��	���B�[�?Ѩ+�����,uY�&*!��Ï���א
K)ѣ����/Dp��@
x��oeݧj�������G��,{@N��/M��S���	4�O��x�`:�+�K�I�%/\-Y���v���C�{'�����Y���\��T|�����|��r��s��D��D4����zi�\MῌtI�MeNŊ*��e��"��1���p5KH���»�ch[�z�V�7�Qf��Z�Z0;�Ȭ��H��/R7p]�&�K9�K<�
�O��S��;U_gE%�i��5��5�X@,E䲡j�H_�Jt�Q"�׿�5�j�Ay)���<qt��:��q�!` _��RF:m�n���v4�'��ǘ�2����1S%M�����D��9��ǯ���5�w+���'��#wArJ\D�Z,!�1�1�V����i��׿H;��	,��������G�<y��²���~:~q��>�\���ϯDv���;	� )�H�	���W������xq#�6���7Á��1[v�co��e�@�7�R`��S��d1�����a鷪|�$ւ�lF��H�[Pŀ����ƴ���0ylY�Cm=��9J�FlG�Sd,�(�]}H�&z��'��x��/a�.�j�D���='���L������S:�l���9~2������}׆�����Fr�M��H9��HY����=�AED��4�R�Z;���#�9��{�4M:�v��NI�T�I���^w�
����bw��&��|�Kis�D�@�F�µkxP��s`�7����?�h&b՝��i��%���@��>�F���m]l��
`�E'�2K�P�7p	f��e.�/m�	�'.��}��ˆ$C��~Ս���w���լ���TF��t�r��nmNV�%q3 ��HF������)��g���{�㖚>�b�e4�3
���m�~�n!�hSr�#�%�jM��G�|wƹ��h2��ɹ�CT���{H�L�v.w�r+�
.��1�%q}w6�'����J�ѝ��X,�qe�V�Q-��Wn$5�<߀V���>��nĩ9�~�REk�����R|R}����6�O�U8R�y�ou������f����Y��ѺS�xF�6k�pb�I�3�9^C��l `���|���dB�8��'g��s�y�ɜ�W�����b�9�@i�U�F��!���v5���V?��A�B3���Q9^ĻS;D��C;[K9�⴩�N=��N�E�|�NG\M�*:��?��_2��n�s�<W-Y�����!�����T��b�J7��F�Nٗ�Wֿz�_�l��:�Sv�#��׏�ɓW�6���Q#�n[�p���]F�J���$!¬Nc
r�MnӁ��T�I_�(i�k7/���[F�߶�|����o+%(m�xj-���E��2��2��4Ǚ�e-���Z4~��� y���޷*"l��_�o��j�g�ܢ�9lLt� �K�05�5����8H��_�7��_1��	�ݚo@�Ŋϲ��%�����@H��nE��DV�>4�����L�*|���[%�p��>�F)w�����Mlq�ݔ.�!J[N����ğ�P�%�i	[͵��%,�!Msp����%�m}r~���ts�jz���	���YU
��J�y���#�uh��m➕��$ދ܃��{J7�Ѐ2�$j�q��'���f�ܭz��TJ�k��� Ӑ�¶��0�p�X��G˲��e�@�),�h�y*�%��1�GL���R��ߐ�I�u߳�nQ/�L�Q��r�=fv�{�!���[E������\#o5�<AClG�e.R�2�Cv�xQ�3�k��~4��7:@|(��U�7"��Cf�h�:8�w��[H�daH3�s�@3��2������pq7n�����p�qJk2t���#"I=t����R��x[�D����-Nˤ�3���vB���\re�8�Π�q��Yt����,��_BQ��u؂��I�W��D��f?n=v�XÄ�xp���5 I=F�z�I��7�0�o�ϋk�J���]z�L���du	�1�'�����ꩳ慅1n^������љUEuDB�����U�h>	GN�xP�hhl����E�jS2�T/4 t�O(3�c'�Ru����i~�:) #τ���_k��1; �x�>'\ƬH�F}��P,�i�f\�Uq�g=�97�׺��ȩ��i�0��3F��=д<:�ZO���=�=^��cHEv9y�+H-��M>�P�Ԑ�s�j@���P���O�����?�L�=n��ϐe`�}�i����QSf���F���nd���pAso�*��E�h����6�4�)�b��%4�O�p�V�����"�L���ZŻ�\���lf�b8�a#@޹H�c���7�uK@�0$ش�G����wq�z��㉸�sф��_W�����g뜊gc���9��B�r�LT��+-2|ņ�l�
����9��?�5A�P��`���/�*���a}y
7©��Y�ͬy{� �5W�k�5�j����8F�i�p�\\-��7t�m��@��y��p� 6ĻxL%m����л-"-e�l�h��
P���T�c���h �|绢pHK��H�w���Rd��?���CMdk�Dc�qO�>;��^�a�����Q;�W��lc�jyݞUԖ2��_D��"eU�B�ns.F~�@Y���)��W��39���|D�V�9��ϊE�Y��F�I��}�s�K�T�5W�ƀ�[?�K�#��'c1����������}ɰ�.e�MD�#���p���\Ʒ��G�\G}��	��@��)Y�2�d�W ��_�� x�G��6��	�������v��&),7Fȭ�'_Or�=�.���k�㶩 �����ļJ%��Lyڬݸ½�8�>�Å�I�{MO�UGJu�#��⽶��(��	� �XS�	��J=�}}D��4`�.���6��D/!)�>�l�L0��x3��ûg���V��2Z��l�4��pH4g����W�ra����;_��]���ܖ����e�{+�X<A��ģ�Xi��������u"y�����Mr�g�p�J�<�`�	b�DF,S�É7�g#���:�q$��]����6 ���㷈���eA	u�k=�XnKZ��u��43B&�q~�����=u�x�79�PEp��JNٺn'�U��}�����?�/a
�	�<�%��M�󜍘�@yy]�I�7"��""��PI����j~�@P$�>c%xB��]jc/��p��6s&�紼xޣy,y�� Z������k#Kn���JB�PM�*zѮ��������P-�*w�<�i��tjo�op}qS&iΪ�R���S��I�O�=2{��5}�T�r�Ϛ�,y!G�}���&��d��b�e��B仍�f]?�*���Rh�f�cӽ�d���l�;���^��Sx][���Q���;�S\��7%�PCT�T�hNg(�s��Z�Uס�����;��
�X�+��1�2j�r�gEu�rU�>m)eBk�"$ʕ�>R�8��/�fߔ�<`���P8yP����%��k�@p#Yl���ݬ�u5;�BY�p����o]��Җ�t<���n����Q��E�lc�>Xq��D��ɣ�Ÿ+�_�6�$���K`��LqG� _�?��|3��I�j��u�&��F5�����/%Zz�h�|>U`u"�;8��B�����(�M���O��:˶[�E1�:�ҕ������<x���ZH���C�D�n��5˒�|��\��1�	[��B/�9����rT
O�����5� q�,U�M�z���j�{����-�M�"��I���������Fh���np�X/���m*�~}���e8+0��!QѴʤq���<6%�@���l�ذ*r�\sn:j�!�\�7�C�a̬[5��0��=�L.䶅�U�E�+�d,V�r_�6��%�g�l���/L�8���e{��
J�.$py��t��9�$,8?�����-#zw��Х�29<k�'����*T{��K� ��э$���2 �b+}V(��콋�Ӑy:bYwS�B#ݨ�Cԥ��R���cM=7ߛl���B���ۛ�/_	Ey����g^%_]_t�Met��{��U�`0u��3r����/�'��/'�����-\�S`E3�jLF5i��g��Y4��"
� �=1N0�~�m�Ǳ_}����A��Y�S�?�:R��]^�L��	C��� X"c���&��5�niMP��y#��֦�X�w"��o$ܺ9D^%hk?�k���B8	_~��t�4Sb���O���éa� F9��Y���l��׮�=9����a����"^`zcR7(q12N����М)D�/T¾�(�p�1�d�n�O�F+���w�~T��Nz�P9�v���-��%��$�<��l_;����j�nx���<[���
���������}����nQ�kr��R�q�	l��(^����4	�5��1Q����k��Ӑ��ƾ��p#�ɭ>6������8E��� ?������ob�����~qz�6>n���������$�;�L��,���P��j�_ea3 #��kv��|?��K"y����Ƅ\fb����'�oץɓ\uR�����0�L�:?���i3�"����lߎ�A1>���^疥6��3���C��c�A����nV-�y)�̪Cx7�;�(����[d��Շg�<8|-SO.в�a=uW�g���2��R��8��_#��6��3��G���L]��'�8��a��Ї'���?�u�1�n��h��C��W�G�V�����1!��m�äy�汯��d^�P�HhY����[�̎�˰�~���}B�v>P��)�
>a�ՙH�y������r.�7^���4��Br�QMmԤ�2�	��/x�u��B}�g�.�'Wζ����*�[:r:������,�'�$��,���]�bRt�~$I	(�=�pߐQ4[Q,�/"I�~$��j*Cpڠ�2գͦ[�Ȳ��}"��R�oK�ik����E,l@�0
n5���yQ��ڜW����?7�Շu݅b��xM��&L�fݞ�6b�+���$�JW*�����!t���L����fO�!T���vh�&Kpd	c�\�Kb.�9��Æ�^Ґ.z '�0�/�}��T/N|E�+��U�|���%��på��rDH�Z|�0 Z'x�p@�(�:���E��x��Vxڛ�^�?���-��G�y��ʠӟ��0��0J��,/������?���[ND�5-<K������<!� -$e*���gy��jiޡ�(T0��_ S��[�0���U?�w������������3�{kX\�\��H��3M�P�������&�"Y�r�>ق%Tq@`m��Q�����kU3M(������rOG��č�TN�2�,�X�؉��ߕ>`@r�S��?��"�脓�B ����x�3����"����t�=a P+���_D����ׄ^7)�����4�+^ �iRע�R�Z]#�y�R��:�V �Ʌ�U8"`r�n�2d�5s�F�}c;ɾ��Ѧ��������k=���::��HO��"�Hc����EЄX�>qG��=ZLZ>V9J�: >~����
/ ]���)�<��� �(�2ۮ-S.	�/dg�N��rCC�����^�'vA�S�J�ж|L�Ѻ�qL��3Wy3��ӊa��!�1�T��ZV�M9�{�����8C�}�*�qK��������	�]�=�B7�Qȳ?��1���T�Z��G`mlGiF�?=��j��]���4��@���r��Ǭ5����b���S��q���;q��l7��8����/iD�;�+8����K�%�
Fs�z{�+<B\2=�J'`�g�4 �~�C\��F뀷 3��,� �!�KĖ2��,顛'�$˼�[�T�>�����J4�,��߿��U�m��t�ޫ:�J�H韛͉/�{�������8�e����?�}΅	FB2Bnt���c�I%��0=�?�H���oz�3/��WI���w��C��*0�vO�/��o���fO�j���	��T3j�'�^:#fWxR��z!���w�S3jQF @��ʝ��i���j>1�!�w�r�XZ��X��#óN.I��*�1�������	h*�'�I�S�� ���h�ߌL��DU��vz�F��Mf7����$q.���zSL4j�o
���BJ}��5�b��̾zߛ��� �3����V�*�ױ��V̍j�w��P�^N�n�oWX��:$�[��ni"U�t��?�0���3���1���q�IÇ�gf�� �sc�O}p�ԯ�xM
��ɘ��m- ������<�'��(Z�������D����X>���n�ܝ}}9�=�s�sC�mUY��ho2�}��<m���[T.,����@�,���B��`�`�4���]3^k蚶�x0���i�!6,Ɏm
��y|o�M��?`��T�CGI�$�x�� �_��R�]��AV����A��׳�����jT���i>�x{Q�8����
g�I;|P�h��~��0\4B�]�O��S?�g�'d��*�ȣ���S��W|�����L5[BI�Yѥg�_�����b�@f+ l7�=ᨦ�8���l.K��m0㼖�ZT�%2�H�.hq[��Ny�tM�眗�7U�6XR�u�X�O)���噑9��&��&$�p;��nܯ(�fG��'᢯y��w�p.Vq��������a�Vh������(�dN�_T�&��nY׼b�6[>"�^}0�i (Ke����eY�y���%=n������/<�v"x�lCB��JqgL��d-��6B��c��[��G�h�%lK�[_&ƿ��M0T׫�&~˿U1��C�^���-!��kU��]P�tC����Z%{�	 �0ϗ�^kWc��	����
ϛI�GJ��Ae�U
(G��&|h�~T�ࡁ����χ�̰�L�W�p�j�1|VF�4�0*�hr+���O3f�EdS�K���T�@�?�[�c�޶+�lN��-��w�(F�?`;�#�#�@��X�ԕ��XG%7��|�U���.�j�*}�Z�G���a�o��+k��=�� ���9	O$z�w���h� *�I/f��u譿A�W�#�Bu:�9��U������c�ښbzJ��h̛;W`��kR�����_��= U��6_,Z5ȍ.j�8���&A8�t
�E�ۊ���&�I���΂���:f�/7';f��ɹYD+=��*3�x����:�����Q[�?1�44��S�"A5��.S/qB1�%711�B���#��̓�+�L�}?#�K�5�Ճ��W��9�~�nƥ�9Ω�c�օŽ�^��� ���������_�b\��5w���WĚb y��]��]���(3�,�v�a�=�㡺�'-LgH@�3�{�UM��"��{`���2���đ�3f�!y����b���&��n9�T�C//;t�ϭc�2��R��!�]���w[�۰72�Ϥ1�p���ѳx�H_U�mꃫ5m�bڥ\�(�}z��3��+��@`Yb0�t]>�n��M�S� ��V�����Xs�Z�'�߽�9��L�eX�W�>���k\0�.&��Xt՘��+i߬�3wg3/@-i�i��hY�P�*��y��1�����\�6Ox"�=��\�M9����_7��hˆ�v���)2��K���S�=�����>a]��1a��4tM�1�=�L�c�%G���
X����}e��: �����5�2k�5>^z�<gL�"�'�WӔ��m��N�c)��,3Κ`0�����
q��rۅ�N,7�N�u�B⦆X��ʕ�{nƻQUB˔����5t�ݶ�e�%��2�j'F�~g�_���\>�C�%`D��7�P,`v`�5(�����ӒVj� O��1�SdlmJh�F.�6-_��Hr����<��k��y�J�������v�4\��Q�I���?hTLF�;�Ru�j%�{0���J�"�a���iF���>J^x��N�;& �������?�Ҁ:\_�@ӏ߱����҇�}�;��N�g'��+�|���<�<���P���#5PKJG�.zc�ɱ1����`oL�c���m�� �;6;�f+1ٛ?*��1���AjPKYi���dt���0���*�������A�)�� �}��p�T+`qe�� ��|M���W�f��,#�c��$ �%��{�Y8��Y6�B�=�K����������r/ڜQmnWfz�|�b�<%9������Y,�W�D$1*7�ō8!�������z0;�*��)ج��#E�
�a݊9�f��V(9��v�SBEQ�}��+��
��O���G�Ͷ'��L`j�8*��]/�����h��l*^�^/Ui�X��G��4|���֎���v�Aw�s7I��S%����Q�bV�!�K� �">�8� �fv���X��m�6w��c�ȁ����`�<�����ɚ�I�6Q��{��$Ot��������Ӆ�&	��h��	x%PљD��h����f	��������M��<)�~�6J�Q)�h��`��(���
�c^g��G�*�P8�r
����q&����8�f�����B3A%��9O� I���P��q~X��-F$I�y�%�G̮�x����(6���Q�]�V�H����F��2ѩx��ǂ��T�u3����t�����>d��1, �@~�<"y����PPWcj��-��7��>��^v*�m��EY�7!N�8���wP�Df�=����[�\ױ^>g���*q)Y�����r���zQ�����BbÕ�k�@Lr�7A���)�!��$챋�����o����n��?idt�v©�H߈���L��I��rg` ���K>>+R�$��_c�[�g��������s������εQUf"�o��/�+y��>>�[l(wX��X�0��ݓ�݃�@�X�Ӧ��|T�����ȳ�?.�sgjTx���X�^Y7���K�Z3��㛰A����ߊ��Wo�Օ�[��Ӟ;� T�.��wJ��50��kjOՈ��{pi�ɭF��<xf�4��Ρ��N��4ɨtW�ĭ`�]�`��+�FS��H�K5�K7:�>.�}v`�!�ը�P��'~-�!l���x��͋J��%�S/\gz���`���*���Rjԥ��m���6J"u�#���C��+p�M��Qh��"*M��S�V�TcE���Uc�2�0*�� �е�����,�얕T't��6;�	�I��y��8١��RA<��)�Xzu�Iř椕�ԯГ�$���Ö����)���^�Zm��mv���l��L(%3`V=�5*g.�����w�3�J�)S�t�M/G'?�<;h_�[E7o/c�Mɪ�#'���.���?1[d��+��C��?G�|U<L�۸�5Ut�_���*� w�(y��2
˷�Lը-��ӨIR�W���٧��?��=��&�ī�ת��U�d%uAw�I͉Qm���)��)`y;j��+�B%e���/ԼO��ɗ�~lX�菵N���V��
N>�����
"_y�D���KA#F.߱�k�mTN��,�'�;�b�,$	��X��*�ԉk=ݷ�D�[�ۆ�t}���ϳM7I�_:gEo���#݅��I����"�֯���L�o1�������z��D([����=Z��@c̀dJUA�����]�Nf4��ޮ!hpg���B1�c�|���=� �e�
͇�p����P���^�Q���� �)zE,��y�(^��o����_r�m�+��/Nu�]�Nk�U���5���E��,�sӭV��a����ݵ�0�~�
4����A&��p�F��:�X721w��5z O	g����3/x��]��㦛m㟪��xq�Td��wQ���[�g2O2qϣ����Lߧb�V ��}���j�
"{i�!^��(��^��i�T�����\��F���eS��3Ib�l(s��q+>����A
�9�ۭr���:ek�{�i���X4���V�%T��Q���R���3�HPz��E�B�g�È4�r����JR�w�+���<��ͥ����T������苪�yg�����������Z��,�ڞZ�SK�;t��dÇ9�\Z� U�����]�n~	�X����iKw-L�`�]���}w�&����f�������.�R�ZٿoU���2�]�����_�n[�=m�h���N3X����>�B^�G�n��o]�f=��$����?P��ʏI|��OS�L��hŤ���`fS�:��Z:��P)����4򦪰QO�9�dk>��?+(��!���N�C�l H��q�<�k,f���ec�
�`Yt,��+��x�
�RD,7��0c�	v(뾲!�HH�sC���9-�vv���Tr�Z$��SG�3#,C�&�Ds�N����g,�&W��dG[����Ai��k��`0�ڏ�j"����-�I���t�y�����5����<�ny֦��Tdv���f-��酣-�{�{�J���
���
X?���NήYg/�RU	j"����zN�Sbp,bE����;D:�O�r�����.�9�.:��>��2�����F��z���n��L����k���c4�(�$
N��@��b<�Mu�hCF�	
2�S�xu	��������A!q�+�fb>�U�]�T~G�<$�W�8F���\gD�۟��1-���CI|��	z�����|���h������-�u�R��95�4�-I�n\F�����},��W�#�;s�L�7'�g����W���̥' ��b�C���Fl0W���\"ɜh`�錉El�v�z^��PP?�--�~V�cǅ�~'[������`i�}�^�u|��U�t`Ӗ�POD�����\/RL�o{�0�E�;���8����;��_YY����%��q�Z���k����ވ�
^�i7�A6�w�"�ޠ���h ��+ɯ�\�����+��DH���)IG�׬�%�	}�;P�i�"��I�rM�r�Z���tK���EA�Z��v:o��T�`��@��������~���jT�k�Ș��_��Jf4ͬ;QvcKė%0�ҷ��,�flկ�r4f>1�� ���V�2�1��`��t�0�^�jRC�t�!�GbH4oژ�[JuɊ�w�,K���g2>Fql�h���)r�w
j�N�Z�1;x�Ы�@��s�h��)��Ȑ�x�^�����0h�D�`G���3;��7�iS[�lٗ}R)a�1�Yu�G[2���I�PQ\ x"%ak:�Zbf)�{���ȸ�m� �{�~i^'��}P�!�ߪ�)���1�<B�k��5�e��T
}�ƌ����������)��x�S�z�_�&�����nT���y���<�d;I	�����)�%	rk��<e�0LM�������M�Q5��i#�ha�v̓KΆ;x�ikVM����c�{��i�v�#��og(y�-��k�ٔ٨:�};Q"�����>�k��:!�V��oa0A0��?��'Rlt6��j�����8����-�Sx`�;�D��|��[�[���gtK$��։|��ۦ����{O�c[�|�{2X@a5��jC�`
� ���C��3vw}`�O�G�!6>����8SR�Jq�vm.��5h��+����f�G,P�7M��6n׫��>�uG!��(�^�G,�Mtd���k�����ws�� �q�c!G�G�~������J�3p��(<�J˃n~#gu+���x�]_Ed��2X`h��^�j���'����a���"%\�T4�K��U�:Ȫ[��A2�TԊц,	�%�����"����}�-����yRdѨ;O r��Z�J�2F"
��
/	�w�]u&�]�-��k0#�����9_���o���������ވ����Mx�V�J�_3�&$�����t��B�010�Y�)�V?sGL��E\	j����3B��SJ' :��DR�QRbmq��cQ���r�P��)�>0G�/�
�� ظ��W�M�h)*�J�,���jq=�ҭ�(�E����t�b��t�c6=���^��N���+)�E� y(��d�U���oU�2䋙��{lǆ��>�J�䅢b�y�4]pc�h"��?���#A����1�\ҕDH� �Ĺ0�������9��"��m�~Q~��rT�`�	���<���7�w䙎����MN	�]��Y��}t9x�LO��W�.���]4a	�L�ZT�9��)v}D��h�Z�Q:��Y6ڝ��<��5�}���N���a�"�?�ط:U`���!�n7�Ҟ���ܠc��X���P~��0ū��l�G3��I�#_6����� �<O���s�;�aS�t d`xN3��i�f[��]��N�4��Iu
�.�=�/WJ��p������1�lU=t�5:���o�8z{@�n><�Io^~ⅻ�Kv���d_{���\F\�7���?O���٨m�Fp�Ua�E��-���W�>��=�s�An��׻���W���J���d�Z��ǭU, 2�4\�6k޻'^-�%3N�6XArĵL�!�Y�!��D �V��>X)ɇ�d�ޟ�c�qR,8kT�ʉ�OϗE7j-��ze��p/F���ۀ�,��S����r��		eEQ���v���$�"�.��9�XTW�R�j��y5D�@�!f�Pj��ϔ��0<%��BQ�Np�����_�����d"��_�N�q�!���P�jUӈ��d�Rɣ�e�T�X&Y2���������p)�m?=��eAPٰ��?�S��(2}	H���ݜo�����Y��AEb
eI�C����r;(�DL+�U)��榤�]M>����ᕪd�!�Y�AT�,�K���s��g�X]�i���A ��������!�Q(ˏ�{���=�A��������s���^��Tլ����ǂ\�m�[*����2��2e���~>�' ���qv�=P؄������1G�Eޏ�,Oh�&�")��9O��s='��h�Mx����Z|�/>L��o�������7�Gny"���z�)�qЌe�`�n�?nܘ��bNr�b���2,��ҏV�V�@���~�6���_(�Z� ��f�����%�՗�Z��,���-�<�ɱ���i�̦ؿ���K��&fp�F}�ۤ%�Ao��|��Uᲇ6�V�sV���<���n_���ו��َ�2_b4�f�� �����Ƥq��#��b���Y�TQ���V��Tُ�WͶ)۔xǛF������]ȸjT��]ʱL|�o��S�!"��W��"퉭���U3�c�@	��!�9�����/1��.fI+xٸGB"��y}?U���Y�����J\����/�O	@�;��٫����aG��~cX�;���b@���ӿ֥@�'�t�<�[�iݸ�*L��c-.8Q�cP�ĳ�e�����{��F`��&�7���#OM�~�q���?�ʶ%��%M@�o:��̔�L̲[��q��{X}�.�O��6������T�̏����K9����������꯲��_�%��W 5�`?TS��L���5�i��2B|�a�ߌҧsW��x�����{=�˖�0MZ��^YLNŋ�Y8����s���\խ�[�v� }�1������V�	c�Q�D�b�=V*3�_K�X�V�T+�l'��$%,9�����/�n�{�-׭�~���j�o�\�#���R�{��
B"?����p�S�~��E�5�z_�c#������NvU!�c]~�mmf_|C1Q��bz��ڰ�w�6͏Zc�V�)����8�>Z#�J��"��`����s�P�U�E� sN����$;[��?��6&n#�*�x�@��c�����c�V�3�OE�Qx�9>?P�A��C��O� <��MW(4.i�^��,�r�%hIfǯ�c�7�g�q���E��
�S��p�1�%�J��������RC�r����e��t����Fs"���(d�2�_��F�����4֎��0P�8����
Ҥ*�����r��kD�g��At�ੳ�M���MQ��4��
�T���*�g���C�RbI����H��e;��l���4d3�,]^L������lq=�Ms��T/���C�T��$�.?t�+�Wk�
eb)�S7�e����n�QmGt����:�rQ��w#���ȾL�C)G�.Ъ��Q�r
�����e�S���΀����S��.'��cqrN<9~N���]:aH���k�;
r��W��Szͼ����T����&��{E�ݰ�?�����˵[�oo��2'�Զu�(f�Z�u�Ђ����Q��0��^>ԥ�>@t"�4 /�1~�A�r�ت�bW�3��a5�;G���̪�A����6�(�Xh�"�OS�C1tr@  ��8��A;=�I��]�<�"�	lO�\��xWDe������w"�/�P)Fl���Z˹��B��N��νbn�[��D!Ur��<&�[?��ۋ�&%M�UY��Ɠ��Ӄ�K� ����ரcsF&�7�5ޏ��v׀�é�"�x��sY��Z'2D߈ރ��:�C��3���\jj@����Ŕ{ҽ����g�u��t}�%��4$��km������x)`����ޜ�K�`��B0����U��|m�]2b1����I�%�6[�S��#'Щ�ԍAP�7>�y�y��P:�5�5����a��6����e8�%{PU�*�?q�4��e�[U��1��PĤ�V�ʶ�6�+f�����GB�w;v�jA4��[���s����O&�'V��UDL�rd�	���̮u ��w���2�ƚ���̡ұ��P�I����gּ{�6���Ε�{i�Ub�Д�o�^��+(��3}R3�05��t"�,r���`L�e'W7���%o��A>6lp4����H��%-�:������~�+��2	�S�WG�Kt'�4;=�}����j��"L:@9���.�K���5x]ſT�]�3��������z�
s^�L_�? b�/7O��jB˚�y��KZ�x��D�s��I��X:��3��������ho�R�hW!gn:�����AJxyt� ���z�0�ٞ8?j~'��زN���;���)�bW�&�HzadW
��Dge����f�p[�D{w��C�f��Q7��q?��zX�������'����+0�����2�.�%���������>@��]��0&��6�������!�ѿ�*�~Wl|o%q+��b�r�4�`�e�C��W���c�MӴ5��(�5�	>S��Б����.�G0@=93��eD���H�`��WP���u��HQ���?�HL#,���xS��DWL��&	�]��L)Ɲ�����*�C���"HOI��*M|X��L�ֻx�x�G�&)p�56y��(\�زmL��?oI�T�3��ݦ$�h_��l qI���k-V����p鍯*�"�Q�O�9ȝ�X�B�-FL萣b[7:W�7�ս_�l�q��ҍ��%��+v��1��R�U�d�ֺ�a���ur�κ9��k���'"��b\{0��,J���K�ұ8����/��N�#�C���<��3�:�{_�������.���	܋��u�%.P�r$6�gI�w��S�J[�ʂ�HO�fO�ML�itR�ź;�A_/���j�*s\�P���#X�w%Ҋ�ze]��f288���ZRm	C�A�VD�!w臠�C�jQh�m��o���T+���v:l��A��Xl�^ �0׼�g��~�n��k��DZT��1B�ԣA��F��#V]�/��I���FK4y|T�+���l2)(y1x�Q摭���"ܑ���3ҏ�\���,��Sܧb_os!��\�?�(�
C/��.y��C��Hiw����a�I��Zz���u4��)rF�ާ����<Q���4��PX���נ�����C�7~?2��)�miZ�"��'����/ͮY7�	1 ��0�&�k�R1]}X�q���i���52u)A�!��$�3���x�u,�����Nx��l�fĪ��b}(Q߱؀kHX9[¶E"Q�����[G)�Mz���m����3���w	�B�0d�CD���(��'������Pu�O�/���дB(�f���!��}}j�Xҧ4*�0�9�8��W	�#G����<���75�k�T�"�"���E��n��<<Gkp�Խ�:�&�g2��x����7�O섖����
X�Y=�M���]@�G����r`��H̷Z�GE�*C��W����F8>�E����(�`єyKp��(��j����(75���h�����vC���TYu�i��s�?m��2�q`ǽ��$�+��e��|���B
��� ��P�}[�h}��r]���$~
�k��`��"+Cx��ڎ��W���zs��G��88,���`~�G�f��ƭ� K�aԫ����>����W\��!_x/��u9#DW2:����1,��D������a������OE�T��ĕrf���ܛ��HY�U6͆VZ���zL�03�P)Pe.��  g���O�K�%�W���K�V�
��5W6NJߔDV�3�A�����+8�\n�@��O���b#7���zV���D,�&'C�r��Й7��/���[�&��L��XH�F�y�`��J�XF�����Ÿ��Vb��ɇ�@��7��'Y���hW����7B�pr}�x�bŨ[A4���D&�N����4��K�M�\���;e
�?6��ג.%C�.`�db;T��Nv�:��['|�/�7��qC�(�`r��Jq��l��|e�*⫵��ܳ�k(�9�&� �j�Q�,��3�[�A�uX�r
	�a��R{�4�,�M*{:��$�q���ql�f�I!L�*�
�Е�xf~Rfu��nO�� 8������\���cj�N���iE� �B�E�>ߙ���\xΛy�$9L�=��W�#q?x�/�o�����u4}��	]wUwCy2b�(�c��F�9QvKҴ����-��if�[p3�6�(�[ʋ�HF�Wnu�'|��b*�`uv�/�;�W_�	!�b��R���<��(�?kO��cɥݗna���1�E������ H�!;��s�q�4�h��&F`h�'̐3�[�%���ywj���Q��py�U S�1l׬Mqڏ�����(�C�dZ1��C��[��Ĵ��ω5�9��j�C2���y8�#�;��n6��H0�`^)h}K��2�� 5x$G����=	�����~F�F�k��+~a$a��k�ҽ��%�ʔ��`h��I{q-�
.^	�o�W5��������Y���ds��;��g�(��7���P���B�}|���H-�пTjr9�H�h�S��0�̷����Z���C#T{���%A�n�-?�g���?�P�6�@�ȋb\d��G���k�&j��ڶg8�0gZ���x��|������n6�|}����?H�շ��ni9.w�c�F_��g�3��&E���������t[I갸/J�5��w��
Sa��ԏld\����_��$��'}�e�"�D8F�Ua���ͳ�����o/���wE|+$Ng4V<�y��n���P�tJ���?����Y+B�jj�n9u��/f�v?�n^2���i3�3�]F�6@��`�m~gf��J�T�Z���1���f�������F��ߛP�$�w�l�wz��nx�ˑ��s���<�������Af���ȴ�Ql�;�Z&�5�EeS	@���≭S:�a!E�MX�l�/z���ߎ�,���ڦ<5�g��Fo��1z���ud�2�"x�(ɹwӉLNk��{'1�����u"v~��F���wL(�h�0.7��	��3.�� n�cT��q7ӥ�|����c��o��u��{I��+�ʉ��ѹ��Rxb�2�(�o��R;Kơۅ����`���N~�3�6(�+�ymm�I�=��q
(�M���V�3����⼹tX�_ܘDu�LWЄ�W9�8�{8�蓭}�b©u�{]�D鶄˽�	~�\}��{ߊ��=��>/�zpI!G�E�TU�2�k��
n������
C�e(0*d6�v9S���R0��o�����V�x�7��=i���ϛ�����eU$(�_vԊ�0vq���+0A�l��^�M�N�y��� �*��݁��6�y^wE�&�t�Fyw�=�\�P!�Z����F�AU%lþ�?&�<@���Yŏ�̨�SUu,��F�\ă1��>d�6b&ݯc�>�Z�#H$]c�v��P�Ce�j[sd���f�G�;��!������%̧g�n�]��Xw4�1�祯0��1f�+�� �	Q*ߘ8~��.�Ef��­�#{��p/Y�\6�ٞq��)��j��Y_�R��E%�;9o����;�OΞ��r�)��Dt���+�&���I�(�ܰ�:� ��Q�;����D�t�D�����@_����w�8�� {���X�:F�<��-�V�_��Ɏ6ى"T��?��<��9�^�<A7��F�_	O��?��u؆�-xwMY��񵀀B��	���LAz_@��߄+x�~b�z�kK�1��*�X�i� �8\(e�����'��oΜ�J�z���J��|�66��a¯zr4�p��.��MO����nR�� �De�때��q����jRL��g��E��� ��!4�_2Tѷ��@Zf} ���?��(콃a��X9��!EË��⤳��8�������~!������.��F5�p��}�+^�]5O���K5`qpZ�}}�A:Z#I�u��苉���M�?�%<I�,�i���6X��r��?�s+g&:f]g;�!Jlc`_�cm#	���dS#��sa��[SܖV���LT�	��4.��������x�'ç܌� !a�}�:"Z>���I&"#3M�^5r�Nɵ�G���v.�*X���u 6�$<@/2E��{�fNn��.?�sQ���4��F�\���DD8�6��)�G!M6�3,�`=����AS�4�]F�5�{�q�ڳi�Iwە�0�(�`ç�6VJȇ��響�D̃M> �FB&�F
[+;CPm��5�U�y��Rmܓ��P�u"CA4?ء�	Y�I|�q�J�q�2s�y�(�Y�ۏ�K����"�&�C�삔�D�uqt6�pFS�0(�����Bֿ�%le\<'��Aٙ�u%���'uQT>�Ytl�FϬV��()�i�:��av�A��L��X�<����`�c�(KV����aG�htSCv�z���d�+L�h��
�1<Ro��4�䖑KQ��G�{K����{��)6X�M�E&8`*���eƜ����,��\����C.���N3J����g�FV��aFI3&�c����Oٮ���R���K:d�F�~ދtM���Ti�O�ɩS��QQlIj��&�(�X�/�t�SИ��ΥZ��� �0Lk��5�q2���Dμ�w:i�P�v�"	��"�4����L���$��C1*�<����[�&��O��:�=
q ���_~�����$UG��#ؾ�Ç[r�(['T����˦�Z��ۇ��xͺ��$ttӖ���̏�-ۿZF��� C�|Lۏ�R��h�.���?��+�e���)d��䔇�CȐ�Ȃ�$[HD�+�������L���J�^�L��:��� }��<Y�]\��&M ;�%@, {{���Խ��Ji^�nTn�@UU^��_H̚�±�5[��|h�����:�)��V��1q��͟U��"0m��.�{^��&.����&��M����'�#m?O.�a��E�ю4����_��{.�SJG�0�d�+'v����#z'/���٠��ݢ~E�E���/D���]`��MN�����3�+�yA�ad��@>��B�I��)�&�%����.Dq[�c����(#.��-�Y�wX����%��S��r&&���b��<�x�(���������C��Ybt%���t	��T���̦}M�~dg�w���ȧET��<�ś
 ���e�u(1�����2��YC]'y�yH�a}]�x��.���2��eٖG�:^��o$2�D���#Z%%�}�䴞R8�*x��M���,f$I	u*0�2;f@,��6V��Y��ԔV�N�$�!�ɞ�]9���ѧ�nhӴ��^��X�n�R�"�:p6K��׎%�%�H]&�ԝ�զK�KEیFj$�,n�,�u�w�k�V��A����ȸU5�2�?	�L��0�ѷn	}���dr3A�Xb�`�#G7r�D�(���Yԩ[~
�b4�H�ȷ��l��2"JɆ�@�o^�n�/�=|F�|�C�HB�~_lN�b�`�d_�t��>�}�,�tS&(��/��E�����-��ј�#8?t��65���o ]�i���X|i�ט���w
�#�߻����sPV��}�q�*��bEt*T��
����ɓM��D�#`�?X�t�9!,����u����tQ:IԲ�B|���,%�'����_�g%4C�d��
��N̟f�@�V�ԗ���G�`С���hMQt�y�m?g�&Im2{6/�iI�!�	t��{����N�mW�ZZ��V��!LB�B��b��?u=8��Ь�F����tD�͜{�2�&��wz\_��1H]w巬��&~�deƇ�1s-�L�+(J�m�E;�k�E�[q"wG?��/+�{S�	��0F���� �[8 ]x��O���w���1��'��8�wȅ�`�=r�	*��.�@֟�Z�/�>#w�ϧ�����E�+�[5YS�\��Ij6�+ҏ����ZB����5b������9銑o8�%�N!�C�%��z���b��6{�N��<aG˘�f}{�c��v(Ɨ�|��C����"�����S9��b��>�d�&�����԰XT�J�(#��W��vg ���f��v�W���S���L��i��Í��͵�²r�~��
�@ocBY���ު}W���A��(���BT}[��Mu�X_D��Z|O�fRgT��Q�j_m�>�:���S�ڂ��\�Ӧ��e�K��&�F)�`�	s���9�0[���p�h��+K�b��;�ד܁�x�5XE���f��Tx���ߡ��� eϤ%l>�n�[�����;%�9ъ����>r�&A���V�Ա��;���Ҋ��z|�֛̜�Ɠ&W�z�����:FSO�å75sROSE�
�RwT��U�)��o'�QW���n"�E~�X���F~(H}�쬑�f���&���&2�H���xHmWa����40�ȷq�s]�Qǔ��dN��0|~b��r^�pE��z�6|g�
Lhڣ{��}�^J�m����������2i�G�l�2ձ��k��8Ǐ���A���l��-J?:ZfJ�T;�}�QP��-�b�@�x��M���U��rԂ���䰱�w���b�[iԫ�W���c ி��?�=@�8�t�*������{s�R�|f��[���]��7L����ؕ>��E̘J�P-����d�Q��4��F�	�)��:D�m�!���2��1 ^�j��#�!��浐{yp�N"�x!��p��\`�)�*ʤ�|��,�`��щz%�|�Yig��'7q�67��W�
��43�r����7�w�?o���Kq��Ö���C[��.����JRf)m;�1',�2�f\�B��k/�����pD���؀���Sy��v. �9�+�0�k�����`/#���F��#��_���ӑ�T��,�����3�^1�(;	^
�(��`�@���1^�L�T[�үZ�i@8�*n�J����?a��D����ۜ_�98U�=����Y�a�h�5��E��^겼��L��xq_-H��Zb�l7<C
&GL1���"U�Np���5鸼�$�� ��
�����}W�Y���ĆwJ�]��[��f�̂��9f�i���CDȫ�f���0J"i��l�@d�ɿ��G��@϶v�u$�x���%W��,�ï��z`�������?�2��"����F��c�HH�m�y���E'k��͓߱/�HJ.Z���V���3��p�b���A�)����
�˶�Z�kõi��� ~l�CR�i�C�b�&:IX({xn�6��ytt����a���\~�r'\W�
�_o�4���{�զ9��c���BI��9<ѤuX�p%)��O����os�<s��=�/��}��uu�u������&~�z��Sdy��Vfd;y��Z��y޷ȝ�R�xE�&9�:�� |�{SO�zZQ �?��K�x����r�U2��*u�^$���%��)r]�tZD�D)ye<(K�>�ޙ��Z,W,SFX�D3�)�6�O���A�~ �s��9�AN��]�]vI�\R3��l�[AZ-��l�J��p�9l# ��;�(f����.9��&��C�F�>��`�� ��"@��]AJ����3�]����W��L)�ݺ�8�~x|��^���%+�q�!�=�A��}C��$H����ݠl"����3�u"��0c���Bc�i��rWT�����(dKME��TI�N�[�Y�p�P��a���\�Ŝ��,~4��`��0)ƙ�=������}[Pg+�9WoPs
��K��e����O�i2��xP�JSY�N�2�����K�/��"LB
�(p?�1�oơem'��vn��8�s�4� �f-:�A�m����jQ����f������օ#�;��'��Yʏ��٦�
H�j@����3�V�~F�į�*�;3�mC^�h�G�S���{�>QS����#��%��y���\�����q���p��S�y2'�����WT H�GyB��zQ����'j���Rtc}s����}���dh�;�	?L�Cy��O/#�ޯ��(�埖������S�mN���מߴۑ�C�l߇LrCڗ�8v�3������	��b�_�;?� v٨��������n����짿�]e���h���9�.aĕ+��T�����Y���jK�K��z��K��9�Sq0��,�+	��1{�qJ���k�������1��J�7+��^C�o� �?�(��*#���4�C�x=�ӳ#&����m&!�+�2xR*l���5��W-���[%�&�}#��y'$UltC	ּS�B�:�+ZPL�W{&���Ƚ�^�b�N�5@	̈́RL<���̩嘹̰�LA�i�1F���!Sm{xpn�=�J��r�<Bx���{�T��d}�����1���A���Ar�?-�%5?��"A|�6�F��Q�y^�wZ����y2V�8e�w�\R'V!� 7q	s"$�]�0q�F��m�U�@>��%Qv4#f����%J��9@�V&=���co�ŝ���4
p�/�H��r�v��L@I�V�p�fr�"��'oz��j'"#����P6�5��@��k͏Q�%�t_2�@}�U�tDȊ�G!G�.R������2.ł�+����0En�+?���д`��qn�.��d�@*�&4�n*P�]!��]!��P�]r^�6 ������s��J�J�����N.��ʄ\������
*���L�	@��(��wwv��1g��"�4%��<{im^�-�<Q���*S������$�#�c�aTHM�T�π����2��Q��q��<nYcY�~�go�؅�a����81�������,ĚL������x�ve0�����]�ם42��
��<�j�F�s�c�d��'���6�ev@-!�|鞊��$�{Ϟ�OÇ�7�����H"@�n?�\L�X6Z3������Q�ae�]!՟9��%�mG�6B��-���� �ȿ
�Q�Ddvo^h��7*[`���g�o�|��b������"&�I�z�U�����C.*��F՟��D�汘i���;�/r�3���̰(���U_�����p˭�ܫ��I���1.�C�ĕ�)�i}��Q���~�!�{�&�/���2��@7O�1�=���w~}��*R�P7�l�8���3����HW���b�:��A�Y�����[A�[��.���S�ڰ5�߁���c�S�c����#�t>��j��i=1�ua��?�c���Y1��`{��?.�2�31��F����JNF/d��9-"<�r�Q�#'@����q7!��
����o�a�d�����́tꘊ8�)���fNEey��^�s(��M��'��UU�B!���M�k	���\uԞƱ~���pcU683F����N�rb���v�Ȋ
��qsfT�ni����&�g/�b��f��
����������Z�5Ꜭ���ǡ�I�V�F��|����(g"�E��F��:����_�U@�#�"�zo���5�AC
��7�>6A�m�IwęYή�Ux�cR�����C&����eT��Q���hϑB2� ��Y6��P�>�>��ⷅ�Q_:��j��XB8�������~�~�[J1�Yފ���j�q!�.4Z�!�Zc7�G������a�iy���"��A��16�"����dQ��|~�F��)7�s�&֐�+ERB�ARz3ǣƬ7B��+A�@ۚ�_�CD��&c�q�F(�p w7�~���AB����2}����_�
!uΟ䑦v�Xr�0����@��! */�����x�}8Z�Oɝ��� ��;�U��?�5?քW���V��gT��hb� �|��
xǫX)hOa�G҂���8O�W��t���I�[��&��mpP�q�j.��rF�0;�$S��m�wCW���S��â��&W�x�J���"��Ȃ]�D.�_��,����b~������vuE�p��E�iU-Y9��b�=�7��rf��A�pWO�C�yϰHl�'�g�z��~�D���z ��b���6R�7�>���㋯dZH��=��+�"��@@S9��@r�}�vņWi-:�`i%�F��+dB�#H�U%�e�Jv��5ЊU���u�-ҙ�Ҷ�b�$�-�`"�,Fw�ؠPO��ʵf#�}%���(M��x��&R9�u�&��&�;Ϝ�!	�+�[�o�,��m_�����T��e9^<lU���t���[]�XK����L�>���^A��B��{3���[_?����m���'z*jN�)�{�y�o��A�.� t�D1�oT���U�O�L}9�X��(�M���+��I��U��m�(�vN��wn0b����+�®��[W�X�]_�Zi"C�����'i�����j8B��'v��"
X��,�n�\�No�	:B��q��1:�T��M+�6�}*.�a1j8��X��_������Q���=C�۳(�#�bk2"~�m3(�9����ٜ�u-Nm#��.t\[�)��\�Ϳ$�f��/������X�k:ӳ`��a�E��maC���͘�2�o��	fP��R�@R�s�<���T��Ew�2?�}g��#_/��޻��鑼��t�� �ޟA��Ej��4�;D���Q��gmr�x2��\
����^�Ͽ��>>�ᅅ�@44y�~���A���� �<UܢK`�l���~���uZ�O�3�BR�/�lu�p�\��{�ƬCux��y�:�k�͞H����w��\��"=��t����?��ƻ�w���}z���"�X3)d�97���+]��ʔq��"9��K6:|��s ��f�����4�c���E�q�J�ҍ�z�ً�J׈ϰF	�l.�4�@j��ʩ#Y�LAg�|Dz3�kP��xo/�g�fKow1?�����~Le%�x�J�脷�
JLY�0$���t�g�Ԭ5�,#���t�{+�Cſ�9A�1��$D�ts�|��DV��.�nG��F����M��,X��e��C&��>��.!'�� �v�:�O��{=t�HTxp���f��նw�>!8*gW>���Yto����t^�6�g�Mm๤3⫡��e��-fS6��}���@�b[�,�B`�1Q�_��5Ei����(~�Fc��s����c�9������l!�q�`̛h~��
�I��O�6�E
5����^ȹ�b/TN�?�5#�����#~�|�<XT���+���c�5�AO�N%��x��i)�?	j�2O�"J{�3a��*�������r�ڋ��b5���2��b��.'n�j�g���U����)�|V�&�.����.O�ĳ�ƕ�|A�&�u��!��r�ٖ��D���v�Ę)�a��!"V����ͯ��R�DT���J�˳��	Ecb�iA{�磙ȵ�?A��R�I!&�9sk���sM��7&Po8q��R��!�\��=�� ���T���X����Gk���1��H>|�鈫�Ȉ����ߚ�.�FV`n ����
H�7�Q4�|���ڸ>_������:��zɕ���Zjz1��HB�l\��$���hY�˪�5)&.�����V��ǔ-Qӵ��/���ߊb�b	�_aT/��wq�U��)�lZІ�fH��}��������tE������ ���\��ĸ\X���E?� 5�%8,��8�m�L��!�ĝ����a�#��Re��䉳��N�y��g���/��=�'�i���13o�	7�/��n�φ�FM�;���ݫ�dD{��u�䈕Ԧ���nѩ̄�^oD"�F��{.7�.G�%m�ȋGw�#Qu�tȪWw&xoqre���2�$��@ۭV��1�X�}U_v����؉�|�h�H����s�]k�,^�GI�`�����)a��:;�0�}�!�gV���]�l���/N��)S?�;-��U5 M�	��sek�M]6���)��Y��d9�Z�Y���!u~Პ(��$`��閱�����؅��x:̤c֮Kӳ�D�!/��jUo2�y�:q^���6��>�A�Ùf�5/j���'-��f>q���x�ʹ�%o`�|!��	�]��_�kռW�z��r�oD�h~P.2��-^ҊE%���d_�s M�<�sJ����+�Jb�xC��r(�/��<�k���n��g� �����{��wʜ���^}�$t0a��؏�Tq��#F���ɛ�O8If�6I�7U}����"9���D[%�0�����y,�j����I�1�H-�V�m��3~f l���J�c�G!����`�T��y],�㞡�l\O�|s�.���{Xj�}%�����*�XB�o�L�%�p!<�]�4�gl2ytYX�"�_�6)̼i�|@��l��{��Q� ����[�m�g�O:���r��� 6R��l�`��QE�e'�L|r�nO^���|�����`57|�M�I���b���T�{���k���팢txj�o�����[d1�5nS�`9]��*][6Xp�m[b�ÿ�JhG��c����[(&�v8B<b����y>Ap��*�r�3���0��|��=�CTR'l��~���� ^���������>B���r�H^�0�OlU���`tC8)��_\"L�Q+�X�G|0IOM�lO�?�
�3I��&�����A�BV�N	[=\���?� ��6G֬g�B,Ӗ���u�Y, �Y��k\v�6>���X*47��W���3b��nn�X��M>�/%ג!�ǷB�a�pUF�a�A��5��؞}�2���Y	'���
g��ޡK;0��W�LpS�B��-#6x����<�f�.E^��=��F� K(���$�� ��G��H�N�,N�m��бI��䤶vWP?�[������E= F�x6XK�����ݲJΤ@@#l�v�S��
�����v7d�g��ΓHk����O2�~F�>|)LU�u�%��t��������`��Ҫ"z�x�KTJY#�\Y��>N���z�4��v�m����	�(Q=�#�=�5xɤY�qM��1�I�P��_����Y��6s���!WE��"�Cv�w���b;����?������,�?�Go�)i�R�JT��-N���'�wJ�)���i�!ވ�O�jH��~r�!f5��^fѺ��qVt]Q�]�,�+a:\u7Xx\w��W�o�a�ՓY5�D�A_����}�+��E
Dֲ�B� ��t_%?�n�q���{���߀�+��{����v]����ꁇ���F�R��FZ��{:�{��J�j�k_��T]�Qj��]����ŔBݝ�k9�g����aY�g���P���S����0q0w/dQ�[@����|g�9��i����]L��I�Z��7[w��j�Ӈ2Ґ녈�{��ҠMҸ���ųB�F���I�;���R�������E��<��g��gk�޳�o�QH\�'r:�04�>�c��?�zK��BU%�pY(�٠���:�Ї�5�%z�D閭��j�{���h���.�CY��9LnWr)�,VJ�JU -$���{U@�$�֘�|#�[֣M1��G��.c�\c�GRt>�J4]`��]�� ��"7�k�E1��'��.~_��d4�D�09�0�'�����mXq�����7���p:��ޘ�qޭ8ќuH~Fz��}�(�10�2�S�� |����ǔ� <q�������w�6Qy%�.��Y�����qF����7!J���u��2��Yl�̧�)� mɲ��i��>�F����1��"���e�����'\��"U��O�Բ�9�;��7�+�~�\IVjS��#6��(m���������Y�7��Vl��W���(AJm�VYY�-A���q�⯱��-D��x�KbF���}rGz~�2Gk:S��� �е��G���t�ڬ����3�q���^�V�X)�?¯�|d����Gw��z~'��LPq���5I���?7P&�4Wا�-�h�!�joD=�a�T3z2��ڗ���w�`)$-*6ƌ���4j@!��%ǀ&K��{:G�V���2�������y
 ���i|"Ť	q�Ā�?�ϖUS�������	Y�,H�?�Ǩn��/k<�cW�p�"O�W})��Ve�u������ٷk`�rT;���wi�ᙔ	�XHFu��I�C�� %��lO����n�\LI�@�l��_W
b@"�N���v��+�_�f�N4j���*N5ZD�ʄ��!����5]JH��uF򦽕�!�2��z�'�t��b�k�s��+;g͇��hA�&B32�Q���l>U��P�/���d:8�8=��>��>V��`�X����R] �RMʯ�҂6ʍ{����a�G{K���?-��j��J�b�^�w�8�������$_��wrŠ6 GP�3r)��o��XZ�i�况��c��0�#�+��W������73��)���.D8x�E�܅Q)��Y.>��槟?���2�t���X3���?:@�x!/TO-)N7@��>`���s�7�zZ�w��0��WC܇?���!�d_�-�y�a藇�-A`2
r���z��N���.���c�!��-�^`�=�Q��P�L�J5xõ����1»<$2dI�Mr�su�����,���ޕ]�y��QբP6.2کV$~��|���֚X�㱥�8�_M��g��>�����)Ez��;/x�g��нMx0Q @��v��^;>-���&��֏��V��P���8pbC����>���2���<1��V� گ�|��K�F���a�p��8`r*IN&�m��BI/�4Յ�񥶉.�*��ski�v���?$n|8k)vRP��K��_�:E��_D�����\J�85��dy�����q�p��-�błI�4T���$�y���\C=ɬ^Z4�ˌ=��/���f�ϔ��bL)�7�s|g��1�]�Cx����LgR�\h��3� ���P7�/K`I8�܁��T�.�X�0"U�$l��@S��n���e��l�i�쐫���,�TMu|>�Ov=�0)����pS��Nk�P\��RCe���Jopi�}����a��1b��Vz[�H"o�R"�D��X�%h;�kՎ�w ;j�Xn�$S���S%NQ�*���ZVp�m�bja�#�
�=���0]�a�ݖp�X}�$���[|g����ڋ�8nc�i&���P�[G{P�Wk�������Pp��a?�l�O}�ȅIU�&�^!��OL�W3i &���˥Q���&�>��='	-�#�'�el�r�3cVFϰ0�^,�wUt��W.��B+�4�0�n�ro�C�^�V�v�횛��[�'�u��Yu3��Qu�?U?�#Q��;��y��.|��6W?"֭� m+�ym�Ts�,�c;�u��~s��[T�އV���g��gG#��/�r�J�7���b�IƏ�{�C}�!G� [ƍ�;=�.]Vd��>td�K��P�:�`1��,�b�z���<� M��\�N��,T������,���q��+��-F��5��H󣁇93%=.ja����2�]�C,ri}�t/ɯ����'ǅ !�ꢜ�Q:��q;��i��?��2����g�SR���9�)W'Ê��o�m~dFo<���p[ҝ?��w� ��҆qa�F�pޓ����uP���.�r��G� (��X��r՗�K
�d=K��F(͉?DX����9l�AШ1/�}T�0�M�v3{N2���NO���$J����q��"y�g�q���ЪЋd�G�Q������$�3}�^S�*���v�eSr�y8Qs�cf�H���5��f�G��Qrd�l���"r���.��ש��a�r^&!%p1�F�e.�.����&w]�A���\�C�A������e��nЏ�����`L��t���ٗ�R�����?ݡ�����J�\)����-qH�|<�# ٴwIcEO�c+c9;�?X_�OCb|�(w�!��������G�}T��W���On��}K���r�5Z��u+Vm��?��'m7�.��^�G�[����1x������4?	w:T�����k��5�����Be��څ�g���:"�b0���
l��n·J�J�@�]�Y0H��`>�Y��"�-�;�UJl&���mwm�oM��D�_T�I$�ٯ[sx��x�Ǫ���[LU���9�� ��v�G�t �hN�*޿f�pQQ�������[-�(`�C���5_\��tYvԅ ��ix]W���@��� ���a��j-���କHG�WG}h����D_Vӳ(����ʧ��;��.T��[gy�n
e�Q�Fq�F.��ؠ[�f�>;�N�]7;O-g��ifiŬ�ߥ���Fd�pZ�O��'~�wJ*t XV T;e���Ǭ/4��w%%��a�龜�~t�m��^�[	&�c��%Щ��'y��2ڵH�0�@���&�᳝��'��T�����������%�d�}a��q�����D�$�����v�#���3,�-d]M]�Tp�����l~P'H�ǔZA6����B��3�#�5��D���a���W(�s͘��K0By�A��=����G�����.����un�iȆn������"uCā]��k�e���r}�O�����[�,l?DESa��QK��fsM�u����S� I(V��O�(��K �#چɈ�_[�aW����`���?������3_��g�*7A|�,��=?�y'��~	KVU���m]�埤�:"c�3&�t���Bկ@��ov5��M\!5�*x-� �\4( ����Oo.�c3�a�")t���;#K���:��c�	.��T�֖�����b?��+�3/�l�G8��P��}hMW(
H15�# �&	�CV�-��q`�l��hn����pŐ;!XY�ni<�����Wkċw�['.�
�Xn���h�?4&��ټ�+)+�	��ȽX��V��t��O�g�z����Ѩ�5ED��%���A �����2q��z�
�����;����W��w~)m��Xq��0������4�n�n��*ds���'���[*� ����H���Q-mXb��N�������w(��/�'�+	T�����g���Z���Ì����!��j�%c;���)ۖ�c`��{��3�����KV����I��4��>�%�k�wWu�e}���[
$`7����-����ܱy�!;ĕl��;��Ƀz�Ґ�dI>��B=�L�5��
�&��)]�6NM�9Q�z
���^��ե�r:��N���ݕ:�g��ݣ;�Q��r��d���>���[��
�b?�_�4n7?�r8��S��c����'Tq�A�A�s���&�!p�7^�?Ԧ�����w���Z�}j�� ��r1�a*��A3z�>u�E�{�	ΰZ���A&��nV6�x�'���a��M�x�H��Փ5i���)�Ѧ�,y��.(�u�ϫ��+�]IY�E�TLe�~˓mQ�k0�V����%}&�����\�E��J	
����[a�
�?jR'���)�	J�<�z�N$t���-#�o��߿dlz��ޯ�v��\N�3CJ�ߘ������������ƀ��{��0L<^��vp(�I���_�>��I�j��!}s�56u�sp�?B�~�K�%T��m��'B�3:u6ߕ�]R��B,�>�4�5�x�� ���=��k(qnBc��T�~��Jy�о=ANwF�W��~��'X��Û�>����~��<�V1�\Ɯ���u�OR1���bΙi�5g���o��1<��{b�aצ�y���KB���e�6Nz��_��t��T��v*v���p��.�+��:UJ�w�B�h2Z�(�^�uX�Y,���*~t(�ؗ� "g%�}����[~Jjz�S�G�����n\7p?�=�k%i�G�@�_ͫ����=ѝ�(����gY�,�:z|����D��ޑj����̿���^ך�8�����]���,�ܥ��p�����ГҐ���v��A��ke�\�NP/^r��I�Ċ���o�g�dk��§*
	W���z�8��.M��B2�m҈�S���	�G�`��?���9��l�>˷3=�M�`��å�0sr�o��7�0y�Q�煣@�q�ܟ����#�f*{���P4L�#^*Ëz���(����d�����=F'j�> �2
��7XBol�kZޚ8J�q鶥}̸�$پI�#�[�H�'�|����E����MؔJu�֞�$ �������e��<����ĩ* ��������͆I>�%���S|����v��4Ջ �������A�r�h0z� �o�������y��c?���V��r�[�*��M`�w ��q�+IA|%x��>g���ŷԇ��C|B�����΃���.�z����F6`f�U�zG�-�2�z�A`n�Ջh��=�а�F��w/r��n9�v������X��"%���&���}`�����:�q7Ύ�%̮Bb�%gv�lRX3-�����n/LylXl<�����-�R>���c�?�Q|����	�d��q�弽 �g[u?�Ğ̇�z��賐#��4�,��.�%ebjs��R>S ҷM�M�gLI	���$��۟hJ��͝�V�<�x�%0c}�����{�2��֧���u( �K4�A���%8IU'�� =��w�����5�xø0��������[�����Q�K:�����l �7�O��?t(�Ӓ�+�7�R~���G�|ۋ%y�ŝh ��aA�>�ߕż[c0I�att�%+�8x>R��l'��.�5��Z��;oJ:�9��W�6Wݼ��@�5^[�1k��V�zV\����� �	���w ;���+f=j��j�����O���T7>�5��Fȼy��[�͹KQ�|��<��'����;쀧2�}��'P�:|*b�g5�K���a.b�80�	�5��=yWީ���� |�POV5H�<��}�~>�Pb�q+�~m���d.N��`�}Yt�=)S��5��Z��ˠx;�h5n,1�,>�����S�W[��'#���i��eڊ%7ڛ��>O�k.��o���5����1�w�b�h�b�C�6b��$ـw.�IN�B��ϺR�����Po��ZB�����9�S�ѣ��y��K_�!�nHL#����������?T�F4��HR\>��>p��"1隣���M�*��I��[A�����X��24�@�{�P����l��F�\D��!�{I��7Ҝ�QԠU��1o[�,H�0��׼�n�7�jh��DV��ʌ����#�c̑�,FI��g��U=��cd�̙4�k�!]|'4ہpF��t�6��p���f�ەI��'�Ĭ;Vc��~��a5���dɽIf@���48��љ�C��Q��7���$��,F������{�]�b�E���mY0��q�u�I���Ω����ߓ��A�S���n�<�
��,6�G��Z{�7Y3Y\�}Mj:�����>L�r;�dWoՌ��֦߻����=j
�Ɣ�w��8�J���7�������/I�f1S-��ڛ�>��=xt ��CƸ��G�Oy33\@{ݾ�7�0%;�j��K���
\����"I�Έ��6��X��\7�ܜ�>�{��	���X��Pc1Ap�O;�k�rsw�a~�:k�K0����7�61R�ú�&br��<X��!���N��NE�������9A�g�t��s0�Y����n&��SӠo�|R�������#���4N���iı���������(���ے�\d���d,Q~�h�髢��]=�`�k���Pw`0����M'���^�	rYt�z�-�6{� �=�LH�J~�K��Йe)�(�R^�
���Yr�+���)?vd��	a�/��ic�;�-4lɐ_j��.����F�M� ��r& ��*�^*�|{���ߋ?&~�G���,�wa�jc|$�]o�Fۯ����GB����;e7�[{HM�Vi�$Ͳ�w��x*��1�|Wqb-ifh�A���=S>��U$u.��X"�	×7�ÿ&*Vi�&w����m=P�j��Ӗ����?=����)S�o=c���^H�{��Kr˻!
Y+��.��H2(V#�?^��0?2C�Y��T��]�kiS���r�#�aE��,U�n����x��t`��=��bpt���>����n3�ib�7b�����, �"O���u�%�#~��7�իF�|��%MʷC��BK=E����ӋN��`�M�*W�Cp|�f���W� Ub�u$�.�7�6-��oګv��x��˒�����o��\�>��-z�jN��y��#��Tt�|�x^)�'��A G�E�p�R����ԅ�O-+�����2[�ȗ0#��{rx0���4i�s|ճA�FŰh�9㺏�'mL�(/�KF�� �oHh5��M�R�T�|!Լ����G� �;��ڲ$F�L3�F��?Rx����8b����K�!�p/��,e����2�<�˗�e�bq48L��G�|��ζ�'��|8�qy�?N���A��՛�5>�N���^# ���[f�4��Zi����A����2�hX	��57�~"U�a�(�yy'�Ѭ]bXO|�L��K��>K���oÛE�>o)|%�>C 7g���>�#�UDM.�Bf2wV��\��C�� C��v�3Z�]��W�����K-y�p#B���8�=cq���' !~�_Kګ���IAM�e��Zv�§���}[�� E\���ʽ��z��:qZ�u�����{�B�*�m�@�|GSj&�oC=�I�9�����&u9�ș�@��gw�N�x��O���L^�@�o
h��j�� ��ڢn^�T�ìՈt$��B��'B_�Qy�QB���_��r,݇�=�"�]��k�-�:�fA0�63�3���ȄI��oe��b�m������AΊ�Lӗf���0M� ��P
�<Ț��x}�X��_�ꅔ_���)~e]]��#.[������W��s���x�Xƿ�
��� �b�Po�&���ڭ�ڬ/�vƐ�3��kN���5f�e?�<���}��n��5P��U�-Jk/�a=��Ub&-OJ.�Ҵ7�֋0���޻�p�?m8K����d�1�I��n=�G-����$� ���L�JH���@�H�7A�vb��+�E�����o����^���×��I=���es.�v`�x/������"w%�d�jV����Hv$�~��А�߁ �?Ѵ�t�\ɯ�#Mꭿ8G�	^�)��-�*S!�rQj.�v~�3��S����,��� ����M,V������I����3�[�y���c�r��nW�[>x'
����ۛ�M� �}�}�kW��d'!�*&�}l�FR0�f�6���F|�Ϋ'��/�Ďo�% eY�����}�^�ei߇��7��;ݞ��u�$B`����[�Y����Ʌ�5 %Ӈ�U��@���2.9�O�Dh��u@����2z���2E���Ӥ��$|`\u!��;$����7���$A#h�*�%i��Tݴ�W�(�\k�ўƝ?Zî��&��c��t��]���UËu�N��������X���M:�j�{A��:�"��Psd��V�H�L
��Rg�������v���7NQ�y{K�x���3��J��S,Z�ˉ^C3?g'�%�Ua)�%���v�C�q�iO)���zҰ����S��P���k���_Nc�7����K�{� TrtO��LK޺CN'�#'_ �u-�<�u��'����]�D�Z;&k"��4��l�h������7(c;ճ�M��z��1�m�@h��^�IG0����4xxf�r�M$��|H8yy6_LG�s�.�8h�~�O�1i�(D�ni����� ������F
-]FN�c��SG��h~�/�c<�Y���#5\+�e��B���t[�~}B܆e�+�bV2}��@�M4RW����!�"��_ ���6�N��&Vk���۶!�9�ǿ�D���8���$m��tZr���`6tE�C��K��Ho�#�.��w�q��db=?�Q������?�ّ#��dh�����l�Й��W	�e�1�7�6M���O�I��k1�>;�5��΂Q���cW�5��Q��W&,>����j�{� G�#����Map�{��F#yd�o�쾱�UK�����ֺ�>nKRꑉ�]�Џ��}� ���辶�<s��͊҉䝙v�g={k��xhJ��X0�l	d�P3IZ	�����q�O��G�|*��SQ�v>��%�㫄{F����n��GЬND�on�zl�J�5՟@�;*�CΈ�Kk�]�~V��
G1բ��8ZA�JZh�;ߺ�,���݉�uWL��m���-S)��:�D�?�/� ���C���gB 5"Γ��&���}��O2 �3�K�{����P.��,߽$fua������	?j��
�/�L���HG)��Fm~��Ga�����'oV��zqu��I������?�{iQ��9$�hQ�_P]jC9%�_l�LA�~Ŋ�x}^�e����]~> ��-s�_���n�o�ۈs��>Ru��C��J�d�}=���	c��`�������"�?{Az����Ӆbi�օ�dI<���<l!U�@']�>�z���������P����ĩE�
m�6��D�g�Q��_���ғ��/N��r�R�ȅ����7�w���v�%��{B7�� Dg	-J�?V�.�8K����viA���׋2�\�V��vm��նG� Xj�C�"�I��θ�pA�����w��&ߌ,7��Js�O�u���c�굷�Wo����}D��D,����h	M��U2��j5Ƣ�"�����&}o.	�v���߲O�"ϼGvd'dٚ������PϞ��\\T��q@i��N�P6Q�� �)(��)�	E_�q켘����L�J0X�<C�ke���'��w���ȫʤ���b�k����|3���|R���c�uԦl̳�@�,n���	�!�,n������s��8
8#�3��ľNҠ���&;���t�ķ�!K�z�*��E��ż�,ﭑ���$��Z����>Ûe�ZS�T�-Ø��1î�<A��|}d�����."��)�AK�z�a�}#�C��
 z@"
7��,U��:�q���I���2��:�ُDԉ�\���nRB9f����'�d�x��ʞo��q�e�O=�͕!\�@yK%B��+#g;���&M;O]S��	�a���z(w�`SvZl�La�O{����|~l���p��{��g�d^��)V���oR�����0�[}E��@1���&V)Q�ج�W*�㓷,����ϝ%z�Yc>�R�����Opڤ�S���[�Բ���n�y��sE������0�m#l�˖�\��f�>3�A^�ku�B`+"���{���ڛ�Y��D��])�wR]S���2����"�:�KpjE#J�0\P=[�B�1Ar��X���b�>T
 ���%���o�C�C�[C
��j7Ͼi�Z�Ӊ�	�<���F�a��w,_��ր'ف�A�����V��R�����x�V�9�s��AC-5%^O9`c�h�6���K�n��mxD��o>��G�c1�v	�iZ�~ҳ���I�C��V���!��V9��]�\"%���S�|������WK��5�#.S���Z�΍{��#�
�_�C���U��Ђ/��l9��9�1��4����Z[�w���ڽ�r�(,X��{�r�0|1bF�X��"ӥt�l�'m���\!�x�ߐ/Wʢ�2�&�_l�뒜e�-Y�,�C;�x �繇稍�d{T M�^"� ��_�D�/9����Zn���v�� =v�Btmْ���-�b7�O�I�zs)����I`8�4�sU���mLF�5��
og��ͺ�g~E���^8r���W�.;2����1���ߑ�
wt�Ặ�e��:��9q;(��i���U�������ͧ{��)���[��x��]?	~N|�+��C�S�=�Kкt^����������p9I�e����;-��
֓�� ��
9˃���$�l4��Tnġ�7���HsSAj�0G��"|7�|h��1z�6'LmT��o#{Hse2����*<�Fg0#4�Je���E���@�� �չ���w���8���ا\�d��m�bb�x��u�TW�<�5*Hڽ���
qȚ&���>�$��b__�Df&��N�"��:�~�q��iR���{J��FEh��Dx��Yi��95����Ovw)�թ���xX��8��9�;�D�gc���L�~:����fx�;�� Ϫ�����+?�@?j,�8����l<-�6��sg��9N���~�mw���+ s��q��``��Ajz7ûuՋ�q`A����*{+���˦�kO��$�fH�ݟQ���A�K�dF���@�\��S*��$*�li��R9V1��3����O��{psi&�ؔ6�n�-O��u +E �{~� �?D���7T�.vX���_�B�+B���f�ZfC؊�ؚ�	Ĉ̘wb�k{a����Z��;��Ur�,�-�\��f�TцRɦ�;��'s��ƹ�o'�ߓ��h�3,�/SW�܌3t�o
�Ye��%��1�k'��|�a�o`Ae��($��Nu��]�L�-i=��^�>�n���Ä�w���=Ƨ�gA�ʹu��߹���ݓ�В��&�_W�$�ވ�Q��US�W��=��|��MN1�Z\8�0ѷLH��7$>

I�1�	�8|�����n �YyKF͖ΙzkO���
o��H\ٽ� �Ex�����H�3ʦ�?]�.���>U�[�'y<N�	�Z�q/� ���Z�d8�����\�	�%�MJ�F�#��<M;�Jw�I���Ҟa�{+��@v�&P��.�e��d���e���Pq�W�y�Pwȫ ��ڱ��7g���Nf�{��(
���\��5�%D� �Cv#ۤ&r]��ʎL�M�J�P�n*�\��Ԍ���_S�_���JD/#i��n|�w��P�냗M�;����e,����GE���n%�8��(�nk��xy��K_.&Qd2���Ȉ!t�+4ҥ{��K�~���������ɏyѳ�ɬYz#�4t�����p�B�.r�~Lb���y�$������Bl��N.�
RGaG������~��� �C?�7���t�*Y!3(v|�A.�f�,�QKO��d�~�WÈ�b���5�[�{�}�5O�С�& ��%��/��ݽ��;���h���u���U�;	Ȭ�N�{�2bj� �J�	�iP��� "���b����;��P����J��@����/�*^�5�� =�"��t��/�/J�L������9]~�KIUQF@&������^���8�����-U�Z"��t|OU���5j3�Z��T�r�R��Lx�P,��J[nhͣ~S-erH���cX�6t�BO�,�(0��r9M�&�vKX��&������f�/ٛ,��OF��C��6�'դ��YY��Or7��#ʋF$F�w�X]�5HQA��Q � �>ײg�y�2�mS})?>�oo"$��*6����lD��'f�<�U$V��˗C&��>3K�}�$��a�2�T@M͎���S�~��C`��Qsch��N�CM�T�j��ؒ@�:(��7ryTq&�d4O��is����[�����rh:��$]r�:j�!��'hS���遙�b�4�դ�P3V8����Y�������h�ӌ�����@R������cX��@�O
�K����߂{�IG����ϼ��E�VV�7�3D=���ҍ���~5`��5F8�A��p[���9����1a�eF�>�����{��R��}�
"�x e�Ƅ���ie���r�,_��
=��C����9=�߸��˅A�Yqǈ�����$����F[����m2{���n�Jg�g�>#�}:��$�m;8�O��I$<��DM&`!�!�$G�,�X_ǆ{S���;f�L}�6��F�/.���DBTe9��4I�v��D"�=�6عK�ˮ����#R*}P�(���'U��<鳫�FiL:�֦�ܿ�S�	���3)b֔^�`cx{���Q^x0&��4%"�!���
� ��'$#���B�+�@=�9��r��w�U��6.҉�1�g��]�o}�����6����A�5&u�H��Z��h��w$%mg��UK	s�\�H9u�H�4��F���B��~Ⱦ�^q��n�:�s!�go�D���4� 	�of��K��dH�m,_�6��G.*����}Q3��Ŭt!�"���WL�]\���	Ɨ��p��I4˘������ڿ�/�������:�ze*�v�e�n����*U�C����`-s��G���?/��K�i~��\Lu
�_o?2�O;�ׄ� �YJ��	�;�ݽ�f���Ϛj�du��<Ma���I��X�w%�w���_�@m��ģA/�����N��r��G��!��?
�3+�pa����TӮ!�I�W���|��>�F%�6�Kg}��^��P�ӜU�02|ƙSѣ�P�)v���ȝ�tQ�_�A=��`�`C.��I+d�8��&����LiB�f��MW �,}&�V�㔝���"mr��҂�c���P���/0�� �֏��)�� �0x�$/�@ֲG�a�*_,Aa>��'�*�q���!��$�~�0�����0��b�l���QۀE�M�*�2��JJߜ�6C���h����%ŎƢ4r]�����N������
=f�hB���v�*7��
SJ'�C���3�@��!�d�����?)�s��KI#Ь�r�r{��#��a�w?:���5��f����|y�q��!�`��/��.��"=��&��m��V�0!�n/
���A�vG�^���$���ZҞ���6g)T�r��E`4�L6Pd�Oy\ lz������4�M�8k�˺�~�f{�㾝�b�b��݊�еHW$[6�e����%f�!�vB,_x��i�;t�r}�Z��IZE/�V�\�ȡ�u��VC���Pg(���J�9a���RY�-�w��=��7
�4��N���J�K��#��^AT����PE|LQ�:J��|�K\{f߁�ۛՒ�)�&Ba�ŦX�����cF?�(���HO;���\�9�D ��(�q����m�pO�P�<�Fo"��-��^�ͪO-T�a9���k��sL�[�����A4�_�a
�}�\��wd�B
3���ha70�BN�Ï	�罬���\k� �YQa�U2�<ä}�!q�^�v%����krCF+lc2�C�{U��?�ױ /�����0�����e�� �7D��F���у?D�g������K�� `�f�u�̯��/sV��'���<�f��Ou#�	�z�`��5���U���NK�hMU��4�!p�*�%+ѓ�q����z��^�w~eX�<��W���ϡG����c�FO�r۟fc��V �BqF�?/	2�a7��J���Ǿ6��q��҆dqf�Y��G��5KoR�o�1�{J ���gM�i�TG7�'T��W`��.���� A���c*g�V��l��y*BҠ+���D��u�A�v8Eh�2}&�[KDr�fc6�s6���E��r�yG��AuUAa���Y�W�fG������ ���u=~������ҷ� �A�.����1P*(��BNܵ9�|x�gб���'�t~U9U�UN[fӒ�Z	��S�]�.�1���Y��V���%Uw���p:���#��/[��ġbm<����U��qJ�{*T�@���3F�K�#�v�%��IG���?"om|$���Qqi��{Ԏ��=z�����"'���Ĕ�� _��Ya�ÁiX���!��F��׾�!�;���^�rRQBI=���dN:��R'�v�1<ޠNY�|�.Ug�G\��G��&>#������Z�-�I�?`o�,F��	�no·�����}��a<O%�m�R����إŦ]8>=E�n���e���<S��D�ջϞ��&#�9�D��m���@8{���k��d��T���H�8�1�_��B�e��L6`R��7Ux�Úd`�I�v�B�Ɋ7G��P�f�	�����Yź����nqy�#R�U�*8��C	�m�Ҫ~�������{� �G;��Ck�4^E�t�O�3������U�8�!'���]����ѐ���7z錛�<�{�����(��n��fR�?N��W.ޯ�<���	%"����ח�C'��;<�I�Y���'�y��3C����X�������9�}�h�r��ͮ�z�,�I�p	&*�Y�%�)Xv�2�5g)X,C�&b6�:��&�v��zr���ԶU��_�j]9���Ӝ�w�/�'2�ȿCD<��1�VD�D㔐�>$
��R�$|�!�v��4��xEr����z�����(�����儦�cF��;�w���[���;�Dj�;�����^A]�K�_����n�F�b�֧���|\�bV���(Mf�OF����i�ai;Y�S:!��t�OƱ �f��i�}#3��v^{3z,��x�9��4P�jux�<����6�U�t�4��*�oK��a��ɂ�l��� HK��;�q%�(B�f�;rד�\�u��Z�z���|�Y�勇4k�֓���ϗ1�W�J�">R��%Zш�}��/qV2ԡQ!ｫ(��w��QE+��w�
$p�����~���iXb'%�h�'?ɐeM,er��x!n�n���7�r��hv[ �f28�lE����zu�2*��l�ߐ���	;Kw��{G���5��b�Tj.�3K$����>eKL�r_.YN��Bb,VX��f���������#
�ZS��7����ضA��o�g6YR���YX���ޖ��P/�>�Lƿy�ȹY`���yMqO���H���ab5@�)���H��NY�)��Sz�T���VD�<q@?b�$5:C?2�6�U*���o�5"�)�Y��CLV妆s�6����d�T����<�Q?fK?�N�gU�K���HA��z��a�؋z�h�����ȴ㦩_��,�e���h�g�dF����č���0 -w�&���$G@�䝑�]g�\�W���Q�|��~����Aq�k\ѫZ�q�nn\�_�B/�4���Єe��>@�}pp��5�]���C&���(5OJ�:{����-�G1���]a&���a-|�9��L�D���pUuƣ:(�ԓ?k�i�V�OцѴhv!���d6�r�U��� �C�Q%����.�I�\JJuؘ�|�~*��"ݑc���:��'�])n8j�~7/B�
e�M�75yY�񽢀����쐼o5�� �$0 D-a�72059��B����Ԉ�$�z�X��A�	� ��{���z��Ru�@^�b][^�f��4���&�^���s��R.�8�����3�|g@e��N#���k�q�Rf���P�k{��Ws�N<y������O
��P�@S�&Y���c�S�ʙ�h�����r߭�c�`|�ޟ�_f�Ԣ�����u� H��k��Rv��Qe�h��p���
<%�X�^jP���y�� �h��ƃ0ėUgӕT�M�;5�[���>Xioծ-C��p��C���°����5�G *��h%ę�w,�>�بO�=A�޵)����~>Pu*N8D�����
�*�V�CCEƂ��';����7�s�զ���Z(^m�>��w�Ԕ���d��z�+�j���c)����7&��h䢀�̠����ףW9��G�\{.���c��~`ޑ^��3;.?��Z��Um�N����Ĳ��� �*P�G�y�Z��������G�����-�m:W�8N��fY2�lN���űW�K+!v��W(y���{�4.�:��;�_���4* OXü��� ���!���\�C���@ɦ�$6�L�%FUW�&�3g�-�dC������C�.�H�RP����"�洛� �R�~�{�-
{����}�ئ�y�S=�)L{�f9�*�B7h98��,$J��Ė�dW5J[:Y�>Ѓ��0��+��Z�Йj��?ZO��$"W�E�C�8w���}�{U��wL ��#�n۰;ڪ�y�T���UkL�rp,�o�����ԑZ v�2�5�����k+�l��'�[�1b����� Ʉ7��.9Q=������AM�;�g}�h���l.��V�����ULL�5�[��C��F����������MXso�S9�L���<�x_g��i��^Ю��h[�3���W|�;����#�}�1�%T��2��?R��n ��V}�ҫ�U��p�������o������º�RG�6�������*x˳�s�Ari���v���U(��<!3�S4C�������D:t?�M,lpuON��1�WA��{�`�=�?�p��F���F^����C��KWjQ[�a�P�Z�Q�c���m���O[7J$�?;�agr�BA��^b����
�|`B���Ga�A����C��gGk�zld��tp�<���u[�z��S�G����n7G���*mrpG�@m}�*? ��h{������
HI�<��G��ʆZ�p?03\�b��ԍ&�������݈\`k)�%a�*X��h�����4"��{S�;(
��є�x��[!�(�#�P��ǁU1�6-
L@��E�>��ŧ���}$[c�3����i�'�B�j�қ)��:�?���ö�^�)��./o�A�.f��4]�H�zl��t��c��Ŝ3~MAQԃ�����aS��cR���Goa��&|���F��3 �q�ꠚ��p�R�@DG��r�h��������M�.K�~"J\	�ϝC^��G�vB�J��ǐz�}F�m̑�E�O��U,��#�s,��C��
�w�f�<gn�J�����Y]�K*g�]��
�R�b \��`��1|1��{�~w��U[�Q�얍E,�Ly�`��XԴ�p�(��Ü��ȁ ��T�a���azYȻI��5>�~eI���ۍK*���PfM�d�g��q�����5�$_�"�} 3l���R��U��69PVOg�w�(Yl�-`聢�/�;�&G����/3
DH�!<ӽnc��":��7�dG�ž���ؕN��4b��^�SD`��SH�z��|�Ү�2�F����C�%��da����-��mx^��L��*��n�>	(��L�B<���{�熟{�I	�$Ԛn���%�f����A���.��68��&��_z*@
������ե��Y�Y���T��Ъ�!'IY��0G���ܽ*�y����/��=(�[G$����i[x�j@fY�,6ai?�"�P�q�mw\O��u�9�O����<׭7��*��W�Ň��OcrN&�}R
qV4��P�G��**-�%w�FW�Wi�ɪc�t�#�%��5ly����)u� �v��h��]]�ē��eô����U`��H��$-[4������@t����7�/���2���߯�t��e��Wř%���I��Z��Γ�xT��� �P-�ރ㱫{�8��'�5?::�� �} �A�p�	<4#�=�-Ϧ�+f;l���Rzڶ��0�Tv<Ua�Ci�@]?�!/^>�p��ޣ|</�X��܂��d"?��Ӡ��HY�s��c��������S�ZՈ��y7�����Oa�F4z�va����|�Ln�����O�b���Lڋk�n{�8�n,c&n��=����E�l����v@ǫ[�8�V�����Y�5�='���� }=�7��SX�Uw��8�Ms������v��z$b������8`#���C���9�LPF_�׆>��^��[mG0@����TalP��pb%%�00Y]FW~�g��2.nhː[���$���T���n�JlV��k��KP�_�9L�!��n�}�.Y!�O���t<��g�I���d䜅|l�DX�Ƥmj�?.�JD�T��D��L�L���D��������,����V����Z�x��c��'zm]�V�L�X�v(�g/��YU#%,����-�gQ����|kʹ;0�"��M�G{`�j���$�J#w~� J	eTv���z�گ���@�-N��~���a�9}��Or�~xi�z'{4��^��Xy_f9��2�i��2��S�7��!8���+\(0M���X�I���M�gg�,��?��qB��ON�j[99��.����읬J�e�њ�T�B[��-H�O�C�=q�cG���U�X��P]�g;��;�U�'%�� �@x�yG���բ��d]<iQθ��B�86�� �KA��c�Eɪ �["�mhB��Q��D7`��%�i�-� �Z�B�j�P� �%,I�öGi�����r/Hs���O6S����D<���ڷ��2J��v��+"��)�J�6��oح��Eb&��%�*��BK��������A��^�Q�s֍���-R���p/u���:b��(�a5C'i�BE�e�5G����},8�x��
���Mk
�`!ھ�\����jǶwwp �LL����
���\!ƴ�3�$ ���4��Z�t���&ǐ�
m͈e�m�`�{�W���(�D��������X�;���>}�N�@�C-�=�J������L����a�#3���g���/=�������,B�U)���x���W<�&��+�Z�"�4��Y�H\$,�(� ��aБ��ƴD^l�fuf�>N6�52!��z�S�#�%�k�cL�'���"��?��DճtU�vʴ��
[�?���� ��hb&��K��@
*u6���b`ts�93'9�t�G)�^[�����<G�E���m���q
�����l�Ӆ�Ž5j���
�~��|P�/������X=�4ޚ����U+�D�O��;	�ѧ���\xc&8�$ć8x����h��݈t��� ğK�-ճ��G��{����,���H�~�nƎ�3�$���� ��S���ϔT|)��X���#�a�h163���J�d�XE�҉��O��EX5�l���/n%����SA$L�sK�,&�YrqX+�5	��!���Q_���P��o�� �����������ס�TM�o�g�y��Ͻ�׮.�xR�^K��o`O�̓��H}%Q�('HI@�v3�����o0yN�&�!|`b�3Nx��ӯx���o��Ϸ~��ƺ��L�T�v�y Ojt��f������rmg��z�\��|��V����l�('�H+�K�{]?��g狠�&�(���#�����;l(poo〘]����"�+��	��U�ܴ��c��r�_R�J�h4�<�Z����Tp���P1Uu�������g7v�1�q����LE�pζNb�flC��*-�w�g��:�Qs
{{��T�<�|+����c�����]�m�{.co�.0�y�-�;��i�9����I�|٨��b�hL`z2���=���%�ax�0����]g!�˿&E�����n��V�&Ys#.�Q�	��G^x>�I��(�kZxH/2�ˍYD����	Utu�G��w"��R���AP�c�)�J4�z\j$
-�ns��*�]��bXܮ^[�:7*q���Q�E�[؂c�
�Hn"}�J����B�jPQ*bB�ı@�]`1c��̐�=P6/hb��~������a��[�o��� Lu[PZ3+��T�FDOdANh|�R���I�[(v�!���:�em5w��~��r.��P��N��Q��e�����>��ƈ�ڴ�mxu�$p�+��Z��ꭷ�ds�Rx�D��Pi�(X�|�SB�6��Geq�D���F#�����p�@uӻ��tz�֪�m��q�!�g"{�H ��[��������w�5'?NL\Qv�@�\�t�'���g=�[�G�����B��c&�v�,E_���P�/�5�6���g	�)�d���j���5r��_y�7��Y�銞T���.��G�P=��"yT�V��l�;G+A�П��n�����7��Y�3��3�,a�E���pQf�UB�*c��b0_�y]=Ѕ�8�=�)Xxq=��S��i��_7�	ʪ��_�rC���۰is�&����4|>n>��=e�ü��	�D��S`������/5?tTx]�h/����0�=�B���T	<�p���{���G1��iǋ�����a��pl�Q�z��F$Ũ1~n��Lp���']ǁm�Q9�RᤒǼm����,�	���W���|��n��g4<��{�ކ�0v��}��qh����<������v���B����T�[;�Y��ۧ�Z*@S�LH@e��{N~/�����/��n�M0���+[�j�ݤ�A=HlȚU�,�ٰm��L7@myy7���H.�T�0�"	��nï�P�C���_V�B5n7_99��4�{/�Z�T�����J�9�C�VN�2rٿ������J��W8�Jӎ%(	i��>���>��3>?8���Ç@�_�@I�6�ϹC
�<�__h�Ѵ�\.m�R�ٙ6��P�_�	�>��&H� $��P�fd�	�ۅ�ј�?rt�=Yk�ǻ��p�����Ӄ���M��Th�2^M��z�(&���x���D��F�� d�8J�ߓ`pb��9=]��<a��%��$$ճ��Hg�.t�Ǉ�'ضmO��q��B�n��\8S�=k�a��j�X4�[y̐@�A�A<VވÂ���;k �v ���̞�u;ہ�W�}����������1��$5A*j�L�V|��L6���s�!�D��?��4�M���f�%�!j�nS����WC�/R�H�I�2�,v�C: ���2��Ŝ��Ǒ\�l��� Dqc4�y�,���j�j�9��ȋM�Q�[3�c=#R��{d�ېG�\�)������ˏ��p�]�QK��u�{;3Ώۣ�����gSƩ����^�5v�n���sbx1���N|;o_���8z#���	�@P<lI�ٔޢ�
E�y�A^<CZ���~��<E��X��f����K<O�-���7�v�c��ؗ��dVF�9���Է�3�(�tb�:�FJ�7c�[�.���]��@�t;fjН�����b����]��&���tQ���'�xx-�T���' "�:����{���`ݗ^W���\2�j��� �؄���F���g�A+��w��G*)�}�sԉ~8�S�P��In�)���h$<|	�r5eM^���=�:Ci��T�u�r�O:��e�@��|U��9�m#��|AV���)FޥWIt�.dG��
p�	�ZOh���=bNk�Q3
����9}X7FTUtfg|�+�_��7蔣�60LM��4d������f��<��/�c_����,�?O ��F�rȵ`�D����HM�`�7II���b����UT2��գx�J[7�,��:�V����ذ���(��3g�}Y��LT�}��/�\� �D���왉��~�=������4N-��l���u�'��N�B*O�z�;m
D5���-�bʄO���X�l��iS���Ad	H�����N�.��^Wk�Bٯ�X����.�y�ȧVNL��S�k>aW>d�S%�=�Զ���&����ۀ{]M���F��90A��@�E��W�?o�5SX"�w��%j8��k�t��X���T��%�N��|yo. �p��r���m�5���w16Ѣ�`�}� ���v��e�h���ku��Nl��~�X&�s�6�U?��sO���xs�"g���:��9m�N[���B��!��w�/ә*ъ �)�D�V�;)�i����~�� `����H���0�崩�Y�%�?�㱘�J��yO)�$����xD��>�9�0��c�\���|��E1��ZL3�\�,Dj1�9�*����=50&DF��!�=Ƈ���8|��O�)r|q�T�p�0��;��~R�s"��d�\t�,���*�1�������F���?�]����T]kP_^�A�$O9F�;l�	ᐽ�����>Ϡ��d~d�)|>LkD�n����s���� �m����{��av��,�T�$K|��gV��Y���-���X�_�M���Z�����S�����r�t� "ﻍ�����O6e܏�Ҍgw묐��t�YY.�] -9�����Gd�N��ݽ5g���=UIM��S�������^wTFt��BU�<�U�TB�k&x�^�fN8�Wx�*z�>l����c�b Gy�d��^�8������y,��]�eЊ�^e�&�*4~q�[����R�>8Xf���ɇ�����$
��W�S�#�x�;��!�ÓOgN!Z�l�!)�k�g��J9��&7#DS��7^�(�h����V�1i� <rX�|��e���4't�v�� S���w��ѹJ��ౌ�Kφ	�˩6�� ����5K�5c��f�?�6�0"�4P�<�y����ʞk�U��,FwȕҴ� i���$�����]��Dk8�%��1��\��F�*%Ȉ&m�X�8�&T�������6�J�l6͟}R�M�-N�j���S�H��H�x8�U` l��i�r�u��&EbɓQ��3a�z0a��_��`^��gt�ڳ��6���2־_��Kj���#]m���?���{To���t
�,�YM��T��y�u�!�LB�6��&Tͥ�nA.[ɓ���2��~T'�!3W�|�P��U����?3����r����pxy4����f��^J�
Q�o�S�c��d@ߋR\��3��\�~r���%w㍎�`;�k��c!g�e��{J!FsN�b6�N8�c�:�f
���f��Q�)�X�\��آC�خ���s�a"P$˒���jx�Z�q˿ኙ�4�m��2�&�-�ϐ�����rASc���x5b3�f�LaA��R�ٖ�nV�����H7� z� m���zp�e���!rG�o�	Aץ�1�IJ�� ��W2+��C�1�2{�aJY����r'ӛ�}O�"�`���J�Fʊ����W��s�@ukYS�C�x(�6�jqB[%xXq�6�t��O��r]�q\��}��H�!Uw]��ڣ��Ѫ�u6�@�����E�d����-��	��Tޭ�gc)#��VNT� ��z�N[�C���\���l�+?�*�j�g�ZS�F����(����V%��\\Jp��� �u����� �H���2@��v_����7� 4�"y�]�v��D�[]�q�e<Ȏ�1T��/8��W��9�P��\r�Q\�>3 �M�C멼���rǥ��ȕ�X�S޻������-nOH���Q���:2d�W��Y�v�n�7���h�V7Ԑq]S$)���z��I��p�^��ԅa�$ۮ Dz
�n����w��U;E�t�
,{A��b���H��&�%�y��rcEݔ�'W#��X��f��y-���8�_������s��:�X��b���-���_9g;y���h���tB,�_p���r�<��}T(��qG��aF�
�+X!*�gi��H���}�TP��1}nq��Tv{\Rwr>#���:p���`W{�E���t�<�F�1�h,��ߍ�5���\Nr���#&�*t�~���sR0��'j��<����w�ŉ�'�R9�>�`�f��2&�$��N{k��\�u���>Y�E9"A���nf�;M{�e�%2�G+ �ó ��R2:������7�iiZm%�F��HQ�AS
����z�}ZY�����37J�B������b�?N q/�
OI�Չ�4 X_rY�9��\o��1Hb����
���L�FT�ԂCO���P����!�cC<�/H�wrM�1�m�TvSrL���GNv(��+��P��0��O���R=U���=!�>���S��.1>$DFQ�-�"�y1��5�:�'P�Ju��
\
��}ݷp�#��س���
��e�(0':F�6T���e���{	�r��z�g.����V�@�t2�� vu�ʒ��t�b��X�-����h�au0�I�0#-���َ���]?&Eb����W�ag<�ĕ��T�e��=�o�7ݰ��*� ��s<A�-���{<���,m�A��X�ˁ(��xķ�b�LtX=q���\Ə
?}�Z�D�ɭe�MǏ�����Х�v��\ǔ�k}��	>���������[�hyVX'9���3%2�[r"a�:���DY@l��s����o�I�g�l%n	Ga�g^�i%by�h��+�v�+�=_�ԍ�e3�^\1�]� Xq���e�N$�Ͼ���M��^�h���&8� 6��[�� 0���VT߄�� �5���e��̈́��H�z�8� *�3��P���x��K�~�M��&�7��6$�Ҿ%���o���0�Jbt7�^;�w�����{��[��HYo`t�9ѝ��.x�����u���C0+
$Lp~K���sR �Ye;��K����������+���݅C�ғӑ�Ή��5h�tO��R���t��O@:d�L��V\��Ÿ_���1ܗ7�� �^q��x� ��ʧf�nV Qz��8��{�o���uL�|��]�u�-q�#�ZNiGVL�9n�U4�D������b��Y���b���K��c�~Dz����s0G���{O(��dZK����׻��q?+ֲ���g5~��M+될~e�?�eC�/��[�C��~oj�'n�ĀL慅�� ad3�,Z���d��[Xr�h�K-��TS)��>ȳz�no5~ڄ�. l���p�̴r���q1D~��S��*��|�jO�1�g"zqe�K c��P����ޭM�S�v�M�;���Q��Q�� ;�Oa�n���絺��BLo�9=;�ViI�z��N�]s�B����;˸�l=>��B�}��XBp�x�N�:����.�Ow��p��i�;�E���}-�o$Mc��x�#wݔh�57�gK-q�żՃ���ŤN7Z���2�!�!}�R�!�aF���g�)�*��+/U��^f�p����!2�,.��{�}#�b�d6|)#��VKwfU�IWF_H��4�(�\\h( |R�j���4�|t�)�����h��&����u�D�8�"�.�9�Cw�ݣ�fl��M��J�]}
v�7�r5U�RcJ����G~o��m�o������!��@H�W*����7V���5�O�4-��}�:�'�`�\�4T���)�
�>?�$mx�2{�̮�<EK��m�]���q�% ��4���a�e�K�o-�����Lk;)c
A����>���a���T���}UP�x)��!~&�?B��
�x���#Pp�m�W�*#my��G�,N���L��7Z����E����ڝH_���UM-�$��<K\\*�y/���l���Y{��]ɜ!���t��H��+���;?)Ս.nĂ��P9g ׼X��$�O�l0W�(a��L�$��7���+��ϻ��f�
�p����r	^�M�C�G��\k�f�?pD)�5���L�������\����Gyh���ʊ�j�q�-ks@�9v�H�:[�6EBR[h�7-=�f�hu��lԇtpR���	�����m�z�P��lc���^���5�!�[�Ϙ��u�VQ͠w�w|�Y]�;��6������HkG��A;N#>��d����M�7�����?L�vq��9"Xt?`VY�K^u�b��?��ecT�Cx�VH:=��P�y� Ͳqfu�ܴZ�ֹ=
��p0f;!�7�77�Jn���m����V�_�W��&��n�Z���@��g�ca!�#L�X�;�P���2�_l� �S�e�V��F�V ��Մj��wyU��CA�����$���J��d�D�u��`��vDZ@��d�[9���L2;� ���X�h��2�"�f�rz~[)j����12��Lxr;��9��#�5P���|s3h� �'�O�x�����uY���������S@&�]��aⰦ2{&`�|ܨ*,GQ�,�7���(I�|�/
nhQ6sJD�^�_}�V�3$7�Q�To$lr�y%��pA��M#�1� ��o��h��L��\{#�����8bm0�y뿒� �7�\�AX�$ ZX/&�����f�幙���G��1b1>u�Z�ZX��)F�	;���>�����_Å����S{v�h{zX6������M�G�2õ8�E7�=U��p�|[�߈"��n�� 0hu��a��o��5+(S!��s�q���7X�7��"���OxI&xg[��Wk��E|]ㄩ�)�ߩ�Mz���X51=J!k*gZw}�&�N�J�q�v��t��z�{�GE�з�^kW��V���5����ݜ�|�ԝ]�]^�� W�f����oH�t�d�~��ZK����o��I�TO|ٚ��0�&�����(	﹫�`{k�P�]^��c����G-Ws	�|~���{��5|�i�ӓ���	jO�������U�d�)����0i�F�G{��m'"���k���V� ����r�j�|ඈ������QL_W\���W�õr�4�p��S��_x�6�y�|,���C���	�N�-�ܨ7��Zi�?�H��a�2�)�[��(kU��[c7� �#�<9����k ��~�ċ�J`s��$��e1�ĳ��LA�?k@�7ܼ0[�Vb�mt�`���U�ԧ	(�v���)������\q����u-]�6kN��N#�O~��W +k4Z2�N�i��\�O�Nc<h���A�Q��.��m�c��@�@�e4=U�x�@�S�hq ؠQP�(�q�����t��oo].��Ly=���NK�Ɯ*P؏���gi��=��0��:/Ĳz1����ms<��䠏Ĺ� :�Ԍ�=/AT9�[�]�e�9�n��b�7Ki�'��(5�(�`��#�+F���/g�Q�x~_E�O��<��fp�EZ��
x	S�O��G�4�'�^�w'-x,��s�����['S�č����'���N��B���&��������>j/�ݾ���������a���U~�ȑ���Fφ��Ƚ�h^h��Pf5�{b�S����t؝M$Ũ ���0#	r5b���E@=G�UU'̷��;��c8T_�8�H�"����ت0�~��=+ϾͮWHS��g�d���*�M/�H���աT6ήjJËibɫ�T��\/�X���(3��O��T�rŻT�zQ�=P���Q,]�eվ.����Yw���YB�*����.���o��3-��h�̧z,(y��8��G�B4��.TF ���1F���9�8'Mv���Bm��B8��o�H裈Ԫ�?X��ƩͳD��.yA��Ic!.�k��D�F@]נ��ˇ}J��O�����W�4?��	�Q�UY�Y��%�bՕ�e��ޡ)��&���:�����ɝi�Gg�sZX�CF�<)3٠�hV��q��2[�(�tF���J�B�6h�b��~�To7?^-o��^� 4�&�hQ�N+X��g�����j�V��.�w@v��dٵ�Ku���z�0Gխ���9_? �'��!6#���%b*C���"�%��B�h��0���c�/�+�C��-�m��5��4M��TEڸөc�p��x�{��K��������V�;f�	���i�E���fV�Bh��4��z�� *Y� �Q�ׄ���|?��h*��<d`R؅�2��N�Y�I��q-Ex��̬�Q0�s�Ѣ��M�����,(��}}}jG�~�D�y6D��V���<!�qyj9Tw譄�
�jK�;p0R
O�X7ۓ��!Ae�DDWm�j��l�wQ�C��o��%x�ү:m�t��_����CU+m� �3U杼jZ)�3�;y����t�%�@�H�,���?�����ǰ���6�2�E"��>Z��=�sفh��rc7���d�.KA�.,ėpl�I�~K_x�s&L�u'��qq�a���9�����)<S��NP�"���+��B)(�����В�I���UG�$���l7^��1��eMio]�r��͌>�m��[N�Z�f 3ئg5ִf(����>L�f��;V��.X=���-	b�9
��Z�m�QwZЮ���5���f��^u�~i�Q�0�� �ruⵚҚ���P�a҅��!G��/�߃�s �����"awm0
�ƞ*,���cٍ
��L�-� ����p%Ք�du���<�׀w��bq^�3XuO��ǖ{�k�(��J�֌�5����"t��V{<�ay�IF��I:��Աe�qj�Ν����˹D#�4n�Y�	gJ��77�<�ٿ�X:�u�j.؅�ւ����q���HyM���'�p$t��k/��4�/��*��X�#�l䳧*�I:Z�����Ø�����5\�3�S{M��}.�d�?;X!(���z��@(
�NyV|?E��#)�����>@�h(��+��*��$V}���ʐ9i�n�b�4N������1�P5�ak���lR+	/�'�>m�ͯ)_��2Jp;��4z��u*�������l58���(��=N&:�>��"r�FǼfa�C
]��u��k� ��bJŹ�Ն�ՆB�^o=���ٚ=��Kw�9�F��;U��~%
#Z�)��n��N5��ᓅ �J�0��L%<����w�ߞ�}l��G��=��_�Η`��7�ݫe���|a>�*��*\���$���}=�e���w��Q�����f��4;軇2�D�Ϩ ��+#L� ���$W��w�2�c��Ѕ�#8���.dF�5��a�Q��gu��<�)�h��mJ��`��oEE{��'6O��U�Z
[���c������CE���[�^X3�"�[�Y�8,��:�H5����,M���J�*y��H�߇h93&�m�{@@�|_C ��T��Y*��o��	�2�;��%~�$�PͯE��b�<�*]��U�b�=�H��:��|�B��6��Y��
3򆻲p.l�3�?Z��t��@��×�]њ"�Bᄌ����'ik�����CA���Z<����A��i�r��&vs�N�ѸQhQ�k;؅���<yL׶W���Ѡo�f�sD/�ڡ�.d㪅6�A�+���y�	���3�VI$��k����B	�HF�IΌ�d\���q�ym+T3P�7WmW��.��g������	`w��o9�v�)A�R�������!X�4ĸ�4�2��⧙30��Y2G�6��ycl���
�U����-52��g��5Kẍ́��YD�T���z�{z.3����<F���<���#kbU���ҩ�Ҹ�e3�H<E����,��y�}�0���l#ҡ�͛_4��iF�MH/�����H�wwaٹI�	�XWjL#�C*t}���pѮ�O�j�k:��8g]0d�1���%<Ѕ�,L�:#�����A ���֛6T��MM?H-���|��l �ղ��U$�V���L����	�VҞ}h2t&/[I/�^�<�!��EE
9L�_t�¸!<I�������g�%y0��G@s>���>.��-��6c�r��r��×q�6�ڈ���LY ;
b����ꐎ��.�#� ��ݳqqvc�*L��+O�ѐ��+(L�6[O�:L��1���2���O���H�Ij�k�,[�%�GMn�}�p�Hob�r��\� ��n�aW}ID �����Num���ӳ�E�/Lǳbv���	%��R�Q%�ųA��m�?N�D0[H��A�,�D<���ɜP���^�m�"�`�o���Z*"��~5��cN��l��|���^�O<�5�c�~�$�"f����\�_Ǐ�������jD�_ӡ1����h7���GC�hᓴ22X`jB��-h��su�ue�tF�D��!��kV�k�xȭ?]g����E�q������#��1��M'����=��[�]�����؊$��K'X��z�r;�DN(9��gY�l�Q�Q��F��Ј1j��=D��0X��ɨi�ڼ�|*�$;y5�{Ů����+8��_k+��߲�ij����ي��c��L��m��ь\������>
"�>��l��؎dj�.�xD:	���Z
����<�:y01�7���w�+��	3��3�� `�`h�E�g{�7/�>�1`_���-i���cD��ϗs��w��S~�mO0wZ��ai���vϹ���8�B��8����,k +�(��^�2ofѤɲ(�x!Zi�-�����C�`VVA��r��zI�ڱ�4�1]h��;��r����m6SI����?��W��Y�N���渡*nKs0����6��e<sM곇�&���-�}���I��b����4��v�6��DX��|�'�Vǡ�oQ^�+��㣅�� ��%�(���<�D�	�ӧT�S��\�F�SH8Kw<Gk�I>���Cu$ɱ��;6K
U���
E�;�QԫI��2;���0��_����XJ���x�yw,�\\J��f�.f&2}�����qՒ�X/D�N��e�Gm��XL~�S}+j4N��J�t�i+��˼v��w��R�%��0Z�S.�����
�����ưN��n;�z���78��8:�/��5}�������bg�+�R��j7�(���G���Z�_L*�F�[��H����ip��������5 Zz�k����% ��������m�P��Q�Э�z~��y�?Z����ҵ��T$��o�[?B)Lo׺�3�=Y�҆���qws/�鈿�!�����@V�͑���U4-�ֲ��Q���������/	�2��J֩��8��Ƿ?3���γ�T��W߳�8cN����O1&vR>��z~�����l�@h1�ع�J�Z�(��M�+�я]�c'�&r�zc�~,鈸@����2��n�׭��eg�W��&G+��Rb�FT�������m��,��q��^ˏ�B��A[
�:�`����G*��@�g8��pmV�S,n�ֻr߭��S��߳Ųk(%J;"��q��N����	���%�h�X����]�h#��;.�K؅r�m��|���,`���`P�G�zW�ծ�D�_M->v��]���hфi���q����*�P�깷�z1�M+�["�
ĝos�t��{,�j#V�g�Y��c���W������Y��m�A%�n���A�
����jC\"�� pD�sAc�q��xK�r3��z֙�I��^<8^�^�����BH��F�����P!�jX�.��2���b���C���+:~I���s2}��LX���6���&����(�4h޻�Ҵ���Z�iNoކ~���������E�1yLքE�5�� �=�Ķ�2Dg�t��|��=�ѭ�s�/�GGTu�Lu
J
;=��/��`vQf�~������\��]x�<ҕ�'"+&q R����7��v��yu�F?�GD���\'�mFL7LC�<���Y�T����>޾c
�}� Mm�(�'GDT�߶��;�͜Jsaq.�-s�ͳ��ZW:�������?{��Rn��m��?W�:�^���+��X��F��Z�?�z������$�	�tSY��AR�s�߇��5�=xn�����T��y��3 L�a����0�o��	x 1I�B�A��g�����b�QC��n���~v�}�]���y�;`�F)�0�}�t愞�,hޚb�~A���)
��1!x17|u�_s���df<
��uۗ���tzN�M��_�{7!��Bnq��F?��	����霁���ԪQ i�"/��S�����f����!�jS;�*V�����ü�#��x��B�;��7u:ѵ�c�t�x�H(3����>5�y�-P�:f�A���/"(�<>�Pb��$�U.��o��j��`�73
5��ކ���8�P�-���L��
IL�6+���Eg݉�Q������~��G�����̛C��&?� ��0�!B��:�A��8"�S��>&�Sj����&)��/l�L��g�F|���-0�*+=������`�G�(Z�hY9��������"1$lD��S�k������7ܼl�(t���Mi��
Mc�[Qx�;/�����Z�%=���Y��f]�hN�Hv��i�̨�x3���_�G�`9�ҡ��E��^|G�`g"���`v<s7ߨ���r^����/�)���O��#�V)0`.�;�*��zm|����zU7 �ؙ�5,8��"ԟ��c�ы��!b�h`��NȤh��*
7�yt��%�����NG����0���x���r�!����ԣ^y-�����j�T�1����
��y�&����� )�L�K�����ٜs����xk�Kj���XX$�3==u~"[̫o��@=d�8�[Z^�t7s��!}h����&M��lLV�qp�KB���"�����U�����P+/�AX#`8D����o�od��~�	��5���ex��k�|����„�[]�t/ng�z���+U="��l=�����+>�\�:CA�`�0e�*��n��qC��^Λ�D����/q��;H<��-�Y/��y�����
��I�@���R*lw�lY[ڌ�O�7n��dC� \�]�����T�`]��]n�lIp��qwĞ��
�aM��Ń_��;�<�t-d�U��O�Z!;�37�A+ QJҩ�vr�%=9/������K-T����1���'3�����H��rߐQ�D�P?t���l�~0!%���+f��YCj@�U�ցE��С���WP�*٢?�Y�Q�}@^���M��:Q�߿Ѧ�^� $
�7`2rM�=���;��'i�2��H��v&R�~z|[k0+������fY�>�����ME"����L�)�����L�Wxo������$~���O'�|�7���}Զ�#G�?|�����y�0X���z�By�,9�1"�����89���\��"�|�����	{x@ܢUg}�9ڭjD��P����Y��X�� l�H�+��Z
�D%[J|�Ϧ�\��fV��c*�(�ؙ�)C���բ:��y::�&�~!���#�tv J����pƅ!j�}�Xe�g"�9]V\�����/~��8��b?4��֢�vN$��o�8%(±VR�/7�S�u�6�ɘ���ae�i7�?w�Rna����&:/;�)9�S�)��n�����-�߽S�w���>���J4�'C�����Z-!�iQ����H��J��I!{t����S�T~Xi���
����'�_�d������p�R6dA*���z�׌{��uL\9[��Աh��g�u�;a�}�o�um�rǛMV˭TѠ��y����M�V� 8����AN#�|gli��������B�#J��Ek{5J��!/��y�$�{�o�q�B��Cn,w�?+ه���~�-�<�OI�5@~`���}j#��{����ڥ�9|�I�⟹��L�A�'�ֲ�]�5�l�����(e��9��.1:j��y��w��� �/� �l��e��okn�M��ҵ�e�
�g��e�-e �%�~��#�y+C�)�2��d�[�:�����\.q�e�D��W����w�J�7N���GL�sK����	�'#�]���dq7O��c������}��yytVl����֨�^V�e{����ޢ�w=����~�zg.��	Zs=�vvA�+��(k�;�C��4��IK�ZϮ�\����3?�fi)sfM�"�^�t��n���V��K n���Hӿ���X.H�`�rH��P���C�\")ny�Z�c���✯�Q��\�������V�Ϡq���Σ��;�X�Ǿr2Vq���a\��ӂ2��s�럋|Ɵhya�T�!${\
4^��/�L��
��T�w���y���k�����p]Sw�k��#�z�`y�x�Xi��������c箣ǜ혌��2��9
�@D��?��|;��n�c�>wXӯ�qf�����'��R�4�s1?)�40(�!�8�0�Wf���L�}j�2�Uڹ?mP�G�E�-,��^D�.�kߏ ��(�/�9l�x��W��3���9�����]�̶P0��w4C5�
����n<t��$��e��.qᗓ��E�F
3T��x3󴃼U%H���}Z�2�')��-:]��<�������.�f��#K���C��n�꒫[x1���n�#���۟�"�3�	�J��=���yagS��Z吉�Id�k��>��~$�ߘ*e�i���QL����&�F4��g��r�66���@}3Q{F��_[�@6�R��T"�z��±�L��q���v!��TXS���XnqWbsF	t��e���E�I���[���ن5oZ&����}\<J�J$>��N
��U�&Rp���c�l�)=���OgͶ�����A�a�%�Ǘ�?��2N�L��;e*@���$�(�B�vΌ�9�c0������� ��W���s���,]�[���@C&s۸[��j��h����F�HSeA�@�9$I��ۧ�{f�|��t6+k(]��na���d�5�fEM�k�g��z�V�C�u��p���:c �:�����E��B���a�w�g	�F֦ˤAw�sM��Pp��)�H������,}�K�%(reFȬX��w�	���'����H
��]�u��Z�׬򗂴z8��VN����lHI3gt�n��7�x���~RtTy��V�>�vu�����2��E
�~cU�3��n�0����ȻJ�-��C�a�����q������Q����Q`v�bQ�10�1x�F;;?Bj1��� ŕ_3vw�����8u�wt)�~@k��T4���^s�p���т(�!'���eDy����cQ#�7�]�����Qw�R�u�<��~F�8W����9+>M�b�)��&��죵��J���N��.�Ж�_��^|�/QS��7#Ic�,�|q��GC��8*��:j+�8�JC; T�b����
f9����ے53^�y����$���CJ1fR�/kb��[�b�����H	��Qu�V'��0����4}fʫ�71�ܞ �]*t�ኛ �5��I@�H�.i�oh7�z�P��Js��eE22ԇڪlf@��yԷg���iU���o�
DG$�찞�^�gr��	5 �,=�YX�RP?R���6�xȐ�H4ѐ��ҹy�@�(ug��G&��Ϧx+�V�t�a3'��ۼŢ�Ï��+VJ�C.�o�Ka�$:$T\oKE��iQz���b�F��Q.�wi��S/�j�4�����.o5WR���3O�9�#f��ܜ���<T� �]�"�Cf�L�K!oN�����k�X2`I�{e)��a�G����/ S]�6u����
*�c�5Wj��5՜�"�E1vl%��i�]{2����;x�s����֖�Y>�pkø̵FU\��u�eW�T(�ţ�;�ˬ4��M=�J���HLN�;|-k<ݷ>�~�kLw6��%�vH5�v� ��\�i����<�/����c����ar�O�~��&-�z�8>�-�ɴ�b߷�~N�P�x,��ƿ
̣B��,�����=���ڍ�~�<�nr���r��� ~�#��C���W�~���j�. ��B�5A���/�+��s�����㯹I��3t��)�rh���/�b�9��Ak�gH�@�����5�Y(T�6���\�����:Fc/�KnWd�x���(yI�{H���!��%y#�`�,�k-��X�#��y�l����%||�8�P p<����Q�aj'��֓�J\��Q.[��K.|6�-ⷮ�(]!]���c��1`�
��w*�50o��qs�JPr�E��/��aL�v���9M�
��|�$��Ø@��&3�$�e#�]MU���>���)����ŦZUJ) �6�Ҏ�6��e%7�M�*���J�7���V=УqC�KvZ��Ȃ�`|C\��Wt��>��<6����L�`����s�2!%��G[�����y��1"���L!!�B=i�Ϭ��/ОW�:xM�t$V���2T~�3�OJ�����S��K�	(�`���yv�q���)	�-��#D����y�q�"Ȟ׌����{�����Q81z!��f�F5ja�yB@�Qax/��fV o�4V�Y�9�e��l��y��HtM�U�k�z��N�@�	��8mKN���rh@�k��CO����/,�OPzi��2]�i�,c�	�_Q������r�ҥQ�2�����8_�o�W���l>���}�: �]M����i��$�lS����m696*�.֩BP����7}f�0|L݆�^�֓s�tzM���B!�f�t�(0���3�_���+b�����+.��IG}� �mv/d���A�dI�3z���B�ޒr%TC=է����0 Z��/���՚k7j��tWv�O�q>���;ay��[��W�w�B�Ӟ�Im�j!�س/
@�c|E��|�R"��1�+�N���:%N�5o�-���1(���9�c-��<f��K	���.�������Q�2L�#L�����h5�4kE�j��^�,���b�H��k�nX�*��0T���2�a:f������$&����{"!�.|��my���D�$�T�� ���5��ĺ2���SDvp2[7����<�}����!l��f��C��%��}w�K94{��;U��O;X��y���w�`��;:� �i߶�0�{�H�RO�]Q��@�솷ؾc����B}����S��Ux��s��+�qm���$��v�i6���0��XI��Z���9�g��I=[I{�k�L'?���B���/T�$]g5�7��'}���]��H=��s��J��KӨ��oi�IJKrE���o\N)�*��G(�F���r�����w�����h�o~�,���#L�	�B2�7H�E+��"���z���t1����J��s��)@s��C�ʣ�b]���e��:�\��l�������ٜ��pT���JCR��/��ө��TK5V����s�ͧZ}�C�y�.������b�����y��f�����u���=Ϸ�_[ͩ�k2p���uB��5e��� {�D#����bx���"`���E0k���}��+`9����U�Bv?�7�:�О���S�<D
�'�W5g���E��|/��C����m%o��ZyC�󶄭o�U���RD��'غ�%�F��c�N�kg�U��>��&�7�N��@B�Ә:0T��x�^���W��oI�9�Ȃ:VU+/G������^��#߇�n\/�[���%���c��I��I�����p�㖝FkCkS^P���e|�SY����.����kr�l�7kU���k�^��<�	�?m�u�3AT�'��A�S d�H8䂰�+�J]�R�����K��!)�|��|�g�u�J�Ag9NL}�m��q��\��#~���
Q��G�-o���Φ璊t_�@6'����w�R�&aw%-6�w-��_�Jjs���>�)k$�p��D_D03w�Tμ'� NSׄ�z(�����������"������Q��L�aF�r�L��e,����F
E�=�bh�UJ�S�rmٲ^{���65�:�W5���3��r����Q�C����n�Q�E5��b��t��FÍ���5�������\�}/��Wg�&��>H���1�����V]�%O����Gj��T&�"�[E�ً#A�0���LMݡ��h ��B$*q��tc���a��;\jR� Sy3���5����_�=]�Dc|�Xw�J���yl�]�$_Uw2g?A�՝�u9�!"���ٳ�{��@�����x>6H|�_��lδo�<����I� 2ؘ#,7��Wc[0^�(�����b/MM��p0�����9/�6�9c�+FP��� ����х�I��T�)����xS�Ŕ��/���=_?S�(���u+qy��_����!�Pqz�3�/�ad�2����)��7��b
3�ڌ�f9շB�H���E�@ ��)�cdVR8<�6�}�x����ڰ�H�-�'��|dDO�ߕ/ʛ���x���������U�(�\�H_��|��d@����9�e��!�3�����O�E +$ç^[��r��u���ב���۸�J�R�@ 9S����
)Wn�r�����k*'���s�!uQr��Awers�eRU_ƃ����,�sx$�-��-ڕl%#���#rt/�����(EO�8�S��/�~�����;� [kPN�I�۰x���=cY`nr���J��ur5c��;1�.��*Q0����OO����)��u�О7�K��A�=乯�����:J �Nh��Y�̰Ǹ�s�(h�2�����[iX���	Pv�W��G��[��4/~��g�Z ,�8��|����T�]�KUY�(*�d�q-E%��"��l5D�w��A�.t�t��D���0�_�'�hpz�i�o���2�������L]	#�����)�ZZ�kx�)����}�n�Y��4Z���<&�2��)����E֮�x�PN/��������"��6*���J�R7��M�t�;1�ꌽD�q,]`�G�
��5ь���Qꨧ�|*)BwHeN1�ND�ߓ?�EA`�>w4&�I��A'�7rh�ѓ�e8�I;���v:+���t��V��/�bE���qՑ7�Ч�F�F2HV�η�s(��	,=;C��Bٳ>.�e�v��k���z{W��u���P/f?���7����;x�����\v@�F�1����(vy� �
�T���X�f��]}=>��;��q���ng�B=�(�'h�8jN�]gL.8�χz���i�_쳳+G��T�-���ڧ���9'��&�<N�b�Z���-L��O���ޝ�n��pd�9�f%�S���&�p�$��b!S���k�{<��;	
M���:���H�QB�����=0=�s�'3�/saNWk3�<&T�mvy3�"�� }6̣��ɲ�� �N�I�X����q#�_RVS�[2X�x&����V�$K����S{�"��g|�|d[��k�j���}(�+(ϗ'jђ�um�80w�j+��_ ��Lu�
�8�cK�z]eB r�R2�]��M�`���1c���0f�[	"�[�U挿_�Z���k��׽�5�����"Z�v�����L��e ��c�F���fM��2z�v@�����\U��>{=1�B9(�,�W�Z��@r�.�3_S��"}��c�T������<cm�k"F&˰��S_�l�kJ����S�ف0bXL9+7Ɓ��L6;J������P;q��޲����@=`���J֭qkj�n'|$v�s���2��}�m!�h�M�EPh
kOÂ�ͯ
��iC��%�Ȋ���瞎�"qJ��{O$A�)iG��G�o|��dUyj���UG�?t,T,����,��k���WӍ3J�-�gS6 3�V|(��ineJiʃj�O�ëV:�Yԗ�6s�7尿�����>�x�u ���
�V�����1�/k���1:VL9����.k�f�a���������ٝ���d��G��<��{~���������I?�`�rw��4E���:da�P͜-��gO!Ͷ�<W@yT�Hy⹐CL��/yO�\n'��ij �m\*�{/�I���t"DE��jή�ak���t,����>e=?�p�؜78��R%��m���-iF3�Q�����.�lm^��-�]�Ӕd]}d�	�S]k��w��/�ZV�4�E���d��S%�-��mD��_*�����PCjr0m�c�_�0��JTp����kj90�Ӵ,I�fr�w��!���{Ѐ�Ϝ�o����^4�uR���sY�m����Ѐ@M��lG��7�t.b���
E�z�����4�����-V�:�\th�E��k}^�oR�P�)�S=�U�x�� g���{B�dS��F)���Ԛ(�r3�}�B��h�ڄ�s�+B'4U����	A)�xE܅��.>Nqf� � ��O� j�D��pQ���2��� ��<q��rsi�F
�3�S��:��<;J��M��Ȼ���][S/|��9�1/&��A�UC�G�<���=�]��E\d��F��=ʰ�L��@i������}�5'{��q8"�T��6�}�fzf%h�2T�Z����<�+҈<�<[*a(Hj_}�	}R@Z{��&뇑��9��� �m���F�ð���ݣ9���~�Mm���&��i#�1,��d(`�����]c��&���ow>�u�u����<l�/��O�r(XF������|����C7�u�����.�.)_�Ґ~;N蔶��
O8�+����0�^y�,��]��!.��2�K@����� L�ba�9��Vq6)"C��a�Ư��X���q�t"�<G��{*�zlY�±&�?A���ݧ��3 !V���#�H���%�=�k�(���;! �p7�jx��I�>ldR�C����(�'r��U�In�����U|� _޶�K;�snq�$dv��K_��SW�袉2{zU"7/���QI<
`�����X���%�5ſVy�����U�8�m�u��	�W ,�� �Ԭ����'��b�Hw�}��I�����_�(��#P��-mG�֚R����3��1�h�x�w:̩���ZF GD=_^H���/O�V ؜)�����DM�|m�0�w����ǅ��L�51`h���l,0��&��	֦/�	��?L�pY�r���/M9N?)k�U������� %yWP]�����Ϣ8�G�d!G��k�))C�����0�8"N!@A`y�q��.��+,~Q�l�4�1<o-���� ����?�1͍n:	��}_��k~�ϻ����+���}�����q�z�d�4X_L�/!t��/8�3%)�/�K:ay!���[�0u�|h�"�|���'��w�$5E���aF�]D��K]�m���4��N_'�]�δj�B�P�Z����InP�8!eX��z� tG �*yp�1D~8n��Fn�@�b��-��[^ʑ��[��W<P7�]/��GRw�w��D�D�# ��#~x�sJ���m0z[}ڀ�Q�EVQ�T�B=���3�j�ၩ�1�~#2�6+f^`>�U��;�WN#~X�m����P�	P��w�D!�Z��\Î�`ƚ�+;'�r_!�q5��c���}� ;6Or^\�:5��1Mn۲=�XZ��J���.�/�R�F���؄,�<�$��_��BVht��!��ĩ�ϕ��E�Eԃ$�p�2��!��^�60#�����=2r J���)��%}C��ȀT�����7I2�Cu������S��]]�)�س$����Ь��0��Qp���VLKh.榊@|&4Η����[Zb-`��*"��,�#AD��H�py���È�E����Y@������|�).ʃk�e�<��u<D�5���
Lw+��(��S>7	{ڤ^����v~ӭquJt�����_l��a������>����wA�Z�� к�zO!ջ�T�KJ��7�IztX��?��v�F���p �e�#MCR$�>ך�&-S�3���OgLh�|�|UƵ.!wyVH��ؚ�ă�2�By���[ki �B�^[���&	�LwuӁ5g(��t�<f�2�%A�W@������(O<N"A�M��vɂ�4U��ס:��,�|���"4�f�t��ڢ-Y�c8v-W�4�NRm§P�*�;�^��.�3H3u��m�^A��i��v
2�!w���*�S��!*�����A3��Qz�1 �^�1���P_v6˪����8;Đ ���-\X�lQ��g�w��W��ҷB���|G%?���� �cU����!�Yh���F=����s6��鿆���8+`���!ܸ���d�"n��*��H��I��_�1sQ{�Z��٠��8�����+}� �c��%�=��v�i�6"�q	:`�J���_f�K;���p*L���nL'�I8J!TJ�/,�SG�ӟĺ�����K+��	��ˡ�TNًޛ�Ւ�fGjf?��3�u��ϡ��<�,[���z�Pr�*�F�񏂡\��4h+	-�q�H��j9��}oi�J��k���(���u=L*~�?,�IDc��*ֺ�p"|_��������@��iM�q¨-�PK}n����.2f��pLk�v���_T��DP��E�)���+���Ӓ �`W{8��y���lG[�w,�Sͣu�ܖ6��	�5*�G\��MO��Gt���h�d��H���>ev��'���m����lۑ�{s��KԑU���DЌ��W�R͒n�b��mA�ԉop ����䅷n'����/L�/<S���Z@���J�yoK��@n��O|����?�ځlS�ж]W���2z�TXC���y�w����]��~�("DT4j�a�;L?2�U�X,B���ߺ���)�:CL�����C �?8߽pm��=�F��η�4��\t�R{�a�����h���g���$����_��y��fH���7�3c�_�1��][X� �իH��ϡ|+�>�l��1e�������BcøTu �K���ugAj+��5@�<h�;����
��*�uwgυ�H�옃J��i������F}N��f���׀�/X/���]���.R`c��y�RO|[pR�%Y�ڊ�;�>����d���345�_�,vb@�����f��(&%�-U�r����[A�j�<�I M�~xr3 �`���=gr�S�S�d?b���N4�cOM&��$�̡�f��W�ݼ'E0N#g�BظD[�H~���S��w5k�d��_s;{�5k��Q�7Q=����o��;��Y����!x�?���1�ZӲ��X�`��3n��5����� �0ث��b�>�$t�?���c�6837��\��:�ۢ0_\\�]l�bJ�O|�X���>|)�K�@���:C�6W��ϴ��#�Ǫ�e�~2p{w�5҃�Tl��'NaI�"�O��-TSx2�
���W_��� �(h�Y�Cpt�Z���-�y���y ���9�	�))��׾!q�]s���;�I���	�kSm2�N�o����+�3@�}�e��5e�5�pa7rs�����ޏ:x���8�%��C7|����סL~n�� �Oc��v��nJ��*bӇ\����~nS��d��	J6�9*ё�$��EHS�+��
��G��� >��X��hDYK�
!"<����PLo�3��վq	���"D�3�S�3�+s����ujRn������^�	hP��tQ �>�C�ds�C��|���2�!�tK�z��"��h�j��]�����)�H�8ĪD�ޫ2��Gţ�c�öi�o�����w��#�`�⍰2�G�#;]��^��"c�(��8'�t㭝h.��>�ݍ�^�:;���f�L�e/a�I>j��Y;�8����@���⛘��Ռ��;��;#�a)lj'Omq��`����%���E�E��d��Һ7?-ƴ�k��UM#�����*�^�I����'1*>�޴1ّ*��q�Vf"9��Z���2�̚9[m�f�29|�@����ݲxΝ8�{"��	�W�����5um.�0��I~g�´S\�T7 �=ܔC˞�1�Y��Q"Q�[��W��@F���񋊰;#F�ē7�I�$����z���X���Tɹ�qL 
�?���
�ڄn��C��*�A�3�\���D�H+YZ��ɸ�� ���6�"j�?{T�L|+�C]o�����	]������a�_�	�)�����>��,r)�j�T�Z�La�#P�)v��:�
�3旱zE`���c(D�:�f��B�9��b趫�RD����ÊD�p��X���i��U���C��];�8}�gr5���Xu_/3��	B:�ʐ���4n�����?�k�hbN��j��9-���ّu�|�p�<F�t�;D�]a8��P��@�3��)��a#G�ӉER����E�m�+��+;�5_8T6eG�S�k��t�n���$������Q��4L�&]�T��%=}�!ap�b�t7�.;B�\;{n	�_|ˍRJq:�}�A'���?�*�\ݏ0�������͒@��:��#���ҭ'�̦pTM���8��>=��W��ɉ��
Ѐ[d%a�� eB�~�b��cݖ��wTfo��4��ߒb�����'f��1f򨸼͕��_z����e�ײ��y$�aj��@j�?���l� n3�c���O� �K�/���L�E�|x �������J�Ml�_�F����s�}���4-#��	u
�-(#�H��ع[��̼mue��Cu�]��sug���K�D�S�A��!���ת�M�d��OSp�+`�����(Y��c����w���+l㥍����P'%�7Z���H�`� ��p���l��@G����K}(l���)y��w9~��TɄ(�1����pD,=~ˎ���yi(�O�k�2Ȳ���m�B����'j@��� ���H��}Q����*�e��J֧��T�+�{Ͱs4Yy��ph��2Ӻ��$�5�������$ 9dô%ʆ8��\�����_*r\[Ċ��Ւa�>mV�Ur�mV7��y{�B�`��)����&������x�ˌ�p_���lJ��I�x���&w�O�$ɉ��㊙�]�@����>��I���n3�v$$Z�b���K)){#ޚ�F����:�CLsP6d��E9����&i~c?��	��$�-0��Y��y~ím�x�O��}���3�=Ivc\�r���'�^h�&qQ�����3�}�"䑵T/�*�P,��8}TYGs	YP�eg�ꙇ�jr�A8���+���Ɩ��Z�r��/�8:�$��g��Y�+�FҎ0����#�M��|� �&;�Y�@��X��l�:���6gf�X{����X��{��h�>�戃���������t.ן~|���s;X"���g�bz7�FՖ=����nR1u=�� �H�# �k:/����d��'	$�C��G���ٿf���g�Ku�%4XQ��>�W��n�h�7����$��g �ix\��C<D5�RVV�{Ҷ5��g�P���W��C�<��l�?��&ʮ6��raC4��X&��4c��*pn0�R��D8�Sm�WN���c��n�]x�4�� (�9�R	\�o����Y��?1殦yL�,SFT�\�W�^�r�E (_�_�����(�ؙ���� ^�՞����l�����8x���a��x5�@¿�����r�6��(ɳ�)w���kd3R.���h��i��P�
v?��uM������2ߜ�)�?�`a��K�����}FJ."�A5`J���P<3|�Nw
_���ñ�1� ���I����]|M���N����{�1�k=��X����rQe�� ��>b�S.B��Փ��;z3��)=k.�Gmgk��r��>_�:���',����hѹ�ur�>m^%���M��e�ʗ9���jU�Z�Ɛ�[����9Z�R�	hk=�t#^N��.k�ܜs�?`�����h�qF�kc$�O��J�:+U��.d %l���G���ks�{�#&�G�I!$����������Y�\�J�?Y�?���Rr��:[�s��c�!�ұfh�n;AJQ7@���0J����@������ݫ������ٜP����m�|`)��`��p�o�h�硘�����rW(�q'���^��YEn�˱�&7����V%,��G��?]a�����N���ֻ�0	�} ���)����7��D n��*�h^6��Z	ʉ�rK�N���� �S�z�.�8�>d.3h5ۋ�Vl���j�`�bvEc�x"�E!�)+UR�5��R1�Y9���K����j�v
�B 铅R�z�E#qsrf��:�����	�Q@�	�sd'��,�2^�O@�xc�r:�55l[G�p�wL������?�|��a_SA(婺�ʾ��~��xu��7�r
-�p�|����a:���{y��N�S�eR�QN����1=e�}��1|Ǉ�q$�A�W�jѥ�Ψ��´�R��Pdi}�I�Я���+A������$c��K�s��].���a�h�3F��nĘT�0���� ����I��"w�I,�+�ޣ��%G��w�+����&�����$���qu�@{�'��i��c�'/��_4�B�%Z��M �����~|+�9<��L��<�1��+�JN�d�PW3J�P&>Z��$�z�8duG��#˳��^��&�>�փ�U��	Ca���7�l}�4���B��c[Az��~|�dR��մ�+�[����*���N@C��\�=B�%��욟Ѭ����[�ք��w=�Gn�X�rBϤ#iC4�I4B�]OWi:*I��Exj�i	Yd.Xl۬X5�6��ާ��(�S��G�m��@��*SU�&�Z�:W�(������k-#B�p�z8�͠�X����z��n�����WNF��.�Ź #�|O&�d�ƃ5Pun�Z��cc�AR�]�W$!�u��P���<��h���ω��W�5����m�� �|ݎB�"/�a4���Q�8�׶���&@E?������U��������C=YGld�h�jn_XJXE�Kꁒ�F.rz|vH/�~�Dn��sn�?�
���'kRf������(����S)��᫸�EZ���%eM��n}��V;�}�I���|�<���Ӽ>��GIɏ4գ檊�m�.2��:�����jvv[����$�;n�14T՝������l0��eژ9|P�xZu�?^�1���XǗ�ῄ�1�^s4@k���j�l8S�U��ڜ��5�-�撞�^s��S�x��'�n���F+?)_�@�Z�<���\�#m���g*�#E}L��X�˃q&�F���l�?�=e��+����3�������{��<B��~�� ���+���]�f���'6ո�S��޽/�����#ELh�)5�wn6�2贒|��!:����H�h��L4�@�Q�z>J��E,�;�=0��9M2�O��?��`���W��[���-�G�BM���;�q,';�y��;�CԀ&�0���C�ma�����k������k*��P+V;�0���8�8�
9��D�v2I��Q���(6�H7����o�� ?������ǐ��n�D������MDB�M����Q7��򺆟�A�d�7��cJW[خ�3���� ����$6�������~{�

e�I���-v�����'W*©�X���e��`���3�:}�����6���iМ¾Ev0/�y�&��r�����\ra2���k���ܤP�-�4�*�q��mb��>�x!�9 �6ǿB6�s):(o�e1�~[v�GTMF���Q�K_v��n��f�8L�"\�1�$���x6��cǿ����A�e�Y��3� ��N̋n��)a�����׮4����vh�C��V7�ƸR,ji,�.6��� �єD����B;��՚��[�w��{U�IO����u�=������?۽8L�5=w��0D(�E�ƀ����C���k<z5�]�!��6CZV\�.�S:2�J�>���3{@ ����!�LQ
`�ӑ�e�0
��d�٣i�`�K����#�P9�ĵE�bʾg�Tek>\�%��3s���fM����u���cu���Jd��-��tX
�@Z���]n/a�ϊm�ٖ@_ۘ����<��=�-�@`�z� �T��f_���WjH2�g��q�8�>�@ݫ͑�5�06�԰ĉ#D��7�fp��<O��}����<϶iZ��ls~�1���8FL����i���<�[Ӊ�tB����/��3T�ω�%�s����67�Ll��2G���S�D��dQ1�U��w�F���}�z�L�|KX2��l���N���g��%+��'$�W5�Y3֭��p	^v�N`ͱ� �L�֢���K*O��Ҡ9ՐfV]���/t�����(fkA\ڡ���T&�']1��%�L����B.�>���r�7�4�Ϧ@K�8U	$v�i x�%M�y/���j�=Z�uS���� �ވ������CwY��O�q[:���0jK�ZB0�g�(����0�C'�B)e����������uDW��ߡ���?��=�:9�أG˰����͎h�;M�@��׫q1A��]��|}���	|�	�fi����9��U9w"G t �FR��j��&
�w>�����jt�`41�4�; ��qj��t��&��W�M��mC׻yN�}��n������DS���r�V@sOl�ќ�#8*賆s׎F�1����#�h�Ib��K)��0?��Ԥ�to�M���(�>5���79���I�����D�t���^=*U�$`f��"�JnV)�L21k��\�f��BPxG�`@�ac�G�#l����[�I�A�%�N�,���NTvi6�[%���A�)�^�#���9פ�aJ�]D|�!�\�s�'c� �R���)ɭ�A���$>xnr��u3o9ڒ�u�=s1{٩ۄԻ�x�`�WU281����B�:�t�<�H ���$���ѣwE�ئ�������c�|�8׾Ƶ{���%:��e\6,N�hlEU�kq���F�ؒE,�����и����`�M=P1��b��MC$�|��CU�3�������sPM4�����н����/-V���Z
��
!>�o��(�^�*��e5t���&��E���cγ��w��*s_P&�����i%�L��s�؋�BLA,����,%�L��S�O!'<K0E]�OXx淈)�� ��g���`[<vz<%��Y�M��H�#�����S7�ρsɯ�5-�MT�w=튜��`-�P5��m/����t��>�'��b�"�[^)C[X�\�ڴ_q
ZX��OKvDOZ�'*�#Ϲ5��M4�lB��J+"��C�T�3<��@�Ϣ�ڌn�~��Ɖ)�x�G{d�Mm�ծX(���N���S��\N|^<ǷOkL�|eN��B�F��aC_������
�F>�� �WZ���oY/�Kz��j���i*�<�$���!��)����9C���7���~���ljC)�kj+e�/݈/�!�0�U��kVF4�_���9v�=�Tq=��bu3���ܤ��~S���65<���(-��S^@$7���!d[���a�c�tm��I#.�K~@e�E^I�"���j����w�q�ܩ�LT�qB���C��N�|Ъ{;���;��A�B�e:����p�������g[E֋�Sl/2�P?���&�ʰ����58N�@�Y=#ۛ�h�#��^�i��+5.��:���s���	�S#ik�۶M��_�pA�Oa,N��z��p�3ǊFAD1��s[j������	�y�!��^X�EĽ�9h!�
��h��>N�bB��l0��w�`��J������\��9���J�͍�q,;ã>�Pe��4�xk�l��1-S ?����A<�� #��vE��Qƞ���]pl7�x����|����J�����M�K��E������O�-	�,A���FUP���t�h��C�WKO�HIK+�cc2Y	�[H� .����p��v~�\�����~���^�׉D�Q����C'*��U�X�B���U��}�}�\�2��Ŵ����#�N�Fl�%Nm}��]�9��n��4��`����J��Q�P�u���L0�gь[|�������|�>KՑ$�^=���L��
i���L�Z�o6i��ue3�8��x�ܔ8F�s�
����>��.�(l�ZRN3������(��GQ��ֻ�SJ��uG�a�irXp�}@�B��r-1�.��$c`�Q��X�}so�K+�����r}���囹�S�z�Zˍ��>aW��bu�|��g
'�*��?��u�{�<ëЋ" ��"a��L-��ñ��˛��J-N�a6#�ң���^9���q��\A��5!���{�=�9�0\�:F�?�~Uo�}�G��b6q��d��}*'Շ���41�Ĕ����+ۻr�&<۫d"~����w
n}�(^]'I=�5�٢}�W�T���\ 0ꊥ�G�\6Q�":x��l��Ej�����(���&	�c�e����q�^����N�@`�
�I��6�e�)�i�R%}���{���}���.?�'JIr=��`U7��ܛ��BX���d(�\N�����`�#���R<{�ܦ+�seK��c?��Tq+yؕGq������Z\bʱv�]��I�u#br}[��&C��K��A�J�6ʹC�e����^G}�����i(ԙJͪN{��l"����4M�O2(��7^>m=KH;�Y:Sh;�]�X:c(��I�X��`t�
��,9h7�:�Y�C�?ɻ��z��o@���
�r�i�9�L:�6#��OL[��oOD'��	^&0����8nu9�T?b� eP8�!]�V��j���>K��c��=	|"N��]4b�z�ͥ����S�STKYyq�K�Cy����"0�ƪ��s#ZQ7<]X}��ٗءsV�3��i H�]�K��B��^�	Ys����B~H�\F��pB^����e�5��9�Η:/��2���9�Uٛh�I�����́���g����� z9+8r�'���g��M���( �)a�;"���f���?����q�<�"��lh [	=�������AO�C:q�NxT���}�qW��.}�΍�-�x�̒!��)�Ro�1Q�1�5[O����-�΋s}�1�d�D� #��3A�����k�d-�n��i�Qz�@c�B��2ށ> �;�QH�_x�HRg���r��o�]_3ցi3����򾎧�	����<z.y����y��z_>!�_�������F�z��_�Ն��đs�OW�KU]��
��(0�g�P��F�x_���Ӫ=���K%�I�VT�{ե3 2 P���N:��^�c����d���BL��T��{Ne4�g��eM�Z�mh��`��wɘ(��_�!����� �� Za�������ę^��2���U����u�(z�_;*K��z�X.� �����UI��o����\<p��H�p���Ds��T�ơr�
bf�
��D��G/���o/�o\t�;�8��4T���[�y|��O�<F8�1{����"�J"���{C"~ڃe��O8� ���GԈi^�G��b�뙅,t]s�������	�
d��GG)�:�x��-xʻ�0~�*����Ҿ��Q�+c��DCK7Ww�����ݥ�۴$�|15��q�~Z��n��p����)�K��e�Fsd{>`M瓝����<s�$&�!�j9�o4T�(r�J���O����9}bc��j�{L���j�~��0^��Эr�&�)$�r���,�Nc��4���R�N~��]ҙ��0�-�a��j�m7��)��=1�U9�d3_i�D�f�>����h?)��,`��W�͹�v+	���*���WV���0����6������@�u~�LcR���6+�ئ�m	�u��G<�� �u
�2j�[�) �t}Bp/4�[���,'�VF�)q��q�ڳV&�\��H�D�1v��a�����`��x��2�g�
�˥�!I��0kޠ�ɛ��Q�|^����ׁ1Ǌ�CJ>�\8���β��;������B��
=����������Y�f�+5z�=���=5���`BjI~o�Ȃg�����o�ˌ$�Y�Z��6S+�Psm5m�u�(	��.gjZ7E+�,��
c��Zx-�~ó_\��nt��D~����ՙ�J[���BE!|FkU�-���t���(�^4�VY?��Z-���ș2O�
kBQ޼��^�9�i۝\�� rF3�!�Q0Ŋ�:>�k{��l%cP�S��Ot���=�fS	1LOp�ۙ0�1��� n�� �Ҧ�(J@�)S\����?6���Υ-@��Ukʂs�/Sf���H���͌+��c�y]a��C��YY�A:$L�����B�v������u9~s��8�&�pE�3Y�f��;ݣ��|	���g�ם�צЉ�:e��xx4��Q�	��t�B�!�9���I.��ƴ�)��.�;�ul��[p�>��,��$���2����E��师�v,~��y����|��r{�u#2�D�p�����5;�]ȩ'��2��%X�x��H���Ҵ�F_���	�O�
N��(��8~�x�� 81g'��jj�ݣ������h��FR�/�KDl�('~4nR��s���^�@��(����{����	�]ˎBܡJ�ѯ��u['�N�Rh��1?��H�	䳠�d��C�RHNͯV�P��A d��q�Ojli�D��y�d����y0�v�r�v˞��aFu1� ��+�wL��[d�)��5Yo�w�욊�Ac�&�U �#ʠcHڳNm9�4��V���#�Le%�ԓ��=3�? X<�s�'�*l-�[%׬�#
�a2��R�� f�`��C����5��l��X!Ycu��Kr'�n�������쳡����I��������Ts�i�K�µoR�Q`|�A;S���gAL����g\�m����.�8�n!�.w$�أ|0�7)��9���H�G&��8����\��;�,zl"��:�*���B<�ŰM[b�+�,��h�]t�@Rxr���6n��`K��.c�@����S�X�� �l5��:��+֌9f�mXN�Ws!=%��Q��=5iџ?�ꞩ���]�,<��2�x����+n|�?�8��9c��gAg|e�BɃh�oEFTN-܌<�2e��®m�F���N�6���%��{_n�8H.�um�6�	j�[����y�7�f��m$��^&j�,P��O�7^iDfԑ�,��������ap� GP|2����HGjВo�o�'�_ҏ93_�Q�r�kn�@��R��O%N^<��GA�֥��4\�kLn��e?ݥ�ӈa�|���=<u�C{L��Dl�h�o���鹦0c�3	������t��8��<eZax�zD(x�#�)��8{u>�m�6��6hZ,-�)��DPz������~�[qjî��t�rX�����萮C=�NSB|%�	c��P�t����6���w�j��5��:����u\>����,|�`1u2:	�z���3H�*�R�E���
�w	�B�W�� W�Ж>����y�ʯ�"x��;n23���bZ�nUa����@"K�x.ҟQ���}�y\����SI9ñSր+�]���<wi'/�ˆp�>"I��!�?�W�����A�d{���>|��KtY[#�W���Uh���}-HKp$�OAS�SMX�M*�X���p�8��~�h�s��l�΍C쪽���~oN��~�D�.<�	�0���n$�F�s���m�d�C�v��j�6[n���W�a2F�i��*
z�U�8�J��L�-����%�x���	���a_���0W��5�)!F��9Y���|�,��1N}�y �-+/���.پ%�P���xmK�JOn�?�[���A�dbI�����:��!"�� ϰ��T�,�K!�(�t�`m��\��1�ӭPե=Z۹��c��#ں�j�|��,���F�J�G_評 )��7�5�`N�6,�͇�#�r�`�kix�P�=3�a��P��j?�1��#Th��� ���M���P+�¼W����ѝ�"�!0-j���c�d���6Z�*��uh�������3]�kjh�f0-���r�r���� ܄��?c�e��hU=B�h�2�խ�OB�/�v!eIh��x�\���|�"�ɨy�>!IB��F:+�53�����5�.���9션�[sYx۷�1h���i{c�����p�l:wY-XU�f$&ޞ@HP@l��F>bfu�>͐��<{��ϸl����k���1oyKѵQ��z��Ng�$��ϗ���`�ǳ���#�N`�Jh�=�]6����&=�g�-���@�~�V*8��a��=�f�,�ʥ"��k�9v�n�=���Nd���8�*�:-S�����:Z�T\���ݛ��8��v{ᆝ�6�~�xX	GQ��.Y]�-ٙ� (J4�c�T<?��U�#�9cL�@�'�ͷ&��0A���5Ŕ�U���ץ���j,�kɋ�x+dށv/����t��q�)�zb�䩱�D>R�3�U�S�;*T�뢄�V���Yf�������P:HNdd>�(D�D�9Ӣ�,W
��8m���"�nC�[����L�����2�R��m����?�\�W��.Spq�Uvg���6�3�*a��	�;F�j��K�f������>�O��7�Ά�P�J۹�R��Jk`^�w��˼�J��%��ǀb�e�g\�ݮ$\e��M8�{�F�����U�rQ>�N�4
e&C`M��]���e��\\� r��	�����o8�z��� ���C��T(�<����:����E����N�Lll<=�ݳ�$K0'F��W�AaF�;3ځ��?
�k�q���tvZ%2��s�L�!.�E�Q'�׮�յ��q%��A���3�k=R飸;Z@��:�� 0M3���}W]�׸<H,D�'�M]���6H�����l%�?����P��F��hp���������<��+�Y.����$�����I�����f_|�Z�{00WMB�U�_F:H^l]K[���s�4�.�!�'E��҈U9�����/i����ڥ�-yŨ���!zަ^�h�ut�f{r��-�.��V0,7�a}����e�}����#�4+�n�]�0�ݻmD��{+���>�7.�:5;���Q�v�r_t�JS�B�
w���k��ЭXKvJ�r�\EԐ�S��6�ؑ�=��3��r�o,��f}cX׵;�Fj��`�9�Â�c	���(�R�^�fX]Z�����		*����Q��l�.4�?G� Bʱ�b�<T��`�e+�Y�%ז�>ņx�� ���\dQ�|ӄ�I����b=Ok#��V2��Hm�%��^o{������D�KZ���T�'(�|&�a�,�a@�w�,L5{A#B����E�G��L�8���j��&f9�k�eR�ߨ��*���Sڌ��32L�xgc(�,ʹ<����M��-����A�4:)��[�{�U"u�1�e��dT�G�����?� /���>� 
�f��j��K897�sQ�~��nT�AAV�f9�_�a�y��yGҺ[7��P#W�@�S�6�ν����$�P$�\�ؐ�m`!�u����<�~���.L[r�n*V�#�8<j��v�1�U���hT��W��9�4ԽL�G"�M��T}T
�٩0��{m �����ߊqcH�����]�Pd�e�F�F��X�t��r��
��{��:���[�_��_�s0�%�(�F%�S�7睤a
�9�Ul�� �1,�ޮ4���� ̣��?�)��
��Qb���B\+˔�
��X��hwnF���`�H�����> ,UG�j!�R��w!딎�U��E�w�8��rv�� ���F�,�g4P�杓 �:7*�g5 O}8��l���h%aW��k�	����dу���wc9D�.�U.mX�8�yh��^����)U�
��0��\�	Z�+��\{�x�k9٬ V�|>������`�4��p��?�YiN�e�r�P�K
UCy�_x�ܕɅ	��E�ڋ���B\\�{oa���ct��H��߉~�U�a�T+m���$4����/�rY�PZn��]pRƉ���zT��5��!������΀�U���\N�6�ͩ��=
�dZ\!���p��!h�;>����A��g��SCs��`��en�C�|,ö���[ʨCY�J���,@�t�/[i)R$R�� ����2�p��5V���|�0m6�r��JJ~G���O>U�'�TѬ,f�,"`)��
�
B����t��mO�@s"i4�v��$M�ͤ���+Ύx%��\c0P�HsO֪���9�:��R�]��(��2\^��EoYz��S���z��=S٪��g�ҏb�܏��^E?��`dj<U�}6`YAHտÊ�Y���8PÐ1 ��0�@.&���mT��h�G;��ke{�Q���3�!m��O'6!+W;AR%�<��LX����e@֥eT�dW�Y�Z~��lx%�o��nw�����)�B1��>��3;a�����8S)ao-V@�Eʅ0`O��p^Y���_�O�D�4�rV T�e^Z['�Xj�P�ߦ����,��\xV�_��9����"�g5p8Û?�;�����PE鸊��v:n��&�6{G��}�<�x���6B~A��S�O��k��Rvj)|��Yt嵒�Z t�g�o#d�?�w+��PY�%��%pe��Ld촸>��_/&ێ��?Q`�&�FMy�u���L2d��))��+x�.d�Y����nDú�����8�2��'4��|x��}~���.z~�Wng�g9�u'3h��0��M��}��ԋ@ٳ ��	�E��e������lf��#f�+�҄t��[v�6���}��+sh	gb<S�7�+ߟy)G�"�DJ��ӺLg�Y���wƷ\�8W�F(G�6[�$� ���j�:���3��j9�
K7�H��k��m�H\�7��5nɻ���s�dh��K�/�'��Y`BL���������_f�>�)����nn$3�E)����/]gt����y�B�+��'Ç��M)�/(��	Y�6�'c���)�!��"����,c��H�=�|�y���� )Uh��8��Ϯ8[�������Spcg�b.��ۆ���L&a�'�|e8Դ� ���I����
�������1�x)V;�5O���8N�a����e�itn�����X-V�`��#<�,If�P!��N��[x�A[J�<BA��o�"�-�����O��$�1�w�a�Xȓ�B���x�훗����� �H�u�ӫ���8��F8Mk%X���)yN�ԣ���7zG��2rɻd�=O�d�kb��|�5뢖�F��`ʸa���� "c��|̺e:`�('\u��W�n�p�XAXlri#x�&%���q��y��KLz�:C��%N<��O!�O�6�|�A�Q�1��d���l.{��\t�O��K���W����:"	L�r�~]��i�]{òN�L\[����4X�8��Xƌ���\O�~p�������q�z^Ƞ[���t������%L#+�B�t�B��Zg�VW�v1B:�EϘ8:�fL��R*�M2ۊ�*Ty�B�Kc��~�zF`/�O	/��S��9���_ߗ���F��~�粨b�K�V�w	&��4�J�p��#NǽӾ���%D�$���`wJ y���5���:aa��R�c��J�wu�P:���IE�{Z���]D�'��y� X�0!j�'�2\��]������9 T��
�A8�<��s�Y؇��9�?�Ԗ�4 ��7E4�f<^-����,W &��2��*l�|@*v�i׻x��[��~�{��f��:8lY��Q�.Bم)X����k.%v���=  ��/y����e}�w�����Xd'�l�j��A�ب�o����5�KzQ��gьS��>�&:A��ʙ���mW�q	��w�tzD�󷨁�0Y����ێ����5�<�O��j��}�x��ť�G'3zV|���8�]p�Y��H.=hn���
����=�)'ٺ-rF�)8=�� ,����+����I2��ryK���� �.5�ў)c���<�T[���#.�J?.�
!l��wr��9��c@�17z=���_���9����h�t� ����Z�M�wb|}Du]r���	ƨ�����S��}�m��*� ��
�C�/)0B�)����Au�����(N=�k����̿<����J�ӠT�p���+���o�Z�V�'W�Mr���� �mdD�~�釜�n'�Vߢgv����g�.@}���'>����@�o�*(i��'�7#�T\�{Q�̃���� A䇳ųA��D���MK�[��a_1�Ʋ_�.˘�Ia�u�`G�5J�Ŀ�@�]7��X��ut-�/�x�<����]�����K
c�GБ\�ڣ�m���y���`mq������ַGM��ٳ�����@��cr̆�jf�q�y��'|#�a�
ͷ�m����F-~�Zp���o� ��o:"-��C髟�%���-�j�x�/�b�\��1�N��l�L�i<��y��b��A�G�u����Ͱ[��T�qn��2�ը��I�TKx�^�����b�#��y΍��\��\ˀ��A�ޫ�9,��9�:�t �mI��Am1X\g��.�>�B�1��s��V�8VP�Ih�Pښ�;%��lC}sH=�1���f�س�u*=nOxO��k����.,����N��At�Z���;��D��cPol"L��V��sI$hW؈1�a'Îw8�Zk�7��#�(���(#ҫ�A�U5P�p�����f>�,c\�S3�̍X�>F�[^g�{�XAԆ:J5���x�R���q:
E�k�h�x�z�2�4��(xZ�/�c�EE蘇��b��u ��T��	�Ma�b3�i�p^�¥3?l?4�����Y�I��rj(�����-`܅ɐ�Uw�z�j#I��/F6��77�г�_��b���5dG�rY�qS��l���&�7�jV�H��w�q3%-Գ%������ �[#ɱ#��x8��X��U��8���UnM.R��'ᙽ�a[�]c�k�j�ͺ?��cae>�)E��n�l��@0����|��_~���	�����9��g������Yt��+��
��hX���C�M���{&eBӚ�;1�H�Gj����3jcK�h.��ZC^O�\4\t܂����b:"n��m⸂�M
��CH����w�w~�J8���m�}�
k8��1,y��6��'r���c���^�,�����|�� ��%Q�Tf�kD����_�M�Si��������Z�(�����͜B�YY�bH:m�rVۅ<-{%���t�|�}��v��W%`�fy,	������v:>�y�3@6�\�۠�߉���la���G�H��sP�$+�\J
v�k�J=o:c�x׽�)�fO�PBa2���&����2���]%��q���KNǣ��	x���wk��*��m2ƽ��'@U�1�2-�̘LEN���ٚ�J�R����vU�̴���uY+�z�J��3��gS�E�t~�$Q:9t����+(���X^��*�|#��7�5��J�h���/S��X�&g��o�
�=��wo=�?��l��*q�t!)v�S��D0'H2� U����8y�
�h3<X��],0�*n�dtS�	���f������3x�U뾠�EX[�����"�b�5/bku@��*'�]���e
�Ef>ո��ö���7��(�;
o���ct�������9i�P�����e�<F[h?l'T���A���w���{ӧB���`�� ��Õ��'�Y,�{�F�	��aD���8G��m��r���>�-��Ǩ�g�+��7<)�:����Iode7��H(&�L A��5C��_��n>��A��qGT皮��<�!�4�ꕞu=��K���	+�-eu�=��W�]�by�8PCS�������!\�͋A30�iF�ZS"����3�XqĝRU����":��X�ڥP:A]�HD�l����E�H��%TU���Q��������~�=R�Ua�i���U=�MKS�5=*��@�p�`<],������.�0g<��Ȗ*���5dv�̠������P#||�+��Gq䜈d�<c%(;�biuAH©�T�8V�B���:�e>γ�Uܢ�u	H���u޷>�Iw-�Ǌ�7�,C�J]K���*!���$��D9(8|�T~j`O��&�`���En�jWY�WO?�F���m>�����m��!N8���U��&��T@ ���Kd
� ���~v�� ^�J�kF��/b�7�<��9!��$�4I�!��gp��rsp�s	:�<l�D�>�0��a|r�{�[$;��nx�VV����r�������!G!֏qb�>Qx�>�S�P�Z�yRh�E\&Óoo�QL�Q��W5AKF1�2�i qF�T�0ۘ�@�:�յ�\��3f���&۽��*D���o�//v�q�R���3�1�XecA�ڛ|2�
)*1�E�7UR�E���ڟXd����+�yxU�[\I�ﻰ��9i�0ǥݮx͵�{�����k0�IO��~����Sc�TѬ����ڪaL�U����9߽��3�QHC������ʭ!�,~�m��%3� ���c�^.���,�z��|a^���+��ʀ$ja!&��bO7�
�0!៉�g�C=3�����26>(VՈ�?W��@����[��(�Kލ2U)_�$�.R@�H��·�N~`O�3�T	����_�'���q*�j�_,%'�x���?��*8 ���6��:���i���L�X�[˕��M0>�lj�K�)�ͫ8�%�f3��FV�/���b��?1�)��M��s�*�\���vg��8CƥaN��z��0���qap�Y�mz�$�CO��fRg�T�n-L�9B�/���p���)%k�NV��t�wc��78'd��������'I��(Ŗ]:g,t}�;E�<��e,&�$��vY�J�ZY�􇛫Q�Z������<V�Y��s�~�h� �� �:�q�d�e�;us�	�!JS����e�i �5g����s�,�x6�����/ΐ�hGe'��KC�~�C�t,[�I��&��p3uWH��(.H�3�D'j?������fV?؞�f���$)�����xq�Ô��]8҅�>g����.�shq����&\=�"��s^����v��{(4�pz*j_��s60(�[s���%�/�Ύ��Q��������W'�׸�-Ԥ�@�NMwe�7���W�Ǝ�U7!�p��k�n���e��y˔{5f�G��ϔ=l/O������"�_ka���eʮ�f���N����~k�T�j܌:��z�8�c��+��v�Z����x�qЂf�D�3���jf����Y���{~�)���Z��$�0���f���ɸ��Z���]J��Ux���"y�ܗ�X��_����9�i�F��R/�bX�]�9i�s��D
��,�%�~n!�N_}���--5�B�3�m�C�*0ID���>���7`��w���*�<r��=<�_J�Q{: ^�Ck	�����!��s�<2 C����'_��"��F��\��qjP��
�,<��AA���]�n0_p!��*z�k��SBL ��m9^�̣S��u��>��i?x�%�nڪ���4.�b�a� c�=F���]�B5��6#Em�4B��B�U#�擰��Q��� ~��� >l�$� &V���5�Xx�k�U��\�eh��?�>Wa��pmD�im&��Pʛ�pxxN�r�@���6c���>H���B6eyW���:�ۑ���ao+��P���a��
�Y�X��j���YTH���oh���#�u�+mnٯj�i��?t�S:�0�s�x�'p��$LΥ���-<Ʉ��U̻d�h���h�X*�,RM�t��M3)L�Һ����TM�%��m���J<m�>�#��)2��L+����ٝ^E����\�b�I��E���M4눕g�.��s�CJ��g$Ʃ
�0'G���e01�Q�V_2�3=���Z�Z���}����|4í�'D����k�K������em�Y ���\��H��=�$��C#z��Bv��w�&���=<���i��J�e�(d*�j��ƕ:)lg�H^�E.�J�(�y���~��Q�K�f�/���,?���<�o����U�w���B3IN�`&ZL#�.D�`"�B������7�\�@g��)����O��