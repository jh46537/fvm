// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:21 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Vd5U6Or2KlKg9PjPC+VmCfDbGG+Ha+npMM381UeVpBbwQJbU49eTq/KMeRP4skG5
2zISOyYMMEqQX+1/TaiMNz1GNiypK1PO5eIYMZdWWKfIk6g9oYbVypIrzhMo/Bm5
6Ym5R3e84XMz8vhzVSJRTsmHWCbynAcQtukaUbKGgk0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8288)
qtrFqTD1bL7+X7HPSaYqSr/CeVO5c9Mtsp0h+60ocyTLEzENjDuJ9xCU6LKFrWen
ZH8GDcT6DAAODwYxj8Hoy6hUPYPOQzJ7r2hYtB9RubviXXV1gUikD83Z/aYYgehP
5FajlKcisi6A4N4IxlzXqyg65uKmm38DsULTgFpGAvtWOLBh0kkSfhG8bmc2lVRB
lbPb7/167aTD6465YnT5jVl6aklwdA+pqV9V/PQxZjt7TKlKzrHQC5DxP/7XroYr
DB+EGbPsU6cvCp7s/Ki4nmj3HIHpyqI5tlEPr6zFYPauvZJVRbrcdqyzSXFAmvqA
XlqjDEhUim3phhwq0IDIiZZjHNbdg4I92skshfnSuN+hs0SaqdblVJwSSuXOJIUQ
fb2JefyEEUJPClARKoKsSvDjDRzLDyTwixj7KRi7yF3ZlYCqQd/Q+qB1t3ARY1Na
1yG4AB5yDw8JEQ+K+nBiC/2BYBZEqFulyqCcnWFEm0L/n26WVDXxiPxcma6Zl8dM
CjFhu1AqqwR0QHGxB0nM2KtiGIsbLiIhOEJxqFNVYYVYNYimHZPE6oXpgisR7a0c
13MYP/m1sHPMWOHx7K3lYBODe0wILz8FOdmtMhX5k9kWOdF4RIfQTVLRhxd0Vxp6
B0fGar7+7XFe+6Ma6rrHUa02RnOOnXbKIw0Uru+ql/E8rzApUMFPHuEDOj3RETez
aEIm4JULgexX3BSc6DFuSI9I+cpTYYAAcvQsBgVwJxZzoOTJSQ2Vc/vTmdHz9QgP
xZHBnx9oVRAYtsBdik0nqenGfRHUt705jx3O+QIRP+Hb0ShnhzXKMIOoqs7JwE1G
LdDStnPXMGLvhIMX5+y8bQOp0uNB3CSES41DICdFabCJ5dfERKVe8tz+hGt/zUum
j04bowHDz1vNR4duSFo07F/PtsII+HOquutGeuCA5WdO/+T9PP9DxARFtSrOpYSi
E9Dnj1b0Q2qjpJ5BuCug/qQ96LqF7xdmGOjI8Q8kO9VpT/s8oEBJq7AeuYixmMYk
hy80gT156Pic560N8klIscNFmfDAm5+AZdhBmkJcCmn7tggQN05U5aKbW41VjFf5
r+PMum6hKZOZTw/d9xmeHgyDfrnMXl8eTwiOyyIT7ADyH57Ptqf6uSoptJ8ClbRi
An1yylstKaoRSfDlpEoVHn729vbJh8Fn9JFF61yKFJpz0Wl97Cute5+5e3RC15BV
DnYwzhTCfNE5GJkfQQ2kchkQ3AABZItLC0dvEkeITEC36ZMrpoi8NcK0gQ0394bo
RrCRdo98KgIIQ/CmwSmYmTtzksJD4itQAXLjiGuZ2z76edA16CaR9ewn02UAntaS
HoWJRQqj7vua89g7e3M7lLsTRXLzdALNP3f4S7J2WiWfrLqSBclKN9EpIGm4zeL6
a8LYoN37AxgxxospzJk6vurRxXUgowU67tx0ZBCFLKT78GyQ4ULXRESKLPds1pFj
0ZmSL4s4p+rxE1p9OqnevqOoPBc70wbDMM+tpnGYqPS5oaergkdq9t6UBNyomhfv
in3HqHS3hX25jiCEwQ5PcbOGtD+aBnlN/arZFbwrhZHqKhX09xO3bsXds43svtme
i+m8yBRvleiu8YEG0zJ6VUujZBd1uMUMiR93rIBMWZf+MQeUA5enF0ZzoOK16dJb
9pCgrKCV7a69ZILHxlbdgOYdnTwBjwa56pIVA8Ckgeu5D58XexKLIggDW/QUwnpR
iotCCieY2N8AsNeTNcPY4exY0Gi9GGKYrhyajyLmvOxlN/ZEjISQNhdGzzR9GtmL
fpc7NkHzV+J5Npq7SvlgkBBoj+6qsfUGW3Kc+KlSKs0ApWDcMQcji6qCaWJMo3Z0
rbsVF2J1Cyoj02cw7FD5seIv5hNtDceaYRvAnYW0xFpaYPGD7tisdQl/GWcZgdPn
+cc+QJV/WtMfZ3/6BSRZs9zDhpjP2G5I650iENJtBSPN3T4U5sq97bvTM8FTwbix
QiNxaJe0FSIf6SOUr94PeOsUj0icW3lafsYKXOMpiyrTaoo67G/4/sx2gsdrOOSS
TF+/gklS1tEIQqVctKJLPEA5Rrm/iqWeyWBk938hr63hE/ggD3BKByUgyKFFhjRI
saDF9uGrj5XOFErHLByRgikEsOoO9AIdEnamPGXAOImFVHdbsXLIg4h2YhqpUWJj
fvr64fcJF0oqjz1SSuKzapFYXrHMxx10kehlwrXY616K/Naol3q8LIynS0jvjKDf
+Gm1E+wp1gFFevKKfj98+0DOTAuzJQKZrs2CNLA8Vw19qzXIQnNMLMZV0HpuA1fw
fjyGgLSEzGdNzBQBVSako6wLfzgyEiZ14rAJy5jZVmjURY8kLEUyY1JIIF8E2GQJ
dl3RWvuggW5jom+tKXMus8D4wZr+xV24brwbxLjvlyHqgfJCiTimCXAsBjJVvMwa
QhH/TG78OiLuWthyu1ZLlzwojBNeToeYZvvF48GJRsEXMlgVTHs8N2lFYPvSX8WC
WXL/zQF8ho6J00Wza6Crz+2W3K8+I857Vf40ZZ0NSrAiKyAlvbbQ/u+40NmZNSWP
3I7oAyWSZsoYudTmnSb2/eeCfysW0lTWvwQiavKDc8OhXESpFKZTp22r6/6YO6WC
VqvwPIaqfx+2xc1QuVBpDEStLdblv4t3iRbrO9ZfRgAouAIu1opRYCNnPKtVDzRi
4o6buadJ4qWrZsRxDkybHMrVmpBZ65qyphH03tQHb80VEJ066ScdvnIOtUk1t19a
w67ZnaU53reHbjutJ8xUaq/dRIc3KnIecORIz1AsGUt+to4J3HHl4DNUa817GoGV
dNddG/+5lgFOKrF3DooO/BRLiTUU8LsSnfx9q5pSxAloxzoLeI8CnbgL4xx1B9jh
xolYfRD9xEMZPJOn7hhotb9TFpDqsYq+FizFO5xsOtkKyRpyG6crWcjteNUhlLHS
6g8s377latKI2gXR0yAd0U5PhvyZGUifUsyzb8v4f8EhPRlGCQVNbC5GSixXsWhO
agPcMaa0YRjcCpOSCaTfauy7RtCFOppGHhsWt0uOj+unW7OSEZDPImSmX5QagxqO
QrKsy+l6M3y0/f0Dsur+VRO8KL+Dmt32autK4j3XIAe5tFqGglJNAcS4HerYNzh1
Gjq3M/kPfiCZu7fK+WyK7s5LJCPxDSGzype66vkJTkZuV4dhjSursLWcPTFrtHiF
zbwdlx980As/yn3ynSA+uSRSGTxChBJScIlWeV1azXpz8s02whaaGUec4hICGHGh
TOq2UgyJh32Rldi2I8kdLpwTual0kW6Qiq5zQ4Mwn9zJ/bLBu0T5Q171C6+O7kru
eooyx/+SJMUVFIipttoAqSR7q8VTCdtbhvZpchfLQ/X5WzKczsa2cJV7NQOF2x8J
ZgbpTjYrxQkZ07CB8EDrecUwqKBef6hOsDn39ngNMIv8qrR5cT0Aaafq6mTSNrOX
TfY/SQHP0GAOCO4X0vNtA2nDdcbpjAJolpUrM0I1GFEYL2zDYS3RdB3hQ3fMynmf
5OiGWzhKcw38n07T7SHSV1uz/hxFf6+a95jA9C5ghzVYs7cKx4jnZlbv1Bdt76q6
G2T0dnuDPfdnNC0m3Y/7J2fxHD+4rUq47q7mdxl73a6IUzMh+lcg6G6kOEWDAmG3
Qer8f5ECdAgvwqO+PL5m9wFGfeodwJXpraFWQidPgucP4Q7znLw4FRaoe7SaLKSw
KlHQK29bVtUXqck6JLAEsyQpGf7yDYJddI/yCg6EII/kqNxY2RtEOhvQ0EvQ3wMc
qWa66VY6RTCwXv3P3uQXkdv8+C990zfEJ0Tb9d1BsDtj+4PzybhAm0gntrzknHRf
KGUn9V4n/zrxstGY4CT0fHR2BUHPjhFeHpgT4eNo0NUYuXimEMIOwlWb/73a2s1E
5rQ1xr9nP6mqU4FxuMqJKs56Vq2Tb+9IPfJaLdInRDlQIwuzu07txif3+fD8o/1K
SooFst78mETi+Wt2wjQG3/nT+FrcjaskUE4Q/42uTNeEQc7ckTUNL0+9+kLxViCL
N1Oi4hTYlMdV29142c1FZ+OyePczb9zK1ZzYAWcJWaFmO0V4gDKAGQjxDPjoF6wb
XhFyzBvq+BfXhLuSUjWJJAQvauXj6kUrT8vkEq7/w9Q35lSqHJrtkTDMSdRa1PIf
UQIRDVCDPbBlc9vFa0CYWzutlFTVoMvT4t62KDCp0/P3sFkvF/iyVvcHpJ5O8qc3
B/JodxqEsvcT4xz2idzM/z3gUk3V+FpAvpE2/e5a9cqSEhJ0PvQHSQwaNloJeTjs
TBUmzka5ivMfiW3SdlAmHe8y2nd354KyU9u2ut4l8xdbbUHBFLQxQbSI93z781Wx
cSOi9i31Ly3gs6epeDPFrev7UUMgKl6LBUhyljXqSI0PT1NzmJFtoVCYvo/yaMZp
C+YvP+cVG6b455P6inPQahPvHnNEXQWHPYy4bmneEQT9Ydjhd8DaQdWElpsXDV0W
sA1yhH00tAfwgG7hQDMj6K5JXn7AWdZqjx2wp8XQ/qLyNfp9lzyNqkqOHLQshsTe
j7RumhF2IRv9Pz/vduBD1rYuk0U3+wRzTxu0RqdJLyuEL+VQDD1/3XECy4FW/Gbd
jIk4+oCitEaoUAJrcOZSVWiK8ww74/+Om/1yGYQUHXRptD1kSG84MIxVhpXc8KIl
cq8CYJVAw5VBgW2JyCLS+DdMwOn0ksWZjxY1a2bO20WINT8aIB53vAtadLgxrBtd
0s429hYbEKfKOxUQmYcDXTpdDBPyV5gFecMhKtZfeK5q87vnBSrh+lGStcYyPoYT
K3huo1Hr3+KgLOavQcfvbjnOIPuShkca4H7v/zkwQzYAyzvSHb9zaV96GwrmqMDu
cjpPH7GYX9Bg+NUAI2DAn7lqd1XwkIOUK7E+3yg709xNZZcb9rQuugJjX2kB4dYM
CGvrkcgcKokm9xkgyXNNYrf6XP2gf/wUd1nJN+CKnDKd7i4Pm+iD9trEcPYG7Pev
vm8FcV6K7XZTBdA/NgdaeufNJs8LN+xMTcEkianS1NJYDWci4s1e8fL9oqoMB7bJ
j9Ughak5TRT0zpiZ1IlNtyLDSo5fmmvBpalmjeu8lxYLHj0hYDKHwcdFk5ecbTiB
DbhzH2Rdd6VEfRdM7Egqvew2zTPXBTptomNZHnYCi/YqzMbzlbz+CRbNlF5Ic2UL
JpVJPyqg6t1vBL0JwnETVasG4D4RBu+G8MHBgjDqQcxzqlUFylfoszTrNx9ZuT4L
Ax2mbDXaH60kmMg/7Ko6Q/eWkujysVEn451g7/c+6RhlmO9dvR+Q1oRewuWNTZwV
Gmlx0T97SDRJMIAF2Q1rK3MIYsU7Y0RHEz0grWSr59JLORUtJR0QBgCowYysuDNF
I3qkUIsHKYrYcGXPHJcg/sInWjLht6dKI/HNietz5NVeF8E7/bxuuzYwvKI9Wl9l
JZzw8/kHJf+z82ugJDWsBnekAQgpO7xwDMV+FdOv/jCxJaIgdlmiNqSAl17CC0EV
I43lq/gpTbJJJqf8nXJn+TxJa+gIuyFp5hAoF3b+MFxlBKsQhUJDWLvXMU2oREuQ
vL8inQexqcDoo8h8+g0turcr/8LeDm3S9HEHEavSc0vfQ2U9TYnOO9DDJfFTM4og
LMuNOA5/mM/3lGEDYZhAihZvSSBlT9K5oPvbJVoMLUMxykDc1VZ9MFeG6V02Z/WK
nuoBLtU/3KnxPNq5F8lQwWgL8eZGFrqspPEflWekTh48rGs51qSwOfa1msb3f8Vl
1+Gx1BeSDcTohOqaO3tnRAyQKaW02CaxpGRqtpRUqg1GDNqg0579vqXDFJtluZ2X
z5QxP3WwN1gcsu7QJ06dC1SpzM5Mo0LnEu+68crsfzqcGtIcEfnTjpLvWa3Zs0Hk
zmJpkyVY7hWcohq6wkviHyX4aiH61sXY98ifrieSlNLeDnSDslV4os/GJl4bMX/g
RXADh1t067eSpw+hlnimYsVXaJoAlahFBwkGLEOjyXyUq8/xhi4AndDa5W4k0PCr
/tM973GXx5z1G4vyh8zLml3jD/+qQwzlw6eivLAx5An3z/7TmLvVfHize1z5Mp8K
ckmv/69Gx0Xd0pBZltV3PJf/+d0RfVF+7vy1+BIUd/1sf4uUk5kmJH6mqXDAD3hm
0gKqDjlhnl3B2X7ZTv8NtO8KN7owUxwtJ8kmf25Agn12jem+oTWx2oSXc7Pj+iXb
sKoEbeCC5hb9cROUPsnT3bD6qon1GZkpNa/VxO7nlTY4D62O8fmkUmIp8KGJTu8B
qXgnEbCE2UMSNhYUXtjinoitQOPBrQWdSFfuZGwLAmlRsOa1xpW84xHJ7iohh1NF
rvlP8FssEOPf0CeqZs4rtvDYKDVg9xwyq34OvLL+t13pUBzF67torN52TZ3pjdvZ
i1NkUMzeQhK17HEWde0qY/r61157xhXgH+q2C6w5Gkoz6P9wqLFKRLWpKYTKy7r5
wxjsZr5egsQypJoI3oLkWUzsIZbrv0im+r9ZZXuQeez3w1cbbOcStUZ7MThANJWB
F39CtALftpOa6dyavvXpRs168RU0wwxNKQPqhpkn9DlcKaHtnPESjo3JcgO4Juu1
pKnuF7n4KsBdSIPb98KNkgATKH1vvDYfmXa8wnlmuStmPNpfUziKtEc7wVqAHKfZ
XpsJfILhLgorgi0/CxuxZZilLkHPlN50wRB/kKcpl1340iRaFWo0JfNOaEQ6MHJv
aCMsxPEfuns7/jJXN2Bv9s7S8yZ5ifyy7lwWYjQqDSi8o7knit3KDGaEw8p/lZnN
HYXZnFM7r2vCbwqszPEs2yDe6a6rab3RlfEQm8aDbYgQjBK8IMNYM+vKGqnu/Qa8
+3ONrD3nFDCO1g2mnNfkqJCdtBa7vzxYJYK54sRhGIzcGGpM7msx1ALkVcYfecaS
oBC1Di2k8nfV0wfF8UH8buN6LMV5vqfgYi1LeTlt9VQIVMqVDpDRoWNciDoNPFus
4bEbNHNXee2oDrphDjDQuDzvzphjfpHeQp7tT/EGN9E/lwtbG1nY2G4DnnqYJXHP
8bpkUJ0AVkDLfxny5tgY7C8egHhgmIDj4pUtgMq0fTTb5TB8NTgbQWMXqA7rhrtG
OEWnDfkr45qUCAizpI6XCxeq67Ca0Pff3sj030yD6wYme+LHSEu8XCIodSMkXcKA
NoIgY5PZXercLMfAGXAraX7S74Yvb9+q1jCRmHmNUyTwlun6HYaV42mloNDAtUZN
8WM2skPEERs7iOyFyBALcRfP46eu1P4K85jmWff8f7CI2t6b/J0jYpxlvyzrlKpv
Ngbad1YOlbROGmhEbuAIUGFWdA3do692h3CDvBOQKjwBKSSYK3v+cOvyJZ69T15V
0KQ5X7zia4BRTpvfqpHOoxgqmJJCg8G8jisolKYm6Nn7QTRwyldMlfa1dH7dbE6n
9ZA42edbMJLivTdOiBtB1+writtFuP1la7iCAHbhTBDjvg7qnV9ovgwpJJsBEiDU
NqEXyVSUy0c21t3AR3pEzmG+IANfwM68uyq3W1rLLBh++GkV1OWbdDmPfrpRRw6R
020Eii9XsHfqC6KZdbY6vANpY1jXD5YUS6Z1+0AKMjfqZ8yp0dwcLWGxXDsV/vmK
CXgBb/6ruZZFcSxSIH7+2C5hFUikId1SCEAnJwwO4hfWElPohrMdcES71WAIaGj2
7GWDLbHrs8G5Qk1ZK/PgCcnp/cEfHlW5464glu8qxpLHdNK1bJGpeP/e1l2/jncC
ash10D7l6bNML2epKAqbDuoTLhtIrhvIw487ABVVhQFVo5rM+uGwDhsEtu6iD7Ld
5LXx7/fCT675EDhOSp32+DcBhJU5haOuSVRKVZ+NFlsBhx9VmpXg4MaiuckQMwWh
2rOofyMIMuWvh2zo+U03kGC/Wz931zmsJ8YZpufGGrbTIp39gk8Nl3AhOj6OkC9S
d2RRrXb9YNf33HhYQ8kViwyGxHEn8wNHF+coEk/jptLxAt8sNR0EASC0FhN+2iiB
hX1lF5v0RrVvZUU+9RXUNABe8H5lQbjEGZ1aXy9ZLfYS2jTssqNbPd6yN2BVz4EI
ongtY3LbJnTUIvgGuVGNGgnm4wE6cliJkR2t0jmxyCH+QNkCuJiTJlCSbST8AAlx
SrYIM7OzxjIovWrUakt8oO5c19K+SXy05FTdtzuyeVjkY8YLu0fMNHQaa/h37/L6
semU+Joxkm1F923ynOSyQxl5yX7iUR0l8rQNTCElimuvE5dWmhCvAS6sAH1GVthF
fHq0cLejDdvXXTS1KIiKQnZd+JNgE+PiVtr1QBJ78BPVZCoAyeGMKaRnrSDAhxjw
Fhditaq2T0+krC5BUE4vSvMcG4SQ2V2MoOHyvz8qmxuFmLGAtAkyBvI+TmDf9H4L
x4fZha/HfKcA0WUzcHAM+5z92i8uzB+uoALAGWZNZJnCatQ1EEkzl+sEmQNC4uEz
eFAI6tkyrm53gIWSG+kAnmRzXXdMbAsRhYM1URXLt/lpft6DIE4TF2AfRpY+mE/H
sI+lae0DXmYD2n1CpHnOoxk0fhv2j14CTmCs2yGlCxG4nuyD5Xv72DxMGRcWdfEe
lbNIdmbt8/4Gt8Y0CQ08zk3GqvJD2aZl6x2cm++N6UveKHou9jnAYNkluFBchVPN
ADLkg0OKorEkcGsj0qpLs1JQUTE55HTnhndemt3Uu1QxffZtpwnA0LVR8Bd4HaQ7
dIgrygkn6u7VwY4L0CAcgCIjYG6jS5+fayO2egU2Sa7+YxRAkH7VwNPPBh9mUt0X
AcPFh9rHLBhvcK0UJaGhbvot+y73cC+Gc3I6yX0nAV330b6xRe1xZKZzpUdE4roB
okVmSIXtaUALJ4ELsGYJY8MQC/1TmxhldiFWW+DH66b5eY5Vhw+vFS9AEzsIFkSd
mKvX8xXrCe4A3BbO32Cu6jZEFk7SF/cYT4BPIuyJGiN1HjVf61/QbiDNjcJ+U9Ml
RWqevPgbaHT1maAuJYsgr3kow9i0Zc14bNObzmzRwP8yyUQggCfz6lpB6Dc7t/sc
9izjw4eDacmPvs6MJZIZeJtsNwb8hJuwrQSDJQqj9qF1kciI99epA2NP+9YXR0ti
nGZ0fMUOhGiK4fZWCycSGcHP2iB9Feb7B70drPBLOLpTrLOcCECBaAcuLeOUnCtq
gfl09q6wrz1zyBMHSAisiVNxsmjtJIk24UGLileW2ulULEwX72/hwv9Zw27hZ+Ne
qDJ36X/L5ws5eWrQVXC5LR7xJ+boKJmmEsIxiHSWBMGpsCZkDCNBdKT4fl/3Tudb
XUaOrmGATT0XNFd7jxtfGGJWAfzeaQ7wj/OBQLQDN6hypjAKQJdrBXJayouH2bdR
QAnv3XP+y3FwETaEg5FyXXa8Nsa76FKePBdBg3QTcyhLTT0dPpArpEtsF/KVy0RE
0T4jCRSoxhm1Iu6k6DzfR4MF4kO6yAeOt0SkH+O5KovjPw9pBbjfC+62zq21uLB0
AmCozu/KGay48LNOM23xDc7pDtHIyv5gUVctA6wHbcd8ED8LFL8wLa9BB14VKN19
bdSyHCDiwthh3GafrD4IvVGOHhIJ0aP/8WAnm7HEYALZ4U1OPiIr7W2syuKnvWMy
0ZoordcU5nOgRq+fV2IHI7jjK2wcKGmwLGUXTyndJKWDUh+i6a8a/3koCsgs2PGt
q4+KnC6uC3zZFb0uNgfMYfDYMy7mK2Nun8G9hH7bPvYwrXan0Jcl3zJk9cPLbudQ
7BEP653u4MwcqPrB1dLdvG8tmUhriwlazzGaKCAL10nO/lq6a1m3Micy6Vz9oE8M
+yodx9OQG6ao5vTQLpxK+504hQibPejCEtU4IZT76fyJ525WniA3K416LNDeVW3E
dVfF3Jk06ghRJAVBVsRY0QwCpodrO/7OYV8BwyRCvJIYylB2tDCVSBRmDKLticBf
q3Gq1WPlDAfmUfRVNN6mlA0o0zyrS+bdppLDRb2iHnRTRUMDC8uxtzUlJyfV64tY
drOt3y9UAl3uoEhnETsG4sEPq4Md0SJ/Xma65pWTW3NiLBnO+ijDQbj88c9Y80dt
oz//RyUCABGBYf2Em/KY1K/xb7bF+bJdB9Bk+hvgxh/LNYrryfOuxCB5W8Ik6yki
gvPoykSg9fuCHwkQrQv0At0f2/nJGeIVjxQP/gNsu6qG0hmItoGSDI63XoHZhKtd
X79rM55OXHgVrbOY06Z6pM+A5co3DrakAIzU0jjKYLRbZw17jdE8CmTUWh+kIvOU
j823MR5hDYI8qoWPqeUYTL2GchFbOvoF/Kj0uY+AUnIslXiuAjV2/1KPq24HuzF2
vCQl0yojIR59xB4lILKXRuuDH271uK4eyU/p6ygp32DNbtnvpUunttm4VWc6N9hG
i/r5+/g/NjAZSGZ8vIJjsHo2ueMfGLDETRWNV00DYzIqYUT4hnnIP47/O2uL6Utk
fnHJ1/3c/l0OY1crFAwLXkWDj78nDmSzzGAoxEUm2yeKEakZmjeq06Pc8CZgqeQh
Ihkc8V5InfixL2np+VcFUg57uAekBi7wswGYHHP7RuK8FzXA2fRSHGzZchHi3E/0
5/MfVCTO2BfjQUPONqSKxr9Ocz58v9DLr9PVCPyV8gBo0KKaS8+q5g31jM3kugYO
kzc7jlab8Dyk/GV9ww4dmAiYheK2HhuST4/ZNN7SU1bdehbGB8KFMaESdkWN37cx
Vf9t3khFQ9t4d3hF1lvbFr+JLhMD8N08qTShyjrauwOUJU8YVe/eA5pPNzEtQM73
yN0gGLY0eJFxC01X1fO9caNsaKjyHvTnhyYIAVrqG8DaQ9eu+m2ZWFcwGyItZ1C0
7oPsAXOaITaqM/LoOwmboPgda/cXKA9jVTYWgBTIfRwZREMRZKKuY/iI3m6hVQm7
c8nhO06zIJfQCm0pq2AnJvxv+hY0O7ikU0pY7R8y03QmX2KXpaIKpbvJRX0atHaa
1EFNTLWZzaH9IRHXWfbu95DvfEvEN3NNWuX65HO3CoRbwHsRfu+vEC1yqG7QUvjP
Vp5GRS/4sfEyzsLhEE1SoRlHBDNw3g02Dr+6vCrPBXc=
`pragma protect end_protected
