��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbж��ъ�e��9p�dP;;F�c������w[���}.�d>̨����P!�*W�=�|QR��t��p���'/����J�;+EnZ�v��&fZk�_;h3���ġ���W�$���ݛ�g0T
�7.�m�����q,��;�j��#����E���rY+�>����ip�ԳsȾ����(��6}���)��o�ZM�� 3�kDlz{��(h�M�ñ*n�:��@��]d�)�$�ff�>��H�o��xgt�N�'Hn�INm���K:�ǈ�R�Nܻ
������e-�8�q��H�]��ذץ�ϗS���<J���ܼ\�|�>J�pհ)���j�(��SOTc�������P��A�5��#G��_��0)3�yyqZ�(p��l�b<l�I7%_���tX��c4JeU�A�G��LPKX-��y�f�D
��xRL�ѧ�k�L%t�>Р;��G{��I�WkA�)9��U�Ra�?�e�����"M��Y"�ӧ��nFu��՘�{L!|h��`>�|bA�߷1d7�8���ұ8��X'�O����?O�Q�Q@'�ԣ�|��( x/��Rځ�����̳u��D�
��ٙv�Ǩ;�T��bo��:��L�0$$�H�r��x������N�dԬh+��y�_͎�]��E�<�A�ٳ�x�L3�~��d�������A]��̓_�Z�u^�!-�� ʟi��Ų?1`ċ��v�NbC��̽��e��a`Ĉ$�z�m��cr�7e���W�o��DF*�����C���g�n�Tz1��	j���_.달y��m1�o��$��^DB��N���/������|���g����L0���^�z��J>�l������-钳^�§��Bܺ�8�V��0��ףA˙�-�A�P��Ϙ7M'�ރ����w'��W�Ľ:��@_2�,5z}��=_%����U��(����dP'��c9����ǚ�7�.�R���l��2��2_�q�;% b�, T�Ή�D+9i�Q� [�l8���)(s��Z1(��4��=c��c�\ Y~=k0�0�Peq�;��¿���ȇZv�+0o䬾��9��D�{`|��HQ:����	����>��hm�L �⿢\�8&���78�&}�g~ �'h�<�o�x�<=��~b'��H �Sx"�a^�>lmV���U�#$����!x�O0�{v��(Lؼ��D���Qi��BH�b꜒W��#���#��v�A�m$1U��y�c=��1�Ț���g��sѱ��tKw���n��F1�=�9�I{,��)��H|^J��f+l;Xη�a�Lm�[X�h˼H�R>F������ح��7??��\kc����>D���hlCԘ)���rav�kE7�j��9�Yݒ�UM�Y�k��JMoT�,n�mE��90�bP��|�hQ��+D�d�7h$^���$�s��Mվ����=竂�N���H��8�=�δe�G�'4�t�eȫ0e���� �}�q\P�֯�I��bM���R�q��s�W��W�����>N�'G�,��D��Z;��r|zA�O��E$0T�}��kC��q�~��X�[�3���T�,�I;'�Ϲ�:� ���� 4��X$O�Xx��;6����sɉ0�&�ׅ�D(es
�fߧ*���3������D�[��A�շ��i�x�ZO���eDE���\��;�kE�=�;;��3;�
�4�%Δ��B8����R��v\��"�|, O���7yY�/,a���IWex�p�z"g�vۮ�H�X��;Nv���c e�[����"�)k�(�+ݶ��	���]Qr�[7�3��c�����QTr>9�2-����Z�&8�l-�S�:!-V0��ª�Ж�~�Lq?B��07�%��W�?���1Pi8 Ă؀��jVԙ3�f��tƴ�;5/}�/�b�]��¢E*+=���lgvVfp͹�9�3���T[+��]�
�FZ�g۩޲_tx�,� �n�����`_4�(���{}N޲;1��&M]��w�b�`ĎĐ���d�@��xw��h)�Mak�o�XA��툙��&�����h�~�y����t�L�h�H"B�V,M[ߏ��K��2����,�,ݩ�yi������ê$B��5i&��)� �\h�u���2��n��a�	Z�_1rU�,���;$�gɡ��}~��!�^�Kʘ��>֯*J�{��א�e	!��X�y��x�9q��a�2,x�%��K�����Y��W�1���J��ؚ�9~J�Iq�:+���� h���N��<-��� ��?jm�c���@��p��Q�b�$�f΋SPg��b�p!�x����
�������Ra�]��z�/�o�����`0	��/v�Mkwh�{r�j g,�j�� ��5'ԗD�"-��N�G;})W@���e8$>;M���>[���h��r�s	��_V0��w�n���b�3�|$*�K���Z�E�l'Ԁ�ZB��}Z)�6��=����T�T��Te�V�_�\Mw���_.j�`¡�J[��uB�����{�մs�-�apK.@�=&=��6� ���w4Y�+AL�x�O�Ao��K��i��
����zT���j��c�^��6�O�)�	��Pϥu���֒S����wԓ��p�.��6Y��AsbSy��q`��<�g���oʗ`i+�m<&���4[A�JE��"���'����nGU:2�Z�vs��ȧȀ��@N ���]k9���v �䜁���Y�R��~Z���E�;���n���>��N�[}�zY��f��a��	�ͭ�/g��S@�ЩT��r��E!�Bq����]��<�L�����?�n7���P|��O������`٣4�5����,�����T2U�^2�z"��t���yi�K��=R��]P�T��X;Ԓ�Z8w2Ln�R_,C�l<FI��:�ޥ�U����QM�{��u�u�������fF)ʲG���/J>�t!��8F�i�	�[����DX������|S;&u��D3K�4;(�gs�xT,1���P�s\³Ԡ <p�%�
PZ˂p9�1Of]ފs������%�33�#Q��ro��A9(�I���3�����{�8�n�d��*<Wh�	!XfȄ���FͲ�%44w�H�� A/8�ꩽA8cΧ�m{&c-���,P��ּ8��;3�d�	����k�*��ǀ6M�������qY��X�UՊ��}�Ж��E�����H�v��nS�����ɳy��COb���&�E�2�|`�m~N��
j�/9�M��iPK�h�$E�M�^4H���E��4�Q���g�_��E!Ć�"��5Q�֫K��'..X�ޒ���]�6��W�:�>�����w� ��T��J��v�5}�m�HҌ(n3��e��՝��wG�L��Z��S����f��7+и\E/uԄ�o�.>�l���.�TD59vQ:ĶgI� U�Ll��զ�vbհ-�J�e��sT�A��Ex�^�t[K�r���Le�� �$!j���sS`J\�կ���L�� ��-ȁ<Ux��H�}�$��Y%5�4�Z\�@4��1�U���J��h�ם���(�y ����(q��;*�G����~�����ѡ�n���N�����v����_��'�%��)�����?M���g���?+hjk�4M��3O�Ox�'�y����7��� ���U&L���@���yy��5P��@��:y5��U�O�����^���,%��PX��"�����k���Uu.y@3m�ܛ~Mm?��/^۸ǡ}�	��@��
vK$�	?����W�<D2-��yi�����O��8�f��7̈́@W�s�Z��W��P�;�oH䍻6cg@�4�<�)�	k2|�=�����'�zp�uv<c�ps,x��1(6O��tq��Y�dW-�n��``	���`�1
�KzS#Rd�P��6��[1r����70 AϜނ�v�g�b 3`�˱�Etܢ >�A90,�Q�.�kg��=�~^���\�w� ��W[V��)���o��?� �Z��n-l�}ulb��n.U#�r�g!I�ڽ���@	�x5���H�<uXI�z1�P�(�4W���_O �ɮ�)�W='�YT�=�m�h�5UQ���)��6X7�&������f]H�7�R�&'v�׽�ӎ�<�Bn���Pu�SD�$����R��=�:v��/}��/$���é��9(�m�M��Q�����>�Wx������lu�^��N,�����t[`�T��,z� >�z\�l�$�G�7;��͟Hg�����.��n��72��,�"��)��Aw�.�T۳wZ(��3ݏ�p���S�O
��Ԁ�iL�z%f�	�ؼ|j�3�l�;�#�������.g�4ӗ7�vĤJC���(�Q%z���)�ܲ����ZX�y�mcR���$�Z�;"�_Mm�Ղ3n_A)<�`���+�V�.	 "�1���÷��}�B�jo�P�쳼hPֻ�a�1p�#�"__�4+�$J����;C�WNhEzQ7w�{��y"����6��e�`�cUx�'Vqjz�����O��'w�{��+9Kq4gqr��.��#�ߋ����-�O6���Rr)�46-��]�č��+�x��LM(��{9�6G/ ��Q�kh�uMX^�}H�k��)�lD��z)^���1���i��`�".,8�ֻx`!�X�a���A���.�<�I�4T��uˑE�7mU:�����n[ΊW�6�&!.�(�N��vA&m�[���<q���xM���cot2�>�-M������=�(u��sD�Qk�# �/�Q�#*�Ѡ$��K~�3i��g:QX���c�)I8��m�(��K�j=��f�5���{��(L�TN9��v����z� �l�q���=�K�ߪ3��d�z���ӗ���*�`.���[z7��^���R9����Q�U�Q����P�S�yE�˛��m勊���Y���K�
"_�0h0��|���������qT۪��|��C *aeb�-������b�Ytg]N�T84uEtۘ�!C,�x��"i�C%�o�}��.�$`�h��T*��f�6�3���RPĕ�QJ'D��<�xT>�	��#�,ۻ��E�YOii\\9��G�Q�qyn(xCϰ�3�&�<f�	^[���1�7-�_J�4�x_9u�z�:�)4��3<��:.W��jg���:������%/��k����os�R�[`}A�'\�|� �υO{ʫ�x?'�1�:���5�S,.��������^�.ɏ��tԲ��cΞ���w�����P;��9]c'�S��:�v�@�����$��{��|=`f��fL�8g���*�$-*l��H��=]�H�Q��ri�C-?l;�0�fx���N񯮆5�Z�S�9w��61ޛx3����Z/�}�jPm��_�r�1b�l�u5J,�p�!\;�����g�9_��&�_������w�7����w[��F�B��\&B:�Y�Ik`VJR�^D��m�!Q"G"ފ����;֥��6�CG)n$&��t߬������Q'����<&���\�v�$9����@�T�z��Yg5 ������jV���5��j�H.�fK~Ǥg{\@�%w���6��Y!A>1xX�_��)������G�UU����lj6Z����2R�V*j��5��]�۷�OS핲
_��I���]����9y�U�W)�����" ���"��ȧ'y�C6w�#:F�W_'�/��������p�?�UK���~\�r.-�/�#�s�|�Ǻ��C����V�C;�L�0���Oi�!��,��3<�'�L�@[4���M8��zyP/g����_��E�<_:!����[p`�QH��5�ߑ��*�G=�b�qF����R�1���? �,�ݰ�C��H$_6�4�����	�6���'��@�SD<����Y_�i����8F�WGD�����1���WP�� ��GkK+��|;Ut%�h�������*Ty�Ch`4�E�w�D	��6�'��E�A���©)+ G�O:9����v��oH�;���j�4�5e21Rhd4[�Syr��$"����w�!������UQhZ�Թ�}�DL`hq'9̈́�RJj�⁖��s3�Vz��Um����eH
�J��O�O���?%�[7�Z�A!LU�n7B.*j�����	:����i� 5��+�LW��"G����O�2]J����w������Y�6�9l�'�C��YihY��~��.ź���]\�y[�U|.�* 4�9`��5ŉܶ�oj��P�*��O2x%�9Zi˪b܏*��`����9r]s�E�eژ8WjA��DPՇ]%�J�:�jN�VM���T9,͟��xޚnG��׃���f�7��k���S�*%�˧r�?F�ʌ7:m���ȷ��d��>C�+8>(CC��g��V�|0�
�gR.���P�Us#��'���;y���ʈV�F��h��X�=���S �3�W/7�����G��1�r����я��3����S�!��Z��U���$x"ɹ���}}�YZ�_0�KI�=J������C�������i{� �Iߒu�Lg����y"�V�T�_����s�����H�C8@�,Wp��Ϡ�����Un�7��@c(��ƈ���dË��C�7˅b�����u�RpR�z��\�LV��� 	�Sz1Iǫ�W5Y]N]��M�$u�iU���5���*Ui�c&�����&�M�
^\�v������֑ )��9YjR�����n�0�Л�Ivz1�����ђ��FB0���^*6-��4�#(��O���"#Ĩ�9��k�i2��T-�h��]�QlO�Co�A�Ʃ�fU�*f�j�a��^�8|�O�Px$�%|��g�:xC[��q	{�\
�j�!���,5���[�Ǔx^	$�%X�6��Õި. b���]N=��� X�Am���?���g��A9���ç�H]��bF<9���M_ٔ��Z������u�*�˸�>a�]�mrX�ҍ(X)W*^"�xb����&���q0g<č�瘗�