��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�^��h�����mb��feE���0�8GI\�VE�|E�T	dݹ._lR<���<ߵ]�uj�x i�(0�|��� 
���{�G�i�S�e�ΨI�K��L���g@RjW���%e��I���+mv<�S�p	�ë^��R`A��-P���(�ᲀپ��Tem��Z#�;�M��`W[y�(4���n�y@V:�+X��6=+=�DJb����eֵ�Y�l:w	�=���7��_����-���� *�����e�K0Ś��}%d�/��wRa�NCd|6� f���������"ѱ7�s��r��N���������l��
�૥ X%m������ �
)z����^+�TB6uܢ�~���%DX��t���o��&�ӑ9��9��pc(~B/�Y�� �q�+��s��n��A���B�.��!��͝9Ar՚�1���#1y�X)Ϧ����b(1H���HJ�29���xf��GI�..����ΦrU�	�3�W��NGM��ߔ���i���o�˞���Q|:!����J���6�~�?����x�R���,IS�IwCY5�̻�%b�b�GW:�r*e�t��Mom�%��
�1�z
��@��/0Rc���W蕺�v���
��R��.��К���xҼW-[���d�ޕ��t	�{u)�/�n�g�Yn�PD�\�4:ud^?ꥤ�|+>�7g�P���P�Z��н�:ހX+�i���;��2�� ��'Z=Q��H0;�&qx��$s,졯*~�L}܅%f�KlrB���I�#>�ܟ�`�v���ۺIC�_�׈�݅�a6Bn-��p�?���l,[�V6Л�`l8�$B�)b�.�������<N�2Ы:^�!}��qv)��8��}W�����
[����:�˓h� "�;y,�ڜT4a�Ҧh���:�9K�T���Mwe��N��8��#��?�^�ӿ�����k�=oR\{�,M0�5AO��ǄJ����Nv���I��r(.V��dT#pߦ�I���Q'��?��g��B)� �â���+/�<$�T�49�vj�p�-�n=�!�3+�/t�i*NUSB ��yI<z�]�I�_^�
u:�z=]qg��8��@O�uS��ilX�$��V
	���8�^� ,����k��lf�,���s�k�JO��4�,�<Č�80:yDX�x"#�x���n�t- %��P������s���Zi5e��o��u|E�!������7��z�H�1ႁ��t�E�M��:c ���0��F�C�m�Dv�&���j����誛��g�!��Uڀͨ"�%��}�2� :��ߧ�; ���:͸�Pi��>����@t�G5����B�oB�N�Ӻ��].1E��Dcȟ��!@2��w۠�2�Ӯ�$�Z�M�nӧ������
��͛�;(zn��g\h�����WQ@$~�U����`
�Z��n`9J/���CT��o��_��"j�J6?�<�H���f�6`,�jk��;��Vc���4B���i��K}�{}�zyVbSv�n�l��rɸ!��Ag�-B�b�)Ks%J�X�%�(IZ�h�N+�`�����k��U��P�G)��t��� gy���>. ��"��������M��*�t�T�QM�#{��D�ᄀ)�(�M�p�
�t��y�j�h��@�Ţy�ρ���26��;"/�7<o01h"��k6Q��e+����n]w��4->O���;l&W5�,9����p������VX��
���5��$!����$mv�Wx��;�7[8�[b�8�ڐ������R��J�qF�f��`͡_5vN��(Ƿq"���	�qt3��^�롚}�@��L��T ӹgcOf���l/�����FO����|
	���c'ց��vp+T]��]��1H�틷��q�ks�T�D���V��on�-�&����K~sI\��#8{<mԵ�9U��������݉C�(͙�U�W�������T!��]��˸��ϖe
�՘o4���[�l�U�Glg����lO�9q��_�
T�����mN�w���o,C.M��ѭ3�X}h?�tV�y��^I�*ە�`Ӿ;Tkg���v���ܐ�Ťe���nK�AE?"�U$�\J]w�Z(�u|��N�ʺ�fJ#�n����G��~�uV�g��;>�Ѱc��K�tПe�9 �. �7�~��,���-�o27���A!�٬S�%ht��z ��_o���U����!CR���1��ke��^d�Gh����z�����Hã_�?Tw3W�s��Zќ[>۷�r���٨���R1���D���|�_�\�1?��@-�w�wDb��U�#v"��� ���������ݕ�[VF��dVN2/z�F6q�����)!�V�̾�2Hrl�w�J2��r�Y���ߦ|��K#!^FT����R�/L�AvB�s�E���E^�B-�&h��ǐ��4���O��� 4Q�-�>�*~y�i���z&�se8����h:��ۑEu�����QEp�|U�hC�����N7(������N!��cO���7�-[�-@��V���Ӏp��,[�����d�{WH��"4�~b;EdɒM����+/'�C�P�x`HJ�B����RP�CW��I\�"FV��y��H�X)k�΀�r���G�u��xk��u�����?)L����[�Ǆw���Ś�r5�A�{oqh׿5��Bl+�`�4��"��T(��p� w�L�$U��9��wʔ� �ݎ��EwPe�f۴i�z�[�Ճ��VƝ�Ȣvǔm����P�V�����y�纫�$�p�ç���'� ��5��,q�ȷ������ic�/��-��^����Ot�Q�]�<]̏��-ཛ�A�Sd\#BzSРxA	f^��	B�A����"�����G.�6�t�p�e�3Ӭ�b	Qڟ�m㋻��w�P��m�h�PB�H�ZDd�dsų��T5���3�$�r3$�"ᯇ�v���wfS�l'�a��^s�����X`�X���^�T��"��h�eKǥ�r�~U$�S����G�I@����?��#:�W��c��C)8Y�I���q�3 1�A/�[>WZ��Al@Kg�#)9Y�^�Hf�Dm>�P{e���Fv\*��DX������th"]�s*25a�]��������`M�ε^����u���>:��+~0���]�|cդ�V�l���i!�f��:��6��2������Z���bp���t -���³'�f��[��.����p�<�wr� 93�X/5���6{9����n_���=���t��.][�AVp�'�|2�N�	X;��Tu�S���H�C�nL��S���ӗ��z&ʾ|�D>����[�j�7v4���B���Y�!���r_j��_�@xGN=�\ONY���À�et_��C[
��
��+��neNyJ���T�ʄ��A��q�~�g_u�����u��CQJ>TB�eA���y�$f�}'C$Ojd�/@ռ̩�%�V��BW�����FȂ�tL�JE�Ma�� _$�e6�/p艷S[	Ff�7␻p�M�S��	حӁ�x��/�����*�&�0���P*�(ssS�/�f����U���U��P���W)| �DX���&x-/ΰ@���+]Ï������y�� ]�Ap���qO�b����|+�$FD*�>对T�d(1�e�^6毹�St0c�LL�c6\X��l�J���֝�g9��g/�Ŵ��ʫ��TM>�?�% E��f���@�(C`s�_���'�%L�d$g|c"xO��rp��P��ķΩ�7b(�t�Ϧ��R���}�:ʹ�wZ��	��>=eh�"$���5���/(m Hv�`d-%%�� v��U��OB�j"��꽐�0�{6m�|8��E���}:v��L73�N���$qK@&-eK����Ԝ�``�j51��s�3e�q���;��8H$'�K9ΗL�Q|�7��s�'|yv[�4DK�:]�m̯$�+񫴬���%2l�a.��r{�N|E(���v?����AM����u��:9�D����=w/rqA�*嫼X�<X^���;!@l��'$��B-��y�D9.�_���VDUn��2�O���|?���g�#B.��^\���R�Pϼl��v�7^�0��H%{��4�U%
��5V��=�1'Qf���	��=V���|�1m����o�m�2L��}����6����� �ooxI�j����{o�[|��p�M�f��g,Wa�̂d�L�H:2Ε6��!��C/)����r����%Nc`��1��H����c޺������D��L>ֺCL��2���3��GM�iQ�+��(5�[��پ��&_Z*QX�����(T����UoB��8���}����:�c�ӆH���W�2�4��/Xh�E��w�|����W�\�JW/�P�0�гe�o!%��$d,�F!��G<�pT���{@��cn�!���\�OS�E(\m���k@�O�~�4.)A���	b��O���[m����3��1�7&���*1Y�.ɟ=���'���J�Af��l����k%��fߠ=>/�� F.�G�V�s��|S8܃H��	�Ko%��o�4t��3��ŵǺe.�w��Ȣ�Z�9�eBD����{"�F~�I�nƔC&CPbXkl��n�<7�j�D��εU��*�6��<llE�*C�8'��"%"�@����>���0*�'4�4��d�{��zʘC�U�&�&l^f q�̛�p�v�я�L��i��ݞ�M��ܸ41�+`�����0�M{�̶������7�db��C���XL�<-%D��3E�lY��x]��=�_N�A| <���6U�8HnH'K��&��۟i��v�n/�c^�܋�8�IՅ�M�� �ZJ6"�,���Ȃ��[( ��;�Pm o�o���ny�M�YhO_b���S�5�gv�Cf\�R�Ā��wUH�b�ևҲ�<��/�&���)���P@��=ޜ��J��¥�����4~���+�_��]U �C��#g����j�� �^q=���.$q+�Z�@X!��2X������K����R�խ;^��5�-�!��t��x�dZ2$���)��*=�X�\��N���<n3pT��Ek�Y���"��Ī�g!򳦙p
;��nk�d���is����z,�-�����ƕ���=k�*��9S��Ijm*T��r��%;�jCoh�b��N y�ྖW��-PU��&`lMⴐc%1I�4�>�����ǀ}�HaU��d��t:��D��X'#s�
<b؃�����NOhw�^Q�s��XQ1�L1#̞p�\��S��\�G���^b�x��շ�K���%�3S�u������bS�J���o��d�wn��"F�W,*�b���5%W%)�.B-uZ�8��p���1���Q8�?Q�N��*N�)E��v��/�[�]���X���Pj�݇q1�zz�E$�Z��DҤ ����M���/����Yȼ����B�����g����!e��,RJ���`P�PQb�@J��E�A���|I�Z��\KKu���e�O3H+Bs��c~����-���E��Za�T�N��\�%�[Ń���ά�;y�ʎ�yl	���f0�������W��y;a)��E:�|�y��)�sZ!'R��`�i�F������@e��47��lau��G�]��̱�m���9��a>]���LH��5�L6�����0�Xn�`�:)[]o�l�'������Q(޳2��F�)�Z��}���\�eA�Ȁb�|G\�.)۰�󋵿�~~�:�;A�۽�������eh�P$#��C�����N[��`�&�,a+]�y�?�uuG��?%�0�zKAQ���bz��?@�Z��6V~���S=X@�ãM� ��,"J�D���g�y�oKӤ��)�9]�F�k����ˮ4@G�g��N|� |�AR���GʩJt���!�����8��H���%y�LF^k8I�AYh!ă�v-�ݘ��։���fy���;�t��T�퉥"������s�}te\3�x`/ܷs��=�3Q���©�ڞ19�5E`��t��	Q��&�(��2p���K�"V5`#�B�?q�{tEl�ҕ�Z W�ÿ.�Ou�J�j-�X]� ���#Hmg-ϙ��k�W���V�([���~;��W���Ʌ�>iQ�6n=��E��Vnݙk��(i[N́�x.#(�`�Ŗ�1bM#
�Ü�Z7�����%_W#w��F�H���ۀ}?\.�z��4�UEW�@}�� �Q��Nj���
6d�La��]��V�I*a�ݺ*k��;��Q�J�f��{�5հ���1z?��Zթ��x��f���X���R�8���A}��LB��au��g@H�HgLE�5�����ǒ&H�FV�E�Ԫ�ԨX�6��[]��.`�C��0��MO���������Sn)P��ve�?fF��JB"9��' �%���ɩ�^ ���'�V'��$�m�3�p��xFh�H}�aЏ��a�d�P�{I��x�K|���?.�!�}�x{(뀔��bI'���90EeuW��"kzj��p¾�6>W�l@;��؛�=}wE��=�X��<%8�7��$݀a�GsD��a��8"��6�)+0Z=ɯ:w�bpz!�b�7i�c�2�BI.Sr٘��
��v`J/V)ggR�[N�����	�:|ƿBJ~�}��RJ`:Ð����SE����IUr�@��h��- Ѵ�V��k���X�ҟ-
�����_R�ji`�*���D����G�?:1w�pG�Z�b�4��'c��������j�!��=^Q���[�BD�S���J-����6�b�e�0���y�r�G��$�۵��7�LP���U��F� �/?=����a�=B w�ir���p�э��ǩ�~���n�2��rN�r���	�ت�>�G7��&�`b�O�Uկn�Io��Br��|x�8]O*���z���D���%9�/*D.V	�0�c�Q�j�Ɯ͚��3�n���,R�e�$P�D�8r�?-��K������8z9�����9���ĬB�e��l���CP�u��N����4��/�G\?�{�u�6��6r�����⼏��P<gJZ���"3��O!9x��KDP	Մ�lE�㾿y�.c�a�����І�[瑌�͐Ph�33I3Sv��w��h���1B��3�d��̲�,�����J�׏B,�x�۲�3U�:yь,ԑ�����O�RPe��H�=Уڹ��P�׋���WF,vZlM(l!�X	R�86������Z+^����n�];�����ؙ�!�&�np�
�OC0��j���쵶������]�v���I�`�P���_�u�v �}�<T-K����8nK(���_�Z��X�-_�*h���Ӏ��}��l���;��ҕn�N��̬��j����q<M����dW�Bm�s��N���<4c�R�A�޺��!�����٨�6(�KQg�[��ԉ�WEZek��i�&���(H_|�g��S��(g3L�m ��]E���!��w�û���*Z�ѓc�O[����rVڡ���N�p�C�����,�� ��,ZV�M�3����Z��j����Ae��v�eA9�����ص�Q7O壷R��P\�� �=�2}�ɫ�w!xÜ|��-~�H���l�!!IA0�6w����3T����Ff���R�c�^�
���m\�ț�4Z�����A��SEy��U��t�&�3�~�7�o��4��l �,Z�ޝ@r�
! �X�B�v{݅���*	���U�~��I��W�bᨥ&�h�f<�����j( ��!j�57=��_�����l���R�4
0Q�}�y���e�#n��k[�K�(B��#d=7��w�b*��{Y��5�Y,dӘ�mg2��MKq,���f�C,��h�~��c*�V���b�"o~�^+�K?���F '{�\9��Jji�����A��K5^f1�+S�hd�1�#M�xE�l��`3:�u2�`!��-����V�G6�ʀ�kWc�/�e��޾�F)����]�@�Y��z6�D�hX7��pn��p�q]�n�ӺQ~i�L�R}gi+%�* �6��Ǻ��ٞ��ڣ!j/�Ɏ+�`�=���V�Slt����*فP��"���?n�C�=�_�i�V����W�/H����:2�b$�J�b�}��l��ζ,\o�;��)���gS���I���$Я�ߧ^�L�����l۫:����D2k(�xE�t���Qg���QNF6�����u�J0"���$�KX�=/����!�9�P����r8|8]_�wIc1`L���ݦV��<���������ˇ\�E�'��Ke�&4�c�L�x~�����!{��G{m�4
zɻ �H�ji<�}�%�G(�
��J
g�%�7���u��5�z�	�4�LJ+���u���j�%�uW!ǩa����+m]�B�&�a�+�_ۘAB@��G�4����-(�:��i�O�QF�GrW�?�9b���:\��~�W�q��I�`Fxz@�3�� hfF�e���_א�d���V��O�M�;XjKVuw���/p/��(C3"���>V~�Z>+�P�L
��/:$��(��)1����el�����砹u���Ɔ?"%+ ƫ̺}|@�ٮ
�^`��%^�΅�+���^t��TX�]��L�2����C��1�J_��¹L�]>�X�:~�-���a�G�#*7���vD��P�/�!��·�k
%;�?���[�&������j�X���F~�`�?..��R�E�#�f��p�����Y#W�Zſ�6�[.Fc�z��2D	���&���+~2���
̐+�?n�<��'o���΍T��e:�|!�S�v�=�e�M-6�g�:�H���I�%�����������\l+9/���B:�Q�:��%��� �ajS�2�����U�<�%��VU�s�[�V4�w�B��Żl�-rV���-���\��uKqJ�+sc�����G�H�\i�^F�bO����� ��) �9�21xN�97��G>g��h4���	h*5���_����L�O�>����dRx�TD�-gg�K�یj$�+E�5��q�(\ٻ׶�X�YM�D��c���?=^��6�U�b�x��=أD�Ktpc����f��|q��Z��r����R��7.^Q$�\�y3d&w�e��ٺd�k����*M��J�B^۸b+]�1�K��
X��I0�0�� hV�w�<.���l.�zO+�*�<mydC�#[=� H���b�Bw��d�$�@��3�Ӑ��+фQ�<o/�([T� >��Xy ��g�1cg)Kzf�A�GE��A�C�g7�9H���r�urb���@V�	(�<7�(c�l�|��<ޣ�-2u5>��M�9i�-�	�t~l��iO�=�B�ş�c��ZA��~����ٳ�n@ݪ�k��Ke����Ӊ1����e��}�����ƾ�E�zw���OZ��T歐#Z�i���X�\��-W��/k.ЈKz��`{l�Xq�P��3Yjvg�ԃz����oO����|���_��(�&�.+��"�#,�J'�|'ϙ�x�gUî԰�N�颂b"�����"���O����~:WIb!�ߤ� �����!~, �Y�ЩXov^.��y�C���14��تI��
����ɱ5��H �u���^�]�0P�O?��a%˝uƟ�;�b�ɳ2����s��ҀY"p�[�7���?'A�i�r����P~��j�u������j�����Sy��'s����xQ�ʌڦ(k�O�G/��!�֣8��68=6l���ܯeu;�q.m-y:c�t��H[x2��*6�8v�I�|c�T��-.j���^��%	���n����)�X ��^���?�\ߗ}�����l-����6�TÈu���ī�p��'�G-�(#↤�?Uzw4�!�!����I��H@�N�y�k�iBXb�2�Ʀ�Ol* �9�B��1��s��T�B8�k���y�IQ�r���� ���\쳛��Lwϯ�����,W_��4ٝ���d��.�J��[��=�c���\T4�,��%Ef1�cے%3hM����g�;�#��L�ڙ�v�!���g��&Q��K��N����(���V���Mi���� ?�m��9��`XYΠ-Sb�W# @�YOg҈�iq�"����P)j��5}�2b�
���ea�y:�n�/7>�ei г:'��U0L�u����_��яa�Z��T�=B�و�s�s�L�V0.��@LNJ
;���_���;��O����j�=���:� ���7�����IS��-=���kۙۯ�.�HD20A6�
F�1�KZ֭��^{P�l,�s�6�/7�u�p��թ@�mU�5�ӂ�	ISz�w���R��5/�p�8��)��
j<��e�T�zH�a-te����ʸ9BŞ0��Λ���f��n�7����vf;o�\�8}�C4\G"$�F�=���t���_(y^�V8-�*w��
Ii]�k�v��+�:�C�`KH��T�lx�Y�8�L��ߺu%��>͓���qc�Z3�7GSMr��SE
�D����m��&+��|��v�h�!C�}�f��r�4۲�7-��
�ٶ܁1����|y$��9����us����M�bR�������~�3F��D&͒�b�;�D�����M�U-���""��M�衩����ոN*`��씈z�eU�y�Dw�-Zs`+���b�!�ho�6@��.�h':A�9�b7�1��RAj�Ǥq-����������h���Z��p����t���%����G���U��C��_󃴟O����
��Es��/Y�&�ܮ���^�Й|O���vZ�K�dRr?��gg�R�N�35���J!9�_jI��ϓ4��4��R?�� ���Ӱ�"�i����629&.�.���=���շ1ey���a��Ob�Ɵϐ�w�OE	�� ����.f:��	�Dچ�k	��%W�?�]���E��!�B"ĊJ�=e�$�6vw��A,\��<���G!�:
9��_a��#�̬-��_��v����)�f�����⌳e�������o�h��+��8�^���7�_�#z���d4C���wr/�,EL���_	0�-W�Uf3���Ղj�}��EI�%�D�9��#Q�9�w��o.���ԑ�Y�Z�q�`{��Q;���H�)crw�u/;��F�D�'��[6�+ZŪ���y
p۰t��g�	[�={�me�E�cr2�%��E�q�T��J����[P?��ƛ
{V����1k�M���ߊ!D��F�K�Ӯ�\��?F��E�GC&���:��q�5���娞��W���D�N�B�J���<[L_"O�a�eC�ʉ3.��U��ݨAdG$�.z��aEH���sh�'�X;�#����$a��z���j���{�s'1�3����b4TO���i�]y
�B�����F�*����B�F��9�O֩�fxC럂6X��������)c'��P�'�������-�[�g�q�ީ������o3��}J��q�n��\7���m�<�`����vH�d&�����O�&�۠�g���2�u�n�:O�{�oi�����(���p&�����i*��Y9ϸ��C���mK-�<��-`��e�-�*T�1O��W?y*�#`v���kB�֞��FŚ��ڧf��M^
�~3�UX����*n5��=�=Q4��7m��d����#N���8�Z3��p�)�r8���k�ݩ�LC	�I��	t��5co�5���T$��I$0��0������(*�	���h&��[�
Hmk���	y,=^�0jp�������wף]�ښ|[�R�i	�=����l��U�fǹN~�zŎ��jz��z�٦��]:�UӘRr5
���`5�ѧ}�=E��$�:@,���5&b�TY�Ѿ�MN2����D Ĥ�TP�~8��^U�<�VIq�Be�r��E(���9��M�n��9Vg�褊�z�'������b�)�V��i������X{��(���f]���FBp�%��}�@(�P�V�ew0�&i�S��:�$B��.�@ڹ��p�����	}u�@T0�v�-"6�*��hN:sρ�&����Q֎;��k�7q�#���Y;!0A�cQ���\wa�ݵ.Sh���9|0,Kc�Z�d���s.��#[A���h���N��IwjH�v&9t&y�ʕ�MLQ_�����j�s�M�bVw����H�Y�柎P��q��T�����t��@N�~0�%5 Iy.�=�L�9.�*>�4�Z��Z۽^���S�*/u텟c��g�p��}�r�0MW_mL����qm���7��=�<������s}!/�q�g�B�����J�0�c/�ƫ��A��<A� �,�G'�3M��'f�<�L�v�*�D.;���`6í���5T�P���O5T�{vo�D{ܛ��,,��p՚~N�g�[���x���keZ�lA�S]x��J,S[�0y�T!�b�e= �T��2k7�|��V��;s��3��
T_r
FR�eA��?�w=TA�lUu/]z|�`����	��?$�^��4\K'%Y��d9<�<tr�3
���j̒�Jk�Q!����.�U�?�Ҩ;�)�35��|��O�?�Izk�h��\�Xb+����SD�Š���PEsxJ;�~��8}��#�Ò,2J�T�4W���(0���k���y��
��/�sy����h5;j�Ed�x�xD�G�4�͑�~�TD^�������҅>%G��1q�����=��S薇��K?5
Q�C��aq�{��,�^����<g7�8�6�>'�p��5H�S��0�>�v��u�d�1�SĨ8.�F�KpOX�Kp�}��G�4�jy�n��B+�Ĝ}���'Q,�)�B��S3�77nR���ΖԎ^Ĺq)�ꤊ�l�-=�L��y���,��3�E�+� �@��H��@Jp��$*K�R�t�f��a�so	����jCP��|Χ�0�f\�����N#a��\G��M5��x������w+Q!��"�!hiv�������_B�����h�;�� ��z
�9I��`Ù��8�Ia���}���Ov)�fKOd��)���Hߙ�uJ�`:�2��*�^�j̖�_��������=y]���8u���x�j�}��*9��a$���SY�?P��� ��b�9�mH�ih	6(5���$��]��뽘�;1�7a�P���;� hFl�����PI�o����G�`���xC�MgJ?�x�7�}�`aU9 �
��U��#ݹ���1��吝-ε��E-wʬ�td�pv�V�h��ʀ�B� VH>4�h��]��0;@x����%q0�l�+����iH��Z��&�Uzͦ:��^������͆�4�`!��N���׈f���͞>�!�i^�hq�=�3Z!迹l�]���t&n>����c~+p�wB����y��^�<��@Ғ�[� ѢpK�i)��� Axp�s/�����������'u���Q�2p�%�ꃈ*�AĚ�$��ڍ��A\w��]NJֱLߚ��$m2˂3{���`M��g�H\�j�'�����i���s�t?���Z�_�|�F�Uۡ�+S�-�)-�Pk���? ��1Q�B�H�]�#�Mҕ��R�8��S����/o��%y@�'Z��`~�r▱����e�����[�fy�.I̟]�Fj��Hg�̭D�`��#��t �Q��	z�73�|%X-|�y�C��Y&��)�u	���{dwȏ��כ�����h�
@2+QrD�?�VV����@?�A��䬖�X�~����ڬF�C���81��i@�gI+�O�K����':��=�@%	���9��y󒫃�n3�U�?:+�˗�$C.�$��e���v{�*�0���ٗdL�Jl���c�,�]Z_�,�p�#l.05~�A��5�.h�,�Kƻ�99,]������q��D|+�����N��dշ��e��oX�Z�E�ո���a^�T�0���bڃ�q6!�U'�Y��,�FPq�}�/\��E�����6B�LW����*P��!�'��z�g6�u΅!�M���&�vBk���(�0X¯����K�_���"p���y�R��g)Hw%�dg�h&�3����f׏$8�s�d�$2���:��B��El]n /�z#�����O��3O�t�O�B�9?�_Z�&1s<�R3�ar�W^�6b�������F:1�0+��w���C�X�e%����A�'/9��Wqm.���"��_�(��/P����u0iQ"����~ъ2]s��_��#m�'�/�Q�>�p0
���;Q¿��B�䩘�5o尘-ڐx|AOm_�Ɏ��!�r��p��PSǕ��,j�S&_{F����3{��"���_�=)75��=Z�>v�114%8g;*���χ:no	�lZ��؍��~��'�@���S(�қ�����SO�W4X�<I��8��I�vB�_B�`�%l�9��-,�缆'r�a�O����<|��8�3"��n�~R6�@�)�[$�����&8�1���P&��^�(B2�>]�q�a6@ܙ��Q�2�������4��r��K����\��V�c��m*L�&է����x�,Y�M���G�|���p�|K�ۆߘ�t�� '�P2O����v�ԻA���A�b�����E��$ 
zU{�{��ids�VK;"������3�M�.�_�f�]^1�K*>b��@.�)�g�H���jIC!�Ii�l5b:+d��ȧv�@KyB
�m�+�]�Ƽb-����/��V+�I��Z�N�$_�(��j������I�N����[V���픾����M��P�y�2b]f�uJk��F<�����\��yS��S{�W�ys�Z�kq�b<nE����o@�q�	�J�}�ܤ��[�#J��r��c��[�C��?S��%�'v�M�"��&�%�w�猌n50K|�a	������R����v�EŕI�l'O�Yw$n�B�$C.e��^J��e�
��ϙ�)�󕚝A���G�w�S����O�7�Ց(P*EX�Hd.���"=K�O�u���g�g��`(�M|+�����O����"�A���(�p�5o5��/�0IY_�~�l8��ZS�@'>T�oMp�Z~�M�G�3��~� �]� ��	[]B1<s���Euo���_�:�����.�S�>��!Q����.��j��O��d�DÊyɐ���^C��B�s�_�+�����e���7s�����X2���Ns�J�,O�½R�*>sZ���VY�	 )#}���+u�y���ǾSa�B��4�K~�5�R�H�@����,c����B�mof2�jZ�Q�
y��J`8ߓK;	6<
-��z	��}��0�q�߰���Q��rsvk3����Sii�MN�BMދ8����j��,z���M�>�����`2e�h�*I��!FH��z����)[4��.�ÛiM�@�4t���=�a"�?�����@����%@?{ށkG]v��|+S�F
�l��oj'.1��F������C��ɜW�������М�PY�ˌ��KNE9)k2��Q�P���Σڭt��-Z!��L��˥���a�rc�O�S��W��P>�������[�"E�C\,B	�#�'�@W����+��ࡾ<�?�u��Ϟ� ����g9�Y��S�w��iݍ�:����J�V3��w=���N��o��o8T$1$�B�3��c�F���%����)�jF#��U�FP�D_���Z�4�nG�!��4��	�G8�c~�k�)�Ŕh���e�1��jmn��raV rDE��vbI]o�d�W/�=�3'���?��pi	����֟��:���D��t#��æ��OZi^p�<��y+��U���:�Ct�:x��g�.���#�BF�q3?�Y[���<��ǎn���7�f�\�����^|;V3�}���6�8�뺋���8gY�h���'2�Ɯ�N��ն`���5�Z�ګ�H$���9�fyS��M]��7_�
��U�A�@���n 0�^�&�)DX^YX��~��j��bn�tb�N��Z�'�������QP�_�Rяx'�bHa�u��Ø�O�QzIs���D,p췱$QS�_`��$ן�ǳ�0�o�(���:��F��H��2�S/��;H�lB�z�~aʽ�R�[�+��d�x��v2*O��?��tC3�"��|3�E�ܨH��w/�O���&15�^���0j��瓈�r	��2��D��-�6�82HF��+dK��?�w/]��%�w���R�9��G���߅�u�_P6�25�%�^��v@��;Z1��8����*G�,LK9�R�ҷYM���r9xUe�]�8���,���Q�$��&�A�7���