��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQG�.�����t�������Y����C�ۋej�'���ᄽH�*F�7o�$�N������D$�K�>�J�w
e$9e.o��U�x��ܩ�����k�g|��Z";�l&S�a��r2R�G��,.[l��Х��6����{.좋�%=�W�yW�^KN��xc��G�#��y���GV��C�θ��~5qf���S�u��Bd.���\��
$�F�������|�/a�%d��!�﮺�4��O���~��nTX��uc@�K �P��J���xZ�W�YXq������j׆�Z�Xx����2T�!�K����a���A��&���o����E=)"�)^3B� /חqJ�o_ù����k���D�*S�˃��)������6�f&����x��x�"���&�=p(���$��F�zV2؇��L�!R�n��]��d�
����>���.�]��XB�'�7r�>-� ()�i>C?�Eް� �L^M}`w�?���y�ni'S[�z>͚��B�7$��&��|f3�$�*$7�p�.��d�հW!�'s&�Ǔ�6��b�A9(�����(z,O�5a�2���䉢�{� Tw��<�O�{���>�o햢Sݻ�E���y��h�J�#�)�AZ�F�7l[Xc����%�� �8��U+[��"�V[�{�:����`��v�yf��6�I�uN��!�(��eh/�]L:�`�w���J]̐=�Th�F�tQ�\�ч�J���r�2/vי��gI߇���J����ߑ��u���}�݊ O���R&�����/I����FRFc���W�o}��a
��� "�2�f�@[1��R�o���%9	����??K�;��8�J�����Sʚ,˘;;�����K=K���B��y󊑭�ʕ;b�Z3;DYZ���I��c�G�����j�8_����4�4��6"�閣\���w�}"���|��W����X�I�.]�5�a~"YdK�/In�14�R�ü�<�^�l�4R[G������S%�X��x���E�Xe�1q�@.��s�9:�� ��qs�fˍ�.��D��v� \)|d�?zj��+U�=!�! *g�+�i ��M��K���r���U�	��ӣL�0.Ӳ�Y#�ir�_Q�C��1���c�9���6MSN�L��4���p�>�)A���yy�۪��q�AW#Ժ]A�F ��<j/��!=���V��	�
�JPY�;�O	��s�i��B������Bf��W�8���c�:t�y �m�Q:C"&F�]*�|%��	��c;Q�3P�Eu�Y���n��$��V��6ƫЕ������>d�6���J��.�x܊G��2;&W����434
$}�c��1+�gc�dk7|���2����XP`����񴹢�t��R�\��^���ˊQr\�˰�+�b'q��s�5����al�\dP�#$t%�7� ��� H�-��2�x^tT&A��9E��@-l��f��o��w/T+`l�1�T�6؂��
�����k���N�#��e� ��Z�Z��T�BÃ$>R�H;/��aҝ&��Ƞ�[��f�o��:�Q���&ֈ��CNA��Y�ef�ڈ4���EU��(���H}x���Us ��㑥m��{G��� ���2�߾��G�qHBd�Uk_؀�=#�o��s��7!Ζo��̸�":��߶\��<2C��z`o/m�f�NH>͡4������m�W|�5"�d+b|�٩��X���=�B�-K�S���{�"G|�lS	�E��B 즢y`8����@ ��,�uL@�) ޾�WiU��0��PN*��Kc����FNC��zY�����N�bC;�Ő~�{vZ���j��=G�dQ|�r�Ā���\I[�0�E��yJ?ݥ;N�T5d����G�Y_�H��D�#E.2XT��&�P�OfT��o7f��gׇ��ؔ��@������V���%��N���I�agА�E��!.��%�L����(��mf�9�s�S�
�)����'wO�1JY4��Z�?�V�^MՌ�ͺג��(�$q p?�F J�����^'hE�G�R��A�CqJ��t��h��fz�~��2��)��D�e�+X�ib.�V���a@\�,�2T�јf6��껔`�K~�����[%ો=�pd6�?Gޑ�ۂ_l-���$:��[�d��"��W�"�{7��P �ub��K+u�X��d���#�;qn,�9�*`g���]��ϕ��l	o���3>Qq<QD��z�<��5jQվ�c�~ï�t>�I-���y<?���&����Y���}�%o!�m�?$���xBD ������Z�M����l��NK����8�ݵ�
���=�އ���kũ�YX�P;"ߵp�(u���Iߑ}~���(ES��t����$��L��l��1:�[fq=2��S�St)����KI��oZ�����}��ә2Ђ ;�)~�n�	�;d��� �.gs^d��������l�6���e�@V*��~5\z6F� �uip\�Q\+yR3��=�&�îtG[V���~�0x�����mwE19��5$�ܸ�ut���
6���H������53^��"���B��ݤ� �^
��L�r��ޘǫt�]�&�Nݍ�'ף����X���"��_���*H��8��~Y��εB�4&�4��ݖ*�3�W�A�K���@��w�e	>��Ģ��دF��U��8?MR�>�V�(c�9�
�n��*����m�fR볦��2%4R�6z����H*����;{�줶�fra}���ⅽ�G�Z'��C���0Zz[�3K�`S����|��f8����GOqA@�([�gE�Di}�͚Sz�n�HM!���.�l�.� �O���i�!�z)��8��0�d�}���ݴ��z�a��פy����}��>Z��2�mb�ڙY7���h<f��#�MAk !��o�!���\/MXP��|����9Ά�_&	���w�����X��m{���,
��~�x��Y�0
Y@m��	V��T�)1.je�@���͈pgSf6Y���%�=	�CHm��~>R��^�Zя�����s����a�?M��q�4�&Q��%�o;�m�ԛ��r���e�7Og���V��3oB��䕴#@O5`YMf�%Kh�smʾ�]�3\$J'�)F��+��P1��D�Y~: ��YlK=Bp�ZW��y^�ḯRG)�I���(��7Z��M�O��d;�e,�ކ�4 &{��X�u���&���(�:���(fĶ{����L�/��Y,���hKIW~��T+�cgx�מ�]b�!�짢B�s�	�[2F�;����{&h��T��{󬱯O���wW/kY��GW�j���G�n����sG�E`���u��8ˎ~��ڪ"��Ֆ�K7b� n�a�2�Q�V�'��T7tX�WcM��A�4��G�_Xq�5���zNq�$�����zjJ<y�.��WT�ЅCt � �	+tjGfO��g�y�'�P�n�]��749C��B$���w��k
u�g��_��]笔�����=�K�7�I_p;�@h�@_M.��̠�9ձ������$m:�<�SC��\P�S5n:�K[`��5�h�O�b`���-��-w!����٧/$���L�.���++��b��1}�H߆�=���e;WfJ3�@r�D��-8{��l7��s#����n�w�"�ƿ��c+\R�5CS���
ru	kc (
?��>�ͼ:�/�� �C�c+��E�����n��}Fx5K�JrNT�]r}^�-E��*po�����7|�EP��͘�X��@����WO�L�Gv�[�g9b�T��k��A����Cd�HY��Ղyc�z��U��j���[�o��������lY�>��y0�ޓ\,b��oK�<�q"ޛ�lى������N*��M߶t�ʓ!n0nҺ���^1Һ���(�K2�N,�P����uQ��Ǖ�� �d�dǺXI��V���e�����Al��d�_����ӊ�}��^l��dT���/D���j�6����|CjӠ��"��oT�6j���!��c��/*{�UDM�/	��p�j���j��>g�~1��3�a�B�
A��r������FQX:��1�iձ�+��ڔ��
HwU��ะ���t����^OU-n�(�zW@��q�pX�S�������� Z`�����|�H+�������]7Ne��K�g\��G?�\��%8z���E����fq�Nŷn�+��Θ�i�]<���|�ب�Ňb�Q�s�1������a���
^!sË��؅|p/N�@U�[���Ɗ�� "���U�X_������]SԢ3e�&���l�Rŉ~^��@�`�(,Ę��eJ<e[�T�Gm��?���wC�ewI��oR��]�7w�Ʈp��N�t�P (�7>X�G������b��,��<�r���`
Y�u�Ӂ*B���c0��H�f���	f4�YS�Й�5�T;쪺.X�ӷv-<2�{C�8����s����JZ�����Ökr�'�"V4[�@�V���^0
ȩ 8����"�[R^7�0H�uڽߦ?
�����M��`b��y�O��NT�+
s�o�t�Dc�\r��w5��1E��x�s�R����Ep�����i���<�)#�ۖ��e��Lo�-���:����*l����� ��	�w���Vb��%ሤ���";��-"/K�.�8VK�_~�a0�_����kp��G<f'��U	��}�Ġ�	?�A��\��2Js6D�#�I�������a���:���s�>����Ԡ�tk��?J<�`��,^�,�����i��\���0�M O5���e�/W9�b�]����r%aB���fq�.6D�wה#:�����g�'�v�pa��ڊf?ݕQ�r���A�5k�/���O.��#j��Ox���I���z�sd��ƹ�~&Z�����+&w;�&�u��*�$y��J�}��RO����|W~I��٢�0��u̖YJ���D0�_T׽�0�ax��d�ߠF�3���w��v�];���<����U��0ǲ�f����Ty3�aB0"|U>���YF�x )ya�ҧ��^�B�d4��B��L�@o����ߘ�!u�nU_T���րc9C�^k�ȅ�ߠ�	Q�5jKy�MF��C/�(%`���o��=�q���)ː:��Cxh��OR蓢�%�v�?�����%�vf�+RO#;s��6��嗂FIЬi�Gso1-�
����ŕB�u~�Bx[�&�����$���EA�cڢ�{K=&ML.0�	� ��,��+Z5��-UU#%jy��F���'a{!�ōq��u�)z0M���7��Р��j(�����D��b\��Z-�p^�� B~��h��5͞���h�>85$�p��;8 ^����fƮ��M�5��0�B�G�b����ԍ�}����_���S#w8p�q1Y����Q����L��0O.KW�K���DK}���#1���0�����>As���#���uD���:4Ƭ;����h,����sW�o��d���P�}�4����c&]��R^���Ui�|���w��ݢb:#2Eǯt�,j0��~C�O1%�	I/G����emfc#�#Vǻ�wM]�J�I�"i��d���@���t#�3���IOc(�:Q�ɿ�F.\�"g10-������/��؅ sA��X��ʳU�N�M�5���y��Ϗ/����
d@�f}�bt2t�Po��\K�\Ӯz4��j*�!�N�b٦H��cEq��X��{4S�x1?5�3e�6
v�'���!�dC��J��ޜ�j�n0�I�I���C(���]!�*��N�᭼Q�x0+O_�2�<�@�D�m�&BбG�ٕ��k�،�/����8_�.r���%\�ew#Djr�l�>�N\Q��ޜ2���Y������_����	����Ƚ���H�W��3�t�~�j�2!�/o���5%�!�A���',-,( ���Җ�c��P<���-��e�{�'1�<��ȷ-
O#�0���7�n��@���~}���!�M��I�[�`_B���]H�D"}�YZ�e30��YV��`�0�p�i������<xC���OL5�Ss�9K�E.Y
��-��zs��Z���~�'ꯩ/q��7U� v�Q��2:khR��c���_�okU������˞��9��=ǀ���8�C�߅eDV�7�oa�5�`E@ÿ)��������a��h����3����K���iԮO�b�A�ӂ��we�h�x|_$�0:���Oy��(�,5V�/�]�E�Ad��E�K:�:g�2�}��br-/վ�ߎ��[Ta ��=H[�1|�H��{�ɑl�r�y��_��wŮnYL�0����ŵ<#/�$���b,K�u�P'�/�D"/W�p����