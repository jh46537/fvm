��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���_���W=1����o �6!�z�O�]E���	Rߗ>���B�e�S�w�m��^UA���0��J���{E���*#'"��x-L4���U�� �
H�"ZC���Ez3S�ē��s���Q�^�Sš���P6�X�~���'<Z���#O$6>2�S$�6��<͸���2
G.�Ja9���bd�J�,�@��σ��q�>��}
���Y�4�	��]I�\K����6î7���h Q��ue��?��|��������0hc@$F�с9iX䠴p��hQ���3/ UO<j婙��ā�?�����#^�?�����_EX$Y,W%��-��8�O׊��`zxw�P^d�\8�����#R�77l�i�doN��qve;N��̋ �T���l$�J�G�hW �D?�
��:�3���Ϩ��[�P�@��O�V��.~�t@�+u�����黫�n�8�uV�>6���+�
�� w����c���\�C�����t�"�A*���V��>T�>�ϐ���Ѯ��ȥ��-I��%��ӥD�[���<@)����[&��*������,�K�n�9�~�[ϯ��6�aɜ2@
��H���m�Q%����J�u���2-PE�0?vrxB�7�QP���d:�:�m(7MR&���bw\f�v2rƦ]���o�r�!�|�ڢ�&�s���ǟ�v�'aP>6�D���\�)�<$��Z_�X��a�Q��6��W@�д?È�!�3�Ji���������Ͻ�N�gN�RV�@�Om@�4-��C���5_���.�Ȇ���2�� PـX�i�^����_e 〿6^MwK�����3w@]o\���A�:���(Zwܐ[��]$�?����z� U9J�D֨w�]l����&3�OJ��C�S
c2�"ha� I�3[�����,�j,�-�Z��"��m�eY�E$>���F�}�����ݕ9���J���� c��cR��~�1����7n^�q)�P�)�R0�/Y(��򆓼���o���jT{|����|�cE��&�c��t��Sٟ"]�-	�߿�����UR�7/a�[�VmX3Je_��r�ڳcdΎ������J�.0>���`#�Y*�|�� ��Ŭ�1��� ���;i�����]�2��q6���>�b�*�*�������<3ؗ=X77��8�J������B7�a� �Vɠd�J�_`�ȧ^�>0o!.�@����J��dc��|�cI��e��l����N\�����AC$٦J!���69_��B|0�u/��W�⧯OX+�L�g&̗�v�(E�x~W�@Rе����]2����<,���I�Y�@�SK���7��w���F�(�{nN�%��?����XK*1��#�m�׶ƹ��E9��2(�a,a�X��~$\�
�%��7�r�8�+97~�B��3ҝ��+(:�[ż�nD?i՝r5�/�H�𽻼*!�0�f��>�GR3�ߨ`�����n��f�� Ij�ǰZ)���;���/N��Ž0��i�niB#B%���Ԫ��~X�b���G�FC*(  D���Y�z^�i�Ǿ1�xQ$Ï��1D7S��}N�
́쓃c'.d�CƠ�ZH��]&�C �����:Cgq�aL�E��\��V���ݓ� ���p˙f��4��I�����;����#3�>xȒNκf$,�n�T^�S�YoH_�渘)q�T��W�țl>m~���G�
kK�E�`��n�껔ߥ�N�* wůO���n'מqa��!՞�S�{�d�!��E-���O!6��cg��6Y��)��sF���u,�5��q��}��=�3�)�����{�*'��[�����e�>�L�VRģ�gx�T`]{]#�`5x��R���QD���4B�O*�� �~(�ls�.�k��cic\�	��iү�wY��>.(A�|;�d�`�P=K- ��)4�O��h$����!	p�:�=3?�O7��j�K	l5/��eb�|�ƬT@ī��0�u��k�<���nD9V��m�h�f������B+1���(��f��=A����N�aAW��+(���8��g�"ؒ`��O�~_�sWdo�~�=�[2�/��g��Bam �=!W��U,7B��4����_^М�7�K�mt�fQd��=�(O��-�VH4=�.GA��u���-l��1&��c6�* 5Ų�3�Ԓ��<���o4���?�o�H�&�Dbp1y�[ێ�(��g���.@$؞cI��V�0���21���-�����^(95�1ţ�_Ѽ������:r��̿n�Ҁ��z�u���ϋ�h[>A���))��#ζ$}GMEH���"���ǒ� ���	m��u� Y��
a���K�e�����<d������^$5��.���ċ?Jb��CP'�Э�95В�W��Yԃ}-��b4�I�s�>'�IG��?��+�+�%�ϵ��[o��S�u4��V�	٫w�ƪ�x�Q~Qp���P��Mz|*Y�u!>[oGsPA�4��hu��	�*_g�x��i�N����A��͟�F������Y��e��&������X������bMâ�3-��ʮ��F����ᮇ��>e��uO��D�c�h_���>g�)I'z�Q�P��U_9��Gvx�(C>�����eYqA3���ߨ�V3 ��V����]�J����/���S�b<,栗���:q?��a����6���p���L���˛^ �T6r�琐��[�j��K���5�� ��m�K\����ɼ����ꟊ&���
oy-!��wm?�Qg�f{)�G�?��]O�����h���h{@�n��+��'*:�/�𕥯p|V��`�[w�]L+�;��ja��eD"S�P�s:C���m�Z[����7(�C�k�����@M
�_tS!�@h�V���<�`p�?��Q�\U��f��RD�_=]5*'d`8'���y~*��-to2>�!��)
DmQs>8Z���M�|�9���<���h.7�{���4,$� $�����\�m!?X��=��@},���f�=�s7�W��(��D�7�`��L��Ѹ��D1�$O��ㄫ~��P���#�Խr��@����/
�4e�8 ����פ̢��1j�Ӭ�/X[�?$G"l ��o�1�������>�Ͱ���8w�F���X�D�C!fK��^���ikkQ�P	��N#]��3�&��P����������.��B?�K���`�����v�F00i3����ܡe�x�-��c��b��{!3o�gN��xv9�d|�(�� �A�xOˢ�2g���P�R1�kN?��^�m�_�IS+�t8�s�4(Z�?xݲ}A`�+��x0$x¤�k�6D�oW*ێ�bp�Y]J! <���ů��]a3�����dQ��-L��Lͤ`���9-oI���৵�P�=a�h`�Y�����)���T$�;Uu�T��O���o�����</m� ���=�zxob�9qN�%�H57�i�w-�+{�7(�2t�u��H��<�ס6%���G�̉/�󝺥�����v]q��)�fU#��Hu��@���7"��nq��|M�l�;+܉O���>�(Vh��XW�c�]2������/	�ȇ��zE@���p����/<�	o5������������4���b�����A�Es��[�����I���\�P�w�q�����Kpcm�W�)6�eY�}x�k�����������)�p	]a��z�D�H\��Kw��Q��SW:Q�2\0!*�[�$ϟ��=��U�kی��S�nr��L{Z7i�/5���ɰ:�ƃ{��?2�l��K]������ٰ�����M���+�;s��x��ur�B���������]��<]n'~f�n�.�9i��F'M9���ꂲ����)�׵%yc�o��T1rqaI9��9��ٿ���}R9��M8�DUD��vMR����Ba<2�I��۔��8���Q���3��/7�Ej̘���A�C�]�!z��xo_HE���F�����AnzЎgA�	�hnC��AB����Gk�<�L�C7�aYE`Kkp�O�b捐��
��UH��G��E�́���rw�o>�.{���p^ˆ�mTf��J�PA�W�I�S�:3ݳ���t쁺b��9#��<ah��4�Ѵ�>c�邧�q6V��/pǌy������\j�}~�ĿAlz�u�b��J�����e�!�=U��$%����xe
p2Fy���#
H�e(N�mD�Ֆ�`cYi�QP�c��A��Cs��YU���#��4)jX;�xUp�>��@ae���]gܓn�5Ae������o2Y�v&ǲ�f9�[~�.`r�n����{���8 9o���]������p2V��Y�W?� ��1�Y"�֟�5;�D^Y���4(	P�}��E�m{4���f�,�	fqӮr"v����
_����=If����w�&��H���v�$�\���+{uH}UT1�͊ 0`�GWx���Ŷ8&��dǯ�S�V�hU`�z&��T)\޹m��<?�����}3C���Q�&*P�%<^��u�A`�p�v�V�l����%������',
�6u�YpE"DTG�r���c�rc;����x�CUH�M4��Y=�D3����[l����e^���za�G��긹�x|՛r@ƆW!L�ߥ�'ۺ��B�;_`D�ag6��:�o�:C�Ҕ�c|���ɘ�@��u9& :3a���0[c�[��%SW���j���ه��u$��h�pl���܉�Ӆ����^������s���6���̢����&�z
�͚ 
��`�)�#|!���QC��������b��r�#XɎ3��2�r�c&�<�r�Ӳ����M��0�we&�AX6�?kVJ��P;"<<3~)�ԩ��ǴMN���ה�/u$���L:q�5��X�I��gIKh�S0P����*o&�}팹i7m�:na��ϫf<���A�q���pX�;��YP��[�����'r��/3��;�"#w:AC��7�WeAg���}�ʄw���L|x�zK�@��H������g.dڿ�d�����;��<1G`�X�8I~��e�JQ�mD�������A0�� ������sPt�0k=�Y�-2Α�N�uct^��?5h��xp��&�N;[���%��=e
���6��Dp��(������Bm}�4H>aI
l)����l�0<�*���H���t��b�K��BCp�������ڏ y���7�K��0(�_`9�`Q�����E��k%����v;�0�A�>���e��-��:KXt}�; +^�w�wT>l~-?PN�aoe���)*y��¢S��LX�S«p�����iX�g$S_�� $���yc����\5������b�u"�����y�>�X�{�{�݆Q��#i�8�P(��b����!G������N�W�VR�5RO��7Ƥ��쮧�!f�Y�0u>[S?��c�fr�4�ح,Ö[^H��ڎ��3�d!�|���Wm0Ak�K��
�,��+��E��5�ܝ���� �{���&���m]\����� B< u)��8;e�k�,N�c�Xk����Vy���L:V�5���zw���X�$���M�܄��P#�X^tݮzKs�	aV�\�rm+��]�ZXEj�]�� 1�zfq�@}疢�Scs��'=� ����E�����S�).ê�1�]=U�rB]�nN'rxx�
FO="���h�^ǅ2�jx����**��
;y6Ќ�o���=��{�S5@��JŇVM�4������y�Q�)EGx���
Oц�*�ط �wJ���TUHu� |2�'�!P�.{T��r�4��R͍���N���u��2ڜ��6����/+��s¥FB*D��������B�~�Bg��S����a����Ac��=��O�YSe~��{�s*	-x��ō4o��j� %®nAV!�$o��0�f�V���
~��1�z�m���f(�^Јev���q���\9��vI�x㍗Y�Z�'�gQ>J3M����-�A�<��R�l2���c�I�o��א�TrUd�rN\;��Eu���=@0$��_���s��~�dn?B.c��ODϻ���N6�W��!��O^�@�@k>�aGM��m:�Cx�N��QZ&��7-��/���5#e8Hp�l��#��o��$v�fa��G%�sD>�G*r�3�2���7�Qʤ[Do����`#�G5z����ԕ�|| pR:���\@� �)�#ۘ-{��5�7E����|��\Y��0�[��Q?.���PKV�u^5O%J
����������i�Y<!�Ds�V����2 =ٴ�ڱ?�M�Ձ؄滇!����M:���㬭�Pn��}�E���?���:�\9|;�mN��x3�G���F\��Ka�N�{�P��j� �ڄ��f��q�aah�m1h�\V�+�y!]
����*��4�ߥ;Ye�����ۘ#�U$R�����	�h`(�&f��mTL�k���`��Ǳ�a���!6�	��=���}�1�W�~oݾr���M�X��G�p}�$���|�ަ�iݽ
�����D�Yj�5��k)�ANoZK���Ŗ�E�p���UU�n��,`2'������<8 �{����ͩa�/�2�.��	���:�OZ�����QU��ah�2.��.G��"Z�H9���x ��p�z6q��-ˏ��C�\�M��8�϶�(�Ã���lX�g�p��2� +}�q��ˉ�����o�L8��!�0����G��=_/v��to<Yn�{4�6�!m�X�#��m�7]�K��F
Y�����#�0T���l�e��hyNat��&�!s��_��E�C~�9D�����d�)LM*~SHf���d��N���PJ1�_Fw~0���h���8An/*�Dp���$D��v�2������,���4�!O�)i�I���T�����^.n��kT ����p�L���n��b�kR��D��̈́��p�5Ӏ�S�wL��h��m��-X����K��;?}��ݨ5q��83�j�͞B%�G�2d�N~U�Z=�`z'g�\Bm�8V��k��!g{�DO����ܥrU
Ne�]o;P`�D�������8B<�b2�0ϱ!��A#�L�]D&�����>�՜�����=��P� �%Gh�]�����]53�V:(% 7KL�d֝#�O�G�+ g[�Y/�u���4.��=�J�'bk0���xv��=�n��Eҟ�����b�s'��3oH6�� ��S��1��LCiG_�V���4��f���Mqe�``�\p�{��[T�<]�Á�Yr�D4I�����@I���I���M��M�,@˘�l�W��e����(l���
�mĥ�-���+���>;v�i���x	n��Ȣ#1e�M]lX�z�^����'c[؇���y���+��b����_7�P�6oz��*`�zSh�n�/Se<�
���ՠG���	K*g�eݮ������k*��!ּ]�"u��Zn�h����YX�w���1��ަ9  �S.���ωe�Uby9��
�G�{�{P���t̥��ӊ�;])7/�({���0��<��}��� p"�M��;3N�~Ɯ�X��AbKe���]s?{���nyv @\��Y��ո���D�)eat汔8�8Y����I(���_����m.�*�!�_�Ԭ���p��'Y����a�r1L�9�{���:��X�I(+Q�٦$��D��wЪs,}�I O+T�a�=��Y�ܭ�%yGK�����|��"��-����$�c�]2w�x#��:/@�#�!���rG�.�)�־o����=�d���/����y3���h��Y�~e ��j}.�+j�p��*���0%8����IH{�$of�Kqlj�\qf�ƭE"4��v	ᕃOE�-ݞ*Z\�e��4a[eU�Z�Ve7����_$K��7.���Ӭ)����7�d/Ң=�^��&�!㌦=LcBD�P�!���C`���,#�A�n�~n�6q{�ȷ=W?pox��6�ClJ�wA7���$�q|�0`��yRR�Y��
$$��G��u�[���z]���w'ZB�$�X�^�oJ�`�aE�\O(�u�M�+�81-W��Ua\��:�Gꐚs��~�NUԢ��-b�ŖjQ�����ea��Ѱ�L�n#���=uG鶇DhF-���ս��'�����x�LR�+��0f&��2C��;`7�a�2��H�(�����|�R��������Ie�0�4ȋ������c����Bf�k�	�G�ʀ�X�j��s���D<uE���������W����=��
��V:2����P��B����9F �!�k�����nR/�����<�Γ�`��;[�[��la�ƴZR�I8'��}�&�+�� �|'%NUّ��؀����(���r��4�3�?Cnv���K2hy�������� ���N?���]^�5=����X�O��%ښ���C6mQ�Lvl�)O��9��d�[�͇��H�ו,�p F�#��U�&-Y���3���Ѽ0
w�����?Fi`�F���~���6NE�ݒ�C:G}m�����Z	d �����߱l�Ԧ�l�����a�nL68&���{�cl���{��e�z87�w�_+�6�k�GHEXo���WxUMWP�6�܈�c�8��^�i8,��w{���ݮ�̀9���LO���g|=���=$�$p��#���D){�-_�)�d��dI�͟���/�\�gR9�,���F:Sݎ�%� �Y��^W	��~_i�	���V��B�3U=L&k����qґ�Bv�$��H�Io�j�K4#�!�����(M�O�jAӅ������*p�iUۊ�H�ι�o����d��e��h��9dC��������QK�L�"�7����~~��d=H��!����Eߧ�֨���Z�A���i���*�ͅ�xd��Ezw��L�4Y�.�uc+�4_�A�%����[��F�t�nS��<s�߲#ʠ�D���JO	{>���Y}�#�ؖ���s��
�Ǉ`�N�͝�,A��-	i�P|���������e��Tw��ap�߆���q���O^&Z����E���S�Dg��b�N)|���5�%�Xp@�'�ֆqa} ���$����'{
����,O�'K㶘�=�R�Ⱦ����P�G��U��*��oh�H�������&gC�s��ώ������W���6A���[J齰���eQ]�DR�)�y�F�+i3� ����h��ă .�C��R�@�t����P�"�d�%vg;�|�f���TM�!�φ'��_.r��BZ���SG7�A}�Yyu�����b��K���]w=������E�������#uwΪ����Ѽ�93�]�"�����5�u�e�t�������8�Z+	���U�1�Z�чn�|��$=8��y̆|�t>#��l៾�� s�W��r{��������"<é�1���:abm�:4���~6��[ȋ���FĎ��ؗ���������R[�?���b�-"T�d�f�s}������7�jxs6n��';Zsj���ae���S=�Ԃ&]���p�E({��X�*��X��K.���lk�j^��r�P"?�U�� ]c��$"��ʎ6�nm�GN8