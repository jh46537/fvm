��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�������s�h�qQ Ҵ�pp%�bs�!F1���|W��ٍi�\��չˇ���7Ge�+��9�*m@Mm��A��/f��XT��݌��GP�s��Ɔ4)c��f6�}jwS�����r��j����Īf�t�8J�gmdD����I��h9EWC0^����T�
�we�g 7H�����2�^/����t��PY��Ivs�b�q@>y�%K�~���*0p�w������
��w��{R�8u-C���_f(ZG��|���/zg��P�sIY+�e���<8%���⌚��8gn*rp,����_{���W���J��fM����D�~ۂx�Q|�hCުŶ�_����[�����������=�՞����6�����o��B�#A�����4��5s�32.�^�`�!c菂Q�h�;�wטvm���Jy�#�d�d��_ǫ&؁�	_�dYй"�����61Eg�;�a�F��)�mw������<�l9��₁7�3��� t0�
�u͟�*������q�J����?�$����~��H�	~5>�+D�q��F�*�&��'�4W)��^̀O	�cN/s��χ��4����M�L��Sƀ��= �_����{cG��^ca�n�"/�l����ڵ�h�Q��a�'�*�៰��E%��F)�&�f����ې
��{��m&4�D>uG�iT����^�e����n	��lWD�B��Hk6����_��-�O����`�ݒ��\ZZ���P�+
a���:y������Y��*d�#u����2��b���7��`'t�f]Z�j� 3�����×��	dx��]\���Qw���<� /l���t�ǍS��:��aM���Jx�s>A�`TZ����e�We���xY	��K25�� ekC{��[h)=���L3�ҵu1&�CR���U��]O's�6Y.�84�`^� :l�J���.�shj��K��z�=�eb`�ߧ+��@"��B�
�5��,~�W1� S���
=�}��V:��[�'��/j��h�� +�"�.��Ƞ�X�d�tCιV]��>�Yw�ZV��b)�Q	Ĵg����C/�]o�'*ڰj�D�^����N���T"���7h4��ɥ����$=+��)T�/�e�@j/7�O�;�vQ�x�:�Š��\� ހ<8B,�[����l�#�a}���b�h֚qJ�@I�A6� )/6&���+ٍF�9d��e��^�v*o������	����J���Yx��tT��T�&Dмa����[�Y�/!溬h�'�ڑf���2|l��?w�Ág#�m�(��k-g������?���[�?nQ�����/v=�/8nh�XXxq��>���9��8k�B�@G��� 2�T�����Ӛ���S��F$c�[��)}�=��8i�m�V����?/�oFތi�"AD�7��+��./�(@�o.�d���y��@P�����=����R�y���n	�	(+I|�%$�
%�J],��E�E5h��x!���]�:f����ZqT�8Ne�G;�W[��H���3��e���ЭP�G�����q:�J=@�Cv�k����=�G�k
����sl|S������������!�Cj�f^�ɺ�hO7��Al��6�!WF�~)h��_+�J����a9�7���Y��F��@����K�3���"��������n~C�ѝ���߂����Mc�_�볘�_#OX�d���0)�h�E�p�@ᥒTa�*�R�ݲ����>V���$Ԇ�-�d~N�'��Y��$5�yMt��.fQ�ĉ �*M�/�eZQ�+�pϼu��鈴8�<��"��Z����D����gqw�(�l ^^)MC�-l*���>ʇ%� I�HV�h�d��#�|kQJ�+@��h@H���}��VS���}ͣMb0�(��D�u����Ԛ��gN�O2�^2�[챙�Z=R��J =j`)8�h�)~���%��mQi�� ��*�k||�)r��s�4�ڢ'y��Q,�yr'X��z��C]P�h�U�#]��$Bj�Qi*uQ���];�4
,�͑�+�Ù�5;Z�ۤ  �S<)̍w"��2�R��!�2#�3C0|"\)�ҙ�X���	�cf��␟�o�0�&��dndL�dގ�᧲Q�}�VI芫z&(���$�V�ùɷ���@���� E2:�3�li��YxQM> �O�%S�E�J��3����6s�8��rh��ڌ�gK�ZR��缗��) �@��<^E�\�X�|�FT�P��E��Ԧ!4������1��W]�!FN�z	
�&�[i*�S�h@��1�*ǔωcB�9�ȥЉ�w]��	&p��L,�k ���L�}6�<)m���¯�y�,���������ɝ|��dӠ���d"��Y�O���U7a9�!�v�c�
����.��'�~j�f�t������Jp��������t� ���bc���V��\�F��^kSW��%��kӏ�%iG |���U���"�8�S��������c���pc�j�zb�ZE ]�����#pK%����:w��	��ɐӊ�̂O���ƾ�R	�~�J�S���M��f��ύJ8 ��*z��을��]JJ'���)�V��p�|,��WRU+�ec�#f����������`}���zP��� }M��H�R�M�8�U���o�3P����P�.=�|�(�Up�uyX6�|W?\���ݣ[���7��ZtmW6�A~�̚���ɏ"tB�*�-~�id�RN����l�O�gB�)��5���u����p�OjY����K��e(�ɈB�^�\7���+�A���U����\5�#�Έ�*6.iC��hJ� i�7�f��ᖩ&)ζ�Ϸ�-^�5��8���/��0xW��A��|/���*�lG��!g�d�!Գ<w�ed���a������;�x0�%IT�C��،�)�+�"��).��](��Q�[oeװ����"�Q���9��	Y��WE���{�pQ,DFA�ڳ��|`nٛce�N�&���h��~����Ib����%�"*.�!��ql�Gv�De+�:d768�\�R�R?�E�X!rR�t��C=�I���+}�}��V/܌H݈�����cj˱��Q����-áG#(OR��F�&�<o�Kl�YNs��Iv��ޫ����&I2[�Ւ�������O`:��yu���(g���j�ߍ�����j��i�]n����j��½V��G�O�p�%U2����t(������*RE�tg�,����b'�m� �YBX�K�06�V:�(/�y��k��G����K��f����t��Ⱦ�Sl]�̮�ێ�X+�!�w�w�A����!3h+`��2�f��_%�5���(���a�sD���	!����G�]��`o�y�"!y�QB��q������T<Z��j�H}��������3��ǵw��a�Kw>8͚��y`B�ʰ�h\-�o8x9jr�I�j^����12����_�r9��F|�҈�w^W�p�5$�u�uxmGT����ϡa��Xi/c���3�;��ZK�PW�����}�#MV��iL�����6)}�(��+Q	!�4�ͯ�F��烼�J���:�JH��f��Q����>�$+`;'\f5�˰����SĄ�U�tH�n�P����6n�k���V* ���T�Nx��U�~w�R�Ѷ3�m�~�g!���k-�/h,�g�����4%ȯE�r3Y��dt��/���a@�6�|��ț�\3�;m�v͍T���� ����_��g�ʥ�� �KE*�E����U� Q�u���Rn�}4��e�q/���1��6`w5�r����h���/��(c�Ҳ�h=}�WA����i
�(��\1��Ŕ�L�)�f�+5��"��9�{/���<+���=o�؁;(.��@L�� �Fb�[�a�4� �r@7	$rE[gq�ev��*�����BE�N���\q��/T!%+5���׳����]�H�G!�.ďY��ض���G��-���-~$r������e�r�#H��/G���yّ��âF}?y�@��
���}���H�|���?s��Ys5a߻<o����E˂�xFC��҈ub����3��oX.:<����#��]����	��\��m?��M�P�PkK����֋u�
V��::ӪL���0����'k�^I����g~]\��kQWf�O�c)[1(�]n�R��5��H4n��>(&~ԗ��p�װ�ek?T�;�6�UvV�'&��I)U�S�F���FZc�$f�q7���m�U��
@o��ҿ��ݕ&\���9�������3�Tl3c���'�9��h>t���]�mu�������k� >��B�W��fR[]������}{/~��\`e\�9�@��}��S���˂۸�tW֥.l�����L]�yW�ɿ�S�V%��K�+!�����,����@	��<����W_�M����߀>w5�fm�A�Wg�c�l�$�k�#�0��̘�BI�/�ޮ�`��P{.�sd�?�q��}X�7�T%]��S�u��_�`�`ͱxY�j�kAt��qnK��-}Q�����"C=ׁ+1���ʲ�C1Gx �e/&p1��V|ey�����Mo�c�U���sW5�Z���,�+Y��i�ڙ��y:�����zN��7h�L�[L����^�8�?��z�"����u��JڙZ{���=����/�;6\nE�yv��aEܐݒ�n���s�t�TT�h��;1�<�����^7!1>H���^�L]�'S"$Ԍbn��l���gt������?S�>q�������]�'$�6ֵl�i�hϔ�Y�x�$ث����k��!�SJ�ױrt��D���=��[�t6��N:����@R�hB)>����y�� ʴ��pszs����K
Ak�V!��Ro�kEA�t4�5d{Lq@�֒T�ȝ��>6o|�-�aH��Z�dT����9,ڙ�K�٧�r��{S�ZY���~R��+?Ʈ��
@�H�!�Mkd��j�D�~�o���$u����Oȡ}�Ee��}��Qܙ	x��>i��y�����^!uN�f?&c������� �
T����	c���Z�|�(�0����e&��zξQ/�*�W�Eq7JӋ�R�V}�	G~D?|xK�\$�����-�VcC��P��(}����BW��J�/�Sg��;1( 1���ՑZׂpP���%#/�㏸��f�����Qw��<~��E�(��kDΨ�� �I�qA=�9R��֟��%�t�#��ý�},q�'�z�ͽ�T/��0)�`
��Y?۸Ѥ"RB��㟒�^���,Ξ�5W��(Qz����1�>N�~qH��Ώ�]m�%+��
56��#?kXf'%��5&���r��9F 2j��0��--6�*(6���4{ n<R�����L�O �t���ȿ�0FB�g�m@��r��:�6o^�d�Xs�
�̏J�>��
��������� ��;��ez̒����� Y'y z��U���e�%WI���D�@u�y�X��p������Ꜫ�k�L9��Ɠu��Z����a i�6 �*��"��g�L�{"C��Cj�&/F9}ua���q�-�l"R�{�塚��:�!�?F�
- �:\P�.���M��V���\E��9�}"=ZX�|��������@��&��:��EY�آ�� ���'z��eN��:�z��lƳr!�3�g�o8#���g��s�χ��Ю=m��N�s��V��dJb'���8zջ�%^��N���J��+{x~�����TY��d�w)e78��ߚ�b�'pG�7��Z���C�-΂)�p��R8�9��ɟ��C�3�/���6�$ݨx"��W)旿����I�DO+���:'�l��햻~8t�]���;���@�}����/�0G����7�*��0rO��Q�6�Ұbi�d�w ���Z�����dO�U4@�$o�:������K�!�� }a
*Ȯ�;6������ ɸ7���p�<񫚖t����|
��Gr��s���F<#����:�%K�1��>�c]!B�Nn��cf���������"�ɪa$��Dפ�������:M����=���P�j,�:ʄ2������D�;�6����B���w�u���@���5X��~�����������
��a��0n���Iʓ,�㟼�4nlP����DӔ��~��W���|*�H� �I���~^��muU�$���[g�����&9��0�A�Ӵ��V� ��1���	1�/Ƹ�I?F�,{5�����+\^�*����E8�������!8Iw�,Pp��-�H��Vl�d�s�upR���6Rώ�(ڗe&����Q���X�{-��9�W�hY���i�&�?�'�vS��l�#����}�yq����b�_f��xu�n���f��Z5�����#��~13$k;��s���f�d�Kٗ���U6�g)�5tQt��O&z����F0�\V
����������-�cm���f�����A#��	��.�쫹v��ԟ�Y��~�4NL kb��@M�76p�����Ƃ� &�ko~�t��څ�Sd��V��TERM^�4�#'�\<!���/���H-���^gq��W�����(�n�E��(c�ΐ!��xi�z� >����+�%��n�'��[�:T���6��=�nS	�wg��%�j<$G�ƣ@��B$��?L��_�/��.��/'�υp�Pī��l,_�$k��'<�"�l}���"cU�i�O��Z�'�$��߆Ƿ�p�	���ջb��h6�F�(�O(/��v)�Ȕ	˦M2��@����D��\�����!���Nw�V`ƺ�7���=ؒR�J�L�y L��J�bʗ`��OVyv0�ps۽.d����6&�g~�*��_����=���UZ����+�n�$���%�U��ߒ��&C����r3�q��t��`7��yO;X{��W��yC��2e��f�\�ID�|ll����M�5S���x������E��;/π��N���QR�$���y ��2����؞�)����M�姠`D�9�X��K����;��T֛�m�����4
�j@�O)"��mj6Tµ��ߩ&s��ud��R������;2���+��"W�Y�&����[zs�TX��������Ju%m��:��4�A����� X��MA�&B���5��3	�����lC�~��ZnS &�P��2hH�S��5b�Dh��qԈ�>$�1ZD7U\�U�����)�+�F����0��vo��ʟ�C"�4os��6C���ю����솕��L$�Q�8�A@�L���e�j��b��<��g�C2�t0�&�l��k0��]��Y� n�#�aB�7ծS��L.`>_�Cr'�\�XBDw�6��r%��4�+�aDT�o�3p'��O蘣���6�� GԿ��P2�Zޢ��U�wg�|��jX8L펳h����&Y�q\���<Ht��<�0���������KquĪ�n��(j�x�*9�tWs]<���n�j�wJ��#{i�87xV�n�w�WD��1z����ۧ�}u~0PS�b�]`��ۯɂ��z�jg�}��2:���[��S	S����v�`(����1 dB
�T����'�5�n�mO�\e�60��5��
�8�g���S�&lO���`\��f�Vc*�;�E2�]o=X>�l��f=>�
=�*��ۂ��X����,o��狷��gH0%:g0��/���m:���tПBI].=_XF�{�p:ѯ�X��!{�!�PҞ�5�<
�G�a���tRj?��o���QX�@�F�����W���p�=�(����t{1�Fgν�+,�'ђͺ�-�t���YrMi��0R]��Ll���ڸ�K	�LΑH�w-����+=�[8��Ͼ,�)��O�nnd���[��"H̡C	��F���W1fYB�a�+NM$��P��&@2����{�-���K��^p��_��.�X6��sd���%\W<>�H��rȱ��$���=g.D�,N^/桥�'�W��k{(�~����hv��� >�j��x���(N�_`����<U0���d�?%��<K8K	�09�s��CT
��`F\�S���d����tS���wg݉=���KW�D_�9J�̳s<s�MSEY��!�����~�H� C�3��c��� ��[AܢFfװ$KSrE��yN�Y�rx����%������NY�1*fye�%)�y}��\`��	Rb�q9��ކ�s��{$d���
�d�3����s�b�z4o��I��?-�ts8���a�rW�AY��c}���,"�{�G1+�a���� ����l*�7���	��C�.j�>цh�WcM�
M���lHaф�[a��]~��l���SI�r.��7h���	�K7�`���d��*v��/-�t6�+9yr�y,�6�х*�y�hFbʏ��#�'7!�kaF��Ս�����(���is�㏃�B ��<�=]�39�c�`-!��5�&�}�̔3(���i���{������ź20�4���ϼ���Ww�0��/�]������*ٮb�	qe�0W�c��~�3�m,x������c��������w�@y�1.�|6Ѱ���������-k\t���ot�2�s6��\' �w��k:�l�)�/���.���J��!�-;!�`8�p寮U�ڞ8�J��J��]{�-�ܫ\>��xx�����3~�=9�@�k������c(j3�-W��#��,I�T�b[��P��r�X�H�N�a��H���<����	��;�g����5R��o���R��g��8�� LUI����4���o2G�<�.GTViT�"�9*�&e+�Az����:����� =8y�Ɠ8�����U�՛� ^Ge��E�U»�ঽ�u���w���8�@��6x�ks��C��A2A~��������wh�.:5������5!X�W�L6� R2؞�&\�Za�������}���b��C"��?��`y#�Iۓ|:��[ �n����Z�����!l"a8�.����_��L]AP���D�=ﴝSg���#�0ei�8��R��M��/�X�t3�!d�����Ϻ{�i0�:��q�!fE������� ���|�����/ɜ����5�h>�Y��?������Ӈ���K?���Q&f��Q�����'�3��1�Њ�B���>�BJ�C���¸{��WJ��&L�Jç���~�����(�X�/�Q����F�E�L�����BΡ�-�b�=`�� �W:�ȭ��v���Xw������]k���/,;/��ӣ����OG(�r{�S���Ͻ�w�-�5o�ȯR݆�˶����g�H���*�Z=��\�.����(_G�g���^-x��(=����=���%��'(�/4	��s+&;� �5����U	<�"}3��Nõ/Z�]��NI[��{���5�"�r��ͺ�v�ՁB�݌���^-:bB-�"y�7���_�Y��(�����^�P̪j�t�0����g�\�����g<��|(>{��2S�)kǪ�ٌ}'�&�I[7=���)�(�E� /餃A�M�8�fT��hXT�ڍ�w\�ж�V�xz�����7�W����G^�B�\��Po)��ᕨ�]S�43^�p������'n���wٸ��kP~�5����@=�����oZ��Sڸ6ϮT��v��8�<=�L5=��/`Mk�	���٬XS���]��j�xq�e
����_g�e$�0�!nQ�����^q�M�46e����Ə�~��~#��rD�\ԅ�Lt��Q>u0cA�+�K"�C�dSh��dN��ru�#���Z��,�C���kO-�%ы�k�$ӰkUf\�7[��ɵ%��� t	[K��k;#D�s�N!�7RCwt��·��_�~ ���93��� �y@�t��>��b��B���'#պ�j�~�#�3�
Y��(�!����Pů�ߐ��.��y�<�F�����{y����d�9,��,�3����;�/�)��Z��8AM��^p?�.�a���s@��+�2(�jdQ�i�}9N
�4��W��i ��s�i�jr��˴	���W(���\>ՃA��|�[��&� �N4�ҵq� ���z��X����h<1s���}_�4X1�R�/e�q����2*�6���ͻ&�4��:�Y0�R٪�(Y��I�8~��t��z��7������
�
�[^�2�:�� �B&�!,+&V�Ù�aR�}�,H;�7�OPQ�G��
�;�ý��ɱ_G��oF�n�I�s>s�w`b�Q�Yn�`{�;e]s�5�f\�4@����(?RҲ�)��4Ҥ__nd|ԩ�����F2��s3��k�	r���lA! �A<9xL�V�OB�����|x�HpP�F��\zhG���7K��6$�����Z���%��w��9����Js�� �BM�r�ݻl�v�W_�Yq]�Ω�z��*11y�ٻJ�o��Y7���5��6e��q��3�{�ϲ>^��(
�>̞S��U�*�t*��`�����\����?����cimYW|��S�s8//��ѽ=�zZ�聇J�)v�ѡp�N��ܨ������;Tr�&�������[*G�--�T��W]�YE`L��"�}�q��P�8��|ފ�g�z�뢰,�/2��8�	 ��(�*xk���[\'�:��V���M�0����!���U�n7II�5�0����=���gA����A@V�H�9�m�V�v�����DlO�cd���QC��'D(X�![*FT,#�o�g;׬rg��^9p���U	c�/u�d"�;+rG0��Ya�×�=���sK<����#0ֺ������%�Lϯ 0����� \�U����PCa��,Bo��(�x%���_��>�u-nf�t���Ng���QQ�(jiE~4�4`��\�_v?�)��G����'DtpD ��i}�o��s�H�w�6#�H#f��g���I���QK�'�qT�G�QM��N��H�x��1�1�pҕ��L�w������� Dϐϛ�.�l�迯B�̰	ZD�G�7)����E��+���Pm&�/d�,<Y�HA�T�v#suE-����U�i=���C�	�E�-7^��޳%���uֆ��{��i4�1}s�
gJ`�6L���+H=��a��7N�1��k|���8,��A��0p��Q&ϥ
gҐ@���Q)��<L�c��'���:�q{W���TT���[�5jO^�v����״`���%�x��g5�k����.��'��Jb��:j����`��W��Y���R�a���Pd3ܻEx
`��0��ֶS�pV�� �w��YS��o}��s[O�T��<N��8hm�ۺ#����3c�y�u@��R��M��7�k�,8L�J�P����\t��7�[���w�ۅ��y:��ժo*��.A���9�{,��PS�G a����|��#���;�O)��-]b>NxS�*]�F$�7,��:aN^fĕc�H���Zs�=��Hi�ȇ���m�@�����1��96�
�%P�Q ϑ�@6p��� �$VA�d�J��:�o��[�?V�t�L�`,(wL���)��]��?������۔NBY�T�w��z���_Б�@.�%�)��O��mtU��W'�łh3�x#���;�4�g�+�O�ҁ����<�����ıS�@��B'�	eHJվ+���U�[�9����U����H1�ġQ��b�B�!Df]i�dߊTz�/����ޏ���/3>��x��}�^W]�iƨ���Z9�o�6�a?��m/*�H?j���y��ُwZ��|�tg^N\�ƿ�	K���Wa/�����ynp$�(�h���l�xOcdN-�9NY{0�t;�-r5 �/�*�Gԫ��ݢ~T/ܫ��+����d���"|���^�vV�j%s�M�����Fԃ>��/	�/exQ�'ܜ*l6��}s�w�P�֟�T��>��4B;����U'��e蹄4�`�_9�����u���rt�H�9�,����x�7&����'_� 句|��g�#v�G#3���6M�'p�=<\ƛC��і̋�]p�՛`l��kD��m���}��6ZeF��@���v|� x�>�y��1�eW8oA�w%��n���P5,�Hf�JRk<"_D�Q�_�Z�v7Rf������L+��Z}r�(���������#~�����(�`@I᳌t��X��g���31'�P����Oð�\6?�ڹ��]r���j��c�8�;��������K,�l��1�WO�}�)�5R��q$S���$�������e���K�v�x��'N�3�S��/ָ����fev��lpA=�`�[�3����w�������;�QW��^*�L���VIN4��U���]��wf���H�^�(!�E�.;V�|z��V���O��Q#Ky�v��R�u.��� V�Q ������/�������ۀ83P�n+�Iz�Y�~?�L-��1}�NL�S�w�&�tg�070��&���k��t���h�Vr��{	~�A�H�/C�bH=Ƕ�Ǣ���#���t^����9Q��K
�}}��R�%̾`{m�'~����N��\��N>��1����ŽF]�ąoN���SuC�V��3��OK�&��xHeOKu���\��(d�Ԯw�di��S��c؏��N�¦k���ld�bt&t�n2#� :=T�	���u�!�SrۅQC����kH���[�=��5wp�*'�MF!�U�L%Tu	:T���8'����Ȳ=uT*D}����y������=�\[��e�TR*��)�،��6��q!���@��2d�?r���,{C���҆�"��W'��\���S\+������t<��M��L鋳����Y��~ϠR�T=�/���4K ,Y\�?�AԄ�6�/�֑/��5?��{��b��R�m%+*���̤D!8z)z��Erx6֫�G ���V�y�l��j���+X�������'��<��t+�ߚ2`}�0�V�:ty�Dd�A�oEYE�X:9Or��pIg�o��KEQ6~Mx�bΒ��X���6ǵwr����u�U�|��7q�D21|*��k_�L;�Л#Dʼ-E.Q�*�`�"!g�:� ��m���+�{S\�&$��sC�V��ٰo�|Ä�L���2r�ۑ:��u�L��g��6�;��}�|I�Ѧ}���㷪�V�P�������d�U
�+�˥i�]ĀW�!q�L�g�|=zZ�G�&�\U{y��#[��M�t�~�N�V�ga��s:��"��m�u�J���JՎ�����2��b3��c�`	�uk�a�����י��|�"��"fB��m=s/��#Z��d�7����F~	t��-��V��64� �u+~Š�r�l#X�!�㪜��*�+o휅C(b2�ǒD7�=Oq���/S�Dg����*��,�1�$i�i"Y`�fk	��7>�O�}�Xv�b.��|a�Y�8Ձ.���@����
۞OsW��1�0�5j�A��	�2.��}.N۴ڀB܁?aR�;�'�j����?f%�X�u �C�;���ǍF��(��Lo�[K�R���St��a��������-�	��ܖ�Ѓ��E��pG�ҧ����#{�,˳j��Ѷ����!��.����F$��տ���N�Tf�����_[#(k��^nn;����B�t;�.EP[,Bd������K%W��˪��˪��J)or�6t�C��%�	Q���aNo����Dr_Dr�4>�*�ʸ�f��T$U�(�{؂'Zt�T�#�Jq
���ú�%�����br�*$	Vl&�(?@��� �`��"�
�>f��К�\�)&[�� S�
�~�������;jA�N���&>��� �y�h��_{�>Y����rg��K���VQ˵�)���)���f�i�(�tڌ��oܰ��MDP���#����+x���y-�֯d��<��U��Ri [�OPԺ���h��(����XёB�nrO����Q>*������jѝ-��$c�gĪycRJt��7$�~�q�#�\�C]!�L(��F�v�岌ɇN��3�3�q|��>$��N���1�C�1�ڸڊ��T|fce�䜅p�Ŧ�y�c�j��pSn�Ht� ���M��4K��l
�icѦ��*����x����In�(��:��g��%�?�@��r�[$X�} wo��	����� �C�Y�O�Ӟ���^tQ��$���' ��X�閬`�/<پ�,̖��S��JB�̮�/7yxQ�T5�E d`v���?_<�?r�:�@�c ��tW� f#�O��/��PJZ!Io
6^��d�ts�Ddf��+�$�ʰ�#�u�z{���	{���·M��	j��C�_�:
�LH�^�'��N8%�*@%Hc����jB8�e�bA�qBb����jP9@��"���z�X|7�^J�Q&�c5~���FS}ؖ�p5����[�}�d°^7���jih�,'���T3��E����S�!N�|CJ��\��3h�Ԯ��aP�@�<�P�0���"�[���^�\�+��R@���/������� ��4�<���l.�"O�j}����/[t�n<>����Z)�!R��6�uؔ�W��s}
KPp�g� �|[�<�"�$�'0q���h7!b��N��1�lR�Ot��@�_'s�'u��ٗ�F�o��P��d�]]�*��U�ו��K��Co�2�,��ˁ��)�f�&�5����y����R���+�H�i�2������OY�u��i���ݬ��mp�$WO�7��n�fᅙ��	��%8���G�
�Qb`�7e>��Ҥ�.��S�CT��,WV�&��I8*''Ζ��U�lp(� !ϯS63�Ix�*ь<"��-�#�4>D��O�~�K����h	]�vSRcLM�O@?w��)Q�w%�����)�K�iv����rYa����N�o��.�4�g�4p��*�^'Ӂ���]j-�K�V0�ެ1;�Gt���Fu�� t��ރ��G�:�o�b���t:�^�_���Mm��v3�Ѕ*�P��K�)螦��+�?j�bo(�m�m�9��h.f?G��0hGs�/�s�����qG��i��ך�&4`���
Ȏ�$ �����!q�T�Z�	�^�e(��.���|��(���Y��0��^eg��H�У��r���� ��h��:8�K�����{J\�G^�2�":Uc;F$j����׮7]T>q��G�vL�CoS�M'p��W}@#Kw��EkM<`t�$�KG ���]�6�0���F����q���Z[�̢�����y2S����m�Y����ʮV��ϛ�gX~�<�Eч�+ݹ!����{�·�$P̋LO�}�6�� ؞�w����������Y]{���1o}ؕ�o��� �RyG뷪SSwC`8y̬��w�Ij&�S��������q�sN6×>�|j��:�k�w�^�CYE�QJ5а�  ��':��zC�9�ǒ��=���`���V��jdq�g�XO�k�7�/3+�?�D\Aё��E�>����[�/Q�Ri�T�<X5��ӗ�3����&c�Q0D�/P.)#ty�[~�f�mY#���l����Cc��c
���S�0m��pR�d�"����*G�ϛ]JE�
A���\n~�p����r5,����.�tXh���2Veݗ���:����OСޠcf��0Z[�4DT����B��!�>��{Lau�L
iYY��Wq,�e�ڗ^�yb��oh��jz�iE �GN
Ĭt��m��WuwF�ږ�SVyn��֓Qsv,�+(�J�:`w�~�dr�<�R�m;d
,K��Y�� 6�u��u-��8��no�&R�>w�vY�����_�m�<��,]{|�J�p�������m��o���xYT*���<@�ـ  !�2�J��*O�A%B��L��K/����w�	�)Q�MׇQ��{�e��C�GH�y�-�㷩m�ZB՝&^�C� ^���Ÿ�c�ʐrʺ-��C�1p�n��ѣ�P<f
�Jݾ�i����BX2A_,�����e{�x���A�׍`Ig<{w-��ՒVt:8,�Ð0��5���AU-�O>}����Yp��:�N�F�k�r�:��/d�_���E�W�j�r#5�$D��ߡ|~^=J9���n�?L���=�4�΃q�aB�:�3��W��i$��h1��[��S�������T]Jq�
"�՜�\�"Ҩ�2g�d�Y�h�^�ݸ+1�����

�W}G�_l�_`��[�B����<n��q�c��IP�MƼ;2d�ո��i��:r�+��sH����J��^񈍳��r���[ ����),?���s�O�MP\�� Fa^S�{ q�A��z�?4��`v_���|Et�K�aP�z��%U��X��d�'�3Fc0�S\�v5�`���`CH~&S�5��_=�n��<�j<(
_w�2���w�I\�~Ef")���'���G�t�)	���[&ep^��l`\����%�����[J�$x���T��Mb�	�n�m��K��ɞ���?p(]QnF�w2x,� T+(�N}l��|U5�/Dм
��U ^�m���T�tu�F���PD��ͤ?�0�y����p`|�S�E��
��+������õ�b����NK*�6_�*� �s9NEbRC=˥��|���=H�Mv�(SZU]x`�C�,�w?g��e*F��ƾ������;�s��d��%}���y�F��2?�Ŷ��%U�J��>�2A�	�ˋ����Օ��C��cd���@ȃX���6�U�J�hK�	�)t��������������S],�:-�I:h=#1+����#*�!>nRA������vjv�������	!j���N�0�����M�7�a�ɍ�&�s��{c��=�V	���AH����ߠ\0�n�2�K��_��ތ�P���r�#CC��l5��3{�ީ8(.��Ǳ�Y�#ɻ�z�m�ڵmi��݆9���P�ک��!g���W���]󀧃�c*g�����b�������_�F�]����}��c�X��W=�3��(7w�m`@�09���C��b���U�I��t��uE��f
x"Wg T|"� ��)�A��Ⱥ�j����8�(B"ٔ2M����Ɩ�]�X
T�P��Z�F��,��{ix,�e�"]M�O*ʣ_UD2x����}3Gg3J4ê0��� ){�p41�dc��A��`���U3��,��0�� �Ƨ�8��6����;����o%a�<��>>)uC�@Wp����Z�z]����+ B��43��TI嘣��Զ	`�����8��y�<mDقY�/7�d��J����4e������tcaK�o�ʙ��n��ZX�]�,
1w��1�ヱS�:ES�*�J&�t?�! c6Q���+鹋7��.b��ЏU��L�{;ҰiN�Y�wh���P���w�������n �@S$�qS�iZ.ۤ���5��D�v�)�͕�� by��	mK�[
�I��t}G��&�8�t]��q�����ZА�K%e��9�p�N�9��!�p� s���=\���u�6�]Nbi���@�:�bOwp%��c��ikm��d�	҅���Q�7'�}U#0����ى2 ��t69�f��'o5Ҙ9[I,��+���R�2V���'�ΨS��I�e�t���(:�@��o)
V�9�N�7�u)A�b'�j���5>����t��8�R�����h5�c�YM�&5�z��>�`C�����67W�c3���jَY,��K&Uu��Zi�����q?�P�l)ף��D����Ă[���p避�20E�k]���$v�ʳ�n��Djl'9fzf���TJ]��g3��)��1��g���1�+�Gg3�>����Xd�(�k˞��۷��J?��<4�Y�y�)�M��}��x2|ǋ3.�0�s����U\�[�sS$r����<�$[B;�L*g����,,�B���ok�J�8��0Vx�	�C\ޝ�F�v�ѝ������.�[m
0���8o��g|�Z��h�,�!��Zt%���2�	o��qT��ܞ9���#��l�Wĳtaf�N�8z��#�M��2��*c�%U���敖w��d�)ࢩ$�=�|��v��1r�U�/�8�~�;t�X@&9��^ED��	0�\��aϖT60$~����=b�g)�dX��0̇�l|8�W9�!߃7�M�G�j{����[�y=��d����Q��1��T����4�z�B�k�h�g�R����7�?׷��/e�ĹpZ{F5�d:`��\�r=��"d�A���~([,�kwŔX�cS���h�)Sڏ��{&��.��|�:���=�Yds�\��X��W�=��1c��1�a@�z�A�puQ�O�O���8�Z����d+Yu�U�R��@m�&��R�&����	�cr�E�Q�-�JF]N���ؠ�gXz8�P*�x���Dp��4�j�@9�Rxo��ER�k6��2!��@���dB?�"�GNB΂�?׳�O���Ձ֚,�M�.�P�fE(cC�+�*����0c��η8�rIw�=�-6&#8;������ӓ�g�F�M��a併/
�2)t������q�H�i
��34���ͬ�9!��@���P-�0�@�����O����}>�U���R�M���Q�Ai�����4/"�RIϚ�A�S��c��o�I���uB#<���D��.��^����%��`?r�Ѫd����z���Q�	@��U�ӟ����Y{��qJ���9i�Z�,�%��>`6��7��i��C�<�cQ2]��dц���ዄ�KІ���(��~�qS�M��)!w?x�B�q�,�ܔs>w�Q	A24�M\u�6����;��ќK����A�Y�!Ymz�/�[��x��r�Z�b��m�n�(֬)�{(�[���n�+wP
��h����䑺
L��|�ٲ'*��xaE��\�L�E��󂻻ףE�F8�5[2���(u0I|)�dN~׊�giK�4 g�v���=.EEW�7-{���#����;����E\8�/E=Mֶ���h4>�O�W50c��YLH��t����
{=��E��'n�f�[<�;g���]���ա�R��|�٩a�:+�=t�}z�S�d�_�+��G��V�����eMy���2� ӑ�����������Gݏ�	P8��0�=B{D�{r=<4ќ+Ji��e2^J�����E��f��I2Z�`u���@5���|�>+̅�>�� r����>Z��Y{�LsXV�Q�W�U��5�q��=�p+bT=���[�~���s5��x��d���ht��tx��
?O5�2	�5z�|�i�߳P�mO�%��s������Q��]��������I��p�	��'�C���fi��[�=���J������-�x�W33�"�����"�P����4�F��e�����	Q!�l�h����ŅRx�)F�_�Z�-�j�x���k@]�"7�^���OH{�N!�K�-�6��X��`�d]¹�vO�Yi�t��OOb�b�L�y/,�}�Q��{w�5 ����P����GK��pg����Z�ݑa��B�����%��`ΕI�
��a�k�� ~�W��WGF�+<,�����ۍ�5CP��OŔ����ϖ��nUq�C"���1�3Kh}_�������&	0&��>�rdj8�Q��y�k��B'D���k�9ʉ� 	��V�����u����W���i��y������E�8ã��qoq|]���9
z7��F��l�N��j��ѯ�Ֆ��R/
�z�K�K��E��S\/}��E/��WG����Q� K{�)��E��`bA�-����˥���	DmX�룳E�ڠ��s�$T�A�~~X�-[�Pr�5������R����@lh�F����~V�Bᖬٞ̃G��ٽ��?|\ߴؕ���D{�T �!�GID0f@S��E�t}�-�s���>�th�T�=��``m|�����M�iJ��i�qέ���O��ިɴ��lt�ߩJ�B��iΕ��*zm]��K�`�-�F���sAЍ|��٧ 9�ue��B�N��a`�&dC"
{��Mi�<�O��j�gf�=����p�8�LT��+˰�oY ��r68��}O�j�(�r�E.Gm�S�q���o����ǡT�g�I��c�[F�{owE��"�,0��x`�O�=�&s��ӵ�9;m��O�
T��SC�;x�R2W��$[Q���4�!$��H�Ս���G4������Lk.�=��}c�Q(�f.����=E8�6��� ��&� �i�s�!�\�tW�B`!�TF��|�;�5rV��QDv���L��C.��,_��5�>
W� 1=�y�l��/\.fK�W$�9�Et��6�?���͖������Ş���2� �"o�}'l!W��1�Kk>���`i,T�� ��87�_�=�n�xb槞�,|� ��,����xM���4�����AU��jQ�#
ړ�����L{;�̛O���2l;�?P��1LL����ѳ:�B�l�V�7�k���2F-���_��L�u��?F=%�X��q�]���^�F���*&�9`�.�\;�� 	.%��F�����a��D�M<h�*�hc�BA�<��2�[�1EU��$o҄�������a���<*C,.�c;�	�*&z�JT����7�x��l �2f����:�����⢨\��+`r�.�d�$9�u2���NZ�Z��w����F��A�J��1_�M���6��Eq,:����۸(�pd�Y�	.ӛ�m@Ȑ�s�trZ?�FN�^�OCu�>��?�݇��7��,�����gn��6�䷈��z��W�Z�V�цۇ�N��y�'��ʖ"4c+��Kb7}�o�`���.M�UB�V<���Mә�T����nnدcqq�k
wC�*-�a���5�����(��V��,\<����>�;��f���.67Py���ׁPP�k�:���Y�Π<h4+�p��D�$�~�"U�9_]t���ǥS���UN��[����څ�dʊ`f�=e��~���x	5��u�)מ$yl6(���xE��(Y�`�*G��nQӍ�
^)|<��Od��Vx8<fF0!���Z|��zڈ'�;:%���͞V�� ���J$+YVsWgNkw-�;b���E��?�O��Mo�t0&�M�4m9hO�Z��$
�i"nE�tG�j�J	N��霷�D�����)9��˿��A��.�37�Th�@����E�K#��F��(�u��ss�pr]��Q���M��������Z��'#���0THݴu���٪L[��xUC�i�J�?`?%������e�Yu�ߓ<tɷ;���/A�p����iJ��#�;�O��œ[��ծp���	�� ���r�d��JUyG�@sƷ;���wTe-Pn*��a�*G��m�ׁ�*���Mwk4��s`/��3 γ���V�����D�����?�F�����$�[�� �A&�׭�;�V�m�������i�r�@�wGΜ|ɦ{���T[�ΉF��#�y[chHX�gƫ.&ƕ���x���(a�<b>*�jl�)H5�����ґY=�_L2Ar�fV�*ѡYgb�~�ѿ����1�_f��B~Ǧ˸R�vo�lL%��{����%�6��C�^�NH��3����Dl��?Q[B��{m.���0 ,O�+��	/�%�Ǚ�O���Tt�XbDm��{�r�������KZGoxDd5L�+�rI(N��f$mW�����K܍�.��e�qM�$l���s�Q���?l�
��y㝢
�j��/����e���0��+P�`:P�@�Y�� �/G�b2��������}�<[���QMP�\D��p����ϖv�(�����R�)"2��F?�<P�͕�oC���X�C��&C�?j"�we������܇!]6q0*O����ԭ�	 p����y�5�o<obx��=������0�
�&�e�R`���;�
3$�b'l��{���$��i�q�$Q�{��@5��N��#���G��l�P�UC_��P�>�����wp�*��yp%-��4e��En!�����R��G���dtZ@�&SXY�0no��0��}�te�8[�S6�N�>�|�Яp��4:GU"-C][@z��Ƅ|۪�����I��1��Ԫ]	D-]A8��Y���F�a� ��J	1���
{u5}LC+�m�i���+�2�%���s��e� }M���3'r��r�J^�P.�9ŰoP���+�ӟ�h�Կ�a㛌FN�2�Й�����,Gͷ�� �U��[�P�!�M�^ן��ye96-�$w0��%�?�3E��Ƈsȼ��%��){cXuN��y��xrlL��%M�/��'�}� ��7?}��_ K_���Tɝ�ʧȅ&)� IW&�w{�������¾���d��KT+;M��	��BY����ϵ�OR��`�v����Kȍ��L��3���{�^��iM��G����II�7�I�*����m�d��o����Ҭ��������n$?;�V��I#�::��>�u�G�,�=+��`��-_�y;����2B-2�Xw�z;�T�PB;~�.��k�D�
�i��c^bv���!�"]�����KF(apJ_mC�+ *�ߨi��"H�|Ǵ����E�Ө��Baj���bF<���9]T�������f<:��^��|T�y����m��i�k���eL8(�o)�a����+�K��kƙ�2��WnQ'�WǤ[^�@����2h����9kފ,F^�/���Ϊ�o��z�U���:0���0SÌ�����e�7�K.��u�2ߣ���÷��Z��'F�H!<0�Q9�l�!1"�>���
���~�Ƹ�#;���
�"�I���Z�
Ɩ����*7#������Id)�H��0dxM��Q����
�1��Ѷ��j{��g��R�����~��-��aꧩ����:�P"������#��c�v���K��+Qh���b��\$����K������x�ƃ<g�H���Mn��
zE�����*o.[�<�bj����x�ь������7/����aZfX���9B�.1��Q�ˉ��<�hНxA�����yS9;p߁��0\ye	~d�cj��5Sk��ɠѝ�w���l�A�@�|�%:���A39��Mޭ"*O��&X�2@y�3j�{�-S�v��仺'0lv�&N�p�:V�6����T0neb�X�
�vA�d�-Eכ����G%A���d�֛l+B��uؕ�z�r25�5������Zb`5��������jX�}��z�-
dL�����Q_�S]}�U�D10(�vh����� �9��}��7��q<���B��w�94���<r�2�5�}�RX2�������ԃR����E�Z�lW*�4I�N�� �
�^�����lٓ��R�Aޛ*��P��"�K�I�K��3!��k�N�+s���@bo��a���2B-�'�̼����w-�rM���w��e~����n���5��[�T<�D(�Dj���\i�'Aļ�H�;�^����҃';it��<_zz��k�De�3�g�^U�����V�����y�a�?]ہ�e���]p!�gz�l"��QuOE�0��{`Z���e����Un �t��
�S&e��J�#u�o�����ۛR�0������Ӽ�{�/�]W\��{'K�br�ty���֠��P���l���V��w:�����\�;r�*�����޶! ݆;0G��C6��o��y)
�����A>�	���T����<U��z�e����/D�:�Q��z�N�gU]ɛOʡ�U�0k����LSH]B��+��[<4�B{,_8��]��3-ES�M�fO�k5']��i���Y�RS�4o�;?�M�)��G;bhj��0g0k%,-G>"��Nl�H�<;�,(�gZⳎfKT}�4�{�ٴә����!"�u�D
��箇�)�Ba�����=(c��������9������@���(�a
f��{{�(�B�ܲE���M�G��� �)�i�Go\�Esq�zG�MÑ���z�5�o�˅fχ-%�ǳ�^L��M�m+�De=����:��Ē��M�%%fF�̎�f�	)���l�����";�%��1Y6E�ř�տ���g��.L�CO�8+,�GK�~�0Ew�g�DX�,�$@:d��aQ]���ڿ�xM�������B$�܀�5��+��k3��"��!ޥ"��DR|����Jݓ��F3��CXy;��c��	/X�J�s>����MsC�q�~=�߾��xn�P�E9nY�u��*�N�Jڹ�G%u;ҹ�;������ؘ��k4$$ ��y��1���k2}�ɨ
�X-���,VJe�:��ޛ�{�z�V�Q�Gs�����ȱ��T�0e3"�E&�p�ӌ�cd=���Ǟ��wzhp��>�F�m�!]>Wa�򋢜��0ѹ6��ufM��rd9oH��y��іD�|�<9@#��Z̮�n�|��WCx`�'W���p�nՙhc��|�.��h܋�7�5��#�˸�5EC��9a�n��W>�mM*��<ߩ�8�YN&���xŬ���H_t4�P��(�	�x��;�x��m	 0���v�|���Hp熣�ؐ��x/,[.l_)�o�}�RR(����΅M�0���<]�4�������&���[_�w�
��8��8*�������a�b��O]��т9��"���J� ���N�v���>.�������F��Da�	���9J�8��i�W�g�
�;�&H1�r2S��L���q��yq�a�xIv�̭a���/}د��qXm�J.�[�R�)Oc?qz���m��x�id�c5�>h�t������Tu�O<G���% �����h��{w�L
q�w��μ�� ٮ0<vV	���[��w#iq�.N�,�;{ܕg�$�:��B+����UI: ~���M����W4�F<T}�[}������%갛�۰XW^������f]��V�ER�J�I	#¼-nݜ�Q�r�r>֥f��n��c�`��t*ܳ�*����2o]^��:�X
�t0v:8���ekSOQ���q8	��E�RC;~��M��o)���5�����WY��n;��' ��������L����v�-�#A��9�)zm�Y�P�g�Ls�c0�c�ύ[�fۉ��V*�K�KM��������+5�_�ׯ�4�؃�W8⻟���`+M-��o@l��d���JI����^#q�IoXea�	zZ�6��[��)?v%x�4!f�����aI��1*S)E��?�:�_�_U��������Yn�^�.
��,�`k�m��Ȩ�O�k�W�qy�r?9�?<.��w���_��[6�WwI3�=����������27Ə���U&;,�m#W�)S�j�M�;Nf,�.��mY~�����p�3"C�)\N���Kh��������*�A%�ɐ�q�X�b�M(G�ҋ��5B&�eo�P� ��tj�#.��>_6�)��i ֝fJޤ���5�o�����y�h�%'���T�D����:0�]���)կ�o�7��O�_V+_� �j��W'�l����1������0v}�w5,]��`[Z�!��j;�����^�{U��b�[(EE�te�w��V>�SF�NY4��!ƥ����[�N�\	u0���mry�M�3� I�����<�1�G	~{|l$�6.É�/��i�oYU��P�WqKRC��j�� }���1~o���k��=y����]ZS8��YӆHM����ڥgˈr�y(r���c!!!M�}�M9!���M��ӎ��ޥ�N򢜷��T��98�JqTOB��@�vPo�P�;*[t_�������o��=����j�M���:&'��N에8���g%"9���a)�]fE��oz`�A�)��+�W )mC�E(�$���y&&������-��]]�2�+<lv��AC''�d�\`�[D�*��jٜ�%-��(e���-�����ޏ�*I-���u���#a�t.w�n�/�0B�ضǟa�E�_��1�W�(3,$mf���0����̵b��k��t���^}M,���_l pSgi��/Z�������A>�	L�5���l��
>j�Xf�{*;��u��*[5�>��v;x�S'�����t���l�C���O�7	MmLh���Za-���K6��uh�p�����y:fM�(�:@=�����d���,5��$*�<Z�i,�Ͼ�`�� NN��?�ZJ��+� Z����~�
�yM��n{1uw�Ћd�;��^r@�]�?PT�q��HQ.+�"�Y%Yڕ��r��C��ए�|()�%/#��J+�?Isl�{�Y��<�Ѳ�.祝t`Z7����Q�xDy����_Ii�LK~��g�]�5���TH�0���2���.A���>��6ssԦi1�;�F$�7Ѧ��
�#Xt&��1" Sƨ�lݤjK�_H��b��o�gǗjݿE(I���:��T�'uڏ͍���Zb&��v(`��Y�p�� %��K<,��6�q_`�5��m�)_��Y�	�+���d��xb}� 	�t�?�(O
Bp�/�Nt��f�wc!��ֶ�C7<���<���ѶI����S�$\�XM����0]�i$�{,F�^�'f�-�����i��y�����.Nk�8�^�qL�#Y�i���c�� �Q$��$>�u;*�u���J�ZǬ���ۏ��f����.\��g�ܯ�[�x_����y��ֶ��	<
�rG�1I�ғ��6C�Y�Z�����x��=���4b�Q��Մ�n5�X�ٴ�U��Eq�	y3 �h�4�>���K냮���WO��ы������η�ڐ�0���Z�*�N�"�y�[�@�'f���0Y���3&�Mo�d�Ī���q�Li�$:8�y�W�u��Iw���dٵ�����o�_����E	ǋ>IR�^��]������B�#&�&Ǐ��s7��}�4�f�b����"�?�ʇ�ci�O��FI��sO\&���4���)��Ak!h&f*��ZȌ ���U��g5�5��N]Q��ڞ�S._ S�?v%pmz��ڐڥ�5q�s�C{,+��]]�U���Gu":�bo/�q��c��E�������o7��W��#T���R5�|�����?~���/@�����d��0��y���9�ߢ�dW�{?�'�9���Jx�I���)�0�j�[��vv?����c��W�O�ۓ�7���V�j�Dϟ��_�ui��~���Ҷ�'���zU�$�yPΤWC��-a�+ݝ�p[�{�vf)5ؿ�ڠk����DG�'8�,�s�T���A�҇�z�B��i4a����EFk���CL��� 9w��6{�H��nI���Y�q�za�9Ҹ���V*a)���}N�s��������3��*[�;S�����w�E��o$cʯ��c��5|��
��'�5?�N�S5��f����pH�2S�-H��p&��~oa�m
� dI�T1ٞ�L�gނ�rވ��{W�����}&B��[�ό[\���}�Sz����B$���a�9g�"�����ߗӠ�1���76���Z.��;G��ؑ^�V�dJ9����ޖ�L޹<���)k$b.�C?at�������1�]��]?���r�rB��A�����I�O�t��ΚV�R��������>3�Y��z���f���EVA��{ڙ��b��t,���\><G1���k
�k�Ȣ��4>O�f��rό�j�������H���s)$�7�m^w!a���ɉ�6kV��q:��4퓿K��p������vBmx~E���/kU`˔<��� �cU�͞��-�[��#8�Z� �t�?��i��3�. �����b<i��eL��ls����=��6�����	��z�g
�P���ЇJ�R����N9�q!T��y����0�p�KЅo�;�B�x�a�W%�d�ؚ��+��V[匏7�:��T*�WH������b)�� �ʾ�i��	���gv�d�UA�~¥W{���//y�j�7�p|M���~buW��`L"8�GS������aK[,=�8O���'
��s�7}�f��Ʃ8)���x�{i�s�ɘ�^+f�f���*]f��ׅ=���L���(��� �Zi�{.��W��$O��JL��]�<;Gb�� V�
s��.����ϡPWqR�y����~��Zv�8�l����W1^1
�&���ۢ�P\�c�S_���������些�+��B��Z���Z�P@h`&��&�����C��lR��?R�$�`Y����Y���S�K&{Ց�տWXk��c�[7V=�����8=��D����U^��=l�<\��:��&o����篺�7)�b��]�ʺ}�����#!��O�~aO�N���� �5�Q�����\z�}%���C��'�T�n���ɭ��X�g��5��I+�8#�@"�]����^�����R����W><?�Ьr�ջ�:W��D�����Sb�SU�-��0W��CUhLXJ_g'����b�qX����xirmn�
[1�������sN�]�Tnp3X]zu{g��⽷3�b������2��S4C#����:��$�>-���<R�r��G��job��)��
ʣE�������.�s������(IHa�h;p7:�1c�#��N�4�u�	��?��� ��1�%E�.Uy�Z�ÅΌѧ�I�^����|�?�c��q_�Z��̠(�'��DKŭB=�:�^qzYiq����mb6��:X`��C /**|Ӊl���� ,����_RW�
�$/�bc���,�]D\���q�����R6a��S���8�(f3���E�IT�,�
��M�����)��({(�8�G�it)V�A��c�Uu/�-"���Ⱥ�c�� E�!�a���cY�)�l�AF�`k�+o7�4�.�F��b#�s`�v�^�9��%1R�~p�xuG8Ssr2�(��ϵ�&�։� �G�� ��F*�"�n����e*�j2�wKZhQ�AAVa��Z[ 	R�cد��A�#�[���(�(p�ll�	��<��B�~^7NJ"�3�u���w���ql�`o��h����汅���U�%��!��
�ڰNȺ&�4ڼc;T>����=T��M6b*A�-aW.�(���0�ڔ�H>�Q�u��4P*������0�0d���.I���	(�*��\hZ�=�戾��:�b��q����*���B���Awhp�=(F�vB]6̕�,˙������3��F|PAŮ�ܓ�ٚ��D��<�.Q�,?�̃-G9􋐥�l��o���o1	zl魆>�,��S�����}C9v�eO���<�A�[�-��v�UP˟w�%0���Jf�b��^�Kq�&z-FZj��^��TD�������HN��$� N.U���Y~e�H-��%�P���Zz��#O��=���M ��Ө�c{��J��PM��~_֬�̀P=����Q������f�B|��>c|�N���e���������I/�0���*XvS[�3��V�,�9nk�5�PuB	U�\[�S&�j�s������ȸ�5rnȍ ��ρZ�^7����]��xúC�8~�q�
gz���Sa����FhCh��/unqEq�=�{�u/���Lyk{7�S8�qw#I��J�L�$�R0�w�N\��F·�pu��.()�H
1s�nY��P��1:|��"Q�ek]�����B�9:�K{�͘؜�Q`
�C	>U��#�{�C;,U��ݱ�ݟ�X���|�)#����7����}̝�tP���:1>pчcHDR:!�cݳz�~��E�*#GK6)�h��p2y���,�e���������Y+-�R�R��;�����R9�g�83�Nm��^4s�������i�e��f��>���?�5Y]?~7����H�˱5�o��8]EJ X,8�rK�&9w>�V���D���&�y�D�RӰ����G�1O����Kr�Fu����Ȼz|M1�RIw�D��[���n&�쪭����x��IFO�N5����T]~���ܤ9]���K1�0�$� �z��Ur�pbY����ۿ(�H
j�;�~m���W|-¦{���υpn�=�����=�<��	� �mͩa(]�z��WF���Oc�+�:����d�W��c��� L��'���>��Q�A�h�1KWi�i���Y�����m%npQ�~�oP�m)�R�:��W5h���PB�L��T�袕��Z��r�P{i��Ā�/�[���0�.n��9ݽ����tK���J��{�۫	=��s�M�*�t���8�j�z�Q��Pz�6���"[ވHB�ox�ڲ3�K���+��b��K�������������E4y
���8�8��h�RF"lം�r��O�b]k��?f=h߿3�v'��,���@���R�~}U����w�W^�G�������|oI�g�n!��`Ln�螬��Q@a��tɹ�Z�e�����^�c�<{�n�+��wL��TF��WRH��KS(A�J)�G�`C�Ȏ�W݋0�`<ZO"�\�%��"��܇���wM��.0�
��B;>�&�t�r�"t�{����+7E����/�w=�;'��%l�y=��;{{�]��@`盭Q�P�~ȒL���x��>&������<���$�F�=�<�?cf	���"��?^5����OO�Z��
�j�(/���	��T�R�l5<%c��W���k;��s,�s'�T���Τ���
�#���X��067eP��@gI����"�9�'�#͘�g�7�h�叒������sK"-f(���Jysk ��]����ӻz����\�e&8FCH�{�뿪���`bc��R��7Į�J\�~{�l��ʾO�S��f��Ш�5�����{���@��dj�&S��~S��Kt|Z�"������#8d��:W��=�γE@g��'.�^KBUE�Id��ihP�a:a�A,`zY�.�a��<�H�L0�E`�������,j���&��q�I�
�[չIR��U}�;� ��c�j�,Uk�.�.�MOB�r>�/�Wp���t�u�tj�]���ʚ�Z���"��$U1��]}���  �xY����[�Zq���8����~f!m(����fxf��`$��3���e���t������ӡwÿ�����s�t�*���>���H����k2����i����p�|H���?v�ɩ�&��r���a�q^�p+���R��r�icu��[?q��gS]u��fr�Uu�C[?���������ϯ��0&>|������rM��uS�j:��n�;�g��4�VՆ�{� W�b�w��1rʺ�����u0QF\n�U��=��>��;�V=(<��Yk����>��s3�d2�M�	"0�K�b����-�1����V��tƖ`��j�I�+��c�_���8V@����[���0�ߓQ�y�M<�HN��'D�m��C'7�X8��r1����:_��s.>N��W�����}������b=şe���>��������,�= R����<���E��w`n��:�6���h��t,�h�;��\���z��J��F��C��2�ÇT��2#>�͛�(Д��)���ϟ�E���ؔD���W��J�E�朕���s?TVPk��%%R���)��.5��O���|Oa�1z��A;����P�[��=Gy*�7�V�i�W��}�W�2��'��f�y+���
��؆�x�<}�ΰ�>���g���]����ݩj7y�#��(���q7�t�����mӒX�x��Hq¦����Op�3�<3�f�z�V�?��T;�7�I az1��=<�I[m����2�O�G)+�F�#�D�.�c�3��O�7���Θj}H?��~N�%U
�^0<v����1�'�פ��}P��-l�>~b��c(s}�� ��/~�}��5�f�y�|&��AL���cW��AS�HF����1ld)��t�A㿊�����Bؼ�&�S��:&t7v+T�q�(�}�t_{�f���E�W��?����C�s�я��ӯ�Kb�mY���ߖ�Rv��K
���[�Uj�ߩ�!K7e��2��o#+-�����%���Z7JГWv���҂˩aK�h��*��7F�������.'��VΰE�.�сLz��G'l<;�x$�R��!VZ��s+��V��f{�p��;�������%5����LMz�8^w��Y_آo�������+1n˧y�U�I�WA�����?�`!B3Լ���L��t�S�V0��^2\�]����D�����钶��G����u�Kg��d8n�*�L͖(�DEyR:����	�ub��8
���',�P�hk��6{-Z���8�vҒ�$�r��X5Ц/��'���'����^7$�������>F �2�B�c�b��Vy[�?�Cn���S��{�$��kL׮�k
Ƥ� �\ᓬ2���5�˹{i4��!�T9�IP-����3����_n{ �|��ؼf 
V}�K��N�p!B�����nSA�D��V�P�۱�Y�Q(�{�Q� �zZI�_H;g��a���� ¼X�1#`B�q/���]CN���b�8
��D�y�����μ�������S�n���c,J����5�vވJ�D+��ī&�:rG�m�4Uv�,��`ɞ)w�mAu���'C�n���[uky�C�$ҰjI.����w�l���$��'0�� � �8hڪi5'���"/���P�4�Ĉ�d��01G�-B��i�c��0���ں��G�R6Wu��y ��uV,x`�!�2�2YR�Q��7^�4�4���q���?�j;j ��	��?�v�9L���(����/@�J*w�~���g�Ѹ��CD��D�"eiy�]m\��c��Lc_$ f�g��.��h�a ��_O�P�z�E�Rxk�r����ji����lXm�H��Y�Y4t�3�d��=����	X��]�UΫ+\��_4�8ZN�҉"��"py����a�q��c�.aLi/sx~�#n�x��G�P�?N+�����*�V�01V�&�S�InǤ�S.S��Q�3�N�}���ެa;B�Hx	CYnyȈ��r'�x Ǒ�ܽ< q+�#t�}�P�6��F�O۽��#�t`����c[WI�Ϲʷ0��.#FzvV�g�6ʮL�;p#&��B}s�#ـ;�v^�����l5
ϪY���i�ʭ]� 7)�=���(�ۇ����9�3$��#�K��|�>�5�ћ�)�p�+�y#>�bmY>�0�c�Ǆ����S���e؁{̃"6h��)�C/�c����i�d�Q�Ip�a���$�y�j(c[M#�CA^��.]����,���m�Kwt%���P�	�WZs�8Qs|��L������ {`*Z �@v��W�W���*�&� � V"HU��r�@р�F>��,�S�ut�l&�|"F��+�>�M��b4����h�J��U��W�Z�Dcq��(�+�ڋO��F9���b|�߮������dv��1�,	ڂڰzR��.���K��xI�;ԡ���3Q������kYk��Cn�I�Ջ��� /�$�k��=O�L8A�G+5��l�|��N��mH9kJ����F��ؒ8�f�kc?�=�A�pG�<�'��������8�vu�켑��襶I�)�b��w[��H�dg�{� �wlC|�aJ��w
��#�:=*�y�E<>��x�#ʈ�+CdE���Au��$�S	�i� ���mU���-�5�`���2�<�9�6?���<Z�E�p%l==��.R�N���e�mDf��f���R9��o�\��`����!U���S`�u7��H��!t�EZ�Bj�,W{����"�D�E�s�����]-�J40��]���3?�:�b1+�~�� �L�\3Yr!�%�֒�S\S�)�a����<+e��=��bv?�f�28�V�)kc�i�ӆ5����B$��}:�\[���M��P�t��[����V~^o^wX�����5��[w��`��@�4T�G�2����Bg��Mݦ��#q�l�'�U�M�����9�n�n��gZ0Q�S���׎��S����X��Z�m5�0Yb� �W�����~�t>�G�N�e#����۹��%�[�r��+&ڜ��]P)����)��� �MD�K%�6SD�U�d��k�к�X���u@����\�N���`t�}�+3� ۤ�p�-Iw�v��	>P�쀫�;C���3sPK!������|��D����&C�V�p-� �C�7�]poռ��2g�J����С ,��	�!H��<��)J��6�n���J��t�䪗OK�G�T���[��Z�V���"Ďl�e���FP�����~.�c�:���m�� {W�D�|�ě*�ȼ� J��B��Z��%J�k;+�֛e�~��~'EP��B]R�l�<��BG�Mх�׃|������~ǩ��D%�Sתܛ����P3RV���V��3M���&ơ���M����Fy/�O�����Ce��6�L+Js$��b\�:9�QT��BW��Tx �$R�� ,/�'��P5�XNt�4j� c[Ͽe���=z� �6-��ɷ�r���Ft�wB��f���B
~���&j�t�E���_v��C3�m�XY&��d萻.��TF!/�*�߅�$�!���u�ٙ�P��b��q����D�:���QY�M�47uG�HW��Q|F�ؾc�!��V��G���-��S�W˒`��Y���ac��B��NJ�P��p�Y�`G�7����5}�
	��������oI���e�ھ�M���w�1~�2A��͔�I.��h�|�	tiQD9e}l'�J���#r>����P��P�z%PK4߃�8E�]{c]��ͼ1VÀ�n8��̦����LО~}a��>=MB�W^3��f_d��Px.�k1,Ĺ9I��*�hF����;,�%xB/�s];�ck�1�mLӄo��#T�-�:���wi�&�"�r�T��@ v��mn^0,��6y�s>�0�3��3vl�G���pi�}�w#5�e��!�x�Հ\��Z���	��N�ٳ��4&��_)�oQ+<���^2]��Y{ۻ��Oto�z�}F���`�Dkl �80)#b�/VU�rb�Qi��W��c��V;��c��m-S��R��E��7�� Y�B��5p�!�4ɋy�a���Զ�Q�X��� ����p��Ooe-��O���ܘ��wR�ƈ��^)�ʴ0��V,iYRν�nϣ��`m���"� �R��91~ek�!�Xu[���\5����Y �o۷'>|�yy�Bĉ�ʧ� S�1t}h��E���/�{4�`��CH�k(g#L������ϵ ᚴ w�΄8h�7n_���=+�m
�,d\��)��󒉑D(^��#0!����7"Q�	,Q�i���0��BS�|e�m���A2ڤ�4�]����e��6��-"3��?#�0�t��[�e��/�5��zU��P��^$-d�d._z�Q�]��;�?q̸�AS��)R`��HW!)���+C=���C8�2�����t��t���J�IT�QHDn�]2��/@�M��j5��$4�!��ݶ@��L��s�N|_<�t�@�1�n��Al��>b���3ΏE��`�È�,5���Y�X�%Dq�K16V�ͥV��\��Y�7��e�5�UW`n؊tJf��җ��s����`���qƁ�tj��B���rf#�m	m2�<�V�?fq5H����J�4���w���b����'dh�=b�.B�=n�qy��%!~�S�7u�Oι�F$g�O>m��5^+oc�q��𛇜Pk��6q㖝>�d_�Q�>�ЗO��@v��03Qs��U$r.���#ԑ�O���)�~9�GCjÛE�gl�j��Sw�b���>]с���d:�A�� �0��U)��J��&A�5��w��
�O_��M��+��`j�IQ�5����u,�Vb���p��;^�%� ��@$��κs���[��B�i�A�����ӧ7�<p�"*�+����E�7����o�0
��y�!�J�5��>cʻ�6V3X���2�"c�Ī[�	X3i?��m�\?&��U
�f��}�8�XܰVe~y��p���'��'8��zKŠ3A!4���:�)f�RK�]��)�(f�U_�r�P���{4���J���+�{�'+:/��������n����yUr��8�.׾��4v��Jt�ş�CF �$��R�.�����Q��9��f��=�pnOet�v(�)��ष?�[)�g-��R��� �@S�����fUt;J����Y�����ޠ��/'�X�b꣟n���~�>��Q���M BC /��i
uɌ%'�&I����vg��As�b~Z��}�\�&�K_L5�/G���*��e����d]�����9¬`r�kR5��5h��Mt����k�yB)�@���Pع;���������V�������U�w�]wL�u���ɫ��}<��1r�I <��ː#&D�.��uM˲K�O���t�]�LV=�D�\��V�ƕM�����#|�p��■J�u��m#��Df��ݒD�:N�/*�N���d��v'���U<Eފ��z�lJ�;�>�y��`����j��U�j)`��)y�$����ou��R�f�ߏ�f�k�����wh͘���h*b���
3s�0��,ò���>"5_�'P%����?0N*WX�6y�|��q���V�l@�m�}�buK��W�#ӕd+1.+,�`���&�}��N,Nz���L!/){ބհ,��E�ȹ�ǹ�K<�'�*w�A���󠰿��8x���saq2MН����<)xe	�i�������pN�\D�;�و^+�vp �jtؕIT݆��9��P��'q@O�Ih^�ZWM�Z�z�+?���6첨Ga'"�zt��X�����v��%������p���7��Od����W�o��N����a`��o��ш��dj�G���.��$bN�5���b��;L���A{��&�O�ѹ2�^<�]��k貶�ą��/�D��	�M�P�Ƙ��㎏�E�[�g\dt3-���D�M���&����>Ҭ�ʅA�Me	����I�mx�Q�]�%����g�*���!FxQ��:Id2�����%�g��j���L}�^�Y�p��U�h[g938d������yo�ǣ,!}{�%�\��e@.E�۰k�D����x.��)�n�T����5��W+�0Zb��R��i��7*�T3��q��&� ��&`��L�Ǐw#�
)%��d|����"�s�ٽ�2hr-&ʷ�m�����$��HS0_[vZaC�� �-���@�.k��
�\�f��٫h����`����r騦��.հ���~�d�3��-GO��/�D�k`��B��-���r@$����.iˀ��6�ޝj�����l֟�߄�7M����p�_7@f�+�Y,V)p��l>��T?�x�� ډo˶H�yh�k��o�d ��
�D�QW�'��#��P����V��r�Kv|H����?����k��6��?
�
�gs!F���|�.��1:+�.g��z��P�jH%S��c��\?����{(��ҥ>4g�6H��C)|�	�R"����r��?���(CZ����~��1	U�����!je?*���r�u�=�/�و�tt�	� �KA�Z��I�ēh�-E�]i<����7�Հ/1lz>1�;�1��T�D]��r�ԩ|?��T�x�~qr2�Qh�ա�x�X����	6R��A����	��l���7�P,ꂁeW�܏�j
 �a���f�6�厂�3 Ņj��!�L&��GF渝J������/M=>�a�NR\��V��7�*nF�_2A�q��ޤ!q�ZN7����[���Z�l�H�n�b���)I6\ћp��,SH�#t���ZZ�?�W������L
����a[��fY�	f_�^��@�ȱ��7��q��4@\�72���=ٚ��_3t�#rcG
6W�$�`4i��F��'=e�7(kƿ��K5 դ0�Eʅn���="������I6�'���l6���n���t9�Nk A@?�W�V��Y���̿}��pf�|e�cU~ `D�!*eTB���0�IB!����a�Zm�;c�
��n{�My�{M�x|��Ͱ`"_�j�9� =� �m�͊��`��1?�a_G���'mc����`�Ew����Dtv��{}tx��z�݃su:o����������ʣ)>g#�b��aҍ�v�\XTg$��ک0�c�
�^|�K;��E0�:""�P{��7�u��h��d%W������}��^&d�I=�������o�:rϩLv�Co� 8}}ti��/K�w:Y����~��.-�?<���������3�ۧ5���K�,{����O*n�΀�h��f�����5�<�c�\����b��;*�v�#[�S2b��i��%�[�k�QuL�oU��(�3�En`��OX��XK2vo������	1Q/ֲ��)YI�8��=�*���t�o��5ԥ��/1��]���k�@Ȱ�e��6 ����7�=IQ�tA���}��W!Mol/����2�������s�.���u��lBp�y��nF��O�H��/�`K����.�N��e�F�n\~�u������4k�m��+�Gs���\h�p�]��b[IL����.��!�T�3��`�o6rA7�3xy�C�����������=jt�,�W�B��xŕ�`g�4�(!7���El��Ͱ�2�n~ ��1�~��['�cG���T����[�.,A�I#q���G�����<ešk������u-�p:P���A����eFȴ!���8U�P2\�܅��iW^��E������~�v���NgO��� �m;����>?�Y�gV�fM,n�V�O����<�9�~�跄�c7LI��ї �E��;�.�:���i����y��h�3+� sI�m*0��tq��.l���Ġnb{��;��Ik_����a�0Cg��71;M8l<�P?}p�f�mGT�$�_Zu@���`��t��WWN��F&��Iw�AL$2�QKB�>B�Jw�F&vg�?�Z���ɣ���{�e�a%e�#�J����,^:���n�xn��c�/��<"���)�E�g_�|�32E�x
�xU�bG��c��o�H�%�;m�	�����F�j�\bTRӣi���wb�K2��3\�q�;-NI��[�Iw.	d0���0�ԁ�*�xH��)�l���G*�Fzz���mO's%)�y��v��D_s�+M�a!��:�z(i%؏�o����U����Mn���"X��Mi�g���B�o�	�W&�y�m	����G�]��;�(���+�x�����
��"�`I�Af��؞SC���
aG���--�Q�94���ǭ>Rҽ��B+LRbN�1���j�0���"�������2F��v%��NB���JjX���u�g�و���%�X���C�rOV��5���D�>?+�/�(�J�{7A�# �,�\3݇r��a|f9>�{�"�i(�,�9�&�S�jXo��	E��]�$�8��ч�D1��["�%2�c���N�-����-	�C��3	��ƣ�$�ݜ!�'N�iN,�Q�_��V���7�j
���\�wrl'24Jq.n[]P���S�;��P��L�Z��yFJ�ߕ
%�E=��&�p�m�$��:Tj��J'��2���V�D����|y�N��k-�j�:K�b�ܒ]p�"F���u+m~y�w���X��ʭ+�T<�2�sw-�|�¶V��m����V�?����*�g�_ �G�k�@�b���Uv�+�>3��*�1��=�A�A���D	�#��zQ\�g�&A5y�Xb7P}~��:&$8~�bD��3/2t(�ϲ�O��:Y¿㢦u#(R(1��Ͽ ��+U��:i9R��١ڜ�6�"�D����q��Lݪw���+��J�M�Ma<:K$;��H��XJ��=g!���"�+�� ���9؃e�W�j��Xk�m/j�aQW����D�
�,��o�3଍�M�ַk�/l�FG�	�,���>�Գy�5�2?=�C0V/I�po�{q�����\�UBh�n�}����WG�)�Xd��	�<o
�L�R`P	���aqE��W�'��%|10cs��W��)K>����k��Or�RJX�6x5M�S��֋s�݄��ǁ��o�9�[�M��+w�O�+M�X���w+��7Pp��d0hx���\ɥ������I9|�����6?�u���h9{�T׍C>�'*d�5*]���J6t8	ǌ��,�/;B�˷��wp����)��2���_��fnQ�I��>/;�.b�j>���P����;��>R�(l�yy[tt�K���/�.$D�*��`��@0/姌�~b����x�v�L�A�'�L��J�B��������;BTxMmN^�����2��c0,)p��w'(p,�����֣4�GlaЦ�Z��P