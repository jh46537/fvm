��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"�.0�у��u���D��@��납\^*�Y��+:?Ăh�g�зdA�O�cjf2��1Jeq�ެ��²gj2��$�Z���k��>�=���ȸ	�~�,t�c i8b׎��$�<7]�,a��;'�c���D�~�9Wg"�zp ����$^1�{쩱�:�����/3�E�{@�P������b+��Ky҂J�F.�F8 3��F8�Z3��}|�3��������_K��K�*i*�j�:�r5Xp�� �>4�ɽ4Iu�bK��Sfm,'�^��#4���0<1������U?OܢY+މ]G������lU����)�.>���w�~�4��7���ȫ��V�]GE�+��(3`���D��Y5����{7i*2:���T~ο�ßy�x��9@��ͪc�'�s �2JX�ꘄ��	��s\WvW��{c����f8��Fu8٘Rm��mDprJH���Dcs�P�h"j5Ժ[��]�!�r�w�k��ބ���{�B�?��[�ӡ��az5i�'1s�:ϒ?]|AN��rkc�:���ނ�r�J�L�I�4Z���I�ﶸe}�[_:���5d���F�EZfO�(N��S}�_Y擅����[�@��|���U�5 82;��"����&�Y�.�)�y@�����&7�$�x"�����w@c_E2w��}4N�UӬ�ȵ�w�W_l�l�{���N�����]����<�[�����h^j�O�[�)9�� ���&0�k�Ux(���0e��}���{i�2k��5*X���T{:�0��;D��utF��t�N��Z}�~E��vt+3592ʩ`�Tm�U�^J_�2Nb�1���G�6c�^Q��5ޑ4���Hӂ��A���=	�ڝr3�`ibL��LЉ��4��"��q��;!��#+�I#a������d!F�
@�%�KX����❞�ƈ���di��%Q1}U�x��_���M�Z)YD���]�F�+]F����q�Q�5����$�l+$�.1��A�YĠN·���!������9g�Fԙ/��+�̔��N�L)xy�m6�l����!)�&$/2�֢�bA���/E���8�[^�H7���'H�as�}S�J�m�Q61R�+*���0$,"�ǥA�l�_�*�)�1�+ùn�0~d."k�7���&q�/w�"�M��:�qUF����l���ܹ���ȧky$�#W<|+�����G��;�߈"�2	��f�/N�ک֋��WNm7Y�?z�X���t ���I��fq��~���]��0�Qa� ,-J/��!4;�O%Ń!G(W˲5�Љ�*ҁ��բ�=�0"��v��QwrG�>�-'�k��R��GP���[""�z~_���rbW%F(� #	z�b�1l�z��@"�b`�da�@�٭�A�FNT�^�<���㖎߹{��������O�e�
N['�C�,���Q����9��R��+<�P��۞>,Ҏݰ����g�uZS�ż��g)k��_��3T�y�l(RoʗLl�w��!i��Ϟ���
#ϋ5#��rV��0� +�6=H���C�߅��<NԲ��.�w�8�'��8p(�W���*,��E���BC}ūY��ň?�~
�]g����р	_�]��Q䛖�Y@F�B?ǆ-0��7}&��7��6D_��]�jx'��Aӹ׽�h���p���](bC{s��\d�� y3�t7&?<0�[��h��d�V?��|�*B�}�;���)���%s`Pj��i/~��`���;��R�`����(��L�^d*�b���dZ�d���<�V�Xz� %����1���}HR�����˦�q=���B� b�o{̟�!���� �F��}�p���<�L�~�q���1��O��]���zb�bqB��a��=��)0@����aЕxsX�ci�S	��>8�����6�/T��n�$ʔ�)2�5�����ڳ�b��.��06�	$(ϊ@���X9��CT|#�.� cK���w�/}���k�����J5������ ��;�/�۱��U���Q�	]ץw��5Й���-��>l3]5&�93(�%r(BM*0D�i�����h`/`oG�Gї�:�Y��"������z���'oy
yņ����-(����=S��ss���o�������G^��4�h^e���f�8ѐ"]]����.K��F��[�ڡ��$�΋U�b�g�oO�H�:鍒�j�c���?�8����s��f�n��t�N�����-��:���q5����'ڽr_�x���٫�\A��l/p��Y��x�B�y��E���k�#]��`���q����nd�B�
�Ռտ�����ڌ���~I�h4q���b����@?���)�i�c=�J_5�;vt~����F�|��&ʶǌѨ���F������ye�1JƤ ��,�"�4qMK���h>���=��|�з�=&�oP$�Y����U�����\��0���N|�����5�v�i57��_;�%�2V����9ڼɌg(k
���D���.N �U?I��C����F��h�F��b�}��1��2��ٟ㚣#I���i_�'��͜>Tw����l\$o���&�����'AC&�
���(��w��=�`�B?c��������9���Ma�	)�p��ҔA��o���{�gv"\��Pjb���a��*/4b��M+���Q�2>!�(Ks�e�J�J<4�E�LB~l���_d�����"T��)T�&�i�ԽcQ:?�O��L��!���a���v���d�&:QE`�a�	�Re��j�6�� $L�F<���g��2&��T�2�̴'����}k���*x��r��w%!z�� �5^o�
=�0���
\�(��Y�"�ȅ�A���.����o�8������	 �M�m��$(�s�~�W��0���)���ܭw;"![�@�?~����#TlC��Z}�-�9��b�O�����L2����[�ڛ�3�*M��V��aF1L��4.���[�\��A7Sۮ�tu	;M`A%��
����k�i�%���&Y9��\�!-/��4�u���]���bc��kKj�}+�g���%�w(���]�97g��i:�.�E�o��8�8?̮'�.,TQy+ivn�Α��U�	)�3nV5��%v���σ�9f�3ޒ`g�C:%�8����q�ɣf��j1n�~�췣�R�������.�c"Xa���׶=.LH�M��� ��C3 �R�l���,إ$�X�9<�d��*���,lБEu����å�$�8@�H�#�Q���3�%�K�k|�&��~xĄ��1�Lw�C�0�"���p�O��|�yL�h�^�������Gq����ʆ� �q�5�u�|�NgJo�@��2�lE~���YoR�������(���O�HX���s�^�P�W��GB�o�]��#p�-��Hpn�/�u�𮯷����#�g����z�{��<�@�u�8l��M��ʇ��B�<o��beH���s��{r����uy�뿝Vn�9i�@[f$א��+�랤eF�&�r�N]*x��r2�����iY��y7�P�}B��p}�\]-7���,���Kڸȑ�)f���S��W�{G��#�c:	:1,���"���W����+��R�84 4��"ACL����U�^E^�)��� m�[�:�W�y�-Op%��5v4�!.	�s@�aF���֘uN�<)E��O/���;m�$c��+)�}�:��r@�ή��{*b�Ia�V�>�*�Ga��
zFBB*����6��
h}d�+�ܛ�K/6Ϝ�}���?¤��K�
�����f��d�T(5���s4��u-�o\
�5V�N>#.y�9O�������Qr+H�'�\1#���٪ݔs�W���i&�u����91��2��r�ɄԦ��~�h��ƥ���؞W���;���6%���U�W�(}3U���$OOJ���ac��q4>�J`*�������dT�9A��LQU���#)����W�n�DQr�i+^1�Rk9��	6��Z��ڸE�=����ʹ���2�ꩦ��@-Y"Ϣ�,���H��"i$i�Tn)j� ��Nn���W�j��sWA�-���`�
 ��##��?@�ho�v�I�511˘��J��kT��Υ��srA&k;)��Y���^�؅��v$jQ����p�B����g��f>v����gV"W��c�����3p��TJ�RV�mCJ�(��.=4a���1;5�7�76����<���Z�F�����5�m��e%y�+i�up���� �P�]Y�\5M�����^�r(���/�2ANK�Z?�r�m�o��:�TM�&�1D"��݄�
=�l�2�s�`�b><�V�,ڏ�.�s���\Qʽ�f.�u'���$B����\��'�H`����<4��x��C%�����سMA4Q�`����pa�W�̫"���d�z�X8������`����x�F�3�ʋ^/��MQL�tJ��޴y����&|��~y��|����n~��(�^iЂ	���2F��Eۂ��$���,p�c��&z���{�zƧU�?T��׺�Ϗ�C;�b!�|��:����H���myFc����?M�ћƟ�`�,�_�_��[ٴ'I�&<��s��s���d3A)���ƅT�4&�[�͐��FZ�]��f���꽺�"O�6�T��#��9��}�����,_A��?����h��|&%y��UF������)&v���;����rC��'�
3�!8��Q�����1�x�[�")�p�!C�0N�Y^�zz���ދ��\�4
�2���R�Ք����Q��X�>���-MH�K�= �D�M*C
�$CF������ �� �t^F&�ՋD�0��X����HfِJg�M�5���cᲅC-!p������S4�,�4|Q�8't�������%(ڮ� "��X��~ODe��h������GWNa��]�?ȋ�K����v|�\��UD�"��I�v^ q�0�G�M�|we�<܄���z��x�{h�#��x�w���~��<8V�����(D-��a����Fn���q"�(��K ���,�R�̝gY���g2��M�~����\oUBq�3���n"@
Y:�jO�`<r=0r�Y��M������6�-l��4aG��Tc��5�����	��\�Y��d6>��L^��7�b�E��_��>ߙ��n�U]���}��7�R�F3m���A��7�����?�g.9����������i�D,��o_p�R��x2N�1�
�3�_� ����r��\�}��<�r/<��+�-X�?\��᳧�Mhy2n�u�5N���6 )R�G��o&!y�A����O�ü]xJ�}o.ֽ�ҫfD8�����t�8@俻���=B�S�[�!<�p?��ڞ��q��I���Xʃh2�	�S-xN"���C�-0��r'Cjsڟ�S1��Zr, ȹ�?����Ҵq����JIFy���
J���f����F�:WVQ5|4��ʝ�5O�H_#����!B��~�8�*�	�Qr`���q�c��S�+����\��p��f�ux�,��px�v�j�m�3��K9�6�y�z_��cZ���4�c�|���w V�{���%1->b\uY��SkҜ�>3ܻ���w�������E��バ���w��C,ɳ�%>ӛֈS L��B���]���O��>���`"o�w�9dr�$�����h��,�a�q�S���7�����_Y�O`�p�B2��|Z1r�"X����H����)�⛬��-���iJ.�K>q��Ok�`�R:��8ǡ=��-���Si0���'���>��ʹǌ��>���vڻ<��9<�x'�C `4iO� е��UH)x���Q�wM�����沬W�"U�\��h� i�H������`��&��(��f�L ���a�]�߉_]�sDt��?����rqh�"6�s�,r���F}�4��/EQŕ���{vNy�v4��(�GN���K�+��0�#6� @��5��}��5���^�&:�.�NF!l"����7��f-<=�N�J PG3l���?�4�5Y����x�W�o[S����
�T}��|�o���J"셸�@iI��x7Z?�����dyȤ��@^(�wL��kH�A_��kOq]���A��d�U�ź��g������	���Q�� ���Í=��#������@J@���{�]� #��!��=�S=��O��O&��<0]@�jM�{��<_ԄH�����Gdy��Z��]ıYOz
=|�u<W9 ]�5���$�C���Qn3_RE4:�,�� I���~��h�5�8�����d���}�"9�>7��;�5�K���\+�m7TMW�5~��
 ��h�vKSOǎ+���*��k���uQE���\����.c�I(g��٬(�N���*�\�k��h������-���xvi��\"�~�ޅ��@�g�t�\V{D�V{/��"�bP�⏣f�ZI��IJH�
x"���NbKȍ��G\���.Oߚ���'5�0]z-]�Y����N{�C�Wv��2���Apf��j�'d`�ʣ�AhZ�K�S���l���'�|��V�g����t4d+[W9�6��f5�� ��@��a�ǌJ?B��ix�B�F���;_b��"9��Z~��sl\�|���''&���C+h^���e����xK$�4!���6)_��Z,6���Q�-N$J ��@���{��2���:��_�'��5'��,��%/(U��cQ�����^�X2I�g�����b�ߛ\\�j�-� ��Z��^X���Y3z��8�*��V"8��"�NX����\�Fu���7"_^�Z���8v]^��<r`�_��eVh%�1�U-�y�{�#��A�/�͈�ak��O���FnC���p%)���c(�L����b���^�/��@�,�;�iW���]�� t�]�\bJG��[E����ku