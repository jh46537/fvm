��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�I�X��a22}�<�����kp��z54���#{B�T�&�(J(�I�}������~�c��l���ċ��h�G������׉����?CH�Nm?�3�,���:
S�?_W?��	혤X{�R�=�FW��oh�,����{cW�F�1T�A�E���������y��q���~ޭe�L�37�gZ�lOEA͹Z�&!w�� ���B_ϫ��E�l��ɜA�Ƴa��%7�W�G�[f�pw��^e��Uu����h{б�D�%�j1�֌8�I;U�B� z��3�r<����kO��Ѯv@ c���CCi�1�KՇ�W@�,��:fQ�����MA�ş���W�i�����E�����DZ�Z�8�-�,�(�p��?2����sNH�����*ͼ��"7�3����f�פ� ��럮k#��ql�8�f����tt��� 6]����Hi�ђ�Dl�i���(��%i�C��$|�&E�v�L�,�u��$��f2�_�G�=�/d��w�@�>o��\lX�Wʀ����hN;)�x����������N!����h�&����Љ�$��B$�В�%@춛V<�������Y�S�)al��u�!�XZ���^N�$(��wiǴk\;�OX�w�� ��d辎v��	�{��P[w��i�ITXhs:w��fwХ+�[9tPI����`ĵ=�4e8leVcw���ֺ��R-WҪ -�ڏ7�sڪ����v�3�p��Ė�	�g5KK8R�vozǡ {.�|F��ڰJ��[9|81�/']E5��J`gh���O���(���0������R��ӭ¸� �gu��<MW�N�`��`��_��־�]� �NS�t���R9m4ď�@��h"�zB�#����v��r'(L��t1,e$gFp��A޵,a���	�K�Y��mq,	^��ee�d�^�r_�^[ �;C7B6[�mqKf��T��B�;YQ�6W�U��#���rp�}��|��FN��l?>L9yp�f��q7��2�Y#�Ti�Y��eC�6
�q��|�O��na	��n-��՛M�mE�$g�����؞���Ԅx�LwS���Ng������+�f6�6wW6�(7�%�=�`�8XK�]���f�8H\ �Me��������˱t��c�w�ZgWEq5�﫡�3��l����c��,����?���2Drnr*��3�Ӱ��Q�V����w�Z�w`y�+8T>,yC�=,ZS�o���Z�L��<�홺��#V}����E�q�+B��۪�Rh8���8D�&��+^��>[����-�8�_V�eL�}��ޝd���!�Sն�a׳������S��f�R:�]C_!��TJ�k}3�V��x��]�	�KQ���n^,=(r|���k`�����9P���;e-)���3%_���O���
u�KOת����&�;�������]�;Q �-נ�A=;�g߈W�,�h��DB8�=Վ����x����Q�ᒹ�{�B0�<h|&����{�I%�S/�k�7�7����r��S����m�d��>Ǵ��4D�g��]��i�HR�$�-�7N�L
P�Hfw�	GǼ���#f��sH����%�e�	���y���{�xW�\��k����' ��v�i�q�0���9�ΖbAH;�@�"�S��L3ϛ��������N����BP�S}��Q��d�JI�!��
L���K�����׸�bTy�VW�Xg����6��c_YM���qx���f�����RW� 2��6r�2	�v:(���J����������L����ZiΖ�E	и5�DE-8�|�0��R:�T������M">�u�O\K�f�-�n����Z�ú&��d�8�٠! hV�F�<}�r2��o����@UMw��7Г��A�GDI����B�F�����W�3�(a������h��Lݐ_�ѓ��}�3�e�:5�ٍj��q�'�_Xs�����������{��O��J�@+�Vr(^�H�p��!��F�(��eC� �?} ��po���f�G�@� f�ño!� �����ܡL:��i���B��'��֞��RQoHා>+B��u�H ��^���2�p����N��f���5Hd��PMb������(^#ө����=/C�c�h��/!/%�$��3��-pV�y���/D2�=�F,k�[�ty[#V�����F�`���o�HF)���m}� �qU�k�	�>G@�8�:�U<'>E�,J""]��w�����)P/=��t�ޞ�:`��~�+]�[�b��:43m�Ϟ�7't4A�f|6�_��Nr����|�n�Ϛ�4�����5@ݤ���o%��L��,��3��-n�����z�(�u9E�'�au�񛧧��.|��P�wwY���ޱ�=�rbH�<0[���
	��R��z������(�5��ձ����}�Ԝ/9��bd5iK
J��ש�)�=�Wц��կz]K=�/4���lk���
�X���b yr�K����x�������o��k������P�=O�з�ˠ�\��v�ȝ�fz��
S>(�{����"��=V8�<X��;:�b�֝�ۣ8�؜ߦLA�\D���{ǎ���y���Di�W�`�-g��Mp-J�GXG	߂�!8���Kh���|�-���w���f71����5g��j��0w8� ���GsG �UC����*���a�?E-C���-S�������(b�׶��t���e�OX���5]�����X0w��㯊�:k�i6�K��]�}�F�:pPG�c�Y�д�r���.���V��o�ն:���zo��&bPw�)��[���@�9����b�H��ʖ���E��	lJ�l_]"!p:���I5�>NX]�n��/�1�ʚ��G9��c'�B�le�d�q�\VR���'�#�0y#��rڢnQ�����1=��B4:�Qeu�-]|Lh�<�ꦷ T�D5|1��K3!<�'F׶JAY@Ւ�*f�PN$�i�Nc����}3\��T����%�
R��'�͝"�[*?R��p�I]A��r�����m�Rk�|�o�h�S�NJٚn=�*�<\l��`�Լ�����SJ�T�7P�Ì! ���d� ߏ����Þ�Kxyb�E��s�2Ա��S<^�L���L|�PNͣ�&<�9d/ha<��jd�v+TE��/�0ǡ���x��n�����|�����IEs��P�gHCjq`#��<4 EU:(^{�Es�tn��r��؞�5J��5�j6VI����/��~8��x�#}�#l�/���4�~�\���Lu`|0�i�K~����x�HB�/���U�K�J�Y��=�M!�j��������a�V���g|�%�]���ٍ�5���hk_�����0�x�O�]��m
�	�@J�)�zg�3*�Ѝ�>Ę����b��?�I�@v@|�b�+wp6����9�QC��Ղ����@q�d�|2��`��[�u�Cũ�ldb�:|(�$E���N���˶H�����ur� 72��`�=� �+�$�>���«���Z�n��=a�W	��$��#tH�Z�����W�0�7���Ɨ�k��S�C�j����k+��~uѹ��w����]�m�U�x�⇋7Nr-L��:�9��7�k�ِ!f��_��ב�`�[/�9HeY���Hk&�D���*�ϋ�qR�@�}��w�p����� �����#Ks��]ʆ�nlݒ�aR�6��ɐuS7ּ	�M~k*_��̸�2tp�Z�����?������.M1�������R�gGwa���$Q��+�5b8H��v�G�UJ�L����_N� ss���P[��#6*L��N��\�~龫:uaZ�	�-�'��t�ڋ��,��ϠI�8��f��6�$=zp&�щ��{�|��yN+�8 ��D1��W�5���'�����a=�j�̏{���c[�@!�����{|XA���^�\�ם�T��F3�͎�+0-8\������ѻe����'�p?�+�<�?�$NY*u坠#���i7�rr���ˇ���B����J�;���l(
�rʞ��ӳ'K����`=1��@
��4�@��TN���ZU�����J��
�:�$L�h��}�bi��ڱ�5YM�$���c'_,u*u^f�s{D"��2T��TB���f٨ɥ�Ţ9/��d�ä���-t&c�^n��ճ���E˦P���Xn�����jM��Ui���Y���߀���f��!z�gwn.�/�4u�j�i�Q�C�{�G�;,"����R���d� �r=5Z�������i�(��㡓 ��7Ա{p� k�5q5?٩*:@|#��"5ynK;�#'B��8�L��Z�N<蕲�$���!����w��Z���zd��z�!r�����C��b_χ ����'��%��֯i��9�u����9��~?Qø�/�gs����o7�kM�TIy�#ElDl�G�9���s8�C��h;�����=�ػ�U\\���I��+W��"�s�h�1��H^Ḗ���y�$)��z��֎	���2;��q�Y����T$��e��-����� Ӯ֩�rN���Ml��E����禡|�HYVe����Y�&�GE��K���h��t�o�x�S�2�+�����,%���G�#yCa��F ����5�8���!T�ߟ�
���Fݞ�%�/G��{�\
��JY��}���U�-���;�_.~�~���95�w���Y���˴VUkfIٲ-��r�=��U�>#���/���H�~�.RYo�� ��1v}5qȝV�\:�\&��?�S��"� ;2�Q��'˹�e��
��A��a�p�,N0a:m�l��$��6�b�6bni*����?�ױ/�#�a1��`��zm��N� Ɛ�Q�A�K�]���.1 U�o���.U��1�X��x�]n���GcP���> *?���4mU���*��B< H"t�u?����4
��2��4��(^�߁�iH4{���Á�`�Э�*����Y�8���֦@�y���Z+����'^���1Z��d����	�6����	Db[A����pf�c��;0��$S]�̸֨�O�2d����e�b�-����[Q�� ���~�uD�Ry��pKl�W�!�ԕ�>