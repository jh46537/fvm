��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{�e���Kb*Y���g@'^��?��_�c�/��o�a�����G���2�˰�:����P��e��	�!��'d9vR��ۺ;8İv�Pm�w�dM����Ə"z�p聾Q������5�)�RP�(ݫjꥦ�t�O)���
���LZ�\Հ���Z^����K���L���=8;�]��RX�5��]�lJ��Gl_��:�E��v��_^�rJ9��(�Jt��.��Ax ������^�"����Li����M�dk�W���7�67U%A��MI|�9X�/�1�!���wZ5e��x?~T�U�}�L�z�sڽޣI�1y��ԩ��P0j>��<���.��l8�a���	�����H���}��0%����K��nO��-}�[����NM����W�����	i����$C��n\��v�S��]�:E.ֿ�d��m;��>$w��;� 3������kSQ��e;Hwm��.8�>�G����q�x����͉��@�΀�~A�p���/'�:7-J\fՁ�t/�P�lQ�1H5|�do�O����c�9�t�!9F����%k��p7u#�~�\�*�!���5��\3�t�e��v�L�,+���#�K����Ib}TW�^���:�(�L}�	3;s�SQ\�k�.�	tpW�4�PE�0�qM���.�\ �~�]����X �n�ɢ(���� �W{�đ�=l�FT!\h=��hީ�E�{^|����]� ��*?;Ыg�����ɞ�Њ�q�|���\��F��;|D��S��e������~ybW���° ��M��^S�5��1��(|Ņ�&�$m]�S�U1����Jfu:h�m����2D}oU��QlZv�?.kq�?>׋Vu����Е�PqC�׃f�fאaD��gh�Y�H3�L�F�X��k(d��3:�'�yE�����3��S��Z�	�3�B>�:��Q�_\�� �(��չ_2�����-׹Dg*���ĻD5�j�R#���)�=��p��7��Ur3rwf�r����,z;2��%:���[�E�)`�Q���:�^�\���r�H90���7=�b��W~}@�;�����1A����r1�{%Ƕ�(���� YM�'y�FQ9A��������y��5	��]W&j)���ݕ�����ɜ�:��ٯ�H�e,��#lXշα�E��wֱ6p��������oZ��+�VJ��Jo���@��f��lbDs���"(��p��� 2��������Q)�k�nJ�x�˔Kq�5��ﭤn�dl��l�h}XA��0^�#���w�A�rM��;�?���!�e�Z���Yҷ��1�Z���_	2�BB���hTw�A�"P�p�x�o�6��ݙN~��������LO���VF��F�!���;��yP�d��@Ƽ�p�4�_��1Jً̿����G��Ul=�u�v�"�z��d��"X��⠼9�$j4����#��jʝY�o��عD�^��E�:*�Ć(���cH����DHv�{�tf�6����e�3���g�q�M.�5��Q�i0dY�o��Sg�sw�c��j�eȤ�*^�K�
��Y{̬Sشo��u=Y1��´�=����[w+�Å�Rψ�iANL�l�C$�����g�D�(wC�Ꮖ�w�7�}��jg�v�����J[~�m��S�0ʦ�����aٽ��J����D�"�!
))eOt��C��]��FoE~��%�؟>�q�Q8��nC�[�&����=��/)�i���n��nL���|�Py���sbI�f�)=a9'_����%W{��>���2��,��j���u�U&oZI�I_3
�F��כO��	��P/�̂�����������`�͆jx+P���k�O(�']������������4>������9�[�ihbQҒ@*XzFT���f�qL*���\{�CJ��Nn�RbBs ��ל��� Ҩ�c����0����蟳%	�s�[E |!�u�[z��=�[}�R��|C�1Rối%��bA^;U]4�W�I��@O�R&�yq��8+?�c��;���mQ�����Ѩ�1otr-b�Ӯf"$$�,���_�¦���t~�+��s�	�4�����|�&�Ƈ�
�]@}�P8"�g~�B�2���Gw����K��0RU��H0D�V���x�����WpQ�1�|�&�fa�'���髯>&�;kV�{�_�xG��u2hS�}َ A�'f��a���g��j*�AՌ�C�r3e���܋e�j��m�\ְ\�}V�%T��_�a�����	a�-��]�[k��}~��:4��W[7a��_��F�T���O,�J���ߡ��T��W=L�Φ���.�W���Yf!���&�K��Ù��h��ߣD�ZL�!ʙa����hs�</{9�w����Hgn��L u�ք��*z��GO(H03e��`�i��Ỵ�Cɺd�<���q'b|�.I��Q���SD�B�Mz��\#dE�fR�� w��1A�Z ��wk�/&����n�,7BAڋ"�>Fr^����aK7ø���"���#��y�K����0�,n��{CA��"��vj��1U>D6�-ǉ��6}_[i�HY�e��%�/Oɷe�Cq�N��d~��I�њ����!%;Z�rRL7���ȕp���\��8��2�.?��E��b��8<4Ӥ*9���@#�ߤ�E�s��R��}�F�)H��_���/b�.Sw�9!������ܲ���Aj��4��)O��ݔ ��Ɠ2JLڅ�K��{�=�R{]�sy;��\�;�)�.���q���.aO	����������ʻ���5�.�^X�k��#�VH/�K�����jCJR3���L ~�X�����t����G�j��)]m �$T��}QT��\#�\#UL#� �����)'����i���`E��� Tœ����O� Et���Hw��g0XWU��NӕR]/��Gt��+ՌTz�y�,u�~?5���M(��Qc�
8ȣ�*GD�jUl��)��{j���ԗ��slT\X�����m���V�cm�E���P�3@Ϻ3M�-�r�(�3��,ذ�ۋ���n���}]KơB��Z�y��h:��.�i�倜�&��]�SYG���`&sl��{{H÷4�r�Ӱ?FFW^��J^���ת�_u��E���?��vE����t�E�0�D�rQ���ڮ��c:迩�H�l1tc��K�8����cva��)M��݋ކn��q͎S)[�-�F�����$����\"3�W��"�#�呟|����5z���:AE��Y�ҿ�1V�d�@�~#>QJ��D5���_z�