��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�×M��������`�X⯰�]<h��� U���o`7Ɋx�!�g���I{H���f�����&1�+)��ڷ����m�/��(�+u@��K
"��?A���yt�tn��@<n>e�q'J1B$\�xG$Pp��(�n�����k���6��[�ھ���K7>wCHYܨY2�d9����\&���~
��z�0�P�`F�����lȭ����>s�jO�aߐ-��>h�Y�x?�p����m�$��l�|�,��*0�J)��$�PC)͜7Wߦ�K�"��i��j/��
�[���IKT&�B��rN��,��<3�FI��;�
�B��Nj�tO.�һ����s\-����3v�l�����Qc�+Q1r�0eP�Z���O���J��c���4�#�bO۟��3�!t��-�j
�~A�̀��e����wo�fͤ��U��P����X*LL`ɝK��4ˌ�s8Ļ)M����W3�*1��lSU�Pj9Uz)�؃���c@�,�2����WDAro�/>R@S��|g��b	v+B�ff �c���~,��ۆ'�?�5���.�yk8�k�IYݢF�x3�vW����g��a\�f'{���跋3'3���ô�� 1	a��fL��&3*"i�x�N�Xӡb�r)]!���Y��T=XQ��s�KUE�h̓��I&��N@R~&����W��ت� �Ä��[W(���p��B~���k���.$YO�H�;�LZ+��l�"�7���G�=v9"�X�/g�j豏H�	,�/�!�p�����	���?�'I����ƅ\�r4K�dB�������Ūa3Dp*3��+�3�Xly!��;�#�]��y�����G�Ąe�~R��F�f;�l:}m��7�i��C�M�k&g�G�@���@l`�1�do�����4oʩB{,�LD�x�4����Ҧ`ek&52A�֪��UM�*�������4i�%�o�FqB�ܦ�9�����x���0��K���	�ʑ9�M
�-�/�Jw�$��� ���;Ozj�U�&�f��	���Ų�-,h���|N�=��:n[��=F#�{S���6;i�I�wAθ���?@�3���hll��6(�U>3t���|�G��K) z��P�j�mlQ�=�e9ȗj訝5nx.�+ �ކ�r��cƣ:�@PP���>�R�љj)PR:\n9�Y�*���`����1� M,o�oJ�ԭ�Ӹh�D�I��g�(���7E��K���թ���>�M��R$�����W�	f��e3���X�i>$ʤn�b�L���]]}�M�Q�jA�w�ķof&�������σ`�-t�x��檟��!r�U�Dlv˶[g���ߦ<�����]���*Vu��ý�0���:��#i�R�>6p�h�<���6!4,��ǜ}__�2g����&Gc�]�#A���nǖ��I�_q̟�e�e��?��Q�T����1ȡ�-8p`�1��	>�kS
E�r�y$pQ�CYt9��o���/������r�p13��5ßY�:P�������?[-:�11b��R)ĝ�ӈ����1��V�k���k����yNH��7@�zVg�w�-gĺ���	դbI`NGDo���S�{��u��RO�_]���V�y���m��P?h{����B+a/�=9죾�/��]:܂������\��+�ӂM+C\�~t�S�%2^<��8*�.��Tior���{�Q�0,��PbE��^�ZN`��7B;-/�WcL�v�@g��=���/����L^��ۛ����QX{3��H��P���#�Co�S�ֹ�7T�N	�3O�ճ�Y��"�J�dzfx�t�=h$F�@�ybw�	MeGWK�8G���.�Hʉ��d��n�k$�vl�KP5��+��O���=f�,Sϒ���5�2��R/�V���]�zP8�N�?qUP��ǘ.��J3_&�_������clK�D��Iy%r�k>K�sY힦�#U�ң���Hf���@ӽ��=�H�k>����E�g��͜��E6��t#�U+gF���0զ�Ay�36As6.JU�Oyx��l�f���>�H��I3CZ��@�6�ʀ~�>Hl9&Ʋ<"Y��x�<���e7b�g���cOEџcL6J{�X����?�2Yʼo�s,�6�?P7mu�n4|��ȋ�6�(I�j6�|�>4��*;{��5y�W;����Tu�w�.'����؉ N��ͮՙ�?p��a-������_�Ѕ�W���Ӿ妗[�������]����,ײ��,�n��/Cz���ۈ5I��/$�,/��Ѿ��g�Nl��JQe�M���/��m���k���tϸϑKx֥_}��u���ci*x� �v�;����ywY��8���u>��i�ZV�-K���oi�]W���驡���v=Yq�Q��aS��d�R$N2�3���K��l���JE]�}�+#Z}�f�S	!��@I��~��XG�	����g .!yƵ��Z�c������)z���)5mE��:�D�:~\�
'���+�JU�x�dv(߳�[O�<k�/�Wf	��r 8��	���A>O�0��	��_���ݮˡ�a�!@�'�= ��Pe�M,�޴ܨ_������s6V<�c���y"�p�t�N�Ke���?|�|Y+:�,=O%\�R���D���!��P��g�ֶ��	+�!����g�nd�	�ϸġ(�(�/��M@�x+���ΛM �nʡ�t���� ���C���)�"�"���>���Ό�E�\�������J��P�[ə	�)�S`����P<������E��7�P��/Q5�rʑ�V��3s�2�!+�`c'���E �X2��x�7�� ]��9Uٯ�� �~���x6Aa�a����~�y��3՞�I4��Q�6����n�^�5:G�!!<8�FzH��BA�<[�k�N��Ո|��˜��q+;�ĭL�P��M6,��x��-�T�t�m�ȯ�P�^�O3xr�ɎUj~F�=��_���p
U,���虙����}+�@��,�k�_cYA�A��eF�-7����[w�VRd
?"�f�[����HV���>���~~$�̔�l��ֻ�����23&�*_V��S�N��C��w����P�.|b�	W��B�Q��F(���͓��(�`���h�����7���t �m1��LP(��f9������1�:�Rn�{�n���D�ymQ��t���V�֝)�_��@�x�~]���Օ�h��ϥ��3(�uKg���n�vBC�sL�F��������6�*5A�ۿ���W5T���UCJ�ɵ�p�*�%��F��X�ݼ1��08�9A��&{Q�!��[J��誁(P٬��k5���I	�ԓ� 冢2�s�B�p�F�O�[�����&׸EV�����ϔ'��[_2-C���y��ؙ��+�ʚӭ�O�.u���1��N�e��N{U^���۩i �l*%A����������X�}���D�m>󋤞ӏ�[�(r�z�T�8)� �b��/mx�7�30=�u�l�mn��(�0S�Ƒ��6n~��^$�r�P��b��W[*'��״ڎ���� ���>R[�r�*������:�2���o��Y��6�][O�,L��k� �{�M�CӤ]UO������S?��1�I_P�k�^:c*S6:��נV�M¤;�v9+�%�H6��X�ó���w�0/����Гk�(�ȗ�I
�Y֕k!�@�ق�-�(�	{\	�c$� X��؎�:���k�氢m�rkS�㕴G�E�`~�A�x��x9p����:V��rRMv�^����j^�ǈN���6{}�o����}�F<��b�M�/�&���:n\8��)�Y���V�
���4�^��!{6C`�3�	����q���?Q�v��D�f�W.xVs��)�R'��3HjQr����0f��|L6�ƍ[��#_q�����P	��'����m�̵>��<��ڗ��T��v�k����z���y��+�Q3^Fl���>m�rP����/Q�N*c3�a,�yH���5<z�}jX*��z���UM6pi�t�.����6(�%�B����_U�\�8�MY�b֯+[=�Oy�g_n%&���%��,��M�#g���hg��a�`"|�����]�t���e�q�\��=o
-��7.WWL�FdS(��M)�#?���D�qg/�&��qpFq��xBPn�>p�A�8c<�����ni1H���է�D���"ՎT ���2N͆�i���dGq�4���<:�	��[����"D���,�i8"��L�K��\���8�<MW��k.���I��Jсt��@��k2}�F�t�:�Ҙ�8͗��a��.�D8]����� �_�7������C��B�f�W^"�E�p�q<��k8�n��zs4ϳ*�N�q� �/�Cާ�������jH�0��/?��Ϩ���*`�cT�LvC<
E(l;Â�T�	��BG��s��^f`��s����o��3�^�T5�u{0ߛ���ӔD�+�ᥩ:�Me�H�����P^��
Ʃ!�O��Ճ����MU���^��qh��`�����[�6R�o(�E�|O���,���K�4�CGѺ�!N�Y}�dgt��)*;<�����~�&qQ�,�e�:�2� ր��K��ݷd.i9��c��݉\t�O���'9#莰�@�g6(�����3����ȏ�9���D��F`��0n��V;����V��$_�Au�j��SM
�F��.��Jy��ߴ�O5-_�a$�x�i6(�#$)�J
S�AsgZd��>-%js��իz�}�K7D�%&�����^lҰn�X��"$U�'w�|���u�x��X	���lƁ��ߡ�{�c����{Tcl�`gul�ّo�Q�xCեV��lkp���} L�������l[DOs��&r�]�lZ�\g�[I/��)��
���=&���Wb���Z=b�Md��]��e�(K�P'X���˂ػ+q�:3��]1�eo ��^u�k��_�ؿ�r�	IuU�|5N(wŉz*/�m�&D���Ϛ��q+"�9V�v�uj�9�`
��T���#䪷����G�:�a�80�}��u��*#����������`�b��D�~�g3;#b�l��|�9�G][<w�m�H���������t�>.-�`I�e��➝��-���׸ס���4F�#��z��H�͐�-�^]�-c1��5���k������>��+�^��&n��Q��m�گ��е�����%)�(s�U��Kc���&�va���t������y��7�G����j�4�Tȭ�bFS����q\�<���VzJ��s6���Q�y t�|�ÂH���@��̾3g���4ʦ�	yt���.|��B����!�?��\�D�T�=o�Yo��?L���$��}`�q�Ξ ����ݒ.N�Q �Թ�"��G�L�B��}J#�&k�����$���qk�VIȥ���4C��`s����Z7i0#Β��������v�ц	M�;!�l��MV�M���[B����ȩF�/ O��l8_�d���w-�P�g�>햏9�wi���t!֥��_��.<���ChS,�W�B�1