��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�Y�f�ʴ��d�m���8P&B�� �� R͝���c�	���)es"[��é�#�‍?t���4�5!S�TP��k�$��  ��y�྄ !��g�?_�'@��-;'
 �eǩ�7�?��8I�3dU�c�G����t���#���v2_Ջ�	�!K��B���W�n1���'ri�ꔹ��jz;ƷWq�kՂ��[)�:�kq���ǋ�h�섙VB�w4�e�9��[P�'��HU���H26�p<��i�x:s��Ο�K�|xD8�	�۱�L�.»Z2��J�8��,:ف��4�ʇT���5uBP�Q��C{�b���u�q"3�?�*�Ivր��q�Q(��g$@�z�]K}��CjI��^Mjm��(�݉�*Y���\�d���v:Q!�
��8���?i-(�uQ^�yX��N��ݰm�{JR��R��3t����Ri�����qZ�e����#��츸����QC�5'[qX����MJ �c��ʧȜ2Ҕ׋�Q�0������ӆ�ND �&�䀐=8�n�-d�;,U��hB��mp$qv���N��uEI�	�P&�fe��rݙ^^�cn=�]������!Ԡ|G<�Χ% 2<�$i��j6��i�:�������,څ����.0-�w����O�(�MFd_�{'1�_w��]��f��U�>ۧ7<i�O��6��¦n@)�����U�m~Z�n}F�ZzԶ���u���Xk��l]��)�	�2n�46O
�$���|*����^�GtoZe���{�$8	<�S���6���ө�_�ש�Ԯ�u`��b���Bh�֯XC1ps�l��AV�?�`֗�(m�<)Z�&3[b��.�M�j�LFa[�����l����R������� p$F�i I�zL8�>�^���UA�ڞ�~�s�o|�gU[��'`�f�M
ͳ��L
�h���Y^mg�5��3�P_��İ!i���,�\�`�F�,4�\K���f��Q�F���>ut�geVZ��*���?��eNz������q_�\}�o�	ۇǚ~N���z��uw$��9Gc�0Y�,3MY���wS�?�s��G Y�hY%��U�:�/���E4R��7&������ڶ�Ѷ�x��QR��Lۼ&�r;������P���V�򘭓pڍ��5 ��H������^��0����$W��"G

xi�3���_��X{�}G�#G��Ok�XT� ="v��O-l�(����\��l��	��G�P���L��}�����r�V)���0��Ɩ]����'7�k�!�̯ �r����lk��%>����/�5%�����2߷�7S�ʻO������Ԟ���OM)���z�4�Y~v�������MK};~�S]��O�C�����0�*g�m5Yo�O�q�O0����k�L�Lӂ��/�	�V*�.ߘ���1Dw�U��s��9�s�������Ci��m܎q��u:�$/��?����L��[lj6�����,�0��ߴjv��z6�ć�������A�x_v�1�5?��K����f�.
�2�9�+�#L�j�gIg��ז̹�<`���*Х�Ȓ�a��j:�*�6�_���5y��4��o^��"=�]Y65���8����0�2���VO`j�������T� ����C��i���h%��i>#�;�I���zKyu*7r�w�o�#JX��� ��7���n�L�F���Fͦٯ׊�3R.�#:塛��d�Z���ڜ��@~ ��U��I+{�.����A;E�P�Ǣ�`:�'Ŭ>����ᓒ�>����*��4��n�K;xU-������Е4�[��PEj2�|!a�,��]=�i`]fc�0�3�P#f�)#��#�.ٻ$�S�Ʋx�o����h�9�`��G�_����)��$�B@q�uy����b��:�3A��N���	Z����� wc(��)���9PA��q������B��+�rѧ��e��,��GV���r���ܛ��#��'�&j=Bn������˪�����2'�T8������OJɁc��>M/p3;;��Q&r
!1��],_��ÑbאA�k|���;%$���a�*jr�2 �6�Cm_�$���F������XK
I!V�g�/б}�sk0�����ԏ�!��l�����yԲ��7�:����ZM��9��W`C߷l�^�6�)0���6��l'1��;6Owƭs���ޗ �t�d��*�2���;qL���d#�_4x��R�:O��#_KZ��^`]��r�Y�l/ Y��#A��E����iN���,F{}^�������MWf����_�ob��cwOW�8��� �!�SpW��n�C�z��}ݯ���6]�"��o�+]4������SL/q�PuMȔ������Q8���A��F�9����B����<mX�T�73��lϝ̱��F�t���K�tራy{t�+��,��3>q��������<+i�"�R�	m����̜`�m�=��?��}nК���\8��Ӿ�tw �\���#�J!r��;gi aB��W�Ns�� 	(@e��8��\�BUߟ
��A���W3ȀF���+�6�8�`�RZzL�V4~|.y��G���8�y!<�H���������C��i9~�l܋�G#S�tCe2��X��Ⱥ�/�O�
ϱ8�/��~�P.��Z��-(����Zv��vѼ`�א\>�~T�Cd%\��Xm��Ȗ�t�фu�#�b)��7���]?v�WC~��h�����g*�~���J�[�W�L�m>|`�`��wF"˟�	Y��־��!�W�7Dsc������^���s	ۍ?��f! ���^����c�r�����x��:M`]���n��p%݄۞�����[�	z&��5G#��g�&��uv�¦�S�k�&V5j1b�6^#B-!��/S�pTO�ܸU
� Xx�ثC�%E��'��n����9}��oB���]�e�7�J1�����ٗ>S|E4"X���6/MY��@i*m�
9���rCݳ���]��2�!����Ɓ��RŚi�e�����d+~�#<f���a�ז���v�.��C�A���:$�4�m�H؅xKT�;������Ϩc�(�
�}�#fU6�X5�-s�!p�8����vA�n(e.'��L��{5��Z��`%����{�j��*#���%
_�	�/��WU܎̿P�=�;��4j+�rut��K���E���Arx���R��m�#���Q�J?U?��)2Tﬤ�Ij�9���G��nr9!M�6x�����[l1���n��8������s6W%�W�P��`�w��ƻ�\I�9����JL��?���]�͍)� ��&c�6>�����y�AΰA�n����A��S��)U��1��l�$L>�L�dě����3F4�o�=�c>b��<��f &�
�BH�P�t]���?���h�	��l�n���]�����i;���Z�nqLr�z�#F�g�p�)ʱi�Ybٮ�X�Q���?O<q�l�~n�6]���r(���Z������D�gI�;�73�)'�a�����'�匒J;����,�x[��%�q�;P'�uZ�f�w1�ND����&�j0�����G����D[�Sw�^D!M�4C�%����\��Eg�����u��b����q���S`�S�ӵhAt�0�%O����6�XN�n�ԓ���s='��9�㈱�Z!�]�y�?�\�~��tj��	�;m�U$�猻
���j��Ly!��� �;
. *)���BTy���_���فS���Vg;
ؽ�a�:�}�=�M57�φv�4sB>�R��r�?x�������*�EF5B-)��ή~���h�b4����<U��>�	�û�>P�s^���e�^���"4���}�!��*�ڕ'�>��>���ܵ{�Ɠ m���Դ{|�1�<�	�	ִ��.���b�m�l�0�BZtY�Ѽ�!p�j2ӪVim�����E��䏊��N�'�-��l�}1`��<����R2/��w�ˋ瑯��hLV���2���DX��;هqDq(�(Ѫ���O�6�2C����[��b���}5x^u�:�#I����fM6
J�
z[+�T�������-`O���V	dW� �-$�Vb4�ƾ��'�����j6r�o��p��<J��,�r%쩨���r�bC˱W�Pf|`#o�}�޺��ӳ+-)߬��-֖�r&2�`1Wy�^7p�;�}Zu��/3L0�2ΰ��$��_�iD�3M+��#MRA��Ũ��V�J��]v�h�~��:�}��K�����u��~�Ɣ.[�'����D��\�ߕ:��F���6����,9A�K��:qƪ|������_�A� �YM\Ug)qPc�)���vN ��w�u�C�a��oOQeDK(u�ڈ����'��m�������$b2��kRX�~�Ʃ�%��7Q�m��`��/Q%�>9N�D�`�y������a��Q��@�Fb9}�y�-� "�		�O���=�޷
����1_�I�}e�'h�!�����R0���
�"�qCgG�_��Ȣ�}�oL(d)�IⳈ��@�D�7�J~�8i�K5�>Ǝ�
tp��PS����y��3-���Is��Irqd��L�RK��~|�>���]�w�$��z�u�G�$~@�6�?�J2vL��>����2�h�d>�We=?���}� D8���|��k�na-BI;�\�s���"�D��⭨B?�0\�F$<�M�m�*,�b9���ҳۨU��35䬨k��1���o��*�pR ���e���c5��Y�/�}$FW@;�4�����[jz������yI��=.�6��s8
��}' ���HP2����ka�n�R�B��dSFdڊ���+^�*׍�/ٛ�F�^r��9%���c�
�E�'Y���XM;D��ʯ_�n���YF�ar��N������y�K�%,@,���1*_3�L&�#p{}��coX�ڏm`���t�J3U������.�wq���'�"���SoX�cOu��y�mo����O0c�[t�sy�R����K�5�+��*�)X��D�ǜe8�e 5�����c��I��YI[p"�(p+���36�kN�� �����	�a�.�/t�C.��R����]�$O���Y�-��������@�Q_��ܑ�v���.Qԯ�E��:^H�I�O�)dr[�
�O\& ���Obu��L�`��ٵ5EEЃ:v�Gǻ�T�>���#��Dfj0�洢5�7�S�/��D�`�^��
��n�֫��'�@�{��7�NY��v?�Q��Ǯ���$a �uU�W�K�p�3�$z�+�c�ϕ�b�U� E��{.�2
�ʝW�O�Uq"� �A6l!'l��ϸ