��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�c���G�J�,=N�{�P.�*�@�&��^[��Ԇ�Ă�#�a��� u!��;*ջ�2��n��:#7��l��8����k�D��"3rd+���]��*�a���7�a�W�Ce�L������ ��5u���#��)�g���=!5�g]4�y��t�/�Y��Kw"������u�J�M&
Rܾ�a=�;�D�.[9>��_2�j)���&��%O���b�R#([��%x�E��8[���i��xh Z�ulN�"m*��5ߡ��!���ʛ(k���=���&�}�n	�i��8�=�(=��>چ�����[��/��#�qĪ�7�������m�훓((IF�YZy�r�z}G,mJ��&���\�}ֲ�n��i���*u#R�c� �zP�Lr�U��]o���� J���Y�\�J��_ա叫�#�/��1��":0jO]�T�F~���?r�c$,����Ti�o^��f���eq�d��U[/���s������h~ߌ�o'�%v�j9���sY����2D� -�'%��Sn��x���}{<
��i���y�+N�i��.�w)B����&�`�ܜ�ۮdA��@���԰g�TF[ņ�Z�W�y��t�3�����jC��� �Ջ����4��S�/s�w�,��b��u�ƶ�>��ґtչ�J���F%��j���`���C�3	��@A�#��|���H�E̚n�s�ワ3.���lrӂ�|Q~�]��]�\!��F0�݁ʃ���Z5�;.Aw�� q���p� V�N#���m�R��6���~���R�t���[�0R�Z�aK&.�>����?f����!?��$:a'�/)�P�~w�@��z�G�g	9a�8�F�!Y����U6�<��#������ş�Y��Gٍ2-F0��eJ���XݓJ�a��dgT������� ��1�!z,�g�
�"��2��1�|�kOEV�TZ��e&S[��n�S��� �d@\�E�3����&w̜E����+^A�9,�)��������.T�^5N��8j��{:/����
�d^��U��N{�{��ҩ��I��Rǀ$Ɯ!�M�b!��~��
��Wy?�g�����[��)���lj]�.f�Q�������(AD"�d�*D5��v��rv��+����B���v��թ��� ��)���9�åCC�!��JfU�%�.1�`����nNf3�Ʉi�=���kH�� ���U��%`
e�R�} v�~Ǐ6��dq��wΤt���.υ���֣���gIM�B�r���I��|��]��0̾F����4r���>�������LS�.��@��NY\��`��d�jL�i��1^#^�d�i��~��NJ�c�VU�y`�*tċ�j9�	kQ<�K5��d�쁟��X�:��6��^}���y{�C��p�.Bi�(j���
,d\�ʏ�KL8� m���F��q\u �䵪��]�"a��~����rJ�*�k}�cy��>:z�5Γ!���?ܔ?vhb��]Qɍ�o�wBlii�}�`e�D>�:�y�rĂ�\�:qn���r��O�>
C�E��⪣���@|���ʎ�օ :���PZ>�~�@9�B�ި&��W�ϕΨc��;i��U@#]Mn�#[�	����&�e[����I\Ѣ��F�<�m��"�@>́����#�¹�߮�QĳT�����������C��̣��7��pL/u�Zvn�[��A�e���Ղ=���^�y{��4��������76
dm�z+!�����j?�퐣S�A��l�E�D�Ge��,4$�7w���2�k21b>&D��Z!�<Y�x���j�Iϯ��B@{d�vĆT���`���}~e�U�{�@�>	�`�{讋8P�@���7��:�u�6-�����y;���cO6֏��F3H��t�t��G�}Z#�שx 9"������՞�69\-^ӡ��R��'No#*P�ÎNOi8���)�!��J<4�]�u����������P'���Nz��L�?Q���ww�H0�E�(V�U�M���Ũnd,V�?d��%e������D%_��y\=����mT�������q�~0Zc~���p����(���I���<i�;s�Hfkx�PH��Š��J�� [�q����ڵUd�i�.f@vԠ�廤U6��`���ciZ�M-���H͢�2�@Kڗ~��?�w�rWV2uֳ�۹���ޢ�6��2�f#ˡ������TL�u7#���Ў./18���p�2!�O������LŚ��G��J{X���7}i~(�E�� �CR����_A�.�#?��,�3�g��m@�s���uNT�Ά	n��Ia}(�=c���/�C���FoiY���kS���>ں�/�[����I�Z �N�x(�/D���>��p����J�4�AKj<��.ը+n�E�<����M!��M!�U�Y�7%��
��t� ��r�𑺤=z?� ��J�����J4��)�N����)��G��=�{�h�u=��bAqڈ�w1$8��̲X�p�����R��X�
���p�z���{�.w
��ی�$�=��kgd�|V+_|G�-�ce��und�\H���+1���ww�!1<H�}�vf�EWd��i���=H�K�e�Sy��"� �Q㏘�T>z�I_ʽi���c�X�OP��`c��}y��/�����R�,aO���>> ezYu�GL��G%U�$BQ��7\px�Аra����_Z4z�j�b��{�ٱ���0���(�O,PF�q{I���*��d��f�2��7w���?���ZQ��0 �sJˏީRY���]e�&B|y��x�m�����*[m$��U��Z�$��Z޷���s	�5n6�'��1xӌ ������l��?�a�ݝt<����勊�1-�8�4�4P��vV6j����3�*�gw8��#�d�6�B��S���5�r�u@���{}���:ьü� ����0l ��p%�Y?�N]�]�
M�<�ȅ�I��)�)ې�v���!�.#��|���v�)�pZ�H:��<~n�u�WGe���W!�i.���B��_h���Ef��u���*�9��b�sn�Y���N6F�r�G��ؽ�K.�CťtЛ��4���F_sW���>��e ,�H�m�m�5��pF٤����$��0��6���e����wII��SP�pg����&���g�!&.��}�&� �-c7�{�8���@���k��9jdi���,���}���D�2a�����x~[���o���Ol���i�Oϻ8� e\}
k^(�7������?�͏Nr�31��5D[ط���Wi���Y�s(�8Of�
L�c'���U��O9������)x+|�O!NH�>U�rS� ���;7�a0�'�Մ�+�UX�px*�b�@
����"f��x�Ox��6�l�͊q&0H/4��y�#x�<�}�YK�6q2L�9ДƩ��v)b�?f��>'܆��X�9�us]�٘_�,��L��� ;�¸���#C!���4O\��j8��$����g��ݥ��W���X��G�q�o�l$��؁OM�ᢹ�fU�����X^}�`vj��7X���6@B��ԩr�������K�)�����%�gs��P�6�[����NG��dee��|� �/$�L�O0=��
���`f}��)�������嘅�>xڃ�������)���Wm�������+"�L�w|�d>����/����h@#��6�V��Fj��tɎ/qˊ�x46c�3׎�+�	j��s�"�3��Q�W��v�:�f�3��x�㱴�Ƈ�J`T@�O���#CI����x&�">��#�,��V&��덍���Ÿ�L�tF�����t�r�"x0W�ka��A��hJ<�%'�Ό�帉9o�	d5���j_�:w��sw,�B)t�g*���kFB��	[1?]�f���^/ 6� ��Lw d��݉�=zך��l��&!ė�����w|�&c��������l�c������h��
�t>����K3�/��}i�U�Y3;X�UjH$g��݆�Y�Z������-��5HФ�����O.�[�}�,�D��9.�K�Q,Dbl�nD�N5�+I�;18g�R��uov���Zv ]Uǹ$�!滃$�6|�����]N�̸mTPڔ3y
Rq5���/��������2>2���Ť����u20S+�hľ�̍����)w�$�w�ya�e�r�	,�����$&�p<�>

x�prI�p�u��H�J꾡Y���2�ӻw���E*-w��ԆM�1LjÎ?�v��k%p�����5&��T>74��T@�<5���Cy#����4�kZ�<��cI�S
e��R��.�1E���󶪨Q���Tc3Ls���� ���6�2胕�v����^f���XJ6q��>6��}�c�k��Ip�^n��̖���;	� ;��!���dωXZ)"��Fr�s��q�2�˷3�tN���L`Ȧ%��bj��H�1����4.�����{bb�Z�B����,�2���%�K�ZR�f!�;ĝ9� ���ω���"@�Br�W�v���8�B�6�80�����s3	ܜ�1�aqUm�-Ȟ"Z8:���"��C�z=?��*Lp���o����ɑ��#x�=wE	��?�ק��5��ό��J^�3���*�(��6��<�W�6U���6c
���[�7�9�����˻�{	?٤p-�"W&��m�yT7��i���\'�|�)�zZ����v\{�Ќ(N��O����vpRPļ��"O�	�����k��ZAY<��g�Ǖ1��r�Lk�/W�[j�֯g���)�B]5������R_�+^&J��3(��.jb�<K�q�H�x/�a����M2V\��#$z�X�!�w�C��юGt+k%/���B�5��TMڴ�P���*@���(��A{쓑;�1��Z���A|�c´�����q��7O����A쁄��`�qi���j��N�� v?9�����	~4MJ
{<�W����<\O�ŧ1�?V����H���M_7�v��Ż!qu)�o��a	���p�m$��iZ<�����36d��&�l(�sLE�Aٱ�x�@�מ6+�U+-J�~�Zʄ,'�Ju1���a�g�|T)�qw5B�!qR����W��r(+�d)�GP���ftU�5�V!��^�_CmZ[���0�<�ק�w�B����!s?n6���:��Wڐ�{�E��b=�`a���	�ږͅ��?�r_t��I�a�	F��Ђo}(�ס�j�Fq�� �sЄͷ��7�z�\�E�G�8�ٰd�X��u��$g�g�4��ٵ½�N�~2����l���$�/FA�C��SyF��0���p%���SMo�S�����W�r�+����B��g�7`K���o���׼�|k���"\)϶�V�{����Q(%��#$��sW��U��T*���P������pבՂ)�$�SVNJ�Ԡ݀��6q�����[�a��2����r�4�?��N䖪�¦�"�Ʋ�l|�0��I^MAR!YDX�/�)�>��R]������ kGʹ�9����D�!kf�!�A"p���a��4&n���ʌ�Y�A��f.��e:���nF&��\Z�\E�5q<\�� bC����$-�ĺu4�6�C6�^���˸^NS�dn�a�1�+�����ם�,N~&�>���^�>I���}����!k���R���XW�X���ŵ�� ��h�@ �\�gy7�{x�r�G��t�}�"z���s��c�:�6���5B�g��� �/�Y*ºqps�1�R ��ȝ���Ї:K��!�4}@�~?/S��q��n׾S�U�0]BzAݧlx��Fu�������s��p>�#v��"�0�X��hrr�~E��c�H"�p����G���̾���a��tC��b#r"�ڐ��&�����1�q�s_O���w*>{b1�}���˅1�:!�n��O�;t����Pk'�f�5�����/)ɟ.�����o���r*����g6��)@Q��P	��)b%q��5���u�:T��8�O#a�"t��L�S����}h�4�b�N2��Et�1SF9�knz��W��P���H��c�@�K��ӆ�*�O���t8�2I�d^!� �C�?�K.+�$�< '�w�!�grË��y�[J�����p�Z7z�9�m�:;��7n[`�C�j��pwO��j�<G"E6�ay7ȳ�1���V��`X�z�TAW�8:y��@��K�����OEΛ��H�O3	�ՉK�_�2�	�Ca�/��d�UNY��Rb������<$�����,W����T�ܧk٪�r��U����:�65rƊ�Y%2�O�0�D��mi8S�����#�f�|�g]N��S�����dj�}�2�$���a�����,��5�y���}L]����"0̷��B �Y�]k� ���^���8aj�"�I�S%�_`V��)������ƹ��#B�����3����|�?i�`��o��{!��ܚ��&�WG�ViHj�R([�;I��@?�����(%I���U�����[c��N՜�t��i����mF�m�<��<���!v�.��0{�m*��><�>�-|Qn��LT��JӦN��n�����G���IT����˖�dZ�	VC�V9l�F�u�I����J����n����FG�L�O����J��|%RYP�U#�&��P�: �8r��K���Nc
qOn���ٶ'q�m0�Zɛc��SV]�͌� �i"�n�dG����BT��-��w\6gaNvi�E����!�S�['��<�՟� !S�z�Gr2+�,ݏ|�ո��/��*¦Y^�[�:��^�`۴E�L?µ��nk\��[��E�����b;�ݰOY{jڏ�'���s��)��p���$�����'��ټ�7�K>GO���xĮ�Dm����'"���B��w�#SZ�=�TRa�5=l.�d�Y+o