��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�����M�+��P4��p�<�� ��L�F9H3�(���>�q=fd@g��������w�u���%/y1]��-�$vC�R$�S�<n4�h�RB��!�u��l;�uXk��#\���{+ !�4��r�����Yj|]�}��qZt/�}9����6�A�5�T߮q�H�7�YK��Y$S��(aZ�O}l�8�z%�&�k��o��sǑ9n��j���=tКU��Ke��{^���>�n;��<��h���+�6)�MT�e��/@u'�������9����1�����Al�!�������<8PΖ��� �)��_['mv�B`~m���~L���""���N�%<6�M�����i�?���Wjk�l�����8O�h�\�q3��%B�	8����T�n�w�`����R�^��]݇sΤ&�*]gv�-��Ȧ̢ԱVN�J0�Wȁ.>�i�Qx��X8̃��K%���u�V�ʋu*�G�]��HU{�6G��Ѡ��s�91U��b�'�`e�2����L�;^�����0~�h~C�$5e�h����q������CL���p�����b��4���e��ak7�c��r�����)�C�n��*���56�ȺPP�s�6|�B����H��؂���eR;l�ag��k�1��Mߨ#^�=�.@6�z �Ii��a�P�Z��k��y�6~�	p���Að��M�����/l,3|+��o&����XC
)L��(y�6j�S>���!@�=>������9���8Ѷ,�g�%��
L�R׷6D���I�}7AF�|y�y��Ui=��L�li&e�u�c�����+J��ۜ��PJ��{��)�h�������8v�?=�i�|
�\�~�"����<��\����������J�zAI��(p��4��i�jD
=�0�HZr^2�
���E�H��Zl�+ˮY<�p�6���5���.m�CPM�v��#%�3��/ӝv����=��� 4¥�l�;~*]WOk&R1�Z�����#��o��JSp�"��V�ٙ�̽�'��(���WuY���� F���+J�)s n�{�.91�9e,��XZ�̹��ɴ`�����f7 �|937/'$ ��υ)�a��ؚٺ��K��j�ʮ\C?&��{�D�����<G�Tm@fL�Ғ؊�X�c��:�)c�юDH(�&(Ǟx��Y�l��W)*y|����,-�;�D����>^SPGUq��Yc������=H"����Dj|��7�����r�Y���,�i��,���sX�zΌ����l)}�a�����<��:���n��HPp;1"��Y�@����Q�׺?��ؐ�-vN��Y@��-(UAD;������0A����[ё�I�p�(��M�y_���2X�u����CH2��f��%(���l��EO��%��I���>$�]�#�������X�+��)��+�Y�B>�A2y�����5�k�$� ߔ&�؉M1?y�J�	w�.vÆ�%&t{�~�-���"��ֆ���tT!�I�|i���'��e�ӝ���N'ޞ/�C �x�����i�[�����v5]R;Ȯ��&_6{�$s�F1�L�iD4��f������n�}��X<��.�w,�;(��ZvX�������n�M��o��5j�sG�����-��qk''�\���8��7���|c�����[].I�i[�tDt���.I�����K�[{�v�8��[�=n�\��ʬ_��!�t5˫�e��`.k~~H�0�������É>0]�x:j�Շ��� 4������ �Ja��_��;5To�a�]�	�}N�f8����^��1�L�ũU\sݳ!Tآ�n[�.�wZ^&`�L�[�l��n���Ó#~t�lkD���<z$)�{6�߫�S#ȥA0�z�^�z��Xfm��{a�� ���-���?�)����H�J���d]��>5~���(?�[��Cl,��k!�GL'���!/P�*�\��p��+Msq\��,��-Z�#��U��gN]��[�[����y���iD��L1�:"u�
�F����mȼ�wtȾt������c,�>HL��ʟ�LVb1G��b������l0��%��L�%�j�57P���.4��B� �ÿ��<�_�$Vs3R@9]�
Y\��qAR��q�9�S>g�Oq��p��x�zd�M�>i�:vg#��V� �+��7E�)�U1ͫs~0"�
�-םs�%d�5���ٲ��cҜ�o��j
��u��u\�����F�4�Z�,N�wV�����t���``��:�ر����S�V�=#�|��8�$y��QL���J~M0��A��7Xu9K�S��V{��1�R'D���eu0�x�f���qeC���w��ɔ�"����`%S) :���x�Y��@N�����A�ᚷ���="�����3 ��N%�z,��c:�e����}����iҪ�2H��;�Y�s&i�3�a ��2ވg=�QX����-z����HN�Jڼ+m���f7�>4�cۉ"�H�C�c����hkmcKְ�S%B�BT(�����l������
�9))�I�wH�|C?�+�g�H�6�U� j���|i��`%��S:ӐT+٘٦�QQj*.|�dK:��� �K,�"�/EU�������j��ˢ��t�B�ȗ��DV$���/���4�]�`�9�ī4�T���K��4#�9��%ޫ>l��QK�2�9*�;"�˩ੈ]j�0
�;ܶ?�g��h]�J $-O���M�U��ۣ�W���>t�����=���P�gJUv��p��c�y<Do��e`�TO�I�2�I���S� �CM��M�&}No4�(��p��k������1CH��&q[�t.�z����E�$�5�� k����L�yf�M��I�W��$������6�|�9�eCz��y�J���N���褃��cSI�8��[N-xe֧�
3�f\������{Ǉ�ݼ�:<qp�)���,S������z�����]�m�RDǋ4��Ȱ��������w��=$�6(�����~������d��P(�q��N���cI���=�EK�KL���n��k��:՜lܐ��l4�/�u[lm)W�@>�vu]7�%�\�ڽX'��R��:��/¥F�Ўf=N8�qm7Y��Qj��EmuA�[�¥�� v�>fF`����]��7#�OF5/$�r�p)׳�1��ʳ0VI�w7�ݰ��*�w�7�!^��S'�G��T4Z)��NE�ʶ��J{.�K���K������U޽lL��N�4�6�"���f0�ۊ�K,�7�ε��!�}�Oެ��l{��t��j�L�XԈL�t����}Ws�Zq��
�,Co ���UgK��u)~�H`O�}��\v�x�_��v,�'�F;g�/u�j�a�/U*��窒�����ۆ,�ٵ,]Y�4^�(�������6��J�e�w���tJc�y�\m�$��	��+^�w�E�(e�%�8�f�&�k򊸐��uj�xh�� 65��f=[q�"��uο�H�T�c��ϥ��7	p��`�L�:0��~m�<��
�*���:�����A����-��no�v
6�`��؊\'϶���(Xs\s��|໿	�S��Z�#GtO'u�)��F+����|qĞ"�]gM�8�-A��(�ż�cx��2�{v�>�o�s�o����:^�z0�]_�C>Q�$���i;쮂aR�!�_���m_nI�4������w��f�V����LF2r�5>[X�
X��d��Io����N�dD� tF8[٢x>���l�����be_(��(�����y��t�T�D�����th{DM2�vdVK��`��(�rzNP���w%J�`��kf:Z�;r���=��;Ɩ�3Ҷ����ih/"�ڴ��E@��L�d%d���M,,1�A͆~���S<�`��$���w��J�0��~�v�8��|����1N"��H�<�"��wX�&�9ci���+6֧��*l- �  ��w(L��N^Y
~)�����F��Ԭ^���8�F��@c�����J3���?M�)��K��K�2l�0Ĵ��sp�1�������םm��o��ͅ��O덮�L�Q`O��7�=1�Z�Ta0���:�l;/���p�`�gr�#�,�t	�b�d�i2����fx��.�lY��'��i�*4n�Tp7f�B~�.�F������|J$_PI���� ͤ57�Ǫ��]�K���L+�#���<,���TK��*�^��-.��˽�N7����!���Zv��1�9�����aML�C�΋�"����'��L�=�_,)�I� �d�S���6]��&x��:��y�V@��YIiFr�A����ĥo%@��##	6#ȣ)Lj���ȣ��]�soRk�Se��g\�t/w8a�3�H�������ˍ늖� �(�Y���pT���ݾ>U:-�X�KJӖ?�Qw ���C��MG"�
�(��I]�����,��>����\��`D���a�-���M��"*8��p�N�,��"s�*V�]�u"0[?�yk
��]�o1��O)I;�:}x��$��.߳�9@��Tj����tu}-.$Vt橃��T�H�+ժ�NTB\i�T#��^!�}2���.��A_?��4fr]�x��L~���@C�;"}Po$l��c:浨��
�����Ց&J�Χ�uw�(�Z!��sP]O_�vkPSQ�61Dw/!�ȳ���8R/ۏ?�狇wW���@m|��G���E��{�ٿD�W3-L4��& ����Y	��1�6Tm2�OJƴ''K(zx�Ǘ(Lp�g�?��%�cK���4B6T��4�>�J����e��m�`�=3r�Tr��N*�9^���M=`#�9S������KO���[�+�DQQ̡�S���x�hK�V�֞C�K@]�c�t�$`�b٣9������~�����0�2*�Q���^���sȜ�
�v�YƤ��Z|//�n.GqFҮ����n5 
7k!>���T�%�CE�`�*��n��0MX���yc�E�������l��S\���i���� �<�&��������_S��(�B�%V��N���_��	m����A�߮D�!�iC�]`�:�N���1��mU΋�]a�a�^��8�NI7�}�\r��G���KϺ�÷U[� �u?#�Rn(e	���Ç/XN{��vdV��m��yB�����_�=��+1��m���ղ���AF���ꇯ��S4=֎��w<�/P6�smw�1�6Ż�I����ɰ���6�!QO�r�0�q�Z!U9��>�Cy���M�A���륍�G�5qtV�x���!2�}�c� �e-N2P T��V�u�pn�Ny�hА�ŐaR��u�7W2�R��Il�W+���<Qh��Z��i��w�-�7[^`�(��`&�n��gJ�Zϵ=I�����XRU��NIO�ǲ�����袑|*��`�ra��,�����xn�d��Mt *:X���X������r��OВ>0�,�Ԟ�'��C �ט�F	�#��E;b�}��0�9����&�uPLH�5}4?BxЧ'���/��j6��
r�������UA-
�
m�HR�Q]EB#5r��;â�b�I�ڝ�1y��6��qYF�M=�p�/�ӗ���ZHw�������>nL����[JQo�2G1��5㩕'�o-��[8!x��%��|#G,ŹM( ����v*�h�DvU���B�>��Hl�23���bV��a��֞�jϖD)�j��'���īp�G���
{����|�v�c��
j��@H����$TG*Y^XV �M�\՚���9҂�*���������H����$�Iz$@#}]RX�.E(�3�0s_kN�-�������*�ʠİ�X)M㰍�H�o���Uc�y6L4 �!�Ѵ�)|2�C+���Ôt�Bl|\Wy-�%׿��y /r4S~r1HM�A>���B�U8�:s�̕90N? ���bjG�ș�T���Ў����T$���qCq�PG� %���O����������Z懐�SX^�Vg9XB��.vV��k��cK}�;Ǚ)�*5e�/�Y��%Liz>h�:h{�Z�$e :��i_�Zc$^Y��3V�,��g�;R}j <����I��*���2�6!��y��܉]~$�1�~�?�ؕ//z��Wۗ���f�J�p��\FX�z��|��D����0� ˴��Y��x�Ŗ�Ӛ*	м���)����&���r���^s�y��t@r�i��q�����4~rj��j�?��Vh�m����7ʆ�g� g% �ƙ
~�����A���}k ��`ܼ�Rx�V�8(�&��O�
]l�4�{M�S�����n~�����}����w��Ֆ��$�zt$"p�x��������O�UP�����[߱'��֌=$ʾf����R ��	eț���^��ĭ�B�� �{��8}'|�d�L��\Rւh��0��۽l�CЃ�ZG���fQ��J&,�gW�m�]!1����7�O���������E��TP�A+o��n�.b�G�Flo���4Jat�k��ç_&�w%�y�R�4���ⰷ"�"E�p�SB{x��j~t�,�Gq�X�봶`f��m�t]ӇYOI��u�OKT��jSr>�O�?�t�S ��p�1��/D�/)�,�\T�+���Zz,!�)٪��w�4��k�1oMj��h��J*'�.��+��ۘ�K��H�˅�P�2�L�H9�i��c@W0�ҭ^��l�<ϟ&�Yn�u@%�D��013��~/u��|tLIKZ�o�(r&��aC��;�c:g�(��� ޣpdk&�9�6==�L��� ��#������Xsi�C��+)�ee�W���[7���h�������p7xz�iU�vk����m9�so���$֢� �4}��I�H�E̔��@���ں)�*��R �֋�Y��ܶ���{]C<����%�}O�L��H{��������Abߐ���)�*���Z�j��y�)x_S���Ee���ly��.��{�'��%'��D��S�F�9�־���C4Ah&�9�A�@.s��)	aд��.���a�^ָcZ��bn�N�=������dv7�����d+&v�b��r�p� :�B�t3���л��<5���_���WjyzX�Q��i�Ip��{3��s"T���;�\��bf��35>H�*���[�'{��AO� c;�u�f	v��-��ȃ��!�w�Ey}�s�CL���u�/�l"���t���cӡ�簊۽[�঻�֍l��[�5|�K>#��W�$p~"�8�s��Յ¶p�P��n�� �&�q�/��k��* yU��)d4�x$��E%S�w�L�mI�|/1��ɕi~�JVnF-�� aX�;�&�?��<_�A�2cy��]*[�gW�h���[��7�v>�A��۝�xVw����ą�Ua��pe�����q�^J����W�i`��Zx�QŚ�װr'� �Է�N?�jb"��-��Eb
H�su~���n�;E�ĳf��0��8��[;yg�g����޴qP<V��Hዴ��MYAR8�+s�W�v����9X�e ��:h|3~����#]���ܜ�m�{d��v@��٨�3���|l���l6s�BH�&�;YK�O�P��D�ߌ��١��[��
y��pzˍi�b���.��H�,�q�{�ɹhn�/1�R�^�k�,8��o��������݄l�O(
�GeܠL���� [V�;[�t4(��ʅ�ۧ�:��^��Z�u�RU^\QC*���U/�E�C/|lŻ��虡T��Eբ�<�B��"Q�޾v� d�O	EjoB�K�僘��'_���]��I�����N��H�Ր���E���󐪶Gʏ uL��r5k�!����U�*bWn�%
\��i�H�~tsozK�R�1�f5����jcշx�0oЎ���jэ�������l7ލ��Zߘ� �U�Q�}\L��?�`�yx�"��t����)J=n舢|ʃ���FG��\���v�r�;!���%�.�RkNP^5V*�(�rN���KAtk�pn���Zw����g�Mxph�D+�`��ӪhP5��S���x:�w�V���ޠ4�����wrڱ�zf|x��
 `]�|u����E���� �]뾳�9����+*ب�"���Oi�:�̖���i������5���Q2�AaQ;�R����ݝk@d/uˊĢ�I2���e���G�H�6�4?��6�����I��
Ȓ��j��;$��d�V7ۆ��E�B���*�s� ��wEtv����{�gW	������edr��s��?F�� U�)iJ��D� �[q�>(��UT���cETM��,�.({�*�i�Y�FH"��(��-D0R����۲�::K侔pP�0@n��_�:�p�EO�f�L�=�1Ӊ�K�f��J5BE�6P�~9v�U/��}��� YbzP�|@��\{]�_�nH{�@S�Mߋ�G/H���<�|[�Q=<%�T.�ЪB'�@�Y&G��ш։��V�V��U�������O�i����W�,����Ϟ�h7T�ȃ�"��๟.�,�G����*w��Z��b {��8���>��_�bVy�j�o�G�E��8�s��Le�N%7�r
�Z�A6{����֊�f+$����5���C�FI��ļ` �����%a�� ��s��	�с>�[��e��*%:���MҊ=��W���lV�%���"��=\+�A���v�����x4V�����ՙ�Ce`@�1~g�oV�h�����S��t	N����/;"��G_��]8*����2�o02�J�1�4���^c���p%��̎�����'�)��k���6]�j9��)]�t����ؗ�]�2趰g�ġ]Ƽ����ы'=@�Pf���m~�u��oz6���CC͟u�g+S��H�ޟ���zV���a�^0bse�[c[�f@�a��L��&%���(�僤����o�f��u5u'�3��
D{����ޭ��M��F��Jj\��oںr9��,��p\�@?��l%��w���נ�|D���2&J�E���H��o[B��1�w����Mm�8��,���8�=܃�q�ҕz�'�[IB���9i5�*���{w+]cM�s��X#���*jz �� �R���]�,��z8���Н<�܈��':N0ɕ�5�F�RH�LXohW1�^2�B�'^�B��S�-��~�i���Λ�k�����l�q��?����H�߽��6P:n��6؋r�Q+c伂3�a|�N=�6<�]���YPB���
�KrM>v���J8OZ 5��젻��6�b�^W&Q�ӗ�羛�i�j��^�0�.Gc���g$�؜�U�����@q#rQ,{��� ��FW4z��G� �f�������/eOcX���`��!��gW��<�!��-g�ė`�.�j�]�煸)�i��<���<�B��E�⎑�|���Ʋ,"�x>�3�:l_м�ah��SR�8�t����^����
�4 z/X�[Bj��',���O.4��Y�%9�즮��w P$K~sD1Zix.RB='�+�2�I}O�{��#���T���n�	_�WR�t��Sڙc�A ��#ےi������QWu"��Z�P����f�2΀��.��������|E��.��v�<1��H��`p�At�\e�m�0��v���V�V0�KG�*70�sX2���4�6������$�R�tף���l7���-w���;Δ��\J�������?�N�>o�G�V���XB��d�؟`�O�`��4}ގ��X�6;!��)��s�1& �A�7�ï�)@�(.ql��R��ee�H:��2>l^·�o�r��g�}#9%�޼��\EH���%��>�e_o�C���y�-�P�%��p�Ed"\z���"��d_���S�EC�$��EK�r)�:��l��8&�� �K���g���<I Fk"^V�R!�q�hFA�ɎI#�oT��k�A	����!��a�!�/d!@��b�PE8��-���U�*��޵�h�<�U�� �x:8?%�g�S�b�����|�˭�T˒j����<`��{U��]B�~5ld�
��9���*k7��0V�5}�-W�.o��kR�֢r�97�!粵�`\Hm��������M".�S^�N�%D�C�;~�Q�맏�wW�3��F�Sh���E܂�^�w�t�M��zH��"�i����|5��ڼ�~�K�eeLjZ
����IK^4�� �$���Z
B+q�ب���m4�*����
+R��=���]�t�T�!�r7��i_	H(�Jn�5����8'�t=��6���`3�ȫ���X8MI+tU��Z�$��N^Wy]2�In��F؆����0N)���B���Nc�(����p��������Z=�q���4��@�&-`�V�9 
z�|���I�����ҕF�I��:�p³ը������ݓ+3�L*�(O��p�y��C���=�)����,�?����'�XuK!�JTf�z��F�>�*9�0��7�0A�c������`4�.ʁJ'����YP�1�<|9��Q�T��1��������P$m�����e�,:M)5���\uY.�>abp���#@�FX#������xA���]��DY��\��r g��Pze*�#������ca�P��u�!F�v�p�O��ƾ8Q��b �w�̚��#������l�u�-t��GK���3_�ը�\��O�^����������6�#�JMRTZXL�p���hS�=�hds�yɈӡO��m��;k�F�`mz\H�0�Xin}h�~���s�f��@��	�L}���{���E��L飺teA�:��OP��X���!�(���ӥy!	���pe�fX�P��b�)�e}��Fh�dB�i��C�݂�c�6�`��-M��ϵ�d�����'�,�v�\Ɗ|�*������ ~9���]��#x}�_>�x]��iM���͊=�z�Ci���i9���&����,�@ј�1��`VV6s���D�j>py7� ��)u���˔���g��Nys[��D�zn�aiR��K4����&C�#��Ҏ%�&�-���o]���v�h�dC� ��ar����}�8�J���to&���)���qwˮW���~��"�H+�X�̏�|����Q��k�����CkR�G�r:D��^�V� �tfA�<`���Z,�p2V�bϛ3&C$�c�� �.j�!	��s�1m��4s� t��ѡ�v��e46 ��_6֩̢-��|�Dm���
g؇�����k$�
�K�^bh��=�S��9���w���cm�}2Ӈh�N=�9Q�P��Z	 �o�*Ɖz�{�;�)�,�kFY����U(��J�8��q�ʜ��)e���D/��Գ�t 75����i;d�X{��R1<���1��N@C9��c�:ff�ǡ��&�ȴ8?�3T���XT���}�Z&;�/ƵV��:�U;�&�Ȗ�}M?t�A�j<a� �K�֫MM�={TL�>��N;ن�t�ݼJN�ɩ��R:=��
�[���_��u�s]��%5�Z���! ���0ތ97���Y1�l;:O�
�E,O��D�p�A���q�m�o�j��U-��c���/\B�����ҩA�E��@Ij�A�KD�5�aE�"u@���>���l�e�ڌaȋ�a>���UU�X�bui�AX�kp�0����H�U���Zz��e��S�5"����(Ӥ\��.���
�m�?���bl�&�R`'/R��˟5��g`a�1��'�dm�Fu��n��oa�}�k.�DG�}�l<��<���4�xY�'i��������`Q�]���j���Cy柣��/�o���U��=`xH$3��'΃�r�	:ۯ>�G��%����e�D>�Y�H!~ع[}.��I�������<�|�"�����ӑ�n�G���U�Y�7�ĩD��Qb��ҍ��[��}D�ʥG����L��>�)�}~�:���vh����<@�����	��Cq�;^D��x��t�<xO��9�L���z	c�B</<��({0�I�Quh�
ZNV��F�
���ԳG�)��̳P}����{W�(xh���Ƥ�z�K����q^O�����R��31�4�);{'�l͛�\m��n#�����d l-|�'m�N�s�m���e�Y�#)a��ۼ��<���^�Z�z�������P�
꘠���|m�Cf�򈞪ɐ�Ye?���+���-,�ɢ�x��I�tt������`�*�Zn��Ľ�d�� Z����	τ�<��	�$t0n�+N��p�K!�W�=�m�M���]tZ�v�G�⋁���6%�ܥ�v�2�G�s��$�}#�������-~�,1[�����q����C������(h}�,��61���l�A�1<W�$YbM�I��]�m�M���.:�(��Bԫd�T�(��pE��k��t��鴴�z�ݧA�ō��m���:��Ƒ��yc�VAqC���)q��-�u�w�.�zt�-$��ͩ���9��Ȼe����X#�(Q���4� �X�QY�����dl��^��[��f?�2
�����0� @3Ƒq
!�a�P>�m�T�-k���T�[���ߕU,E7���ǁ�����/�~�J�C]{�����q�i;�t0hi*2~�#�7��h.s�Uh�^��:P�:�}V�ba�H���pq�4�v�U�;P� �*���t�9h��`����EfF�@�%SPvů�KZzǬ P61ک��?���Ж���늂%Le��1|��D�;�u<��lD�ؠ��E6���Ȍ8�T���6=@�� *��mA�Yf��/�h�fGu|�]��q����Hʅ"��zHy��} ���@�ے��K��l7>�����Vi�F��#����:l�3�޵:3!��$��ߓ7�*�ͤA�"n�s�D,%XA�.U�r���W��#S9C{�|�������u@ga}\��I����j]�ڼH �d	���yd�`Q6�)
X�	�r��@�E�UsA�JZ��v�_�����eK�F��n��p���jd_a힥z��L��S����մ<��:z�n���|,��:����0͵��Vi�.�
-���+�riH3(8���x)ma�#.Tx���h��T���P!��G��ƶ6�1s�_r[@K�-:/]j08
�4��5�w��0�L�⟎� ���Z�/TO>?>+�^~�/n<O�_�:���b@F���G6�~S<{v9��.�s�x�@CA�ɀ�*u_�F�~թ��8�|3^Jb�{�O�^�	zsu%�{W���^9�fO�Ђ��_-%:�x��A>�p���8^Bt�	���c3^��6���\v��U�_%]�Ϸ�vط.Sh�P��\�
�ԾR�3�1�>�-~��{�k�D����������7���o� Q� �H8���+}g�s�T��F1;u'؇�2���ޭ˦��-����[�������)�/�v�a��׼NX	�V��<�D�v��O��SmV�P kӊ�Ȓ�`��u�S1��{(E�\&[Ғ���`��e�7�Kd��[�<��JD�7���n�pB׻N��r�v�sm�i�H]_�b1sD�iJ<�s�������`/�i�6�ڀC���v���}���7~��.���fD�-Z�5x��.u��ѹ��>�[MO�������["*~����+�Wd��w��|�"dЦ� �����d��Bݮp8�gJ�?��Zރ�\�D>'N������k�1�%J�ef;�T�q�?}U*����!�p9�¸W�Sz7Lb]���QuV�5s;�)�q`2�J�Ⱥc�пj�"iX>�����<�^�LI���Ig9<�Co���WەG��P�L]�M���w4�[��{�W�
=�ޞ�8���^� kǷ��Hӱ��_�K1�9��a �<��>�FB����Tʸ�ݫ��ҕ��Tj&���;&0���gj�M˵�h'�e�$+���!�����g[ц(q$�KRs�g�v��W�^��.�![h�q��S��o�X[�e7��%�'@!<�F������ ���(���H�K�J� aZ��s[���_��La졢m�DsK��/�yQɶ���rAJ���^�_zm�km�9�g���-��O�tO���/:��&f�z�T�Պ���Ǳ��ږ�M(����	/��8�`�|ȵ�>��d�C��Hm�W9�1��}��1��fM <�^�~jb}�O���Bʹ��I1��1<�! ψ��7��d,�ae���'۱ԱLG���\kp��2�
�J�	�/���͗V��=�b�h�����/���Fk�fm4�-q(GJ&d]��C�$L�Fi[�&���Y6Y�ОPM��gN�ƾ���268�m��gAg�T�G?V����E�12��A�߅%���4��(�<[���p���͎�S0�z,�@�8�3	��M��L�$��
}�ގA�~�aE��d�Z���PS�����.����\Q���u�N���t���Ϯ�X��d)�!��T��J�,��`�޸q���(�-9�5E�tFJ)a�=����� V>��y��8�6�@��y�u�}A���/%!�@�|y��1��`��	��r�?qs.ǯ�zv���B������[�!V�-���1���Á:ͨ��t���k�S1r�Sj �{Z��aA^�݋
�$�wa��o�7tZ����7��)���άU��\�):�Զ��+�V?(4(��wJ?���,^�-i�T/���S|�g�{*�6��D�=.D�L�tKS���>�x�?�q����/jA���a��VD��p��$<$����:�B��7�3��4��q�C�܆��fTj�9@��Ղ�n�E�V��2���?�÷l�z��u(Y\��mf���p&�yJ'��0	���D��ң�h���㡍�q&_�Ƣ�@��z<����Ϩ9^jB�V���l�z�_���;k �8P���e��T@i�m�^J�q���!*e(N@C�"`�MZ6�׹�j6�~���L�v������@�}L?��ZM�afovB*�L�TN�u��!�O����A���>\�;Jy=B�zߠ���T�D���bx�6i[
�V:����d��f1���?�;ϝ�E���� v�j׭Y5�{ob�Ev4Q;�71e'P���{�/^��7��mHa��7c|wi��. ��/v�ߋ!L��3AJ�Ν���P�:�r5T�4)�B���#���V�Y�Uy�f���j.m�C*�d�6�R'6F��p��@�� ������B �4"�tCz\��
�h��qL:L?f[������0Pfԧ���o@y�BQ��>�}�<�׾g�u��S��ʓ�yь�D��~6�P)<�?_*p�m�ǰ��4�Q�~��#5�m�(m� &�S�t�Fi�X���ti�j�C���J���N�'�U)��h����ޭ��CT�մe�_���afݨ�m�v1|�߿��=_����n��ƕ�u�;����m������3����
�{�Zvx�n�����	��:��f ��Y<�r�����`�*�,=���E���P{�xJ���2��z�!�B ���aa3gAƕ�+)�$��q�O���:}󶦓���>(;��]i�
��T�Ov$f����6���w��T�����m�b@���h�G[ʥ���q���	xB���y�rԈo�B����n:8l�S`R���n��c���R�Y����O���;F�t�˨��G��_�OF^��
-����ca���@3k��:u4d��S\,�|ގu���L-p�į�k��R1}j�/$��C�>�u�5[d�0�C�W�-�ȟ���_��Y��;��&�nǞ��߮Q�����E�>G�5��#!n��{<5�<�{�0I�w�r6,�3�HJҋm�"pKwȔ:�L7�3O�c��W�88�$qSӧqgΦ�SF<^�s3OU��S^˘(������!8j�ذc�!���cybj�m�G��?��7��xV!D��P�?ҍ��n�����i�PM���,��9ʎ���kw!��F:NS9��~���]���[��)�^w8���o~�"��!E�qx�(������ZT� h����]���xV+��r�tv��qo���X�����J<23�I���+{��	<�L㪄��3,Pݍ�o9_�G��⇩zR6�>�X��`��_��/JS(�=⍩ae��F{�8�W�� .�/5U � �(��4�m�U�л�����L��ڰ׬�N��#V�j�F���^\��4��A�QqB!�5G.��9�ҰsJ@�,��� >1�B��68�y��fa�J_d�n�M��m�~�K�?XG�j�Rjx���<^N3�8�.xMc�q�Ϲ_�|4�gy�bu� 2��w�*�+�� ����ѢN<;�4�
A����WžY������t9������D�����CC��!֢�c��r)���\\��9P��J\��e��,Ɏ�E�m,O��<��B�'��j�q�c�{rJƮ?W�d��=5Z�h|���s	p4�K�/�"��b3�n��8�y���S� �˯���C�%܋_�=� ���q
�e'�r�|P#Z��' �������pK����nl �BW�}f
��p
�?��M���� 5��V��o_��5�a��&����L������i}�@q)����@�Ý�?q�X�\W���u�R�@�[`ڈq�o'&�*��l$��ԚJH�x�
_����������t*H>���;���~��H}��o-8$�a�M#
>b��S���H8{�@_�iT�M�C�9
7ĳy�jNry�}��Ig>Ȳ��ǆS������XQ�/삨�qJ� ��Q?+9��;��{�׉�.��A��bI��t��B�T!m$�$��CiQ_g��uB�1U,�=O���Km ��	�E��ց�S��i��F��ɘ���r\�~8E��D�X�,'��KY�K'��O�}v�T�<�N��u9�Y�>�5��ۨ����W"���س�0��T�rW��K�85%��g��;�Ώ�w,ϣ"��>K!�S�&�r�b�T�o&�pw1N����=r>��9� �P�x�܏?�,{�.o)L�"u����j�������Yo��m��i������/�.�?((v�<��dC ���P�������c@ b�bHN��tyj<kJ;Tyؚ�]!����ZÔZd.x�����Q/�ߓA2�����`�7:b�m�{u��<5Om�,@�H���Ɗ uop3���@��*��f�עof���<$���T:�鷂��E�����O�`e@�74&�V���9kЦ��G]�%vF�>c����N�	Q:�C¬������Q",�؞ʣ����[v#P躊?nS�k����k�Wn5?<��֋(U*GY�Gۋ��̹����+���u�������kRq��Ĉ)�ٍ �$p���&M�L�7�\G<������V��Qgn9$��)4ݠ־�Q^�,�4���`���f61��6����FRBFj�ܝ��1���SIju��i���0�٨��b/����䓯�*�l�zr;�W9�������]H�BX�=��Wȧܾca%��[˞ب)��<�>���9�@�2���3���ޥ՟�l���s2lV�#0�I��������R�d�\0�� ����e�&)�F�~�ׄ��#T��$knr=	��"(��̤ҋ���l5R�Ӕ���.LU ������WvNs��݋T��G���I���#��T<j��
4OQ��M����3�6_�F��B�CS������|���uzv��S����*Y5��4SS&$�X��d8��F�%i@b\?+�CSh�s���5��C���S+�f+���~�x]��Q������@M�^Hb���G��ܱy�'K<�Af�WL�G�0׼�Fy/��0̏Me�$�z�p�#-�z�!rM��?�I
�'�t��`�ٔ����K6ϟ��3��.�"�s'�Y���ߵ��^�{,�_���=����2'ٓ��vM��%�"�Fa�C.&H�z��V��5�o�+>��O���l��TQFߚ���v����g.D��*����Z�3�}��]�$`i/�J*уJ�9��=����3���XmQ3~�OǫY�Y�$J��2�GE���X"�$�	{�3���1��h��\������M�n���{��C�"�[�cc���IQH(~�W�9��F��<�8��C��\ 1�aw����,���]�?E-�h/�H�i����:���R��qt���[a���LР[�~�5J��ƠFJ]�U� u�{fr��Mt"k��9�������w ��"������3L�U�䟮�uL
��� o�H!��.~��6dy�}�o1�Xv�N�;lϦ>A ��ȮۖbG�3�A,�<"q�����(R���U�S�*�.�p��b5�$����d
h �݅�}O�M��;�b�QN�+JC�trz�$���V�����
�_ͫM�-���o[�K
��^��Nz���Il�=2��ך>�\
���J!�"?[���{�]���(^�}n�H[�?��BT�-�|�LQu�A��;ƨ���!�N��s�$�=�m�����t�
vD��KV�o1=NyM 1�6��0��y'����� �j�H�_k�kqtD�����g��3��s��0/�@A�R��g}��b5e�j��[ۛU�)�2*t��A�7A��Q��U���al9L��vӌY�qq�O)��7�)E1�s��(��B�E�J���Y^T���Yլ��:��cϫ���@G��Љ�j���C¡��./K��,���-�tw&�S!7��q�^g�c"8��T��ݚD�0��m��	�s��rY�$����۵�	l���:8�GPM`������VJo6w�G�5=�/	�L�̶��11J[�p��Vd-�pVݵ	�w��S_���[x� &��K��FzM���޼醐�O`w�&y>��#�vk��~ߟ��%Io9�g��9�ل���<�^{�rU�;� my~2�>k[��������]�3�ݔg=-����-9��z�?�ES	�N��-����/K��gczJo
���3��4��n�92���>��z��.�vP5*5��8{������h`�/��p0���XA�����f;E�	��g=N�����0E��ݞ�c��[��ygѭ-(f�������~�X�� ��I��0�f�RECneH�h
�w�ӻ��.��
O���Z6�ܝzьhv���*# O�02`+���r�e4�ܛg�#O{,"N�P��
/@��O7�p|Z�b�,���^{L�y��L�_T��=v�����Y;8�H��Z8��ؐ��SH\����WZk���F���bb�/�9�j�9����Zȷ�Y��MP��#32w^n�,^ř1A>smh����$;����'�ʉ0L���#�
���ߴ$.?FO{�Hc� n�k��v=V�]Y�2�bU^M!�]�xfv$��K�����XT�kҼ2��w+d�Ģ0�48��J��N��7�u�
�������t�,CV��qN%�K�ڲX�	^��LD�Q!4jt ]����b�o���HJ�]��ĵ�A%I�f���$������s�t��u�飅J���e�%�L)Bk�A%�����i�Y���\>wH�f���g*���(aN��ꍬ%g�>'��y<���9�=�M��+�t����ǿh���'G��nGX�+���y�#�Z3;��D�p@u'�/vN�.�������_&�Vy�2U����*ڍ�魧P��|. �3�?�`-74M���D��P�w]��R�#(��"7z�s�C]���j�4TƮ��(���jl�ux�u��]��2P<�~T;�뱸\�p�*��w���&{*F�M�ݏ7Чu��qCjuK�k�̫��E����g��**pߥ w~;b*T��:��Z���G�[�x+�7R:-$Fa�<��]t�3%Ή���1�n�lҋ埂2�*B�o����ש;�d�N�"z���m��NZ b�z�z|S�sx$�-�~K[��i4�D�>�sV,ܑ�-�	����,֊FckW��|����K�ۀ}*:�� e�g�-`h�����k��	�,����42|g싗Kg��"U�3��JϢ:O�b�B�i���[�H�@U�KV ߫m��k ��i���7d4yoJF��P ˎ�{�<zI������i>���4Smij��Lk����g4[���ٜp�qɁT]R�n췋(	*���ZǢ<�����XrШ}},����HsR�G`����c[^�q�����<E{q��[%X��q��Bӆ�<�_^ٔ� ��`XH6�>�s��p�1i��/4L��\q�D<@�����a��m{�m��#Ty���1U�<���%n�릒&���-��z��j�z���u,(u@A�u?v2LL�-q��]N�Fj�"Ez�#������N��� )e� ƾ
�>@|<��+*�l7x�ִ!�����\c�&I���s*G��,P��Nűς����a���g��sa�EfM�&m�`�К�fT@�h@�0�|xɿ�ѧ���� �ߛ�nT��x�����5���W�}�j���s�AT��=�����2>݇��7�7����2J�#��L)_�d��1u��(��8�8�([�;I(��QO�;�6Y���{���,c�1W��0�ٱ	
=N���ܺH�)��o��=����p���?���x֚2Iy�����r����*���s���+����n�AW4�{���5ȢL�����h�0W��N�e:��x��]�w���N��9�
TLg"R�ǺΧ�}]5߱�u����d�k8l�@2�cr��9[�gK�Qe�|��-�w�Gy�eI5�]y녒��CxͲ��&<����+*XS�y<7����o�Y��R̆ݖ���AYZ���W�3���j���� x\��^M���>3z�����v)N5�e�������2�)}ܕ���H�h����f����1��(�(�=Ӯ4��C�`����DJԆ `Vv9�>;4�����K����P�����"
,��C�;Z����u킾�o&�2�����Er@�)9��7!�.��.d��{/aƙ��[�@/�mL�Z�/�?�W@!�v^�;�X�OCj��O>�Q#��WF{�K���O���P��65MK����R�pg�����5��7�@�{.����
�~ƕU���L>g���'O[�1�J X�S�cb�b*R�c��N�\`}V%5�!��NOm�WR����P�#��#1(��W.߉"�[�KL:�kb��c�'Ya�Zo0�5�pߝ?�aG�g��5�a,����}ڡ�k�� �Ux����J�˼>)�G�h� oy���'���K���G*��}�U�������c��;4�� U�;�z��`��55�
g����WJ�9��Ե{�3e��f]�ýU�5�vq�& 72ټQ6�		���םռ��b��_*bb`�~V�-�a8Q����0%�4;�1x!w��N�=9։lUfW�H�E� �����&&���TF����;�l��/y�Xo�(_<�����4�cY����-�*p�5'�v1LM�&�6f��a72[����,�@��X/�񫙔�;�<$�"��IU(��[%���]'U�7#����m*t��U9dT�`7�Qq"[R��*A෯�6d�دhE;h)���H��r�����m
5Т_�ɘ���ֿK���i������s1[gS�<��C�Ĳ�j��NB�fS�<�Xd�f�q��B���P�B����^�`�bsSd|�!��¾=9`ꂇOB#��K��Qϭ�p"Y�~厗:=��R�(�w*���S?j�㴫 �$yy��W��g]������²-��R/D��2*u�2��Z��˴��>(��n>�J��̩��"X�8V� 80���1%2%� C�&De���딱nڰ��A���c�S3l���y=�#�4�6�[5��o��n��	�h����h~���Ad_�i��k����%��&�9޴�,�)#��U���p���	�F:�@ږ�����h����s\��y�zє+S�F�O�4�5�� ��-�����c~��?��t�biw���c����Î@^&}��e6x�L}�.��~s���u��O2�8�p����̦�?(��[�1��q$�&i�N�����F�RO�	ЅG(`Oms[�����I;<y0Pd`�k�a��dE(�Y�o�V��K�]��ks��������pp�G�
�|����t��q3��c��𗁿�ԏ�����
�$�����pGQ��	�����li�
���1,+&j��~�z�(@np1��!���_��ֳ��Nњ��zU+��@��Ҙ���'ʂ:'l�#�*M@Ƙ��/>M*����v~eo���2� }Y�m�m�ԵY[B���A8�@� 4�8;�R�$;6�3+�SL+�4YG+�R��D����S�ɔ�Z]tLXD�'\��$�'W�$+008�wO��� ��<ڎ\#jU������g�[��o�En��,�������b |�ٺ[ �t�0�ߚ��ŕ�ɫ��G�v��ͶF�O�������b n2�&ٻy� �][#� ��/�w��bb��F�A������!b�S~�����r��@2���/����&N�	nσH�"
�Y)? M-,��H����))Y0��&.�r݋���AE�ʎ
Ị-V�67.7/���}X���#H����49IS�g�z��c�,���_�ϗ�ٛTqn����v��B��'/�),e�t�����-H��,Kg6�����F�.��~�q��mpͅ Gv�U(���CRd��&��x�� k��H�~���"F��T�I�����^���o�¢(x�TY����%s䘇f�9����|4ub� ��]��1��B�o��I��Q��#2�h�4�o�A?+eQѻ�� p��<�^�`��j�WRo"P�+n��r���ר�?�*�<;��:pZ����j)Q�=ī�����B��js�D�#{�
�	_�y�֧�/�vgM�`����y�SϾMWJ1�4���Ϋ@��@�o@54M,-��?�����M��t���>1����>J�O��u� N/,�t���V=��Y���ɗ~@bU�n' 	��F[��M��8���px����dC!��Ǽ�q�7y��g{��Q�-P?�ky�Tj&Q#�b�Edڎ�4-���E�b�b�i)8ӗ ��=L��<�S0Rh8
?�XI�2,خ�(�{C<I�W9e홐h���Vg�gxZq��u�\�%�5[�=RF�=��3|f�+�5�'��� �7	�,xo��D����rJT��ѩ�o��e)goR;������0B'mhc&�~�D��%4'G�7e�?�W�-�fZ�_��nmc@�9q��
�1�2Ѧ���3�U2��#������'GT-�c�cMƬyJ5�{��ĭ��]nuE�m�{�]7������"�a<��5������Y��l�O*���Y���Oin��1_����/��=�A��JW���ĻR�����}�Q�7���JyM=�X�#�����'*�T�:���U?��qMϖ���Q��茤.V��f�������r����H������2~���]���zI�8�xⲒ��u=R~��8��út�c0�0A1|�S>�u{��F���2�=�/�Խp�2��D�������:]�;3��ٿO|Q5��B��Jm�r��k��M�胁�%��ϣ�_��xqP�

��hh�2~�p4f���1=.~��_ˋ>]!�@�M��4�v��m�4�e��Jp�ɼhU�����5�B�v̍:&f �|�,�k�Se"�9ǌ�Z��e;n؝��]n�����6!�&h�xg���_�Ѡ�!�m���9m��;�#�t��?o�<����͑̓o��`�Hs�~f�L*e��G��HNt��ĝPQ��C��h��F�+�\�^�[��6&jϠCO�Q�nhu`�����3�{`x"��V���ޘ[&E�S�֞'�	��#\����ov��5p����ؐ��^�R#�*X��-�3u��n�eˢˌ�r@�����l=n^���'��.�E��&]����[	.��UY��S]Ϯ]ϵ���6.���ֺ��t�,a��ۜ��D�vo
�N�/ 9撦i�ċC*!�FtT��Q��,����{};�bl�ـH�	�>�2���A��[x2�<��e�0����xe*q��Q�Z��Յi���w�#�D��]#�G �̄�f*��"#��c��m�Z��f��X��Rsd̋�K���aj�*V�Js5V����&S�T�,i����F)���>O#ߤm�h�;���R��)������P=%[�0ƹ%�����~�����[,�&��Iff�c6����% )չu���=-V�E�u�/v��H��-nvѣ���ïK(��M��ݛ����dG����`1:���hc-,ʺ�(Eh���D��D����{)��*�I��QM�[���H�y��U���N�m��^�+]���Z�
g���]�V*�t�Z���P��p1>��n<f@�b �$���e+"be��N�U���:8���2�3����~��V6����M۱�14s�m!jʵCi6 �C)��� Y�rm�!??����@O�p~(�z�6�5*ٶD�tFfa�.��O�0jn��ڋ%e !/tE�ѭ����hg9]�,&�|����PK_Ѯ�	�sfzs!Xk#��l.YݵB+͟�'��p*'�,�Y���R@/�����y��5��x3�}�>��_7ݰ��.����`B%5���n�w�旼Y�	ޏ�'W�w4�.��/W�a���H��c�R.�a�O��*�O�u*膛�fF�+k�^�f*�9vݓy��ԑd]o]�����_����@/��\������#!|�u���rk�F�q�/�n8�\=���c�s�6�Q�>ꄠ��Mu������E[J��n��̝ܪ��J 3���o��C'	��O�|�����d�V����3���`��R��U�`\�$aEK;��f��W�	�.����P&Ɉ֯#ŲΩD��>	�i{��]��R�$������ݷ�$d"߀}}is몦�����bX%��2��n�y�n��7b�!����6�L��մ.ۇW��Ň�
�}�ND���6����I����p��n���[�RR�(�����n������ւ�ӳ�R�����a�ۜ��iޥ	�����@f�ҭ�Om�-�a���'f�	m�D~�V�
_�����Nh�@')�)�~����EL԰@E��)D�EG4H4����^HoI!��6,E�E{o��+�����WF �u�u�]ل�`��R�c�����
�O!�i{{tQ��7#��岙nXS��ό�z���s�_k& ��F9�pZ��Uew�gd��i��}<{M��Zӷ{ߘ�ɜ0�Pߦ��_��nz�˩��Y�8�uY�]M��iW�?��t��R&�mI��iq$U���X��J@�F�7�Ҳs�Z��y41NH<�ߞ:,��F��/ �5�Ϥe9�5Eh�*N�u��c��mH�&��iD��U��lE�ݞm
��F�祘Dfq5m�e���c8�'/��?�¤,���D`j�AH�A0�6i��O'�JY��#���\F�적�iOP6d[�dT�,��#�-D�>xm ��Q�$9�Gf��DAۯ�ɡ{ς�^���y��J����ߣ��Ғ���b<�EQ*��O�-�q��T	�eQ��`�2�GQ�M����q��,�u�W �A��D<�h���)A:ә���Ƨo3�'���]�@�'aco�ۛT-(ƭ�X�=��5�*8��#�Vt\�h�i�EMa�8��#��W�1�!�}4�_뷺d����?�@0�B'"J�+�w�E��`e�[H�!sWͥ���1�w�I>BחbB�9�Z��c��EHƲ��P�Kx�-&�����p�a��H���$G&\�w
y�s:������3��&IWs/Y>��2����Y4>μ���҃�KV�AZ���@�����3�0��-cn��8�4��n`���N�ܚ.p��5U����YW�o{�_y5����g��	����"=�ʂt��:��{�D�T�hQ=
^i�e��xXBhF���e�Q��nWi?�%�;���
�p�ˍ������Ʃ�"O^���^�$��w8i��?�A��u��j��&D]._D_(й  k��9Q��|��
�!H��7��ve;��ɖR���
ӑ�d��4���{�^�%�@���epP�퇽��GGD;6��v�]i@����.��P�m�X������S�B�=!\�����	 a���\��i9�Q�\7X�Ҁyj�~����١��e�� }g<Qn�zA��o��!�vg��l�1/�[n�1U�bK"F�d��|�oM�=�%�O&e�}��T���x^l��G]�J��+/��fi�@Fsr�:<�V�I�l]�u#.c$Ew���1Ǔ1ѫߏ�o��
'�D|A�? ��? K2_Rt��}���.���8�N2�����5i�K�0K'2��V��29G�+Im�DY~�Q:Wx�oZ�x �Jcׅ�ɜ�����364[L��<���d!�^kͽ^L��`��o)M���Y��
�~/���	�>+���������*LP��j�Շ)�&�V��t���>��㘎��jɬ�Xލ�-W�2�v?����Ǩ C�<��.:�=�~��b`R��v>�heb��T[�$V�~%��W�np��A#���=R�^J�+�s/���ȢY�:��C˦0�c+�S�����9���gޱ(�=�j��'�4eY�ȏB��V�L��+�Ms��W��i���L����6ٮ�kCJ���)t �%(m4�T����_#1{��롵���[^e���\z��~�P���x�,)������žl10�3ׁ���X�Ƙ����A'A�(�fH���O�mj��䩘B�k���[����߹��Kw\hZ35��*'��=sFL0��yqk�ľ&��>��|��W`NPK@�!$MD�N��y��ԁ+���h��[4S�۠I�3e���V�Ҵ�=��9f�a܂�g�7��#C���*\��k����V��o��__�|dt�H�"�7�������Xݍt��ܔ��Ωk
5��`�L����8�|2�&^�/W'$���ݖW�7�7���-�HO�4!O75�K����G���P���"�ۓ�H���=�C��j����q��.�M�����c����vC�3T[^:��,^����U���p����7���}v2�G��1���+^�*��, �M��m��{�_I����uR�0x���E��Me1����]jp�:�̉",�m����{�[����|BjK:̓&��v�� c��N{��.��PXӡ���?3��r�g�� f�3�qbO���I �$+ �1Jl�+�����nt�.��Y(9��b�%�(#��A�O@�@JD�����=PIR��D19[K����<���������"I���\M�P��׳<	�E2�~Z���W_h��ռ���x��V�J��[�)R9�
�|��Qg�Ԟ��/s�7�#ķX��W�Εc���:�.|B w���'\F�fM�!ު���[_���!����A�knE�5A/�!\���4����!Ց�,�9�W��ٞ�Wh�����'tߘpW����Hܴ���ZZz�~ʔY�j��ևU��Җ~:�4���Kh���:����Et�U��(�=��f���>��/I�9�'�|}�����z�`T���;����ܳ��X�e��+�����Ĩу��'C�Y���@��e���ѯ%���[!A����U<�N�G��@��}���+s�-x0����?pc��ݷK#A`��XMEV��4dnz�X-��H�|�\>��73K[Clv�Ϸ��@)��
YT4fxZ�+A�[EP&��wb��T��[��*�K��EHx����d�U+��@Z���7�<_��~�4q]b�N���ұ< d�$O�����m|mgP����4-n�ƠE3�!Q��k����3��t�m������'�[o���0�C�$����-"%�Ǡ�P�Tn��B2:Y^��g	�C��H�Nȫ��m�?D�P�v'g��*�l��,��j�i���4	P~[Q��کh���搆û8@I��H>ct�T�uh	M���e�^l�Q��I!|lH��_w�W��(N����~�G�Yܝ $c:�t�)ڮw��$�~�~7/�_�z���q�P��߹��t`��(~�;�c�C＄(��ܠ��G�fĹ�i�
5
�\p?d��E��2E܇{�[<�8�r�����i�+X�IHWL�z�8�ͬ���Y�cS���ݙ�����$�u��շJڶ�/��Dg���X��a3�l6Df� 2�����Eh�'�i�K�P�(����=����4>�sZ� �Y�ס�eq����!u0�c�֋"#1�Q|ѝ��l����
Q+���VY��%"a���m
�Xk`�+��55^����5��e��zd<���4�����q��!o��K�흓2�^�2�)W?bg�	l͉��]��'Dg�����t ����aW��2c⛊iD��f2�Ȍ7*����$)�t���O\���9R�2E��=��.3��̱�GK/�o������Y}���9@8��/LO�MJ����pR��B�dui/x2~\���������{���M����Au���Sl�E,�9y{O��3�|�|�jq;��ƻF7b���G�_g`bh�+�+�qM쐈
�AT�ȺTxI�D���U�eX�ld�<�	���Qj�\NvٌӅ��_��	�Z�Q�r>�X2~�����r6�''9���4!�=a�R��5�T��[n�K&8��_�MN>�qX6����EJ�7gVN#68�:��\fq�a�Ȭ���i�I;�y��A�UL��4���{f�Q��j�Z
ǟGp�w�
	t�����A]]��;�R��ΰ,�9kX��.��LgB��P��X�Y�ޔ�Zs\Z�Q������/������k�%y¾$�p_���!�CX���t�Lc���V�oyK�=��Js����q�E�!F��1����[7P��5{W����2$F�ˊ�cp�/z(JJ�/�ߦQ�$�fB	���ø����\۟�St!k�O9Q�;(FEż�X�iD��i`D��1��J]&�,�?��Y4�07�W���$�k� ����s����%6I���~���Dg����JgߕK}�T����!C:ʰ
vt"�>�B| ���l�.X�, ��>��:��;�VW�~jѸ�Ԟ��`�q�	��B2&ܼ[����k�8���g:&��ҩ 
���l8R݃���r�m�7�$n���<p���Pk��{���f�R[�����7�:(Q�q�ʓ�m���N�԰4G|�3�4p���pc�2�<���$��sUJ5����3#YTԌ�vCQ+��D^~d	m�%ď�L3.5t���h	9�8_}@R�|��e�~S\����=r�P`@���k�t6���9��7��t9.e��q�.�����/v���ʹ�H��N w������ܖ-
6�rGi�p���I~:��d�v]���N�M
�~�{�(?�|5�B�ijgpr3R'Q�����^�9i��+7?��RKl�)�4�˗S2sJ@�hV�{��/�!���Q!"�@��Z��٩=;$��b�#���1F�,%��6�li#L�}�����}Nyj��xՀ�m�ky������B�̎��,#B�ݩ�x�es���&�ث�~)0��?;�x9=�]��ÙR(�6u��Δ&�"p'b%��3�������f���'����XI콿�j�81�mYT>�L���Ru�:8'K�����x�{MT�;�����l�$���
�43��P�*�b���TC�M��!	?T�CY�G�!�#9=z�S!G}�>!.G�l��{�Z�Z ��_�\3)!�GQ{@�	�C��&��e6�L?�"�'�K8F��yo��<�y�V��h���s��+SE�U!����0?�'S�v��P!�L�n: b�tvω�%�7�A�K���E�^T���y--���=k�0{:�������eW���8*5%<�P�)���!ӄ�!��9��+�Y���z�C�-j�2:�d\����$s��s �߈��n�f|l�h������KӰTG8�`:F�|"�M^��>���7�b�ҽN��S�й���"@�u0�pS����8*���Er #�˦D<�U�B䲞-�4~�o�(Y
ҤTY�)�ל�t�|�{�x��Ǜ�	%eS�޹)4���%�9���]�pTo�(]�Fߕu��Lpnͩ��Ӥ`�&���I��(��	�罨�&����m6�̓_Ů���%!�ʐ���;�dġ�C�kƜJ&�c8+>w�p-jH��4[��, ��j*/[iM&{��P(�]��e~i��� A��*?�9���6��b1{aSLzk��b_-��HeN,������g�ܼ�\~���ռbf�1z�@�M���� dO��@��a�Dô��P��q�_�t\r�.!�:�{�D�u��������	�ie&��7W+� �L��0}�=1!'������)>�`�C����Z�_�W���A�;K94f![�2r1K��+�HgoT����o	��՗��0��&:)D&�H�Sׂ.	,��	���^W�	S��[45�E^8������8��$��6���J7�������u�ݵ2X�A$X�Ak�X�B�,ڨ����?�&�&���]����N�B���aew�(&+���w.����p�$�/y,���˓�蕬�����U2���� ����\#�:@pu�^m���\n�<��ӫ�9��0J��#]*����̿օ��S9ř��!z�"B=L D����O���d�G)�Z���PS��ql�|��"q��p۳ԥ�V-�S����ϣۥ�S�/����=�+{B����"�5�F� 8EV=Q��˃��4"��S�gTޭ�����+Glo�	��>&\�VbΪ�iӃХ�ԏ�+�ȼP����}���N�%EhJ��i��l���̗Ś� ّ;�M���hJI� 4��<���|�_���8��Sb�#�����F1�~��P�R/��QP0�Ņ9S(�JW#�_�)��Di�$!?Q�ˇ�"��(I"��&�y�ܣ$�)[ue���˵pN�o���4,vD���x� Z�F2�	�T$?sJ��Ge�潚r��Dӥ��T:��tL3�S�cn,��U�����e�#+�C�y�}�r��#\�Ϊ��"ix�: ���4
5�9�/Mgw��	�"H7�LE"���Xe�$��E'؉��o��58x�/�<ć?σ*p������woSQ1�`��T���qJ�n�*zVgR�)�u�ׯ���Z����'#�X���i��B��hO�q��y��hWG�XJ�n�ҕy��&:�84D��ԗ�����G�gm�[�sR�
p(�Z|l��"��U<�oq��k"d�2M �$w$�^�AY3�HyGC�C�ybe.���՟j�-�O�+��Ce��Z��&(��
J�pX"NG��"DlG-�r�� �A�]hh#�A)3�˪m1`���#t���bG����T��y?���"�t��LՓ*;�+2�pR���h�CSn2��,��C7�u�]xp\!;3q\	�!I��%���!��\~9�J2������[rl��i�c.-�tp����|Q�+�tp�����V
u�C��P�P�9O=����7b��}�u�a\v2�mXL	�Մ!�q�������Y���3�K3�u�L��;��kp�m"2�1	�sC~>�[�܂Q�_�D0�;��W�0H;e���x_0���-��N�)����΋62=�J��qò�� fJ������/.1F��M��;�Xu!K���W�;����Q�㪨cz�N`�z�� �	\%�.�>�r=��!����Żh�0��2(�^m�3-p��ZEܰ�򟃟������G#b��j�iSz��Etvs'�}�x�k��^�3We2�v�\M~SB����}('�+�@��]RIzə� @2�at����ok��R`�_@���˦q����	�?m�	�0Q2B�<���m�\p��ԡ7���D!0�6yK��Nu��M_P�~^�V�S�#A$��W�Gl��L�yr"�2��ҹ�e�HQ~��������W�:�u�P9�h�C�ö�!��=����sA�\��c
Qv7SgAv��թ%�VyT�Ç�6�O�ַW;�,7�n�#VoF`���k�T�<�-��T3��N�'~2����D��%�e��
[$ܸue+G�2=�ӓx����3d��ץ���M	xBT*4�K
VP��~]�M����cp�0x/D�1'����f��TAS�$>C�����*�|�#�� �5F���q̳b���O~W�lw�:ϓ��:C��RI�^�.��ebV�6o3tL�B���R���##sp�[|�6���ry�fo���9��Uܻr��֕r�ֵE�G��N��q�(y��۽�^Z��Vx�1Q��m���v�=�ϔ
.Rڢ2!��]�{4��*��VN�QB��U�Z�%�)z/��q/^i~��Wj��+P��óF�j���;�]_,��n��ӳYbvja%~J�������P��Y�%��f��9�O[�B��3ƙ,{��!+�<��<Ĺ���P�V�/%���P[�f�ڦ�%�L�w�j�^�!�O>�\��5�1��r��:|6��)ufޒ����'�1E���`ڿR�:��3�sT��V.rȩS��k�LG
�e#��e�:g��Ź�̔b�c�w��^+��GJ7��L�FSxw�hi�K�LT|��Y��,��C����f~{B�w�{@�t�����YX���J5��s�Jh�� B���  f��5��
�҂d�R%#*�\����-yZ�~�qu�ӏ���i�#mf�z����O��k3��Ä��¸�}��:�G���`v3�H��D�l-s��+q���+ �ޣ�mEX���=��d�;�)�$d2�yʟ���/
lz8���r�v�5�gs�����ӽA�%Ȫ^���VUk-���3�_+�%����.���͝�H�GD�ߒ�ʕ`�wd��c4�׃�oV�����<2?�}[X�����!E��+�\oB��<��d��
Hr��r�(�NT��U�|����jUE�*o���RY�Y���J��T�D��P�C�2��=�;:�oR�X�A�f�����h���9(�E9���	�Ω�s�1�]�<6�RJ��1Mk`$Ki��P��oഉ��x�H����]{�>с�Ln��Dg�qpd�
AYcFPf�B�Uǳ�ܠ�<k�&1�XN�z� ��}i�}S�>4�$�XeӬ~��$�R�?�|#c"�o#;�'gn�}̃�%6O���S��1^tPW<�v�M,9R������$��>7�����e�/S�� �
 �֪����;��]H�oTw��u�E���W���bk��P4����?��tyX��}�x�a��G����7G� ���U�r��T��# �38�&�Į�Q�b�.f�z�v-!1�*��^=�L�	��.���/�M� g��D�$���C���<�ԁg�^&�)|�3&��Z9�fͅ�ui�k�8�_�>]���ҍ�1�$*�|H�B5��e������>��n�_����+�}t�ΐ�������K�Aϓ4 �, �u�b�9=���J(�c$O����I��/���#S�|$�w'���_�G_��U  �Q��@�wk�p�A
|�a�=�،�A���p\q�mo�5=�}BZ3�����R���m'r����|��]d!��ԇ�L���qc>_�xd[���(�6�Du�,r3��e�7������ى���F�V5b�f�؈҂� F���c%�b�?��HM���T�W�TiQȄ��v�ڒt�a�Wm�:��orW�e�U����ln�W1�.dJ��w�MfL ɫ^
��6�J�#a	�<D���1����;���`�t����
���*4ނ�Y���}��|m���ۇ1l�)gL�en�(�Q�Ҙ�~e4�<�s�L�!�/!W��2zj����JPc�Z(�o	������j!�h�ru&���ᑵ5�X�y��1"|�@�3�65�P����=���3WK௩({�� qX�Hv�Yܩ�$y�]��� FQ��7z�ǭ,	a5cL��v�ڣ%�<�75�*��!��h�2mxI�
7-������� %�m��㼇>��Q�ߍ,�F��ʗ>������@���������I�(�NTsJ{p��}y����[��m{b�e�$��;X�H�j�R|*ZK��Yf�~O4��#����M!��\��?$xrL6��^�;I #�+�ӦmTf�m���<8�8~;��59
��c�A���s�-�;�T3�4Czw�2.ض� T>פ�d�@�����r)����˽(�'0Ѕl.����3#� ,����{�\7!BJ�|��Ffw��Wv����|gI����bLg]��-��QTƘ�O���\��-���N�G��Y��+�8-D��OlhX��J��{,=S~xO��
�50�,"_��S�b,ڝ�Y�=(>���a:�m��F@��{ܓ�۳vC�qU�N!�'T6]굋�ߒBH��M7BZ���L��h&��;�`���:��~�M�s����g�a�uɖ������@f��/!�=�k�'8R��ţlL^l�����[�G5��G�PI~p���_q�$�O0��iiM+����P��{��\4 ��E��D;�Uz���"Bd�������&e*j�Ү���)�8̗~��8��W7�!u���wLuS�ܡ��Y!��3�[�P��4û���t��6���Fq򲷠�&�ar���|���:>ȳ�����6^�f��N:���F!ȡw������e�
���LQ����"�[ʏpm�C$ �2�B���漭��[����y}��^��[���>U����$���[���q
o�:��9�slM]�[�EǄ��7��X[>B^y{
���!���-`�B�e�ٗy�J@�( ���:rd����Ȑ}4����vYl�������g�/Q��a�ǫ|�j���+�b�hD>�8�� .�>U�q�Qk�x������V�qrM���Ű���G ��_�<]�"�7����N��ݒ}�:���:9�Z��\! '�&���}{2�\'b�@,k0����f�Q�-�����6"������]�r�ב��hu����G�Ok��L�u�gE��z"t���^*�7�pM/w;�dw�x�%��.�;�-l�	PZ�_��aB�,�`��=_O]������JFNh�Teۗ>V�>|�"$���y�i�uŎg�[�Ǒ&���L�j�W=��Z�X��I����ټ^����l%��0��,����hѫ��sN����c��ݞ�_����UBǐ��N!n���j����*F�U�LM�`V$-a��r��J���p��>��p�^)��1g>�2����Xi�NY���G��KҰ�Fww�ֹ���4* {����lC�ָ��i�ki����Hʻgԋ95ț�PN�k�2L$Z��DŇ�$"�'��Ҧ3�F:)LH�A��U��j���Q6�ՍU�T%��>&��>%��;��}�Ƌ�e�ֻ�df)��t����ߚ�Q�!6y�v�J����i�!��az�b7���$�v��W�*g��	T���̙�O��1�aZQ^}�@�"��jԲ<���i����ʎL�pj��d��x3~X}�l����:�2��c�d�l���w��}6o.37덕E��A[F��<��qm^��y�2
��.�N���[wo��C-t���w����E�kٷ��� �vR�o1�ĶԎ�j4�To�V�z�=�9�k�$����]��7�8O!�5|=���F7	x�GA��[T���͸
iq�}����,�U	'2��:L]��{�� J�(�CO<VDh���"šq|�e��2j�V[���k��r����Nb�h8y>j�$�}g�)�XG@PC�ݐi��ܦ�� �}O�~��)�*<s�$�_�lQq8D����	Ef���-�N4��U9fp�\��X�0+�~�8RZ����v�T67�i�#�w�3��)[���s��@r���I<��p֯P�x%b��n>kܙ��yg�����$�����k�V�D��9�4��Ŏ5���#}�U��D\�D�Y���|ߊ_�#V�yx����Ftr��QP�.R����yz��_��J���@j��Aw"��Df��K�h��)��:�I�Q���MnW�1�9[;L�RƋ�w)ƽ����8�;��`��v��7�a���)-��ng��Rǈc̘�)*\8�2	vŚ�7�[R��H�ħ�]�8�"�꤫��
p�uwjǾ3>f�;�p���{���}������s0g���GOi��mP���U̴��.�Gg�ٜ�wi�l/�I�q!�'P�k��>�dѽ�:�`k��9E#�X^J�z�;zii�؈N�^�=#L[�|���Tǁ����(L"���3e�P-,�PK���C,OE��\�a+�<��	iXMK�V��򏆺g�!�}��ّ
\��7��Qi�PqH��d�f��R��Qv�
�2�޸��J�*�N��i}9������P����S\����$]Ӹ+�m���k$'Z�w>Cpg�;�dc�A\�j����s��4�h�*����1�������݀��uj��Ǘf�}�g��}%W��y����q#rN�k���Dib��*��~���ӟ��vA۷��$-w�Qg�ts�{І�]��V�X��6m�����c���u�
|c)�����y܆�60k���A��"�y]�R���q�NSw<z-jW��$�l����RѭY=��Z��CZ���}�5ŽMU�_g2���bBǖ
�}��ٶ|	�&��g�>A]hE��ZQ/����g�fR�� �U�Td"�ƢV�v�����)�އ�vu>���>�!QL|f:���i��損z�-��2�������P���al����:�%%Z�"�����z.zK )y�L�ڿDOw+��ln�v#��O�����[Xe\A�i!�YxvI�t�2	]uĸ>Ӑ7d(���J�[9��L1�4<������<'I����K<��M�VJ��5��c�m�3��Y��-�6�t��<&mԡzEc�R�@�^�Ixy<&�g������]��3��k��]�d���%6���~T�~��^����ebѓ_�	�N&0+�i���o�D���/^~�9�*m�'	���'K�������C��>餂��<��X�(V�mIQq���l�ǿ��c� �6"�wh~�w��Ԃ9y�i�l�7u$?����c��/���B�q����\��+m�ءE������:�H�l�6�l`���V���7�T�}�}���ʅ��2weqK��q��*�P	5�97mLʪ���}�Y㕤h�T�|3> �HC���E���=�L�IK�77T����F��7�_Y�0,��O@�1�\>��ٵ��	Ժ�Z�H�7�+y9��:-����@KEڒ�"��puLiu�FG4`\�z�7�aq��G�yK�H7@B�(�$~:�oʺU&}��ɸ���/E��[�MZ�����Z��f�=�.��0�����K�ũhG��g����� �d��E1{x�촽y�����_E9��L��k�S~u;�QՔZ~���v�z�
�r��Qy^̃��$2A̵`A�6<v��h����y�L�<f���l[>+��d��	|��7�`|e6��p��v9�t"�A�>)�S�,���;��v�`=�?��R+�!��G���4ߔ�
j�/�%��������?p<57�Q�v{���C��X8�[z���-�/Ю�΀�,���"5'��Q�������FN2�s�-�*��X�m�Yv�@>Z����{��e��)C0� kCg�^0��g6ۨ{$�>�lw�0	�L��
 ��R���O��*�kRC�Jy�ե~����������$/3�*�}m]0��#�s�T=U4|\���r`h��5c��!�9�`R|�$"���,��y���\�g�<���n*#'��Л�m�N
�b������1C<&#@w�qnu��+����H���|B�?|&B;'Dd9��|Mԇ�R��H�/������I�ز@��?^a?�f��o����N�銊#����-�Y�l^�N�tz��f��h�j&&��?��@R�����`�v�q%*X��c1v�Oѕ���>mכc\����.{t�*҆F��� [c����7����_C)�՛Lv*Ӌ�#�1�2\>�Wh�������_�=G����`6v�77��X`*ݯ���d�g�!ƃ��]�������N�R�c�A6����O� c�+f���`�Zk�#feML����EI]�du|�3�ҹ�G�v�>#�vd�N������k�Ώ)�O~���A��Xn���"��'�9X������DK����$�*]��8)
�a����m�7���n�,����P��}�.?��Rط�f�)*�2��0���*��o"m��ʊ�I].�*�
r���-y��T{�+��)d��Í��)S��9\A�i�,��+����fz�}��OoU�8�5�D��p���ہ\B�8ƠOl��6Ғۚ@P��]��:���n��%�3a��U>1�|�dF�)� �ݚ�@L.[f][�v�uc�t^c��$r�Dɹ~L�
�Vϔ?�o����L}�$L��a�OԆ��
˂ V[�H4l6tJy������A���ZŘ�Ͳŀf�f���񶁱F(XQQ|��_�%<C�"G�K�`����,xv���ñU��WU�`a�А/��V%��	�i7�����������?.?�՞L���0)Z� l�a��/���NϾ̜i����M���ԕ<��(W?�C�xt�	5�P#}-�,;֑��3��o1�`0C�&�^��tw�&����*���M�&�FC_���$·�N�����:���a�������9T	��~`���*dvwKv� ݡ�qv��e]p�4E⩓Z�p$��UnJ.��d�ar��E����w�S75K!%�5�~�ě;�`���5�.�E��Iš�I�<��:����5j���N�����)aH#~[�#V��:uhRRAol͸������MIvD�������(�v�7�ұ�M��4,V����1aܬ��P��|P.`C��×����1�&�:�~��V��Vl�z��F~i; ��\k�@ia��qwm�t�=��(�ϝ���8%��;��&銆CY�;V��{n��s�'ӞF_E]1E$B'��6�ӝ�-�}��m�\�"��_��a�P�`Cd�0?�:���ۣ*�*&�R4(��G���I�j�|��d�:��=���t���Z���Qr��k	ˑ���;�?�f�l�G�s^�AdY��>J@�ka���mH�{w�8_&�Z^�|!����;�~L���-ug�F�m� �^x�7��`�+i>����/�����"C`�cz�Q�J���ٗ�m��$Xܾ5����I���������x�Z��W���0�e�z)6����wPU����He��i�߮x���i_������ZR��6%Sq����v��b�����M�t�(��n���8a�2$d��NSzv@0w�u�����QҸ��0O
t�'.�O
ߦ�*���`����
1��_t��?��f��� �/���%���_�X\�6*b�]dJ"V��Z�A��6�(l��,��Bl,b�J�K�L���̔-mt���E�h��;�\�w/B_����L-B
��IXOJkJ��囘�0��5R�
c��]�H�mS�N	]!�ӧZ��қ�2�v��0u��<P%�G��ݥ	-���iֵ`i��
�;�j���Ɔ��Uķ�!��Dokl�/�� 4�?�ӻ@_$���D�=Ⴖ�[ZLk�(����C+���Yڄ�����|9��.�<)�
(=Xe���k��m���mŦ�>���Øڈߩ�.I���!�x��-_��P��^���[J.E���P�.����H��y�W ��d��)cl�Wb�;��8j��ջ@������K؏-����|U���V�7�%O��-��j_���:R#�!n�=A��Ya�p���_�`����'f���B��;�=.��xs%^B�r�-o��e�Z�����1��+�ފ����7�"�V?:��k���ñ����{퍊ij.�?$Ҭ ���S�T��C����C[*lnU&�����m$ώk�q��ml�>�����ė����Q��cLOF/�!��>-�î�l�2q��YS��$zǾIf�sgv1:#�Eg1I4������r���O褽�˷"H�U���Ph����5�<�7I5�2G���\�\b���kZ�������YW�����Gw�YK'1s�#��DM����D��*��x���^/�S����W0$�����zᒻr킺ZGש��0�q1r��J=M7��X晑{���>�h��1�A��V���+0�ϵ�zCz�f�5K �i��[�t_�[���2B��r�HJ�'�[�G����,��\�.G��خk��Y��k���nyg�u��Ϳ��aXb�m�'�}��`�2�'��m��^�V�V0��L�K4�f`j6����F]���a�Ͻَ^#%s�Ѽ���$� �D��0�9��"���&��Ы��..W�'Y;��{B���o�n?�����VXaJвƞT]<O�R4(Q�&�i�m����mo��,�	���'/�8v��k܈�@��X7'd�_A��wW������E����Ψ�=�L��!��b��)lS��S���A|��Q���ni��O���7��tr���u�s��bB���o~��l�Z�p��"�0�E�q�@��~����:A�Nձ���M���HB�����=��*F���[͖�`��9KK���HQ�z��`��LYj��5p�w�����zw��Ī�-���yVj�F��A�}�����&5i���i���~�"��?���2�h&7a�1dA���ciѪ��g�B��p2+b�_�>P��������'�>��D��k�������E�F:���.��v``B{ bZ��"�?P�M],]�[#�b&�l��1T��f<�|�mƮ�õhj� �mj�H�ps��$���<��dSns��i��2��z.�{F�uCƫ����׺�)`Dj�P��(:�Bfs��f�6��t�k@�Ҹ�nAܡh͠|/�'�ҿ�r�t)�QvP6K4a��;e(@���Tg��k��d����F�Zj��D�� �3F3['4��*�3�W]���ߟ,{�nq�M���O]#"N�!]2�t��Gb��'���>��Z�5K'bxb��`�"��)�
4��=�&C�� J���g���&O�����d�B�G�q�'&^uՁٛ���B�.�^3��h=zT3�S[`�����*S��|{Ili�O��%�5��"�Z����Z��w������H�����_�u��Ƿ+-Z��[��s�(BD�L���J� �C]��G���5��T�_��`�:&A��h4!����D�'���qm��5Id;�U�V�^Y3%��pd�U��oȖ�"1�{I��־a���I��fw����=*[;�1�R3���m���-O�b��q��n5�[[7MyyeB=�h�O�66!��$ܰt8K�[,���`/��ƀ��"&�w�s�B�-�O���ޡμ]١����g%i�jܱ�*��t
�3&�����R�˞�vm������O(:�ն��CA��j�p��e_�o�R�O(�n�hw�!-n�~��R(m6�+*
���r�K�޶��蔱E�O ӽ�o�ѳ���Tg��A�
�4�xըe��b#���an��j�#�asP�L ~e�K�OH)�s1������=�x����H�J��65ߩ�s�m���SU�wZ��5A�����a��Gz�s��Z=7E��5���ǿ6���C�ux�M*�N `In	�4��5=�%[,�����5����k%��!�)�U�r�Vg6��֜A��nn9�G�H���_~�?��{\d���U�̠�#�B�P� �i'���rE�������}PGԷSD�H��֕E[Tb��ʋx(h����Cu��9�e��"ЧhdV�&0�8x-P��s@��^,�4ׁ��5L)2�2��>!��H��$?Pb���-�os�P>.F��!c�urco�e�d�ŝ� #�#CP�`��&���()Êe(I�8�� �