��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ5,��kF��#��o`�Y�7W�?Z���;В�vm�
�ǡ�Zw�Nһ���띰"����H.���W,�ލ�¡mWA����EA>��;�JG���)�҆�xٱ����=޷�s�a�jӻQ	�ܿ�_l)�2�NW����xM]g���A�s ����S��u�Հ��Y�_�5)P��Cg�M�x|�P�.��u�p0��&H����I���\�zl�
D��vi���{�F��*�M�~~�?"2�2L�y�����2*�������9;:d�xw���r��)������12C9q��2�VwT{J�������l�Uc�+�����.�}�y'��5%�!"�uȩ�Nz�A�^�m��S�@S����l��㤐03BR+�[yA%��*x����R�=�ӎ�*"�a�ߝ�^�:��C����G�d�:����%P/`�MQ��\y�μ;N�x}�ڤL#x��\
����aMZ����Ӭ����KC�S�_;� - ��Lj��6X��4�^t}��~���&o"d��CQs�g����e�Շr�t	�E@�"��CX0�����%jW�ܞK
���p��ͪةGM��sCF�@1�lHa�m�zfe�\�c0'W�h� -��R�=š`��R�&�z�h*n_��c@�h�����șK!��G��Nc��B�y^�������S K����<+��CM�4��_V�
Del1�P��-�O�;��a3w`�����������k�hx7�q�����p�%�|�?����ҧ��c�U7�=�L���Syh�ۯș/T�/��%��6Q�\m�R�[�������DI���#��$�x?�[�P���֮����?����0Y���«\��..�=N�nr�Fa��J"
J߭�[��/4?# E�d�V`?v�.:��o��d��AF�ĸ�F��l�[_�I��c�Xg�vn:R�Z�������n���N�V1�=�M���:�\�V�40^���~P�c��>H�<R
倰��ʥ�c��K��rq�;m�Qb��hf47��-2��Ja�A$N���o�������p��	"�a���ɞ%�Fw�s���@!�Cr���7�'�|L7!�:�0�=L��^)zw���#&���)�.D�]������ȡX,e��Ҋ���my��x��t ~�f� ��q ��K{͓0���@�:�+�5_p~���y��ጀb�%�hS� ��2<ｸ ���n�^�l��x�8"������T���0����jK�N5�_%�-��0��1$N��2GɸGZ�Wk�7ay�&��a
3O�ĭ��uʝ��!k�(��>��D��7,;�m!�=�l�-pL��<�$�+���^$~�����|�֜m�.#��4YTTE\l�a�)��h4;�]�p��:ic�0�Ԅg�:{v�����D������ҧ���+P��7$�^|@�鿍 �?/�1�if�c�PW�i��0�����{�PPsB	����N�������E�!���+5S8��̓
��Y��f'�Gxdvo�H�����g���6�9ц`�������A����t�QǦ�)1õZ���ma)p#-!��L!��(���}9T4��ޫh�[�T��iX^l�`߀]�0x�R�V��ǚ6�3�S~��X�.^b��