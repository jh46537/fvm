��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨס�>�6a�
�Ys����'Gc�$��@	[��%EO��D/�ѯ�S�B���&Kc�:M��xD~@�����]B� �j2ʘU�������������v�oҸ����0Vk̃pW�#�}L���"�u��,L�92b#��mu&T�9;�O?݄-!\��T��m�6��L��o�o�Dɇʡ��\ƴ����q���S�q�,?�U?cgK| =S�2d�
м�6��+"t�M!%����*��e�R�;v6'�l�1��k��hDu�.�/5;T���ʣ�����8nAQ�Pf��&ֆ��V�9o�&[Rk4Ƃ;������Z��������z1���*GQ՞��Z��'���3�g��"����@ȝ��}��>Π��x�r��e��,�w��1�`�m}��5]���6K����T�����PV~�.����������[����!jd�����_�ao$�R���ٮ&��!�%�NS7��[ZNuh����@=d~% ׁ�8�sC+A�q$�Y	<�n�N�nLR�-`4]�$�Jiq��xo%���ּY��:2�=#A- �~�ѕ���:	�"f�����%�u��ᗽ�5�^�,Cv��k�0\���q��uu>(ԱDx)	�t�X@�cx��6A?�{E���/���k�S����tu��G��������Z}O�X$�߁ IKi���W<X�'��Je�4Ƚe����G�m�۷�9��w�ֹ
GR�5�W�P�q��(�)1k��ި��gɛ�c�E	5n���~e�>�z���/Ǜ8� q��މ�?�m oO.��ڊ܈O� �O��CW�n��\���b��X$�1'V{:߸ %�^��j�PG�"C���^��$�4A��׾I�����4���B���aX!�8�Q�t�֎�?u?gG[Z�i����ӯ��s�"�$x�]�[��s]�3>L^���A��z��)K/��#c�t�)&iF�������,[B�\|?�)���&�u�ў�^���q�<�<��k��!4��ꄻԍM2D�}�	�Z�;6�;6�C�oۮɼ��x������;LΤ��Ά;�a9�v	L�x˳w֛�]F�gF�{<_�9~+'Ł����tr&#d�`�>䆚���`u�탌`4��T����޷bERwʟv��#S��}��5d�Yy��b�ûIh������y�\{+EK�|>Z�x!���{�Ѻ��"�Ħfv����>�e'BI�F|���&��!U�Βs�ԯ��QK���b^dYi��n��������5�"���㤙���q��l��ղ���Oi�ݯ�%��*f[Z̆��*�?w��ق�h: e�G�b�@&/����(�0ě`�
�N��%����ֆ��
�2��Y�D`_��c��� �)��+~�i~�ދ���<���j6��fV�{}�����:z��\T��l��7�ëv��R�=��'
�Ɵ��8��^/Ǿ%[�~(A��d���\�ˋ����H��5��K� (dK՟�rJVX2Ԝ�
,�듏a?�]1V{�Y�~��L/(�J��YP�v7D���+U���("������g����c�%��9;����`u�&'�%�z�~s]�<��I�"Ĳ9��B쎣]��A�	m��FޢjW�R�@�w����黔4װ)=bq^��UF���@)�5���6��:��{�@�潄XE;l�Ә��M+%dS����︭^�-3x���a߯q�����]h�AY��D�U�5:�ocvF�ER���o�B��ц��nQ�Ov:��?����Ԧ��ܚr��yq����O&��ޞn!<���� B��n��.\Ġ�����:�mR�L[�kG�9�ӯ\�A�gqಮ�X82�-����^�\(_*Qo9�č�)]����o�6�H{��;��mU��k�y"	>i/Q����W*�e�:�"}0��Qu����Z�ZP�g@7�� "�k0���_��BƀP��a�2�j;�W'��N~�I�L�E��uf���q��;s�ƙ2)����~�`�y���1	Rҿ��[��u-a�9�}���|�y���ң��
�e!wݟA��͐���jۻ9��g����g�+l��qڞ��pJ���2K�7�{ �\��׺쨌K�����i}-�o��D>�r(���4�@o�nV�ң��V��C����b
�j
*LM�?���T�������g��MǞ����zdA����xe="(O���Ʃ�I��+@a��l�EȘ��x��݋x���]��-��@�O3�@28���~�C��/xv�_�����+�P��}^{���۽��WB(����#Du���K��|<P ��} ߕ�]�_��u/���BwV�����LC��"48�M@g5�U!��$�aJ�:�Gf�+�Ya �	���aSk�ꪶ�o�ԟt�WZ��|n�[�-�i�U8��q0@�t&_
ʒ�A�4
�����,�� ]NY�g��qy�'��/�e�܁�-�嗤���I:�#�\R��߿Mӷ�>�Ċ���������|�铚V2�� �)6�����������̇�rݧ]�w��]�|{��r�^�c{&�uyj�tRF���8G����^������o�(�����R5�2�2g�-��d�^��oaQv��iq5
��G��E��p���q�"j����7��\{b�� )��=�%ʪ�{g	�[���T��"^�V�,���0x�|����H�!��+�I�~w;]�. �+��M�};�:_7?����}Z�[q�Q)((��9i�Z,tW�n����wHN���~��`_�=�&(QL��Z��\[��MԪyA$�3g�O&W;�ueŚ
1�%6��{�D�0b��*`�D�n��+-�E����Y��xW��(B�A��F�������Ѝ����Fz47��N_�|_�0!��.��X�:��XﱯG����v��1�:90ap�V�Tc��-f�\b.,�2cg}�%MY.�o�;?�����=>��c�&�NOJK�M�}}�4u�+�YM�޳FH��R�@g<���Z2s���-�sm��ԩ��!�]$����;��;���(�3w�λ�"�үtsM[����0�[���*F_mޒ��J��'h�,l��Ⱐ1X�l�/���n�R-����6���ы�ڞ6��c���m[(���8��Elh5��$��H�o/�]��ޥ�סZ���3Ci@��~��)/&e�:���k�o+h��AVqL,Ɉ�*]��8MW-��R>tЧd.ke�$BVz#.����<�����V�g}zK�Ur����Ҭ���Կ�鲏�E�w2�0�tԱ4G�q�tJ|�i1�I��P��q�{�������b�D��aV����9��{C�$�v�ޛ��۰mR��U�Q�+°>n��k�KUw9���o=	�@ՠ��:_Lg����q�Ɔ@�ʋ\�r+yi����'k�����9Z����,���:"���k��-���H���߶�,����s��s�������dg�.l��;��0�����k���u��2횝�j�YM�bi�l��T�+`;�J2wo���,7�WdI��i��3�M��t4���e�Q�Y`����Ӂ��e�n6Dz�l�-���/��'V%#{'��ˇD�E}����A�x��ՙ(@��o~_o�Q����JXU��TU���*ȕ��j�u�����r{hމ��#��,[,O��]�����l�*�Q*�@�xj�I.����r4��xe~lԉ��8�nl<Б? �Y�@b��w���(�18r�ӣaN�Og���"�<O�i��k.g�<7W�1=�]@���y����ª�F�~*�b�g��A^4�^�䎃L���&�k�2�`�'��Mj!U�G�Xrw���uF���R����Oa`�G�͒���ͫ�Y�;?g��w�n����=�e��Rw� ��H��Ds)9{�~ tk�j�{��	=5�uj�\�jH���{�h���b���0��s/�Y�<��דX��o��H��Oåzߴ��lxs���
y��U�;F?��Ζ+0���b����pl�T�!9&��B�/���Y�<V�c];���I9��r�f�j�ld��2����8�b���2�۝z�$�������b�����X[?l��_8u���3;�r���=p�Ly���q\փfSH�X�Q=�wZ����J��0+ENT�{E�'��l������Ĝ���.�a
�J���X`( \�C��1�)��1B��e��O��?�L��KJ��ꮋ7��T��E-`��o�������G-sᣢ��dBz�2
iv�t�3��V����?���UK$��>��Y�$-e�dn��lFq˦����%��ym.�Ӣ.OWhXyR����˯�X�q�ЎI� ��C~1<:}�|0k����^x���
[_��~q
�6�9�@�~l�<�6��w0 �XF�b0�U�yRC�)��H��%M�<]l�Y���RQҺ�-���X	����%���t���� 탫���C�<�eU��v����9B4'�b�G��]����ڍ.���Ns���8\�~wM��tu�n5��t	B��ĭ\̑��ET�~�K��I��	$��xQ-���za4j 16]�lC�u�5���!dz�*��x+A����m��n��Z��H���͛'y�zas��LG*d�T�*��`��U�}#)� �6�I7�Sh	�Y�@(�6,��>ݓ���G
�s����ˤ,��p��A��N��Gw��H$圝�4�`�h�-m��_}���28�������!�E�]M	lF��f,aW��`�^q%vvP7=ZIsj��*���C?T�\?D{ �\���d旺��B��l�
f�{��G�IH?:���{���S�	���O��4|߈k�p
��cɲ�wc�d�ATn��ʲ��Z'$�S>�D��<�E�j`n"M'�!|��Y������C9�J��4�ԓ��3Ao}��R���1t0�{�42��{شX���٬?Td��,��X"����[����~�7��f*[�	^=�o.��d�xNʺ$�%NQИ�r����?vjΊ�X���ĺ.\�� ���9�6>T�㨑E~BL��ʐ �_��>�UT[��-0����Q�9����������2��d%v�t��WQ�R�	�p�%yH;�J'v��8V&(�`"B{���8x��E�f����M��z�ה��N鯟���|�"��]��b�!��l�qTC�wX�u���C9m�W 8�"0|�� s7���������\��=�"%<����V���5�Tdb�'
/u�5�䢜N��5^�>�J��-���9�E�M�+}w����:
�`
�و��c@�T�̓��ݜ���l�ICc`9�!-������_�[��
�)�V< ��/�Y��R���'��ׄi+���3T� ˬ�mTH/�nc