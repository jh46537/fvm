��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���9�{RԱ[ж�8�����������/a��:��#Շrb�,��Y�)n��M��Ӡ�5H�������w�� �Gx� �Vg~�r�5�t���5�Ш>@�t���57�s�f}U�������2'�k�l�E�g�ܒL�������(B`#�%��ǩ��b�y�ّ��o�ka�0��4�~u���͸c"�x���3_�XlB���J\f��E�W����	�]��8� HI{�s�zq ���s,=�G�:F�V����Y�e>�V4e�i��_�F`�mg�_}j��&���\���B�꼗5�%_����^��Q��q�o
|�zyFB	�9{i������ag�rʲ5Fe��Eó?T6��}��K����JN>Cgc��Ӛ�cH�`��(B�� �l��j�*���gjdų���\fٙG�%���$�����tXS)�N�����f�td���kt��*ؽ3��t�����-w��^XY���L��K@�Y<&��F���F7=��g���=�p41�z�Y~��%dh~��5���$/_,���\d���b�J�Jc�i)vs�L��]�U�Z4~,��7E,�~�<�bЄ��
c�B�(/��kЇ�6+���?'��X-%��,*Cd\�H�QJw��Y��)�>d*5Jy/�����֌��%�G(�^`��R0hL�U����v�A�k�3uNh��V�3SIK9�X2D+�����ٟ�`3ѝ�6&�
*��G�ӗBLc ��0n���m�:Ҵ|�Srv��?�Ь��P�[-�?��MW>!Oq�#���gXݤ��>�Ҩ���lWj�z��'e<j4��̂���:�1���
YM����<�'o��'���������$�Y����i`c3�Z����?��ɼU��,I&���wx/�j�#�MY���k�#� ��м&�"��J$��PZC&^����XN�ʏ�6B���'���Nlp6l��(80H;+��N���cm����7�[��G�� Bq)kސ��Y�g>�y�����sc��ԇ����vS^ì�<-L@]y�ٷ��r.�2!���^̵��$+3H�呣8/0^(&9@�"x�3�Rt0�n��ה��hjg)q�qܣZ!��OK/��.�8�~&h@cL���ժ}�pv�;P����,���<��^Y'[��P�5��
��y�i�D��p��S�.�v���r+�92���N���ȋ��3�HB��4WG( 4��ɮ7T���8��Y8���"�R��`]x������<
�
��R�ױ�X3�KP�.�Dc�"׍����e�N��.^�e�`n�4O�1�i���{�n�������^���[��zp�P��>,����[�Y�x��HC�XPI�>e[Z�l�4�%�Z��b���>u�dA�_��#<w��$;�(e{��8�Q|���9؂��E4���Nq�ENu���k"�B��a]�W��.n�HմT����G͈v�JG3i��  v��W��Qs��HCo�.L_��:�x��D������Ҟ��k�y"Y�)��o(���!_U�QLmcQq�c�6v�k�vG
(-�4>�r���w�����OTI��"\Ж�����aZ��{C#H���s"��z��<>$�5`��t���+��נH��βp:Fd���'&�;�/�D�������oАdk�8����%��U���N��tkɁ8:-1E�4�4�w�LAW��+T*E`ʡPm��!�/)v6g3�g�N6r��2ק����18�*pM�Q֢%�!c5s�(��aU�m�����T��+Uh-�$�,�rO�\l̍�CbXMC���)݌{���C���v���������};�::3t�4%��N���TR(ص�)*d��݊����p�{E}�i�{����
����9�5����Fs+c�DwTϹ�-j��{�z4V�\MP$��e����;�鑚���Û���E�PҢXX��Q�p������iv|*rx7����*3܌�f8�y���`gNh�����*ǥ)���C2R�K.s'�f��iN���+4|�f	��g�0�� ����[�oP���Z��M���kqi:c�b|+\5�\
.ozƪH�DX2ߒ�V<d�j��/U�c ��iB=�eN#��j��t8B�h�T��'�"-IU�͠�~��_l7�I�[ ��3�z�'����pnn1�Y� �;��!��2Cb!�[T�1��;hF�l�c�;u�2A�X�A�>z�F7I�����Y�Mo?,�=I��[����>� �n~��T�Y�ur>�F��MA�O�/І�~�W�N>�\�],ͤ�81C�DO�)ش���ݙ�^ݍ�-��a0����Խ ����,#{�u��ٓ�����\-��ڀk`�3L1����(����{�D%�7����* �������ȥ]��3U���PD���R�����z5h��s��Z^�W�sI��,�Hh*�,�4c���d�:=���v�j�&�菫��i�<|Y=����k��N2�Fn��;"~U,Ec���{Z��}�Gx�{�rL셼#�`앾O6���%���g�$�k4���?��w@�^O�Wʓ�-�>��� {?9��[eRJHa�S"q�CcI1�I.���?M]�qe��7�fF���}�F�,���e�h�3'���aM2쉾o7�IJ�=q,��
�8�6+�^��13{Qkg&��vSL�T�F;D�'Zr��2.�>S�m�v�6ğ; ��N��rl�
o���`��� @t�_�3vVJ��l��T�z���:5M���9%͕	@e�O�dl$�jO��k�l=�r�YH�^'-EjioҌo|�R_�ӷ�Is7��s�܃"m�}F%�/�٫c_d�[��/��@�y�O�R��`fS�#F��5�˪�� 7%	Cl��B�~���j�7�H���TΏe�y���v�Y����`�6!�����D;m�h�q��]��k����B!�X�8Y����i=SƷf��fgaR<i��Nx}E�����.qe�<s�N��ee'9J;��"�Y�b���;���%	��NFo:L�W��o�IF�\�`��V>�<���q�[�S�^%�:b �Q�6u�0+��NF�b��!@`<p	8;&7�)�K�v�[��PP����¬�&@�P@��c�W@�X����]oIIo���=Փf���D��w��PE_�����RV40�k~�<�W�l-=H�]�GΫ�����k|AQO2~ξ�x�R����+9�	Z�$Oe�jo9�0��^Jq|�'.䎒���n^���,gS�j�5Eh��!��u�S)�TA��%9`U����#O�b���;�� s��\�{Z��ވ}ǡl�dw�=M�-8T�v��@�w��D����˹ĞXm���'���5/���&�bo ��<Ƶ�z�bX�m�>��F��q�}�������8��a/�6e�ce�t^fo&6*|.���{vh
:1�\7�oC󷿭x�>�)<�+�F�f ?�x���pVS?�+<�����G�z�����0�Ǻ�=P����/�)A�Si�H`�Q���a@�����֞vj�؅��4�I���{��S�Z�'�OH��GzF(�s{0�.	:)m>�|�+|��b�[n2�]�&����r+�]�>�C
�#b(ׂ�̪������3�Ь0s��At 0yb�X��z0*�㱚�Į���Q{��v�1�;�A8����jss"����g}���yc�J��7�}�߯���4�P*>��
��b��C�wN���#%�R6V��&��z=�V�����+��)��X;Q�E�'�j�L9-���y#�&d�-�/���"h��`�o����^l��<�����p.ě"��%�΀5��{-�`�hZl|=����@/8Ʊ���W��Uˤ�5��<���9ǳF{�;	��&����(ꀤ�.�"Y�a�ԝ�$�@eB��)5���[B�J�57VLQEa����0u:�`Pն����_�[v�Ϭ\50ƕ���8Ʊn�8�v?��o����J��`z��;����"A�|xr�<����T&0/%��<0=����G��|���r����xA��H��B�	+K˖]�ͦQEbI��1�U/�A�R���Bl�O�������h֊F��D+��Y� ���~ׅ�����֝)Q{���c���__�y�0��C1����I�4��x��l�ˋb!־��
��{N�N����!�^���ӡ��ߓEs�iⅆ�q2MuG��<�bQ]a�X�R��G�x��'C�'�x �ȝ��+[pz2��p4�?���^�����4�x�hHĉ**:i�vբ,s��Y��]�S��~�qH;�^�G4���;A�+�V�����8�;o���l��D)��O���j;(���LG����q�+v�n?��w�7RZ��G��a�� �I�`�`�,ϐ&L*��˗���軠�T�tğ��ϻ� �pZ!w���7���Y>����u�ⷀ�%e�p�u�(��C��K�0��<�ʩ��Ux��%r�ǆ��}����w�U��Ɵ�0�N���/fx�ц�	Yp�`��n��me^�����	�]䬵h�~o �'��m�nc&}P����^wQ��Z��Ds5(�Sw�^��7yq}.�ɪ@!S��Ak���#�"cn�#2��->�"! �������#ji(�*�}�QJ�%�%]�܂^��p�Vc��l��i��j-��NE��^�u���&!�=���$�v{���2hښ����hXPп~�l���:�/-�"��:1U��5�˪�>M)�s���_�~rdv尿�DǇ�!R�y�����3������1:��{6˅��7,��[6�����2��7�TJ�LP���ӄ#WPi��0t�h�0��i���hZ�qM�Iv����yc�z\�6�������Rp{5<%����oY'�Uf�>�@�/�1�1�[��uٱ���Z���:c��\�[��Z:��ոK�٘��h�Mx[�r3N�����W�%�n��"��ۉ]�9��.�I�c R I$�����e��1X�u�}
]�.5�`�ja���h׬9~���J�� ��{���	Xh��i�sŀFc��:�\ms3���PtF{��M��z�OJ ����eR�Rꏋ���'&�ViPC�
�!Ie�����魀B��x��T%�E��N����^����d��EZa�f����!ǳ�x���[��1�NO+�oD���
�<L��6�U�d"�_�t&_[2�4vO:���1l��9¯'¡���k�e��3��F�I}O�[ku�_�ޚq#�J���Uwf;��ۥb��?���lH�@���Ó�+$D2�;�Z���u��v������!(�����f�Y�J�ӻ�"<M�����*��3�j<���l^��?������6?Ӽ�Q�̰��d���;W���5�V4RCփ�!�
�w��3��M�8����'��D���T��AM�>�}4�aW��+:[��(�a�~'�Z���l�ۍ=nlM�yW�"i�8�ci��U��\�8��X/YL��rޭw��|��#����Z��-�*�@�R���!�G��Q��8�B�{���=��ɥ:��V� ��6Z&�P$k�?��G��*��P˶��l����v`.(�.��\�tz���_w�x�/����`3S&��[��K�h����=�a_��%�g�����]���d�)��ch�)%;�:���6G꼾��J6y�K������YZ�0� �}u"@f�3��|��K��܁B]�e�T���P�M�����h����@U?3����w+G�1^.jIj�����H�`$�X\K���@�ȫ6�u�����$�᭒~"-O����|�n�}�0�(Fn��u`�	�W����M��gW�z�j��D�HތI�L�;7oܤ�(�n{�c�'EZO�9�
�h� �we/��'k�tW���^q
��Y#�%�&�(�R����d�2>_M!�W�g�uFr�꜑f���F�qZ҃�ա~nc�x�>�n-���r?�/�%�!�F*G	^#���B���k�>��m�VU�M�F��b>���\�m�+��rN?����XzZ�j���!j�Z��\���YZ$���j�>�P�+u;N�IV��}Q� ����
�"s�0,R �;�,	�Z�xu��|ܴO�Tw��&p$�O��7�2�����cӮ�/°=�0�&f��T�cS'��W�cW��l��9W��y*讆gd��ڂ��XL��
���ҳ��nm��������?��SȖ�@���b�RB�3O���ɗS۵�wz��3���c/g}�/���[�\������]������2�&O�pzmr/@���r4�{�@}IL1�H�����! qʳ�Zl���GaA�����:���V���O���CN�m�x�����K�����9����'�\h�W�؂�Ώ��Ga*>�30I`�u>���ܹ���@�-�Ԓ.�%G��[�Yd�W���VK9����b<ZcY'��������ø8L����������+Q9<��V�A���%�iD�uyI�{���E&��dd�{Ã�Or�f���*�[��:wMcs���M)�g�V/���檘5��#F�ћR�Rz/D��E�`g
���c3�ƫ˧���'9�X.ɠx6��ߴ��ܞ�"��4��r�	sۿ	�o6�(��<�ٛ*E���0�tN�Ddn,����d���V�K9\0\���)����+v%H̷'ڨ�#�Z���^�