��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�c���G�J�,=N�{�P.�*�@�&��^[��Ԇ�Ă�#�a��� u!��;*ջ�2��n��:#7��l��8����k�D��"3rd+���]��*�a���7�a�W�Ce�L������ ��5u���#��)�g���=!5�g]4�y��t�/�Y��Kw"������u�J�M&
Rܾ�a=�;�D�.[9>��_2�j)���&��%O���b�R#([��%x�E��8[���i��xh Z�ulN�"m*��5ߡ��!���ʛ(k���=���&�}�n	�i��8�=�(=��>چ�����[��/��#�qĪ�7�������m�훓((IF�YZy�r�z}G,mJ��&���\�}ֲ�n��i���*u#R�c� �zP�Lr�U��]o���� J���Y�\�J��_ա叫�#�/��1��":0jO]�T�F~���?r�c$,����Ti�o^��f���eq�d��U[/���s������h~ߌ�o'�%v�j9���sY����2D� -�'%��Sn��x���}{<
��i���y�+N�i��.�w)B����&�`�ܜ�ۮdA��@���԰g�TF[ņ�Z�W�y��t�3�����jC��� �Ջ����4��S�/s�w�,��b��u�ƶ�>��ґtչ�J���F%��j���`���C�3	��@A�#��|���H�E̚n�s�ワ3.���lrӂ�|Q~�]��]�\!��F0�݁ʃ���Z5�;.Aw�� q���p� V�N#���m�R��6���~���R�t���[�0R�Z�aK&.�>����?f����!?��$:a'�/)�P�~w�@��z�G�g	9a�8�F�!Y����U6�<��#������ş�Y��Gٍ2-F0��eJ���XݓJ�a��dgT������� ��1�!z,�g�
�"��2��1�|�kOEV�TZ��e&S[��n�S��� �d@\�E�3����&w̜E����+^A�9,�)��������.T�^5N��8j��{:/����
�d^��U��N{�{��ҩ��I��Rǀ$Ɯ!�M�b!��~��
��Wy?�g�����[��)���lj]�.f�Q�������(AD"�d�*D5��v��rv��+����B���v��թ��� ��)���9�åCC�!��JfU�%�.1�`����nNf3�Ʉi�=���kH�� ���U��%`
e�R�} v�~Ǐ6��dq��wΤt���.υ���֣���gIM�B�r���I��|��ֹ����C��1�8�)�F1�JE�~�N�RӖ��A˿�p�Z�X�3�u�o�ed���-S��a3c@���y�k���>�$������M�|s.��;#�:}�\ga=���o��!���m�j���hr�N�?�x[�l�8��/�G���j���_Be�6Ķ��ɏ#�wcr]@��
0�#Kq�E��X�//���TA}t�?Ǒ�2���^�wP�D�\M͝�l���8_e.oCB�#�� �#٨��OW�A�>�4�xo~�dgBΘc�88��7���<�`�;Xa��^�[�X�S��H�X������z���{��Jw!����uR���o���1ע��T0��y?5<k}�'j�x�V��f��^��$Ǯ|��������;-&�|?��(���i�%���?Z}߃UjQS�~Y����5#�T����TX@�ܡ��>��.E�d�R�|��;��-b���h�=|�F�T.��� �W��j��o{c0�5�΃;tM���F���~ʕ��;�b��nV��~Y"�g��A�D��&}�B��|�x�D^��r Im2�f�o0Nb�ۜM�7G��&ׁyv��s�v�טG��ܿH����k�?��Xr���a5��8C�)^�QL>M�17"�N���z��2����x(+ .�����Dͷ�q�KnGL�#%7���G@�"r��bcM��@��;=Q����:��'ד5���B��R�d�T�!ߠex	�F�u[�d��P�袥�������\ؖ�=�������dk�����E�
73R�����x|���/�S��?S�H�{R����^L���T#N�*�MT?*�+��VX8"G��*����˧�Oم��x�ٷ���u��
3O�@�Jo�F�c��:c�T\2�;*v���i�)�޻،����cDC��H����EL���$k-E�t�E��`�/LE!aV�c3���u�� �����/,)�Nb&���FM�[[��խ�bhTQ����)|P�րф/��zWtgsm��ᗩ��ǐ�����d�LVGӀ&�5�g	*�
M���H�߾p=�; �͹~.��ݨGW�1Pf�/��Β6�߱W��� u��^aWa����������U�C��k|_�k�=HLd�(H.,T�W���yĊ%��Zl���Q+6��ױp1��Q���7��8`)`m�=��V�A����,<���G2	=�ϴ����Jx���R�����ǭt;"{�D��˟�Edx/��]�,�N�z����U��Hߔ��!I�+7.�����q��\+j~�̦��o��	 �3Y�ARWQʃ����mMa=����!��.�@��#�@� ˋ�s,� #̝n��/ ������&�H ��'ԛ��z�Qv���CZ��H���ȑ0E8B0��\x���ƺ�p���6�S�r��:�S:�E���ح�� u� 5?��~�oy69qGo�GFvMƂ�٢5� ��S~a�nc�|��6�t�ip��N�����(3Ps1D&����2��qŉ`.9˄�;C!<Tq������u.��ҩ�U�PbGp?C��`P"��c��4��'�. )�J����{X����j�E�b�#+Rj'�oG���d"Y�L��=�DD����x��??��	�u�b�QӾ�T����d�xr\5(�v�y��F��{24^S�;0C��v[%��niZ��S��{�c.�����b��EG6US�n+p!I_�8x���X�@Ҕ�g�#���l>鷰��=4'���ѓNǋ$�Yjؙ!�'�P-���ә�����1�iy��t�'�e��ߔ����cw��$s�:8Z1G	n���7�꓍�����`�������Y�TѪ7v��4��6���X5
tDyTᶁ��Ah��_w[.�	�^� �����:r�����kH�\��J��_�����R�r0Ͼ��<��� ��:iy_�%���cС�����8vu�3Ythn�A�2;���D��g+�]:	{��6q3�|I��:��q�B�7T���N���T,B%�Bk��U�ht]�{��}t{��JQ<y{3\�4ه�<)!���+�1%�ڰti8 6�y�	t� ͟����M>��τ���6���ݱg��=/b?>��x��ܹ �(n��(�e��@9�|�<喇�����Jv�|f��WC���u���D ��/���@R��]K-�-�a'Kz#�_H��E?_v�I���Y�&��V�b�j�c��ż� ������K��.��S!��u֔�q����L�a�~N43KѤ#��>ۻP������|Bֹ#����i�I�%��B	�0�](�3v�~yC���3�xW�Rc#�SlUQ�:)�<����Bw}��w����>߼�iK���RR)�-��z�
+A�h�����#��o�,��=��A��W��Kҫ��^r�K�< 39��<g'z@.X��v7X��dF%t@^l3ʡf�e��B�<~[F̏0�+v����@6JIr<�l�����r'�B{���V��j�l��"h�P}�[�	�����9�G���,�������p��C	s`�yڮ�T����J�l��|{�AVk����R�� ����[xSe(>��l�s�P�Bѓ��oM}����"�a�����G���so�l��Ƨe��t�ꐞe�}��-�I��E� ��箹~qQN�۰���Ύ�&�Π�Fc=����:Ԭ\�8]��Ә��:�M&�MASp�M��ο��Y˴��ˤ�Y_��Eo{w[��J��`��U��v}�s�U��:����mt+���B	}�Ӭ��"�/���f�'�d������8l��u��P�&d����'^rE���WhtreB���|��R O��m�3��2"��ani%���I�<�nD%�v����b��@��<��Ȗs[�2W��ŻS�'���p�M�D:�w�C�pK�����x���ܨʾ��3ȃ- =n��a2=\�O���Y��Xv�-�^�e�>��RV/�(V� �⥫{zh�)C㢿_�ny��=�-���p��숒͘M� ���)) �\ݘ�ҿ����Q��L��1wxK�IG1X�Q����>��|@�]���U����v.��.b���X�|ֳM�g����<�s�!�@O<���Io�"�;�*u"���I�(��G0��g�W�Bk�ib���W�,�����Ce�U5��7Ѧdbm��rg9%*��l���30
�$w����L�J,s�����(ޔ葚@�x�G��{�%-
U��G.�#O�Ap����]���M�i��N�c���6y���:q�����HI�I��ֆu>x��������f5��2��X&̝L�Ԉp����7���}xt1� cu<��Դ�z�	��N��z���b�l�Ċ�wkȕ)>�렰���@Bc]�ߵ[���.����W�RY��Q��hz�I�]��O5����&�||���-?���ZJeX��%dX	�����S��8&�25�zl����j��@Ś�%�:�2v%c5�wήITh^�[Tw+C�)�`Q��'�D�=]���?�y��.���6:QG̺�����˾�8B�7Cv��&!�x1v�[-!�� F)��ѮaMy+���~�Tn9�G�Uڷ��M~hv~�G	��T7���m3k}k��1e��=^Js��7��l�yu�y�ѭm�^5x���ь���pw0d��om�F( W]"l?&�0��-1V���UM�6��D����x�����X68}|��t��CfQD�Z���zk���qJ���:˲2kn!�����U���|O�k��˓���"�@WQD�|�c<��Ƕ��/�ф��$�1�H5�\��T��pٖ��� r�ӆп���En=c�މ:T�v9��S��˷�^+ik�0��|�k� l��-O������=�*�-����d��m�SYfHׂ�����J��H�L��R+{��vJO�	��&�q��&��|��P�T�S�T���Oω��^O��d�ᾅ�������u��Q��������d�����2錕`*t��[,i�>⑯U���:�I:I�g��\6VxmKHH����B�q~Xj�(�q�#���ċ]����-R�!�����8��uR��yN��{~3�`�{� ͳ�ch���k�S��]��9��)e>ؼ鿰��k-�|o1M���`N��c�'&����=�l�����u���I�,L�פmo���c�!,��o���N��[�L�sm���&)\�4&u�������Y+��c��>D��~��s��b$�u�)�%�tt�g�R��5�B�`8={�@�:��2xh@���^�HE��Œ#7�ܨ��t��Ԉk�І�n;���ܓjN��}'��r�r��e��0�=][�A��U�)��Q�����{O
a�[L�H��1���?��y�>�q�!WQ�c��Vg��� .�rt.��#~%f��6�^i|�����c�a����&�R!��	����Az��k�>y�r��vp�6a�H8`~�n�X�q
������2YO���>
iI�8�C�� �#D��:�h�#��M�Awc]4����P�e�w��|D%!g��r�j��ʟ�̶P����cgl6@��Y����4��W�y�~"Xr��|T���/�����ٖU�c 1ld;>d��aę�%`�$�Z	!Å�vD���Hm�!�S�����o�<g%���c@CT�M=������z&�#������^~�AZ+�}na�n4���<�Y�^�4��WvTI�3�wt���=�a~^#���Wsl�bOf�<C�׊�T_�V0����ɽ$�����(��䎍��� �z�:%@�h2��a	^R�l�5��!&��hJ��"a��w"�G��7���Dad��H��yc��~56D �xiY~���� �`��ϡ��b����?cy�|� ��q��u�^QV��Yg8r^ͦ�	�����>����c�ۭH1޺$�,��iITC2�(&���(?v2C���W�&����)���H�c<�'�b�.���l䴟��6�D%F�6R�0�ͬ�s�D��m�a��(�o5ym�`?8M�dvu6|�Kd�(q�:H|����8q�PV��*��<�o�S���Z�c�o��C