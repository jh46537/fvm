��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�;��I�0�y���Q�&H���I�q�TlA�<�ЗJd���� �P����@��	�d�?��ҧ�iw�MԼ�k���A	Dsd�M��T�wY���׏�1�M���H�e��-�BZD�V���ȫ(_㨟���"��M\5��"�J�g�<X.,mc:�'�A������:_�+�**Ẕ.Q�~�c�0aTdF�qME��t��7��x��V�?�`$�U��'"𩔠��������q�����H��\>Cɦ�C�x���5�g��#�[�PFL�3O����֝fc�;�t�í��ρ]Wo�sU2i�*~�)h����v�b�tTOJ��.�%Pp�5�T���i]!��I��<�>.k�u�2v�����L՜�e�+��iܾ�0�������B�d���̓MwD�D�L�;0�"V��GV�f�/ni/E��7�|P}�zbY2L�(��+����C�����Zϊ���&���;q�4����b������&b=P��3��J��f��Һ�	E���B��nsu���v`��C�˷J������}Iٖ�Ǌ�ZQ®W��\m� �亓f?!�w�yd��nK�#��b�-u.~ZK�lk��Dy�c'� �|�j���R���Kw:�cDU�Q��V猇����_>��[1ˋE���E�����@�q��p�� D��~��l����ȣu���Dd̈́^7�ĵ֔2A�K�/�G�wo_BȚ�G�i�y>n,�N�P`��q�v����hq8��6���9�oz�pLPb��'Z�]����7�����2q�D�T�_��*�zj�s�����2�֩V�S�A J���d�_�`� ��~i�O���i��bk�ÅBm_��dx�b@U���� ��v��;��/���~��������΃rZù�)�6����7�Lmc��,}��|�PMH��4�����~lF��`A�#��$�:��t�wf�`8`I_���jE�J|������o�u/\%*� h<������pQ���J��a�ɷ&2XI_?��s��m�~�X���6��'�N��� T�~�ȝI+�g��u�9%`��N�̘&���H ���[����X&�+���JMUZ���-��u��A]e����5Zp1|��b�q�3/���8W(���z�O�������W�Şh��N;�k1��L���U�%�*U%�b�|��TE�~~Oc��c�� �Y1Ōا�#�)��ˤу�x�O�̼�*(U�]������ Iz��71V]�(��^[a��N�N���d�ؓ�+8��\h��_�Ѣ�)9���֟/�\����+fZ�Sg��<�,�Ui$ۥ�ʩ#���{�ғ��my���w���E���7�՛��ݾ�3�+j�drG�&�j���&0!��j'�Y;d�t;O�u�}9�`�&	I�+��f"���m��g�9�w�)�i_�����)�Io<)�V)"Ȣ䷗A�9�*1^�]ǽex>Y�I*	��������@a���K�w^�,�ed����� y5�Q3<x	0-�c��!i���:�6߈����NrW#@t��l������Qd�:���5�th�:̑+�`�*Y���~n�5d������~���7Oc��lR�\�zM֙�L�"]/:PO��J��HY�Ʒ��X��Mo,��5	zd�Ь��禣W1J2�^�8��Ă[<G- �@t]����`�P�E�ׯ/0/4$�~�w�\�U��h��������8(QV�Ѳ��m��'ܿ
�x�E�*�\���NB��H�ڿ�����������Eg�u{��7"|Pգj���>o�3���� wO����T|OvZ���(�dʯ�k�x=�ިtԕȧ���q�b�c"�/�sͥM���n�p���B~�����;vP �rIJQ� /{?e>�	t�8G�H�F�t&��
����q��!w[w"A]~p�'e��o�&,@��O��nO��65�`�OKc�(�8��)&��=�ϐ�%$u�sy��t �_]E������#mKQ�� H��a!V�ʄ�s�Kv�ra�e�_����vD�߂��a@�]��%T����bR�N���b��!�R[�U=z��!� @�����?@���-�q8���5M4
mGou��k�{(��%�.v5a��2m
 ��țQħN�ؐ��$"wI1�EM
�[J�,�Lů�8&���� ����3`Y�)},j9 �"_ѷm,��d+L�u�
©mA4n�+�x�K��l:=�۸z����˦�e�~ �:.�M�)Tϲ�ƿ�(����*����j6���e`r�'�g�x��!��򭞲(8�`D-�	�H�j��
�y�� #>�K���P�C�'i�7:�N�T56;�5��5��З��؀�f�k5~1����}�љ��"�ǿC&c�3F�rb����	N�т�o�؂1*4�H�����@FQ�����D�6h˷�"K�'s��>���JS��f1�h�N�'�_)�w�?�Y&�	ҳ�2R[^|�`�#�V;�"��tg��r@_��x���� x��a�~
v�1�be��X�����\�h�r���gV|}��2�D�+����R�-BGD���A˖gM�Ā��&+�EV��$��;�Q��h��%�ta'���J��<�3�c]��?j�tʯ-�	�b�ld� ����[!*8����8aJ}�ȭY�����/�60}��A�/4e�[�m7���}\9*w���h0���;��3xb� �I�E�ʔ��[����0̮��И�X����v0��v:�P3|���|�$��G�Sp�{�Z*15h��qp���r/QT��ݔ(+�J}���#	E�!�J�-�;�*3seT�XIi�Ư�p�Gm�����<N�t�H��U��d�J5��'��k�!�>эk_�(��2�#�5�W�����|onO���c�D��v�xFI-��,����9;�S'�Ɉ�}�ê�^��z�4�h �~�ֶ,���'#̪Ճ�nv�֥���Y���MW��:/����˙K��G���!{�(�>��M���@�c!�Q8[�0���^L��zF�a�V�Z6�����W_p�8�+ׯ�A����϶�,$,����Y�f����(^kcO���&�'��=��x�����n��_�}P��qs)ε���3'j�����4�� �� sB�+�Y�"��#)�`�Td����z�Tvᨳ�����m~��S�$YFik	T}-H�}j�+0C�0Q��/TX:�'�c�̚��_o��	��ۧ��1�>���Fr&�}��D��I��*zvCi1�л��W�)2��N�����)�+���`�Ι��a���u(�����p��|��E���נ��j�
%��{ Ӭ�brS�	V�!�!�j�>ci�-Q�љ��?����S��X3J�r�������{_bg�W��~�s;�+`#u�_��3���fO������e�w�\��M����c�ѵ�{ɶ����{���2j�sS�+�]� ��KHH��/AD,Ú�X~
7�Yh��g�3W՗�X�A�dWy׵GF#�\���"%7a�e�pLD���KL8\�1"�����pk<�����=�{c���po_B;8 tb(zXl��;r�'�U�. 
iѢ�B����G�M�j���]���2R���^���١���3ɇ��2/.IsH�G�GV��!m<�<�#�>��-K�R��>��6�Yy��<�I<�#&�^SR�v�z���?#Q��U
��IG�ÈM 5�@ӏ*�I��"_H�XC)ѯT��9�����M��{k�� �\��4yAk: �=P�T����/O;���4���I]�����}'iQ�f�Z�hDM��+!�f^�*���}����1�b����d�J�o��n)2���)�{���}d��r:��1.�g��r�W��q�1&�`@��r֩�������'�������O:M2U&v�����W��r�d��E�cI���#3�h�4ȟ]W�cؘ^���oN��� 墶%��FT28s��A,JB\q_SF���<���ӧ�5��'^���W��*���b���^�#�6�B�y/�ÕN����ޢ��|"_ӃŹ e�D�#x�1e�֗�!��D'�����U N�[��Fv:@�[�o������d����+*���I$s!��>1��
�K7ć2y�느���9�:h�����;d}r޻~�	K��q���4*��5���\�o�-j�~rN`jY--&�4������Xl�}�����:���N�����ݛN��6`��y��Y,��]S6sz�#�p�2t;��'��`W&�ִ3"Iy�mt�Ǚ����.�r�IA�n������1q�"�_�I	S���'\!�?J/�҈�����*M^A�ZX�
u�j�>������؄���p�2���+�¯ B��jze$��(��$�EU<�tĂ�N��L<;u�
��W隹x��
���C��A��/K���vM�fҤd������������E�J�ej�I���g^��y�9U��*�� �G��_H�+�>mM���<�4�l��+!��݊_L���Iip�ᰔ$��u�ÛQ������HE�fG��HX�u��u�.���&p��#��zj�}yy���*����>,�'a���rM�^�� 3{?֏�T[}[1tX��KQ���T��;F�akg�6�X����ʬ~qSR�����ss��H@=*����jF����/C����
��{p�[��(����'�|�W��o�aaʏ"�w�$�+�U��̌�>暬��&�U
;��: ��U~�Y��d��b�c;έ�"�9�Ğ��x�D5���nt!���Q �u����4�n7GX������<���K�?�Ō�|6���������ɦl׷%�<[S7��,jt��;���qz"f�;>�7�iY^d��S�T)5��>��0jJ�rQ"�����T�ƕ��cc���'��CԿ��A]��!9��'<WP�̀��"���n?�O��/W������FReOc�����bU6�i9���b�y�;)��#Fj�k� Cǡ�O��Y�9���s��2ɯ�}�����