// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:20 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
X1sDQZD8alE/Qsa6J/kbwWW2lbiZkwugz2ifgWgeetjJiJObGzWmLGkcASnYhOMZ
5yCWOdnubeTORF+8MbDdOHpMuTnK5zYteg0IfPOZSUFSRxANvqYYtwPksnm8z+DZ
OaQsX7/WgihNtiBaeoGlk2kcdvoUpda08s31BwlZQ6w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9344)
SfH5jnMWrciRT4djCsV5cElPqLvSbXcwAwgUbD5Ogf2P1N3gKRaMOnYxZVfllCKO
CHASwc0uBazvcMao3o5xhFD7kkJiu8JwXW9GWAiK+x9RmzajRl7CIIl5XsNXnpTE
NdosKzebpoocpguTtszGXVvGbY36YVR8g/+l7G1kGvHVKKKRsGNdYLRtTd59GrLN
8HjpDKuUBV623+SDdKJx9exngC6Hc3PgoSJ+evp71i7wNsbM3O2yXcV/oIXrV//e
LrD2kb6nYfuhaqy6xQMebTEcqlCOSTNc362d5g7ECkSQILEeW5sUJK1KXkKFU9D2
aMjeRm2keSfh0hIk4ClwXC2a3jloFyPELIKIZ4Gi+c/UJ1JZ0QXNx4yZmQ9M+jwi
Xjhis2vQJS2XNSBcm3aE+tID/DA57XDwG0cwZBIwm3tl+cMFI1WWwCYG455cT2nU
dKJO5KP2DK0CVgIn3B3fyXdu963sCwxeKReN12GDG1ARwLrdhHxPyQom3u3pxPaW
YexinydQpiFuihU4yq31syfF3qiIZ1E3GTb9o7tem15zSMg+o5XHIrOrxP/oCUbv
sbLrmi8zXLb1SDMt/YlviAjwOykeeG5EAZ32xYHLm33w7X0OMVL3DEs5n8ttzGIh
c0muhfCM1WEj2YDUOUJhGP6lFl89ieCmkVXAym6fBC+nn80IApOazCZMzUHzbajK
YEjFXN8wv3M22hQFEnYt1DcKdgGR/LzGcdxYpQ7N9jS35Xojooy7HilLpbDX0ok3
F6goB6opLJGvYTr8/uD5CbSPuUC8eIENiq0pa5EFBjuhrQdv4rmlXAVlbhOnROjx
Ojxhzs7DAC94c/FrYf0sAMp+sNGMo/0i40zvdDAzil15HYw8ANldmypJ0nl2NdPT
JoboTHHpPcJ8E7zizpJBZn04qwtWCJM/YTeER4Q9em5D6jBOFQsiJA4roekpCUU/
IPbaYG7WYDt2WQt02n/ed+2HTX73GXMDdwoGTH2GSTxGbaDEaGNSQV6zJ7P5u6y2
NkRLzW3ErsfkzBWRbQLeMT6JI3OzbA76BwbRnlquLtfVmzjoN8c16V1Tk+KYX9mO
45CYtw+P4scWuusKF6st+4pVzwxpLADLWx6lomh9Iz8egRzYVBVE5aySTkSb8iRv
Pdh7TyPdj+2wW1lx5qLAv7+D9uiSIzqcs/onIMXvnqdqh+jfH5WQKQs045dq8bcG
qfE7e60gzWoj8nRiDXynVm16BdIN1ocZaEIP+iNYjVJH6bXCrNpK4KYeMpDbzVPp
KO2MBAqcB7yZfPX6mwI4d+5LVlp/mPgAoirgWm8dSSA6LZn6ugiWI5mpeSaoeeJc
SNWq+2sSiP2mUbnEgoMowanvbtf+9zG00zVhoOJ0mF2uLVXdhcwFDMazyVdDDBoa
FfpzwCWhYN+5F/JQTLqj3qYjRHqtDqnAfndexMo0CcNFlLoL3fJOtA8ZGseMhys3
V8P7/0NiGs/Wfooudkvy5NtBQFKudKY4bK5F0tYd+aIi59Sir7cw2cy1V6d5vw8r
vgfYVTi8qettthcrh3ampfc4wQzE7opxpQ0kt7yjzvcMZo7Zz4BO4DfKI/OpHhwN
ZmuONTlVABaXvM4CwNGWTAWoggcEyqrfAJM7XASmGrJjYjCpRUKNIUJge4siEv09
vSLVfYNBQFeGHL8xjF19VW7ckC5eBUtH37cqmqNQXkUGinQAbWJfzv88hZ4qm1Pq
+2IFrSyK7ZC8dsbbcr8aRgBHD7XAWIy5YEi4MZNfQk2EItyRz4Glotv3ps3wUQvj
Xr9ULzJ8DAWm5p+Q5Wp0JIc2af5RKA64XvZPyvcIERwwibbuOhZwuwucEG9na7rG
dR1UiLRrgU2XFRekJKLbMftU2dWBiUv0VQRkOi4m7BlDzhF0b4RxxUO1susOBJWJ
1IAYmBj3qHsQFXjFaXiPrpnvwcmyzg+LuNfQMs0iPB8cyPPKJ0kPKyd1rLyTsJG+
DX5GT2YXB3YxU10Uys05r3UPZ4hatNKnmzYHLyeXrzorSKKade/3kx1PFX6U6d2f
FdH6RLtN0dvB6znZg36Ba5kTJeKKTuM/AMsrKtHYarUPg22goj+tGjisxOCX6AZI
v7I09j6766CQ0DJunspa+6fr26AEpjPk9wLlhd5W+81jJEZ31pAgtTezIvuhpOU6
1+uSbmxm1NNJoMS8VFUL04zjMkw0w2T49sI3lW9oOfuKOa297+1ebgU4zh7C1+Ho
GMZC1w2gD0ceqr2ITDPKhz+T9sJpatjJCTCYmnd/21lOjOBqD/rXHINdIHeD+IY+
rnWO7YU3bFHyC7anO/xMDY+A3NkTsCGfPJ596uRd+sXwgrHNQebp0cLnMXW8Qe0g
VqtBYUSHlzzlqvMuWiVOwwb+yRhN0dVV8cFez+aFHFBNotzKTv2xRDT0DZr9Rek7
L+witQxwF0fgqk68xaS7X57zok4B37QKZiGyHjvdeV4vmf5w0d5v1i7SoP/ZEJVq
OHWu6j+9Fuxv0NLWN26KDnrKsOdcv+2ceD65Olqz/daHu+GPwjKPgCWNy2ZipzLn
XfD5iohs8wPjJdINyln4AgzW3w4opM1JjMsefxLhhPdaHr9N0XNkgQrR/Te0pshd
pPJtqAVMNCI0V0Nkbx9cSSh0FoavqL8hxzSjGhMzevZpvwVufsZvXvHza134IaCv
j8bmVhoi9YzSIVdOiXE2riEYkHIL0AHCp7ChXjxq5P+v19yPxxDWB0jv18y0El0r
KZSkIdeFpbv3y3bzRtH37s41xGGvAYgh0Tov3euu9mRwCA3leL4qMIP+68y8wa5e
j1oZ4EtbiyFVLEPADaROqAlpaLYiP3479iIwZcht+p+cNUvMaLhLZNlwMSLswEYW
Yx8Ighrz9XvGuVegbo3UcL9HtKtlw1egUacTa5G+CZVoXwHtUnc85wkcxYR6knYT
d8idcJlGE4cFIpTxgz3doxoqmdnyaNA8SKSIVAMD/5g1G1MMOpf+E+CjaR6vvm81
EdSWD1fhRFXe9Siuqsn7FJX6HUjh3uC43F/iRWnowQF5L5WrpV2ZmVuuYlIDVHSF
YYSJ6qFJbLSX2MTJddyZA/AtbM63QktpI1JTbcG03pG4uAxNY4Lu8zkOEjuNUbhX
5tzehwbjEpFX6YT9fbTbk661wESovVrzn+1es5qhR1NwMrWST03koT3EmWUB0Cfb
jbIYgZ6nVnNi3wbH6iAyE0vVfRwYCYVqpvGJT9PucMTcd2cG6POKU6DERNUGCcFV
WypMNKIsIGC4PDrfckHyRe5xyVefK+Sgx8YkVV+oiwL+MkBTzCGdMcS7X5GsCwTp
D9bL+GzHf9iyliOM1IQ3mu0SYGk9S4NZlqQs/QbZynRDPPw8dTAGtNo1ZHfwT21n
7n+Nh3d18Vv4x53WiX/93o+Dz1Lf1rxa6cEskAXx/OIJoAAq4MVT0pcxrIuj5KBU
ojvt7j4/ANRKvFa5EwPEspqybE9nupx+AMI+mKm++/1f7ILAoIWcn3anXF9/L1bm
BCbKExMEWA69MwdmlssdROOKNEIUMHOTt3dQ9T0lyppkde3ZbdwFnIjB0ouzr5Ci
tm3rmEpbHwu+wQwcPURykDMtf75hIEZLlxOPGwL4mswn8C/hViIdYyw+sLQB0mXv
vb8bk5gJivkUmoPKYqAp+RKWgPKvTVjpTTvdXMeP79z1cDUV3pCtD3U9r5a4SDkL
+i1FTVn2LNGBjwoPQNmeyLDi0ZOr/YlRXxZe5bzxNRhat1sPfjImYIkeGV1TM/2I
xIZoTErA3+WlpOWIRZOTvg4rm8VVeXGC6fXJ5YxtrM9ED0gFcxqCPi+HndcSJvDa
By38xu0j2AOf+hllkv2+kSgZ0HPnv62GoP4++lujGI8K8XuPW53645dCCPr+lCTJ
RE9sZmqEMENUFWVnvNqniVN34THPxGy1YG5zRpqitkCTON1GZngXZWB0DgO2SyK4
GSTr4bi5vJsh9u5kDjY9phRddwDVxDq95tRZaV7iy6kTOE9HXvOed87hGlBqoMRm
FnjH/fxC9H1/yImFLmb+hOniEBr7rwbnR1zhIi3zzEqMPOGgw7IDFpnKAZsolEer
FhWzapIDYEZNQBJLgfNb7SchaOsviV8BvAt/WALGjitXjij41JsEgXAAMeIBAX+u
YdqWHz3gma9Yvvz+gC8MIMCqES85xGwrlunutEHrv7Ylq89jgqu5HIdDVKjNrrJk
Q/P1G7OJmpkqvRpK/6kVaY0E5xLOgN5x8l0Wj4z3SBm1w+S3Dn6h6y5XkZ2DjICI
2hLjJ3UJq4kgy49E00aNWHdUqxAcJmYP/47DVEZu1fsvGo6ik2j8j6pIuDHH9gtW
j0o6vpNBLRil5hqRhwx4VtwBUaEbFRbqwwaYoIdXfQJCXOf3PyoSh4fmUwoWKKBf
nBGTYz5H1yIvEsTNxTZmWAFvHnOJhOjoCm4BURHRs+tG2hsclWloU3K1+Tj4cApT
L5PFFXQRhKRtYUQ1ytZPC2AlxYRLaFM8abBkZB4BxOSax3evwZcsCY70Byrx9OVu
D/4bA4C1r28QnM8KqJaKTGYvcUhjJc4NDig84dlpphlAr4A0fOI0JsIcFLE0e/oN
ZAZygfuzKC44TQ4skdMQO3EAYZa4YS7Tbb2AGiH854Bjpg9WyiBZtAjddG2dTfJv
Ui9Fpuq+56/Fa7CnzRO3fjuQ07RqcabMj/Z91QT6I6MmJHSjTsE2hUUH0SOfjAjp
eVzOb1nK2LUbLpbEIxIrl/rL8QgGAWRwVA/M4pFQlyGrJeBJhVFKV/XuAuz2qAzC
xvzEBEkDVPMnZAJF8T+RSU1CRgfpNIDG1xZWD7BDxdLx3+3KosW0Pen5p8NPFPAy
asesH2GoyHzJ5FhgTcbPdN7i7rveq1g7b0q9zX8DngFKJl9BQAERxq6eS5aprESM
UW+ZMydpytDG3KKziJgp/KViTfus2rg0lSTuMLe0T1uTz9Gn8Xngh5pW5vk5m/IL
vIZnNXy5EZE68IbDUYKd2rWkaBfKYvG4pQofjM8WeRU6DnlEumpu0YelOdeh6rJT
KAyUe58p9mjRhjlM+ZVUsDTP9hatqBcDWA7sCw2F5FSlAsR+meQPx6/09J/usAV5
j4vcY5KWzfsAZD4Urt65Iv+rpME20I/Lw7buvqE/7T/BkpaIONhCN/Mv6gbqRGmv
feqfEI6HX5jHKXoloLVlOo50Jzyb2cAuXQK62LOGMM/H469NPunXWMa6I/Spc8/7
6KnCGQ4xAXNXwsuc1qFaWobry2NbtAK8Nu57CBBuJm0ts/O3M5naQ+ZYk0ghBeYY
cVYND8Fl7EjKt44PHqOeSUZHSsj9wz5u96KmX7u73IK5n4Jxbyd1+9ZwyNcLaAEj
gG2l+AgZ8ur/ky/OFdYuEiTJjhb/IMXXNABVc1qJGHtJH9pOLHvqHnrVOc+SZ+b3
VBEZRY5vggE2QCLxJFcU2QIiyJPICZmJHGYo40q2xkGUfoPjfHT9rcUtkRyVS29/
ogfY+3zhM3bJCabb1S7sXbi6pcTtD7kfNEgkgiEgUapUju6vPLv7Yooc85ADEjcl
PLeLFnF3/thonQacwQEMdilDDj+kYaqUuOLohe+l30jQRWfvPRNjamva42PNbtu3
ABHEovw6SZ9wZJWSYnp3XiKVxBMHZoHPWHzOnU46329Fg2V96ioWw5mySpp5WHoR
WBHNS1yiPDbVNcGrvde3w1w2GKwbBr7+Br0S1BF3PHgj0Oxn997wlbJbgYzMzH8V
YcEC4e6q1ciUW7NAKRysxiBBhUZ306MSUeLJUOw62ohUF7n6MDFm6jaV1TMW0D8e
fyfWJIyWNLXsMNTlZstovxD/FA8fCEuBAcXF/aToowDZeB/SZ35BrclLfPKswTzx
6anz1pGCix3R/KjkHBe2LThav9xIqxj4XLScF1GdJqW48JJ4VQWkZ7N9vJAMHgiV
MEAyfXtlBaWBTkAR8B/ugRplBbZZ20zZKoPKiqjsm/U5y/zPVgiNXoERjzRNAfsJ
5T/VW149WVjwW0nmR+uD4s5sUtOhFptCIQVhUb9I4DsJ0pM3MsK1gwS2JryI4Ew8
jwomiQkWVRdvTinxs1p2f76gG3v1+whIDt7V/+P1db5lXaJH39HKq4OZ6lHdCYL5
aJloaNXnEmpVCLpWSzij7BxFk9MYdFfbHVU2HvDFxHh7i/agRVy0fUfPYR7w2YYF
mhacv3erwkV42FGzvkw0iI1cX59hx+3+dPHJtxWABcFFEBqxgEFu3i2eGACJL02e
cboFDYvpGLagIIV8ih0aKvZ7To/jl7G1RNyhxjGk9SnjTMJxt3Ldl6YoD6wr8fsD
SnSGVFsQzzoYSVE/HKyesRckVAPUttUFdC0NjoX6WY9gok2uC5bfBebAMQ0aNmm5
Af43IU0e4QRod7tb7k3b4/0BOoZABa7l+sujx/XZqq2AKjMlpbX1P3zfOU8nwarR
Y+mUKBZjSa381VVpBfd7Bd2IaA0j4162IiycrADsAFfnpOWBEvWKrcT1vD6qjU8C
f3r3CBd/ibvnE0nf3HaqiQ4X9s0kwGW6l8uZ7uGYU56EAtgU/xqyqb0ji7RXv5HQ
mEpa5ORtNsQe3PcBYnKywOTjgAi2G26f1ui1PPJ9E2lc1TMynxmXkUllTa8qmEDi
MHzytCxqcEXg7kbY6HTsKcvMlZ3N9WwsI2dYgBdxRlB7kaljuolxMZ8JZPD2XQ5q
0hJwi0dCu0zPZ1GcAGIXGc9Cpq6o+jxZSJJx3pRzfm9uofpZhfujrKhFDtePavmP
RN8KjVvGIZYnCzvJPpNMTbiWMaC4YapLgHexfETrRXfYYZNVZ/M8BHnJWq0/owZs
bjKmMHMtSAiRe63Ucc+N902rwIkOq+rKr2NXdHnNJC3DTc1jFyNvtwll/nI2OCQm
L4C9QM0BoPAY+GCex99Ho5zdEVlfD5tJ9lfbdFR3GgumlYnbSA5MLw5BBOmvRs7U
6MjYCvMd7wn7sZb96NzAv2kp0lHsD24FKvLhwJFj/1tvS9BNfj/8oGHU0Xoh0GMO
LdjD6Xb8R4naxcpZ21W0VRXYRgKeS+JZT+G67awl61ZdHDsw2visJy6A9Zvuikdl
YWfeud0bhDEAfYRCnL09nP136O6UH9gck5bvC/hoqlJcjOjFOksk4/nQ2Q1wh7IM
bJ8LTJQ/yhxX7Ec4+WKOU40PFM7k7XhhI1JPLmbHjFVMBS+ADrtw1OG4DpLMNn86
uuzdxyHT/3gHdHoslr/XlSqUsvcurQkCFPu00dskQA4EQ0I7voJiyB253SSACeiw
lfsU8E893YC5AuAcJKiuLOl6cljgoowu1HN7gupvjkf+KTX2Fez+LdCqkL9xsCxb
/crI7wcSu2TA7/Dy8Q9c7KUIgB2iAi4m1qY24f/nuYsCgA65iOG06TDwxCjNH0Ps
sF19XkryhCdlPiCn2hxLbgJct6NBp/9mJZd1k7Lw0uS8Dh/mFtJMCrt1SoV7Y4h4
W+GahIXwsZHAmxzrS2prmiDIeSn3jnj6W89w2ji21/7XYq8cGuh26892+TQUOYeJ
XX0LZR5ZODnMmTLgQpII3ji0sqvUGvKgPlOGToT2QBKmSaTqmkNDC3z+DWnyQi/C
AzCsZ+W7TTKof473MgFrQkQl9Sa0UP3jLXZyLwTNWKzoQXWqFrgDGREFgx/9jXiI
Fo7VKdq4iLpYL6qwgsIz3s2s+13NBDWH0mO0mGZgaVYp1j/fARxPyc5zqjfq+tIK
E6Sa5oC/OZN7aLExr3dY9TtrapsA1l9ln/XdMvCkpccecgPeqUw10mN59gGgtdhB
xW5haJpEQfDnsNpaFyjkxmUjEgv7tQGFhJC4PaBM8Em1cdwP/gb/6XnBm/B9wfbk
Ga67xuVG1V143Z9rBbhJLAVZGR3PJTFw1VlfcNLJA0BCzv5x14uQGh8fRJiO1vEp
2d0tlxYOswMkoJfxJmBrIEjCAEbFfTW3J3Jo+wZKXVotZUBYz59nj1miQR2MH7PM
E8u6fmqvAGlyF6cEtswhg6QT1UF4grHYBAiKia0AgWzqgSrscNU89AU+EBQFdxL9
vWV6bNJuSmQNpsnvP52sZ5FQiWRNB9JFs8GaJMduh/moXWJU0ujdbhRm/qhWZ0rq
aqnBS/DGnQNmKEgIDjRxexAr7x8K06EerbMuStkuKjn9mabdJjp3EyMfBRLNYCtF
g6JT4wJCEGZ8M+HqZB5pLXcDt5ovu04Y7SL83+KPuc8INmktXYedy4+7ofJxZkWQ
PN4bPSktU7qBjsEBXqtYrzr3mA4kcEtg17NBOrZjx1zb5u43wrbMc3De7f8ojymY
m/dotka8gAfZjuwbCl7jALpq/B6oq63GBwLJDZ5igGfbBP8BblMM4zZPS/VfYWwP
5+EG0r3P73xHuRubmFK1RVCA9pf5Xm3eSqno9+AM6gVSjmPvjDZezDTSqyf9HE+M
y0dkkzZJ8RICGYMuihmtXgDz8whNZvLRLXs/c/ZqRYteYvAUbq0lcW3d7VULvqZ5
FwAB7gJdmFDIogUeYDv+2tex2Cpjmy2jx5wTvedwNZi8fF/MvawrTdzsZ91MIixK
ruklQlb4K+IpoEpsrAL8Wvd3zlW5Ganr6iDQ9Frs63En9sN+BWydYEtDA5/dtXM6
q6VrL/PRuGuWRvqLbj9a2/3QXfNDAYJdXNuLYBKaigGJ4gEhIioSRRzUXjApi0ZF
LqrAmVg/lfBcvtBk06VPne0Bnr6FCyz5KKLA0LtWYp3x6ZdqtSw0FbXl9AMaveQU
ILxNPTHx27ZhtRqcJdQeEE48A7Pe5VZxll1iP9dE1mWw3OMwylijZ95O8LL64UEW
bsh0dRqX9EEct6wIQ929lwW8V9uaXNVoZeGLWhhWuQMhX8s4P5REHrbHUhGbWDzi
JjVcCCD8AYJ2vJUjleyOUy/9srCcBH2wXtUR9p/wXO9/l3eNDH46D4V5BLVJars8
zta8YJpivp7g21V98D6w2CvWgwrpczawAgmvymn4Ouc6H0mtSRTKZgAPnlfUgEpw
+g3BW4Gms15zeoJ1PzaU3G7kKuZHiFR5KRTOzND2oKkHA8an/aSK7YvwGTfdyQuq
YRPKsbTwogUqH/N56J28P4UYl3nt8u/EWeqxkuYOpkSgERzMGTO1++EsRBab9L+r
77HxmYmwdjzTiEojytjoo/9UBDgEXLkzv/ZigYkro9YmMLqXdeaDaQv1PrrffuPD
2UBgEc+HPFD2gFBBq+qxiAbGqTj9YrJik3WJWQ1Uj2jHIX0k1/3RCrfTiqJ+2AAw
NDMTiM1zhms0j1vU4v25sNzx7HOEnX9HaZ72KDDRV95rzjxnw/HGeqk5c3qqhDM4
iXohjl6HiMf/rh3oIR2/8S2wjmWJZczAT0q9uTSZHFVGB+4gFa9sCmJZ4ll7j8dc
jsq/cZIWFPyk7VLTEEYP/VePxG2Dit1I8iHGUn0VNqXtNVZW7g4UQfds7Yl8/UeR
ImkmJuHMS3r4LXnC+ZTxd4YaDNuWq/q84ITYqhnE52lkVoO/DPQs/4Em+arh7QaG
+kKXvcSEeefrstPuP8QSTYmVtg1A6Wwt5z2xL7x1oFQSMx/MzsoHGXDRIxkEKcIe
UoWrt/QhfaqQfLB0goheUnZC9dOgImx3bly+CTZi3yeA7HQyLC9qJhqf2yvO5G7h
+XYWWj2zOErdG+DFE+Ssybm19kwzNV8gFMr56MyBMCQ5gvmsd3YPGcfUQ11NetGd
8BbicaKZlIvlEZaFNRybtUpufO0dUZw/JojAztBl1xG37lIojw0YaUlfQWgmea7J
UGIeYKzxrsnwJClAupYYdppY112nnvqQvz7rTMlre5YtJcb/WRLZLI0ja9ev/xfy
blS7w1xONlOMJzsqAfH545TEgNqXIFFwR6U7FyYEMQJ8E/A3x7wY4qY/jAbGliQv
JxZutvy068E2UfLw1+vRujc0zQPgJeTGPXrr3sgmKxtuZoWrsMGh+XqqiAPE+Pkr
RAhyKkJ43Aerrbe+koGTdfjC+L7v5IQSawLZod/jmjoBNZCjUVanEeAsZjgL59QA
+f0VOXfChIGiYgdE4lgU76dcgKZOMBc5TbD6Rq541cn3dTTZV7nWE5PJl5Mc/EDj
DzNUmLUJ1a5Q+OHbUcVNnNHFCeI4u+u87FPuca5IK2oTXAtD4BXEiVJRW1n9r233
yC8iitL9bDtrjuMrTwO6R7o8OuFx1xCmYy4U1wjnxCwgdDim/qCvLh98sKCvyfGW
nMXDBncAsB8x96CafHHYZAZa+YB2l/U8c1Xv0gQkEy7WCeMA9HLbFmhoYknqdFqd
rRibUKVSMQc5LXiyo0LK8y9Ic7kjY672+7PDeiYSqWhMV+vVDwBw93h09TUBqUFn
gPU84a6gj0BtENApebomhiUB69YR0JHQw95SHtcPPv22GOE65B2jl+/46xAB9Dem
Chq3uI2fpz7Nx49Etlu7mYkydawKbzW9orb94cgIiGFk28S3MGs0LfBAmLZzHn7H
SU2eYOVDZ3LaMXI24irIzMw6CUeHiY+ukMthCzME9VSn6z0K/AwtN2SVJW0+Jp8d
11ZwgWLP/W881P8acxT7wBG+kW9LBq/FexvzA/P0cUbohZsZT5JiVX541p97rqi+
zauABt1Lt0MWpmmEHlR/p7CZcrVspmQvPK/kCxye1EisRIJFPVmAKgDA5uityxX7
IyXsD9QaYn9Y23x4stgConuOnYjuvjZnkejm9GC4O82xyCkx48iFm1WJGm+Uk7Gq
3bH5qRWDcg9WL6YxCAKAyIPI/miTit5RkUGHdBD1qeyjnuEW8vf+cGGVNWN+nQbl
uf5Tg5BaFCP7M0/pX0HIxRGpLsYxmf7bwln5HfJEwB5M3L65J9tYZA9wLTpAyK5K
mwiNz3baPVNIgoX1Oc7aC7EVXQXUswPAlL+KJshX1TbkJeFdCRX1BVWNJ9NUfZ2i
dQNztUhgECWVGx9AWd/9BQmXbY08uvh79D9MwgAgSvtMZKle2jxb3MQrHVtjuMSQ
ZAwag8HOO8AtcyKW0I0P5P9RF71Bx2KusTOOgh7hFEu/1rAheNCKK+ZLuD2xM+B3
C7VAREhgqZ3UuMnGq9Xbt0dJ2htshXQ/BWGcScrbBLWkWlxPQFnFm8ImMFQDckO3
8vH7WQPK7OZGDaGLppLwxf52wGlm0Wi7gFq68+kRSWKX5y8tNUJUldgVwmFKO0VT
TL131OiI/LmW/z0NHhpWZc5MNwK+aRn6Ymj4+7s15ubqUc3zYY6AbldwqYpsQGBK
KOT/osSSLppD1iXVD6ElTyh3KcHd8u9OgfQb7hJp8dFspWj+HzK6TUOjHnWcGA2i
csE1xBSoEbQMVJ/lEXT5/1LZc3G/bMR6dtMXSAuOCLouXEjHi0Yp95gsWUP5D0LY
Dicmh+kFIeqQk720OJAQzq9L6PxtbM9B5XpGYcSXHl2NiDGtQglNGimviO7KIckB
gDOE1Cuz5Uy3k6KMtk96c1MfFi1qYvwSQmM63Kp0QbNI5A0XdqaqOCK56znBJAzM
I4ymgFJOPtE2JIyq9aNd6QIC4dX4bo9GFH6s5KlqXm3He3jkKdgc2MJyCBYiWVrb
5R0nW4v0tQUtUqehkncKIb5+tYXuT2BZART1W8xd7jmDClOTFOzAtfldpqUHyanZ
654QfSJu6R78S6PryeQ1JDE3JNd6Auk+WVesLdegC7CqbZrAvccAQ/uCx2/Az9EX
V15fEUVgF24oyGUHPDBj2rJRpOsAlgpn3fowAOFMyHzTpSggm/jTk7FvZiiV4ak5
UkkLubnN6MP61GyO6qEg1yELOhMYPR9EoJ+KTtKWaOn486l13e2yMkxdREdS9z1Z
PLREmVzmd2UboR4HC89XxKp0I0uDFfKvsgvecC+jqcGa3ag2SyUbyMjSfyfeKm1u
sEvzL7u2z0LhDoCRMHAbUqPPtGJ3jXGz3UNcUuSklbjzFs8gVSvqo9zombHXWmog
Yl2y9noHiUK/dCy9+qh4lx5+chGgIxomhXaEh6HFwj758TV02Jg3gAx1hE7sq/yc
KiHLGeZMuUrabnoWh2ywGk2a5X6giAftE9botijlDAn6Se9/p5B4YZQTllrUWG/n
R4s5YjVw9Ny54T/MGHw9fA/NVAYo5z0aG5ZYzSAuJMesG4gK9z+LkJRhRTikk1VO
Jl4VOGtG/NH9/aojLYV29NJdU6SCeyfjGUansZCOOWRzkdGHjjZakCM1ty2xQ+JO
RwI4IXbnsd1dFdBTRyY3W/LIpgLRgNTGluLeLUx3L99RO4k+eh8/LIRDzZMSp+8G
LYgfCb0kHa456zhcrEcADaA9CfSm4nzsAe4fNE0DhLB9tGakglyTiBJncLxeLR5R
230NojfH50JjspeZtwvkzelgVPNtULOh5QT1nPUd2qCA43euTzC5RXnsXZxDjfZe
6eFW1PD7dQfG4bzMhMvunJu7wYqqgob+bm7Cb6v93hY=
`pragma protect end_protected
