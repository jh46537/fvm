��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���Ⓞ,B�$t�{����c�,�-��� k�4�	��[%��B�?���4��\�@e-��� ���u����'᣸߬Hӣmy� q�`L�S�L��-|�,���Ξ�<j�����̨O��f��U�,ﭵ�h���voҭOu���[�)n�g*k�<l��p�l�O
?7�""I�ŗ;�óR*�w��!��c�Z'�5�i�K�N_�P�2j��_�[Xz�q����'�&_��-JXk�ǝ��=�e�H5p���ʛ��ڙ��2�Ḍh��t=�*..�^�h�Oo��rn��5�Ħ�K��ec��D�D���R��V�t���w_]M��v]�v��n��NF�+_�|�}��T��n#�<�1V��9�\�
�s]�d)�Ͽ�Mvɑ��!��,2<�:v���2MwM7@�PK���{�cI�4����L;?��������p�����ɬ�'/q� ��o}I�����dp��C)�����8�CJV��$���_������Te�����|��A�!~�5�·���a3�qHӤS1]��d�lsg�-V�����C6��G12�%�/��U˦�\���G� ����?Vl��TH��~U�\(;�dS��u!O=��o�IoR�4�9�Jj��*�~�q��#���v���so(5�W~��(�/K�Xj&�=��V�Ք�S�Y�n�Ep��e''� M�i�`>2l|��Ku� ��2������:zG�?t��W�dېa(y��-��;o�Ym���*���R��sm#�v*%>�l� �Q�lG2<m�p^I� v��D�����#�*"�!S�VRi�5<��;E���]������N��q�;ܣ]�1V���DW��<�����*|p] N�O�Bm��% �]	v�(�za:9
�f�/�������H�afڢ�4;
��bh�4���2�96&x���dat>� F��6�!�7^�^\� �������Q�j�ɢ�_�3DM���↽�817h|��;7oϑBVeA0�j�_{���*�<x�Z�6k}� m���[d��P�n�@Q�v��[�D̎���J��H�y��S��x���:�=X졐�'���Dͩqrw��w�
O��47�p	+͐y`pЄ��y�k��0{�	H�PvÚ���c�6�Բ< xB���#������)�F,o�ڮ��R����^��;k����e�ԃ�S��A���Ny�lal���|�������2����ݜ��E;_�z2G#5U=�3a�.�=�Saw�r�݇>�Ƽ�V�'O�|ֶp�Jǻ+��> �٦Å���֠�e��p��xr��؀b�N�Z	UD Z�^0��T��������^F&�F0�)�D"��瑄�������Q��lIF��_gb��h-����L���dE��m��=(k.��w֢hI����{�ٜ�p���&'�*_|��YX�t�Z��vy�*�I�"��6u��"��g�����Q§�\�4d�
c�8�,?�g���>j�}�vS�����A@�A��� �T���7N�![t"�[c�qv�1?w�la�.A�<7{�q�x����엚�NX��'?\pޯ
��!�ҏ[ s���
Q�qhދ"��ym���˯~�n�c��Ԉ�<�Y�<��V��=�����t�{�2��ߞ����p����!���������@?;������]QZ߬�|�Br"��VU��6�6��쫢��݊�9�8q���#�t
1�)�Sw��a�UZ��A@������i*����R�-��#���L�J�F@|�]����	�=U�?������X�h�آ�V�G���nE�PYu�����=&�3��������m� �����)��J/+�f�.r�`���|���H��`漵aE�|�8#�X1v��g�l�/�W�?��|����P��%���c�F������G�g&M�%R�|�xL�L�q��.Q*�����r�5 �_O�O�T��Ts���iC�M����y��i����d寡�-Ɩ�^�F���Y�ɫ��<�ޟ�[������5�R�;��+u��Ä��"f5D��E�4����=1�#gz �� ���2d��"�J9:%�����*F�����X���$�
��>qُ��vJ"�!v�r\����͘����@�5Yr�P؝��*�{���vI��,����	rIl�N!�]R���,5	����u�zxW�*\6q.G�/�z�߾,�\95%�wBz�DB�?[b���H�f�N���۫����I�qf;�������HQ��n�4D�)I�W-~�?Zq}�N	����i��[�1ʇf V��3f�:�_�ۆƕXdsw`���66�MVk��g:�R�U�5֣�� .�	���\��8�G�(^�=����h��?�5P��)��馾K+/���oN��r��Bt��ԭ	��B�("A�?G`��uf�Fa$��_	��A���GvΠy8�M�8,�el3�~���/��k�2_Ӧ�}Ȓ�ڃ�D8�~V���t�V�B,�G�j �� �&0�SW�FG�\A�1V�o���(x�wT$/������r�x�K�[�S��9��t�'�2}�q���[=�6kx�)�r�WC�L)2�}�5��%ս� ���&��]pI��Y�*�s����&�	�?�*7�V�4/�\�q�{&�L�p�R;�2��� 9��1Bd�S�D�HJh�[d�W�ȥ��\��+���������?���M	���s�X[�^~��~�Z����Gݬ\���Z_m���"nm����P-��*=a�`���j
��n���q�MK�O�sV8[�	��]����l���3�7���k&���ӯST^��ޅOMW�[5���	C��"C���w���I���o��t��Bg�+ş�ퟸf
V���c��*�zUѴ�
ǘ"��3BS����1�Yޥ�H$H�zg�Mv�6({�9��i5ȖmQi��"�iK�.�����]Tn7K��vܘ��ٶ�nEj��oZϸ+���Kͩ��DT�~��*�
8SCtgH�)��y���������6~'����q����^����͗�Ps��K�����k㱣<l��m.1D{��(���j �uǭ���]����NuJY_�Q!���8-c�D��F� ��0��Ҁ�r�n��F�ľ�u+vڡ$������!Qs��W��{|Va�*���`��d?x,�<YDBR	v���4��C�~ec�L}��a�H�?`,�_D�j�R�*Z���EuM{M����W�x�1�C�~�zvF2'Fu�Pa������W02$a�j�J���%6]E���I^�_�+�#����K�N�"�7��:F��+U�P���Ԩ�r��c,�I�I�������~��Td����>���/��g�TH2���%�O}�Q#�����tZ`}~+��}cU��C+�s�Y3�*�jL8�_�hƑ��D[O��������m�������V^ԟV,�#�
�j���4����7�Rw��w��bZ����8�5�z�)���3���o�ߛ�91�{֔2����I�,��x�VV����E&�����<�iBqD�1jj ��a��G}Y�l���� W�����M�:��-�H�R����!z'jȒ�b
�88(��S
v�?#��̒��f�T	!�J��8X,�5�FqG�G�� c$����(6	/[�ڛbmk��7�c�����9�$d�'�x�[WX*�5��0D��c�2T"Y�P�lk�%E��bR��3<�/�ca��5�����+� H�&��Q��m}i�z�t��h�=H�o� ��E�(9��l�¦�؍��!��{[�ӫ}�?�a�"$�-S���)q]t^��ΏYA�\y[�3*~Ցݬ�`nH���}������e���u� ���b�l��ՠA���s��`�l��_����|�4�C���X%~�iV�Wʌ�9�܀��i@��c�Dk6I��)�G�y�O�-[�f��bl��>�*R9k��6떊�L��	�˝�3��U��+4�!m;+�3 	NVM"�J=��VC���78x�䪂�2�@Z�0�i�BwV1����?�F�Ǖ����� ��g:�Eo��^�8!M�>z�[;
���j�"��*>֛�
<Q�	�=�reԮ�H�q���*��B�L􉘑�[�Dw�Ġ�ɾ°�_}a�k2(r�:>y@��a���Z�d6��0s'�!3aG�8�<�ތ}�(3�""N��3A]\���gN��%�Ƞ&Pi"��MFX�>t����_nI)f�qCD|c|[�]t��p�j.�n��Y��L���/,�ai�3W�ro�1���9�L�Ld��O��$sj�F`�Q�q�Z�j#�P���$�J|��/HV$� q[�Q/���b�>�7�Ӛ��dy��]El�v��KI�?��Z��;V
<���&��V����Z ����:�����| /��_6����%	���܂
W�V*�>�y-iLV?J�{|��/�-�\R�Іø�B��g����*�!H����S�XA� )R\X��Wt&�b{�_�pKׅ��7Vpѣ��k%���[�DA̺Տ�9%�����~H� ����H��Gq��$n
pa��P\�ݏ�8��o�B����>Rj������r�M���sT�Ӧ(=�77�ls��@�<2��N]��*"�͚�G�K����Y�0RG�:å{#on#Ⱥ���h�I*��o��~���Au��x��\���+��k��5\�q`��z	�˰{�;��n���>��X肐��U�R�W{�P� .2��OE
U��#l� &+?S��LU��X�ZY���g;�4�����~w9g��w�����:]s��E^�)2rl@g�F��K�:���܇�΍���KG����Eϯ�'@Ь$���^��!B�]A},8v�tѪԁݜ��źoO�)~�>�����H������A��]���:��p}o]��G}�����}q��R�����u��o�ۧ��H�>g3�"y[��_l�b2
?M?$߷u��k�'j���x�p	�*���dp�Y>��[o4�K���nM� T��s�rA2���eA���e��8!�R���������;z�l�°�s 2���ɗ�vj�'���o%l��^(NE��'��"�l�CƩ6���D9lz�@��r����|P;0�Hǉ"��UG�2�H�H.��[��C����G�* �� �Ъ4��bm�#mnS
���c>�.�pa��n��'o��s�d?�I�C{#���S��C

e�{����0�o��3����F|m�AU.�:��(���fX����F~�$]�"ԬyNM7{�>Ѕ7e~v�@|^�P6rˈ��@uv�m��T�Vӎ_`����Y�puP�.��y��X4R������u����ж�E�a��4;�@�4T{@���f��u�3�"�w����M�eēߝ�� U�Bk8ᡘ)�\�B��j�"�x�&�麾�=w�7��pl}#Y�(��_M4��aA���A��"4Ľ�Z�A�_��.�|a{�Ss��$O-�3܎m�ʃNĝ��)��aR<������6���Wr3ڮs�@�\�Xہ��4�@��X�� 1�!����HF� ����w�_��`��٤�h�dO� �FrC��<��j������li��@�����Ƀ�}X���+ݻ�OV:�$�5���8�7��"�0j,�
���"���X{-�g9,��6�[Z0د^�̃ls>��bf�]>��w���f;��3i�rĒ���v�	H'�T�a�77���[��kA`F��t;�?��x�9B2�aK��|�^��0�r��$n����@�+�wWxo&K�1�I}�aL���F���7�X=Cxa����,�M�����a�0�yi��(6}�`��X�r��.�u6c-K��fD"�����������~��i�o���Q���� 1kq�k|�%�� 8WI�MyǠҁ���hȦ�����ǿA���Տ	1Y��\����q�?�]o��G�my�*SNq���j(���ӡ<z�X�J�Bb�tL��{[e��kT����<'�Y��!
���I��s�tu �E%3����R�^4���V���$�0j�M���Qb��H=k��ӽ�="6{��qr��SlnOG�^��puG}��)�ͳ`��^��z�IIR���К�̞A{K_?����1�i����A8a&�
���(d���Ct �ȹ+��X�c������2#�j�)SI&�L�4+{�L�m&y�>�����}��E~g{��|1��,��'�D�Z1��q�ܪ�V�L��г#ST'8����
�pfU���@:Bf*Z�n�1��vK�Y���^ZK��� ���D�2�)�KC?�ߘ��&��P	Y���H�91*�����u8�r2AEuK�Z�P�r����Pp�/�h�3D�x�PA��C��O��N��Q8�%���	p6	�/��W��J�E|�:�u�fh'��<�Il�Bj8\_���<k�] ��:�4���qdYa�"NtG�m�a���r���a�u��)��N�[E�`���c�׃����pp�p�9؋$t2=?^9�3�AN{Hw�Pĥ�1��y������[koA\�r�c�Kw���4�Im��&÷E;���Ypan����L�K'G��b���2}`��ae�!���U��@y����|wG��*������c�{:�1�+�fμ�Z�W�͏H�%Н��G��.�z7�Ƚk�MtY��h�L�j����0�^n�~U��4`�)w�O�)�<�$stT��-E�)Q
��R�l��\����x�N����X��10�U9k1�fn%
�����8!�y�Dq�d#��sQ��mh�����VS,0@"5�		{I��v��N]h��B�2�ϷMU�rjڐь.Hj��H1l�!��cB.��I��/�1l�Rۣb��1�k���Z�����R�}�><Iuk�,\Ϊ2ٖEh����e��c͔B�.�\�ko�w�T�p�M�Vk;�w����7Na���H�p�"���W��?޶��E����G��>�3��y�你��r�&�\������P���"�ʷ�;;o�(�o�W�4��e�ּV"-#lf=~�ڧF M�&r��J��"!���m���"���v�v�z�����#c��JK:kV��]��WW}����H�旖NW�>/Ϥ��7W�^*�D6�GI# ��챩������Q ٲ :�����9Y0B�.9	���N��Ύ�5E��DC{ܴ'����79��S~|WKy�V;�7�_
AK���&!o���'���p��1��9�ʝP�l�%���^p"�ѵ�e�R�������)�s����pB�x{}������G'Jޤ������-��3����ɞ�m@��]`��)�չZ����[��E_{á��X)�-�VWF8�����5O��5�"�T-�+�l���cKǷ �P��Nٶ0���υ��hh�đ:�$�0�\�� w��^_�,�|"�J�H�/S/#/���\!*r�|��sȌ%��=_!X:˳�ƅ�Z�(E�Į�Ι_����:Q2���dG�B�v�>3݉���l�m�b3�A��N[0l��+��r^�����2?ī3l��l��Yc��*�i��v�(s�W�8��tW�?L�TF�ٴ�x�ӂ�M�ͺ��3����Q��-�Տ�m���뙜��Y�7�+���˥*AZ��:k%�`��O*x�i9��=��nVKݯV*�����_�o)�e��&j�9:�kʳ,�%�~"F�&�j�Ps�:9s��������:�,��uUPx!��Z�Zk��0�I�l��V#`��8�@����J��}��� B��Ж�/0pz#��J�1�1!\4�q�x�F�^3|�' �r7���-׬H�;#PQ���u���}��������(ծ��a0K ���v?���;��*:Q����(�L�Z_��:�����G�<���˝�S���}��u��L������`S���HC�n<J�����V[O�:��՛.'�~4��;/��|A3����C�~�7s4?��������bdʙyA�5��e��
�Hzm��8�l�Dm�7�g������PEi�8�T�2�;*������Oʃ���>���0o���ŏ�v{L��S1f�l8=S����i�x$قeN������+K���Ϫ�*H����s�0�X�*,,W�'��a!(R���@�y8Mބ��t��l44�Ҁ�X���|p��O���\�K1��<Z�cRҢ�d�DG�d�@ dR����qyhC#aȨ������0�>q���	��	�zv�Z^���	f�]H����[����B����.�<}��-C�'��	w�K]�쑉�&�5!rJa��2�*Gh+���X]O�8���˙��Zm*�$$!)���v��D�Q �fIEPe�n@:V�ar����k���ؼ���𡃥M�8��E���Zh�3� ""�B9�������_��a2ـ"�� d���G�����g=U�I	��M@���1��
�i��q���M	a�>]����z���k�4o1��^�|�O����h�s�fn����l8�������6	?X,2�[unυ1��^�θ����w���F�s���f�ڿ��߰UFB�ۤ��	���_�ⳍV��B�&�Ş��7_"񝻿%����c��n�?T@i���Al�͂��������~_�h���*/�þ�l}6��{n�]���H����T'ɏ)� ~��y�7(%�T��jY#i\!8Z%�˥�a�G�Q�Cs1�C镒n�;���3.�=���w~�O�,&���rÕy��E���t2brQ+q�gH<R�$R�k%�a2�xipb�����s@��j)X.9���!]l+�NdV�Lޣ�+�=��<*��l�&P�aݿ��vܭ&0��J�F�x���=��Q���f&S��`�ب8?�_q�f����m���$@�T#&d���f��4~�h�_O�t��E�1�QP������J$"�5R��Β��Uf��V���hVJ�!�N��br�R�{�˧�����{V�W�w����84 �"�tN��� p�#-�@�v ��o֦�#�9��\v�#�ܞ��+�f�Ǜ��eE����ہg���f;*ĩ7��5� ���l��&�?�{��C����`B���D���;���7*� Gh��eҭ?�H�BQ۳"�k�C<A��fB4.�_��ĪD�������Z};8�=��@^X֧.��x�?W
c"�-�Xu ��v�{��K����0�Ԫ��
�_GՊk����4in�=]_������VM*�j�ZF��+���C{�����\�lԿ�m-7��3�֊۞�?Y;��Z���e	j��;�'_NEe�c�����?_�ݺ�����0|t��|�p����9C �B�_
���]ЃZ��+vw!�}�q7��<)řͺU�!����L谬�8ok
�Q@����ۨ��%��Ī�d[E�3W�&��&B/D-�v���/t���6�3�&܇w��Tr�
�{�b���p���5 ^�R*;~�8*�Jt�j��S��mH���}����gHKO�,���Ov��Wp��{�d�|�z*#g����T�\ٽ�%��qw��S7���%����eZ��;��Y1�V�����J@4}�ζ�}�2�(`��@Ӡ��'k�C�߂:#=�1CS��߷R���\x�����J{�2���2���]����ɕ�$�V�q�AaSi[x{���X5"��6���_���b]h�>�р�n�`�Cm��X)��gT\5p%V�S�A�ih�%���"R�QJ�\����}�z�>�Y��aS��Ғ�B���M'V;��7�)�����*~"nZ��I)t���J�Ȉ�f�Â�-��D*W'�d���:A�{aP@���w�0\<jp�n*���?�\�����2�/V����h|��
δ+���w��l�{w�N�xo�D�s!>���0R���=���(����&�����:趋=����^���ha �L�q7u��2�3���
�*qR���S�����2��{�g��8�,m�tj�l�5KVUMX�T7�'�D��wrV��?�2����#��r��M�䇌�G���������~ k�S�u�Cj�x��������SgV�<<K�v|��Z�ۗ��*f�#��{��%b3"�|b(���l��l9]10v~����M�M�/�o�" ̑���:�hZ���J�XͰN�'.�����l��{��8̻��rr�ؗM)^l�n��@֍4Z	�^,��
��b��c�]5এ�9�S��1_)�=�cv��lNK����t5�ix��ޭ �G�-�9�?B���.��[���1_���x����+�>_Ϲ�B�p�mB�}���3�˧�eh}��6+��Z����M>�(�8��� ������Q�@�U�������1}�`$=3ۤ��V�Y^�9��y�V�d/j��m1�n:'3�Fٞ��&�k;�2�ˠ8��˿�ѻ�!r��u�{y�XӠ��(�Uu�v��P�I�X�Ҕ�"���^\��C�}`o{"�_�u�6���I��g�4Ugg�3\k�;�������IR��l궩,����M��q�iY�8����#W���w�������^̮���wC�.v�/�\d�Y:Ҷ(�!&����^-^U����|S�`�T�����$���#����5�n���t���e��Haی���,��I��97TN!5MO���������If=*��wQE4�*P-�u*�6`A,���i��~��/S��u��E���b�g��dn`��G���A�JS؜^�+ڐ'�f+QI.z��:���!h.IQ�?�lW^q}۷x�Kj�xs5�����A�K%���8�5�T�"����~��]I��KJo�C�b2�[V6�q�tg��?��������ڸL�8p�up�6U�` �~�O����_7Ɔx��+9QS>��<���oa�4 �@��������+��2�#6@=�^3G������ӌ*tGX@��L'����0�S�z���"`��m��7��a��͏�,��C���� Td醀?UAtA�YO}u���b��F���űq����젳k_�y�P��G���Cʒ�b�����ұh�o)B,]opq(�Ԯ����������/Jj��x~m�圏)#* ���	"�j�.�S�� �I��X(�+���Z�ǹ7���S�T+
s.�d��
o���8�N�����g��?>�h�P��|8^����V�ʖ}�dČ� �-����дLu��%d	��bs�p1�s]�'����������D=���[�j���)u�$����~�C�%b8�;���l�kПh��D�m����[�i�7�ܙ�}�5��Jj���IAZ _� ��K�?�W���3k��D��k�1��8��:�]Pv��&��Վ��?��e�n;e[����G/=L��0�5��ǧ?n�gw��4�á�ٳdl0}��=��gq�S�{��u������83"+��(���ʩE�s��X���*-�%�������2�[�<6\#���]�BS�3Hcu4�U����a�n�K]`S���Y5'nC�ϋ̿�.�J{��Q�њm3���vf�����U6w4�s�e��\�H �o^���=w�������22�3<�,��/��d(`Z2���9OU�Δ�5��6�sZx�nL�bU��I�@	�L����1��On白B;��ﴎ�Ŀx�Pi��b!$�?A���I@L$L/�`I��*�O!�=�Ձ�m��_z�<�-��洲H�ckr'���w��WP���[Yڙ��M���\*�ie��[d�]H�}�wB�\�r��C�l�ɭ�x@3�,Qg���t�����+z��?.��?�ql�C���MէQ�%�f^�/t�NN��x3�?U�I�c��&�`5���h�ͩ��yV�o]JF�&T��V3	f��B>(�j?�#KN5n8��wLV1�!���'�A��E���ms�M;�lN�#�/�+dB)3�£wz�u eEx�46P�qъ�ޣ��b���Q��e@k��#�-��qV�so#8�u�?��t���Uz���xӸ�� �©���a�����)�w���V�`�q 5"U҃����K�q��ّC����KEm�QP,i���>�� ��N�j���SQ�3��F���.����cP �{B�׌�׼V�K'	Pu�?�7j񾵔�C�5��PT
 ��Fq��~��J�S&�8��R&�L���63�$-/A�~-�ci�[4���[��Q�B�f'9ه�\���~�%��gM�����o^��T�O.þ~@���J2��]���]d��)9��P�$W~G����/">YCs�r�Xk�q��<b�+���u�	��k`u�7KΖ�^:��D1'�s��C�F���Ĉϴx.kԫ��*���*�f��#���j@jӥ�pL�c��{sG1`�#����^<o�����'��`0Y�$ �Nۣ�Y6�GN�0�kX&1��}]����H*!����|9� �"��V`{�n���?��
¿F�Yn�W����l�}J��ǃ��&}2�:�e�����K[�I$�?�Tx�?;���!y�IU�XaǑgb�A0�Y�H�c�m7&O,D�ڃ�j�)	�&A���	x�h����tf�tЍ�3_A�Q��6��?�=Ԫ�OƎ����36�đA����x�{�^j�nܶX�C.��ɏ彤Ya��H���� ���D��d.����:m�`b��=l,=��@d�f4���%ζ@��b �ʟ�
���$�xq63�7i�}D�yIY��?Hyș�Tb��yA)�o�v�8�U}�z7_��Ww��̌��,�c�`B�HS�N�iu�B�d���gy6_<���}�S�8���|�vÄ Ζ�K�<�����?�0���ESNc ���6�?��:�]� �_���0l�㚥�}�v��:�v�ܚ}G���_���� =��(kR�N��+�*������=�:Ē~��s:ZT��!��f��rֆxa�̫;7%��9�Z����c�AzO��6�Qn�nw��A�➒&��|�s����� 4z��_0<C�9`tz����D�/�S��T{ܟ=�]k/R�"0|q�sR������=}������Ӎ%�a�!����@�����H�cu�X_�ܨ�&�u�c��o����G&C�O�ЃG�B&�֢k��لm��XՎI���%�h�7�*v==��J�<,1cd�Z;����u����r��ubS���?:]gOM��|���FX;ǞA�1KŃ��S���5ZU�8'��P�2��
�&�u���{��YxR[6F���ax�S+��cDˌ�îA5���w8�c�m�;h�����7�6+��Yk�Nq�v����q/��+ɯݧ!�q�����3`סy�J(v�t�h�'\!���xy�r�s�u�L槚�f��Nc�O�F5GL	J&�,�k�kǀ��}Y*[1u�$>�"X�D�&�޾�n��a�|՘�h/u55����?{7z5�HFD� ���ߧ䤉��&O=�]T��CTk�(�q�� �&�?w:jͯ�H�`�¢ew������t]�8$8�jl��� X�b#ŷ�*!� &��	����E����z��M^�UhG	h�m�HG�:ٜ�T���9�-Z@���I	�}�9�|��[i�Ro��:��zը9��E.�T�FuTy'�̊;�!�g�R�I�o���G?�Gh�1�����	�|�q#�i��3ҶG4q��Z�~�cJ�c]f�,y���+��D�eD���U�9�ku!�*I��G
�/�9�ML�ZR� t%�F��Bt_�ڲ���5��e�GҬD��7jZ�P�mc~�y�V�q��3-�X)��ve�f���Z'S<s`�}Y�B�\ŋV�l�iJ�r��U�[o2A4@W��:#�{����K4S���hL�ď��6:�\��[�����^#��r)�
l(#�]��_ja�j$(�̹sx_[���Y4+��V�'�fZ��Pך�ʘ~��&��qq�b����9�:���<@	���u��ς�	�N>�!8m�v�k�-��J1��Zw�ܿ��q����>������?�c��0�'`뻥x���!q��U�m�-N�������� p�>ĳ��%�(6?n�b?):��%���aI�8�4��%W��q9��Z
/��׭G�R�2�2���@j��W�_3������c ��KN���e��nZ+��\i���C;E����7�B ؇o+���s�������b7a	�Y$�}�_T��p��h�U��H�T�T BǮ�<�t��N�y�3c[�K��=d�\�7
��Lc޸C�C�T��g"�Gv5ƽ�B��_�ǵܦg�F��$��acL�h4����*�{���"���M�]hF{}��P�b�q�GܜI@o~\_0V��;��Ӫ�9�CBcǅ��Cq�3f�|��(������D��/�3��>���cf�?`MiFH�{-l��N��0�"CA���Y����յ67�����P��:?Kx��nj�Z�<��ݯ��{7~7WB�s8�ó:)�vd����nB���Q��������������w�0�Q���ոиl��9�Cv8(���ދ&���m��0RC, �;+2�r�vaŨ���R��x��;e�I�ۥ�d/�銷_}�+���ۋ+ɯX������*�,��nˍ�0X�4!�S�SZ�겘U�Lɩևa������c����)(�j�Ȇ�'�^_�20�w�Iޖ���R�;���͘w��7�'v�u��W�7���;�7��M���Tj@�����Fd��_#%i �_yv�S�m��h��Ld��&�m-�蕑e�j%��e)!~%营4v7q��VF,o�>yoa�`�-$�*t`�x;f�� ��A7�^��.
��p�Ґ�1ȱ�*Eiu��T�sr7czc͎��(9$~�����-����$�o��9��?�c�ϓ���˵�ֻ;�=s����ߌ&��N�؈���F�H 
t�����Ѿ�-�U�ڱ+H&�f4�}hھA�|����L�"X.�P�%)��&���+O����H�
���'(Z9��y����oU�M ]׽��@A�/�%�Q�3G����c3ZR	[k�S��A)�o|��|�N5E~:�U�|�x�JѶ�vi7y��g�Q�ᛔ�PҝO��EI$���.^w�A��ݼ������T�����.��+�dQ��/'���Og�W'RU��4Ḵd
��(ȫa�=PK�	��(�G������4��)]V�!:�x U��O������:T��~\��9�2�L��?U��_t�P�Hp2q�&UE�m�K�.��;���%����
�ۣ_�7�ސ�<;s����Ln��a@�����f4�[LsZ��d�Nԣⱬ7>�]{"�����V�~lܨ��8|��Q�Z���6�5����C���9񠩄^7��q�v�eM�T�<|����0��iM9��Z��X�p�;��]����
1�3@�{9�y�r>M�������[m��!v����:U�h��"6jPzg�A�G��:)���5E_�y]�!�TF�����v��س+����M	�'�xC��I�	�����5�g�Yvnÿ�w�d����-`�[%�7?(�J��q�?{0���Ŝm��f��Y4��9��.E?��>!�B��FR_�m���� A�\�po�xh~���`r� W��
��?���]�9z/
���	T����Ѹ>3#�9oD_���[�R�@q\��c)���NR	l&٩���w���+G��M4E�ݞ�C+N��KQ�$�&e��v�V��C�с�I �9,k.B X��yM�WHy3�/�. X�\u+���&��(.��2��Z�y��[����Zq{�0G�tJ�z��}�&��/`�S'-�/J�[�F�`�*.��ij1km����ne}_r���U�z����\r%�2�i��Je���������%������ovC�\Z�b�ķ`�rǳ�W�Ko5b�J�����Ǯr[�T��l��6������/c�����puy@����F�$��{aC;������x���bE�7��;뙜���2��wM��ò�8�+Er��Y��"��<1$ϔ���cGhe�����<J43 ��z�ݑX��z�E�"Q��!�첛U�џv��rTZ=�� XB5�TL��3,�ؓ���A֕jg����9��b�]1�Vo�|[N�X�\�a�l���8��[��s�߄nc�4�B����� �E�ǰ��Hh�Hg+��C���nJ#�	�BaLj�3�&K?Ѽ�]����(#��o�1�b���v��N� ���VדdϬ�G`g�{A�٠A���B)�9��ir���"y9W����U�j�ȷ���r5���5���+�ņ��5����?m ���}�I�L�2��h:����W��n�@���-�`�ټ
�`�Q6%�ݣRt��JS��m�ߡ�<Kq�?��_�.�&L�ԭ�:u�����A6qN�q�g-{#,�Y��,�i:�C�BJ�^bz�w��<V.^}�T�;u���3	� � m�Js�On����{�D�L���ŸGR�|���S��Wms���G�֠B�h���wk}���w7MS�=��M]��@�Xى$M�A��s�
a��j(찱L�`:�f�,��.^1��]"�=Bb�+�%Eq���&�� zM=Iz{XX����G�l���f "o5�]���H	��҇��ƣ�	b~������N����$
h�����Xx{0��#	�cW&�'iLӈ�G������PDe?�Hb���LC{V#K�F�.��BՄ���p�ߴ1�]1`�=�!�i��g�Q-��l���8�V���= ��9Tn�v�A�	C���ͅ�Пy�����q�s����M���Xi�*M�'���T�)b�W�^h��چ�IU�ZUۋ^�D7,
{;�j��@bF��
-��O��J��3Ҋq�q���-^��XZ2Z���u$n�# 䏋B�n�b������ؼ�ݓ����P#���A {�d<��x�����.��ITXͥ�ǁ��Nt�bڿ4uD��:0�D�9ay�A,9�Â3G@]�07�n�ٻt�gm;Z ��N�.nN����$�N�W�����%�i��@0XrǷ��F����;�H"^H���-i�o�9N�.��,=h���"��S+�vQu�\3������͔��\�h���_/z>=a�>SMOc�@
�j�H�o��-��Ng��~�O�]<U9�8���u0	����PEÃ���S�d[f߶�L}L�}��C}{x�����!��t}O�_�e}�"_&#�5n$�RX>�3��� P��)�/�1�uzc.cق!�P ����^�JA�J^=h�J��4H��c��<N�����V �.c�BEw�@�4��	O��i�%d��,�3�vM�΁v	��@����p�3;dìak�m�p"[Jv�.�L�'���ʼ�#�����Ϡ.�i2�����E��	>OU�� �.{��eD�E���������d���ߡb�(l�<�B�X������^+&�2�Q�1��N��j�Y�u�.�ň���G���)��*�@�)�+ᚏGN�s0�[E�"x���exS�� Sl����"����b�[bęM��C��B����E��SIfV��ԅy��_���uG�p��4-���0N As�.�"�8�WŸ�3�c?�����p�_8BYMb��q��7X�d\P��� �GT4|l��U��>Z�&���7]��}��	��C}�m�Y�<R�atN%�>1�I[�:���f��:�ث�eZ����?1F�b�Ck!��¹�X�m56�2Ѷ�z��n^�+|�'��H�_���E	eO̐!��cB������i����Wk3ꐊ��2��%���קD���p��9+&�&�c5�����`
���9Ƿ�s���و�2�r6��m�����8��jo�kՆ�k���3{%7�s�&}a�^r]H��d��uɲ�]q<� |���d�CO��.W���ְQ{Y�LM��
�"��9F��|Z��D��I��.4{��y�u:��C�1v�p�>i2���`�ͬ�_	6�1�m���&$�7k�����,���S�v�A�+�M��T)�,��<��D�]�K�i����E�{U�,��.� ����6g1��[%,����۔���#�*{�L��r��+���ӂ���`E-�4��i2�Y��]!��=A�(��S~�+�>��G��E�R�T_D�u�k��E{�t~44�^�����n8�_ϔ��Lg��B�#��T7B+������=�˚��~D�,	^27�i��C[�����t�d�� 9 ��ŗ��	)� ��DfS�SI��x�~�L�&׍�V���Z��-�&�f���H��l�;���Ax���쭽�2��ʖ�4[|KS�Y�����uo܅:��яRg!-�a