��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&Y�%�ddؐ�ပb���p@}y�| ݀'�2��DuE����qs���E�);s2�>t�c��L�/r�L*T�4X��O(fV���,��㳒d�<靷�2.��],eK����w���Pn�Z,�!cN�iN�ɰˎB���\	!�g��JlI��@� �Oi]�W�?�v����DL��,�M󊩘BJL����d��-�I6��o�]lɓ�3%yx}��+���l���,��%��pB���D�t�B���� �\���f��n	�o��ᵗ��?��,�nq�Eq�yp�m%E��8Ɂ�r'��[��,�kHL��oE��$;��|���Ii�t}k��(�e�� ˪%ׅ���y�o
��>�x�1��{VJA�d���t=���VVtF7�iRb�=6
k�>���<��oq�����r�F��a��_{��3L_?�B�dV�@�7(<֤dXsVڕ������f�6�mX���'sq�y��|x�[w*����ƍ�x!��#�'������3��.y����!�g^qI���wħ�ׂg�'dA4�w9�u�z���]�7tiZ�`��z��+�Y���'���rc#�%�M�:�J9AN����ȓjB�8��O��*������Յ�ּf`\�x%�ע��i� ����c�M�]X���w��2ۏ���ʅ��F�w.Glz�s'�HB6����1M��K��l�q�%س=��iN��O�#��N,��I�]�?/�79���O+��.\`�T�jzWC�
�@�3�%�|����^d���$�y�����9A�����I�I�2=�1%B��<�,��$�� ���LyQ��~�Eg\�ALO���" ��/���t��%�~��\q}N�1�n����f�[��Ee,�goY]�`
���`7Pp�Ͱ)��D�W4���4�������7)P*8����d�$Z	:���& 7���Gצ��<�=%���$q��x��(���E��Z�5�`�"@eVX[׿*��:�Ui����q�֌��G�ND�ۮX �a�?fL�TJ�4�]��J����4�n"��L��v�9v��+�;��IuM�ψC��㬴D6��`h֓w�7'��պ˾z��V��F�e� �?���A&	ew�(⃰�F�q"�.��t9����y�f{�(���d���! )0��O<��ht���O�G��"9�Q}mP�����:h���f�������v�d:Z�CQ�#.���ŭs�	LvT|��}Edy�kS����-�q�=�9���я���<	���k=j��iTo�������=�m��* 3)�n�M��xf͖T�����_���dZ����~������JP�u��0|�fŸ�(�jN�8b���cZ��y��𲢰訝:�l=�'8���AnW"ό-O�M��<c`.��κ]A��dZY� mQ]�Q����w[9K�h��Ƿgi��z"l�n����'��7]<���ґ����Ǡ��"���Sdx�5��rJH����Q�郭N�4�S7��~�.����y�X�T����b1a$��P<���|3��C�j�@]z��� ����P#&(V�4�������>Yz�r#׼>T��`�Y���̉�nM�%S�`��Åw�l�����n��.��!��v�r/
Gf�R���d��&m���3<����r����vv�q|�5��w	d{ؓl�,�^c4�W�x�J�z)q�%̫�9�1�wW�KAVP������������e��Cl*������b���fM��߻g�
��d�*W��b��~,f��Ȕ��_������ yV�	Cj4��4����рϕj �6Ko�0V���K�3O¨� m}v��=G�&�s�3�-�y�ȣ�-��!YVk��u�%%u�6��Ѯ�ݸb�\G~�����A�?��wo0~:�Uuf����Ƃ㥝���}e�iV@�z!���.��ʍ�y��-��lk�e}�{�@Q�_���E��9�&�3r@�S#4w�p*H��jZ����6�����6�|L7�W���aT�i���J���E7^&a�Y5�c��8��$�O�P�-�i����*����^�#*�P��suM�FQ�D���i��m����(C!)� �2��ҳcIQ�{����WH9����5p6R�����!�r����/�3m>o����\���"@'�<w�]��%�"��\��Pqb-u�ޏ�>P*�lH8��_��%���H�eq��7���N�&�\E����G]mdf�$ڛvхl��?w������[i#Ny�k/���,���9�ziv ���B��WwB��<�4Y�� �H��|�����2g��P�J��Z����4��|��$���[��m�F�����O�2fQ�%1`]���K�yi�����470������
hR7����M��5��wJI�����7H�)Q<������o��ԉ�ԖB��@W��y����D"��#�Z~KG񾚡q�NR�O{ ���˫�}����d��]9O�H�Xf;�M�T���;Ɠ����6���^���6�j�1LD*�O��4�f��#����`L�vP�� ����>n�E�2:<���]�#K��}����=�h����
c�X�����Ma�5XBn�����ʦ[�� `㣀��,hdp�����_�^7B=�kn)���o�ǭ�m�K4B��.�meҚ+�͍�o��v¹��T|��I�2��y���v�>qx�:��H%U��qW�Hѡ�cl80z�8V��#'��@�,-C?�j�=�sSh���K�[�CQ�c"It�~��K���sd)+R���v�V�I�c���9m��[�*~��8m�v�ym��5���RN��r�:�|'�f|3���l�s�-Cd��/���hf?#o3v��#�?놓�����'���(��e���0�H?0��2 �Qi#2����0�)'���,�ꂝ��^�=r~�0"��G�@d��{*|χ���&�\�P�^��ji���b���h���ӭ-h����y/�����lﳖ�d��@�w�A��vGU��Z�?�;�"ה���F��S(�r�]��:����N�y�׌]U3�����lB��l�����gw�̔p5%�,����F����7�ѐ�q��rk�u�k-�v.% ,";@�e�߫n�<YTqIf�f�k,kelǬM���~q��΢�4���K�Г�l<õ����'ܣ+^ISV����;_=5
&��}v��C���w�~-��}�F� ��ҢB��L���O@��B�*5���!	&"�ߠ~M�MZ�9'4��j�^���B���tի�?hE
�h�<l���Ք 4�{�v�ǜ�q+�3Һ�Z��S�v�9L"$��H�d�
J�b���\
���Z�#)� �5f�|�7�TL���m��f(s\��9Yk�� ���H]8��h��]
v"ct|���m3�b�z>��f��H�ph��g���7t�Pc$�hdMO�*_���vYD&�Y|�����m}O�����.%·���jM��;�oZ����å-�bژ��H�<�;� 9P�#@�5����^�"}}���<���H%l�T�=_u�
��C�jg,�sP��$4�!��>`����/u�XS��J1��R$Y��W�N
J��ެZ���$W� ����zXTЖB��P���C�b��0k!oi?�B��T���x���鵙h�XJ�����!r�ՙEX���95L`/A�ة�y�f��'��~.m��,3wL(�������op�{�AG�R<�#�|\{�0p8�P�a'�z��MNY9Ԃ2�xC���y���f*�JFt,(H��=(q��)���L���2�' �S���X�8�=_��������HSy&�;o~3���Z����u�b�0���$q����Q�Yz�s�Te��];��� ?��4�|��#eS��Q�x:�)�7tp`�{�����tn��S86���w���N�Bg�e
Z����6��s%#�G�4�J��
f��8�H��D����c|�y�,��E1��@�d�u�oN�W��g�A_��0З�Tbټ3T1BJjkn��%��x�r�d�� ���_(�G`�O��j�2o�^
F^BW���zN�
�f|ء@��\js"�v	^^���G�9�a�Ҟ�1�)�ALҜo��2��ݎ����c�$u���,�u�1��[��TS���7ClӠhe4袞�.���-�ĭp�ԄR�<
��*�3R�f��]�zok��aw�k�lMߠt����۷��s���=�B��=/�\�w�?�8�
Bǚ��\Ԋ�,��N�3�����O��&��N��ˉ�Vꥎ�{^�㝦C��5�|���"��~���sq�D<D���f��g�p����q��B8˚��>����zX	�4y[R�N�?�U>\���"�#�*���Z��6�#o��#�����RJjڑt!Y�T #?n�Ni�t�z1Z�{6
�	h��R��D:A�hhURgY+\���&�� M�wr4��|*+��Q��G�ݕ�)��WP=��= ������*a�C<��]����Eb��ūw��_����d���ev��Q^�f���S[�I��XV�� b�K��X�Iun�?��6��]�gk�&-�q oR�9�� ;o�Q  S�Qm��-��pY�aQ�Y~�t��`J��ǩ&��{B��u@�.^�;��&�=�	��BϪID��x�]�����w%���1t�C���AU��Q�]Z|����V�+�tZ�`�DP����s�`E%!��:��wv�%��?�v}U!H'��ͮ��	Ο��x|$���9!(;w�^�����w���j�,�rUϫ}���T7_�2��'6�^)A���T/�MJl��*N}+j
E:5��C�%&:��Z�D�q>κ�HE#)����%C����� .�P.]�>�Mߨ{�A,���B�ٰE���1i@F����:VR� 6wU����Y�?@��)����'KPV�N3��? v��C���`Jn������7����Etr���l��'-?�h<WM6��p?�����0�����ݳ�//w=BHOOZ��%0ݐy�`ժ�UԞ������:���+����GY�w���EX�	�;��m %�ťV�+IS��92 �N{�haK�r��e�d%�m�ζ�=l��x�@ ��-�nM��E�}� ��O�7�Ϟ�ns�D��EDM2��ޤ�����G�l���,"3M�	��)��;�P1
�K�]R��b��ܜD�.<\8�!r� �.�i	b�G����F��
i�� �l>��Vp�V