��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQG�.�����=����y��Q�{� ȑӵF��� [Lq9��C[�KI�l��Cq���>y�B�%:̴>o/mw�5�'�H���%uc�]�c��oI �1:�Y�:��N)"q8E��]���O�l7;���|u*���?��$�,e:®��~���A�q�_N]�Nye��eIJ�3�݈����e�4~��z���
��NS�����+.ߓ&M�b}�6ڣ�L�o���1�T�u%��y��-G!�Bj�ry�J��(Gn��}���'�e�:����颹�A0b���&�j�=��PǿR�`�2%>��dD��َ��F������$�tU@������'�H]LY08~I-��䓝�9y��2�Ք��h*�Ktb��bJ����x�|�[���TN�K��k�PŌcA�B��P�!��uiߎ��L6]'����f�X�=��D�6���:����h�������X1�B�����M�Wo�S�m�"?`e�_�6�߼���uC�>O��P��r��h{�̵�c
}����=i7��43J����}�JT�*/��F�C��?{!�ȯ�h$�4Qn0�����NN|PxY�f�%V�E���(�g(�eG�ܕ�y�#$K�j��<k�5gpl6�v��<P3v8"5��PZ/�+Uq��H��2y~����ٺQw��Y��'��Dl����s�f�s3��ڃd%^�k���4�ZGM�g�x�-�վ{�et1�)��ǟGV1��I[�a"8�<��:-8�*'T����<YJIr�W}s:8DB����H�����]��Z�@#��f	�IH��;q���Mf�/�[G�h�`��}��J01Ϲ��rR+!�;:h5T�ٵU
��'z�2<��˲��U��:R"J#�7 �(��bYL�xs��U�jA�u��RgOy��Xb��'E!�Ҝ����{63��m1����Kt�u�Q�%S���M��T0��In�x��k�˷$�p��6���wc�:t��	������hoi�h����~!?8��YuB�^�y�sAC�͔�[9N����(�6e�l��$��&��gi\�'A����Z�fWi���z�z�=6y�œ58	��Q4�� \����V_5�%u��U���|.;��T}\J^�YU�!�[�J�n�a�{�o���*�I_ѐ�f)�$Y�_�5+H�q����ܻL�l� F��:䍓�^�$�a�x���ip+S�3�T@W�r⇂�Lt�O�bJq�8Bo��C��ƕ�1L@��݀�*g���F�N�HW���sG��CVf�h���"Xԕ.��8f!���<���2��C��:��O$.]KW�`bۖ�������O�ֹD���O�o�^���T1p�J�\��6,�v�2Bm"��kU���Bn�Ϻ{v;�������ǉW��x��䔔�`�t3c#���n�!���C�F_~й���8���!>Y�yXK�k�?T�Jb}��b�r3�03�����BuR��<�m����"TXR��T<̓�!��A%�'3GI����f�fue���a��������&\*�Kq����[:�R�J�k.�s���K��<�/p4e�3&_��Mkh2-�� �
��HxW���.O��˰�4Cu��~��c�~�Ș�b9~[����=��"��h<.�5��Ubx�v($����x8�Li)����/�X!ٶ�����z�cXן��3fT,�UH#%��)=�h�05�I�NJ���io�""�4��1(5�&)�*�f��?�������;�Z�(Uġsb��U���s�a\�w��/�� �v��l�j�ǁ�Y���>���O����6~�:[���-��y(-�Y�9�(��Wln�; ��_�а_�V�3�A�T�M ��qQ�=,��F��G���!g���;�3�M���`_@�v�.2�;@���1)(����ʽ�.5T�nQx����5#���X��ȇmv��"�)	���%q0�G�D�*�����v�l�2��uyo��3��WW��:AZ��J#�3=�[̮a��Y��2?|`4���}qfI�y��@Q��W��/m���+��%�w�~>r�qz4�u����=� `I�ub�g���
+�P�΃:#6ljLfJ3�'K��'%ͫ��z�u�%�	d��~xJl+2;��	M��}�˂5�+�ȀP��gmQ��)�_��/��Ēc,�	�ث|8{��
j�z�	����}]���)�*Pa��%X���w��<{�ƥY`8c�]@U�!Q��6����I�-�/w~V�.�n6Yڵ)��!��bz�:��{�x�Z�%#��Hg���"9�S�����xV�<��:�ڻ��;�j�	�d��w{vV����n���v"�v[�"7��ad�S�0�1u���dD�\�s�~�z��> ������}�o����1�B>t��h�������[bR�����S!"��l�*���E:1AbQZ��~��UM���z���%���,�����6_�JuME~��7��M�i��?JeÆ� ^�����Xϭa���,ȓb2�w(SlY��}k�h� F�V�h��D)���g��oi���lj����0�VŰ�>J����&�:��B���uҵ5���l�g�3J�$V�?�79�)ӉȒ�H׃�wEĄ��w�Г"��q��{~�fX���j��qR�'��T{����5�Db�)Bh,�}�LW�@���X���^��E���sG
��Y ��>v���u e�7��5xKf���0D��x��ۧOpF�����&�0�0�@��aǏ.�7swB��BS�7�O���"�1^4�o�����+�ԇ��aA���j�U�R��Wp� Zd����Y��q�bn�!��������ݬ�����(�!
<��-ý��m+j�HmN���s���Z�P�68`�or��;n�@��[ږ�
>�������$=�����on#�_����n����C����u�믉_�i4�i�27�El5��ߤ�I ��`O�Ó�ҭ!�ܼxB%1�Ɠ�6L��$mYA�(_X�z��,��ڮfgK�q��|�"���Ź������^Y�SQgر�&����?�4`�U�GO3���`��syIg�CY��S@�u�!;�8�y2�S:L�o����~"P,���pֶv�9��b份�mF�w$	~���-/QdC{�wq�-��͌U6�f��
&x�:�q�P�SM� N����۠����ե�,I?䕰��73�<�T��
FW�#觿
���'�	"�r-���m�����jT9ХⳚ��H�6f���H����BV�?���*)f�����<�-�}��[����U��S����ea:����������)�����{��2h��*�X>\ck`����\r�L!�L`�����a)�����!R}#�2'�!��k��%��d�)���`r3ì�fL� Y~	Z��k<︹���a��b. @;{=Ȱ#�N�Z�ɿ�^T���+.��H��*	\�?`Rg�kj>�������ҹ=:ggj�Zvɇ3��V-��m~dD�R�\�=#8�b���B�N�B:�����A�-3�����+���p�1��n�':Au���AI5/�e�3�hۈ	�g��)M��Ơ�5}�/φhc��msnݍ�\���۳��h��5��]mf�b�F�z�7�,me�2l�/��ߗ�18��N���hu/��rcu`2v�e]3H�wS��-�|Y�a�%�(�I�n!pZƚ�Wl��������+#ª��V`��![0���OՕ��fqs���Ē��&���VB�?�D{)F��eޑ0��ۯ�3���YSؖ�Da�̽�N� S�"+�02�P�[U�dP��مD��h��Cv�+����h�1F�O� ��N���@C�8��$@��B�S��76���Bb�nd(�'�!�C�p~�K���/I�n�����3Aޒ@)m�.z:-5��o��Ď双�@����@|=4�x��ݞQ��g�βh�)$ƦŘ�3B�����\���&�����%��F���҄�����g�̙��8��ÿ�1�P�4�Jq��_>�M�R��QGl;]V7��qc~c���FdjY����� TT���足ɓ�U��]+$�}��_���&��!J��dL��GdL��i\X.8T� u6=m+�@�gQ���������%�w}� �:��{���եK,"��A�ƒ���V��3F��+�%�����Dv9��:@߷
�t�E�B�I�n/��:�T�N���R@67�����z�}�����!:ړױ����U�i��F����48	3y��(���6�3��.	6����& c�V�+*{tr�N�v(���,ó҆����l�\�E	��8���s�'`�p�������H���ј��g�a�`�������o@�J��ͧX���Lv�޻n#JK��g琒~�d�$|�������K߃��*%�Q�F8��G!�P�r�Mwv~�I^[N��9��j�jD٢PV� 	�B�9���p�٢�W���ֲJ�p�x�\�-{#_1 �s{|�"Y����ƕ��������%��R�ٺ���|z�s�/,��D�{�/Ӆ�Mb��m�Y��A��6����3iaF�Uk=�I��Ŵ��RT��)o'��v^��?2�'+��'�:*���]s�"���l"K̕,��d��&�j��a0��Eڹ�������
�g���:V�.#�'���³�I�I0�C�]��D���������!�N����p#�{�q�$@�A0���Iv���o���)S5����͓s5p�����!�j�q��(�'�<K�ډ)=�C�<]Z�L�W g�ڊ)<]MW�As%	v��������3�$��]�Z����Q&h�t�0�K�����GD4�"-D��GZ�K��2#�	���M�!XCn�/��[@�����5yO�^m2��M��%w�6