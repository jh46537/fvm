��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��_)��%%�.��D�ֹʮ��������7@��=�y���fA-krT������&)���N)������&���8Ol.4��^�t�9��Ai�����q>��*�sv�_٪����qT������\��=�"�R2
�D��Y�$�c���]�c}��Ă",=�Dm�@ B�Ňm� �o�2����c��o9 c�)B�wy��~&�N"x��#�wE�>�J��$������% �YdT^�#���Ϫ	� � cY���A���Ѐ�w:� ��fg&�7���HE�(��L������7agzI�x�ZU��qo3���z�FĽ��%fy�'g�3�Nuq����R7l�}-P��xv���+n� #D�d��b�p�c%�������C��9^-G�w%��-e9I�G�g���|�9ғ�H_�<	�Q&����C�y�z��2�����(��j���տ��oQ�S����Bm�>�m�"���5{��� �U�^�QϮ��'֟��
g����D-AR�Ə�d8�z<z�X`��a�����8�L��e����=�þ��׍��_� ���8x/�(-!d��;3;1��r���}2/Yx1��4�{v�(��&����Kl���a�� �AV\�� 4�x�4�DT��sj'h/��]��Xc�M��
�l/N��O�wr�d3��)��p��5�CCk4�˵�и�惭�m�tԋ��M���o�JWJ�~R�H�k���`�b�(�o���u&z���]���Ȫ`�Y*+]A�������>�M�U>vD��z�X��!�4�e[
p_�&����&�[I&�z���5���ݪ"�k�!�Gw���P��2�=��Q+�4�ނ�eH,��?���8�#0��?R��꣚t�И��8����#3�ZU8�s����\���HL�F��X���A�E��g<S���SsΨ��L<���٤��/~��
��OJ&XA�i�j���d�b��f�`��=bE��c��� �z%���+��|Q�T��k_e�ǻ��c�&S`$� ȓpǧT�PN�	+��&;��Z<)p	Uu��0�c��Wc��,������ucf)k���_ue���u��3D��n՘(nؤ�Ww�*:���l�c������/��(��5t�;"�<�������4�����e��WR��0�cB6(>�f�0O9qf��D�:*E4��E��;�w�*H���+�5�-�C��a����lɽ����b��wc�����7�c;�Y�;�/²�M�$%���*(1�mm�7���n*N��
&�/Wj�����?���+�RS~�����u�z�W�:�U�S�HA�r����[3�n [�t��I�q���e�IW����l��Kz�xD1�sPV"�"rҏ}d#��S�2a��	E�3;zݘ�5��2@`l�][�0�:~	:wtX�b+�T)�"�6�ԇ�}���+q���T�\��~`!_!4�/�`R�*Z5�0}#%�R��hlnxH�E4�q��0��_>ot�[":);��p���9�����S��Z�&W�:j��aa��$ß��*�$oR��+޵w����)�:%4F�v�yUu���	�OJ�{cu�r�5�y�_���G���/�MS���;)��og'�M�X�q�w+�(>!�
�3���q~����@���� zύ4�������H�\�j�_�r^&/a�':��s`����e�^* n.��^U}eĸr俹~2<=������lH8x3���+2jĽ�@cŃ�D��g�e@F� N����`�N��-��.i\�goy�v�KZ���V��b����W�(|�/R� �Cn^@�oF{+�Ҷ{�tG�7��cqл�x�����)��eY$����=:�y�9���8�s�{x�=;Vi����������AI�ȇ���_�iuc��ǃ=R+�H�J�ITs O�4)j&q¿Ch�Ǭ����_�&��SZ��~�������I׼2��hA�HS+�T�� +�;Qm��i0[u3do�Մ�(��*��P��<9~�/��zLX���(�p�S�Q)��*�\uG���Z��%'�\���{�~`��a o��a�'fO�~�����=�[��2e�@��!�@ ���*~o�k�0x�G���Wov�:��
������n�w�|�Q����7�&/9M���Ih[:�q�l�f5̗�:]�BG6�#������z���{$!�W�\�B�T�
7������@�;�̠��\�E�a�< ���0��1�:ڀ��~D���D�C  �F�A��ާ��33��o����1,��* e����C�K\�],��_�MW�^�6�7�[�A,��V��%1��@�F4�'���9mkA�CT���������H^-��cC@�o(�W�C�;��=�;����H��I�M]��E9�`�Q�VqZӼ��9�PMl�E�k�DI�����k@�ӳ�q<���z�&hyx�\`��rb��\6��=Aj������J�~y}*y����y�
�~�T��ͮ��*D;�\��eY��T(Y&hA46�
�3��Xk;���Wv:�A�pf�X���6}�E6�r�t��h�C��i��(�Q�.��p��o��1����%�����`������eRS{W��]Zr�Ff$$�b���KUgE��W�N����	7��D�r6MDȉ����2��6���k"ʮbQ�nI"Ӝe�uS=�0�w��#�$�Hcy",���t1��<��;��?m�c�,�P���4��8�]�����Rbd�������)�L�Α� p\;g��ŗ#�G�%�����x�]*���;i̴�{��M~oS\|��,��b�`_%���Te\����O�	�'��s��9�m;�Ǒq�C7�B��A.}cg��Vu@o*�~ڒ!�5���A �vb�mDT	{>����'+)\�|����������Ï��2`٦�aF�T���'#CO?�g�(���aR�2ǭ>Ω�{����_���yd��|�l��21 ����_���=��5��	h}< X�T�=�׍�8M���	�-?T�|h��!��`��"���s#pn�'�>툗%WF�+ր%6���.Ji�4x�VЖ�!Ŀ��Î��?.�(��cM�f6�=��\��cxc�lF�(F�h��ݑ�[���"[9=�w+9��dR���{*�GG�w\� ,wc���'�Bj4 ����i�5 ��uO��N�r��ؚ��΄Li{�b�u���4)^^x`�<�
�k'�d�qs�{���ojo2m�ag�`�@2�oMgz��LF߶��>����(H� g���i9HxLO~�n8�@߻ �����f�^nι�w��]zܭk׸Y?���gJzl8���L�2
n�����eC���~o��f�S������z��'��AĪI�
b�Ǳ����!3e�d|�e=g�����[h�Z���X��:.Q�b�<�l�y3���T�B�Q����tҖJY����h�#�>�3�O�$�r_��fz��!3����hA?�ežrvZ�(ů�2w ������e<>&}w,��ܲ|\�*lЊ��H��=��+vM�7+T{��b�?Y�ώ��W12F�����_�_��yZ���ד0G��1����)�Yj��K��-ގ�i�9�O�{?����L4�\��,=����j��͞�C��������**1>�^���
X��M��0~�V�������)偑�E=_c0��M�9�zgW��TR�|k���1;԰pxg@.ZN������"��Ah�+��0�Z�"v�<巂��x��Q���)5h8���|�-��={����hլd ��UxW]���;;�~���PMnoJ5���b0os�o��)��HS���[��~1�AY���\���(�˷	�=R�K�_Ӝ��`���8V2|��vñkq3�#_�t���^�*9����uL�tqjE�3��+�eb�5��E�l�.[<ش�L_�J�|>)���o��J��G`zxQ��5˾F�HR�%�_���:ru�$��F"�}6��A�����l�HU��JΩ��M�U�^� �}'��r����' �2���S笸9X���^m�ֲ7���	��>�5�P��ַ�B�Ύ���(�G&�~��j&�n�͟v�9���%�������~�ߥ+p�N����j8ɤ�O9Kn�KD2��Bkƈ{�86��O�(Ҿ��]�v��!%$7�z�Kv�ͦy A�y	�j����wǩ'n�h���,(B*vE�4��k�� �zh��,j��_��;�-�ww����rIv��0��Gj��UzP�3*�Ț��w��O����\#�g��8q�׍��կ�Y�S�W��.f��PVw�GO�WB��[�`��U˧L�������l�>����="\ʁ�|
_�id���&��d���D�eO�!��2e�(QnBak���f��c*wS����8�j�.A�w�#/�)���Q��r�/�uV<�h9���;���_>�
�}����_���fB��򅙳�-|�~7��h~�����a9[ֿ1�s�}��Ҁ�"����a]|^	s87^K�9`.�?ڃ�N��+#V��k�v!#8�E�k�3�4X]��1����	�%~�XΌY�B?�)��W����#(���N�Y�/-�(�r���'v�?�«���4
�Hl2?٠N���O�W��(�M������2����G�ޖ����7�^�������-��n�ƫgC���>�f.B�w�r�4TC:���\�EB��Te�{S�5�XEt�w���;�������Βz�kx7hx�j�+6��Գ��X)�=�+��G���y�ſ�P��?�`�����i���É�Z�� �R�+Q_���Y˯��oE��+�Q��E=��Gkȯ�q�W�`La�|�6�or�&|Z�N�$m���]k�����Ӕ�R��b�h�-i+�ťb'v"�;H��Mh��uZa�E���u������`:��$lh�x8VX�F[��	Dv�h���f��;��{\9�c�_ٟ����F�оn`dw��i�}��-�[L!�͂ژ�B&SS����!5��gY����i��o�gt����L�J��L��p��n�����t-:�R��=�<���Dŏ/6��l��[x;u�/R}�:;o���9�������LuCX�i��I%��F��3XP�(ߓ���h�S�4��\:=�b�Ѱ;Ij����1(9��A��p9SL���C�[8Ns�d0˞F ���s�D��C��-Υ�c;5�T�_��v����A 
!�N�_%ZL���m�C��3��V���/ũ�M`a]%2ALm���f��}���Rv@�G^��}��`��(��U]�(�p��8N�S�D���O@���
0E�������W�����֬͌�b�(B_A�ޭF;�X������TxX�'�Z��kUXL�S^c��#�����|A�SǎS�E�O5)"�&Hk;�ǩ�""u��+wc�(v�D�{gX�:"�S�v��c<��n�Dj����|�e�I���{�Z�pε3np�J��?����\V�(��*�i~kĩ�&�oV�`����ck�NQQk�D�������|���mӥ���u�M0k*6�Ǭb'��Z�����i���@�4=ǉG$�X;�c�WV:GR�4_F�G�i2�C�!�t�I�<E)���^��r^������K#(A����d�Q��A���I6I�� �Ha���
��"�2{y�\�#��}�� �o^為	 ��4zm i!���Iіƞo�2$ͅD��[��1]V��zLGܤc�Q���4Q4y�R�
lg�O��֐��������S4�WM��`m�5O�}l�׊�!��I:%�R� w�����	��r�qa�x����m��#l�׍�����8Q{K_��t]�nC�ف�]���	��O����V��������+7c���<&R��:k�-�����J��l�W��ߘ�WoL�s5�8�C��/g�l��oJlt���x?�\˟:�[ֿ3�A�H�EnY��k�9_�5iƷϏ��3
��������D�9�������P�mW�ndݗ��r}�t���\���L��{dp�I��8��U�Id闎e�x��F��.�ʦ�������:m�%���_�f�vIz�#�Q�r�px�QJ�	��!�����D��������*]83yz��Κ�aWr�W��]hv'�#���o|�Y��ɺ(�(�bG��[}eC���T$����|�Olh�W��蹡%["FV���Ҙ�V��HW��mq��ut[�y̨,�6�� k8\������>���9(�vkH^|�~�:zf�U鷧vP[-��e+�C����x?,�b��6|�!�)�����mp����8�` �Zc�6��p=���t❪ԫ9�SrR��wF�\gt�M0M���D n��n���U]�w͢0�z ��)��h�+�!�'wk����&����җ�Mr�G��4% ����Gii.�Y�D^�}7�*��zXq"v�S\p򁢏���,,��/�[zJ��u�k�J��l���}s�.��|?y��]�Y���X�bP�h?�7��>�R܁��Z��) ���$wm�'W�K81�b�R�bg	�!st=�3����D��<��#��ZTEn�0Im{[-�&y��v����8�Aꕾ�نW%�$U�@\xX�;��ŭ��؏�k�R(�-A��m]��sv���D���MI�XO��WcA"k�~Y'��%��1؇��d6Z��5k2^8w���ʎ��,��g�.�Ui�>q�R�.3L�?H�����{�$�o�C�r��;����#c���"Q �-�L�Xbn"!L�hZ��\������Wa6���e�nJ�#jo�R��m�I�gwp���U�����PD���Kյ�0^*$�*���]����yC�|�"���k�N�����w�]q���u��7��Y4��`Pݣ��nGvR�@���R�����P�xrϩM�h@}鯡|��1���A����b۔���T���;3鯧�����6�#{�p`��'
Z6����X��s��I� �e'�6�I!�a=�^�YF�[��t)�׹��V��E�/Ih9|2���!$,gi��ޅ�� �L�=u}����	l�{�f'߳7��[�R@��)����ĉ}�YY�s ���>��]�A=�lJ��Ȣ,ܶe��oU(2mД`���5��ުK�����j�y��s���B%�A�P���ʟ��T�����Ymf���}Q\k0�1Q�e�v��?[�a�p|���:�;�{MD��[�t@3�&ֈ�0GW�jZ��J�-*װ�'�j����r%�����Ҏ�m��I�ev<!�Ed�:��Ut�������/3)���{�W^���4Q������{��c�\WV������'"ӤV��i�I���uO�?�P������eC|t(@J���>�MQk߃�	��V_.�_
��wX<��C����-Aɭ��.�؛2�V���E�=�aM�v���ǟ��"�auJ銏�"St����j�$H��u�����{�/�"���~������m��5gMhy���HI�NۣU���pL�����&\T�
������l�jA�9O�ϳ�j>E����6���~��<�egG��`6[cl��8����LFl�*�̫טbD�ibՉ<�(_H_��r�_֟����-D�7��ì��mP�[�M/<w�S�ା�W~��B�O�#q��e(�(q��;w�,� K��3d�h�8� �d�]�N4&�RL�>��d����݉�;"S"��$X���=NI���v��͜��֮�&��s>J��w?���4� S�.]�.Oxo�OE>���~���^�^f@��l� ʨ���*Ș��v[�`�G���D��Cy��@��
|�U˃�Ŭ�A�rNt!�$״@S��L�Z���g�2��c��0 �9=��(�qzZNf�����_�lc~B���n�?\��%�ض3�x�"���pC4Sy{��	����դ�^��?����<f%��.�ǂ�ܝGF#ǎ���{�{�9E<�yZT.H��:E[�v���:��ƚ{ʵ�����h8���,�=M��ER���O2і�����ڜA���[��j�Pȿ�#�R/�
���t�k}*e����]�M���Td(�'W�ʛ�,�+?_��Q�р+��X��vY`��Yʍ˺���L�B���{Q ��I���cgCT����]=�&\���}��x����F�^J8��X_Io�.�A��I.��l]@8m�_\��s4�0u��O�_�֢ܲ͹�۪��[0������e��_vM2�DX�+=z�GX���3�w���$srP�x>�L���� 1qf�Qф�²���Y�	���c���I��i=��jAn��҉�o�?p�0fջ�nm0��l����d�q�n�*���s�l�Ѡ�Y+��CAD����,+�o�����s���liy��#p�5���LK�/�J��Cǡ�MYr�s�{������zqw@�8�D��˙xa�y\����M �Q����J��;���n1����$V�
q�I�<ؽ&�`N�C�>|�<����J9�7�+��c�N��K7��$��H�P����,�!>�Z\~0 ;Z�L;ڄm3��X���K��52���8�l_E��gO�E���g�+�4K�h�*��F><������u�
@o鲷���Yhl��w�<-�7cO�n��d����ا���l"�0��~�]��z���b��<|����+�á�gU����\a�єLB��G-�����F���{�ବ�U���S�s�G���gG�Mn�ԑ�*�6�k5��HGԬ5>� �o�� �^zƋ�+�gȹ�Fj�S�z�`�B����p)^ښ�<�6��@����h�0�;o�|�Z>�5l�A�H(z�<����+�ԧ3��[�Up�d������`+�q�}����S�"���2cA(�䕩���<@"�s+�,�f��f���A3�Fn�+Y��f'��vЄ]�Iy!&�su��ͣq͢���"t�WF;�y�Y�	�h�ueL��;Ф�2~r���o�����,Y��w��������b�%P�}�4�0�mE��jTqȈ+"o��4H'�����A�TwԺ\���d�XT�8R�I^,����Y����T!��Ã�Q�
��U��Q�����p�ںa������-Z�N&��z�l�
��(K���;"ӞJsm90�tdL���,?��#�	��E�
W zD�C�;\��m�*���n]�A}� �#�K����=tz �X����w~�<�8S>�u� Rq��ą�t�4!�p�9A>����+-Y��$l;�61��Gh�XP�$v@��
L��J�#���)<��D�b��ʩ�%�>y�C�P�4؈_��[���5��MXa���?(07���s�̪��^�:x���6�}����%���g`�K�('}�h4h6iB/��};���3��hS��_p����i���j��쎱��pQ����7ܒ����w|���X#�!�[V*�c����
�ӷ�͢��~՝3ĝ��v�D�e|�O7��c�P���Q5�׎dk���gR�p(p��J
��g��#�6c��؀�J[��py&��$C��b6���=S&��&Y&m2�����.��l�Ѩ�}s�yR����~�U��c��f��D��l�����t:���:��"�=2��Dh>��O�������(�D�L�0��^���d�(�����H�s �-s^���n[m�V�S8ۊ�&��¢��cE5X+�r��M	%Q��FB�REK��J~(_lh	݀3`�������*����)�i +�Ӫ��G��rx����Tva�e��Ɨs�8i+T�OE�y"�Cs���V#��B�y���-�v�g��Ρ�ڽ/ێ�^!�i5�1�f4�6.#SZt�?�e�����#��C]v�a[@�����QGT�Թ��*r���o:��j��	�[rdvrZ����3l|Y��g�7���%��<�m��ݾ�����I�M��n�O����	�
֔��_�%����~dz���!�u�T W�d�{���U`:p"�a<�GB:�ےm(��:|'����ӛ�V҇:�0��H��9�Б}䮸54��('�*�.pl�P�#��$J~
��X��@���� ¦nǹ�}�2��i��&`]�;�����n�d��e��=>�~6���u2���̊�̘s)�Ty��"I�)�?НU�E���j�Sek�l��Ҝ�׾��W�ӧ>x��	.��p��E�N_�1xH����b��ԳRX,���k��n,]h+����gF���3�sv;�^KO���]��Y�O�,qm��W��4y�7w;cF�f���g;�xҸ,�3+q1���߅�18v�$�B^4�|��{e��<Õ�.��V�&�<7�:�Ǔ�r���
�Z���xν$͔8�c>�Y��A
��4Mf���lx����nTR7�$�6m q�%t��#?��L��� �)�#�(V��1�Z��x4
ơ���/�3��7eˊD��w�hi[�Rq�}EhxӠ��=s	0D[Ҕɪ��#�z�N�4:v�kI���呏�ҏ����4A�2�|P�]T�lI�Lk�c��vV��)a݈�J�:M/l�p�K��çg�����
N����7L K�<PA�}��QT����v-��X�}�j1$vb�P���t�M�� 9B^��{6:���	�]i
�}���C�� �r{��85i���+�ig%�R!3���V��rJO�&�;��4)������1���:�Q
���Շ`2 &a�Ϡ5L/����֧jس�H
س<T�����`�2�Y�ZGp��?X�k"��Ϩ�&�_)^V�.�e�������s�:�.�-J�zt��:6�Ma� �\��	��1�Ps08zc���M�6�u���!(�zz72iG ����&��<��h%�X@��o���L?`-0	��7���V4�Ͳ��{@;>�����!��%�?��,(>��}v�;�������U�W�9:�R!d��wh�бnf�7[ ��ln:���&C;71&��iX�L:hF7k�#}��2[�[ہ�dg}I6L{�d�;3�@z�� YZ��ey<�C�͟�����.2�@z�8�t"�ts�%CR&��r������$����TY�"�X13t��F�����VS�Si�&/�-���qv�|((�(�w>�8W��u��ˈ0�K{�GA1[xEcȚ�5I�r#_Mnw�`a��,�xžUtܴ0�M�j��� ����^xs��z�gdo�#�l�\�O��2���yIM��pOz>�
\Rz)RF���<�cu��wl �(�W)R���?(!�c��o�o����`0�a�Ӹ�cD"��i/QŌ@(��^�?�d�䩩�������AA�8z�3"oe� %	��ء��w�;�Q8�>"?�i��Ψ#��ƻ/��b .�������NxS�^��#q��� �+jԇ�Q;��f�� y�,}��'�r��:5⳦���{%b�\�h��]]G�pw�$�'��T��"�U�8�,l�}i����ы��A��p�`���WaJw�����7x�i	���G�4����\�0�����r��	VF$=��	9������#ۤ���f�2��&�8.����M-�F� �j%@�K)��p)�z.g�L��w�X�i|4���Us���������^|NG�d����ﮞޑ�9/�����::U-�XC�^�\�Dޣq�]��4���$�*2���P��Zb�x�B�o����gmS8 �b�o��:����T�&T퍽�������%�ѻ��F\��������`W�Z�fɈ�Ѫsݻ�Y��w1�u]`Q�����i�Z�4�>¢B㔓�����%ӗ���1y,��fY��=V�kX����(rT��$6�a�z<S��!�m>��kd�=ހ��.�2�� ٩	x��=ot�Y�U���"� �M%�����hFƕ�Bb�ʁ��8�V]AY{ܜW���@���[e`��ܹ��B,�)Ou��'�1��P��ԅ���wT�	>y��L@+^���Zd�J,P��X'����D� 뙵��^������b�u�ծ���0ڪ���T��<��U�6y}C��?v+M�"��w���,�vW���P�)�z�����o���U��7[z6p�&Aj��R�x#)�(]W���]%�_E�'�]P�\+�u�nK�e�1�,�ӡ&3������M�r���ͫ�����;�bk=jR1������]�Ml;~d��-��-��TII�Ӗ~�J����ځ
�\d�P|��D������H|p���+����M%��#��]œLnr,��CʉD��Α�3�9twJ�P�~�����Q�g[8���0�U����9�\ʆ��ۤw2�3�u;@̠K�w!��w�VR=�B��Z&1�qѮ������..p���4d�3���>ä�k�sp��RJNY�W,���ѫ�@{��:�$��I��B]#�̜�˘��4o��e}����FL�9#yzr�Uo�+ޭ��c�� ��T��γ\�j]�ICp�_6��6���~F²�Ӷa��χ1����>L��sF�IH��G�o�^��YO�xh���4u�Z�ֆA^)�D��PZw&��s{+0	��rLaS,�����L��� ��e��K�8�VM����_�ͥ��<�����L�R؍�S[��B�ؾ?�0�ѱ�+ΪR�5���>��_��7����V;ao��8��2�k���ɯSo�N��c@i�m2�kE� �t���c�`�,�/׍?�����LT8����?V'���W;K�jT8�I������n�/`�/�Oʭ%�@�ژ �%����1���LX��Q������0M�ѽY�N�a�P𑊇�C"�(A����U��_I�\
��s=�������{���B�=`۪؇�k�d��RZ�6�b���
2�N�Wc��WЃ�I�i��nS'rH%���w��%�t�����pk0�"�#�N�Hc\���7�g�~�����魝}��&w�b�UV��+���=l�c�;c�ą�B��~��Da�^~�_�y�m	l��p�f���n��BS�\��-�l�>��cE�aѓ��8hz�ݞ���i��	�,���oSG��NTA�z<{��"U��"��8~�k��j���*���b��-.���w��P�I7w:7Z4e����P+;�X;��2����F���6�D��=�Ch�%�}�'gj1(�\���+~�~~�m�P��FR���|+pt���6w.z���cr�����4Y�-�%��dgj��}�a��"҇&"��`4�{�����m�j�%�rpLo���A^�+���音�K���TgY�U�ň�X�I{�s^0���M�Ϣ�X�TS6@�����in�V�y�<,O�$LՅb>~�<�x7�ʫ��ӯ�,PO��j���>�S���Ʃ[ 1(��	����F%0`΋-R��3��1�m$�Z�yi�X��s�����R9�a�"'{��W��j�}�,��"X��0�!`h�mݵ0�啞w�o���)i�09+p;��i����\V�S�8��Z�&(�\gN.9KI?�;ڔ�.VQ�<���?M"KH6Wp��m#�����$�Y�h���^�O��^�	J�W�����_Q����&}���d�pj�pfQpE�C쪉<�Ye�È��.�e��pU��OwU��x���YT����!�s���f&W�P.�ᑦZ�bX�,Mɬ�Rn\vo��?x,o��Ţ	����.�7v[�*�������0��Y9y;���m��}�����&cl��pp4��Hg��4	�W�>LG[������p��:���n���q[f�JV5�Z��8 G���OcS\��֜�oU�����'e��]�Q�$8RB���&g�,-L�ǜb�R-f3����\�����TA끣����QW����⑾�&���=dq�s��բ���^#4w�Ą�ţ�������Lgo�8��x�������p�a*4���~��Z�`N<T=�3�$ۜ�� 󬼠��{�6��4���U��IJr\#�����Boz� �0�HpݾL�
K���x4@O'�Y�d�ť�W��lǎ�Gy�zF�ꏼ!��,�,^c�� ��8�Ӳx�qފH���N��j��rY'C��|d�n�������6`�i�v����b�o��ܾ����Î���w�n�x��M���g=��v������UV�N�!�D�aj
�<h|L��q/J���5~K���$ר]�C��i7���� �(��^�6a��z�n;�
ӊd��oD����\�ܷ%��u���IߠG')�ʸ-�r�k`L��`����lJ�����0sq�D
dǵpx=�J� �3o��2@]�^G^�3[���Q�w$D'��;�����<wv���N����M�t_���]e����܁��� R��P���Aw�Ql��իo#�؆h(�*s��!9�|ևA��.3� U����b��rc�tF�H��f�]U�����if��`��2�!C�����hFb���@�6�eza�O�6��z�RA��'��xUg��;\�xmy��\����ް 	c��hsm6ɼ��sɰ1��ݢr��f� ڜK�T�X5�*�djg���)y�
PR]R���k��������Ӹ�/gn,��@��h�	�@tC���-Z�œ��V��Mlf�Y�L0�q�K����x�5��fB���	�w�r�T�9aa��F��w�:o��| ��b&��E&����� @A]{P�ག���Wۥ��j�(� �,�]as���h1�p![=� ,��F$������pk̪8���� �F	��/|��4��5����}��ތ/)���gC�d=���k�U�����޻Z	��pAn�k"�U���+�6��_|�s��1��������L�D�����u���
�SI1oS
|�S�/��ߩ�A��t��|~�ʘ��}s{���{����Zk"�Z>a'��a�% Jl�����6C�v����R�ڟ����Ɲ��[�3Jx�/�Ǻ�������9kқ9��j�!��pZ{�����,�W6�d�7s���??�q^^�=�B�/ h�f'�4=�h
``du�]�y���jh�z̑��`2}8�`IXf�U,�ɫ�)����!�;	����P�h3�R��2�e� X��5_&��3�����h:T�.3���5�@��$%0B9����򎯲C�W��&�k
ik����F+;OӇӚ�0��?>�>kx���sr7���{�5c.�Z�T>��j\m�-�:
̯�a%��Mh3���Au"���r	����W)�]nA9�\1g�4R�� w��� Rܜ������-D��h�:�1t���X��˛���Kf	����Rc
?��WF�2H7��Q�뜊��bK6~�=14+ѽ���H�V0{6�x��:��f^|�y�q�<2�5�FɜO�﷕(☓�������r dg��{�*b��y*'��� ���c���˧���b�����1�q�S��X��M�l����v�*�-���B1�7l�I���^�[K�化A<��m܏�_c>��<A�b��:hY�kUpBSA��N<���'G!d�k����K�g�Nx}��GɁ�V�{�C�Ԁ�\'\�9�2�lا�������e�[��MIE��|�)����,���!U��Wo���?��].���$%�������Ȝ������m$v�r1�������l�5=�C��J�`/|�)�	Ѩ�����bH9�ey%����8��7����������7&@�e����.�q'��;��ۜ�#���`�򋀦e6�:Ƨ�9P�1���@nC��-�z���D�=�t�:�j��M:�ǒ�8kFE��R�g�u��X`��L}	NG�m<:M���N�c$��4���V�����������wT���f �b�S��?d�6�+7�-kj�R��=��}t�@�Ra��I�FB�З�/���˵�<zx��-;y�H�?{N�WM�x��l'Ǹ�k�`.!D T�����5����[��B�a8���	�y���Ur=.�4!�Ζ�w�jd66$>�R�	�F1 �]I{��`C��а��l6>�D�q�nqW�7�DW 4*���y\�Ұ\ �{�p������xo2���p����{R��h���0B�so ^�V���ͻU��O�qk<[.�@���	7���`�eB����n?����RG!Z�T��ol�I�W#"��Q��~� 1�����/X#�4O�Z+t,+)3.�3v�C�����q5~�� b�i�ә�_+�+�_�y�N��þ�����K��$W�i�B*�{��	.�]J�F6x9[��Yf�c�V7i]#��ͽ��f,������m�����k����Mq�*�3,t`�3���J%M��T��H���æ�׵��
�Y`;�X�D���b��
�@�[�*��$�M}2ϗ�I.
u�A�Е8F&�j��ak����<()����, b)��׆�+���ͮ��=�7+�ֺ��A!�`�6Ș�y�d�3��ik�@`��mQ#��H�='04�k�������I��fjr �Cks�c|�|��Ck��SW���~?ġ�@���|�o��:v���[Y�S���	����{*4�X����>�-?�B�#Tg�F�(V�Q�[���hNO��	�kxN�崵�q<c_��}�֌�˝o��p���S�[~�f[ƧD;�N�M��>���&>yWԶ�$�њQQ^sMeg�Swv�GT'����>��H���ss�1Q�t�<�e�?v�}�և�O;V��٣�@1"���`}ݗ��8(�]��Njx����EN2�R���h�� A<�S~n�5����f]�R���͞�L�����da���+���O>0O]uDA� }My�|�2?��a����&l���]K�[Y��/DW`�7<�@-M�dǷ�B��&]�Ap/MO����>?:���m��I�&�O�O/��d��2��-� X��Q8�D�{��&A�1��9�?K�%�fKB�����R���,�T�S`A:���[�˔�P�!����MCm�C���Q�O:�3M�g	/Kwk줵|p�~/��D�/��n;|�j<F�d}h�Qш��u������q"��26-��&*_UZ�*�
�~:�Db�^��ʤiho*���T�D�1?u3F4ڮ(��GlZ��S�B����nZ��A�C a��;�'��Y�w�sP�fV�aX �;w�<�����E�V�i�#��}V ��_x�d���i��r��A���V�<�N<-���I��ͥp<�v���������a�@���kx-R(�|��C~�}F���}�]��p�I��c�[N�S ��X�D!k{�s��x�v"�����_��p��K����(u�m<R�y�4#U"���C ]�~f8�p��C��Si�^�a<c�K#�����j�D;��snd~ljv��n��E��ߒ��:�me�ng8�4�fə�w�l.�9��$��Q��D'�܆��.�J-�Z���Y��l����E��l�����Dd��!�-k�u�WѫvjBg�D�0���#1u�HXg���+�$ޚK����`�ǔ��"�;_̀O��j rz��R�q�V)=�4wßc�=����O8)%O�ADe�׿���,_�H���^1�z���:�,��z�>ۄ�d}	�����n̽����)1b����"�i!�ݜ�ޜ�/�4�*�W���L�yZ ��dX�,"����󱁂=���]¨�t�l�3(�b�q�c������qB/0,.�M�[�:���9��ԧK��B�0��zdc���S�?$�w�V��$jq(��$$���ڜN�˘W�[3&���R���]��%��2sC%����+04�_�g�XT���������%���)ӄ�������Y�k4���S<>M��8;���d?�1/��}���Q�U-�nU�����r�b���mH6�S���r��X��rݭ,�
��$��E*�j�װ�8]�gp�	��
(J�m h\Oqvm��҃s��W��9h�M�$�����<�Yw�.���&jYyE]ͱ��@I�����;�1}v4v)W[U��,��x(��G�T���Ǿ��&��9ɸ��2 �j�%����^��l*���i���x�!����6��r �z@�+��@�H�����%TrM��AE޵�0�i�L<�ݒW�����|�V�D�h;���R��l�^Y(�(�$_O$�����������P�qx���b�{+Î�]`��K>�B�~��܅��-J��i�{f���v�Y1IԘ��� �Z$m��Z���P���+m<h�f��V�%�f���:�P�U�x<�Ej�d�J�%� f0��2��I� �V�g��� ��g����3�H�oc"���º4�%1 ���T]�T�T:��3��>
8�:�6t>�o�֖�)2R�l^|L-���p��X@�҉y�ޡf��S(���z��߰�)7�D�[�-;��@��w9ȑ_u(-�o=�.�#�~2:Dɺ��؏Uh����Hm��p<Xb(/��ac�r�f�q�2�8��3�F�b��O�]u�'q��	��R���.� ��·��8`��#��sO��\Ȣ;���'L<�@�_��X�r-˂�]ҩw=Y���qRb�P��[ ^ɮ���I��If�9B��|�=�S��[��W:E+ȯV�o���f�}>0��������H,z�'�V��PrG������s8�@�U7r�x���6b���$RI@��<c�*q=�x����nO�Oǲc@]G$EQY����x��!�+E�b0���Ț��@�����+K������_���GNZ"Z��`��m���nD�����%z�~�.i�E��Íoʓ�~c
u�Ч����B��!��T	G�>���)�z��I��Û�[S-����a�=��keI�5��ൔR�U)���q�'���ȫit�O���b��h�-R���W5e�^��F+'@ �SA��e_�QK�:���$`��Qtn�u��7|�~��S��$?�4��\�F�yN�L������ߡKӹ�1���g̯���p`��2 �Wv&K[��Ju��.}���da�K}hH���op�}E1��Y<��v�7��g�Ͳ�x;R��Y�]Y�a�=Yʾl���`�d������"�d~���n��n�^�&s_A��5&�;{cDZ
�7w~�ܰ��mynwH
���
�t@�#B^�r�n�e�����a(S�97(u����U�g�Ho�r�g�����
���¼�E�%L�����X�p?�z��5+,�lA�tu�lL����辧9�z�t�<��ȤE��P^H���.���`�Bn	�Cq���bp񄠣��qG`-�=�
����*�f*�"<7��Y6��\ף]� [�SF,�ah��#g�j�4�������S6��q��O�j*ސѺ�vڄ��+;�����"Q�{z��:X��̛�{WgN����/T�G4�G���,>t����B�=[7�?�3���A�D���@����E�;�ұ+6�j�~?	�O7��a$�vig��B���(�>W�����	L�����w�����3T�r6��k�ل��?�$�G,�ʍu%0ګjd���5�>'��]�_�B��r�r�d�&��pGș�Ώ-��0�ݷ����Зڥ�	�S��5��5�D�&|��ؕ�D�~ߺ�%^F�/Ő�^u�\��?�p���c�l	��=�@�n��� 5����ȯN��.䄯!P�K�a�1��F�FڳqF��=K�Z��� �B�����Yi��諫�@��8���ͺ�8GyX�m��l@X���c��VR��]�/�&�nu��)�iH�x�%�g��p�`�z�k璏�ܿ��(	���6s����,�bȃ�s�w���Z����'ד�z����d�vv��Փ��aѭs�[�8�`3��I�"���kua��Lu��sWz�S�]�{J����,tH<n��@3�}�:��q���鿰2yn�03�ʑa�P�jWC���:������昅_e-F� ������s��o��c�={L5�Â���Z���H!�	�D;%j�C�I���Q�v�诚-�3+�A��X�r�Q]��K)!x�1Wx+j0����g���-����2��M�C�"v���5Ga%�C�gf)�4�|�҅'l�^<?�E���;��_�Mr	 eUg�_�}t���M�<,JB�r�`D�w�2�4�2.��8n?x+��z�P+���Oe�H�i][���:�$�� R0��7��n�k4A38&������Y�I4;���t��Z�G'i�w����F�Yva�&WO}��6]V~܁/� �k5τ�r�sZ���W�b@"_PDt$���"׼���׈zaz$;(�]'U��K�]�$`(
%�a�9Ył��.!y�f�ՠ��=�:�?1��Z���)��+�i��dbS;�52t��utXl������D�D޿V� *����p���%/\�ŋE���jA����{�s�$��8�s��`70����$	lЏ\���+�����g���"����~q=RZ����J�#H��VGc��]�0`� R��i�L���H��l*�B(�0�k~h����K� ���=w[c�2�_�H�Z�	�`13��H���K��꣝���hT�˨*|��JY�/_�Z��riMu�l3ib�"N�1�q]���'�	�w�ٕ�w�ڎ��bXk��҆�\�M얚j<�4���I�2j�B�ܹFZ0�߀�*�^-�]Þ,���7Z=�I�|�������/�E̳�&7��U��b�nx��]��D%F��(4�@���d�3U������ܫ}�H������I6���d���\���6L��(����΁3�`=�=/�~:�4z�$�Ǯ������{�ʶ �H��%IX�K�/�G�8�B��.B�QB��*f�`�( gQ���A�(Æ�	ˍ� ��I����6���3b�s
,˙VN���tbr�:��h#����ѽG��#4ԎN���{�����{�,�,��xaj%p���x���^���(ɨ�E0�ؠ oi*�<��ڱ�� SM�V��u�P����Hn�AR�i�^?$�QP���>�����m�� �ڑ�վ�����^�f?-w#��t�����4Ѣj�[�;N����#�*��HW]V*�pnD�=-q�ӫ2 L�ª ��E�7e}B	�Z��b\�,эF�ݓ�M��w���a,;�6#X����o5�/�N��R�rY��H9�_R�����Ȇ���A6�~a��H\�ʈ�C�3��E͏VQ@S���Z�/lV�Ш����r^%����9�5�5�(�ix���^�go��#r�Ζ(���MfGř��ˁ�}�xbV�#$0&��z9%��H��t���®���i��L��:L,T� ��3��tK��<�~#��Ñ퓅82 ��}��r��t�3�W(o,��#�-|���M�+kI[sOt�%���c�ڂa9�
q�ub�Yp���Y1O�F��o����eBߺ�%�\�����~��5�?��법/����S/���:|��-+-4������sDd��}�.�҉�Q��ڻoܳ`ݸ����w�+���h����/w#�(�R�s���n�lHX�-�a۴��h����y���4=����%�T�0�N}����hvCl���7� ��^׳�G�n���t)C��XX�����Hr�BV�砸�;ʙvf�ݹ�L!r�`�(�c[U��]A�x��K���f��?��,�l_�l�0��h&X�,� ffH��M�B9N*{g�x[��iq�G8ki0պ����q{��g�9Dm��9e]����H�>��#���t܌�.�z��SԢ��=tE!2����M��D��f�=�5�.�tao��5T9�-�R�U���<�*��ۨ^u��}A[�0�4e�Z�ݚQT���ʄ��^P�`� 1�˨;���H�5���sJ̏��]{ۚ�:�,�R��Fq
�|�_�i�BFs�������/��w�z�����aj�n�~UbM��m$u�P�����|�̈́/��zB�9��a�
F�D8�گ�e���2��u.@�$�*�N�B��
��݈(���x)N9�fYu �}��]\7wc�b0 r���H��fj���j�эU��g6w�y�T))'�0%��0)rA`��Hڽ��'��o�+i�=�ڟ�97��i�K�%��g����i���	�W��P�
`��}�w�Z�_����Sk�6�ؚ����o�������B�A�AH�q(���Ë{��`>ݢ���[2�ηv�F�-Pȷ�d$d�c}�!^�T2�K��8�>���m��ŗQW⭬Tl���:����Ͷ�4B5U��T!�j���T����Y��T6�sr�'�W�|V'��0���MZ�z�s��%�-D���}��G� cIx�g><ڥ9e���w�j��ޯ���"F&�s��7:���M�|�!��;fF,TjC̛Y�a����9ULZ+b�;�֍�ʣ_<Y��Ȭ�(�V�@˼�:��6�?)��wL����Ͳ��*�h�Fǒ��5�j�v�{��ŋ-| ���%�U��P���ǒ�"��ev��7�RO�Q%+b~�?`jU�N����~g^��y�滢y�o��߿��;���3��f�l��UI1�Y�7��6����H)�(u3F��zV�L�%�i�ǒߍ��y�$��ߙ%��J��◣5�,�\��>2B}�.H�>�~�@n�%���=�^y�m$"r���Q�΢o�c���`��v�����Մ)�0�A�C7
AcX��P�kh���6� TO��4D���l�E�zLB=�N�9x���W���P[��ώC���d�W�s*���N�����k�[���,D�Ũ�s
&PZ��#�`+|�/r��^s*Y�Dn�[ ���w������S�5dH�I$�8�د���:Z���MxĖ "�Y�&�?c,�V�?[ ������y�18���f��.��4��ݡ�/uNA� K��'� W��a��6������n
�J���9'�����BnC ����'�5�bPYp�V�}�&fʃ��/	����#v�k 5XJ~���������4�a�6���=�r�-tY��c
ƶ6��P�G�yᩙx����\�̗A['dPK���>e n���Q��L ��_�r�Q�>���&>�i~���'C6e�Ae^�Z��:��T'n~�<�DC�oX�q�o֪M�R�yF�?�[�ԯ�R��yA��$����!��bs��0�mZ�֫���y��؃C��EM�CW�UZ_uK�^�+&�h��Y2��9c0(?�ƜH���\ j��x�%#dj�o}xQ��$��ܷb�'9|���Z����9�$˂�+�@+c~9*�{|9��Iv�Ny�${SA˙��H��!�+Y�U_>dW*��Y@?7I�޸�%r��sg���Y_�W��� iC٭N	�AJ��86�mR6��O[n�����9���6S���r��=�)���C� �:.Ǆ�g���z_1����f��U��nR���[H�B@��+eA�ʭ��ө��iJ�i�4̇�h[ٰA� OK���f�[�N)��tv��P����L�������ɣ��C��JKi�o����[�Q�?��8�p���=��(&�G��Õa�]�3mI��Vȇ@�͟����mrZ2�O@)�k1�,�Ǒ�-�Afk���9`(��P�G��]vr��u0�l,�%3$ #f��\�j��D�!�|�>2ʕ���H�NJ�\j�]�\o��"�2
��q/�O��� �[]��(����i}��ID�����6ry�Zft(�����'b��OxL��X|�����O�H�t���.����3[�YIB	?|b�*���MtW�Q ��@��T2*x�?ؕ"�� I�#�P􁴕�Q�c}��Q2Nb�f!;�bչu!ڲ�����ݫ������Q��<ӵ��iL��ҫ��+
�
���.���I+!#<���\������-��ܛ�C7E�^+2h���-�H͢�k�:ߋ]����ց�H#l�_g���.Ӏ]�������1�"�|7x��d��9+db?p4(T]Ʋ�7C�"�3�8�h�{��U����
U�Ig�Wqz:!�>2Ip�$&3r��� /c�.T��S�1/�k
�[�|&���@-��SX?ȱW�EI������������O�-�*(������q�n�yҩ�b�WU���߯�t��#P�1�Kb׮�F��~o�P(K񘋃&�0Utc�!�<���#Zt��I���)U�b2���9�4SB��o�����Y^�k��00ȵ��O�5��Ee��e�!N����h����2�\�N�����ݍæXG�v�60`�
�t�����H���D5��F�Pg5�l©�N[q�f����?X��~pڶ�����tN�-���`�:�y�Eo_�zr�����ʰ����h��X�,�y�6iz]yFp�ڍ^{�/����9lz+�,^��1�^Jw����a�(Mr�!is�^8c�v9��Rw>Ҙ�FL>��e6��њ*��%A�����f_28�Uī?-�n]��{�m��[�� d<�c�#�VW(�Ms˒�;/WF9��}�Ν'�m�+AW�$�)>�2��L�ԱT;4NR ?S0���HU�.\X�Qp�n����bD��ͼ-lLVO����_�ư��i3n	�Ϛ���@�
�b	��ɍj�M�W*�`j#��]�����у�`C*�t`'���'���!dZ~�\7��� Љ��>�9�0T��~<]���C�]��p�~��\�
��3��zc��� ���w����a�g>�'�~�R�G'5�%�!>1/Gf������xi����$_+e����OL�����QW&z7��2jMR*@��╳A�/���W��׹>s��<@g�4���*�<�P��j��w������9��֒���#�KA(�q�}�0�,�4�F���#-lG �����o�c�ztQq�n}sV��35x�����-mj������]�A��2	��L03��w��U��@���2vjV���n�	����㤏�j��5� \��*�C�ם47<px��5�7.M�x�cf��n~�oZ��9BJ	�-G�i����P@��s�)Q��h/������a�E�'��,�J�o��:�(���:��ނ��4u�@�O���Sw=��70�4(��>0��P]�{ORv��֧��'fw�sY��G���ԋ����<ߍ3A��m^�~�T���-�Gcc2I!���jy?�����xX���� �(�a߉;��&��ۨ1��`��n�9X��V�t.d�'��t��D`����?���ܠ��^}��Ϧq�6̲k��~I��۽�� ��v����86�?T��K�=���)xT��q�)�)'JܪYN�P}}&�EmZ�ǆԘM2ұ43��,����ҍ�@�+�:�4�-W������I֚�EZn�0�G~M��د�����ne�&��\�b��Ħx�P�S�Q�'��ʧ��a -=4h�*������QR(\1�F^������_vfR?ԢI��{�5���L�w��
i�=!�u.�Rm12�fa
�`�,��l�qG�j_߿�����"ܣ�����7�k֝��F�k�q�l+�h�Ԩ.�v-I+*�ʣmz	�v.i#�f���a�ڸjX4N�+�1K�ATM<�����ȚmpE�2OY�.�ϯ)����ř���(5�}f������ #�N:C �����8�W��Ft�}� �C���O��`n<��p���7a�
˸�&�8�?�$_�z+�
��D��܀;�`�+��}����i������I?_�v�O��%}�{ow��µ�
*�*=���իU��!��`<�}����Q�x5�g��/� �m���8#r�a����rU_��DTFm�t��4CE�'@M�ڙoyT��e_�x�s��ֿ\z.�����#�s�gMk��f<_��＜\��~81���h����Si:O����օ}�>��¾��f�g�g�:O!����^O�E�Q{-\�!��K�X���S���}0C������s_I�>n��j̝��
�-����h����r�2�Zv�)W�w>�ݧIB�u����&���^�l���Α�8��1j�0mk8 ��6 �)>q�DH_*��� ̐��UI�	؏�|���II��7�#������!��N�<���c����s%ǉ�*���l�� u����@�vĲ�Q�b�ѩ�>�%����]ɨt:�O��/�~F>9��[�k��2J��ag�)�]�cn�����࿰�c3״\��Z��8�:d�<O��3饶��<u��<�{�����VJ1Y������Ϛޡ��T��Q�i�A{sA��ئ�"��eü/ڊ,4�qJ]�����@�f����ֶkB�B=�;��x��;ò����YM ��f>4�W���Y1�j�$S�� ��s*<��u���b�O��I'IQ��i�FC��Z��$z��i��h/v��̛����ó5�<,^���j܊��v���,u�ª�Ƥ��r��>��Y����u�&M��5(�MC	u�Vׯ?�α�d��2H&J�F1��>��[�폏�:R���Y���w�̎C��1��
i�ƅ~o�o�{�fs�9���(�a�3��Bx�-�"����"P�7E�����P���l���gK�ک���������L�E�P���aǴ��st�mB?K�Z�Q�9�;s��g�=^uC�IA���z䂳��qLt3f$�TM�D�"���y�s|;�[B�S��P�������@Cɰ��)�!t�������t.y��[��1�̿��)Et�b|�Q�Vje�_�\
_�^T?rK+1h��I����	?���0��F >��,�c�e�`�M�Q�FP- p4��'wVU������*V��;�_vI�&�*-xB>�Mk�H]�A�k,����~���q�����kE�JR�v�Cǒ|%<V�,�U$�8徺:jF�e���e#�� \����1������?�غ���i�L�qI	2r3�P;.��n��n�JT�Nm���Ha����4x����S���W
�������HS`ڧw,g�J���qf5��-��
�rV.�=L_"�8# ~,��;v��L\1�n�J �:bn��|G�R��#1Q@���;|���"��i�Y��Fs�Je�E�� ��|# �PkbX��%���R�?Ő�k�*@M��0 �.OJ8D2��ϕ��>o����YC�:q,b���=<�j�}~G��^ڣ'g�g�w�>5�A�h,���������X#!��}0J�˦�+}�v�1 �fQ���@�ym�.9������x7�[9�EoSr/�9�h�rz���Z`��#���@��S��t8i�M)��q��3�ߐ�'`���ߔ���#���ت!�T��7����:΅��G�c�$gø��?�cԂt1��gdB@�m[�e_�o��o���h���$���ٔ�6���.R�ϭ,�����a�>V�`�`a���h�[�Q?/������54�7E��+�kK�믪�1aIZ� �G��d�:�s��J�&����jnn#f@8gw�Z2[����Q���"�eUEěsNQe�lPL��pZQl9v	�S�tu:���� �c +���} m�d��V��۵�ؿ��\'��6�f߅]�,:�!t�/�0J��Icr��Ub"` ���-O�᭸��r�{덗]Ue�ʣR;p���̺����XU���g|&�K`P�a/&2�M>�
I_@��@������zY��O:9}�����Jǅ��
�p��W9��,�Fa��o�1���`��i��=&�%_\�)�&q&ƐP?�_rs��T-z���q~I��&*@�t�꼶\��+��^�3�/��G B�S`�1��:�7�����ę��~��1#�����f��
i��]Ճ���f6I�u�{��{����G?��@*eD�Y�'�\&�./{A��+�Z�yY�dm�ё���J�h/A�}˹�ˎe�;qU�o�'�5��L��D����20Yb2��ى�E ��#d^�;���힬����ɶK������/U�
U!����ǎ�{��B��-o_;��Tr�.�{t  *��͟�#�H�cH�l����9����'jϋ�s%���Бϐѽ��Rȭ�Ul7�6�0����$��$�9)@���%A^~�"G��7���V�|nHc���{��OP\���F*��q|v����w�_��s�oUo��t.��h,xcM��<�焋�i��-R�\÷>`d�����{(�e��3\�v��Âl|�й��F�GG�E��3�M߭�M�^t����!�a�}yoTwP4�Q.쾗�iȟ$]v)҇��ѯ,i�;*B�g>0�/D�> ml�kx���}!�B�gL#4aA�BoW�o�X~��W��Lʘ���[��W��X�5���L���q���>�'�/�(�fj2�)k8���ΡD�+�e��~)�0��y�H"�O�P��J�5?�G�q�m����n�sZ�|"���S��{aLS��ȵn��Kg]��͙~W�i�]|!�/���$�ܝ��<������`(oJn��q.焏bH$�	�(?-����A��~;M��t��I3�]'X���{��!s�v �)w�MW�^��ΐ!&���a�`^�N	}�KP������C�sc��,�`�)��b}a1�W���kt��=8����&�^���=R�6 ��K�3��<�2k�&7��	�WR�=��n��،5J���}}��7n��cP`.f�eD�HHu���1�$�6:�k��zK�M��:��sQƝbGj�D��ӻ�/�%��c�9��0l���׎�>�j���`{���A;�	�RQ�fJ�i��Mk��@�xӘ�p;�C�R6�"��f����H� �"p8��~,�S/�^��8҅9�ID�Kg�x���#���2��+����O�mEjtc�w��2x|\�F9m��@����tH�]���^�5���@a��YC�
�㨬F��x���҃����?��ڗߨ��D��M����^8�o�Jw�+<�K&�F+�2�_�Z\�ϰvф���Co5X֩�@ ˬB���Z�8|�Jr_��3R�1��uj`Q�:#���ʡ���Ȳ��7��e~AD�``������oe�~��e��l���IS�z��=�w�N:C�P@��e�H;?��A3)�X�hE���1�;堑Yk2w4��у�6p�����09��;�p�E��Z���Y4�� ���qI�5k�����Y.�����卂�Tmt]�v�3./2��(1;P����&p��N����(�/�_O�,:-�<�k�aD���D�E��5�<��/�iI�a��H2��#�^��za�#�R���f}N#�l_v���qc:�����p#(Rլ���]��hi�WN�J�ė�*��[b̂VmN��Ϧ۟Dg!]��p���+'0&���[xвpf��H�K(����	1�0v
m��9�o���!]�TVV�;�R-�X���
{�9�� �fSHiq(n��B�틎���rÓkC�P��7xQ@u����ur@��;j�M�q�쪥��QF
	�D��52�1���ؘ_��љ�*i��Z$��yx~�|<���J ��$9l�ܒ�L���z[�\���h�eli/�8���������}&�����\*8��*aZբ�Kʊ$��B��_g}�� ~3P�]lg��5�rH�$YQ)����N�؊�uU�a=��-�\Lb�>�[D�c"
?Z�Ϝ�o�򐕬���-by�䐠Y�%<L�g D-S���(aگ.	�����%�\��A`0#Yi�l�������FX��rywnu�@�\�C��ؕ�i_P��� �M���1��
yِ-fy�B�u&���S�W��Q�4x3b��Sv�dS'���r�&2�3�aY��aE� �<�s��0ܥ!��<lm��@vD8�������UH{Vi���QG����'��e��lJ�p���k ��Q\���a��N��� ��H����C�r04�ЩDT۱�}�7���B�}}���8�C�|���m� ��ѡ���cm��Z��x��Ff�s�QM���M}]?�{��e@'k��)`B��ap�zxp�;V�`Sd����w�ۗ�d�
�m��13��BGҬ��,��.=�,t�7��\�V�E��
�Ɋ�f��=�D�p�q���M��c�	�oWSFf�N� > !��w���J\o��� 4��CzÄκ������l��W��k���m��&�)p�_8�#w��q4C��4h.��DT;��C��2'�rJ����5��%���:��f��q��B
�/�u{J��s[�n���^�M�5DX1�����X\���l�(@��g5�`}C_+?�Ύi	nYA~,��55�*�(�׍#X�JɂaY�9����.���W �e$cm�߿+?��ڵ��N�R.,���ߠm�	8��n��0Z}�V��ɛ�-�v$��3P�9�涄�}�t�ߞ�}��y�Z���m��s�с{�2p�3�o�
������ߋ`��%xe�]�1_���@T�@���W�{ӱ�F(C���b�$<�H�O�I�n�08����r�`R\>��2�N�h�A�K���w�1U&�
l"' J���\|���AfG�߀��&\u�Dg�h>y����M2�,���T�܌�gHFÜH�A���48��K� ESՄfD�t���[1.J2Y糇�
���=Uf�7���-a��N �N�����E���������ʕ�*�������`�A"���u�8�&�P�━Z
�u��ih�����;�j�Ҁ;f����]��!��J�A}��U�����.Ў�go�%���-��/�\�+܁w�En��5�B,�g��엂Cj��i��B-�]��Rn�[h�$���*h�C���VJ)��_��b���_ȍbj�q�U6�C��B�����y�gZvqTA��F�L��V���H��fe����S�r���߆�	P��G�Ms!~�?�������a�T�z���
t7����7��d���g�p˵�t��z�/�p1x�#dqpK	� E�h��������;��	�ט��a
�SdL��T�^\�����n�Dՠo��v��^=�(��Wn�,o���=]�ڦ��=kn1��\���I�Z�u�Y��EZ���5�y��0���0?�oc2*[6�@��i��Wc#m���M)���p}����'�wh��o L��/ �ل!3���B��Uݦ�ٹ� q��I���� S8���߂G2���W���4�p�S�KT�:�yI
m=��p� J���M��fVF��o�'�>QK6�������&��Q	*�{�?����d��<��:6
���{���|�=aCo#�Ts��Y&�����}!.�y@Q�~���½kBc���^4U��x��0�ɲ�o�t���*.��&�ߗhr;T8?Lu%�g��}�xu�tdA�%R����D'%p���'$؋��*�:.R'�6o;;΋E¿�  ���|�.�4��!�4���p���ʨ�U���{'x�N�	�%آ�5"0,8/D����x������^[t�k����oLõ�����1Ϯ��`��q�&��K��t��W+h��\��Y������d�>� @a�h�V�[۞���8�0(��)��6}�e}�/3:���]9�ƽm�,<�4r^�6]�<�}�J"�Gc��FהÍ5�`���?m'��ǲ�rJ(��8l���L!Xw[�(�3l=�}>�$W��[U��PR*o2^n1� �?):3�ZD$5H���׿�$�u�͌/���Q1U`�M;+�
EoH��gX��pY0}�^S!В�|RH"Ȗ��������]����$u3_��-%���.��	�
�!=��OT�?8�h��ԅ�ʹ���*Cb���2C hⷝ%�v}Xi϶8��k|P��.`�
/U.�	�R�
����� ��}b?�����9�͚$�iz�,r��&��/X����js蜅c�'N���!;��%Ono=�.���Pw!Q;�s��-�W�J�Z.��#yc$‒�"��W,��u>M�Z��s�n攃i���D��d"a	�\P����d]p:(>[!(\�;	li?]|�K谥�k�%�4��a~�nĹ�U���Б{�D��8���&�Ǣ���4�K���|e�����y�C(�"���]���O1QLk�|?v���f~��*A���t��Cb��ঘ|QD7ģ��e�CrH�y�k��zr~�;>�)���3���3�����{2��Y*o�\���0���!f�U{<��4�-�v���7��E�;I�E�w��&�0�:>x�k���Y�f�7��h�6�<��4��'+� ����jgǥ�U��'P�櫤̜�.h;N|�F�!X	&ǶBQ[4A-��qq�K��H�7�Ӧ�膗�L�����fŧ�}���>' `�e.�'�
'���_O�N+�imל�8�$i����JK�#�f�ޡ2\�������2ɼ� �R�)"�[�a9v��~�ٺ�
�O��󙖈���k�hma����煭Zfi�b`�6s�pX�kO�ٙ8�@�;�i����z�.�s�?����lmgt`�/e؎Z4Kp�_MD|Ԍ|��9z\�֞��²�d�!��BZ!:��V�J:�4"߮Q��3a�Wx��km/��F����UF8���C�|�8+���1�9)+�vn1�+�K�'���%��\x�h��$C�G�9 ���;��o3 #nߏi�C!#~�����$OQT$>H���n:�2���g0cw�Yk&��k[x����
:U��fnn�w�;2�I�~��_0�c����{tBi� 	cnq8���6^_���u$7�M�=����`�K5+�c(������^�\Dn~��q��/L,|,ىOp�Ӿ�o�?�Ŵ�o7�s,���Ʋ+���L2�J��"�zM�@��\�U"�cʊ�Ot�E�%���������a��,�;'��12�/�Iܞ���o�S{�wx)ot�<G��ּ�&��wm��D[C\�*=zUݗ~��h��f�C�� ��C0�����\
!�H��!�;��Id�p��rG�s�AîH:%����ѕٯJD:�]����<
����*��/��VG+�!�NU��aՓ�CS�
I���E'�X@J��u���j������^j+�j��s���q�zc~��0A�y..�̲�$��*v�/Ϯ�C����A�?��J����s� �~�$�`����h�����>c6����_��1�c}�'���@jwSYOL`į�+5?��nkkp]� $�D�Y����o� �`�u�E(��	>����t�X�,IHWjPԛ���p���2$z�C�ȧ1�Ѱf��38�{̸�ࡌ�O�iU�z��=@ u�O��S�x��:���x�15���:!����W���#�!�y��T_�`�~6��f��o{���LX�a���-q?�J*�kv�3��k琲�7W���F;Ci_�Ls�\���VW�D��D?��:ɰ�-]�r_���N�t'�%(��%����y������@�ƀT�x |�Lɛ����_�K��6v���^:�n��ʆ��۩!�O��0Z�����+��f`��N0���ܤҫ����^�����qDe�p��C�Yz�Vni2*;�I$��1?� ��~kKl>���>ɷ&�뾤OJ�* uVä�UZ2�'>�C�'�ֽ��w|PO�CY>w�:����ĩ��)�?��R�s���J@cTGPk� g���@�`���mj�`X*Ǳ IyCxz�I�k��5��KVғ'͌m���H�����w�_g��Z"M�>*5�Ӄ+0��K,Z�Y�@��䟶����?�����	���SKzB��9,���BRXH!2�⯟����[���s8����e�AC������"��a�C�8Se��U�ը+�H	�Z�J�Y�qe棺��Ά� ���NT'а �=Q1:�R��9��«f�����gB�X-��ac�.��N�?tP�|�K��5sA�|�u�dm��ҙ�7��}���u5�!��_��f�N��V	m�=wA2Il8SG�;�P��1y��N�&�|�+:] m��/@Ȱ%%��cŲ�q�t`u��3R�Xpuv9es�Ýfƍ6�X��~&+t��7����ݳd����+H�J���Y��򼒜Z���q�NoZ�.b�@r�]�)���*�w=�%����Y>�ji�����1vĝ�}��1�Z.�����[��5��U�����jL�4�P���b�Z -�	F�~��f$�SuF��N;ەt�Y@'E�Ѩ O/r��LEA���.\���7P��v4�g2�in��#���ʂ�FN�Z��6�<zV_w��k��'6RDt_�6�N�z�mϙ~m<�I�n�;]Bh"��'����{}kh%�U�837��v�\�imh���@��"A-�`��}�f]g�2
�[��A�*I��[��B��9"H�v������Z��F���G������޳L+�՛�ŝ���9БB��I&SI!<o�%��"_+�e�I=��RZ���b1��%aJ���p`� n�=�;~yH����Q"�B-�'!fY�0�2��2���͌*���t�?��(5@��2v�"V�`���[�8�<���۬���d��st}�ǚ�N��Y|��Q��vK���?a�!�ղvJ�� (�Al�Sf����"�7Ӕ�r�!��9�x	J����f\:�����_�6<���R)MDVj-���}����ę�&�[�4��.�Y�Ml���4+�:��E�V�x�Q�-�6I�z闯�~(lO�U�_�9����jf9�/�A_s'����/���Mw
�%���v�׾�H0��GU"'{,r.V�9k�����D�	Ô�ϯ�&��8�M�H�2���B�l	�25�\�~���NaϬ���g�j�欇�͏�H\��@I0x  ����~q�7��R�ȡ���lG��8gvAZCHj�ښ��Y��gWbY *�W;�Gw�=P����ik�{��Pݟ�8���JG��U3x¾p��M�$��}i&2�m�ة�f�q��Yf�"��lذ�VQ��v�d� l{���
Y����5yT=.�s<�j9�x>�¿/�D�S@�@���u�(FW[Sp�����:�4��vR�r��<�fe��y�_	��ѱe\���;���k��nVڭ>�e�$ϔM��	��ve3Z�.�}��e�e��	WXԵe�-��Lu�C��D�T'�����&;
�����L�h���%�,��P�H4U *������{c.M��``ʷ��nl1��G2� x���a�'�����θ
dR�χ��ΌF3�/�a���F~�/��t��=���i͔'�
��h6VU���s#R)Ί���E0S�^-{��
9
���2�SgT��~��(ސ�G�M�B�mp�C:�W�� R���/�ޥ0nk4�^����8�P=雧�QKS��;���.��p��놂\�ˍ�
��Tnz�������]Ֆ�?�s�w\;`	�;W��Za��s( �6o�8
���g������6"�)���fI��&���FO2L�遤�օ����pjxr�]��gn�����@W>�
l2sC�+^�r$������Ԏ2i�N�`�i�^�E�ko��%چ� ƽXε��A
MDJ�V�dTH�t�o���� զy�PlbR�C�Jd���_�9�!<n��i���	B�YQBT���X�
M|si���J3jv�JW�יЩ��U���8\�GD��ݏ�{&į���H�4;U[ZtV���׌�r���$f�����M<#�O�?�vX�ti ��bD�3�lY��M8�bG���$��I~��|?�3�d�I��G�:.�a��\��x�l������Qx�"6��y��s/5��+�N>������w�A
ш�������J��r#ɩ��(�y�zh"��Wּ����,��M��{����_�i��3)ɥ@<��fϽQp�p��P���h����Q�N/vl�j���m�E�m�kc"��=͌�Ʉ�dSK~a�D#g�E�_�Ex��>���^{�˯�Rur������U�}�x1f�Ū�I��h� �z�q������%�Gj9X�m��&B���@�װ��
_|���vq�nR����qܺd;�ۛ��Xg�:G"�{2ĩ1�D�,��<%m�o�˗�V���D3_��.���r�]XJ����4�>N�'G�l�������P�+|d)zڑ�L�dV`Cc'� 0\��!��|g
y}�Ĉ����{�i;E�ö���T3LM«-� ��d���q��5����M�۞����7H6���T�����[��ʈ!�BxI�s/O_�^�:�'��ȯ R��1��$�H�F`�x
J�������ק�(�t�
���11����1.Ē������d:%9����{�گ�B�y�RGʋiɰ��R���K�cPd��ZPƠS�F�4�#)=��P���cF�&�BR��B:���o���lIY���d�&������`�D�}�x@s���Y[��¼99*:D��gl2�]��_8��v��Pse�n��:ea+�6�"Jx��P}�FǢMn��Q�ς'��E��������lG���Tf~�+4$�䬱��?����]5j�Qt1�_NRװ���j����N5���������P���2%��ߚ�������p�!�?�CZy�S/�m:w}�籰F�J�B���߭7s�c~�E0��SI�1sy�|p�>q_u��\8#T�3[�BU�D�$�R�igR�ҔǶlP�
��u~	�n�\�#*57y���҆3�f�:ѼKE��z�lYOΪ��I>�f�t8��R@�Q����a� u/��/���u{ 37Q:������������/42��S���"D��q��m�Fԟ;Ү�8z"��P3��{�E��? �2yi���K�֚�����;��X�>\�y�L3�4s�p?��m���:�]��ڊ\T|��n?�WrL�ėn���A�sʡ����!�X�"���%���JT/���T\@�6�t�k�]��A��ޙo�Ɉ	�����G兲�ʘop�,�����R�j���13�s-���*�۬g��h�[!���s?�	�J�l%t�d�:����fȖ��m�'y܃�T��%��\X�	�H�_��Zݣ�-����9�y���1:��X=� "%��>P�79ͺ6C���D�n�k�F���J�ؖ>�T����u��9�Vy�_ W&8*R'y*s*�?��;]t�-�q���4>;�U�W�� ���KG���zm�*n�g��u�>(��������^�f}7�M�HQ|s'�<���F/����m���:D-Y��!�5����h�l��Ql�J
�G	�����^�Y�����⣂weKs���Ӯn��ړXO6	�5~�eH�XJ-6V��S+#�D�:7�"֨[ ��N�7���[%��x�������v/{4~h8�HLIC�{�>��oE<U9�i��ۨ�ހw�9l��5�b��Ko��s"�5P���Ü5݅UI�y~��~����W:�]4̸��:�I��G���\������|e��[���9Jhx��u��
�2���9�է��5�D�|!�V�vx���T�3��u��@PS�AƋ[�9��f�]U�㵼X6G_K�r�5o���8�\Kڇpb��� �#�z�l�[,�r�15� �]�HV�n�a�聲98���ހ؛L?R�Y���X�](����/}X+��V%� �B�2(�ј�ii��3M^1$b�֖�G9�MsV�2l��Sм@�ޥ�s�*r]Jߏ5�@&��0l4�*pr�U�����t�s�P0�UtY� ٞ�V����1l�<�6bF��z��=m��7|+�NԶc��V��,_8R�_ ����o���L��h_�=RC��[��G/�y�{c�mduu��o�,E���ݜKkw�ʦ��"2P���8���b��N��w5-��,�5��M�xX줦M;�5�n���9tz�S �My���ɘ����i������X&{��0u#eAs�Į�v�wΣ4�RA�|]�.	[��@}ZE46���A#sL)\�L+�AP���1{&�����2�W�lȫ0 'i�%�s�+�=�Y��.)?�e6�p��s���O�0�W9s\�J�\�ߴ�������O/W�륺H4q�z$��<��]R0�P�Z��i�\�lF�G1�K`Yu\����{W�d�Ε�u��30���a��+!&Sf����4���K� �2����5���=�F3���u�,:�����abl��6�_a�G={�E$����9�t���=EM~aN24��>�6��,�Wq�!��D����I��7�q��7�zr`��at2u� �I/ѕ3������u�aF���C2"�?�h�1�t8CcY/����Q`O��(���9v���+��� _�(V������Ð�����˜�ޒIŊY�sm����a-ҽ�qOGg��a�Ws��$�wN�G
sl�ۦ�/�Ԟe��o�P���6/�k(SJ!{ObJۼ�Q�
���Ώ�Wt��V��lY B�
��;��Ь!-_�8��h�,Ca�-��d�a���W>-8@����(�6�l�9LM=9o�}�����g(�x��Ne�#��8�x�x����-�A�����[�� r�������������ݰ��|DG`RyB�����.���mƽUմ?0i��i٪P��k�ţ��Q'mJ�2/��y�~�y���i���f7��!��aB}��c-^'e��C7�cY�T���6���� �����&��Y�z2y�����jT����}Ә�� �9��3	.�(�S���w��`�s&ҝ���s���[��Ӑ�����-?Կ���P�[ #�`�CVI���q��Xk�GY}���K`���j=��1̦�E��eh��
4������G���o��j���U���@��?-e�H�XU^
�{;��"��l��B���'�ih��-��Qp��=NbT	�����	+cVPa�\�A�S#�ޣ��.��.dx2�l���؝��}w$��&>Z��������R�]8�{�x�%���I\\QX+�I,D�@��!�1��4��5��웶��nsMY=HC�	�J)�1֘����4���3I�uf5�,\t�^J&���0�g���T~��Ͷc0�X������0K���m�y�-��$��+ra"�/�ég1��A����O,f�S�F[���	J6˅�۷��C����.%�*yJ��!����,2e���W�G~����~]���*��E�
������[	B? X�}��>�\#�
��g\��Ff�A\S�9 =�	^V�������V�+�xlK��Zgm<JD��n�2k�R�f��۵�[�]TS�]��l��ϐ|}y�ȓd�*�*GK$�gv�!�������)l@m>��v��嶵������%��	P���
��59vz�<<K6�)�������r�¥�+Y�	"k.��l���~�Mq�������Z���Y��lkH��߼�����EW���{�����G��v���7捓\h�(!��?�s��g6B���lY�R�˵d]m���υlO�P~\��/!N�������u�'G۞�d�%�9kj"�~ZZ�M�˂+�0��	��:l���sza���L?��Pj��Rm��iď�k��|��XJ�4j?���P���λ��"�|	�����n�|p����8�G
�!�r"eq>23�� ��3IUFDD��j�7s7$��1�а�|.,����a��	#�Ah����'Ϣ�f�Ur&�zE��W'Rp��֧Eh �t��=�=���+2�F4N��ҧ��7�%z�=�j�RU���G3ړ�A���.e�>4�F����������3�]Χ����+C����pO����P@8Wt��0�	p?�{U�oy7�}:�9�A�êī�V�iޥ}��a�~6,T~�͙J��DH ����k��zg�������W'���A�G��.I#L�R��\���H��j؋nW�g-��[F-���}��^*�]�J�1B�k<�h� � V}pK�r�$�Σ)�Y��Ɔc����i�!W|�}4f�+ث�%~�������p*���Nα?�	p�e��D��2k�n�/��)��B�-g냒��:w�m{@&r�G�O���0�'�����v �f�.8�%�ݥ��Ǌ�]��v���|s��c#FX�D�m�\�ת�x�F~)pj_�-�"PQp�.�~h{��Y���<-�[L����\e�
�����|,�]7gO71f�2�/����q�A���f��싣B	�R�����H���H��:ݢ-M�7�4z��b5X�5���@ߙ=Qٮ���#�#l�e�]��Z�!�5,��m��+�����p�D9Al�fS��~��S˥I����?Q�I<��O;�{�މ�w���� ���kv�	d��YiG�i�iA�V��¥R1c���;�27�ܝ	�9��3��b�!��^'I�]���#�#aܶ��͖8�����.��ý��r�I��h�I|��t}� �Ѱ��[��a��UTċ�H�!�j/a�2uX����t*�����r��3��|Uu�>7��9�:	L���|�A;c����6���YC�S@���[{��!C�Jy;��[�p�|�o�/�\��ߕV���꒓)�l�6oU�)J�p`{߄7�k����1L��R��Â;\ݑ:��a*�z4�(��1iJ\\� O8�6,���C�:�}7����^I��r<�im�7_�I���x@��n�R�i�?�!BID�s[Q3��B���g?7*��V��Oh�y�W�(z|U>��g�D3����sq�u4fG�3��$+�V5Tt��R�����r���BM@��k����#<	a�Le:��N�۷������2bc�<�k=JC����81&|5,��{�R��r�rǍ�^�Vse��� ��Q�WE��~����X�emƁ�[)�����|�M��kf��"���kƠs�1��<UV/q�٫�	1��o���'�6m�`��5=4����P"��F̩��-Ͻ���/w��ލ�<��b�B�q�г�6q�_�'����� �l�hu�`V�䉱M�3A���EkM#BePpQ����(2�xZ[KÕY%�`��q�F���4?�i?ͱJ<JPJ��k��~E���W��7��B
�e2v�%t.x|?�E��R�Eb���(��tg�C08�ܠ��i�5�T8I�k�#Xp�
c";?��[I�m����O�֪��D�6t��3��b����YF��"M�[�`d�.	t�YY���P�E<.!��ڷ�����*w�i,h�d��u�։GlZ�ݮ�<�1�H����a���-l�S�+N�y.DGF��!�Y���1JQ�=?2����]|'&�������d���Dy��V��5����������[%p('�`�F�D�.}r�fv�<�Gld�r��k�2I���MŎ��k)�r<��;K��%Ϋw���7�{sr����-�<�� �0�p7�QB踩�������M���2z�	�jU��-m]���}���W���b���|12 +�~r��"i�ci�I ��xR��>g�H����8�2�bRS��cd�b�}Hr�����a�{�BZ��k&�̮�ˢ�IXm�LmF�ԅ�ly���8Sn6�%v3�R��I1]���E0��͞ʶhd�j��Ճ}6�%��T�<J;��Q:;.���KU�$X�� K��Ȯ�~�S�m���: ���ǽ.���A�7Mr�%�P��
V�V͐�ە��۱*f�N$�� �εIPP�����8TsҤ��c9����-�����@o�������}�)hK�0Q�n�����Y��IY�i�l��L�,X��ӕ`�Q�;Lu����e:��x��C!���eo��K�}J�@�j��NC6����L�X]��6���qb}p�'*^;4qh�D��RK�qhY$I��J%��ؖ�Ƭ��^��K�g��pO��eo�Z��r�?4!Ov:�����gG������cl����fI}��Ѿ��GІ� p�6�v��ZȺic�ϑ苳��b����\���ӨmV��O�� �1ђ��Q���1���}��)�Κ�R�������Z�_�g��1EN�bb���|&��i�F�כ��'�$ETș�[PAcњ����f8�JR*�f�H�HN>e-�̲��;�cֹ����[������jJ�[o��\�}`b�U$�!�cT\ğ�$�sM�&V9�* dhe�K����y��v���qJM{�
����jy��Ӹ-��UK�"[�s�.�5H��m�7f� A4�e�u�l���?�����z�sBx��#`�61[��߀����<"W$Ť2��0E��3$�n� ����e����t4tq���=����	L�v�N
r�{Pˎ��D �;�M��iA�ҼPZ}��}���3��oXύ�1¬���.���D���cǎ!A�	u��B�6l͘d���x*� ���)l�B\ ��&m+��	��!1,� :ZG�n�1E�T�^�A��2��n D]Ԕ[�����yd�A�gM�NA��wW�H�-r��*��O����7�g*���4�J��3B�Οp�ۋ���U�M���`��fD�R��KW#`�����%ъ��q�@ϟ8$�:lG{ <;�lS�!���Utݗ�J�7�t��ɷ^ԅ�-%󑽓���-J" ����=_��x�>ߍ�`L���U!����a��¼B�aw!)+ v�J��Q��b18׋R� }��f�� ��(tgw�z�������.g�.������O�c���/{M���#F�Tt� ����FL�H�dbT�I����t����|p#�F4#A�4��~g��2B��1���g �̔ ]���q�U�96�G'����.Ă+��؝l���>�q�g��A���/[7�?��HV����b��vk�	g����8/T;�d�Ak�ny�,�e���͎��/����tp������ <�i
U�:���|�I9eW2���-Da�>Nq�UI�P�wF>���A�Q-��0S� ��qAߨ����9�SF�sO@gDO�P���t�c�nS����RkY�:�p���Ŀ}|'�n#��6mm����y�K���5�p�S��c�ǀ��@.�q�q@��t�������}|V+��y�ڒ+���@}J����:2��{F�O�����D����{$a��wp�p��#�tc��KSxk�G�G!��F�3��h�g*l%[�%>�E'�'�}o�.F��S�hF�����B���i�}W~�H@�&�;r �d�Q��$�2%�E�
N�Ύ���x/H�ْ�G�CcIǁg��bE�Ut�i��=荁�1�Rdaŉ��*n �m���a�C�$MS��K����o�u��w0.%�4t�e.U&XIĜ��k��  �zB�޼{���&��6�{�>��/���k0�m��m*~�Е�D����8w�1�Ēc�#M�qX��m����>~��S��,��X���r+���A(j�ǡ\��nӠ�jﳉ�������i&(wC��$���\̾��}������0�ֳ�O�mt�6�� �^�7�T����N��nH\�r��s	�I�F4��2!/|��InP�
��w$�·��u}+��c7���i�,�ƜrZ��Ig�6�'��q�#fx�"�[n�["�}�
ΧO�I�@c���0����	���\m�T��'�,�\pP��S`�s�Ø����u�F�d�u���<_	���e��ǫ �x`��U���߇Wݓ��X]�Iڱ�֘�m��+���BH��iq����[�7{����k���J���_�i���ʋo�"w)>w��<�+������uƫ��p�p*YV���B�@�����3ä>з��t�uR��#�ʗ�x-�.�e��4�Ԯ��d�2��<�&�n#,Q�IC-�!�i���g7�f-���T��~5�E3g�L�FI�{
�A��"O��NG1|��TQ��K*-#2=�t�7y� '��w��΋��D��RaC/��!}�N2g� O��T^:���wd�/���h��Y-�J�Pu�RH<�H�-�`�PW.�����νWa<b&�6+�9��Q�hH�|:]��.lv��^����so��N�!DrĘA����=D��:�]���q�y��gW���j�L�K�|5��vl5Α#�w����u\�pV���x�R r���0i�s �Ea<����$í�X�T��s~�;�![z���zW�������1����֊GqN� /z� ��B�9ϗh���8��q?�]�̌/c'���XH[V%�uT1�:W�)��k��;�s�E#�=8'N�����v��q�qc|���&����v�]#h�E�Ѕ�D�D�����+�߃