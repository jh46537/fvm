��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O!) ���Y�Q΄�O��*Ȣy�dsuQ���`�Q}SA[�.���(��<
vɼ��;4���͋s1D[
�f�T�[��h�K�"HO�¤�TwƜ|�J�tR:����p�#��;������A&�K��HȮ�!!@<Ȍ��VV ��k��ko窿ae����ZS(�F�FO��2�;Z=��t�)W�{yo��r��(�K�StcN.�����s{P�8��AN�C�/��~Y����[#�z�bEB97�'���?�$'�����ِ��ǰ[�'�d�X�������%��`r��`���8D�]�At���w	V�򴴌���R����F8[4Nj7�-���ιFUEp�]c��$W��9P�|�Ԝ��L�?�9�8	^rA�Ƿ���.�He���n0�u�+}@I�2��P%p���-���6��f�8Џb̝h����喥e n/&ρ�1��ue��Fw�����s���Sܿq󀷀�	�~��ݒ�-i�Ȳ�G���S1	�g��<�ד��f�t0-I���:oۼQ gD1M隬it�;y����4_���TB�چ���thh�bL0���]q~�����4�Pw��Du,��8n�,�045��u�3`G��볮��"�W����`�hR�u��yI&n��xc���&����7���W>=���Ű��T��+�ς7
�73�ȥP#�lm��"8:�K4�j��c��<��d�eA����
���&c.�nP�	�hy�Q� ��l54ꓭ��ٶ���j'bz~�������,��������&l$� �+��D}�4j̢�0��)z���#ef �2)AuO�3�ۉ��p���s�l,��p�J\W?��sk\���k��}�a�.�.i]�q��W���o��9�����^+@���T�ӷ1m�$�X��<�j更�UGk�y��b��}���8uw�h�R�b"㕑I`}�0B���B��v��u0ۇ���A@��D����N�Zۊ5&] ����I��-�K���_å��HҚlL#��^�p�wo�O!�`'����^6y1^��m��7���s�5���"����BM�&+��#��_����'k.�A�$ʎ����ąI�4Nj�^��Ⱦ��4�e�zg�J �Ty�hL�%� 桐e�L��ɏ3�jyBh��ߕtͼA+�)Y-��Ż��/�xf4����c��tBn5m*�:-�Ξ&,��*��%��EϹ�Qp��������C���R{Z�"��]>�������$)}�Dy��QU��U>�[�x��QQZp�\i�K+���iչ~J��nԲ�19���y��%7�#�]ԫP%c�����DF���
������yc�^AlmXD�$��P_�W�� k�g���Z��(g��P�e�k�b�����٪��=N�1��+�)Ȥ��E�<Cwr^��<��h�U�74P�Qvq�x�%�}ӡ2����fkH����=c6z���Զu[�zk����v@ٚsF�A{��v��V�מ"� �3k(U)"9VӼ���}A�6*�ҊX(�	l��[��3���E��N⦜���n���iOɫ}q���,ދ�	gЉ��6ï�n	mvNw6�wނ�A���w��k�W�|�0�v�k=�Ö���s�kW�ر�LǶ,��$%Qi���Ʋ�R,�y�
|k=���2H�p$&��"RRvw�,x�S���Y�����]51�=f>!��R������v�ܝ��h�0k~q>�ߓ��S���M��%ޣ'�2�U��V+��T} `m��3�Y����ŦȮ���{%�4�3�%���^�<j���0WG�Y-��Vp��G�B�ٮ6�ZxL�I XCV���pzM���ڃ6f���Z7
M�~Ƞg�]�Ê���� b��������׃J��Yh��pBz!7LS��V-�`���"��C����JEl���qJ������nY��WzUK�na��c��5�:	�r|�p��Q���]���C4� p|�g�r��xo<)ւT�x�8ѮL�w&�C`���Ok�{�D�%ޱ{�&�)�5��H&e��Ha=�B�� 6�|7n�n�ɭعű���@_���ڡ���Ǎ�
�|���ⱟ�����j��$�Y�{r�*��O�}�c�KzwL?ҥb������e�Չ�گ�E����d����X��`��s�,�cXC�A����s�댟t��T"3�����2>ǋ������R�
�j��4�(+(�(�M
[�$.���i��m}0���yC�˯�b���0� �=���s5I;���{i����l�I�$�D�!����;��-I~��S�:���i�,!��{	�_3��3Eo.裝RN���.�v�($��Y�_5�w��d�$rNj*���FM�E����%X|��\��P��RuT�*t��-�J�5���X�w�$��[�n�Ϲ��ʓ�t�j!౾�a�i�.wp�6)bx	"��46�X��Y{��m1-� �椈���ޠ7~�*R�����\1[�����p�e�
Q\��TNwF*����ip�Rs����r*r�J��*�bWJ�7����=sSw�� ?am�(7@��O��mO}��V��l��5�����̬z����
}�j��=0�0�����K�x�ik������KWJ���A�]B��Y'���{�ߗ��M��(@�33T��=�����fr��g�N�Q�\@%�����&I9�� &�[�ZG���,}ȆǓf6��(�Y;G�i��]F/2	g֎�l*��nG�D���K��n!�*��t��ʴ*����%��"�R���Z�B��[T�s�O��t^�?����������	�3&& ����𳁏4n�gD�M�"���Bێ���tx����/F���%
��ӆ�	�{�V�&⟙���ެ����I�}�F˜x��+i�i ��z�+�
S�Š9�y�9�����t+���I��~o��B��0�O�w1�,�A(��^�l�O�R0���1e�R](�d�}��6^�YJz'2�����H�[��-z&�j�#b���ջ��f~��WNb��L_iŦ���ݯ��q��� 2��g�H �f���}2��ד�V�2���]�I�z@�]<6�y�ݑ�6��I��X�Gy%�ko�8��n����y�a� v���G��ѳ?��2+q�
UEJgS�r�+�O)R(8NR�K]��2{��m���	��b$<mRc<��#�<u�s�
":�*J��3�ddz�%��ۢ��.H����ŰM2���k�-�z�Xv��ɧ�k �{-�J)om�cT�������av��+��%h�ke9�̀�zhtw�9��~ol&p��൓�O�O����ڟ7�Qa�En�=!<.7��.x��E��������	����y)�@/��{�����$��o��d� 
�Ƒ:%��O��[ΞC���n���=�AVF󉬖��HVhjCӮ:�-����J��5��Y$�R�q��=�+i �~~Ȕ�Fo�>f�`�0��'m4�?o)z��(im�BC��+��/-.}�G��[5M��q��ʤA��v5�^$��x�UQs�6C:�$BAb��Uk�ڕl���|  M��Ԃ�eWr�}�D�C�I×1\�4��Ej$��2����32Ӻ�v '��!�Ez������rk2�*k����)���X�h�a
K�9�/B��.��3CM8��Mj$ާ���{Kn�z��U9,=�!�����ժ�M	$\.��x��m�X�#0�K�/¾�	1J ���K��9X�2�u
���8�`{�I��A9��)k��N�]��ET��0���e6�
�#�3掶��y�{aP4�'k�	)^����FS�����+M�E.kq�7�`��0�wcf��ރ�}'��-�ƼV�ب���;v*�?�~�pJ�����&�<z�����HB/���f�l�ehh����,����x9��~5�w��H�v�O:���f*���= Mo�%���ap�tXM��=�9A��=}+C�q��|к5]:�vɴ�v������_|�
� �Di������h� �Q^�U�vG-c��)�sU�)��@�<mwXüt���|�y�q��ѲL� �?H�xux�Rk"����Q[�YE�Ǌ6C�5�����ۆQ#F
���#N�u�mo)�����]�6���)�W�	�����G��\�̆�1D���u�_�>йw_N���*ho2��e��[��C�?��r����t��u�5�,�'�oF��-�!����3����t��q�p%�OY(G�E]iC���0Q�
������矞;�;a��:�g��|���)��Jx�c<g��y�6�6��9�S�q���B-0ǘ.6��7H��9\]{�(�齀��0E3@�H�j�!�3��J��#Җ�\�[;\9
���`tD�$�锧'�Zd�8��I�n��~��g���rO͋Zq��l9�DJ(Mb�û�@��(�'��4��B�W���w����$.�.a��%��zX���
%�\k�o$X�\"�)����7~=�4D�dWɮ��M���}h�b������4B�����`��`+����q�
j-�~hx����,5)�Sg|�^���S�~��Mo}���3)�j�z!C�P�,S�[x�����N^�",)}��l��SC����^Uphg�xϿ�W�*�O�_�z�Ç�Mg*�vsC�-�վ�L�s��Re�3����o��B�ݶʲP���4�[�Ԣͮ���f�qA�T���z>�?�q�x��Y����lj�N>paT_�+MqP��1����J��Cn[�G8���ڐ����a���+��l����;d��ݎ%���"��ezW���q<NHS�J,t�at�BĮFT�K����D�FU��o<�7l�����q�rW��"YO]�{��T�˧cS�Z�����y*��cDD�UB��5�����q z�q�H����鰊�ܵ�IJ��=�����V�e�<Y���+҄�<U�!�At�cM�6��$��m�
��w�-�!5^yJkeR�{�^?����`�$�oT�y���Y Q��YL|�+gI*�#�~��8��E윦I��N�-�m�e+��N�p5iX�T�b�RjE�ES�o1.%'�G̖�]~jCS4��u�ag�2.�CA�� Ė����W{�$��ˉ���}ڰ �'"���Gt��
�6ݮA�FnP�V�c���9�-Ђ��x�&����h�8��(,�sȲ-7%�������N�]�v�0�	�])O�(��qY���p�IH�r�z����X���5�}�`������=/��1ݖ��F�?F�	e�B]��l�Dc\ѰL��h���vNx���J�����`%'�@(u�i
��|a���Pѳaz�~}�n2�����9�!j�'M�ڑ������P�C�5L��1{��}��0��2:���H����AI^"�\f4D<�[*q�i����k���	b5=1��]�I_�ܨ��2�����������PNw�A��ݼ�{Y	�����
3�d���Π�"��m�c��i���@��Y۹:�:�so���@Zk��O�����!7 8��\V��(��$�����W/�թv龉����*BvQ3%���Ϟ��~Z&����yH`ڢj�v��a�IGe�kZ&����P�C0��l����ӹ�c��-!�jo
hu� �ɬ5��?�0r ���ˠ���+w���8^#�,��h�c��>�}7� b?(8r�c�Q�}J��FjEs9|�|��J��4��q�S�8���}�`|DGH���<!'Nu�'M��q�ֿ�a/'*������?o����0��E̙��Wj��F���n�1
����2�kmw88/o	��5�a�.��@��*ح#�:��7�|{�AQ�Ieӑ17�{����p^����n�2�uz��o_ly5�q���R��J \x�ZٿDt��b�lɞ�.fӂ)+�5���V�ܑ�p�4iV���݇�;@�n(��s5^��Tx~�"�Y��z���"|�Ŋ�㤎�I/f�=ILU��a﯋�|��mM�l&����cLPx"���T��E+
�%+~B�h���u[մ�<e���El9?\K��(���w���8���.d!'�n}�Qt`P"`�t��`RB�[�U^9�%=	k	�����OTe��|[aj�C-�\%��ʉ|�����e�V,�%�3x-�RC{�hu��f�w6�M�StZ��p[$� ��ƛ��㡴�z.�󯏋t���>�[�[��瀙��'�I�=���7c�+������<�&��=��I}7�ǎ�9�Ytˤ���>!�a��1�	[1�{�=c��׸G�l����<z	F�ˍ�>*Ȗ��t)��E+Ph�i�������2$&����L�G�[!��n���铵���Ϗ[���ێԘ�W'�����Ʈ�]p��l	���()�r�9�%��_�\v��#�  �'���[�XX����Z�BZ�n䠩�ODL�v���B�˂�o��(�"-�H�_e�����"Y�}�B 뎭�6�I�J'�ݳs������~k4'm�ꠢ5�2
�GM!:���ef�n���/r��ڝ�*;0~g+�X�iO�(�o+�2�4`:㒝���!�{ֳ}��;&-���iF��m�z7#�?�(���g�uq'��i);\�J���3ϝf�F-L����Q�OYS���x�$4�M��4��8��\����>�/�t"�۵O�$���-&�f(�)Bَ-y��+��8�������,�9fw2�?d`�}j��eۍ�ckI��^I�K�q���KmgJ�s+:QX�>LC����o`U(SR���&�� ��3�,xƩ��fYӰcJ�A:� ��!	���d�\�*Zp#p0� ��#�Ȕi��蒔�Z[X��r���
q
'�c�|���R)	dt���A�w�!tˈ�mw�)YhC�n�L{!.��==c��ˍI9΢�ʏ[�K�
�[�g������-tgw��v5Eq��f����"~�В���� �D�vcq4&��O�$/f4���/������j��J�sׄ���<��v���I1�h��ؿu�,�{�)�X>6�~޽A��!ڟM)�*�$���r:�o}��,���Pl^�Rd�?��;2���Y���X*�Æ���)&m��+��Aq)���2@Ԧ�ta2<2��b%Fw��h�v7���̴vqy�T���K"�\�W}Y��������G�Cۤ�AJ���)��Dg��3U�C`��@����a�1\�M{6�Z"���]+=J���K������e�H>H��v�P�"s�6�r��?S�H�e��Q9�֘ۑ�dz�-�߽���G��^�0uFA���R�gx">z�w�8��}|�b�5��I�X�b���S��K;ڻJ�`K}vG܋Y�]��N���I�{�K!��R"xɋȳ���h����H:1�≂� CeO�G�3=�����qY6����O��%tK�^F�	;���d\�2���N� ���aw�<=z0�ѕwT�K�Û�W�����ο���Q�=�ޛ㦂����򿺟3n��?-'�e��!��ObVm+��gEڪ�"V�'`?\�xP�3!G���_���C����,�,)��݇���X&��#�7���M`wX���ѵ��P/�)�`�\��Z�{n���k��i��b�=�����reY ����5I)��h�I{�,��)��^{�&�	�Ҹ�B@M�n=CY�jߔ
�R�4o�oa�d�|�/C޹�����%�hy	B�
�ۆ�,$w�݋���1%� �Z°����U����\���qA����?��Ӄ��#���s� o��c��5�M٧^�z-b��꤭pˌ� ��I�o�s��͙;$l���� �h�D����?��d!Ё]��r���p����L`�����OBF�Y���m��&n�2GA��=^�ՖY5��Kʸ�CSO& ����. ���h'��ۇ4�w�"ι��+�,�	�k�����8���^��.o�@�{�A^3!=���V$���n�x�p����߳pƺmZ����t.�5tȺ�����26������c�%��!t�7��
�r���_�F�;ˇ�ƍ��m�i��tJ��w�HGT<�k�Uq޻5[���5���t��8�^��w�7�A�9|�Q�S���VK>�d�t����'���Ć+��k�h�Z� �3M:변w�6�ת�肌m�u��wO���=e��rG[c7���d����+w�k�nI�G�{�Q���%E�}�p]=e"����ꖋpn{WQ\�����ڥ���j��QωO;w�$��/��\|�8��r/ ��?4O�>+.�-��~�WxU)��Tmqp�����t���TͶ}��s�O�B ���$��v�:�4��>U �٩��S�o�,�c�65-���)�V���l6}Y"�����nR�'s����œ܄ڊ˓ �:���X�+"��ᱽ?ΞRHZ�)F?S�ސ�x���]�����ϲ����s$�l����S�����*�H��M���^�4�#��3���$������.3�+���|o�8BqB<�Ɣ����FݦՃc�OXY�P7�7���..���VH�	�L[JǋC��FOB�ߴ�^/_��aa�ʙ��X�d8�!���R���N�*�$���|�6�=>#�9��7݉I}Vͪ�I~!  �t��i ~?�ͮ�p��0������@�)R�2َճuLg��d���U�8y���Y*�zA�=}���O�_���������it��Ƿ3�c6o�(g���!�/Q"<ad)����g5P��OϺg#���*�'
�p3L%r7�����!��;��NZMr���7����]6�����e*f�G:�諝�	������+�\'�{Y�=��]>��O8s~������l��h�9�"��D,a�P�����Ov�b��g-ˬM6cA,͕�3UpSƸ��%��
YQa?�1&��Id������d����GL{t,Q����QH!�$\0��j��5;����r	���K[ ��/����<o�h��zp+*�f���f�tM.q�X���(#Ѵ��RW0���TS���P�� ����(h�e�	a=K���Ta�Ă �`�?h��B)���V������]�m*$"w�a�/�xh��� {���[S�؋i�<ϥ7@�ZPKy�Ci^���}�o�:�ؑ�Py"��T��JE�� )5.��jWJ��]�5��@�(��IJSX�B7}�ݼ_��,���}�qzf�X�Lc�m�x��"")��Ȁ�V�g =��)U�F��W\W亩��U�0+[֏����I.��W���x�����{�.�[?a;���P_^���<`������l0;�u��l!~�̢{�<}w���C���\RJJx H��ۮd!�ވ�xt!gY����/�̃��EK^Woّ<m��m�Q-X�ڋd���^��p� *�&M�߭�<:Y 5��Ciq2+���[��ׂ���tu�ZH���j�X��k�����\������U��3
��������]jg�X 07��}2�=x����۽�]?��%�@�9�=��;�D��S� ��֋�:gr�1A��B�]]h����RD��MƶiY��2��}�Z�@:ښ���"�Ĺ��8?�d��Xl���*�~Ax�� x%��(���q
yQ��dQ�ȒP�3ß�<������
�~4�?��s�}N	G���C_Bݑ ���
�|�������=��Pc�Ik��M�>a���R��d���YB`�@36Zd�zh1d�:�����4�^8 'V�y���8��sa�W-94E������ѣ�đ� ��>�3��^�HX&��_Ny9V��A�*�����-E��t��!dwd����뗜/ҷ�%��q'�"�@@�3������n�ID��b�C��Z�J�c ��`�0@!9x�%�@�d�L�,�qe!�;4���X,�!=Q3��k���j��T}��c-�;ȑ%������ �L���3�1Z��\�pKG��F����=z��*�A������t}���л�sٖe2�k�| �4ʬU|귘GIk���<�����9Bqޏ�|�����ܪk���!-�^�.I'�N���B�Z�k3�ϾO['�������&>�G|T�վv�z�{��:�C�z�O�^֔�M��9&u�=�����r�d�+Q֠+_&�e(�_�b$�5��L�E�E�����9^��*��~f;E1����� ��}��M	~�m7 `:�.J����m��D��pp�Q]���
gޓ4��w�N�#��߰�E�~N��_��6�E��"�UN�8)��K�7�$��7ˮv�K�aks^ԇ �����/ֵ��Odm �o:�~�#���q(��|�����`��4�&]h�_�?�����
�	'��d]��a�N���3��\c����̐8�l(X��u�[ V�Q�,�ć�Qb��W��:b{��#���C1�ٚ(��hL"�n�G�181���b<1����QAkV���rQ�Ue)(���=�`���L|�m8QR��-�f�b���\K�&��Ż�xB���V�6@�}K�@��i�� ��+�Au�.�zb.;��-�3�(2�;�Q��8w����L�q�<�