��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�Y�f�ʴ��d�m���8P&B�� e��#1��O��+}��F)%"k�+�o��>��5�T����S�bM"�d�J3����40wG�;G��H�WKjU끊���Fô��ơ�%�X�`���/,
+�$p�$�s4�s҂}�*�T� ��Dkz\�3������1Y�q4��t	Vf��'arK�re�,:n����6��A^�.>S������fP��/	�r
�V���P��nhX�k ��ʙɇD����P�i܈j��%r�3����v�pQVSp0���X���4?�`ݠ:� o�-�9}"啻���,�T�~�������k�T6���O�����ͺ�'�~]�k$BI�V����y��\|��G�r��?wG�Id�5�����-�ܘ��k��
��"3�����XV���!�߹̵�� Nu_��\X�֫��K֖�jD��1�@�xc�ފ�^5Pw���觜dpΕ2$l�i�kKex0�m��/��%&�`�I�����-��}R�mLl�""M���X����+da�o?��L�l���6$��>s���`�K�|�,��Y&KA�~F4�����K2�X]��Woz�[X�;P�����
����,�B� Y�Q�b��X�vk��ȕ9���aKM4�I�:����0�v�d�4��^�_��q�f3���F����[��l-���ʅ#0"ƭ��#�K$��N����x��V����[�k>��g�/7�៳	xN_�Uu�#%�d!�a�x��h<�����_Dd���+kĂ��1��R3�떻
x7M98Y��a�L���B\Q���*��e�$��u���@�8\���☍&�4yi�r�RC}+����fU����q�r�w�е��xԦ��a*a1i`rUXIY��}M��z�|1d.b_��-W�-8�i2���R�Q�~���P!ř�i�</CBw�q�"�%��'���%l�n��Ο�#S2vT\͸�GH�!��,UN�	�2C�W0�X���U4j#������@Y�/�>���@5�!���R�r�[H��w�|���F�ӅT�X��}�Ӹ��n2	@v0�4�]�P�{u[�z�7� ]���`i���f����p���e�7Οe�Lw˓V|/nE�5���J�
f��`���w"<�`�9�����6�8�L�^���!�Ϧu���}ϡ����'۔���k,�N6�(�Ŗ�[`����,�?d<���$��"G���#�W�h�Ͷ�t���Y��� %p �*����(�6 }e�����E��9'���c�ְ�\J{B��-s����GR5��$m����gșYҤ�?AS%.���@:��`�(��o�p�f�8�����xX���ɑ�������Iik����`��� �y��Bm �hHU�L�+"��B�q�8�g�|�h�좇��\)���M��]�<�B�ۚ��k3��e���-����v'3Z+HF�S�n���p�sۏ�X�GZ�I-V��2�����b��;��ō%��9_ƈ��؂d