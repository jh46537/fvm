��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	zON�0sǏ�袭@���4C�;>��ʛ�a��Aؾ�lW�x�ғ-s1D����HR�uFSM�����2���=��ĆC��1������\����g�@��u�I͡�+��T���gc�H�*Z��H��C��p��@�g��b��yH�Zj�a���r.�C�J��5@M�q���nc�E���h�g�A�9���禫4���0��>��i����Ѫ����[l2�)��7mE��~��$}����������:���z �Db��oW*��GE�u}Ȑ�����ba�4�g�����{�`k;.[,����j�d@?�r��K�i����>�;�i�t��çQ��2��3��ej�b� �paL��i�6#��KQ�r�y�,�����"$����JP�m��g�i�!#��Pܧ@ &&p'��Z:�F䩿���*��v
�͸ 	ȹ�ZβP�]�� �UGe�ow��z$D�j�w�y�
�ϱ{�|K�SP�9!��LE���a'{�8Ϧ���vGf�����(E�>(��4�R��ʹ?��|ڨ1a�@�}Q�8J2�LO�����b���Ι�Cu���`Qp9~ �����i�����=�b�������n��~"x�@��{-ރVa8B����m�H�8��"p�q��q5k$�-������F�bi�~nb$Y�f�HZ�6m�]Y~T��7�'�w(���.������6]gkͽ��Ed�Q�0���p�U�K���%3��Q
��|�2�e�-�fG�XUq�ao�tC� Rt���Ƴ���!!�����_�I�п��\�L�CbdP����"����b� Cj��������av������)��2dJt�j��'��W#ޱ�h�*q�2�4Qz<:w��[�6/ �ؼ\���A���b��K�T�u�e���nf��XRZ�g�"`0�C�ǡ���I���.� ��5��T���|�/�Q�EN�w�����sP5�0�+~�0>Gۖ�ϫi�ʣ$�AR��]"��D���`ց�A�.��O�L�|���X��Q.��z{�����BܣĖ1���m�H��r�h��@Eoi���^KC5
#���
�$��ҊHY��H�t|͸�i���d�=P�)�+=�F����<��3���f�6|�xm�(�l�\K_��~@/��3�����#!��~V�j��b+'�����9�V��mİ�����>>�ƚ�wA�4g���������*;��[� ,J}���<.ڵ�=	ye�X��m�a�M-����:)�JZ�	�J��c��
�Vɍ*3���ſS�(�m�k\������xT:|!}�?8Jn�� �R�L�����n�!w7]������u{֒����l�2F/T�!���:�/���tҝT��D^�����2
�JH�-H\�W��Ŭ9N���y�{�Ĭ����/i�*{����q�I �?Z��${� �ɨx�+��4��޺�� �Or���ˀ�!T�n���5�'��~:5B^ka���o\��r@C�h�Y�ʎp�bS4�'{��O��=�P���ҙ��ZC4(�	��_����:T�y�T����]�=����߸�rO�iu*�c�F�s�
q`�M�;���j�ofj�N�p#�k�����s�aL��wЬ+�eB�]�V�'�W�@gS�l�3v�u\T�D� �ΰ��v&M~��'��� ={�kkU
�d�hS��;7�y�)�����%v���� ��S��CْC�^�dB\w�Bd���e���Ic�{E@�%�w��U�#��>m�q
�pݤ|��H�1��4�p���z]�ۛ�'4�9�$�d�64^�;#��n�"�𢼙�×���a��? 9 2��g[�r�c9CʟV�4Ռs���c����8~Ȓ�^M����
��L J�A�36�	��.Ǝ��}{����N��w}sջ�Vv�5�
�������S?�4�Nz*���B��)�a�b���z�D��X���07|�i�^��^�"l0�g�I�PS� �ؿ	R_
���6��y��̹.�t�;_������r���j�[ք���Sm
׷we�Q�N|�H�?�,���	��:��֠>�x�$7Z���`,ơ��h�|��S���6f��"z�X��}J��Y�l�{/��}EW�>\D瀫�	)9�n�K����q�#K�$���4�))b�97<�C��ų4(/u�26��:�v��ѥ�U^*kȽ��M�в��	H��jw7i�.�@ϝnfz!��>�_-�MWD��aJ�ѓI��.i-"&��+��@���&;�DW0��A�3}�1+�JL7�2�?	Lް��Bb���rk�}9tr�g�ְ*�,��>�3�����fO&��?,�L�T
��[�`/��t1�P(�z�<��i]�$��G�L�n
\e��j�byN_�xu�}�0��Ԯ>_h� ��I��u�%g���S^�����j%�Fh�$to5��������ǲ�0�ʡO�<S��?��r����N3>�DU�(_7����^� N��}����a_��j.���o�TtJoܬ�[e����e�ʉ������;8��R�����j$����HG�pz:���y�^����iS��	��wY9���N�̤��<Ayͣ�3*�yqp\ŷ�~��B��U̴jz#{��X�����"����AQY��)Ա!W�-ۃV��7q��Ca�5���fp�a��M�.�tT;C��}j-��lqBm�#�`O#*��׮�2��=�|����{���a��D���� H�B m��d�"�>?ꉪ.���-���e�pXc�&?1�o���co�_�����S�<=�lE<�>MJOEQc�W���r���e��٦�	�VρF�*Y`%��¥P.��='=���`_0��E�k3��У�~'���h]; �8Kt�%�k��v|�|δ��$J�&�����������@mgR�(i�����/mpQ�sE]�
���v�$\Le���JzEEȄ��z�8�u�!]~���`�Ay"I�F��ϼ���s�v��l�!��e�k��{�JᯈL��Ȃ�)�(�O�����T�אE��|�1e�Wl�㑙.�w�6��AH��rm�4?*^��90{�nD�NSGwe�lMH�q� ��r�0#O_�dm��;�Mr��s�d~���&�d�4[�+5��e,Z˾����4�5m���E%lQ!���u&*�D�����S1��YΉ��Q<h&u[��rm������C�A�L�9� ֛O?5��`h�U�c9���ВR.}����OmU{�q�ʾe����/4=F=?�4^oL�<����2� ��A>�ô� w���-$���^Ĥzۂ^�Mm��E8�{l�mX��WI9�I��+�72�:�H	��y�SK��;(*�n��x8�rM�jp�[Ac6�k�W[5/�8���m@:��)�v��Q��@�ߕ��?(W��p��0�V��u�!��{�I	��G�(�C����M��"��O�l�z_N�Ƿ�z�
KB	��\��'����Wa�韜\��Jt�2�&�C�:��T�exo��Y���5�EY	e�$4�Io�a�I��52��IE��{��S�90�Y��s��Fc$��������Cͳo��6%��ZE��H��]����_h �i̜ѻpd�8��[�IU�8pL�K��rw�VxӇ(�wW͒b[}͞�&�����N$[a+zp�~Vu�}��"8a[X����'�S��x�}�\(�pg�ZC�9��f1�*��0`b`�Gݰ�hd��<�kϑ��j���r�����D�=��5�Zp��Nuq�g��_h���?�˒:�o}!��u�|e+�7�^X��D>`�b$u�U?"\�+�m�i�Ԋ��Z3��6K��v1�q���I$? 8�^+�V��h��K�`��#s�Pn�ύJ��E�^���D�;�I2cr�~���{�n[�!"��k�g�a�
iI��R�R���/;(�)P�^t�8�˯���Q`A��j�+٢�אּ!j��ڤ���Z�a3�ˉy�҂Cj��h����/x��O�F�|fD� �����e�,i�/����St��xcs-�����1�+lW��#�����ޢ'���W(���S��	������+�`h���&��и��`�M�d`�Ђ��l��Ř;{."j�0��=`��E���e�E�Q|��e��������ܛ?����zOov�KţL)Q��M�U|<Rю�j�����������RaJX,�̧��ϯ�=DtM��EO-�`�4��(���4.���-!�H�x��3��h��8���Sldj$�7	�U�ػQ������z/� ��s��`�dd�E�B�6������;4�GO���[VE��i�]n|H���"k;!A} �n��t��\���̄&�l�RF�c�>ȹ)�t�u	��%a�F�b���˽�b���M	*���],H�V�Rd���q�1̃�X�?I��²�����!�|�zn8�չБSG̓��5D�V����p�t#�5�Y���BI�xt�OE�1�s��"��I%	7%��m�ݬ��H`Jr;����Juz��41[j��0�ԥō-JMJ�öqg�-i�m�o`�'�9+��ܪ���ru�	�o��}t��)������)A�o��gR	U����hl��>w[���2,C��h�xe��F�A�k 4�
1'�)���iv�!�ٛC�vY6M ���U� �����u�Q����v�T���xL9��7KiS\�[�t�*���m��D����>˛���_a��A#�O;ߍ�>v6�^�����B��9��
��
���o���_��`��',D���;z�m�]s�G��E�k�\<�1xa�3�!�ht��'�<�4%cr|��jR9�/o�Z!}ʂt��k>�Ovn����.i��4Á��y��8�|��-��������N(y
azV$�^��N��bp_�� I/�m�񽻷sɸ#ˬﷃ=L��@7#�_[!�=��&c	:N� �ZL�.��X0�E!��U����-��B�?U8dSo����Rɿ�4)�AMd'�O���v�ݓuqN�SѓhT����v$�3Q� !�	�-���r/ �޽�?K]�b��^U�����1W����fǅ�/O��QQ���}����t��*�Y��j�<S�H����Y?Rlx�W37�䱍(�� Iti�ŉߛ^�.ؐ;`��ss��쨻ɺ��Mz��b ��֪�jJ��m��F����V�da��-�>YJ�㠹$�kUay���n���}_#=����U:	�yr�娭:�z��WT&��L����sX�9uT^3*�86�<`�)Dh���Y`]�F��ٯ�4����7Q�ޟ�r�f��^5��6*IO�L>OT�pNٞ�����Gbm�)Xi��G�^�	SN��W2�Xv��}�J��|�F1i�C������O�;�T�-��:�Z��SJ�e�����$���zT��� V�v����X��Y����6+���$�kvg7���tR;���<��t�Ǥamɋoq-4��crOD!�*1 x������QL�F7�cמ�)w���n%J�=��Ê��!���/�x��p�P�3������P��&�?SR�狓��tN&�0��#%��#��І) �T�qF��2 ��ٿDU��M�8�+M��ߜX�(5?mCz��8�2�*X���~��OqU�ʇ�YF�c@��� �d`8��z�W�&�<uuw�#MB%q�vsؚ�dY]��1<���	(SQ��+�� +4�G:�>l�A�.�Z^%q�y��ivѻ�e�=���dff�.��%Np�����e�nhme ���WYd��������!�v�4�>=���~��D-���ê*��m5Y��uS��1����㯓T�5�D��3R
x�ޅ&h��s ީ�PiJ�K$�0�@�D�@�Re��s2]fqeE�ə��{ x2ي�䌡[8C��ѶՆ�ɡ~�":��"��Y?X�Yr�st�E�ᯈV�⣩���N�&�
��7{��,���CL�n��X��ΛE�"��噢��Ů�@ݛ��s���VKm^��6�8k�4��mW���;cΨ,���+����TH�I��QB�d�6�U]��� ���
�dc��
>���%-xDcp��"Ӧ˾N<οFx���4xq@��.+������R�^�47�K:`م�]ûI�l�=��c9���b�qIn��AE��3JI���n)P@��u�}���<B�U\���=$c�����%�������u��e�?������$�Р�v8;���	�/Ms ��N_�pF��P�� ���K��d��|Q�ݚ#���z=�y�΃�1`�
J���'�%���U�5�n*O�*e�����0��V��HH�U8���j�S#�b�ra�"�P��۽x�Jȉ�-u➥�e�)��w)3vF4�������y����``dKcE���C��s�+\O��v�r������f�Dx�q젠��[k��}Y�j �n�>��2�	Ȏu M9�-��fk�ݳ��.S@�mJ-�x��tgAR+�ܸ�1�!��Ʌ�LB�JW�D�G~�ٞ��f�%ٕ���@��(4��~�vh=	��~E���[�9굪k~a�(�1ꑶ�����g{%e�Rg\�5�f
hd�zӏ���j'��M�5!�
�;,S~Ŀ�d7x����GA�w��gѱ�=V�������% �fC=�:Da���Un�wc&���2^����;Q��X9LP)Ff=�d��Vo�(9nxj�!�L
lۨ�x��<����z`RSp���\������.Oe����n|�J��H:�l�0��sI�<!�?LƘ�f-�ƝA�u�#`Ž�P�V���$[(_e�����x=��'N��w��$���7��{�u���i乖(���=Y���t����o�T�1�������T��H�kp ��-��5�����v�SQ�pd	�ͳ��h�Z�p�&���^�s;��f������幔��@Ç���2?�:g�p��&�Q�p�J����6�����9���ҏ/���z���a;�Ti,s<q<d~��:y�Z����	�q� ��o��/���q��>�ڄ����qȊ);%���xa�ӏ�u�l�7]�a7��-�ԉvL(����լ��V��ߡ��t9f/��\'yix��g~�����]y��3�����R�Tj��r��s`!`.V�C�ĻD򋫾XI9�������y% 6���'%��؀N�V����z=�hԩ�l�8�1Z�����78���4(�R�ݼ����i�S�3�v���֟��SH�z�[%�C~34����t�_::���i��X�Q;��e\y
�1�7�7��ԍ���#���y��> 6ru]�?j
z���c�-�t��Od���#Z?��Q��~d��Ͱ�)گҺ��=j�qŤ�D��ܰ��!y(��3sM����k�M}�_�0vg�}����+�:)��w�P��kaaV�ި.�=]Yj�Z�[���W9U˵�b�K�Y�Ƃ���3ў������֊��老�>D%���Ȭ��Q��e���wͿ�����?�]cM�C�I�u���<{mB����rO�#�`���-�b�����ޒ̙�lh�i���^b7-!֓l��}z{����	��"EN��M�PَoX�8}��.��`��J>��>{Fa'�R%{D�ciz����Y�p���ws4]/���ܪfvؔ��_��~j�����yg;�����8�������	�wM_���hNQ;��~���8���W��4�ؽ�h(�9MZﺡD�����vǗO��T7�3����ݾ���	�G�:�L��J���~��3���ۊ��=k�6LI���x��ɋ(X���M(�]c(�����e
� &N��{+iweu<�L�XB���^��u����7��i�>��c-<T3߿S�񍢆{[�ѢZ�]�dzڎ��0|���+_�cf�}%W�MT8��)�~��$ʱR:����P���A���+&�"RQ��S �m�-��J����"�,cF�թV�=gXz�63�����;wQ��K߀j�k!?@ps�9fAn����2���t���Q�� �_��Oƙ��ԛˈ�W����	���̱�BԒ0�2\g�;��X淄lǇ�;��Xe¹_n��<[�C���.'�-O:�!d��d����.Moi/r&N!��f���l�K�ZC�2<�#_��o���i���wC<�PL�뗶�������І��BSo�bL���R#� 3#�Hp����!�v��Rϝ?3Q�5upy��ȫЊ��S��O�� ���P��MLnN�$���X�I�G��W�����k(���p�k����pH�W3%	0�p_�ƶ�X�}�y̙��R���3뺜.�J��4S�/ׅ�H^g��R�r�L�(���4���XG?�j�����e`37�f�\�d9��uނ1�B9�����֧�Z���URZ�d|�Ϯe�m 5�.�"�u�O����� ��J��{�[�����7�3���7��~+������`�ͺ�Ы�;���ù�'� �[}�H5�?_}�9]�ZN1I\���C �D���Q����q�� 13�'=9���) @췂�1GJ��������!�>�5��Ѿ�qG$"���bi@�LOLb<pf �)����Q���9��F8�	�GG�g}�Bp������b�������n]�9�y� Q�����Ƌ0��@.硅��XWP��7@�,)놂��b�,s������.�����x���.����!Lo�i��
7��"��:��a�w���9�i��(� RFW��F{��~���,�� �m�׼g�
��?#�)�GB�u��Y�%=���6M��w��ԏ Ս��C�e�g�ɬ+@}�D�4�t-��h	'>����]4�(���<����3��F32<1��eCK~�R�~�~J� O4�{�ѶA�8��ܺ���,���������^���Is`_A!�呏���������bz�k$�04\JFx�V��I�a���f8��3j��%��zΦ3�|�]��_n752��M��p���v��io%6����@Q���?�ՔnI���������1h/2�Nv��Ŀ�=���r����{��+�Bh��ǒxd]65��!��_�o\^�<5��m�!� I�l���0��[������2	�
h]�DS���6v��������ʣ�� �	j������D��!x*�s��o�<�������`���+��SLO%�?�A�Hg��_��f]>τ�.����R�#Z JZ$7���y�q���6�I���<(�/�'WS ���pf"��Y�+�h�<��-ц���f'ލb7;�Z�F���:�28��C,]E�NyE&̍eU��v�R%}2DBL� �&���1 dt!0��3����x�1NQ�w��T�}�����G%���"�����L6��hҙw<�W�?��`�%G엏a�oz�4@�@���Q2e!����=�<�am|VՕ�ͦ;���5���i�RZ~�!�Ԇr�]hc{U1u�,7��u��;Z\Q+�+ �,�\�@�:���"��2��1$���.�.�n�p��&�������K���%%��R�CݡX�\`O?���R�Hl�����+�+�,��"�v�4N5�~��5�� ��̾�T��Ν1סRI�a"� #&+�[kI�K���!.��B+ץq?>��!�#��(4=������U��#M?;�+*ya+)�$+p�81%���~�@���X�dvH}��B�Ne|�K�}<��P���J��g�%-�|_��i=��e�3�Y���~&���-S	�ò��r	�#����c�ɮ���x�
�3i~3w�z��y��Gʛ�L���ϣ`3�br�kG��E�o�D�b����I�!|�8ĝH�f����G�ɗ[%�{)�_@~�zYu��nH��K�p]���~Cc.e�@Hʣ���>�9h�+�Z��r-JN"X����Nc�4�ùFN��em鄮X�l��a։o�Fe�m6B<��V^Գ]��c|��ʲGpO���T���R݉�7~��@[��9O��fp,�I��g�U>.g\��X:i�&��om8��9���n,�6 ��h�{�ȟ11��������&�U�H�D2���,i��-�6�9�*A oZ��H�}"q	4�  ���7}��ֱ[��N�8�N 3in��#|�:��o]�,n3��sQ7͸���!���	s���l�]hs��i�q ��j��`��4VȤ�����!�ɬ���Ğ����g�j����#���%�+�^����!���{M���Ō�gWZ��ҿ&���������\,4�"v�aU��Dq^��͓ /�z+�<�fnI)Z�w�ѓ�A��
$����PZ(b�?�������~5�.g���s�ڮ'<�ht`ρ{�13�N��\��}'�|TSv�S��n���S���̓�7^N�3\������r߉��G��y�����b���p��o��,�^yӇ��p⺜�$�7P���^C�'�*�Ű‎�Y#�{uV�a���ߤ'��]��q*�D���7J	�9�p�����t�w����=kC�b7�`��)�f���n���}$��j'�����rH�Y:�P
9�;:�����v�oӦ�^�g�4�7�9ho��� �=F��ng��gs$zD�{ԛ��l�U'l�S]��[\�>���8�R�5�{����?��i��
z�:��n*w���i�����T�:�'�|1��EkQ^#���Y����+��F�i�@f�1L�k p�%�[�7A�0�f����������6��aB-蟳� �+�/���$��{o��'G5���]�>ƭ�i:�Ǒ�x���t�W"8�D%�߯�����lr�RRy_E(z�j����OY�vv�.R�-)�L �>�d[��Ɖ��3�����)4���Ϙ�8��� ]��#�w@/n��z���}r�.����i��/�?��R�F�͜�uhEX+�r��!�@,�.�{���9�����f;^@T�|�����I��,�D�A���ۣ����F��*O���L��K�����z��8S)�e��{�i��uct��d��K`<O�_�gR"�6�d��G�ο�����A>q^Z��Zg?gM���S�Ōu�:�U�d!�jv�4B6��,�ia}���k`t�%;!?��������IXc�:�_��C��/�pEph�S{	'K�������6���?�Lﾻ��;�y�⹍��mʁ�2��q��n'N��97�2�i�%o�O.7W�'GR�d�XA��N��y�e����ĳR�2�D�ӯd�!���k�l��~������cl'I�8H_8bq�:��±�G4�}^i҃�yL�Mw80�ĵ��)'�D S�)*��Ռ �l�t��GȐ���x��9�F0v]a��Q��D���,�>��>c5١��u���� �:��]�D6��}ݡ�6�5L���o�\nmU��6��x�s��ǆ��R����5�l��M�k�|�U�	��}K~q�f�H��{�k�L�����!G!̧ ٗ���#H�[�F4����ћ�%�����2����0��ÓJ�c&�ȭ���,�FڅB�9oG����F��i%����&�ğ��®@p��"�d�&�j��@�n!���$�Ya�~�L�-��:Yy�X��D��D�#�Г����&��1&u�K2*9�rŮ(f��y(�C(��h�x�ϰ��҇UF ��*ag��<�:S5��k��0���i��8[��W6�!�z�ʃ#�Ź}��m�7_�0~ 1�b�m�B,��/-��U���U��舖���&���Z��L"�Ā�@�[�\<uL�e�i��ϥ��|�s".��4����N�]�q�ғ���E��7);��^S9Ì6H��d�q�?r����>Π�Y=�
���ʙ�4]h���[��N̉V>�̪����mo���8)X9܏��э��	��Ԑ�3����4�|pJ��Y�?�Qe$��8��'�3Y축�ʩ�A���BEQ|]�k�,�-�aW)�0���@)�Hj����XA!O:?����t0ht���n�='�_���k��ʌN!��ݺ�)h�$(��� j�y�a�x��8~č���`���&A��x6�R����_u=E}��t8��=��=�핉����2��_?�)��o��1ߺ`�`v���֘���u����8�l�E9�M�xtA�ݜ��Q���5^Io�25�.w��)�ɦp.�S`WQ���G�@����K��ڶ��x����4�.<����r�/�@�=����	��s��&�-w��)6����0��Vlen�X���VY�q��l�@��wu��^-�3�6̓�BC���s�����c��Rm؀;���>��0mސ�h!�B1�E��?�v��t�Ἕ*Y���i�6�,����7B.�̭&^_W5���63wa&�iL�oIc�����}"��J�Mz7˼�!a��j� �lx��B�C�g��'���!�Ǧ�=p�S@?�g-�⣭�:�S���p�e�D�FbP��)n�p}��Vbt�j��Bi��d;/X�N�l1��s)����e��죝D�
��b�>GL��L���:�7�H��D�T�Bܹ�\���dǫO�����5?��	l&֋,�@���O����m���L��]��>�yhP=X�8���I���ޚ���v�Վ���?b��Q��YJ�>��cp�i��%�+W/�/�3������ �=��D��Z3R�v�.y�r���A)q�d�
��'����"�P�Yz$'i�*�H��&ϭ��$ �i�bs* ���%O��À��UI����3K<�чm�:�����qq5�U����x�.�Z{ңVB(qee7���$?Saݝt�r�`~��*��z�#���d��r��M��W9ѢC�'.�B(>����1�h����Z�+O���G�.�K��QQ~�?]�r�	PS�˷
>���j�j�F�J�F%�*��ү��N��"z>��h�/t/*���}�������3M���:V(ߨɶԼ"���6�W)��SK���]@T���d�}0�<l]��0Y��N�2��
u�2,ZY\l��A³O������ '-��t�U�Ƚ�іv���oj�co-�<�$�3o����fOy�0��wJ�^9Lr��[���:�D�,Z��	��C��Ǚw�F�S<m\C�xb���oB�����y�����ݪ�ȥ�Y�q<�2�Wf9Ʃ����B���9�XE�˄j1wV7��0͵�<̐��󙶑��� �>:�f���S)װ4=��[%r��y��:��U)���]|=����ԯ�o����-��7$ŷ�"�g����.e��A�l8b��;�gudZ�|�~ !V���d�4����Z�肧�fn�h���E�y���4�K�PN�����wZ����.`[�0�F� �kLd\�#Cz���B�ɡ
���T��˯����ĸ	��|@̜��� �:j*���kS��;1��؋��?~�	t�Gu��NQ�1�-Dւ4�E�~��Ƥ�Q~��:������O�x��Y��){���T����~�~J���<���MA?t{
+�Ա�y��ò`����u��Ǌ�7y��L�8O�(�צI�1��#C]�V&<�I)�"p��>��d�}=Է�x��$��C�L'yƀ�U,�����+�5
�E�z&�`U`Kc3�t�5��7�H��,nFoqI���QFZ�SM���&k��|$������G�Ca��wf�������%a���AS�]�����De+��e�_lp�����T =�rn���3$R��7Ir�%�P��ۡ���dZ�;��qG�b��(�/g�=��D{\X#Re�X�g.Q��ӫ(qo� �E�"�*a߰�M��0!_W��lk}. �����)خ�4���|�uֆAG����e]i�t�vxQ��Ġ8*a�|J�Ӥ��h�3����N-&��l)����0p'ӧ�O�'�L�T�d���W�k�\:�oE��Z��Ʊ(ٝ��c%�R��J4^��F���O?���.\	8����?p��`boIcBw��+�(�.a�%nOP����yb�~�#ptC�����w��IȘ�2�0f"�9�aD��P�E[�#AQ�)ϐ�P�f���N`��}"�f��JԹ��5/⫻��InI��R���Q^�z���M�����ZO�%�@Ũ�η$K��6�G�]O�g)�I�שVly�]���^Řmp�
�V7��gp@�N�'c�-�g��?�eG&0�&8s�5];�B����
�$��/爓��O���(�����C.�D�s	Bf3+q��޼��D�e�[��ߕ�J)��R�VM%[�w6�ZÔx�PY��{�=�~`��haR��:����^�`�~gd�ke�zgn�{� ���-��]LG;�!]3%��` 'U�L���#�f��/�SL�m.���Cӷ��g�A�ʭ�!�ln:��5�d	{�_UbD��
�M��O�͚�����?+>/O=�mRl�ZU!�
ڠu��|��mfD҅�?t��N�6��6��5z�ͧ*��O�����#��[tB���0�@�ϐ{ޓ?�F:?*�	�P=D ��;�_�އ����MI'�?|���D���罖�#f�|�{�Z�{T)�<נR`RylɷM��_Ѵ=�i<�CzT.p�-��*��\6�Y0�qG_Ȥ~!?n	���Ä��Z��f��K%JPiA����L�F�}<��0� ���|��l�E1sh��~w�mϯ���40�?��3��`�tٕ�����n�o7��wVP]ڻDhF V,��@��'|�Tɢ��M4�!y��	�d'�G�hpT�4��v�GR������8���k)q��m�#��oM�ay��&X�kJ&�f__��f< � �.���-�(�Kzk�Ap
�J�-�y�
?߶i���BU��rؿ��sD�,P��kc8I�
W!���� ��2�
�u Q�e��t�k$���	5�Ԧe"�̏I �	D�kn��m���s�'3���S�\�t4�����.! ����dL�X���i�ѯeS��U~V�>�jm�}��T��t����C�?�~���p�Z�����4[(OJ'h�zP���"]B����%�:2q�j�8#D:}��ҽH���ђ�x���'c@i��U��y���ͫ��֪����
qZ��I��ST��ȕ�eI�����A4�|)��"|v�#x��6����"M�4|�K~�y��k���E��e���m�����,:M4;7UqF����H�Šr��=�Ga�`s�8������ %+n�/����LاM�����v?�OAe�E��'�ǙQ�#o�jǓcI&����@I>h8%OԾ����O��J�6�K�`�������&8�ṳZ��.�~a��!=3�_�j�+��#�)db\�%�y���qR��]�޶#���(����<��[iսW�y�FP�����	�m���m�l��f���NM#�E+ʼ��[�q�J��iv�Ό��V�n�0�O��Q�O�Xa���l}�<�U�*3_E�юT]����(5("��k��)V2�S=c���'�v�?����dO�Ɗ�/m���X��d�8w
i��;Ui ߸�g��팪�E_��S�/����{�ޝ�a��4l� |U����=��A�w��i�0Fؠq�|P�H��ct���JP��-՞ T��!�P�>�,�b�ư��n��7�88Dl�i�����ˌyE�W0��$�������=Z�O�˙;�kӶ�H�%"m�Q��"���9�p�{�-k?DV����Wem%B0f��u�2�D��9u���|������eM�t'I�!�<
qZc>��<�L{���)K��f��9�ߪG[��SH��ԘW]Η���2�z�f�h>^D�����e��=	3n4�P�Tx�F�-~�����P�R�c�mἾ	%>U�VS4����#����^��z��~�{ʭ��Q��ؕ��"���V��8�
Z�]� ���Rxfl|L����,Sh����Pϒ�S��>�m�o�%]oTt�1j\���B�_�$:�f;Tß'�������sř�]���4��(AĢ�[�`
ʱ)a��3Qi��v���zA2˭}��I������5�v���mT��{��1l3�@>x�6�IYe���sk�7(G:�����I����f-��f�7�a
%�X����5�+nQ L��)�H�[�.�߿. �/���P�Mn�2�C�'���N���ˇ��T�tDeڗ��h'��-C�Y9}�7����&ХT㶥1%���&>һT���Z�^��vo�'���@����ag�3�
z�:�S�L���0y�}����C)*Ie�An��B�g�����BW&J�����vD�3sPK�k�T�z]B`\�ΰd�M|K<^��DK��7���=6�N�ZI�X$�^}T/���ɶ���L����*owZ(b�zr���!�)�[���Z�J�G����7�����'N�C!�h��][�H�W]M��]b`<Έ����	��JR'fc5��1�����p%X,�q�	��&��39ל��B�p�� �L�#����IcD	otѼ�+*q�Iv΅��T������$����θ���c�m|,5Bۜ�܄ph&<7��������/=��#���v�I�\D����!�󝙵:<�W���`,B�]�
M,<���[��_=4�b�[�b�:6�a,���-���\�	������G�2�8�������z���6ݪ߄�0\c\\^V�ӥ���7���l"��iZ��>�%����ɠ��sx��:�w�T�?��C����kҘ���k.��hS��e4"ŅQ]%�1'��@|����I�EͣvL�uf���[HtN��ri�T��2P��V6/'t�2�Q/�����㌈�]�Ǒ��_���?㓉��w��lń��2���Ż�m��g��ڝp*ep�C��T��8�V��p��"1�&����E�~����d���ο[xٟW���R��`S���r��g��d��*����Xj��9��~��Z&	?J�¹�/5&�� "���yh>%���V�mՇ�o� X6�v-�~D^��h�Q�i7��z��'RI2Cv#��Z:��T�v���x���U3ȣ�iCc_�`��8�2�^̧��߳�^�)%M��B�_�v�e��_wUn��f���?��y� �h�{�Q��a}/]�(����U׆���h`V����m>�O���e�Ɗ�tB��[:"����h/M�pѐ�3��`��:H���T�q�D:CZ�X=H8f�J{@\�+��߰dD�z�}f��L��(J����5�Ÿ2���$�:<pjQi�S⡧�#ŐG)��gZ�8ٱ��x8��q�/Gdɉ��Vz��C�j\��c�Z18�����݊K%o�?>V���ns������0�<�3�H���2�<v�^�9f�UG8�y찍[܄�y�൬GT�B0�����O�1�I�㗾��"�/js{�C�j�0�;oz$�ڌG�4zK�����1����ZR��b:T�E�|@����������kG�R�*W`���ŜZ��QH��Y�>�߻�M�l�y��$GwI�O�
<I�6`J��QSM%��{�Jq��Y�`ObW;&C�[(��ŮE����Ď�/�UH�Xcc`C��� f�3�����m�ƛ�������y�DzĘ�r��ڤZ�A>ғ/�@�ƴ�ܘ�VG���~V4���T���^����.,x���'Q�����1V�4����ӳGg,(@G �m(�䀜cao.6�K��b�g��t��U�	�ȁ��'�w���~�+@4��";|�p������_�=�8�l��P�ER�ތO	Ԗ�,�r�U<�i0�W�B�����{�Xb�ʵ��U�
�G#�1Js��	bË�����nz�c8L�oJv��y9@3�u����B�[l݊�ą\���Z�N��
���%��fL�m�)�<Z)�C�'��MŽ�uG����j��6�+w!�����x��*���H�uLF}���ZW��J�R���ƫ�S��1��!�"ډd]SJ-"fJ�X�~��#(Z�6Ϟ�!*��E�N¿%#�Ml�7v��^8��!���nC�h�n�_��$�B%�׳�B y�Е�ޗ���J����ΚR%`>D[ �F���^_�]&W�aXn8�-h�����ܜ�w�����@�/?y���.Q<�H~�2Fh
�����D�Mo�$D�ޖ�)��%��q"
����>2����Ń��$*�[:ʎ�A��!q�)s
-y=UKI,��%Ԫ͌9�����FW��_k�l�v����-� ��k�����M����$��g�mye���#zf��q��	��P���U䑶����v��`�x�
���=ir*(`@�,aL2�^C��'6)KE������KAۗ��}KA)���_��şx�U��s�\^��`�