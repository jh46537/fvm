��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7]�s��^TC#�yM�g,�%kڅHе6��&E��1�A� �uc��&"1��
�"&j�/�Ax�L r��=r4(l٘�uL�}�B���?H�ҝth����5�Ә�FØ���\�V������]��Y���'��\�;�j��P [D�m݉�Q��凟j�1�� ^�������0�¶��X�֜SM';O���+�d?2鵄��]L��>+�ee*�������RM̷LY�L;Aj�p����Wey�S��eO!#�;���q,��f��وS:������0Y�1���w������0tBgL̣��g�^5aI��GA�-��i@E�%�����Q(>��ah���#�B+�˛� `-@lS+GnuEO��oPQ�/��^o0n >��M�r�~�%]�f�7Cb,����g����Q���r�{������)��-h��{��WI���R!k�3i}��wµ@��lĂa�bӰ�CAk�ll;RI��fU\JX�a�K�dI�	-c�a`�x�$C�k��w��i��|B�}ا]~�(�K�,��3^� �ݨ��%R��W[���w��7��;)�-��v*�Nh�(��)̶����a�`�x_�C�� ����Z����4��4��'���w=LH�U��7�)r,�H�?[�Cfk)�:k�л�J�cđ�ɨ?��;[���s����_ORJY�J�!{tb��]�R�l�ųCy�AQ�x���^a��7o�ce^�wq$�Ʉv��oʳ(����8 5�.u�)��g��%c��;�Sp���n䬫�&�ѷ����+��s���bzA�4u�}�^mp�H8��o��P��ۚ�%�zk��,����*�N�� H�c���M���x�ENv���wto�k~j���^I��9�?�����t�|�)�W��E���W��lM99��Χ�kN`aeLp4���cI����BZ���}; s�Fb4�a�q !͡'#�)�m�Q:M�eS�M��>B��P*�!Lc�-��*�?�^�Y
��ږO.B�{�s�T�ʢ<��`�vۊ�p��Aa��̋�!�����NG݀�o���O1�� ���J��}XIa�Z8��wGb���f�g~@���9�f|��Cwp�Zq������;_�!�p��wz���Ufe��g�1d� [A�D�T�f_VQ�v�Y�
r�0$k��q΃�-�mb�Xm
o�c�����#|��j� �.T5�f儒ݶ�&���]��@��-�Q�;�4�������~2����"E������t֡P��Y�`�7D��9ة�p*�� X7�LovVPޒNK�m��y0�ԥ�Y����E����3wY�YX�phBl� ��=Fj��^1�Ѻ��5DWQ��7�bF����(Ś���b��P����Q���s���v�b�e�xVUù'��ġ��}�����J�P�i�=q��Wز�D؛�̦���^[>y'��u�`�J�>�o�&	��bt��K�`$��s��߽�A��Y	B��L�B�M���{�Q#r�21���t5�d/�!;�,�iG���,��')��	lA�=k���O@Yy�J��%��D4�>��W,��[�q�+�]1&��.π�ۼ�<�L͖aݯ��ti�������Lh��K�bѣ��9J���N�A��V�j'�-͈qj܌T�:$	��{A�f��V����*]�K���Dgd���HM��l�y[�R��t��^��{���p����yL��cZ���f�d�O2��e^�n�	��iguܪ!��`�I��D.�J��,�i�[V�7�r���?��Mŵ����������d�����S�Z�muYG{p�*��VaЋ��w[��N��Ws����nش.hK���K&�8/ܗ)�6��]>G�>��0�w�����<ջ���<5,�?B�ZQ��q�ѣ����h�zA�.n�\d�?\��_�k��ب8^c�F!H��d/v�j6|p-�9�೧)�z��,�I�}5U��O��D<X��^�c;�k"�H ���̮l�����Ě>���ĸ;<��#n�u��e����km\x���4~����E������x��&-�p�>4Eס����|\\y,�zZQ�tpf]�{��G����|�b2-�;��,�"305F)���W΋,a5$-O<W/�5���]�77��-��K����]�rAV���SW�
�����u�nwz���wDl���e�����������w1}���G��.%?�;�xVDs����J�:�Ah��jwň�WL��Ʊ�pF���*�;E�N�pٲ_7���کD������`z�o�_����[����h�>�ݴ���s�e�2��Mc�[.}ջ[�3j���i�ezp1�a��<�k{vB$}�P"2��n�t!,���p�zz0�����)>%iQ�Tr�oγn�c.�4��L�	hE3/�o�H�[������e�6/��Z�y���0�,�td�ڲ�s�� f���aG^���U���>�g���qY5rMYҒ�a&K�\��xt�����Mg9�<�m�) wa�vD���C��gL� ��$�ߢ��(`�����IrB�6��/۟��l�M6��������NQ�$�:�}��w���8�]�w����]�l[���P�;C|}����ޙ�*�	B)զ�۸By�V�D�W��A��C�F��/w6�d�;�<�����ФD��OZ_�z\����'ur	ͧ��C�0W����d���(^e[��򻷘�cl�fMbMq��Nłɵ�N�Z(@�/�B���:�\�?���{��]��)lAh'��kO���Ü`e�{����^�[�;�tfp��pب��׽����q{�dy�^>2L�Z4�������;��}m�	���X��x��<^1��'B�o-�'N�F0�̨���Zl�[\����&D������T�"!��-��n�������pp�!�"� =��f�4��>iĭ�^�Ά�U�a	<�r��]罈�Āլ_�~;�Y��nB㑕a�[S����{��G�yf�B �)�q����yy��<��r�cZ�/���54u��!�A|�Fl @���1�=�����?�b$?(�Wᚢ���a��&�����	�%�Tt��l�sh�m\�	�Y�P���U���)!e(������Xh~F���×R��o����X�22jM#�Eb�T�)���ų�� �n8�>�UIƮ�%�O=�� �ٱ�KN�3��:(�C�\+Nt��e�V���O�^�A�b$v��Ĭ>�n�^�v��l�>O3�.��;Ee�� ��G�^;�Q��`s���=�N��٩��
Â���%��:S�0�;\���ђ'���f@w�D�:?K)H���
��|Dn�j��dr<�wpo����~�~S��|M�ᚤs
ڌ�M@G�6dq�3��2�&^x�=�N�}�Z8.�jNaR����@�w�@�mw�� Db�}`��&C�RրN��(0\�82���q�@�xq��y���q6E��z���T��~1U��l(�
,��oƄ��Z~��²���c�3�AZ�9�R<��N���PZ� D�`҂�����6�lS���%��`%�
�5b�&�n�B�nL����>�%�7��j�^S?�r��L�B^�+����v]�� ,�}��;��Ҙ]���`>O��K��S���+q�fO~�0�f���ن�3�S���8���v�D�T*�/&.!_���XIe�=����ك�3�� Z���.ȉ�d����v;��\\��Mx�]H���d��1KV�`�7��?���~V�J�[<
N�T�~�T�J�
ۻ
	��rE[2�c����j侨3��F���`���&'�M!Ag���1�\ypx���w7+��p����*�����ZT7G�tw��-��t��>䨺�I?��WJU)\��}`������=6X�K�E�{r�K�|��[��3xI�ĂG�-���?e��K�f=��Ԁ 8%>8���j[h���,L�|��k���_�]޵�\���и����J=b���-K�Z�����IW��ᔂ���p�yI��K/�m��l z�#U9䰞�P$RaISp:�!�Z=v��mvc��I��.7��艂�\����ba_�V ��E��Zk���tu j�"�����],B$.�$7���)���:�)�&�nZC>VlЪ�S��˨�PpJǵu|�b��0h;��L�2�2�9�GM���<�t�Y���A���7ΰ2��d.o;8{�Gvh8@!�j�{���i�Z�C�q,4	��$}���n��uy 5ԧ����6ȫ�O�ܯ����&zX����2b��d��v(Y�h���_a|�[,��0�u#�Ť�����L�²���J]v��hP�����k��٫J8_�����+�Y�M#�c�\To"ai )]lŰ��l�r@-�:�/CE�@�����9'ٜ��'z�������� ��=��6,~���.�������i��:��Ve9�Qv}
]Q
4yUE��.H�ay.��^;"�B����15/F)�~@'�mF�b���;|�N�=�����k�R����A���l6�w�d���e��ݗ��E�ev(C��dܲq�i�܆�i�Z�S��"���ȟ�^�B�ߋ����';�vJE��0�p���>EI+1�ׇ��0�"Q� |e��,I:��m"M{����{���q!�:	@�X�RuRw&�b.���T�/ˆ�LF����,�vgB��!�Ĩ8@䈽�%��;�\��u{b�W��w������(�
�Wd!죋��k<S�h�	��J������_��<߆(�8�=L�ر@^����s%����\M&�O�F�|Z04U���7��nX���-u��ˀIC-*A�;�	+��E��1��z�-=$..�Y_��R2���}�n�+06���r�"V0O��"\_��ʬf���#CT�E'"c)�p׎��{�=pD���V��Ёd�.�Ν]W�fQ�a ���ɼ|�2�uE��w�b<w/tuf	��&V͸w��E�k�0>5 M�eջ��	F��Ҭn���v���D��9�^F��(�x�;yIztK-���=/�|��'��,Evq��n0�Z��C�hΫ���j�^E��,��Ж�J���K�"�t0^����} ��4�n��cwjm	W���6�еYo[Ò;�6�۟}s>��iSŉL�J: