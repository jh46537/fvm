��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK�Q���L�OX]B�Ј���}DO���!"$
0���l�Zy�@�Q�䎁�1�;7gF�%}�����Z���MI'l|&��Vߪ�^\�Q��EsGF��	�M�|��Ӗ���'��T5^�] ��S�3����':���gm���k�R�Fo�m����>S���xvS����#��T;"�4���ů���]�٭<?��߃������O�!k�^ �B-4�u+�S;w��4@-Ra�Ӊ�D� ��'Fj[@*1Sֶ�{b =�S豮z-�G\����#rAn�G��Z�W~��q��m�#��	X%�߳>~W�c5��v�ǋj��\����Fi��;��{�ԁ��,>?�g/�0V:R�E�nO��ƅ�gg��)P,�ر<��A�����8'�=��P�.l����s��.��!��]?��������OD����G<�Hpk#���ժ�Y�;޽� �����v���A4^;��=U�g}k��N�+K��]��U7@�ק �W���{��"Z^� ޹"Ԙ ���N�L�me�7>���hw)��7�2�Q�����>�m6�=���eg���k8>�ć�N`sѭ�zpe*l�2PL ��|rs�&-.'2@�MNdv���;.P������A�!�*���W��E�>�,��W󴉶㯔��iw�K�5���ӑO�iH�4�ԃe1Wڸ]a���9��U%3n?{�����M�L�b�~���L��
��"ڪ�����u!
ϿMx�S���-�sB�BA��Eԭ��
��x6�f���s��[GjL��N5��6N������1[�j���P-�3����7�0�!Jk0<��ez]p\�]	�w=^$���	��<�iy�o|��)�=]}^C�����z�i����HLU��&痯�c	���q�H7�J$Ԧ;��%zI:� Xa��TƗ��	�k��x�������
 ��� }I���ϔ�]�;�̏V�!��{L�����3<�����]���.�xǑ_%x��¾i�鎗�e��rCCu��;X7�Z���p��p�t�	=��uH�|��q�
�2�%F�/Rƫ�ktSr0SuN zg��⽓��c*��k�f��{A���дe��#�/J��s2D{+��=��A�K~g�(s`�6�s�߯M*/<�Ua���,b������	pd9���c4���z��U�+|�2E�/	�D�cN�����qxUV
�����q*�����|DG�ZDZb�{�R���#�Ǉ@\�h������2�wob�Qe� {��U�+Ϥ?�畸�?v����^j\ɕ4,&������X֝'z�zl�/��E�"LCp'ܴ1cn�:W�E������37�������"�Ķ���߀��c���/d��m;���R����1�//;�b*1%c^���o�c3�Hm����X1
H�Z��%1^^��c�F;���l*
�w��/�*D����;��5UF�.l����"��!A��ݢTz��k�k�q�����^���{���.��J<aͧ[�!���8���Z-"{#Y7��1�-EM+ ���CZ+�L_o4Pa��X�bîr��uU�N����*�3�f=@�}�-��� Q��mF����/�&��D$귱hZ=���*D#�>)���b!CR����]!�zYb��l�壅��}zÔnY齍�g��'d��n`����p�YB��3>����Zz&v���=�'�N����-@�L\���U����O�ή���6�ɻ��64�!I�e`�	}L0�͞�8�$r����|�#E�45��SM%X��&[f����[V�̌V����扝R�1n���W�P��ruR}T�4�o���;!qɍӐzzm`�GE}`qE��r<R�zFmb��σ�0Q�Ͷz���$�w-1zJ4�����a� 
h#��̨�+s�%�E��s�����&͹$�bK���S
�Ys���g��v� ���F�X�?�hߎ$JV���rt����(:m"��s<����:X�*�l^4j�{[D���ҟ0�>]��GNzSK�fK\�o��n^Ʈ�%��n�j�<2"���~a�,�37�e9F2���Q������or��5�ˎI0����v"	��t(w� v�!��n��6,\'(E��/*�4�qp�����.���b�9h8��_�:&��|�������w�ea�K�INlб��T��EP�����&�ɴ5�?m0M�Խo�������JĨl�g܂F
r�㺰��V���9hIAl).pc10�D�w8;Ⴧp,���9U��"�)�ߤK�ɡ�*�7nH�<B�$,O�:��Mo%1��+A�-f,v���*���B~�iz�Y�:a\5k��@`x�-���L	�(H����56���Bp?-��!,���ݩ��M֦96��1��r-��r�Bz��Iy��c���slY�Dr�3��T�⮱��f}�-\M��LZen�?���A8���Kxv��Ⱥ�wɒO�d֥q�P�a���y|t,?�u�5�Z���]���+�y",p������M��{:�L$(֥��o;��x��TӇ6<�z��1bL>���ۖsMʫ�7��o�	ST��cj	�2ce�6&`uΡ{�R��3h(���^CT��LU�d���d���H��P'�4�Z��l�8����cw�Fи�J��0O�tM�f��&���
�'��y��Jb��\�\�^���n��fD�H��� $r��[�/dhzh���dԲ���E ρsA���>���E0E�V� ��y��s��D�m�1�mڟ장I��^̒�^��H��ܚjL|z,�4Ԋ"�cMUpX�m�Q@����R�Z���|��I�
��4�@���r$k,�-���z�6��J*�	脸ۺ�E�NME�\�ؼ`�f�q:wI���-��(4�/�Ȝu x0"I����9�z�vVG�f6���GX	�X��q�b���0Cf4��L;p���ve��gGb���X&�7�=����`��z2�P��6�����I�ͭ�"7�v3Ƣ����8�X{ң7������������L�q�@8�����h|O~i���F5����Q���7Z�#{������ ��X��N���>�K5T���)ǩ� �՛�^��Y���������p��* �zr�Q�\1,��X_B��? �ʆ�ક��/�[!�Z�K�A�����,"B�%���s�=�>@팻 �	���岱��W�v�p��O2�x�6��j����q�9�Bl��{��U��t�l\饤�'x�E�hB�Y�"c���fP�gs+m�v4�uK7W�d�nV��fA�J\���V�x=Bk��z�	٠&
_K�H����¥���;Nɐ��#���^+
߬A���ID(��}H�������z椩$�8��8S>�\4,G����p��Ӱ�{Wu`�=1�����a0"�������H9>�{���P�V}� ��XR),]n��Z���M�m�΁�KY4R�~�g�u�	�VQS]1z�B+[	����.B7��?�ޝ��8�*kC�ՉkC�UrKU)�[�b��?���n���Q|�r[������o"�3��"4dö3��p���*��|��ɗ+#�����*$}k�xT��K�"z��3��b�P�	�{i�:�=}�TU5RJH�a��Z�t�}��x}\	���_����6#�߸����P�-��N���'L�����K˩ZQ��m�������%��*v)>;=���V�t[�}�L��U�Z�\�FZ���,�u#W�z�d��Su�Es�5S` ��ZJ��5�R[3��t�h��ۮ5�[��y�qXs?�#���|�[��8D��O�!��ڳ��>r`[w]z�þ�G�0�_]L��b�',O�R9s���R���}��aL8`k8��{�u���ބWۣ]R��A�-]�b<SP�k5{�KZ	�/?�k�n����S�6���}i8'I��ɦ�ъ�#fd%&!lU*�Y�����s��Hsh��ʻ��@֧������I?:\=��4@�'����@������@��O>z��+���5x���pږ���e��mY��䅰gn��^�����(�`r�s��nzn%�*an�p]c���Bj��s@{�Ñ�(FUw]I�Z]���@݉юk&�&A��W������L���R���Ƶ/lƈc�KΗ�������wi���}RS�~��30���ȐMZ+��\�17k�S8[���������.�}C_��2$/2�6O@]�7`x0?7�Ҙ+���F�֨���xYp���D��Y�����^�yO�
�9�����Է2�("H[�>�4i�{?�,�����q�{1�38�F0�Z�X0-����r�۷�%fň�����w�*n�C�O��@x�ߝ���'%�u��l9V�`h�!���}��%Hq�v"������V�l�����7���	.���kuY��
����w��8
�z���$4����x�����(�1P~�q3ޝ�$��*�C� ����N�'�9H�e�W�X`֬!�RD�{F����&?&Ϣ�^��<gr�2�u�fY!��%v�a�Z�O����Z4�{����ܕ�������uA]��x��ր���;�r?�6��\ek.���˝��w�N�eI��Po+|X_���<t}#��)�|��G�T��YN�8�U:���`�<��Yu6�15�㶱�/�ʗ�m���~|#
-$�Ԏ{e�H()��_f0�� ��
��8���5m�Y�煄�jAk�J�W#&�?F����Y�ٴ�i�$��#�?�|�yY��Af1Lgh�3��~4��&.��5� lJ��K�}%�����e����L�k_f��nFM(�
1]s}�H�v�M�ʽ臽'\s�dw�NF�Gfk`�tցl�5uJ6)z���&_�c,���:���3�7���B(EM�(�6������%�����(�����g�e��#��P$iF`0���0~0�`p�D$�	��6��G��<�/h��6��I�%G��y�������e�;h���K;��_F{�����}���n��[�&	�B��a �	���t�8j����5]@�E�||	���a4ga\�k��q$����K�lƀ�+��Ŧ�*/;��9y+��B��`.�ehM���;(K���w,F7�٩׸Md�\���K� �� ���صCxwg��E��zKy�z�%s��h��1��HgU9ؐ�n/q��9�Bw�X%!U~C��
*���&�ˑ�f!+d����jg�V<�s�!���Gk�\|$1wҋ/�$��`V��J��;�0��#Y!�3F�:Sպ�[)IgK���у��܂i3A@� �+��>9��I�()h<D���nt��:Ô z1< ��b�����)W�+�}\�h;�X�F��X�����`���P����u�s-&c�b���U��,�'�ݠ�鯢l�$Q&%sG���fc���^h����~+��a���p���xv�������kG���ʻ�3E���5��Ǥ�OZ��F&y"�eNi�/ߔ������8tXo0���)�)j�yq�߬J��6�S�v1բ��D�q�C�xN���6��qC�,i��m�?,�w�-9��f���ǰEOR��J���E<�R[9'��HLJ�C��h_ЁcPwN�E`�[h�S�r����`TBeU�à��XF��hj�_��$���5��@�~��7r��;X���.��Jr�I��H4��%�/W��-��y"�����gr&ܙ���M:�=S�L�2c��G�UƩ���4�U
aMGv��|U܁�<ш)=�����ԇ#��\d�����g��d\�ȴe�Y����NeoJ�K΍'U���JS�#