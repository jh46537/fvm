// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k5heBrY6jXe3/GqXFHefSZmaEEGKziCUUu1efYb5c0WJN0yoQF8pk4pVmkUQk4Cg
OQUfA7fHxrl7Ro1rLh/vGZ7dxh3R8pYnK9SQhTujUvaKa98T2+P0Kl8Ku8UN6wrQ
mbqpDvIkc7CVUjujrG3AJ0AJcgMYSbYdiVJj7zR2t+Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 93456)
TfSBrB7OMRxrHFFflSHncDBoI1DIs97t/hLtUx9PKtweSDa7TSRQMRv88hHcfgCF
f9el9zvI6ZvtOu1zu4uslQzxiXd77XmUXzmCnKoTqj0pEFPFdjdLgu69uf8ZJKkH
cAd3VXQwZKie/eckC2gQ2ThQ30Hl38/GsElfU7X5oVFGBuBDPyyQTSJ1LBE87BFZ
3+gLoTWBzRDkopcP27ooC7Ps9hbmgKCbsmgbfnqCTZxfhJ9/sGRnZ9piqZoU1MUm
E1rTInJ8jlo54PbmubK6dHTuL1x0gIoNnpSoWvCu/UlJvczV0PkqoKJOGFIFmiQ8
YulVM4f9AGboCP4vPxLAupKhTfi5yimVaOp9oIIeZqzHLA1hLJ50WEmNvHVxuzsu
5+QWpsXnAB1VwbpoupbU2bIEM03JXBRfnAefddzya2m5/idbaJ09Sc8qy1v/YxRg
mGC3YBBMFKXQ5WEJPk+EjuPi132S+YifsUvf8hxE/5CEzc+8It43DZnJQrIADZMm
xiWM2xpMyR2gu+jrKLWLmrmBWLTNVbHNUDdRt67pVasaewXT2tjHXVpai38nTQ6X
jTT5zycZCvS2kbn1Nh7ei5WUxr1aiclEql3ZmfF3FK5C/lbFyHnWSgv2/Vj7pU4V
TxnspEgtlb8Ik30rGADCFv6D6s5bDy21QkCAR6ZV+5u3zutaQXH2R8daYnOBAlA1
WSY0JsxFWQtAo+heIjn03RcA9ZWT8cCDw+f8CU68YqRWJzEXBk3rkz9JfP95B8OK
gtWJAQAk8WtmndJGgZQJUfqHyVrI7ZmgPlds8G/i1kksrXzUxttHoh9QqB0JJG7/
u9aPba6+TLRStc21trxwmuyMashaTw9oDHqKJI5KHGDf+5BTrQK34KYSVnvc+NmC
wxXmIsatnQlJlQKhFSMlM+29WamSiFxkzRYpbKxAKLSPEy0H8tIO+8cqVY4IOZ95
i4p5TWzi965SUXQCBY1nSbeh11b5MOERYIR/1WDL/lSyov7PCLOURk3+3ENZSFtM
2SHaXeeAZx/V6uPPsTU0+e7Ws1MShKjUa3eTF5G0i5mob+d/SwZ0vKeiBhPkCCGY
bcZKuLW+xQzCuVgLtWEFLKDNbLkpQqyU82x1f2wYXmr7yQZ4dT7ls+jNIpGb+RiN
yD5DbQqKuo0VRngfAD5fSRKmZXZ88blRR+wZ7UYfGfR0aM7N2aXEWNYzm6vdaeid
VkwCDh7ve+MGiKSo1VRJ1BAwEm/sQDDLx5PosuGBCZkAV0pe/tEZf8kJ2D9Xlh6J
Bj2pPGDjYMob4VfnGhAO7XLpWDCysjOCj43fmgJk2xzQ0itcNNuOdsgaTte9SAvN
JUwGhMiVbcJ+ZdvpPj/LtP8n2/MOjfucYylqRHVIOBb2XVDCDr+b3uHBi5u00v92
p1s0nMzA/FrAjs12kxN4TGLNLiPxFoopCffLD1/taEnKlxYHqv5Ay0rTxoxdQ3T9
nYTg648SUP5VE7NmhK7UMAGj/17katd2+nA/FklHnUrJQjBP0mSFOy6OD936Z9qg
WnKdYriGu4Q+EeHKB4VfsW0BYE0JzL830kfLR+Hfh2Y8wC6pnPCjcBAMDlZmHTvr
ORyp2BCbu1crswFJ4PYjar9BeCqso4OLU4YUjXSgabPxHiKDPcLBLRbWr+Lj9ig+
1vXATVH1J7dvv58wHBxwih1mIXYfiMvoq/j1KO/Xg6E70ZPjOy0XYArTKCcfCPkY
vYyu1Oa1ycXsMnGatn84iA1hlLcC0356Qm7CzPmdoAGRJ2TfOuti7umqNLt9IaGf
ghet1ebzw30iA62cii3SHtzVLychEByf/85zoscTv08cELAlB8jksB88HbmwULTx
FvxcKpykGkL4DrsbYv183MrIsQ5TAEXyJcZTjDfgEINNWVrA6vpNnfk4K9p3nAZG
WOdpCATb4Gyswdx/AiuHKX1osusH7zkrVRGV5+xt6clfRmytx42oDIZ7TwFMhWnJ
VsWm1PhW5jbYLsdGeqTPBVJ6WZoPx1tuLWi1ATUryNSXGRnX8Ghakyyz1YyehXyG
zNe4xLm0x7Nvkw0kUUzWep0MNSEOrxXWj6rs/mBFYaCFvsjgHsfBSdmKMiXVFG+d
cmDw7sBydArrqhqIorJpuveBz1vwpTqw5V/AxUi7DqHSEcrSgLk8Ff+yvO8dbaAQ
pf7x2CXOUPNxuTtP8GFmJHMGPAPYPEJoIyaWB76ZpPAxFoSwvTbZK9c60weAe6OV
fT237Vb+wXEzZmtHw+030Bzhow4LBNVuccDYSWPez/LX01POnYjLRnXMIzz6kHrP
G4Oz+jHPpACx0qCVHEJDkmjVjA6UJtbBwDAEHSCaRrLf/6vEFNJmbp7KjixfjliW
Kn2wsFdKMqCz/do3rLzj7yVU+OU1eTgDU73FLzfAoRvllHqt9JYEBFPymyO25ZzB
XmvHB5m+EoWp89u08N4m81AtoTzBA3bS9ygdL93yLn3P9xaW0KW9jHmzKuCn6sCt
6xH79Pxzb7EDUlXY0LxVmjrfq1JQvjRQGM4ca91DJT4BpSYRSq4ClThnMjl10eN3
GyioYfTguQHTYc3kM+TacgP/5nhZVsMwoyQugYSSPPKSa5CWhiaYdSKilBAy1V6H
qmJqZqT0AfQVlF91nEpU/02pPiYShCBnjbQegFUs7o5X2bxvwsx7U/axO0Aqh4sn
pm/E2FMI9ZgaIm0htfpAbnYO/gIoc709NE1oiPOovFXKkqPPjGQaii1J2k3MkSOW
yNjCyf3KYw9zQr5ic4gmHnk5JGAVvPJ0iZWQCdIZWKVqO6IjnyB8v6ecErDfBmFB
HWaIOWvLVRprJ/EZp1JYGOsaEBC/gIaQJ9ZmrizGR8rDSkrApLQnRFT5lPrJSJyu
tQF7mhWmynE+GiNjsTTjwv9CxSozWHHx7RatfKbKoWtkiWQ77Cu3JBtW+ee09HFv
tCYiAlqs44tdFVcNvSaQm2nnuP+LTqx2fF86OOtk1+PSJIAl/EiZWHnR0mqkDBhm
JT63Cun3j/+zrvzZWaXsrPAUnVLLKuOOqK10mlZJ73PVr1r0ZvVNiaB/zh70izDm
1i3xLFGzuayKINVcOlJflAc8pkqmhFPmswwJeJiql2KHipNwVyFAtlyN+yhvu+4L
zw4Q5aVi4arWLapzKqzwyR21YxwvhMTJ+xT+iWNUT0IZ/UsjdpTsvg6JPf1V3Hrn
qt4Ne17wCIJlg5Okep+SBJ8+/s+ZzNmwvCRcwf3AjLjH2oWbR3+zGLSHem8QHL3w
YoSYy6yWwMnziQNP94/qM8tfDDv5mJzdJfYVJmFw6P+lfOyE0gMwDtM9iAuN0gLu
aqSM7ZTqHpIq6l0jTy+FJbw24pjX9SbzluzSDG/FjeHIWQrl2Om5cQDJb6kGp3S5
t9V6lFHko97gBMH4lOkUBTXyWzw/GZfGLhZXjoeVWjFWl39RTbm7kBhr9C6SE8Re
jFwB+uvyh59boJhlfQ1UOHmNSF6Z911kTrcxF9ZZLWXKk5gLRGoX4CATJ0X4lkrc
13HeHZXmH/2KEh0XA8WyX9DaGIirBa7a8/MkPyY7+VmZrT/DvtOg9z7EqctbSZFe
38KNhLPb4tut3OTDSJap3Uoc5Ub1XavSA2Y8ASMwIaNjCT16hu9/CYQk8LlwE52z
C+mohr4U+9B9NWDko7pZVrvkSBy1iAGJvrpSx3e1yGyB6zjaNPw6sPaU0bT7GVUY
30AM9FgfHq7XhIpslnbiRo2870+BH7a/VmYZhxmga+bI0XAy0iTovnk02YhctlLg
I+nHbJtinqLKjLJZiLrCADOOAHLeskqz9tFANsWLAYEg234nxKJHHl7Mf+uX8O/F
KAbGBln6IRocROID7m3hhHR2kSnGM9E6mUpQFpZPzmo0hJ80OhG6nBDrOzIUsfFY
3CUySTI5OOWj0MaOdb6GePghIRBqg5BKIFZC3PzzlbnExQV7cyAOsebCAOwwVHJO
3U9Fh6RkSFtjdRZMaWlEbcUOCFX2gHXiknlJWitKhxSBnobaLNmE1i/K4WqpUd4h
h2sOR9qbXdgYIOjjZLgYHsMaWi12MQGemgSNBvhGJ0LIk6AS3gcdi4fZullsIhW4
7J9nMfActkjDTmoKtCS+ks1T55O6bInXPO3xZqHiO/mJunInIoIenKPQ45WbrzcO
SVnVBNKyDCeO0TJh0IfIYRyODpbQmMTrsM+OlZCEsK5t+LP7JhSYnkcxVXCIpVuB
cs6thsK3hgEZS2GfWwBX952Jwk73/5Ok5nqn30/GZJkuSjBiFsBIKhjWw5dWm12U
cUV9y9C4EbW35fZK3g32BHJ0fDZc1GNAB/rxuD2U/ze2QOnJ5q9TUr3zSd2n45qV
zeNe1+L7JGUI+Iqgk8wnKF4rf6s1OX5ZD/8p3SM6uHISenPPy2+awokUOzGLGR1I
A/w1vWEUMzgQVSuUrBkukE2E4u8NaC82O8UYwLf5K3rRwp0ZA1SilnqIy5l/l0cZ
gSJopI9dsaeGlzfc7MbUbpqHeZ+vUj40fiT4VB2Qz7Bzen3o0QsCCiR8qmMevAVS
Xq75Nsqe3f5xdzXJ1hnw6MeLR/oq8jkGGUGgMahMph/rofwSdiJT1SuvoNKH01yO
xGMbEpn1XUbfFbrC8qKj+jWFj21/VlDWOcATyl2mGtp9PXXVNMKi0c7gh6DrDUYp
hIZbU1uOIuGREmk8AyHLZv5I9renaouqo8tV0LEMUTJUCpL+qx+upwOkrtLaRfx8
vjc+Zn9WvwMOBBafTlZwYxiANNkIe/M41M9zLNHsJ6SYHhRRcru07V6CE97s1Jw4
Jawkm+MvyeLTUttU4jHQ5KpnmAyxfQeN645/GiZhr/O+Lsw4jMgZhnymMTK2b6Wq
8LX5PoYeNCAlc6UGaHmZ2crFnPgdBq9KBj5I0YEP1fClNXquBX5cYzxS7yOTp8C+
yQ4nkb2dTTSsfzKPdOov0SRsrnHD+joYM4ueunCI12Wq/MZgcN0Q6ORr7+1Q1HXX
RUWySvm6+gPm3XdRiPLkIPrfr5B/xGDoVaGJmCflc9lEVILnMNOOopsIPWz6jp53
ME57eS4Aq7De30Ym1RJCpT/CoxFfqPZC0kySALYbIarjUc15NaWaUAgjUZTltpOc
ayYVpZQCLfocKALUWnQdUAMYFuorfJlUaLgm5aFBlLlaVYY+zlx5RKD9pId2y9Kw
Yrwgxfin/AZNT1K0+DqtkZXtvV7UZbMCgMVHVCT3+QBbzeRbwEN0xUxDgh/bqOsW
kdk2YjF8UqRd5ouIvJbkFULT0+XOW2paYtkGM9+4kkLvUs2/apRF3TbIui8/jN9u
Nui0IMQ6eX8n2WT/j4+r2kkTad43sqbjEimH+u55OikzmxxJQYZTLYGH31tmaLZK
ZHktIY/OPPHPOORE43ArP6DrA3Q08Ypj+NWyQTPMh1BlbH0sHuIIRH4rc+SkQcOC
VHTB291eiXflRYVI/3Ea2c+ctLaIzHc+xldZARKIKuBaro9e/g8JGC7VimsYGQHc
Jd3I8Kxd/+2XGm/hgRpRYb1rQEyISqah/we8r/o6H7qmPqHoQjJfq/0Mpmhp57qB
Ua+yMsios1SnS2VUeVjFtDDAmurJA6xc/3E2BRqtrQsAgQnabJNRHfV7irhwafcK
JOVoLfOOI8szmbDuFqf/Lr4m5OewYk3FFKu5VFQWOo4ev8NaTjt/iTIf04zzFa6v
z8OiEok81k+OsflaEuE0kLTRyIQu+P40TXG2FDnMgiu0bbgSfutzUpsZ60O+tnAA
FuF70gofvcu54+vEpghwW2fW7prZ/sBxUDLu/YOmFCOkwE9EeaOXRpxikgcbKvek
DimzGs0a3eiyTORmnVoNpfWYEqPi2m6qqnCpl+MKeoyRLmWCr7eiuz2Zibcou1JQ
6zOh8uViep4P9iF1YlQHCnJRwiXF/48kWU4FI6Gf/2niW8BuqH+Se1Tbn0e24GYH
ALGlrcbidp/7jWK1w690s7RwKDLm5j7Sa0NKZhasFK5kVoEfS2LIrsaTwSob2h6Y
OeaoG253vzJ/nknHOn4vZHMYZZXCMezfoio4rbe1+OkEU5op+y8/8YI88HfkHygb
oOo4hsFPQILvyN9JhgrSprmc5CMng+ce152SVctLIxvseniAphCq7k2IoS7Dwiq5
nf6fHlWqMZnYear69jnPuYL6USxJ4V0HttoWED0fnvRbll1BlNfB8IKuNxx6TcyC
8KQ3T+gk2rkBl5aRfUo4U/osR8IRqJhZqPGlQOaIPyz+xk73RUs2GCR2UvJgfkCb
bN3NpLmApSp/9XpjMqKYyijzYRwPEcymFDOitovKiz6VHJukZJ1aIKyRfCKPP2RK
LDYGAc2DY9QovFxPONCMDiyIagO9DT7ObLGXpGDa2nommgj0P8VCadXnuJK5zGik
ZEZmxiKch8F3586afUC6CQ+xZPEFg1ycegcW8YtAwHdYCB+VyEYOMLCZF0UJ7h7L
pWs/4GHchoDVRZdcMPAGTKsdf9ztUopdgSrZmdRi9PQx0Uz+RaDt4ykNgObKa0PI
KbTlXR/WctMTADMKyKku0vMvnei3Z5R4LeOUyZn69Z9KMuG7MkkBsUxiNvJEThhD
D0q2tq+vMfBe4TzbTKpVPHuCNKhpsPhPE1KwwICJuXZbnZaWTccwJBotG57/wqwq
R8kDI/O223WLWfPSHCg6Ycu63tJXFjExna8kc38sAV6gkBS4BC3F7RZyrjeXf04G
RTF8pv5HRTUIAyB7lzKQPPELsLh5TAYO+uZrh7gpwPSVoceOo4RkzXLGFGQt44Qa
asPtCNMsf94xLMY4h7pawk/hs5rQwW3D4VXstXhH1AQlIGRDH5ePWCKeDrJw76Fk
TCXHIlVGtlFWY3E48pF6Pa4z06hOrW39L18why7Jwgxc5ymgNaHgHMLmhTP9zBEN
wrPgqTQrQAV4SrGTIzQv7hpc4HnBKXHxh5qX1lJ44EH611DEvypKD3ATgm0bxUcT
xitzguhjGKFHx7E+W0yiSWQYlMGrGiYeaQ8DubmKHtLTqacqrSJwNTVDnh5LaOOW
pR4ZzZegL0hgFg1pbU8dFYsaV16cD7IRpgjYgt1fTHcCP5DGtX6PeCDG3clFKHvy
nI2FVv/9JQ2gSvsy4z3Wjazug9YW4oLBZ83T0UFJzhpcUm++WKjAMYdhz79ig4De
ZpPMgmJPaAZXPz8vEAtHgX7Ku/sFTHyXVPIGV28CjnFjjQ43Eia+YCSIfm4i8NKO
IbRaqJBFmuCb08bE4NFcyubSlfTseFsi8EEOLsivKaoW7gdYgjpzy+BnpvdMtDBs
Nk/Enp1oPKRBPQnLpaL47Qr3MRYRReBCKz7rnOzOrVw5g8Ru2OdWuEtu1OCBahxt
sV9TpkKKdaUgQb9EdKBjTOzq7MgzqeM/Z1h0eq5VT+VYuYy1XQxRdP9lhMJVT6cT
EfbxbRwb3deSFQ0lEl0SE+u7TNPEsvTsoIVJTcUdFGmqIOnQPSjPVKmzkIH/EirI
uuyjPP5T5/hGkPv/ubWin3z4GfgHA2FIEcgchGbFbuYg/4yThpkFtFnw84Ihdbui
OYqtO2PacwSZnGi/MUeRgjSbJ6waH18CfGubGA7gyXiCubt/iB2xrYA61PG6IkNc
cPuYMdNL5lJYyT6i9kdEd6iANcRrB9rGeSUie9hHlshk8jsv5ztCFKnf3SAYtFOT
jT2YvN1DSAMKmELWENDQd7yd5qny0ZRQ1J2C97EeVjaBixizjGupCsfFuM2oHUqB
y43o06nR/12aJKJaaDkQdV+Cgc43lDZg4VGlE6je25ZxjBpYeKZnli4+TYJtmBay
Xvp+zK8e1YIeLKkwgawm1omI9tO+9k1EVXVmb17vYOIYAmYdf0k7MAZXqgxGynJZ
Zq9yX4+UhhO6saQAGK3DQu8P4XWXlJcKBMEcwDxjyt9XoYSVlSnk/B02C7O2Av3M
HVxr4JH69J08V0EerqaRD3G6JDyLmAsta9sINYSlC6JMRYbEReKLoN+ESCKgyesC
gO4apXm9g4EC3rpZ/Hk+p+03Ji9a0hksY6VC69bsI4enHkJkogEqMWR1ny2gAbta
SNp/0SxZHDrG0Ws/55gWbgXFqdBUxSo2DvsOyKLRrHcaoXh4fo3/KfpESZ70qlBb
Sg7KBBj1SBcJE2boWFNiKEvNrFSY0JeA9+bHkbLCnD/TTAOAV6IIrBtu4OPM9blP
2hULpomd133wqH78ZDKi+QAESahLQvgs1S+wwB+tHrNKlsaeegXVAmXSs7UrLh0f
FO6J7v9TPrPpRwE27kki2YH2WrH2U4Z2ZYwZRqKFp3UlB9EbLEYsPKtNV5Tx1D7L
mp6MRA08ybD23s0oP6FC6ct515CTUGYAFfZAtKh1dpBYOMC5+xsA8DSTQNHBRblM
W3cVnHpo5ZSGBXoJdiQxHcNVv4L4aI0UlmehBtyMtkrvOITHdYRDliWlZke0FR/O
orbMIWmCfXiX7O/1Nvr9pFurAB1Jdkm0XDe0i/ebidr8R47wp869ER7N6DKDihJM
ibi1nX1varE83PTIRJO65zjH7QYusEyXrL+7wjXBGdpu5Wjykkfxc/g83CZn6kks
NRaL/mDvxRFyTfZoNlR6VJkQbeUEyRMAO8lgLIfdCyf5cAN4MMupUdg0nG3P636D
7jEYtcqNUumQXvtvzmE6L9DMFb1+Fy63lQ/S9saAOGYOPeA2H1X47NBOZ7EO8Q4C
LLfMjAuld2qYo08KEz7C8TQYVlHZIPA0YqyaIy2D/XJZDdrcigRncxSmC9ShzHAo
yNQVtEu4AuhYOk0PAmAeBH2819JZAv2UywWSy6igoSrai3RdY3zMviS+OIAxNV3R
j1BplGMMJkXXl+HjPFzwUtfX5+EEJsTCaNQC5Fzc5ySM5GcshP5yVauOW5ht5+wz
cAl5ONiWgsmywJZs5KISXK2jIr4IlTEoctkm4Dmq2g75h5DptDL+SBDf6Y4Z4x17
tVCJJe20rSWqBCoc9Y0utq0WrmGT/sb5J9QC4XE6RawyNUuz/whyKp4YAjRJP3p/
hWmFKkX3+Yuw2gZkDYxwjj9nBBXDuOyPwBy7jUCLYQo9JMg+iEF3ENpBw0HQn2VG
LOnBKvPUq3v7ORUT3YBJeEuF69AYUxZZA3O1med+oJaxctAaI5k4AjoU8lXbf2Fi
bghxMCehfyqlUIM3DmfK9mWNhU1zr0t4QHSkSCNEOO/Ar636mK02/4dRJKgq978i
xzSWGymaN0yNokH8V3f7Ubtwv+0SdZvWVQSj1qphRwAmVCQpVEZ5JvoaTxdcJ6GS
uRoU/XrbXtmtfXCZDCf+xgo/cP5w7DempwmrNDc/ZxgG3f5SM6nRVN2tc5CB/8j3
GxAWSYrhEUGYtgIyy7IWrsyJ0mbQIcd4ImeWLnFCPzWglFZuPa43jRSdK6L3vm83
0eJjt76s+RATPUHbwJGPpl5v+E0KrYxMHRL7SEVCELxZmzWZMwNspoNnIVlAvDAD
/nJugHKx4XpEs1J0A2N+NTsCaKJUX6iEwaFDFbl+ty5toYC+0qKtaqhRYyznvnat
Bkzkz37r+GejJ2t67ZxMHdGHgFDqDWcAF/0HcHPTEH1i+NbCCI/T0H/FUMMoOVf2
qUfdBGjY3JqHhrsZAWb5HbsegCEgURTeoIAd3oKVC5rh3ZWVHzEo95qihH+hQMmO
MvQDFz4jGgJ9tTsrU/budLjU6+yrXOEw/UVRiHrLD0APrkDIZWUs3RaLzYhPUZt8
qWAKsggwgXfzCSMTXX3EmvN4IGjCAAl4VSB7NCID5au8i7CEbbNqKC/DoB2BLm/i
ZUdAq22cg1WCbU5f5FMUqdayW6JfukzUg1VgEMEBhhmve3KeLuHsWqZsO9JDlNHq
nIXRBooKtKvJYW+JJIO0uUGNeVk/t7PPy2PC5VJ69+/lxSN8OLHMr3eqC/EmMiyS
Wx84QtgD6u2W/FngTq0m+qBvx0Mg2yjmIFzqlMcbBAGfLgLICuTzgwIWFhdWRL1j
AMAo17lU3Cbk6hheyuudJ55CwW6EtZIkaKofrfpQWyLM8iwaDuKpO0p90qxyPYti
Tm4TJE4b+ArSYnyTm5s0lu9rAnSXmtvfbM2bl9WuQWBLI4N83RpfhEWvnu2g4zwy
2+OVyIGcwAj7xfjcH8aEJ+kz3mqjVrXlQ3rHfpfFVoFKtGugFjVx5TtWeqtP3v4N
9cWFzi0i1/zT7MqIuWu9pCzGHRo6f5tLL5yWGNO5MHaBFAhj/NBCva/qeB04X/nn
Qrug/Iss+neklB2VRZJnpBJIMXi8aRMAvsW9fD07nSZUVsHJpOJxhwgVKA3xQvpF
poIImC4rB3tRGQATuztCsIxxHC7/Tc1BJkqTBzTYxBD7krvQVQDcIXqJsYXYg8yO
IJ5l6ukhYlRFI2gHnKDqGVMXk3ESIXw9Z1ovbITb/8YTZaU6Wq9IPdy/r8Tj2FLi
W6yJUllksjeGnKIEVMaaT4jw8tivZmD1NoW+VPfhnUYXLh57si2/3WgXnjMaR0To
f2spW8fRVeehPH6tzV7++GtS93urwWIkIwjNrLC2sviKuRj96QPY+u7K3OE7NO7F
nbluj+5zOCuXaobggHhRdWSkExkXEoB+jOZc0QQJNQJpXBh3Kb788KuYWlgYALUl
l9IfWL1lFIvkzTDkdhTmTyhXcpi0yH8hQjZtKk3qseXhq+TaxM6OXUcVtnHIfTVh
41xOqMKzDKpBlDQ+RhV4Z6uC3ksiEapU/AVarUfeI5OOSBM80G8OHR9RBmTQedU+
OloYtv9vu0sgfWconKRwKkt/th42yfv8Ae12/WMo3qAiyhkQwbVDKey/IYLvJytP
MnYRpowZU6Yr7Rx5kgwPf/118PHf+rMMs5q2QHGxBdir/eOvyc8yDou4sXtGKklj
2kDY6F/tQKpq38Kr/KDbXa+EMxLHyD2FwE+RRAIEgY9JlOoyUfHjHyCbVtQaUMDw
2qJvXBYOYx52EzPKJ7uXLfs+rZb7fEf1QbP1o0WRoWuHsMifFs4oAe2wMggyWIHL
TT8gGJn9pKTSUR21CRrIZ2JyKkbl4GktrnbGD3i+xY6dXpA9xyfqlzFQu+cP48M/
EiVql4D8BWUmeK5YvoYj+2xVQy4osqTDJqJNry+qxRjuIY6Hbk51bfhU8QFIw4qE
EwJnUn6N8QB4BrM8F/WpwKzteqk7AOmbQvZ2vrzv9wSYxFo03y4MWLggUwyiQxjA
E5mhV3FRJGljlUorFnxeA2xrz5JGHn50shFaVfhOlYmvjAQKw0m8awNQE+ZHi9Ip
2WazMMteSYB/QmIlfVfcGjRA+a77WDtXxzov59v8AH1MTVR681fGSTqS8HSulVvS
BIqBYbrGQA5kRYz1YbNRfwND4NojwlYQj0TNP/i+LsKoqlkBvPWSeqf02vk+dDzR
pts38QFxwq62sgxP+f0RmFtmoFNT9x9RezHPd+7BiIAjZz55vaDH1z4b2RSToBHe
p852HH8ll7zl1SKS7NLUtiVecJ3jpCggp2/EcvvkLISeshU8QK2QAwkRfFquZq3+
Q4yg78Fvs9Uv/TRp8pZSJYNStO2gHmbv4knTn5zJsCSbX0OFRyTN37JT0itOzgSd
cMFxQNh8FKNPvl/0261MXUtp+xvdbuXA8f2knj1r2myEIuy8yeW4kAhpCG96Fyda
MLSzHmfAakVK3f/gMXMTPyS97LihCPQUOvZpGGo819QIkQHGclqdTg3m5hk7ngyi
lbXQLasP1TtlPRaqeMPqJEhgRuDgFeEeuAG+O24NPTFUlIe2wqUzBZt78DFqgozg
vB70kuE/iCX8lrsCXOHGFXD9WCSoWqmA1eU9lbYbPEtkLQkkdSuFpc0+53xk3+4A
Ocwpw618KNybik3n2Qot2Gf66V0AOyA6Y96g188UdpTKxUaI9m9HfReX6EZ1/os+
CpRQky6bJve/cmlPkSe6aqAvvW8LLfoVz46dfKAuOPnzmG9NGFcrAUChkPusfKXj
jxLMm9bx9iH51+X9Gh8oJEj80ozlt/aY8ZhsR1uYLBJ90qkB6GCZwrmkoEJcDBAK
+FUC2uQmU8MhHUOFr1tniyVNHA8yR4KfV5qk9soKowk7mf+QsuVCAlnIskt4bkKy
kKcciBCiON7IYD2xG45iMzOy7+j5D6j9wDlKVLxIPE36J1UHbywvkqTIg9X6jXAQ
3CElGccYImjvdmPQ0P2++d/SCq3Us1FdCjGver8oUa2qKDWnpFCunY0NGPa0bA0c
BFvagHX7E2THkugUh7Ca22pGYCmn4Nw9Q2uCIl5ExVpfRgRsTvkbB8q/ICVz1qpJ
qnIr3m2ehWpHSdl6KyZNPT80jHoC/+PpSJTqHKH2pAFxNH7LL1Bb+8AkqxKKzbiG
uRDlD4Rwq1zJY3FLRlurDxbxyzT1+VIEZFsG3nAy036zw9Vtz5PH7maIElNOSD4Y
JwPr40C0OkWErGHR61JKBBNWQTAN99pkr8Yt3I8lFTdOfsuyEkR564ZuqpCA/vKP
eb+ecthzvmTe+X/HeBM5FxW6C4G2KQmm6MQN36K1P9MuHJy212wPwHSGfHdyZl83
g7RdTbmW1DFTD9MMW1GOv2r8Zj6EekM2EFCZU8xt51ewI9qA9atbk9gj6CIpEXyc
8WUEqeFcczOX/hlw/dlkattcGa7vw3W21YqhYlxBuqmiU7QesBnlYeHSdqabLtp4
wZPqqRgf1+NqofJ8uGqyqxragqqgmv5lO8D44vdNO7bSytWunomdW6hXywiPfRdP
CnsyXTnCrB2Ebh/hq9zZ3iaJ502EBY8ZTdACYodRM826IUsNFnrUrmkJahawfihK
RuD9h2+f+ks0SeOyQEuyMT9F1sBOoB4wgJ1nAjYLiIp9Op7kzAi2G/Z0IH3P/oVm
GVMAEyyIVPG4TbCbHCaXcscE80CLbG9LjbWw6PeznqJ/LnQndZAfnx7i4nSv+60V
oDA9Zx4/+e903AYtVx0IOaUMw+Is2+YkEZWpKkhO/fCA3fK/zf6mXZ6+GqXNhrpz
Bbw3Ev2NNIsdqHwpCT5y36tcFXvVauEivlwTTtoZV+z39lf+jSCOkoFJkogyVWZh
UnKpG4TRh00GfRK+5G8iagnauYbhMGHgOcOb8bBdq3jlIlrYB1e6Xaidpbx5j1E5
SFK4gKaRsvYUybsz3/IYN/eSbRb5yHRi+Vz4dfLmFXMIqdHNLa+uI6ZJJLfeVD9i
sCB3SHaXWdhrOdv4/xOvhbr8eqcig7nIYdFlvOjdHKjxEDx64ipLE0TZggP9i9Hz
v7mdlqeJck0xs+1EeLT12U5pl0djXPdkwpQiIcfAAm3MPWlEFuOJoXOwulYRHXSD
z9BAWwj55tDQYn83ZgHL1LfvWNb8sbOb1aqe2sv1X0fuHwOsSqR/1OoTRCyl3hXq
OZIt0BBfXyWlHtKVMAX9rBwzo7N60yDDkVqyPI1VxkrJA5h6JzOtryBUjxTyWxOp
zawFCcPfpEldbJI/kGp27O1ErvOaPmZ8n1hqpNqjLoSa2miwOLBZZORFZNUvUE2P
gXmmWJB0OTp4FyiWRmPylf0WJQDlA+Cv54tNR+df8TXrhWrZ/K+HJTQ1ikRsXLC9
PO//QBhUqK+VTZcDhxGW2gAzA5FhwQ6uCJLVh+RtfqUaMK5TyQLAM7jTwNjXHNZS
f1hcHoGAG+JZ0tlI05wZ9WLgPenvjDgpEEGxn3oPRtHS4X41NZoqZtD8jI/paNxY
HZp1m3x1mqsyk2WPUbUf+7kvE9nvsqFTR4j9AocyLmXDsyTk/jbAfKgJgJhXPe8i
HNDWSYJVVd5Qv0qmLhDg117Af6ZlRVMiVMsmrWc4GF3aWlaAFT5p3kqagkiNRnXU
miZmwCXgymgRTp03427kXqfT2Iyx6oEDegFcYD0PJjbLoa31+DpnXMffw9emHN+w
BFR1mND9lZkkevNdqZ0Su+xJr70tuYvA2WbgMlX/jop97URWWuLMajkSBNVgr2yI
NhP8mpUptSTg21Uao7U7MCjO073LdPT9Towucjx2EnsrraY/rMVE3BAHfV8CLwA6
yK0ZElcQy4ioHR3BiKkGklHhi37J3qBOV6dU12EQQU+lcLL5EwKM3ZU80kXXUOX+
aNppFIpC5Q/1+AN/Y38+HMtHOoMG5H/rEFruX5eXGv/1elN47zs6MrfC4x/YANJe
izCxcr6wZPM+BCIoTirApkyIcCq4CH0sP1Gsi0ypK2jLED0dUYJTKEvAb1h/4oiG
atdxr2Pcbg8DapA9rfIjm+WIUM98BDBCOxCT7guG9O5gHD30ZGwQEVhhqFJkj2vH
rMGHj8FzTI2+7a6HrLvX64wj/y4tbCReQqdmykfzAElaRw/RulmE/+3wda+IvLec
FdJbAKzAJU4s4hJkIGh85Pxp14OJuda5MAWt1uOCMcSjhA7NYDrFk8P83WlLJh1G
Vh+SaurGYCemXF3Tl4U2toiKX9z6scZllc2+9Ol6RNtggD7ALwInNEaNnIWYi82V
8vaR8O2FwHXB9a11csoVImmaGuao8sc3pdLslq5J2Bw2vQ5tjuIAGzuqAD+TlGZD
fGWAO7gATy/AJ3I4E+yC2Si82/R3ZXQ0JoZbi3WZMIrBmQTVFVHlq0dJeSAZHmJq
eGA494xJ328wQcDimTP/AKSL4Vrzk6dwST1ngq4o4YWNOcyTDwprMk6XbGW8L5CO
wLzOaiIb81kA9WK/pZBYZLlF4LHcWjNVh+o+2xSxTd4jNW3kh2yi4/0Pm1ViqDSy
iB+7nG4RxVtAHpoQqyeBKwuMkRE8d+b+RTIu7/8Lt2Glc+ZVC13Gf04pM0o4mJEa
9HHxA80jTWpCxuBTeAyzNIJ57/p/Ge1dAvodS6AnZfB5kLGwFWmGQctkvu/fTxjE
Tm3czzYtkNwxiydWFdLtEWLflk+kX0d9H8dbyiuF1j13h/1lUEasYJ929N8asVI7
mNEQ1Lf71N6StAcExz8NzSvlELkITxhaWYL+VxUBy47MKNPbynB1d8tEzasqe6Z+
EH5HVt8FQlnVjwZSqkvck48IMjzIfZuYUsFI5fHQy/WzM+psWZbmwXVFFmwWJtHm
rIP5DWaJfjF/E9YB1ksoF0eo+hJdNwuujb0sa2bteutUaxON3mbXu4qKxemhz9R6
VdlYC/tTcioeTVQ8sRsUBnb4f6B2xKDSk880wfquSDmrNqQCUelLIZADn8oLiDkk
rWB4Uwy5AkD3lrPRCmbk4Coy9n3pEYTRcT6BrALT/m9kJ5d9oJMjXHfJ6Ub/DFeo
Wg9aAvMyxFYn8walt+ErQBRhy6Wxe3zUP0psLr68HGeO131jtmtijg/gbTbEUDcy
pOn+uNmamn6700S1XIRJl4+EqXRQXF5y+OO8KIRWjxb2RUy4a+CvtZILAkt2k1vX
94JkskjAeZF0NfDxQqG8CjjL9c5esr040D9FRyra39JzWCrRZRuoAc0vsiHOLsLk
m9EomgQIpTOQtqP7GNwTG+aolaMnglgtWP+8DgzGxe6xjmL7URv+1YwADbYF++iC
AvAjFgUfSFmi0iMM3k6ayp96Gw1AXsdYyuGGgUHvR2JH2RiNqTaNJIwoffcKvdFf
MdVOu3B+JoQNl6jGL6UvaZdwsAZL4k6Oiwpgt8lH2nimgXALa+BT7qwGLPLyAE+U
Oix9IOR0/vwu+P84xVbQUEdK7QpUrmXhCNJ4Z3MBLz6ex0kpm9hdTYPmMLRQU3Fj
vHrkZAUtfb7l6G52v39UflNiN7qgdVoxS2gz3AeAFLV14mC+oOO7ZLFq8dyCnfke
DFnqGDRbVB3Aokg0fDbFMSsUksaBHJ8sqYOVIeqI2wQR7/ciBkOO50kXBsKdNQni
zRKIOjqihnfisiMQ0qDu6xMqkBhCxFZD64PhvrrB/LPsQuMEcziLceEPXnaxYi+i
7bXDdpmlZevSq/rDdyEMOOxMTpZml0+TCC5wNE4zo+hhmnWmXOBS/xsLqUptN/9+
RtsHFsVCmY9r60R8uHD+QXzbbzL+49PnmXSMNjX/RxEvEa+PphLXvnRnpd47tqAG
pSLyCMZ8o/tcDyi/KaIbFDf90qPyPbN89vjuOd9kQbS1BkiOiqfQPp4TTHcCv8Ll
RNcRM0mTgCvdximpWRB2t4iMwTJedKkMIFP2DDoK2jA6D981hphIF3dtBPGNFZNX
wN0JLxnBP/8Wq2nx0n4oqh7FaIiNlP7iR6q/LQtK2hFQkV3raLU/JpPW0pi0z99L
pry6z6+bvcx8GWFoZLfrunJN3r4IdMZBeOn3oBRY4rj+NY4sAjt5fX+6OHo9J61k
fbxf+NSeYuoEU/XKNWT97JmXhCJs+yj3Ce9eB7eZRBFUe85KekhPs9S9PEDPfjEA
cGQNfRm9k/csQjmBgM4kv5uBJSg/aXsfElJJ12i7612eT00n8htyoDb5faIRdf7D
vleHPsgSXLl1cwqL4HWv/KLTTo/HxnDkSRRQp4J4rmb9JNrJ+scavUtxKrOYMmES
MBswG4Qg8xJzukMIkbBEG+9jO3d5BN+bxzLFc0aZwUwK+YWkTDuns257fsvajBwE
v0V3gXqVJN4C9QiKcXcGXUJe8CVjGmeiY6txAX7aiu1e/oP3mvwQAu8vRxT2CiEm
dXQlhp5J4mmuYBxoIAY1PGJzrR3eglomE3qK74wIPL5wBBIXL3DyAbH7iIeNb/9m
C+SeESIGT+OGGzJlo/Z7nSiksR/1wGFjk9UNwjXftM4VPPwJHG6SxS1I7mC3FR1v
WFYiAtQ0zSHzjQsnmcWOxyX7BI7mfmz4R2MY64RnQhZ+TGmIn8tyw3KplYAfqqzF
nAqDVPO1VoOWLYL5SVguauk8Ltl0WmnJvCclSOltI7yvIqBavb0Oi97hejk9mwUO
3Em35iKM8uYprDULjUfno6jvk+Vau85MRH79XX75uJQm2lUeiBXwjrNqr0or9CF2
E+O75yjqhHYg4IlgFxYofHCyDSATHtcF9EpN8ryfsDbE1vBUnUUCMDA/xOHGiisG
oLsmIYchGQhHr3gGLDdG9mANtiwPOV9/Vq3aY3blNRjdVxgvOWKGzeN/JZZxdvf5
xgtsTLnMt/l6ssj8Om8ARW2H/gP1xSZRnyQWeZXPpRcaFAXlHEfxlZc7Aa67DF6N
xVCVbZUi78coUgHgV+/HAjmOnuMMtCH/kBzKrHzsyp27YyOjxb7FwDO0QnuTH+el
G1xwVjvfle/+u3Txu8AcljHNV004WL3QtYtEMocf9dyu4v3vgl2EqG3v3mIvdvtA
KoaVMTQ5/CO5yrnzVpquXUQ5/4sJNj5YhUuWGjQjOs9kML9L5Oa/2RnLC1RPFzAu
rFZXfBf8PX2nqxVh7OKrD0D9ZvxfsYxNNSWiPkgFdV0ksN2oB1gFlgMczIkiLOjW
iYBSdZV7uPGi41byTwyipEjwmBLBPdW+OFS7RRGCYq1vXQDvmJb96rtyvsYH5v3F
VB6NJB2ob8fy/JU/1wPZMTToOEl89Vqf2SVQp3tVYvTB2LSfvWTQ1leN/4QMfFUt
WQTZrd1Z4owiBtfVqTZwetxMFzhzVdrG1Q6ZBFYn3SVux6VlQ+77Up4neodsnqve
v4mOvLH5yVgxlFQHFQPhHyOT+0Pd/NBnpSsQIBF/+4zvMrs+sOIybCFIdwuTtKcq
3zDLBUDVViX5Sf9+Kz0OQUNiFT6/q3ubuB4rkFSrOAdkWfpHQDn41BSVDsmdnng6
sAuwHckk94CC/519am0Lxmbj+OxU+voy8JoNvQn/5Qffb1hbUnM1UjPgo8cn0OzH
iMMH0DRcD9BOg22WMKxMeSyCgfAOBknid7megDnfl97vw7IPBR/I6gZCtHERWrdi
nZHHqRCekZtSD8+LpSkyLV7f4xUBVlEue8aFEU13+bA9zIBoFePsFW0ggb/uYew3
AbGlNnJLvpopBpaQyAuvGXMv37I9vGgP/oXPK58PCREbE2E6QWyRV8TCr5dcyfRL
ZqHIEh13z64HWgNq3rlf8ye1m5mh+Sx3wu5Lo1Y6z3na1GdYVx3g8h/kG4pW406P
ZC1Nde32FCxggJAQunQlulPdBWmd1HmBLyc+FXMwyMFe96TSXcp2XZXnjMQBp5N0
givGcMgc0ho59W4mOwVipk7XgmOLYWSUNaTvMmLKRjE4pMJM5GoC13+btHELWd5M
SRT37XXt4tBHwNwKSuP92IrB6EfiH7mpT4jRwLNoAD3af7BoKFAL2V5Hz0O4vXKp
7hH3Emufjf5h2zkmaLgwil+xR/7qNoduHOZlsjc8oQ6X3xePjte/fwNlZkn6pT41
3U06YvWT08ySQSHXsU5IlNO0DPNcZ4wRwEc/hf0FpFpj54dzq8jtXZrZPuqiD2vR
wClrbAmakahBc/73Xh0WlBSDB327sNYd0Qrtu1nm/KhRsSlLV0gXZ1Qgs1pDW5DL
jLMNPhj4ZQ3STZHfu5Pd8SSkzqaIXnbPgoTfeMMOqpssxy6Qgk0YqaQxwtvZLnir
IPDKNKiYJgAV8oZBnyphILsEMGKiXEJ4CwaeazbWG+YVwZC8W8V1nKJX35MFcFw9
QrMxRho15bRACUC4dQ8d4R9Gf3YuTYMsB+TaXgnS+XVUgL0byo2qCrFox+VEbYlO
Ne5Upx/CQdumiwtXDDzBMct2pz0VX10c0RqeDPlxdHKQ8ZhkhVDOuUKW3vmZO/FH
LPtnYBSZHSxbQl6sRric8n/tsINUnaMV4arK1/qFWnC1zRz51I2NWJHt3NiVewNq
WcFhxYztsHP3/5aLBc1HAxVBEYNGuUW0jiuQM8NNL1e/Hz4u3gRBKVXje1PaqjeB
sBOGB6D5SBwnPRlx+eiS6M5hVIcw6H8+UXTlyX23kbOqrebVCJXBX+wCsXze9ZwI
XmLw5gtMx8RWvCa3GmWzc2nzaH/EnnpadNmjVVcwJASAWSIV05z3Y5gUt97pm5Rz
lwu6pF0IsZvBcdAQLtcmLTFHGE0iIbs68XOUP1COBRvzxntPT3E412NS02HPG9hD
TWHEkasYPPeIlCmy8WtukVU8w7bKs72Xfpt0jRaBP2tdNdE/4sNESmJ+TxOWywTc
pxtg4SVFcqyG4O36xLGoRnUpNOZxEC0ByjWwS5UbkFo39I3EuQgXZFquhOYEo24z
GQnN5tBIbOW70pFfwb8WAzEjBCT+IMSu/1iboTYOtZSooU/1SbgyK3mrU5XDLERG
mmbXxQdV59AAqLeILMstZXgSAL2bDS8tY2Ci5ffFn+K46vuXRWl89fDIb3wqVUjA
MG5e2YeVlB1Hf3Rge7zZYA/kRYGSVmlTwdCoVeXvQVXnLsZ3xqrwP5KqGWkIIur8
CiWHrqkcQ8tqePioOez8HDfBKJ65tj3B5rCWmao69dGuIh4E77p7S61JmC+MUpHu
YtSCZHSSPw4GYlXuAvsx+mRnogOAYx8Sx+PGaGmiPlKxPVqGDE+RLA/icyvQRxGn
oiDkYP7NYjVf5uJBSWe92TFKe/Hk8Q5QagzCaoi5svXlkA7pO6yba/tb2F5MGyMT
68ZDrVl6nCvHhb5oWDfkIXyUrqZ4VTtsIYaz78usvHjSG/Ign3o29g+zsfLoKF0M
TTEQJkPci539OPZhwkShSfov0EC+sLTbKlrnYH7lraiOQxJqepypYl3xGSPX+++M
+ekvXwVMfytodz5HL5a+Au7wRwxarXJdeCZ1USux/Uxzj8dbod1eccAoF88YpkT4
WsJaljyb5I7RhVmCo/Iz8rpAQS2tXM0CxxxsIC3BQ9f1S98pHaHPQDHX+0ESbRDO
zqBPkLLToTaBx4qSk3wDU3254/iikMQXlD4QFD+FH4zC9qzhdEeChXExkTrWcT6t
nFVVR2YJJ7XHcyNb6McruQsHMbWLIQAPWkt6TFIuOobs0qAhLY5vpPKVwTWgS1xk
rCzUkyFpzztJX3vTutITUDf5ZEes8pGNDrfq7AhHXjxkMyqnZbPL+U2nCWR/5p07
jXtIoRatqNkyETfOwF7XcC35ds9XyLw60pZEBQ5B0oW0Mm8kdrv0fijeWEskS8ew
+kHozvokvt/nYa7PTyi7Rfw2e5+pGzfirBA1RDseBPwDHRir2+C+OOci3zsyddl4
NNfx3sHsJkQ8Ia8ChLGc9dWYVTSL1ys8KlR1TiRHzIgQzHArs5HZU5M2DaAwpnCR
He8a/olQmo8hu9CtuSOxkU25Hr6kiEWLJp7gYnUYr92fi9EWCqmmmBqhhyIosIR3
gBuj8edhH4CNE0kEVnZcUos61XSjOOWhWZYQjqiY2m2v8PXruzJ9EJdDpJZL+Tfq
vvqqez/j1aFN8eV9eDdlaKGJV9RHdL59sXnZpiuEYmht3t+lIBTpQyBSPv0eQIq1
A7qeB61JhalBe/1RL0+/ZJJVqojC+nuNNINzX0OvJTIsspOdPRHgMPuGZqg5xBqn
BvJOY9GTOMSXPcgi1MkILhKK6dLg5fqCMNJxVUT8T/nc8UHxV0uKTTdsdzHplMKj
Ip9QgVbla9BRnkkK3XLI0isWXFT+pNBeEyisaHwMnLgaQAhCAnLdYUNPBXnqoUJZ
PlSoXoxF3hf1RmzjCC6KnSzmj9i5tRpUOWmUrWn6PzJuLhAJAvi3U6MdRfu+VS86
fRZ9pW4e9vDW/C85UrkE6Ccu2FT/9UQOYbfv+Nm8Vvv+ytRc8sFi/8fTUkOD0iJt
p0jSQi/7pcNHnp+l/vVGbIK1wSxD0EnpBpSS6eLYIvE51yGGzlM1gaiBrI3XoB6v
eLHYG+VmfTeObBIgYQ1OnMz5giduaTcYlC2JNUU+YgN4z6S4Leuc3KWXDIQRuhUJ
hi6A52IQrJF6ylUGHNfPs5fXgNFvUWjQWq28Gzmwg3hKXZRoH1mIFXJJayd54RIg
BeT0z3SkZ6G2b84UxCFNsFTmo0nnh40fESXLZvJ4Rv0/ujIwa6bxDpNlmfD1lmPC
Hfe4HZJ/TdYne8VvICQ03iymOeyVQungGzYiI43e1p0YBD4yNCXnD5f+diKMd6lC
d7PelmmbLazkOaap8u+o5w/wvZZgdxUr/GWbhR8jglkRS6O7sBl18tQBgHPnKjpM
d6Z3/LnN00+zy7HO2u+kzlfuOS31MwBxFt150CxNMRbqHxl4ipuXKYSxQQpZcqpw
SeYQTkwx52pscLPfeIlzpVlBGbUb4kUt8jdL+Gne8WejLI5Sqb3tDJLxn0iX49uC
V35MIGg0Cd4x2WcraWO/eiOfiPfmKB5Y09zP6XF6TvRX3Xk29Uq/kptNify5A4pt
tAEDM4uAJmg9tQO/i0LuEULIJf1Uw7pIWNhF98duPRZZeSaXxOu2wSxfz3q8XDSk
nXrCaWTyudlN1gckZsNdZjyPMG5SXFj9yLBO1mlkMjQ4Cy/ldWAdU6LHDoaWo/Qx
c7L46FC8Z9nkI5Yp+Hfgauco7A4YHcIFsA1gY3CX3di1iZT2nKlrWnRZnU+qKSqp
R1C+37Pkavxo+8aLxSS5srQXDINnHGZ28Q+He9X8kJF16d4cYBt5V0wTB1/14RCm
IYXNArSvyBVQo87CjwVCRFjuqfCv8b0AuNOSg6chowvF7uJBwWq9RUcXW+edZ9CJ
nWJDEPSsao3uRw9gNsgSJz++9Q2OWXWgQjIJ+cykzYNmZQcnOdSp/lM9wKJn3fhG
Un3oIXlxm6ufbVTkcT1NucnYr+eLdIAW7/HoiElELGvueV8NhWY7DdrFhGdnm+s9
7tZAhdryjSYunV3M8qp3cNStVcuoybIdmqGmousvUun/+bv4WHhyN3xDiV2d+T7z
uEuAgLaqUNmB/vXDQwuSUUeZX26n/IQjBz5SVzvZ5sS16b4dAjuzpFoflep5KlO7
0QgHb9q8iE3KyPBVaeTwTRfKoQ/gOFJbPVZB1S/0nZRzFwSe0g1xQqR12gOQQ8uX
DWBFXtnd4yDzvl+jTRepnXqN7kIlgygfazFalTm0RZM4K2ldzeaCdPdnIMzQYskk
lBvtUloho+wYurif/DF78vP210pfa9L+2sGQaX0okWJlG+zfbEjWSwF7PQ7L8jN2
NUDB7QH3vMlnCN9ZoO/lnJj7AL4mrLsRNe2SkU5w3BflCJlRnL7CbOktJHl4LKFs
YdnzLtW6lUFHhf5u80cGppMmJdBTdsYZdV7XEoYDdOXY69q1DrWe/Yt/+Q3nuSSH
E0tAn46QyLJchT2xnUwLIohAqQu0e5SWYa7xCFyLSBcPWL2rzyRsDhaY3Hxc3s10
pp0Wev0eL3TGkZ091S8FSUOlAvurfNqsMjXNa32fGhjbOfrwF4A4AIs+h+bLLiu9
Yuu4Ru+7WfcxBjqTWakDy2geT2DTHrJ5k03oHAH3CUctRMzF2yip7/hQ8uVxiyW9
aCEOJvtFYtw0KUo7EX3BfILiulB6Jefuta2uLoCwK7XiYlu3E6du+17Bt0SVAmkj
31yryLQMskWdq1aILRMm1cP8gYPf+HZx1Yb/Tedw1ymy1wTt2WuGni+svtpwPHPl
d71gpm0GIQ85dibg/84k2Ll3CoUhV1rQNVTNFBhpr0AGWPKaAS0Oem4Ip4L4nBz+
mdKDT5oFkSQQJqa2khCsqwzpP8o86exbc2jr28zGslB7uj9BQsheOwjsnee0BFmL
1uIO1B6+D5OrRrWVIX5wFuZWa06A8eWWUg1x3KH1qNDUtOV2zLrF02PCBT/tnJOu
TG6KsF7+mmMlDt70Wi0Lt/LBTrHvWkoa2uLWYGlkIvjv5TK+ms2Xyi1VWNi4eBbr
KX+xX2bvynwtFNveQPxxqXsGaeJ7Bzxsr6ab+otQ4QGPYsGGtnMFyy8EGO9sYj+O
TJZrxFA5EMN6vvPcfRdfPxDYuYCZn9P1hxmKhwdk81NSA7ldMCIpcpb7wm3cTX0F
ou9w0l3aAOaHOb9Mz2Vb0rpT+3pZ14WxmroUu9HfZiObUd9PWe7S4+2zAXlkN/nw
mYqAV3Sd253My8lP2qniC4A7NHJigbkPRoeQMh/Ga2B3YUq48l0fuzdKxeTs32ms
Vs7QRPMeOPgZiS0BGlqfYEvufDHMnXuKe9jkZQ3o9WtDfrPauFzZ4d9PfYYlfRdu
P32PlkmRlevS8yti2eeAeKvqSBvw0IAiye/ZR8jxPWEx6Ph8AVIxYPTDJrWJbhIK
qVzYqJKBymjzraMMn72I72NijPU4wOm0nzB6wMUH7C7+nBzWe2vdYcFOoHwLqQOT
99657iOlx5UaySrfF2aTHWMiMfTQBmeRrT6ZE2Z078zBJwa1gSSnYbSyGPBbqgoT
T10SJq2iBFJV4i/szKFKgkOOMgvmRmHBUslp0XI7DwlB97WOPtS9kHtBnhtbmXp5
07RhEbKZNkzNf1Ykm65U4uX1mFOMbVR0YGOmHB8+chdStm3bC7LPEak1Ga5mhBmv
zSJwaRUifMOzjAa45usC7WpNsRFeREzs3xQrpPXgFAgsKwa+0ZKvK3eZJ0ifZGiU
FKxW22sZpkX4ZLJ+IPmrZVS0+O2Q+LJZd4wVH7/WcEaNBmpV53COvrgPgYZF+ANP
xYKR9cMrGoHalG1Gca53RsDWDeOEJb9oUbgBdlVS1sEyys476TsgLJK4ArSiLNzW
jkZVa/4aPnSOK1GEFp37gAcaH2phf/cbcrI9b2+mZ3BycEXuAnRb1ZWNzExjXr+9
f6zxqIO0DjIKjwJYXl8k5Q3JDSkC25yLJZFQ85oLOtgeGAMRwBcv0GyUNFveo2Ur
NzBxTJS/GvGkrHf/iS02mwiDRhJ/mlyKvQhpwUTWzum/XcgKbYaEIaEq5qAnXwse
+JnGspMUpcB/ZBtV9wBJi8swc40xU3HeYjgWSgvdOZ1IDhXA+WUV94rCJAzFa5jE
kePqu+ujnesckUrIhO30jXpVkYEMWi2c0Bdw6sNz0axEIAb6PmvzccJL7hj0Gifp
hBK5pSxEG4j7mOGa4SJ8xgOk/OOVrS9gs9pLqyQUthta4eQMnRg0dxtTgltamh9Q
5BLfEUIFe8uiDLUaQKIUtHUp884LhzvN2Lg0zHz9I6QA4MQOUXtf1958equnyNwH
VrsgHCgXnCksXFpEGBQye41t9gT8v8yw+Mpil7f95c61Z9+6TfBMaXItm1lHCfl7
bfBDqJJVU3N1d7FZMwvep1eWGDFSjfrS1baanezhbBMDp6Dkm+OBmiO5CVQVwXCv
1LbXEqQBYvVd1HQ0prD51/ZIQYbAKBq9TAt64myiT42/HRy7OFaMvq8CEnUcmwn9
noX09ux7GV8HHhwvVtWQ9Bj7v3H62Qk2V+hmUVAeqblg5oxWzZDZQDzE9f4BT2CW
qrTC6NRBnm26SwpNg5W7fDS0EwJqaVP0eq3uShvwBiQsRSkllqQnPztShG41Duuk
jhaa95tigZj6wD+LNX3jjLD8yIxxydLCGMa82Ebj3oDML2RpOquwoGfRjZ5TgqpM
yQK/HVSdH0SBj+bHeKzL5A8QR+SHXjnISMDqUy0s3yuweUWUpIHd8PdFgTicNCSJ
ovbwzgJekar2b8WalVEfiKY4yYI8tUlqXqN/umqu2hofh22kSFRyH5iProjtXjT0
qAYDbzXQpewTLr94MOHbGse6zccfmmnGDfXNfLhxiybpqqjKnyOLmfidy2kAOR0K
TFz/EwFMm+J3kqFe9oHW4MAK+soNE4j3/W8tO/pQjko1+ABeFNP2USoYi8SdBnam
aVVqNcffaBF3cEPunEgUl8AJ8OzF4aiOE21DKiB5eShRInb1wtojGnCDDTt+Uxlx
iozmX28EQ1wd7ZNmlBRXNwzyU9e05vMqoELXUUdrxFxe912nSxSXOthcaMCzO+ve
wBlyhAtnEVUrdZHd7nmC8G4FrfxP1s73FdPl7n4kepocPDqI6hz6ipQAbucVSU8b
xt4IhJPGPaBC8yPfIGs/KIJLdfOwSF/xLQ1Aw5s5Szvl416F5yhTQytVwCnrWuuc
juRouZ8jlXGoA7XUc5lCl6DevyGBV7zddpHRWszleGAlP3ds7wEdGp1a1ioa9mqu
XbbEd3L4KuQJj+WsH91VzppItkcfk0mbNkX41rndrw/UwHz5l2/maW2d+baGF9Si
J0HQS+PB+ozsol7FA9dqBwwxFHeFY2qPI0yp6PtSHLnEupntWgCb/7/c7t5ReSt8
TmL03GVWivPJM6SufeMQPMcwgGwxfRSDbUlGCMzNyhCS03vb9TZe0T5BY4m3cP9Z
r50cx2o9RjYz4Fas0isqbyYI+2zmRJ0iqViM0+gKAXDesld/s4n6DmrEXmVj4KnH
8MpeUNdxhwVXCKavjdNinmU3Kqf98Kz8Ad112nag8+V2dgxK9unLNOtzYCmtbLfW
Udr66QQ5x+x8zi8rvFnYoyWKXSx5zz5aMNGx+ltXP5LHNYvwbPO6wJIkLf4yIuMh
iTicmpUfpj4XeMCCU0qyu+s+n0cv6zW/zwdIiHHCAFnmXa5k9J54xVqgIFuNmmFg
B77BVrRG9w4LWQE1pZmlD1EsPbzB6S4xp0+oCqZKz7PwyFNxt4/sc60Tne2N8Qaf
qML8bZSQjV4D9Zg54ZJeyuPRp0B7I7S3To2hlbtDqoDlsDytKvsETyRJy49ODTOL
PlXjukPFCpSy2MZgMKJropw15WW4K9ODfopHNHfBloFV6UaoWM/JWkCvpQRKWGR8
6A2GEU1JLVbWSGViPBHwJ8txEmYmrx+sHp3o1oZxvTrhaCgy+Vtje5UYeymy0AIn
H+dScAPi316NK52dCaJqhYEows9sGdX7yzODVFtG9jMHc4VjdmJd7X/KORPgnwb/
0xXYDwwd/cZstulrEUBUmbV/Wl3GDJ5oVOE28SOx9RHEb9Lq3Pzfz48TgHSVEElI
GBxtAji8prygtlbp1l7pW6jz0jGvrynCWUGFPamFnk1zEtNJt+xLs7SDq9Obalym
m3KGwv+HNjqIVj7r10Di2kUF9JUjU28xupOq0wsevLbh8gZekoPd82eACDm4eDM5
SLh/vYYc2fZDIuL3no3OIg0bMsUPTKBEibHQ+A+Q0u+uoBGmaY7irSjgTOJm4nw1
+ndi5WXBolYA4223lzUfjOBivWm/emmqkQqK35332zBSyh5jHR3bBaSf8uzpZa/n
Q2L4DSG0l+5/8VQu6k2WyI0y9zfRVkSfSthnEfeS5DMa37gko31/NybJuNCUn9Ia
ile/sdjPsJGbaB2DHQ2AWSuXyzW93E/Nh1MeHJPBNzuE8Y+MaHGTiSfTKnm9KIEl
rTkBazLL++S11rYSBX+z6GMzwasFVHOeDd5PBDUNhYg5blZXssIKCKAfg2jVao9v
mUi3pJMRxFG2t/D+WOVMZIPWspdwXYGloiCxQOvdcQj4HMabced2e05cCiv+llUy
1GviTxx25XXcyClXFuoEfJr/0fj9J3RcFvQESojR2SRzLs+KoDqML1Cf3eWN4yhP
gL8reck765M8tAQifyYFH9cPourDxfXQBN04//YQsPo5MHFp/XNXA+9I38nd6omh
lA9fxGWd8GrGdhkBptmWigEwt5i/R+PWTjcskDuUDSJkXvpbiQFrqjdxC/tvPWx8
hAmLWy77PrFw03L4kPW1NGZyS8MLgGUY5EX0VjRisduXj3q8r+ftpcQTefFjcNMI
/lJDQL1lZgVyjAc5LF5CZpznCBTgVZYNUGgghrutpFyKgocdIsJQkMR9RCI0joJy
CKAg0PiPfn/t9cXfnpbpuJlTfWK6x8MdcoAtXaxqi5CDIOJpeSS8YS9/bDfpIHYD
nOrl2TyydKsMUVYTclgkV5XFUkOxQdiTjr59ryoJEQyGCypawyQztBjzE30Nh+dQ
TVywo+fYOGb7eOgeP4RuIDN0S4e0KteroHHVKIOeAEA8fVzRjDIHWQ+XazPimjjt
ofwnHV/W/O5jfvMhR3JID+9sH2d9beHnFNRNhY6LSf5efK3/BC/ajPptpE9RLtqr
Skk3c6/OdHQwwZ1/lMR1EnNMm+YQTfZpvpq2qxJNdCxHYnI2r2oWKUCCzAv1ng2E
doIUaQ2m/Gr/V3pSfj4Pc8ZmO6Dk2vj0nBG6APGqGBED2uCS44Ih+NfHLAAVywk+
jT5/9lWNUGMEcEush8UXRQpQWo2AB1rMnT9/aCNPYTdUnvQpKsq0YM2A+fDdUMeW
cMGRaX+uC5DEDbiBNdvp4rxZaZVj/sJfaU0BQqLY4+CfKJB+KqvuwgwgpxljBTD9
P6XlZt0Qo/rIoFezPtqtLfqrDE7bquV99se/R2nCG4i4Q1v+HfS+xro2rF1GyZMD
SwIcAP0WzlDDz7bMtHUMLciygcWlYHFwAvE8fe/z12/sn42vWabMCukP5Gtue4t2
Zx1tZuYdkUy5E0tqbBVjgWiaxF7lmtiEIZIeJxPHcAOpQZ+2ZTABm/L2bImOJJRN
vO85nrusw5/sWE56Z5UfANgzSBl+gU47o6cijwIYADiiYRT1w+gffn8862waLkKm
6JCT1OS3/eybqGLwPjOI7NBRTQpZng4Mg2QrWyNuCMkLnw1J/2cALaMN9Klw3d07
K9su4kZ3hxuPKuHiDNZKujeokW5uHzNgB5XX7MbXDMB/kcBDuvy3zq9sN3+om4Sp
JtUojv2xG1pxA0nygWGIO5cdDZIzGM/YkIEM8bG/Fzo+9On/R2P67FoLDtZMZCOq
LKTjfTr1oeymLEiksVuPM/8c7ek213WmQ431O759VkKd1v8leT1POQsV5Cne2oPM
aTM1NmXvANIHBU6G4DPGRXntsbOZTEA40f5Nc+gyMrKcSvCoRjZM0vv33iesKkfu
oJ86ATywv652L1+xxp7qSTL80r4oknIkruC2ZvRXZIL10rRTkLjBd688qMvGDk58
+qIaQScgMw3fFGj9gtKtrbdhKXxdpj8a7bwkN+D9dvg1sMxbYvVqReQe5ZNfT/GZ
oYU8nzcxP8/61kLMCFvlA9mlACNW3hZ0IWTjRouYwZcD69tCpcRsrdPbk4NARu8K
s16/Xt6VXNqcv3CGivFTK5d1Aq0DtEiSP2O6upUQaN4mj3nqMAUN/eIeu0GkL8+v
1FKUCYYwsDuHATaEysKtmlW00vqCq32BM7wb6MsummB8e8+53+ynqotvFHB+zSvv
G1cMXrnHpbceQPkVuP0dHlULERdvd2i5A4870n2/001EuCY5pfq57PLhyMOkqRrl
4G94oluadcp1jtrPaDPuWvug+XBGTYJf+KvwNr/xr2HQHIkyBPmrw3lONrtPyl9/
xrH8viUo+EA3vdbhS9LhbvoYVYGLUrK7T7ttpiJE/JIjrACfJ4T1ayUnGzg15sCM
nwEPoZ0RPoK0FpAG75pR9k87FjH6pz7CEpqEznUhb+6CSWFBpDbZssh5QLuCC0sC
vrK3sFip2GleaWLd7c35EHPrU20ivkAD25LkJZyx2emQiJdT2ENwE4GQGCvzUxoi
ZnnNHd//ZQZFHeHOSYIY9YWnzIdGV3nHimNSyM5Uo1BctLId/KeK7TtUTNPiNfk1
psE1N+h7B/UnXhbuP1/J6/1FecqrZ9c7LJT62bHg6dAUskaWgbAH9Vd1NEk8x/iC
L//ckl1fMJAgTpsw8TJjoASRARXwlSdNyg8YFvT6aEduN2DvOLUc9YfPRJ8UhSBW
nZZvROZreev7WTSI6huamzOxe1otv7aYXMh1DFPy3WuA0rRgWGYcSMJUgo4s0+sp
3nzXAnfiOgLBoIz2hd26+I7OU9TsZqrlKaoy35+i99SymTRe3KJebMiQzloV90Qb
5Gd+Gte7ZiLmWu8tI3Ak/KFtDLUQbZL6xi6D4ThFWxUohNZG+44qDA4rktnIeiO2
F8rYB8fqjgefijSE226bYHNIsLuB97hMLy058ksc2RlijcaTImzZqu+uAxMp75i+
H+BZVRGOgx9Yo0dKH6okc0uNCGsxi+3aR2GFUN0Lpz/MMEOs3iDo4U2blDmALONn
i6AhGK0/u+7pFicGjCPaQDjj00ZWiQEf0cVGUBB6Ilb2n9GqZYA615pmUtRxrg7U
1ug/y7XpqIABc7h2CkdQRk3/cFVXnCTlcjKJ/yL6A9aEeZeZK15dxY5FCidAUyO8
tluqqWusXhOMuO2mIP2PQ/TP8Diy+PdpZrb8SbSLadIHzFogxj9SlJKTd830dGsW
Wo/7w1TKkP0ouzbMsKnyFz4YE/ylp0H6kT6qdnqfRwX8Umw7l7v9IiBiEhbi48aq
Mr6GKr1ZkA6ImVt8z+DCRzNFJQuGZDgZdzmPYGgceFL4Uj3shqDXa+xbiajQtkjj
oGMdlnPINSK457a4zenmXV4Oi8JUwXsXk+VTVER6LJQxjRcGCPWtDJc9A8keZ48L
aLLoRI2eN+/BJANfveI6zYfsxRCyxOJ5+0lUskAIxv/PpSJROhVBOLrwbbiLWyxW
RQhgn4TCVKdMd4lJamT08vNmtxwGw8dmDA5ocjbGUe1S4wJS0VWtcdQuUkPIBp6c
NQ+VQmurlGjFuxXGLGsi5b6cCrzvYdjfE1kRGcOmJ3DSO73TGTki5e/NRZSGEx+B
TyMxXnHiCBOXj2/GQRCRUbA4kRo+MavtGJBJ0FYPR1gD1qwwwA0ulIb4S2XpFrCc
ri8wT4qutnRoPhxsCRD9o2ojEKARhqRfrPVrtb27JHh/HEGSdDQvEPLwYLcbh4SJ
mOOVqI6Swk1A+CNfnejzULvyHj8o4Nm9QbsOB3y6ucssxPk6OoOTATH2NfWZYXpm
YvrrOiaW4wAMqICNbruuqo4TgKm0f+LctSLDg6O550jlQJgSjtPHHqZN27JGrZq1
BJMzzxTj7NOSynXHMneNXsBxniV9knZ1IxM83TqXNh9bzRkw3r9wahtPQjQTxras
qxZBBkMrm9sj3K4P0H7vNCSIto+//QdGb/LMev/xLcgdqoDrWsRopEjiIIsEwJnC
7JIMALcHJJkQv/m1IrgwrE4uoxKQh8+ICkpeFOiAyWJbb37DHZwjYuXuF4sK+3JR
knpNUYSsW6qoLWla93N507I6uPtm34QvWK2MNW/FVfE91TblINa1dtNZXHhx7Z63
sgKe4mKKRgTxZI3RiRUJtrwShbp+9NLbt14ZeHP9UG0CxhSZIT1k1b1sDtcghJwY
LwUYwMv0/SqVP6/VStlB7hkRrW4Dfc0TiTCe2O6FqGim1q+hnENKngtmMo6+ZQNb
FcLT+86Yz+rRTdXEafh+DfD+wMc6ba7c2Jb2H70ZJtdyTWXF8y4vLTkMCbwfbN2G
HYvN+Z1R9gKD10hWd2ek/GDLkIXnl4qOcvgtH1XZJBbHdH115Nr3olVf9ntPh++c
aEeMnpksGcB+DGyRuHUVSDcCEH1zdF0XUV3U9C8DzSlzC9qEF8WLlw7F3Eyd3Tnf
ke7fU2z7QG4qKUGEFThy4+zr1dNb9WHRoi3g0ICvlHV1c9igqMy5IcyPeT4BRB+w
dOyVQ6pq3D3XI12tsXJQ7VO+aS1S7+mXnLZ51vWMh8fjRzXJ3GfYIsa7EmCz2aBF
d0vm/Lht2oHdhaVZx4Kg8uVu2szXq8yktpDIJ3SJfKEJTnhy6zKIb3j4pM1EZQb4
Sts5OSGAgdoOs0h0hmgzlxzCCUb+4VdPzYF06ef4UaXUYw7JPu9accgTsscmEewX
iuSIa8SSe9B/78gOSgPtvmcpq5Q/zOFGCdZnA7HUrcFxJ+QWWZetSts/6Wy9AExS
m0wVg24EMVPkCwlIVBR/Kl4AykjdZpHsUVZ17cRGzq52eKnsrBsYpv3D2zVocX2Q
6kn4+Yfo001Dkbx7JcNjOmWTSOe1l+cFGmL4Xs8XdWPB1OLG4ud1I6w1HU5+WSSe
0qCBGaWdPYR4AhuX+OEYUv4XQj7HRvwP4CoGptdV20xxXyFE4QuEo8wUge5UA9Uf
4riNE6vZCsG2UkWfiV7CjA6nG0zDkURwZq2xD2LxAREnRG4/pI0SLzt0sHpXjLtT
E70dna2/stM4Lx9hFRtcswSy72fyHimz49QBb/1ay7RcN9fKMLiNpLqj4kzb7Rjt
Ex0mvKG3wHGG3pCqWnWxk1dCellBry5xJ9U8VmoenY7yW5aATuWYeAB0kjt/mn7k
PP0/Rh+RUIx6OdeoH8TXrznof8aF984wh72zxhKewNX3iGkmTy/7PRJmiEZpbQP+
ROl1MkWnXdp6EFTFvqT8Fy7zWRBHBanolKE5j9SfSR6lqPy6IN/ZZ5UScrBM56BO
363vwPAIaa2pPzhSKIs/rxkUe4Am3sQhMjdzT3+vy4Y3yeEKXuyMAsLx3jnmcLy4
xd5WPU/JjG6V37L/rpPCyUdXnRtunUMwTxohYF6eKVmwNea6NCtxC1EoAk+N6SZE
aV06uRPqbwOKoZ9LHPfnkdQQ50UELWezpu9ADjljuDra9c4AKu6CenSUMi+t1AfF
LtzD5fjjgnpqoBBzWiZWRdjqnVIyBvx/szpj0ryw0D9eQfPiuQ2YLBFlh16R8Yap
6+2Wt7d8Yk20qSSnjWbs1U5UdPACpQMX09JgwYHDlH9DX2tEeCAOgkkJnUb/nJ9Y
pWFxnHt8tziAs3n7D6jR2Mwu7ZqrnGFXwyuVBR7xY5sExFInrpLml0/Hgcqt5zSU
csYkKjzszj2n+GWHkpZASsV8I+Dz713TA6VMU14rRd4+vx/13UWPKx1SbVUoqafu
uOrvzFN9BSNGn2ppgNnxiYU2MuayXmXMvCnm52kHSFySMOTzw5vvbKrzgl8VKSx0
mgPVh3OZibCZklxaDiUXzJPQb99884fzTiEBAp4zNbla+kjwKIfPTiHsQ61F1+HJ
SmG+b43UA/l0d11C1P1GLvAqePPglej6hYI35s3bjxkr/bBk3Hom87ubUDPf0jqH
QvmXpjbsYXkq9AdGbbmzZxCxUMnqUMfbZaIV4AepKmN4KzRo3Sv0K3rtis09ktT3
S7bI+I7qklgsitZgEjoqGi19iV7J1u89mItl0pFjkGHBnJZL6KYoK1Voy4UzT4Zx
7kBjkayhWE4+gzrTWbgLCUey6JK98KZfXjoCWjntXOWhXapSPDsOrZKK8tEbZSrk
bbng12pulwfwJaszRML+0tnOzh+u2wPrfYRUvCUhly0CSi7IpD9j0uca4y2fzDC9
fXu95BHXK+++8sZHac9cPJn2TwEJ4DBbk9s9jdlcQ08kJYJP2eC5XUqeBsZSGPAG
aFE6FXpIFP56h/nJYbNaGDzY1Qn4H1WOutvMMbZdfcSzpVFF2onpkBi3E/WVkntn
FlkSdr41MJwqA9VVu28cwYXDkZQG0QqlII3eAQIl9G2OwFqPfVceBFejr4VlblzP
dPkc6aZZPkp6AKeWwM+zlFJmVs1oTy7rYW/qGAXS1UtKmI7VA1GYIcH2H9iOVy2m
oC7F7B/brjZ8ThTG2ZqCQlLqlm/yaM73IZDfCd1HqomHY8omlWY38teExFuo85sB
Qw7n3bT5nmivrPBhsul8wsdH0p+Y2j+Pt00aWFdCxY/tlmiFKKcg5jOS/bcd9Pnv
JNA1pAhSVwmKh/lBwlIrxkQFYF0QPDcl5yCUS6ntUGl0ZNI2WjhtJ/Nv5fyP8ljz
2PMfRkSEJbmhhUVazbndjVG/sEdZx7Jc84gRejIalcBt8xE9r+mKU+ZEMyuS8htK
XLTLP9eTksQdMCU5edpJgBaKh3OuAtniJBxiVBuoz6YKT4nM920YsBVvLxsCY43f
YiVR7E3pG31M6p939CtsRvY0AYMdX2UDlEGGwqv4AQOhr274Wyndbv5+RwmIOT0x
HSRvS5uPy1tFduuzvWy8vkNopX4LFaC5zL1qXxCI6BLnCemNRrf/iunI5VvEXFxu
cOgQI5MwsDAuoTucG0Uzkfi05Y8+Yk/Fw3CYCM2PHq8Du3yso9/uc2v1AOjNYCQ3
91k1rLTsnt+tFU9BPSPvT8mkKPP4k2IwoN1YJ8xIRSopsU/D7SOarpcdyO/zu4Yf
KUO048SiYGL/6SlhZ7fsgMC47KjMR8huCEsXOzdiQk3S+EDGzLFiscq4ySGHqila
ms+hdYzhRfaQogTqYDu9N+WeqyRRaQyKWiSGoQ6tbdU7h9bSh9aeOMD9qeRDDUtl
yO4zlXlRVSQhSWOfxTRD/Qcuuo6NxkZFKaVZ7u9+GQjs+kArVPn/KMhZGOx2ns2B
v5vQ12MNQUHDYtgB4JyP+jyKhD4RfTiSOZutAyrGh0og1NghuMlO3naKyyNeMHLg
/VG/t8jgdhL/pv+PxdqCXK4c7lDssZtxAXpyBxsF5lU5bKsH6SSRQV0Vve72QQzy
E7YiMx7KX5fbjBHJlRuidPJaNDxMKog/knCNY0ZVSh244qCHTclnQjEdoU9DWahj
VFkzBc7bhWpPTW0GQ5I4kFBVIOSJK/xAfiEj9PpeVsOWEUucqwAz51Ufnp8kvng9
r45zjaZRQCfJVR6uA4YjVetAxHW055wBQ6vApwqAf4OaffCeVJy8OUAda477cwrd
RZJfdZGh6QY8+7fq3l7JqfjbQBA3XGoT1hqDcs2DgnhMzCWNtcVCh0XuTOTAaZOc
P2ZPmhvEWhnyW6XJsE9TMm64eWW0aDNoUE3i2j4Uk2AssQExYPclDEurcLFtIknx
4KCwUUyou85V/u5wNTlLdRTC9yQJZfmov4zbMCberhdkxYozxNodIFjnYa0xaA+n
P7nd4zu5vflmb8RIVmo2SoZjrs3gg3VlRKJM0RjbDaINqhm4odTSClJgCsgV826g
Y+kf8MPHMfeuj/uQpijDAxIJ+Hykuu5WdmX3UOJoMxWNfsNBNk73LQt/OPJxqhHe
8HQcX/Cu2D697CQUdC5B0fIfqx7SqMIeDBr13mUf6dxF6bo980bDITffMtxZ51Ag
mjg8IiP7c/o03MqVonxaprUKFKFF+JADF5kUSOOvhUi8JsEMhQc9ULyNK+6mx2ui
kpPduskKOqJu0CcZrWv8OOOGEpvKPA5v/e+0u0SxkTu5SqaTDbPJHAOgvH1Th+8b
z+G6o+nyX0K8UfMQQDw84yXPTIe1mwxoa22XR0OcBImJjXkg+E+qDe/7+oBftnER
fGMsdmJOzf80pS3bIx1n8zGBldJ2NGI/IbvAGdBlBecIR2RKvYA8zKQpePjcI1e+
Xahj0YInnc6ETtCPtbrJ39+zTVW1KkN3TCzzIwwnAvUaIFAHIivky73+Q/swpHGE
CqiVVgPQNvf538REobAY0FdFbZWA9g7UGl49g0GG3QubDXLsYDS2cnbUh4WuWhdG
IK6rQxdeUmGlcF7lZvOJrCh/fOhbw0ui8+xxI/ViqqCpdzATCxPIL4+0JKFakX4J
Gs+yRugo+VfAMSQrRf+I6WYpXFR9s3FDferiBCl1NiEbZUPv4Tk+sh/Mw7JYCCQb
ugQQVhRPeTydeuFm3nCESedKqtnFgkgENkuqjPl01M8EexPHhvt+71EQ6O2nzKPS
FilQ87htCidPbIFKYb33JqCP2zfc66pI+LO4AMrNBdnUZ6HIGv6RSNZAYQbig+7b
k/8r4CxrTFNFwrycG7Tmt2yvNd5Jr9EPZwK7/mlju28Z+c9N5D4QWAAigKw0HltN
D4OQcWvH3RtoqVxz5FzKkYhW7clK32MtEs0/dfhGZzYwrG+EMlM85H4TLnCvIxc0
lmZZM7Fpcz8XFtO+eLfqvJ94HsJLp7lScpexsm5vBP6b1VYEotG1oprf12UnExkf
lvZi9YTEX5TiL8ol5SXZT3vK6pHQpr6SSLcymQPRx0YNqd1P1Z0k15N3pL+1mpVI
3y+C/BJVsDS5oAjFJ6Bf1UCh2ooiGvCwKksAjyuiMVHf8Vgk6YsabqvDNjpbQcgy
5qUdt9BboTgWVvJYnfsE/13PCRYG1ulTS3UHJplJbDUhUD3w3MUBKhguBhnGdA6d
RcIfEzot8JjzR68nGFdzQL+D2xTRcCqWOdumDkETYcRhdgQ+PqcyqnCdkmdqdiag
cSCHy2IYao3l5EmDzLgdH9cl+me/VMSvzb49YUtPpbyWC5tmxbXI0NcCLagAo+RW
QlQTjucR6JLxHch+8xXLR1/OXV3C67N/KiKXbrdw3IXVn95jtyaB+VV6Qt62LrgI
ODF8cKl4vrmT6E1UP8N8shtDuQDYNi9ZgEq65WGy8jFM+xSIF/FQU7FtuBNgo5aO
fH0LCOxEd3o6eUpoerCSbfybUeF+20kuBf+IeI5f1xcW2mMb0Ic5+84LgYWd4F/r
Ir1wnERA0nBCzsXtEi+gitAUu4FxC8KIl2FI1u5ECsdwj4sAXKEh9iD6Cx1QeZm6
Spp1il5Z8e6tOBZBTJvieK9w9T97kuNlNe865p+UIq3bACccZoceORoNZaG+GtRa
62hc+8Xc0ryzH8ASFW06/HHpudZSxeHLarA3W7hwRaPGPb7BvaM2MN3rQuu8fuCg
Hwm+260gVqzpSpAqzXcHRrtSOBOOPjbP2MwwpQy0S9GlCv4p0f75PIKt9ZUZnENk
9uxF3geoKnSiKnJBRS7tOFjEpXg/abjS1nv2UOzIue2GSkUTchUPyNF82fcxC7/u
XEOuQB/2QW7OLS091ycHzxU+o9CdygA3H5kPcNH96tD9kt4lKG6cCU0e7qb1gF7a
JFL1kZNFqtJHpVCb2BUKs2pCJq3u/jLNTdSICVVmqUPqKwRx58hrKsjVVQsYG+kS
EbPjYuPUmN7yjSHtD2G9n+L/+bt4wa2bXaRPMGRqpIiNQC8b16w+DTZnnd1H0/A9
gusyq8qdbuc8Sn87a+zyfpjk6ej1zELtf9GRAPiRxRTOy3fxUdpmdOc0OnO8h+Sc
fKkGffnnCGwN/l0WuK9bjaXBtglwtOXyUAYqGXJ5b3xOoJB32vBQ5ZXIiqc5hIvh
ZS56RJp+vGGD+B1bc7iszqDfIXuZWy0aaHezlHjMNYB/4qepRkUNDszy/+WWXqHR
dEJRIfOaPTFU8UD6KVbqRP4/uqP3rX+FudvLGqt9qUZ56ufEHrywyy0qAVRmZpR6
5u0AJr6tN5RFelsC2fn5LsvxeRPTzsrQ/a8dlNvYxcgFbaVDE1q5rfyqRmvDo6lu
Gm+TZTsQcMzIZDOCKw3SlnNlcpieem/STsiGOL4Q61elP12L58k0hUv817vX5oEA
GG92xR9Hn/lFnTrdADUZbKMfT1bfWJVGlCJ+taYgxHxf6xQATqF4TzWgXvrjkjF6
t9edmvXivJTVKUF30LmmcxyoaY1FQDvw5Z7i82k7CfQXUCa4ABpncYkcRiws5JXO
KKhITxGv7qEgEGlzkYwTjiWihc0qych8/E4oJBjVIvx8PMqddBEj+qJHee/uJza9
dRbO7Bb733hve7ohJif5pmbUXiEMW7ZfCyUZ5altrs7gm48R1JuGd9cKWP6Kt6Ur
Or98ASDC/KG1sLiNkvCfUh6WHL/n/4NFBqBCyK8IpOoLVilZoAQ73phdsngjUEUW
5Y1uoXvtwcptU0y9niesPs21hfX4J9rQvct2UnlTsVvr4cm7MZ1vPtQ9+7Yau8rQ
+ge3LkeHwFZv+jlZlT74tqQSVuxNyEVgUnuEEh2+93wjk3eJU087EmWWm+31jd/b
RABpu/e1pTuy3ivZ5cvZAo6/ilxsRfNbo57yaKJaXW2d+6uUCfbDtpvNZFBG30au
F/ClR4aNDdYFOxpY2/mUJ6M/DqN0pioShxL5N51aFE5f5tNbmrZzY6oc5HVLv22l
aBin+JqOijtX+JD1mnTxRXVwT3v8NZseCL6+dgFjF5ed3VTr0fkeLN6nJvf0GddI
rkigKq8FhY42X+ytomM2qw+f/a9MQf54ms+Ii/htRabniiLk4h9UW948ziKVNEdr
kfz11tJGXdxrPSD9M6+OaPsN/+kLw0NdRr2MjGOFx6KzvNvykNYH77DWJ3Oq+lGp
fTZEHwtiDm/0De+VwBR/z3jk8kT3ObQv4eGwW0JJV9C3CV16v+JHrrKwMjCDH47x
cYXxhLJ8TCVkEnUq0BRZg8NuH1T4jytJC+U7whiMDkTrZpHoTe8tBHaZVHqM7Smm
AQE46Bs2DTkEDE4jkjsPYZmieb8eu68s1PTNJAVd+3toS4YBBjktt2agnnKxf81G
AmMkuleqmP4NrAUZBHVxlhgEwnSpeHqfK+iYvZ/vJ0PdMauBycjn4neuqQxWNTWE
3TVe7++BvbfYiU8F6Rh7RZCqRXFV1+psIl/xfTRH+M6/aY9ESRfMI17bw3sTaPKO
34UOP47MVClmqaPcpNlv6gE74sqgot0+fu97uiLy6iwdhcRqH/bEzcjXZHdLYg9U
cpBKnmbKDi0SoVr9P2odEC2MZkpPAVC74/DHfX67kYyPdbO7w/saV6SSw5O6PR9x
BDgvh6T7+YmpPLxnjfzOeQJ4yd/7Y3B5EMIQkuyclNJRY3XawDf5PMYKx/qU88qM
UBqEfGyJRbpnPTJQqCRR/mOrljEBc5fb6UrDilxuV4c9de9PPvRxCjEJShM8K9fj
8fIGOVf4ly7qgSftGw6cMnn1wVWElZTLCHvDdiGXna7vsdlc2JNDWVP8hT343FTS
2s4rj+Ko49LlO5XSbOilcE1tVXGgfrcQVGX/2KMj2XcJGfCSqzgq0hgH5hwQAO7E
E3rd258IK5b0pX1GZffSIRfmjI0SJJEdRSm7xavJN6YLk9fy0eHCXWgywDlq6CEk
XT9eCn2sLAdd1Ygckp38AsLaiAjQOkhTqmk5mrvdPSE8TbfYgitlAm388V6Ir3q1
wb4GBc0KcGMz0lOo177oEhehjlKmBl1+ITXlHA/uLdNIKqsaZp9ZHsSE26eWrwC9
f/WYw9TngJ09njsxEMGCqM5lUf3BkqkAXa1vGUJQIH5bV/APLAzolkdanVINxwep
9zmLk2vyLGVgn7xPmw34x4cM0xKfBNemPQddyGkUr6Xe14osd0a/AkM7T7HXlsXx
Q5AbbWKGVQkNDwQ4903h2aD5PyFl7vBfW3GrRuyvRGQvd3j02FXFMg2XKfYTPG2P
oh8mZmg/gPeo6phoi7SI1dgNcSBe3KZtTmALJjb+EXuoeh86eKbllJwi64R+WbU6
BiTuF3k99FzoBSOkTYMQW7kIdly8+21OlhK68SkKn0o/2BI8UlywKgb61yS8E0Dm
BraesSEvCNiwsgaaZ3comIvCTQFCiACtJpzPSRRmhTJEVTaY2LF2JqcyrJ2+3RRe
YToITIemPOnQcP0Texmk2bc5penxQX6/vy8uOxvPnolVJejZaBThZp+S6WpP7Gbn
illnpaHxcQHrm7Wte9Eq1yyeamTOgjgQGp+LMW+RZzjAwYiYYLNhAS78xrwR9DRW
XkZs2aNjGQnQV0NgYy8Jv/sm+yywIfc2fRTHtbw+a1xzjRVtSyFmLpqLDcxXl8lE
S3QItpdPB7iIKtHnblFciATRhG4fyBaoVheaiRhyVSnmeaAqGw/rjFKPRlliCNn1
vFK1943DuBOQVu9nWEjPnxTTtGC63eUV36ljsmrvOkyadKvKwlJ4v+eaCru//Op4
6mo4mSuLX/bzsflghrfA3UrePY+MUlOSIFBS/8pPvXgLY0Ar6E5UQsy7nV+PaPA3
SUCFof6RQDivaxZznxV2a2gszr0IQkKySoX3FjkxscFKRlDth5TTjnlqNlTCfVbl
W54A6I6hP3RxW3A8mT8nBYHcg3hmz4zm4vL1EB0dECekkQO8i8hkqgFUFYvrMAAx
GS6EAEL2ZnoIJs7GhcPwraALR8HJG2RZ5k1DWRVRkixmMzgHq8QJo8BlzltzDWYT
7OubdApy6tDoB+NF406zAvZsIJuQ4haDeTvVl2zlJ3vEUFqIVy4VIWnBRnQkrkCi
jxKTPXeTCU0HTPUJu6ZEiVJU1BS4qTeUrWCf6HMELyz17KYhpZWE1IzEbncIJBlu
3PBVERtET9AX8igwRY7FeIzPs5PHovBPJkGj5Pzq+wlREmMgABwSigoyMwxbDCqV
EpFTtEQNdqRb8sZwDRm7r/uUtHtMLjoAbGeqP9YZv+Rny9AhDBJNOJ5H0Uo0dZuX
zkaOA4Hrp76Ob7IUS2Va7TiwyPCTFyoQ+NFqts6NdWhgUhPHQDhWHSYEFBLaojHW
iAoDf4AYoh8KPkj83cpmBDaekGuDpYKTAuVS4p3lmkDXi/wdfauaxBnaf6+tG2WK
AbcUK5mfFLmgWOVWNJT7RWpMDBbg0yM21L8jsvrMuBeIzn3EGLRjOZBHILhG7oKU
Vl7ywIyq+wpxaJ9WMfIl6kFYuW7TxJYPKc4UskKmNhPrZVFTd1e7Owd1DOAOVSep
A6Zl3UXxHEbaFzMT7AsO6U+BD8b7eK/dYZLLcHG7xxFe1hn63tMEvwkmtuFe80TY
z+UXB9V81VUvj4I7dUBkxSBZ1rSDod/lZAdx+H5tGyfXVvIN81jbVaO+2MkccxEo
ml5wiEE6MGqvZGdXk+4xTk1V76tphszJ3/DBuJAv4kEJUl+rWGIUro1i35fK0bmC
ptbpZwuogBvkod01iTUBJ3qmTJWF7jqnhS04QFChky08sqPuHufkU+Ugnf4Zf6zK
1RjwB07lYYrFu6WqvbCawoIudfP5WyGfvPjlhwi25rv6be2WT3Taq0NkdXsqjK5u
oDLIX7vB3++n9tweIwywd+D4Mhefchl5Sgqp5bkKwAltyc/pJPi9eQOie0uv50ti
124vg4XiJnRf7FF6EGEltIaDHzYgkX8FtW40ArjcDmXEtyNwtx77kYn7ij3WHaz/
IgF/AQ1wThbHLltvpvkivMGjnK2yf5a3/ET7hDpHh4ZqPgPDqFZc099qt7u5pDvZ
NymqMb1ftBq+WjKPefRPnRz9B0Nm9K6CMjK86EzKREb5HONl7Ce0EK1BWTbqgxVz
l9QNcVUAmwr6EYiB2x2S39faX0AiNRktABtWNU9GmTHToh9tZv3YiWMQgQWfEKtq
u6jyIJE7BBAderNQtVpM4erBRgIvNoFyirZ02HYIzoCYpr5aD4OiNX9nW02tTDwG
ceIIr6yXf65nl3r/DxMB2+xtVGjCISYq6Fdcmdqrp0+r5y8uheW9MDHuLFVNuRdc
qhxL5bH+y782/7PaNNuBWz/x8a1gSRxzYY7UTIsehf9vIk8TJh7gv5v1yMcs5WIc
W2lgegj0i8J2Tw3P73BDN4GCS1WUvfl1DBd+4eYLRbxvZOhJdK0G63sNCGWoL2j9
+jd7rfNV9616i5t36WGeJHn2+tr0udL3O1yHpXv+66HgpTgjnAaXpF8D6qDSim5y
C8vDBXA+9NroC0cgXmdGQd4ml7CW4AGwSXQa4NS+H5WctKpZU7FyR4K5na1TYeP+
44CDAsTE5FhrXSyGIfr/34f8pfLR69pi2ZkzV6pcw9X/q1BH2ewmmuSI8JazMHR0
iqKj3Y5HD3r6kTSGVyogglXWakFmyBGNB5XotCdNBoYWAp9ZOV74rW5TDH7AE6G8
PYTCFnoiW+fUfHUzXWaDBjegmP6c9ZH5/kF+spagZcuECKONqwV8r7h+eFcJGAwk
MHH53LdCC1Xj5Onr+Y6/r7/AdyxKYUZTL99AWSBNatOh7clJWKpXpOz8K0SMskwF
6ONDTOU8wZu1MTOLNWJZoX/Ha5vd8IidafLqrpeZvb09NzkHLCt00nbysX7zenRZ
Jdyc1z00uKw5TVeSuh2GpU0p4/KGq3hL9ARpAtkpkYuuU/1n1Hj/VsHP1BAGEpXB
q0qUuMzKyAyFk3aj8phSr+k+zB43HCoDVVOpSvYikVcMVKI5UtzQYf0/ZKBhzbtF
YLIrKJw0Rx1EujAcIpksRkapoVB7ym48P1fgq+amnOCYHOabGMphAb+pnLSjgq4U
aM1bW94TfygQguPIbBLysMVV4XIp+ynM9Gg/RdkI3X+1s82JpaJ9OTJ1ZTQPWAD4
p3LWPxY0SlRyweKSpZkIsPDWPz5xSieSNI5InvX+GZ4E5YvN4HqcCLCO081yWtR6
X9nIIshD9YlUuuHD0+jYvF9ISsjO2s/nu8QsYCphEONFrifp/KV4cdWhIvkrw4lw
VfkcrWrmW6eUI1FTKG9mfXm1Cq5WaGcFEPSP8fwOkxG+CxQ5Y1BA37f6V8vYMD09
vJYjhaE2UtKfXwZbjqciv7mMtOM8SG3tM7CkbC4A0pgUJI28b+TgbM9lr5Tl5OLN
ccUAGsciPu1Romg9gcYLsCeAZkY8XFpYlT2qsCeU9fK91X7r734tvTVLaMMa4PKK
JZ8O+IyIQo0a1reGQbGxcMqKHjw/FvHq9WBx9I39zkh1LHEWzZO2xafgak68JCoR
8swcp+E+S2jbv8h6P3LWO/eZIghsrqBbaxFSWIQnvSfsAhD0zzMi6Yu7rClUMn4u
qVzZM2at3j5waZKUobSmXMsWk8pcWqjje8dQl5b+HlNKq5csIfpcfvhLWZMTBN0H
MQqT1c5dXwY6hvP1KZMmVx98hx4/1v3DHJy5GOruxrrboz7eg+jETZCRZL0tF6CG
qcEYzK5Ef2WSFhgVYTCBzo9Z0SOnD2m/uylsmDDI0H2W/jb/LwOTV4xwvS4MaXRb
/T7W2h5AXCYPL7yTUnQuVNTF/60eWq676hcozzUPNm3b012WBGhdpm0Gi4FS+8h+
HYX2FHFm8Qw6aSxqZHVPGsozpccB+R+kK4M9Hx7Qgern617GLkirXdfWdOOxOhRa
s0U/W4z7A4BikO8qjgPXnFh+mMGeHhlLx5PDMEVsnlhJNcMQzqFFKy89t0U/s98i
ll093T48EIgssujGujzNMs0DbnoVa/9iwlLTamj4NrUUkRorVPQe6u5pS7BCLR1b
ARQbNpYJppkr3E988aMwCWUfEEbXl6DHLy+puRpkf04lKB8JcmyY5HoyUVJVbUX3
3Rmr4SRcXvj8HTznWPH4W8oNcfhDxNN8HYi8HMQ6O10K3AiAp1rNZhGtv97svWVQ
GRNl4JMa6/SPxtqH5xCZ0sGxUD2e+ZVIzWZTrg1eJ0Xz3FoVWPESLJ7iTd+xkmeq
ktc60HmISjvV5wFbFgdZP7O+1WIP/n7Ndfgx2zE8SFEcPBXWGbxmHFvCCkdTdEgI
pBiPYdczecwmO8rld3tuFJxe948hh6l2bW7JC8HvyTpqNZVSgh1JbfhQSnqBGel/
ymfB5WFFa6JZFAMmu5oKFLPwbLsqC1zkcF5UA3eRXNh37/au1wqFVr2rzFode64e
gmPTKfHa+GT4X1CuHHp8Tgv6BVNzm7/+BsANLNmfJXzpXyvQ/zeZT5A/sZe2XcpJ
nxXjEPZPBComV4b1rDtaK22JWAifDF+rX2ofslTRTSsDYp+qkpbYGIvPJ6I4pwyO
ztpNRhlaVV32dkdD9uNf8LNabGYVYVmEbj4d6CE6zYxyiSo906Wv7SG16+H4usIN
NaH1nYUHNeCMx/9+Hk5QxprRjUlsYixDSmll5wOPO1wZyUmpl+3egIGZLB7iMy60
e4CxZC8WC+MGlPNYwGrL4NvJyN8/PF8aBiFs8OIdxPFbF+fBeWc8gwV+EmCbXof2
8os6zfQQtLj9ehA7HHW5z1FsIpGBSj8VNu1kZyXfcxD700+h9YfOHT+1PXUC7BvR
GHVnLZ1a99KtTK8cPOfjPuujH7U/rKWL+/SEJkjDEyxhzqWqP92bsdsJ4Be739YF
Xw3BJhBRkgSWFE+H2ZmZRZlxfKwmlWhudWDNIu0ZEVQcOzLZdUCkGDZYigMi1Ed+
C23OBzCOd8LriBwZuwzPB8O/HKpxZD1fdAvuB8eameuI1Qjxvtx4EPKmgle9/RKy
5/8dJDMaySHQMDX5Sis2To69h65F3bxCMnBAwkkd73WWumKcTg79ebK5BHIjOs6K
5k1Uh3w8iHE1BQjOY0LG773FmoyVG+V1jzRdzz7I5tDcAT2k8tSxb6sXiXfr2xK5
OU3VV4MnkT8xGdME+3P65RkynrfkVSnzhgOr5xbR5CF16CO6yHPOG56Du8k3Agu/
/D1bCsyvVE/hu4Z6vkE2XSN9bG7ZJ/zarY1LSDEZ/HnNgB2bpztHWVIXYas6DIxd
zIf6aKI7T7TTZ1n9InZSjY93zIb9dwJLai1fT6b3tEmf1DuOD68+F3pv2QDPChHJ
idzwv35yAK+tyUj8RVXVEUclB+PmFCfUDdVvaI9AHJQ+Q9PkrJeE+t9umBOKVlV0
sddjzsCRZaV68ZF0bVbqhq4FsOzhvPpTVxdVg53jJmYTjvfN3mekjsoztpMSqikm
dhXeyZ3RhRbX7QOM1s7WFutzAJPJ6CXVybNAf1csmGBFa94V6Xd8N/IvEoPjK6Le
rEg3WFpAzD4fjw8TqyVzUAcu5M4mvhwzUalUPwisaRwJf9uZehqCJv9PymMMYqYB
ajnTlOL8OHcnjum6QDC86hGLg6Gj5maoO1xHrr3ERDjmIzrSFqRmsNdhJTOrzZ9t
yzVHvyuTDOC3JcV3OLYLXJ+7NeMtCofadtc1qF//uPqIOTh7ON44KfMl4hHh1QaE
lfkakcbrYqurAQN8T583TzuI2sPB0EYlgaXeKheYUPwnb4XgX9iTHN70vWfrJriZ
p1UKyS9+ZgWX+/GteZmA+Tkumxdj75qMr9aqNfUZGLyhvNVtwIRMz1foUEfbDNrv
jan/v2q72OVhVJXOCSXoewZmECreg7fkBddxYiCKVYOKCkD5AWLwqw4HpVQ5SeI4
ey5vM1OUwJBSOepM1I2yJgkllKLrtL4qPylHIoxKjhSW7blUKGrgbDfmC9haMFr2
CNrGW/13QDx5yoGHfwCexP6CC+CM8/SVhB0Jlie/AX1AXNJ73DtmJ/j3iQwh6RFz
DvSr6eLcU+1xbnMndTZzoEqJV4voDXGUnclrEJreNJf3k1sMWVpEekJxp2ohCOB4
IO7UnI8+yGal7WLWKVBRXQPofFaRrbSPbTW6RLRKohmAfaijb6i6Iba0Liy+HVtp
l/yUCLIz9orRrTIwBJqUs0BreRJHKvSsspETgyuxuyoWKSEVxsupcH+QP473ZnZ3
nhwnx0hF70lBr1ROUuuUe9lZnI2dudKZ/ffJNmhXyBUL+zq7/EXSnbfGX2vgy4Da
Zk74bzvqLAkBYYXkzkXIhxAUcane54pmEJPi/b0TbRxiyD3Ch0gl2FtC/ZKxtnyH
44K8FzKK0/xfhlsbq4gkrQgLjCaiYfilOG0DH8eiOsZxvfeSr4raR7OW3aVOQN5s
bfvjXFjBtjZ+dO8Khdxs79rlhubWhKg5ajb3+T9auEfuE8l5+MNzHtgSesB8p6f3
cngxwwY2FMAKVL53oBLYpGfTyO8Fuv8AT16/dV+05zGaKsLwozFvBUWRJ3YKYDiQ
vzOYMuHzjlsM4WGHMksnxdXo9PJTlESJ/SQLoX+MSMrXUZM5KTMb7eOGazRSnvtI
3CR2gpDEZLLha4abWubnLhiRBO9bvpcPSoAKunYhGYxg0F11eCYHEc6Wq3KuQ4Mn
dPxc+uT/b3fYVjINIyXez++LgdIMtaz8GaqvEAdC2y+tU9rpRtJHuuBeJc3zM/OQ
4SmxwrgtV2hVDfrD2G9I+/lmxh9wKn2EDwPvXJ9MsAZfvDl1Wcxozicp/dkupkWy
8v67CPeII3BESPmICi7KX7c/KsoOYtDf6ihFU6EAD0X8s8I3oyNzqv25iAscZ1PI
2nUbLFoGyrIeCN5kX30cYg6q1NGk3DPe6AUNA4mMakO9a+EOUho1QO0MO64GrkYS
AWTiQSfFZumLX4OnTYYeagJqORDWt/9n9nWwfBVdtwCSWkfkyU5y7KxIrul2s6Qv
lDS1CekRhRVX3KyuKlJqDj2Vl5XcOiaI7JY+DAdz/r6MIcAM7WAbYbuPMmkuCg5Q
Y3rqNW99xImOZXdhr7G+xBo9cNtDAaifTZMliK3G1p/DdLJCwDCfpFtldV+3BQ6n
QUAK5YMMPrd5CPB99Vbr6aqjjEB96hZvwG2vtR29H2cNz+FP0nKTJOUCJSTYUKS1
xLxFuMKvYO+2cke8lvEenW0v9//cc5PcJHODXDOolUpgfMusKlqxE9qJpeYPhrWp
3UGuoABZuV7v2gXH5kkjVq7/GNV3RoP6K/sHIoFoCe1pij30xmJl3YOGcqgbeQDP
i5WMzYKZFZ4Cgbm0f/mYplivBQymqn8GEbl/b9f2MTYCoVrs7vQpI78cXNKjuIxg
/xWrZtgU01iBLtBm86dZRYi+5HtAIRaKM+S8geU6lAkwypIA0+B3pRwOmJa+ajZz
TbgAH0SL3NMMkrFYNXualisQcNzUQmmHYbnkXagtcD+Gq2QZ195z1n/VujXa2UnA
4dFGjly73y76W6RvFBZ7xPImeJwCJtSmdNrssrKiiDzy61UQDSP5Ltf4Wj1OB0nH
keV47+yiQ9tZiBvQ7Uqzp4Vc7QjmaugMbFC1YW45Ls40zCM44sQZGX0kiBCsEvr9
HRdzcflCBI4NziShTtPZ83fzEFLDc8TJS6z1DKgRyrRLU0VgjiRHuILeEoM6QHgH
+/LkbDUIK7VOZXd/3Vn40YBaTJpvUkYtgAFvpZlX6T2WXZZy0jzZnmG2vCX5N+tp
/P8w1t0TkOY+ZS+aiaQOWAtuVNN66yrhWTjEWGY9s4dAn1vGV15Dxa6RX4WSoDzK
AHmxHcE5udDC4Q1OKBYTgw0a5kKjk4Ows/AabdIMJx0lE+VfL0Ij8gM+fmAXa1EP
ZubeBOU0+Ifd5bkm94sDCZIC+qgafHgmLOoSbLpusUn/xafvi2W7HSe+OIjDT6tu
7ooxDFCzen39Fl2q1+QJILMp7HHEzrnODg0AdWBUVYbOnS4brSZfHiPxDw2hwhFy
9eW7gdJsGGA/xuF6KR2M3jsIJFd+JEZZvGOEgfyyRG1kzMswkTWbofq/R18joYtb
QUI2GDSJTXYRHEierpciVXowUNVu98WB6sn4IEHGvTAScQcdHrhTVHAgHySxmq1K
j7Zh1S+PIYTH+JS5G68PUWsJWLpLgLzimOCbYpbgZEAmnV5igwWFPjW5Jn3QcEZA
JF5l4I7dcSXuLV5oLB6Pt420TibZ7UGeW06/tx2HHB6U2lv5MLABQ9GBfTSS2OMw
p/1pk5J319MtRdCamzG0UMWrRflOeaV8SIpk/DBHtM27GeOcXoftRhvMRmN1HK2r
sQJj3YgjrZ/UUwVi/UW4gBpc/3EcqWWtYGGOm5aZ4equ8daZn0gEKwn3zvmcX9lx
jRkb9NItOA+3/SSly7YiD0h2Vrf9tWZsyVGW2rmnLP14nnO2XYRDYeQuqI9buT65
O+G4iB1PC7N3WQtzv+KIktcXKZOlasT+LDn/z4dA4hYUPc++roqSfZGeGP/a8zw3
g2RuOYxaVcFnvDbF97wlT5XuW2YNIe4Zyies6pNitNys3n7VCCIYr0mTbvIvOtLB
K9NdHU0J7UODi0JsYUz+eWuSMeaK6q/vC5GOv/e3zZEETQyNik96xk5Q+dRT475s
ru0XlhkbBcFcC+fkNK14Ymv6Q54D440YQSjyVhFHebDi0dGdkGQ7NhVnEGZ+ZHt6
oBAo9DlqlaZX0/sjLiFhJ6AfLX0XSYavkDtZprhxYfFnI1Al3XsuyAdQcmbqhBMI
WEn9lxxdkByXMiM+Wq2GRW6/6RcuviKHaKC5ABAYOZJS6hXy5Ab6HJYl7W5uuSMd
a8ueK3ri3mk6t+Y6x5TW13NJV/I7FcrWDCseHsGDd1eh7G/82ZkoRsegEpOhSgn5
pNScoOSfyuPjqxg9md5lu/jeW2eXut7gXov3e5quUiQX8FxfPKT6+UdW7Ofkhzcu
qBHtCF1bnUu2srvpI0KMI1rnrXb4C9U9EIU3F8r8wr/m9FU1Y8CIC7fb4J233N1N
75NNz6ljG5xSCAFsEWeCiJXeeifrozF7fQaUTyAcIpi0CPj5KMY5IOcq2htc1LDV
vuvjUy5nrFtZdhLhj6DDH0rtFjqDVzF8AW/xO2Ub9X4Lp2GkpNY8Kg5U9SBPv/5L
1/4nb7ZIPqMTRTcYVdEd/AgsAKb7CSkV7lSjYgRUo+MaW3xE+pDZdrAH3SU/FXpH
AEAmLBTjF7Fwwh2tdJ/ROL85u7GDsCbNhLDHzIb26bTM27OkoES8SNqu8DXJq9nS
HJtjda2alffxgiK4K0/VDQ56VKYmPnMUeFJGHZKix3vMfd2cHuobPj5B0YRX+scR
cc48IyOiSjgzCHUe2zWyVu6zn6dbPGgYG8lbvDBZjETra21HVbYYq5Deyfu+zgv9
dYb2AXK7ha8eNXDSiJxfr3ezxnvspkyw+u983wLd8oqvd7LcAiNq3ZmZSBflo7MS
L99G0kSy3I7X/B8c7vHzNmmMkFDPqTWgm7K56PKSJh1JtRNkaskLNNkeb+xrI7K5
5PDxuStdQzgComiZChFcOryKzaC/sHIzjDp9Xe9ryAXZRt6K7rSZKNLhDsK103Ej
ywTd4wn7IufVloz72dwqsY+3Er89wVG21XZolA58FIxVC2YFKB5diCZgqWOHTFab
mzEQM9m/+mGxrX/L3YAxtkQT2JYdiAdt9Wz+zPO2ixSfb7m2HecMG6tSnHomYQtN
1HyAWG7iMxdahb6yCf6a5KWysYVSRfu2YCUioPNdni/RvSZvkT13X//3odPwHIr7
Omtrney/dwM3B9HZLJTro0j5uPyViEje3Arm4gWhtvRcT5qfzatvlw1wybYxBj+k
bpuir0qbgKxdz121O4GL9pXR+08h1LkPdHyXhzuAh/Y99tX3syc7iWmQxUHR5Oic
q/Vpbt/oQM5TOqI/qCfFRmQ9GBnsUxyZKejlxNKGTE1YoMZMxyREMNyByi8jj52Z
A58gf8+GuP6sQyjxcRBWtApxPyO0cTM+WuYj9S6+7y8Q+nsra7SjZLZOR6hBymW2
MHnZYPfU6TIiv7YKd/AUYmBL73onPype/gZKZ2aeFan3vD6yAQZuS3/iaf6meOv4
vmAq8vsG5Jx78OzrqNAwZNERI3RAvDLN1WInoytZ5LMmIARA2E/DrB0pXDOuATnQ
ZE3l7HFgoAtTWKwailMkPDNMd+YNfzIj2oD6qKbq1D0OK4VWQ7988TR2GsN29I4I
+5gdIHmJ2j8jTEeq/E8wk4Ew+PECEfL7HQzWSk4QN7UMWRCt1SYbrc4r7UFlnyHt
s9o1N2qIlNqn6Rrw5fy/tIuP3hxUXPC5PNs7Z7GrJHtViDZyrEVLL0aL7sXP88mr
lrQ58UBAug4C89Q+hselxfOHSmKPQYQ9u2mjEwpuEu/gREMe2hiLxMf7CCOthu//
3FdalQBg1OL6ws603LW9XSMd7srXuR2fTLNHAF9j+XxIWJYXdY+bbatjVX/CTvWM
vK6M9W3CArjjSoLyWK4RoeH6N+lb69VOutwhuAJMwNPngqQ3XcwRpSroQUGExRGf
okzE+ly2x/NkwX4xOjJEsQxRDHv5BDaVt1AIDMHZdFhtCBULuSYZbQzHhfiauqrW
iNDPAj2xOgZ7Sv/ZvWRmNXZk59mFLB50koBiMNlJpggUbxm8A4NsOKOY/gdS1M9Z
0kAjcPTU7uqHLZTVhx5fLJ/xVNsqJ9LsTh1DUDDQZq/sRoLEwtzdpGz5PguuwI6T
ofTqqC6VdsCihJ4BtZ9yAvhRxymEZLskELrbsCvfMR8EF1DXvFFsFNSaOIPkD/rA
YOTtjqWxgciOkUsjlpjF+dW9C/Rc49AsNBEmyodIoZSG1n9vHxhd9aEH2yxKAfOR
ez4+jgghMcG41Z6hA5EQdC2V+6dRnQjaCjmzRRNVmw4EZeQKK+gHx+Wf98oAxrkY
oxYoo4i+xQJ2WYRpVjumM/6NkYNTbr1iSzurXR930p0uYFDkMLc3eMVlcEHWJT+t
L9b4OQ4C49MElzseidj/OOHmZpfLabBPxSwZRDyD4TYxM7GR3VReknOCnLskrGLR
AeNrbP3uKLyDlyeU/YR10WoDp8O0ynvraX9yqMvfEVRi9sWJCojEMfwb3rF0/sI0
CvhN6RZQYzXWtad3vKAKfTPlrBNJHOhCTdXwNyhAI0mF1HY8EI9p7f6fZ2JOvr8W
JfXmhDZMpvQClzbHtdpTNRp/mMPseRclldOmaGBTbodL1vAP9lHoL0J+iqh8Cqgf
NsenuC2NFlocPwv2cx3q18tOExBQe12wzsHZ1fnz6QV1G/xbzfJPFjC9DKiBO4he
52G/Vzo5Na/AQgJf00ZwL1D2de+G72Ha2fuAcLOjiy6maHfGmX5QOOkg+I/be+lH
Zf15KKumyJcsLiR/1aVljfrxTpDkcG8LzD8VfB/7HqZsRMH6H5Gv27lyi1N7ejEV
tKFchFVOueATDdJM/uL0sXyrmc48U2v9yW1tJx3B3ozpIfLta+lTK+WG8QpAdc94
7sHcLOf2IkFxmitwPqndDTwwLOQ4npEDEWCW4d6dgSNLMLPnlsof9uLchcnnglAm
g7JHgDZIkvPLbfnqKroR0WJC6u15uzpfghgLTD5V23K9b97M0Cc4EJHGWVgVXwJO
kRyhSaTL/yhdznQOKGaPhw3FQvWxQBqkuUA7i6h0MTetIxVyWSGeLDHqXo3tw6sM
U8sfrh5iDv5FjOlFifTswLItM9oZ6VRYej0duGOTi0T7GKVx0oLQtWldHPIqDrgh
T8msyGFOfhjWj8XUQBuIhmVphPhuDOn0zkuiMdRMxcdSc6wPu7RM7maGCzG9DgpC
2MTuWzIMNwhIBt1ZA72cwTGl2V6Mk+pDln7ffa9KDPIApqUp9lKM3hB5X0itETlW
5m0fV92oRT+3Qj6aHFdYkeANQRIXpbg3H5+m7jxIJ3eHpMXqBB9Tv6dRgYxtA+xg
cC5HYX3I4bCIF2FBnOc2VyCmY2qbh5Q9cjUsknH8AqjX5mDC0F8OyNQKDvNTa7z5
r97PK7v7iDCoQn2qVzr/yC2FOLl5xI9KZXRgyeSphpppNBh0NSXlVQQ2kiYpHZN1
z4bzwR4iGKSWtwILM/zp4qp2TFPlVkwkm/405UDhaZDej/uikqKEHcgTO3x0mmdU
G4vDrueatVMUj/bI8fMEbQmVHNgKw+HgbTICM2Im2W/7LTuOd5N1M/zLLeGGtGYD
7xiZgRBdPiYZ/o0ypb0VjDSVuq32eoBFcnPFFUJ+tlwQr2PB2ztbtoEH1rRZQ9H/
tJmt+d50TGXJvmg4mjn8hOkTLaIDKiLgZWeerzNxNKpr0f+ZqniFY/OCp58Hl8mg
kX1OdyxGIGhks3sm3y9EJSEXxuHu7cxrLAgroE/rLV/vAkuIQxVF6Vr7ki36ZXhm
4PfIyOutJeQ8GGUMgdJarj1MfpcQJ31JhzDQq52QhPFsXWDWzcUj8g84bk2pgSYf
kEczVRqgI2WVo+PmLcFWzfmptU5LjYZYdAHvWSajn8I+vpFvK4j1Dv/kNZIBKkzD
yPHN1ImLS5Tj6iVoQy1Uir9eX12dYGSUmMEr67FZi+N15l9ZAl9mhTZLHcKioWMs
YALGgszIytAtafBWYksbyeIynpL1E2+z9vWyaKHyQDJsntOM90/p+/uAUq2yFDYH
pdJPaWy5vMIZuCrVy01WZ4sNEwMHYpGRbEULWfnIizdODvrwr9ZnMK7nu55NLDvp
RXho/B6g6hvbHqFdqoM4I/w8urNbyx6+dWwslHc5QX60DIEEFNep/SIt5W4M4QSL
Kf34hdsDIjy4ZhsdcMcv4J1e9dzYpW9XzvG393OfJ6UCe2mMhfruFqGEazJXtYpc
tqtdg7MCQsc8jWZR3mkkBGJqbDOayIjZQ8J/sU/uFWEm1rbo/HEfWFfuK4VUHc2D
dqaWkU1fC/kXk+yAnKLa5v+PPTCNSnkR6rdy1htJ16fIV3rbkQk4CLW47E/sZ6hv
POjNNIGJM5l0SNmag1yWXtJ3KLQJxiYGjs3hIQVHe89fPsmxdI2DD5F0/+wMTOSE
XcI9BhMMWaNJiV+QB8KvgkeRRuhEHULywg6zop2x8mSxJCUXfYddJpY4f001E7Nj
ysvGBHSOub7qTvbfQiu7ETXIixuT5XGAKPXGTp/JPJ62aaY6uuCEGmjueYPLJmbn
svwNZ+VgP2nbgINWbGiLy5ntnZ6wsbG4GyiMAIshtaViiQ5Bw7qRJfA6Dv3WVpwX
tsUftSxMcgtNsM8PBntxhbG05AkzyKkOjk4Utcds11wuB1P4S0ETaleQjlBubf4Z
6ROZeWLg3y0HmPClVLWiwN/j9buswhCstytVjOaxGGVAAfLcmIFpErj1eT8I5g0f
j8S3tDOk7pCLQUXnpo3Hb7x2mI8fbcjPr5wz+Kx7ufvGigutHic1IRy2G+0qNUaK
QKc+zyT93kS9KHLlImpe2NEb5u5ZBBkR6jG208SaVo2eEqfLJyfWvMN7aUTnf4L/
Zwut9h1S2DYK5meD7ym9/FwSPVVeEgp9Jy1FfS+cUu7DB1AJCHsSeka8spybkVLJ
Dwjx9k75VkWwQNKRe0JvKfn0XcwJaP/jdDg7v24IbH78E9v1VpAbRzKJIfDHpi2L
pCdf3vckaTI7wO8Vb8/VZn88skfaBs9YQ8PiyVjfuKwfFR1Kl8Qpd1Bqg9pCzwnO
0zspfR9lXLFD7Vvr6+MBPc7ySlw2Rztyw3N1YfrJSgibejGh747AMRAAqUjFzipu
fmdebFmmhb0dTE1ZhJ20dBTDB36NNvtv5ebdY5BqKmjlQYyPwYGGqDeO8rlfAOyP
DE2Hr84Qt5WQOolffTW+4rUBS6u164s5b4581U+4hEr+0OLUAdAFNHDG4Ozen21H
EB/zswvBlZM3aD2j3tjbdT29ZFxjh7h3sd1SDbz1DzwvDO1/bolr+01vQBSRfkwT
XcPulvDtOkJV9UEyh8hHaTFSTe2t9ypS++nmLgqxDWSLVA2W0r0cmGbKlo4tFZEp
nMHuuqPhlS+9OcyJ/hQwUvOB3PuMGCj2zxGH8qK8/1J58NZLJ0Qf69cRpcjV/B3I
2EBkb/iIeiUbebzOLX9BH0ai3KXeTcNgvk9tFUKNpNOYHTIzWYdOKL1BiwHJH7u9
cmXEZWxuzjfx2xOQTCfmiyoKub+IBKAn8mV2N7LgPHSqrqSIfWDi5pT+OQMoDFFa
Uv0XtWG8cJsDHSmgbYtCgE51L4E6aC0NMjns5rUVNC5ZTHWyVV2nGvGrq2tJFRlu
lM+kKfOhwdInV4MxpvKnY8AcjN0O7U4maLSAWR30/23DMLbuvfnd/JHKgu+XUdcU
R7Aow8BipPEg/I8KEVWsJSo1I6S6hzw+tbIaWwXJaIw9NJXS2wlQtpY4pMbQLNPm
XuYr6SDVPb0tbfhQeJMeGqmZkeIkr5IssXQoFgFKUTTCQQ3wRyQDFoHXCPduJnSn
hNNd5tksNAkNSwr5FS6dVmKlSOXYYen5nGqH2MEnnm7B1kXAz8INPxgwDnBOq5ry
66aZ5UKaotjDiiX8NeCQvpDTucHUbxfPkB2qNgroECim+ZXVKzhLqROeWC7dKLc7
ISJMtK/nbBEgWBWr5IStFcu0W34tb7udkr/Bf7DKtijJ/tdniQu2Hg+rPc9jZRX/
bBU8FUdhVBl+bG8uaCmJkMccjiyEu7FmfkdCpVHRe7ZqcsiAWjcFsf5KFqkUlPWV
64bFkGf5zE95s2+m/vBJ0jmy5anIcEr13dxPhJt5kvOgmWxpCHq7zGiMPRYqlHrB
olPaqNOIXtRAB/58ariDJ1scbit37R7qgKM0qsVByflVGVXPLTn6VvanruBq5nYy
Pj5/RVAp4y/KQ7q33391skTkTNt9VLfwJeEr/K82yvThPmfjRByG7j/jv/8uzect
4VMHiUm251noubOKRLz/xFAYUcuS/br1SBaVLEeDcIeD64KsF1ilsKFw8a+xxl2d
z+aEnO07//iT6LCTpzj41bx4GTj3uVCpdR3BIsZlTRnPlBzfdBxaqR0WGg7mNxXP
MghutAtxNGFMDAml5ZOb/i1CvzrBeRFZDY3JPtwTYcTUEl3b3RWuUcwh/lLQU0mC
9QzxGgwy6Rj/Uh+yBZ2R2TXkeVEvIngtc4lDryOwMr52d8eXY8016FBqrmHppnat
HTgEqOPpdvhSP10yRyyZxe12wkXMaJY5VdffcalAQV7pb3XQFvLdPN3jNUq1tBtn
I5OTMnjh1+RfwtmegCG5JZcQMy59IW353FMYuurTGhJbC5CGyYn4Ij3ufl/R3RmX
Qyhah0/Rb9J7nFWYQzj73T+jGwYDxf8UBW7HzyKBtvMM8xC60sVp2IcpiOdMOtQa
gVxhWeOfkPSed8+3km28CLiZED28tGwdAWEewbc7A2fYKtfP+W9msPrFjour7U3R
ubcSxFsRZedTwd8ouN82Pt0kXJNmh1gcMRkVkkm8uU3VkkjBHz++h3+i0ORn9ySp
yvGlLLkCcYOq7y/lpCVgAE1evjoK7qgdWjhkMH1reZaUV7negn3ydcnPViv/vcN6
7XvpFS9lUcPF2o1mVZICB5Kg7WF6NegRR+e1Iu9yZG/Ts0KrMNTVBEDwRoHCDKEE
lU8qBrnB6+ccaKWd4x+0LwwtArkhwoIEjuORZopi6WsrIVecHFYAnRXN5bg4FO81
vSlyv7JOgmzhjBdaR3bNalj0RCr6BAJHHiaRyMUOrH2iP1g6DslNSL83yLRndWGR
X9NcSAx6OuXijWU8vUhfPAeOz54+jX2lHIqIW9uSaHbXCO7+4cb/1OnXjljm+ibm
Ha71RH4pFDb3gQTBCykmtfUhyEih3MZjVMIRuAbQsZuDmXNYgFTocGXAaFYJ6IIk
clc1KEV40GZ4TbFK4SvlbpAGPNh4Roqv2iJE7YIKkJqR+ZfBnkQVT53Hs1nBFNYT
yIAFOksYuWZzvAhgkpbT089Es3iXdm4w2jQlLdfNol2gTu8ImUj7tJKklhAGRozT
cNrbqATjZZ+EdDbnEC03qHXXfhm8mN3Y4VQZOiUtDH0nJ1cVJShuDNIwcKj3kR1R
Ex0+tRyEl9OGXGPNsU2kPeUC91XcgcdL6IB6mun/kvw9kNzanj1t2c+oVBMkQPg+
MxQHoPpU4e0nQxSEfRfOXgDy5EPhqZonNJ5QGBYcBqjS0llVUH9pnmbaFMz9gF8b
8cVD9p/4ZcsROlZITYFXSHl2edG1h8Sv2swGXHvEDvGDBb8zCPTbvmzqVf5rfUmA
OrL1dO7DYvau0+UfDNfX9lxySULwaP3J2SzuCFTud+aiCR43dTNOMep1laQjAzji
OX/oQJC8f57je9pii9aIf3JqaWlXS4qy/NmV2vbGUSo6LNiD+EyfUyV+lOVfQoq3
Ie+L6HIp2a6mEGsSp4N6Tzfb1oX8kR+DrKYqXiXmvzKHlmxI/wQHGczjJ1X5iC4n
QRDcsR7OCoQK+Bw9od461qNtAR+oJP3YZNNhD6vrjoPYRRxcC9L7fCedPqAYtXUI
mM34Swp6e4WdtDyt+VGrsG4ADcqI/iayj4Sr8DilTeDys0dqxfTYWnl3Oz+FHAok
qPYUFu1Kbtis/+8cGJuhcNit5qQAvsDSRPvjQhYup3rRedST6+6UPhfDndPPoJD6
k/rWTltOeRoDR7EoM9Oa+tRGfclxeFvtDc8uSlWnBt6DLiapUYN6yAZgXOLpMxim
Ut8w5PqSnINTnXAQ46iszLbFD5g/YAvO0+YG/8Yj3UF7ssJ4ivZpohPhbkUafK7e
4k1uVSvFl5WD/kI7gfTuGp5fbAJGkXvk43QXhT6iLrd/THlGGfB8tzSrYwntj8aA
Py3ATeZzl5CtkNjSBnwUM95apBgoGIICl951QmwE8rQQfwgRTRpaP0A56q4UHAGs
iNI1YyIJYOaOh+10VJymfta3tjwsClAou8o52m4G7k2saK1khDYdkX60tjZB7vED
KNzD3IqkpbzFYeKKLhBu2+L1mFAkjDeY47TB+TNQSQfehpHpjEI9f8ut2P5OENeB
8ayUJWIrrb7TiVaZNMKMTAI39Qm5n49SlkKzSZ9NTeXC/MhsXGz9GmfcMRcRCCEL
sU7w5OmoZTtXiEDJKMyYArYwqdD9hkRVHpjKiZ+FseeqMBITHxAr1xgRyZnHyGaj
u/nJSVrpJ7/i56dqfNIv5K/hHW3UNobUJ9sUdJmTwd8TbIuXyEXox8lzrm7ifSnz
N6+U0bcETS3ew08XcMQUBVt34O8IEYl2NLurZ4EGW3yITqhQQ/beyni12xaYXK1J
KWigmgXGcGMrnBqeZPF90qr8udGgHqyoqrO9fymk+Ndc3DXPpHI7yxtCkbPO7aaR
4s16Gj4AIZXvywbfxaf/l+r2m/0N/HjvifwM4stfHRvuxOMA1e4WDLzqT8Z/H/BZ
0notxD/EzB3kK7vNCdiVyxHFAwUjblEO6fT19QePyRRh2OvHE6eV42N0qkDE1IEG
/+JAT0b4LNWV01IFJI6PceVJjOG95PqBYHOHvM8JadCZ2eN3CZ0/GebRuw53IeVp
CCAle6A+8q6TRtOfRVgSihRRr+bOJEyqp765Q4V+uxMKTPP11R0MQCkZEp7miR9N
22CXMOSMxbd8yYOn2HtMtYP2RA8NCSACT9xbw3EhYOeitvXd/WSQt7bjz/tVHZoe
wVVhnNQB2FDJlygYE4H4AbY2VUxr7UpKCvOROOi9wXPxTouoP8Whqu8OSbGdjPtp
fVDthcAXDO6zA/FXKfWFrLvrpx9zZ1BwO/mMiqKpyWhey/YptMaMeawXCtAEoWxP
p0Fp89e13D9nV0Ke4abG6Up2CtvXTuyA7KOJ5dxF7JfVDrPPusM7ELVtwZeSIrvW
UffDH13lmwnZzkRYIzPzEzfMHTUQuNs97xi1gJQEHLPv+5Wol2oY+T7sHmM7gttt
6K/Spa5YrOT3hDShwpLIlV+H7uAycgRu8/FETe6A/LJ1/WYP36LlzdY2N0l2G4oe
qeznpqeGIOnTzWXa3L1Qsfg7bElA8af0jShXWA3ZyxmxpJNf9xWXUeuJhFe7OpsF
CuscB3i60JRe2AbiXNojUhtMTw67euq0NcgRDbDa8bR8smTXFQASK/jXx467neo4
vxhLhlLc1eGCa2Hl760meMdouHejH2KxPEkYwfrIIUCv+YaeibMp1DW0B8oHzVzw
E2SUr+/APaQGAHmwpp0T7vwke7Qx0ekxhCTZDNPtXAf4tAKEYSRIuDymGhP5o42/
TP8Nfa80XAL7b5GEs9g43MqIPoH93YTDtnwvuHbF5VqeocT1FjC1TI309WHKSDry
E13uSolxKRmP1oKof04o8LTDk8g+5Y3YRiY90xKcwHKMgbJgsgTVfCkvh7vkcdmH
lAKmz+ZZhrECTLc5xWnSgtgZ2Gd3nv4ON/GhX8H0o7AdhTZos+nJEGarJhn9RT3m
PzZXQtBodx+A9o7xR1EPzk5sxtzXVzuz4gAreFcUaI7L1ij8tbCNNPl/OcmmT0n4
lsiMlKDZMQven/Vtpjy34pa8M4u4lJzGwsvsOCGVJZPHaZfwWj07tDhPGhmc/gp5
GwXRuj9ny1C4/QBxNpDxotfu13GKhKthw3LVJMdjFKVq7eau5PVLNuOEvD2k6gLI
PoEr6rFQFy+px1f7o1kUCczJgr+v4DglFzAhlk0N5bsmSttRQuihFsURG2Yj9lEv
+m1FQVOAfny9WjthvA9sIlBLf+N977lZtd/UE0iYk/lVJCPjhY1SGiBSp/PSlylm
HbYyKJUWHutFeuFE6lZBLIS5Jzy5iPwiJAnv3SMCFtML3pJON8YgB3FOyFQW7QmS
64nwM6ROvOyfpg59ww6CZm1BbjvRIINB0R0y18K0oZGS2+DQo9yN8QaASkxPR9Mo
8WnRuUZgIKMWVCKRg9hypJ5f0X6O3SAX6aSC1vZFDQVaXCIgoW7vGMDc4T08TAiX
545TmO2AFpgcHURocrfKYrmhcB2ZNZ8SObfzBsIJJ0shc2KdDF2X4husIMrQyQNm
9IOTVZpV5mcpYD4O1ILxZTrONPoF76JA14UfF+I/Uh2LjVvOd4bxn+FuhpfKMN1k
RtsUxsudYdeTYJm0GHv2z/vcRum0paW0yzpTND32bCmy9ZpVTI/F41DBiv2yNmqy
Tb6cQRtYLfcdFeyQPNlSJT2WdQqZzJZBSXqlrmAzQ0LCxMDhsNlho41NHD1jPoft
sMWd3n2alkLumUPCUiwYb6Bo6L98G3b6o0FQsGbf0bjb0roDOxyRSrERdF9EGaSA
S4tVpH54yhS9X26cBA6APdCWl41mekkB9RxL18xiY+iZwTXzFn/rFUS0K1lKuzB0
z/gIqB5EX9qv0uaw3S88YO0I3NRRTW3Q0A1uycsBKmZv8GgDkyWa2FWgZFmIgjXd
xZ2Op8O3DXUXWRtYWlamW+y4MqKX5cslh8k1m6i07O2NheFjQa/0A220MsrWVsiC
AxYDN30CggTy9/QOJpkKqYxm3UhYRia2VRdiwtGI6Qsjj/2C9N+L4lAMXsGLapMI
aOHPBmjNCYMsG/gBLKWVfWLt/VnGgEwd1/ALKhVcht/x+nixmmK2D6HlC9dPmC4h
mVrxcXA4l2o2QEk42GQiVyQbHw01vEQ3bPOSyv3/luW2AH+PK0SmSLqXjREsy4Kc
R+LCwEJzluyNkmERMENrL/A0QKt4nDCp9EZIgfaUx1ZTo4uUAP4qpqpTDU0PsRAX
tAmOPwBkLDzfV88OIj68NFLyEVw2fBq2GcAjMVFc/DmmSP5x1kKKp0AUj+o/xzfY
e3d52GVeY53luJe1EeZyl6ri3GfeD4ri8kfg1nmWKtI7TCdW4iiP2BsmNxKVcwPH
rzZn1Ik75FoO3d5zQV+3bXb1GlCFKEq5RONiMT5GhUEds4m+w+gpRrI26cb6MTHC
G877EJ2qgnbK8rY/nlZ/1tnJbzofm58r4ozdBl9CW2c3eW/aEuimzeuWPjV/dnwe
vqyO7ebUGS0ldxxfOZD0asVZsZSv4J5+BpPtegUhHa9R5kG4A3l6gIO+ezw9JtYY
UDkzNwXN85rkbt+I3LKSextqQXdHT/bck5JfRx0SbZ2LrH5/tC2Q99OmBxF2/Bw1
/926Q1vBsRnitY+Csj03JlHvs7EgJM9SDk/o9LyAUd+iXIDvyxwwjh1yX/hZVkAD
Ams8zScR0ga7OSGNUc+pYhADrI39WJlrBQtc0mj3fFOHqGn6uVHGLEHde8oH7gtI
Yd8HQfnsEhfsOLDbKWUZUgci5v1XPhtvI50Jou7n1TceKCthWgq8LbjLC83TfTcp
gP88VVIiFdX//icyjc18X5aW7Yal99nYeFrGkszJ4ZqI1kQ21XaNIo/+1zVVMxtc
ylMYgXMJHhbZiwa2OsQHLntmsDqWH6fUgb0kY0hEc4ZfR2JWKObFP/xUPsCZtXun
cZA76rAIBqYz+bgpeHpKAF5J0mtJj0m5m9BmvosOX5AAAX2FCHi23VNTtOm8Hhmt
6aagHn0dHU83LOJSPJuvui5Cj3obJMJyor3JN/NpFIKckSuyhXjUV6ieNddWcqDF
/osovSXO1DBLG/HY7Sv9HspPqLjlcPV/lWSjA1BAA2KAlU9gNmRsDugMzwV5IJKO
36fRe992vUhGz13EPl8lqYt69/MPKaH+g/9FibrUDDRCEcNX7o72s1ysDBqXTVLB
OmrgO4M/2ShQRDpNlE0WNHPikADD/Ho2+ZJXR3ft+7E4TljY9coW/M78DSCjyy3+
vW8ytIxX6182dHoeue5W+Jq/P+TyxXneuxkWs+Z1Kz8TCgWYEuMWNV2zx4B7j2/y
LWV4xOwH8cjavKOQQ397qa5W+cLljSc7O3272y7P/VR9meZfRJ/7YaIPTAkkETN6
S18dQmyjkdhujLBEDM6qdK8NUmonzS3c2xWpg6XkUNnmybb6SQKRSU4I6PikVq7D
wpCGRQgN9Qisd20pb3Dttdd2uohRxJ4watmZYIy0eUX+9l3fhcf2WhvnntgFGl+a
XWI5e1BqD7NTTXDOJMQ7pbov17lmlzjOrbOnUoI2B3sqUttTuQ8vKnJ0rYD76ejv
DpZy2UmpkXroexq04YY3bbll/8hDbJsYvZAH7qkrMXlIgJaZV0uI98mR5yU0wdg3
X9wJq5wh7kbKNXAvTOmjSBJ0dAUxod+qpr0pOiBTdtfBC1kE/HONdGOxbluxjLVm
BPuVraAP+ok84QurK3ut9XPk6ES+ofLRUbSlu1lFNBvBbULQ3e7NI5onQ5f4GQqD
uAfHxvbYFdOaEjb+QD31yJY3U2N/f4QWRThWYyNzH5u2NEskahcgmXW8OIfun1cK
MgvCWzi5f0t7TyAAZZ3AP8eFIW0yfKvh4CdmRejZAzwzOFdOq7TF5tKqWZM2mwOo
6QHUe4JfTxQH9cPfS1LX1c0p6loAAhv5JQPbYhrMXg/LgBRIfI0FWg9TvNrBMRRM
A3fJPtY2Nq+BuvUaP4EcFxh+QKLpOp8Mi6nO6kQSCYZktg6Roy1oxwhW3RzimXM/
I3OX99DSXzT6BRk1jnw/UKkp70m1AethBKDPf5dwtdveCMIypjD8V+r7oFX59zj5
Q13Hst+6A/MoGRoWsfMbMzAQYnxTXsXK2Rx87v1BXp3dPFTvfq47FeM/BVfvwQro
0aYgRyAZHBJCyjXAd2Du2fNxa8T2Vw04+VxisBOmUJGxsnKmnk/6dnktqZ9aGL64
GmnS8Tdu5caoDmQGUZZskiyzxvSJAM+OS0npvw3x5/vgJTh/68Kb8yhCiOH/ahd7
khBpG08+rqwSzysm0LCE9YcPg/oAPM3N9id836pUdY/cS/FlGqh06xhTpIlOkLF5
QIKIZZsNTF4FvyShs6hPitSQc1hyLjdseLc3v8utpAM5RkRYZb5uxIKAyksxsiTW
YFZaP5FujSunmUD3py87E/PzXlARLMLEJsgY04Fww6nl9L9SR4p50s7bzNmibqCQ
mo6lu5iKgkaxyYwIHrWgUNFo0YycVhTYVPKyfC7Q6L8/7407RRRdW5aMPD/6KCIm
1oWng7qA1SKHcZ0Hh+DPr/rkPxW8ad6Pgb47Lzbbwg5xYNfaPMrKYcO3N6oHxwW9
MAlHSXsinFCY7c1dlZ3VzCtkUI7+/o0LgXaEO1uDlyCzWcCrqyQscej/wS+fVy6Y
iNrR0y8vca0dUQFBHAdOwsUpkvesv1c/fAk/bthlA2aMT6sKFzkc3wZRFRH4uBDM
SDmZ3PmIUnAFDCXTuiwDuO+4gk5q6UUW8xHv0p2RpwV8yRNj1LHMaKQjpKr3sPVU
FxOarQ4ouJqyxnPPNT525a7/U7J0sExn8QYbnFRYiAbYS8Hna5OaICqptf2Sbdo2
QGDeyTAPDwF/QPcPBGclNvlzAU4rE/d6pvuspoHBoDTbS4XIDYjrzuxMdE0o1LkW
v54wMo/eNfSSxChDlwEli8uhUsWnf4PtMbYCqWHDaONWWuFO+xI5j2W8g6GK/P94
qf4BfrWiHq8y7p7gy4AVOUkjvV0JCMGw0k0VZGHa6A+bPRxQcFl/fheaDVwmQfoF
Emk7IRnp6MMhsurplqovWOytPtlS182iZFvyHtA9hD1DaepjoS3rTZKcEmbfHBoE
JNfw6rl9fvarN8WO6biC3qeqK8XOrTNrOb3RPJHhR9/AW1AvLamzdeHytXGOOakd
wMyUEgdHzMLhvQHlm5tMh5d7mjKjb176AAdHhl1MNxWUm23ycOP5cqMbL6uL5u3x
12wXCG48QDt/Owwo9mf7DXRFXt6w/7tGFRiIyyPr9FCXKzgHdprYCl70RQSdBYq7
D6E5Zdrs992v0kYWnjNyzSmSWus3m7QyM7T7M88QLIenn3H9KAwFGo8gUdiRu0jK
V3v2vzSeyC5zLxiLSHxsWiScsm2VsBaI8ekUmrVMuj70JoFpsUOjoNnNdwlb2+Bu
a3U3FBzv9BUZ67M8SPdfk/sE7FRqej44Tsujg0D4q9ZSWyO2Uc7jgIXHy6wwMH2g
JBPU2GqyRE9OwrCFGGYaF/tRhSfNsMxqKO67hmj+C7BDK81WLvAQamJm9a9bmIZz
Wc8RZex50wX+PONZN1OXuZTgPZ5lZMjJg5LVfhdgF4SX6lc4ExnMlCavzE9Yml0d
QsIg5+8e8eSlxIXB9C3L/5zre13V6o/LfGfX38vSWA6PEqXn03Eww4o8vtehQAxP
vHH9c+q2YHBWEcpL5Mb/wPe2R9qqs/kAlRZNYaTfqNyZYxkMkUQfpuuZ0IVRgVwk
9jiHFr6mQV6YooqO2bppy5+btnSFplKavSXNR4EOVDZjk+DqjE/N6i+u9ToS2lUx
S1pgUMQ6XA4cmsIxD48goTb+QNO1LaYAFaE+4QmJ2sySfeorBYFsvNdJVmLiTW8W
2riVrfsb5o9HVOt6bIs66mvniZybyKj7J5RcKTJv6W7sXVsrDBvZtGdZ28i1wcrG
qD6IScTYJNJoiUmvug22TPFJA+snO1TVAWG1yOGV5QmNLaKJ7EZQQy6TDG+8ZasU
N7/HUKgsik1y3dbCuGpROUK0RWkvn1dnZXPTykL+kKvaY36KJQsf8RUAwdpPgpGi
c+SWzwEn9K7HVI1SYmz7ePayw+9d/2wn8Ox6+zl7TZ5M2oRPZDdrwpmA9lxK8Hio
MIBITyzkjOEkBSdZs8UzywqW+bucwva+Q5MLkxqpTPvTYrj8OzCvsXfkoygRXvbQ
sgqGUryL9mxtpV7kqnepGSy0SGZalKw8abnJTtXQ5xJJDqyxO8u6h+/Ylq9qgZqC
Q1Z303MjfL220d6T8kn5L5BOfwK6URC0ywVARIo6sPeGlZKW2T31PHDlBM/i5Jwy
ZpcDJFK86whfgS1YpmTI74KQf+dmOF5aaob9LtIbx1njAOOvRRB/YRegeFvGx+kC
YqA2nI813lkYS/YxjWAc81Pil3ywF75r3vwmCC77S/cnGG++O3W2nKs6/VZJpcx2
1k8NpnPVnrgFCUeJcUTzviodVnZY3QO70rAlK8rR+K2KTUe/yCmFBa0c7ELDKf6O
Yy8LXj0xZcylzGA56arHxseTfKsTopxo3jwTBjdCiJt5LbQhXG5f1v/38kO4sdpA
y97a5GkU15zgJ7a5OLjPpIV2Rk90P8980y71gJDIILRJtZ2JyGJi4ktYRPF8BmgF
SyfSB8CyF7jiveedY414W4dUIrBEIB+rylbBcCMqJ1pIvHNFpEDC+vfAJA4xpXaT
z74au7DDuzFXMMcZIK3MNPW4Ad9c6BcbLhhleL9O355gYC4e0o5RfltePB+ki7zy
2A/4d/5SL/n71vf0hxJbSTFzQxzf+8rhD4DEDuO+v7qYpqHqwp8C6SOZz+yr0Dcc
nWUZO3iVwQz2RoAj1LeVyu9o53W0EgKqvPvkJp6cvzAe0oIR2Z6PsGnp5T/bcrU6
ZbK8mH8Qqb8tqU/Dz2wJu+G9vHssmkeKeF2lcpTzMDE65GvqreI0r392AMhZuKKl
Nf3jb2IPCs8m3rxr/QPe0PuPjK8KBhKAMhjaCNLrZNpGmAniUuoZdkKdhAIYWWpl
aH3QlnXpXIuyGr1nEdmf2gRt87R/dvd6hChBEFNPC4/3ZeL1FhQixr1oVCLGAkMY
N3o3tbJ2U5TtcpNZ6Vg/10xPquMsWPheQqj9Nib/Cv/1NIF+R5LdyhE5gnP3yu6v
lf4n3oxJaMAbuKU8Wu9Hw09Fn6eeVzkq3siznvntFGYkBbasMa8xfxUCTt8g61Zw
e2HXu1Bs6Y3DqqWDbWSbRRD36aWPSIGFdZjnGEzLdKiYFrrh1etv9UZlu96CjrMZ
SNh/hemzyJCqn4EXQ6pM1LJXLqKYs+zRUc8UTE7anEuu+xbGF1R+vqlf1hS0PS1C
lH8UueBx8uIQctaJAgJ9PQQfZ+HvOkpcQPOi5EmQuIpRVLp0vf/kfXc7S/9dnAFG
/WNJ0qQw3Bd+1LZyvE3/JFlkQ3ru66/0eSg66Pnt3YViJctZ0RrNk2zAssweaZm3
BhWXwqit5vBvHi2+S2leyccDZbkVIoKHrrKdxdrI53ir8vSjtWA1dCnSpiTiIBby
TNHxB9CQLWwAdN3nHmegrjM17DNWLYscL1u8kEUSnZt6O3AFZ05+bkAkmk3PutLt
Zs0cAubNRFlOQjXsZZqQXOBYdMdWNMz+T5GZl8pQuQvi5tH7WbtQ5QoqozT+xY4H
vP6eGYf97/r1ICEmdBDTmm7Qk/H/uvDTpZ7A6EnFcOYvTJjKY8Q5myqxyBlQ1RLh
C0OGMsuLxr2z5XCZ6+/aUH+mxmUqcyh1vwb9Jm/4DECKCTVPUb2VBlRFxYh6heON
7JPplGNj+xfwCzC8KJPK5yLlEzIxByNZfg3FpS+D7UPL+UC+RI5osQdI8uky1HsO
cJMUgIsal9Dur+Llz2y744lZ++3GSCrQ2mmy2I/CQa3hyLuwCq7momqZhfQ9i/Zi
AOTK8iWOygCOLDpv79pdoXIt9jMWk66wQ5kJ+E2eZvUjqHq+ZpE0kSmA7Mjy37dl
UXZPnOiLmbS6Ber9r1CsGh6bNGMkawg9SoMumd7gwpW95xugMy7NICHVyJOaqfK5
TdQm3KJI1kP/B1xMeYtObY3z59e//UK9jsfhZK5GeCiniAVWOvHYZQjCo0lZW8yh
EJih850Wx94ev8l5sBxM4AhPKNNEHPkLLX9ZmYyMRZCNgQLw+2VEjQaeBfdzNPQ9
vN85UXfMlwtBVZqhhmWkAap6l/aTVqfHIhoPe+/eCBQyX78/1X+3F0Yj/2WPO2GN
mCnCbAZgXULgRBigiB3WxgBSGNnx5OboSFj2Bkjc3of9eaae00eEk+CG0y+DAWQo
CKcg3uLV05aFmTzcJtepVQ1hzziu9NcbkdtPyerWBk41rzLUt/2mkrQnbinnZuf1
nzU1sSerPxCpPWwB+N99/wg0u6Y7YHBVSSo5ui6Lyxg/EFWFXxDeKvFWUrswPMjY
ZJrHUqYdNnAbR0suYi1PuXQUlht+zfJdDX+n5OGgRzWIuH5WLgKhntRSIQ7uP6V5
XLq3GctPxbOlIV4A9g1xWgYVP1gIe8f4Xv3+lCGz2s9nX/P3lQTI8kAEfmOHIe7p
zoDMKznEcgATI2JLXc9YHZpayTe4/+Ek1gKfJTDq7/zEGgTQQ++MDQkgDksU5oFW
yDzGXsSFnJ0jgAoSj1PNCr2O1Nojw3Pjjq7PWRyISOKbvUnoD7Dl2hRq9skipKHv
NPcilFn2y+mNnxzq1I5d+/Vc0MsLth9Sz0Fc3xCpcgv8QArPKQAzELerDyaIFoO4
E4tzydEuGrkYcKX8SxB3nCMtqDZMUTCEvkeG386cCfQ21SE5aBNlnmw8OpdB7N4A
+AOvEmxzqgt4GNdU9iaeIhsiWTcmcHZjZ5tD32rJnam7k/xDUspwk0tNWHd72Bxe
/3NhbTRZUy/F072Ed2ptr589G7DaWB7oKzZu08LT3Hn/8947ENmm/KM+yYZVX9P0
5lgRJq1KCe9MsoyrloV+NK7BFQt3MO6BkAjKE9qzQfVapNn0nVxLDowKklkvdZyZ
1BVdBscLrWK3P0ggcyfXpeHdRLJ0zWkpxHMqcZjMf1XtR4oySMakwbngKjso6NtD
NvYvW99+Woyznd0C6KsasL8wgI4cGgiZRdtbz6fRakpSxq+vCX/ViS4tz7AFOgKu
NbOtvru+EKjtYkzFWMGwhX2nYfmKrTsZJp1saGEsUU+9E32DNgqJA5020DWIFZoT
mdGpSksxVizsUNplV/qNrShfvZWSRu0+VngMGXG0Tn3silDIQy9T4W4uCrdtJHZj
GHzaZIegTrmtsKiit/Gpjeo9B7/cD05LHKUumod2Db2OMq8OglEQuUQ0VRW+PEiF
pzIPkDyZw6sGT2PaVx7vGJqw/AWgWrXtdM2HQfsj7oAZJD1LjA+72TqyEMLPXqDz
sNguZWOL02Mi0LEHa0GLiIWy91iLovQtKj2DXw8LymdDtHssRRJzJzybtybw8Ye/
UNlYlpkXn+qqwdOHK5bSnDHM2V4x8IutViBfNdRs3ZX/+3rT9nJYkm3g1bIbN7qb
qI1m84U2VTiC3TsVaddYpPrUM1bQz3y2iczZwhRXlk//UO6LzzdWB3aMpoFOS0DD
aqQrnZC3yoq/E1NCeIZM0WhFGPAI2JvNUwhaJdYLM46LqqExMnGHN1E2IHYt5Zh3
fy21WlI6NdxgIQiItoDh5SUYrep04UUBYA36jkg1Omh4KRmlIUAZkJLTKpw8zmYY
cAy7LIEfufaUY6gzIJxPLMi89yBwxRM7v5x6JyzeQ2woFf2IfE/yCfbxKG6XKWFK
zaYRsmTH5kb55S/jXgO7mKNR/HVcsntjhBgXs/5xMabcTvlB1vBvnanA6RyqXOIg
14ys/nhHPgyi2lK4+Uknq3TgkCvscAit1mqm+Ojh5b0goakpQP2N2/4cxyR5dTkw
/ph1CcRxKETf1kVd9229Nj0RN5vAEll0GFnqGNgkneXM7WijUKqOIarcnhOo7s11
ksYW+DurHgYmCGe2CSBUHnOoe5CFgNm453LzSYmzd80JdRuMHf7crlVcETPZrdNz
/vkk66m/HVQdX8erBtdkWXBOx0mNhZdG/CAb7q2UtvOoLxIm562cmypHkNJFUpLg
zxbkBdR8nYi6wmjHYf0aIBHD7vqykzCvqVRZIfAo/MTxv9altPYnR/MxEx0byxPi
5bBNt9N2wAQcOO4A3gS9P6y7qKK2t8EaoEMiJvFskdpwPpGknGywUhah8M58m6X8
AaoQev+POshp0YEVuAgAk2b64v62kWUFpaVRiur9IfqdEhgIirNkgoVNKHJZcrgY
YVejIsA0WgxptMsEIIpp0rJr38S973js59/2omTzKwTrWz6Azvd49nI2CU7FTJl4
A2BkMfRjzlON4ueuZdv+lq4HD50ITAQZ2OQhXBb61BXfXWC2aAb6ptVdFT90keUC
TGkzi1a5luszdxZH/gAJ/Tlw2kjgQQVh+c2waR+cbi4Es/io0C7ncUsjO6yFMzXn
cRzEZ+Qv2XdOn0zpqy5CS8jYtjgM5BaQxW+JqYQsXVZ8/3DXinrwNgpjCztxtdwX
M+M3HkbeDAwxdsneZkJBjKh7xl34AW7HcVhp9x/V8AWqeFx1CSI/n5lswRzyo1kU
s/Fjrmf92aSaL8di2Wfc0+iPmUWLRLqHVECGF0ApXr33c01QZfrSmSG0gRMAU3mU
ficvdbbengeCy+pLTsxLkvh6xLCmGLIyuuZasiXCks1SnoH08AbHVkOfufnrR8db
G6TIsztKT4DKQ1N/VDQQ2GlZmmChXE8TdtJWfpK6XZ8tcUGHAW9n0auk76PxIMym
Pgx1rDTCgt2MY8w2/x+/mT7Zw6pGKZWq1fsOWs9fir67Ba7UwM/YUlpsdW2Q6PX0
Gp2h859H6unG1dHpLoB6/EboRC+dAi+2RPQxcPWattlOeO/TaWMjf7GG/ZI4cXdH
SKTyeigShJSsi612Gd9PV+FbwlEmJrUmUM23eXtsohA0PcufLWkdEUBdefIoG+tA
Hut1JpV3VpCNTLl+bjnY0EiV2/vC9M2GZBvnn0nr5qFOiUa3hgpHPlhRj5Clunyl
7IvjnZ1+/0DY8mghG0IJHyOSlaASeM8ctVHBl7+jkLicMATYMj8gBjXujmgC8lIc
d/pWjCZOXo+mXstmxrJD7Jm10Bo45eWFj5LFSNIP57lP2R/ZlpkmKWpclXR9YYTJ
eMR9PwQo94E6QyL7rKSKeo//wD0yWymvXebpS1FzzyDpu1wsPHqFlKzGiQdc5mTi
3LvAr8/NpDTdYBDoRD2TnYHL3cL0ArvuPiyAHpMfdjdw3kFhzMLGYsj4sOwZEw/O
8nF/soJ6a5znqwuCkNZggxuT7Q0+6ZNobhHrw6PXhDLqbFJCa4sTiz0+UCh4lZIC
VBdGxw3sxijVqAGyj/1Soizjqq+YgoIGqXDx0usPEtF13taVrlXhVT/9aTNKGfWn
iPl6FC4b1Rgj1NEHsXU84M4qXKqac9Ai2c8bKMl2cYXwuE+32Wgde8JDUOF1eimG
ykVAiu1v/QaT33346Td9F76pbGS62G5+3oTM5iQSiAoaXMA1Y/NX+ar44WmFPMzS
s7V1SscZgDzShLP0hyL6j+A7BFi/xykdQTkUEPp+iutf7pzduxInMPYS0xj19f1d
COmINd8ePfL2FWfs+UafFFsZL3E1jrubXWiRJGhMVD9ru6/7JjQmWbcZ58PGuBU4
2sq3IFJgLOEyuk2lkzukK3vpiHnIEHeHjc2MXFw/lAgc6sSHL2XEOjBplDWKLp6U
UrL8dFjMTunYYmvlFHwCJAKt/ZQpJiY5Mh51M9cnfmugrJhzdXHC5OcAVSU2xYS9
MgTxT8qliWItpYavUlK3vTHh1E0FsSGpr7T3Te9ITXIc7zzdBM4eHA1wEKnTrMyA
a0xoA/03dgmp/JlLdzp7kOcFzWQGrSNIBI10VXtqBUvnU/CSac6O27K1MzAiQtwS
WTboLODHWx1fgGtHB4NKf6D+5ekH9RqzFfaQMWqkaS2KHkd5Bu57RTLLA6+a6uZU
2sgvsierH7nIysu0anMaZrlmuzAZpfu9pjSYGu8Brt0IbrngJ/SGIpjlayRtagrs
iqB8soVFsc9txemFwtkTG0WUJPNgGf+URyP6rCWGpOXADYTOV3szGzu3l2oY0ITM
FtpNR1b4+eatJ1ObBCJmUYI6S0maIssKN5HXWVThMfh3GBMmxgwNktlOfrUp/sLD
5xwwaEWEbDWYJ6AdqjnYWAsekdiDINLV9WEG0T2jpexqeiu7nQGcnU/o4qg9WD4H
CQfeUlvTThEHhpeBAcV7rtqzczQJtRX6GfWnb5/jYH1sAJYqV6lODestiyigZtNc
mFA9r4QP5YqATIDoLx1LWH9PQVdT17cY2xWV6qQJkcSb7ArDrX91q2hQdEP8UUPx
Cpm5fgp8YrWo9XMaQABWREcBTvvL2auwWyP3JI1kcFfU1Z1baU0HDrw+B9y8FD9B
LhyGj0HHlnzQ+2ZpnXyi5UrgDaXG0pB9YfRo3g8gqKIHkxwVtEj3lHycnk1MuZm1
Ap2Sjzj7FB1DY7pSuB9zE0kXhOfryxtH9pwbTShVpPSU3505v5cwhWD/7aeBaR9Z
NHgS1ssr2QNoDqCXZfPU4fI3ydLRU1DqFClmbUYpGFfPKYAsakXPVKKB7ZUjlFVY
vaPbe1TlU9uWK9pHbx8BzwkLd/AvyUoVIMoFCuY0tU3YISPS377nPWdtuALJWzSC
OcH+zghMevMR+02ZGC2yZ4sG6W5O6+0HdB/NfupRpYir4D+X8D3IJ1wiOfWp3TOz
b3Ij6NamHkSpbPkqIHOMFP4VHtU1p2iedtxacGwyGbBb0rQau9re62Ipm1LPsVPf
dp1PmD1o57paORmODTck6sBMB7Qgy3CiadhusXi43g3G5oIFURP6/zamdfdTZXLR
my279M83eDIrpbcFBfRO/auvDdfeyBWGRU8otv2cPb2w8BjvLPPWLjJziRoRj5FI
4P5Zo+dNskp4G8oAh40SENWvakW2gp6hvTzGVPprytB1S9calPkf+fWfeLhp1rB3
/qQKVBMGwkvdrduwRVymSfMb2VDa2yfOxtaRkaUKq2hFtg4OYXYqVs9NmGLOuqaX
Dz0Mo+Z9Xy/FHRAoH4opDywzIwkmHeS1rO3TQ+3qjkMd9m/2qDn/Lhhouc73a2o6
ZTTlM28mChicXTtmiB3o0ZwL2OWv+dMQv1GNBaIVyQSsW6LZvpT1iV4ejDvYqEsf
WUPAB43LK+9wMXycHZ2jS0jA0JrvZ9qYnaAnG0sOpH1YVkzN+oY4FGniSAuqE9kt
hM1RuF0V0sPvffgpeJQ91sFV+ycEofdY87q1Dj7y8q+s713tv7JTyMhA/oat80O1
G/gmQe1A0yqXMM0KfCCg/Km9DedDYcBjz592b3/EWYu9zhWbb6f6BNUdspMz+2rM
sGoxfo/eikhQ8Jz9R4nfNonDSRgxkD0Wha89jx9fk78Jx1QBdbdB0qDSioqLCcDy
BzXpqhfozpTPPZbJvMCPot62aXQ82BArppUB8IZ/FpW8KEFkDKwvtuoow1jZYs7E
7CNj1kEfp2Q5NyzbdkqGq0gi+U7pF2OgkiRTDtnbuCjTqbRfNqGGf4K6QA4tzyc/
VNSb6HyqQQJ9/LqV0GODo2twa4Cpy4wq+D2FgBpX584+n5bqxDvSo/GmudKxczLy
STtRfKRJtVpyEuoAIehAWI2ppr9Vk/+d051r07+OqyvaQddQ0S8B7xa9K0pis3gJ
SdLkNK+b1naWQ/cU47ElBhfW9fizQHKNjx0JtQv4VEJ4KYv33l1cUl3JhFZQ/6Sy
S2zqQBeP5S61Ky4cYdghdiNAkApvQZjEbjScppZgbpn2Edm0Vq0q+ZfRfVb9z/se
LhGI0kNxKQIWRrYIkN63HRkaKjNO2UFEPVJUQaMddr6rEB3FgZlVJ1lEDbEn5OCf
mRwtH7JECapwEcfyKKkcG9qZvcJBw91gVbtz7jVtPRhC/2MIY1tF32z4U7oGkMvt
atlBOUK+FrKgPvHGELAowDc0zbB05Oru2UKn7iqapti+rPaMu5I4pcnvjWkW2eni
nUv+A7RbntifLppWHh2cJbagx2HjPUl/p86XXIKWs0/cARtDBzPSLB4/CNzFdl/l
TCeBWihLga3IM3u6D5gD+0d0xkKmtCARLb/AdjsZKYYl3MaBoTPB1GIie4UxVtnw
YXI6sNXfSL6csZd5KCJLeABUs56kmbGg/agCEkjbrNo9qnaYqMW5YP7/2qQ1bK61
ymJ4oXWkFVB+giScXj5Pxg1XtnifPOkSrKSG9sxsC20mNnXCt3CnzboWaOZjY15O
yScA8oTOFxWwCEx0EKkGqZsUeqqeG+MM2bCf1rEZXCUXKq07yLA9o5VvZmdwODXN
6sLiruF1HwBiVL2zFLFk/e0GjCq/y1D1C2QHP3xAlZoX7/1n2ycF9exgy9Jho/fU
AIZHgdeztZU5hBdZxFx1SPwt9BZh1sv28b37WK8rtPHeTwa9htqwhf51WOzdIrnG
9vuCmQsfDWr3xxDBK+tPeZjKlxvwK/vUEQRAyObAm3WfmHg/FtWB+Aeq286TXI5I
ly2MsKzKyjWC2fmYh2o0T68Dux9oaZltNgglnPTM35knGRZj9tVJmeil921WwVzJ
gFmbFrRdRbl7E56CAuS3Gam57unl0G1VIMCz0EJ19BU7XAUP8Uf2azqLq1UvU/v0
x4VrN5VR+epVzA7FpiSqBtSPTl1b6/o2PjsJn+pfzfUR1ZpJrVI98Y1vB2FU2lgm
VgDGLATpyrC3t3KIodYRdxcdaZhBf7YL7ckGKw9VEWHgtzMQLUwlKisqkfXuyuXL
En3WzBIE2V/9tCZDCvMOJV7BPFflvkjv+IpQFtktXEgJFkNfxnmosAgOFP+Kfjwu
S2vsMtayxn6B70BI4PnnXZ7fKafNbaNsAzmzlLUTl+sHBs9WtEOR1dpuiaTCYoHT
cR6EuRBNPLPXSuin77ALe1AipgLvLXs76Aghw6LedOKE8RxSJCFUc0b+NzWwEzN8
ox5Um/LSlgiHsotluyFx8iSOAoYmZS2oJncLaoTE2mjoGgPnllBsp44ozEkwBEjm
KvpgEzkVnS861+pn5T/m1JMQlq+kEzFazMkL2nZY5GkGcyXSAXLMCpoIXz3cdybu
Kkv3+v22oR9CWmevd/V5sKVlvVQuayMTD03RLGhGuJBuAS+gLNKHZs0zZecFtnay
Mq6IOXYy/kyMBj5rN/n3XVGNSfdxGfPkxgxy+KCjzJzKGmBmqcZlGUR3MuF/0a4R
fOdH7GA/NbRtqKuOkaZ/DewcYn3jlVIZTvDnNNVQlF7bRvwp41DFKWFHQVJdPSe/
7IBKhTO4zhaFJp4DDnD/bdpaKWONKWXfnS85ZNeZvbgReIlC9WRyKhOcnE/oLbqC
TjxKjkk1ChiTAeShcgToRrMnzdhgFzNyepX6OSSxE5qovbk76gD4H1nhs2EPtG3G
4kjxSO09a55wHgAmdnCEfMCH5A67grhP+fpMIvPIfcf85jRd98PmNawPRYQMEhcE
HThuMTr6Fgjbru9PA/3U5LafXOEgXhD/pa9WXCzkYez+gDuPIzpYqYmq+8MbMC4G
QqQlx3wP24iakE/QW7U7oKM018MhIBDgioYMVuFrYLZjw2Ll4aTGifYkFsClPUev
E4CyS6DmX/UThJnb9biXTCD/e375TJgMpSXPPg6xDG/ydOGMrgZPjoqmxse7N6Vt
U5Ukg8b5I+Y0AIJf94Yl+0vRr+oDd3vf672a3VTmQiD5QCIWTaTi/qrmM4bu38Sh
tqtqOI0MVm1jHxVMDxvsn3/BZhy/ZX/HyVH88+PtCkqdrlRkFuCGIF1/Uq8pLE5c
zIZFE3sxUqkH+Vf7BkcN657kdDL9pwC/tkt7KpB/3w+/9NezkAiglKxx9tGzpyLk
Xiz8UVUO3dKmaEdPkrX5eIbHwHLJ+SLykbCrCb40SWMZxlfLywqIR/ABi6VjpcT1
vMWr9VBi9/qi6ygF04BJQT2cPDM2N+MUl6F8Q5QAJhh/kSxmP+Vz/sHkyoJJr0pf
BsPauiu/TfzKX2u0ETvvaZ8UN9uob5vOJcOYC/8OAOvpmq7XLrN88fVWEIj2MYB2
3t4+Kgmf98hO1442JpHHVCOBWzgaPZMuYnrtcjM186yI1KLQZMumZfC8KLnYMJSD
LSDf23brUKhKQazfdVg8Y32QVX/khVqIJHjnJZdYvL4Dst6n/626lFXHxR7sSUUt
+1/4D2HzNY85Br4jnOdYgYlEtFhp+OGUULCcXOsa+cyS25fSGE17I6RdvFBH7Gh7
jUzIAA5bIMSQambIJoj+pYguKE0VzdVXyvj/A4lzQq6lFsgbK6Z6cIcjd6mTtIZb
Hk+FSCrQJ9mSHv431FjzAK8ZI6tA28h+Hh5ycJJHWRHQ1I5Y3T42mti3G+CHd2ek
Q1y9tScniSfEcoj7MWcAPbBLQuNoAuqdFo7YxCMVcRCr+XFqKVjHLra76yM2XdI1
UTkqEeFFxxi777aU+kDcP3xQcCVwkN48KawhQLU0sZ2u666y7SQV4cZr4b9SH+AF
hT/ztX0e+vBNjCYWss7bBF1xaiq2HB7tmHI1UBGSOEylEpkE3WnKbFYf+u0OkbBG
Qyq0x7TtbBPWXtIUQ2OzNsb3mK6SH00iBeaNXbami77KWglPp6m9FbB+q0zY3obr
BgRr91nFfUQRMswAWVEOlRg0ItzmhyvUBYdWbbaUzVIEQ2zm0dBHCfGTFoiwd26S
MNJwXq48PZewQZ3T5wUPq3R9p2QlcvLQ4cPr+Fcf+tM9bFQWqeH0JKXxuFsuwQvN
LPYt/OvgMcC4OJ1nzOknuOxkOwUt1D+AWRar2pXEwQR7WAV5iCdebHCWY2Kdi/yU
R1ZvlsT7fKwlsKtNplceHbX81iQ2MywTz2GrcZ3t/aHIXUxlqRJuNEMBzkp/JzkQ
DFmhQNVQ8vR09CT6IgowH7HXMk1enqK622FbN6JllrLxd0wSKOT6od1GvV6FeTLK
N9ZsFAGgdLXM3Gs03yBmnHAeDGGxgh9z+mD8OT61SHMe/Lf85/X5l2b2AGgs/qMl
m+kT4M/JokSlqdsDA2mMsvzBZBvzaHD+qe/REgKCHpleGqTIU6v/OmgJILE6xqZC
V53r98ZXeUUZ+BGr8y0jUzFcVSyWhWu2oOgfiADHg9plVdPCnKJOB2ROa+HhPkUV
/9PL/xDX48myUeBNcvEtyzIUBr+6OtYAPa6IB63Bt5ZlIFdPR3ysHyizVx2Gf9xX
UZ64J7gdwV65PJg2oHi/p/TjtCzAWGO7hpKQC5vDtR/abAG+rZJzfgS0zCfCWz4c
21oyQsQRry+sLHOff9ynyQhHuzhqKio9A0FQTxYaF2ftkrYk786DRbTlqtT2/n4n
KWHcnzqxWxQkATOxyEf9nXwug//oGkPxWmjXH24GQYAxWxFckadFyMK0p13a3VoH
g3EYQxW0GJ5ToKYAST7+yVSOMzWZ5Ri26bfHQn7wTdvUQWSKyN2jC4TSVo0djc+a
+25BDbqNmgQBRSLgO8YkOYSFDGEh3lhuoAmaZFipJoFrxPwwi9mPFOfqk8DzBxDe
O5tJgvgZtgn6kEz6ey7319VGyDMj1uv88FIVjc1xFXEJ5Qtb9yXr9Py43z15rpiK
Uxak28aZMPKtPUR3f/Fq6kgYFIUjHxQvsu+0Ove8vDljnJEK6b0aE8jUAhtrThDB
jkLQ6fshdIOGwbeKcFZGEs9cH3soR11H4ttySi6SV9b4Mz8LtIfhdHcQM/GekM16
Xv0GXUZYoA89lriNOXtQ4LUFnMG0I+jwVby3xRlxApM7kaZblzUkFrjVeR2y2qJG
nwquJkT30BLEYEhF1XEKKorXGdo2u0bfdnDghj3/ASZxwgdYNCVjKqK5hI+NbFBB
d8nrib+W8iMx36AZS/OTZvP73tOGso4HX+D9P8TMwlsxiUL0w/QSZX/EqRNA/KB0
JoS0g4Z/2rT+Gx3TpwpSr5A9hck5AaUSd8yGv85dpKkh2NHj9GJzXNL0qMgRLWib
uzzUY+7DVchZKBBDsyozZJaXxsRlNVj3HvLhQSzSCRSt22G7ofoUwKzKnHCR4KF4
QZnPC7F6VXoQcwLFuE80IZF0mZIgCA8/O5M3PWVef4yD+E8kVyPNKwAYjAmdt8x9
Huot5P7Qt4WkG51UlkSNbj1eJK9pLwTmR1inyXIb7zTzscMa0ZW0kpXKn9gNKuAQ
HQJQAzysc8gbrSaMGJDcQsSGI6E2BseVx6978g9PjwfhG6tzjd8ZTu1HMoAWVFsx
9aPxt6huXkUcn45rPKQ+IsdZ3YcCc8MKnqfFsqKstUoQZMVNs0T4+sLpmLVnsrty
0uYTLP3ElEAsAajFThTBVuRITMMwY/KGHvfiaXebpJPS34EsqZI5uXscKJiUvXS5
0SDkDX84ax6eXtQmbLFrcbWY3ycGqR/w1bszRoFA9uM+ZA5Medi/LxBSl9d5IjsA
nDnSGHzciCCuq4kjr6gnh99Io0kjPezGTobt95nSDGmc+lyeeE1j+Q7BGLmRQVmT
+ZZMH52i8D05VhYzmTcFMtgeOSLXwvNDj4rD7+Vu34N6cjqsfRQ/2/ZwBFT+FfOI
U3kxmj+srcTny8K/AKS2iAOvh2lR/41Fm+ykbQz7ng2JwPLIRRScylY1yKYgOEdE
zry6Z4EOd1W9NPfdRkecPWvpXok/OtF8LUH94CTp0bi4gRduRvM2H9qW5ItXepfn
vjwrGi9ZEeggFPeFf2Zhk34iXUpC6FAOF0N/KnVQ28nLzxXb2a3kX0c3aFWYM7RQ
iDlfbvVsoBjgbIdJGKRQmifJsICOOSXawg5YkOTV0asXBaRCxvNpVHpeWpeAxkjO
lYrBgcjx47E1UiOs7XEgc8f78fEoBSOHexgQg8XL249A//asvvSvkWiBFKzyVLuD
ZJ9bUorEf0LAxPL3j702Mg00SXO44EamjggGMOwKMxf0crqWQZ85muPCj7JScsvF
9pQYlrv6A2j4wdtujGWyKvX7sivb5c8el3gkSQJp4tApxMTn7cJufADbVVG1D6Bx
phJ3cP5SuSm4ECLJwLF9QdfCOOq09bhXhoO2mhTKdaUXTk1qLTDhZIEB3mqrWVn8
kb8SiByUiXIST1BCrMjBlRBXxTnjuSrXAGbwQVlWerwHUn8+sX0DrPAmXlIrn7TB
bBolxM2dTbbZehxc1faGd0pW2/qvzHfobB8SFt6QXAIPJoxbv0XC2JTMgwqBX1PD
P2BuR8YWUz6hlyId6rHs74Itq9DPsdNvAyWniBNpYjtIH1xJjbyXxy9zbqmj9skl
mPkF+5O4Ri1Sv2eZ1dwjbosjt4lRnht8o00I+GwdzV9rmzaifyyFjcv/blvi1X8f
EI8TdcTIloTQ/zUqiQhnDh1J0pophYWDjD8Sg+BEVE6WyWqCnxq09DuH+3E/KGgE
RFnQdDlUv4gZQDgOEQg0kOJXWR/W6ew/RnUtGSTypvdDPXdVhosxxqipNvIYZF3f
HRcreydR95zR4lIH43qWsxanu4EZo/RwfODc+gw1zo44KyrLkfJiMDAu47zWZOF9
ZLYa+K24yWCajrLxOepfRkVEz5heAEgmxNd1pbOnoEwJwniwYVMraxND0fchA5Xw
uFFla3hOEmwMYYdcIwmtPj+xaGaxT7zi2g7DDrVEpP/EwwFUPSRAtVCxEnVNj/U0
0DpAVkbw6GRctMskSCrKPXZjKeQ/8KMqjWx1CDtdUCQ/VBJabDz1q0aKtVjL+REO
lppXM0cCjoNVtBIhxhWJF5LCTACgwsk3oxBZN70aTdmEE4ajeYjcD12+47RNTLPi
xmL37QlBa6ui/zmM/xKXePHbvHgDaM8i18QbbnZqRF8fhFPJAsawxPZO46FSnuov
tn0rruzfKgmc0XOoRF3uRzUT5y6UdnF0AS2T/lo/u4uf3GO1+kvAiM2am20IqsB6
paW5K3d9IvADHLumQmUp8SnIbRzJlWSuSepd2wHIfUGREsLGlTmU6yfHqh/tmI/n
nJqUWlWG4W5sl0i/ka6bNk6dSMCUA+9WqGZe8dUBwsZF3SQVJqXXXDeMFQ9kS6Bs
hZbT//PHaytKY6vYi2MeFXCUOvjxwRncSDZL0B/i3YxH6P6ZKr54ySJ1nAwacOlB
Y4L9tEIlbFMTvJ2OkYe6VofuUeSsW/bSddvTy4iVR50XY8ooyDOIKlfuIRmBvyda
3wgITaNjjmCAetfdtdb/MPSPk8eMbt3PrxKnQM+hiB0fxJD4vX0veLF0/qYNI9HU
MZY0nyB0GF/f6uaFNLvyEM5qp+HLgwOhdNgcZfr6XvpOuh5By6R4HBhdNZJ9V0vM
YZTUobtU46ItDue7qyMQfS1aVSKZtpLzn3QVZtRujDsxzFzCji0XpFMgXUfku6rD
4ersYUGMCnqj7kqDLsGec+WQYsoZ+bV/BVqKV5m3nqhsWXSSccKBNkPQMr/kgfvj
6waEzmCFJEvCtZVsDRaN2H4MpqMtdvz7SGk0myMrg2yPYislkAhOc5j1ScRQc2Q3
PI2ini9xTsd5nNnXMUQRig5NGOK3/7yg6XB40sALibSn0ZIPXWKfRHn6/qbdxdil
uCqDsDYs1+oFK0li8wcMzOTQzFSXz+4GoImNl68TVA6R87trBvzuU9tG3dI9QHgl
IxDy8dGITSkSxN2m+aywHI1dEkDIlkVs2ar9qEzEm/x0va8Ko7wEzvZrh0otV/zu
NQvLQ2irzStT8Yq8LjhCju+Y6lMfdB5sZNFhxOlISzpqjcWnxrqj7qy3fPg6AS/3
3iHi9kNIezRADC9+tjjVCBLklWvw/Fn6tGly47WY8qkB0s1hksW7m/Y6hHP9dWkb
czTFbkjUrXb/HMKob7k0ONbKl+sE8mPdscYGuz2onPA3wZ3bG1EmS37aN0BZ8tlQ
fI/LY5K42rrOerRfgK8JbRarRZdLr1tJ8tAPEw9+BfAQqojSNdfy2LbmvVxZwHY8
1fpCQk6WS2WaRpTZaDy1vM5gp7dzJEEeo9RbzeYlnNnW0d/5Tnm4HMd7FvKABCw5
JHgf0glRSS+yafwqaonvSMpC9uaXmBXre0JmI9Es71WOIqB8gqqbimOGM3/Io9Nk
u7yTJaLFws06IZTrEFYhXWfY16ciMGHzbac+zsTYJHW6VrGaSSg9iwwqYWau9E6m
wFsofdW5PjFE/84c+u3NvEEZvbXFf6wiBTcCKgGmk/Ny1ji6EuA3U6iG25FmUlap
IShZ3q9SHQOqwsd3M8vKcrisD5fanL52/LEHQH38TtJL+LRJd0/W4VqXVid7NqE4
/fHL6jn9npW1LdicYgYucEgqBNmHci/TwBSYKujESpVGezw1uyC3Y79z8dyFFD51
DSNuKbmW98VGgPgsSRMNTNAMBSMwuvKer0yg0hqAFwnhqto0a6AHFEt6RfjVZXSP
i8agjvbuh4SEyjcAFQe+vVcppXdP+RQiNZrqqlsMOPaUlfNLYOuOPAHkbij6eqdA
QhH2fru+sm5I/ogeYN71pWKr6kfcMzEcGVlKyCIa9T+SyqcSc47Ia2GqbXLJvtO7
y6nj6eFkdFbYO6Ps9NOZK8LKDo69SfLrY3ePTvZpIgyLGM6P6ob7745HbihVdHE1
C8WlycYpP9LYyyynWsU+QnlVrrtwotg1PFW2dSlqQSpegujaVkgcoQ211wKGN5Yw
VEpkCBREcE3pxWnaJGbZ/wjcI9x1VaLkXZKZYbxLsxrf693kE/YU4RSMQZhIZ+LU
O6RxB5LtKmA7QzmjZ3UirNKYWkG4vB6HU2km2LIoGY+rOqA6klO5lVeuD/i8Ggv5
OOYOXycgBGz+0IjOrHeDFijh4QCYU+qmkU6eAxso+RpV8/4Jqv2WatnhWVZ0T3gM
cC2Tf+NI3Gs3GJlROYc0sZ97t15rO3T70jCcbyCr5f5EIl+v7PBgWl1xBI/bG5fk
NrTNpNxHpkLQY3ji2djnBJZk1HIy0oPWrOM95qIpo36fGr+WZ2qobUdgfVQ1aHFe
5p589LbLZ5DU9BrrjPAhtQMdoLNYyXTa4brrt8qhx9r+lfM1GCvkT0OU6t1YPUHQ
G+27wUxtFAaP+lFjVVS1atEqoIZi+d/83tAhBjwk7ScIvm7IGpcmzLfB6tRuzNya
Wt8k4oBz0Y3hhik3zIg9OijjYe5YqkkD0M1TNUx+uKqpMCFO0+wMZJ0OrZehkYMO
8jzMtssf67oqtdouLnAP8KCW4BnzB/L0PcXM4L0udmsr7PsK05yTVo7UpcHqf3sT
RgdjdfvuF9ELt1CiEifzwLA7v3x72q2aOj8z8rLIiq2HK1ZBPD85AJwgsu6khPko
Q8Lm0lgw/hfkxvyo3afEs16ZsXPwNcAfW4lnuUUohRcN+j6gF4MsqTi0axi5hsLT
ZbkUsrgyijXMA0fn0IkjumIxl3HEC/dQNbklKkuW6SMtXGr/OS4i6M/cHcmOJlcm
wxs8hyxHbUTqkr5Limidr1phvDLr4JsaxLLEPh9SLr6yd7QGX4/QrIhBvsxqFD7F
Y2NT6edMYi8G4m5Nw2OMBP8BDqcHqFstrIYIHLdvpiy79qxf0Vse5N1pcQRowdEL
Cqq+or6Ryi5PJ6hdOJYkFLhHeck8CS/GE4IqcpdomtBml4pMj+/ziBNk60gKoGRm
Q4ncSEpwBfgckfnWEn5i4vkGx3Ct3DOol0EXhfRZZ8YwCZjBBsJkDC1lTbhy1hsp
FsAgLuGkuViFOhCyLBZNmWLDyat/o1Kvb/BFpiCwnwt3Y+FuwZa+2Uz8vKs1nF9c
Cf1W51F2gy/+BavjFoHyXo5aE9A9YNIoHFif3MIJEJliz7OiK0Vqgz9KLJZoLwsF
fMbeXMv1mtcJlkvghGk188J6gWlS/fG03uc/4pDzRS6flHYwt3NbdtrDdQN4J3sL
okKgAY4/POFrIDhR4hJs2qKebsLQD6n8FQ8P/4VgsvaZ3/C21TpXs0iytlHMogPF
yu0A7rvAwmwBuv56j/kLaSBYz1Zw2GhH6I7dx/IUnopGmL+Wh5Mhpy1T2M0v5kyu
m3yBY8L4E0shxBT/A8Tror4a78QROaTHfzzZ/CeTyVMIIJzc0eUq80Cle1hwUski
kItw+BUq8QkdHSPSXl0vNQ5yOJgu/VgdVbEo8mBrrm43Ywh1a/lARd5nhKasWFf+
CjDnZUXTIV1NHsGJWRRm2Z3iMe9VoxtyDW9KzHsPCJzOSkQbpgPu1CUWj/vZiH1X
9Vnmq6wpR2f/gPbYPZVG2NbNvSjqEehIYNFBWxLtugO0q7sezbpNEzrRRUBzqeYz
coSUPSeOzoIQjmglZXstgHkv5t9Xj7WdgBUKZulDVuvceR/vkMElymtD8in6Fl/A
3q8HlAKhjfnpJ3LmGeNEfT1EcVcrI2YDvq/fharn5NxSSp58SoZ2IzSAbmgu7yJj
Q6XOXwW/b+3API2BAWjs726J4/Y/eEzVacQyfXKfzwfNzgMKvVp9QmSMWd68XjJ0
iIktwba0caFfyOt9a8/marBjH5pTtHySIZpoW4wMEN5zQXGwK7Tuz+es5rvgfjwJ
QLyitu1/YuX5oqIJ39YOCFgImeFvO3m3Z0pCH0UjP9C2PG1yKZ/C10m1AeMOc2a0
8dFtCVAmi+lR+4KmwjxOdvi6AVsw+pJxhRXpDYa3EG1W+ORzbsskF9rjODaOsOFE
jNvi+k+O9heMBlGqJapROAO9RfBzMiZFpsM00mXgQlnikjdhgvApkYDMppltyYEO
qOH5dJCW/sqs5LecHxDEubN3jhnebQrQ5TtlBJ7cp50+HrBJr+68nea4eEdUCS4F
f4K+TPK3Y8nF81hVQCqQJRta3y2OniADJwfTGRiL4ZLV8yW5hoJncVmBAko+Qe61
QAj4QM9g4BJl6vyAo48+jTtbcafxNGDcbJe0PQqnmdRzF0Y1iBivgGS3AtO2ex3F
w5dmY74wi0x6/efY0Yj5/2IKBWwazPMYND2I9NOWKp8KcZXTbjDZ1Oa1rTM95aIi
oEyl1CDXHxuEpNTLgfkZFSJ47uN1PXT1TkKlR0fV4ZYeoYJux7tc//pNmBnE8Tgw
02916AP/OpZKRXzW6d+xGsuqK9NdWvqKXTX7DV2hN1VUI8CFqo7tINZVra9tDs8Y
TLldw8Ii5POs3HKhyCJReR3jha3katdBOUAMiTL2l2yt29/sSogAg9A9KuZJJsYC
J8eq2XW0c+GeeOx9svxF6y3k1k2VioMpHY8HUQu6YcOvSPOdxUPe2zNjJmM7vMHT
LSqrGNklrAIV8fEA2vgYoAcSAofX5/8jx+XIyFG02B241u9GPVa8E58CFrLxbrZU
TLLjW6MpQSDmj1vtwbuZX5ZLkFsKECtTCniC+3VOgm3dJEHIG9FveF5DaZf/DmPC
OqQFJTGH7hzw1YBvHmWfrsojAHgqlcFp092OcdxB9LcgLiO+qIYezHQOCrq+5H3r
9FtF9yt3TQw6P4EYLztybTA9vV4TCd1kqweblOuzrcFOKBIFeS3XXLRvE3w8vEW0
DkepFB7TxoU2fBW6CvFNWocGk54144Zt+7CV7hI6xpx8g/ZbNEWFwj5T313GuagF
KEdPe5YMR+hg6FQdkfA32Hi9tGLtqCOha7VWGskOBUWF/G6y4vRySEqOG45YRA8T
j6PAJzqcNy2RLT4knxqgMI0mYmmQSl0Y0q/5lhWs4Ii5xqPCFtAFjLaiSUG4S3DP
F4hdRlJUSDJlSMAL6/HRS7FyKYtjGSD9xIt5rfpEMHXTzQZLb8cCpJIXQEdj0MFc
zYh1cnT//JorpBKZV1jvPoafeTTvGy7FkqnnlADz5rfioOsLOv0/OCJlkFunHIA6
B/yRFm99+DzceOtLvyBDLYo81d6Izna0G5HJreIki2nWSh6mMvrcj2asbongTs7z
/URP8kbW82UFlZ8araMRBp/9cvhGb7uIluUkj0ytaiQAxdv06dibOvgObIZouAwy
yI+uPROS+xP0nuQmQeLdbvHCXw4Tup4pBAhMXQX6fISgoO6J3owmnhqDspPotlGr
AvmbGULrYnJXygH8fEBe/Wex3DecGkedwjGUuz7Im/Pr9aHhIXr8GrAEWgnaxniS
8sE5/kDlCKfWWwCHB2NmcQ283bqB13vUUBHgZAyJnbzrxWZwIuEEb8aB1kTP+yam
KCKLAdqJj2F+GND4W3PHZ26f0/MclI3KejPpKMmBTvmAW2mzHbox8EkDmzJHTA88
TT0u2rfhGJhh8kCNHHIEA9+lacv71BkgeX/Csmk6nAQN3Zn0eKaUsVMJQ4T0dC7U
WwhVuC3I5Gf4adCTihD2skaqS4Pe2yH72gjRmvbigYD69e5lluUkHeeVQ4JpGNMw
4z4qEIjv3C7G8SaUEGZRfCq3utXxKYGDaEKAeGvst+w8vHidk+wJChKVfi+GqhzE
T0hyp6G93ww1HeWSR3CgAqoUberQqb/T1tXnborfoFi4IUSrovB0W6CdQA9DVlCA
OmukVN1o3hTSZZ0RLWJz6dwzlGtKYPU1siQnEZOlB3HCWurdTgmeYai76rGT/z3d
scjg/Om/l1izaS+7mn4HhR9zau+pBSfmsrFVX8uoa4Dli7KyMHWwrU83HRm7dR4W
itzOsvwiBW1PxWQRQVejpfHs44M4gIh4PqVKiQv1FzY97B/lDUzSbJ8L4TcMNV1j
A/TURCfYySReetL0tnwbzTHdQ+18Yrb1//uM620swC5KGOYfbfHF46Q5cwaBOXei
MzbQibwjFHVpZq4ZoJd5KoRRRviFVj2Wg3aSuToxX9/NDcckP5M82jOjpoyvbwzc
jSX4tzG9JKxhkF8wArtDPhjCffShsNJM3Yp1394pTwgP/bT5SYAqdhw6dUOK7mQj
/JmaaZj94VwAbU/G3jJC3dQCH2OqQvsGtrfzKG+tt736Jp02JAzQZx4w3fpgAJm1
0IW1UTtmMpVM992lfEJZZZ3t9QpH8Q75PEcivHPeEkt6SpmqpxPKwAdWNPGTCgbg
YTG7lvfe2lZl8bwJXnRd8uU6vbeLA+sUCf8su2BZffRpCRH5W89P5qemnw17kR+b
CdqbyJCmE21nCUeB3PxFIGmP3vsDqhbMDVBUeCdZ29DmnUWD7Rd12yBIW6C8SpG+
IDShh0151QVq/qWPjpNGrJUEc36Nr4WQ6bKn4PMUSx/7QFCKzjn6yctAZGw24IrP
Pr5Sd79z+c/pvRSd399rA+vOcSXwjNGl/u/R00qh31a7H3kGmoT/RA3g1GHrIbDG
eqv+3lpHKAbXbUIKMVdVtvCTqxc8pFy7haryEan14glbo4Ij/4l+5dQrZgbnI1zt
CShgnheuqYZcemNA+UXhLu2cMQhb9swKt5Vgvix4SGQDJisY7+BOfM3bYVbg1teU
OUissv9WR5pfOdLQFOC/lzxaKQyvWygTfU/beCzjiiDxWvHf5mJ48l9UQwpXf8r4
a7gZiG405OVpSz2GF4CJ6RCeiuqZUFQlMs4f14pfbJYf5qC1lJbt1Oe5S7nNl7xx
RehHKbpSNSLm6elKe04brzsetN6RkFgJl5+G39SVXFFA4mWqL0SCO7QOHyXoz7h+
/4P+Rfo9vqr+nSCZVzP60WIN7xXYQFvBMFmmHfwvxEhswc8fsJjDncAQwwdz81xr
rkiZjcZWjZ0szZOAG0nwOrtaTVTbBUOznZH8+Z9YYnvv9hXYlUj4kRnGvCKVz0kW
ofSPwNcDQTtSw1sYJyVpz8nCPrUagE3hP+nRKogCMAv0S9vDaEINQ2VazSHb56kR
jinN2n4dPFzcKMJmBEEchNfB5gKNboBATQ3rnVEy8eRkIAbdaHnjeu+Ppe3TN38Y
7DybpDQpetTUcvPCuZ5cl1rFNgImaea1F6Rgau+OY5dNOI3fuqWK0g9YVSiKIiGH
9Ra2lcx4dXFmh8Nunftd0BjBS+WtLsRZhke8jrcS68E514tU+17/CLXkzv9PLrhs
dGLr/he+lPr4IxVmPegyAg/Lm/nfwHiMQ7ykchOGURYpcgbB60Kr1ex+a/eVQq2y
tMEQKGoJHsziu9R7wOvqzSMCHSdfmhCl9YFGDqckdCruYfuUdb0duppbik+zwSr6
eJiuZ/GTsSeV84THJSllzi7/z3ta+32RJ7EQzQrWfggArzXJcFrG2x0jaTTNKTbL
XTA2jpMtVSBthM5yKHTvZLDxRML+rTxsKUmpyiSp/q3C7L3JiKHHrCWQoLIubTBT
wwfWZzmFY8zcJWrZOywFlJCpMH1bO/1GUVpNwOmYmOikpW2QOW+Sqjq9lCtml37G
fBNXGz1+5DotpKkrX39Ksq3PzL9d2mRSpgseiG7ttCuv4dGw7lLXAjLUZKKKLiPo
MkXBLD9shOUmvT06qR6M8f3ZTbptwUvtEBVdad0LmnGIJU+ZKbvt/xnCMsQzQx9D
c95CvatcJC7opNviUnQtLKDnZt/KZsBTFCXnsqQMvOKPhSaMfyNtPWpnO6gwq4pw
63mBWecN/5Zdclh1+bzTLUdPSl3io+vuaNzG9WLAhgcTGbJGgTzFpCB3iIDi1/u5
qun2FTjHvAxZGyePbPfRVQ9IvVI1TrcNmUThzJFZeKVAuQXI5peM5Hvg7TdpMsLe
thWidawBOB/MlxUoJetaAnpCwY+3IN2UB7IsxbLl+5kBjmzDxuuntYk8JEfrbE2G
TjEhjSbnl3X3Nq4uU/ZeAq0T5eCopG06IZAJrEv3IckQXl1RqylE3BED4IX1I++6
HKXGhqjEx8eNqCBiiUizzfcgs4B/eyIPWJk0sH2vlSTSAdDY3Xl9o9tnQ6gF3wO3
6BC43p67wfBStrIHSqqOh3JIHjHo4Ar77J3sC4VtUjChl7ApLGeaEdaLI3tktPdv
gP7fzpa3czDKkucmMFWuRK9l1enAJ1EJn0Le4t3GBt1cl0u4l+bdLsOkmd8aqGDs
hUoO2uFl+DGHDuWpxqYx2zdC26SPIy30dE7fOSYV1G5LrZ1m7dauaf08KQBgtjgD
zp2utyrSSKuggwhvdhSTidC03h9S5Z9hBv/JfoRifUNkS5S7NfNSACdRETLvk9AS
T+mIYfMuch9rulcf4hf5RwVUZ90FoVB+WfMwOEpolN7IBgV/ARxj/oJHbKvp/1Cm
5bcrEUDeM6j3sxx8JRhALrEuWPyiWbzmXIB0yL3tHrQl7Ji4TeFWJKnSZHA7dSDH
XqPN6Pd0VsPhxB0r0IOYvw1KjnTVEM7dgfJ2gh4YCjI/3pp+9aD5EFqRftU8+T0B
e/kRI8pHPkBtfP9h/9h2Dxjv9hSUwkXJqGTZS0jmQDhGxEInp+Q4AMhlC/MewBiT
WnfF28l3lj0pL1SgNhsdrLPjPmrz+o5EydxTtCl/aHcvh6nPZCNrfb63xjvDyLHC
3yxsGz+1fMDhAi6WHUM4D3XyojSGFf2G1oRbP0fGuL49lnRJ28gla+ncNcw7kTg4
qrKqxXNf7XXAAU1vPkbb4+n7A4sGr2ghQuBb5zwur2rXSh6TuWAWcV+Jc60LVJn/
jk7TKlM6h3peFfGe9RRelebPFMFYu9KPSV+4bcNKDyRNxyrv+vjz0C21MJ5t3l83
TrvnXjrFUdJ8TnDqrOqKBspKkOW9Y+YTIH/N9dCOzPZ4yFT5Nv8zGnfxHYGijAEY
6RGrw1Qm21/iPmcs7yDTJ2NdM6Wsr3cBoVNSMoqQwsuHCLILMvVUysB1Nd91IG7h
YHAPcl8MoRhE8HYHVxJHNfWrxApdsMdLoBQLnCOMzyOMhaA4QeAtlHv6CH8Zb8MC
w5BHwaT4RsWUV12PxU4/e2NUEJwbBRnE6drcjWZc7zT+nPTy+rzQm0BEWYcb5YIW
aauzFlsXRKfLZv3hEevd7zeJNtFoSa/5sF05NWbRX1vrKDoaK778qLbEuVz2z0ZU
5R3MRnYDgHZs/2SQ8frM4TCUqt0pCxsLa+oYa11AdnSa+qu5t5C/BHLUTSyYMnT7
f7qpWNLfnmgUhW0TnoVjoMHg9BZeaA+uCrq64p77yPVWkzeWqnpcSiOmxn6pkJOg
s1RCi5WxTdM+KXNeAj8Rj7EkSfyH/DfoiMcK39Kxc0fToMKDcdu7JL9WK2BLB+jm
TD3+C4k0kx2eekGuLBMcLHry16gXoDiHPRjieP5lRigK77hoboHUJDkh/4N8TeBE
2sLLR0if3aHz7ixRhZDkhicoo5lpXegT5k0DdBuV0yYArRA9Gzz+IP9kL4ubI7oo
0Mzo4l1CGGjUOY2rl1Zu0gUEeMCk1cbT/ybnTSS4MsscTjKkCPkSmv7g/kppc7p4
Ej6BiatQwdkzz1mmDBKMQYKpZ+k98UOzaQExvWgtZD3TYX0cojon80DG+S+FAOWK
jcjqVgiHODM3vK9WiP+Z7vCxf5ukKazOSdjMgdIxUOhQaquvvrVscEDC3TfuhJVz
6QRTKLrD/E/tRGCOQ0P/CFIj2EEC3aIdUpooCef88+UGdhpb5MPNPil0zpjF7adc
dFXdseSgL2qH/NxcL1bxz6SnFXnZ4lcm9nCPf3UhR0Pd9CYrEWE6owvhR9zdg65O
taSSz8oiXHjGhq5j2SKIpJ4h/tms4Tof93pKRUzUdAP5r+4nT5AwYy07m9fMN1+x
IJ6w/U7p3bp1JUacPKIfV2XnlxwfS9BFCQvwhWEfMR+2vERP1rPMYYW8Qpt/3xSF
HiAR6jiKzORpoWYTuPnXiC0tK0+0Ynk4hjVtaf1FL10VLeERs1y1L5Yg7a9iQrds
urhQC4ITxgajQ4EmlMIr8nFTGrm+tzFYRftqkQWJIWamQPnnP30GqnJ7yC56e3Wj
CxYIHOKxt7/quaFqle0B+wkA/47G+AOs8Yk48Cpy+wFmIm8XXbIF/NfX8RNh/ahH
TO3x3h7djgElj8XGMUhD9xj96iodmfcC1qV0lgcho3UYv3UiXLzb3yHtnD2trmOc
XIyV385wmZ79I4qSQiAMRA5DYfiiQKuEvtVNoFNX84H6hmidti1gHgcxaBxHn/Bl
Ctu1ZMp61RZPv+wjGNH4ihmjNpe/jNn7DbYuwif7GUVp4JOAdNEGSv5QUr2ckCWz
k58f99L5PAOpuLZkCCG+DH9V451+4zQJfF9aL82HbQmh1Dx/+CUInllU6mYhsAzs
76wv/7LLBNTdveWzErLzRpFUrlciWkxhakdmnGz6qPpdseefTJzqJsxDtTF/jReM
cESYhKhmqDkekvCiOUlDKPN7RkLKXQQ1mJcSaw1CILLl066pwZQaYj9T5f8ZfGRa
DtwmY2ZlE51MxgDAR19xBpMVY4jjl96OErxXs+a22UQyo1QRyjQ+ci6AjY5ygpiG
Qie5kP0ZY0ZhghWnLhg7ugbtVSvwi5XHyuyvnq7dCjxajOmF2do+hwXXAUgMUFOt
W3KnM1r1vnoQVIRSi5WLqsxDfqk/oRMWgEr6Hi1mz8KQ92QaJBi9qFE110sFHJnU
6ljlz9289MhQj0pDSDcuErXP43bts2xN9wG4xxn1GP+1msF5pKIEOZw89VFoA+AG
GxXD1zGMdcWJeWRtWPG/qpgYZOar3GXyWhrggdgnJ1i4nz59OFT+Vxqw5m+SRG9H
yFvpeNWIQKhDfgK1+0fLcWg+XrJjT4JC5Y/tZ7tEGvJxJTo4jZV6VeZ/waSN9jc8
tzQl1yyB+s2CMlfnIxGpEhA87QXnr8qgd4x06EB8wgUKe4np4q+KGhR7f0EHX35k
slJZ+MIsRUS09M2aP8O5MFsKJVyg0t2VNztnGFHwKYlIjeNXAQqU8y84+IuvN94X
cnDUyzREiy/KpfbHF4F2f7ttGke85Vds1f3A1n8Mzx0/TmmJA7EUTxVFo/anSQuB
M3S0vxLxlI0Zrj+/Ubv2TXtvrJCKu1NKoICDFqG4h18fizZ6JJ7r2vFlHGc3pHW2
9pbyxM+4wDDbZK5BtHpa86Q7myyGj3P0UojdAlYdcbzEPiOBgTVi/BFO7eM/Bmr5
V9yupeAQQC5WoV448X9bcoFmUa7cDsiIJ2PMqRDARs30roA/CzpH9kJectxyk2mv
cjzgj0AeKrvYl4M4c7qxhYmu8hHwQYDLiAMCf6IQHxXa6xNo4Y2oUDQf9ttE3s4u
PS2l8b5skMMmvrugAWzJGwLnvVHz0kTO3tRhK6WzEC4l9LSdfxb4IJT68TytsepS
zmBR8Fq9qQoFx6vArGy+lHma4Beh/LX26gi99D2gNar1RaVq1mEFSWl7HIZp9wsn
5kFz4xcK77ZkIgyvDNcUEeoYgJdGuWVQchJaAmGjXcJaBT7/gD49hTrY157BjWRz
xLP08t2qXbaBc7ANNsLWEXNAJxarYGNczPzjIsYlKDn7gjTfsSXLpqf3BktiQLAS
f5j0yiKDSHdjNGBHTswqv8Eude4BNxF4XfRP6vUI+fKDeVCbPwWeT0QNcnPzB9rE
dR34BL3FfDZ8m3thbxn+iXw2786Cu3xgtV2meTowB4MV0WPzfUSrbqviu4rC99Ha
tG0mUFh9S8+7Kgh2AURLPdl20XDMJM7UCayMx+f8qY1+oUQ76w3u3G8l73eIfXHX
MnV8kPELb1LUBL4a1U8pgV0PEXeZMakktlNURlEdRR4232hSBYDh7R64NunPT8hJ
gfr90ZYPCcoc83qRghXFHlHgGLUQBfpNiIvzqBExFB+ZzGoK21busMtd4LJWrexk
0xfjrLzAkF30qjNhkC5DQMMfPZJ6RJrVEFJhL0VP4MV1M5A/xSeMJ6UYplZu9F/A
1xF/baQU8pObn+Ib9UQs5XivlfE2VQSP/zcxiF9aegs15SjyiILxudLy15x274Lx
7R56IAXYGCcekqdv4UqQGGzj/kWt+5pbd7H6icwsTbXvsvesI0gIRSMdo7IZbLOT
iu+aWYI3HCDre0kYjIUGayeDc28MT0lRSAq1vXlDU62279iN2/RSjCrUYn1aWwx/
GY2X83KQEjzgHbFxTTHCujgo3NoetBJtXhVgO1JcUZqqVsMxwkwRZ89Z3dARFtGc
L8yAEUelgIrNYFU9LRGTjzeyodr5ZK3XehhFfgAjXGXYqY3UKXdRoY71DYzh3M3e
sHldUHVHGUpoSCUpkTpZe9aGMhNvbEc9LLqnZ83wJy5vz62ALkRfYkq8Dg1d+gyo
Lp+k5qfpHX1U7nQ9lYLCFXPkZwFDGNhw4hDnQiHPFK31MByx6QL0JerwB9fhor8n
YG4vfzdLr9oI1LPV0ykBt6gqRCfM4p6l1RYIv6Gq4via4rIkTqv5OOk0D0cQnwhS
dGbQCv4vH8g6zknGjETrW6N7GWNyJuYF4H+4LbCbVT3gX3rfymt4QhzETZVpgbpB
T1gQA4WZRL8unqDrU14AYRbEdo//y86LETIMXH3f4jUUWIxibu7MBoFruWppw08x
PIxzK0MaFK4oxFSsYSt1DTp54485lDW03OGOAD9q1/iiKbM7beY9AJ3Ylq4vZZbG
GduAzwNaNJTZ1ICbObu5UzhVjiXcnRHZ3Q4Il4kXv7hdeGaxhHWQ25NdkebAXglg
7GQnwX2J1EWp6AtOe2LNeT9MuLmeswmNgQ5OQwOt7cCtxhKo+jNdjwB8cvSzCVsl
EfKoW3tu3FZowhA/hTwxygTTyX9ukQbUwSx3u6DNWY+PaEKEHbIe3HGQNGaXqYMC
Ys02pzXFipCV9wI1K86JeGSEn6JC+G4MCbmMwRQdUgk41WKyAFxOmOyUP7rkobi3
MhItDt3loatlEn1fLYyLrNhAxYvRH+5teArfF1F7shc79JWwJvNhhQth/1VwfWHc
eZF4B53kTkcj0M1jMukRimIG9Z4LZMTT5OsphXrGYP/MAFO0b+ZABU1xbIMl17vi
27bOQN2EeVpHl298ldLUMgTi2IRqixiIfUwBgSZJRV8py2eM6NmRFJ0LiUJ1iM+i
wpBgyKSbIoxQ6fMI5KVGstLoEg+dyoDgiFjyPYThOp6tlNIiCwTm9QiYIEcrRSTq
5jm/wvm5wtAv31V++PqArBfqzAfLydwLnVhvOJ3kb7S0MmObNwHO6HFxCMZbUX2b
2eduDD5Cc0MRACQtLGufLNIuytcAfXUrVyWsgRvNCAG9jG8ST36Yfdusw8j0XSuT
sZMMjFybc8i178wtzVBRhEVSxGm0hByVV67Ti83Qza0L3/6if6c5BjZrdE+csTQ5
tpjCXwt7Mhf8jxU4X8uIQexPz7orN/dIABLoYmAONSSJR07Ucsv0z2lcDKazLfS8
G8oNw5CxWIxvpmCNXAEey1XdVP+VSxgdFt503yNRfpSUxbbTL++YBMB8OzfLsOKR
w3qYQ+BOOckQcdmEJzHgm7tDV11nXnA2/U+zvu4A804mIaDzACqmELJHFLmiVhuj
BpjqNkurmnd058gN9cz91VD6eqBWBAnAF7Cp7maq6SwndzsrpzjfrOR2tryQWxoB
WA30P/CfipOC/SCtLH6QsaLD1DPYSMFIZK21rUF1PYXt5jlzdfQOb06t4Q4f+3mG
TKVMclVYQklmxWUFuZIaqKLt4HlqSTV+lWkmbNHCOvZYObYQiqoAqfuZnXKd2XR+
XpjGKSzkcnEQBZOkGLRrMJLQedo28hQ4JBxa78E7p1DQUJVsbezk5plLi6H0iUYZ
JWsuDhrBWQvn/vHkCBCJQtqkCe9ILCXZMgONIAszNT5hIB3kJF6pyalmjc/qEgkt
BCcr/zDwBICvmb0Y5wVmSGlVA0zD9lTAo0n39UEMQ7qHUREQqVUhyzAlU23fmtpn
PCd5kLLXolBzemFur83Dkym4gJ6SeVeLsaEcN84he5ake+JqspK4G9bXWdNC9I+s
MfG0J6pyyJPFVR8kszWLPy0LLPhCpE2UXumMM+mtaeOySTdbCglV9GLYFgJb/wTj
o+PWgYZ836BzTn5Fm8gwFxv/x9JHEUHeu7LGfq4Kx4lkCj0wIGnLK9VVxv57kxK3
vbsQeaX8/TrfeUdqokhUxMNrHCGl1mKfcPYIZ6q2yo15hWe8DLqlMnY4OcJWBX6X
HMMIkwXxm414EL0YPr5dNSt3u9Cf1WBe5+PAqks+IzgCb3Rez1hdBW5VasePTozk
cOK5YwSbX+CkDD98OyoaDS8JFLLDM8IffNSgh5jo0rkYAzT1q5NM5yQxYccbLZoP
r2mhhDDsy3NtU2J5/uR2Cao/AFXujIThml68AC9UjFGSwek1UAgEgXQXwqECGww2
xq6B0634ES06g1S5T7nrxTAKk1WTk2eh+i2MWxdisjLQXcl1CWrCMPVoQzWshRUB
mETyMoxwA3ROJUBh9H413r9StxKKsKhaEqVVFpy8okTruwEu93A9QGToOzGCwMv+
46HTF0agDu69yu1SviNzs3f1Ujy9Lyn6WvexO0ghaERthaUcUQz3Eo6Eg4D6oSQG
yMaKN+6Aae9PtF2YHFsDO62cbMdVxy9AylV1DwEBnvzhvIBnDqie6XieLgWgyU5l
bOpcf7U1Rdh6lwIAIGMdp4P4tqmhOR9FDIxfrhhjjtvVX9fhzqU8tS+pcRU5scYK
/kXYQPXhbGBwnExLcrzWaPgo19yAusDYYG7N/m3wAJ5mgLW4P8ZyXrsGHRgYUPNY
6pQKMvlepI2i2sW4ftwm5vSIJaoUZwoTnCbQBG7uD4NZWPODMaF9sszsgU7krey4
09GSoVct1hLxIbb9Ey4303vxZLb9OXiRjhsFoust5WSL30jSo4Xh/GYdwHQbnaWr
vn1ihXarb+t9kVnzCTtO+RdhCAdXAz/wXod5oqrZaixYtgmSMdlA6jAQ7yrjf0/3
ol2pK2X4K8zXBpGK0Ah2wWYZkpQJArqBd6Uj3/GwCyNBFbWQxXLe8cgZgBYXoI0j
Ej7/Kse3D3oXSxwO/WQkhfDfEA6y9O38Fmn28I+rNcaqjh8QTFAqUf5elCn7ar5s
NYnpRVJs4Vq2CuHBQqHgTCQVJjMKZstooBo0YKyDiOqEMdxAiBPcMWVcW3JAau9k
EKappqJsQyFzA5oyiKpj9mYyZNezrDCrbVi/NkSaMQHJpMBs0y8WXjeweZSdsjFt
kLnDbfN3WygwRHnJrbxv/3sQvqjhodnY+CByNVoPDRVgeIsBzTkj2MLJvGsYKDmr
CDAeocaBuTaXSBLhITpiKTPo9zjGSws097q4Tz9ZXaKCRMgHTQEgM1hSGLyqcr7n
FgL5gKgJ6tuc9ae1An3uAl8yVMhkLs3xz6wROq5UyQaW6xzMxpqeNPxdLXOaxFAK
yLNarm5EC/dI6FkHDJvVbC0MkxBHAfzkv7TS0yGDVfB6ixQl/UCcVzcdXwvC9fA/
7z1HkdAkAfpA24aZoKKc+mXeJYmzIUu4ZM+tPmyGx6iOAe8lJbFe5t4zlWLa+PU2
SSv4vsWmSSjSaRYsoBhpfw3PLZZgoaTE0fwgd2HaU5dUjk+UucPAZrC7RkMYXUJh
EUOlKt2MSnk0ZkTDYTYBMYHdis+yrtjfWIblZDb0S3WqFnTMpZPs7t8S/RCMZfj4
Q6H8rHzNeaIiJVwOsmW/G0Lj2j2ySdQHDY99zWiAp8/UyysWcTCqL3SMug0+0An6
jRKzAubnn/m0DgORqbIiUNmaNZja8ouXZI542nogK+uQSeK34YzPXYavd5ygvOpv
yEbrpwxmtZVoS/4dYtzOIIfrEy1EOWPxJRQZgKeh30heHYtrGwumAVnzk2ZQlw7T
Mq1A0FgVlH32Wvk4YBXRfnnhUQYvmzwj83ggqOE0bR2AoNUEukaSGqcEXRYzMNd+
GqdcF2vxulCn1Z8t6C3c/M+1d9lz2GXuPsjds5BRtOOTnKNYRzo/9WLIbGgVM9YJ
s6cHOaLhGs+Ir9eNljOoVDlGrtdWo6gNhaneiTEAsq5KHZQZWhVWwBzUZKMB4JBw
OGqlKV2bX3nqjiRtEprHP8Dyf78x0wJonfXFn6Y5BCJLQ+NbuijR+Pc9DOXotY6h
J2BciaWbcb4vTGKd0S0qQcnXgiq4qZ8WA8XiyGe1CoUo7KGCCQMeJmB0xLRzuaeU
NKtvnruRKbqLbQyBMgO2URhCanIAZZt7NeH5GMB8NgxC/wSGhvsrChZt7R25dRvv
UUoupziWAYUxCvjVYxGWRjtEZADvJ9E0Gs2J7DTpM5rFq/wDlkoviqQAoHDLDAa8
5+1zqh8vvYHrtp0ty1POMPeeV0orZYmSbH2AnNDPj/TP/0vaY6Vqj25K77ZRXjGg
GIbpdxcWru4N1n42rbR/sINxFptABQ+7v5xobn00K2KjcVG6GZww6xIxWBFjzSU+
8t9n0AacJUYaDn2jrSGomNKvmYd98F4/WqWt32xMQkQxvNlX93U09hSoPs44Ba6h
ypgMf3q8SaciaiaWboFncqh/jaB1zzInNN1GadmuS2Xlj57SX2MnqZblx4kQFU5I
qD7pxRn9hrOp8x4cExYwjBLqzi3/XAJ7R7WNf3nznb6rXZdgX848JD23PWCyG6Oh
YkWb7G9+Ds373s+kCLkg8ptXAyQFBN3M180QdYL194dWdELwTMIVWssQyqVdjhQH
YJpyXt+nbdsW8L+n8FJ/FnR8p7QatT/fAxhElYsg08tAa+a1mEfSISzEcX3gthq+
JenpSSj6nuZKr9A7qWhsblRkwsiDCGZ+XRFoPwKplf28WH0EbYfNgM7RcRDmkYIB
KWURL8UDzS2g963EUovLk8iOHabiPXfumgyAJ24vmNrXQAq4bTFRh3hAqj/uBKWN
QEHqO4GYRxmZ/BFoESSrLLqNaRkj6kCW+KrmuElyflIQ/XybsrIVMGecDSVEJ/MV
JEzmWlRaBBU2Jz7/xbjcjMfQ90ogGp02cXUEJhBfakOwfSoMDaklY5f8aOhRt674
p9ED3Eo2iG+AGAEZmujcMk587FyeLVtxKwMEikQs+hZihp2Yyjywh4fJMRPLXUw3
usttp57W7ETxnbAr88pBND09SWodW12vPKPhfe2yM3nIcYjLmsBKYARG4WwqAteL
CfaydDTKyMC3ofeo/bzVShaM99HUqEwwIp90mu20MVWcw5xXMjo4LXrfBpPu33pE
xpnqG6SFmQQ9em85MjZFF6LSTPCmKckDvES2pTw+N7BlkpnyM16c3DfiHEhl9Wve
ToFaElVNUmNk7ApCHAPS7amM9h+D9i9etFwWMLjoj0p+tpKrC/s3y+e658hQ6aJh
0ENE+urYbVuF7egS4ep/EKtvM3RQgLV+eDXzFSlgQ9wEXMF2NRvuL5Ur5nRGFIkK
C3J3ejvF6kYAYPcIYKjf81t9RUp2soX3aS3I53dSl7bvQyC/8Oqiw2r7K2Ywpt9M
eicVLljwwVETniChBv4U1aoCVoMyDpqDIhsS/Oa29DazYtV8eZi6FFnSpCCWkpgw
gJjPCk1Orm9uvtJozOa3H2cwtOox35Ca2g7icBFMPn3pawpjFqnJ3dAMhV42gsdu
zR/mg/a5rq+PZh9Ybct8Zhm47J88z0VP3OMvPLIjNnsScH6dPgHtGjl8mcnXv++/
4lbseOQJKSTCWYVDq2f9oZZC/5bHm6oyabFaD0juzskx39nru7xwKd8sUogHf1oS
5lq29/EUgvw/31vkXq7zQsyQ3wGxwc8aWRYTOTbEjtDHUgXeC5RWvteZUicfBooA
6gIJhvo4IcvCaNIxHWzwSNg3a5sZuJ2vKi/WRNRjEIs8glK9dAq0YK8MZhXy3jRN
wA5jWjDOoEg4BDrnHlxogXzOnEfmTI9DpeHXhLmApNR+YJZpFXlePydX5ASMq3Su
HVZCErZNsVdgPC6Xk1yvdHHP7/xgzGfZOn450US6RiN86RzQJZYztA2Z4GOBUw0+
9jRU1qCCGTVMFGYDO3bccWmAfkbHERYlaBw5fDSzESDtR+AK3Na9ioDHFTP7P0U8
FueDyJbeZjdIbXqg9IiIxptvfTg60WKdpDnbjPXbWMUjP/e4ByZnz0zWzT9ZGI2d
Z75D0jSHU7RF2lyLgTqmLbqbN3CmDJEGkdSdf6GTmdP3hEy1cD8P0Oq7netD6lDa
yKIKfSGqWPqDltkILwo1bMyPwNEzdh7si7221RiMbTUuJq9JXDx4uRXXuD0NwCUq
2y5cosanjpemT3bmxQaVyqD5Jl9yYVUX7Kkb7fsHRkyR1wHJPH/hGdEODQlM9CUz
rJjor6ZNmxlBd1zUMyGD+YFdrV/6EBcvIMcIdgy/EL/UBPMdt4DNrivfFd+XinJ5
374nCOex+EZUOsMB0UCyQNooCFLh+MmBIFIoWdfh9qFFr4qSlIPvJPa09t+lzmdS
TbXxMfH+r5Pnl//ohQlvWMSvhERF12HczdR4mUu3MQcEuEJLLBWq+nXteyB1oZgf
Aqtdi+3N9jQcW3iM+7o2pPA/XEQkS3sC2Awj10q87skCq5895clwks/dmRbrN/cY
KE4JhLfDn2rZv7TZofMTWp1CNjgfkjJejbiiWZDzsvBZ8EbqnkhwnxaDu9fuurUK
ppSGGtgaiQx5zXCJUD7/ww+SfZV9nz2ZJjmv0RdLVvgOe2QjPlwfTEJmgJ5x447o
pfIft2fdBj0bEAFCTTzvSAwhPS3/DV21o5wsfAdyZpDHx3Ml6A5mB0Y5K4aLegwP
vf4x4FWfSwpdutvEr0WdvByX65GNX/GJaU8T1YVPehppO7OHfCBKooV55ugd4CHx
RjUAxAvliCoYvd4VslQ/Mb3/AFf7o8YjMmTdFuzFEO92T9KUSBihGxe6OVNFKPOc
OWiCHejpHPXAzdgd8/JTA5oT6QQg5iCXDevXVx838HMDxnZ4g954LkOTSTW6mJ95
t098lbg7pGlnRA029Rry6715PV47tWBadHs+VTTC5AUbXBVOmRttz/zbQqxN2+aD
0w9DTsh8O5AlOC1ps0xwplr1s/rLz/9jOAG3ytjsLM5BDjlmoaOloWATMk4tOZlM
bWi+D76sj223nM/EWFjX+kbR72j/7VtWS9DZONxCnXOSUUnwxuTDBngmuxNpjHEw
q/JDO932LJi9Yp4qAA0evJccoiXgHxbKggMWGHZsy2be7haFZenAlZ1SMnML2B6T
vRvC3hxoR04XsWs5A8fiYgkm/ta75qgOgRjAG5Qqj/7hEjH3XNT5cHsHpaBT7kyC
6Rg1cBmuH+Q+5EA9WzSQO4TOUkzVtOth8uXvnakBQkjS8414WwUXuPyMn3atR7Ee
LfkbrjUyOplPNGMPPdU9tiY9DHeqhVQCd+HmWgLZQgIDDDdzBsVJvx87nvOkE/3Y
xRJb0Y/jmJ/EjM5/EQtV4oD+QUHwhoAfScLL92a6oIpsvm95/GGwpwvEYL1dnP06
zO0nYs+P0ATSHLHZBKlwAFlp5+rOkOR5lL2WmtNOyKwU9BpmeBxKNFCtSQFwLWsD
nMCs+itYS+GMdVABlmlfYc1x0JV+p9yZ/2hqmE91z/JggH5GIZFHO1nwqN4j2Z2t
s6K4x/8SU4gsSVwJCepeRNYYyB3n9NOIYGWlZIDbiMUJEnUgGOfFL0mnzyNPvAL0
q83jV/E8C5se0tJ44Cz9rqXufoKRVynYUSb0YYcOPadOICrgko8NXzv1U3z9zxID
jKV9yEH1r+Hu1wWnCoQkgYihatHZ45fNXBVKwe2BDWrg2YeXwnMibDiF4p54j4qz
ZjEVDHjr8ygBTVBdbsBCnYXY5DsLAWQUZM/tKsXwGVldflT41BBjAQzOI/ngdk6S
eCUXTDsLOmBTnMgRSDwRE2U0QLQ3s2QJu+3KxeKDDKdBg6b/yDsd1J7V5dJz/K6P
ZjnrSc0iVBA9YZ1DU7/yzfcsJM0V6Hwg/yTxScSFuujw8rG1Nmdjrdiazi8yDlGi
cPhs+/WPPnfH0LPKp46gCqBLV/xjImtVKFdzGXLgP0EKguAWbNepyncnbB+SRuZD
XfPicR0P4F36JOOp2VgaKbKxDI5wCTdhTzlifLZFHIXfk5kUbRpV1a2lP1C8bEJW
I53srQ0p9WH/yY3d6/kBXkZjhiDdCT8K+0b+2Zx9q1LT5ElZk7hRUQ1ovA5C2TR/
CQccWy/48jBBf3Kxoj2/jAK5lDFh5mCmk4cuPyD7T4NuVmTb5GfT9SvBMVg/Zw3V
3CdOIcyYLWynSqxFMg52pesQoH9EbMb+iBS4AeHuviHjg0JpY2/NzN31yFkdQ2OQ
6TgbCsL4cgDWyJtfc8pSbchuycQwVTQ6ACh9NXeHZPJ15QYngAM5Gj8uYLVtxQ0P
Wo3rsHCEKIC7TZE16HLpI41cl4LnqC5xwMQ+SjK3GLCza2MTusp9L8ROWajjgouC
mq15x2oeF0qWMsjyXE3seRVhv1iUR/n9wai4mfisIdA7mx416yeYydJ2rSm3DYPA
J2BS0GeMu+QLsi30rtRoFTPyF9vCveMgSdL6xMHyE3vn2rkqJg5uLwUDfh/uN5m9
5PBgL+Qdc58Pbgsk/kt6weQPfGHt8z6g1gWmB6Oo122uN1gesMZNES/PLCCJhSU5
DXTUYzth/Rk3TzvNjCJhIvi6+nRK+wQE0QPbXmECaAkmhKtscnUIgiuVAc316iGU
WalXGVSifwDDE8LIRSYabuaV9+nQuA7pLfhhuVe2maCOA9VPv91qtkHPW5uYTGLq
OpcsgCvgO2lGebX0hdHkcSAeTV7v9hLD8dWWK6l5Yuyrn8SyDI4BrCE8inZlqtFT
1tXiKB0VNzEoYAidqEF/kT9lgb7jVK/Auj9h+IF9af+QRw/XAbVP+vwSDxblShoR
oiBldguBIOzbiYvk8iO1XOnisnpCu/pDPg11yoiX+0Zd8PlG5Kq9MwQoSB58hmmi
efuZB3PkS02SWPWS2eXj12yjAtbQwAbUknYeJXoP+hCux+8WjDqZ//TnO12Rdyel
Sl6WhJGoQt1gzp2WpiNv1wlY6u0hf5l0GJQLLN+E/21pZRB6HUS646UxADqy1byk
7MeqWEAtgX6lrLjl6V+JIEhTOIhaNZsAHabL3WOAsYrQ89iqj19vgNyQ4StgkSws
WUV9MkpnVU9xinUdp8cowsO2tT6G9T9TxN+LtyHWwifvwxCeAIO+ZZIT9I0fQep5
YOyWpmb0i+JdXJTCCaDl0eq972Z1x3SK8SJDzOP5CT4xtYCZK2Fsl5JpqiVCK8ho
sy3IWDBc/Jo9uFeeJbIsBTS7MbLSk+xQYxzM08RshboMcbRWXfLx6lxgnBpImudt
0oOQVAo12C+UtuSPBvhaR0vx0b6vncHtOYvJp/m0mQqPp7WVOzJdM7ut2FZR2L2H
zT/WdjOeGkLpp8ALoxtiw35wm1ZOqc4uX5gvp6o8svYVqHh72a6pNXYt8fek70Xf
l4YO4oQ/t6VrT1xTfcUvmO4jFWOKrZohT3z/62NxojRPu2v53TJWCwPizmYiKDhK
BFVaD13mYtgyQXXsn1v91WcimZM43DZl5Xi354i+i2AGPHRZX+kF/Vr9J2iG8jb3
T611h3Avrws+WssNGp8UBiHf9YO8Z13owKhSmgZQFaDhPHEx1kQuWkCIAn+KUjK1
fb0RCJxM8FMhtAwPvahEYB5Y0UX2iGYBvShRXWNGRTQ22MEqu6ug3xKYSuZolvHb
ntEBSHNyHIQ4gjDubcEQpzmlv95ddjzmxqeyoJtdhE6Wxm1ppAuJzR2aUPTefvsW
IhtHLmjibmKiU4K2q+iYjE86dfC4bspPnPrI+WRn3ngMDIig7HdZ1BbdlQd4grjj
MLwIWV+5TYm3DMKEsaMKqIx9dH10Yagtu/Lz64XNa8SDlNnT0tccHJVB0QvEz518
9UZLvdKLOvJx4ZS9rWe9McRK8dfHunT8AiRdRKDkGCxBGL92Z15vNns+WfTBRe28
X7j5u3sWiYcOMJspJ+lk1/HHWO9gaEUxZnbu8JnVaWBS0mCOSY45YUTBu3exKskb
tWc8zWQBxWFCX/igEgyPUoIuALrcD6qvS10bVgVRFKyTlQeEl+Vgs97elXZJOrqf
d2SSvY+vHZ+ZInYVAgvKbWwBaIXxxwy9xM7TJQyuOuvfmAx0zflsFjh6j4uQEf3X
/x3iQUv+W/4MaorAxOnJs2v6IkpR32pG06rmuERSlrWZ02DyxqmY/2g0cSJUjY+Z
quxVcJez4L+lMW0fXjW2nC1GYAmkd25pl+0kj4uUAkBHPgbsSvsMoWG2sWRTx2S0
zTqYhQ/QmTsLx4TgWXWIeDM2EJbz/llK7lcPYBJRwoT6XLVR9q+jCsYlCyXoQNt4
gGvdlGHHiwMxMPhE5oLPUUaFh0zQwiM/lXM7XQHoYijtu82i+bwVOv6dUT1Qe5qJ
OE9SPYVrUwJJyBym+TR+pZQkZL4PVK8vQzKVfNQ1R5cQnT8NkrBt3xjvAq1HzDWu
DY0QFOG1mbHC2X0CdWrsgGOGtuz+c/Tq4Xh+bMt3PnUGk/UptQgY7Pq6FyCpiSCb
VITvInCsD2uY5KgDdBKoq4BwqKDH+rJob7RgyC/VLHsy+eCzskNjQ3PAeoXhLdKw
XazOYmw8kg/3jBQ25gbtIOB4SbG/zNwudz4/cQdI9pssaZwHCXTkHhbfYGcmLjkV
F1F4/s0x2DxIY9wRKC3b6gdlqFjPMm2ckCUFqK3ILnSTg0Cb/04nc54EQrUxfkq2
mpxkcYtXG57XtDCYPkWWm41eS4WrXMq5tIwfnvCjUBLw8NQ5bFUKup9GTD9+4crI
EjLDzAWR9II74msTPuNAyvROocoj+FRhC3WQKsKfhTv7D7VN/2Bi8N/w+YD9cVPN
/SGfQKRAXDVCQxvowLdYkAcocr9TZzNBpq+vw0dIv4DTnyPWQWwAlFI0jFniUOpd
+5cEiK/FLhACj1su68LhPZvI90J+BteimIdODORvKlMRp74c4kKcu7pXtLdEXpTC
dyNlpJZa/a56VDID9lReSftGDBJeMmXr326dfQK5VwiwJxL+rAKcrmsdQmQOoQEc
y4/15h9zexf8Xuu0y3okRgCJC/47M8AkKNDMlvZmqZ9vjycpRpEh7UclUvU+WUoO
o+Devp67E9Tsfnk906FG+/PRKQWzg7WREnb4dd4HHZhGfUQHunvKWd2JTAzur6bb
4uSuMkI3ydl3AnAX9WVgFYnsO7bGtWFdbDHpxKIEeVOS9i2lDMV+9psNeUIzo2sE
ptEg5Yj+v83t4Upy66s4p3uc08pZt0aHaFZyeG6+gJEX/BxuU8iM6tiAhVTvSkxA
Vk1rtrnLP8OFCJiOodji/5BWKs2E0dcVEDvnrqiCw6VhMg2GYCwVZBtKcIlpv6yT
dhcraEINr1ML9He8gbRTyGk4dZCI74jZaZ8flNLUL7c0dYEeJDmAa+vRzRwmzyzL
OyCido5OktNnir2no9zPKlPsfeT1wy5GK87FxHEa6wGVrGZFqWCooIRe0X0WusMI
j6s/BDSQ2O0wwvmfjKGVfWIg3wMYtLETAQGPVF9mbbPImiWT4P2cmhmw6hWcAKCU
79q6X1gZbsQ3HGnfwu19fd2y6wtkmU5tmUOp6oZegNY0sW+fCAjW6T5/Ar5bffbs
+9MZuX8tlMmAHjJMIdwQxLhkjBb5vNlUlVZu/MvvY4W59KGwK04zhP4GWRnHUvmo
iMJxsTe5Wtf/XBuTgabI9Je54r3wdoG/O0OL3RmO+AYVciOgHNzEyIdRvkS57kr8
xRm2vZ+mfpFVR7PgrzfgpcxY5sigGFL/6Y4mOoDhyC6aEkPfs8J+wOhXtk+9nGy9
Dhefr9vZef5tL58ikZIpGQbJMYaN06+kndGq3+LrP7h/98vaaXdnGroLorbfUQN7
IupHcX7ezpuAH6PV5pg3BRywH24aYv2+qFkSCo7C77Jz4siyBNWy1a9tfmgkKtb+
4qP7kWpfI63MPuRQ54V0o7KHwqHVlojf2qo+Qj5J39JWI+aGHaEuwsC0s83fTg4Q
gW+/dfbF0Kk6h2UQZXsVkxJ5pcjxHg/GSAs7d3Sn+Q3cQGjtnHru3l73JIwbZUwm
MDDXr9ErrRXnU6R/HMtXundyvJ1L6rUu7f3iG4nqpwlFfADOciiK5mvFHzoYa1fA
g0oIXZwltDHtVTZiEOdYLraPRmrNQgShN4NkthRX/StFWV54decmQqkuU984qUkN
KwHALv+2TUBofC7grZL2bTjfNxkrbFB/+OtEVhWGvKeSMiHsoMAz0cWSqWxQoUEk
V+6BeF+1gNjZKuR3bw9Hj20Py6Ea6qGfLrQlm1lV2xaPonLmuXzAG0/XEqxKP4oq
c5s9RGZGHo51H51xTHY4T9dMYj7ltVWh9OHotG8GvCCJp1sAxdbH0MUxLSxYn2Ce
1/xb6jEB6XVFTQqjJ/9EZW+01lk7gbB6PBPmwO4m5mYQwdUUHPweYfwdwbk0zkmS
ekwzDmHfGu+GyQpxXWFJ0uaUv05WcN4Avrwj8pzEHCvTCtXJEiiyBZk/R6FNEuKY
k30RlgZxLprXcwkoU6Bw9B+2e7vtbGNe0PsMKxMLUuZOO+maUaYh6owo+DprSbbw
PIn0hbLSe8Q2lT02ewJJ/cmEtocmPqjpmaiO0sAVSn1DbSLeBvKq4vFhyrIsS46B
bk8i2N+efq+MV0gSXrZBG9DIHP5fBWabMT2m7gH3IHBsoyxJy3/rT9nfw/qEuE1h
6DO0SDo73Yp60e/GtQHdpxRDLGQZhViF6tinLpZxxVDmOwARClCD1mHUUrO1I5/o
5oin+6GjnzewIs6Dl6LG77yJMToDMT96hDY/axFUYDw9/SLJAa18++wTV8akvsRB
Ze9M61oFAAwSAKd0dPCGGgCC/mnB83Bz8P8Ku/mVIX1OL4cJFCrSwb6h4qig3L5W
CT69M0LcuEMgimECv0ir0ztv9Yaat3uysb9B7q2I3tqla5Df3mk1nY3pkCWOMTcW
rNkF0mnutOWOHvsnId8iwwRxGzJtk28p/qHC6pQ6hOfJtauwnUICC+CkW/DP4AvY
BU3aOQsIxikfHF37X9d7AKvTz13UiVT5VsbwRF55bmdp+kEbcOEZOIrAnmI3Yrd6
t5Yl/rFFeuBqWAuVAujCmlO7jqosr4Babka66AijQ3fqYjaQG+24jrR6dZ5ID8qE
4LnT69XImPxDwDwqlSQpyUTm6t36Aj8KPui9KqJCQpuaIGx+zXTl8VN9mtDvygGT
c4dQWAEneYgw4flk7P1rkdnpeMr8xoGIZjFpa1DmJ+s2Hpx79Zlb/BQDvtrwFbpl
hSEg68CSOdT0deyYvNxSK0du25oJOFs1HFn4pBLwSCxLaJWqHGH/c5iQcj4UKAZj
NrehogBKmC8TtVb0+fYBvE9YHmSnM6mlykeZ0KQ3Wq0V3jEVn5vO3v+REyOoEIwN
kdWp/ACZpcI9+dwI+bN119dXFFJcikP+eP4uhHP63BnjLtx1VgbtUcVfEU5IrARY
UZcoCZzSypryYiaSv7LbTmI2yGGLjkp6ELtnKBgIg7Gg+9hLOtjvAIGxuEdsgeCz
kik5BtSp0vKSUB5mZELhcnKRvvYf5AX+fySYHi4WdMjUoT3RgW5a8UoPkUweO0xH
/TibXuTk8yhYdCxD2foTLRgin7vjKuAv7vVLBQutWbyjuMc1DADY0er3xDujnpid
zd+eXn8O8Cw77yYbBhkAAXGRYtuCBvOoC5BTEbJjNvQq+WVO7mjxfrC12zUJoP5q
aUZJaTNH2bBV/Qs5LEJS1EFGdV7rubrzBYkoxJhquy9ML7wssW9LLTgLdB0+VA2S
4dfEBCy4QfpT0kK6zthelI39wxU7AEdCxnJuX57EZxgVfWkBOs4kL1GPhQ4dZ8CZ
PfcrRqAk1pp29juqU+9qzSsXPHOO5soASs+I/8ZmvxF901rHyUkKfgQsiUYagQt/
PliaR3EdvvmHrzINhHTnQ1rdSU9ZF4Bnxay3o09W1sP0u05dek/ZB+JJVCBnaNM+
d7VTJszSdGPknyF8DAvz4uFffVhxLtc43fR2xQ/DvIVxNicdWBxyPEhqANQjEBIZ
uji7AuEqrBHs5YQh+9qNE7GSfDeIz/QMAmBzRsnco4mw/F82XANnOu4uOOk0qr/y
SukdkGoYaWP/5BWGPfLsz1dhfRoKIiPuA4YN8FBpxSh8oLPY5yusl2C9IW3V4YAy
qNKs0MmspGmM6WHu5GM9WKfZoGNpiyQwrtE9hVpHzllKd9zhvUR0R1oN+5VVbij0
dcnI/gWO7W0WbEWXVlihIP25BdTzhlT9tljTWWYv6b3WRqYDlpbKqWZaZF8pivqt
GxGZVyj27XrxVXZpHyo7/XEjtFgGA/bdv7bwOZtwlDwE16VijHo3YHVDQ57jFJij
GlCr8Yl3t/rNHsFiu9QJ49rbicFLAQ1m7YddquTWQht/2LeUhnCtppwv30diEVKi
w+9TKvsiR9r/66fzeKIYfKYRCNhdhQ0MfhO+SRonK9PaFB4w6s3MbIBFeT97jzB9
G7yybzXyujIxZumuqnbq2f4t7mUFP07iGch11qYbSs0ZA63lvvVBx4OVXjBjtVnO
q0PBaSmlOCJ4pcIt4a2WdSE18rdAe4HIcbVguqZW5S6/aGcGJk8dkmD/QyDlpwdb
Zb0NwnXnHG6footp00aj1rdjVMaIMv3f1JHgaZl+Kf4+A5X5ADxWYWg53rrCeXfI
c3+W/0BuHle9aDUuiI8O+PFh7rY3GxZhiWH9pmkCnWUPfJfsvShqvvA/yzCO+aCH
oZ1Q8JqRFrOzNg05R9kRG9ZiPrXE37PWGueiPFPgp01XrWjhaYufgQw5cef2MBBJ
G7fDMNgAc2cONXkqU4RAHqlZotazGfnZzrPqZag0EAtVjx1nQ9xz89dOMrvOaTjZ
aDwPRcKb/pQbikYG2/ttQfLAAphlcLTwc52aoSdwg8znfOPsVQjaqyOsLkRhEsst
bcRVKNYpD/LgtuE5VAI2o6riPxLV7/HB8aM+8QKmIbk5uVX62z31StOJZJtp3+/q
gsu7go50ptLxWWqEFJvm+Nejos//D/LZjWfAGCWC+D7nOR7M1g50mOqXjiGNxUAQ
GDf1DSRGYZSZo0S31RBzSczoGA5rIY+E91pPgIyIhDsDjMxCPeTw5keVQpiBX8f3
CdYswBdcukjFDEsGaTBKFiUhKazQQv7YvUBnQqhZRLNz2usvdUV92vaRJqMioSLN
ksiWpuBIR02Reu6ptcUJaS+T7rujNrPteBVpmriOraTtfOaIrj8O/mhjWuG9HedP
Ba5q28eVjI5UE2xXhSCa2sFubvWHd4Dpf2ysgP4YCc5HI47F6tu7sZt7BTnVSGUv
I49jkWoj6Pr5RbBpZlBu0sDmLR9MhCM1r42haTdp6wYLGRFt58dn4kw5v4XY0sY0
Tu7go4DX2roJxJdjEoAExBG7G4s5ruLb5N1DBhEgTGH1dezg+daLZwOCferLIWWh
VQIMctdEis8fC927cclzgG9RvomL/SxP3CCVj3OA6Q34csTRq73aeH+L2Dlsz2gM
/3D52HRe9GMjVLzS3XjEWNujJ50mf6272hg7zpRaozdqxlF7Brxp4hmKzrPShOmy
hHCBwdsA39KcVbi6nLD9tu4gE192mQSOVqb4sKYyz/TskIIgjnJF7N5tyxmcl5in
n++bWlbR9xNqwZVZTQsU5aD05Jn54fw+ZiTh18DgNMEd7ifJH23l8do6/tBLC1bZ
URZXWYCuV/VCX4Q4IZwjDHschbaS88LGagboZ6X92v/BvfHBeGaYG0oq7tvUjKjL
LmvbvaMly8IpYHkmt3MXo5Dx1DlUhpi+Dsii7DPP33zccBiu/FR4O+/oNc4wuJJG
CFimRqk9clLSz+MD/SjOU0f0lyqtfKUSeH5fg+HqwvsPm7PCbD1c5tapk2u4r6N/
wUwgwQg59EZqKNgjgVv/tei47fbeJN8sxyOGPFiQYZ2GDRpP0z0TcBo/2f6eJTVj
DqsnO+6eFUx5W/0E1JBeZkxpMIdpgYPf0RmUPLEKTls3zsgGfU0DhIHjTYJwNgex
l8Pk7Rg6pC1K/p9kKVI6AE0FDNSWpgVg6gumpbjssI8kC5TVpqY70tugDNRfLjCX
5hakjQh9gOocX2N+tIGX5M27IGltT1ruwolzMMCytzQLhqnvS0gprV6FrC61hZwr
zX+OqZxpwUOtK3DnzSdzvvE2c6aBhz8MeFK2waQSJe+tR1U+6T2MSSlkTKjqLqFL
jrBTSGgDz+pObnSMcu90jYLUFMyD8kVS4ygVheqhpdI3xqpFmYQhZ0AfWBhcO9XM
8k7bFwfucSXYkv/YkPH3PkVmJ16aOLS6jt80kI0+Il/NvCGT9/wu6BQl2ZU1Mljf
p7M2GriMgsAbkfOvL2sm2wTN/hw0Pgnjy2e2yJBg7WnXHkOa4JEd6Ijqciz75mCV
2qRm1L9hbRGEY/cvLVDaSqcDwSdh+JkTKjAqY8sE2GaZVQe4WJ1sJ6rJBmoO13z5
dx9DuM25BmQQvlSD6ABHjp8xv27Xuv6I5g8oE4ANoMhe8F6i5aXa6Xc3ySG9+dR2
+sifa/gBhvzXnDJ3ksN6HmBRmFmWVG3w74b+fW+QsZAArX3o3NkDlgsvwqskA3fX
t55Nmu/Qmyq5hhWL6qIgZveCk1pkbfvtm5OrJvvAYif+GFW939NNsjGVGIieJijh
t4A4+KMsiwydsec+JM4MQtOq89Ofe+K6QG7FyZrhvEj/zZvZFZVpRyQprHWyhwr3
/2sgWW/ck/Fx8S43fSIPYPkg8toCO0OtmimyP1jZl5pg9r8OZN9vqQD4iokv2mZw
Z+CMLTaIqvFCL0ud0YbRi0WBpMW0vazRiW3JpN8RuS++Ejd2qtoGx/+TywpZqF1V
fmKPqYyYODeFEYP+tXGXmS2WVYOScq4f+ULkcTCYWKZzxYyQohmd4tZphiCjCD4q
P7zX1zBMOjglkyC2RDvKd4kwuY0hbY1HfSFZYroziuDPKn2FGwAQ4p9roScqTIci
BIIjAnAP5PHr8/hmSt1W8AOPxgqNxvZfC2G69WMs+NK2Qvrqm5BG6OQx0Jw0f6fg
iDZhlWJmNtNzdjqZSki/B1iWAmr7h2pK3CrfN4ESK68XnUQ5yS2NSIA8TtWHw+SU
lkmqZHZWK/aA7PX6pN7R44vyi9YwLKf5L8cGqZO+PkY7zr8SJuzUlRJZyjOKL83J
t3LziMvk2e6a8du6Hyo3k/hnyrg6Ad338XimDVURdiDdEUy2eee5lL58ezYDuBfM
tarzUidicB/xeQ1iUz4Q5WGk4tRPSxrzK2jLJziUmjx0IKNiv+HWmlag7XIC8TZ/
llNGL0HiMV1frHq2r0Vh1JXNe/vRLRsyggEqlDz0HFXagglHMpjhF29zSXtowbhX
FaMISyuPzmf3P/dZ4MzgJSn+KFvIH75YJ86Ni7lmvZT6cf4XwIcu9w9gEEpJXQME
Rj7Hlhe7SRBMdGluPFoGx7TE08wSSoZMzWEpej6xMkK00j/xLNYQceooDr6uL7gy
fw6hfPmi3ppzVnOB5UoEHSeC7Nc5ULYl583TfSG8qEpGhEZdshlxp+1ju8PNsLYP
9BNlTvcinRbltjeozEsrBqvqEm707NMpjey/g7jKcPOisKHHTqPclTPVlzFMlME/
uAA9zKcCAmMllujOWZOQ769M3UGEepWJdfsUeBvxtm7BaUt7ZGbRzFe0XYINNUxp
zYedzem1WEeNnmL2koyKDFg0S/yUyQoIqBZMMvLsl01kHenUfEZ7zmjDMAT22GKa
6yleiZatS5rVO2FWVVmh3bnkuU2fH8OhOvqiFpiepdasAiUUZ7tfkgl9OQR62Ubl
7tPoF+8000GYSehhA5Q/mgNOWE8pp4RW9Mlxmi2hM71Wy/hj3fCYw/VH1VK53Vz5
xHKXys+9yMJRruin4+5D9V/prjL3aNvXaHNTSXkAi/KFDQSlzlSqL+jlTTNTqqOo
fE6RfYaOtq2v8zdEX318KX0PCxgMIwrG2Wdh6Y6tRk72QVbNYiErlYg3lxo72sBZ
X88TKfxJqTtJdVNzVwHvnKn+jM+MQv/LwuyzBTmiaeAg6kwT/mXWP7dPZaVGQ8gD
0yGVqpoPwl5tJjMSDRpfpUWmJoc9TxwSGgZ0/uHPSSm1FGS122sBKMknuDy32rJq
wxkviKgH2owlN4iIuOuG9Yl0dk4ytJchFO9W7Kfd0GqRLEVYRfVTFXYI93oy/Quw
Fw5QZ46LMSIhpGISO5laBKKBOjtW4GHPZch+R5J0gWhh1bhbutIhcw1aYnISrxKZ
2kcljNZzTONKUJDuCZugx4ArQtEgA4TD07MUSHgNSd+DHE7c4nGrSij5R8tfVFR6
AlLMgjPlI5mOWVub7TajG50ogoXq5t+bmxAJGXL62MJBJlgp2/CoGspf4mXBwoEm
vWR3uh6s9mrk8Nuo6paEihWDyQgyqC1+oCOm9RgAXWKcroKX6cKXkIi8SW3W9+ax
SiGc1j2zwGQ6RnDqKM9w04MAq4ejYeynwRe9Y17CtHv4n1AEvWBn6uluxRPmTGHa
Ep3Z6QxFO3pwOMnqOUaYOukQc3yg1XT56TVRdL5hv2v4ZJ96J4AwORWjVX6UD2SS
neOnMfQruox+VIu0qetzGsv2N4iBIUhQu3kzEzrpwj95JLhq0P+MJXrHTCfiZRTq
e7O7/8+VLauve0hLq8UoCOZ/+kJxoAlpffZ2YF0lpg1Q3Bts3lImefei88NajEJJ
mz8vcmr8eoKwE+3WPfhsFCLP/Jw9VjOniJCie0+/91flKqX4GMLwggaOo26xHrTa
GoOu8ShPwqvsJapBCXUpVZGeeMMt5Bpsc1VJtIsaXcDTesvvMFK47XPFvaPF++fR
LhwMo1prDYoPsA0VyYs0/G/m0VJ8kL5aUMSC1K8htpvBKsd4u5qGxBbmmWO+dPpQ
JYWA5mQXroKouU1ny/nBqoCQb9QAgFoOzCNMhIbrQhLO72sf0bGke7dPMDtcTV6y
W6kPPjXw0krW8KJpT7VCbKYheI3nDpT67aCHBgcv9r+Wae+LunLrfhKKL3Y0VgmH
2lspnIJM9Mr6+PrrLz/P368TixVykeIMUtBQVZcK9uKleXNVJwjdObaG03pmd+WK
khsUCGXRftVxgMtxk1nfZsa8cTv4WFBVpV2EI3qPEYMa5LinGupJHOLl4Ru/QJ1l
6V1lwFYhOV42NF+m8FjTS8drDwHTW+aiM0/7NbK8odVRWyfBgVEB6Gsha9JiUgZ8
JoiYhH2Zl2gDzJpRz/dMSQQEh8XsMDaADa6tdh0I0BX9e8qvdFK0ISU1ChvGQj+s
hTRcH25IJ75GkqwQyXtSXf6I0iJecmGizpA/99OHMfMVWVqKy4BjSRNljDK1NMJE
YqVO5ymZfvOL7OQUf/JJ72dWlKkSfNGgN54/gZDkNA8L4+cigJhT0PpcegpusSfD
wdzebdowFiw5KNrXcfC93CAQpY7PIzyuHYuaD6ezPSncP81hh9WSpshbdtVMW3qA
1+sZPIyouYDIT746gAgJEX195Wq2akNVorYSY+Empf8G8DYDV6IJAOLnerI0KUSF
wFeAszmEjXMnZmkAeffn5ptmz3nATcn1nwaHj8C+AlNC9lkYXEBoujg3NY+ePCY8
dx94Jta5EsEZNFiqBO7ZEnbFh2S0oF0Isx2ejqfmphzkmOssjZVhDda12BlTPrD0
oXPnDPewUAGIdIPGhPhzt/hXX4t2JQR0IMbVzoTS6wpr3g4VFy0l67+tna0PO2iv
aErffTpnnKfVnpD9cBaEx5IYFJODSnk+EtW14kOMbqZTLkNxRXg+TbMAfKr5SMd4
VPQBFwxWlxH2PkgcFteVk/5t1AG/b7hALuRO1MmnyyioIfXJUlMHmCeW8nvHgZRB
+7lMAJkALBN9Mkilnh6MALbRojNNclbJ3aZUe+90r+gviWOvMrA1zDlfsDAkRS95
gAlmuNAAG3qohOoXxT2PZAXvIE1MuiK7rNP/AcAdWR1Um8jN+1sHOi4Hus5TYQAp
xywxSyLpyCtndZb8+T3E2KFtruhoTUI0TCktrPDigaAe7JDUEAr8dZjzXVj+cuQq
vUVeV4oOkCSyOIae1qZC0D7PfaV4cxsfDJrPN5Zo8hiGFjLJg/d8DWbUMvVgrnl6
jyos0Fo6g4Cd2/+jKlfArWkYd0dbfyqQwvr3n2CL3/FUECrWu8RMv6+Qwq+vWmd5
GWPKmVNjySYqjpbDIdmmUC23mHMXAs2zOLEq7c1nsnwQcqGvl06lAuC9Z8WCL6pO
OmK7rAtCPnnoSiZcJR8P5/hC5GEqcCCtZ7hs5qH/Cbp9vsEyZd33W561L3icM9Rb
QwJqgQWNxxfGjVCvj610ErzBsxM4bAY/4O5ju1YuC26aaybuhkmk65pU+zkwUeQJ
EUMUxmjYqWKqFX+buga3nW9GooqJPr0C/wqzyqr/AQCoI3TU616vdo5ktDvI6+n9
BbpBSkHtJYAAqmxscC/ftZjqWD4mqRP5aq9wGDPcHAek4R3vyGG6m+dQTOaL7sFe
FuWJ60Ueq1SQRl7GnzYDT7ex73+QX9wVZOh1at3nF61iLRxeMqDhpz/z9RCPaEAJ
P6RoIulWxDn3K6kHUbSnQ23s5GUWwwUp3FAgE9AvjB5gK43Pn3qPQneK9N7+JDVj
L+AMLNHM6Kt66gVJEqt7T5ao7bTvgYKZ8mDKk3dpbZkj+YMk9Lx4sgubcw8cHyv/
zgLogXwSn+Qmhbu0TFXiapvdl3Df3W8fMkHjch6ZjWSzuchuTSCmSDta96QKNjxf
6QxhsE1I2dEvvaUxY67PIlbUeI7f3DYmpzMcHXI67MTx53NBfUvjPaT/IhTc1WL3
NDf0zqgZ3xDTUPyDZc8+YIIGEDtsU4b4P6i9tJaBL/gFxoYM6+wXOKaBHgt2K4KR
kNaA053Rvf0jkBVzYNS68VR26DjxCknz45ry/vbZd81TbXevEYJEmbACyzJ+wh51
j37meIyw4KsrRPT00FM6AXFq9tkNXdGyrY8zfKtrGvXkUXBxHX4BM6I4+kpUA+OH
pULPjhXCAc0a+sBVqOzgdaMZHTFK+HVTigLOlqaQFzPfruj94/yFoL+6FcBadNfB
euOqZ+gKm1+xgUDbZfl9lY/cQLrCBVVlAxlSKPuykQp1e1eBJI0RY8eIOt02KlKb
etA/aSFywoWOCfHMFLrHeDmlt4aUmg7QG8Xl1KZhAnnP10TleElaKoctaTSIlFeo
kmJquEECNh8XLpPFHvxnBeYypp8m7QAyrxAzlfgxVXsGxq7Cg8O15zIZKg2Mehhe
fuGO83zo4gVVKZvGM7/YYnm2mqe0aHbPoDd9iRGa1FeHYCu0HnAVO7NNm/6bq4Sz
7dyGPlvooOHlkGn4ZPmv96Tynb8ctCjV64EDdqWRmCqqBCaT8d91cF8Vb3KcL4SM
nUMdFYMq3saymaX5FRTwk4Q5I9yBD9xDsqcxC+/il7neOAzUSkXB3sc6X1MM5tzP
Ia3Pv9xPH2ntgCKdTDuXUGQawO6jIlNZAgc8T+rlgmBUawHNfY4YCjQ6lt8CT+OW
cvtxdWTtPG82e+kVhknspK/QDnFVPcftAM7XPnUQFjREyuKAIXCIWXf+o0H2IiJR
FtJTNXWO/3+X/kJueiM/TSbvFSqtT0drcYr5W82llWa4+R20rDyJyWktmmYnxJq7
hIrPFDxSrqticP86NuQhwcP1EyWijS3/QqP6YjjxlDSedmGVIDKxeT/4joggG5q/
W/XrQcNUjWDW5Su6xhPmSHXJc/Qo+yvcLhUaAh4/8ny4J0qxTBOXchxtTwrq/6WY
mSFC3fBVehOWEP16wsgrXkjbgtlqg0VXn4LB9fxhkvW0RWNis596xE0updxLh4BT
88mu7yUEGkkVFEXKVdilYC4RBvQPgcj5P9FBfpj1QDIijWdT91X1MfQItY1ghlP0
n6QKTUeGRL5rZh0THfkm+oMOYJ2wsMjswGYyi6fBjR6rTXz3MUzbLoaS7GOL5mML
qcHNyDd5xn1OVZkExEZuLpTw8RCyNHKRONp02Vielm0Z3inK9QOwAdAAS28NtIuL
mbDKXOsR5CEu73FtkpPbK/xceIgGLPUHHPQZgIOe0RyvS+XUBJCkSTjVVzlSSyqf
PXtpNMutFk5JUQecAaMtk57wfeCT9kfIwc1/UgUhZTPFXusnPWJaPLo4fn3ZAqnu
d8qp0Vg5+uAQ/thhUC4ov6WEN/Ji06+ooO6RKljfnqjrHpzUmtekNnAmKpdtMIau
B+ycTuo9qd92TinNJO6fAVBQBvPKi/AEFtoyN/GtBRWz4ZP+UPxVGa9beWrynuyL
9b9HJp6UExaluiIkdUQaciyRafaG78cfzgW3fnk22alzCfQZvXklVBeKDL+NJEFy
kfyPTPvQq4v61oNOI++1N0ht2xR6QadP9Q0wg7voPy2zW0CPpE3j95G/3nExhqPy
6rrDcnvVTECy7hTPwwelv58+tkPCbGa9egAYYjbghb3sJpPMWmn391T3G+8d+0Oi
Cr6ItQ6NCigLW2kkY0lr7dnfVZ7RmsSLysnnQxdlIfqH6WcDg0uMCg0D1aouPoV0
go5VVUbK4BoznUfqV/38bII9sStbf37LkD8H8BgT5QcWyCLOJ4B4FH9aGjBsuO19
IuJPEeMfTrOtdpf1IbjlJu8AfOXHtpIrc+tTc1Fe7iq7OSWtB2OgcozrEBolitXd
48hbK9I48Uvls1GyRTrR9gU8rJIy/vXIbobUguH53A7Hq6iOoFw9Wo1nGI9L7kgD
7JcFVRw7YpIaZ9yJ1Xa/cFmZL2HWN+MdJPfocPkbbepONkGvJRCqikSEsk6qWHzo
Fdexl6SYeK4EQ52mg4cVmll3kfSD3um8JoDUZWEGQixO1kSaREKXyn8Ka61TInVx
Zn8tvPKtFREZKiT2uZuYUlB660zTlOUEUljjDC0KMpvzCzN1IIfnRbNNg3NCBNh4
73MHNvhHi5sLPJn3+C6UEHnIpOeROiDTaiKPzz1BDDWiuytgqE3dXPI62ET+xOnM
F/yjZAmJBILcvtuPcZJiDGpaK435eRWa3O7Zv+oucRT38sNPiLEKTc8yULVl1z2s
CXnckGN9IvSPoj+XvJ9W8hCeOroc1QIQSbkaAdJfnk1JQ8pGmHch30G5B7iYEyfL
L4CIOxhyrHbzsY8AiCpe74QLE4ScJUi+VkWdKBNTFvyOfIrHNWLkjPn2RsR0S+TC
hndXi+vZLEJnjvYShJxsaBq5KGkdZ2oh3/G1BQSZpmTdBr0gv8FB3guPcZkih2vY
6vq9f8q0c7eIDkETSdMONm3BlSUmx45kjPwfDfVlySEaNSwn8fhTY26C4TmHqsSM
8jlR8KwKd+2QY6Wh9dJ0p/1iNG7+zt2bxAFSCBaLGfgTxXrHEioJtr82/ikhBbgW
i4TapJ+0POKr+32ycUBghNV5PNJ9agBudkS4uuXsM2WDKpc9NPopBdPWwSPScu4o
BxIJWrADazxdy3Z57bmaz4raJyTwYBn/4kTGMtluXMEUUoliR3pgOZ+4oOJOHjXB
u5ltW/yAOjFnDT41xCStOI/65IrRztZvETouQYMzM3kDXUmKnkkpd1Dtom9X7Xt7
k1SGngEwaO5mLV0fy0itIFq86I2VwSyUdPQX3WAb5ZZ/hwV6AHzuhzcyBVkANzRN
EfcVf8G64kMVnoP5fvW7UERi0pEL+FercwzX3tGtx9KCuhnynkwjsTbCoaNTfxJ6
FJH94LGCKHDNF15YqVI1NNl5J20K4wJ4brJBSWgkUIhTtLlRqElWHQSS8sAcQEHm
sXkEGH+0B5/s2a84SmlqVOh7KP9CyCV93NLi0RkOKIPfEi3IF58o6JHDGdpOnMMo
S5gyDvHqcqvIHdbd+qunf4D+wOdOZGq1hJDLactg9XUUt53iAtJZRSOME1zsmlhF
IYfbYSgGYOgdJWaGzeizEWUm+8eT2nTKl05lhE6RqGMFi98Fwv/DhH/1mQPOSxBw
Jl0wKFpcNqw2hVF3AZJbIQ41tWmCq2COpC2OHa4crDCbDB5KvtgQjvsT/uX8tBLB
59AaFquC+dWFfa79O1FrKdizczfyPqRUBsrVR3j1lJXVP59za5c2VZT7MG90F39O
IT57BnSA04oz3IDr3/8PE6ty2yU50sIvryHodq0Hb6Fg4zvaTaky7l4ZJNJ9lzhd
kQRtJWVVdZ8x4c9Yina5Zvao41ygbC8jBiv9wdpiWGGJX9zY1TJPxSqSGIiyWGD0
LxPMmD3SSQl+0A+ocJYVhkaPcCHiXIdxX8oX9KG6shwunSMnIf+p412PhgrXsAWU
D5myjlnQRjsYVldrAmR8YkEyF8SLIs9TrIqgfMsDc3qGv1PbTGE7fKgrY3tY1cqJ
G7pHsUjrnXBzKbv96BxS7vU+B5opBEw6DbGUWOD4h5Oy1bCKc9mWV7H4GElMfNa3
JP10rJzicXSudX/RUIIvhvP/uIKrau9y4fV3Yl3//4p9ysbcN2EY5r0t3GRxr+1v
dtPNc39g8dY7aqO8KaTYShsy6mE5OEQLyzhXZdRt1NRJAsgKPQ45aEgT21zQuy/p
4BeygrDXxWbFmvsC/UKsalNV8+mO+kIz9GywAmPoVP3vT4nXTjSh/YP+3uN/YPEF
b6nZYsazcFUE26cZyYHp1KMo5I2Cw8EImKX4WMCd8PRH68/2o0HTd9wFnwQ5HFGl
4kHrNhpM/+Q2uTI8CxCh7VIW7xuo7JtCyewHY3xxQM1t887F2Tv2BTN1lfCjY7M5
/1TMPa75gZBa/+E6Xo6jJ3dZGVHKtXwoRXsz3uSG7jbtoqW/vvMazLHHg4hBSF/X
zWALrcfr+fr0wGc6vcBpJ6t7asaQrzPXFenaZhsUvFfE/boSvCUj3W5NFBGpR7iY
Uqcc3sXKyChDL8LQNSf7j/PMiseQoYl2ybXzOoMPO6FnXhsSs9rnCuJo12Dh4piZ
axzVFnUwPZq2c5cbu4pNTORvyaK6qnd1qq9+giDEcMrvap8Wa59g6e4FNl4YS7zw
Fevhm7DL2y/KXHpYty+HcLPayHfbhwCWsOcB4r7n6daWMmJra6kAZWKgA/IaUjGG
n4+v98TJzEbR6hbYY1h9PZtic29c+DrBpTYVErZEZmDG9TTB+q6YWiqk1uclooOo
eW2eTQmI/x+4j/k2ky4pXwfEcggRvKS/kxqV6RR+bgA1Rgh3oe7+o3DPioaB9yzx
wzMJlYebeulEi33AqIF2PU/aVq9BsfouEIy3D4xWxDPrLoS2SwS17c0czkmrBq1N
lP/btVZ2SGzOhZ0JeOQ6tINdAh8dA8kn8vycnn6IKGN/UhdrueUQopGkTNhv6kCV
vSxMyt3YyH5JRSiGnSwhkc/g4W2citXNExb5HgYiwAw8endRwAVzuR6Cj24eN6gJ
HNKNPrtfuZna2DQy4she1PyyerWuKWS0UgV7xihNH5BH2Wp0V+N1ADrJUKHuw/oT
nZvff5/3RhEQnzlpeFD1d8Y2t54zSyRQ89c4DYvI7HY6cB+Vfzp1k5TeV0FOAlNq
R8WickcvQvRXfcbBf081k8B2EHGSm+BlSK2V6zCCKdb3SDc+PUxKgEDcsKGKNgVP
mZNqfORnggMEHNHWgOEwkPFY0lhJzLlsCZKBx5V96zvx+WGgijQSmMsIEmPhS1rg
Zo1IOUzJzYdRKJXfwTM9cWELM1JdQ/OhxCQ2vaMNzTFtKkB1A3URyl8QWdJwE7cS
llnr0up+SvZeZ1Gh0WFjIZ5stRpYlfxd04IjpmusV6ZztZAiYo904TXRY5efsak9
lHy3WC1ek6kMoyuTiC6UJtTBbb070p6Zx699V/Nr97TzxYtltqd1E2cvZQ3C2iBj
hDX43FGlPvoB3pE8LeDtZplze9NhU6PNhbOEH3xxlaMjWbmRq8eRxvvaKARDiviA
EGH+Dd59awtCA+QTwgd5/LdMiyjB2qJjrsKh6P6Kw02BNBPHGKlImxurQHKfxLxi
+55OkYOkshCzWNW3iAX5/QzkuDTM9irjcYcQYhVMQnATufdcVtGr3A35CLUAkqPE
3551xlYGJfGBqLLl3/kuR0Alj9JUs/IouIhPSx0Ls8c7g6k27bRNI73HV/sku3sF
OEcm9F5n92dqsd50QJdZzuq7SMv8nPzBMD9pHMIVS+RRZgfir3gMhg3IzX7SjQLY
kuNaVElGnU9XptJwqIvYZJn0t7pKTAgwEi5XBZ3x2btmugzoikH6Vf7VOmw0s79Y
9Ksn4KBAb0IHkKaVctP7kS7jI6EHu55pgSD5zcQmOJJitL283PL+pHQmGggXOdBJ
3p9YoNkevxJYQrYR2NzXIPSdMDOs7VOuNie689DKpuTdiUOT7JCHd/JtB1Af9+N2
0R1ADM1HB4xmmz101mvJvZqoZgA/yMb/RlRuVfM4ZTo8iSFxyjFI9zAZ2xI7tuqW
+DWoVxGGfS4JLZD1iWWGVS8yEwbuMZNnwJKBBglUlBHgg91kdSsNBkT76xvpLkNC
ERqC1MCAh7NtK/HG8gT7lK9ikMJnRDiE/zO1TGVX7rJSwuVIDnB7VLnOudR2M/bd
WIGS58oGmT7aOEv9QjnQc4MYam+ii6Ru5+4yqW3qC5XpiGEEi7o+Qi8IbwhnA+YP
blqlCW7+Gltwmq0sH9/fqFhvgjAWNyKUYZ2iI4CRpIv9MshO3bl3yHlyl8J9PpnW
Fr147qRd/pVeqBrhZZrnH37cL5IoYG7a1AuN4SeSU8eoX1gmWbYyoDc17PR6uq/h
nrczK4HRlh1d+1SL6ETdggkwXYMqS3WKS7vX2NhLHVjZi2mT8bRUjImp+gsfnTXn
mu17HOL7pT4KDM/mZvssjvKyGkgWSeBH1VjGpik41eb6vvZyeqEzFt2U+97Nf0u8
/48U2GfOjf3wRfUy3V50Uu7KKalvFUQmt20my93efHzJqtlt1IXMxy9Yc5SfMGIa
7RhqEBAMC4aIgEe7mY+PqCJD01g4w8TvdR3xTT6qYY/5njV6d5QWe0kNcNte4lVU
iOxQNxPI1z90jWZj2w6zN9fliklXMEqzhd3ZDU1vPGHwm97/RCu1HvULFK5B5zC/
gWmxrq+leH0S4eO9wH27IJy5u/vSMncx9FK8ZgbnNDOX9a2vkh6pEQ7QS1tn63Zf
V2+1ClIEtQaBrbQK2R4TcvVfRM8y2ESi4kTuQdviz/YdzwyPZPqIAGzXmEn6DlXh
NxKMA/j18QEeQnQiQexYJfWf4CEfUMjTbKDolPvFTeQ3cfwHaJr/dz2RoIw0wFcj
IFzs/w0UlX928gKZ+QXFz9TgEfqlUYErwclBJvxw/97b60ckwhXqY7p9JPQdR+Tk
iuFGutnMHZAGfUYt9F4XnSmsZU6H7VSOWOs7KjBoykGMwikR4MW0neFsbYGD+S/i
eR3I7BwNmh1sLzuKJMVu1QIlPBT6JaFoDjyZSb447bf3g8pmJ57CVrPpPR5RAHNa
4oojUEPWzwgfDGUbUFyw2YsdtWjlsMTjB1UFCBLrwEKa6LeA40UdVzjGvKaWeI/H
XZMiH9fOH3BOx3pYv7TpRG5llUgGXfdqPqMWIPgLHmlkqNI7oP2n50bvlg3UnYXF
DVmD0tijEeZSSdBVaZS7tqTaDBBBN3p693QzP6IYrWNP017IxGXnSPp4EMJ7FDry
HV9V2SR+YN5PCUWmoa6TdSNRbvAtAhjhdhcYZ1zpUqjEWSAVCN321WNIio747PF9
j8/fYo7g5uDk0WtIfORTcRb8pXSA+glGpOrEky5UuA9yDkfltXRZywX2swjiWGkZ
bzJ3eVEMas2GUNnk750N8Ise8Q9bKXLuzHqkNbwhtpZvy9Scp/vY++KyknSedHOi
lF0qngRxn3h2oAeVaQEM3PrmGOgjWiB6upw1s9ZEkr0eciflGYAqRjRG7TlytZ3t
ZlAJ6K9Cfzy88MSIZtL5wHm7Q74Ipy+6bd8M1I9rV3Fd/7WOqj8C+5mbM4G5BncT
ZpL59LPEuPWd/UPb2zuzn0SjWNMQaQ7zJzlpJsTznIHDxFPqsVVOCux+Gjnje+ml
uKk6HvsWAIJooFebctkYYlEOWqH87OazjpFgwL9RvPGk7nTU5RdvjYRMICncWKIC
DmodEFj0WQ0DaOT3fvBvhbXOZKMQDVHG/hCq5VAYV269AQdmcb78jajqqxi6hBzJ
iqFAR22otKqrp56W4aKiiPDlRAleLdNAkgdyc8Q+9ukTtOH0mC1cPx2/zGLi05pw
B5IZ7TpCqCAM9/9CRJb145O+gA0jZ2CvZ9jwJlS5mWCWInITh76M4DNzUhulyroc
rv7b2lVj7XIkr+ZDtAItJOCnv5kIHhhb14SyxyY789xPASQEyCFZHjIxbT9y991M
NLkm1+G/arGzQ4O5gCZTgjXCp3Muiv2Qczltn1NGcOZgJoCZdXvoGh+xNKmZanCA
Mhqb1rLXoZnh5mUQYJ32rlNbEm5jm4s3PTKBf1YKe16HRk//KlSG90sPzkZ6SUEm
KdppiwB0sC0BL0aAPcMbZxk/OUvLEc9Ye+cNdTM8AT9m/+hBxBuqaZHoXPIvIZfd
A3CyhNnEhdyliTe5ItWLY12cXqIOYDh5nWe2/y4UoLQPrusKSIr8lwt/uFCP94Z0
4bz5eCb0GM/00ed3cUWx1FG2BbgIos1e4IWSgIxrYuBHS/Dr/QxFa0QRFrtIs9jD
Ep8br6a2k1RU6IBvE4sjjAFZXm1l9MZOisQTgKeRjjkC8sbqvj8DfxLjQh7zQl0T
XiwpGy6Sj23EnSrDHfX3tBsfO9Ynrs8kx1hRGDzpHCjjVJ7FZEpBd5I0xnNDbjuN
xJXxKZJZWD+JmqWq1858SZo2IPTNYvMRgBNA1SjohkDchi3qCllgR9Cs5opY2PLv
cbqg9c1ST2AwZ/B1vJqfZ9Tc0KYAhfwONJf3SuOpmAwodB9zpx6o0afUOxcdFcs9
S3XfZ/wmnQQfOu6s9kGRZfYhR8czW0oXfZplAB8HubZih2l3kSQuU86V25jG43rV
q2zLqSUuL/anFoye5v8geHO01gGNmcVgRw/2MPLdHPUDLOM4csEKApit1HKA6Skg
BF1OWoexl8a9057JhqrMk2fcwsVHy5+O53FrSLp85iVuuGQH6uzZ+lqMHuTHpCMd
xDQs6r1arqpGWqW3XkIANocoJNplQaTgebvLoetizFOUf5Byb3ckJhCxWxXM7+F4
Nm0QvCQ0ytxTZiZgH1lPXaZMPnDC0d0CWM7EfFr56gHukCG8e9ljLytG2m4RVfPH
ZP+Kb3sbpw6w+eljCcyBckjiQqiE5ni2P2NfVg7FPpvnMTvOvM+0OpBomhH1f0Wn
DH4OICjtxCESK96pTjki+XgXpeTpSytIhLCRfUPxU2q41kGlx8frdSKTXURTI8yx
MmhweDzV8LIxCytXKvaOvba+iXE0LpXGJTYff7VckrpCjxYikmwRSIVqfee6IJyx
yVQwCMrLX4fRp/ZdU7OTj7GE4JHem0ZDgYeCrD/ooWE+AON0Ov/QrFLAkNLOUCnt
JpOZI1huii31fhKNwVOeYM9PK7Gi6AiuJ+5GP8QYcO3pSd5OpPUFaEPhVBzKLUBY
X3Loxy8zrFlFS7URIRlrT77BQ4522cpuc38P+Dv2Q/9ClSiAVJ0efxS77IpNW/cJ
osY7EPGAZBvcUMx/hQCwDgwwC5DkGh4FdQjpApMuRSUmw/j1fw4tijB/Fl1t2SUC
cfZIvqvGCJYdce3HguVoLViRddttiXCmBGeNd25e4TtwWaGzZyb71sQSpC0u7Sog
MXbAHfyR/tUd7AF5d/R5w80JZ6h9dW9HwqEKeBDMsRIS1HsAY2NCNt9pQkxwxCPS
H4cy7uzCnVg0NXTjN+uI9/s5zvHTC01TobvVyQsEhc6MM8OANmPbRGNjiObWU4aA
wOowlQYjPIvnwXWNlWVmsg5YJMeqeY6zpas5uSK9u9dLqtNDrWaTA+owK8dIyhv2
BmnHUKb8Bh6cO41CJcrR33xklhhajjjA9g2FBmPPne5dS7T7NWBQeqHa7OjzQ5X6
FJMpcPmcQMjEffh9zhgDWgihqMLCSCMu3BMBqR8u/eq5bKBLBwugGryiKvUMJ3RD
OMqRwWOlkIH6boVNpihCzDXXOmYPiU//p9g1QBLBu8kI+Om7FXLyNA0bvulfsCsX
5Oe6JziO9IP0ihSUGB5oUYm8xmk4eOzP7iC+x0eGETx8p5z5DvxgsbxPJQOeu2Jy
/zuQ4TI75bm21N2GM4ClxItpSr1WPlEN11S4leOO6/0nFx9DhrOHtJNcrg2WlsQO
PxzS15KJ4NpjTuKyFWBK115J8QNXLDZkB+NYQ2F9nuNPghVLiMaODYa2crwsmjwZ
l9JcTi22aCDzjqy9jKA9nNNR5YFxm+b0I0WAPyXyEypx9sV8XT2HAahylkNSAMgI
9UqQuFGT/2sNDt0rme5eIn0xMsqKLPWbRXCRb2GV+gka8yHH6bZcwp7cA6YRpcVm
Vmg/7auQO9dP9OuTP0K+CQhuV6LfSjpU82KKhsA5CYas+vPXyeMzt2xEp3+B/DFM
PnMK82ZKFjSF9S1rtSibOXNz+JmQQsxTrkEjMuZe3n+jfgSvqabJa3uws5WOtiXz
HT1AOP1HKwBOSocnoWdEi5BTIxaJNqGFkIZp5Ue5EyvgFkY5NJrk8uceeJw7TsCK
6vpP1WByqpJ1OxDELcJDP+F/bpAtcXliTH2UzFJCEHmCP3rtY3LcVJWmGPoFCyl+
rSG6k2SGx3eFXw1Mkt0TqQDxjXEwJbNK56hcvosdKHulsrMBciJQQOMACGRTi9mW
9PmBrURAwuvk7jWJM5qjG+hU4JZfsg/GGzBYjew2vnsBrtBiR80Ub6TleUWW13i0
3W/NKLBRw5UOeycmjT9Xjz1taDwFSAzqdhccP9cFGp7J6d3h70kilLNZ5EtNTaAc
cVV3053FX1hW192CZP3U/hWM0Yb2bF4PM3Boao4GpJMDpAeArZu7HU7pnT5n2MTK
C3fztS89oNl2eYP7ni2u0h/CYSiM7gWy2nHjHBXJhqLxjIjyreCn2Ko6n2ZtpwXV
H5XBpnz7z6oubnt3/WBFw2AgJvXeZ846Rot6lC8Bc7MmsSuz7eaietFxDoxG2nC6
RR298c9/1PKWb/L0z782q+NAOAmLZfKDFWBqUvu6gv9969V5fuluxc+nP3DLAdcL
4hAU4ofF52v+cnA0pZhbsRr6v9bTsvzMUQJdqrLSGq6uOEuk/BkRrriJ3U+zPtj5
47R9M1o9QM7oF10p1C71HgfYprxXrqK3h4kZ3bo+Nd1VDgE8u2sycojcNHLFnF1T
+jMPptnMSyRHB0HyinqNllhkj60a0st3i4KwSQHooSYWvCbWK4kU6HURN4sf3uJQ
3crJnj4ab0wNYOWzBsSmXmtkRqo1wEei1ACT+kdYxmkDGQvC29yDa+cFTB+964Xv
QKmcB5yaTqX5uRfTrNxjK91GlIWJHVYyf8y9/mIegR4CRv5mGsKk94JB9WA0eZ8U
/Ov0qIxR7ZVSnw2PJS3B25e63jVB2Q9cJf78pMwa+0cyAi7EBi1lav/j356YOFUg
E6KaBBQOve7Y9p/Lwx+qjSxJXvRYrG8IbH2XKLEZ4E6WAK8AGYS8R8OnsONjMCPw
Yo1RDP9iSVWh6oPQ7rWYr4eeTa+tYdKR7UevTXGzyvsI0JoJm9TSqkqjkO81Vpap
eQCWVM9aOxJzUOoQRQcYUWm7n+kwRj669q6XxW0s65c//PBUPx6eCDcXoDlrSJ7G
7gPP7kSGaQlh6oBIr/DlxkJo41QcLYfcKYVp+vfj2i8tzhlR1Vb77DCrTJ3PeCN7
eXaVTgKGEjTQNviOaWeTByVT/0JtslKD7c5oBOeXgQCkfUa4znEz0lmhASQXjaZn
RRnPsll0aorkcE2ZDmTxauY7jeWKhpUYG8B3J/azNQ0og6gPrlW9KCwr+y8IgDdu
oeL6a1eKsUyoty3G4joYgjwuFDZlfwB2A4dHrLKHWmtez+mmu2AiAZOzrpp1YpAY
GBiGAoGzcDnBZBd7PZzNE78COgOUGy3dS2ByyDQYoNXbgmvOAxp4T7Phmcwsokgo
4KKvJibKI9nnt8uLljDpcAP309JMtQI4C39Ef8FsxVcQiEs93NhKj6elJavyolt/
PMzn/PaoLSOLVKbGwcE0bHlq8Xf6J8VvHJPrQzkjnwHGeXMJklKGvu4MlrqEO8mL
hftg9e+YhFhP8JeVOmYwB18caCAgsDqLetqyimB+PVnySW0JrABrmrLcRkF0/Wjw
oO9C+TbgZ6dNrYBLrZQPp/bGQw5OSZ6wwC3HbkGBMAFlOB0zWGVHlf4rDba+2GT/
A6DipR4PMEm/QfN862FyU6bq4NCJGR3cWASZT5+N4wIbH5oj1reVAyM/re06J51p
hl6BsiBLujF1KEu5YcpQFiHFoqbQ7gJW2VJ+V1dR0UXri5D1gSlxtzxeaRR74276
fVwgva/Pgjbfj5i5Pst+jnM2d1pfmN34mRDYugGUBiaytQziNcRGX200w+0QNOAS
CfdwUHgR1Ds5PsRgRVQkXNkoM8CNflW5rYfjYN1exTz3GOkJXXzRdLszVm4sb0ko
Y9R3ff+3OtDMWwlrZHjmS/ghwYCUUGr4h/ThjvxtnAoVZpUmba7m7Jq+H0lUu7xL
WQGist2pINAz1In18LoyE0RBc0yHjBap0MICmcz3MSGfDtQPTjLlF74dteu2i0Oa
jvHfQzd1t7ZHyhsWjkf6eh0L5E3AuP0wz60+SsuIISLhIePNlmgWTAoAtXGTWzt1
LQLvUyGBMoHwELvy3beBGClgJA577UTyyKQr4+denPdkkkM3FReMZgXIkcngXPrs
yYnZ1mDmm0sifNrHoptTh2jcTcpr0WS1FbUtOygqyDA5I7+np4mLjJPouTODPkXA
0CDMcuGbWXlvZzI0zT4ySEWscG6/95qmAPGl/aQEo/vYpaoJB2L5rF+vtHj+9dkF
t4rDpxBhWMYnOt1uaJFFnb+R5ohq7oQGCz7KZlGkVT/J7WKNtuPcdhLs1Bk2bY1Q
0Es5TW35s0MAPnfpw1DMEyDonzkKAtJk7Ws/JK68d1OTYft2OpzwYWjiOMqd8BtI
UtWIeFd1xLODqnVgPlJQEhkX412Ix4KIbTth3pc09uS1iy28RUBtCZYN9q/RbqQ2
WUeBZtjaDc/DJOnrPxStEOo7/5LMWjfHoDvPcAO3mJVdxHkQ3uo3nvaqPEjg9L++
OwSDcFIhVvGJoFv5DZLSZS1ubI7cpWbH29B+ukh+fUPMqF8yKGofrTppqXHa3u6X
eSpi69sQag5zc2SbnhKlzB06d7LvVws2cp6VexN/mgVYuyhYyNtwGTpbBzTfL4E9
zX/qgtxd3SVGSgW6bvNVhBqkhOBjDRJg/dV374B32WjToyf6tE7qyE1w0pn3O/3Y
d99a+NgGdc2i5SKBxIhQkJrbbOfnba6P8pSXR/R1JSKI+3DxKZPPAjwRF2sAtpn6
YgNYHqBzhT873NCrtUny51JwIxNBMbzXU/MdcDjogNoYjLZhJ3EUPYzncSOjfVXj
a2WpdWQ5P5gpthv2kvcO11oDVnxeB1PEdzHky8FmkJrQSkB7HgDH+0RJneUu7h20
49Tx68AUed3nqfV9FeYn1NTI8pPFMC97I44VhMcctivzu9D1fVskuvdjxPcqfFuK
Th72E6h+z3QG26ac1Fv3KVXERCSqdkcfMZ/eALLQn3+QwBqmFUQJ+cP4Dvz/njhd
TZCU4bn5NzIdckK/mkBVo8VEuvYkqebTaRZO+Yfo1zAwByYPG2hgBZh+onqe0GHY
2t+SPW/gWQGU+RB5GxVHkVXxACn0PVbOI8EVaHXYxN+PAWqgfNeirJIwA1aSbNSh
A64NwZpK+gkCoHwvYLG1fF6tQMMShMYnjYKa4JpEy30veZToZrRi+yVHgw4zgjh2
khp0fScoXHq+xrxz/z8WujQuWNI6CEnV1OT5tTrhyCkSjd8PYK9fADSF0EBK781J
UuqDKSbWLMJcMsV6S0eM+qIrW1yfEC2y6RJBkW/k9VLxyMik1NLyIvDdjZdXgQGo
UCFzXpZ5TsPfeCuVJ8RSrq9oIq/oH80jMYHOJkvKrMb8tYWc1i12+ftoZOYcWTQk
n2BPnDDYeGgYrUU2rB5Dc2w7sCEwjo9qOr0iTfvgQoIujR9i7e1ZuGnL2bRmdd8d
4k980yoiFtOlj8EhXOweiXmV1GXyZQL+n3jcbwFdEpFeKkkB6jVy1ZahIXVTnLPJ
KfWfYtoSUKxBo7SzOOjZW0/bSEUg5DtUAf+gziSQSnBE5WWWJrVdoiGTWB3/ZZzj
8vbir5mGfdGYoZmPvEJW551c6qx+HvP1xs291Kx+rtC+msxvLAaNS4DbCCV3RFku
1CiN+VX1Ma+FHnFL2LDGCO+UBmu6kQMj+4KZYD7oLdW4zY4vyYKDo/dy24fr1itR
vICwipqcOL0Fc8dfZL2GIMvC2e4VswIYaV+cNTl3Lou9G1Q3uE69jolKFBUnZcvV
c/UstVFC4YYltwDodHksQHsGvf/aHoLMOD8H/sh1EFJk8BmDKyPpBhVB1/OqfjtC
R7lEAaUETFNj4Smooe6q4NDrravR+Om0qtd1jxjzLVMjX1oneigF25mT882UDVjB
dz9htNR5tu2hWr8Dm/i5nCYIoYqxKVgH95WHCBA7xJZF0v7AB1Kc7C/jN4HsnWvn
E0ZV7cTRWPnIeFGlg6IZnJE1il2lFNd/ANrBXxatRxud4DPZTYPY5jA7jcMHhbi3
Nu49sttzoHsPBqPuuz43aJItqyMny/vSQQsWmJKvij5Yop+VrTHFW9d1c9T6Wunk
27QbdTBC8Fxd8HZXuN2gRWVevuAeUdFiWR73dA/M+QZic7Jtwk5HuT/96pSUVCtI
xVOarYTiptKdcC/CObmhVVULNFzHHoBJVDc+6X3Ka6IrLAHVCndrsnk8qaz4yzN6
dLS5BKrmSf7vEKOr8q1YCf6me+so7gECebRhWYlJN60RIpblEP7jjspOG0drjm6O
Tl5ihJ8u0hPwBqdiQLnHtdL70AvB8zgvgCrgRG9nnvGm50mQmGA99JGnOoCfo7Uj
Nz5TquUnW7foyz1xXRai8k4m40vPsr3mLTAb+scKvOj0sXOyP3xXrv0VG+EWFCMS
hT5lupK1ECQFFkjHKhxlbsV8w8hFsWWIENaqUgzudA02WQ7ud+UjOgQ+ho0TZF0U
k9ONBcAqoIVtEfK2c/L4fYqj5dW6fqZfmQdML3Lrvh+Ht8pX54uVnyoEYDIOfPmD
4+XxEu8Jj6Yr+JPaELY/DP/zvWFHyp/VMUogctE5IGcvn660IRkeJnUrgGA/rEGq
BaBKIZYcYyvMxy9TILGZqmienCwzdhDlx9plxtC9bs42loTIP3asfwlvZY+NnyiB
NPK8dh5JcOZTODfKHKVbWewX2LIsz8mkosj9JPtToAYQORD3FUZ6aGYBUQi5gyVf
qBG5kd9gj5/1nlnF2DjsuyuwJ4WElMTN5FNb5anLvNz9qufjNf4anPpOhj3pczgp
Gao+eW7rXuMxT17Wa+BvbyCWgaUITyuxkOpOoxMPOTj81uLwkBmG/8r2H/z2/AGy
tP2yZSBCdwTt6e9SkgJJuw9Pi9IO7CBrV/zHNIsaadq7c1TBqh6LjOPgFgFLcMdE
OAZwDe1MHMJb2EtTVZzoSANvK0Lz5scSCaWAvgj8RuZhUFwZdKk144FHm52hpsSz
4Yh5ND3u+20wPl/i4SWewvGOZbMSXmRrxd/ypYr0qSgjlEnZy0nafgIaUt5rXQnR
xMC1NtmH4EqS3pPVDU+KeLqlAbRZxtBvQI7GyHBxB67YZiBgvgtow9ngZdlKIjxO
lRyqmyjGDdbMNf0BElq1Z07hu9ffiePPycTqfAiBjvKI4O20M4jgrhMf9g5VUrtN
jMT8VpU3if4aaWg6QMeIq1BYZB9cZunGyHlOHQFtrYyyMFArZsm2qylEpS4lPlXH
FmBW2lSGSlzwC7o6sk5h6gP8U5dOKTxORahHzY/U2VdnyLjy6zXzCumbYfoAvp1W
y/I81s2y3bNf1Mu5X/54MVkp679PDbm+12Q+0EbAhMjMhcv17Qvbn1uTSmbgQoVe
EDOjeOA25u4hcn2/LzvbuVPtXNltjuUz19TkXVjJXzRLQ3Vml4Q0hcFmsr02pURo
nxzQ8NEjehJrZic8clIw4OEBR/YwPG9CW9ZcMi+53Fy7LuvZIAzP5SeJCatxrHtt
VjL7F5SYkMbIww0/A4IAFzNKAeXP0+HDGr6vXRGQy0g0vYKxxaQ/j5vVimmvDeUb
x0b9fwGMaaDeEGZ/Me7+Nz8OXMpVLcSlxoyt6/Ev5bCoRrUju53EebQB23RqJfRo
xUrq7S5T0bPya6nIb3ktpI07ZWnymt5JmMEKci03UZCkIrBaKdjDOSF9aiXdWk9m
RQZn99djtZTuwncpNKQRgrva/JFZ7SRI+DDaAzkZQgWWYB+TBhBtUZ916xEBwmCN
N1pXNwCrbrM9npFUf6qBow+62j2RfAxGHllkHFXkJ7sj/XNQAGn31uVy2b5m8k2E
Q0qwsQ2B7fTC/4cSr0vINpIMEoXtw54jGpURGg3eHf4TJYfC660UeuiJmFuteXAv
+l49Oc+4NtHX8snl6qMoc5beM6zd8tj55iXruE9OLX1N2wQokFuLfL5db0cNgY4C
bEaYuvpyD39c0aMljACmgSKmcrKiyCu7hkiJmsLngVbiJgUZISidaDTr9RDLztNf
Nr1kfsmdhyQRGHbpCT+wmpz782c3jK3oJcVeSmCuvEBtBStOtKNE7On9p2yfSOBN
+6xtK4F9pzPeDVZ9MWN9t3xikSiHLE6IXh4b4Tsf29/haoknsJOAjlE3AJrR85xg
5UO/MXZU+zeYVSVpwWheXCmHEMutSJtTyv9YlvV94m8cNrnedi87xsv66zjGT7tr
/HuV/8l9MpXgngN7n7BviDKj1bj3R6KIJcHT+e16vHmYYQVTLwD+dPS47+hFNwmK
pRfOcemqP2qqp7IxD0MpgziHvZfVGIM07IQNqgLtqJnc7H+byMAFewUbR5c0Fu91
eYGhca85E6+VKCeZY5CufD/VArjQfWSsNwR9/yLO8j7cRgIRvdjlk1qPD5xFxRX/
0mqdaRzLXNLNPcAzquwoDTezza1ezLsGI/SyITqOkOP0tJsn4hh+dmXCPS9zkC88
Q45PPWPWMdD0JTcWAH7MKuApcyHTk69Her5npVRWWGidm2yF3dsvHr0EVvzfLyyy
6W4FKdr8ic2yZw6546n5cK46zjF8cUa3UIQxc+XIJ+4Sl9Us/eEaBx5jw9ZTGsjq
cV95f4E4674ijKBM0+GCh/VyDTLc78Q4+1JOi+/tXth1PJ30Bjrva5nL3n202xG6
D7e+NOTlXkTO0j6nXNKN2Ar4sf9erSxbTwbSiWAfkNzpNFlMeBPeJCOgqneqfh42
GoY/Iv8NIWi5bEMZLKAa0vrJQd5fxwci1hGvgu9jJ8ZaRUExV5LwfHTI0h2KSNeQ
ZcoHXCmt9bxZWxt2iEIur/rv2luXzb2CTBmRb766Fr4XmGcdPE6qZn394g2xgW7l
DfAboVyq+atwf2sP32LyE0W2i4J+BjqBoeOgUg07P1MeA3dNTXuN99T5f4RGyXTC
/oygeEpVEh5SG1wslaf37i0AaIq/AYuXmptcu2+fWVzsMBflE1Kkh5OA4fYu/Fc4
GZAZm+RJDZpnAqVbLBfaHgk712EjAY7cvnMBWqUJ7XKgsLVRmNjvQv1C+xOAro77
4Tm9RIR2hZcJ53H7xJ/fnVpf8b0W1S3iDh92znKDAVx652ELbvFSAk0lbZrNsarf
gXg4L8E9TkcrYnDBkZD7HcFiKnFDuv8CJMqYXCFH8yzWNG8M7E1R4Af14gM3FqEL
4yA+taSV9hHgdz5LPI+MZmuigj/8D8L+/wkgIHQ8E5mrd61bUZBlVlQ+vFfDDT3B
`pragma protect end_protected
