��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbYIҚtؙR4U�y���u	�����pQ��8(�p��5*�4Y ����r�S>0��Õ�!��(�au��#'�7�A@=̓S/��NN�5o�1�*���P��ɬ�7����qv��d��. �i�o�x�����w���-�_��~7V���y��(�&e����՗t��O�G���J���%3Aj�̭m��Oa�J��*���}g['nE��t7|U��@=XZ��|�STK��f�+뷎4:=Aop��
��s��V��U
��n*��Xh��\Kb��	����q��T2�H�<�\�5�ǘ���x6�y�����%�n�ӝ+�;Gi�UX�TH1#�0��2��@��ԑ��t��T*WG����v��K����u	�ai���O�S��3��a���{��a�*.y�oа�RF���'ff�"S�:�h�N��7��r�gC@�3=�q�jj�Ӯ%�g~��nw�%g���Xд���=�p�y��̡�~4���}�Ɔ�I
��0r�w{����t�e�$_��c
ޠR*�ɿj��2n{tW�gf�&)SU=L�&���'I��ٍ8��h�}bc�S�|��Z�u�E���/ǊU����`�
��WR ��F�b�"zXoO�����{����qW�K��\������&�
�C��.�� �J̫�J�
)u�[w�__�q���Ez��c���u˳��g×䔰E���acMJ����  O�� Lѻ��3ؘ5c^����v��ɻ���a7kŐ����T�w�"|ʁ*H]Ŭ0�|�����9�8�$MBH,bّ�\���3yP<���O�F`�.33:��5 ��<�����Ε~C����ҬEn�nLQQS�`)�,`4{�7ڠ�{�аֳۉ:E�7�����G�j�d����]�	p���)�fX27��e���S` ��o�0Q��e2�z�	ύ���ڠ��	��!lS3gG�2zyԳ&��%᢬�m�^V0+�w]�n��m49�HRVd8B)��b+<vI����"C��v��xz<�|��rG�?ڈ�U
p��R��S:yΎ�=�/�,�L���!� �ꮇe
m�fX}u��$�.L��<3�P{�`/h�̻�V�/�/ f
%;WNX�+��]虦��-�Z[�E`phq�Q�L�&�<u��Jۻ�s�)��Bz�9�y��,9�B� K�����\��ߜ����	E͞�Y��aU	P�u��F?_n)QhN�U�lB�)�iچ4`�L�`{��o�"3+.�Ȣ��#������x�NF���`1�3� �d��`��7\�R�3��D9	�b��t����R����Q?�-��p�p��aA@�=I"�.N�aK����VԀ�R��.����(��Q�41�����D����gn1�����,�̡�.���q��2�ߞ5"L%|8"H��ܲ ��vi󬿰�]�ǋ�-�Dg wM�Ez
��e-k�>��|���M&��3�=���_����λN~W�21*��|�[������g��d�6X���Kj�^��Q�
ϗ��>M9��`�4y�8�S��|����d\k:���Gǣ?�� q���$�q� �f��Cs��T�m�U�Ұ~���rk���NƘ�h_��'j����;���)Dv:�ԛ &
�pDLx��?�8�꽏�p�t���NJ�_zbܨy<��u�D��=1��K�=!A���Ե�$�]������"��gF����4���k��L�Mm%6�ð�(��#	���:qQ��8���B��C0	u��DƦؠJ�l�x��T��í��ߌ�.���y�k( �b�s4W���9�5��INd����B�,7��\,:8e�b(5yR�G��8!tk9g)���0_�ئ<ܻ�G��;��`�OYM�$�r��v*}I]�v1o�Wc���ޛ%I�v�wW��3ū��B�m�C|r�D������U�s��L�9�%l}��B��M��z����t�+��V���g�M��y���~����\b���K���Kݻ�>4P���h�<*e�,|����έ��������&4��o���e�H���o��|-��j9di�H�W���8u�ϣ��g'��ʏ� KX	�ON46+��}����x�<H�D���WR*\c�U��Jf��H��yt^�;=v���	y��G�4�/3Csc���	�����ci�)������u�* Ě\rٖ���o\�R�'�9����Y�"u!g�����Aĝ����;��졫0�I�{D3jc!)k��p�y�y�tB%�� ٹ���Ø|g�W-0/�Y�7����J*C�������ɶ�}�yզ���䳅�=���U =�tkO$-ܿ�Z��(�;�YX�)�]x���_��u.[�N>���6�B�$�w�l(�H�+����y$��M#�<tb}k!�CA�,$a@��(�?B�5�l��4�?�҉Ig�(���?���>U�W��d)�N+�#�y�J���HJ�h$5��ެܚ�^N�O�d�5%�@KX��D͈�"�5��,�$O��	��`����gȊ*��cí/�<BA��1D��\/,
6_C��i�
�M
`R#_c�˪��p֮q�^M�+��:�W����@r���dүJ>�?�����K2,p���tc��8i7���~̱@�����ˇ�w�AM<9Z;&�H�?�ru.E��ܙ$���1�Ϊ�+;�fu��1_ +!�x�J[�۶��ka��;�.}x��9;2D:ZԁH�RV$%��&T������{���$�I��f�)�}�=m	e���9lA��&~;S0[q���ЏGQt�����w�b��U���a��m�mێ4r���zw�b�!�� | �cŰ��1|��s���)9��I��|���5���wv��EJ�3�5Z���'����A
�G|�x��P�����l��we�],�8<<��;V��W���*"q�s�s�nCmv#Cdw��$�K�C~A�zW�{7�]�y�"#�F�Ux`{�Wp&��Ŀ��w[}\n���!R�+oH]�S���Az�r��]�)\w㏿*�����}�������בc����m4(��*o�Zв�E�j��^ �1�!�:����3����M�((��|2�:�!�>=�` ��t��7��IЌ�&k�3ĉ��4k3�Կ�����5��(�t�a�$�H�_�{SLl����|W�J�Ut�������A&[�[KZq44``��Ϧ=�?o�<���Ҧ	��9��cZ巈�K��������A��]�<����V3x��ǲ{��jh/��i�f�����➂�*��]�ft��bg��l�l��o�1�R>B��������r�'��m����4� 퍉z7MBr��E���E� z� )�I�d];�Pr^Ԭmu©7a��B�k�"����-������7�#����cN�����*�0G�i+�n�/ϩ0y���޿*o&>�%h�(��b��v݉&�X��M/e�I� ��jOd �B��	u3�+*���H
y
ʤ�u,�����]�	��H�l�h$+[8��(g�D�*m�_��Jز��<�靘N�|u�;�B7A�$��]�hOV\�!q��'�)�EKԲ��ea�������A�s��e&V*ʹ;��%F�BR{hvٖ�,���Z�k�b1��w$�8�_��+� ?��.Sߏ�1�k�S��Y��E�}?A�Q�)ִ�t���y������1�]V�_�x]�w����*��[k-*|bx�RӾ5Wx���1�����ju�u�DȠZk��؁�%�?6X���o��Rs�h(*��ںIóP������h-��\p���UDtAs��9.�g�C44!ܫ��1�w�Ě<��	�M�vF�+����e�P�A�xO1�]`��ul'�z���*�w��k���Q��ՒN)l�l⽕�������u�l�(��� [�hҕ��}���\y�H�S|e���_��N�FO/�-ǲt«��J��&3��+F ��R=M0\�(��I�>>u�|�Ǻ���@p��0�k0�(�n�jƒ��6M�y�b��།+�x02��W��ch�d\kT���6��>�T��������Oԡ骖����Q$��}�o.�Dr����{[���ыV����io��i�:��́kF�cS cb�6r�J�k���Ԉ�6��� ���m`~�擽�<���bb�PV�,"��%�7o"(C���5�F��'�0��C�5���#B6��z�:�dO�����<��9����D�E�rF�+IN�hYf(�+�:P15�L.�eI��Ai�D��iJ�'���K����Z��ߥh~�íۅ�}Z@�SN�֔��[]a[����N���.:Q'sl���o�1���TF�+`��'Dvr}�G����"�\����4b�1G�]ꭖre�h�N�!�I|�r$��x�:xej N��9��C�U����r�NA
�3⟋s\��I7��<��;u���f1���G�Q
�1����<t�7a����x��NM�6�g���du���,�)�֝���C�0��=�|�e�������[X��Y�����3ة���9��~�a�c��.�N�*��mB�QE��nc��  X�z�� ������0 �|)S�����U��z7�!_��Bky�D�����'���Y�t싈�uS6�0���ZA���Ϻu�&n�2=}�٪��%<�+���a�(��C!��Q0f��%[_J4�Ìp���~�a-�_}�3S���9���k��V�!AW�O@\O�^:�M���h��+B`1�q`r\ƶҕ���ZvE�]� 4�#\i����R��@�q�=B��@Y��q"I�� ��a%��k7�\7 ;x��9)�5@���?�����3V��N��@������G���e 0�'��C�S�� ��v��A�����b�A��V�Q���S���h��BZon��9!H��b�4V�X�^_\��&Ȑ�jDU�m"��N@�G�]�:�����>sک�="�ΐ������lF�j_�.;�ɦ�<ֱ��A�ys{�jX#���k�G���!A��
��f
�sN�z�i;h�k�[d�Q>i�?j����XK@���uG� TD3��5��)�-O��ĲJOJ���gv�F��L�V��ô��<�H��P�Z��P�5���C5x�\�7�c&ԗ���&�ޡRP�����H �e��R'�Z��EQX���.:���[N�y�-��g�k<�N��#��.�7w�/8��Ӥ@F�f���j��ܭV[��������vM6�	�Z/01?��#Wr��^����L�
P����D]�-�.��%��Ư���j|:-6vR"�)�ޖ��c)R����7��t�#� ��2¸r&f����J;fd�*|��7{�w�RT�	�I� �TX/�n{ez��I��K,����U�zcg3��F����fm�1��iCz��gm~��OX$崕v��JA{a��O���U�`�p��y�^-._2}�pUL���a�9_���q���++W�gk�I,���X+��߭q�����9,ϲPѣ*:��åY�}��=z�!�h�K�$��q���S�Kl(�>����TN$�`�x�HE����V@�YT�^.<֊��)� ��'��/����>\�
a_sa�]к�o��C�l[}��1f�Fpmq�	Ȗ��u�/W���)���]zOS6,uN�R��'-������4�Z����[�D.-@Һ��("/v��|WK|���R��)n��CBk����ޱq����?�b����Ƥ��� %Z�a[iފ�_�F�Lg��h�z�W�'ɽ�PU�Zl3Đ��q�|�wJ ���J-�K�;���
���&u�k]k%��`&��)��X����5���J�"-���O@�*�8 ֨��W7���h����:k�
`Xh=�g)�A���T�[5�T�se�#����$'�[ht�)mW��g����Պ���r��b����f,p�΂�Bn��g�,�h��l`��Ku��_�[$�m���"��'w��N�9$n�b$�4�*)��iH���#�K:	����s�٬�?�r�R�R�1A�Θ�̫v�>%8��iV�ƛ4�D08c����{mbRE�V���{HG�,bU��ٮ�e݊u�������,4����Q��W�
̃�÷��X���*#-gE@n���G# E?ɇ�p2�;�@�Ah��pTW���XjLJ����$�ԍ��	�] �h'#��C����ZdIi͆-���V\�'��o�\�|�;���v]G��G\ɛ�,�M�Aƾ�{p��±ೋ^�����"����ޓ�9�!�o.�锞sH^7qp���O�j�c/�A%���X�S���l�M��+�����f�`k�ОsX"�����5��T��'��
����V�ZϦ<K>�Z�DqO�k�/ z%t+Dy�v>�w���m�U�W8�<�r�pB�v��s�S|:5ï�9����=�%p��Ր�B�e� !O6���ձ��\ $��@[�1PK� ����*v�u���ۏ�"}!G�oC!1p�����xB��<�����' �Nh� �8v.2��a�����bLD8�Y��f��	�{<"ă�xl Es��~e�b�w gO{`إ����[Z9��������&��W�Q��.E��y,p������j�i
��p߿7Y�ڙ�'�A
�-��]K�f���r���%eoOT6�df��V�R>�~���ڽ��E�!���v}��#3�or<��]�%ml:?={h�ݛ��:r1��N����Dr��q{��=<̌��x�X`X���s�n�beD�U��~���wWb�ހ*�1 ����������|:�} 1P�`�D-�~��C������n����ȡJ�|�x��� ������{�X�=�Yן�(ř��_t���4h������a�h�_��ï��/��w��|�`χ�����M.c��ϪkL�����UAc{ɗ�{4$v*��9-R� ���~�[�L)_�F�s��ɩ}EDX��v\���Rx��&G��{���i���K�n1�h3��[�Xґ�}�$C9A����D6�W�\��j�<�(�ƪ��)���@}�,�Y=�Js笺\a�ЩT������<ubp[�����"x
8�<Ӗ����U0��}P�5o1�^�MSc#�d%�c�?�-��}�=�a!�5~ꂶ����)�D5]�����JYؿgℶ����yq�~w�vz�I�-5���!�^`��F��:'�X�C{�!Y�\�� z�Y�,er�1�Ew�گ�:�~2��J�5<��N��_~�%h"�_D��7�~���hS�F�f�,NW�FR�c]Bv���Ha=�d��;�k��2N2�*e��H�L�zl���1?�H��G�,'�0�����Ύ̥��#g��"���y��S�J��@9�bɊ�`��m�ֲdZa	{�;�Yg��" h�v���^�9��|'�RVXu�|�=�	���N����B�5U���� F�x&0�pmU�y��I�>�����\�a�hә�A��9��x�R�(Zp�[�����`s*� ʆl�N}�L�F�C���$�fw�C��x}�p���#����Y�Z��l���e۰} '��!r�T���n�uS�S �sf<Gc���ؤ�8�܆M�E�\5���vX��w��g�:Au8��Ѝ�j��^j�ML�$�!�_@DQ�ARYOS�gIeUL5Ӑ�7� ���\2�+[���x� -z��R��3^Ŵ�'����{l�A�La�%p(����"z��g�]v���'n�����b�S�
���P�Uz���1�7��� �#M$׹�H�^�F���2�~P�2��[�P���)�'�l	�ȷ%R6����nEB�����N��$�F:\�B���z�N�B�HO��E�\�9̾Y�)�����ȉ*���6!ua�|q�/#����b$�E�c�U���|R� ٴ�5�`������>s�˲��:+[5�k�������㿨�PT~3}�ؐR���'#��>7�R����H����6v}
~&��!��y ;�d�aƪ����x�����2&U��+[b�� ���1{��Q4��%��-"1�g6�Y�z `#��Ol^�)6�Q�(ī���(E��A��S&���~�5:�e�kK?Ф=�7���9�T�+V�D�۔3�k�$ѥhQ	��$/����C�XAm��Gǳ{��9p� #�v��u�5���iG 
E&e�V$O��C\�O]S3r�!:,�	љ<i���;G2�N�.�݃�����ʆ�����5���q)��B
ĴH���k\��
��C$��s�c{s_�S{��KcM�A6����������Y�����u4L����������<�[Ld�H!v�J=�f��k ��I=n�#=��K�Gܻ��w�j��^en�(NB����߮)I��-�?L���Z��A]��c2��N3t�1��W�]�<��|�Z�-mU�,��4�e�WV$�hYU��崕"l�e�#��сs"9�/=��b=����zaXO���;��v�����C��`�S�nؓ��]Q��ԙ��{!/�7�D"f�����i������,��"��1���8� ��=����J��9<�T猃����8B�(޳*�]E��XD���I����f��Mˏ�CE��I����Y�e;]�qͅ���nG�'3<���K����� \��'��D��W�q����ӡ�1�Ṛf�P�0$���'�U&�]ˉX�����C��$��,��k]��o֌S'(����':�KA;�3���;��=�m�M�W���<�}�5�]��L��o�~�mnwn���[�s��o30F.��������\qY1Op)�L�s���J�/���]�I'N�&c$�ރ&a=��U����w6��4R����W�uh�E��P�dTt8�������g�J��!���F�kЭ�+�[$Q[���o�DD؈��`���.~}��Eo�Y��hJP�;����
��`Gj��%�S�v�4S�����*YB�ZB�R)�זJ<)��;�1��9�2�#4��<�{��)4Ǯ�� Iw�-����BK��CYtļP��b���\la�4�9�cZ�ŀ 8�l�T�o:�O�������3���X�5J'��4����鐀�fV*4�n��6��M87Y�0d�k:�zÙnff��X~��U�l9a�Ty���~yT�2��e�Z޻��zз%;}�r�G��F\]�*�<}S�G�YB,ߟ�؇�м�q�t���y��6���d[�p��>�K\��ȍ�������ʲ� V���Nۙߞ�'�-f��[1�(���VPzJ�q��y5�ׁn�J ��Ggt�Z�V@�8��\��He�p�r��k�g-��=R�v��=(T�(|�/J�iM��ڿML؄���2�D��_�D��vE��P|�]`�x��T86����-��+����l��%�i�b�~Q,�K�H��8�~�P��@#V��"��%���]�1�0��d?&$��lc�)-���9��!O�&U���;���@�t���7ֿ�7�;�W��5	6ǣ�	����?b�>�ly�Y������F�?���HΚj��6!Q�켑�f`�Vԫ-��[�9ߠ�IcIi�x�w��_����<R|&|*�(p2(]Kw'��өv��J�s+!�m�ޔ|��)�
D*àY$��7�bb(��ː:#�ʗ�dԖ�q�<`f5��m�I�ݲ:Z+SKsjN�o�e�J�C��� VtV�^�kQ�	���7~<r��3c�Fm����:���p:����14/!��.n����C&�ZOf�2��$�/���b��q�K0檥�����݂�e���qs�d��p(%��a�T�b섩�D=I��]�r� 桡�4{�Xbơ��yuV�;?ח�U��If�6Ң�l-t���(��+������oY�s �J�eL���4	NMl �H��z��S���5+�?p��A�Ғ<kd�7���2��O7F�o�o�A��v��������Y�S�%�R&�q���s�g6I?-o�w������k5B@l�{�"���!��em�Ah�H�_�l.��EN� �P�����͂9L�r��XI�I�Cg����#����j� x�[�[��o$%���:��2��]��"$�p�)��J��\"�e1�B:!�4��z�^g[ݑ'R9��8RX�dYQEi���h�����a��7D����F�w�t	>E�T��m[����ˌ��Gr 3V�
8潘*}���5��B���J���Ѧ������J�XF���fz[Uҥ�`���W�A_�ISފ\ƥxMx�@5!��[�+J�h�~D��t�0kQ�u{�)�{Y@�&z{���U}��`.��w>��zRd4$7�1۱���p��V�i���n�CSVtU�3FYaD�
*O���at��-`;�32V��b�<,�w�z2"���s-��K)�6�4�$�'ĭ�dJ+��ώaz4�d�a�hݣ�pZ��N*�48�N|�B�i���>�P޺�/��_�h����-6�͡D�}��g�XG����E$���J�(���#�(I�}3="��#m�m�bf�u����ָ�����[@g���P��%o�@�F�:�3n�4+�-��$�m���aZ��y�XC�ـ/5Q�\Z����5�'�%]�C����%�Mg:����)���W�ijyR]N���q83:����ki�2��2g��*�KS��0���Ŋ��^v6P8D��޺_ֱX�m�v���/��}Q����t|�S�Q�?��|U����F��AZI���y}B#zXw��X���׿lE�E�Ӡg�� �y-	�S��̉���nR�.�j�*����q�DO����Ib�LZ�I���&dW��}���ۮ}�����(�|�n�C��b��C�xrD��U{�)[BD����}j��1�j5��D���l�LKz��y8����`��Z��r���P�(w��@��S�w����ES�5:%��A� �جpK��7��9.��'��+�D�Yz���e�x{���Cb�%�'���Gw2�g��,��I
DY��=)�>�&�؍��OL�p\`}�kEb�_4����+-B��
������0ϛ���Lw�'��͡�I��|��D�@��1j�Ή�X�Fm�����Eu-�7�ד;�T]�7A��C�3����'w\��;^�BH2���ߊ1ȗ�p�?���eb�u�~@-��&����N�7րh�K�bJbMYkQ�/��A�|��(!~��~��']5����C���U�x!/����3��e���1o(�V.Od��WƟ��热
,�� Aa�|���4�!����T��.ˬ�5&�w��%ͦ���� n!+��Lh�I_��d�^��x�V��ʓ�A}C��7�J�GHlgD�.j˧�D"=��O�'��&�������יA�=g��q�0�y��Gӹ�|�|��J���|�jb�6�NR,8]'f���v�"���������jΐ��GK��I[�b��)���4F*�wql����oq��tU�#�$�
�x�R:�k���:��#rtc�w_H�(� ���G�H�ծҐS�d��I#�~�r� ����Kj=Ȉh�[��<����f�;Q#UJ4�7�B90�*+u5i.&&�h�\u�#*'�OX��*d�Zr3c�N-�^�Fд���Ė�4���C���l(I�B�5�pd�B�E�O֡~�s׭�� K�`E���P�ù�)L[����>���Ϥ�55'���� �&�yS-�v�4���*|rZ�ж(wi}LN m>����i���M�	�Y�������Zͻb�eu9� o�߁�W�7h)��K6�)d��;2���Z1��~?�:�7{�X����	�H��fi�B�8��W�ϵ���h1��;-��c5�9�Ȕ�P�D�{4^g�+���L5��s�ŵ���#��!�m��qIAr7�d��"��Y]���*�*�2�o$f]�y�٥Oa�ֈL6+e�Y��hhU�����Ȓ�����&\������J�K�pN�Z�jR#�i��	��姚M%���,4;М��/x��b������K-�L�cj��q7�%�["T���G�4#ɶ@�6�dH������q��/u���;f؝�U29��´�ɝe���t[��?m�Nf�Y#i1��!�]Q���vS}�����ß��Jr���4��h�J@͜{M�`k�O��^�*F29g|�?���5Yw*�@EZ¯�ҪHie�!]���g@�\�*q�ʜ�)Y��R�� %R�[��JWg�f_�i�ͽ�L��O�B�\�q���5YӓU쥰 G�䡸�nL����|n�	}\i����.(�Z`��"���8�4X)H^!��x�i�$�?C�����.��|j��w��Fhݼ�1�O�K��Ȏ�V�"gw���b�'�&N@�}��M��е�:�t�Fj�/z[X�t���I��^���F�[8��<�i������֩-�k�=-��! H�;��̒a	P�ǳ��������,����ƙ�����Tv-�\di��؍>�%��M��d�͋��7��I�z��6U��%�?}�YNq�I�����V������Al�ʱ���6M���$�﷤�Fװ:��g�t�.��y+��p�:k�B|�@����`�es~�FӞ�]¡��T�Tt��l�	2Vb$ncnf�B�[��/F|h��{,�����%	�Y\�<[�u�h�]N܁����+��>�1�-I�����$���.0�ThFN6e��쎞7��F@��К{�Ƚ��@4����@&R߹.�HyD1 �X�)Y��G.��˽�	N�AQ�\+��W��	�.�?�F�U�Se�#@`�\����k-�<�Tw��F����<�X�:�Ɔ���}&_+���%�Z��c�5	$�%�e|3g)���k)|m��UqC�T6�\�D�����^�[�>*�]˻0^�A�\$[�e�/�Y{����t��"?�flZ��d�d� �	x��Q�*{�4�Dq�0F0���5�_|u��f���>��]�F��HqS|��
�4}�v�ƾ�V���D]l5%s�v��zI�+����BH�f��$�"/��Ok}q��dB�]���QtM�3Y?U*h˖��,��}�
����fFp��5ڊ�Jx���\oӘ(e��$=s	��n}��+�G	�8�~�u
V5U���� B���R�mH�}�AR3��1��kmxVY_�o�z!'|}���#�4O]�YP����h�E�;;+�"�>	j��������hm	L�^�D�;^��F�
x��T�	�+�吞;��r��uB-��9�]=c�^v�Yٲ�<*�C��A�`��ծ�&j�j�2ef��)�Q����1�I$�%9����Z�w�?�-����q�N�;�t�5ꢽg!�:�`:�����R�#�`2�M�lX!�ݏ�_��یlR2l�s����=Q����P0�l븒"�r{�˙�����jY�J!�b7r���b������H�+U�65��|\���|n��K�$�ē��Xу{���	��9#޽�����"��@��z�	5�B~y|��par�꺒HA�9K%�x����ݓ�_~P/ew�DЏ��C�w.1��=Y��i�Ns���Kݛ*]{��&���sb��Cnj>���f��e&g�o^��-��Wr��w�������y��q_��6�6Qс��#�>���,�~�	�I��g_Y�+:6�Jp�O�cxh��ԗ'�EI��(�H�5
*�QC�DH��8Z%<�__c�ϳ&;�h͸���!aA�P�Ɔ����n���k�7g܈ �=���,�7��1)�h��xi�ݮ,��M�,*����4��"�pTo^��`�D�l�=,y���3�x�tE���9����Q�Y����T`EH8�?��	�Px�)�/���ـ�f���օ�e]��=��Z���uFLo`�<�J�l�b�c"9}���;��S���Ng<�����S�I���IT']��a���j��Zl�t���߼ڏ�2n����
����_`�j���Y�c1��G��)Ԝ��.������Yѻ���A��?@O�nQ���/P�F>%�"��+~ܛ ��Wn�����3Sw�Mu-���a{#�~ޭ���&�6;��>a/.���j���GL��V��]�#R[g��խ�7X�{\�̬�ߔ)���Y��UHϓ�4�w�>HN
�;�C�����D@�!�V`��?�l�DX�j��x��s[��qQ�p�
Z ����^���Q�q>��fO���<k�f�����%uVU�޻������9!��R}n��ڷ&�]��?)7�ځ��|O'��W�wM�@�ec�L*�]��;b�ˤr�aᵰ<+8t�Vu��.�w1��Ҧ������KApq��c��,D,�%]�a<w(�������Z�1&�PxZ�����	�B%��|��q-���P712���((Nk��i�I���2ƛi��R"ax��y¾�HX��&C-V7��Jν�Jn�I-�cGU��]"�3�<���K�`�{8iV��_�wP9{��>�em�Hؔ�J43"޼�n�����E�:�M^���<�d��l5e�}���g�b���Z�������xl�u֚o⩇��G=Q��e�> {q��������C�
J�{��Cɶ�C��b��s��r*�G�M��mƶ:�RS���R�QB�� �������\�X�{*�|�Id}?P��<zm�&��$B%?}�@���?+�z�­��Ԩ���F#���S�_"���4��ݳ� ;.&.̴�������V=�,S�N�5���3r�ڄ7�ã�d�O���0�;�f�> un;:��o�j���@�Ju�K��Q(�<��Z��3nQ�KM�asV{�D��*@��R���5�o�9����LUl7=!���x�x� zQ|2���^#�
Pɲ/2��ƅL��8�a�G<����#�����p�揖FW��xg� D��-����ĭ�m���!DY9�5ْ��HBN6{hT��N'(b�k�NA-{ @#�/&�d��
m)�CwJ�� 9��f�gW�D�_Щ
1k�^d.,�ɢ�]��ԗ�p�!�K&)�
�m�in"�#���W�:A��\�͎*y�ٙh��>�HX��k��-�J����F�rY����"G�p�((���К��m���tK�`��� OyI�P>n��VHWu�c��
%o��)�hm��u�k4�>�Z����|�a�`��:��R`�LDt��e���D��D�^%��I-��"�)���SO>G�ɔ���\RU_.Y!�����|��R�Eg�jf/ka�8y�ue����E��}M̂?��8�2�B������^�J��E�H8�IU�$�������4@�������o���@|��Y�g�ħ|���@��`ӹ�]�;�/4|$eg䟵H=0?~ī�ұr;���/pղ
�#%�:�Y�
�F��Ruƍ� =x˕'�:��Ǥ�S״T�r�+�݃:H�/H@�Z+���m6��,�Z��%�P���@��=�ʨ�����Nf/�Dut�Çc��:-����;J���Gt�T��K��<`�:}��jw���RR�#���f� ��f`Kr��Q���A��k�s�N;�l*D�3HO
x����H�عG��zb��<��m�
��d�M+k.���?C�Q�K
�Io�57��q�W��\�~BVˠs�*\��hs���g����;��*���Q�D���� uhɼ�Rk���M2%r�)��A�E!w�Y��>Ia�����<q��P�S�����%�$%�^����f;휞<!����i�4�Y�?ȳq���V�h4�!���AFQ��a�>gFL���vͅRh5�t����WFZ��U�u������:�u�&�>ߩ/S;�S#���KB���MU��Dɽ]�������}�aʉꝫ%����л3^:0���X�f�`~�v���N}����IA*����N�=�k�T}�B��G�O|~f4Q��D�(K�$ח�0H dE������K�O�J���G&��3�{EQ�#~�r�M�ۊfx��g�� x������"�ш�S��-=��`�y�B��1�0Q���A����[�P�2��̵V�〖"��/�-�Yx�Q�� �T�5��7�U�IT6Ņ�.���-����S%��0X=�*�X�j!�T<�"��П���5����$�Jn��pH��nY�v�D2�4e,�@�|J�Q7�޳�K��T��'1G�_�����4#0�.��J�Achj:���lG��H��Ylvo��wQ�u�zj!ԭ=�c��ȕo���Ժ����ߺj	��R<���њ�`g�x����?��f�(ݼA6}r
n� k��>�m��z�׾���&�~[y�W󯽃��j���H�o�E.⦈}�"��p�
����;�'���z��+esC>\O�F�����T�8��& d�a�/1�j��g,�C��W2�\�$&�{o�T�B&v��c=ߔԫ�]v��`t���Ϛ��_/�tX��ּs�^rS�ih�ӋP%e�n�*{��٫X�o�	��ig��1r	>Tç����0YTpA�J7*ԥ;���Q�L#��j��+"�-��%�*��[N<�`�@ �s���,�j����+_����M�yK����1\橬��^ g� B���]7�ĥQ��@{�m̎�ouB^��7zY��p���(63_�!���Mg\���\�ƉZ��olT4L8i�Y�8�ѼE�qBAk��
'v�����ax���ܣ���X��T4��1@*�襹�BEy5��QF)[ՙ3F���$� �X���/���8:_�o�8<��!�i��J�d���`}ȭ�w�δ�������`	'�����2����q�@��[L�˷�F�y J��Ğ�7Yd�d����g�1 Y����$��3T��T�{�����OG;Q;�@�;%_�C&������C��\׏��(�,V���.�l(�!3�ǿ��C�E���6h%,�4��g�T/��Kha� ^Cį u	�����*��9�����&p�:�<Ap�,�]5��MP�>8*��NQ�9V�>1�{:R�X��AXŢ��z��1`O�����r�y�rW飼Ǆ�-�.���'�.Tufa��d�HX��A/��V�����}�=a��2�,���moe[�����-1�7�	��Q ��N }@������r�k�zT�����B��/&R���ILX�Vf+ڦC�����ѝG�	Ŵ����;r�FV�m�F'丙�����0�g�������"�Es�����]�Yx�F �՝�����ܘ�2�G�V�W��H?5���N�b�v�~��2�1����h�� �6�YTo���Z�iB�8'u*&%�_��k�G�2�Y������0[���J|j�q�m�%3�Z�b�xO-���BG�����Z��@���{eΚ_�
�V����v(�v�}���'�LD����5C������Ҵ��PN#��~�B��BM^s�~��iU���"/}H����Ƈƺ�Y�_�re����	%eX���a~E{��,��bF|�̄��8���H���W'�f��� W� �O��SD��ަ�Oϫ�|�v�k��������"r!r��'��&���)��WyH�H�q���R缷�I=����57<$�"�����3�u{�?���}�޶���\���}��|��AP��<�DtV��>xm�0Yd�4Ү��=Cl�����uX��`P|�D�í���-���`�e�D��JS�&1nM"������y2}����C��:-J��<�U��l�79��U �?�5U|4��1����S9$UA�=��s?�wO6K�k/<��,ML3�o2=N�#�Ƕq9k�`r�����m
��P#:�����)������U^c�«�+����0e��d^Y�d*:���c{+I`q;�"�;1Fus���ӣ�)��U�gDX�5	�[��Q���0ڸ.���G�!`[�ƓxuD�e�<��)ʖdAW�}��%���/��"�n*��H�Q��}s,}a���y@ff�<Վt�+�h��֞��|.�����N?4.�m$��¥�b�h��܄y6&׺P�+����3=���ǾK�ֿ���Ef(�B�v��`XO��waJN�"���7?���v��q�!Xm�Uf��죑ۜ4�M�����������Z+y�6T�(�c��4�Q󔂾�Xʞ�cx����#qzٷj>��I���C�#N�5��q�̑�>>��X$����f��Hz��<�/���':��!������5}��]�� ��=w����k�%Z�F�efJ�W�qk��b������7�zL	��h�vr�%�~���+����G�z��q�W�R������F�d�����pJ�?hV��qG���,b�,=�]>���Vߘ}u����*L#���q����Gq|^��Vؽ�d�Bs�� ,,�J|+׌�c������ԉ���oF �ध&�V�����Ʀ��5t��"�֢����c�M���R�O���Nڃ��)��ii�����@�G�@�T,�����;*(����ED�S~Bk�>���]u�T�}s�����ɥoOu��/��G%�q(:�&��0���D�S���qc���o�_c#�I����:
��,��zQq�4u�x�QV�鵴G��
ݰ�(\�M�j9�G��slR��VD%�D.������m��2�s����i�Z���h���si�wK��Ej�0)88͈�(��kW��U�T���.ܬ �¨R,���z��M�����O�h����H��L,5�:��4<`,�K�;tJ�_ނ��u�QF휗��;��5y��F�-zcT ��	08�c�/�Z�J^��==lާ�L@�#2u��-��gB�m�X�N�^����