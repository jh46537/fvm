��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���Ⓞ,B�$t�{����c�,�-��� k�4�	��[%��B�?���4��\������y�0ֻ4M��'��&[�A�2��~P �i�)Ԧ�%'A�R�t�t �*�?��v���Pu��G�� m��C�I3�_DF��(l��EO���Y��*��=�S�-W�Q����Ge�E+�>�ěz\����>s9��!�M!���m���ne�&()3�N| /׾r�ƙ��Sr9�`b�	���J�O¡B�J��WaK���2�����(��_C���q#g�sr>�@cF�S�]�"���qpRC�u]9�Q6�)_-Kҿ�3��6q�沿�E�<�����b�����  f�@{;ʰgLZ��x;r���
 �P��\B��"2�yP�#�]0w���
�%
�fE����=i�|�c]T�@l����Ẁ�N�/�(��Ѱy �
B��ќ��è��ā�/���g9x�!C/��P�U4���qł/��0ߢ���.����<��s�:QD����e��,KB��C��W|"n��\ӣ��]
z}7��K�|�)�	F�&!���e*8���f��'�� �fD'9%�5wk:�/j��q�?�/�̩�e���	�u���X�=��B�W5t������i�^�`���.����%�v�@�*��> �^9�kI��f�M߄2.e1�u�e��8ҸY��xw���>N��*w}N_�x{��V���=��9�J���]!	����(�o2����YBl���� �������KT`�#To�Gv��]�f��5%������P
u\Uk�m�چs-��EO�w�H�����Z�V�,���}gnخ���" �%���3&V�
]��]r��zt�b_(z��j/X��>Ϩ7D��Q�P����j��`sS���0Sl�U����d׵R��P�C�:O�<v�IF�b���]�R���bO���s�W�����m�>70
o���;_ǝ�L֟�2z���W�}���";	���� m\՛Ïu#*�:\��X|1u&�7���㝐ק�P���-)g���0x!��6l�EB��.�	/�I詏���L�v�ڂ\�i��z�}*�.U~�fa.�jdHn��Ր�� "aa�W�	AՃ�Z��S��Z��9���V�����))�o,3A�HF�Վh�^(��D".#�G�����A�0��p�T���x�|u_����񚤇�\�](��ؖE���$��h�b��~���S����;�K4A���Ӣ��N�*� �ulFs�B�L�E�g-���uT��c��!���D�����L�ʾ���j+�RĤ[��j�8��5�=���>^�J�=�,�6&�!��Y����Mj��׀���з�͞e���[k���$x�V�C���<{�b���c=-)&M𕹇�����
^�n;�5���\�oR������L�X�6���)܅�P\�%]\��q����  Aq�IKp��;��N���^�c�֌go��q��D"$��������+;�X,Q�@�4��X<�i����Q��
Щ�X�x��p�\��O;��5"�DQ��*���~*(�w`��JF��(Λu�a�<L��o�3�*rb�$^\$F\]�+����l���ҥ������@W�9�R;�w���3IyP���k-@v!C���	i����W�:zӽD����;�F��3��٩�{�[��'����u������_#��K3W7�s�S���1�m���Sf��6��k�Gz����(�q��ŝ�u��:���Ώߵ�6Ba�V2-74���Q{�G�{�{X��꡶mYNrf�|�L	L�5�#���vUv�<����I�E�Sl��J��DlR��(;:Tz�1�|d�slK�?��͠��p��?/9�t-!�"�j ?���=�n�A��_���!'k��"a���׸/o^H֠ޮ�_��~��k��k��H��M&?���T������C4Inʒ)r��'��1��}y]\��f��Y��;�]���u�Z��o�{����G���Hē8К�W���z���-`J�Ui��f5��-���~0ەG']��.+��i��f�z1�HL���;��j�����ZJ:��JG�\��l�:יLǵ�h�4�k3�54ײ���V�dM@5������,}:���R~Sosҽ�����@���.���~���L	  :�Cx�����n^7��{�a5��f���d/,oo�����P���7��vH7��1%}�yiP��[��� O�f���A���-��nԍ#��ꏞ@��T(�"6>�����83��o㭝�gj�{z�9#v�q��EF���7"zȥ���c���{P��{tE�vQf���j���	����[z�%]���sX-��2��/ޤ>
7���-U�����<�¤l��������������|yp�4���#���Ɵ���!@(;��f�|��}����O�4v-}�����B���vc�����A,�"L�^��KW*�SP�A�4�X���0+�V�����LCe�ܸ\c($6ߋ�S�LQȝ���**�UP$��i�!��� M�~Ԣ��W��K2��U�T��=>��)�F[O���{���1���7�j����o��b���V�a�:"�f9v���]���zŊ*CMǜpgD��9)X�v�0�>�j�nu_r(l3?I8"�s
rD�2EJefJ��mf��[�7�qEN:���`0����m*M�9�'�.0��֯�Du����^1��_;e�C���J5=,m7�f�=��|��	����7��q�R'JH�t��"��Wd)U5�����+n��y�zJt��J��W�s=m��Vh��Kd��UIRᒯ���4�خ�eN>���D�l�c�ŵ��ĵ�0�=����f&�I�,Q>{ � W�(���r�oR=7�[C�>���H3�6����nt+��"�%].Ls'ܝ/��w���o�5v�Uϣ�e#Ǒ��Nq1�ҋĝ� A#�a��� �9^�u��$n>�p�l*?�!���s�mM@E�5��<(�����(��$*�v�2�a� Pk!P^!f�� %�)
��Bn����������'I�ߢ�?��)39y�W� Y*�������*�a����7R� ���)��SNAMRHH!T����K�$W��(ܔ�m}�8₮_�d\\۩u}�����cf�t��IhF������LY/%��^$�m�#Rpx5v5��!ບ�]�C^a��2�Lq͊�$�"g��"r��BLZ�٨�m���	勒��ĲV*�f��F����^�V@� y�L��vB�=��'1�;��"�)�Bų�o�'ys8L" �*z�	��}�P�O�dMCGmZx�&[�]Qh��K�'�ޤV����nrw��/
�UO�ng�'b*��iv-� ?A{���y�,�H�h�}o��f^v�ݳ7�s���ؖ$�5Oy^>��-<��RY���u#��N���Z��w5�4T3��������(t�hc"�w���D�^���q�����nl�0�9��]'A��<j|��sqä;��r�̮:���vk!|f���奥�q�-��ĕ���6�ex����sV�˲��Tً����g�J��1q:`��Q���>�v��NĶ�ʏ뜩�o�H1LߑMf�� ���E�Fx�F�+��q��gA���Vy}J-v6�=�K��S#<�L�̠>H��<�ν�l�{n=O/�r ��ǔ�}����H����/.ڣ�ΣH�Ս;{�<"?�r��ځlӺ�n�tW3�`Z>T߻r�n�%j�Q���}��w���pR���?_������7Ɵ���n�x
*:�4T�[�� �^[�dK�Pk�ɨJ��:�ȟ��[��&� 4��F�[�������7�����o@ }y��Ũp
T�J6���YL X�r�mgY�:H�":ZQLE�M��!mx yZndcv�~�Ц����S�$i�f*�U�z�����Bg?����yU268�O�^�+�S��d�%hG?2�U>����ݤ�US�iPu^9)����zpO\�Z��Ҡ@N�Z�O����~�٣���aL��Ȳʘ�N�Q�m�2>��q�F��֐�Q��˱�/⫡�g����ϰa���/����-Њ�A!��
����2B� G�� ;�O���/���!�IH�Dv
l|��T�2��U\�q�>`Q|�L�d� ��o}�j�(�� ��Y��@�`�S#�w�f!0�����L.�
Ja�\�%��Uf^-��Ƭ�U8fw��A]&{�Dt����w��,S�|�bbl�:���k᳆�ue#�h�~�id�m=�~�bt�����#Ɣ��O���EHPk��K��e6��t�3�_>�����4z�J�n�yK1`#�/�����
{8<���Af�;����=�9!����v�֍�r%�l$�+������F"�:�b�6E�ӃЌ&�C��T���jD�o�LK�;�IĽ�1��m�o�^7C���e��Q�g�{^�-���`X�,�/#I�U;/h�U����<�b�L���v�i2������0��1��������F*M�y��PC���Q� %v�>�ԡތӏe2rt2���a�_�u�'�'~{��gT�q{>2v�I�f�?v�e� )��m�(l���@��W��Y|W�����g <�\���{'Z�$ �W��N���끧7nƎnc�凎,���u�A��ܫ�E��(��	���2���Zy�hc(�hff���MP�5���T����l���>����H2���l�M��J�s`8w�"9�ۭA3�Q�L0����_
"9�s�R�%%W+b!O �����L_��~R�F V"�y�����H�{q���q�z�������yzs^r��%�_��;�;��KA��^ZC�o��d��թ |���Xa�d��,�P�E*oE͗׏�Pi`w�o�7���d��K?FC���U&F\׆����~�}�nLG�M\Y9Z����Y�8���G��D/-;X�I�a���˯ܱо�=��8B�5�� h�]�͆�+�tH�]���vfq�� �ƠIM5��Π;e̩\��������3��-�1�������6��r��a5Dw[�5����[��G�G�bw�ӌ&���p���U�������!��yZ���v�c�,(OS�4���N�Y�݅�r	N�����GTy�w�o�Ob�b�0�S�����v�?؞]fR��J>a�v �{��~�hvqy��G�F�<�d[�9$<��h�:���CX������h�_�m��;>��?	Ķ��?!�Y">ʍA������>�Xs�%��6����QN���YˠgH�	IE��} ����ר�\�I��	�V�)Q��̓)rm�d�.��g?/�!o ��U%�`E{�n��٬(��f27k9�@�=]�.-�T��B+���H}�/
���)ӥ��Vjg�ֺ���Tᆈn�BNC�ᭃFj?$��c�/����'+Vi.��:BGrD�^�Xs���n�d��PM����?�<G�-��"���x�mG:6u��5m�F� �Ӆ~���E�a��@��\�.o�%�=��VW�N�[6�\��h/e�Q�|zr��H�M|炽DMl��\���V��ˬ��IA�N�:;QN��T|J,Iջ0��h��	R,�e1y�'su�������hy.Ĥp��MF���Fհ���r�*+�����O�w/#�cX�'���'�A�B�_�%��7 ��`|�ώK�9𫝔���b��F� #�Zq��/�Ip�)��q��d0>W�61[������:Ӿ������y@��mҘ�[��f3�G���|�����Zk�v����V���;�ۣ�@�o�-�Th��^^b���Z|�1ţ���xx���3̶��a��4�dT�!��j)���v�c�Pt�
Ã>�.��[����"�~��D��/NA�י��Ic�ǒ��0`4&��kY�[���+�'�_�X(�ڈ���"�DeO�4�1*x߹��.��Q�q�ω��$��BT�vK�0C�+�6�lc'8]P0X����2yu����w�׊~�fˍZT���̾7�	�1d%���NNz����e���O{:X �F5���\��yLfeNq޳������E�&3L�X��d������J���d�CDt٫y;
m�:֟����}��?Am�&W�wcڬN_�	"�ޢ90֬���Xfy����]��*Hsr�{"�.��]�[�����W�n�ò�0О
��5�W�#��J1���-��w�}�}f&�__���^�+�=ՑY��P�ם�)~,����ZH	a��!b¿�����������)���Z;���A����.��6�H�y��Kx����e~ޱ�*�o
��YTf(:���I~�yu���dY�@� �S�vTWDj�%�
!��p�7���������}W68��V�	\J��'��)�RA�X��u2;2������a��qk���L�y�7��&-�9��.���ŁyC��i��Q��;H�M�r�搪��07.��� 6��\��R�pp��ނ� ��54�p��\G�-Ƥ�whT6`���D���	5���Az����L�ªZd2��ȔV�Y�ݫ�2cVX
l�`���4���p�����E܉Q7�|��I3�F����{Y�����=����+������ȋ�����XyW7�\����Gp�K7��:G��wqK�Rl�[�M���AL�GM(��q��t�'���>M �3uh6��#���{�}]�Po��:�����W�U�1޼5d�y�P��D�;�����ߌ"������n���| p঎qm��k�PQ��M	 �)��W���X�N�x�[�9��裁����I�˾=�!aI�V����q���Ǖ站0}����'VO����[��@��"	}�3��"j� ����G�A>���漯�f�>�#��sL�A�W(�,[�(:� ��%vS�%{��-<�ã���N����ض��B	x��ݷ��
8���wVW6N~�̠�	��Ԍ�5�B�L�*�_K�)T��F�Ryе�f���Q�~�Z��{�Y*.�Z�#�����m���,�{E[� ���؏�e ��u4>��eԗ���ȩ�n� ti�}qs����Cy���"�'D���{�D��\��g��D��*4 �7x�R"�lt��� �.�O���.ְ�,	����X'h��1�Z�/��0��^մ��Qo@_�z=����gѶ��T� ���ù�������N3
��2 ��i! �6�3�oYy��j�
]�������]�.�p	�);z�i/G/�*���.h낗��ˑ��Id�]h��?��n,OaD�$�qaUm�Q���<�xY�e/�9LF��_Wc״��?����uh�0ė.5��_�n�G���@��|ؼtDc�M�)dy�O��B~V>��za�L�)	�+hQ�8ĕ#�]"H
�t#�v\o�.ܨ,#�*!q2�	�w$XS�G8W���o��R�E~ԫo*�J}�I�\D7�����/�>����	f�s3j�-��@�иS����r�Z�|���M���Fc�Fm�<��p�R��.�\�x������w�Tf�JG)�n��<��-x;JX�<� o.�DT�C������w���#0�@/��ࢲ�l������4��عU$29�;u��&&1��׭�ט�̉?zi>D2�x�|��W�x7�X2�B�c�F.�>9�z޲ݦ~�֣�W�R��E�^�(��.C�
�pKt_b_��P� �UԆ8g��&�����iR�*�2��{s��9�6���n5ʨ��zۂ�f
��+�Z��N>6z��S�.Ka""��:��G0|`5i��#��K��jf�3���j��.G#�u+���̭ ���:m93ö�5�����g���2K�X-���K����I!����>�upI������t�/I��]7�&�C͗{�
����1�)�[c&��6㌬��F�VS*K�J2��Z^X��AY��̝��Q\{��4\1<q|f�w#|
�M�Ep&�^v��	
�  !�^s�@	����@ tP�#�UN��i��ąI�"Ir��h��R D���3 >}��_�a��SW��ζH1���A�V:$�؈��}�︬agh�37g��rU�����U}U ���4�69�D8�^��䃇Q�Z%A�)2�2��G�/�{��=�n��3!q1W��K�U�;�uy�� Y��n�uJ/�	fG"M�%�T�
����� ��<z��y3V2o�3��NQk����eޙ�(���F�>�]|q���Er�Ll�7F�v�����w� DKJ���#��?��iv�.s���MI�P�+IԶ����n`>1�7����~�Aǹ����Нpx#��k�
���S�0׭�O�urL/>7��6�wf��n�GZZ�0�x�9�֛��Wz�f菱��et5��,�9�����B'��͑?[	�8�E��+���?Z�Xw�j�(������7��
zf�WGL��ާ\t�������!�2��	����o�~�F��B3��Y�]w̔�AŌ9�d��9�4�*�B ��E0�au���PM��CA�2(��`��T�e���p�yòG,[��˧k�V�:
���C}���͸Ȩ@�`,���lHt��Aca?|��M���jw	�0�Ԃ1��P�ޕ{n�Q��q,�uh�
�pr���	Y�y�0<������R
�0��-ᾅl��s9ù�H_mc]�
�����~�f�s�Uf���#s�-��ӧ�Z����񄑋���&�,*�)�4M9޼�2_��o��`|/�1���W��.�J�k��J疑��LK ���� �-xԫ_@��fw Y�� �� -Ap��\C�:�5<���S�[�~�@�|c�/�E"�W�8t��6��N'�D�A�fI�r�(S��N�m�(��v�0$�P��"�SۡI�>���0���HΎ�Hn�ZǏ	lj�}�X��mt?\��O��H�\����~�f,L�l<q5}�IHp��`�E���0�]�O����g��1��kMp�C�'��]7�ۙ͢��Фh����Ť�[����MI#�f�E#	���\e(�Lk���uos�A�n5P�6Q~_������!�r�:�(c�p� ع��<�o�s��_�R���<kJ�+|����>ť����5KQ�HX�DM6j
9�Tn��ȡ��|[A��z����@tA!��dE��Ѩ*
i=�<�H5�����7�k��v�t૳)�w��f콴���W�r�%n��j��{����X���	�j���w�/*F�u�'kxr�s��R�)�"y�f������ӫC���f�n1�S��X�qY��r���Kk���č9�2o�A�O�j#4>Y�c��!��Ef�ξ�
-��h�'���ֈ-�	�'U�H���������)�O�9,�%~����p�Ү��ޡ�A1~���,y3����H)���0���
��pc���"�Fd%m���"���K�b�����_��Bu�h�s,#�����
�ͼ`]�|�gh��9���U�㫶*j!?9���&@>x��_Y�-��w��K�3���Q!����8��܉e��W;�4�7�E�ROj��cfT�Z^���n2��(чK�j���a5��4}��Ɓ4�К��{��>z�"D�Y��0(�Ud���"��[��J��Z#S��2>��b}뼖���/��j��H��5��.�:�?�l�8�P���xv��p]1I2عӧa�7*�ҸA��Smߨ/,����dT������i�Y!P��MљN�_����o�w<�������[��y�c�!i,��R
:%�gQ?2=P����]x�_���-`��kH�w��(�$,����{}��0�.�¬qA��\b��uz���G�I+�'�S=4_U{8���Ǜ9�AwaX�M�&�`~;�Ùē1�j����h��Eʓ�\�W���B�W.��ȎC��j�-hq��-K�3OM�(�=ɽ��Lz,A����c�R�4\Ԙ��O��]ҷd�:e*{\�y���%�&Y6�د���+Ӛ��H�;�e�@� �(��-P��7�� S'��S�(���U�EÖ�؍�ų��n�j�b���y��@<�$�,à�V��L>������U�aoT�-����.M.�e+��/�����q��� R��[]���U�=,��}Z[�ؓ4�`�@
��R�lX��ߏ���>���"������"��������\Nmc�|^��T�mS�wfl����?��n��/r��&
�7Zl�}5ol���D�;��0�ʰ
�ݗG
�y�xfަPF�	J�$�A��`.ݯ�w��z�92k�mA_9�)pQ>�/Q���*e���`���LN���~�فӖKM��?>� z�������a{kf<E�dnܟ��J���U�M ��_�lW�gT'����x�K�O3�#�(��1���2[��-@����,�� ܋v��J�l�S�k�4�ŕU�;&Ѫ�f�!r*�����h8%V�*ճ���D����e�/RT.�+&��ث����c��-��7+�������Y�\�����:���������xz�Ǵl�E~�X5	1-=¶��w�KR�ɤi]nv&�Ƶ6��;��K*-₤'���ĵfw��3���<񮇠1���`�M��b���h�u��ui�����`�3�:��l�g�}*:�{�4�.�Ḵ��(˪<�j6�1D�JdlȬ^x�?���k�FDAo�?]�mj|�֮����
QZf��g熚�����[u;â��TT?A.���8��{�s�����\�3^�	"B���;� 2�)��׎äӓ���;S�.�o��2KՎ�5�c�r��jH�"0�����)%�z��Ew���?`A;r%����.K�_u-'Vjm�M�I��T�u�[tv=N���V��7��G��H�p�Hr�ȑ���b�8�߸GPF՞�x[�k�;��'IbW��ys?If�{W����l��'����(���v�7z��}���!d���L2�6)컬�j��� �����ݸ?2�[MPS��Xh�~�a��Vފ�M���)�=�T1/l�.�G��-kbSq�eF�!i����QjI�=&�����V(c 1�s]�?��?�pW��c�wP��V����B)a,��q�0���?t��C�j0΁^�b0C%w�M�QG�S�݊�f���ej����mZ·V�i���6y�
8�|"�K$+J�Y1�{˨�U}7�	���%�F�`��U}/��1�Q���d�≖�0|�`g}H�q�@�6������o��R�����G��/GǶ�?\��} �JF6$��T2� �ӑJ�(�g΢~8��rЙ|[��e�٢��F_Q�+%�֋1lz�Y�\�MJյ�},Y�O�CM��V5�/B%����b�L�O�Hi-����D}6"Oo�ӛ���o}�d[��ߜ\���9)��H���j'�p�G�*��DB}�4�9�,�f��PO�w�1�V5k_�d��؅�y�C�*�{�C9X%X-EN�l|������l;��X��/V@1l�
ɴxb��9���!&�nyX9o/)�\Ig���Jq�㵂�9�n����(^�v^�u�c����6ޚv��q�b/#(y��8qy��pS|]R��rǗ�f��Ն��LW�KOr�P��s���R���gY�P��W#�[��E�����~�n�l-J��������
.e�B,���kN�F�H>%����Ꮷ�][J��ܽ���)��2���X�F=����9ew�ӊ�K�,Y|�3pUk���m�����7�>�zʐ�
��f��l��R#2�R>�0���s Ve��#�/6���=��C ����<Yʽ�Cx�MLe���>K��O,	zc���-9��@?(Kc��u�%�����L�ԍS��b�p���	]&W�+V:�gP͑G�%{ƞ�xw�c��0[�퀀?Ĳm�X5���f�@�5��5��N��3�l���q��3��g�Q @Y�Uݿ3����J>��T�ÜX�˖�	�rD;��f��	�>XJ�]�c�N���Bs�pwT.��sb/�����\�`�DN,ث���`D4컮G��>a(|����Ǭ+�9T;�}^��?�X��[���y0�./�g�<�#��f/������Lm!* y�4'�`m�o��\���Q伯��nj$!(y ����-��#�k� 5������9���	G����������)�J1�4"",�j�nY/����ڧ��I*� �
�B��V&���Ց�^�y�v�A���7� ~`d�}�,Z�0�����&/5�ƍ�Q�^}R5yw�%�0p���+�Y�[�jLzZ��>��u���5�d#3���eK<��"�Z
k@��DB�J/7�	kF�0?c�| ����T_�TsN<z�o%�c��<�[��"y?<����U�=��#1��Ʈ9��S�O8��P(w���%��bN�A�[��g)K<�$T�H O>�dW�z���I(��a�?�����	L�~�Q?+J��[g�3"1٥���K�4�GŤg�m��% ����i��-�̌��r���^�f����J�Yao�E��4[I-:_^&̪���Y��d]�x�g������T6uȟ2A��܃|�/y�u@�x���|(��&Hn��-yJ����!�����U�f'��k�/�r�uɮ��[G���S��(&�}�{?+3� ����Z8���^�h,�u,0��@:�QxM��CH�Xc��ᚚ��p9%Ա�WIq���-�+aa���UO�W�	8g8�����4��'���jƐĭ�?�R�����jOX��?w�N�Ԅ5��+�?��<W��/0�xA�Oiyg�%��Md��sgA#@iT���2뮈�Fj(�x���E��n�Tc��4�x���Œ*�t?���@�)��:a���������Iy9�Xm6�eM�ݝ����-gQЭ}B>��)�ٚB�5'vHp5��mI�x�#�6�*��en�E���7���z�����#��do�$	��r� J��|�X4
n��D��^�>�	ч��r��b!��i��SI[3�MMd����ǡ3Y��P�-&�\r���^@�W��;��X���+����G��%v����Ǥ��Y�֜U�t�e3�/f7Xsu���~Q��Q�VhH�������~Q?��H�ӿ�{<LHV[��V��i� NG,�m���a�8��6t����(J^;�N��O���V`�Έ<s�X�a���]oL��^��� ���*4�Nb~�3�,BUQ��@��؏��R����fٖ�~��l��.���	�6vBB��<����@�+x�����b9���G��|.���m	x-��FV0��c8�<ߥ�p��2�vrf+�O��Uai�Y:�5�'j׭���:�P��vm�A�Kq
Ǐ�`�m&{}rQ�_�Ő��2}����;�sT]�+���.���
y��9A�G%�g���@�����.��m����{]��C�ĥs��\\+QECE`k����R)9��7�m��>�&�z4ֳE>:��%o���q>0��N׳��V���YT��#[��(5a�s6\j�M:�kh�(T��Y��0Vt��e�7�b2)~�ʝ\��\dnm��?A�M��"��Ľ�Ħ�֘��y�N�'qi�"�8��PR���(W^\�=	�g�}�s"Q�v}W������ǺM�q�E(��y7�ɿꄬ�e���K��� /��������� C����1�!y�Z;�X�3i�Dk!�K�*��&��h���9U�?��"�Y����VSy8sњ��C;��R��v�E����*�>�@�t�J����j{��*�|C�#ƞ�Oo���S�E��K���t��c*�(�o������d��Yo1�v�dJ�ļ�	��b.p�7d+%��|�MC��4.�.ʽ�P�@�/0�W�t�PX{, ��ff#i������?_��<Z��L}��A̹����1��P	WS�<���ޱyȥ��$�L��{C�^i�m��3�~_�ڢ�JUl�� /u b&��[{8�m�V[<yć2�6�~�:I,�r,�ԟ�Q���5�74��yU�{/�	2)�������Bk�����N
�O��,�
�)�疹r:ʒ8we%!�H�u�/ף����Ȇ���{��M �_\DA��:n�"��n5���X��x^@RH��N� Ƹ�i�gC�h�=\��:ߑT��;r�$���ð�� �$�L�Bt�AV�n���X�ы������7D`Z��?z��#a�"�9u?�G�K�	�2[DV��(_,�z�����}�i2ԍ�t_ӈ��Xu����݄���E9���V������B��8q��]ݙt[5'NVT�G,�X%��9��k���l_��Tug���	f1�@v�<v冃�W[�-����A�;��~m��6\�@�?O8�R���4�I�����
�N�*���UD�n�ߓ��퍺$��T�|�Ga�C}Æ�H���v��!j�n�R�����v�H�P&�A�/!� �K.��6���2�U$:~�C��Ќ�}��JC`����C*��=�k�6ek�T��/H�sR�s��i]����÷��z:���*��+�?�;¾�a��T���R��d���
�3	�Ԫ����8�Y#2�sh�R͍�[� ���^K�;X�����=����Hi�����S�8���f��q�и����=}s*|��1DG�e�a&8��郈��!���m��W�@5�4� �7���{�=k��r?�¦�D@r\����pKQ��&Vo8������xZ�!����nV�-�c�����M�!�< ��X�I���r��qp����tT�4t4'a��Gm	�W*��h�n�\]�沜^!�V�+;	��Vv����/���9��!�8�?��{�{vC�f��=Çm�VF;��y�o��A�R�idu���P�W0�|�z�׳yߟ�Y�{��I�?���~�ۭ�*G1`�������"T�0D:�g�Tj������jN�qBg �ۧ+�pL�����b
��c�P�rsA� �;��s�c�g��Mq�~BG���|��Q��[�^|.`VX��?���2�Y悚�:=Iy��B�HC|i�*��d��K�5��QN��9��K% '�Ї��G�����s��p/����si��Zo?�wǶhl��}p��\�U��ˌ �]�B�Q�8��v�TIb��H�TK��S��z�;9��d��.rB/�t:K>Etč0��I?v��P@��t&���&֙�3�R�
�Rt��%;��8���]���[�|����b�H���N}},T�_���im�mv��0`t�d��;?��̾?I�e״���ߟ�������l�6�hS��̄�\��$�0e���)�$�N���Ϡ��$Af����Z��y�������ug~ƽ��)�I�@׬8�q��Ԕ�ۚ��=ORT�]�U޺������US��:��y��U6������`h2�� ��s"()�<���1l���1t1s����ύ.4�4�{Q�z��A�o ��uO/���h �[��w�
��n�'��Φ�5�
����zmh�D��5m��9?��K��*"X�ٗ]-[)M���S���+?[���$�7z|�4'/�XG��Ab�j��:I��'[K*�X�6��$ܙN�_o�C$���o�e����4�I���ҕ����ի:ӫq;�hO������i?'��kΧ�h��DM,{Y]�2�)߾~��X�\��`qte�>���4R�#u�)����VQB�W�/�{��9��C���*��}{��\��=	�3��G�
x�B�ͻ��R����-���Ө/����7i���k�A�$b���LҀX���/���&�\�m�`i�b�\}Z �IZF8�x��A�v�y�M��d���� ^O�_!�7�9XS��(��zNBk�<���c�vx��I��C�k9�^���>Cdķ� �J�<X��z���G"�w��xV �t�L4���[9���i��Jo��[=�E%g�M܅3VU�:�'�3UО�s79~�w�N���q�.�L���7Sk"�_�l�:#�A��5ܧ�L�N�=�(�T�Wě�_\������l�Nϻ�$iT��|�A$���\�\nTA��/�k�M~L2w��z�V��Q�NMs*���TWc�����Ě���6���
���kEҀI�A��e���MB���<�2N
�a�|?�L��I�/|#��G-2O��Oc�#d��or_՝>�{r��A?R��ݬ�jSQ|�($=ڨMyN�z)tM��׹�#F�/�|����O�aS� Nh���r���W���;����Z.����>.gN2#('�ځ�t�xU7v��-�+W�|�W@x���3:��6���^�j��1�'M�Y���#U 38��T[F�Ec8�N�c�7�� >�bV13�̾WOa��_��^N����Ն5�\3���܌�?&1*���h��|�����<�"�e���r�:bf������9w����NP�Do2���z�(����|Y����S�Bc�C'��_��r�)v��54|'�jI�&2��I9�������u�ϐ��n�E4rF��A���V��~nI&t'��|t1��T(��m�w�����닂j���>�O�13�ÚPHd�w����ה�jΛ=)��Y	]����izxE	��������ݒ3'tkY��I��9J�v��\m�A��qz����U2A��o�2%c�I�,�:��~�z�#G�]7r��CT��m��H"��J@\�Bwϗ�W����6�ܖ���\E��=�5��"�����/,H@�f�1�4���G�{[r�sl�)�$eOZ���l]~z�C���Ө�4 ��D	q:�GIq��E������}�؛?���%^p��i�ŵ;」��aw�_n�h�ܴ_d�	]��ǌ�~��y��T�.cŧ4e�6�L��l��I���ث%Y�Ġvz[��ũ� �y���&�W�~cx�0(���O�����rv�{b|�0�u�A+�sW�R��K|�f:��P��9w'�d�Ie� ��K��zg�%N�b�M��K��R��a�I�8r��GR�e\è:vh�>��S`�p�q�B�|�s��Ƃ.Eq-�d&)�w��{�������x�b�FU���@LX��<_����"�����̈́�����T��Q�NZv�yBI�j7-���(2��� a�lnbS����,+�a�_/������Q��sz��������^���܎�T}ޠ���-�ʈ ��t\)�2��zR$������r�%s��dv������!`q5�~W<����Z�۴m*g����p~)x:�
��x�M�d�6l%���5)�|�~���#�b��G��с�cpw��E	���A,�o�����j9�S��m��`�������2�ʦ$� �o �,k��w��&~��o���G�Z��.&��&;"�����b����nȭ�?+�.�'.� �0�+V~�g�J��l�\�]�fŏ�b��k�1>�Lv�:�0�� �N�E�Jw�~�2R�3;%�QF�e����*���Z�I<�
��"=���h���6/��v��Sګ�A,A	�]�y�&�@꟠M�T�Z�s���( 8JV==CK��C�h<�h>@�9-��\�<�3���ok	�'+<NZ���
 ���t��,��X@�gAm})[�Lke�l���@���]�J������-Hˬ�"oʉåBe�+Zb�j�M�?׉�~�OJ9VՐ���H벎�$�c�ӹ�ç�I�=<��Â���%L��k�l8�����ns�pRbI[�)A���g����H��L-vaM#�W�'s�#V�	П�Xg��ψ���`�_I���|���ry�,g�����a�
�~�pF�a�K�Lg۾���ps��0�SQZ����6JEh['��д�s�K´��{�E(�d������	k�\��n I3۟m���+����.{L��2)ؼ�Z������k{����ud��M������Ty ���6���N=#���vE�(Ȑ��r~�B�c+�E��xKD�tO��H�1��*�7 �q�ǜ�?�_s9�"G�6ƥ2����0��^HE��y�{�d��3�B�(�C�3B�0�_7��J����;���>�5 ���o�mD���݈�r%�\��O�N[&�h�����ghqRO��g�^����,^cs1O.s������'�\��[���Y��Q�O�h��K�����#M�R��8j�VL����"��[R7NR�
?�s���i�,IcDM��`���I��u4�	�9^�ѓPy��g�#4�D&�8�y��D��x�5�U��i=�.��< ��ݝ���lW��;w� 4s�,y�vҩS��7O;�R�q)��0����+�d�mc#�����o��]1�=zX`��hx>ۏ�:����5�������z,�+�>?O�m���3���fY���íum3Z,h�K�I�Ú��N ����1<��!��
N�u��A��{�<Br��"�r��������������+&yK���v|iX��@b�7���������`A�&%t:'�I������*�'�	Dv��������Z �şp������b��U� �)3��gkY�\.��[�����
���@�p#���1h\��&�.9��x���g������m"�'�U��ozn�J���7̃ ���G���g*�pB�;���~���A/�Nӑ��P8�1@2�5�_�t��o�0?�JN/��|:ș�8FK[��J�v�)�a��.���&$ue�_L~v �쿅-�l���6�8�ky��f��k�'������	Y��Sa��l���M�����c7����cg-,Q��S����>r;���Z.�r��
UGZ���5� E�؂�#�{�d
��RՉ�9�Ƚ��<�h=�7��Z�ա��
t &"6��#��xZ�פ��]P�V�j��	�s~8)�>�^ �y�7�dk���B�縯�bdX�tL�E*HߑZ�1��&b��7��i�@��7���c�Dü�P���I�	>�#���C�6u�*��1���������$`�����{�|B$P�CN̳�> e!���~��y�IB�%T���[��K�m����2���MIgb7�븸٤t_``���ƘS����V���>Svk��D5��+��TN��z�����>���U��@	PH��z���C� ��'>6����������x�)������ƸYz�y��5-��,�!�v���Hk#�[i�G���ܖހ�
B=��&iU�I�p�;�߄�J�noy]?����ƥ�>$J�Ef�L�"�|��IC䘵7������)"���N�~F��WR�h r��Y�����>�~Ь2rf
���6-�B ��CڗC��oL�`�_�@���`8$s��/+��>���M�f+��c7�w�J�d�!!���yK�����;��a�Z��c�"ɂ"��u 9����7b<\|����V�$��9�1���Q����ب�ǵ�����roas]6����	(\���0b�>2�7�2��c��H���%�D.˟YLA��苳Um���"'e��\����K�e��O�4VS���4>�#�d�wL��x0���!%��L��vf���p�ge���Ɍ��[6EQ���$���li�f��kd7�a� ܶ����' ���ˑ�N��I�N���5DQ��Ձ���s�/Sr�nf�E3���t����3AMj�3�M9�!��K2h%?�d�p�j�̴�����~���/kkי���؟����"BY�#I��@&��-��3w(U嗹Js��X�>�z��AsέdV�͒D,3l��t��i�#�c� :����*C�uz�`-ՒF��'����5���1��K:�.Z��G�q�G�n�=��PQ~�gԷ|n�߉����6������,FݧI�kx�I�t��W���ž�O�4/��	�r0.�'���pÇ~K��4(qb��J֛)�$R"p�u�7�����FR��/�e����,ujj��ӎ��+��9�E{"`��^��:k�Ґf��d�3u��+Y�y�Z�8:H$52�{�0E�R���R�!G�l&�՚��P�9��F ����*鐴2Ŭe��7DAT� T��=��bôL5L�끙�(%�1�;�c�������ߵ�@�ű4�{v��x%���Ġ8�ʪG��N�_K
{���j��Y�.@�¬AEg=���}3�'U:����T���z�G�^��fYo�D�jS�s���mV4�
��B�s]�[�p�V�|8k�E:�!��/��� `8��ڇ�9��|�������q0S��H��3ױ|��^EՂ�~0��S#f����Aq�k*��/�:W�d4��m����i�����	�n"��t�H8��m�ᴾ�]`�V2]��hj����l��e0��B���'TB�	���-�8�����x�H�x9�F�xZ*@�<g�2��&�_�;� ����i�}&��69�]� e�������G�V�x6���j�R���N�6�>�'�����O����f˞��JA)o2d�W��!ꃐ�LU����q���U���-u l��Xa���^�0e\F񀯶���^�tj�?�Y!�st~~Ϲ4z�cȀ��>Ɯ� ���{vP�Z����Mt�c��<,�� |�����!E̸�R@6��2?���-����8]��5���q�~�n�G�L���yp)L�u���-��\S��.B
dԙt� -��sW����C$|G�Y�����l
�9I�=՞��	Ӵ���T��
�WKɐ�+! �Z��)��]w���sY �������,��m���ҽ�.��n��UךS!G���T��� +�$3ȵ*�{��n[bxu!.Q�yS��c�ގ������������/�3�[(�N��@��M���8��k����84�*���=��Xм�4��EJ�Ϳe��l�p����ER��صg΃k���]�Xڌ�ea1��z��2\��`~���Ps��%��d���_}H��+�MXeFS��P �EJ|��5�u�����~�����o׳�� �zZ��|4)a�5��N���	��{\��+O��V2>k4U[a�󓽼r��~+zG����4���[�4m^����2��g��1O��y��_C+ݏ�W��/R�x�/O�F�N�3���=@��L`!Ԏ%P��?����^~�{"�.�PQ6���2��q����f��j�wk;o�ј��n���恔�6�g}pB_�����9�B���U��� ��7/�ȐV���{$_�5a�;mշ�I�u@���D~�͇�/:G�j��}#'�۝��D�5�th��G�^�!w�Z=(k�t�DAcO3VB�y�;������K��x�%� ��T7�9�d��������7�7��F�Q�=)	'=b�ܹ�G/��U��]��9&��=�#_��( ����ҟ�<^ݫ���5ٍH�^
b���ã;��0��9���xa��(-�ږ�\?=����`�y=b"��'͇K^�;�{4�o����.-��{4E�2�s	a�~ �-��o� ��m��뱣Y΀~MZ���~�vW>�<�n:�CW�H���eG���I��@�3Cd�9ɯ�>��ܢl�:�y�o���dtE�c�s��{�Νl���w#�>o�G��b \!�q��/u��a�8�]-�I�#�|m��F?CT����%����]3�v��7Ԩ�+P����
�v:�G�����)9��R�a���X�|-��۹{(T� �ˠ��r����|�vO�*~��?wGL��:�Ed���I���}Ɓ�ЈB
,��6�O���U�L��������(���Cl������H�")�
oi�om� PT��#B�`��5��'�>�>%yH�3Ǜt�0)��6������Q����V��E6U�I�����W(�ƶ^�@� 7��dT�����t��e{�:٧#���������^Wsb
51[���������=�����������wo�Hwl��U@���̲���[��$zA�ks�D��5��1u� 0I�$�-���e���gI�bmQ�]8�ɀI�Q,�EC���Q(/B�k���Wvj��|�h$@l�ӡh�C���ڳ��㞜�<[Ȉ��0�����'����|!ڽ�0�j�g�+�d8��9J n�[7!���q)�e�f��EˇЌ情��� ��o͛1tĸLSܜ˨	�+���\��Mw���1�w��
UJެ��l�,�4V�|
���u&/��lTc� :^�'����=���V~�إ� "��S=a�b'�B\ǟa|Q�-�p�~(�a*,���@������zs3?���� 12pzK$�%�?��=C�����3��y0W���6r%go��9m?���#^׋z�-�Z�~6{n��f}6��pZ���6�_�ʈ���/ր�w��1B��Οf��t.�է�֡7�\0x�|��I�X�Vh?sOK���䠣f�Nz6s�-��3��_������y�qT����f�5ڧ������ء�{մ|����˓��5A�T0�������IG�z�1���4�u)(�>3�����d�>��({��g���\[��6�\��c�bpe,�.ÚC�i�-�S�s�����3�-t)A�Mޔ�Wi\�&Bv�ǅǒ���J���.&���Es*x�ϱLk�E�51.BH�%���D4M%@F�!��=6$u'X�?�&�� �������o�a�  ��k3��~�u�2���F%����7?�kb�0��b�XK�%h�
Lt.�p���͘{�����5�x�p���/q��6���R��P!����;����3}r\&�$nѨ�<���ZT��]�cK(�8�T
E�o�꺢Tٰ��;�ퟟ�v�1����i`(˄p!�"�������ѺsQD^�� ����|���u!C	C(�M���*��	�@	Q�q�	�#a�;>�K�������QD�v,�S�N��v���,5�:�p�]�^�9�µ���YX(�|�1�q�[���ݍ�1w����x`q ��S��# �#����A���HG�F�,���eV���͍RSp�S��gT��"��J���$�;x\nD
�3(���A��v1o&�򤉩Y��lQ���H!�F<+��Z���p��� X��!��()�K"�u+��W�%߃~�3���Ks>ft�Ě�ns�d	b	�p��[vf�ճ.��A�Z����Wz�PE���"�(��$����;��6#��A��,����-(�Z(��?�'��PrG���{�W�_��r�����=2�^�1�:�,��!���}x��K�f�4�����?��k��c�썁��#�!���W��U��No�S�p�}I���fo Z�T�	J*͇%bvz{A��*["e�S����]X�����8�B�m58�H�N���FR+|�oW�J��k��8�&�T�PXH�l8!<ڱV�:ZBh̜�E?�b_�G��'�d� ��ۍ�����!�I"b_�۾��-��/	��yүۺ��[��Z�����`��73]��w\���̮��aږ�N��@����
]t�3i�.�$�Z
{�VX��ZL��`\j�Nfݰ����i�}���J��~A=���]�,8��D{��/ɐ�'_�~��~��*���gƢ�4�*�>�IZ�}��J^mW\�H�H�tPd�K�����f�X�Εݐ�O̫��*�DV�y��Z&Jx���;�pŪ�ɽk��ٲ>�Z�-/���T�9�9�nݷ�4�r7��]w�4&�G>s���=��-̜�a�?Ye5΋}�O��ʯ�ԡU2�M��u���5/M�͢1o�KJ���"��7s	ČmH�� s��,��Cy����r����7�s v�-0I�{2T�n^l�Љk���L�,��x���-Gm���!I�45����<�������y���!���T,�y�̀�P�c�)�9�*��6�ې1|�r�\���#W��
����!�X*���4��.VV�nTub����Jw{QO�p-��g�W	�pN��3؅��cf�r�0�n;ԶA��RO�S�y�^��2���n͚����G�"���y�kN�z�AVJ��"G#���DҤ�Ǘ@�O6���`�	����X�'����/��U�T;���Z��=�<�1wz��L+��p�[�C�0�P�hn:��iE��;V̰�F��+��0�ʹ�fU%O�C霽�j}0�q�Dl���(u^W��Y�wuϬ��(�~'�%��t7��f(O� I���fMd��8������\��������x]���'`g;qU�K��ӊ�޻ƙ3]OIB��4)|0�f	����Ҩ�T��"ƺ�	���(���>̀x�%r"MFhL.<���-A��A�8�6Pl���,;;+�d��&c�]�j�+ &��^u[xj�C2�����{'y�0t�W����;�T�ݥ������A����#ڲ��稹�(���9+^j`֤�(�L��y��L�����=��B��rk:�nE0�������zh���[-0��F�f�O�)X����l�'�# h�nz` �n���Y����C��$6E���5��9������3�9��S1/u�e���T�1}�O���~��� ��{_a9'ۋ�h��9�ߙs'���&�^>r67�#�ܣ*?�y0?���d(�|0D�׸�}�r?�Ƹ��"+g
QJ2�J^��K1�Q/��{؈��dxVs�`ɲ���h�,:��M\�Q:Z|Vx!��}M����,��v<.�1�A��T䋕���kބt���#��6t/4��xg�/`�N���R�X�=�j��{?R0�U�[~�	���I�o͈�B[zƴY�
u�AT���a��Z92�
����6)��ir�7����	�Ԛ��^|qd�@������Y�N�S�Ϳ�z����Okv�qxbf�qf�cE�9���m������nW�v��-O+�8�W��Om�����-@�r��Z��A@��'1�SQ1�U�4�_�@@JB��܇�H R+|��oC�!F����3�A
 n���-B�U���`�� �iZ"����ó ��m����̒�t/;⭋�K��Z*�I4�ZnҖN� uN6�=�Mq�{����
A�����c���sB����+�sx��YDB��`���J�K�gsN��$?���G��7�~d���z����p�ؐh�Mt�x�'қ�qw�QY�؈ᔽ2اf6�[=N�왗��ׇ%��4��� �*�>~>�&Ď�q�����K����b�=�e���a?s���)����q�ϻY����s9��~�4׎�.�u|����SL&���;������ʈ.�O�!}����Ä D���&V�]�-������������Uf�5�=�%��ϭ����bhˬ(����9�8
�	���zrV� C���VK5�,H�7��u�_�k�Ծ5AaN_��qϸw�c}��!��:��;q8G�[?b�T����yx5O���`d��HUk�?�O�DEN#>"�8x� �5�-��tv�\��I���H׳��YS����"N�SQ� K��XV
����)�Z�[|��H��]H\Y��a7��3�(�<׎-���6��?��y�Ս��g�"���r�Ϸ�0�^nw9�U@�ҝ�����R�Җ��(�����t��_�3���������KI���w��rm궥*/�6�|r����A��=���$I����ٕ̀�ݕ�������-7��[�u�T��gUG#	C����玄�$X���������N�����ͤ�����(,j�s[���#�ry.X屯&���vJ�Ň�n��zǓ-= )����I�ç[^�۞�PzR[<��l�+�d��J[%%i����#��!����o�q�iNT�؂�	�YP�4�'���{�^B<���?j3�;7�{S��C�$�7Ԛ��Q8���n�Y�tG&�B�tץ1(��y~=e�$:�4��¨�́}E��Nh���cό^�����x~X�^e�6�3��5nS�b�Ais��On�' �?
������պ>!k<���$ J�{�\}��̃��F]�(�ы���p�	�I~$���V}���>�b?u�T��O��N�o�g�0C��!t)$�v�no$_>i�io;TvD7X�&�WE��-��!h"���06v�����f��/`�J��������9�Z��J��-$���uO%�<M�:�d!�6��ݛ�e����%���&M���X�
 Զ-�Iz6H���H�UĊ��E.�q�����N�Wշ|��I����X���F�$zG�a�˔<��$y�]$6tQ���CC��Ӎ��l�/aU�

��|�_7B����w��
+��ll��+Bt�^4O���s4��@����Yu�S��n�9�65-4�Ѽ��U�����Qj<���u	�.9���۶U]�wI31�z�*�^�{�.}�����0�]�!�TBY}�nD���lZc{�����JE�Q}b�g��ޅ��GZ��&��G-�O� ���2[�S��'�y�)ӿ�3=�^�:~���!$�~��8���������F�C�1���$��[����2�x�����*[�D�4��Q�n,����/�>F�}���j��9
1�1>&]X�T���U��-��j�?P��@���|�V�q�w����æo��^u��rV�_foT]m0(��Q��C�vV)i�=y�"<����8_1�n���C���+��KC]�q��������qǘ�Ƴ����/F�K�u՗�d�ᮺ��H��&U�F����7EdQ�X���NT#Ϡ�Q��W^�L��P�L*���c_�f��~	�������P��O�tп� �^���x�5-��ax����xx�%����N4~n����D����}a�l��|�>�)�0P�]/�Z�L�l��7��m`H)������o3Yi��Gy���`*^��DR{Q�i����h/�NY@Ȧ҈�dL�9�{�~�0�P�O�sS�٣��G�e�j+f��F����:�������*:ݜ�A���}Y�s�x?:0��:R�φ�1q��@Z~�u�漲��6��2ז���#��G�9�hF�8�H���JtE�G���r��h#��bH�]��*F�5������V5�f!o�<6_��F]��B*��@�J�ki��� (4˻�A��-a������;w\�UX�>���1C�dC\���~Ϳj�6�� Q�`�	<Nj�y��g�$J|�lʕ2�(B"���PbL}�X�q!��D�
�9�x㚮iD$��J;,��w�zΝ���<7/L��x}'�9(�b��>)n<Q�8������av��N��"��O�)>��5�$V�2AU(~վ������U^�sPAd�Ʒ�􈔗��?�)��۰M�m�/�m^����=�v?��L	s����h�h0�7G7�R��*��U�rJ�G�6�1#L�wVVi�#�[5���N�3�Uv�id��b���2���!�S������"�j��4Ħ�ӝ��#�dl��[9F�ʆj�Y��� UӣA������L�`�{��������M,�#�S+Z�݆f�	����]�}et.��U���<���'l^z���X^s�#����aa7�^���E3=U�cቋzz��1�!����b�@c�U5q̗�Y�y�U�w �I�}�;b��lri��d=�t�9�=�yK/�TJZ`����?:�i'��#2��ں/��?p�rа�kl�i��� z���8C��7S���­q�H���I4���{	�mp�?Rv�z�n��Jf�����fSFNӔ�����r�n����Zr��^�����QDUwZ��
��7i�x�c��\��א���2�Ie5��LL�ݮ�}�9i!&U�8�!be�Kv��f�0a����ڽo�gN�xŌ�Sb�neטnVW�8K1�x��\'(9��m� a�M��i�|tߵ*R��᧕�������@Bk���^���3�$K�اHα�R��V=�6�����=�c���(VK��~�`B �'
2��A�!���g�����hӐF�BǀG��t1M���u��2&cI�x�ICWw��S=�l$3��D h���y��h����N���E��o�gaii3��Gp�z"WQ���=���(*��XJųl<���D��~\.�P�h[�Ȇ�B�䯙���L<��R����[�4����U��ܑ�I�_{kӏ���݈�87��鶳"\�C�P���.��S*k=A��h��@��Z���	x�s�V�ac� ��id��l���Q��O�� �L�ɱ���F�CLtic�%B�P^���4�[�+R�J�o;��7g{���?�D7�O���3�+OGLo�=5㨆Np�$ؐ�=�#�ˌΙ�50�sЧ\=�K�����2EK�ǲ���������58)����=�����fϨ�vH��J�O�݌�p^T3y��Ԋd�x�����mT�u�2@Ư`譥�W�{%�$�v��G�<e������h��.,eH5D#7��7iRϟ���uT�)�
�m���/Q��<,�@6��̈́8"���*`1H�F����qa�Ӌ!�5�Z��Lw�Ӛ��%�F��?2�Q1_uG?�ќD�����{Y%hw���F��������@Y�i�<����(^�CEL31b��I��)8���&3�
]2	�3�צ�M�"��oY�����_�!�<�u_��OK�G���ݨT����K�� 
�?M�����g2رr.Y �}��y�(K"_����j�������dx%��������*ޯlpW�u{�"݅-wT�"�ߌQP��DB,�n�>Wۏ&�/����s��8��r�O F}�pv�|���7:R1�Yŵ�8�ٕNrcr�!��P�A^kƮ����9�g׋�3�_〽.�����V���-3v8�Q���pw�飼p��R�õsl9��������;j����Z<��U�N�H�~U�~B���l���c�~9��k/������<c�77�a)X^��(�mK����OL�h����!���m��^[5׳���� {Z��r��Fޖ�# -�3ޟ{������o0�zp\�;�n�`�Ty�m?���x	��g�7�	