��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(|����	t!����YXRe�������U݈�NׂI��h� cw����X�`��\���� �o�H�RLҹ�%��!��*�}�\���&�!Ԃ�0�K�~�B&�p'�=y�wV<'���PH�y\�^'��Y�����������D�x� :
�$�<�W�%�������=\IX�xTSa�n���3�q���$��H�k�X�������(V(U��L���ٲެQCE�v�6�m�C��7�䬷iW�E_߬Z¸�f��G=��E;��Qc�dg�clE{��#�c�T��DV3[�=� ���w�	��,���̏��i�׷�^�v�/��t�rM#�5{S��pͤZ�66&-�º�E8��GhE��Z ^����V�x�)I(���y�y�*����J]@�r�������n+~]��k�b|6� Ӑٿ*)L�4��cx�/������e"ѝ�1
@��>�`�\/l�Y��bYt�M�s)­?>>ɦA{��>���Q�V����^qհ["&p�v���	�HU�Y���|q�&&.o��d�G��vV�7E����W���0��~^�_�D*�����
Z��pСh1<7Y�[\ɀ�<��C2^m��EOܲ`�w�A9c)H���CF3�v��%�'�� ٝ�l��l�m,FfA,���Ҕ�!]k@�~"עHZ\qE|�5���BM\?3�tg�E��	k(|��YM�v�m��S���D\�B��L�M� k�=(VB��?R���vbL��	�^�,��h�U�>��9�ֳW|4r�g�R����d>ߧ�kg��:��Ht9��L������+!�RN�;�M��ѥO������F�g��%֗����7�U+̔�<�K�O��?�(�e�1h�A��vI��j�����d�(!��Y�q�}c5)J�5Vs�zGaIA��R8�?G�|,�K�AkJq�����h�]�"9�Rbf�g5] 7@�neD�N��B&��ʰ��hM��"�|��T��:)�DB�;g�5��vؘܱq���K��O-��j�}�O5�[1:���@�ԙ�X�u���Q�h(5DE�@+�'�ŹŃT�h��H��ymT{��"�lZ���v��O����F�aΪ}힐ˎ�97�P}����9�Ʉ��?QBp|ӿQ�*��+vo�4��`�ù@�������q�4٧��bd��Zk]3�Ĕ�K��Lu����n�K0�V7�B/��i:�q�n;Ouw��ߝ��z��/�����-y��i��y&���lKm���a�L���bz��7�s��d�����^:�7�{�N���}���4���L.7]��ɒ����։Ͳ�&�@s��^�����f�ԉ�����OE���-�����&�2>��3��c�t�"�{�1�/ʨd���tjkI���A6iX�/�=���:	K��e�Rl��U��iEҋ#�0�ٵ��lxy괹(PN�(�hj�В�t�Sӫ`����~�`^�H�m���`�w_Q���g�e�nH���1��,�.��x�b]���k�[�K��,����?����+q�y�=��r���M��Iވ�pL`�6:Pe��z}Á�'��:ɔw�ު���;�;0��N����8��k� �ǲ�JV��4&��Êb{� d��Fp�ax�<��H?���K��b���kuH�	t��AT@�H��5ds�:ߪ����Z�)Jל"�T;��%�b�����X�Vk�U����
ϰ;^UZ�`�b��R��Oo�[��G:l�
�.P�8n�-�s�2HX�g�(@��Ή�R�֗�S؄X��r��ޫhnMC�td�Zq5�&��Jwq�g5&��u��2Zl)K!��_�f�Ǘ5�"t���̞�����G��6uk�V�E8��Mt�b��$�2���(��J��-̺��հ��j�D�e����W[rQ)��d0b��eoSV.�#�Q![M��� >� ��S>�*��q"�w�Q���z��(�<��,�J�pG��H "�;7&8Qڝ�AF=��Y����4�h�l��s%���$R��3ᒊ��,~5��hU��x��}�o�+��(<7�i����i	Sv��`Z��� po���
HE���.��0�a����QSݹ�
7k�R�e���j�u /D</��<�.�{o��9DL��	x�,PL���B�_�����2Xyڃ�ܥ�O�j:à+���(	KqlRy{Ev�6��-������d������<A���6U�m~p�jr".RW��L��7�b ^�K�Tos��[�"�\��0U��������o�`���N+������o�'���LF�<���"�CG�!���Ei����_�?
�#P�"~������-/�Hp��h"i��?��d�مq��¡�Ø>��u��[�*���D8���P�i�y\�>�,�t�9;ng�d�K����Z�2���X��tP���I�%p��y&�A?�~wo�a0�����6s�il)�n%ؾL��Kӆ��y�ɘ�y��Y�-qă{�Ca�I�����B��w�Xԥi�=e�8�A恱����rv�r�/+�$+�6�4���0Oe�쥵���p���f�O�Ђ.�aŶ;�,��)�K��E���S/�~�� +QM�1iۥ�~�/�U9�l�a6^�jZ0v�� �udا�F.��ɕ����az�g���'3Z��vٺ�E����:������|,�>��l�N�˗�˼74�$�S�pƑ�s &ބޘ�Iz�>��Xc��>爦b��ư�60�X�5�֜�&��O��T1Z�N��b�=��b�y;��)浨g�Qk=M�1ACʨ����30ְ�gD���G7��n)�{�2�c&��$��<��z�ϓ��΄v׶�%T�<�lL 5��4�����iU4����Y�/"�☜��`Y����υ���3������߯�{��%65����Pń˘�P8%q�>:ϑ%d�B){���ef�[K�; B�kHЀ C�;��`�X�TO��m�׿�:4�Yp��\���Uѱ��	����p֮�fJc���we�z9!�樸�g��a��!�&�	�V���5�`1Y����}A8�"���+<�%d�x�Z\���^�1X��7���8�T%n�s$.$zL(��)�Y**ό���H�^���x㵬04,����}`��bJ�oL�,�K��T��`1c����&2��ѧI�X<��ͯ��B���R��Iٲq�A�����S��(��;.Z����C�>�B�rnR��Sp�ѫI����O ~�ub]��w�l5��Q������&�Ǻ~�/�^���������m4����$���o !��8:	������ޱC�L-�L&˛���:db�����ׅɴ�Â�H�!���>��u�ʧ�V= ��l}c%Nϐ�ZA�Z��/�_O��Z�����;?�;m!��e��{��*,�H���˻���m� ;��{�L��~��9��m���k9u��,Au�xɃ~1��h>%|V��C�x����jj�	V�A.�B����I��3b�H���9�7�>i>�:5������x6F�
`v�GM������ǧ�dg⋖�/�J�T�g�ۼL�������-�b���UY*�#�`�>��k��H�+R܌���j#���$�{5��<c���, ����9�?	A�n֌��~DUԎt�w�<�Q&���s`�� �Z׮vVA��>��C��;hC�l/�F5�\4ɍ6���y(,���?��;|�"I3B��G�@�9�upJ��U����N�pXdJ���&0�� Q~Ia�A�v������=�����T�6�o��l��u_Mܠ��M*�zm����?��ː�7T���-x\���N�̻����Yɳ+���P��OfF&P�6��h`р_?Qْ��KR�HYA�l_�.s��6�x2
��cF��^ "�(N0�ۣ �����>x�VR'(D�-b!�s�A��7��%��W�k_���:[~�N?u�꠯UVS��s��e���b勜�/��\�v�3\�p�z-�/���o�O