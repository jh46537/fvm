��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�O*�!e��B��K8H����O���vD|��tyP��n�~��W0N����,�����Grs��!���d�3�ٚ�;�Id N~��ZX���p�*���,�@��f�l?Ζ��H�A�i)h�,K�[m/����mi�|S7s�{5���m8=�{I|l��O�ɠ�"ē�q0�}5���
�h�B�c�{0T,t�P��ǥ�Z /zlL(�n+�ѓwRּ����Ҽ��_�L���Ҕ�2�9�����@�7�y;cR%9.�L���wi��	�_w2%!�bP��u�28
Aey	L����^D�_c���&�>�TFd�����75g/%'b�
��")H�)�Tl����FC�{�	q�[۱@���b��Y�ݟ��@3X�%-<��H�.�H�a�-��J.�'#xa[oT4�U>���7�BLK������T�q�46�����ץ�3u��{?L ��y�ogl˳	{�n3��g��L�j��[�yD�A9 Bm��96U,��I����Gioi�H�*����Q��z���Cb�f$�����NX���U�4Ir+�y��M;G��~���T�AQy�].ЀK�p,e�r�p3&�=7�7#"�����ƛX���-�y��2QRN��B6��{�Z<�ʆ�{E�$��lbۦ`�<����4�)�^��r����\�h��r|��4da7�-|kv���QԞ?cfMu\N��w1���{�lJ�y�=�WmRq���`��䂽�
Q�YW�Q]�Sߖ:CW�X����7�+�'5����<�a��]%gު�x<?�Qm>,�GaLF	�Qn�%�Lt�@�"UkG���9�;��^�Zژ}� ������)�$�B�B`D��Y��(�ζl
��e,9��U���C�1BR`�'��o\�x@��(˵e!?eM���J%-gk 0�dX���.&?��8`�����f��m}He�>j$!�<ov�������Y[��%'�Qq�)�VW�������ȅ���L�՝幅�Bw�ȱ6gE8K�p�!�5�5&�;�NѶ�*	JY�10��o��U�U�y�	������.�2��aH���ʮ�`��g.f� ��ܭ��.N�0��:��B:b�쀡�ޅ��p��IE��j�/M�Ry�&JJsJ�DR�g�ZV��:����0s�*Y ���Y�C�m?m���3M�)p��ݠ56/�EF",:Դ�""�X�	jg�S�t'C��7������Ô���ŕ�S�v]	��o��H�[S�eXPV�K8~I�&۹��ؒ�,3k_�K�q��!�P��~�pq���,��g��#&�3�0^�c �}'tz/��]�^�h\`��3��S\Vm[ܟ0�H��y��Tn�S���R�мb��7�6Md����K���l+:��~�,i��&�?�2�f�=�SQB@��z�O6}�X{o9(P��'����J��i/DQ���u�O+��u)&���$�3��B	U�p�q���V�m������ׁ	� M=u�GC>�ѝ�r�yʻ��˂^�^��CW{�>���N:��[T[j���;�4-�mN�4�^���FlR����������"�k����6��ϭAs���9ſ"����B!zv]�����ƴG���oS'�ٔ�`L�7!�\��'�(��?��':9��_M���.v$�a��IK	�zK%����F4!�(���v$1��&�D%�_�Y�3��٨#�c�n���sU��+�uP�j�I�>�s ���Z䗫���uf�N����	5g}�v?��V*��h`�B5�W�4��9��}�QYous�!�h�ɽ���W���ܣh6,��(���a���ց�@:;{��X��:��
g㫚 �OU+��ZSIzI=S�s}}>ܖA�U첤�L�.���X�ӗ[ɷ�q�-��H~���c��R�ۇ�+Kϟ��:���B/�<G��Q@�@aږ�fw�ƨ� h��R1U+�
>]��r����rU��Y�]Vu��� �U�GI.���\Oo޿
��PZ�p��#0l�]lXt��&CSu�`b�8����������,��O���[���x����X{�gҋ&6*��U���5��"�G�{*ag�r}�;�?"�^���:�ؼ66M��R�F1����ܡ&H��%��ہU�Ea/j�M�qǭ��\pD�3ޫ&�����Pʵ$�x!ޣ�|9)�dŎ��BJ�tM!xI�~p2Mh�v6A���䉀jV�vׯ����.�u�Uuh#t���
=�&�����w�w����6t�J�r��JrW�ql��ݓ�wt` �֑M�P+e��_�����o}�®�j�w�Y��}}�v�l:s
�X�Q�����*�-�ս-~xoIԺ����ܸN�"HD-�X�����&�eR�����a�-L�������5����AjjU3y}V��-�����ʥc$�#�՞3~�~c�R��.�-���5>.��j.+���?!FN��[��X-��~�	�'q�e؛5L�`,��Y��T<гH��f1X�uӾ�jD�ð�Y>�#����e~�m)�AJ����(��f?�q�=	*ѳ�atVD�aV�9�z8ǋ�o-K|���؍e��pLd�5WB�[A�E
��âKD��� q8'��g!��l&0]�H$�:�+B]ʆ�υ��S���8�mr��Ϙ�pH�.��qx�� 5�{�!��r@LDn�\uAj� Tw�tu*٤�2J�!˵���}��g`_�C�c��׋��%}�>�WB>wt>�}dv�h�ݎ�V���֛#)-^��Qw��I���.9`>z&�3���� ]Zޅ	?}T�7f��eg�U�X���R� 8dN�(�Ƨ��&3��a�b��Ơ�<ݺo9d����iZ�Y^j��]��f�A��}����~ݝ�K��~�|��0������Hr����
`A:K�.�Hu�/�ZnՖ~L����vUE��hF,�M�?ރ�M>�&��N����ʡ_��e���W���%��l�@�ȵ�:��ύ�K&\����U��R:�9��.����`V��J[U�3�	1/{��|�pBTϽz�"4�d+���	�K�dp�(,����w��kD����OQ(0F�7|��^'���):5)�K��,*�˪�C�YF�	>G �H�&P�<֏��$;��q�Q��I����� ��.vE�Mo�|v._ۘh��z�@�����t|~����=�N���yW�*>��y�����ޙ>�g���ݓj�9��ڪ]��'1Ƭ�&�v�s���&Ɛ%nޠ��<5���OMs��O���X>�k�=�z:]CN�{z}9!kdM�Zl�V�94�w���Ny�O�?ݣ�co#Ur�;�_��5�G��8��������T�5�1��S)~�,8�f
�x�o��Pظ9Ƥ�����*��2��������,�>�YT��#=��H:n�� �ioE��>ݽ^��:����	�h�h��ڀ�V�US����h6�_�{��qV岛T��y,�\B?�["]�W{�^��@=O�o�A��7W}��(pVN�����q[��*���Ƕ1	�$|���2�|����R�8�O녿�n7�S��k�~H�C�/C|���������j&�8貼Z �;�\5���F��`d�r*�S(�Zg�)V��ײ$�O���.#��K�����L����\����;��U�$`�U�)�%�i����e�$����C��Zg���W_X���v9�� V=�<��U"|*#{r�M��͟k���;��F�\4��?�uR>�W���
��h�6�ɵYz������"1gg�ҋ�?J��*񕇳ﲾ���w����i���1�R@b���'��0�ҭ	�M2o�xvz����:��S.��(���X�#o�A�� t�_�L��ԾOt�E1̘+B�s��)�xK��2=.l%-9Eu���n�/;�P)��-/!��D$  5�g��"�/�QB�BaʊL���pŢy��2�C[�/^s��}���u���6��8����X�"3`Xt���ѽ8Wv�o3����W�M���c�	/DW;F�X��	`fB��o+I��rVP���ڮX�ERYp��j� �ށ�����	$��N��o����x/������>YBS��yX�w�� �|�E9����we*N��^�Zͳ��8�W��A�<�p�i�=B#������������ڃ`�����(S>�,%�1t�{�j2��C;�ï��0�|?%ע��aM������(�Aaw�M�f���	�/��?�_4�r�����+!$���o�֞��'(��@�;���\������c�1d�C�us0�/�r!��G.��w�':�=®OA�Ǖ]T��V/�V��^V35;��B��Z F.Ն����\:��jU!�'e�o�Fk+(܊�N��J�FE��Z�у��7z���z<x���H�O뷎(��[�H���'Th7Q�G����s3A_���6q�d,*�9��#7�<�%.�N5pZxh�g�o�8��%�2���0��l���~�(C�z�\�5� <j>Ylj��]������@�q�kxڙ�-hE*�$cݛA����5�4C�j�9{G��{f���$6`뚈��0���,M>��"��+�1�S_X��pϬ�ĭ���lɣ�hz_yj*w��N�mp
1�G/�p(9պ"y�RbPQgM�-�7Q�fF�R�,wzoyI�ٞ����:\`U���I��W�?�y1�Q��o4�,3�]?3��{���0P�F��w����oҎ��~Gq�5>�AjO��s޽��l����Z.�M�&���B�d��d��C��134���?�5�hy.�a��凞�{��a9�؝;4H��2P�t��~�������Co���XR� ��F��7Zz̤j�n�����| ["׶	�M&�zL ���1VZ�� ��]�����ۜ��K�!��Y�4��B;J<�~��0jپpG['n���We�1׾U���j�:z�O`�<�=]�vE�O�bw�W��7g�MM�jY���ڬWV��#2!�>R�W��7C�,�R��MK�F-��E��rՖb�Xн�Ff�r�
�^�h�M
l�H�Z�E��Qf~���8^�F�?�&W�U�#��.5�t\gj7��eে�'ֿn�h�L��9^:|8��-��ů��f�������+��ˆE����x�VD��TMm���@&��ݤ��w|��� O������+Y(�Pӛ?�&���X� ��UB��/�Ʈb�K��dY�`{N򘴅�B|��s����]n⩇ �!hOnn����MEТ۱W,)kR�B�/]]$�lN�.�:V�S������~_���y�i ��x�3N6���(��նV�����@�55!���趘�}-�z�		-/#>~�#�~�6sw�d��u�lR�#��ټ&v]Nk����A�����zj<��;q��@n?()��ĵ����+�����a▋���u�>�&� x��}����Z�(����d��A-d�E	��'��Zx�ᦦ�Q�!�X��s=��%�=A��BC2�B��D3�_����ki����*�I�$�E�rT_8@-�D�Z����9�3��,�D@"�IC�˳)�Y�h���wM��me�/3�������4�{��D���NYFG.�2��q�
�v�N&�����g)�=2���j��qW8U�h������5�?Ĭ*ZJ�RFLnj�Y0�I&�7}p�~��-��׻40BJ"�ǠzU]5�r��-��H��q]�v��D�=��eq�0l�#��(jQ�����s�D.�ܲ���E�禉�2�g�&+��x.�`�e�0��hr̛C�H��I��c�1�i�w[r�����=��uZ�%�|�����J�X�o|Y�Rw7h���<J/�U�f>Yz�W����O�r��,T;�����?�>#�>�h�F-X� ��>˾(��0��f`5D�3䉖�T񍫦omu����C�W>�5�5D�/�Ea�U���=ښ���08���Kߓ�:��S�,G�Ph��2�Uy��);�.��n� �k^����	rN���Cy���/�4Ѕ�êÓ-'WG�	B�́(�?�������	�\~��5 ����i�֨A���s����,��a�N�����!n8�Ip�a7���ϔ[�_�@!x�&�O�1v��B���}S��f�I&3�޿p��4� v�F�-�? \|�DJ�^=��wU�.6�=��	�5o�+�y�Jz6���	>��_������Ɇ����I���aa��	֚��e��44���j?/���>��!��qK�cٚ��	��!��o�)���h���~qͮ�0��M��q�riO�$��2�C���К忷���B=H*���B�����^)��	���^��C�¥�T���� \D�� ��Yb`��������W�|�=��l)��&<~�����W������CQ]��3o�wh2�,��X2Q>�y��]��c�S^b�� ���/9����(�0��F��m��>�CQd�x� ��*`ܶN���yT)~`�jg��$;� ,�(%�V\����9=A��챴� �eq��X����H�R���
��7�u9�[`@L������G9hK^s�-Jw��X���:ɴ�Ⓔ��{���޷<kD�1f�&�]WΒ��Z��]ЋA"1M� ���\!�1��?q�ݳ�*����h//F�
���7?	m��D����\h+�Sq�WG͊F�W/��õ>��\�����*�������kk�\�6�%�+�G�CK>�:I���o���T��-gY��*��b?;��8�T&�xg3�h�c��q�б�3�>х<������n���2h��\7'��O;[��4�};�ymk{�`��9ONzK����-Ȋ���W%�Y�^g��&�M�^�����r-5ߔy��y(����>��F���!b88J���&���Q1���1������]�ۺ���mIq05�7��d���wt�?d?"|�@�^x�]k�l)�rw�<j�t�E|�e+���$��	�8xʀ�dwa�^i�0�gX5����hą�;�!r�S���.]`��(�K�����'�T��y��r�H�������#�����}�|ܣg�`�m"��X	 ���H܊F$��P�}���Ó�*P���w�g��Y�����Pv/9T5��v�oޘq#�t�-�i:�I��P���r������4�2���EB�{vj���332Y&��.�@�D.F%����)����AoU<뮉�CO[�+����
����9JJ�?�Z*��n;��Z!v<3��k-�o>��|�����l$./��.�A/�:�6c�8�����:Fl��R����p/�������:0�I{�`�ʿ	�?��9��F��W�i?k�[��xYG�$N�ݺٕ���PsBI)\w�Ϧ�U���+3i�iXj�@.+��6�%�MZ���vT�^�X�Y���}��m8G�I�(���)4{�5Ç?!Ԋ��coq�k�R)���Q�x.2;���b��?����v����c6��B�&@���U��tBq���}ʇ���^��s�+�ل��:�x��N���:CƓ#d� ���F5G�k`�)`�#W\�IV0�%3��v���]P��NՑ�]J�LHy���&*�-�;`��~�w��~��-04o��60��
c�-&�7��"�I���|9NrG�~�KH�
�V�[�uQi)(�sJ��q ٙ�Ɍ� ck�"�� �Cn��Z)�Zv�|���lJ��p@�ݒ��밡���:~���� �lo-��%�k$RS���_��f�����G��j`���k�ץ�Ɛ��>=�l�&��%�ٳ������.k� �����e�L���i��j���t��S�*�yg���	�<��Q��S�@~1�ͪ�Q�;^��Q�NO��\!,7e<t����'���� v=�_�2N���K�YU�o�|���5�Z�>F�E�X���`��� e��q�C�(�=CÛ�v������rRC�[9��^��g�aʺ�9B��eT�r��<����r窯��P.��Ɗ�گK`�OD������.Z4\�5���[Z��u_q��5ӫ����o'b�d*�3n+��6l{���O��$B������w���M���_�y�owK��)�0�2Gý����oү�%!K�v�F��U�/��E�횶�ѡ�IMә��ʥ��!B�Z�:C&���H��ʀP�ZN��.Vx/�V	�XRY 3t�Z�� ��D���ה;�aO�Q���R�)M�
	V�y��▷�t_�c��9/,&s6����}`l��R���M\�(Wgd��#ExS4
��o�R�M�.H�/��ˆ�R��>�?I���z��#yeD�7��A9ǠC#j򂬣�̩����'���D�������$�G�!���bH�y����|��k��h��M�k�E��K��A�%��'������8g(S����cH
��:K\��G*��ȑ5n� *X4� �<#m�ShA�+ot���K2��1�0H[6P@�/B�`���_�8 ��/ږ�KF�>�� __�k>^s�&�K%��z�r��}���Y+|;�q��>���1�E�<Ӡ
@$�P���>8������h�@�d�_��թ�ӡ(G�a`���k_�M�l�66'trDPwa�������喖����Q�7A�,�����\�aV Ya-��1�$ZH�e���L�^��}p�`L����D�ɖg�2DC&�.���k*�t����T�
�aP��Xa=l��4�ɡ�����������]��J�^e �a��I6� ��8�s�O�v��p�g�J��t1���J�hd�̶���Ew�y����
x{�my�F�3ty�"��؛�7���]�b�q����P�20���ѥ��k]ܯav#�v����'c���+��b��A���W�5J�[�9&86����F�`y�Q�n���ʫ�@�<+���a)k�Y��ʲ�a�����4�QK�l��3m� ��F�o�]�38F1���>!�&��	�d۠���g↯�����堖(���"��F��ۧ���Y��H�z\�QKf����Q'�
vt��6)'��y�������O�a�g�Sݵ�;2D��åM�y���l8�~����7��uÁi�E��/n'챳�� ��������t�f*�|G%��N0���:������6�\O�-�@0�����<wћb��}�G�
��c5�̍K�I�������C��"���3��x1(��
3x�[J��s�ۘ�Wg�0��dl,sY0tm���,˄>�����K�����VY�+�+���q6u�2�KMgEvz�on���~@����$P��,r�P�j�(J g6�����j�4��f��1�&8`���p��gd(5�܊����nv��j��`�u�~��MS?�xÙU�)��",4�kM�e���V|��m��u��ż+��x�<է��q�C�<�X<!4��.;n G��'�a_K�n%��A_�W�����j!���2L�c�$��* [��xۜu�,�&A�V���r�d�D�і�x���M�s�r�/w�G�� �5��@|׹�����A�л�9�D��F��ov�