��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"��Ia�W���n*���x	�`�|����m��"m}��S���-f��t<G1���e���P\TS�V}y��HHC2è�k?@z2���b��W�����Pb#�<�@֭����s���yyٽ�vv����;)��6� z�J��a��W�a��"ʡ�" G�a:���>H~>��d�~�mU���>�	�_��g.*�H�Q˕��WK��B�A�O�����I����Ì
RW� ƍ���PeZ�\����}���j���0A�(�$z��S�0	�čP��7f�?M�!����ֶ���';��"|!^��⹊	���ttɺZV�Ӽ���"3։�E���K�FWi�H�J�d�Og��f��l�m�]^���й�/ ~�v��E����"����}��j9u�]X"¢��H@Ȕ���ځa����RolN���Kރ0��;��q���߽�<ʜ!>=���>�Gm=�*����@Z!����d[�}�1�M�4W�٘u���6;w�ض��s�%�dyj��m��\��h ,�K���H>]��[��Cd�5ơK�����B�t� �;�~�����Of�w �J*�g�tR�i��NV>k�m/#/�F#������$��Uߣ���_5�1��c�pl�HM���/�;���zb�4��:�<����Ī��mG�%��8��\$0 =@��� 5������)C�3�+��6 (0ѳ�T���$	O�m�ߌD\��}�J��Ml��|qϴ��%��_To|�5)p�t^��q@w;y#[I	��𭮠��Y}�Q3a���@&�~�,�p���x�8�S�����}�|��r���dL&b#�J2D��}��k.E�':����5xHER���]cϊQȜu����`����/�~��ת�7g���o�9o6H�e�D����g'�^Ű�
���I���64�0����o0y�1�����x~���������Gj1�9�/�l�8�^!��
w��'&�øIEv�lC���>��LZS�ru�4�v���m���s1�p>�N6`r�DT���Ae�����>'X������H����*� lB+�/J*D������?Et��;r��E��#">��2y�Dbq�{�wk;{đ�Fc(���v��4�.�/�N�pFz�ުq�%ep\�$#:1�W�oh-�y�
���~KO"�q���1��)%�H��ܵ�0�2I�^9#[{
Z��?	���,yL�����% ,Έ=����i�iq��H���C>��dr���ʟ���`�?�D��3�i=�<͛Sz��]LMU�Q�w�4����0@��{������p���%� ��ҊPIۛ�D��ۊyL	;ʵ���thb��kei�+)|���8E�
�q�|�^���g%:��������ߚ�����j0�-��'A��	�����q�>��8$�&��sk_h%���a[XRhs�L��x/Y8}�j疪�[5��9�gկ*���OG���y�w����4�-T0)[/"����^m[T>�H�C�5<�@dň;��hMx�Wv��