��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�Y֢�08)�	�SX����J��;|����EhI�Y/feLv����w�Zޭ��Ɣsk�sxG��?Na���<��᪜�ȺB	�fb"���:>ۋ�sm���y���ESԑ�qi��˱=����֚�D޲��e�r�P�$U]޴���{��-�S�/PQ�h�cXmj�x�@�k��3�2�1tx?y��1,pS'?ho/@^}��əG=�F���5�/�Ø�0'�Z��KD�A��``K�c���9�\�LKK���͡GTg8�y��-Y~��M݃� `��[l��*w�(C���ޱvj�ST��5�&{�N��gwr���7��\�^3if�!�k�3��!^�&g�HY��}⣓ae�Ժ�d}X�LF�i`|�T߳!�#�S��n���cUdh!��W� ԓ5�T].���zy��sC�� ��Ay��|��:ܐ�^W�#��^	CD^^������}4u�i��z�PX�y �^/����#)'��E������Y�Jۭ@�� �	��C�F� ��`s���N�5/�@��3�jN5��)��[R#��J���	�V8yUy��1U)�m%e
��߿c|���]A[ƛ�j�"ɺ���=�"�-��
�*B�2z�{�g��@V���4Zl�>M�Ukt��n|��3�X����*�y�F����&��|��2���+
��|t ~����&k�����U/���--}1�f:9u����N��Pnl�u���N}�]kg�h�Þ����)��Xr5y�o,%$���m�_?���=`�6R/�AX$��m�[k�]?r��$U�Ljo1��ܬ��Y���ެ18̄���K2��5Jj'�5�X\PnI�(��L���dw��oHds�4�V�=R��pd�2��[H�qa;N=p~?J@�"�����[XW��D/�#���.3K�YZ�S�>֣-f7�/G��s��<����YMYО�S�l�I�P�{b�1%���$�1�}�JAjE�Ea&}ð"�ܔ �ur���Q�2O��E]��� mCI�{�U����q�%"ʜ���_*���Ie��_7��h�1��K��v�f_[�H�ތ�r��$WT\��ˣ��f|oZ�F{��������:�����cw/]_�o���\�cg�:��of����h̰Ԫ�w*(�,�GUDwRs����/�����8�$x�2�zw]s�����} DE�8�-Q�$ ���_%{U�O�`� ��}�*c]Bp���9'd���	�}u�.
{(�������mĂb���s�@}����/OέYX����.pmEw{����m-�MpDm:���f ���2�VH�1�����A�, �G@��M%�Hf�l��6}>k����3?����6!L���e�H/`>���F�U*hx3������TіguG�|��j�y7Gâ���6����1�� 73BP&�`#�ݧ@;2~�Oi�d����ڝ�R�q�c���E��taRs]>�����������0�
}���Q�4SG��	?���Jb���B�����Bh�����r�"h�U�"~��9m�/@��^7J׆0xC�c��a*v� 1���Ľ�,P�a[:�n>���rvi��`p���܍r�M�9Z�+�g�f{��:Ԛ�vtb�˥7[��%��K7�Aղ�sHԐL?Qq�H�/�M�P pѷ�&�WW�q��
�X*8=�KdzxZEJR\Vg��3L����W:@��c\=?��B�@m� S^`�%�9Q�A�b]��4fW��B�_�P�$�LX���K V���m��{��kqC���
��~~\-v%��x�+v)i&$��~GT��h�ݡ͠�E�j}`n�����+~_�j��
,�5���}�25���/W�R%���Ll�@Faa���0��6_a;>u�iW�&�I#��ria��{ Blߜ oX��S���p����n����
\�������>LB���(K�^)��� &ݍ�-f?��퀒g�ǘ�c,瞡1�dK[@�4��4�ϓ�w��'��Ⱥ'v#!���f��XY1t]l��@�Ԝ,�c$���f��z���%b��������s7J����:����|�h�^]�tu+n\�D�k�Z��<3���}�g}�!w�	��O>��G�����Z�j2ӵ=^N��;�4����N�m|�$�j���I���}_�|X��?	^��7U��f��[?�ј���$���x��P�K���n���y��d�N�ܸ\�^��Uٻ�A{j@%騾'o�y������e2��Oe��Ը�
�-=�g3��e���N3��-�.s������Yp5����zhSW�: �p۫��%6�����_qr�&�:��e���|5�x +/�soۂ�DJ�������� ��),��S�Յ��r�Q0^�
>n�ݩEGɋ�HLxn��l_�����?�홵�F��f�H�"O���S1�xf���x��羹/���E��/5v�T#w���婩�B\�����|�gf�߀V�ע�T\s׃	6�o���ᤧ)!Ǐ��w5G�R$<�m󕊍h��w�Ѝ,A-�yee�'F�G���`*{G^#��L����8��Oѽc�?�j�5��R��X���6��<��"LU���JiE�H�ͣ�e����bϓ/�.���M�1X?��M���$�-�4�S`����@Y�llI�XЋ�*��&���,$���E%���!؃��8Xj��R*�a�ly,«c?����.x_�k�\���yb1�h�݌֓���"2�C��G���J5�~ڴ�{����Ć�-�J�. c��	�]��7ވ1S̓��]��G,�W�/�1� ��<�ry�o��b�:D�qF����SF�w�71>l�o4�Z�Sn9�wg��+�Э��5WG�w��O`�,��c�X�;Xl���0u��N�eR�ZY���Q��f��-V��aG�$`���G��T%2>��}Otb���u3�%��w���Qs�x�oQ��z�R�2�ݔRY�)�j�ʹ5�����z�m6;>,Յ��-s���Nv�2�zY8��Q�L4[��/~f�JPͲ��B��`�mˡ��5�;��5b��GM
���ڍ���b�'?A�.��<��+Qh��ه?�r�'��R|ZG`�����r�Z��e�л.:�V��&�t�cÑ��p���:M�F��:~��8{��i �/���#m5Θ+x���q7��S0V-<����FNG��h��=����YM�T�����?:v��j��>�"���j��x�ñ�l~��\������]����l+��Q�3IQ�o����RО���h��v,qR�Ҳ�?P=��*�NM�x��j�ފ�*F^��lXM��/<.����S�&�Y��p��=3�����s�ہȣBj��I��'p�!^U ��9+)Bl7�G���ޛ�ϝ}sc�ǹN>ra��ݢ@�D������l;.cJ���c%>����Q�aRT�^͋|�?�Z�z
���{���B)8C!�5��	S�/���$$:H���X8L�w�nQǥ����E�������J�+�$�̌A�\o��&�����]H~����],��4&|C����\��P�p�YI޽�" g8�368�U]�C;r��j6�������^��
(�/�r�T�62�Q#0��`��P)����������\�J��(�A�a�Yj�i9k��u٘���B�ֱ��揘�V��N�)�/<��wt�"騌tLH�X�x	u�$��y^k#Ή��_����kи�u&'ACD�:$z���Y������N.h����E���5��A b�����=k}���K�VBJ�a��/�諄]d��M[���t
܄fT�)^��)S��{���6�a)��ɲk���	&W��Y6�B��� b/]��TCQ>�"��,"�zI���Y5�9��NP,FF��2����넠�4�]�M��e�R����k2�TA��E�1�7ֵӧp;���̟�ᢌ�]�,L���jw[�|2� �������@?{�3���[�g���]ξBNw������õ�	=��}xJ}�ڎ]�2h��)���)��@sjp~�����כt��^.�h��	֛xu�C4����*5g���UI��e��df�a�m$5�?�e����2�:@�GS���!����l(+T;�t�n"��V�r�����#f����2N�'� ���fA[*��v��k�a v.��fEc��ېe@B�4��OLaWV���M>|�e��=��	�������.�""[|P��`���g�[i2�umqYϊ���Dt4��V���3����'Mf��t4�-g��É܌n���t
ׇ̩��`"�FfA�������Q!'`���l[P�u���3�y�v�^w�M�aԩC_�����kO�U[����/�\A�\ʛ/�:
t�����e���f�|A>Q~ ���7&�wǕ��r�k\�=�K���:]��Z܋
�v�i3�ͥm�FcA������ZR��+�7���4�2�)��Q�#(��]~)���_Q@�nד7�i@C<����kh���i[��,�b a�>��E�	l�hy}��&.}H1K4��O��/�Fcy*s�Xׂ۔.�{����?�,�;��Ǖ��s����CQ�=�&U��՞�@F�ǆWF�]˨���,�,ȝ�iJ"R�R���/�B�jM
����l*,q���1)�B#)\��7/֊��k��#eb���G����&��}Ð���L[�����U���E�'��"R�]]�ޅ�~a7����5�t�`�,��J
��LX��Xt�������L���^#g��.�U�g| ����KU��b���Ծ��F8(�ܤA�@b-'�Q[�FV&��A(PqZ �t��)Cۿ�)l�w����`���*W ���ߧ5&tb�g@�Oe��'ɖ����B��ڰ
���+�G���^ᴥ���
��)'cة�*q�aE���}��p�X�6��.(%�ʍ��m�����zdC��Ɲ����1+]��/W�'y��:�o�t4E��L���p�����RI�d��=R�3��%����e<�W
8@o��R�rtD� ��8ÈGj)#�OE<�]���'oy�K���Λ�n��X����3x���sp%=