��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�/�CZ�0 �^r��s��<��v�Ba�ҧ'@����:@���^�q��Wy�v���e:���v;���bL����ȫ�Of�3a!Ӈ(���
M��&���b٬׷*��Q;�bMl��Q��y=i
�;�������VQ�=��-͐���s	˩\h0��"�mV���3}��Ih m�^IE6��a�<~���MZ�$�{�p��K����c׽��]|q�f���t�������X�)���j#�'�F7�=��L�8|������g����G+ی��@��C/�ќf�!WuZ�x�L1�.�v�s���|�s���΁���R�(��>���,�t/d)$�c��ڸ����,�
��Mֹ�y~K�10�H�嚓��+
�'*��7�]�J��BO�-��#R\������,=�^�
+��?��2�C
��` jՂS�	���v��8n�Cȩyҕ��1=P���t[���v����@v�K&:~��{�v�GY����O�� ��EÂ���s�53�W|�t�^Q�3@i8?��jn1g1�$��Wo��Ԭu�4����+�Rf�}\؝��z�ۍ����L�R���(�V"·Df�Lʖƕ�}��6�	;̠�s�����;��٠�<�x����2�@6��]�/n���\o�������JqVϼ�}�}���잰�� ��"$�"`M��Dg��^u���<}3�B\USR"1���5�;R���v��4�r-�\� fX%Hj�A����f\����l)ֽ�2;��2Z�y9ĩgg�bl��:-q��Q��`?v�W�Y�.s��鲟=�Ʊ��W��6[��{��'%��q+~��`����q��e%�IlO.�1�?/�H�Jni�D.G��9�K_�Т;�3fyZK "�xJ>A�5�)�BUR��e���?�i1A�𮆑� �f���`�˰��$jU����9����ϴ�a�k�-U%ϵ�v*A]�~��]E?7�b)�⡑�F��FJ�`�|�~C0i�!U����GO�@I������ ~�ʯ�ڮ�GE�@���p�.��FR��%w��=�B�U/oZg�i[�g���P1�� �J��"�4�V_8I$yĮD;�����v�����H�S�u���hc��dFҘa�7Q���*5-��3aQ`�- �.�١zǓ�X>{���W�W�o"D�K]Y)l��6�5�'y�i3"�H]��ƹ�� 1���#`O^��3D���m�o�@�႞�
C�"vʏt�/��
��C�tl�/�ܤ�{�Ŋe�*������nќi����7 �?���הkr�k4Y��LOթ6|�П�Y�:@�VR|��:��&6�
����X�������`������kmO�p�������~K��d���t�&
�1���ˑ	h����A�"��)p��c��lʟ��U��Œ{ͼ*�gZ��[�9�w��B�U��3�=!�P�gё���>�[�1x�wu�=",�aBc,cP*�B����V�-*���bk���FG2&�?���i�)�!_�^W�.�Ey�����Cs?AӚ�Af��[[�çxs��*̱J|���x�Ew�އ��|]�H�&�*Y¡zX���������:PK�&d�e8�z���W�=srY�bȝ<����t&9)H};s�H� ����-��X<��Y�q��?�������ig ��RD��H�ӣ4�]�X-.�|�,b:�=q�@����řK��XPj���\�^�s?"%B�n��!��:�,�¨�!T*���AH�)3h(�ɚ׺B�w.�n��ᡐ]�D+�k��X�
�څ�"�W�/u���Ì�oM�oA3��U����%ς���+���VB��Q��tU%�޴�(=�;$�[����E��6|�ex/\���<���ȭ����"�ڎ@��9ec,����-�'M���f�M<�e�	�t�I��O@L���:�6���:ڒ���==�}T�>�73�\N}Q\�?yjɨ�ғ5&������s�	��蛵�X�2�;�$�wz(�4<{����� 1i5N�;� �x��^d����tq��D*/�{p e�	\��Ɖ �s�Ce$S���kz���ٰ���B��ma�ٖ�˵����&���Ӎ%n�,�~{�v�Cg	��g,�?�b*xrI�6>͉,=�*���:��~kt �G��|qIDuL(+8�oH�������/
UY6���~��j���k��I*C]�C���U�b}�.,m{�G{�#Yϳ$�������&ᬎ(g�W�=IH�1ߤ�����w�h�����j*�^�Y�2�yi;~ّ
��/�$���c@O�vFf����!8�s'��uM;�hSe�'R�o��^�!һ�4��ɊYK����^#�Bj��<���Z��`���x�"n�r)�HTU'Vʞ>D˔��F�w��K�N����C�w6o�)K�<X{@"�NgN�PM�{�
%}���aL��8K1KvY���l=�b�Kh(�	��~�(Stl��S�ϯ{���*��	�ՙ��u��Ndjkr���Q�~�.S��[6�M�����(i���2�LE�,������l���KN�V��mwK鍢l��\>beL@]��+#�6�u8�J�z}W� EDoY��Ѕ�8q��9��ᛧ�ٻ&V��40�2n$A3�Ȱm�Um��k�7jyTl��u=F9�7b��T��ulŕ����oԠ��{1T��礢 ?z�m���j63���NҤ)~�a�)˼��i	�X��vS>83��5�iAN<2���±A�Y�,(�f�[6)aWD�S������Hq������>P���V�;T*Mϓ+dtP�A������ I�P�H�೘ѳʓL2�Z�v��m�ˊ�d���d��i�8�M.cĦ�T����֚��co`��p�(�c~u粒������2�8;��R��M3K�Jȫ�x��&�ʕr�Z)�[�~@(;��ln$���#N�8�7���߉�Wf��e^S�s-]���Bi%XnI�����j@�e��X�ɦ���HL������#Av�&�V[8��\G2��"�\�-�n�ܙ�����fþȫ��zҷN�j=
M��J��4�H��HbX��S٠o'����*��@>��a<@���t�H�����aH� 0u��UTۗjd�9��/������U�����fZs<�	��ŉ.�k�[�3�G��,])�����.�\���uW���|�s��s�g��&�l ��T|����:�=�5Q�t��
n�&h�V�]��'���SZ�i����p�:<P�8�.�4*,�!A��s��6�凴�(���FYm��2�}
A�w�
�|�Bx�s{ O��ڴ���fpOӃV�L���%ׇϫڌZR��