��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw���Q5��xj�ΐn*�b��ɖv�WArC�7-,p�:q��V� j��$M#h*���=^����0� l���'�J��l�^wf�_GdѠ2v����5�_ml��8]�D�F����~+��;�g&�jf+�2b����,�����e@�|��c��� Nh��� ��誏����Q�˕q2����@�l�����N���+!��?�>�-�C����"c.z�y/J<Ƀ�ٟ�"m�w�:�3��|*a���ckW��q��\Xr|�%�/��/O�2QƸ�պEW�q����-X�)�?'q�l��]�Q��W�@�kG��00M�gm)U�"�huO�����x'��\JZ��qfzuPx{<u��"ݛ*1b�-!	�*Nn#a�S���	�����ߢ<<�*͛�"t��OˆF�S���U��pv5��椁��!�B݂EqL�sg�!m��ۂ�f��"��QlG�}�6v�1*Zrv´Zs��|�rHq��3��YoJK1�f�#�I{:�T8�`�?+q���$C���넃T7�����ނ����Ecg�f�*��D�}�Ø�e����hlѹ�P��l_�Y/mc8�G��n%�;
��>�=���i�y�Z�?�N��0>F�f��0����h_���gP�;����^�EaA���ޟ-���9doXB<J��Rlv��!�ߖ�+��c�Fa6��ɃO���> ������zh$��sR�_�
&C��~I���2C�4�͞�"-�D/��O�����}���Һ3��P�v$V`j�����Ñ
@�U{]x��-�O���k󱓳����r�������7G�-����Z`1Z���������н���v��r�]$ۤnɑ�ŏ6�78��U7vm��R� ��.�gQ��WKN�@n��cf���M7?2�Iwo�LR���Ю�At��QE��Ȁm�ⓒ֚�Y�����j:���rb�
�0�!�n�,��d�0\���FJ�+�2(��C����fA����o��y^�G&䜬]�lc��0���>�8< L�������'���q%�VR4�W��0�����s"�@��q*�`/;�lp
;ȣ	D 6��Xf�?'���UB.Y���w�@�@� ��T
Ʌ򅹚����n��J��Tm�q�.���:����wN֜Y��S��[]�:�g4�V�ci�m+�F3�z�s�����J�9�)v/ڰ��C�T�^�Fʌ�.%?�7�8�kB�NX�B�T���6H[�SB�F%�� z	�"��t"���ϚD�;�f���7�&�Knt���唄�;�t���l�&�>/A���BE�&,���J)����R��b��ZFs�o;i,�s�-2��_�/)������X0oO�|<�S�4Md��w�fvQ}����+_w^=VF��0$����j����JB���yZ�y���Dm����M�%���̍w�ȃByJ8x�"	>dv�aL���Aη1�ȸD�@J�����?t��w��!��^��
E¢��y�"��t ]�����bb��GWw�?������� ܑ�"�T`+L��}'k0R�E뙀"|���AZA+��~g� ��W��D�oW�7.�呂�]���ZR��m�Y2�Ƽ�|GF�J-�4@�56��?�"3$�8vKx�I̚}>rv�f�ִ7%��܁Z��bm��*���;�xG��ӎ}9kh�T�^���L��ũk�a���
�a��ñ�O�ǜ�����_C�
�{r /궕b���9'Q�z[�m�F���Fjn-=H����h�IS��ҹ��WOW&�x�r>�| �c�)��=��Jr�A�/�e�-9:�<��>� ���6�<��Tp��u�M�TO�.����>�3��4�H���qO�SS�K8@p���鋨>h Y������[UIx�Κ7�EyH��1�+Z���r�R��׃A��aZ�w�"d���_��r4Qy�]��G��^��K���S�U%9j>0Ϻl���q���/S��G��8��.n�_.x"ػd��S7����:A�����hꪓ����`x���;Y$�u�7fF� ,�'҄WLB Mp$ZTWD!Gǁ�f�9�ҹ�������k\ơ��k	d�'�)��x��2?�In�d$v=�c�Ϝe�	7��E�e�_�t��L��a[�-i�e�A��*H"������l���H��J� �V�;��~��-�%78o]
�ͻ�#���x/��,�!S��l��zs%��Ơ���*�-�IJ!=�UW��O:�$fb��Kx~�	��p��Sη�g���Hl2C^�i-�LE�_�yw�uz�O���+�p��_������a��"�;�V�O�j)�:|�K?��M'-�gp�O�^����ѱP��wh%��C�C�Mɿ\�
�,G�ͺ��O�e�bC�:����@b�Y7��}+��u�#�C��duM���&����~���U�X��nEG�����ѽ�0W_O��wV��͗	H��\;��<[�����'��'t�a<Մ��Ks�*3�˾�(e�V�E+� h�m�C/ƼW��J7��HH8㲣ЀZk�/��R��țTP�luK}�uΰ�3��kv.��we�oø�潣غ"����&
4�-�t��p���X-V��7T�`���贍��D�zH�Ι��{��t�d]�3B&1Q��3̐S�WWM�㙅$�[�i+{��ޚ7����{�OF��A�B�-���f_�QlCR
�w�3qۻm�PȆ ��y���%��U�nG��~��K�'~]l2z��a�M9<�`JT�������y�Ox�AC����sa+Oʌn\MA��+�{G
[�}�zoӇ҈P>M�pǨ���?_�p� �L�5]p�#�g`4��e	g�Ж�z�(=X�h}D# 8�2��VJ���-wA1I�V�?��$(������j��|��mg�p.��}9�Bm�{W�J��M��j��c������':fR"��M=5�؂Wve�>7H�+�꨾���gSS�Xx5��������,�Me�Z3J�]I�"��a�lD�S˭9�럶�G?�ٸ>An�g[j��%y[�w��@�IZ5������H1͞�%�K=�&�:�e�$R�4��\�"�X�&td,�7cs�D�c"Y�o1פ�L��Ddw�)�[��)c��J�tP����� $.�J���I�����Ѩ�~�U� ;����~r Ȱ1�F�%-R5қ�,��Q�
���Gag吲\�det���������+Q�2�/HU��Y��fTI��3���WVf��u�2�z��zn�'����b.n���P�����I����t�Q�5.J��5', ��َ�қ�͹���m�2Y�ԃ����b�(]��ո�G<A0������+$��%���957�Q�6S��
�Y�!N����,fW!R����SP��s����͙������Cr3V?G�{_�2���ڑ��X��,`4���LUrj���K_��G�LEJ�õ�N�ߐ��A�/P���ݙ��|'C n/���F��6��}԰T���[xt�M�}� �rs#�-�x�&��.�kG����OX�����p�?8�lx�<��Ly��D�	�jߢ 
SA����m��W8<W�p������E~���2_
dC�7�DL\��m�Ň;��i�q�>g�P#�_����l��!�D��,d_M6���?v#I�8,v���f4%2��H���U9�dm�����^k��e��}g�ƌ`3Vk�ɂ1ؠ���
���7G?�����"�ᬗƄ��J[JV�`8�1?���m��۴9㽤�f�!d#�-0}4xI��6�� @4]�3�l��@f��	��v�|��FV���p�����ɵQ�e�|c�gc���7mxCb��������߃�{q�,����nShUF?�v�)參���m,�j��T�)���m^�st �Iq;����;-�$zS��&C_,��1~��vD��C���-4�I����%H`k�nZ��U���uXF'��"��	���hw�^��Yǭ�-ד�8�&��Ou�	L�o92�������K?|�2j�㸉���&�옢����h5�rеc�M���,�~/� �N"M���A�����{lVV���_�;�җ#{�9_q���D�m����Y�,����,~v�0n9o��bn�%�16��A��,��N�����al>�Jp܃JvvS?ݟ��S��������B.���Bjy&�^[��fx�	�h�N�6��%��Cfű��K@���7I�^x��kp#|��u�����t���1�I��{�,��
w���q<��\M%	݄�tX�	}��������
0�,����S���rK�t�,��ݹ6�|�˪�Wʏ��Ӈ��}��P6��.�P0�g�ܕ)]i�m��#�g���C!m@��>�\�������^�|�m�ή>��ŗ'�|��ޏԺ)���eS��Q��V�]Z��0r
o�q�;qo��vM^(,���;	ԛ�~�2��?��h�b��6$�p�@�'qaXQz{���ɲ�I#J-S��>��}[Q�z�k�9�쏻m�݄�+o|p��JE*��2��k�2\�w��:��~��>_�?ͭ?S��Y(+K����{x�A6"�_sP]L��mfQ�u�{,։):����Ⱥ6����A�����\�2��4)As�s��k����L�����HOC1�&]⌤ +Q��Ƞ�$p^�si_Y�j�NX�Q�=��0[ßS;OX>���ڽ%�8_��DG;Tug��X�<T��dnfUl��PW�T�,[)mˊϭ���x�
{ay+�������C��qFaZn�<ޣU�S3.8B�I8I���E��X@[�C{~b-��㌭���+�&��K#�ܤ�R�����),"�c}sNG��G�w⬆����<u���x>��g�~� �k��%f�����}���u���ߪ��4���0�[��W%�kw�m����w7Qfz����9}zJ�9:yȐ3їW�m5�-��c�c��o��;�m������}䌺���������e�[��>���,��g��{ݞ���f%��`yMg�k���q��e�Dk�Î>4͇�
�	ԆI��hUE��˽�Yߵ��S�Z~rP�r  ����88�Gz�)���
&��P�S�6��v�6p�)�"W�{/��a�SR��wm�ΒU-�r��y���L/�w���g�M=���G�gA��#���R����DYLq�|�Z�4�ۅFn��v !3�sytU�>
)EG�eb��S$���}X�\6��_�ߖӎM4�H�y
1	��7.EEN��(Ϸ<���~}�)�����b��4h#�����A&���"���u��ݗ[�y�Zu�H����5�_���9��G��"��JUf��S<(ǋ.,h?��ˆY�t�9}��JV�eF���F J^�h^2dE��o>�Q���B�Q(°N�py0xǪZ���>�����=}Vy��\�ǃX��'>=�=	y|V�ZRB�G?}-�|�j������h�c>�8���W��ƚ�lZ���N�M:p�;��9<�f-*Pw-�F� O�S(�����R G��@�d�fo��uE ��D��V��uI��8�*lsL3�w�nѢ)P��L��f&�
�	O�݉��m<�xD�bC����G���[ƕ���� E4��bVͲ���rQ�n)�}�2�d��C����f4����P	?��e���<�>��gl�F"�;?��b�q$[�{��0_�vJ��ρЁM\٦A� �.*$@f��w�(�l.'S&D�����2h��w�W���Q��Ƙ7����,�U;�ΰdb�\.���˂���l	=�e��V�P�$���*�,�θ}G'4撦��A���0V��s��>*(6G$�gD�y�G@�o�� b%�$ �lR.�gO~׍��n���>��8��W�1+�HX-��B�iYIƷ,<��!7�+��(Rk@��=�o��N8��i�S��啧����������2r���;$?�Q�m��w�I@����	�vhn��|�_�0չ�-�_�m�r�M��P��<���Y�s���"�L�P�p$��{\�Ӽ��F�<�C��X�{=��_�Ow�S

�f�d���E3���W�����qr��&��z@�غ�=v5+�J���~�QE_D���>��*wq&�#��~j>��>��r��JQ�����+�(��V4�#�H�lۆ�|��w�ہ��]�:�v�4�������*3@��^�t�^��-��}�b���.�׏@t�������Kv{��cb���ƀ��f��0��Zn�%S�5���N�K�b����o^-M~
$�$#�:V�w�+:^�hc�I�+�XPZ$;�>"����۵��,NWvT=-	#���#f69�|}��^۫�Y�"L=�������7K,���Uq�u��^'n���s�-lړ�Ǖ�<׭���F��a��G�k�HGq����Q���j���.�qy�q�6� ª|i"�-�y:�8�,�?���V��Q�(������p��C��H@��#�/�K	�C�����;U�_�{�ԅI�w�F#<;�垺	�?�T�A�c�BP����(w�A�7�oF�,Pz�Z��EC��L�B��aN��M���*?zD�#3[}ʀ4���ѣ'��Hd]��
%�J��!��
�r�w�;�U*U�,U1�3Z���p���?V��W#6���`#I?�
vY�n�6��_�Z��;M�0�$*����};U���|7�e�DBu�໶'�:�]��ʆ�[���-E9q���hew�}CZ��;�_�r�Y������3O^���T���������;y���M�A�1�Ų�^��{���ez#�Q�g9.������u�υ�9q��8"Q@u�,�΃����(�_��A	B�ys�yl2t&���jh�-���O0<����+��6p�0��KV��+�I,,�8���zUS�쮖�����[���$2N��YD�% ��̏z�2��|�FAC���ӓ�[��%㵸��,4Z�;� <�\@+iV�ڙX���v�5�_%�e�u*�T�9ٚ\JH�(��A�k23����r48[)��1A[>M��c�a"aƷ��A姢��_�g�Kb8B+e���Ѿ��9����=��=Ev�񽢎��o4{��[˾�m�R]�s*D?o�\��W��~���U��Z�Y�6������Js�9�Q���9���Lו��* ���Yan+�]i ��;W�'zz�ۆRm@��lۍ]�Tw�w�KS�ҿl��miSJ%<��c<�����������RTѳ(;�[?�c�x�?<�v+�D-uܱi��QM�O�&����o�8 �G�<��֭�����q㫗Im2{	/33�p�D��;��K|I�ؐ��a�����Xv{��������������f�odLH�Q�����]�y7?<�5��w5�4dT�h$��@�Ѐ�~�8{���|.�z~S�e� %dz�ơT��hI�hFV�ev��3䕤��ӡ�e���鯠 ?�u帲�4�y�����e@ڦ�������JYjA=/��\�g v,��`m�`��R�jZ�ק�AO3Y�R�4��k�#�A�����?��n�Q�OEvDQ����9��:�U��:l'��pXO��w�+�wɖ��a�98�Do^:U� Щn��y7�@K|i �ş�C�P%���I�H]3*d�Qؖ��8�j�� �ׄ���x��ܑ���<+��h��Wxi?GH�$?mb��PP�|--�5q����Ƒؚ�=��m����cM]X�N�?c����h2P�Y����j���?QBN�-b/��`���(�<�)g��Y,$Ud6��̹	n���f]m��n��J���`�������/R��l�M��)����
WQ��[��K��9@���9����)J�㞴r�ϣ���`ô:s[@O�.�3d{֢d��ǹ_�'�	 ��	�+���HT��������|*�T����D��x_}�Ĵ/bb��h��F^l�-񶊄�I���@vL�{cf��NH|���d�x~�'$BC�7���v��	���n%���
�l)�꿳^0K��T�A���<i���";?�g�J 0J%�=T�����Y>�Á�)I}^������J�D�-���4�^��;�W�I�!4x�oH) W��p�e*���j�,��YK�eYq��N��d�����FTT��3�ࡿ9{�_F&,8�d���s�i�ݞ��y �8&[��	ҙ����ͩ���'�������Y��p�Q�M���̓&�o� !U�-�̧�~O;h�3��+�$B� ��3Ǐ���@NYǚ��ؠ2��*�Ք��&� nyw|WRİ��u7��8?���Ƌ���+�F�n��l0Wn�w=W'�!'0��*�/z��̪zk���J�b}�Ҵ�a<��UpGi'~o��B�^�PXR
�Mv��ExF�S��0��U|��;�J�5��J�A�l�B{}����"��$��۲E�t�I�Z�4T��?��V:�hE��2J��4Jh�<��-t�rY��[�@����!��з۹�8皲����ay�U�e߃�M��(�@�*��5xS��{}Fv��U���U'B"ç�|e���S��k�*k�j�}BU�M�9���
��4>��W)�Q�=�N^v§�k�)z$7`��_Q��v�<������ғ7�e���A��Y�boY'�V^(�xP�%���Ɖ+E�lq�x;�~��K�6K��s�.n-e}�R�� �@��9����v8��;��������zu�����M�bT��pl�<�e��w�b����8ވ��h^�~�����]�� �Q�OQ5lo�}����)4\S�#���XM��Q��5�qG�C���:�&6��39�ŊeBw����$-��U,��sQ��E��0aV�U�;t�uQ���B���_��[t���)�HFqv�S�]"<�䞬;%<�)�c���봧3Թw�)��;5��"�|[�u>/��u���O�GumR������幎�`Q�\�%�c�Ŗ���
L��fH.a6>��,� E��9�)�s]2���n���yy���U��D��n�;����b���jE@l��-�j�x�k�h���}(4"��Xg�w�%3j@�q�J�KHY|��u3�.�Ŭ,�d�/0�~���M�^���y�������g��甝�ΤI���Dp\�*{p�Sp��ۄ�fq�ou��U���zb�\�ѻĥY���~_?~-�j �2c��>l������wC��C*uO��S��ATƕ����QדIb�)��x9�Uq ����8 ��.��~1'bX/Q=�^�)���B*� BYZ�⻞�:��6[uq`��0�f�
&�&`���;���޸xv`��Q�����ƿ1���y���^����x��j\�^V{|?���O�C����Ɩ�ME0�I�WJ��c簩�ʞ�*�c���ח^�Mq��0�:��N]�j˒Jt>����t��k_�A��Qh���6���%~����eeb�<�8��jჷ�_{��듅�R�t�s㵬2���9�-��^k��5r���lPaT�K���qc\%��Ng�^t�S8BCw�/@:�7��CZ���9.^�e'p�֋�^SO���L��E��Y1�	����H�����a�	�º}p�*�Q��Df!�$��@.�QY�x(HO|cOع�#���8�	�zE$(
lF�AZL�6��K���:�D7\
���(& �f�|(IƯ9�{s!o�*ԮW3�r jx��5a��s�x�zx����N&��CS�K^%X\R,I� ��\��������	&Q�E_�ھ��^��ߥ�S�\5����EP���ֽ��e�Ȥ���TFyU詅*lٵW����)�F�H��5�s1��E]��V%:��z?Rg�����|�ymp����9�r1�[�_�<���'�$�� 2�L���hk��d�����7[��YL^�����yI���.UݐF]�+,k!���r�~�M6��M �IsɅ;-��e4g-@9!��@����s�E�'�em�q8b2Չ`��ؗ.u*0�=L�<FQ���.��ϒ]Vqћ#a�g\�AJ�y��EV��aҥ�ܛ4�gڏ}�w�p�^���2^���N�w��$��C�^6%*�п^.��C���if��U}��ɂJ�v;6�վ'��,��uMa��1�{��U�����`��P�	.����0�R���Hld�F�B�b��Bqp���AD#>P� �ٲ�}��,��k���{����y��[6LR�h�Q(���ɇ��x�:m�{�I(s�o>7�a<��ᄤ_�w�2�N���y�6*6,�t�5����Q�.����PP5=^��+�xo�I�r�^��`AG��c��3ё%���)�9c�~��hPuN���*@}d�V�������_��W �1��U�|�N�
s���X�Z����>�-7��+t%6ZKT,6�	م����W��d,��g�^�����M�L��d���mD(%08��*o�T��?G�w�Q�X˱��8f�B�.��R8Ё�
a������߯.$l�sjc7��m��9|R~g���:k�d]������H�TxM�L������\�˝Y���/�k�ʄ�D�&��/��Y������4�Vp�i*rk�B"��-	4����|�/}B���P�zvm�nÒ�a��M�W��T�;�$o�K��}cH�so�E<�G���]���Qژ�Z�1��x�&�Y�&��~��Vk}�:9}f��|�fj��������m�a(x�2uG4��ڗ$3iic�����@�f�t� P�M
�>�Rۗ*�|�zپ����)\�CY��m�)�.�����r�Y��a����&�ڟ�����(�&f	,8�H�w�\<��4�~g��>�c��Þx��S���7#`�Ø�]'��
{��*�'e�%]i��:S����+����^�Ť�V �@ulAn�<+򑩷��������E�@���QI����˰�����K�s1P�q��`:�a�}W/�4��]{�&�tɰ� ����W�a��s�X���N�U�(g�����V� ^�tup�Տ��=r7*u9��R�' ��d��T�w8>?�[k�,Ɵ�r��{�5I�u�N�@BV	���f@?�R½!"��B�6b
O���9�,��{�q&GE������K��z��I�S�N�e�qx�I��
�'�P8 �4F�l�Qd�{�;{�fUw��}��¨0M���{�qNV6ڇ\�=[������y�{��07����ځ�@V��7�S�EQ�>񾵈].����F�{S}�I��ΐs�sF	���jvHf�^��P�ɸ`�<\�K<L�2��`��< ��1f� ��.�B��@ �B���D����<p�}nB���v���׮U��? ��O�3&vf��+��9�/x�ߗ:�0��ZF;VX��e�����(��^��l�M���ci.�ؑKI�]@��^��qT�J��uBr��oL��������=���[�*�u ���2�ya��7Mx (��[K���ֺ�D���
���+�!)G}�!�����f�in��{�N�jl[-z���V���Ĵ������z/H$.j^2���9���<�]�_���n��x��}�/����J
3WN6=���6h<� ���7��%q�o�n/�Y������HݎRQa�J��Ѻ#-�m����r����LD&T��G:��L�V���iK\�ƞu���eDx�Z���U��wEŶ9�;0���	�Q�@��X�|cZN~�9����I7�/��qt�T�G�6��Et&�Q:�z���{ѮbĖ,��ep9� `�.�h���D(H��k�N��&�7oc�b%��_U�aγ�:���?~�ߜ���K����)��unp�x���fɐ�Ẉu�xl�f�d*��6�"w� �����s^;���_d#����0#���܃�Du�� �J���@��S|�r]0tJ,�5�M#�J�"a�)&R[/җ�@�Q���y*�A�8*P�ӯ�mL6�1�Ocu�ڕ4�\�B�;S	("��)�u���Z���c�XՌ6�����7،�����Z�������g�B�_C��8��o<n��<� �1**�\#�y	N+ laM������}#.y>\�cm�"��4s�?Z������O�v�JR	��F� %�V��	��b�@N�������ku��k7�o��C�<�$+%U��6���:B���>x�p�b7
,:yվ<�N�UҴ����V%�>t�!Q��ц����j�e�:�������#B��9��31��:��ճ^K�;�L=y#8"��l��Y��;2��!^Mԑw2йU�����Y��n�뤝�ͺ/����{�\V��<��6I���)��\���ƛ����p�;�/(�lށ���2z�wí�^n޲#MW21�0<��;獥�Õ�-g���B��ʛ���HV��e��Z�Iː��1Mz�U�}J���`��'e�G�Ə��v��\�z���ݵS8�z��0_�>��t�X�뮼>�2�y�:1%4�T���R����g����c�]��؂m5}��RK���Q�!�t�<�%o�r?����IHb@�9~؀�����O�)!�����K�(�������BAh"(z���uS�Rh̽��#��N�><sw
��C��<��H���te� ��h���H��V��U>�G��a��$Z�o� $�F��nqG��t��2������0m�b�NY�4�??�xX3o3��}��hk\{qi��P^��;%*f��n�n����Le�[�8���s�/�PdX�Q��M�$��4w�)�ǀS$��y�C�0a??W�PbnI?Xn~=��<i��4���j˪�ݲ�(a�þP�~ca��IsҴ�&~�5	y`B[6QQς\�>E7�Fa��vŏ&�o�+��*i@0(���L���`+�;a�<^����W�5Զ�a�"�ˠ�J����*�TF��`�Gؗ���?ܒܪ�������KB,�����p+L^b���T��`�2+I*�E� �so�6x�W�O���!���c��BP2���䍉�2�+%�p$T:q�4��P'B��rl�w���_��^Z���=�c2މ��b	�1��R�9j*��h��X`|I"�{/G��kNP�#�⣇��Inaގv}6��$ ������6}i����ͤQ�s��K.CP�&KT��om�r.c�b���vz� �Z�j@)���0�<y�7O
2�x�9|�����v}��g+��b�ۘ�o�����v4�9	��,!��X�=转�bff�z��\
�	�?u�Mf��_�5�!UK�
�8�����B�x!��t�W�V[����4)�T/�A��&BP�mvND�5���*G����"�����Lׇ��t�~ˊ�����U���I#-^����(p��z��-�%b
�-��N$��l}��%'�\��@�;����%�g^��Uד5�0�,�t��Q*�[����V3F�1��b���J��t$�u0�-i6H�޶a5�����g��g�B�XA����/��8�fJ�˽A�w���|�[�'��M�iP!��akC��͸�`Fkk�7E��9㐟nm1֬�z�95���q�l���� ǭr��t�����#8+��?�?ak5a)	2�i՜�Y�P���V����ol�zs<]ј��7}ͯB�~�~���'e7�M�����_WTc�/��+D(�}�A�r���0o1�օ���g�2�� �&��!H�kE�Ұ��-@��؋���.��o��R���V#��9���ߓ;�#2SC��%��a�w���ѢڎA�+��L��J�}=�.V�xs���-]��"؅ЛxD���Azk�zJ�y�0tG�<~�:�k���*� ���<HE�~���e@wUUb&Ǜ�����Zr/�&D)�#γ����-�ZP��dn��զ����߂5�v�:sw�a@j5�ڛ�^�~�n��9gUc��-�b�#k�7����m���Xɫ�F�QB��:�2*lK0��n�xH��D�;V�JQ�m�A����w`i�yQ?�ƌBy�]b��Be�����=;�CQH�����'���=I(q�F1m�8��t{�/�:6������.٭�������<�=ql㒘N���~{�L��?�D�^ϯ�nVk������|MRMDG��y��v�䧂žG��͟�z)�||����zO��gr8&?�0�o=�U:_g��"�?�ªZ뿉�5ж������E�ǯ��PTjA�̫�'�����ʵ5�,�ф+Rx�N��QB��r%S>`�����E�����,~�3�ò�ng4��%��*�3X%@��S��e&8�&�q����r�g0$8
�,���X�_�kf�N#�4H�:�{z~[�k(���������@��>�k"����u�v</��&�.�K�=��&���l�͞����j�[$�t�b,��nQ��լ�GqI�b�܁Ld@��_�[5\p�� �wb�Ir%~�р�a�il�6�T��˼�(܍<�/��+�`Q� �Y��5�j>���<|��$cw��	Vu�zH|�.�N_�'��g�'>�X�d�G���a\y���ϕ��&�ǻ��\8�hfD�ZNnH��x�:�^�P %�<G��%����.j~��kO���5���ր�Ԟ��6 ���_Q�h�>�q11���h�>m��#���ߟ^3������Ż"B����H��e�͚:����Æ9�+T���s��ہ�4��K�щ�w������fAzMNw��ǃ�@%��A`¡�>�C�hz\�KS�4	�;����tħ�1ͣ�����g���_��+q��Á�IO����: �ɖ�μ|�=�m=�-x8��p�����oR��TSnwQ%G䨖-�W���c+D�@m3����>]Z�N�tM�
L0��L�t[GU��0x`�-&5�p=��n���*�[��Pɰ��gQ:��I�h1L�F��<<�^	�@Q�t�gT�:@Lj�jA������?*¿%[�X�(��+O(�����!��u #�o�g�=�VS��f�7ب�]R�E7e��Q�O�Wq�������
���h���.����&����4i6X��� DoGHm��Մ=.çu �o�F�GmY{).�:��1�ni����U*�%K_\�@C�b�T>q�i�g240�W��I��!�{����{{D*��-~�B�Yw��PҴS���� 
5��}�&m��V���7�6e�����ˡG|�3-l�[fw�&��{���հ��v�(�!����U?���5O�(�ۆ+Έ=$�k�@�`FH� 
K@K��C����̎�+�WEu�厘v�>�A���UaQ��j':�����g$L��x��5�k.D�g�>�����M�L��&p�������2�c���k|������p)��i��i2&5��g:(+Qi1��H�Z����f)Ե#���y�!j�-w0��@i����.�!l��4��SOq^ů�c�����L��PUX>���(�=z[~`�X�5���� !37%��.�����-v�1.�7މ�n�?�3��6�"9�N#�P@F�� ����}/&)u�Q@ML�MӃ�g|�Lp���տij �Ʉ������+�)�T@�+��V�ʷ�J����TV���E��;9|.__e���\�l��4�'�����P,е�Ar����u�����B1�Tb��M���j�U�V��$������q鋷3|9@�䡾bL��N���%zV{�-�����_u���o��C���%W���?W�W8��oB�ZB��pEC�Z�:=6w��D?z˽��9=����U����x���e��QĒ�[��٢�@ଽ4�(V{*�B�l��7|"]Ou�-R�v�K����Dۓ�J[��+�Vu�r�<��`;9\Ŋ�����&Ю���+60�ɣp��τ�C1�4W�ꎭ��� ���<��[*ro[Φ��y[DaGZ@L(�.T�/W�����u� �JJ�<���>�=�P������9�J�ɇ����p���T�k^�)����X��!ș�a������Х��� p�x�rb��ri���KY��>,ĸ�%Oꨊ|��� �*-a��{���L�u-����~���B��k�RIpc���	�:Xj��/���z�Z�5�T3��/��8��-��j�.�j>a��U5"��'��RV�'`����F_Ӿ�i�v��Uf��f/��(���D��8�6�����&xj{�%Vݑ|ʄΈxL����A�"Qup�6[FL�����$��!��< gG���==HpXP�4��Aܾ��?\�.i�r�嶇�Mwt.�`E���5�Y*JL37
W�V��4�"�ˀS (I���Ä[�!�GM��/X�A���m�q����2�l�͡�,Y������f�w"�:s�L�~Wk����@
�PڰX���� ���A젖��GBl���5]=���Gl��g㷨���3?K�D�1���px���v8�/�A`H}���"�s�.��҉�_P�K+�~ﱩK�St��*�	Z��{xaEn\�ZzzTuh�����T���z�G�X�X�TU1˦g��L��� �p���.�H��6'#��,*`jC:9�d���g����dL��!4&���3gȓ}m�ƕ~����fY`�4D��9r�m�ƦO":G��BQ��`����dxR?����G�ɂ O�������A�m%0s�}QƨF�����p�߮�=���r����L��I�t ��V1�xG���i�?T�����7���[=��[�i`�{I��'��,U|�z^ؘ�?!B"�#��{[e�ћ���'ʅHWȪ �w�u��DD#i&�d0ͭ?�y���|�,f�1��h�>�]'Y@���/o��)��;}�_P������+G�40�n��X,��f��[6��]�b���K4+S�XΤG"�҅��#���,��6n�"�4����!�H�$P
���VP ��z��>fcB/�H�ۂ(�і�$\ ��`�}A�|
h-u?�~�`Ș=\2��"�x^�a��w� �|x���H=U)/�+mK�V��ls��2��pu�S�ͻ^0j���4�-���*��,D�Ǭ��w��UhR����67+}�T	ͨ�*��.鮄3�OSS�?c����)�������_RU�FAFNym�� ���o���Yi/��P��t�"\�����Y>3��L9 MG�}1�lq�I%c���.�uҧ���e*6SE���bo\iUgR�r�vk���@���rl$xB(N����̫�B�@�oQ�1i��� ��3ͦ� ��i��a��7s8X#�E�[� d��+������SW1=�'�b���u�����s�>�f��<��wJ^O���<Sl��.��M�)"� �<:ɖ���g����e���{��f8mY�8���90���p� pP����Ȥ�;�6Ep�@Au��wNt�)����N'�����O�k�l7�z��Ɛ��Y��1�NU��{�mE��_Rg�Z���!�ng�]�3���T�A����9p@|}�=��E�	<I��k��y�;�(�����
*�z��t��%�[.���|J��0�)�]#^	W^F/Aw�(�ϛ$7����9w�}�7�|zf7Q�YS�G+@��XG%D9�n3u	�����-�0�y��?�.�4���w���U_������w�eY5,�	���K^]�H��~����%t��ӛ�����`�������{(���2��B��]�(�a�J�1mb����םQ��!��'16P��Pod3�\dg�cϑ�_��H��0�w=������Y���B��`�t����\m6]��8c�,�3q����Y-^Q����w�/j��nU�r"sECԔ�}}��=�<��������w$S��I������0���3�węG^�����c���7ŚM��T� KS��{���Ѽ��ZAkꮷ|�%H��	�ຖ������d���6*ه��Y �&\��X͙���G4��X���EA䛻o�dYˊ
`a���9����4$����rz�Te��b�1'ƻjlOfO�`k5�Gh� �X�Y�]A'�� .��:!яkCgq-i�c��>�W����y^��s}�x�����µ�������/��Oɥ^��?������g�&�E�ˤw'�0 ����Po]c�*9����1r԰Bu����)�jt�~{���y�bO=\���w{+?�-1�VH�F���*�}*�z�#���)�Tߎ�\~q��d	_l6 �SK���\^���J�����ط½O��p]w����8��!��B[��1@fB�*(�
e���_�6GX�k욢R��V����&GP2;Y�I�u����piBD{ł�9Q��v??i�W�4�����g���Εu���M�}f�n�Q;-��FilJ*c�M�Q�ׇ(��'��I_Ӄ���T ��V���̾0К�˭ʉ��J �  	DN��G�]D��>z%`DPj>�)a�_G���&�*iI�a������u��m�C,�)�w.c���r^_Q�B��"W��
h�r�*�B���!i� .��3<o�n�V�=YI�I��~��Q�Rk�_-�����%�:g�=�BGY�0��S)���S\����v�c�s�����B'�%���s�\�O�]�����,Z�	\��T]BNA���^1��j�6i���9�mRC5�1�!Up�y�v����r��7)��Xl�c`l�|;3��r���{�R�f����TO��1��Z���*k(β��֔Q�ҁ�h:8�+"�a���7�S�d���H�@)��%�r������$\k��*_e'ݣJ�oóQ�\X����8W�6�W�q�i�Y��C�	3�w�I�>�B��+ܙ���h҂Gp>Փ�V8T\���)z��?�bZ�jT�M��ַ�^��Ն�2����i9����z���>7�1���{(��v
�u(�L��%2��T�f[e%G��h����$r�槟(��]&?�y'�2M��� !O̳�lDz�;�k�`
Q��Y~b�[�ֱ�/�[��0��l $# .��	��~�4�6������ê�b��_��ν�fHM~ %��`�t,Pԯ���ʆ���G����]`{K�3���M�Be�f�]��.��8���Á0����z_�nD����)s���MΙ��n�"����ӯ9w
����+)�Nk�\�ʲ����nS�#D{`��t��8�H!���V�b?!͡]�
+L��B>�)��S��\,N� ܥ&���=y0��Z��[Q�w���2XB?�yY	W���P�K��Z�cw�S+�w��+��Pp��c����¤�B�����6e�X%����ɹmdQ��r�4v(����P+�:Ye:�`uC�`3TY���B.Ge�_Q}s#;k'�4MGk�=�.<2Q�,5}3m,^��Qa�۴��v�1�Y�}��T������t��ƻ��-B>�,R�nW^��J�x
����{����æ���n��ǉ;>Z/)������i��蒝���(�%�k&���/��v*%���q�~S����)`�̱�-E7)�/��+���!a���(�:�(�~!GW