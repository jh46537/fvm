��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	zON�0sǏ�7o�J~[�;�FLP�; �����~�+���ȗSXc���v����B-W��}��ڠ'�e���U�f���_G��De�K� k@� �� ����.`Z.�����F��Z�}=��}λ�>Sq��g��?�R�ӧ3Y�7r@�v��.8#�]���xvo$��ixㄾ�@�d��{" 5�@z��I�q:I�۠gy����b��W�,��c�luf$EꝢeq�l�A�z�X9@Û�<A��$Ѫ��%�@ߦ
Z�s9W[N�}Kb*9;�ې�����,l�Pw��A�E�52��Q��5��(�b=UC�x�z������:#�W��c\���GYY7��d ��a%?�l�=N�%�_�oE��sd6_�&��@���(�w�Zp�˻�D����B�qw� �4��N%�WM�Դ��З�C�=U~�����df����>��_�*�'��b��c�d�J�;)#���g+��*��}�c~ͦ5kz�ݽ{=�X��9&u��$p9�W,�xd�kc3��X�ӛ�fA*6�p[������`` BBX4s?s8����������i#�1��.Ok�D�rf��������j(P��[�*��ަm��N�ٱ|"�5�o��C/l4�����)�[�0Dk��"�M���+;f��$j����ޔ ׄ���3n���{�mH�rR-Fc?߯���j�|����BNf�Pc�fZ[�/\Tᐦ2�3�y�%�G8T�X�$�����cߚ��_�?�;t�� ƈh�Pv���!���r�y?�lպ= �<ڐ�.�K����h@m�/9�������r�PU0޳�=�8V���=N��#L��K�Y2�;����~��$^��+����dd���7>F���Fk3K��P͙����Ʋ$T�'ֶ�Dk�jhO/�bACB�?ˍ��JhVls�h��E�����=|��j���:�&����ϝ�{dj���ȧ���
3ŇB���3b	_���I�ub��Ƽ���p�Y����;�p9�Ǩ� ��L�F�晹?����*S�)O������'�6�l@LR�D+�n�ɲQ��Ra#��Y�������;�(������M+oCт��Fh�.��("���������&g��f�u�8%��ki����L{�$]��H �^�R�`��6ݫ�m��p����YDnP��F�~AMM���mZ���|�,��i��=�	�b�#�g(�B!������]h�cS����F�$|����ς�Q=�&{^�5�5��@r�����d</�Q(n�}H�]��μ�S�2.o�LeJ}6UP5��<)�1K�-�#��,�K�Bt;��5t��	���6x�A�^6t6c�#%�f%>���,$F�/{G�`tљ��w�:Ik�1��9��cuޝ�|71䉖쾫���{����qs	���CUMmǸʭ�4:����ꮷ��_���q�025�n���p93�3�Pa�� j���&��]�rޡ��������Ȍ�<����II5֊� %�BR�c5_kݐ�rb���!N�izةվ�~���]-,
Z�"4������8T�5 O�2D���a�A��'�+\�����}W�kA�+�J��ӿ�]���o����@�Q,����z2=�#^��i���.d!:M{�hX��8��LƏ��C�������g}}���������o�U�G������r�#�CM�Ug��H��$Y���9��Ȕ����~�1o�d��>kBS��N���Q�4y�x��C�檡����ؖ����U@Y�d0zE?^�1r�fm����O��Ցr�����lL�lܐ>bی ej͍�X<�å@y�z�J������b���Ʉ�^0���>+:��{`]���ש!+jt�*-�B�P����l�A�e��,�Xiq;�.Qԍض���#n��$��p�(��������jK��c�x(dx<�;���ÙLDc"8�nCHD%�O�|ZPw���
i�d}�7����Ɂ�wB��),���8�ږ[a��S�L��r���0yE(�R���Ň]X*6C�j�����Nd���ޭ\g�Q�HC�O��o&�����SG�,Q��	o����	��7UQF���~7�0�0�.]��C���}����.zR�J�1n�%��F���Nk���j��Jh#	�/�$vy��.?�l�`=��o�����&g�'ՖC���a�wC�[�~&d��J���x0���;�pfg*�;(G�X4ַ�Ԑ��jP�o�(�5��iT���W9��"�]���e�[�}�\��;��M�D����>,r]���`)"Uz��h��g]��{��Ar��8ʠ���64[Nދ�GA�< &>Nϻ���/+,�j��� ����B��s�g�M�O-A��Ğ�6�5%�Q��+6�� A��:G�`@�X�����'��ӯ�6P�Yi����&�Ĉ�C���_�olfD���:Pxv���z{��̲F��2<��=/P���(T��oG��0����p�d��x��M�*�:8>SJ��ԬL��u8D&�fA6�҈U̷0���$ě8JK�Myk����Zds���X�E/��<��W�*��j�c�n��P@��u���������֥�3����
L�]`�;���E��dQR6���`�$��~*�
L�~	���%�8������~�<:��5	�Ǣ��ux�Rb����
���,��oޗw�紱V���FJ2*B���Ud*��?�x�lL�6��Q+��N�E�ꭄr�K[��ouh��%�_�4Y�h=XC�̃&���5��g9oJyئ�vs��&'�5@�*�=>�<Uu�nA�����o�u�(.�a1�� `Y�.(�f}� :� �MD� �ˤ�k/�W��%y�W��J��k��~'��*H�������l��o.D��D�����H�#�t�Y�|����?I�]i�>��5�$R��>�l��K�KʸN,X)�=�=��:PK�V_��>�gHo{���uD� �׳v�jG��I���'M�yR&.+�1&���s坞+��)	�=�Ɖ/�?l�ԋ��}����ư�|FS�8h�'mYn��=�!(E�Yׅb��Ǆ�M܋a�W5c�.!,�T��_��6~X{��S;��� Е={&�}M���"������)�&Pϋͷ�.����f�!9R�U��pG%�u%v���Q�����&�f�$��}ª����K~~*��9��t|%��M`��)%M/W�e��^��1����Uh�s(�t�.3�nH��$�1����j��N��	2m�E�;�G$��N���`u��}m�����B�H<p��}S{�3�=�J��w��&M��^Y)$�x��y�Qҗ�����aG���c�U��e	\��Z`�6]�|K���-�}Ŧt�5B�e���`l/�Mk���j�Q�l#�*�e�e�[�z�g8G�h̚+S�&��o\��RŵV���&ǒ㹥B1�� ��^%�A%d�'q h`���l���ԗ:�����t��M�{��EW��
��;���2�]6�x ��%Umo����sR���N$�G����� @�﨔5��m�����B�����U`��.�j��c�m^g���)-��N�*Y�TÄ�2$ �3*]x%��Y���LAo���C�'�+�O�Q�L����9h0e�ܴ�|w|�ѯmѱ
�l ��H�̮��H�~�����c��tq��t�O'OO/|�-cD�m��8�^"��ңW�xE���]��;���,!� �O^�Qc�N�LTM;F/��0�-4��p����?�Lk~�xK�Au���D�M��s�R�:-��¡䵮�t�;����%��J$A�ރ$Mk�2�|�7/T�7�a �R-�s�R�#`X�Q�ٵ�ņFU
i&4:�j����^ޑW=��5��[�G�~�$�{�˟5�S}�	��)�'�`'����.��.z�`�2�7�����#�Y�+�*�T����Gl���N�������2�_���>�M����x�mah.��\���'��~Y��38ɿz 'W���}N��W$����U�-��1h���1�tI[��Z,a96�T'��P��j�t��2���N�UHL�kO�`�-K�������[P�μ=�f4��D�r��a88���5[T/B�8;�W�Oë���ك˺�l�.��|S��������͜+HU����(Ѱd���q��s�e����ʫk%�CP�}�P����l���\�Q�S�+hj�&�T��Wd�����aU^��E�X|)�c���������F9��ڻ���椳.B�y��N�wkG��2Mшx��-� 65�AQ�"6u�j|�ۖv�*�"C��e�����ֲ�A����eh��h�����!��-���_��\����z���mW�l��;�I����e�?g*~bң,~�Z�C���$�\L#�<��a>�fk(����/��`%���83��`�*��1Z}Q� ��U0�~~���Աz�"x+1�2���yX �4�7M�"��^"8�!�ӳ���E�OCx@�-��(�Ǘ�O:m�?e���Z����;�۷jr�TvJ)�;��V���n&`��Ȟt��\"���\�� ��_��7��fS�(�}�O�����d��[Uc�B��#w���.ܲ�	2�:Q������v��d��SԯL�^����'�D;>���w`��y�� ŷ
�슏� ���d	7$U Z�{D�%���r�],N�xޛ�;b��\�OW�_��H��k�MZ��2H(�*`*1|��fK�Ƹǒ}K�/dqh�2��z�[p׏Ŷ����Ց�m����op@;>	G�d֭�G�\���6v]�.j�����ݾ�z��93zV&K���pd<Z`k����	�~���b�h�f_���� �|2��~�ax��T(虇	��!Q~r]5[����q���/0�0�f�Y̷-G���{�"X.���"��n��#���#T�z�4��,u��J |6�Q���F������LW��'ݜ$>Qx�-yhr��'P�u�EF9�0�]hO���}ϣ��"�9=���N5���avDL�,�|��k��h���	�W�1W�����s�� �7���"�*EAm_YJ x��TQ� t��i�uR�����k���'6�t���%8�Q|��A0t΢����2Z�11�������U �G��2�~NP��r?c�w͵٥:\¢�`ߪ��߸���X��<z�?a�l}�_\���GE�`��_�ca�]�P6��+1U6)�ts+����'�]�"I���*��yHS�8G��t1��bM�e>=[@6=��z��ҟ`15�>4�/Ԁ�K��Af�2�ĂevG�d$G�t�	,�h���\$�?�f��G�u�5?Kq��ߣ���T��:��!v��*j����o� ���_�� �Z�!.V�2,ǌ[4GӆQ����k8�'B��)�c+�hh���՟�R��� ��bj��O�Zt���r�3�����E�r��,���*�e���y��-�e.�?n�R������$F	b�W�����Ėx��[������B)��w��"0BImf-	c�Љ�H�ն$����]1�E�:�92��6�iI,�A(C�*���)��"ث������%���+J1�=�iD.��� ���/U��ɝ���0��l ;Hč�2I�`M��~�� ���GҌ�Ǣ �0�(M�9�ZF_,Kޯ��,���\��ғЫD��<oɌ� 4j��lNIaN��������+e���)aAɥ2����Y,R~���o�^?d�I@y�=oն/���t!)�|�Y1pD�Me53�����o��n��2�����/f߄(���#P��w���{�q�8Vk�i�W�fHW��R��7w�gw�(w˸�1Į�����ku^0iX�ϐ�U���1�"@��[M��a��{��k[~p��H���i.�^����J����ӠZ<�ff&�qΧy������"�t7E3]�M��\��>L�j�c
Hlc*�� !j����Vre�)}��L��C��c��G[A�o�՟���%F�6�P��m��L�ށ���}��߇��_X���1s%�"l�'��ޤ[x�~o�|�8��:��o�~k�ң
L��D���m�3f�^+z}�ֈ�� Q}e>cn�+Xym<�(Uͥ����?f$!~NX������C��i�ƻ�$��t�7���j���=hò���[����
�_���(�KO	d�/gL|@�%x<F�x�����;��\q҈|�K��S��;�0�Ύp�p;��ɇ��`�4Pl��<XZp��"�j�p�~�3�>�r+�������`�Plk��n��lD+�7(]�������}�.�Bze�7�c��Z^i�|��@��Y�m`�)�>\�ٲ>0|5}��R�=����
�����[O�`q#�*�=��h�W���e�'g�t�sm��]8�FlJ|R��ΨJ�;�멟�v冋F�f���8������8���4�dy�E�\dN�XD=G֗��������3 n5
a�Б�����Y�p�\�i��޵���p��n�2�V{�^M~�!�V�H~3T�[��a4��D�^4��=�ʫ�_���x L�]�����9���@�z��c���A}��Qz�چ�*U�B���Ay[{U�����یu8�)�99s.߰ Pݐ«��FZSY��/X�#J��Λ��OB�!N�Y���b���4�T�>�I4�a��<���K�F�.-��`LQ�w�qe@�ZW�+2����X����8|͂=�1)�P�c���JhSR����QͰ��Lf���O�j �Kgά5������n�8����l�#���S�������쉽��:ir�%Ux��A��9 ���И��K�ZPs9�����׎ݐ��K<�Q�}�y-����.`�|E�֙�J���ޛ�B,Ϝ+��d\�(*X�b:hp���wK��E���
Q1(������J��'}����$�x��,��ӤkI���JZ�F�F�p��ҩ|H��@r�.�Y�x!zK���"Kh?��u�����q��H�s�z[XY��Wf`��e�!�;я{�N�W��p�����@<gvn�/��K���]��v8�$���_ݚ�~���fcn�"���y���`��]�`5kK���]܃&8&�3����� �u(�#Y�U��J�����s�_�)�d�rn��L�Y�@���Nٯ>��V囍f������Vj��=S�!7-����XeS��J�c����;�jG2���'�T�����nZ�"W �:���WiQ���NE�g��wV����x��SV:����o�YZ�Zu�Ϛ/�]��N���ñ���4/ӡ�ƣ ���f�m����<�*�RT�13�z��������1��qRݲ�0��g��~7�"��%?!i������m�5�OR�D���W4# �:�[~=���c���R�7���i�)�5Ug���fl���9�"^�{�j/��f�^?(�]0pC.��{������͍AnAX�4�0l��)��r��������-�Ł�0r&BWdk��o�t��.�6�ۋ��%9� z%,�5s��}E��w�ו4 .�"��HD�ef�����w���m��6<6j��O�ߩ,�c�Gp$�(Գ���h�*�&im�K� �8���𷹙Kޗ'+��1�D[kuSe�ebM=M�T��ɶB�Ӆ3�Ď��h�,F=��I~'R���CX�6�0��u���yl�5��#�t�8p�g �����ACxd<��]z�Z��zE;�S��{���o�ds!>���zu��=W��O�v#��@i�`���w�f�:sε<��Fd�D��S|H�Q�$�� ���8��һ�W�ݽ�"z6/�E}�*��qH"�KBD:-+t���"�e�kC�XNi��hXq���mVv2A����pA1�Ĝ��.$����d�p}L�?5��PV46��Ǫ�o����*���+��Tt��㞴���,�ױ\�y�߳_���yc�8�ޝ ������rsoG����~�!�m�s��&ݗ�elX����|p�z��x�:S�;<>�$��oK�T8����̰^�-��|J�Z�{�ཐ� �4߀�n�<Y��l� kbt��tM�V��� ��H�K�5^����+�-C�� 0q����8J�a�O�Q~K�"�>V�����[�o�
�(�'��w_< �Fb��0���^���Ks%*ff=Qm��q���	<W0�m5���Y��bǤ�R�lU�/aV|�t/|uV���N�N���|h�m'vh��,��U��	9�PJI�) ��g��pn�b�M�4�*�H�]��܈K������ߌℰ���>�R�X�w�[ʮb����P�	U�k�˦�A�1���c���Ȭ��o
��
�WK ��y�H^b*o�w��$ULJ3���U��f:�	S�I����{J�[�GH�	V�u��"`;�k>K��v}^��f��4���J���.������\�Frb�ZN�~�X���	����d��}D�V/&r����� ��[M>����
��	��b�d���1���ř�&Ԛp02�xUK�8~�WW<��.�R2�<0����u��̀��w���$���J@��S�7f�@�|�x���)1]�A�hf�ϟ��2�X뽉���b��4%~@�'x� �y,��ս�b@N.0����e��|7"�K��G��H� ,�ƥ35bi}⚽\�A��<kܤh��WV���f�j.#�ڄ:�u[��T`�N�<���kN�.��/ٚ�埕P3�Ƀ3�\~F�juկ^�^�L���}�!���`��,V��;I�}�P���E;��z�H��|��ܤ#�G$#:mQ�R���^��+]���Q^���a��q�:FQ�����D�Ky�{��K�t��`c]����j�q��w���
���HD�C�G�1��[P�����w�~$%(���ZV���N! i�6wX��x}@z�sw�0P�gr��yb��D���K��FϤ,�R�pŵ焛�괝 ��,������J�Ⱦ���yV���4���Ū�����7�QA9zs%�������p	Nh�MR���c�~��C�jTb&R�N����ŸH�xG�T~��Kv����b�o�a#��qԕgӭ3~g� �O�ȩf��X�)��N���
�z�V/ﻖ&e6��M�Y�u��Ԥ^���A=�Eg����qL�EN*��|��Y׬���Zc�C�����}	���_q�jY$��0`�eY��Qʳ��8�9����ũI@���z�o�V6�"����E�a��l��J�@��l��Lq��P�m�㟈Bmнz�5<�!%��� s�&V�}ѹ,�z�9����V����4��׵��u���F:��<QG9�/j�T[Tk�U��[l���:����N.tғ��L�uQ�up������w�>���V^�����U�f�k��0��]e�Ǆ�#�.�v/�j�.�4�L��O�v�����I�G���XoTZl���c~�|-.� P���L�&`��NK��ׇI�AW�> !Z��ãK��U��ˍ/�Kvu���go��r�.�7�z�
`L�7��iޗ+Ny@"<[o��M&��Ѕ�:�W�SK7��	���y��6�tj�c7ypN����ԁOࣛ�!E3jh4[��p�j��M���Nvy����q�r��3�0�u����!�%��˯�T��a9�~J��a;cq0�Y	x�)�K�m�c�
.�:Ej������|����Gh&NH�y�6�b�t1E"��{�$_oyZA��˙!�_Q��[�T��&��nƘQ�;�f+G71�r��(`)εJ3u�,�b���8�DCd�D�<�Gb�ү�ia!M䒵Bj>������%���D���a��� 60i���́}�Af�g��J��X�ed�-S'���r��o��}y��߾`\���;H��;��6r��z�c�w���U�+�ż���b��j�N��'ml�ڊ��{w��@X6~��e�]�G8Pʞ�"l|
4�g��VT'�n��EjB��8;3(ɾ�|��u�!������/��nVM,`���(M9��w�ю���iU�2/��:�K2�^k��F'�o��f�{-���V(P���]��M���ҙ�h�:+u~GOTE�c	�=�&�+*�U���T����I�%f�]%�a����^��L�Fnw�_;�@1=3�ls�^�g*cѳT����\E�z�.�T�ȥ��"�ʻ���Ѣut5�A/�d��s�\@��U3��]�=���r��gnyH..?�ط�2�t;�n��n�	��f��y^�����68��˾��#`[�h���6{�m�m�,�=@8�)w��)������&9�|-�T�Ń��X�mdL#k`�Bڜ���2�i�Bʹi|v	����.�+k�w�����L�U~D�������W����Ud��hy.���%U�|�D��C�������m_@o���#�'-����fF2���{��!$�O��Ϙ(��c�@�;���c�s{�����YEvg tEn�$�,�����)��ay�Z���b�עj3'0v�����s��m�a����!MD.b%'"����82��V�"A{�3�"��)���B�$��zF�@y��1lh	@�"��{_��A֣J|j5����B�$�@�����۔q�2�Q>�B����l����eC�9
:Hb}�gKMz��@[�:���(���vm�?�7SG��������x�0���䗜u��1"��1���0��I�P��,@�&}�������4���!�lR���y���	0�$"���$�K���N�NM�;�N��G�z����]_������L� �{�h�ohs%�:h�Sq`��8{��t��J���/#T�|P��|����ռ{"Xz��u��;	��_�;�˔�8$����_��b��%W��<��Dޔ����B�=�c�b�b��a��D����QE-��g��n�qc�
�\9�b�VǏ<i�w^b���rl?��4��┶x�A�������3o��$����j�O|���U�Zl����q��ؠ�)N�O����8�t�>�H��z,���028����;��<��$�ݳ�"���qcP=��*R�?ȲxZw<���X�x�w�4���Yˌ}�T^���l /����u��A��q�N@^Ҕ=5FS�k?C�H�P>7�r��������-y�$�2�.p�%~�*5Y��mC �X�Ɖ�@�#L��h��ɑ���XVбL�6Vt�>5����Q�l���ټ�K�W.��V�(�84��"m/�O��AO�=!q�DP�t!'��0|�Ն�94���`��͠&q��V�TY��X;����G�=uPNs�P����ɚ.2م�F�)ߐ� i����o��|�^�Z}�zM���9��lHF��pS
�dK�s 3�MT��}#���iN�c*�
�OP���I���ڣ�HfF��J��!_� ֽi]��K�RY��N�xp]KpX�]XW���"��e�HW���鰆&��v��ޗ޺L�OE8�)��L�M�`Ȧ�rN�yY[���C�Β�Y������Pf��`����T���Ȣ�0:��(U�y����`~,�l�&���bA :��Z*Ec1��/AN��h-@ǈc�����iΛ$��	3]�8W� ֢Dq�.��u{�xK�jmk-��)��� �#�m���W���>���T|�� �A+-��(K^a|��ɭ ���`�rG��/����u;�5~U�RJ��K?K������?�$���J��w��E��$|�]����b�r'GW\tL��i1�7V]�T~�ySL�F+�������
v̓�_��C����m�,��� ����W|W�Aq���n���.�[�|�_-db�Q�hP�Ъ���%���O�Y��l���}7�,b�$�^*?�R�S%����Ox6Ɠ8��D�(�Y��8m���X�E���ű*�s*1ka����MH)��f���I�����	z�N�
�����z��A'�忨��Lak��:}�R���C�"ۣ&q�`v��LԛA+s<d�6�Q�hx����	C�MP[,����ν��>������y��-B��{��<�ԍk�}Ё��m{���D��.w��I\g��`,���\����o���b��p�ŀ�g��D���g/���?t��7��R�g���`ʛ�'A���Dp�s��=�s��	3̣ѻrm�6�R�|����|6�]��:�t��� HL��$�v��hy
vB�)�?�V%�3�P�Qe�!xEOie�n����,."���?wH���gOrx��9���h=��n�r�0C~Y���D��E+�}�Ak��0���'�Q�"���_5����2�+aF^PEs$fK~�����5�P�`p�'F�p�E`��Y6\F7�����;�j<m�W�� ��Q��{c �@�ਙ�ؖ6#���(�у���5�Y{���{8`ݦ`���G���do��ueP����%}�ֿz���,��p���]�����ji���j��{mq��z���<�V�p�ml,B�(��@Jk� �-8���#�A$�)�т��2<�kM!#�&��e����~�s���1�a435&W�,9%�N�� ��E;*��b�5��"���5�n�q�)+3h/�C�6�����m��c��J�TL�����R����.U�N�X�p�8a߅l�2�6�P�E���a-Q�7�Ay:���K}J�Ы�_j�/�?�P�K�K}�&?fE �! w B��9-�4���f�� ����J%7U���v8>8�_KK����&�B}�y�p��.f, �3���d�R�R��!�}�'��l��䪆Ե܍I��'|�s�_��-���[�x��mh
�;%0� �C(<�Ч���a�W���� �B�������ԓ9*�c��jP���+�L��>Zޞ����J��i��:�(.�fzb�JE�t_��b�q )8e&�6�����	Te�`��
�p�@EM�F�K�q�d�?���X��1��>���|�y�9�i˪*�
�fר�U%y�kM,��XX8���sǱс��zU�L�&�[ք��U��r�5p�=
�F��NO��]AHD����R�p:ӥ�a�d9q�	.<'T�9\�4�b�%��(���9/�/����AQ�.�13C�^J�Y�-2W����TN�̦��ZH�-��_K�'�V�1����oB�If�^�-WW�i|h[n��;��ݚ��셐�6��	��A��VW��4`E/�0��G��Scp8�s��:���ͽ�1���~�:�0^��W�táIÓ|�䙚�%�Č.0�iR*����#�H��I��m��)u�=�����(�3Dя���^�y��*h@����Y���� ���:�i�Zs��~�u�
��^}�ϸ��zq���yqo�5��}~�H5��[*L|~�nc�~���W��e6A[� Y��$�N�@s6"eguO�=/7K������J�	!�S����ܥf��
�q��n�ՙ
����ZINd�;}�>�݉�!���6xf��EDEx��`dW��F��Y��3�:٧�hd���&e&[۶�[�}�[q��A�]��5�u�+i�����?ӂV�C�M�=7�O�6/lo�O�+��g��-�?��9��Tv�.|pG+8?8p�U�Vر��u�~����Y��x�u-�+Ey���{� ���ABM��&�C�zU�����=���<�;ݎ�^\���Zv��,͏s;����PB*/O۪�,�6�
zĸ*oyEJi�����@e2Q��I~o�҃װ���V!�D���=���t!���-�vK�e�\j}��O��T%�
�����Xw����z�`���=��V:z�X����]Y����5eRVG��ź�+�.G+�m%2؛ݱ��EͤI@�}����؏�|?)�W�U��Ge>���s/K��GZ����9�ə�S�It+VƸ��p)���C��V��\$6P��JD�>f,Q���SmIH �̾��7�q��k�p�[���*U�tG� @�_JS�{D%{�h�X����������X=Wz�	���ގq\���Gζ����Z�>���9��V�c�V&�IUDu(�����q���$we�o���Nf!�]�zQ������*�� ���ٷ�=�f�b>��jd�&�9'����G�y�	�t��vdc�G"�fs�_�Oc��Ԏ��{�9Ha�^��ݨ{U�m�6���ei�R�z�f�UM���s���Q�ϳF�4����,�1���GO;��r��Z������wY�^�	����O�v�ze�4Ϳ�f���a
�X׽�4��r[�Q@�'z�6pl�i��sg�8�@p(��{�X���Y-�[t,�]�r�(�$�Iܠ�W��fl�w�l��0|�#<V]���BL��������rH�'Q��y%��!��FQ@"����vͶ3�hFBMD���W�jv3���Y?*Tj�a4���_�R��`W:�;��p=���������=��璸˧��Xh�5�C��V�<��溗X���7�V HP��_��,#,S���[��^���VC�!�Џ������1I^MP�L\6]�nZ��vZ�?gP98��l~���C��;��?(Cf��r�՚W��A���0�f�_>�zh)�(ǆ�+3�2@'n�ǣ]�O�[M��b�NkLYM���hH���!�&��1��bR�x�(�~ߝa\x�f9�6�XJ�t��� ��`����bGp|w=x��ak�{���O;��U[�M��f���E��iZ_E�l��j�먠�ݎ�'�腵�d�M7��z��I��T� �m,��Qn�M�^xq�!�����9��H�>*	t}
��o�u�:;F�P���!we+�!0H�\ Q��&��3nqG�@fO�,�G��B��FL����7m�C���r/�U ܔ�~>\��=3����S��%KF������B�[��"$vH�2y_˟WzIy����7v�ު�4��-�p��}���AB�M�}Ur����
��/}��p'���)؁g'2��\��aOһEqYd@*�ol_zRAm/e���+��^�g0�>�+��f6�53��Q�{RMi�\�"�S�|�s���Q�y�f�\g�h˳��X��;_���&�>�.ɜ��ff�-��|�ڶ�cC���_�B����� m��m3&0'
a��*����k��<���o���ܨX�x2sU�rV�
5��v�Q���^�B�'Jg8� ����L&��IG~f�c�-���>x��<o$��������Ҋ"�B]TXv���z�*������!0Y�l��a�Ц�7�����&Zvx-Z�8��~T��~���
��D��H0.b�b��ӿi�.|\���q�����1~�`�B?KLY&4�l2��K�[�!|��|���_��.QV�V�o'4�y��@�0���-66�>6i���RН�f���b'bh�$ï� A�\�N��?�_l��E�56}T���uN�L�b�t��?�:C����2)CD�2Á�����a�g�Qu����ˉ(p���/�5u��@vp�&��6f~�����Os'��\
�xd�K�FNH�VT�,W��Ŷ�G��(Oz����z�E���ӈ�;���כb�9r�f'0�xݟR�D󭺅��l$t� ��-�6N�����`F����`�?@�����I����UE�q����Q�/)�s����fv�>eCJ��#"��h�D��1�jZ[3�<�b0�m��FY쐔�l�-\a�>�1˴&$��
)n2�4�7���I�� ዆��"j{�酥J�W�>��t�.��h��T�n�H�߽�3��<?p�t�_���E�`Z9'��#�DRАu~�t�!��� �ѹ��C��\bQ��Bn�OVoR���ƶ��GJ7q[��8�:�G��˄�(v�.����#��ˁ�V�c��*��ް�7���k9�{��΍@�@�{U����25�:dE`jqQ�ƒwy��v� 5t���>u"�|c!v�i�*n1,��w����m(�XH
��9` ��Ѐ���q��J���js�@����a0X���+l��oW~�Y%�P}v�7����!�K	�O`l�dd��\�W�?HQ@eB���݆q�^�b�X���-D)���KEV��~��1[�_�W���ށl�G|����/��W�vv�2�}����H�#��p1Ȝ?�oo�,	|�U-;[wy HQPd!��֙`4�L���8���[���i�kv�9��IKC���7�C����4H�^�U�֑.�A�E��[�R�э�l�^�3g̘��I�?�+�����Ĺz���R�4�����
	�<�\+�@��)��Q-?HR-��(;q~�zt�����ݘ���%S�\��܈��s���}^~뎡!:X�S�)P��Tćd]"芫�=��H=bj���m�F�.Vr�x$#׎Ӊk���{��{���Dh�4q�f�Ums�T�*و=$�]m�^x��g�X��Z����6����[��L���t��]���(�O�m ���ͥ���W��'�>ȼ�Q�b�'�;�1xO!����"җ�I.(��8`K�)l��^������ea��c]i���g���zO�P�|π�����\pT�qb褰���~�<��M?t��W����D�I���x�d���
U��ͱ�S�!#��s�Y-�'�*P/�%�_#}رk������r5K{B���2X�̀{:T�j3F����}�ڏ�� !rHӏ!���#�`��h�)�x��4S���GT��<��bYj��Zvg���{;���P�B�#c��9����!�h��.ό�W�W��oB�p�0�I'��ϻ�t�����[��������yO�V�E�4�]�/S�ŗa���3�4�d��*�H��1�R����M��S������Y�����e���G� �>�C��G����N��
~[v\��O����K�ٸ�<��n1�[:�@ھx񥔄Vi�	gs�w�L_4�K�<���G}��U��\�������A1Ɯ�#�Mm��1-\�2-fV�9v$����K���>}�U���"ײ�I�>�e����M�:��=���G+��V�ҿ��o�j0������h|9�N�M���w g-��鏃�'�h`��S������(JE��JFq�i�7�d��\co� ���o��I�]Jz�b�������&xrQ����Ap�Sh�*v��N]����.��vE��tuk�1z:�:��N^�B5�3yi�N)��W(�a�2"0ǵ��eQҔap0.T��3�PI��(�C(�)h���y�"�WC���s3#RB�}����G���g�|�%��Ղa��h�rbf��) �0�bf�J�ڇ���u	�Ƴ�b�oc��"_�� L�e�w5�uW�N2{;�2rGԪ����N5�f��A+��������n �c���6�z5t{U��`��f�hPf�,~f&o2���x��m�PI<^��N�u��8R]�����/��(�ʗ`z��ϩ~H�>rl�Iy��®�_NXX'k,�6�Yý��H��ؚ�?�l`�'���OO/.���E.��^����]�����,�L�e��&K���G����{�Ō=�k��(U��Y|tvG	,]`�k���l�a�	p� �cE�+�*x��s}\H���t���u>���!��1E�VrH�o�9������=P9ɩIvs�_W�`�)5��^����쥐>��
��~T��~�����ތ�a��	�m���E��A8ܵ���:��nd�IG0T��� �҇"����,�0R��C1G�ɇ.�T���T��R��� <�z����S�)��:iP*8��z�hN:$�]v�jZ9\L��O�<m�`���u��_4�w�M>���u��DJ���G���>��,��PqN����Yx6hO�|�����MB� Fz��UT/� �F(��o�*�W�#�49Z�c�����|��;sL'��읙`rR�O@P�ڜp2�Z���h��~\cA��Ԑu�8/�BW�<i�i��j�-�9��h�9A>Q��h�3>�������-L���'��L�r��#/�/9s�p��c�1=Q�q0%��&���ҏ ����Yo�VQ5����GA��}^q�Z�����}�*͘��J�]oҍ���6�`p�ʚU��v��v�c�N�j�UN>ꔧ�^�UBuzT/�Y�%��D:��N�@���J��'oUX$d뉢hc����bG�N�Or/QMڝX�t�eaO����~��9��Ӵ�`����,�2� �:j*T�"O�r�$�&2���>E�����%u�)��R��42�k$r�q�[\-<U�|	T1��|�ƀ��uسFjo�[��W~�3z���yBG����y�z/j����6;ӣ�f4��:�bt���x5���t ��]��o�g�ާ�R�Q���R2��yO�$�3���յU�����L�;��>Ói[��8���& �*�f��*�v�"�Ҍ��䤣��#�"&�e���㻩&(N]�~0�����K:�������k��4fk� �gg���p7Q�ҙ���A~Ԕ���,YqC�5.����JŔ÷��1�秝y���@m�{�0�����E�;�U�_�x���tV���]������XU����[i�/L�V�F�y�~{2.���Z�ƪBq�3ɷ�1�����䨌���i
%T�썌�`]X�s��A�4-34U	����&y(f�BE���>C��>z_��S��FAO�N��,/�kT�^�i��=>�C@<��>4��׶�z��{�.����$a�-LQ�j��.Q%t�};a ���V���,���oU��N͙��݋��V�p�2��w�P͐�0�5�O0|9���6�JlG�����.�"�=a@��G��UNf���)��ˍ���*���?`�]U6J�kǜ�T )آ���*�ɑ�B`�d��#�o`Ɋ��椐�!���jC�5����(�1�x��~@�=r���h�f�'=�\v�
(��Jw)�E�O�GKD����T��h��h/T��"E��8�[K���q�{	~y$��z�g̒z��o���p��3�7,���g�6�R��|Le(�7�O�'��Ѫ��|^ C�ӷ���z�:�!�b�>�,�iOw!��7z+�D�)#�c��dP��2����H*���Ȁ5�4��5g|����*Fq�,C�5�����0��/��e=0Y+�{�L?D����K�{F"lG���͡j7t>�Y��gw.&g`������W��]�	�tf��(Ȑ��	?��gp'�O�B(��Y_V�JN+Iw=B��	j#nU��g�GO{�=(ET��}�6�^��9� ��T��?�J��u!.3����D�ǵ�VnԜ�<r��(E�*��\�Z��R�p�59 *�b̏U�<e�T��	���lX|���N�>��5�x4n=��|ջ.��Dz�Z���'�(�Qs�ފs�5��DYOQ��,���l�VHy���?��㑰�Y��e��n�ܖ��x�7�0��/�w��G��!�����zV�\)�E����1+D���~1^�����O���9�*��T����y��5�tr�'$ζ}��i@��V�;��h�Ԃ�8�]b�..��$պe�_�t��ۺ�@�E{+�Z��[Η����H꘴��DL�H<?�LcJ/.�6g�OHI�!�n� �h�m�x oe����5܊�5׍hoh�� �c�g�u_�i�q�+�Z�Dyfy�動`v[�U�x.��������P�7�{܆xV�r���:z\&$sN�\�A��L��l��ݻ�^��Ùъj�yj�DQ⮌1��	�چ���� �ׯ��¹�'���$�B{�el8�)�EW�T[%��p@xs��YD��zr�~#���f60K�]2����5-��VK_0�<@߱SI��J{��l��8êiG�����0'�?A$�qH�B�T��G6��:��{���K�����4ҏu��L��mګ'9�^[B)@a�4Tˠ`EG�ƴȧ���9�>������&��{>%խ.�CP�a��ǔ��E�v��ޓ[��n2;ә��zY|i�A�:Ř�.Z vIXQ�΂����s��I3c@%aw8����5��	��nv��uv��qx1�q���AS���<a�EA2�fc��CPq�N����x_ �|6b+�
���E�w��V��(���RLu�">����d�����Z!��W	�pq)#=���9M}��.V��ӣ��C�(6�ڍ��̒���Nv��L#�`u�}�`�2	R�y������ب2�~��yO�	5���p8�i�uYS�����t�p�?*���#糒�׉&B��+ҙ�ړ�GBX82���`�#	��U�dXy�
�9g�6E&��k��C�:� ���~��_̓�R�_��;o2�̵ܵ����M��8c��P	6��{Ohj�E�gϭ�*�p�%����1O|��>ɱ� ��� ��#ũ7�
"�a�v�|NY���Q��^k*�������� h7�����Һ���'�ꉽ��ْϽt�J���v��>�>);_[��_����k�ީK`�ֆ����U�d������lS�x2����F��
ܕ�������N�%*���A�&W{JC�[Y@�������J�
}YD�Nr�1�"�9���E����v�g����m��o!tI�	�;�g/ ��`O�y[�pCOcs�;�,k�+���qEG?I�w���$aSnnٞn����o\d���v��qI�Z���c-�[�ţ`�l��_l�0Gt?1[iF?�$Pk���j̪��#�?�ź�,��igP.��}��gD�v#f��^/�}��Y|�{��\ه�E��n!�5�����N�����j+�
e"k�^VЯ�=���Hz#Q\_t���MLKi�)�G����QK!��e+�p�O̜�'n:���z_�6�Q�Iqc�-����0?t���B�5j�'��!���{�u:����3��lA}!�(�8"�w-��c�H���LP��cg�(�����:X�AF�!��h3Oe9�רtWr�n�yh����T�c6�u��Uܮ�zM:��E�/���|�k�RM��B�r��9��QId�ß�YD���͖b�H�Ř2��Z�Y5�bZ��c'ts"r�A�g8�)N'�{m�dጹ<�&e!(ȍ�����i����Y�,��mh��DDk?�#��K�:��y������l�Y/�f��h#�d�@J�k��s�����coz��b�t%p�!X�d����Ӡ"���d6��h!���6DB ����۱+�z�c���J�[�5��I�?�u#|��l�rtA��|���� ���I���d4k� fW�bA	K��өG^rAa�����D����I��x��B��S�W������:��1A�n�ʔ��߹"B�\��<	����<!}}�(?�FҾ͉�������¾.�����-﹄��J8����f���g�z��#yt�W<;� >���|�B������Ɠ��S���6 N�#��R)w�Q���Ci�ڀ�ZQ:?�*cc[��5L���J�b@`���H3���d��a��� ;vG�-K2����g:�?*rqk\
�(���T�-!�H�\��m�޸P���ҁ�03�l���bk�rK{���Z_9�c-�R��|yifPnl�c��8eh=C�Δ��&"��[~t�st¹�e�+�)��ǹ���?#̮*?c�o�o��DW�G����T�$i�sO�uq�r4u��eE1�;��p��#�:�2��L�+��@Դ�ek��{�	kނ�)Ii����5r�w��q�Bd����D_�חL�~Њ|_�!��UГ>��v4�&�D�|N|u�j��8���
������LI�.��~/�_~�31�i]���e�Ź�e�#!�/��0���;��l��A�C A$�ȶtg�g���YhO`{�r�D�W����x+hw�Dy�]�k���lJI��Z�s�
B�޲�gw�n�(���N$�E5�(�&Ho�:�~�ߋ�&��m ?Z�����?����7f5)D��i}dƁ�V-�e�I%��v�Y����թ�5�O�,�N{ �?�q�i�2؛
ٔ��o��� ��g�6�3�q���Up�պ�(1��s{O�}�`���+!�� i{�qC�z�P���YM6��\j0�������}��[������AvG������̟HdT��W�?^GE��^E����҂H"V��F�N}���	uUL$���o�>l�P,$����Q5�h#�=������s���i�.�P̟T⩛��#m�L��暟��f�H!������)�g|%�����I7ez��Q~1��,O�L�!	xZ��C��3\ї�&j�&�%� ��0���K�s4f�[��1+�\��(�o�L�$!��t�q��SGq�Fo��S�A8�.�O�?Bhޟ���i�$��r�3Ϯ#�61�`�VX~vozf�Ջ?OXZ��q=����4P�s�(�!8�$e��1���ޡ<0�<^�x�m�PE�fN:���L�3�ّ傿D��\��:�o(�{�����ɤq�xC���.	����^GʳpZ 	bc8��t��.s9O*k4�"�q����a'�A�+��^~����Q��X+�S<o^H0@碉ʌ���.W230iwg��4�")դ�_6��$܂�}I���vyF��b��a��K�D�cê�+>T*�|�`����a� �6�h�YX��"��~�
�|d=`Nq���#�87	-��劻���6?��VC�Eșj{���T�t3�:o��-� t7j���p�oJږ6M���G%2�e?���?B���5��<x
�X)��)��H6���T �b��/1+���?���������ڧ�U��'��u��4�0KC���2��s���8Ǉ"s�uD�HE3EE&�jluoJ���Cc��cp�z��rT���@+Ɋa��.o�@{4U�5&�
J���.퇻���$0��.��(�i��!�|�d����2�>j/J���鞹��[�!(�J{��$�xr�1	������A�R�j��I~�sbX�gLk��}������q/��F!g��fK�;l�>��TY�O|��p2)�9y05��+��l���4uA~�4�m�C��Q��p�)�N�)ʉ�������:��]��O�2��U�����c�*���0�!�ю~�1��,�ّ���g<}9%���+D$���HLv��0l�-3��n�����N#��s��Ӿ'�M��$��qD��'�ȉ������p��f��h�o�aK�&q_nú�t��l�y��w��qb�Y�ı�_���LIb�~��w�s_`Hj a������3ŕ��i�^n�bz �y�/(�񲑅S�H���6����\m�0�6x��$5J�V�.���[+�9�,?�[���N����)Z��V�~�L�t݊,��O�׹_����.<`a(�q.��
3����E?���os��[a)�,��h%�#�=L�I�q|�2�{�R+�{���5�%,l(ܲ{6������-,��]�0���G���yBa�ᛶ�(�M��Y���O�>Ǯ�`Bw�.����젃� v�F��Ѩ(Ͻ�����O�g�z�S*AS��2!���F8�W�Aa,M�H���Wi�]�v��]�%#Ǖ
D4~!a*$,a���x�����F��H�i x���:.!�V��-�ж1J��� ��'��/�F�K�7#wA1}r�n�|�>ݣ%�9��" �=��o���ːd��_��� w� =��L��\doGq�A)a�C��.�Ns_5Y-��w=��WΉe���j���k�l$�K��Uܹ��؟������<&7uߪ1 ?+oB���Mr-�h��'Vi�C{!I�w��7e��u:Rk=����
��6�q|Fg�dK�`� ��hݴ�|O���:v5���Uz_�!)O�I��4I�2Չ6���Y��&���W�\���}N�>P55��ԩ�GO�:�BKs6i���߀�k��fP�����W���:�F�z�ÎH�����-i�[�k�v$�'xmZ�=��R���K�\��R�p�Ə�<��k����O�̿\�����R(�9�i��v6t����8�8@,��]5,E��pz&�E�(�֜��˼����	T���Pt傀a�О��	�{]����h� /{�~"�xw���V,���L�$��п|_��U4p�`cܐ�D~�AL+Jz}����d����-Q��xHo>�l�s�g'������4�� �fv(����o�(���JkQ-�ٯ��� dz w3�_�V��ź��g�R8�+j#����$j�����)E�����OP�sp�'�hJ]���.L4�nX���n-���5��C}������U^b���� 7��yi�����8���ғo��ZW1��Q��m]}������[j,7sI3=��������&��*�J�l�~�����Y��4b랟�o0�/�������-0$]^��9$�rB�7�fyC")�?c���A����U����$ݯ�3m�``1	��~-N����K&�R��KⰚ�<�==���6;u�;�>^�HB��6 ��)�	 ����&�<AfכS�����xU"0 hR�2��D��h���6����W���hKUS'�m:
4������X�:Jl�sb���G<S.
�P^|R>#�'oC�����zF�.�O23U�}&@�`M��X�ǌ^���?�l��ͥ���x@���-�?N��v�K��{b��+w�ٯ_=az)г�,���V�/�Cu%����fg���&�&�����o��_@��|���Ǌ$4�u��kh���&p.� �'�z�=���A-�*�����G��*
����z�A�&���?���<w��Շ�����Ǥr���H%��j��Ӓ疱k��}��5j� ��֯�R=άv�Eo�2����G�{a�x�.��a��?갟������Y�td��)��a������Y����JQ��:����n��H����`���N���Ͻ�)��S� =������n������_����7��}��z+�=���۔Q��d�'j/l
��9R�������@�{6/L|��d���fuB���M�2۴���p������mr�'���혴��7p>-ڂ��h �q�d��*P8`���Q����;�gru,���P�9�����X�N�Z�����_��Z�s)P�ͮ<��H�*,�k�7۫��4q���}9��j��~8���\T/G3���7��|0H��_V}�{�dP2����D�px�#m�2��2kn��xxK>�5�M�1��q[�&TZ�*��������5_���ƭo���ҳ��� !4m
S�4kqr��P�G�}x�z�����{�����=7�[�n�c��ӑ��=A
��rU�3D��p�Ċȱ����?��jdrrx��l�u��wn�I�{�u����C*%�)�T#��w!�G�HQ�z�7=#��&Rr����@��0��wm�+<�u��,��F�N�KT���@���pQ~�����z�L�D/@1w��Nc�q�C�G�*;�I�x�(s��;����c�+~_����3�+�j�i�f��Gɰ��g���TQ��� �����x�32��ț"���8���RǨ9r�u`��Tm��WhW�i�o�ui��V&�i��qC=�F�fevy	mڌ�x ���w2� �_�s'#gɘ�'b�d����".�`/[e� �?�귈�%����pg��~�����̑��彨�I���-�ڳ'������m�M/��|��,��� $�\��w��	Gi�L���jgǂ�c�Bl�{�DH�Tu�����5i+O�7���b�,W8A�X��R:øsW���l��^'�
�*��҄K�J�֖ZȢ�攝�]zp��`t��g��9�d5�zQ���¡ab%�ى��!MaJ4
��*�tV�|���I�+�l���\x�5��*�F)���P"YG�*�tER�<"$m����yע���W����hJւ��EQ�|�8�Q��FH��>��:ЎP��`����=�D��❩�����*"��H�����h2Q: g1�Vd������zF}?)���]eB�m��V��|��q� U�D�w(�v
s�����L������L'����W�;�L�r�VEi��U'}����#��B}5����De�[��#��L��ꄌ`�?�[3_(����M)�\�,��T׿�P@W��P�t�}���46o��\�G����e[x]D��>�Px76� ��M�$���_����'��f�8ꗝϭ���9�'z >�y�b��{�l�8ծ���W]�y滮e�.tyu�S�M ��9�=fػGF����e�b��D"����a��(-g�}#ԥ���b�1x.Q��@7F����%�m}i�����i�m��ly��SS8���V�O�`���b�����C��`��R.W�M������D?�bi����z>�ۜxJ/3�D�nd"�Ҹ�OY�UN����V�y��˥&�!�P�
��1����uY#��1<� z�h�v� S��yÿ+��~)�˅ډ=�[V��g��-X��/q���}մ�+��<r@p�����z(�ްs*��9Y�.b���b3�q�9�bL������+��Q��6��]K�����$�ɤPU�
�`�����9�.�+Kc�p��F� > ^�i%��H�R�% ^��9�h��G=����LD�	Fu�`jR_4#�߅y�*Ԋ$��]���z�t���*Eʢ/��'�k�oJ�Dk�(1�<�=�j�@ST٪����nK*pp�/�u$�s��˧�e�>�ԏ�{va�bv$'�����:$��2�&sz [av�e��J;E�5Y�8Of�Ej���0�]�$c��}��H�v��;��T��/,wRڑ��oK��6v�YF$%�tt�>]�.�٤�3�h,�6�'�	�t�#��q��s��R� \|9l �Ύ(��]i&H�Iʝ˼Z��)B�y� ��<P��Y��a]^+ˮ2�9m���|����6a�������N��Bz�!q�je��^�:�� XhXD�GI=\�1�fBA�}������+믚S~D��T�i�6i2�#C)�e;q֗@.��>�ٴ�k�e���e|�nr��7۵����e1YZEu�j�iL�N$�2��Y0꧞�p�l�������1�Uu�7i�֍����g��MI�`9
��%c��Jy����9��1b􀺬��.t`<�)�Ņ��2{M�ĺ�~����[��H�a0��XKX;�١�Ϸ
=��-r����e���g����7'Gq�=ȏb��ۦ[_lVסM%w�L��i�cA� ߖ�\_�"�Rg�׾D�T0X���
�OW��ƚ4E"�7&wu�R��$<�.G�:�(��H[�����C'��jg�:�F��;T�3�QɶAp~]K�[%C���#�X�����D@u��5ॹ1�ކr!/F�G���y.�BS"I*%c�1Iԋ�q��{�1w�W�-PA]�?�Ɇ
�*2�1x:�,GD|��ؙ2�}_����T�w[���>V���N.!�_yPA=���heeeC�9��4����/�k�[mF:S]��ǵ�AJ�~��l����y�i����~�7�D���b����ux�̂珡�� 4�擄����"6�^Y�2�J]v�~5��G�RU��j�m;h��"�.��=��D�����c^�r=�������T�;��9d�_@ ��+�O�\�Q0O�`8������q����ĶQ�U6U��?�^�A��ϣp��q,&ZIN�f ���Aʦ,�08��Ml���n�ύ���n?��. `���`�ׯi
��g��G�W'؜�����;8�Ɗ��2�4���9�6 �<��F'�ubq�v��E*{.VJ{5�_|��)0^�b���p�oȌ�k�\�9��4��&�\'��Y�;順�����aa����I��:���DY��d���1�!��S�}�oc[5���L:���Hn�˹��Z�t?ЕxP���7��ɐau�V~�-��W�:�ƞ \�if�`�l��Ѡ9n������a
g��"G|7�c�};fg��=SR�h��q����U�-�-��!�WO�(��'��_x7��.::��%��e�x�ݴ���]������mg��RF����+����� �2�Iid��0�1(�� @�H��Z�Ä/|ʆ�e<������/p�"�q�SY�:�/F��}8��l��כ"��nǔ�c��5펕����G2uR��s43�Mi�q���]e��?�}\W����2�V-���:� ���i�$#@ECN�|F��Y�6^l��^*�;����Q�|��l ~�+Ba&��-{$�֦���\��38o�l�%	�¥��^h2Jɨ4�]0��Rd%^ N�a8��RY~"�]Ӝn/����6�?��	&�w�3������7����@�������gP�.N�����Gw�>w��i��{�!������!/+�R;�>o��Z'�0겲����y�m-���ymd�!	��:�����#�Ά��f����;A��ٖ*T�vt���4������0�O��,���lؚK�B͖�M=��B���Yw�qHMGD�(K4��W��t= /���o[�R�M���s��A��pFQp�(���|0���RI�f>��P��@-�u�d��'�B����`_�6���4�E4���ݪ?��0���9��24td�$C�����J]k4��pķ �°��l���P�@^��g �9b��FP\^�����v�$[6��c��b{�޲�y8l2	��핺	������W]ˌ{�j�7%�|�K��ȭ�A�R^����C���āҲ�Q�9�Ki��	U�ѡK�
��M�����c,Bk0��m��Č����MZ[�x�޸8� S6�/���8��U�	S`9 h뮆kl�$<������b}y:��X���G�|�'�G&8g�@_:�yde��5Å�Pת���]�Jjk��N�y��(X:|���D��;�;s~�
�0$9����g��z
r�ۉ���*��rx�&dךcr[�ǅ��U�nԿ��=T�_��TV�>SâȞ,:��f�S%�o�H;S���_���`��I\4 !O��2�������q
��dy ���'ɤYl�ZVI܄z%���4������§�k�,o}(X��l��#����w'0�:�Y*u�¾;�n��s\CM#��㠶��׍�1��ʧ�QBcR�F����E�D
az���@J�K8>��]��p�<�`�%�&����#8������3�"yE��1dYcV��,�v)��p]Q庍E��Z\5Ŝ5�WcTc������Hv��H1C����iZ������C�����زln>@�X��O�7�@�)^	��pڤ��m���}�[�i�}k@*�9*J��o��L#�a&*k٠�i�A���6�	��N��%kM3�.E�i�(1A�LZ���ŏ�|eӎ����� �yõ���.ZPTw��-181G��ĺH������K���]�����;_][��p��L+Ag.��m�t0�`Q�J��"4*D��da�e+P�M�&f�jxH���|C�Didif��3����v�|�ʖPɉ��V=��smk�v���!R[OS�s��丝y�O�$�+`�r�^�}UiR3���L!>a�,��/D��WJ-�� ��KeT�뒳��.�WV�7�7��~6J�]/Bp�+J]l��;g�X�P?�ް�%�+m�J��<������-��6�u�뼇"�r8AuQ�����y��NgO����[.9��T����aQ+ςB�6#�Y��6���8H!d�Q���@�4C��+�gSaۘ��wY�"']a�e²1''���
꧆���Ek�6�9hp~ �p-k�*��L�>��]%*��w��*5��c��z�d�5�[�o���y���ԣ���F:��
G��v�#�QK&�@��o�&u}����Z�7<ۄP9�x�A�@�D�O����J��J`�z����9B&�Q��H�
��8����`2p	Hm.�ǝF W}'�D(�r�Ӟ�Zl/IԔ8��g��'����&�L҅����agv�1D�A~֋��19��	��S����?�ig��E�.�h�MK>�ܻw��y�O�`��Uy�6u��+��B)B+�A�Y�1�T�N�Hk)rU���_8՜q�E���W!B\�1.�>o�����?�C۹��L4��U��
l*�B{�O���$��8�o�E�Mk�9����fp�0�T8K�.VIǈ�Gc�� e���\���.jo�.P��t�WWJ^����
"z�R�փܮX�rށ�a|���R�\:7��l��6�'�ӟ��S1���F�b�v���s�#�F֪�8P�4ʥ���jX����+1)Jk�纝�o{��5\EB/����4����+읰����nv�(���ݿ��I@9u�;�	*Ref�`aŕ5Ѕ�l�\��څջ�e,�@f*�WBn����\kP�e֎G¼���QH�^,&PQX�O#�#W7���z���%��b\�iO�����:���w�<��x+�9��?v!R����N�W2b�v�"_�T��Pa�t�YM''�yΐUSF��^a��*�W{�:,��%���f��C���k��)������~���C��L*�F�vk�������֟Syf�gN/�?�Nm�<i�:&}����)q�|6jU�M�u���Wc���3!$i�<�=$��[��=��	��=>��j�SS �x{�����pᄶl\m��jiY���R� ��o�1;7Nа���h�� :���i�E��u�,��&-��a����$�'��z�ɣ�(����Gz�{��/�)���` ]iM����i��/k��u�����/X�{R���׍�T����W[��A�-im�%�Qh��\!�=��_%��n������2X��^�~��G<��,�-�ь���:M�૆�c�v�Э�����N<�uKm��X�[g!<	4ޢ���?Y��p�.���O���`>m:�:Ә�Gz"Tqb�@m�����~� ƹ�<�*?�$��AL����J�����:^�WȮrn�^		Ϣc���}�@&7�^�v��cH�,A������3?�� t�ҫRz�2��[$��6pGs�yz	�� ��ޤ�23\ b�5��f�k���4��=�k+��=Zf���v�2w8룂/Jb�|���V��u�g�:j�Nh�%�ab�扝*�J���Cw�D�����(�j��]Ug����V2&=l�˺0���AX�˵G�E�褭<����������GLs
>Pu��rf.��k�\�@�g�v�6�Ms<h�	'B������m�c�b�2����P�t����\!Ϣ��6��3�Е,�2W�m�E��c��H��V����^
\h(� ��� ���s"�I��FŜ);��W/�B�wL�->�c�Q�9f��-2�"�A�禎��0'&����#[6]��,���Y	���T�QiY��%y���^#��(���3���� -*R��>��������l��B1��~ki%�\��\7^�W��l�Gb-s4mٱ��޾[\	p�)�G�����;ф�M���E2g�a��bۖ��I�$�֩����Դ�����4عi�T�q:�L$$��(~�w/|޾:��s����)Bo��x�.`C��1EAw�pť$j�)�
J�;�9��)�nT�����09zү'�h����v�$xt�ztSp�y��α���K?��G��k�g�|l��q�6�Ĭ�EVv�v��=(�?���"����Ȑ�9��_���D���FԀ���?!��g�{�}":�a{�VcW���Ͳ��є��¯ه�.��]�N���`$٪k�s��K��g�&F�&�&��s��%-��2�T�Bt�6;̇�*�Zd&�r�����C)u��yicO�HƘD|���C>��\K�	������TW�p����U�jF�=��~e��.n�`�e���ԡV�r?�!�*&q���M��l|Q���v�\0��u�� ���}�fŬ��ii��Y!/ɐ�wC���hg��m�h	�7>ʞ ��	uE,班�{E��{�ۻ��W�	C��kc��]�\6(��I������ݖ����#C�U�{��u`o�z=2z��l�"'g۟�x��$�ꊹ]\3����Z�/�����(�ɋ�� 9��o{}}���"F�byT�'w��,��Rz���B ��X�[5ͷ�Pa1�Pk���$ SCΏ�5�c��֫�؈ PGCM*�p�FVߟۙ�w���34a���e��d��P�2���5o������l������'�F:xծ!���,��
4�훺��t�B�7��(7�.��<4��,��
�;�ܭU��NYK1姀��F)bCpȧ���J)ǐ���
����'֢�u#��E�vG&C�-g��f����&ܠ�rc����B"{�ӭ��EuP�lA�yʥ�m���-�h��\_��O���;�bGU�`
����� ���;@r�^�7'TC�9`�E�N��������Ɇ�ul�CR�d�IǊD:PIFr~C����~��;?f�Y��cv�!����v�IL^��2rNs��S��f<	�N��W�@r����I�;X#U�Íi�Ez?t��G9���+X���D6у��I�nR�Y~�Y�x���2�e����ý���E�k�T�(�G%5�P|J��\����GM�0�QE)"fd��|돸�"��*@�?��-� �	�[w-3B8?uQ�ṣ��h�{��e
BO�(�*��7G�@��}f�ACV�!!�LLY����	��[G3�R-�cA�!��U�!?6R"4�t��`�������c`t	��,���V��Hit����ne��]B/��6C1uM�P6�]Xv$��ExixT9M��չɮP�ϬX:�����K�z���4�B���*	H���*�o�@hB�<_K��\XD��l��"�����DL�ߴ!�:ICc�)�F�l�'7���X��K��K��(	�]e��X�>|�"�5`ْ�ɕ)M��pH��e������9Ua��vr��5�s��^ZyL���%������:��3e�<�VJ	L��r ȥ˾x��a�fM���N� �2L�T¬I��~�Z^#�3�M��� 2E�d��;�Mp���)��}��T��F��f<	!4��Z������镭��m�᜶�F�|����#���F�R����ni�|�k�
��0E=�]�JC�	�H\��B���5��4�f�:pHІ���]S�ҍ�'[�&�C0~/r������Н�V���i	��e)�9�. �ׯi����㰩q�"ԟ(M��gո�@n��O��;�r�h}یr0�ö/�������5�5v�ۙf����!;I*���uQf�o��@G���Qc�Ǘ�Ģ�S�P֝6�K~�Kq�c�W�s�̨[�J��a�Gt%�/-��{f�3R`Z�Y
���c�.ǌ��<����<M��p���jp�j��w�-�~и����\�!V���K>R��ۋ��׈#Te�<�3�^[��B@�'!��c�*�Nj�6�?\ڪ8!r�>i�Tji�ʂ�m�ݥ���i�������{ F���ک�7tG����0��d�?���w	g��9���j \�̌�:�Z�ȕ�PdC���l���9V�Фp��Y�am͖s��[��<h��è2���_R�rwqʶ�7XL�,�wIo�E�����.�_����uk���<��̕��r ��#Ǧ��F��t�"��;?c�z�������ԡ�C�C��ٜfz�|���R��uϙpu����7R�X�UOk�MC~���y�)�^� M����Q�Q�MM ;Tb��'���u�U�o�r*����L$�2��wC������I�������bc*�#6�A�M��]�Xtx���k�����/$�U�+��-%���3ؓ�.b �%o�����2P���jHo���]Q:4�[3�\�}�n0���0.��M0���p!��{(z>�,2=}͞���j�msA��Q5�3�6��gq�_^�8�AU�h �ड़9�(Dؙ��k0�UGl���kq�pA="_����I#�A{9�
8��b�XB�JC��KlӠ���={��׹H^h���Ⲣo��������s
��u}΂�,�4\�=�kѣ�Gh�гZ)Yx����k��^����u��	&��9���� �Z���c�w�UG\�:\���Mt;TK�����T�l=�T�4���w ��"��'�(�l��iY���|r{��V3�_�V�c�:�)�� �_ӫ�Q*&U��Ȋ^r�J�����q�W�!����@��)s-Y6fn����=�������Pu�\SƋdY����a���g�'z���w$�
�.�r2���Ms�	b�+��U�u���6�+/^;W,�P��n�B�K�˅p���#����ëʳ���Њ�jV��rK줊%Jm����V&��[�"oU-�x�9tD��W6�p>�:����؞��_�i�Ds��S��b"��13�yl��'�G ����-�4j�J�S׺�*\ �W��e7���jJo��Z����#�hI��"r>\�^��PT6���5>�*\;��7Y���)��Ǌ��y�R����|�-�+�9�^�R���T��ߥ����e��Rmm&��Z�rd���r��5�i�9�zjs�;�%O����l�V^K�\���}'(���ߑ/w{��fMP�U��x�H�{�ۤL1h��뮸�0!_=���	abt���s 9]����q���x�<*.���d�c3�c�d��*�!��(��De��AK"�E�FV?�G���M5��8���jy���U�Mg����qE�K�n����<�0�]/�6���D�m6���po��T-tGo&x��%S�
)J��IS<ϩ����CW����8��q+e����@V���dE���E�����{�x^*�h;,�#ܛ��d�G������L(�K�V�Q��t�*��BҨ���:A�"����KclݕZ��q@�Em��!D��Q����Y���y:���S����q0,���q������Y�n��4�2"6�]'C�*Y�t�q��Z.����k�3>}Z�'�9���A�ae��I__���� �G|��gD�}hW(ɯ�I���y�X���OB��p�8MgRȏ�9�8���s�YYڿ���^�~��(�ι�t�U/�J�H0�}��qCD���EV�D��1TS煑�"zΪ�3u����'G�'Y\�ۢ�b��JQ�)g/��]�h����\.s�mTS;�$��:kimmʚ<7[_�<�R�Qr��T�r����lݞ�����o4��L7^�r򡐞�&�q��#��Zƞx�&o��qx�s��;��!PT���~*�Q��^�ڼ}BX;�n{L۬ �L��x�u�UO�bN�جo�T���ߪ�?��V��wƴ���D���=�:�e�w�՟w?��@KS>�q��"Օ��pi$�s�U��}�V(����\"^��1
w) ���;�P�a^Ee��pɵ�:���yb �F pu�/gN����|��oK��00��G�A�L�4İ�z���&[�`o��h�\%dBa|z'ư$[�כ���lhC3�aQb04{��t��@����YsoX�uX��������Ia�\��3<@������� N:թ�T��)_)��ӯ�z0������`�8D�!K#�2�a�5�F��m��I���|=HS���XV!��q8DCs1U|8�������[7��T�UɰE���äDe{h�2#nB�p�P"�~����G�j� 1^ڝ���c�K}�b�G�!-� a�}�m)�[��s���O������x &�����%KG�S?%j�	Չ�O�<X:t�7��ˈ���#l�f(bv�V��$i��ȷe�ru	xDɃ6�؆l�A�����p#�7
ݨ3��n��oR*��Z3?���>[��\D* ����ɟ<�_ھ[�h���˫��͕wd։Iw��֏nBEm�G�)&;�5�С�Hx�	��_�}�2�9�A6�F\k�e�Jl.�&#�A3*`�?l��iA�B�ɲO����E�/��H���Qă4�{zAQ︝ϼ)�x��"zBw��"�RD��v7B�u�{�O �Nf�E��$����4����l����̡�~2";p 6j����Td�E�Ұ@��H)��v����g�HJ�p��i�6�J�K��*�)n;�Ј[2SN
���(��̻!�vt��Z�����]�xe�W�)[�Yo$�9�	%ALCx@�t\W�*��l���Q �n�*�n\�;��~D�vY }����bŲ���l������A��*���S|�����+٬����n� 1�5�/Τ�%��G���1�T�Xa y��^O�S��A*�V�o�;�L��tWI���xj V0�s�¥��J*:�&���L�1�CF�� �X�6 ��@��[az���O�(D5f-�?Q�q��,f��xH�2u����w"���xP[jz��b���9��F_�}/:���a.@6�UI�
����'�I���8F��dΎ%Y��Ӽ� NM2��oN���^�Vx��BO���M>++����	A�Ƌ�N�L�wc-���n�׬�At ӈ+&��&�)�|�iфM�3z�3=�6�-�'�|�a���#������^iD?۟r�V��1����r
M	n�q�v�2�+r"��k~�) KX�?s:�����aPeu$��D�k�/����K����E�ӌ���(Q/���=q� rt��B[����M�w�w��@�A��cx�����|!�/��q�̾�hP���E�U��QB�e{ܬyA��6V�3g7C\��I9swc>�N�����2Y��J���:��Σe���-��ꫩ�P$�w�밍3z�^�������y��dLN�Ү�"� h=$-�A7�/v>�>���UJ�����E�0��R�5���a�ౌ�o��c:�ݪ��`u+�`(�����F�kjcai�Q�klFwnr��X��{�s���c���\/�}Q�ҁ-��#�y���Yj�'�V��JU	h&u�O�B��ِ�����`�@#��w�"�?*_�g���KG��	�}9�����A?��.3nV2 ���g��ě�h y��O+��:�dU`|���{k޴�C�@鴕�/��²����'�YlE�,``��2���z�i��A�J����'3g�T�I��!.���)v��hj8�e�aΤ��n^1"Kz���(��EǄE�rg�� �qZ�}�"c��S�\*�uSr]�:�`��u�K�.��L��V����(T|��{�� ���[+����)1S��Οt�.�ld�i	�"Ϳ�-�޳J*�JN#�a�DIx2��b��o�cr)���;Y@	���M��^] ''l�*[d���$�B�k�+,d���%�~��ß-�{��QܟCX�8�-*�7�Vي�4Uxz�t #W��ֻ	k�"+AB��2R:�Nt��BB���T��$ꏶ�<;�d�a#��K��G�(}�@U���w�>��yUXQ�S���e��Hr���J�U�G��F����L� )aC-و����1]��
g�G��B�4�ԭF�@�	�m�x��_�c�m�o��XY@[H(�mmm<�E*� �w�=�D�#�Tr�^�o�f�ls':Z�wo�w�ͅM�5h.��I7g$�tG´�632y���I�6��x�QJ?����F��lZC�33�ʒ5����+�g�tC��s��ȿ�aPcn�_@����d��T?I������n��&�1�=�({&� �zW\g�I�̣�8H:17;����t#����Fl\h�Q�C/� �@ػ��Xq�C3�t!t��N�K��U��T�|l#A�m�eL5�Du[�1�oI����Y!���	=��j��R�~�כ�s����ݡ�zH/и����sJ��Z����}9e�����X@/d}���۔���T�4lVA�.l�)�
Q) ��_��+*@�@��_�#�~~�E�N;L�w�;�,��9�������6jF��� SW��H����' -u/g�Sm�S|��T���:��ZK�@�:A��>	�)��Ta^��ր�Y�%��n�{J9�SqM!{��Yʏ"��~+�d
,xj�#�(>d{ u�&���N��Ÿm���=�VIֽ����k���C�G���3�5U̔	A��w/o*6�Cxg�@�}^ʚ&_6#|Y�T���
�ore#_jY��<mw�Ѵp"�j�5.7:�g���⟝�(E�����S�Њn�?��M7.�Ub�ަa����W�H�3�����������iD�}�z5��2��'2���|t���4U/&�N9��v�l�o��	O
�.м�%�V�m���̅f����Z�G��Ū�T�'yo�f��/����ߖ��k�;����RE��P��B5�1r~�ּ��!��~�a3o�չ�}����ap:m:Oڲ��b�⌤�NV�T�S97́i�{&��ty{c���[�⿴���<��g7:��DL��s� �\=�f�.嚪�{����6���
�fN�����a�	%T�vz䚕Ԥ<RJav^+�����ʋf�k"���?->�&�a:���R����ԉ�n��i�Of���Xe�&�b�d�á��eu�Z/"�����VM��SJ�{�G=��ܹ�5�Yo�CT ��*�3q\��6ςIfP��%�(~�n0�n�4�eS��h
'��[��a��"�z�����33���e��H�����/2K+�J����iN�����$��jp,����P�
~��G�H� 0ȴ�v1r/S�h�"[y��Xv{)�#4��$�>sٜ�k�!���c�Q4�壝��Inn����������d��؟�֚�<�7D=������X"7g�F2�(ڋl{���t�u9P��i��U��0���Z�?|��ê�`}��xw����,�z(�}��`_W?&ZP�!r5T^��IV�Ok!7���M�&��b����t��U,��;��7'��7yϘ	�w6���Ke~�ά����Nۯ�&]�����rX�$P_��8-�|{�~�?�\l�U�+#z�p�Dp��������t����)����w%�#\�B��TW���qb�k �Gq�Ǚ�o�2��ĖN3}�u釁y���"��#OYN>� ���h9N#����Y�7��#�8k��q�(�<lq��l���`�:���K�����A�-�cH{م�j��d�	jɌ9D�av��()Wޣ`咭/G��`��MV1If[�Z�\�}�O8�^� ��B?�ƌ�������S�k��y���[çZ=P�x8W~Q��b@��	���t���p�y#����T��܄�͖)%D��'�����*J	�+����H�t�0���ɍ�s��s�Ψ�\T�U�+
�U��f��2�j`����вMx�<�JA�%O����G!P�'<U���':zpM�����݈��<�n�ui"���1��ڭH\����8����"k�>zdθ�S������Y��P�`:��>1W{˲�^b���|��M����&��ӄEE��r:Ŵx+�0�R�3�S`~��J�� _]��,㚘�=(Ѓ�RY;�����=�bF��[��u��Y�{�w����vXf��k"���'P��Z�xƢ!A��`p�@�:m'��������p�W��`�D����_�K*�f1xZO[[�5�#�ţnJ��s�.����M��4�����k�W��n��8P�j�1� �Hm۪��]�B��QMwyWĘ����(�H��8G^�D [��YHP��.�A��WS�%R�'����9�����x���+�fE*�u�C>�t,=6���!�t܅����#�ma�^r���9��Q������1%����<�I\qV��\(q��<xҦ �'���[1�P- S�-L�Ш}� E"�g|����/���1���-��/՞:1���ޡ�����'_p������Pq�M���īg�,aeyZ�N��`n�n�W�<���m�8�B��d�j��r"%��;P}��U�+���!�
�CKʒ������ ���D3��'�b�A�Q/�u;A-���ýk,r�Y�	 ������y�H�U9�v�翠�8Dk}�B��Hߕa~��2���ʉM[x�C�N�zI7d)�|��mN��l���i�[%\�8y���\�����3��9�q��!�U[�5�5��^5�T�Ъ���g��YPKD+ڛ֒{�t��N�D�Ffg�T�����xy�H�R��aB�H��I��F���M�R�W���1�-(��62L7V�~ViMy�.-,F�1���i��pt�'8�9W{w^��Id]4�]��I���P}O:{H���+����\�
��ҿwbT��|d���{B1����}��lJ�q
]�̨��QՌ�����wѧ����\6�4w䈢?�s �:��� �Erځr���G��m�1�!v|�p��?qI��<�\��D���`<��vn�Q��[/�&Z���7�MF��2#��6Q���cZ�1�<M?�2�1�Ci�{�( �B�^�5���V�V>̜eϜb�R|�f�FԿ/����u�gd`b��g2�
\��b��R�a���)�}i�hn�NͲ_��Q�-6 M����+�F
����	�X6 )A������i@6��]7v���x~��t��ܢg�q
�|�4J�fgP��9C��<=���kG��2�� Rá�x�ub?���c�ԖU�ք�͡>��� ��~�-Û��EF�h��s�jaq�/taD)�5Һ(2H�teOh!�҂ ����>�����g�2��Wv;f.����F�L�c�D�߇z���KO!�s��+`j}E�1M���yup�32�>!���j��B�N궳Ӿՙ��"9P,��ƅ�n,3�����7?j�#[P�ÿ}Z�(Tt����$2�s�Sa�Dy�RL)̲��rm������f�	ū�\"�9�;,�㯀�2�٬�,lI(�{�#0�)�MT9��!�T�뇯���n�3[�p����s��
ݹ�jJ܆��}�t�7��\F�`��/	�}Ϝ�"����1ba��H�O,�~�?&7�x��f��cTi�(�6�͜����e �x��^�΢�F"�P�vYk�Uf�˽�	>6�+�/)ΟȀFD��Z���
}-����h���w��-ĖKP��=���\q��B��N
��X������l`�6��h�?�O�Kj�c��9�hL��V�ŻR����H�����������Pxj�u���z��*�xh�2����9���[x�fZ�`ޱ���!F��K��Tcn� ��̦\XHf�����6���ա���[�~��眡p�������_È�1`��ⰽʁ懍�n�.�?P��S�z7�8'�d9�^r$6k�^�#\@\����2\X��x�f�Jz�٠��K8a֘��S����gu�67r�*�
��\�	Bp��>̽�+g1����D��R�?!�4�C��>���}�ߠ�ljz2�[j�B=��sR�\�[-z�����N��u�y;���J�\��`�nn�
�JA;D&;�f�%(T��r�&oy�=�U��	�N�o���/rz����lT+�7X0��A���}���$�e������a�+1(pJ}�a�7��d�ʛ�C{uu����j	�MM!vܿ�`g+�~����Lj��|	_7W<!�J�XX���[���S$�<-dH�~�-WF�|��_��{Y#I sJ�<5��o���1�O7(g���y@�h �%�Q,(]��N�F��~`]~�%F���X�����]7�2Uc��lؖ��Ί�'�hU���w7A���!��+V4��}�S���˽]C�����(�t$��(��>9)2~��9�)v#ϭ�� ѳ�D��B����AqE-9"V�⻙ Ķ�g撠��΃'���y�09�ȿ�s>�[�=���ʴH���Y�&5��6�I�?�<�������֬aQ��I��j5ME��+�S�p��FU$(�w�hK�ft���&@����\G�2�c쿣G�3���S'<�%�FR�o1�e��Te�,M�4C�ٲ@P�IL��K����kjaT\D��1;�����f���b �*��e+6�
N��ߙw��۳	2L��>�OGrz�"�g����z�YV�kw�.��|WAM�=Ah_���
b�4����H�w���8����9�@��k�o�}��P����]���#�t��^ ~����y] $�a�R�>�(hM(����Y�r߶#3�w~r�����;�Mc@�h�A���Q."��>x�Ao�����C`�Cѓ�5l�Ca�7�e8zs1iRB5���M�#��D�\�V&ysʝ�:�e%��!-�$���n汘�5��숶D`@�az��}���rI���7�N����lH�u�_�������ʜ��ۧѬ���;�,f��t�{Lm����M�籨���-Kj�~�,���=
�f�u���rGm
F�����TA���k^�uf�_���u�LM�L�����*�Q�oe����2>U���,�j*�O�����\��]#L����3�4e��$c�>E��T1*Bfro4��H�ו���Q��=A�I���Q��!"r}����`��9���za��(����;���
��_���]�&����̗� ���O�Y���~n��[Nl��©��X��Ů���S~`�C�Xmx�$��Ã6?���ћz�2�{�`�$�||կN��.=�0(��������)m��2�6	�ܷ���KV!�(��݃f�P���pjY�8d?�B�H1��

�xE�n���=��e{L�^�H��k�a�Z���=P��M�$�P_�/��N}\	n��<�8�+�\J�M�Um��LRUыt����y�\��5���W���c�{ �0�.�aR�����Eڽ�i9�u�$��'Ӱ�{��� ⦷ȂѰ�5��l���;[�`�V�7&� ����@�\�W�+��W�H�+��UJUx���:'�J.��1�z����I��,��"�=��ؗ(f��Vɫ3�z����,��M��dp�~��ε�̻�<L�3s�OA^���@�|�pτB����Z��|���w�W���Ӑ��-J����N�(_�6�����8��;��6�b�y��������+�6����iN�T̺(�����|qn���}t-�5����KE�q|o��%�QK+�f�=<G�x:��^�S˕`]�ӯ�Q���Y�?]ݯ���O�C���m����οW׸���r�����钎��؏)x�@V��5X�bd�%��oʮC$S��@��/�7=�����{���5027n�0�7��n81K\҅q��p�`P���"[���A��V 1��W�U]��B���j���7�:����h�%>����0�ʆ��cr��=Q�E�c ��1i�g�h���u�
!!�H�B���[a+�����б�e��+6�J*r9E����(��1�R����L�잰�[P�ȳg?!}�����q��|?��"׀�Ŵ%ȱ���!����g�!>�~Xc�+(A&'E�p���v���pm��d#�Ps�a Iկ���|������kPJ�	ѕ�)���'���1�������[�/;_?lsz�LO�L_����ܱ�	���GM�5���8�U�;��~G�c�0Q�:���ߎ;�]?#0�j�*�Y8�R�d��0����t����I��U3�L�Y�Bo¾#pqܥ�,˳d��;��N��΋ub�x�����0�/]UؖZ�#a=:��|V��k���)2ѽ}���/�r}X;��%`�[�1̺I���cjd�Dj����� ��F*�Z!u�_�ӡ���"�D���Nd��`qy��XO�k��+���1TŴ�{�\��ԪT��3hL��-��8�D���=�+����e�$Uih|���:R����.����0��CpkY"�)�r)f!xK�,������<��pSB��Y����
UBj�]\���2��ԭ�����SwW��\���>Q��*����:�30҇F;���m��������>"fPBl�ɛ�ʪf��]�E�K)� ��U�m�ko��vMg�ۡ��T����Q�,��Uw�a7p���ֶ1��ܕ�=�l�Z-qR��️�my��7��(a���D�4���?����Z@.�3S��z����;m���2�vy�+a: pt'��Y�Yq�p��יִ+�`���{)�W�S�&�d- ���Sf�������I��6��נּ������_2�h|���Ib8挖��y�ݼ�){D���e
_��RIj/A���W�G�aC_�Ӧ��%�~KӅf����;I��c���t�c�G� R�%'2t	�P��q��Dq�e(͚���ǒd�ꨝi`��^a%����G�6����	�S_��O	�_1���29T��o��v�֏2�Q�y�P������GV�^S)Y	��^�Ak�Im�
�M4d\�$�~��nk��_���	�<�Kc~6���>�r��3,M���^���*x�M;����%��N�����ה%�Y�LW����,����|�Q/���Sw,\��Z�M1�N�="E[�M xR�MJs+�J�"U /��n��ǋ���W6zBזN�My��[���>*�1Ol.���lI�z(T���W����-
i���y+Rߤ���~mK�7�P���Q$U�]��5w��׳׫Y���,�ks��Cߠz7�M�����ǣ�t��j��H��^Cbk�OY�! Gb/���� v���`e��8���3d4�}G?ƥ�W������1Lm��oR�(ԫ�:��J����;���F �$��+*T^�Y3s��()w�`��Q�g��HA���̢��>s�By�@���a�@��C��#%m�?�MM���P:���y�������u�9+9�{���wS_����
�gֽ��gZ��ȹE!���hEabG�_�_�0�떌�e�.Y�zaA���/�c41@��k�6��jP���aBˏM����y���,F�U`Y��PE���Ś������@�C.RZ�S���"ɑ�X�$����3���� " �5��i�h��^[�9�	M��;)���p)�����'u�jgcZ� �����6���y8���Fy�����Z�I��5���Y)@�VW�~;��Tc�}��Hc#ۚ-B�L�L7>��fv���J�VG\jy=:���sk8On���z$��5���]�EAВ}ٯ�r|����[�7�v�P�Z��]�#��I^�
A�J���Qt7���m3�ky��XV�]�8����@��=���4#c� ��2s��h�>h�/{��qC(&���Ү־��6�Ҧ����Hp��e*3[���5����1{��;��]��Iئ���ۼ�u�On��y����6M@\Gb��*I�4���FWWn,Y7�����C������6@=��)���	`�5it�+��%0J�ȼ��bY���Q�W���whĘ���M
�dPCk��8b&�B_���e�b��=����]��g%0�5���ߠ�4'7���Ak*R��鲗����9@�g�?.��⿳|q�z�R9U��vR�a`�uK݁,{�}#b��Q�A�k��N��q3�K���@4����&T3`�T�[$z1N�Q�uěq�o�"$��/G�;Q����m-ʀ>��%QJ�m�0�Ƙ�x�/H�#;k��i'�a��ލ�䨄!�4A��C���f��Q�f��3�@�!�d_�m2���,~������}��OG�
����&���X��\��7�"j�'ι��PCT�0�ြ���>�%�)���c�F�RQH������rY~��%��3�땵Z�;`'v^Κlx_ �GM"��i���s�:��_�yS]|}f0��������W{V������5K�p*�s��U��oM�ek>����0��'�'��l>>,�8Oj؊g;�=�B���dY|s�d�DW�B�q�NL����2��@��sd���HƑ����Y調 �dFYw����1�ux�寿�Sk�kb;�,$�P=A�ܩL���x�97�9%J�C� �Y-p�|rOvR���,'�ͦ�B7�7{��	'm�~D#����u*{{��M�/�����F����s!�~�i=�D�i����R�;H��S����K�:���1~R���n��ִ���H���S��í�Q��3{��^��,�A9�)�|��a��U�`�w�:�tP��U�W�X<����k������Q�*�)�W�XU?ӛ^h|6@F!;ö�a4 IT!qC�ԉ@���H��i�#��ژ[���y�G3�I_��0��ª���W�0?�`$�%$�?4���f���]��5�U�Q�k�ZL�� �V��`?y��".7b����)�|��z��*�	(i���E����;���!f+� �%��?���|��FyQnI���눹�XʴU�p�Dy;	M��M��Ƃ���|�JUׅ��J����f�4��㬭��:��"�c79'U-��s�;����� 6f�f�]](И)��b��Ӹ�d���+c�Q����mt��d�[e&kl��`���)���y��� �qH�W0E�M4���Q���N��۳��Rړ����6��S��!�0�SW�
^���K�i%�9���%�
r�'1f��bMNc��7�b��1���Xa`�G�G�X�S_PkWj�l95��D$/�3��� ]��6o{vmY�>2B�x_��7ڇ�g�w2�sU�:�O�<+����c����r�%���?jP�{vp�_9��9,��I
/m�s��M4�F|i�Jx��f;b��г#&������-���B� �Ǟ���|�K`�0��l�=����6�����.x�?��6��1�A4�����I�w�I��
j��B^�7��09�Y��.X~�D��~�v��ї.]�x"t䛘�����S�"S�m'�<s28�f[pnի%nռ���5ޠ�+w*����6�XBtؽ�T�ծκ�>l=�v�ru������~��{���(�J�w��4؜��H/���g�܊s�5���#R�෴֔�P/��m��\�~u58͟��"�t� ��҅w������>�z�:hL��\OuS���ʸ�Ɏ�3 �r^����#�qx���]���o�`�����>�2]¼�ea�6���8�)@ZO�i��e�i�3���# ػH��D���qq��X6���i/��k�%ׂܵu����S{�K�0�B(f��[���TK>A����:�P�
�v��6�*�obn�������k