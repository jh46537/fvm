��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<a�J��Z���=U�5e�h1��=~kY��b�6���a5��M8摞�
B�F�Ԅ3_�̜H� �Y�~�
��yuY��̾��6�E%�6M��m�B�e�v�Aѝ8
E��&��G�f���o	�K�+�:�'V
Y|����:nt�ӿȉ���`؊�\�v��Xr��$�<�$�	�'P�~e�_��V�,�#GyP���(9tК(�p]����m���hw��=��
��;��������^�!�X��Ċ0�ͥ��2)�����d ��tK�g����t�K��o�1�6E���QT�]aKQ��e��Ր��j<�{�g�e��ČB3�7�,�^��}��gԩ��������#)w&!���0���}Yg��w���y��d�SPk�拼��}���p����3��G�*2h�/�s���zyx��G��
�~��;B9�D�7|י����E��`&�����I>�=e����2u��;��j��@Upkξ�*6\���7a��"_k�������i�G�cJl~��bF��I^8x�c�ŅW��ɚ�t��A-��x��$M�N"2�'@�N\��̀��+���e��gcY����3.�E�wSBhX����P>�[>���L�ZA��Bx��"m��X�r�-�nw�J�v�3�L^���c��(�������{6E���T:�����&�	��O�J�B8]���D�|a�:�d��a�ߕ�n��x�����Bku�sZ52��ϫE���k�NG��LT�Tm� [�v�+�N��a×��ee���ivW�N���jL�
�GYA�S�ѯb+iJ��./�)����!�;M�{�V�p�$X��� 2���	�U�@��@W�ޘY�m�O���7��Ug!m���  Zо0fM�p>Q�����E����� �N�%��.ޔ�Rs2�ujIuB���=ʯHH�BV�k�j"�rp����E�Ϥ9���١����������9?�����G&ۃ��Ci�	��t�dY~����"-ϠP�-*ZN�,�
�`�zQ(��V*@���~;���.#���V�{5��,kՅh�G�Nw��S�ag�T�)��@��J���j�����䱚�e�)Cr�=.(�4��5̈R��w�),
ȿ�k� �3��3sWt�.$�N��B`���]��ί��s9�P�o�H�K�	3����_[��#m��v�W��Ӗ's�ʑ�}��t��-6j	��r$�,a��!�'o���)���v0�z�O���U�A���2M�+�Ͼ�j�l/�!�L©����$�|=�����~�ٳ���"V����)� pA�N䗨$�j����1����x-:�8e����kG�¯^�y���c����_Oהvw�AL���Vy���l ���W舛jsJx����[�V���!���Q�8Y0|-���Gi�>P�f�ѯ�ob�|�O ΐ��$a^+�_Ħ!
a,Zb��K�;�O؛�3�����i���<w�u���.=�3�c�k�����"G�q��1t�>�����i�K��W�����'���
��i�ә�cJ(>�'�@� �u�UxFe�B"m���� �_��͜�G�L�E��h�:7�Y��2�XF���Yda���o�(��mF��}�4��i���A�S�N�XYj��� 6� �i
>]X�Au|�]p` 'COT�١���5���ҟuA!��޻�u��s�R�����FE��So���݉k:i�5�\Äy^X5Ч�,���D�X47���]�)�z�*ӬwY�RWq���#����b���h�m:���'�zL���MDM͕KtWB�W�=��\b�<vpo�B�������a!� 3�|�#�Gю+�0��N���4_����&-�T��:G�L�g�IA��z6b�-�E��?��vW����F0��$�� #��4��ЄaN��?w��Ӻ�v��>!�j60^�j�Y�(.V���%����[#��	�l�+w"j�ب '�٠��m?��<�G��K�ɤ,-9eBS\ǐ�-H�p���E	���P�PEb�V���}bҖ"3jW�,er��P���>���YSw�SZ$�U��
�i,V]̹[�������G��v�VcS5�mU����Q.�gC���%l�xC��>�#m�yg�"�~�~ D\��FE:��|w��#�k�Jɴ|����0��"��t4�4k�i����դ"e).J�Z��'XXP�ǍM<\�HS� �����#�G�HM��2�Gג���%�ش�#]������\��[��4������ӧl�mN��b)��s�"d�e��4�<"�G`���GC;w3�t���7fIA[*G�TY���9���<�Y��Q,{a/a#뤙�Ut�j�(8��6P�dKm?S m��2?�]�V��=�� 0���O��/�<�#>>�P�}⡰��Һ;J��*��*�x}�ɚ`�ǌ�̎���'��<�4u��"�'5OWU�[�k
	x)K��ᢋ��ڈ*�A>��F�`���مZ��or��K�l�`�s�!+���V-gZh�mHK�}�g�j�JC�祥VC����u�5��Go��Y�4G�L��go�h�$U�;܈V%+P��v�r*�!��/����m�e�t������TIC�Q�U��$� -p:5.�)P�4���вn"[�&x]XKAJB��_�b?�u'#�V"�#�M���;�r�ӊ�x4�a����^����j:Q�~�-֊z�|*x3��Ŵr�R�W������[ �/�<�M��ΌN}3�R��7�>��7��u�}e8N�EC.�C*bG{h�8�.
��!K^󾝍7/��k(�UK�_*e�-�H�L5�% Ѧ���}aB�sz�J�^?^i������m��-�߻r�[�2� %�a���17-�QTi�#
�w�]�v�'���m������Jts�~d)��{��^҇;�k��j�2�/*!Wǜbсr��P��^'3͖`6@Cq�,��"��bڂea��?��%tm�S�wK�A��1Y������^\�.�u� Q�̱��1��i�I̠Zp���Ѝ�z���U5v���J�[l�7��Ku�aF�w^��e�=��5���&ĴQ���91�"s�s�+��ӂGFW�W�|�OMu:*g2m�3}������4O��p���X�˫����G�PRg�N�*f��ͦ�.4�֢yʗ$"��~��L�码�aqH�Ѽ"`�%i�.)����,��&QU��'o�\�\(�i�|r:J�����6�T	>Bٻ���p���-9\.�*/ڍi�w�� fP&�ڠs�s���NauPK#�>:��d�m����R{�&l`69�@:���v>3Ԕ5�/�em��©"�dd2�W|+\5�BoE8�ׅ[��$���C�D��&@]J56��tKG�����t�V*�C"�u ����YrՉ�/�=Y
�1/C�QЬD�~}¿��ܲU��ⳖSI�<0V:y��"<���ՔN4ۊL��n�֞<gR���2�����Q��6J�Aʤ�qbt�R�ܺ�(�%���h�.5͋b����v5�����c"%8��Bry-�0����܄�mu��b{��nǜ��F�m�*�Zw| ;��7�-8�*9LQ5_��*u���3+2�tp�챨���,�U��LP����li�u^���'�3�56�������IR�Z�� &;�œ��O�����F3-TBn�'&��>d�ڶܙ���#X
M\\V�tx�������a|���^�����@�&ڿ��A��u?�:2`/w3��ol���z��1 �\3� ���Y`������u4=>�0~`�ɔ	KS*p�Ro��; "������䉄���!����kGhʫ�ۖ��dRdg"'s@Z��<�8��HOa֐�b�����޴�,����[���9�&U�"�;�b��%3�1�U��װ�x6x,u�^@����&�b��[��˂}��"Z��~�����"�|� 1d5(%�L�? J;�\2��|�
�]�*�d��r0����54��j�a��|L3�C�"���w��6�H�]u�0��'nLV��/�{��N��B;U�<� ����I�uj�u�DV�>Kt�
�w����Z�Lc���*k�jBA?C�xj`^Q�H�G��ݥ�xT�ATH�(��v�?�Z�NI��\���ns'�ߌ�)%:U3��XD@�f7Wd7���}��˾�0�K��q!�C��M�p���D}�\�K�Qb֎W��M��~�F	d��b��i�g�.�ɑ��u�)䲅a�Hy�9&��ӳnZ�4^.@��v_�[$���|��l�;�M_Cfb>H䪭f´	�1���L��#v�&r"J�?����E�'!�N�=���4�[�"�.`���gRWLE����PB�m](\�l�E6��~���`��J,HA� ���^`��=P�y�r�'�ur�қn��(`ezِw�Y̅Lw3��� �'�!5�ʥ$��?���E�~�CB�Ӫv�1���?�<�̫���yYL(=Ύ�H`���Ey�:�^�V4{9�X�]P��h�u��˵5f���h��b��;�/�L'Q�u3ng/����%�9�oka��^�>���d�H�}X�܇;m��g���t��ا�f�n�H�+��ǒ��N����6��q?J�-�(���)�fK�Wd��.5npc�7����S�ra�xn�� �_���Be�LR��|]����1����q9aY�k��S��i�y���7ȼ��0r�o\�9�x�̉�Ћ��T�?eipw�0�-\��Nޥ{��B"�$��%���Խ�h��$�9p�hL��t���K!q�`;���]�g�5K�^yY���~�V��^R;�G��~�>R�1��?��?Y��;0%\<����x�G.���r�ݭ�p�+Z�81Ƌ�G�֋������O���v~$��tG�� ߺR�0�'��K��G/�R��e�;C��A�Gg��X�G����t� K�S	N��	D�w�y���>�>���VG����5ӝi_Q�|7~��QPn�o7�a��\��.�8��e˼;_���k�%���$��(A�j����tI+�9�f���+Z	�'s܌�m��v&%�&�O�b��}MÊ?�����%�5o �J�B��+������jd�H�S���cw���6/��F���S��%��0�Ɖy#q�%N/>>��4S����;��ËR4��S��Ϲ.���Jq*
kU1�r�"2*�Z���ގ����:6}`���2l$%Nu[�Z�!��m��jp��8�F�^�S��(�%�B������w4����	�~ ;$�J�NMOe���k	8Z��cS\ҥ���W�X�"�[/�ZI ��A7���6�̀-�t/���f}�Vo��)/;ӡuP����{����*�ZDq�,�S�a"��O���OL�Y�[���!��r(r8W��Sq��2�n@O�H�*�r9�����p+�k���$y���?��-~��F��@Y��3��G��e���	�w�b���E�G�zMf(�Li����9N��Do+i�>��č���z@�C��>���Leвf��$�4��Ol��jL�)L��.s�d�M�?.�s6���\ � -�
x_�������{�d���q��B �?�z|����NT�U�E�Cq�h<W=����G�J���\��b�)��X��O�|^�(s�X��%;��J�Yn����W�f�&^�~��,�:�/�F�A	����ܵ��4�0��Qp*���iK�Q�7H��f+���|�%p���m�(i���56�]���٭�<�Ͳ����w�f��k��}ۺ��")�}5�`�hvb<�}�W�F�]��r$��?�E-���Xr�G����l��VY��ޔV�c]��6�>����	�����檣@�'6��i�J�
�LF1��a	[��az�s�X��6�-9\�Ǘ���W���o��2~2ɔ�h�K��s�[��),80/#�Oָ��b�yzI�[��}
�um���鳫Ip.[Fd�*bύzv{bd�=�������e��O��qi�f86��bי�����ޚ��s��'[%�.?�
�ξ�c׻	��f%\h������g������:w��*vB�"^�@������<X7�Ђ]t��C�>��0�%��p�'����V|nE�j)ik�#We���4kt��-�f���p׀<W�B�jwFV�\A�������9�3f�"�Rbc�4�k|3kޠ--f�Q�!�G����i�d�:��:]{�޴)C
�e|��a���@�B��0�X}���y���[O�ku���}������'��#`�bد�!��_K����SD�\�<Qdhi¤�r�E�̠�+e�FS��p��h�:o����LQ(q>��`��|@P���Cgt�k���8�\ab�4���'��I08`��
�ҷ�����=8iC����zޡ��'��o���6���=]Iw�R\}�1��`�úQ�&�ˠ�S>,�%��0/J̋�.���fVՁ��cR���6]}:g�IK��A|]���9*o�f��Y7�+�)��v��s� �Ȕ��m8g�D���N5f:��� @��M�oI�a�����h��S�����o �j�#80���:A��9 �=�B}*�B��	��96�<϶�"�� �+^�P.g�9��9��6Ȟ�.(�����L�/K^�A_I�8y��T���h�����J&MM��>�|��CV��K�������}ƛ�@�=�:�c�i1��ɋxy����<û3�,�����&ve��	�\��t��J���L*yY?���30M�KT9����Z�q�V?E����'���$� �0:pt9$�9v���p��@=M+pj
̆D#�*�Z�&/����m���=������k"�iC7���X�;��]�A�{��7�f8)n`����P��@��?��s;[%́k�>������R%�֭x@K��G~\:������4��U�sXz��`�i^5�� �j���Լ����@Q�G͔��%P���3�s�`8�hW���x�X���W�b�a��(]w��!��6�8���!/���~!��^`�4�Ƀ1�ĤƢ����D����o8'�q�Й�z�â�M�C@O^��ѩ��ǷN���cx^�1�B�U�E�� 9��g��i�d�L��q���B��� M�<U�L���$�Uค��N��)@�W��1ج�"��6�7mTO���>a���r)��lo|	z<ׅ(�}�`���ķjY��{=�
���_Ǡ����6�&��v�SH���D~a�>:#<�m�NH׊M����
���KtBb��P�/vkl{�aX���%W���ؕ��ZEF��t�y��� U�IZ�f�iH�G����)H蠣.6{�@ �ږJYQ$c�5��N�=(q/���kG�)�-g8�g�0G���e�%��_������lB�t8ၧ�n/�-��3������H���r�����mP�Rg⓽6jeV�) ���M�F���b}�����uٙ�u�爩=l����U!�-B�ĬT�Ʉ�a����Z;��a��X�_c�U��ӏ�=G���f��Z�����+S7'v{#��P}��4Sc���c�p�ZH�']Z��/��y!FH~9U�\~���QX����[����K �|�"�}�;�D<�͍�l�>�
�F4�^�����i��)��J��1c�/�@ʗ͉��`�7X�(�,^wd�TXo����������/���K_�@���;�b*Fec���8� �W\�!�Q�D�uGh��� ⋺�j)�t�C^i��^��8�
�yH���{ui%^r�%%������I	�Օ/?!f��P�U+�6��$!K"���#�`��8�����7`Y�.��1�bW�_�"�L˄C�Λ&��U�f���/p"5��D���L;�D��1���5��-��7)yj�XD��Yo���]�L6bգb�� �����2��=�t��7(c����
&�~�7�w�f(�x�����N��еF�50%���w�p_����j$��9�aޘБeŌ�&��J�1�:U�"���*�K�2)���l+&X1*����"3\�hK1�~���m�J�M�l*/&Q�J�����+� �|�*�p1������.q_�Yx������۽G\,F�;:���u��Y>��f� ��4��Բ����0=6���Z���)r%	�&7꒶a=���$,�q�������M>�) |L�b�7M�8	E�d:�&�>�/��or�¢zi�'fQ��7��e��z���3�j����a�m0�/�	�[��,0$k�/M<n!
�L������V�C!�u���Dk��n�OB^�(�U\Y9A�,"�܋\�����4հ��wˋ�! �w��"�-)��X��C�� B�Wn�;��5���}��HĆ��)�򗭿oD
��ြ�~s��k���F����Au���s�r����,��%��Ԛ�1�[��F���  4�uqW_9���mj�'�K]O��gM���#������V+�p
r@�f�qYo����Yp^H!yj5z�Qb��`"|,�	5zݾ�$t2��|�A�w�K�TȠ�n�3�lb:lO��s`#9���+*6^�b��F�1�\):Fuɑ���E�[��M��y�&H)��P�jP���bg��5��v��<�q=�pY���i�Z	��K���H��P��i/K��4U���,�����*��b��,RO�����_�P�⪉������do��#5�Mf����z����2��N_�aa�B��Ɏn�@OY���n���>S������fm ����̨�erbSo9���j��_�]�_f�1>�ۓSZ@�r�Ȣv���zm�b!a lZ��)�D�
*�z�0LJ��w&p	�%��6�����!9K,S��}�y����5}��}̭�MN������*���Me:q@��}��ּQ;��g�D���z3�8V���m�3p�V�����;��p���]E�2C�NaB�4�4����#T�T�nOxs7�+T�y�h_LnBݓ�O=5̾|���3X�&wM��	�K;�,>���S����)��{}�u�'�:��3[)L�Gh�h����Q��7�~�3D� >8C�4tQ���l�R�xd'{ba̓���4Ʊ�$=N�^���5s�~o�M���������Z���Sn��n�hL#���t����g�����g0/���^���jTf��۽���D�� �׸��<�]�/�(; ������ȥs�� C�W7+��A��&;@(�@K�NE�HjH�S�Ǽ$R��'(���6L�M��@u�~l��4v��&w$������{�}��䛧�r��S�al.�I���opE�AA؏�����yo�cǡcK�fu������Tq5jXI�a���;Ԁ{_��;	 �ݴ�bk�Y���5K$�2	��D6��č��0�B�VR�����1�6�=�7�,}���c��p�u�(C��;������[�h?����x��V���;W�)L6�爍��E)Ͳ��#E��;@��V�1u�36H`��؅aa �`Mŉ�=݆��2�T�Ŭ4M�Ɍf�*qZ�X~V
Ĝ�"�i���f��v��pDJo�J�Zqھ��. Tfx��HW�!����6��c.vY����P�����p��e��j���F�ʣE:z3c#���*���ǉ��kU��\�E�U����V&(��M[63k4��-�5^^�'t˽�*���";�b넨q�Z�3��G���^�����g�����)I ٪k2"��smѹ#%Nk�D��V�[j&lD��"@#O>/v���aU��U�	��օ�Z��N_(�]�:�w����;��:�U{����Y�d���b�Sq-Sh=L���t�]��_�(���:χ�s#{gVo��Į���Qn��&��_;r� vS�x'{u3s����[`�on��DQ�tgék�>��a��W��^�;J�实f:l�ᓮNF����ĩ8@�S=A"I���v������h��xˤw,	�����KI���z�Ć����[�F�N	��];	�ٴt�	OT!3W:<Bu�R벭`0�mk�>�f߄�8g���������'��Z+Q�c�{��� 4��c'��Ŵ�`�<��$����cN�pR�KW�B��JP�UW�7+�i�4}j��w�s�r9\�[Fv=~���I%p�Y�^߇Q�H��o2�JD��7��h�����Z�%�)�G��5撪�DP���˅�?��o��;��f�C��MTѵ��@ݏ�78�gC�DJ�\��$�U�
ҙc�;�Ҽ��]#|\pbp6'�*"dxY�h�Vm��p�L����C�Q|�	�.� \���q���E�vkka��`���\�G�Rl���6��Ǎ���R�z�'��d+��0��ϼ��!`!Mi�� }>�[z�q=�[h�%]�O<�&���f�æ:�������$V�$+�0`�ę{ʳ� ����~�0v ��Lց������Fđ|�`i6������'`I�A
]=d=�IU�Z�a��"�l4V��J�-��J�BS�wF���eMU̐�uv�O� ���Z�sG5x8��,���H��o1z6�'?|��Ɵ���N�g�eaq����^=o����)HO��յ{�A�A��2��t8�&�.�C󘆪�;�]4A�ɛ���o-h?�Ӓ�̨f�΃�ڝh2E\�wz�C�@
;#�lI��#�Os�������w��BT`Q	�~�G���1�AgZF`S�an�Ϊ�M�4'wf��s�0�%ӮZ����'R_ZUyU�|)'X�����K5��MYƤN��r�+����,�\N$(�q�.i0b���q�f��&q���q�U��Si��)��^��l�+
1�AfU2��n�i�"��r\.��3-׻� ��|ʠ���b�~�M/8���gIY�t���ͦTԉۖ{��m����ּ)Vp�Jz���ct��.�,K����gNQ�$���I7U��P��)�O����Ibfo��x�KK`���L�Ww����4��P�葅	�7<��x������I4=K#�K_�"B���y�@<�O]i�K���̽~Z��Tq(�����D]��*X_����]m�Ê��ZM�L���S .^�DԆ�ɖr��DD���sUdŒ^X��E��M.��R6K+�A)��W���X0ې��d������~��9*�H��i8���
~���.���'�׶�����{ivҠ�y��W+]�
������*�?yI�5�(�ٴ�B-�� ܪ�MZU���IV'Q��e��_˾X�͏{���+m��5�$����|�ngL�7�i9�P��D���b�\�I=�`�5֩����jT�`UL?�Y�r�,D9�t�ݰ�O��L�m^.3<��gC�$�N�o��BD\}��oAX��PK'sA{�S��f�.�+rۚl�d�(��F��L�R�N���w��9���#��\�\�t���e��EV$6���?�u�c��!���vfw����c��p��1S�0
&Q�ef�t��kX
a�����!v�0�S��K�B��SU0igV��/K3���rl��s��C��UDQ@�,���L��==`�����Z�jH� �YMU�:���r1��\�鼴��d&�ߘB��tzO\�ZQ*����T-�pi�`oq����G'c#����4��f�(3U�ɸT���`���zB�����`NCcj�ճ�cG��Z������
�:KyJE?
�	s��|j���7_���X�w�$,�+�q�+�'�D�O
���	Q���\���F5�N�����!��JN�A!C{:ݧ&�u�s��� m�:��N#���/v����x��wX��Зf��$+�,G��٧_�������5[݋����)��f����"����yXR��Gb�q�87 ����5t�Cŝ1���6(/M����$�ݶ���I�����L`�lW.��h:D��?c}ZU;�>���tb���"��d?��Y�\��c!	���JH�~$��+>FWI���o����I�}W��oy���m�4v�2�Zb
���M�`���zY���}��vv0.���Ѷ=F�8��󦖙#�EpV}�٥�!�Ph��/��&������PL�
�x�Jbۿ 骆+���'�J�}�m,�'y-`�ԛi�%��O��q�K9
[ʅϷ��j��������c}�6D1E��S|��z��?�s'�� �?}Vɲ��2�풬Rt�b�0)9�O�{�r��d���19������l�2�Bo�P����twt��@��*M1�S&�v��I;FL18�|�b���rVE��uV�|!��d3ErA*m��u)��Ο�WL���!�=�3
u�f��}QB'�x�~t4���3��q�wMF�,A�3c�L��6�vnզ�X���'3�D\T��;��T��'��T���I�YV{}N�g5T�8�ǝg�4������X��(-7rY:���u0�1�98�:���	!+S����U���_0��Z��W���0G�z��QϦ���v�/P�7B6�!�tt
t��U��R�f�eZ��� br^��%��0p{Bo��6�Hh���8@�'�X~�C��F\�ջ�73l��#�����=LS_��S�z������\�,,p��+;n�Gx��Lr.H�V2P�T�c�����;X��],�wi�@xv���<~ؠЦ錩��ڽ_Cش�D��T��o2uHdl���@�0$ʁg���\:��гp ��G49*P�^>Y۰𺶉E������K$�g�L&|�۹�ɀV��dB����8=�s�I�7�Ҁ��B�`⟯Dn�D������m�Zq�Ld���n����'�ɤk��NZܨ�����͓�;T;�}ϝ�]�c��H9��);O��Rb�'{�dt\*��%��4��C\}_�N�E������'�~񺪥Aٛf&���tȑ�r!�ay�|��0�<2��5��{����ܴ|��һ�Q/����ߘ"k�2��Q�<�Z���5�n��Y�F�yz6�&�����ع��k*�!�A��f;z����ξN��{�HOq���FQ ��r��&y�y��
1�~Iu~oQt��}齥�Pս�<L����p���.]�GF��a���6[¹���_3A��y�O��u� M��'�uvɬBt��ͣ)4��v�@,�nmB�t.h��U�g�]������c�%Ȃ��R�>F���F�5; '�MQ F����vr����C�
YaH��Ж��rU�����ز"��eNF�DJ�=eBGm3fۇ�>�2��c�p��c����C���ɐ�4�`�)���"&;���\w����7/����������\΍�y�`��a_�|bD�7�S@��_3�%��[7��4Q�TH��͎��+]�	Mo� e�{�pS�߀�J�$��c���ȭ��9�s��/l>h���V}W���RB�Z퉯a'LW]b���6=$r��o�'Z�"�#��i�I�BH����\z� /�O�;+��FY�$s���c901Yڭ�ه��֭2��65�V8�&����8_9s9�/��{�\�I�V2T�t��E�UP�P��'p悐��RUr�3	�E���[2�G��'ŌL������@׫x��9�i'f	#z�k0��b7G��^Jw�5�ЫR<R�TN�V��/#�6�p%�2�S�I�3�5A>����鈮Dߡ����.ӧA�`���l��6�Ed�1;a�vXL3hF�u��kt�
z�����}L%��¥�c�/7��W�'lI������SXyl���8�"����~��y/��h��J�d�4�����ќ␙˒)�"uV� )����� �_�J (�۝F��~��9֤�B��8��P�T���+J.�*( &��F�.|���'���E��D5��E�"=���������G�E�5����.��gJ~�d����Xnf��I��x�x��d(B�泍T�e�C�3����Q�G)kjT׈�*2���`3���#��WE��O���YBO5W���u�����Nn*[��&R5�.vw���
�bv��\�݆�@����j'�=(�;4ӍD�