��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���q��՛������@�oa�R��Iz1A�#`�ԀP��Iqh�3��F�`�ҥ����c�
K4#����ge��T5��G�z�4��R��\3jU�;Ѫ.Xq��d���D��nmac��V�ܕ�;�)=�(?0�י+�k�襮=�%�YO������鏷w��>�s]��6�t�u�;]��4���!����q��
1�xF!b������.����\�2�X���`���~���4�k2Y�a�w�7=�E�u��#��_f�g�:�S|.�� �֞/^���J���,\*��p�#�0k�|
]c(��7��ȩ�'�Q�	�kR-`~���Zk8�$'��x��A1����Ko�� _'-l_���\��
+*�q�k�����V�LZ\?rŮ5�xwpP�V�22m��w�j�{!��;�Fs����]U�ӂt0���� �d��l�F)2+!}�]�RB�7��ɰT�O����"g�yl�����y��b�V����!c?3�4��������%TD�������)F�p�8�DcKD�Z��f�X��,�EK����:gY����/0��E!ѡ���mr����g*��M��H\"_�R�P����'0x���YJ��Ȕb��Fd�%^�H����&/Z��,3�׷��?��"3�׆��$X�����G�"��_P��	C^-�6�s�T�X�j��p�i'�:c���
����.g�<(��-�*�~�0p��ɽk"�;��ɒ�]�x|{�6��xbu������)LO�̛̚�U�3��o�ޣ�U�D86��iN=oq�m Ѧug�p?�y��)�o��$G����?7��3āh�s�J1+�m�+�g���t{�s��,��K�NZj�PG}ܴ��Gp w+2�W~��9uT���{c�
�ķ&��2J���\^J�XS�V�¢��1$hJ1�L��Z���'�����!oD�1^V�S��t��l����s��Ӫ���
Y��re�H�8A���W��#(����?4,u��$'8\d.������Q;������@��n���O������V#�(�(�0*�n����j@H׍�3d�i�A?*݂ Q&�T���X���В�̟y��	�#n�e�'�I @t�Q�rU^D	R8{�~�mX�C�*1��O�0����2՝�.+K�g��5O�j�[Ͻ� ��\R�1���Z͝��b�ʞ h��5�"�������3��<76�p��)\x�JQ�C�<��u�w������G�0Ɗ�Ӈ�%�Ťe���`BhF�d0�HeuV�8��8Ξ�؏�b:�<��Xg�E��"Vڪ�_����Ħ��y���}M&˼�|�8$�4�$t~�Qw�]��7Ɏ2;r��,)����I�)R�?˖��J�3�K��2pĵ��)�]Z��N�]}S�hâ9�U����]hQ7>9���[Ffψ[���,���\��w�G��'��h']s�;�x�u�%R�'N�їx��,ME3�8�Wַ�����/�E��
�����X�����Z@s"AH4Qq�5�\���槪>p�1�q��}�E|Q���Un�mY�����H�R�(Ԍ�����~j�sYx��|-����顗t�C��� ��R��}{t�~�n����_�Rv�AY��P.��RiO���~=eRE5V5@�ƢK�>�LK}��&
�K���	b��3_q0F,���$$	�6�ܜ��=�֪��$;����HJxX������%����k+��iW��>��V�P���.�m�E%�e��YqZB(}��
�7L!�,e�n�
Q	��K��2"��0ۮ�RGGQ�b��%�r�\O��u����J���gs�cK��'g^;c�-m�#`L���`"2�i%s$ݍ ���b�ptBiH
Mx��|�SL�sqS�F�fY�ӳ��^�(�o'0�
��}�8�O���LC�,]�09���,��t�%�nMlG[GW�
l3�0��FX��1�[7C��T�F�?�aU���0_�7���3|$M��\g�o`y��Ʃ�3�+�S���"���wW������\��CM@x��uH��>�׆B�ɿmǷ��?O$h��s<���JL����6u>?L�T`3��������|����#��t�'�OA��W:�4Ķ��C�J����K���q���6���_):_B�UŻ�����cg�<.?;}�^Y�<�8�z�Ɍ� {��4b��hC݈`��
����hY�x��4c��"o$`%o���������-n��NwC�:_��/�{}Ul=U��L7���pr�.�1Vo�$�`���h�>Ǳta��jp���`���2�UHxLX����y�,��0�Њ�=F����8_��]J��啹(����G�佀!9��>�0U�D�l���/[֗Y���SPw\�^�/�G��q�;к$y���D7ֱBu|�U)H�fޅ����_�Wݤ����������Q��+�-�gﺄh��}w�������g*�u���d;|�k��5|�6����Z�����!.�G!�#�"B�&�A @ӲJr�i�bu��!�~{>��<rr#�Xγ��iXZC�̇�l�r���䎬ji�ϖl� �>:#�2�>���~�ʈ<H�R��.˛�r��UCnCw�U�����2g��(�-t�K�@�f��[i>�ǘ/;�ۘi�@�A�t�n�`�EQw��kh�F8�T(�ݘ}l&Q"��6X��!���'��_zT���T"f@����@�6p��D���5�%�@L�[.SmD����R jR��!���C]k�X�%|,\@��M�J�`(m,�Ww=���I���%;�aosC'+~��hN^�sȩ�|=]�c�9�A�~a��`�sT�)x�.�ň󺣨�3�J�\Sq�������O��-�A)��k�q-�DAu@&'s�q� A�&k��sC��9��_=�5���xcă���t��&�Y��Y��"����S��$��%*�2������$�i��?�R?��3,��Sj��%���Kzߺ���# 1ѹh����%�K�awK�\ѫ�w��W5N�џ4���� E!��������"��������K`׮%�L��n�t+.($���.o���.��� ��a��[���f �Q	���_HJ�t�]{/�]r�F�;��J�Cg#�=�[?$���B�Q� �^�<*Ss���nij�&(��ul���� �^��n����pN �N���!r=.'o�y�b+c��:%{������+Zl��r���Բ�#��H�S���ح8����H��~�ۿ@;�U=j.�ݶ	�����4�������z|�B9���Q�%��e=XW���ڡ��vRb��`}��������L�'m\N�l'`�A�=P]	�`o�g;�f��� u��R���b��h�J�}=Y ��B�m�j�,i5+Ť�����fԹ�0��"���Ÿ|��EIų%�g�U�� *��tX�K�K�O=L�<�|�L� X��g���0��n��.�iv�j�ѸZd�=�wԞ�L�J�]!�Yc�]��a8�#�����]o>}��a�b}4}#��7܆ǛH
���;�#&��ͭ�ci�I����m����9�=��'T����wli)��7���s az�R���5)`wO$�KԱ�]��
�6���G��=i��rVm��@g"�-�̦є=�4ڐeg�N��X]���*\����K�k*��9����?�<��gJ�(@K�� ^�P�Q����u �Y��M���ٓ��&�W�����ی6�0��}��}#���8���+31�
���'��4�Z%�Cmu����	v�K~w�
Ʋ\�*�6�{$�.����/_�Li@l��	wP�����SS���e�k�,���!��rwH�jSwP��[�y@�;Z��	���`/>�(��v�uG�zK�	b�n�ཀt+�"�*���� y����[I�Я�,��������?tu���"�4Q�F�NT��I犢�1�85aG
��2��q`�G��S�hB�&������nr�j����҆!�p��Y��1j7f�W����ۣ����}CCqlЮ��Q��7wf8��1�����g-!��ʎ��,(5S[���ߖ!���Z\NJ�\}����u[s!1��ԧ��&��씱r���S�!�����e�3��/w�^q�].N�P�=��:��h4$��M�)���ܻ���0I�Gg Zf�B� ׳n����Y����W�?�s��-�|�C��M�
%�H���_�O%�M�Md͉�$������1.�B_��<���w���Ʊ��V=�e���G\�21�p���ı��KD��'��%aga�g�(��P�MÚ���1ot�d���x�z��o���	�7��	 A�u>�������<���l�~܂���w�p$���NB�Z5&8�#�$�������褹���\X!�O���)�R�NR[%{���F0ox72�QvB��;O\A�!`��[GJR�`b�-_G%o�J�,ݪ�61iL�{McM���}�A]�嗇m�*�{��"�1��\��c��s���n�K[M��E_�������Ϻ�_0�!�����0���ɏ{��T��eΖ�e�Yh�&VD�>J9m�?<��.�57T-ҮΓm�
ei_c)=6�`EJU��Ԑ�M�on�b�׃�˯J `Z�P�J"�|:�UiA�tɼ�~m#��J?w�+0��A"Ԛ%mظ0ܩh�Ɏ�g(���d�Q��C��$ ����`��ބNT7�~&�ؼү��ܨ�,�O��v�0�gDKQ�V���Шj6�夆�
6s�-����-_	�N��m�G����]�G�=	���3
��6s��
|�2���vo3GL*Y�ɢJ�����T!�P�Kf���ià����y���rEQ"l(��cC����0v��aGQ�JkjԀ����:�Y��9�$\�B]�}��j^q�;kg�ƙ[��uM�2�7^�:P�P�Пg0з�[6È�#K�xa�d�B�)�8�=k[-U�L�e��\�V��Dp����lIY�mF)��ֈ�;V<>U/H+|��B�QEO�)��~�N��4�UYy �綘ƨ�2�"j`$�0r �k�U�H��Ỷ�DQ
|�+�t��G��5A�<f��}���Dm�P!`F�?��ʡ���A�߾�x3l��Գꀍ��+�P�]Yѧ�D.�E�-��u���΢O1ϑ���[��8�F�ϗ������c�[�A1���
#��h���{B�����>�X��"��Ԣ��V9krf�ޓ�N���5�	��H�?ə�={��%��x�Pl�*�+�'3�&�jh�� ==�&>[�SQ�_JҼY1i�_�����%�c� �1F>�ϭ���W���i�� F���Q|�c�����B 	��0h[w�e�$�t�����j���B�Žh�}f����Ǝ�N��X��]	}��^S���E(���h���x~�A���s�,�� �>��wR+j��Ձ� tK&��5j��PuiS��D�Y�Pu���	��l���/N[f��^��{�nU�`������(�C��6iZ ��@]5�3i�W��K��C��7��7b5`>,e�k<�w���@�0��l�ʸ���������^�� ����מmX���KG3nD�L�YlN�������6DG�YT�L^Tm��x���l��E��BCeg�g��Ǟz�Է��"!����d��?�{�GY��q]Hw��Sp���ԛc�\6j�""��,�c�U�~t���H.)h�'�j��1y�&��9�=�mw!ϥ\�/r��(��ԅ����@A?^z,0y�+� ��Z�kz��汦Ն5m��D,��:���%ٶ�ӸH,r�Z���S�t�o3�6?�ΪZ%�]�3��z\�˾W_9��<C���~ ̵��}��E�g6����>����|�h^#�b�4�Y��|P	����۔W��׀K�����s~j���;����i��p�8��[x���<�:�������߉G�Eʔ�9y^�L���Q�R  ��܅��"�p��K5l��ܬ�6B��b�.��4�[���1��k��0�[l�kKO|�̂����W~;��<��F�Z���8��=�ds�z�H �Xu%��pp�K��0g��S��
�ѐf4��+^}��)0W[Qf<�& ���)�6�����Q�ִ��2Z���np�D���f�����k��kE�UN�9s4��Je?�A^�H�J�9ؔFv��>�6񀧉լ��A1\���w�<X�E'��t͂yd|�� ����xr�8���C���';�������Vzruz}q�;H�]ßV�ގg����ѱkXg��S�2�z.�X�`űYI�+������%�)=��[��&$[�X�(�WF�"��>������9��^/`9D��]~b0H��H%�h��H�gW��C�c�?�4�Q��e~ď0�W�l�`�F�X����,p�}��H�EM7����,UX͹�Ϛ��?,l�_�'i�����&�u e��J,��M�zeᐌ.4Iᲂ��*x�aXM�����2Gf���"0�mT���u;B������?T�t�W�&\�uL�yԲz6��,h "8����NN�v���&�%eQ��*�a�D�NH��v�)(�r��p޼��O�wW
�m��'x:�4����pU�L�����ܩ����o�~����Q�!^}1�� <�C�LQ��G��w�HZ�-A�By��=��Ρ��Ƕ# c��0��,P�����B%UܳXy�Xg#V�p��g�6č�&~K˥d1;�������@��\�����5�QF�]�k�u��CV�U�Š�U��o�`������:���ә*ė��F\x��dr��u$�,ʍ� /.9 ���KR������$����q��t�<Z	σ'��l����7P��5R+��_=��΋0k�@֔������
�a��J�{�1{�[yM
Υz��%ę��(� ��.���:�Cы�V� 	�#8�(Ϯ^lv3��.*��b��cu�OVl�4�f�����-;�k�����T+��݉	�vk�:��yIs�H:3܅E���q��f�/SP���/�.�isZ�s3�V	����9�ˡ3�����(�w�:��ʤI�n�(�J�/�`�(Q`B2+���{"Q�Qn�y�ɀ��Ϙ���p�Lؠ���
�&Ջs(A��ڈ$���/�\Ł����Y��?����P0�k�˽!]@\M+?8�M��T�3� |Ca~	��&|Kv������Nk�ba<��) �cȣC��-l�p2 ���;3
t<goz�9�T�6,Ψ�-<�E�Ë���(���X����%{aS����;�]�g��Q��8�E(il�`Y�h���/�:~���%�|#irN�y�H:����F󘒒��;�O�zg'�/�U����Q��p��::� �3��ݴ������TZ:5֠Ab��m\�_����`�/o�j���������A�g�����X�y3:nt$gy�h��܏���4�R�&E�I��~��蓍@C���e��I�s��ޙ3Dx�u�[�^�W�Qnq'�}��
�Ox���@��s�k����*�zָM�0�B�����_W
V�Zf�ۍ��D��V�� D1�T��G'�~.��[Ȳ����%Fa��2�-&�f�ڍ��&��!d�����t ^!�巠���Y�	�	�ӐP��������:��Bf�/R[_-Oz@F4�������S{��_*�C.'������^����o?�����������@!K�9�����+�!WV�9I�m�d(�=�����m���"Ai�5��]7����B�@��g������>ՁoE�xt?�k��&(Q�KD�t*k�3h(��7���y����\�j���A�3aX�D��.�Xc�s%�ɸ!�l-D4އ��!��ȷ��0����K5��=�OCQ;��j���̽	<��s�����I7s������*3�X��ᲊ4p�u��2�P4�~I�o���^�~f��w=�`�0Wd�Ѹĸ2E28Mڭ�%%�����U�ua%�e�ҳ�ys�S��	4�s|�u�E#�V2��ky�_�������z8zD��*c��J�iF�ѐ���������鯩&� ��"� �p�K��ɱ-`������P�����>`:���G|�(}7ĕeV�kx��g�GN�7\a����gW?v�5�Թ>�o�GߩQkHX��{lc�ة�E"E��b�C��H�Pދ�Re����	~�5�k;��E��N�3s�brN�Ji	y����!~���iwJd)���G�)߅k���Q*��(Oe#�,A?�=
�PDz��M�nV4��Z���|K�S^p�(w��#����}%0h6��ksC�A�pP�x�q��i�I����pu7&�V޴��dy�W��C����<����nI�Y�i�N*��7���b�I��Tm	ԭ	{�ɕ'��g@qV6k�PpS=���	���/�"
��� ;���d�D�,�Z�آ����B$/�QXg%c[�*aN�����z U�1cB2���b����,5f��Ų���]���>mo�7>n&>����߷�P{m�-Ҫ�Xd;� l��I-�T��29�}C��ս�����֓z4}]ӏ��j6:�}�ağ	.3]�d��,�*̍�����\^�\�oxʵ|z���Ы����H#��.���B|A4�1�=TV���kåؔC�iBD����m=ÊA7Z�;��Xu�T*]��N���?�<a��٥��?�ɱ�̆�w�N;�TF5A˰xY��w9�4�lc>��VZ؊K����X�/�z�H��MB}��D�����Q�t(p]�c��w��Ǵ�%�1!:�y��UzSh��7%�]�\���c��e��(��|L��{ �
�^�n�Cŕ_b_a�I�[�N�:١��7�/s��@��]}<�>��ޕ҄���<���!��2��c�M3ȝῷ��#P��, ��-s� ;ۡ�\�	>N{�b�P%,�7�qXm��g"�t�r���?��D����)�Yez⨗>�Qs�W��m��?�Q$�{Wg��?JX�N$��U��1�=�MDG�#�*R#�i�	űj��q2��'<������!A��D=��56w��{��Hu	��s&/�^�ur�������^U�}�%rj�v@T�4�6 p fn�/_#x6�R���
퀽S�����0F���4�̾��0�����_�P�:V����M�s��:C��4A'9��G��z���+p��677�[���h�#��x&/I��OQ۾�1���N��m�.��ڦ��u�qreJ�g�G�cu�~AFM�ו̻Y��H��{ \:�Q[|˓�n��^��O˷��!�p:�0�L�ةz�7tM▏\���ثE�C1�a�U��X�z�z���n�Q>��A�w}Y�V���FvP�!+<�.�n���Nx�P����*��'cUW�R#xE����.a,<��rO~Y~���ĸ	>Ƞe�KG�J�@�H�J�%篌������X�=1X�7M&xa+���L,?"�P͊S��=����� b֘��vT���齬d�>�}���Erk�����y��#%R�x�է6�W��K,�"i0	�������B�:5XhǊ7f&�_`28qx��ـ)p"���^v=AY�����]P�8#
D�6+���[i�$
�o�7oT(@V�IV㹄a�N�64��=e��l<&�zȠ�/�}G�5�uy^�!����B
���rZ��Q`�f�j��54c�O�`Ⱦ��"g�ڏ�+���y+	���,�[�C����sD���W����p��)iޫ�=�H�G��-�*�O��	z��"v���R���b+���O��R>����9�GK�.�1��bҔYzjf��Pha�����F6����*@��P��K�ٙ�,��S��<���0�=	�e0�m��{f�&�Y6~YfJU'�{����¥[�$��,kT*#��!J�Ji��±P��5m{ X����gl^6S�B�D1Y��g�8;P~�=˫��!Ž��Ў��K�'�(�4,v���[��B�;��O�>i\0����Wr&�y���bxԽ 	~u�|�[����A���Q��[��L����R^��H�Ҏʑ�o��Ʃ�jW�f ��ޒ��Ŏ�X�2�
�8tXq����z*��-b�� K� �p�F��	.@%��jgԫ�65��3OI�_JvA�|x��yQ,g�uP%C$�L�"G%�%@MTněϙ�F+i��Kx�5X�5(�Ǥ֌ᧄd�n���oP��l��7 5ӄ��|mY��4h+�����QD�L����`����v�b����/	��{C�Q� Q�d���ޫo�4L�-���U�k^��j�]�|����_�,�6��;�Co�h/�l�R�&�>WU�f(��[NU�/�J1�%�/̻걭g�d��� �imG%bJ�M5����Gcl�K�t��%C[�U�#��3���U4��Έhk��oCH}
��T��_pfW�V