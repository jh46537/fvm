��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨס�>�6a�
�Ys����'Gc�$��@	[��%���D����7����ӣ�h�m)��@q-�M��v4��䆗�g�})о�v�z����w]�V��-���;�s[+�+�C�Ks��H���,gjHN����24h�n�#	~��E!�5�����q�TK�=�IN��
U
�D������
�K����bS��j�mrVG�������xw��փ����U�ӵ�+�dr7c�)�J*H��Wv�'j�̒����.X��/�3�( Ɔe
.� �+��GwvUkY!=�'�k ���d�����4��ޭ�����)�y�f37c�d��N�O�P��Ц�j߄!���b7]��=5
���r�q���$zu�V�2����U=A:��r���&( 4`��A�,�x]U��j�ֳ����a�t��4Y7"�>�����}ȷjgLy'(�rS��ڃ�!Ύ�pH+�ܥ1�4
�Ax��oh��+Gꏵ���c@b_
��GC K`���tx��ZP
����2\��7���1Ȑ�<�fY�U�>�n����\��v����p�d�TT~���六Y�����ki���U�f-4m�+�."��㿿M���\�e7�x��|~"Хm�#*�r{�I�^�<� �x�]��݂Ȗߐ�mFEU�[�[*�o�1l�ǩ��+�ծ�G6g

}ښ�3����Z�hv5k��!V��� �B� ]y3�Р���Ÿ�i�T�E�#�Vj⼉^v �z���^�M���N�]+��x���ڔm)��V����q
C�@�o��H_rp��Xe��KT�\	�-.����Qy������7q�����ZV�tf��q �W�цS�qb+������2*5j��>��p�ӗ����.�5�j�K=ō~_Cm��}�`�F��5Me`u2�tY[�T�1r|�߼�)��`t"V�� ���.�0���
��1�gלLL^���QQ��^���Z ">��TuV`&��Q�����1�&j�Y�JL�7�oh�����[
n�%G�����x���j=vs�[�g�]�����f@<jf�Ԡ�[�}��ǩP"�,W۠���n��Н�<�	d�2��˵<����琉hx��]��!��9�XZ�^dMt8[_���N]f�k%Q���:���ʊI�|ó�C���p)�#V}{�|?7��el��d�<M�~�]��ՔpR�0W<]��
TE-�~�5(	�l\_Vƿ�ſ�0 ��L���A��krxB�"��X��6����US��CBz����Uߛ�:6�О�?�s�����ܢG��!�H����	,؉62+9�
=���n!��jI"����5���������us<?�J4��Kw3�6��6E֞�T�`lλ�>��}�Z:CgK��^a��)wP����^T�+{YÞV�=��1B�Uڬ���A�Y�l���ŨN�c��X�K>�N����������$�UO�����	�^Fi�|]����z��<'�po�p��D;���-���J'Ǭ��G�9(�	�hOW`/�
(5�ӨФa�q����-_pS�$dғi�x͝�RTMLu��z�uT�Ko�m!�6� gI
l�>��X�5�h�Dt�֝�s�Y�4`�%ͯ	�l�����S�D]?�-���X���Y��H��d=�6��x���1%��
�ݫ.��]
����Gp����Q�P��ĄV��*��郶f�tF���s'�{�2��Z�Lx#\
���9r�mk�c�������]��ǋ���O�]�p�`Ҿ��2 �g�HY�2�s[�6L`���ϵ�!��U�$�d��mgF��9j�t�J�(��GF&�#�K���$���ւ���'����!�/=���;	��{�bܼ{���-P�0|Bѐ'U]�w�6N.��Ѕ��:U��5/�b�}����N`��g�rUz	42�>��g;M���O�)m�+�ք-��5�?b�lmi�''���Ǝ�(61[�*e9Y��#�>_b����k=F�)\�o�(o$�M�S����G�D��.��g6o2�$�q̶\Px�r��^Wݯ���K�p��a���Ƶ����ӽ�[_m�Xˏ��FGЖ�		w~�/�*Kr�ؼ8m{��<�2��A�rhW3I�- Pg��yvP<w����ҬC�as�L7"~�D�P]i�'�Z���E����5��լ#o�`��)7XR�=�B ��E[4�$��aXqI1��I'H�}u������Y'��s1�6�����uvkSҬ���Wt����TJ�� ��M�R�o.��;\>��f�����g3Q�;���;��?y�S�Ċp/L���i3׬ur��S�����Hr��������#��� �+o��Ē<+V������Z�Z�"��(����,
�����T �� �s���%��!���xҿ�8����Ւ	�}x�O����h�ρ%M��2�:45�D��@��K�!��]�:�k��lЖ���x���)��m�kj�0�h8��Yõ�7~�g�\�fGL�9K������w�b��u!��B��;�~9�咙>�e�L�nI7��`����?P�|>su貛�Py������-�!�7�]N�-�d�[��	�[��H��!��cT�/��KCe8�}�rWL�p���Q�.�.�������fs�0[^oNL0�˷�Ŗ���!?L�un72������k�k�ϧZKG�lT����^B��������
~�'��FTw1wک�'WMtL�h!9�Uy��� �.�/�(�����e�k`�a����N�u�8���pY=����x�M����t�U��{W��}[׊�G�Q���aJ1�I� ���ѣ�4{��I�~RÂ���6V�[��|��0�ͫ�硂
1'к�h�x@D�!.��/�b�S�,�!^�Dڵ�ο)	7�R�K��@��F�����]��h2�˰������N�:�]$L�W�H\՘�7.�Ux�'�v�W�D�})3�TY�qAE3o��X���VCT(^13֭#��I�j������BV��i� 3�e\rS����U��c��6Z�w�Y$ �<N8B�.����q�:<m�$d��O�r��%F����f�d�
sܨ���|�^3	{�@G�q��yp #`IY���U��p����kge�R����l��I�������q�3X��&g�٤~ג�Ke���B��|�<��74(Q���U�.młioa�>���C#���i]���A�Uq�m�?�<X�L��s��<աCJ�Nv�:��ᖒ��)tϾWg�,_MGD�D���V)t�|Q�@T�cо�$���� "���`y]�~e�h^u��<��՝Q���H2��o5��GL�A#W����g�8%[:bTنF�m1�_9��
�7�+#Z�Ef�§�p�y���Yn�s"}�.v�	7`҇SK3_�����.s`�� ���F����*?�޿��&ܢP��D�1�]��{V��}�׫\��|�sq�Y��U7��	��,O/�:���r�*s�h΃~2��5����x����[��6 �,hY��a�OX�	?K\kr�;!�_���W�u�*[k7�Ԍ���%�N
+]�@�o�B�g�R� ��� ѡ����0&u���݄%7�v��Z|���ͩi
Q�sQ"�Z���ެ]��w��6�������u1t��Cl	"	�����I��'�:+F ���h������BE�:�Yn{���{'q9[k�.�dN�)UL�Q��O�k�i��Tn&����+Mb*6��A{O8�cE{�5��I��}��� ;�L=�օ}de���̌⼐ҍk5iB��\NO����k�p���a��&=�:��vĸ��N�L���|4�Ӻ��VŖ.�M����]��i�M��@��SP������÷��C}�9l0C�;rҷ��L"?�;)`��-�m�ĝ�C:�Cu2	n�e�@C���!H����Y��*�r@����?G�]�W�O��]�
�#�]�o�F ����up���p��J@)��vޜ-��C\K�L~gUCVq���7U^�䳷��W��u�c������F-���}�Mx�T�ɪZKn��z��#�������������J��߁t��"��������p\Wg�%��z\�+��VD�9��v����l옒n^8��<2x����-�m�F��	�!Qr�66h��$ÍS�}�	�*`���P�M��R^�����4E��rR��/pE������ǎ��bnֽf����L�����I�����DSԬ:����t�Y0`���]��L
�X^4�W�r��&�/eOm�*�|Rv�>Æn�WB*��mҔ��&ٸ��ģHm���w2;~���wKKG�t�*�,��mFF)T������kyB5y����q��0}>�GS�������qH�ݏ$�j���V�:����ɷ6NtE-�Zq��V��kw��q�r��I%C�m�����:6�EJ��~����ť�2E�[��$/뙽�Tfѯ.��qiGs�����n�%�F�/�B��4�$l~�p�#�]z0sʾbG8�wiVʪ��K$0�İA�YO��˝�u��s�{3#/t�9����(`�
�~�{e܂���!O�p5�>\І�C�,�����.DcK r����P9�z,Q��y<:�۸k�O�H��I>k<�|F���HuvW4�?�s��CGҽT��j�,u���h�֏2�`�{F7�=��ts<��*+f��7������W�rX��%�����6�kYo~o~�%���~�4$\O�j�zH���C�h\�E�������	qo��ٰ��1h���cƣ�����p>V��K�葀h�e�Q�[�4��O�HSҞ�<G��0]֗-��^���i����W�vO�[+�}������Y_k���Ϧ\���Z�[�:���
mM3������+�u���!��`4�)��@v�ՠՍ��'M�!�����B5
^�g����/�p�����7�R��3�