��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[��Y�PZJ�O�e-H�E�".�h�Eo��$w���I+6~~ɷ�Œˉ��r�s���o?#�;���G\�iv<3&�罟Qq���%:Q�q$O}m��ط?7��
����(GӦ�0�ɋ���N��V@����� ��(ׂ\�򃛧'�쾌˃��%#��8}��0O����|�S�P��0�������K�'�����3]q���L{V4&����w�AZ�y�0F6+�kD�d�����T�R\S�c
z8��1������l���\�x�'Β�O��5h��\��g��0������֊~�cX��c}�ZK72W���X��*}HhG�js��9��u@���rG���ڌ�:��3p����8��+�`\붱�a���Փ��;ҿ��h�T^kf��+�,)�ac˗�-,N���׾mS#��Y	�׭�H��#>褍��蜫UX�u��e�G��*�4�a��I	qU�yp���_S�Lg�6pk�'��v��C6�9՟�����`�� v������D5��g�0ʝ�Mu��]�G�?#F�	�'�Y3��l6�M��g�ۡ.�m�#(%�k��Ϳ��}x��*A��wX���vB������H�NM��E<�#G+�S~�=�Q/�W�X�+;���q��	K676;��<��,A�W�sR�8��c��딂�7�������ҩ8�;��)��wA�],���6Y��|�g!}\䓧�FW���Q���y���vmp��� n]-�rX#�#22�/N�I�$({�@܋;{8��a� m����i�wg~*d�	.�p*3f�1�������z���G�7��yV")�]�.�v�6��R��}+��dy��ٵ�hრqI-�oť
?�](��i��u�u@Vt'��@ �bbD�W�YJ��&�����}+M�M�MS�A��x�����q���/1V�4wYf/�}�]6<V>*t�ى�/��$�˩S�=��b�(
��V�oIb���o�@b&��u�i�\�|cD�L���{WF]�!�u�VT�֘��� hZ�F�3����S�E��X���S�8��R����@�2fv�n~�-�IJ3�W�6.ib���j�v5LO�H^[��h���.f��32\@Cۇ�������ڱ�褙��k�[��J?�J��q*�Hc-O��i������w �����qL���}Rи�*4���vY�|@e��hy7n,P!Y�^�:�}kqx�kmE�fbU��\�EN�;�?�'�$I1�ݶ��De�5����Xr2i�S4����@��FH�`����i��Y�<��@+����ջ�DC��k҉ߨ�,�J�0��e���D �+�x�Д�<��ѓ(��>='��Em�eU�]���%�A���qQ���H� ��,�A�؝\���!�x��_a�	ɢ�6Vi�Tn&��d�z��
.�U#˔��;ttK-�S�^�/S�C!f ��"����c�P�2"���
�U��]��ؒ����E��/�)�0CY���&,/�׮^7�=�@#��хb��C�SeG�ՠ?h3`�|�8��v �S���?���^Z�J�Z;�egr�4����d�޻� n���m�k*-br�b������-�`k�R�6��-&�Њu+'���J�B#����و�q�q'��ƅ#`Q��`.�w�o��<˛��ݘ�E�h᳏,�Gr՟^òѸP=?A���� '��-<8PX��~�;��CaT��"�� ���Q���+W2:��iϣ�jj��F|�Jt�;�I�a��1|���o(R�fA�1������(Kݠ@D��\��sB�Og;�Ѧc�Ϟh���z�Q����)HZ�<i�q�5��z�Ԉ�_�2bk#c*4`�G�\]�OO)�V=��	V8CL�0��G�x�_(��fq���-u����̧��z�2���u�O[e�!��h6gύ��U�U�aΤ�78�J����.��կ^���7� 7�@x��8	�r�A���j��D�5��v%ܚnjҗe�k�u��{�Aj���	���
)�a�P��i0��e-x
jd9�Ȳ�N[��T��aܐz�ds�N�O�����lN������{,_��+O���� �wB�#-꧉|� ��T�ko ;a0q�֦�2�����HC,y�fp7��̝*Q��8堕�6��[#Õ�1�E~�yi�X��@x�R�p�G'��X���~ -1%��[j�3BJM�^~���6�T�)�����A�^%J��x�����x���<KiVno��?˂~2	�{��j�,u��>K��c|M��~�[��@�PP��s�59��!B�����Ԓ���S����c纜S{��z<�X��hRoθCF5I@-�@�q9�N�t@�͕.�2�����c4�V�lwƍZ��H����j�0����K1��#^��`�f�>���|���E��?�y���=�������i:����pgDM�����O	n,��>b�����$ ��m��^�IQi gK�"���F������+0n�8e;�K4���X�,���4�qH�ǜ ��g8�HW�hيݫ�j��� ������f!��^D�ȇ�M���n�Z��ܬإ�:k�̖]�U`�,��1�r�-��D�r�y�'Σ���Ӿkq9_�Tr�Ҁ��2����lF'K���T���` �i�Ј`s�|���z$��%$3ɞ�!�`)o���gnܯ�:��$E�3iLVYƲK�@�g��c�~�CzabY�A��*�����tf� 1<#���|�d��m_6L�=��J0��B����+W(*dW��S���������^ɒ�5�`mI��W�������}P<���>מ���``��A�7� �p�PC,��槭?�s��Î߹����F�J����PE�	b3��i�1��{���UGR�i���2�
����E��p�J�c}����MWѿ��+��ې �/�6:��PY��[�����^��@D�}&^X�Sӹ��Ң�	h$L�� �|쵅���;lLIۣ��;�1�pKc�?�a�NS2�қD��+f�@V##��X���U�����1���,c��\�<pIC�Vu��O���i��a�J:kw������7�_=���T'��Tg��A��w��|�`�g=��%��Q�H�
��yl�D��g���T�**�ɚa�@%g�(T�r��h�\$�(��F]�)���zI�g����vu}%u6���R{�;�_�\��W�q�pӠ���u��s7�e8uիJ:"Z����f@u�0e8���{ǃ��E��t�����{<�g9oz��p-���G��ڐ�U�(%���HRJ�����B8D�}�����ml���lU��Q���N���4����`��X���Y�������"=�E"�Ukqhj�gu�s�D�nf ��eޣ�6(A%x4����AbI�
x�������L�?ƌ20���5>�+c�cW$Ip�)A�L>|� ��{)� ]4EO���S9o,�$%VĤiĥ�/�>8��:���:c�ӧ�X'�(a�,02W���p�m��a][W�{ e�����7��}��<YK���k���r	cĕ�g�HM�bC\�Ŋ�7o�p�*Ee�8�L-�8>�g���aD�.�^�����q�,���>��.�b�X�����$�,����{���w8g� |L�Ɉ�ڞ:"O'�M+
D,L���8���/<��\B���jq��	����{G؆d		�
@4��o�����,��:+��_�_A,t(�)��T��LaZ;��it�T>�.�O/���|F� �;EC��<����BLb���:������ԋ��6]=@F��- ґr��l~t�ݬږ >�;hN���7���L��9���ؔ�P��)�7��
���Ѣ&�aFS�i�ceM®����	�9Z��0�k;��Z��k������`B�#�~=צB��tL�%c?�J�E�eƀ�{�f����GM���J ����.��` �y��SYZa<Kh�5A愦2��Km�wȀ�;��~���<�5�:�CHt)
�	�5��H�:6lM���1g���?��k�s��7��0W=�O��q�/�^��o
�c�2e�d&%�9���2_%7Ϸ��0�u]@�����vh�C��@Bp��2��K�48�l��3�{��mqѓ���XǴ$��?���a�;,yD`�k}%sC����<�R-��A��
�[Z���lʌ���W�,0�1�b SDm���~��Td����X-7����ځj�1tj��n;b�����'a��F�ڕA��Iz��G\Æ��V���o�D�ˣ;����3VkP�m���t7��N
a���(ˤ�T'��s��1/K�AL�4��t �K�2�+�(\T��JJJ���nq���Yr��fF����d���{rSu�ý&mM��6⬌{M�ߵz|���3����.^2u㶴�qf���
�T���f�SrJX��,Z�V��`�l?/LsU4�]�� ����[]���`dt��d'[|xab�����@+�N��~O�]��B��t��� |�i�X�����ذ�k��с6��,���T9ek������o��,NX�i�f7hO�)|��YLd@���#t�|ʗ�r���.ݹ 7ۂ��|Ggkג,@��"81+?��'d�� ��@�k���V���%$����:iƆ���z��n�c/bC�	Z�q̈R��.�j(-|�)V@���bM�_��t���*��j]�4��n�&l�{(J�x�U�0���3u���zI�7o�������e��a��[���[:n�E�.1�H�9�2���m�Q;;(�X$���/Hd�W?�
��ֆ���~�y0b�7�X�m�I��� a���+�qʂ����f]��A!�08����W%�q#�w����8�����ҷYL��v�&�Dti����H��$$S��jSM��_%���66 ݏ��*�[z
K��-(�R������7�k[�,�"g_���Pn
��y�����A8�B�S� �xM���UbB��1��_8 Ď �k��gRk��#���S'U�.�'_eޘOq��?�#�'N�~�1n�H{��z����an}��7��\���3=cX�ߔe�Ql��M�������-:�Y?�'�U��B�'<�����R9a��8J���F��Z9���A K��mMt�yS�m��h�N�l/�}t��V�j�϶�F���W,����<��ԃ]o �l���D0��ϋ��Oː��y��q��Z�kD?�s�@���OU��VC_��^J}���2��c&IE��'�ӽw���c)A�`�}��@�{9S�8�PP��~͖���ōmT2����VLB$5/�^��њ��'�者�mL
�}x��ܨ�����]ië���������վ�+���O��k;��p�{ �zF�de��t�W#�3#�֒�~���0���a9 51,٤���N��o��֯���	N[���i�	B�t(���o�qD[�y[�����q��8\=��������/����7 _@�qMԺ�X�䪇c�:X���j��=��r����R��	�s6\[�D���è.V�!�FRBa���~�μnp�N[��v� �Nmxx�$-�f�F���Hdy�gz4���ƟR��]k
�,��T5���m��b��oZ��r-� ��Sm��Oa���}���I�y��i�AH���ǧ�<sF����x� @IjՑ(j��VI�W�-t��Z��X���ey3 ��b�<���4��3�W���V��=|�Yn �����Ey��l���%��(��sF��g��B�s�d����{a�j���>�t��v*����^<�䌾2�(���r�y��wf�xi�!/������H���Nh���ڜ�h�+�����`VWD"C?����
��÷Nj-���k�>D-�k�C��Tޛ�g�"����-*�^���όO�Hd����ܣ&���zlD��%	����k��}<����*��u�@��#���&/\��]�?z(||�!�>��_&��p3��=lW2;ck0Bs�ݴ;0�ݥ���vvXX.��E-4,}�����|p����Y6�ZJ�!�8�.�S�� �K�E] 52�t5�kyE�[�T\^����N%��Vjyg��KC�"��y6]SGXW޿O��0Rm#5ï��Z3l�(m�:�P�[kL��C������F�ӹ
�od�BJ�m�,�b�/N������h�@4\�5ұ#2�wg�����
$��8�;�Z���p��x�	>RR{z�Ke�������kG+�@�#���L���IQP"���Vt8INч
�W!�FF���ca��M=>,�ڊzZV��`dUK��\�(NqV2S�]2�:�?��\�^E��Cq}���J�DA6��v=��?7M'١`e�ߔ-�#��U��%��0_nG)�vɄMw+���'i4Q�G�_K��:[�P4�S�+t�Q����)��Qgq%�	1J���2�h�GjV>b��S���'�6�R8��C���7����|�_bt\��WM�-�$���B{@l���:���0r���3�yLE|"+������'���*����B�Chn�r>�e�,�4D%�����Q�-4i g��Le6�A14J��iz��Y�|�qm�df!��G����exEYzU�l���"\r89�|��g���(iWZZ����4��Ӌ��p~�E��}I~-Ujdm��[�\,�dL�{�i��o���M)�+�2<�(�a����1:9P���]�/Y0Ak>�k ��WV"8I��f�ߝ��BN��rOK�.�V"0��<��f�;�|�l2��~���S$�XPFiD�Q����)�=F�:?웳��8����OE���XhCwk���|Ҫ6���V�������u����F���)�<�B:*�V�c�g���N������c.�з�G?Q���ɮ-���q|K�H�|*qLJJ�8V�yљ5�f�F/xe��|�l8��J��X7�#��X�:�� 1�m�1_���ǲ�˂8����L	7�]�����t?�ܩ��w�s�+\U���d�=����&�­�,f���h��vN�Twn�/Z����l�+�W��Ԡ�YRv���}��I��R��j��k8B�����^�-6�J���T��X��C�CTAu ?�c%,mP��@��TyW��?J�VX�>*=0xD!�pѸ8彐�\NcG	�� ԡ���=��=���W���&dX��TK���X|�G��zbXŃ�Z�ϲ����+��v�$���#YWE	FK�G#����a����s���r�#/�6���2>G� G��<o:+��/���[p��7��-���	�Џ�F��p���$��k��S�E�EEs7�e���oC��~߲U:k�����G�r�?�9k�_����}Ȓ� J���_Á�z�-��O:Z+���P����V|P��f���ɍ$;�������&b�ipA�@5ŏ��
�:�� v����qyw�xC��ͼ~P|!E�TH�Vů�$يŲP�/'���4G�q%g.�d�[���Ь߁��x@������bn�)X0�w�^�xXT�LK\V;�¥K-DՏ/����p}��|��������Lͦ�J��7[7_��ŵ|*U�T0*9��15�D{��h�#<��{t�"8����
�zs-j'������\���
��#��cУ��;�&��^�������1R�oz�+�3񎚾���r��s��+��!��������N���S����U�4�4����R�.b�w2�fz���T����J� %�u>y�|���}(�-���ҟM#5;f��TR	�=O�k����2�@����.��F�Q3��G3�O�����-h����_�b��&���\�eb�f\�%�B�|
�� ��Vmf�u�'f�1D�@Ԓ�W��:$E8P�����q�̟�р��
A��9��c|e����mwAjz�����a5eT��c?! ��(�@3o;��p�1T��>�l�����v�הO$w�l�S!��>>l��kP����τصpS��pS����5��7ը�����1M�W�]Կ��OE=F���{"kUN�Be����;!I���.z���M�[آ��:�pB�s�ޝ�x)G�Ch2)�1��M�����f� l1�8/��NZ����]?��bi�//�k�|�|�|���s3Rm�ޫB�K�P�r�n�S~H�1mG˰�8(�M�!�Tݸ��kT��f�-���V����%B'/����&�Sv}�U��;�p�EOU�sl<[h��˖�N��k���[�WXkC����FJ����?tۀ��rN�I\]��=�*�#�X�������-M�Zb�N������G�Т�b7��Q��/`��#E�F�>!�m�3R��Wn8�Z�!�.��������7GNR�w���˄���}��Ѧٷ�n�o�_y�Ə� ���cD���
�i��`F�3��v��*Q/��%3��P�zr;��e?p�cB`g����X�@�;V���`�,�"#+�jO�ܜ���M��@�����[:X\��q4\��A,bh���/����?��N��:q�/B4Lb�B�?s<�=ys�	FdUP��=/�~	�{_g
��L�J\�tY!^��21(�(O�;z����|���E������<(�� ���Jn�9pi�ӔعzǞ�Z�Ǫ�:���!$w�R�B��Wf�5$xV�$��C��3?2.��]�t.7�`�8��B�x�8I�v����@ŷ�a����ɖt\��v䗨�x�|�u�L�;� X~�	�S� ��Ҳ��p4Q	e`���ht����2�i}�E��~��]���\������m
 ��N��!,�&����Q?G��;f'%!�A+��Pa�;�Y~V�"���m?�|��2�}�����(�Y�y���T��2JXQ���_�����0����T��D�ȕk���[4�B��y�u����%lކ'$�4��6$xT��n:�ޛ�G��]���j����/��(��v��O9�u�]׈u�Ab3��d,>^�	�C�R1��r�sQ$�A��[
9*�EV�J�ϋn�6���]�ol����+���,����>��٩�����u���6�H�_���TT�L6����f�U>g��K��@�΋����L��"������v��!Җ�SOr��E��+���%�hW1X�Нf�9#�1������lټ�{�츜�cy��1��Ҋ�K�Q�w_� <��`�e��%�����m"�Y=[i�Z:��S�H���ע�
��Q���V%��k>�.���b9�iI��W�V*�e'ߣ�H�h1���h�GCh�C�$J5ǥ�z���(OXW�?��o$���$�{�e���V�L���JS ���/Z�h+���n����E�K,�`��]ܻ��el�p�ے�& �i�R�~¥��#6�$%�.��������k���o��G&*̉�)]R�>�J[�6�ѐ�2��dP���a��4~(\��h�@l�h�#U ��Qr�KvK��q�%��"2&W,�f8"N��Q���-�IY��l9�8��i������fDƶ>99<c�n[K�}�0�=�a�Ό� ������ ��s)�U6X�/��z���UkO���e�9��ȹ�=�z���0����u�y�EK�ز�Hm���ؿ�[O�i�=��y��R.,����B�A��tv�����3"����\���7J��R	�n�K���)]��5�A�s�샫�����d)X�@����;dDrS9]lAa�	lG<L܊�<4	1�.�q��ˈ,I��9�0�o��aG��,�R����x�{U���0���]M����gAN��$5��eM�A�#ۊa�:�U�Y7"���z"\�
��U�U��k���T���J&�(�O�RJ�߯�ДX'�����fl���q�V��	4D�6����L32w��������n�i�O(M��P�1�7B%��a�j�ʦ7��V{�\��N�0w�'�mjħ��[5;�*fq��đ���˹�8W�^W/�x2�&I��b���K�j��D�?Y+�>{��-�ә�M����vS�@B�&�VQE#;�%(LУ\������vI�
�W�,:���`��&�W]0!�f�xG������ґ�O[��餌݃��l�ͪ=�����n��ny5�� m3�dmL
��d���H<]�1j�bi'�����!��(���]������'6),r;�#/�D%�����!�(�y������a�֬Z�������D��2�!�\����̖s��H�3�Pl��m'�W#�<XG�V4����1Mt��:@�}�Dw�VL�^z�V�@_I�]��2�SE����w��Ϯ��h3O�}��@�_v|�i"�f��2\n���;�H�����nK႘�g(���hb�uF�҂�K��À��5��b�6�]�c]U�]�-:F�lg��A��WΑ!٪5rH�{#͓���M�T�h_���w�LH����+W�ws��H(7Nf5t�'����	�U�EyZ������'�bC��
/@�����^�E�n�(�Y����ͻ$O��$q&/5��޹�.��9��ʡ��Gߌ0� ��L�?e��TIF��\���������H�`�ق���V�Vŏ1�V#N_�'i�|�{[�P�4���EW�|u���pC�5��|K�cG�iH9&�.����$G��+��^�1�z?���x�c���[�1xwIiB�t�su��a�0^`�M�Y9BY���!2j�lU� z�jˏhA`"�[��[fwӟ�U�0_8��E|@�;�mC�0�y� ��� ����C�$I�/�����Ir9���R�-�Y_( -נ7W���敢�^��HP���c�+[1՛�����H����mM���1ĺ�yz;���M��������ء +9�8�'����n+�h�_揄Q��X�~���Qg�����4�('.׃���Ř4�R�ڐ�����b�H}�� *�S=2Ι��M�^�^��zؾoe��D�����
ř�:,_/�B)�7��}?��j�?!��"P���w�_h������Ӳw�f�hr��R
�{��\���bg����k�
ڏ!Or�G�$�d&3��!8lf*յ�;ݜ�6��=��H�y�)�Z�;?w�6����ߩ�T�s�LIV����K �AR2���F�y(�1۠r�%U�fqy���of�'�J����+D�J�T�����l�G���t�.�fHr�3�Ps����hَӢ�H&��6�6�U���:�@����3�kڥ�+��V���b�5�q�i�ǅ龰(��J(Χ���-,����'0���A�)�&���q����$�a�y��H^����!Q�0��w��#`J���"��j^�`]������`ī�xg�*��Qu~4���PT����:MX���Ff̕(�!G���,t���n�[�2s_&A�ڌ�eC0J��y2�H���ȧ����0�~t��~��kT�[٤'�4c�L�Jz��)�Z� �:O����f~~P��S��������z��[��̧�g߃"��r-]"�E�dj4����3�w�����lJ1���a׵���s�`u��:�C�;Z��d҇���#���������]xߊ"��@Y��!Mf���P1"�#��E|,�T�@E���&�}si�P!���y�!tI'�g�I&��̈K�tx����V�D�� S�XK��"Q^��o��� z�{ܵ᥀�ԞF��?M�5)
V�W40\��8I81���}�=���CU0+�S�RWa������.�Wi��5"T��6��!�7����q��^pQo�9��qcF���"Lr^ڊ��p��^%��'Y[�1���VU��-��[M\C��L_Y��D!;�	����uCS���qK�a��t�?iǶ�<�l �ۂo�|:	rm;��%vQk9r����I<�W�g���M�w&	��h�k��Е���ʻ�е�R��4W��Gnj0ݣ�aK����x�X�1�v�3'�7{�~��JP��>*���h9��s&�jߤyV�@#bG+?����������M��{����}W����Z���jDIc����ub)!8��]�v ����%�� ��6�Z���N���T��y~�Y�	���RE���h��Hz�f	�{xp��ȩ���?�m����ȭ��I�(���� u٦�G�8��N�o�r�?�n��/��`�M-gtt+1ڷ����[k�����ayE�
����u��g�y*th��Q���/�f��b���B��a%p9�"_�.&q�e��'�JT�S���t�7Ԙ��yq)&��ⵍT�d�=�qQ��7�kԂ�ܵ�\$}�k'6�7<pVy'������w�������Sbo��3n�h'՝c1�p��4N9?A���a��E�^�C��w��A�{O���k�8	��^���0�_�6J<_Q��y�$����*�5�����>ͦ�u��Z��NŠϡ'�{N��KM��O��^���õ��<�Z1�)�����_(�n6��r o+&f�uh�i�T��ep��H�4���ڏ��
�2�*��ݠ����&n��9�a�e/k�EI��r��Wl��E�c(T�B��� �vJ���d�C�]�A �A�n�}!v%���4�$W�I}���K�}b�B��R߭�}6[�������r-~Pf���K �;?�v���x<��L�r�x�u|�\Ρ6�y����xŗ�ڼ�E`Y�"#�̋v%�F2OqD=Ƚ�5 c$�_�Յ
�)�"a�&����&)0��"�A��vu�`�w��y��)�l1��0�m��]��'�~�}�u����sm踷vN`y]-E���،�j���㙀$ԝ��Yn�s�ɾX�(�o�zxpb���?|�	a�Ӻ��s�%�����3��>|$o��(����P��U�i��j2f���|9g̻>�<�@�\�I�7l:5���)N�j\F�_�ȹb����'�t��I�:d����E��Bs���&�4p��IJ@f.̮���\�&9"����i鬥��-��d]� ��^��$� s�`�����o���j8r�$���M*2�%�s�a_`%�Z���u	��qӖ��˅��ժ����h�G�˛
c�0r�U�Gx0�u�=v��<��퟿7��*8+lA_�|���_y�PnHu�3���Q+Q��(�賱,�4�#fP��$��+{�0T�$|nc{�ӆ˜�it��=d�b�9�Cq��'���߷70Z�e����!�/BY�%� o��͡��Ϥ����\q�����Ym��T�h4Kp>��t<��
4��8�*[(�߱��w�4*�n�[T\u|���0����sO7���#�Ӣ5&5d�r��;1�?~�����aN�\�]̀~�����yvx^��\��Z�_s����T8�c��-��\̣�X�(q�)��E���9#�V��'+jx1xJ���7��h(��d��)O��>��"��j��]����l�3z�����Zu�a%�O��>�O�~;���5iͿ���D*��4�.&��P׍���\���Yy
�`8\k�l����l�%�笐�`:! ����U�@i�kC{"шg�$&O�6v��n`�����~K���ͽj(y@>G�/bI�T2O���RE��tJbbBF�����IB
��;_�������9=��PP�oI�+;<��#���r�;*:����5��h	�F�����F8��T ��������'`����,��ER��?x{�Y&;9���3�_�t��'p89�Z&dfGY�	NU�.g��pf���j9���#,A\w5 ���˶�*y�)^]�������$�]�*��jJk�]��xyGN���R>��'�CU�^w4��؃��1�� �bǫ��f|�B�i��v����/�W������^�����eNT����Y֣�[?<�Uȵ���x�/�ԈRe�[��؝k`�g�C����H������I^���\���x���RP�T\悵�`�3��}�S��-��ρ��+��!@#�9�g�:�T��t�����X\���T�L���l�]ς~.h���d�o��>� 5h�����H��c�C����\�"%�J�x��6^(�>�r�D�F�[��_�<[�й����r@��>Y��ƋV���I�'{�,�=P$n���յb�>un��E#Dih.�L�� nw��CP�S�%�Bݬ�A���[g{:�ҵl#SkX�B���s�<�6A��sg{w"5C��p�<�[�g8�u~mi<J �gI~ޜ6�q_D����դ�*?>2�x�k��e���|�J��I�`���>��{4I0�㼐��Ͱ:���WGib�#��ct��r��ι�eZ�e�����v}Uw�#uϳ��4��1��@�?R�㓬��J�&�^0p�/S��-���u�)d�zA�j��ǟ:oq�bR�e���R��m���A���&��A0���P^�=�7�أ��6�=������	qk�+����
�7�.a��i�++2tZ=E_�����}�Mӈ���� c�V�W ��Ԧ�o/ί	��d�P�+���ΊU���{����z�x���������1�ǩ��m�w��\i� ��_xAuLGP؀FQ�9~yhc}8.&A�E���݈�|�w�l�vlp��P��!�cw��o�Zғb��������iWS�! ���GA8&#�Tn֮�ǅA��38�e �ұ���!n�iz���w��"\��x�D,w9���h8�~���rY��:����;�.��ˑ̤�d�\e�+R;ZJrW�F8�� ;�7%�0�4M���r�k">��[k*�n�����w4ҫ�kg�=\on*Pαv��^�� w�c�Z����Z2���$h��fXT��B�C�h����Ұ�#/\�;�����r�-f���]ZԪ~i�� ,ND�KU3d�3�mQr�6%�m���T�E���{�˚�oy�H2��-��z�"�yg�n:���ڂb�	���I�8:��O�j��B�n]����oL����o��`�~��}�Ac�$���i����cJ������<���8�$���L
�~����Cw�(Qs�5��YHt����ô|Z�6]*m_pT�j:�mRK]@���%����Ǥ%"�����u׶3�f}�� =˓Z7:z���̝�yάd:������ǃ�Y���� �U���n���P�6�=&NQ���K�B���������.�׾J�٥o��v��6�@��qI]���u������������A
��J95�l6!���Pԟ��3ۯ%ot<��R"��E���`-�z�{�އ����hY�``���Ӑ�I@����
]X����u���ęN��`\cg�9�D�3���	�\i��������	f���I��nd8K���q�' �����H!����(�����06�����f�_ib��V���?l��Oʞ4�ҍ�vuI�Q!�m�V�W@�Y`~��蟀��G�o��,T{]���� Ɛp��k
�P�@�8�i}6Y�/��֩�3��ڧӇj�I��R��4/*}�:l�E��<�[���$������9҈j�bJq���OJ��.]|C��+�����;��m�L������D�������������|4���[��ᛞ�L�k�`C�eJ*�C�0��@�}��f�TjZ1��/}D��-B�;��������><B�s彸'���~0���2�~�-+�_o<a2qQ84�������s]S��V$�o��Fd��i��Vd�̛��ɦ`.����ج����ȇ���Q�!�¢Z��T�+�(F�wIqT�	�ԙʓqb$��' �����i�,�Ɩ�%��p�$��o��W����ɰ����X�����
�V@���\��<��r�AK6wL�D���eF�I]���w~R6�
Yc� �� z�������+�'.}!�&�X�;;��BJ��'���=NX����8����3���6h?'��!�k�أ���j\���}�Ň[�_�P9�A����oF)R��xP��QU�T8U��݈�\�}wZASr�a�`�MGVЌ�)�w��yw@�YAӎX��fL:`,�m�]G)T����j�6����Z��5䃀��ңQo��b��%��-��8	5'�II�>T($ZP{Ц�6��HԳr�U�\Yc���,3z���8��Xe������y�%�v��i���9�Wl�*��+�,���0n���x���M��/�*i�uc��p$�-����:�5uy?�8i��s���ߵ~0<R�����;�&�,�2� ��y0Q��P"�j�#iC]i&�w+���ZrU���� ߭�C6�t�ؙ�W*h�������S�������ueDF�����J[ <՛W4�6����(���d�W|s�h[��z���7��	q VT
&�]�Zc������6j��)U
1� �nOg�vɎ��<Y\M�e�������.��1�]���ߦ�.�J�)�9C������;�T�Ei�}Q��/�E�7?d�S��1�����f��+����(ễ��y�ᑒ�D�ȫD�9��Y��'��2*�v(�=�H�|��{M��fD~�va�xu���z��:hb�?q�v
����=W��DC��2ڵ��J6Uܡ�)���5��J��8�}��c;�4��	������ E?���9S`��gȆ~��6�a��ᣎ#�/��Ѩ���r�d.b딨���s�W:Rщ����(uIt�������C��h���/�ih��9{A�p,���0�mc#?^��$���6��d�I����6M�QB�b<K�BQ�����'$>S��YI����aw�f"s�����7Z�א�X,j�~��6�X��.r�� 9?uHX�8�	�����94��fSS(7����yԃ�F�2-�Й�'ʝ(�D�=�ҫ'$�7�
��d���_Ή8&b?a&���7�� ��a;,#�^��[UAV�0:H�k�6�D3�c˯umB\i6��AY�I�+ayf�Lf7V��g��=��Xa�F���Ȩr�����WHù�s���fQiү R4y��V<&z8O��l�S��p��2�R��$p���D��ڰ��vHℎ���VYAE�����q�L��ꂫ��a�w�S*�ϋ�(چVk�:�}��h^t���OD%*>xNE�����a��+a��H�:D���P�.w�g���ލ��%{fu�ؕS;��s'"���1a�ӵ�V�֋����w�\���X�C�?����l��D%�[}�z/�����6wctt�8��=�X]y*�B���Y���Yn�¢�g��}y#~���
�/��15�����B�Me��/��`Z�t�1LtG	Ah2��lg����H<�h��3��`������*�#x�6iKU7��<�S�������S X�e�s�TN{���*J,SG�w'��`�)�Bm�h��PHF���R̨���;ˡ�6���2	n���38g�g�MSr�y����g-��f�v��+�s��A24C���� 6t&���6���U$��~�l�&�h����ڻ��g���5�ɧ���Q)_����r5Y�Q�.-R��~�0�reB�������+�i�1����o��]E&�6�
�����/
�s�H�T�-����GC��1�$�=�5X!��ߚ��"���G`�)/Lښ{����FV�ZW4t�m��{��+�{��|�ó yf
M����i�3�3v�� 8,��_�(ʱ�\�bҷP�i�Ҡ�4�'uJ�4m������b�<^/;���P�b�;|W#��M�Z��m����z>{��i���%��XT&��=�[<�࣊�Jf��Pw�i�J�7���pS��۽� ���cԝ�hQ�_чM�o#��`ls㑠>/��/ѐr	)W����	慩_�s༢���;�e���{,�����'�����4<�����W�&�[�O/*s����Mm5�q��'�n��?������e��-L��r	M�7MxzG~����y��4�h\�M�lcT�0��G�R��O�Ƥ��E9Ë��=����6��S��$�n���1p��g�a	�����R