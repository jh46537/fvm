��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�����:��=3�J�r	=�� M@Q �:���!+��?kC6U�T/���&��	�bK����V��D�Db������V��yfʀIG�D�Cs㠆�.�`OI"��\��L'1dA_���%��:��c���'P���G��4BS�_VW�#�6����ZT�v�O�! Q1�fX�<o��3���x4��̢�!i}���IZ���C} ���ӣ��L�l�,��Z���#)GO2��ׁ0 ���_y��7�����m��n��tGo$�=x:�U���������3�YX�"}�ۋF1�0� �-3��{^Yt_-����W1�>_��M�-�����������&9�^�?�ʄ�BϦ�s�V�gW��ĉ�Y@B��9`wg������t�I���Y�<���A�T�L�Z5p�C3Y���D��N<�;�n6��y��S�s�ok�2d�����G7��~!���e�}L#<�x�lm�'!�� ]q�����p�G��wi�p���^7�L$1B�.��� [�9������7�l�K�Ժ�߁�����1���� cI�W��~񃅩J�i����u�Α��o���/|�rӫ�� �^�K��PT��8�?�6���TSk�-^� �h�:��yc�pR�4��&t@������h�	�>�Lh3�蠊u�F���ak'P_���(Y����ꢪb�e����6�ޜe*=�s�m��+�����H�q����iz��}ͤ��?��e�/�W-ĥW�����2��*]���sM՘�a�7!�Uށ;��4_ ��:i?��_�0�m�y�לy~�{�n?��}�'b|�H�>�0_k�>��o4v�i���d�oR��QE�~��;��P��h���R_���{H��t���+a][�ᶢ�/�J���_��z�K����E�z�+v�U����2����MA�ֆ"ރ���*��2V�Us�Q��=�xh�uJ��Ԇxj���5K����.St�X<��������W��G���3���\��KBbH6.\��Ѫ�NYF�f�h!G!!/��. ��K���]r���%�9|,a���'�7�٫UF�w*J�=�〯�ז�a�M��ګ��VPZF���� k�h����W1vG�|!���<��f������-��xv�#�h���$�(Y+��E���rOV�!�߲!�o;ld+b����!si��%̉��F+ Tp/7:fײ>x�3���|���)e�$'���|l������c�ڶ[Di��U�Ϻ�A ������a���-Y_���5[
�(��_��Z0�˺��1 K��_4��EU`�\�����R�aј4O���.iMKy�Uھ!��-G-��ɶdv�#�����^t��MהI�F:8ѓ�Bo�RϕsC�����f�2ӹ�[� /Nl��>c�5��==D���0����';�;��3�3F�u��o7nq�h	���Cg�f�X#	$H!r��?�}���� #|/(n������3�5�g���ۙo�[�/�Y'GB�zV���t���p���MM;%��Kꘫ��ά��+���勇�l@BJ�H��ڬ�E��@�{���~��O  �k��t��e{�ĩ	���:�����S��?��u���&Lx����ŗ&~E���
rs��9V��*%�1�3>�>�C�m@#8�x�!�q (�����*�[
:�C=������������J��~�01x�!�N�~��K��*�ĉ�����k6\G�m�\ȶ'V�vY�/�G���rxUV1d�ﮭ��J�n|��)�^�v����q��3=�#���r7#���u�*�� ��ɛq` �`EA�����V�Fh���+U������{��|��JX;�1�\[v,J�yO�,�>8Y��qn�	�\�R(:T�"�1-�N�3T� ]9�e�>J�H#������Y��Y�~u�a�X���5�Z�~�3�dTc�����e^�ϬmG�]�UO��.`�Ǫڇ�tSq�>r��g�E��T��=Wo��ȋIm�-xĤ���h�UnD�XYXh�/_S���jeHtW]�qx����xq#O(	��&;�*ƫz�����~�'�F�~�V�����C�gG�	t
� ��0=�������RΈږ1��4����2�rO%��!|��KP�N�GC���>��{h�� ]D� ̄��pb�2>�S5�נ6ؕR�F�'�30>��x���g�Z�8�'TΡA���M�5��Mi�?i�a�e��%��90�a�������I���4�3x,ͧ{��io�Od��`+�}\�����>3�S����h��=���_ԡp��It卮`]���v$�j2�����r�?tӶ��fxu�m���5��4CdD�VT��v\�d&����栀�m�\�Յ�R�4oD�@�4���2�-@��C�]�!�1)�(����{e������1K��j������"ą��a�7XL��]��s<z~���ػ��k��8���tF�"�P���}�[,;_��蹊�� �P~��^%7��@{��Ji�5
84j^��Q�{�!-���x�~>��I���>�;��gh��6�gV��LN� J�@��V#-����z�t��=v+�w݌��M5o�-�xl�%��^D�r���bx(��kw��B:�7дC�=�d��p��Ckhg�q������*�?��{�\���r;�H
R>l<O���C�aP�F�=/Á��,�h��-Kŵ�	�LA9)Յ���F�����2���{�=���!y��m��m(7�kC"۲���۝�����	�,�c�+��P:$�:�~p'[�,&�Ť��Ÿ`���`��=2�H1��4~�ܘ��&�_��FA�?�=Ի^�w��B��><�%�>h�u=���7XEi�wiNi�q����]׶� 8,����U��c��d�p���:����D�<�m@6�d4�o+j�V��N}(�QE�4Uy�a�}g��ܓS��@?��R�z���P$;ŵ�c�|�_o�W6���,V�4��+����H%0����r'���xR{8�hS<�c�:|n8��vgNק�c�Y`�_���\�x���!����l,�
��r"��<=�a��֯L�2��C�H�q]@q}0�K�Q�����0#�qg�D�ݡ�yX�Gg�HrG��{����Ƈ��5Y��emL.g�FG��-�x�Ӌ��S�El���}��1yp����1k{����\;h�/���W��	�')�}�t���U��m\�;���JZ��g(�U+)���ϊ���F6���lT��2����'r�e>%?s���k�����.���;d�F9�a*���;�b�>���*������x���FS:�)�|�=\�4,��(�@�T ��Ɉ~�2�9��c��Q韜�
��Jv����D��~	�w�덴|���n��-��V�8*��3�퇸���_�뵖��9��x?��-���L��
卟��AS���F����m�,Q�a�m鳠Mb��&2.�ȳ�RY7H�t�_)t)��[� *N�XM�@���W������͎k���	��k��Zu����_�a�)��!_��< ǜ~�q�!R�f>�ud�
"�k�,o�s\�Қ�/��7��N"��_�cH���~%ҧ~�.��5׊J�ˤ u�KK��Y͏ܲwQ1;yarh\Cn^XO��*�[I��,�?�}.�4�up����"�I�b���ĭ�*�&a�K]z��YЅ��!5� K�yB���űc<ϭ��^�;l�L
���kk��} "����6�ՑN<P��yV7�u������$�ꮌ�'SE��"AnR��C��Q_FC7�n�{�_����h�t;�h�IUΐ��`YD���tX�A^}iA�cdtDJ�������vF�i5R;�Sq�R6q����H��֧Ayj������-X�����qW
��Am�خҶ��V�l �QQV���Ҏp�@3�;Mz1�&���>�[�4�ōC����r;'���\�++x���c�8+�)̌& ���TZ�LȽ���4
�l�d��Y&�Z�gh
�iE;�*�Ȉ�@A�c's�A!�G-J�S�
)8rY4��>d+np���)�ag8�I�G��A���K|��(�{�6�	�˔U06���/�TV;"� �m�xf
(u��1T���&��~瓹���0(��MP��RFT &3L�����U�B���6X�C����qt���`�N��]�d�Iu�{ov�w�H�~�h^�}a5�$9,7x���m~ޯ>"��3{�i�"���+��{Gd�z���W�zU5�G�L��:�c��T�_2 �PH���h�[��=ɸ.)�J�OR�|����T�樂��������������"���W] u]�n��%��"oģf��aQx{�2Z�l�)���{� ���UD+	BXu�8T��^�uХ��h��}U��/N�\& ��$����	���I�C$��X����2�A|�ǥ�O��=R�dJ�`��fƚ�"g��J�e6pk~��H���~�OA���t�O\J��O�����}K�~u�n�5�wl\�3��{78�NF��y+r g�����'�D$��q�\+��&\C$�٭�0�HKn�%����MO�~�it�
�P'P������-u[-t(p	�����{��εue��#�ca�ѹA��>1\��3��[G�WfC���Z�a�V�HL$��,/~ӱ���'�:���7B�a���|-��Ȳ��l�K6���yK�u^���8?���@�G�^�?[����v��s�8r�F!�I�$1��5�vۖ`�kW0��9f��$vOGEB��۹��s��{\��Op��+l<��Io/d1�	n��X0���8�(���ˣ#~�����'���֡��t��>?sL!���wɲ�f�ߞ�=� 9����P��� LLi['�n��b��h.M�v��Ċ�cwu�~&A2�O/���9z��G�T�t&%M��U
_��vR�\]��̋���z�aSo��_�A�͟Y߷2��=9������l����w�wA*W0���j�/	(]v��لHGC��Qh�)�'z�!�z�ȵ�TV�Ȼ�CRx��y��ҳ�����]�o!6db(M��4��O�#J�2$�\����*h'-�d9`WQO����X���FU�yӫK;���}!E��&��}����D��]�5(6�h��{ϋ���МJ�Lx��)�Q���r��k`���QB�s�m��C脖=|��`��ѣVG`��V�(?W�)+�"�-�蟅������s5�Z�97��,ǡ����{ʢ�ʫ���6�]�BY���~���ڇ�u���(���pC�%��b���>��M�=죦ʿG�А��	�X`h8o�
�W�L�l+�1���
�7.�<%up<O�>��4K�������);���*��"A z��ٽ�0dU�ߋ����w�\�+����K�gnSA=c�K1tL�PzU�R��6t[����̏C+�M��B�����'L�Kz��q�4M�s� s�#?'���~��Z���p�����!���ƻTW��/w�D������I�,ۭ����॰�A�*�n�t����D��i���z�J�$���Ns����6�^}��,��H�PD�4�c���H�2��z�=����@[Fe�-܏6B}�Yi�V*(�xKp��Ev�G��0�S�I�_Uz���ZD�:n�K�?5�et�gh�VQ�F�;F&�����}��U�������]���AS���rZ�~�dc� �7+��ݚq�^��`��Ěr�Oi� 2��>kĮ��MzgN���n^�~7���m��dߙVwnc�l�+�`J�������#�T��z��~�	�)������*� O�g%
���W�F}�YpjI�C�@���O�8��@���>`mC(T��� H~��g�	���""���F�$�my{�א<����o�S#�h{Qv�V:y�� �vh�d�ղտ���0�x�������倚̏81��-�4����z����j���b�� [3,�Kh��3%���z�J����-�����Ya�j������r��`�(ggm�Q�^܀bˇ۩�^����	aD:��24�H��됌���p �.�w��6��}�!@����qef~K�I�]2�����w��JW��&5�x���_��] @w���o��&(���β��Ժ^*ނy��I�g�v�3YA�/ܿ�h7��.�Ƨ�&��n�C�~����O[ZߵUk��c���0���_�G�����&ש�lU��wr�JaO���C�H2�0[�_S���r��rǸ@>�R@�ÃI~������d����Ϥ���,�ܴKL�+3oE�ܥk\+4�Յct���~���>���Hg�����S����~q��lC��>f�ZD�(��<�`7 ��lͻ5fm�g�[x��v��y U�����y����N��JU/-�*�"�wId�X�i'�n:(�A�׻��`g�˘�؀�r 迆(�Q�]q��ǜ�-:�%v��A,���r��53r5���A��c�&�~c��_sU)��R�:��r�F���d��<���KyNYCć���C�'�� ��f�������,ꕐQ��)��~,Lb�G��(DO ��~��
`S#�/�Ww��]�� t����r���pg���A��$g��j�m�.����7�z�Ѡ$�1��B>�n��x�J�_�jE�T�z���wOg'q�c�`73���p�Z�Ꟗ���O F���RsSfʔ�A��M�{�Q��y�M#n�Bl.~m��,��Q�t&�BڂG���4:���H�h�^&����ԛ|�Á�����R����褐��,'�N��[�y9�ND�P�U3t�C�
YJ$�{��9{�<�J�5s~Z���o<LI�ep�z��E�h��MH-�4	�B�C��ϟ���]�ӲMxA��:&t�dl�jzI�PqY��dF�ה��b�J \\��Hi�W�E�'`)�ر�:��@���s$���{�.�r����&_f�e�b���1�?~�Z#�I�:�@���$�����`����|�"��&�F"��չ�ѹM9�|���gPo���@��.��H1��)�#���齻\��'�՝��{'\1�x���᱈j���j47�����%�9n"^7���_�?e(�6IQ�,����_��R�j���w��{<��	���e�y��*�P���ވ'P[xiez�>���g7�����b�@:�X?�k�p�.�Oy�����I���̻���w��7�q��$�a��j��4��fT�ǈ�qBF�ѝ?EZR�}�p��G��n��6�Щ�c}�L�V�XҶ�����с�t��Y0\�����ܟ������F��#�x��̤&<`JiԪtd&��-~��$�+���f�5���Q��$����-=�i��vp���ڈ�Qj�9�P̡�6��j�L{�<�4�9�B?����J������01�h5�R4�2�|S{�&+z�8b%��,�;�6��/��l�Ѣ���Q���"{i"��2���K�Kg[^LrU<�(�$-���������
)�k+������̡�w����9:����S��A�Vߊ��S@�Hkэafʏ�@3a:��ѭݢ(bS]/p��1g;�A��I:�Dvv�gK��p�M3��d�r4R���p��B�������3�:�d���pr^�I���vΜ,�[n����uخ���&��.z�Ɓ��%#���Vgzl1*�7���E:v}Nl
fD1*/�U5!� 6����z4f��a�E�nm;svJ��f�
��}fr0�2J��}���4
X�I-�j�'�~�����/*���oɔ�#&*� % ��L����h�cm��m�q�PK�Eh$�B֭��k��u�bc�ɪ�+��`���ÃΡ!.����*m�AU2��]����9_8c��d��[ڟ�I#*������OE+	I�[�gG 5B=�.�����]���"!�C��)��l��X�4���a �0�/�����I���Is��Uk~�z�>�V�5�}�rS�j�R�i�1>��,�7�F���h��T��w�	@#h�7���n�7C�͆ؠ�lʓޭ.���6�_2)�4"���L���0.�ۍ1�*BK���<G�h�(g�d1��	�dNB��IF������}^�ߦ�7`���-jB��Ľ;��L/,�|[|!�V`�M�f�(DB��}.���}�!�/�l�W���@o�P�ʁ����w�>�^k�P�97� S06�[�~uHW���v�K�<�r|��U����UZM��Tt�P����ph��e��q�%XJ���B���]�'�>�O�7��_�"�"9^Ð��ߏ05�m��Z�S ��2}�E)d�{���<��cT���&N�SN:�u�W���W��1Ch�w��43�g�;S �$m�>�������Fa���M�.uɧ�H �h�e��i{�r�?Z4@s�.&A�/T)�[�G}K4>��˚L�k{ہ���-c#�1���=���E8y�����gjgF�xt 3x�_��zC��v�\�~�[`��;���M;9rՍ�?bjӤMq����d��%,�q��l@w��9������`�I��� Q���Vӳ������T�R��G��VTUS2��Jvؖ
�b9&^y�=�
��#?�J�Z�������]1�=�4ǔ�f �x��ycɿޚ� ��.v��x�^l:� m�l�᤼��E��_괭�\�_�r������.~�����J�aa|C����k���ؐ�i��*R����a[�]�Fx��;�aǠ�-��~w6'����\�������ܹ�`N�
�b�R>�o���c���H�=\*:�{��SpbZ~�`��55I���+;�+��6�l�|�u�x��,"o����_�X�#�fE�i����LT��w*�*��6�:��Z�Tu�`8T��vM8��=;}5�o
#q/W��y���㓟s�|�zT�Ӱ�%��!�;�)i��/���LvDx���,��]׳�oK�?��"��L'u� �gw�,�65�*��5|�5�d�0�w����iF��jN�뙛�����]O5���-�1�㑆��7O��ie�ZgAڐ�m_6�;WUL�k&�����]7�2�+@"
 �6�պGW-D�aSf9޷�eG��njc��<?���t�)��5�Ϳw�L��e��)��Rf��-
8���v�"��	T��)�vR���Er���Qͦ����K��i4���-��c6�de�PcK\z�}./m A
!�2 !d(q�W�Zu�s�+�'���FY��.Ly�8�~z]������sf��=������t�����]�]���ݞ,�
�[+X+�=�|r���șL�~j��kZ�'�\ܒ�ev�Z{���Xh�� b���ܕ�i�`�`Ed@K~5�Ui@Q��y�.�}�� _��t]l���������h=y�ҤʰM�X�q�<~lPy�X�w$$�v%k��'�3���"iģ�>8�GKM�{PnY�C�tE,�5���?]�Sk;Y�hwQe��q�3l�?@d��?t��	���EO�8��KH�d��]�,�44X��>�\������(@ƚ��M���6]�/�=��ʟ@_I�SN�ANrV����=���T�e� =��2�EDJO��J�X	pW��.Tݳ�n�	u�H�2�S���*خK��G���V�UD��/  a�A��﷼<nW_��u��U�;1�렉?���o�І"��
�@��8t�?���e�CK�����\�<Vb�7��mgf?�'��9�2��>P�ݭ?t�2Q��5o>�����.=���dWM�$$"�4�/3+�o��[sy���cr0t㍵�#ԇ[�\`�Gi��FbrV"�
�F���kϰ�(įx��WG�uȳ)alB���0_E%6r�?�Q��h\�o/ϧ?�v�!��K��>�O�`�v΃��� %n�x5�/���d�])������z���r~�|��,A��D�(l/|��Ft{*��
���y֨� �����`�H�騔�W�|��5v��p�'��ϱ�S�D�^��4O"��9M}�;´k�)���Scii!(�Ņ@u1���?�8.P��C� ?��/��dRJ�#����j2	:V�$	����P3bڤˍ�Q��R�u�7:X]b��u��:!�R�%q���J�4����P_���i��8p�*�2������c6?�V��=W��i�6�<���;�U%��yP�0���K�M�#g>LH�`�}Q�k���a���8M�N��	���?8C���T/���g��R��Y��ՈpX��O���Ngs	o[}��t�@�����!���C^b։�]p>�Uo����-��Nx
P��պ��t�A���B�N�Wwk�v�c�����C��L��\F6���-������^�:ކ��q�Z��!G)Ҧe������&�N�B�$���ߨ킰���z��\� G��e�
�X��Uٍ���jZ\)k%���Y�VY
s�E��尔�L��)t���!�3;� �'�NQ�ђ������Xk�o��X�Sg��0����Kۂ4�L�Y�&9�#���5h��`�������3�U��K�T�����,˸�$�U��'m"v����1R����'j����-�,&��Cr�x����sxa}�TL�~�W6�b1$TI�gX��>���6�I8�2>Q4mU���@��Jo�Y�V�3A�t{��.|�?���6���e&�`}Li�P�vT|�d:�.�.'���2�6޲��9�Px#]��}��7_F@}W���l��F$�p3d���9�v�:S���Z�<xJ��A�w�#�j =0mlC4��z;�����X���ɊcФP�3SH��d�
��;��dU�j�R��	�I�b�KJ9�g����_&9�{4�ʆ���S��=�@�?�;T�;r	���H+ec�MO��t�JW/��	���w��H:�G��=���c�^A�,";8��e�E��\�o��*!����d�;BV���p{��!�~o��,w.7A����(��7C���kp�Jș<�n�8T�lҢgq�WZP� �ݤ��G�|;�ʯ�z5��#"��$k�;�Gy�qh�!O��i��Lʊ.�;�0��Vq�� 꺱�Eԁ��B��5��Eu�e�=��k�ߓk�'A�w��1[_J��":@����r�͏�F��0E5�>�M�XQ���vRH���O���ru��ݱ#�S ��'W�����bF]9��W+����P8V���<��}���|yu��s����c �P�#�X�z��* %w�Hf�����IJ���O�����
g��k��[7�n����E{5ȓ�Z2䃮��]"�~߂Ӏ�!:���7�o�2�y5�Q�At���.���b��������h�"o�+|�ɗ���#��#/g8%6p�L�	ɤ��EaI=0_an>Tޅ~�Hҵ��J�3�B�Q���B �O�VS;Ƣ���/t�&����t񿺼@�W�waͯ���N�]K�і}ߑ��'���vzcY�v�|�'!����C��g���e�>a���voOY8����wSbɴu��UƏ���)!������P��oc�s�������E]B�}r���0D�徧td��]gJ���7~�']V5�ӑaͽ�t�S�m�Q̨=�)�C3�N�ϭC���}S}�����*!� |rcFG�T���Y�v�Q���զ��g��]#��na@�k�\y]�m��m���� ���"E��Ԁ���D�=3e���5���?����&W���w� n�.w�v���;	�Հc"M{sĦ��"����s;��r�wq���}�Umj. r@§��ހ���*@-��=.��<Ш�e�^l�W���e�6r��j��;4�����$���:����	�S�X*HX掘���u����5,�r�L��p��C��r��K���.H�� z��/� $sYt_#�?V,��Nj��Ǵ�k�(��������o	��>��z�/5��T{u��]i������@�t��C�$Xur��x^�y���n>�X����
Ue<I���yowD�b!��jd1X�Ư��qVn��~�&�s:(5?��4ָ<"���&4��$�o�b �3F�g�w�QJ�)1���*h���v�D�O�ևX��ًӤ����6���������j�oUJg�4႐��
�����ƯP2j���'��;����z���3\/ ��:�Bcm��3��C�f���ޯN��oa_���o)�H��f1~��6��3d���<77��s����mk��!?�BC��?���?���V�dIo�j�yV"9����pl�̀��zU/��e�C"=�>�o-��!PW�O���:C�$�]��;�d�g7Y�m�8μp�"��V�x^�\��b��:�-,��a唉V�x�KlH絁��񎱼=�}7�' Yo��C��ƌv���-��3�̏w���ٗ���1���1���_�����(
q�M���I�w��զf�ۿG�b;F��G?7��5O�"�&1��F�)�ѵ���܄���]wQ�c!Di��	5���;�⚚
;x-�PnE�B�a�٧�2�;m�p��Й%��֗�]�n�`�8�l��Q��D��WK݈�`�{������N���G��*���)����B[1���?\R�I�q}4�?�:(�����>`}�:oBK̉��ˠ�ź��Ċ�AU���h�:�B�����|Ƴ��ޘh��KB���7�l�N�W
i��W�5��Q��DQ�d?�&�>Ϛ1�CP��]ҟ��m�&��Ծ�M��{�u��iWѼ8�5ؿ@��)�s�n��/��7B��u��'�:�}�T�:e� 3����'�����e�&�O�(�hf�e�B�f�*e8,9�xS8����<�J&`h(	�k�e��ڮ�'��M�|5Ƅsl_Є�
�Oe�݌P"��U���qWڝ�_�^��,{�1s���a�Z�s�f(��'4١ctr�l�@��@T�&��I�Iw�˄�X�
��'Yu��igF_7��RQC����o=�z[�.S�
y��.��HF�<��e�(A�pP�y�?�L�'��S3TU,T��@��e��?cu���H�|��t�-m�|�2p�՝���Ƿ׳�0q4����r@p��o�����~\g�r`��z ����qQ�m���D��Nr���@�91Jr�W$���������z���(���U��B�t���R�ܣb���A�}��C��T��)�m�)���'�ϵ�-r�#=ꟃQp)���4o�K���+�)��;|G���EU��z)�5����c�V�sW�y�"���aI�����~tRil!����BO���aL3�O���bh�YdԤ�;js6"S�7��G��~G묜a��uj b3�uG1�����n���EEA|dtc����ѽ�s�?�����r (�0�P�����.k��/�t>�!2@Dyv���� �ޥ��������E�xm}��]�o�ĩ��mEn@����%�����Ǵ��\V"�<��MnFJu��������*�y�	a��;�<;��-�	2`@�\B�h����}GA���Q����^��(`U9���\�:b:���O9�0�4*3���mW��cp6g��N|�G����ؓ/V5��p �*�#�Q ����:��+iYF��o �M�r��c����������#SK�p�F�r��+e~6*����<[c�p<������_[�T��PK���3Ѱ����H.6�ϗO2Bw�,���I建gJ�����v«��`���]�8�����}�m�w�7�k+F�!�#Ҁq6zM/���M�`y�NU��r�"���=K�O	*�^��(n�BD]�O��eq�C��H�L���P~eHUb�ٜř4�?�֙;���1�Uu�Cd��%�T��Z�l\w��8�o�KY�+�AZ����$��h�%沘�KM��57[I��ȿ�a=
��"��f����=��Z��A�QZRJ�&m����?`KL`�F��	�}�{æ��kZ�v����4S}I!At�@��P�}<��۪��QY��C�Uz4�-T�_�����t��bT(_杏�+T���K�(��?�S���I5L&�q$�6��M8;*�T`_�}�٣��*��_�S��54CLh���͟)�
�(x�ͩ٦ˇ	��Gi�*�D��ω���xe�~�������oI M�_�rS�'L8���׫��ߎo���/M��F���ҁ�'侈	�X<����:�8w�����y:�V�-�Az��^��|�嗺�zX�b����Aq�٪@&�]`�u�8W-8^�6 m��%��'��P� ��Veh��M�����G�~(Ə�b�x��*�i��5��/g��ņ�?�vj���w~m��]��Zk�b�A�����r��K�c�&&�/��}�I�|�TE]��j�1��>�S�E��u��StȨw�+�,�[��.�g]n~v2~p&{���c�M��8Ġ�9�* ���W�`O�u��n���:~����4z���4�X����l�T�LY �.�V�z�6�� �7އ �������8�U48������e��Ȝ��ǖ�[��~Hf�Wi1Ѽ�NuӅ�����:Y��l� g��ʔ\��ԏ#���gH����]�R0x�g�H�\�ǳ��2\�I�8:�w�gaǧ��E�,�nR.}�u��X��'��l�_-�$Гg�\,��&�֐� �����T-��`α�K՗�!��KQ��L�?�i�ۼV�n��o΋����x��̘�~Pgm�yb�<3�)�{;�i��U6/�`TK�B_<�B� ���{0t��w6�����E�E��m-�%6�LX�5T�0N����Tn�W�����v���	��.��O�H�?w��a.Oy�V�m��oz�G������S��(}Y�j/>2ʻ6	 ����݃���d2ތ���s����Ί.o��t��`��"Z�W�_�������ײ��f����q�����a?bq?݁	�ٹ��r�����LV9��C/���d>�=e9o��Fj���%\�^?��,g��|fB
�"Q�:�+�@
Ҝ����L���>TU]���.�����F�ʞ-��9�=��}2!���nI�:L��lTl!�%)�����?�ͷ����/��C5:u𫣧J�fP��~˘� \h�-����m�Y�R��"�M������0��=�{���//��qK�MD�ѧ�*�^XBQ�����0?�az?�n������"b���Cܨ�=/�}-h�CD9�<wf���iD
� �
����`�)��D�/}�K�#B�ͻ��V��U��eU�C�*�p5�5
��2 ��w��C(��0f�����d��zp��Eom�n�-؈����C�\�A[+h��\�צ��EWS:3{*�rg`*Q�ٴX沆j�}+�ݦ�g�<�3>~|d���I׊��ѫ�8fc��D��^H"� �OT_�M^ݾ���8U[���?���F���B�
M) �ģ�殖��zģN:�W���:έ%�h:�ez�=��ɖ�"N_��~��"ݧQ�o��O��E�" Y��1h-!���亯�q[�n =.��|<P"�5У����8M2\���g���@��@{�9UP���	j�5Dl���no.�/��#<��r�<G��?X��O��I��
�6K�mvI�9W���$M �A�$����� ��>>�h�HO��N'��;8��8���7A��z6oh��x��X]����w%� )E�L�ݣG�?�r9�1�4'RoQ6|���V�LH��66�؆�����H]�)��8��n^ϖ�J�_�e2 ����GY�;��r��8HZi�����S���]������ ��K	M���	th��g/;fV����v}*�lVB�-�r�"�F�U�
���k�	r��o����jE�H���ޥ��n�y�iC�%����q��;ӆ�mB���y~&��7��>�=&"��K���f��˪�q	K,���E�?$e���l�eڱ�r���c2p�<A���B�@7�A����ӱ).����@��`�ܽfnn���pĘ�0f�P^ٻ�
����I�� i��9��2ޞc�g�K
����2`ls&ꐽ��bx4������M�_�FYU}�[��	��d�-�j�jPJ�\���wB�Q�F}�Z7DHJ�͠x���A�Ĥ�G�A_��,�buqp����LP�Q�y?�:�S�ɑ��I:���L��0ny����5i�-����ձ�J�Yq9��i�R�]!��5��uŇ$��G���L�
Koz ���f���J%�NV����YT��	������/��͊��5�	�pǒ�����ݕ��ؘ�o�����b�k7H�+�e���ڽG_��\��T&ά�?�S�F}�b��'�������8��McL�����WB�=?���6
�u��C��������ǭ�L�-�P���v���6�?��͏6�F�NI���Ο�fb{O}7��@�T�}]��M������܍j��˘IB�w���+
N��F	��	�Yt�p�TO5G�7ygJƄx��@���X�GMd�X��l����� ����ዜJI�U��u�v�	�O�C���Kqd���3�|����'�s��^��9-S=9h�H�߃���f'�6&'MP��E?���-+�a�l �җ|{�X���yM��V�*�*1k���K���dv �|��k�a���U����?���.��I�D=W����������]�A��̇����f�@k��ey�]�"ExN�� �B[����g⃈���=�(P/ɾ
^���8�+�7��q���\�z�Mk���9�Nqb�2I���c� ��+JI������~)u%Ű����a���F�5�%Q�@ؑ�Ů�@�;͚�Cw�Kե@���c.-�8��'a4t�k~\�v$�*�O��D~��z@ġ0��-d�� �h�2��g!�����ғ��_��}�a�
	��zxܡ;ի��-�ߤ&�'�\wAL��щ�dk�Ɏ^�lX�t���$ �ղ�L�ޟ`�7cb���݄4����P�_eH�3�Ҟ�W�懗 �Vd�ǂ�Dh��c*�!h[δ��f�&�V��}�<dE"g�3�����4q�a�RZ�lіK����t�au���A��pBʘ��橱��������R5��AB&β���a�.���/-��i��h�VH>ݶpӠ13}4L<�2��M|h��������"rƙ�̞
~���Y߿�Gc���*>(�0�� (ĿD������_�`*]�7�5�A[��pк:�پb�G��B!�9��[�Jj�#^|���u�$-1Y�Z6�5�9���ж���]F�[����	8|X�.OV v)c#n[]݀hM�pw���0ĳ��H��PN����j�S���t�D�RjŶn�I�:��Z���a�5�0]^� �5(�z��f�x�@��L�c�[zG��2����Fk%Yc�"SofZ�B�L��)��X2����2��c�D�K�c���<�%�&��C�l1[.�6-�d�Lu�N���?[�0l�~�j��&�(�'o���qYsPrh���J�/��n�K�^�+���1үIG\C<;DV�n؈/ʆQ��'�nu��>�!�����էi��m��>Ԁw./�g�G�{�he�K��*�^	��3(�Q�A�ϙ9�[%���!�J��m�eM���BE%�7h�o0r��xx��m)�ٙHa��̰��)�+�W�)T�o����h��^yo�ĽP�Q�
�ҹ�;�{�}�$�#�\;��vF��XT��~]`��ai��}�^.z�oI�r�'��U�(gf���4+�v�8�9ي{͞���\���I�`������i�r�wd�P�/���d�e�@�y$pj,�Zf�k5v���7$1�x�<y�]L]1��\f�˲:���.�B۸��f6�C���xi%�kxc����r�Lm����1�x�:	�.H���UY�q`V��%��ԣdֺ������s,xB�=�M��J������/�dﴗ��^�TFO�"4ߠ�a1cں��=3T)ϫ�P��l�Bc�+e��vΆt���P�ɶZm��yE���M�B�N v����4?m�qϦ�l�)A�@���H��tk�p��(��:Za�S�hɴޖ�y�;	�{���P�.Jި���#�ݐQ�e����&�F_� V�\e�T��J��+�:��2�{^aN�|����*�������"@�=Ԕ������eqh��x@oMKS�|T�RL�$&�I�Zf@{AR>@kD!��J:~>mx�A8�r|!g�q���Af�o�������##Zjf>�Q=����\GK�@ut�p�ga6��}��=q���J-��]"o�:�!�;K��.�+s��wYm|������aO�ޫ�$�?�Nse�R�5�3ύI$������A�HlC�{{�Q~��MwCZˬ���_�43�6p�A
1�pXeQ�~�+(^�b�}�"�:��z0i7��r��g���vS��3� �4�����q�}�ie3�h�:�Pe���������j9���S1��(1��QÛ���O��k/kV+�;�i���{Fm�x�:v�T:*��U�9�[<�^m?&e]_�x�%�lU"M�)_܉�/�Ջ��9�2.!���y(�;r�x�a;#�ng����H_ub�>6hcܔ�=? ��`�t���$f�=Ö ��6�E���ƹ�Tv�(����
T]1�9�C"�&�6#D�[�	��EҧR�^5c�*�'	�>G�|H�Ge�6���+t�U.�3'��_�%A�p�lm�z�¦
������<��ƶ@;�u;��tѫ�L+\�%��2hR���������eD��<�%����ے�_��2���NP����x���������q�{�6�.�1e�� �T N�D�PCS&��Oy�{�G�o�M���:�{���U�M�UK�#�j�N�R/c̑d�'
׾��3���?�>��ᢡ�7FUW�W�J}�M.�,�+1����}��;���3JI!.��7 �*���=o�Gl�U�JC�a@D�Nii�M �j���ߴ��ݵeE��"p�Ey7��S���e�jI����CE����Ф����.��F&�����B"zL$/��<[$L^���'u�G�n����:���E���FV�[M���ļG���,x���c}z6�1<Y�=_^νO���V�;����i�K�9pҨA!�c�Ia�!C�jp�Z� ���&<�;�2BP(����Iӧ
H�I
.�)��j`����҄j$��z�M�h����\�i�	�!��:��b%��3��/��LK8��G`��P�\�v����|��[r �Gp���OU0�J�"L�+��+`8E����L����j��2[[���íR�ڮ{HgN�U���/� �S�F�j�}
.	U1�%{�+����IO`6vP �L��*�E�-����z~Y4���$�'��l-�T Wz@_/�[ΨOĦlSWxqS��l�Ս-n���ӎ45�=��B���]�r�/�����{�#9��ب�4.�Ա�����6�6q�Vp��,�1S�߼Ɉ�em4̣��^:�uz��ƣlY�O`g��ط�j�Xi&�L�܀�ڽ�YlO���x�ۡḥ���d\�Y��2J�� @�E_�Z�q�vYWSj���1�{��F��$2�ɣ�~���Wʞ��*�IX"�`��b���L+��(��˅_�6F�粦�J��y�7���ns��I� Evc���sU�<�h��Z	b����R�O_�`�$����6��������
�+D�Î]H�y��~O��r���ސ3z\��ϊp�J�T��_6w����ׂY��>�C�Y{������F~��-Up���?���3�u��ef�]�]H%��?FwqΌW7\[/�WaD��%=<��q}{�'�?Y{�x��$�X��e'"���.h�G|:o�=��� lrn� �?�>��wC�Qv��r��Q� ��#�ؽ����@�����VY�;b����vsQ���B܉�r�9k��7�F��u�`R�� ���_ҽhW��;���G���f���aä:MN�+�������଻O}�,����S��)�0�t��]-.ۃ�A��#�S��X�pQw�C��1ڽr�v@�Ԡ��9a��ㆧ�AH�P�MҖNf<noI*��y�f��RF�@�{�w�p��(9m���3D�K‘�W����rٞ�T�v_�a ���'>M+`ifI�����TS�IJ���~��5�����Ȩ2�������_��U�H��Rϧ-�s�>�NiZ�*��,�2�qi�mXW��sZˋ��x�w���Aɘ����C���m��N�>x�V�
�*�0��x9=?���좡��gy����s>���4�	@�]�x��jcn)Kߕy<T�я�6�<��̧=/	a����ΓT�/��� �#� %��φ���[��æ���ID�0�؆�·H�Ɗ6?h]�`l��p>֟ɟ�䰲̮7,��64����[\a�ς���:0��F��$I�񺞴�n�� ��Vʛ���p�ݽ��WI�S�Y�[�U3-������O���tIsԛ�ŝT��k��dx_QL� Z�QK��4}���4<��4�|�p�a�N���F��4���D94|B�fl��^����?`z_�7А�Y/�؆��E��\չ�t#��d<��I��/C��K����/]�'�ï��x3�9��l�z�R��|t�q�/�Ae�3�8�}��g8`Ym��h�S{t�Ф8h8.pƏ0�6j�d�v{�4�_M��y�<xS����?vwJ;) g�S/NHc�o5�#���y��[#�Y��4����ʽ���{����{��.�������SKQ«Pׄ��F �8ŤS�F-���e8sc�C�ߝ�a��NImh�>�{ؗ,��GFXޢZ�u��㲔������)s�o� 4��Q���E�S����b���C�:����{��{��,����xNl�ek�A�
�`Ϝav)5�J�����ϩq�{�a��"O�`�-�M�6;!C���:��Ǉ��Nt$8�c�О��66�ۤ3�% W=�?�_s-���"]��@���O��=ֆqse�[�v}��ig�.�u���5tϤ|࢓>�b^��h�I���WW93��{��hs�/�.�IYE����7uH��@��:�;��C�(Z5���"�:6S��%iy���*�������H������p �y*$�i��.+Ty���;7�1沐�IƔ��Lo�m{�"nФ�˷�n.�`���7�h�ST�}��%��^��Z���FӸxt�*����Z:���9�"���}�������mm�ۗ����,xɦ-�*�T�ϣ�*���2Fz����6B��B���vZU'�d�5T�~-�(X��%�G���!S�
W� �w#�Ѣd��s�&_kZ-뗃���&0�M�%�d(����'����2�j ��W�}�m��%�[�����U��j
�`U�(�b9-.+pY�׮�y�$��1Q�>L��Q��PFS�7�{|�yz�F{��i7|�&F�زoxY��څƕŋ$�)QhOVo��E<�av�T�EC�'5CM�^=&&���Y�Xyl�|Qw�{nPxƨ�0 9�~����i�N?��V)����N@f۰�k��?Z@c��n�V�wk��Ġb6x�eT{]�8p,q���[t&����l�,J[��3��3�����/pv�3 �Hh/Ғ�((�hϭl�(H���B�E�a�$�r�� �t5?5��?�>�ױl�������p���	8� ���E�&�*i����3�h�~ד�r��1N؞
���%Cu�L��f*k "�'��v�:*��Zơ������[=���?:4�>k/C\��/{q�r�.���y`g���Mm��l�ÝGӷS�/�����ڶ��	�]ƭ�z�3upx}8A�����'&.$F#�_�Y�q?ӌ�QQ��q���uu~�r������1ܙA��Kf��>��,���aE��/��cx��(,����A&�:�P45	fȜzk�!�K&/1���ԫ"ʇJ�����$4p��r'�b�XO�24Q~c��鳭�fp��b/kJ�+U��������L��Ef.�Sc^�����T�K#�nl��ͻ����_�а�nJʁ3|]}��82���磊�BϾ��Լ��f�7Z�ђ�����?�ֽS6�}c'�Z�R�XEx/����uD;�L��:�|t���W�_��4ee*����%e�=�����S湴,��o���5%�`ݯ�I@9i��!z�,�ܷ4��*>|a%e�f��bB�y�@�'],r8�./��$C�*Q�����n��,��Cݠ�A9���g�e�I���t�T.��#3�Ƕ�,V=J&S�t�Znw��ŉ�yu�3��+�����69L�R�
��m��.W5��ǖR���,��R�ߪ͍�s���ͧe��aw��� 3;�AF��ݼ�Jn�k"�<��/U�I�!�������DZR7?��]�m`�N���Q8��4���z�����Xq04҇/*nk�|�gg�Ѽ��R�����+F4H�;>��Ύ���F�VSv���eR����>�ؑV�KA)LШQ�~���3�Q�U�^g�2�u��	�N^O��RH+�#��%|�͜�aa��xI��a�N�E X�]�RH�����.fa�*�)�8���7ѻb֡ȁ%I�k��MD�~*O�q�׈hѸn��
�Ó���33���25<啰���������2,�<���V�0�ݔ�w���a�ơF&��{�$�� ��R�@�B�T��T��(��y�=�}0&�ͤ?U���ۢ�U8��o�m7��s�����B�>�I���k︀͖��;WK���K@��=����_]0�8�}?��TN����oXХ5e?c�b�x�[Aw�K�c��=�:�`��L���R����+��j�c���GY@����>�݃�cL}�Y?����B����j�zE%���!>bUe������w��lSPw��_T*��E�F�y�sA��d�/����M�&^V,�:9θ�Dh��&��jJ�qߎIy#u��#����	�Ƣ���F���j���hF|����������H�?U��i3VOT��p�m�wG��m��PIR~��k)���ne-_!�j�,T�����e�Ό����(�^jB�?Ytֳ�YR�tl1��tn�G��d�'��
��l@Z���Dje~�d*��Yb��S��P�b&�y�D[��w hpG�~��ȷ�� ����R+�R&3�O%���@��TG����ъȈ���.���W��f�@�0Xu"����A�F-���������ljS�x��74O˕\th���	��?Q��eD�0X��.��it�|�}[��?)=�.H���Ht��w���]h�$a	Q���ǭG�;�l�Rs(�9�A/�Z�>_g�+6t4�s�����﷝7��چJEyRWgh������ܮ�yO�f8���ͺ[ڥaӈ%�l75�T{�����G�aY2Nb�FqG �����]U����ٓ�*2ڐ��u���'a�In����9Uy2BKPˣ2�����j��ٛ��nl�����=f��r�W��]rhp�!>��
rt}��KI��k!���|$�T�n{��������䐮G��_g�gD���3\�;��zĝ��c��b��0<q�L�����Y !�`�e����a{� Xk�\(��ը��T!�#��݊%hLC5�<���衉���/F<�o仞�F�C���e�:�P,�O�wk[e�%�}zd/Ն�M��3�Ql���)��OQ���̐��ɟF��a���;�� ��3ü^⇋W�Z0¢D}��C'�"��r�W@$Є˯���=�v;�Q$pE��m��sL���s�-�L���/éy�/�a�!��2�w)xx�$���1b�t�5��2Q��8)*B� �o�"aU2١�Z1� ��kv-~�a��05skH;����0��W?��l��䵍�Y�p�i��ʚ�`���ņ8g�&4Ш��1w�qT�c��ܲ�S��ϯR�w���fEF4����~HkMո�晊��t藮�r��
�Ƚ�u4�c����!�s���0%48Km���`�YW�A��l�4��<g모���
:��W��@�^b$�^�XK��l��L��y���53�\��ЊCD�6�UAGg��BG��d���R����כ���f.����(����MA�34��,ݡ���[!�b4�t�b���3z�S��MF��1��·��f�� ��*��K�3=�U]&I�=:C4 QZ"��za��T(�N1�o�ȉR\e}m[�B_J��[�O���<-p�Ϗ��+3wQ��|��=��ˈ~���Z)�,��u_`�S:TG��ґ)�A�fg�:d4�� Ʋޘ5;S���~KR,��a��.�����T*�=�����������XZ'�p�|��q����5��!��VX�dվ��z(8��q��8������Cԅ�(~����g�L���@J>/o.�-���������� �V�6�ӥV�V���{����!D�:;|=�,i�����xNz�Z#p���O�
u��z(Ŀ��gZ�N�	�{���8��/d4���+�nc���	������{�{�+��Mz6V\�^���2����bZ��F���b����p��g��$!1J;6~Y2Xz�p�&����]I3��jp�J/d�7k�q�u�A��fYT��l3�N���fw{�V�K�����H�B����5���*�X�:���d�WC�Wt��}jx��XS��a���`�}�_����n;l��{�m%x��/�,1{}TV��SC��oAh��4�=�9���AZnu'���!����r^���wǅ��������&n�l���a���N@{�`�#���~��z����g��Y�[��$4_� �W@-Di����T%L��g� �Ø*k���� r'.��D��!QC��25��X\�c���1u�]Y�BO�E�ɀbEJ��[?�M����;.ԫ�*V��xt�\���o���rO�p�5~L!��UZ܇$���C/��}���an���}�a�T�(�?'�gzF�l/�-�F��9�l�w�*wWȊn��
\/��������{n����#����:ET��vP4��� �ʉ'� �<�� N�G�+�07 �W�X^a���]�d�'jia/���?j��DM�ݓ�ʉZ� �^T���g�i�iH���p�o-c���1�XD$��k*��<�1�z�|�L��)LZh�]M�EG�/�>6���`sX
6�(b�%RF���j�jy�T.Ɯ���:�"�.Kfac�9�i+�456��8V)`��Tٖ�@���V]R,��Q�p���^��^VU�2Y9L�i�qx����P���>P:u�ꐗP�0ɸ�}c+���z���iqVL�`!��: P�AZ�wNI��P~�&���QC�`���&�A�ȩ�Ӣ�;��,��Z+=���&"���"y�J�r�f��ܓ�A��¡�3n�h]!�>��a��5BZ_1��i��oR&=��dO�Iص��/��k�+q "Aэ���59��U�|^Q��̋.�,�<&y1�!_v�K9��k닗��h��2�_�gT�K'9b8�Yex� d�Qm,���wfR"��ӤS�)���� ����슇�d����?YϺ�N-���k%���Q��/b%�����NF1�_�8o�g�c�!��wB�0jG��>[e;c�A��p�M�K�x�}�	��m��Mʏ��֔#AwAG6m�]moT�^����fmv;��`���U��ʁ���t<<�s�P�)�|zЎa$	W�4?`����� y|����!Ɉ'm�����2C`Y�b�BS��+�b�
������?vz�n�T��`pP����j��#�G��t���w�[�G��O�����P�������C��1���"�%�Ȍ4p�<9@*TG2sdiY�8�ث}��O���;ʜ�) ���`��tb9��kM����f��]�}��)��� �Jm�-��`F°�4��ȹ������X/��[������I>���Y	x~ ����ǅ���MA
p��"�'���je�6T��낄�Z��u�0�bW,P'e��^��� 7��xȦw������i�n'� ��"�Մ��oѸSM����ooI�G Y���b�����o�ԉ�Eʭ�
V3�#���Wݹ8��.������b�ޥX;e(�����T��f)��椻�� ���.�rQ<���M��Y aQ�,|A~=x�N�9O Vnk�+n����U�fs���cT���`#$<�8>�/�4��9Zoha7D���o�g��{�rw����8����:�O|�~���F��=��qb��3��B� H���)yj1q֧����y@���h��sm����kj��`��)\qV�f�S�d�e_:�+����+^�+��� �����7~,������Z̹��ZL�HW�
�M�֨�5؋���d�<$���ys?@l��D��G,.H�6�"@Hu��y�.{=9�������\����^ĤIN��N�J��P[/�H���G�S] t��%�sq�IK��S���T%�.��hF �Q=A�_�K!�'	���U��`9 Ox���% �j��t�[׼��Zk��=7���
j"�N/��Q�v!�y�>(�-Q]'�DR��.Yv_�;���>�/�EQ}�'�]��9q��G�TdF�qn�d����>8��L�{Q��Ρ=�Wd�C���zۨ�S�~�@V%7�;b�Pi2O�G.�Q�C�����n ���;�B�f}:����7�.�A���`I�J_�=TXF���0�J�8�n�L�U����mCIRO���W¶�<��ЃLQܘ�bѓ�t�ԧL�d"��@���(���^Lņ~ak\#LȔ�o�멓is,��ayv�<7�25/������5���;ݍX��m�|5����ǿ���${}Mlm�]�E�1mIvf���pf��ڹ�N���N�D��P�A���u�Q�s۰(+.M>�x��2d�H�u���'FO�zܞ�B��x�'&�A D^N���W3������J��5$��T�Ķ�����>&٪A��dԲ��N.�d:�'�q��F-j,^���T���B���D8o���&n��� @��5V�����W�;3����Дd�)C݀��׌����!{��L*�RR�A��9l�\bC=B���cĥ��O��r���E���&��|���Y�1���\g#��҅��0*��	�ӽ{ɓ���$�60E}n��O�9��LI�"��������Ur�Bsl0�I�����eZv�x��q�h�(6�B0�^�s��u�E�$�kS^a��{���c驔� ҁӳԵ�?^W��<�גM�8�;wR9��ek�{� "�2������s�����Y����g�� ��M���{0� Q��t5�����v�.B���z{SQ�Q����fE�ח�'0���}*��w�1�H��(�g1I1��Gh��p�2�d�Ƴ��g�Al�b���gv(��D�f������B��ò���/�?9]6A����V�c�H'��6X4Yt�<�B樹�W*���P���{A�z?p*�/��/*�}%��:G��3�A�)�~��<����5�oVS�1����ݜ�73�A�+��Y{Kn���7���_D7t�&�k'�A}
U�۠�҆��6�H?z.��^{M��B��=�M%��O��D��	 �\R/�k7`�L	_���f�yɱ{@~��ca�î�M��L2��5ݦ���<;���>��|U����'I�(�֚�sƘ��Gs� Kd�BI�!�xb��5é������������l4e�z
��(oW�>:�۔�iC�)I��:�|~o<�ٷx���#	�ϥ��X��e7��Oc_��u�b������{��[f2���]����=R���0~���S��	�v�Pe�&ZTad���� 9>�<}r�`���n�Y{�{��b^�`��� 	���	n�=ɺ�~��������"�2\N���t&�}$�Ha�� �-���s�Ǯ��Нvn?�yد<ZZ��ҵ�c���� �&��[ �B���Yoξʔ�����O��M�!ew����=�%�a�/q�oU�Y8S�K�n]���fc�O׭r��7�N`L��2R8������L�ݥ�@�qך�+ܱ]�}�OU��W~v�0�*��v��*D�����g�62D6!\�BP�����%.��׹QPs�Ԑ���J�j��j��{3cĐ�Mk���u�T�y����W{�8P�$Ei���c@&������N��X{=��U�;�M�ω�nnK�E3�ć%���22�c�VE`!��S]����"h���a��x��f��#�o׎b]Lu,�f��t��Pt^���^ޮb+�m� �9�-��*&Sl��^ F�t��X���XT�D�z-,y73ܩkv�twO?�)�_��,�BW�F��rU�QQ=��X�c-�-[����̳�=�m�)W�g%x�H~*:�2!�-���'�Y4���#a�C��7'O@�'�i̺Ck�y��c$�h���'F��%@Lt���g�GûiA$Ì��%%���ѿ)���/��Jp���Ȕy��ͦr[U�f2Rڟ���바���d�/K(�	�VC*�Ip�]"��lS,Ϣؚ|�Ϥ��΢��i��E�}6N�n�r��u��yA�ݎ�uv��z2{���ב.���O��:�l���T������ˠř��H .�+�,��8�q����وу'>��n�CU�첚��]����v�F����~<�x__��ҹa��Cѓ�C9�n� %�0>��G��8�u��zdK~�%��2����{w�]�/	�/V���SpYU��ج�T&�n&���a%�����b ��^ܬ?�珩q{��(0�������4���k5�cpe�����4!����Q����d������,�N�BSK��>uWS5��� 6ƻ�ȧ"�yva!E��n*�X%�@~gĶmu���rb8��h�P���m4�}�� ���؆p^91�r9ȗ��K�#_'i��|<\UQ��[{tU1���K*@��:�c�b����J�ǦjV�:�o�R�N�q�y�����Q�h��ӓQ ���׏?�.5C!�NQeH��}(g��T�7�|��F�),��MJܲ8���W�B����}qJ!䣝BS�����f���,���ī��í'	�zj���Y���v �DR|�i)VQTrq�Z7�v�~D+�E�;�t�b~i� �.+�u|\�������ܯ��Jn�<
X�i�hkD�L�Ы�7f=b����<���X������9%K[m���83�ٵ�����t�E@:(�H>���B�!�����ߐ�lZ��s�H���&g�O��.@�2��ۭND�,ۅ6eT������`���Βi��J�� l/i���Cs�_m���T���ޏ12F�z�GѴ94��*��a�3 OW�3�3H�a�!���O�,�XI,��듒�[US���s��C�rY�5��C��`���}��"r�L';l�}=�����/�j'"������H������NnS���Q ���DyGC{N�n��7�P�.�`}ʔ�")���T(�/���M )nK1r��q�|�q���n�Dd��PV��ٌ�Ŗ��p��UK$��Q&���T���R�^o�kO���5h�Q�32@�	�)��{�nm]u
��p�TѤ�*���N��:)7S�f�AZ��k���	N���.7��O�1����Ƀ�Ji��\b���^+z��7�^f����b-f;#8���P�a�<�|�� <P�U&煈�ĕ-��8�͠� #=f����*�ܙ�W3�>�61��m�Ԡ�\2�����Ž��+�6��SGC���c�`�Oy�⤎fR�y�� �|\�����
ߜ�IC���Y?`��Ͻ$�}8��_'&lA=�	���m�ͺ�<�C���`�]�˳��T$��o
�s���6�G'�����k�Z�P��.�lutE��y[ba?�^��y�s	�1�'�@�I�}{/�Ds���3�0�\gn���|7	��/� p���=0u��`�E�7�o�P�Mz/�V켃��W ��������ޥ-)hw,����`��̠�b+M6�YѼK�Xo�[d_	XF�*����o��8�v�? �e��}��CZ�]\W��d�<�iR`�l�c��jU�@;E]�>-l�=��2��J������ޕc��o^�t����5����:�|q���w�D����y����w�U�"x#��k�G[���o�`���$�)V���y�Y�"��E�0d�8K;fUK#��M�/-/��1�;��/�������W|�Փ�Ǜ�)�8ݰ?��"��\�7�1(ZDeL;!�v���Xn<������軽G�y��jE��lg��8~b��b^���s�P*C�Q�ۇ��0r�U�����2���<y[���h�.�E�](�x��{��HC*6�\� 7�A����O�6I��ks�`-p6���ThM+eO<Kb�'�[���hO���͚
n��N{�Uh��}���nQ�9E��uL�����>�v�,��c��]*�1u��W�05r�������{B��yt�E����8b�,��� �k����t�e��T
��l~�l��/��g)���_�
B6d��G[ev���P+�W�n$�n�=T�����Y�\�T��p�U���#4��0�ŉK��ݍ�Cfۙm �&�CqKPy���� ~�u
6j��?�v�)���������6�M|�7��,$��K��U<�a��ג���ǉ���t܀s�n�H-s~1v��!��N��O�{FY�������9�7(�,�W�颜R����ZG]��3�JKa3[z����������G-^��O���G�ް���(Ɩ�~���]��+�A©���p��wF{C�F�dLl�Z�$U͏B3�c��q�:��ߏ��	��+@b�����9��[�,z��+m�a[�}5�|�&ͣkn��4!u����APs��"���c�����.zEsep��e��1G�l��ou��_�S�9v!H�x�Qa�?�J��A�c8�Ͻ���T�h ɛU-0�,�g�O�!h��j�{k9�=���� ����	 8�T�tp���wK*���������m�#����7��BK��ki�U��+��S���1Za�kW���2�<��\����`;�$m}G���<�K�P�o�c+�Z�x�.3�KUL"M���mYa�B��0��r�M�L�=�*��#����o��z��:�T�'ή��&��;
2��N�<�L����8ѱm �.J|{�l12����^MR�%�YN��V?�~>6���)�o�Ɓd���/�Q9�k`�K��A5w�u�C�n��J�v[ڪ�������J��OÆ@{+�y{T^��� �C��JMQ�������D+N�G=��9�m��ٕAi^�13�'D]1|_����bw�++d��978J�N��=��K��k�5kUU|Fs�=�P �'
AE���꒤ra�����y�U���c���.
�NAQY+0]�&7uз$������%+mY�Ak��db�Gf�I�5<4���Y�J����#��:.^ŷ��U���ʴo��!�:D��~�?
�|maB�����|�4��s虬G�H�L�_	���~τe۱�N�[@��m�J��m��9A1  �!�V�u��D�-bVTW
��G<�ݗ�T�J5#�m��1	!��O4����E�����>Gmͼ�D1��:.>��Y�_��"Ⱥ�����4�W5�U�XD�����3�)������/ã�Np�ק�a�	�N����i��"�7Y�Fp���M3e�y��W�߂����F��[GeE$w��*�Aug?~E��Q����V|�P�����Yma �������ݿ���O��N�ҿ'_8�ɵ���w@�^��^��~�c�f�8wYl���Fb�~���&��63�J\N�H7����^�,�3A�K[X�	��X%u �Ѽ�7p@Y�Wm�͌��E#6��O_>Љs�yrn���6�>x袶�U���{�Q�1�!��~�0�5�	�6���4˚��ç���ܳ�DM�Hk��kȴ֣1V���`��^�kk��]�ml�R�B9�6���Y��z�ww���)��_{ZWT2!<[�}��TXh4�2	5�jO����Δ)��G@���X]�/�⣧��5�t�f�Ō��;ɪ�D��r�q�o�W��b�� Pن/���	dW봌9�����4�1�)r��s]L0��6l�����p)q��5 �Y�[�J���s��Y��{J��!�͟Q���sr*@J��!��"x�DڭJ1<�:�6Q�H���n�G��C˸���N%��@=�c�"���t4�����x������q%�r��8b�R�!lx���V�Ă�YyvwM҂f�0��%�����7s�G�)�=8Y{�A�+���O �����}r굼9��p'­_ZJ� ��X����G�6��r)p �d�rT�3%�R�S�?�h/���(x�L�U���������"
��c3�)DC~i��QS �ø1��QY����
? �9x[<F%�o�<�0�~r�̎� 3"B
L'7��Uv��H�Z�0zH$�f�"�z�1
yp�u��(�NN�~�>���Zfxm@AD�9�%�w8RK��xo@�5�#_���]�����$����+�_�?wZ��EN�w�����{X���$�y� �OW��'���!Fh
�y���n�Z �c��v_��n�ɈKn8�Lg������l3j�KT��c�xZ�]��дǍ��u�u����N�xq�<�)A|���{�L*��d��:�J�ݕ���N������}�D1����]�e8r�m�,��-����W�(tb+�hRT�C�T���dY�3.��:���Y�ޯ�ɡ0<63�9�d7>/k'��M�q�0D�(r�;�A���ݽ�6M��'� ^*��Q��o'W%7�}����_�h.�7b|�`��j�)��5�p\�>�t��F�2��V\i� gv�!��Ť{7�7�D8�3�Y��Vf\��4v��N�e�,iܒ{� 2t�i�%�t�'2��o�1����qE$�-�����A��țH{U١�d��������恚s氶8<���j���P��� �5��]Ι�|K��?0�T!{�ɧE�7/(�k����ڹA��{okF*���ʋ:/	�����7Aa7�X��	7O���;�h���O��\��-�\��A-�-���\ ɥZa2���|�4���l�Qt�X�ي���w��0B���P'��=��M*�b�iA���3X�lC���)uZ����Z�C�b������(]��J��V6[�~��*�7��O��gX�9�#��9ę8@�Auі �5�U4Vr�J�L�[�D��~4х��sPga��i�װ�{/p��+�Uz��ϕ�v��
@d��߻���I�U�J������Ǹ��0��V�WC!ҫ��r�tİ�֙<�������A������&���$��cHG0�(��]�/�� �[��V�-��]�e���}xHx���Z�a�*�����1o{ʦ:x}���v.�������d�y��j3�#�����N��W�?O`@~�r�N4p�f�A`31�;��.C۾��)g���L}��T�=�?K*}tm�˗�$+�ZS��d�w��������F���r~�-��FCێt��N���-lCG�YqL�"���xh� i������I@o���y_�x��%���\0��&� �a:򔶿Ԑ�n�ٍ��0���x���X�XP$Ɨ���,H���@���J�r�1����N~�a� ��"Z��D�*�ꋷ��7_�9���oe^��h��<ޡ���|�M����Ȗ�1�`��M'��S���l�b��(��>S׺�(R���;�4��Jeu�r��a���uA�fۭ�y`��e�Z8r<�l�Ď��̋�+��n3 	ՙ�����wS)�̦RL5kY,�+z�_����h��-_}��	Δ��xO:<3|��}���N	!��� �����m}���?piP�J,���ޜCq	���@���K��}�y6�$�	*�g���鿳�^��"����.�C�P��㮙|����N:��Ωz��lb���(���/��vX'K�{e�tq���� +/�?p��c�$����^������~rd�I	�j@fk>�ٯ�G��t��Ć4<3_Џ�ޔ��۫�H?�f.k��_�~G��ͦո��n�_n���鼐��Y�z�ύ���HҞ)�ݩ�0�,a_2i��Rp�C�/����ć7�"��+dv��>��$T���AKu}Sa+E����PBJ�zW� e$�wV�p���+FP@E���b$�K�Zo=N�%%�4I������y��^�x�s^�%��q`/�e�"���?_M,t!ё��x,���!娦he

g��蝌����;; ����1��8��>���6�Fz�)�9%�=a�*���d�&A���k�]yÀ����'AoF~�OE�w�~/��s��䚽pP�d�Z'��g�!e��"�<V�5�;l �j��wp��m�h���/i�k�F2�nV�ܦ�������r[�.�����gre�4u۶ɜ�Nh�&wz1�\��􊦊[WZ���8n�)�C/���!�*|�kR�8��������Ȯs�<[�AY��;��c��[��N�#J���
;��xL����s�*X������Y��J@��sl�$�e�F�������l_��Sq�EGyH�h�_B>�D�}?� �\(���?U#��Cw�6}�B��x���i�̂�Ѥ���AP/�#���B��a:�y��:��*�C&Gg���2@�O�����"}XR�][������2Q�/��6E�{��^�9�yVټ�"��O� 2�`HY��xcDj�p6�ݰ>��~�ݨj(�I
�:���e�!� �W�I�b?���=Ƙ)K9�lK�Ir2a��fUd��
~Ө[���ڕ�'���(�}2�-.��б���A8��x���+`�b�Ӥ��̈́ŝ��&|�/� ����i�oX �M�A�U�Re�8��@�O����SL6�I���[�
NQj��W�j�����S6}\�lk��W����J���{Ǳ�=� e�Z�m��s&nJdU�ϡ�E�H�r���-�H�ګ�R�/^�W���W'�a���F v�K$o��S��մW�r�����T��@\�|��V_���n0�d�WF(H���ܢ�i�׺��Ǯ������s����Mb�Y�F;�(�y[��~]#��Rb�p���z:��[ۤ�r�:�Yc�M�ӳ�p
Ӆ<wF�_p����Y�(W�^\�l�Z܁���d	�թ1�� G
^'��l�]�aoơm��$�x������j?ye��iʡ;�)ٔ��K�n����~��U!��E�O<������Ꟙ�S�х�#v�!l�l�P���	��3�
>�0̃ᷳ�P�a\�Oo��^�6uO�(J��q�?/��t�~���.T�5���N�M�W�������khG����"�,r�hrba�jV�1d[!D��	�X��^ر����W���)!撒���$�Y��� L1nM�
�MJ$#�7�ߡ�ֱb��Gf<����C%l�c��y~`�̳X��|�-��w��dzJ�<�t�"��#@�Vjg���v��PE'���̴�ʟ2�ߛ8���ޡ��;���+?`��e@�ޚh�>tW,[�a1N�<+��Em�����/�c#3@��Ɲ����l���
�$8˘�so�!E��n�o�UATBԚ�� Ƴ�U9�L��w��=��i��!�^� p!���':?�w5{�艦���̫Y�}"���)c��ñke���vj��h���E5�z&#
����k�~?6BEދ���k����֪?Y"��#�ڤ)���ՠ
qTA���NѼ���_�@�]��; $psp9�u���Gv�w{��U���1n��C@c�q��.h�u���쥷��ʾؚ�xP t�:ulz-�*�<�w-��@�0�-US�I���?��(1k��N �ؕ�z�d�AǼ��%VZU���H��P�H�pځy�O�����\Hk�c��W ����o��p�]uCV{�|>PS!��4�P�<Rg��v�5�K��{lKAS�*΁7�����v &������zA�n�EfR6hn]���*��/]I 7�G����E�G�{��7���q�d�ϫ�ؕ+���"�������QL��1�A�F����VҰ�'A
��V�`6���Wr��F�_�^��K�zq\D��]�׌���Y�1�~���IU������۬e�#!���ufs	BK�8j�!�}^�0h����ΣH���0�/E�g�Ԁu�n�)��L�4`�����j{e�&�;([h� *��H��d,q3>�,A�lv����djڈ�����v��u3�{1#���c��f1���������)�n�d"A���˘�*���)���O�AZ��� ]������WN'U�B�i��X����;���C�]����j��Uo|�2�����mA�"͞�ϫ�u��3;�2{-jR�,#�7�J�m�eP�����z�N�����ح/4쑣���D���+h�;T���s�=&=XA�~0��A���<�d5�ͦ������Zv��:I�D@�����'=IRd_�G�G�}d��~�ص+��q�p��h�W���S�������Pf�z��GgK�VԈٝݒ]ʛ�;��`t��|�V�9�n��p�:��ܒW^5	(�%"|��IN�q{�l���1uqt&�g1a����c��A�?ئ��z$h�K��1'q߃�ر�ϒ�Z�A�7@��^�b�}3�/�d �~��g.��&h<���2���%Й�`!'a�V}�w'�	���ܑ�b�r��?�H�El�.i�����.s�ګkd�����������~l�������������\���7vo��븁�J�,Dl'MG꿑ڄ�^ϕޮ�>I�z��!ʍ�}��l�
����B*��,D�s��jB�čG�	Q�Pm270"3L����fl'��X2��!\7v��eI9ӥ��%TeF`�\���q���ZCAu����h���|�U����&�:,�ƋG�/���W�&��=Qy(S\Ş���9�0�X�
�NҸCp�u�h���E�=2��Ջ%�/� X%���7�u?V02�ADG�/��$�L�X�vD�0R� $a�.��w�7�X��I0*4Ӽ�-�����o�q�Ed�Ʈ��D�G�����N7E�#������j�ި�pZ�>�!_��wB+�b��R��J���Z0O(,U{&o	wq���+�MTq��
����3��3@k�Wui,����x��ua�;����k˃��/{��\;��*Y蚕���%$au�!���
J!h�q$9;�1�������c��K�PxsA���Io�}�	uog8Vo/N��*\
b�wf�=������>��ا o�o{CWູ1�Ӑ�9W�R��by����i{iW�o��~�O����׳%���G����io���)1�Un�!�����Ct��L����:J�*��h� �|
i�/6�X�)��3pQj=��6
J ��o$(�-��ze�M����!su�jR��iA����}3�*@��"�L�A4S����(r�v���+3��^���^�b�v��E���$�E!�3I�H 1�~܇�e������7M~���9,eўr�t2#�0'�	H��#��/�LG}a����8�<?F[�s�@���,a	�ĳ�A�k
z�"_�}\q�[5J�g��h�V�ۣo�^Q�'?#ײPiUǴ�d������l��8�8JǠ�sw�=�7tc-/j͟�0�u�L�F��K���1r��o�[�g�&M*8Fz4AT峗�m :�t��o�����+aGT���N���h�.��3�	��7��oφ�%��!��@ �@���E�񪔑�]�����@~���~=~9�i�.�칏��u`�%��H�&�����s�m�0��c��J��C;�`��S��ֵ��	�����uZ��Emo�q������"9W^�;rd����.��@��n��U=�nl �R��U���

3�pB��{�%R!���M ��3��X����y�Z��'w�+*����E�H���g (o��ۅ�և�7*'8�M���@�,ׅ�}_��}g�́��Uy2�Z�ɒ/㣛�&�E2����R�j�t���8�(d�� ��Oh� 9�Cl�����T�v���P��%�6tq�=�a*�:�M+z�b���}�.���O'C�R�cJp3���z*e��#�l�;b|E�����/��š)��,@qK���h���|&��6��w{{���(}��+��mTW��O�n�8�co�s���W^�G���:\�A���N��D�����HX`�֏v��
�jJ��r>��*%S����t0S�6��v����¹�������a��&�^vdҩ|�[w��4S0J ���e�>PG�w)�-���h�u��5�B^U�߉^��1���hF^�C���aI	N�Ne[�H��!���Oo6�x�`Cy.�B{�ڪ���`Z��~,p�9�쳢!�&�ZkJ&G6�Ax}d�wp,�{Y���3��z%��a}�	DS���@���8��q%�
rgu�"�"u8���!���S�X=��!��[�O,m��J��$3�Υ�u�B�b<;	��\j}�T{�YX *������b�i#ҥ�f�x����Ϩ*��Q�Xv
y�JBO��n���z:�֦�\�.�vђ�ك�����x>������^xX5����J��}l��;#@y6�GdB~;�{��Q�ೢ��h�f�&\�'$#/ǘ��y,��g[��A�-��0�!ќ<��v2���������ML�L�&� ���G�2$���W��q�jv�8�ԾP����bT��םtI$��\ՈtfZtu`7u8p�8~-�k������+�^�\������5�<뉔�g��|Y�%��̈p�d���'f���w���=@C�a>2r�n�9%@�}b3��a���s��[�lCU	wD)�����@��P�;��>�‵�HD���Z���aLl��6���j٬&
�������~z��f:�a���c'��s�t����T�~5o�o�Y��{M���ԟ�� .IB>c��
���l1B֝u��u�܉t�T^glFg��7������lpA2Gh�vA\g�����8�E�e�'��$�	}{;�H��F�0(���z������jO�Ii.J�X{�'HY�~yR��yY�3��f%�� -]?����� J��x�ږZ&�j�Ky�{�c	��� �Na��ܢ��n���~���qZ`Wt�T�����8��x�1b����)T�
A�X\�H*QC'��W;g>��!���0��M �>!��Q������S,����X���A��M2��4�}���u�$�!���8�OD(!��^�<\Z�m�	ww�L���vx��S2�iKD�]�~!PA�"6Z���(r�8�$���H�!��7�P_�B��JI��T��L�&r��Ӝ���y�z?܏�F���^�U5�N��Ĭ���1���OM�I��Iy#�L�X�h���Ҙ�B�]Z�3�|�.��Y���9�H0/�-��.�z	u{<Ε�;bXv��=@�oBD5�;>)y{�qeo����)+a��m��)o��:2Li D�U,��R�[��\�����U(��\����]K��OڳA!F	_��*
s'71�$w-T1�4�/\�`�>�!%��C���T?INS����P~{�p!�yP�2v�'h�8����l	� �&\��n֪�������U������S�ȍ@���@J��]�~��>� ��a�������%�*�e�^Ծfx� �=�cTS���ˇz�D�\�:�kI��)��e�!ɋ2�2#���N"��b�(/��Rs΢�Q�&)����-	�K��^q�~���Z�v�l��^Le�J4��1���$����W�)��4���*��s|m�L�3j�ۄ���k�!��})*���D>�Yk!"�8L�(�GD�+�&i��h�Q����{�S�{%�:p�Ɯ�묡zDL���r��NP��l"!|��I�=I�\)%Ry��`�R�p�El��|�tq�7:qJ�
Q�W7���&d�S�Q�-ZޞW����@��C��C�լ���[�����������~8������Œ���"�"�ov0�_�bHS��_����7U(4ciw���B�b��'���L@��[��&�Z����#?"���cC&z{�]�@�q�sJU������s�;�x��0]�7���Ւ��Q�e:|c�hE��w2�U%k�����eS�����ꌉ��wҽ">`?��k�{�w1<{�?�"<�"��RP��l�F��Y���a��LCgV^[u�h��U��,;$ه���er R��7(g�망��*�L2)����b"H�D�W�
*�� ��Sqz>J���I�&A��.q �������0��J� O� ��zUF�GtHJ�G5M��Z=�O�L�^�6ul�k�);���<����������&8FRwd#󩠕9�K�k!�+YM���ͭt�$WY�["�kQP��s@"[=d��ob�������o��ֱ�_�+�F����ub6%�����y8�a�P��s.��v{�<rY�=
�_:��;�4�U!�~F�|
ՏH��0x��eVa�[Jm���!ߡ�XBc� '�t����
;�8c<�ǈ�r�S�E��������q`
z�[�����mn'�PDO�Qs��i�����Y'#����<V�9 �m] �t����\��|���|�-��׍c�=D���L��y"� ,��.��hR��E@�����b[��Tj4��E�>F��4�|Xze���7S��Vf���>������.�����=�[���}��1�r�St�!F����\K��(�B�a5$���F�����g3����A|�G�UN���/���	$^�=�V����h��R�i�t�
vě�6`�6��>�oW�o��$�֛�P1O���5"MWF�+��&
G}U�?�-��v���=7]krm��k����{8��%WY4����\�)��Ǧ������]w&�.3M�y��/T�����|F㗚���	l��Q��;�_5y�G���<�z�aA�f�K�6�Z~Ѵ��¿a����[�o��w���&l���`7_� _���UW�Ԧ4E���&�k�h�j2�t����R���%ȴ�n�M�9�{y�z�yB�[��Ţy�U��[D60������F"����h��KբT�dcR��BP�H���)��OóB9���������(�K?��t��/�x�����~���Df\6��\dɎ�w.����&�B:d>�Fװ����З �	D]?��i���o��!u�_�V�s�Bv��ɠ\�Z�y�I�ȓ,l�]�����=���#��d����ڦ��{N#72�.�s��u�����,dX�E4��y�3Բ$���0��>݌ZE���%I��:,f��7D*J3$�[�WxU�-����F�U��R��F+�f�~w's�O�~,�m�/v�~�}ee�:	�B�U%��܇>,����/߫�y��4m� L}C�*B�y��6?e=�B��J^\K�/fZ6b�K�OL�*�[������\�r%���o���!�M:p��L�fɅ�[w΋��ׯ	i^��y��@�[^�Nޔ��c2�U*�c�vV�����6ߣ�2�ق�ݨ�������Y���,r�!����%�|�ww���1��G�����,�s��\(Ұ�E�|�����xb�:f���ʫ�ϫ��xq���>�~6O�r �� ��O���0pW�F����\@y��J��C�|m%���o�PF�7����2T�"��%N��/��bu����t�l��U�np[+	O�"��א��V'w�A j�w������:���I��u��rD�3�tZr]~�<�7z��*�]��P�͠e�=I��ћ�K�!g�v�8@�B��&S���ݒ�#-`w��^�6�q3>[�D��]��e���F� W����牬���wk|ߧ��AC�_��N�H�갑��4J74v�AP�0�,%�Y��#��8$^��z�jg]��e2rJl�e$N�/��t#�m�M �(�r|���?mÄ�)������<GL���Ǜ��!T��<L�����]	�̸�VJtة��ˮ�C�:4_]�R �4�Bj����H�J��Gy���A+sV��_��'��~Wg*[�Ǔz�r���C|M�!���G�C�%8&�E���_�gv�2�*νB�c��n�*;���Z:)���UC	�q�/�s�l1�+�Gc{&�r�kS\߽�����ȹ3��&#ޥ���'�-��n/m!v�g�s�X�5+��r��E����7O�^����'X-hJ덜�%���)M������e1����6]�ͦٺ`���L����n�dx��;2�R� ��'��g��y��on�@��+#8�F��v��*���M���W`uX�k��ƛ-� ���O�)�s��O�M�61��l?}��.
��z�JA1;��������6�*��������kO]*3in2�i�"��p��*�Rv�f����t�m�
CLF�խ��u!�ͣ�>�)��pLWBF�w�z���m٨`�(|F�ڰ~z�XG	���!T'�\��o�j����9�؈�ʟ��.�{�A�p�4�iL�w����e��0�&.}�7�-oW)���R5�>�uz_�'҂ �s�F>Nؑ�T2�r�уƣߪ�_�Uښ�硸�,h ���N��é3���y��#�/�PB���B;2B�`�]�}I���uF1������C/f�������=r�q��6��bтKn��F�������2<Z����8 ?`��<	Ar����W,U�CIa)�ߙ��F3�<��`�g>nBc8������~��y�&
c�'gLKD<+�c&���&u �R ����ԉ��7�R�y_&O�8�Mt��&�s;��59@#�2�]�"w���Q�FSV�ܒEW�D`�#��X|\n�s56]E�2����} ��7�Aя����gF@/�5q$1�h�.\p��|�`Zm��9�@�R�#ɽ��Q����pQ���}L[���,�?���zlrxB"���û�Klq�S�0����|C�6"Sxϡ�06Á��d�\�����[�q 	q�B�	���yZrjkG:Ä��͉� r�S~�6��{sN��ݍz�/7��Yg�O.�Ի��*�9���(� ��EMH�͓�\�񛠧��*�DA���.����
N��?��_�{�� t͖��:̩>�7.{���C���Cq$�;J,3����tw�m�+�1^�Q��7�p~LF�	�Mc�.	i3T�|Wi@���)�)�d(3�S�����Xi`�-�_&�m�$�'��/� `�)T�4:]k�ʦ�М�y*��kh\H��!e��/}����<b���@/*e%�=*.\�]N��.F-x�i3���Ή�q,��.DM�K�;X �G\`t6k�i���c�H��d�7�J���S��cig�Шݸ��%|�4���O.�k��IoJ�Q*�w�[0 S��L���
ve�
��	Ik��\rFhg���js'g�߿�I���YS��K\Ҁ�2����1���ͩw�X���mY�F�g�q�R.Ɣ�rW���إŊI��V�S��5�x�n�����b'�.l�(�xwpE;��r5����88�bB���Ot_��j��^ߊ?��3M�S�쌅Yc��ZG۶P˥3;���A�R�`Z����^�<��z�[2?��B�&��xҸ�3D��ţw�Ӣx{�\���oE�~���ч���w�au�<%htF�,
���-�v�G�6� �U��j�!����5={���X�.x(�ZS$~aNC)Nl�x�+���w�-c��Ҍc��X@l
/JD���$FL=�| ���Tqu�>�F�a4_�,��\�H�-P�D��${�d� 3J��[���#}�sP�_b��iE�ϗ���v�^�n��>�v�o�%ejZ>	&*mcܭ�x`������$�'�hw2h|�"A� ��S;9@��_�����vMT����ǵ0����4`~�\1E��e
�t=�Í���J��I#�?Գ;*�f<l����"����=�kg���6�'ͮ��)�-�0e}��u�M �g��Nhq�e~u�����oՈ��7�=��a̗b/��s�Qa���}�/::?��Z�~�3P�?ͱ�E�q��R��Gd�<fV���;��c���A��}3�����n�@2 �=���7�
M�7�3C��?#I�=��+�5�by9��L�s��*��M����j�h:~������i_����T��B�ji#}g N���^	d���/��ߧz}��4%a�5�O_�+ �[��Ҝ�.�~�1�u���H�u�L�@�ק�?�1���M@�c�jY_ ����X�n�y����&����/�~�����U�u�����R�t��q�n��=K���*cW�R&	9�z�{�ۆ�Ї��x5S,,a�#���~��������K��-�z���ii^��F�P[%O�Ah/�S)Tm�"�2�e�Z�՗Uֽ{~"��x<@�Ȉ�ee���T�R/��#a/ݧ����`��-k��V,�r���4�Qc�<0��t�Ż�\��N4E��n�꒡Lԇ��O�$g2i5���; A����c͐��yJ�c�@�߄%�!���e~���̜%Н�t����3��D�t��5�v_�z�x�/��j�d-��q���K�<Mȓ��ιn�5ڊ2��ƕ{��`��K�Ke��1XR���H?8��I_hd�ѮF���Sv�W��x�ٚ��^JS�`��a��'#Se<��G�~{Ǉ���P,�%oA�p�p42&�͍�
�'1>6��8&zJ��G,b���I��{4\��l���(	�6#bL/�׸�'>����,�\����4��/$��C�^IV�qDZQ�¤;���E!�>�+2/k�bY��"K�ѩ�m_�Ҙ��K��Wk�x�� /�N�_���9X3}����w���{��s&�GٯI�4�.h�H�+�5
� 7$<'q����94���F��+�$I�����=$m[��̝�*=��=��� ��9e�-/=��$����ܙ�jÓ��٪k�ʗ\�;|�m5���]�&�>t��4��h9�િǥ�e"�pJ�X���8��(>�Ԛ[j:!0+��9�v*h�R	�zZ���Q��?AD�d_��&�.�`�\.�nnŀ�^\�O�|K��N����0ʄ"{O/V��k�p/�PGm�v����E��ٹU���H��KS�zn*-qxL�k�`�x<�F��*�|K5�����hʃ�E�	�Xy�(�'�hBuՔ�n��Tf.p%��^$�F?q�w���627�Z[�?��&.Z�pC�s�.�A��ۭ�A�0��擮������������3t���9�CU+ꝮE/�p�!E�#S��� u���5vR������'a�m@ȤX�U5bDg$ez3T,䤫�����쌕+��&��>
)[t�5�Eٶ�$os��8;�*����&���ն�S�I�Pz�J�t�B����ظ�̢�1)}�
ʑ�G���Gz��r�
ĺ _e�I9R�����s�!	��0ˇmK.���ݒ�'�DRIfUe�O�7m��#��Z��c濴`���!Ya:�.29��]̾�΀^8�� �%���#�쯥�&�]-��5$RM%x=��9:���p�o� )&���o��8CI>�~�ރ��w��KzD�Q�b]�L<t����m$]*N�J��:?9?e�۟�s��N�5�GZ�S�2�qapd���Ã�'�ZƴI ىHp/�NS�zQ�T�!ݚ�aF��0�|��6eMlAژ�;x��ST�A�Ɉ�֯�,�\��4Ƙ/��r�E��Ыnܽܺz~?�%� Ҡ,��_�U�Ho�1�ܲ��V�3a Q��]��I�4���#A{�ɽ�K�l)���N��ת��*Z;k�g�G�&�['g̥�w7Tg���u!����rk�f!C��'��7�iy��{XI��"�]�$\y�U���s��R���k��g-����>e���'�2�y�9-]��sn����\�S��e��u�w�e�x�Q�-���V��IK��?(n~�#F�f�'�k2pą?�J\��F&(�x�n}��8�:�gP�w����*�ʓ��J�(�c�+1*�]{n~��He^3e�����'P�nȘ����-� ^���jɤ�q�K��m�<f���o1�Ѯ�B�:1��D�U���Vm%M[��2�euj{bbQ�V��m~C=�SI�1pQ��� t���7�{g���J�����K�4� ?|J�?��%�U�����$D����&Ib(��{�>>T����Wd3�S�OKv	f0�ua![ߕ��6�L�-�9�0HĆt���2!�#��T�,����(�Vz=C�[�6sL��R�dZ��f	U��g���Қ6��^@��>��V�$Z�ч�J�_]�x`X��O.ѳ�g[����@y��g|��p)Z?�KBa�p�j\���[*n ��M����<0���_Ħ�뀅�q����X�q4��g9�*���9��x���pU���f*f"%��BD��i��,aZS§1�+IY�Q��$��1�@	����zI��&����p	2(dsm���������G@dƒLl��O� ?�gnz�:m3&۟9��6<�U��d)\��tdR���}���jƇ��8sm�z8�tv����G~�VRN0�2��Su��i"�+K�a����¾g�+T+���iP�D�˚}Ȑ ,�)>�R.�p���.b�Ǟ�G�f����Ֆ�p�r��b�\�V3�q�m�A>ŎbK�t��[5���؁ְb�0ˑr���vd� ;>��0Ӫ��o\�$��[�IN'�E9k���P�lW����C��M'��nʔ�^�J�z[�����u��S��C��>���^}W���?�xv_�C���2+g�_.�i��-��]$��Ø�{@Ȳ&�����F|��:o�A{�ܵ1����!6�%��B8+���ꋅ7�2l{�p�ômbU��GҌ�Gr����Q��Ջ���d'��L�^��]8��J#��Ia8T���2 �R�#[*�u� ��n�R.�e�� ���'��5����`d���D�� ���s��8��Z$�S�5%�fv����ָ��������6����,9�3Ƕ�\��CU����N��T��	��Wn�ޯ x�ցB2!)��IC��P��F���YP���BTLZ�p�d��C��[�3/0��	 �Z��&ɻn��zu�~���8 h��C��K��<�����ux��Kpؼ�k?|p��J���
/�#�x�2��Mm��E�ކ	T��5�*�+�WfB��we��4���Y�ӝ��p�*���U�r:�>��\�4"f��n��9x�)��_���[����{kSfFCN��y1-��2��mu��0Y���n�IM9.���Ӭa�n���rҺ�Kb~\�ğ��[5����"0��NƉLC)�kҊٲ��2�s�#b�OL�c>k��}��{��t��.M��%�<?A��~2I�[�g���%r��}�d�,�w��Ep���Ԓ޺�Ԃ��	6�Y�?�V{AY{�����uvp��In#p���������tg� ���>��SLG0������������=ts�'G��pȝ������@?�dY�A�%n҉��\k�L�Gv��T��ş�0�ȟ�<�]JV�F�%�(��Y�?tc<����mv-��)�0j�מʵY&�w��;G���'�ĊxTT�H��Uє�Z�>9ng�rR�6se�H�`��*�������Z{� ��4A��(�t�!�����2x�fV`rz���zf�34R�n�@��w�Md�E��5�v�i����wD���lHl�ou�j2*U�z��mMA�Z���Dx������IXΛ�g3����&9�ڡf�^g?��dI��m�����^p3c�����ȶIN{׆�"*����C]HV��=�5�x��νl��7�Ѫd���ď鈾�aԁ)�l�n�q �_��F�fs�s�>jY��I�Ͼ�V2�|�bQ]=��:�>1���-|��zZz�e���Ue��J�۵_4�������.�� н�b7���͡�-�p�K$o<,y�M�@c��h�_4Y�{h�6x�W+�x4����v�D99^U��хm3l��ֲ�	RBu��K��ҟ�\�3��ԗ�FQ"�f����h|�0�M+��P�ok�	�����d�A�~�Et�*[�ڿ�D#��g�^��f$v�T��:Q����7�{=�hyX>T\�����5v��pV48``Lt|)���r�F� ƃ�o���8u�UǆѕB�0�/7�x0�7v4b�[��������J�Z�9P_ș1P1տ�ԛ�Y����t�#��2.���֔uW����K*m�'ވ�(�g�.�g�Id``λ�4zd������g<8�@<�I2�jN���n.͔�EK��_\��V�� �.���&��L��qld�Y�g��I��3nh���q���S��f�+�-o�݌�D`�cQ[��\��	�\۵Z��$u?�J�p��l�N`IY+�o-ty·��[�Yƌ���L�O>F�Y_5�}�^w�z�_y�� br-��4�s��.���k\�I�N�"��&���4P����Ѯ��:�w�����&�dD�'�9��g&~(����7�x��E�k��@+űs׎Z�F&�NZn�W�ÔͻҌ��@E�x"�=�$��P�v>)t�d9�6�{f���P�BPM��~����trW�XQc4w�^�mi���FM��.t��ՁF���T�&����:��D�Î7鬓���ƠS	������ږ���r��s�Lʂ��%I�)=�7�vD�W�^Nt�����s�.w��&�������	����X�Qn[�ųUz:]�����$+<i.�a6gM�ef���*�;E�M|kÒ����J!ޥ����xu�g��dQ�l�t"�{� �]2h"b^>C�a��a�������ʤ÷Z6����>L�����ӳ��Wb�mFS��Nɡ�6�Q�zB0Јc��TD��2!W�覽,jI���Ƨ�X�*�%��(s��s��:��^����@�I�_ Rb�2S��nr�jh�,��:�H$1�����54��q�c�ݏ����a�XF����d6n���8�O1���9p��}eJ^�<Ċ"�-�K�t�5;�"�)Cqn[��Ĉ��c^�n[o�5��tܨ��?6w�~
�ͪ�e0UQfrژp%u,[
	�CYYhc=�D��+΀����,\��2���qeb�\��7���rHW@C� '�3�j�Ῥy�<��/�o湖sY��/��̩�v�<�e�E��)̺3�\6�<�a�d����3�Vp�3Z�kU�����0�z^1�LlI�gk�0��"��ZQ�2��^�����Kc�P�՛�䵚����!�{A��"�����L��m@����1៸�H����u�>�uzKӍ*���"���H}�u�0��C:ŮD�Z�U�^��æ�$��䫜����%��=3�C�10�����D���y���*V�H&�)�� -��*K<���3�]MԾ���Q�ٝE�QE�>����lpR���7��5*IT����l�^v����������������RmHUsh厦	��G�j�s4�²�D�s
^H����ь�7���5EǊu�(�X��ќ��|��spv~����3�4� ��t�h����T���K�iu�%��%�{�kwI%�9w�C,>����F��*�~� �1�$�]|{F]�Ǻ_�ڙ�����GG?�q�,��R��G�評%+���U�Db������w�ނ���6��d%v���JΞ�)�\~��~��ֲ��l�0�� �xa���N��u��0G��Ç��9q$�����ۋ��9��/=s(����,¹��H��10E@@('_�J 'zd�VͥL�yd'��ʰC�o�P5;�2�+��]�aX�mĵ`;p:y��|��QE�嗰o8L���t������GA�a{I�A� � Fi�Em̒�e���Ѧ�o\����_cQ�U��J��Vk��@ߣy�ؿ����<}8�a���}�^��L�n���I�����|�n~'��U}ɧ�U�q�W+5�H��M�ߨ$\�r���Tzv9�@��)�����I�Ÿ��h�uϣ"���W0��Y���4�8Vj�+���L�7]y͖���FV���`a���y���j�/�5��9K��)�_�qz�p���u7�u��{�记U��IG�a��F윹.f�8�Yhy�W~M|����2��~IZXT �����T�kU��6b�}�}��r���K1��y �t�Qԅ����&�"��s��CZ��J����|�Ȯֻ��%lɈ�
����|.Pٻ#�@�ćt�q�>�k����1u����[���'ҴL��K����'
��{�(�ut,`�F�[��)��nd���j"Y�ϐK廝�6-?�OT���$dV��a��=:��Y��t�Lx�`����2��M�/��er�Xo���}z�j�`Q�B�i��� Ty*������^G�R�S��H�9�����ce-\'��|`���i1�t�t�C����A���Ɩ�盌{��L��|�(:aR���z���u44�(�Ȩ��R@t�Yy��'Z;�;A�ta^���O�̕As�'��J��^���M��-@��v$�
��%Ps�a�Gš�@��7�&ѭϡ��QOg!:Q{ų)��DƄ+�˿������(�����z�8����-	ΏgAϦFK\A�Yŝ���hg�3"�s]-Mi���	.��:o���/�g�^����ot���vrW��_F�-��`l�0d���R��\F�K?%0��\��^��oT-�x�Ƚ�sS��i�ж��U���T(�&���r���J�&�]c��Ԕr��F�A�uc/%�!�����#b�H		T<��[NZ�9�M�)Xˊ.x���<ݝ;���,�o� ���vpr��$�g^�-�z�c-��\�T6I��7ٛK��LO��:0_F�hp�#B�u�^9g��sJ��-s��z��5��E�x<�4gp0����4����AAK���Y���FO�X���I�q�G����U��3�A����Gu��,Ք!8�?��o�p�ɶE�I�9q>5D��:ا �Z�^^g�y�(����F1?��:��E�?���3�P�G����5�-c�ot�qb��?hn��Ȓ�e0ב6T�>3-��=�;���1���4�fn���XX��}� �td)�<� 9�B1�oL-)[�6�?<�B#i���F�=4�'h�̈́��Ej��o��Ch{3�/q�Ϟ��������G�YEdo&���}�PSo���\�[���#G���1""Ɂ��C�r;�bo�F{�o�_�J��a�·�kOɎ�-�*���l�����&��t�o����Ϙ�E C�7�:{�Xk ^�s%�HKǭ�*1y���.��O���Z�>vC���t^�bN�|A����i� �����`~�f!?N��RѰ�vLEB?���m���+���8"�m&@-��R0�uh錎�t�߳��AX�(�*�D����g�¦�td׈�F���i��?C�"�RÈ��{P�;��ա�:4gW�*�q�HQ�ڌ_�B��)�M|l��`f�1����G���V+I��� �����R��Y8��DZ�L�]�i��Ŵ������OA^,�d)��p��@�w��gn0>+Bns�I�W���t���j5�'ßӓ��ʧ�ryn}��S}�#C ���b��d�>���E1�6�j����WU/E@>�� ����Ժ���W GM��&�X�\��|�,���a�V4l�F������rlX
F����I��CҼ��.YOѓ��3��s�25>ؿ=3�T�e#�U��iV�{��4��Y�f��I\ٖ���V�+~0'UC=�N�,��A���CE	B��	��6,{�A��#�ԝT�o���Vs�B�=*$�Ӵ���f�Ie�Pd��L��gmr`�=�4��}/�S�R�	�
hI5@�eV�halL6c�����FQ�Uv�u�g����i|�,g4�\H�.��5���-�F�b����
���A�:B�[+ѫ;�!���n�y���z2&ɋo�Od�>T̮��5��	>�iF�`�O�?�s��"z|�Rŋ�'=�������Z��J�a��.������ �¾�+mM����"z=���D1�$��Y��5�{9p�Gw������&Q/Rʬ��l~�hi�?�E���4�_,���eɸz��#~�^|�����j��xe�;KmB�#�"u�Cw�vh�Ә��Pi�|�,�O�Qj��f$q@y�D��3���*nn��%"͊h��z^��Y(��fb.��ӫc_q�}qOVF?T4�H�QjN��<R��r	޶���6>J������jb��D��K֞n|D�_��2������ۭ\���c����3���I^.8�E�XN�نL���[��]�����4G�"��EpČF��b"��ǔ���.I�߃�[�/�T����˲,����t��&�]7�d�x
���e��˛Q54�|].�ś�ö����M���{�0��ġ�͑pn���4[���NV28gf��?��E'���J����H�Vvo���mu���vF����Q�`5@��\\���AY�q
�',�Đ/+a��{�V�VZ�Z0p��.��܆��^W����i���/���%�`D���}�岢n�������˛`�O���&hT�/ ��z<$�=�S�����`���8��I�A�Te�_�xGl;�
H�g
��i���.�`��7dr������^Q��p��K5ZZ��~#Rk��Ӄ*��ވ�Ğ�՝�ʎ�,�0��?�#�1��Z̓%EY��Yk,oy0,�WYWw\�D����-�ȍ�,A��J��#��9G��i�AC�RWje{���QFࣱ�Vr�X?�o��ĵ
'K�`�a�������6��z����*
��Í�,��c�X�W'}�/8���E:�=<O���_u�r��r2M�KX��1d�Ol/�Ό���;4]��/*xU����d_g�Sr�׳���qx P��HpZ�'�JkY� T���H�eZ����d�a��;�Lu#	�����>>G�,}>^�TQsP��:���rN깝�\�$4�UZ��� Pc唝QU����Q�є��=-�*��bsT�#�l�M�Jr\���t����ɔ]:I���eh���&'�Ϧ ۦ,��V�k��Q��z(�/4Q����T���˲5r:���~��&T��E�Tn���%�ʐw��Er(�7�57�ݿ�� G�Q�����H}J��F��PoA�sA�o�h��Y2��Im������4 `@�o9xE��!��IWG#�b�m�]Mb�/ڢ�8��O]L��,ziJ��2��B
z[���aϰ�~��3�)�-п ���6U�������� �>��K�S�.��^"
��<��g]�&΅4GF� c�?lY�1���@h ��оo�����A��PI�,^�6%e�H�n���A�%גlI_���g���sH�qcG*Q����"D���$*R]���Ӟ����_ׯ!yR7�TԜ���t����-(#��D�E��]��\\�j`���^9�X���i_O_��&��^��l?�"X�Ehp�#B�;�So���4<���+�	�S�(���i�M�eT�x�& �+���U^����`�Z�*�Ң�F������YuL����A����=2OZV�lQ
�]����2K���\�jN��]c #�y�U�,
�o��$�H��WG���`�<\z�
)d@�T��r�Y���)��H������O{�����i�n�7_����o ���/���%{!t�lVw�''ly�)���	؇�܊�k����	�)�w�r�@��J������͹Ǽۻ�:�B��N}�L�B0#������=�D��n��ڳi�q�(�\{1-8�(1�Y��o�����˷��р C�v�_	�(E����) h����NPp��%����&��w�R�F-��:�)�Y�<0�·����r2f@`?�w;i;��O�^��)0m��4���q����0�i�S'V��X3\D��$1c\k�� ���V�������MQ"��> [��s�b�$�py����#=�L*8s�`j?��4,�!��d���^�?�F�E̵+���
��,�R�iSt��]��wq{�r2z�5����v�J��	��u�
�Q������j��Ց� �v���9�B���眩ن��ě�} D��y��N��S�!��oG&�.F�D����-13�0b`o��[5�����;��W
���t�g���+��پ_1�yz�uޥ��/�s|!uN}@W�Z���_R"�\��W
#������4�eR�\]�*_[�n��y+^DoT�l��@X��B3��N������u[@bj��%O}5����<�$�����F绥�~̷�ie�éy��#Py\�u_H�L�;
��� 9��2YV��3Y���O��MJ���u�7���8������U`��h����q(�,nJ�BX_K�q(�ȐQT�fH{�(��+�h\xt۔rU��Z�zݓ�7sK�BLǯD���9jP:[����'B�h�>A���B�S�ݮ�Yb�5�|��D��\,�������*@���(�jY����۩xؽ���c�QK�B�ࣜBN����v�(�y���ȣ n�S�ZXU�9��B�i�fXtݗfo��@�����i���Ё*�- ��j�%�˲Y7i���+��/�k�'�σa|�&)5@�������a�R�i���9N,{������u\!2�XMT{��(y��WÄaص+բT�$�3FO���>}�Ǌ���ڶO�(�zfse|k��9[�^�%�+@��C��c�(���w��׃�[�k����m��)�/��0�������@�p	r�ðt�"?��2�jtO1��Y��u�LdD:��2�r�2~ l_�Za�����X��X,�X���d*����8�o�����S��#%���� ���7ux>��<vp���aP���+�r���;A$��A�7�=Mf����|�7FQṘ;�>:_��Q4*S�q���r�1-��r�q�<���I��|%��;�$=��K�������sm�ک7�Uxb���Y�y���@����>M+7i�p�m���O[OjZիD����iL�~�>GUdp\��x�Z�	��%\�$���2x��͡r$O��.KԥMWG�!q�IWI��dĒ9cKu'�����R�:&6sQ����U�&3�AGǛ/�7�
�ǽg�q�w�lu
������W�� �-����
F��ΕŪ��b���w��
��O�-����♶P��V���2"s�����7m0��Rr�.rKZc������v?�� }�E��#����S�vCv�^�˩X�J�/v��1Ͼ��TR��֚��r#�ҡ�OD;4��0�]�9�<�P�E��CNm�Z�Nn��S���k��2�[�P�8�}?��*	�lz�AG��u�֧�f�:ƈ�t
B�H�{���Ck@J��ϗ)��_�j>ZN~�F��,5�'�s1UF�%@������Ʒ:p q�u������ggŖ��>"�RL�A��<MY=A�`ջB]�jg{ޢ�Myy:�P3�T�6H��G�� �qQ���DG�N�����ː���[,&����93`��+�c������9NILf��?��Z���{� z���K*qʴ�Şǚ�,��|�Z\�@ ��k��K'NO��GJ���qk�2s+	qgQ�1W\�A!J  y�r)r`�d�w`y�r��C x=�/BC��hs���b?_}���E)�E�����h�G���{ ��N?.	Fv���Ę	��q�./�0Yjc3�#��]B�G
�Ep�%�13���؂�~�8W�{X��&e^���Y�3��[N�2U���brC��o��F�$�Q�"����Q�E�J���פ˥��Ӻ��j�k:���{�0���x�*�8s_z�W�2�B����ZsJ%�X��<?�d���߼?�;�#�����3�!��i/��0"b �Uf�5N�ו��PS$�z��t{��K���*E8ӱ�'pbF�+b�XNj8nR:���Y&���v�������ѣ�?�;i9\H�Q��З��<������*�G]s�!J�� ���N��� ʇ�a3�Ol��f��/��>.+����L�qNUڮ��k��t�
�,������Fc�g��24���%��D���"���~`������|�v���f{.}
�J�$\��g};�K+_r1!�?d�����i^+==3h��vd,t���F�Mуøx�ё�2&~��vK�=�-(r[�!�,�asY��)@�y>-`46���/��y'�^Y"�	�\Q�c<�8���_�Y/�q��ݮ7~ʮ��2��F1�A�jxhs0�Y�����?�6qf��
eڥ��58��G;�̍���`�KC�
�W�n	1���{���&n��6�*��);ȠxH�KW7"��`9�tP9�nB)"��X�x?����<i�	�e3���Q�,�<:.�_�*�;<�x�؊��愾�P.:5=�;�eF�`�O�} �ee�n���TLY{:C�<Ձ�i��<�kDľ�đPP��	�}2��b�Q�aD�o%�J��kϯC��FnT�Sd��] ��Y��8�M��|��\eϾ���#�� �b뮓�9M���:CO�hM�]�:�G�)��E��d����kXV��\��}������ �Ug��Q:�a�}?�$&t���mkl�6��=~�/����b��CH�
#N Y&*��Lo�t�Z]����_ e������:���O�@��)�v�����i�\=�����w��ó�@�t�*L���2�=�]9K�߂ㆤ�w�!w	��Ȼq��e6�쾮�2����K��Yz��fP��j����#xnKK�G5�����}��D��Y4ր��aP�*Æ����`d�?�n��P��F�2���DV��Xd��t?QnUv��S�����˙��/�0����6\_�S�yD���?���Ŧ떵W� �i����0�
.��S�[�8��.yLl��t���<� q��4`����7`k?���Ρ*�,�	���
lbt��	$����*�>��ؼ�͹^�8���5����-j�2ej�����Z�R��0p�1N�[Fۗ�r@'~���lh�y3���L�/���w��c���<��-| b��6$�� H��{���'�=�j!�f�?�ލ ʀ�?x��t|a#��͎����e�\�`�y?�5�n3Yo����&gN��$�£�;it�z�M�/4��xmwt�j�%�׌t#���y�H��rr+��V:�lT�r�7�����*5&���a�|I���
(�^U�F�(^q���
m%X����Nn�gR���B]F!�@����@����a@�H�_��Ƣ|��=9t��w��	�z�)J�j�@.H��^���$rtV��W@N�������{�����8�}Y��71e�(O�ٟ0i�*�m��>%#����Eΰ��d�t��Q5�<[wؓ��51�$���F=V�Ҝ�ľ���>�}%$C��eT�%���IY���=����5��w8��F��=&">��/��?��YT��^,��#���	5
����HA��2���������7�J;��F������ϲ�3�^+@V��{�`w�J�g>��+���Y�(��M�d�SL��3N�m�Ѯ�e�9��Ze
���������6*&�v*4si�WmE��_?��Y�08��tn���-�A��a�O���Pڞ5c��b��@К���}V"��Ƈ3fz�9���z��`r�vl�?�x(މf�󎚍S-��YV	ۆ���]9Tt�j�Ψ����Y7t��h]�J/��lBd���]��L�)�R�e�c}ha3�Ym�q%��Q!���-��z{���q|��<|>�*�2%y8�Wܿ�ޏ
��$M�a�ɳVh��?U�̓�'r���D��mC&�����z{��rJ����ь��Ն�� �4�o��z��	4��$�b�^R�`Q��9��|��-a�Z7�3��;-1��qt�8��څ��Kd�0�*�`�Ը]�w�K(����."X?A'/a����s���2�ϩ~�K�Ď�g���T�S�Q����ѝ5�W\�t�o�.��Y������|�nYX����S��nT�*��qf�8u��n�y�9�����DEu~�}�_�����}���j-`�`����]m��d
R|�A?` %�y����NcZ�O\x������^�~k��]}�ɋ��)�gT8����gl�WP�s�q(.���	�`�p�9,OШ[��d�R~�� �n8��.�h��N����C��_���>�r-`�s=q�0��������-#iI���H�ns!M�������E#���q���U�ߟ��}���?7�y�.�i�^Ç�H�"�q�m�	��*$)�hI���^�3����T?$�R�YL%<���-`y�D������
ۄ���)���W"*M3����73�2 %l�.d�O��y����T�{�����5̀�)���V�[��￩ǿ[ԧ��&BB�������P��&��Ol�uF�TR����R��5�#c��M��֩x�B��'�,�t�X�6�^�Ki�c:h���i�ܫ����:�҆O)�8X|��PO��[���;j�(���`=~u+���
���Q��1C��Q� �p P�C�J��׷�q �l�]�����	C�l;���%���,~�4�3`"�Bq2c���?XZ��Tm`>	��e< �h���8�LyT'�F25�����3U���{�r�L�_�����͗V��9�+!�������웻�)�)3WX�Z�ф���}�q����'�"q|��L�[�y@!��	�ꠀj��S����EA�X ;_4���d8�&+��w���<a��E�hC'��@:z.��`}�Y����*#�����mT=�fr�\U3��1oJ��$L��iM�p�LZ�~����Mf5�3ո\M�i�	�����]5��"�*��c����??%���%�5	!v�:���,�KX�3�G�;o�;Ϣ�Qsh4x;E���)7s�^IG$5�Q���rp��:�P���5�����T���C�a�f��G�k$�D٣3��������f������ݏƔ�o�:���B�ۅ�n�z=A���Æ��S.�9�sLf�\P߻#>��^��(��\��U'�7�)/KK��#{���3�`���x�oN;�lci͂� �G��a��x�0=���Bn����@K�$_8(52W�$�fo�;H��1h���Ӎ�pۥ�S�?���cʇP7��$ɩ-�i���f���X(������NB�1���^z�R �r�f�K��,���wiAdu����,`L">���:q6��W&�G@,�.pϕv���`�)�T��3��P��o������q��FpU�|!s(%���!��4�F���)/�������S^v1�f�f�]	n�B����Go\�^��ΗY�>u�|��#���k���1�Dy���,
[�"R%�����ӧch����(�(����zv�<j�6_B�Q~:���/���{����Q��![BU@��W���ϙjضe���cbx�f6�4N	+I9B2���:��/K���#�hʐ|*�b#{#tF#*�D��"��p�ϸ$��Ԡ���u����*Mo�2j�
�}n�#8��o���@Z��z2�:���:���,5}᷆�e�����G��֧����u��:4���`;�qJ!����؆� (t�:@^u� 쇳EQC�܍�}���o��˹��⣱�J9Y�C<�|0��$�C@��*���D�G�+�*=%�	*�m����دx�r8&)�F��"$�O"��h�scȐ��o/���u�[7��g��AZ�mu�[�0r���@�[+Eey�kdff+h !҇�]V1�z�ɡE����
Ɉ�bF�>Y�e%;�{�eN���=l6"���i�:�Y]��Q�J�!?�.2�v �ܴ��$ȷA�� ����j�^?�lV�9hk����%ӫcm��$K�X	*q���7L�y\xu#M�B +E68`礸Մ����(����Z��d^i�̸
�$[����4$��������tyC�L��'6�O߁���>_�2	jӫ�a��\� ���V��i/��eJ��?-)z��kM֏���,����ԡyv\�Oֳ�����=���-s�a�E��,�i��`�+��S�h���g��GφlI6u?V%s̊Ό`E���a�(�{V�����h�=�>J�OQ�lH?a�5��#"/�sY��{�:=P?�C��2�J�`�$�F��;^c����A���b�P�}���q�#�h��H���Y����^5Ѹ�Ydr�%?� 1�Z����T,!|�I��y����Z]nC˗���K�vQ@9z�3tը�@7�3Pŷ�b���i"A��7�u���oFn|��	m���+F'�O�L�L|���� �=l����7匟�jO�h��oɚ6Z��N�M��{���!�j���He���+F�@­�Z?��F�x�lI�26OS!ٳu�E��<��Vq����z�x�Ak��L!��/�)�U�>4�A������
hu��FX��j�U����1M^bX�ҤI�=:����r��Z����Y=!ꇤg�x�Ƀ$��q�n�!��`P�ꂥ-�'XM���~v>��e!�4M�-���Y��J�}!7�c-���e 8��[>�͇���m����d/��X~�P��r�C>��S>��ʆ&�D����!h(��h�~&)��1Fp���U�"q*dS��B��t��[�4;�G�>h��y�;m����@Pc�����G�)=#�'q���я��ԓ�f��!r?�=��Vy��)����A�d)�6��3����^��>�rU`!Y�i2(�����$�&f�W�J�h'6]*���1���',b���w��/`���]	�h�M�ű�9��f�L3�¬���������3�����h"��T�" �H}�>�����~�)pq\M���́L�@`DOv"}�6C\b�����D�(�Y�5��Z��`�@?q4�rc��N(���mq�5Yi񣻖�6Z�)�hܴz�N2�7�HE�~[��\z��:�4��p1�S3�B��7���������{vs	�bZ������zT^=7g!�6�51ۡ6�:�H�8�o���7�Z�����?����D�ߛ�KX��ӹ(L��;jfxc�G�3�6���o��+�( �i�S��t}"I]�&��Ci'�MT��Y��1�>��+�ږ��x|��/~J+C)6�x3�f��D o��+�SW���
-�+ͣ�|�b�)&_?8���rC�2W<�T1�(��%N�d�mF��&���S�[nS���'W|�Җ$Rవ��E���Wh3+wx�R;�uxTEq#�VS�ꪾ�xq[3Z2�>LHk."�	
��V��A��Zb�Xp��&�_���r��ge`�O�@-q�@�y���vU� ���ˢ���>���y�J� ��F�� ��T��yĔ����7�v��<�}���׎�!�D��迖?���t-Y
�G;EM9ys-�W��m�Ot0���%��ѝt/d����P���ػ2�F�Fh>*ĥ���u���<F��5���K���4��Nb�x�����A��5�%P6��!=:n{�!T�Kġ�k'8�T�#�t{�o)����즗a�����=��e&��p�1ָ�O�q�i�P��K�vZ*[�W\��Pd�|*��$��Cba�U#�[.���X	nx�4�`��GH�WbT��%
��jS_|4=r��EtK�mfN�(tsg����p��.��\�Hx^Vq^ ,y9�qc�F�.J}��Eq��pS	ջH:���r�b�BC8�oa<HgZX��/�.ƍx�f!�b}���X�=��g��5�n�=h@�����z�)�ǿ\���,��
��Յ��f�.�t�L�i��NNL�i�G�,�\��6L�O9���֣����D�l��=�h��>@3|8���W�^#M$F!謖��b[���:
����'{]�c��/x�]sv9r��Z��9��M�'�I�U�65�D9[�wEtX�����
*=��h�J\�]o����w�]��
-�a�tqǧO%ؠ�bJ�0m�[W�")t��c���9W��A��jș�;��U�-#�~�ٚ�J�|;�MȎ~����:fa<û䅠y�8�Q=�����x�;mz�*�4zW(�8��\�;&�Ƽ|�\�e*ݣٽ%7�g��g�o���ҋ�e����m�t����H��#����9	�%�:g�f��*���{�T����q�cG���x��7��5U��a�?Bc���Pu�)�~KP�g1u�)7�+"Eso-�tݚ	Oֶ��>2��E-�u&˼�E���T��UX���7Y>Fѹ�'���6���y�.0A��2���M�"��}��sg&�N0˻9�����H�	��A�\�U����+���xZv�/��ĝ�1�}�us!�o;X�����P��!@��#SQ &#+9<C����,J 2����q��:��=�m�#��<ә�[�rO���������~j�2#y6��{@���`U��b�)RA��Q�.Lu�1at!.� �Ь�Qx�Z��2��;|Xw��f���ne%n&�Ѽ�����=dz�1%��W�8� ��DQ��
g៺Bn�8����+@��Ć%��t�'.���L��6�y
�%�֥ێ9mL������L���*H�r^�(wq�d�-D�x\<��B��u�Y�ns�����wѤ.{~��� ´��Y�~L�z�sڋ2�����7��3����se��c�|�OI]B���܅��̞ĨY�̹vJ<��4�?��k�s�wV������J�d�p�$x�	U��l2�1.[\���������1`�+	���k���v`��s>�׮U�rЅG��~��^�y{ﴈ�H��T-
�Eq����'=��4=�?����ʼ�+�ٓ�@ԯN�rY4���k='|�������^g��T�(:IH��xMӜx�\<X�J��@�0a��Mz��k����1"3�(Gwy������� &;KT�6��]�'�3�v�Q �wP�,��!㪻�@ٟu+<c�W���<Q�|���J1L�Lk�F9 ���_0��x��i0Ye�Ά�Z�j�h��Jď�g���-�x`cIo�J"])�#R��b)���ċr(���#r�._ϖ'�Ic,�Q�`����$��<����2�YE�p���k��y���3��8���͆8�ú������o�#��>~q���m�d�ͩww���<Tr�G��OS�~w�%���*��t`.�2�?�6pH�#�|�5��|"�!�J��Ne����t1C��=$g�m֊��=8�5O80@׃0`[b��^�5�����H9pљ�sy�bc���<O�Gk���Y����^24x2��a��5�6Ѿ��~�'���(�<��2���A�ܚ�'�ז����?�2��JpK�⎚=]H��0�XIο�6x�Bx+�AV�K�.�Y���Y-��7A����k�a�aV]�u�7��]~/����䭫j�Q¿O�	FA*�Y9����G��?m�gV!2u%Ą�_k.�q����<��s١�P��g)� nP��wY�����AE�Y��on�F{��4*������y/
'W�f�_��ǋ��=��cğ ߦA(��µ.8�T�̳��'B^�����
��o7���$�⦒�Y���s���Q�`�E	��M�VzeQ��~U�++9���Q������G!RpW�4�����i�V�i��gW��0�NP��(^�r��I�:�]J����o��D������.e me��l�/��-{?��GmF����,�E\�)UuW��Gz��B'F��%�^|��Vg����ѾHwU'�]%@�.%o�uDT��0UEc��&$� ��Ym�7d�>��*��Ǻtg��"Έ�qvHY?}.f|E��l��DA�i���M���x��|��uZ6���:)N�p����,�C�әb����}�������t3���}�������<���׍wH�5�/�)�x	��Ȁ~n�X��[���-ЦO�=^l�Z�x�5d����� ��*�|Zo)z$�̾Dk�9,yZ��d0�gB?Ʊ>�����m9�M?�'��V'>���m���rp��� (�jຸ	�U9���Q��ѱe�r:���:T�7*�N�2E/fy�U����̜�#)�B��n�s�M� �a�����(7�!v�q��k�-��K$L�MEl�1;�*���.Ɓ�S�,\�/����
IÔx���J��F��NQ���{���X�/Ry���	�Ǳ��y��O^�/�g
�t��X�]
�zD3�ֱ[���X��g E�ŜT�
�&��Oȩї-+bI����)��L��'�-��^S�d9-���w���AF�L�kn�I�A��ʣ	ĤZ��� �0�Ǜ@�d�"��:)~������h`0d���I��_T8W��]ҏ�������=C�ds���
���������/�M����:,3�t���&N�b_+Q_3B�Y4���S*�S�p:|j0ù5���٬v�@3R�-�O ;8(�L(�r������-�i��p�����}� 6J{
i�LB:�eI��X��h>3c���<����(6P� ���hK��ѩ3�^�>op�ȴ �����8:Y?� �KO堕&�p���k�tO���4���1m%�w䙷>	���?`�z�>Z{��&�c���	���+)l+R%a��BP��Ztu���a�7����h��J*$>��X���p�dIΰ�2�K�{T+�#�b4�:�����ZU�m�V�{6=|}�緌�*���ӗ���r��a�c{�\
��dJ�{3��K�~�U3K��������j��lȂG�ј���U��ؕ%P
�k�$f������ޤ�)�C����=��h�԰UǪ�W��x�$щJf�bT4����E�|J�5V �Q9+=�ٶ澷m�ə���5�+�"�h�ƲR�����/���Z��5pM8��l��? �P>�3h1>������`�wR�lBL)��`���T/й��Ş�x����v=&�,'���Q�'���@:t��lݮO�y�	|�,h�qqf�`'`9���s�y�=����/�p"I��"H>������M���]���&�d�2���O���A��Wek�iKJb?�1�OHWy��Ls �1��񇢗W�:i������M�7�����_;�p�����@�ŷQ������ڡ*K�6�,�Pk.�v�1B�+��k�G�1��̆#�X3�l0kĒ�Ac�A�bE�o�HV"Q�-�$:���	!������Y�u�&�xn
i4xH8�՚���_�[|�6��������m�z�H�4���,�_����$�D�*�}��*��qv�h�Z��" esEk#�
�#Tb��������z�>�L�>�S�q�\XF���ntz�'���kT�Hk�F��w��]��'�m����� ��8kg��Ru�0B;а�X�߮��o�������}�oN�I��	_��`�>S?�̤A��6|uS��;��e�$f1cO��uKc^ǈM_��AD������[��#��N�L{���Uڄ�ٌ�>�J)�J�˳`7������P|�5��h��r�>��"^~�e���t���Д.�����d`�=F��S`���nb�ب��;�����+�A�V��c�ޓe7M�a �� ��X�N�A�a����5�Gc�w�6��Ȫʥ��'7��CJ����wݒ�����F
�V���C4��_:�aE�H���$j�����s��mR0Ѡ��,;�QY��%��ИO�[��-Ga��$4]haI��p�m�w�Jwwh�+GT,�~xK��<�De�m�蹈1v���ы�Ɵ:�_F�a*�g~m��|��3:���gk��e�s@�~�5���sCՉ����=幝�
�W���Ԍz�H<�u\�#Yu	�V7�U��6ȱ�m�(9�������}s����ӗ�v*u2�yI\��܍�����'쉄$�+\ܟ ��~�ʩ7,y݊(���*o*��[��ͺ���
Tkn��C�۵�0>���)�]�����K�r\�v��������U;��7�0c���oCT@l���A���JC&��EӢ��)�B�\�E����6��Tp+ C<6~l��a���0Cd��6�~xP9�c�|]��&p���^ĸ�(X$��!~}� ��T8􆅢��20J͟Y1��_ �S�W��ɝ���Zl��/c���!���呓!��=;� z�����#BD��Fݗ̏�A�eƝ�E�9�����a=�����jA9mc5� �w�6d$�>��WRp��Ϧ��7/'4�!*;�)�ѭ������6������Fjn(��hd��%�����g��̊0ŊDH��u/�<���!S���ܼ[�	���� ~�C�j�]�1)u_*�3~����������oEE�h}���4��7!7<\�f�C!���k1]�޿1�R�Q�pY�l	��0X%�E�k��uk��	
|qR��F\���A@�� �^�l��[%��K��A��K[n2�nF4=@6���uj�,lp�|Q�(>��E��Pq&\�i���3`�E����)<��IJ����4��
Y����o��(l��,��ŵֿ�Er�P��h��7g��+*rG�,��S�øsV�Uh�w[1 ~�a���\��(��\�,���O�y�E`�uA��{@�<BM{N��~4yb���P7���L�&wZ���%�[^�������qJ��Ό���|n�n?������"y�5�@�j�{�͛��/�X�"q�-�h��6�F�;5ؘ��X �˥�/����2m3�����G���O��Ρ����\�Xkt�&(+o�!ٖ��b>nD��e�=�Đs�P�a�q*��	�2��_n�\�Dh��1�%|��1��_%���6�^�d�Hp)�w��U��j+�3�w8�6O�����V�X�ָk��6+U��U]a��*�&��<.}	˔��Y�+l�a��x�7 �n����Ͻ#������~���z0���ܢ&�^�~U�	���&��Xv�s�M�J8�YQVT���2t(���wd��D���z{�:���!��ˌ�X�d����p��L�l����'�L�+8L��UU�Ȝ]G����hhX��h'�/���RECp,�
�
{g�)e�5�4buuVϠ�q4Ҥ� �,�d�w^��׾�7��c��.h^M'��φ�{��=C�G�M����E��LI>1\��=�J�r�D�n�~t�[|�h�������r7���Sd����O�{����V���y�]&M��k�[P'!(����E/����*�=��s�P@�>�I�P��U�
��޶X~_�o��XH�k�U�2LX��b f�g��߽�faS�M�|�h���|�0��� ���W~��0��1ǔ�%� o@��@��]A?������vߐM�Y\_O��.y�:��ŸqC/�w�Z	��*�G�ي�j}���e�$�*��e0�����VT�u��a�;v�٣��< ؃��O�P�>1#�zgV�3��W��giP3y�ga^&����㥗|V_�k�V�f� �Gf��/Nl�\����u���puі��[�_?^g�l���C*�F��~i�'P+i�b��
x-N�]��XW�P7B�Kv/��$�OH$?��9kst���j JM�?s�Bfq��v�8w��VwQm�â���	}��)�f��q-���7�?����H+i���QoH�sF5������MyGߙ��<8��L�R�q9L8fB�'�`1����S������}���SK����#�d��7 t10z��#��蜬D+]2[���"L�p�`N,��qcŊq� �c��C�5 �Q�&-��F祑?D��G��b1����6>��vܶ�ָ(�m-�o�6���:7<��<B>+k��;e/����R�S5a�}��qHB�Y�#!vzĭEH¨�2�N?�F�ỽ�*��L���z�H����
�ǻ%X�IM����`�Q�`{��p��?8�ۅ5C��rj�	�e�;�ف����0qEB�dh˙�o ��z^k5\u�ƾ�K�6��$�}��w�FK�Y��Oy���JX6h[j�w`��r�h��Xfݐ�i�گl�E��J.n?���n�`6,ߖ���:��|��4�l%�U<�@ғ<�h�����Gk��p��LLU�Va^��?Kfp�����G^%��ny��Fh7�1?�⭐���$c��g6���M��[��+h �ef����M���1���cL�@��Q�3q�x/к���9�����1����,�̆~ �v�q�Hn��L���}�"�(�����x p@_�g����"�q<}������0ӀJ����xї��!�"tl�'4�����#E�:x
6��N�~8]?�7�|�˸����y:��R��[.�������Yi)���y�>$��Y�"h����»H�=01.]:��~���/�Ӱos�⑕7Be�fc�������̥kq�^��g04��%0Y��%�@W>����(�-�5׵)��ª*%���(�d�v���x�����#h��\�$;�����<����f�����^�.n?z��&��݀z ���{���I9\"�n���T>�h�Vȿo&���Y"(S *��)�����/�3�뛏�T��"}+ �1�<���j���z��jc��y��='p�љ�zB%P�^��k\7Pv	�J4M263_W�93���w�`'<�y��}s��W:�Й��A��S�t��|c[u�!�b���x��o���&���%ȌI*K�d=��J��$���:�tԧ��l7E�����r�#xYа�B��X� �ც��˸���d��D�^[	X���Ɠ�0�`�[�+�#���H���� F�<�'@}w���^?1Ef��a�d��4�β���v�>(/��[���㽄���{-�'��3Kٷ�S��g�)��t ECt��r���ΎH��˼�����y[6cU�5V�uI%6}���NO˗]�*�����N�g�$IO�]�&���k !�ЙZ�����^�Z1gͮ��������a�;i�𗉆FV��f�9�[�y��~܋�֢�5�.��d��y�.E<�Z�0p�� �d���c_�����$SW� ����a\� �փ���B/����"f�+�$���fM�}��IѾ���P�����R���L�P���q�J�-.�{Ev�&t�C�O�����d^��Q5�7U��5��M-���#�E˖��N������k��x����+�!�ʅ@�viQ���X�G[7���x��U:�Y*%�d%j�� ��j��zk�ǎv�%���7�[���s�>( `�
/���dv�:a����l㾫�w�;a��+
3��[���$՘�R���Q�= U������A� �k�d���P��`؉�\X+����G�����d�`�T�8U?t\�K[��eJ9�=!$�57�p�V��.�UF`1cQ6[��H�oF��e��E�k���ؑ��C��Y�u��2#�����Rl�P�"$S<�w��ܯ`#CC9���Osb��mۡ����~��#���_`�	� z_�CP��1\4�)x{�*^�f^���Hs���(+S(��B��I�Z=Xr���,�4�j�������2�Ջ��N��N����I+���=�@�O:���Ҹ�<j	��!��`e/D�� ��ZE�y��w>��&��Ew0)2�)C�첋(w8�ֶ��a�ܫR�Rq�Ц1��L:��0�̟c��z���K�W��Mo���I�&Z��� 锖.��K��-%����m�,ǤZ�im�4͢o`G$��iD4�[0Lc�6L;8�|
I3�P�Óel)�zT��&msK���}�ɟ�O���E��(/��&�?{�l���爇�z}jf�xY��+���^�P��s7K�{v��`��B��q� ā:2ȩ4�,��jS��I���5mA�*Ib��S�	������&��H�ʞ�?�����&�0����n3M��h�i�!����D�^\0˳�ayx$����o����C��U/�N^�����7[w��hp4�a�k&g�6��")5G�G{:]e��9?��E,��>�}8Y�p 3�ܭN����࿢�W���J�po0�p�4<m��6����:�`�R���0����;���8�<��
�lNC�z<�1���KZ�!7�rS� �1e<��m�R�p}��a4�w�[���Yq4HU��3���S<؛h�T���XM���-�gj1�Q��)8p��RDS�9�y��w����h���ҟ�/�1��B�\�͊�^�kede�Lp�<	���a�/^bH���x;9�����w�Yݲój)��h��p����b� *�3�~�t1Ě+[���?��zj�I0�ȝ�QMTR\%`�~"�Ts�L���5ȭeO��nE��Rf谢u/3�X����%�f1��8��N[�>j��E+J	�؀s��M� ��f��o�}͉͜�ìo��DPx>t9(��q�o0�\^VL	o��>�(��S�EA�C�n�J��\#���a6�h,�.�c�tz���Ы ˘?S��H�P��;/���7�%+Bސ�ߘ��$.a���҆�g�^0���[��[��?��^e��}��C+_���������ߟ�X���|C&'߬�Y���e4+l�:"uLߜZ~�c�w��(�wf�?K�����NRn�� |�+D�%s�N�=~J\<��2ˋ#�e^���3	�������dp��FTTE�KX0�������b��	\<�]dӀC�A4��p@��T��=��)���0.��>?�_)�����¡,T�,�S����M��l��	e����܂����;���_O�
Ke�������a�N�\M�Ѻ�O�4LU�x�|���ʮ�&���e��6�����|�}]*\E�ʂ
c�N���mJ������g-6�ó��!Y/	X�@����N�g`ư��%4�}���C%���Y�ƨų����f���.W������l.�*4s���y�6jT�
��ֳ���:��#���J��5p���UȲQ����م��H�|�d'�ُ��+j71������|�1�sG�����P���#��ˍqP�{�8,�݅�� �=�[�~���A#����N*\'N� }���̾�"�svex�j�x�.z����n!x󀋟r�+|Į0��-�'��]�ʺ�xS���~��s�Bbk�=���.ߔ����Dއ�@.9'��+/���Si�MQ�i|�$Ǫ�MZˈƔ�Kx����l7ޛh�&T�%���ߗcv@D��3��%a��J@��7^&x3���ZO���"��]�"�N#��8L4�A,7!�]���w�����~�[��s�ACX��__�;��
=Jh���%��g����n�:C�:����D�J(t��ۏ_������/�/S0I��p��"�IuW��a��3��9��w�g��l�V._F�t�H��EP��X�ΰ��1jml��d�k9
g��b�
㉉�cw�����[�Fw����.0P�H��i��1�`�h�7�mB����
�uY��Wb%iuL]�(��>���,��KV�{��ڶ���O�"g����u~����5�����aj!�?IG��~R�X�X�ID�J�q)G�]����l<<a5�u�-��}����U[Hh�
ų���۰/w^ǘ�+��}p������'�Q7���Rj}�cI*�q�\��"��,3(������V�Xusþ����j�pcĦ!�j�*�)2Իe�ĝV[!�I�=�;����b}�|ҋ���+��n�����`�G�䤲������9�ώ���9(�$9��W��Z���eiǴ:F�$ܽ�f����Y�I��n��f;�,wvr^�c�n�{�mYz eԺ߁b6���׏i���:Ƶ^�#�N�ݒ#j�gi$����r�.mܤ�s��/% ��HpK�]z�U��{�еۆ"SMƜ�2����d�p�I�|	��r�ڑTq��"���i6�%L������K�P	IZ����!R��Ba�����Z{�x2�0D�R�f�2�&�K��M{��<���d39���`Y"��)��Ex�=p�t3/_l�]�6����?�u�gl���Tx<+q�{m%C��	UC��L�_D54�ZbH�g�_x>�z,����Uu[`n��4G!���.H}�Br�:��8�T��3�O���m�f7j��nVPq��H[b�����?��!��ܳ}�@�U�g�b�ĄI��v��>���I���S����Wi��ޝ����N�A/I��GÍ���I���l�x�������� -j��������������Ѵ���ڮ^��O�sP/A9(Iaw��U�q�ۑ)��z�搰I��t��sb@�=OD��C���N���!��� e�7{����e��oNq0�⛖�	��s)?�lN��㱵�+��Xo:*_7o>����O��#EYhp}��Zc�k��Z�kwz��D�/�ܟ������]�7�-@t:n�v`�mD��m���⬜�\�1��ݨ0��&�,2�m����t�w���pV��l�J�[�v�w(�J��j�EW�2Ԟ�jFc?9Q���!����h�pἒdg����ʠ�U���gݜ5�X�Km�B�*<=���~=���\X�`�v^�!�G��|��@~�Q�Yv[�Hg���
})n344��q�	���0FO����Q?t�nB�ƞ���N�\ޓ�k�;��p�n�8�?��+��Q(�-�K�<vL���Dá��]��!8]�R���J�FP,�o,Jd9�O@,o$a`�.ER]O(�/̙��c֯6R�8����'��௥Z4i=��ͭ7�{cM|8�����ڔ���Q�1$r�	ԉE�4��aƉgA�j!눈iq��v4�o�<��Q�U:9#�e�j��t�V�ҋ�Rb��-�_чoj�=��Gi�@��C����4���y�FQV����s/�1�j%Ū�t(���M;3��{Hg]�)�Xr�3�I����]P�'��<���JT�.�F�!� �Q.�T��=-&��S/e��P�λ��Xwo�Ӣ�y�8��c	�)tto���4=o�'�D��\PZ@�����r�X(|�VEւ�_�.��Ehu� ����f/L#���z.�.)�"��ex�H>�y,yk(�}ʤ�V#DwuI��&�Å�>��IPYT�}�/�KHJ�� ��Ԁp5.���G)|���Yȃm���Mȁ:A�!��?XK�R�bZ�q9�u���O&�k"�պ�g����d���E�!�8}��&�ڱ*�}��:e��v@㖰���Vf���)(�^�'��46܊?)ٴ��b̈Og����m������t���{��EFx�W�"'Rb}��S�-��
p�S)��Z$��Ź߇4��_��l�C������n��}��$�e������NY������Ig-{��*�I�*2���Ϲc6�����2�2���b�,nسO+�ފ�v�By7��y �WⓓZFHM�����B�[�Q#1ӱO
!cn?����z�S�8E�/�>j׵�$�{w���;`]���
�#$��/������.!���`<���c�6��9��'��e������yJ-���9(;V�F�/�^�l���J2 o���_Ʊ��S�L�<L�Ѩt*�B"�������>�r=%%����}{
�gp�vQ�Z�؄��44��P. �*������r{A�t�em|��\��a2��_����W�m�`�
�a�&�zA��^�a����x>���4H6�aX��5<=��!�sl�8�JK[��SRI*���JK��9��X�X�4�K˗v�ŵ6q���,]��e]�������g� �y��;�Ifʇ�n%"��{�U�cKf8�� �����+�o�y��7&�1%����
&/_�k� L���(�gw�=�rν<�i�i���3t�n7�5��`��%��B�p���e4���^���T]���9�2곢��F "WO���þ\%�9�r��~,g�S���`dn}|Wӥ�\ �}�+|ƥ��6�(��Em�rdŉh�'{���L�����~�:��1���R"C������[��j\��`5���v��h�z�Qu^��k�0�X��L��(�U�H��v;���7���#T��R�8�n���p�x��R<-�t���7�d�E���e~����
.�$9'�MU姶��r/��Ϧ�ŭ��!d۔)W��^�0b���=Dp�jtl8A�#�^}���= � �v�7�;�M�T�b��R�m4���y�HViG��XUX�ӽT���n�����kA��dh>}S��<���4^պ����/47�}��fq�c�}S���pï|�)��2��R
���oE'��RD�*�.����j4�Gk�A�;�/�H�ʼ�S�9�CPm����������F�-Y�=��E�B�9������H55�Ec��F��Vl!��]0^�A���#�L�<`V����گd�bA�?�S�p8=܂�Y�K:���^��]��G۴�M�{|�J©��?XG�`�6�+%7��:W\�&�L���p����t���瑢-z�h�2��A�������.����h��:���?�6w	�@�8:1��논��U}E��5���)>�c,�>�9i�tq�^��N�z�D�Ik�M$xlE8���~�/�"�޽9ƹZ���N:!�3�6|w��&��Γ�?2={@�:�X+ׁ�*��K�mq���j(}�X�X����oF��~g���bّ0U���'`ę�J��;�O̒��}z�]��n7;d��`��^{��ߐE�X�ؗ�	9��wt�� '���x"���%�\��oQ��0�[�KKE�*����G��n�!�0�Z���qLb��Nٺ$��W�a\�O�T����6��mE�&��:_��GU��&����E�'U���]�S��]74RY��׿��<�����t��T����Խ�ֶH��V��
Ѕ ��k*L�2�gΣnF��<�T�>�b[�*r�X�u&��}C�]�yi놏
3�%W��|Ԩ�цq��4�hT��y��g_]�;����ق�V&�(�DFr�`�b�-�PADJ$5�~~�U��x.����y�����F���MG��F*�Լ��Au�fG�!h����v`��-,�YHfT�s�AM��[��ر�R/� �Ly9�i��]�'�F���Gx�+_�)�8����Ф�����dq[������]�y?�c���M�಑���&���#����Y�U���i ���v�ጁ�;������_��и�r��;��y�O󰗝P!,W���}��؎�/��4g�.��u~_�؋�\���֢p���RbFE���]�d�H�b��Q}L2��NN舑���	��HK跼9��b�w
8�1��ie�8������>��H�`���d̵�H"��Ԇ��N:���Y��|l{g�H�҂n�Օ�A+G���p���D�m�D�YIK��1�k��n,���;QM���\N��IC�D X���
r��
�k�	�Z���ka&�#�dZ=w���z����7���48�M��Ҥ�*ӸX�?4h�4[�s�5��Q	r�k&F��c>a�<0n	��~X���ɞʁ�?���x������*+��3�g5�"��2z�ms�\Ǟn	6���������NC?߬J��sc[��oX-�@dR�83����k$c/�!J�����m�&(��鱘&���6u��p�T���{~�~�N�E>qJ- �ljgĨ�Y�à9�lV0[���ܒޑ.З+rJ1G����ϠzIs���к��\�^0������}�sc�lBH�ȲS���p5�H��A�7�';�����X��~��v��@�؈y���D��cMț��Ǣ%��||�F�m5������8�eYy/��	@7�t~�Qtk��T���3� ��P��p:�n�s�`�su�WV��ѻ'UG�"}bEm��q�:���`YQo��
�� 6V2�f�j#�w!�C�%���H�a�o_��W���j[�zt�b�8��#�cg�)�V�v�����f�X��O �tX��>hL�� �A�2���If�A���Bb����)߯Q��f-C%|�;�&~n����.��
�����Hz�Y�,���~	��J���C�6ٕ� E!�X׎M�Ng᷺�ۼ���f����6���q�;S�!�)yƲW���L��=�bH�r�r��^���-��,?U<�����x�r�jƒ�)��~2��u���/2�Jɕbrσ�>�����"�zuۂ�|�ey�ÌwCe����$�f�/�:���򤼔�Lj��X���T��pקfTLZ�y��rh?�Ǐ����20�N%���VM5@�'}Q�7u7��s�%��y�ꆏ+�Ow���J' v�"�Z.x�41M��Z̰���Dwx4\�|�FK�	)z�N���l�XX�2�&���f1���eV$s$�AjR�8\��7^�ګ�KIDAL�[S��>k��~ڵ�Kz��������l��K@����`Vq��/��6�T�Տ#���≟���w��9�����F�Zg|1�Hi#�;Fs�jA�T�P���Ű�gd�<�M8���cDNEz+�$K�,�
�H�lo�i��/1;�q�$����|=��s;��j�YHJJ�ga�5a�_��dx�=�9:	[d㝳�c Nё��W ��v�!T�O�>A���4�ȑ�,F.0�_�(��`���,}믭��ְ�.9^"$I�E��x��N��{u��!z��nA7��=LZ�dx7n���"=r�Ԥ5˾}�@����+������0�0�U���A�-2�k���M��>�������1���~��;I��e���eg�G;��˃E�+�����@��������n}5������t��[�u�ւ%�g���W��`1�ovyon��F>�<�4]��d����t��\o�M�I�� k\��@b�7�d7��K���a���@�l����h�f�ڱ��R��
u�7Ԯ�<�7�����2��	�=���U0D9�����8��_���11�������wڡ�9��?�D�����+'C�2��}\Px���y�@N�n�ә�kXW�&Hձ
E��@�!�4	Q�V�.r'�-����k+<�2O�3��U1��w���K(�nP���Kˈgwp/�`���^VQ�����]��9����-R��2�ݟ6�p�(����|�����p���A(XD��~�����'�wp��@�24�N�X��)H�^w���zi`5X�8� X��S>(�<��I�}�"�v�c6{~�Q�S� �OX�;���9`z�XQ,S|��%�-�Gv*$�y��/ ���N����c�� K_U��C5�ø��Tp�U���( A����z4��n���
��r;N$�)<�A{aG�T��Ϗ�'��~�8��88�C:5ܨ��;��롌���Z�췆�t�2�VQ�ء�ȸ1�g;pSίg %�=�39�iblN�'�ߢ.��@�[�[´��tR�C���GͿ�ZᆬFE�&
�W!�ϙ�[-��"�8F7�ظWxk
�^#b�	��N۳��J0��*���砯%�l��Ĝ�/1���$�`��%I�5D3DB��g���"��:���\BHл�1å�d|�#�,���_1I��i�P6!->s�`Ξ������C;1eT�a�(R*L.�ȭ�n����kٲw�<z"������Q_��T�H$���^��/�9=¯���N��R��Ƹطop�D�|SP��O�c��[�q1�V�Њx�6e,;�tg9�� }�g9��@7W���o2V �v衢�����Z&�.�uJW<��c�W�E�Դ�Y	ZƐq���v�┨�I3��%�;\QӨ_�K6�l~h) ',CJc���R�u��1F���f;���e�e
^���U�^�F?lo`_�|88�a�7렐�/%of��Z@���S�'���i��(��F���t���$���G&�o�(!>��fMC_���sY��6��]&���A(:�CSR�5P���(��B�}�
�?��?�B[��7|J�$q�� T�|um�����1���Q-,\ݖ�3�BH��xƐ��
�NG[�Q6��nB�k��tQ� �<���cDӁ�L���V���7�����~˃mTj���!�Ay�����X�_o4�X(��W��!�3�,��,��j�Fy!�:����
.s͓-`r� %�/R%j��[o��A.�r+�aRϖt�d(����:ǳrV����)��J0k����������P�4noN���Iy��2L�:�F���J�L�� �qu��!���-��E9��|d�3�E^�X/\����6$-2r��c�S�O�Gz��e��5Q��ҔauEeOu��S���־���5S�=�ŏ�i�]	��zB-��e����tBx�o��`8� 7
�C�>�G� ���vTzy��_`��V��1)���t�ѡ�/NvS��m>�Ձ�5U�bc��}����$�� Fx�T�<'33�:{A|�j:�2%��4�a�Z^��m����)%�M�ZB'�r��HP�Da�	������p.��.����p�P��^`�NВ�kk%
z��}%��]�T5㕪�i���k�w�z��f�r^	.HB\^{����Z�c���A��u�o�_3tk�c_Y��I����"|-	.R�Ze��/�VxP��ɾ���T���/;�!Ή6�WR�!ma��a ��h��}����5�Qt��8b@�,=����O�zMI��1q�jgg�u�b��hU��ek"��D�M:�����p;N|B���ջ<��gDf�{#\P��)�΢
9y�OM�wV{X�rW�<Iy
��iIա6�^��?M�4Y�`��6�U�S�u6�?�	�����&�ec��n���Y<�w����	B��}���l�*װE���@���ǻ\�)"�#��.߭i�\4��W.��,�B���ѫ[d�P����f'cX
~��e����/�]S`�o7H�����
�=��,��w��%*��)��W�%n�����J4̭O�7�g~?!�����9v0s�45s�(��+���vG%H=`^" ���D��W����׺\b<$l��Nb�qm�4f\���,�0F*jR��m)0��}�<�)�ֽ,�(h��G��G��o}Wo���x8P��ҽ��=f��3,*}�E/���VdZC�� �f�M�n��Ǫ�)xJNzo&�5 }Hnm���0mhB�TN��Hzi��[F ����i3�hP�dc"�H-�{}}G�f|e)>C<F���y�_�r�����]_B�y���|�v2e���ѡ�n�a�'FJ]gJK����"�n�������7Џ�|��	X,���m�<��V�=��qG��?���}�Bj�}r��۫V��}� � ���4M���4���/��J�0z����g���-R��WQDӔ1>%��mF��.�̡�LN夆��)�*�9 l�؂��ɩ�f����n���%�����;"�s�̬��ڎ�
��w��_������SI2 	�@+\����~M1��i���ة����"���8����ﲂ�٧q�sl;K��c"2�pMi���2ր2�r\��q�r3����9���r����/�Lt�Q��n�u{�X8��&Nz}R]�<����Zl�z�8�tH}�y�J����|�c�S�8S����O�M{p^.��Nl�/�;�v��g@0c	`aq무���$n�XkY
p:��1����P�{�u$m&��HW�����N$\��s�oQ���tZ^U�KT�Z��e����m�o�!iw'�(xG�p�r��ϫ8ReR��N���w,�Չ�)���taY��49<�E���:ջ��iRc��g0EY�.K��U˘(�k����ْ�VV��t!%�)�8��Y;�ۇ%%��>�TWܫ�4��!�=��k�i5����f�<��-�:r�:�`-9f�SY<@��9)�-�C�����z��N��aAe���c3����p�Ս� ��?�m�X����EԗJ�|Eh�%��$fᛒ#�$L\3i>]j�
`>��P�Ż�q��l��s��cA�Z[O��������)����Q�ъ�����}�i�'��zj�[���.FY�b���W�s�As���k
�h"h��|�h��)s��8(�u��2,T���q�޾�Zr ��G���r�W�@��x��j���s�5(���|S�.\���TW�=6�Ype_Rz���HJ�9�W'"����QWM��9��驗�!��aO/��,�s|�X�_5��\m��(�yq��n$��J�����?��������6щ2�hI��l:�(E��C����LL�q>��~�Wj'<Y��u���9~7쮲 ��_�֠�w���氁0��JO�P� ����اD���~zN�Bhmu�f*f��Z4�~�������D�O4�(#���/�������4�ޮ�^�8�{�$��]���pa��6g�K�eW,WB��̩}ET;����͵�����N�X���*�K^��F�s��h�D(�I�f��'H�Gm2�֬HD�ў��o L���7.�=I�>��\32U�D�	��9E}��4,�q�G3�~��ݚX
��(�E���q���qf�����݂<�7���,ʥ	^B�'%Ve��=12Kcl1��Tr�G��Dދ.�~*[���G��U��%xX �hϵ�vܮ�-P���"�q�[�MNe1w{Q�,n0@dyIk�Hr6G�pЄǵ�]o�rz|��5�c�H�cjå	u�����X ���]Y�|�N�N��������t�<�w��A9�?�c95��wU2�D0�W��/>�-� �ݭk�I~�g`=�-i�����q�2�`eg �RI�mM�n��X�Лh� �]����f���bR�לm:}a�:���@��g�M�7~arW�tA '8�υ�(��� b��I��m�ioȇ�a8��R��y��Q�Xk�N��p7�Eh���s�Hx�4���pOӗJ��ӷ�*s�O����G��9"�&]���:�
�zw�7_0�鉈�eMkkT�yg�H8��4Ak֛xF�&=����>l�J2������S<��g������Σ>��c���L#���6�g/8���Z��Ї��k �n~A����M�ܼ����,����Z���`o�T��gʪ�Cv�|�@�3Q�^xt�R"�»�ё�d�����V����P7�r֪.���ç�q�>�5Q6��{B$`иN#e*c��$��ʨ��Y^ҵ��?d�h��m�����%�^�nr�`��;�&�A���DRk�d��x��Y�Ė"AB�6�~��μ���3_���O� H�C^�@�Z�+�C��n��",���b���d�k5��I&=ta|� ���]"P[)^����$�i�z@H��")�������MD6+6�+c.�ɝ_�$���x����E�}�=�Q����7C{6�S����«**�Q�<͎x��S��2KN��y{Y�
hK2|�	�k�\DK�Ƚ��P?��K�o�3��cj.���J_F�g���I�͹P(y�f]�=[����e�xf������g�*�u�ݹ��|^�����6�7#^C�`��^��_ Ư@"������Rr�|�|�g�@�V����s�����d��3N_�b4�R�M�/i=�������1B��cO2���)%��\�ԧ��-�XG��[=�Z����\#a�"Z[���]�k>7�S�H�#'�	5���SR�ܦ'A	�oć���^�J���ϓ�k[	��<Ug�'ۂ6��^�`���F��>��?�쑅r	c�4*�W��ʿ�W�К�����N���ȥ�����5E�w�#r��7\�J�7��
2������O��n��)r�M<Ћ����;^)��؅�����<�9�������I�j�O���R׌��sS�!ᑐT:��=����{��m�ނ������ }����|��D��RȠ]{1F��C�xtj�r��K�o`�K4#�}J��i�z�<�BqZ<�s�O[tg:u��4-fB��A��la���Z���@LA
qc1J!ʫZ%�Zd����>%����IL�3d��Z��G���ۻgs���B.�Px�&��,����_�45��J���G��~3��H�\1Ƨ�Ep:�Ƅ�ب�o�a�ت�C��{���1M���;ilG~)�BeUlx�d����Z��;���\t Mwi��n�I\�ձ�lnI��}$yX�s�����?̩ܾ-�-�����m�������}�`��ԯ�C�4���B�����?	p��
h"�L��փ���<�,k���AX��`>B���'���p�!�M��f��Z�`B�*ɋ�<	������#=$�Q�d�ɔ-S�y���6-��!k����l���o]�)���W��3��K�%B4�y9*y��Ж|��)���$�n�ȾH:@����h����W�rs�!���(+�@���
G�����'<}^��i������6[&]��@D��dJKǷV��e��?�������ќ��x�=�佤�9�'����vN-C��6��F!�K�u��cg�����}fȹ<���fM�,z���Dy!o��U+?�Z�o�x/Y��d��+:�Ye9\U*8���(�Ov!-�������hӶڬ��I$'^kKu3 �X��5�Ny�Z�.�9U�t��O!�mQ�-%"��i�I��cs��ɧ�I�u ���u�u�@3��Y`��C;{����Vu6�@W���x��v�0%ف"G����5:�V�%��j�z���t�J�*�����.M�)P\�y����������5*)���%1ä��v��A��l���'����,'�J8��jʑ!���]��S�`H�0�����3�/O+l����!b�V��3����9%p���6��P��l⡣��r�-���/$+��WH]��E�� b6�Zi�Pt:���}�u#:[t���mph��W|�Il1��e���ٱ���$��dv�<�QkB���f��1q�.X��!|��$��o��/6�5�Pr�pj���_��xq�%�.�+Ƥu 9M#s(�<�#S�?��=�)�ݷ�������e�2me���J� �Ƽ���k��������YA\�/*�#���0�t���(��:���.:�/�\Ov����2��Z�Ky�~�ԛ"�60vCL���Iko~QƦ��;�wTؑ�"��/kvg�Ӄ�V��}a���]��ű�s��Α����}���L����A�g��y62�IMJ߯%3i\-�@9U1T!�Ľ�'�tەxOD�ʑ�̠5����tV@EV���z���42��H ~n�EB6�*�]�1Z\@B��S��T�� ��Z�ܣs�&�S�B��Q�^���05fʲ����K�N݋ԑW�O~u�k�� YJ��)��?����t]���Y^o~��P�^vr��G��бן����/�tJv� �_��_�*K���d�A
F�z�,Izk�a ,W��A�j�Hۤ܎��hy�Le'q�߲,�[�/�?E�C`<��H ��o~"D>��mKXl�c݇��.��M&��T�_JjZ��L.�x��#��#�R�G-u8G�;�%kװ.ğ�N�e˥B�#��Ъ�I��i�Ŭ�^�q�T�N
���{���îZ�"Ϭ�u��(O~-'�ڹ��C���^��/:r�2�q~دb�2A�����g�d]9��a[���U�@[8��zI����YΎ�>�]�2bO �(�׀�I��hA�x�[n�j��h�N8HG����5u7�o������ �k��]� ��u.y��ǀ�G/`8��O�9Xq^�mq�:���U��6�QR�Q���`���e,~���N����	�F�ھ�SuX.�����Ac&�E���u���|�[(:)�:��`@)$��A�;h*3àtÖ$�4��Jx�6��P;�܌�*�q&��T���U`ؐP�I"�cS¤D���8��c� �]h{�Ha'#�g�U�k�	͈	�o9 ��] ����xwU���j7b���<�@�m�B{y�0���=w�Z��i!��nZ�k�1m%�3����FD���:�*�Ɯ��e�u��b���੃0��x��Q&v�qFǝ� M����Ht��f�+�
wM�֔k�4�K9��Aɐ� �ģ^����LJ�(0��S@ރ�e�bYR��A��+�MyI���,��o>IH�cz�Z�R̩-o<�FW�ڰ��#�՟[�3��跄�d�(�8�P[8G|������F>4(�-��� @�^2/�V����^m"R�0I2��ۨy��Q���	�.�%T٢�q�h�i�NeΏ���nB���(�y�~3[*����5�ʝ�3	�
�<bފξ�_0^��G�B7}�> �>υ[���Tl��_�N��-���:n��1�jW*	xؾQFkH���������P�����/:��W|�b�'���g�	��C-��-C�N�<v�s�O� Ա����b3��b�J�Fثiyh-���q�GZ�
�r���tM:ʳ�� 8I"�������4��'P��t��m��1���R�x�Qbs���Cy��'i�E)Yi\�$��%�k�g�'�j5o����ja	8�c��"���v�Y�ɅE 69��ʜazə-�_�Z��+�[�]R����u��6l>!"J�$X�E�53�A�#F�L�BE���K���F�+|�����Gٖ�2]�X���[�v��i�1��6v=���Y��Y��MC~��q� 3�F�s/X���-:��N��)��d�a�2O�גq8�S���BA�9��:E,�I)����,S�T�^i��B&)�e�+�gF���x�ח��j�F�X�>:rWooT��ռGo@�fO��B�����j����6�(�'\�c>-�l�G�5 ��1����X}64<n�%��KNn8ǁ���YIܴ��M�9>5����"C�9ud�ϫ�����U��F�
�������]���{��@�P�����(�:�����H�dv�	��u�
��]E��kٜ>���m�h?�О�w~�`0!�'�*�����c����ӰVl�-��ZP�ogɵ�=��ՠ~��*�z���V�%p%1W>�4�.��0_��{&�b�Ogj�v�C�ŗC��{ط;�m��`��1��|`�̌�0�[%/Y�K�]*x��}"�0�m:�V�����}9-3޵;!�H�P�p�~||m��k-��vW��� ��L�\%��-Ж�,k́�݁c���� 3�aIB�r*�5k<�35���ۡ�=�&[t~�z�b��ґ7�|Yo-��zc��������,�Q���`1�J�����d��jC��!#��V��U�8E:�����pz���%���+��O4u���Gye��%�T�l�׷� ��dKxi�tZ�?��^a�ǭx�\f1{( ��u2.�U����A�|jK���G���@8Ӡ��\�
���.%����XrUb�I8یD/:��[KQ� �C����S�:�G��K���3��X\ut�f�չo���h��@n/��
�$��� �9��%�ב�!L���[_�=�ߐ�.ƀ�{�FG\S���ڏ���!�BsJ�7ܰ�� ��Ь���ǝ��ŴbmaMD����i�$�w���q�H�C1T�1��fZPV���Mxx���tV+�E��٢(�H4�E�&��D:��/qZUDJ�;�~Z1�����)�{�D�����jJ]�;�Vg������xf�����a_p;yR:7�s���HUۍs�*ر˃����n�� 1Э�N]�o��v��b��p�H;��n����@��Ѷ�k�[��͚�q�{1|�k����]*��*F�vM�X �_,`2�>0Z��/Qx��nQup*��ob���+�D���X�;�Χ�O�6sЇUb�!�DN]��-�F�G��l�N�*<s�+.`m����B.M�f� �^��Ȳ�JK�x�fc��S6?���CJ]�`�m��fy(}D.��
�P$Dzfq<T#\ߛ]=�行gE{O�d�/��A�K���Fr�7}��}GJ$��2I��l�14��.�;�RF64=�ݲ�އ��`��䚋��˰#��K
9�M'�b�.P����QV1�G�%E�H��᠅\�Kc��V�3f��6�L��),e��}6o����m*�Q@�`�wv'��0kR�b�%�O\� �aH�ן���ܲ�P�_����Ӕ�eXw�Y^b�T��2VJ�R_���Š(!Jg�vK�������%Ox�������q�T	A�0�-��،�G�^��A�@XA-��-ձ�Z��%�(��GA=jD).�{}r�U.d#�S{xX��c�_b�(9�/c��XXz���h��^rT����=N(�/��P؟L���NK?�F��C�'i�~1�A�b!���@2:������G�i����~�o�'��#��������Cv�[J�1���a�ߟ*g�_��V^�ӗ#����&�[�L
W����	M�K�+���iT�ҫ� �	��ʧ����<�;$�L�X�!c���&��]HN�0}k�����xݹ2�PlU{�9�����<Ó�����4�H��
��T��T��0o���8â�i��FH�Y�>�r"�7�������8��B���FV���3�㒪��jH8���:�)�8���'A�{�Z_W*D	�R:|�՟I�X�?o������:��+���V�=!Y�s���b�5��"��r�z��7 ����v�,�e�JLg<��n�A) �݉�fh����ֵ�X����}�1�N�фfd*Wf������I3��Fw�{Eh�/#6�*(�Ć��6��Nb�<�ș\I����� '�;u�Y�R��W���~�T�!�7L�V� }O��q�ߑW�	���ɩ�%���q��2�T�����2���=��4��Ҏ��P��4dUE{s�A���ϯ)ˎ��V�������T@�f$�J�-�(��o��SjAG���q�Lr7�(s�z���}�Dp�c�9�q�\��%k.�F�Az����e��\���`
}M��s��Q���$tM`؄]2�f48�lA ���4� y�-5ʽr��`v�v��`G���B�Wv2��\ZH=`�?")�J��'-E����&L��ZH��=�鏽����W@��W�&ϵ�]�%g
�hasY�+�v�����(�&�0H�ٳr�_)*��"6	f%����`�Y�Þ\Dw!i'��4Kj`Ro�����"���wo��;81֋���%�i�!��W�TlV��sRp�&�Ju(6�Z:�&�'�̽�dڡ�,�s�^��撺	i����F�b���^',�N "���D�?įy��%I��k���_�� S	L���O݄�B�6ԅ��|��L�F�!-p@�J�c�(�c�ڒ�m�X@�#(�C%��-��,�dD�X�(L̏^/ƿ�O?!�4�/xJ>�{��%e�ށW~� �I�B�(�AϞ��Od��=��{���׮�*m����h(xڲ�/�G!��)�|)����$�Ԃ�l��bҬ�?�O�d�7���Dls�ʇ�I8v��5�|�Fjp�ݨ�EW������Dux�f���!F�9�VXhr�����,�P��_�S�M&ΔC�k�����^f�ZP����w���p���H�J�=Ys<�X��+"6j!���R�H������-p2;�D%�n�	FZs;���JF&�@��[b�,|�5i܈R��z��[��l�5��#k���bH\\ �"�ahòmk�R�ck隷d�<�tUM}����3Q-��d�����'��;��Gs�k!�!��5Y��*0 Q�����L^�b7�H���(�m���_^<~�|}덪�D� �D���M�gh70���	rB��|��r�ηB�,D9]��e=�ȏ��-�N���O���'�+qgR4+��y����
-k�^b���D1����{ק�ZJ��eu��EBw�1(�#�O�+��2�����i���5�Ad*��E�/,!�-�a<�
���%�p��dW-0��M�1��2���ݫ��� ��&vZ�|�O��)A�z�h�ȍ�JOtdJ�Q#S$��j���qUЯ��<e͍]C��w���sS���p��im�3^�K���>n�ڧ�XO�֍�|�+�[�c��;!�ǞH�������#��4C��.��ƻ���A>�}����_gdFPd�]Y����#:�|�i]����	�Tcc-�����ĂƆ��[�JhG��T������ꌦa�@���.��B�$˭���6zp��z��^X�A>�������G���X
s���~���)T�s��Qr��R�R�%La�FqZ��i� ��nC��ؒK�0�*�"��'N[Qws�ٯ�ha(�y(�]|��]&L*��&[ނu��h������?��0��X�tm܍F�;�)*iЉ�r�a�>���fAϬ!�[Jېe��=�a��f1]�<������{��?�������X�,q������9�:H���w%^�od���z�6��f�	��@&��쏅$����C���ǌ�ހT�/���[\��I�C�1�ޅu���Tid�:�aO&9��t��2�(q��s��[�-�T夂�� 5����~YYC��4ttw��O��`M��D; K������h�(P�U��X'��U(���FwD��1��B���X��o�J��3�x�q�����+7������1�\OB��Yupʆ��Q��B�Ô
;v�˞��y��c�{��,�j����g
�'��3�I��ET��~�z���ܳ����k�Ą�xz5���Z��p�a0�ӝ8E�!�4�1����Ŏ���:V��!}AY�����3�V����:�s:T�_y��UMJ@2����U�~^�@_w����0��O��#���I�V�H@4���6���:�@�m����6W�ܺp�x�_�O�f��U��]s�Wv�ޥ,�EX�Y����P�����Tx����<{�~�����'�q�#��_h��[�6)���V$��C���$7LSv¾���F)wh`m(����dV`,�|͜���[e;�s ��p��HW�8mv��	KxU4@.�����w�Z7���M�G�pwG�F4-���$|R���\����7=�"�1$I��LH�+,�W��H]����� c(�m����[�K�OY& �w{/�䠣_��_��",Ԛ�`D�e<���|�I�V�.���:ö)j�<�1a)ڊ��+k��	B��3:�B��Ob�M��w}�Pa������>�x`�v̹����DW��iF��6���
�9���91��ut^�8B�1;Ԩ�A���~���N�����ͯڛ�P��"���T=����R��|�I-���n��X,0'�HQ[���.���2ł���-h��>.��61�Ҋ�����&�e��.O~�	+�j�2Rm1���b�}�]h�A�\&�Dh�ݗ�4áWZ)%9{.�D����,�oX@R�<�y��Uj�� ��^/^F�U+gv?[%���H�Azĥm������{o�v��e^ |)��3�+��A\����2�-l�����Ȼ5�E
��6KxP9J��:��5�)�W6!,�Aa��ķ�wA���H��`�{�@��<�ph&IWh�'p��֚FfxA���2�?�,� sJ?䘒dU�\����R��]�@�iu�,6�7J�$�0�	m�-8�4�0^������H�{x��[ź�"�b�A���-���m�ox�m��s6~�l��w&Si��p��r8��U3a�/f�?RO��GD�
x�`��$���M��ubm}�%��L9yb���������]��p�M���1qʴ<� ��d�ڙ������ ���6F�D�������k�+d/%zD�  �#3�� Ia{OG����~�h)u��L#�<��Ǐg"���>k�}-W�����N;�J[�u�H������ѭ�Zɰ�{6"'���LbЈ����#��X�Q����+V�sv'�Y�̠Z�Q�3 ���a����rZqO��rQ]=���+S�O��X�%H���o/��]^}�����li�L|����Vϱ�c@���	(P�7x?N���z��v��>��o�'��Z>>f�z`�N�
(@P����ʜ~�Jo]�\'X�G&��
r���w� mn#=�X@J-H��5�>X�&��=�u8%��7���9��X���K4�f�FԖ�p��\>[X���G�I	'{� ��KO!W�l�������
ڸj���!���oe�� ��t�G�HZ$��(F���Y3K(8%�pU�Od��,7�O}pQ"�d����v	78�ЋZ�G+jFy�5Ǟ�ݶ�$}{�"!תW�)�1�sg�|��������,�T��F-�:)@wcJf�Y��//��e��Ł_���Ɩ�R��%%�HBߤc���;`7�c58?�-
O
����`W`1QE�%�$����>F]�ͮ�R��}�L���n,@���E;*�|�^����˛���t���d��,Qg�=��w���yѫ����[�_�d�Y3xY���@ʪX�!��"��}2�oz�\@o���X:b�F�&�E�Xl���<�Gb6���K1,�jZ����W#QHyVd�~�iL�s>|��9�.�c��}�M�7�-�]`����4�>���`�)	c6�My�'v4�
T�^]:W���^���/ݵ����p(�97��ڕ�v�|Y��0�`�2�y[���A�k�K���_���I<��dy�����E%dƎ�y�7��J��Wt�#1ݴ�<q��(_{e�ނq�B�,쟬�!��d^���Xm����i�^��tM��2S��H� .r�{��T����w�uO���^���%�J;	RloU�B�ٟ%\t�A�r���i��W��]u�˪�(�!���ϝ���zNr�̃�U��U<D�h�fP��I�[A[�P[��\�3��U�u�Fw�H�Ė�I���l���Z6R7?'��\X*�G;��y�Q��lH����`�
OJ�)��Z��V�+�{�����>t��J��>ۋ���qE v�F�J"@L�ƴN� ����Jtp���A�����XI&ۅ���U�i5�/1"=9FxQl`��b*j'TΟ��J�H������]��RE��x��<s��F�f��0���[e?��C��Yڄ�p���֠�2��?!��V��-"o�]�CX�w�8�c.'~0���N�i�H��RA��/��F���K�?w�6� w#L��k����d���*����|;��TGKbE�2�<?�*1Yb��@����R�Q���W�1sP��b�w�Z6C	kڮ�J� ��tֲ���6����z"��Ӳ�E,��������]�(nǅ�|CG������%3�*������C���g�2�ۇOx�S@�DŇ�
�&�Z BPp|f��^�Cm+7?+M$�ň| �8t�@nzuH��4�<��x�Q���p?�4�0Bm���u6�<:����щ��^q�Wk�g��#�C���^ px���^!���W5�=����R�3M�@n�;ت����ҝpJ��\��J�ϻ���ðZ(�*L7PNt��QN��-��bV+ʚ��s�=��!$�3��_݀��I��bq�l�`���=�3w=G8-�(3&jC�ѕm_5K����;З0��⋥�η%:�٨P`����a�B����,3!N �����{��7��W#rM�eF����U�v���E�?��UU���>�ٳ^�Mp�x����E/a����X:en0����'�Y�$	��Q��HS�Wz�K�1���p�n�SM�u �0�a�
O�9�VgŔ�W�&ŭ��M�[���I�6��K�ʔ�=����B���wM�����q,ۧ���l�\�^[�s���B���F�����z��V���2��7�BZz���*��
���!�XK�b�c�5Qrz�Y<A�љ� ���d{�i�`����J=�T>�ۤk��MBߠz�X��Wʘ�������#�OF���pL��ZP&���=�IG$��n��D)W�DX�ϛ7?*��o2gw�DБ�gP�ed�۔�ЉS�v�T&�)��I�wR��q5#�S���J+���Òz�.�@kI�}�H��X7"�-.�/�V:�/�2\G��U�Z@�齒ҕP*��}�p�!��W �v=t+���)Oa���͚��:Rb�&��ۿ}j�Y�����_��֣�X���uR�s#��3B��~��G�#�u������q+m�K�X�s����:76�����d�-r���Z��oH�h�gK��i+�l���SE�b��s��)ia�����9�PҾ�<ѹ
0�ȑ�!]�Sܖ���}�3]s�(��
�[x)�.�%���]y$�	�!`����SOw
|ܲ~�6}e�؋B��O2Bگ�����7/��(K��� V����[�����wJTqJя�/���6{��#���3� �d�5A��A~�i�8�b�k����\�� ۧ���D`g��gja��==]+����ߞ�闈�G���{�n������z ~���b=��=,p�	���RI��*�^���� Lh	p|ȪP��� @f��q-	Zr�Ў2!���@`��������eՌ/o�G�@_R_.:����L��Aݷ��<����b��A�$R�ܞ��r��r�\u��4�F�`�����	�و��5W�v�y*�F�3�?���;\:�6�*7 �d�
������7,_�F��T݊�
�:!+��3b��ke��gB�_譳AC=�h�(/�O��YU9�D�藓S�y���H�w���!p0Rd!�"Y�Y�VPG�Va��Ö_.;�#���t�.�)�Ǘ�D�$�H�gd����/�&W�,h�˯��W������@m ��
�]v�/�$,f?����>���{ζ���)$��/4�E�\|�����,�~��D����h�x��0���r�:���A�Fy��N<8'��G�A&���,է��Xaə<-���ؒ}�`�3.l���q����JLp�IMO��&~��5j��O)�}�'���\�{�#�����;�s��hY{
� "@v\c�}mb%�����tH��ץJ;C��O|y�3%�G�l4�n��_��m��@���>��
2�$d,̆U>{���v�lqu ���eϜ�eiT�m�?'��:�,�;N4���j8����x���	_���AZG��2$����� �[ɚ�eߏ�ww.?��O|������e��1d��ɱh�;�)\Rҩ}ȟ�����Nje�v��O|y�z93���q�D���~���� .	�:������$��r������M�b���\}�5�\,�����u��1 Q��Dn��)2���4�s�Mz�d�.�E1���_%ƪ���Aq�g�/#��@��&�,b3h�<�
ՙ����4|)'�x[�I��
��	�p,��"��E<{���cH���!JPq���le�Pm(hr�K�(t�2
I`��.��}�cY$��%�E�����xQ��{��s����V��8�!|����c�s@���&7�&�+|�bG`�
�NG"��
�p"s�{��]��4����fڋ�f�k�9[�xe1��$�k_�q����Ii���8�<�DN�IC�#3�t;���Lmƥ�����b�X�҇V�7�rM~��mE�~��zU�L���Q�u�DV�bd��o� �?Lק���`7�������mG0�����XH��i��V�w�"98s[�f��IZ��Mw��ag%=0ֱ�Ul�-S,B�(β����OF��=	�)�h��lQ3Y�<@��Ⱥ���TA�� .���{,�HϠV�2h^�%l�
��f^����|�ΐa��t�d�@Vg��$eA���#|�9Č���ρn�T�F�>���hgl�(��p�U��x��O����ra�2�j_��n��#��?1pG����V��J){�ճ���
��F�*�2�����h�M��sy"�,���<�e�tV�^�=�3}B�=P��:ZD�d6�w�R�3vw���r��<fW0�<�/� �l�8=��E2D4����)�"\���^h) z������]n��R�kF�}��_PT ��h/3	�p�m�~�nY��V2af�n:��mB�������&N"�+�� �4j���˹RT��y�
�f$ϡw�� �.�P��zd$$=ƜxC��*��+���к��)�&��4VC�)�~�k��(����8�\�P�8�;9G�9�4UU=\�>`[�=��]Q��z��r>)��,#��2-~;���?fsY\��*�T�]�N.�f����D�Gm'�7���V���n���:��A2fk��nݪ�����B�L��Aoz�u���t뾊��	7<����SW
���0i���]b�a	�~�Hm�9�B��y4UqV����c>���I�@Z��ދ���m�O�oY��dX�@*-���bɝ�Έ�k=��<5Y4lgbP�~��H��+C��Y�/?-���\��H
�r��5yL_�je�����+��G�lc�w�qE��x@�o�=ˤ\}W�Ko�H��?y���sv���[ ��'�H��S��|�i���^�pԃç�a��㪹-�;1��&�5Vl|�,C}������H�q���POc�A6î��P��q`a�Y��5^J5hB����9K)�뱍�V�8Do�5����ŝ��~���qu���c�;�Oy�GC
L1Hu��z��
q9��h��k,0-y$������o�֮��P����^��B�E��.�$��&w���^��/�kn�o�������W9h�}����NK�^^+i��`J�9�F�d���k5 �Cև�,�����^w\�bO�����<��P���GF�Q�Gȋr
��7$Zy{Ǒ_X�<�|۲�LU�fX�B���#�X�ӗn*��7���,Ңe�5*{F�o��˳�X��a���G ��9�A2��W4д@��i~��c�A,���0�H�Ai�]��#�z&�9܆����!��)�~��z�\o��㤦F�9�>=}G ���	�*��f0�8 	�����N�}�I�� �l��	��~���=�J�&�A���e�a�}�q8(`��7�/"��Р�V^���2�;_�j\_���B�
]�;j��`�?���������1w�C�3
�hݪ�V�K���ͼa�ƒ�����B�t�����U�i�0�Ю�;E�J%kO06�۰�̇�6[ʣGq��{ȉvir�4d2����X�����F��N"���r��~��v��,\�x��5rƃ��!��G���._i�sh �A\;�d���'i1�����􇎮��D ��������V�zJ�?QÔA1�����v�J~�$�[;'��`n��ߨ{��P����������F!_�,�A�1~�L]mQ�v��)=�?��N(�𫚟1F����`�5s�k�IH'��Z/�xíH�.Rv�����,���_��^�G�pA�(*�p	����^߰���gc��^\M;� � ���@i�<&_�Cu��..���v������N���`'D��i��U؊9�稜�P'O�z����Į8���l�",�[���Gc.yN��f*�-(fL5]���R�AU{��
�d�!����)���$���}�_�%M�~}ʋ�V)k|O���ԣH9HtN!��­8�����ě��ʨ&&��n��#��w��s�	�,|�Ƙ��դ
o"���&�Q��g�i���o.�&״�>7Wy�b���p8�-՜v��*��4��6Oȃ�����5f��^m(��sl�d���s���G%�=1��VF(�!5M�r��R[�.�Ֆ`�k"�a�%\ b���������	�ǫ@����A&_�^ec6f���i4��-ܚ�7ߪd@� ��!��ctQf�ߚ>Yw��;o0�ڭHZ�����ڥ�V\0A�В~��[Kif�b�{n#c.���"�h"��(^�nFc�,�r�K,�YJ���Y�I���W��M�A@^*P�� �< �b�#�{���5F����pØa����	L��d��̊�k��,��z�6��pOm�S�y�b4��<v�Z�y%�1r3T�k�56q�G��nW�Z��Ce����2�aU���.c���8�>n��Ig|!�G��`=���$3�Ȼ���9)`V+���P3 �'Ȭ��/�g�!�7�(H$�k�v`\]���f*��,�S橧,?���'��1��9��m�)���� ��i]��7d�������1����&
�X�]n�p��.��f�k�:�B��>�C'cR�o�%��إ��3��(Q���رk���i���g�Vp��1�6'��[w��gV�]{y"���!��a2c`�h�3�6Ob�������P� ���"7*��=䷓��T���n�E�L�W$���ӜOc#J��8i���>�π�n&}V��=��O�DvqR�z[x	�{���Ǿ��LQ��n/��4@�{J
l8I�׮}z��|C�C4��U����JR�ȸsu���Yj?����x�?�q�X+�ixKd W����ս�ٍ��
O�o[؁��G�$&���.�� ��!1�%l�9N���0���b��`O�/B�J������Oy���R������0�^�nc�R�(���t񳥦�3+������J�M�� �;<A���T�eTߒS�ٹ�(vElg�J�[G)͇m�%�k�]q�v����p�b_��8t����Ñ[��V�}��+6.��}�C��V�%(k��� e/l������	��$�d��
�u�K���Ў���ν�/�;���4* g�)s� �1^+\ʉ�ӄ�:���ץko)_uV�L_��8���Pi,�sB��'����$���Z������șK�\���O�K�#q �����\V�S@gO
>��$�**góV[�~'P�,/��>�dCeJ�`H�t���E��r���({{f۽�_D���,�bF��5 \����k��GP��ږ�U�e������=7RC�T"�r�x���mx��[��hR'r���Q�1=��1�Vi�S��)ijY�gLN��V�7����4RQ䳖�8(R��y��?��:���3�]�B. ���	�%w�����Ҹn�ϱ���D�E�G3�B�|�lB��]I�6QS��f��~�t����/ Em%�R@��#ܘ\���f�GF��g�:l�hi�#g�w7A�.��'����Vg��L�o��k��
7,$�Garm��	��#tڼ�����8XatAW�ŵY���
M�1����@2��	�]�a?�:�<=.�I�;&k��Q	u�E�1���+��T���}`N4I�U�9�����ݏ����$�3���$��0XMhR�c�@R�.LESՠlі!4�c%���^�I2"HǳJ�kwr����J�rn��0ڟ>ǂOm&��[�c���^�G��C&Y�ќ�5v>�#ԋ��kQ�\�K���,�(�eJ�S��dn
�����ρ]'&G����p*��]�E#m+Q�����2�"��3_�ﬄ�^i�J��UQz�����3A`A��&t���PS��'�~4��c;3�P����B.[�F�n"lk�+N��9-�AII����V��z1 �Z�L�N�ҏRzrxAfMW7Rݰ|LI�l�D��=@c	OK�,+�rV�L��E�4����`�]���e�AA�%�� t�����l�{��u�kAF"o���7)�j�o��u9D��ذ�-Fu�W�*!�|ޣ��7��`���
��+������M��<��6�+.�; �I�N-��^Ss/R8����H�)mXZ*z�'�;5�~i}���k��?�X����2!|���Z�{�VdB�ӳ����������H��c�R��'��f֩�S�v�쓺[+
X}/����"�L�o__��A�aC��#�����̷n4����&����+�����M����>�aP��j���[n�ee���Q鿐�J�N���̸s~�6{e�$�s����E��[�z�a�[�J��@ϴ����	
�W��W�q��,�F�����l�*
����	`�=���>�~���܀:��8��q� 4�������D@39�*���G���;�qUI^
���k��[9��M���$��Fp�e@���&N�e .˓��L�h�o�w����H ,>U����)f�3oD ��A'L�o���T���߸��3<��F���LGuY�@d}/7�՝=��?�0W��г�J�P��ڒ������J�tI{�>�#����`�ų��Ҕ��o6��9��hJP�!�ٶ�0�㌧eK1@__���u��\��cX���*�r���ʗ�ti�ŵ�{�BЀ���z�f�Q��嵴h�'��5����5D[g4�޷��������U6}��'�0^��<T�ڗ>sgC��h��&������D��k��j�����5%㍆
�b��8!��.��YЄܰI���4����R�P���;��f�E5O���s��� �: �$.�2��ے�|/~|2L/`��W�H"6Dُ���
��8�V�H�L��l�C��P�,�\=��0��R���`���Azwi\�|���v�+%��	����� j�
��5y9��끫�&7�����o6&�:��h�F� p[�KZe1e�J��P�kh*��)�a��u�@v����(t�i�c�%
En8 �
X��x�#-�j�Zy(���$;'?�U��p����Q����	�=o���ml��F�c.棉�sqƆ�`���t`l�Q��;�bL:�v@|��B��FW�a��1��(�3D�W��k|��7ہ������1;.L�yB��6WzQ�8n��p���[�x!"d_4W����67�?Ch�I٪�F��zR����n��4*<o7��h�|�=��oVFqhU��=k�_��?O���da� {��} x��߽6�01W�ula��V�����0R��UXˆ��,��Ц]�mB �e��l���1c��N/�,bY���hs�W$��Iޟ,ަ�=U�Ù{gb���!��\�J �K1�ee<������!�����&߰�!E.?�a[���oF��2���I�A�޷�1Vj ����ְL��RP����p]d�G��g�}j����_������
�2��L��9q�ޭq��#��BK��b"!X�d���b�c���p�` ���kSC�j�i��x�ڬ����*��0 h���iTl�̺֫C�!OZr��F�\��Ԙ�:�b�w ���4�y_G�R��R5tV���x;B=���q�͗H,}�V���L{_��Kg���-�1\-�����5q��r��Ӫ��hd�T���7Hz�"O�!O���Eh	���=��"L�r�-=�x�0/4��\��ͣ�i��_$I3�u�kR�E���R36�HL���I�7�'V��e�Z8�g�eD���D�B�k�i@�܍�O�:��6�姆�Y�{A�F�G�S� 	��ʁ+w������1Tck���9�(�����_RΙ����K;�F�r�򠧆�ɚ�����20��3b�]�5��,L�?>�����{���#��Vbq)���%7!�#�E����}7w�����@,�;��M�#ܨ���`�F���o�����|�����w�ֵ3�`x�R�u�&�(��ܪ����@k��ʧ��VQ����� �t|�%>4E�3��2��Lbb�ދ�����H˜9��E��>����I5�i����	�D��w�V�a��b�Tϣi�dl7m�Ь��%)�p�}�BR��t�h�ƽDX�?`Y�$��]>��)9@�:���rU;����=�Ѩ('�~�~�pp)iت?�V��;XCo���@\��N,^���^i-�X�M�9���	��.Gh�ˬ�-���Qf��������H쓯��>,'�T���џ�C��B��eFH�[�z8PF��.8�y��A�![�^���'.�YAO��vނ�0*s��jwE�
[�<"�bb���ܡf������]���I�s~+TL�14-|x�K,�����h*޾~QB,ѓ�����Ep0��!����>R��ݤU_�K���9�y�YuS�ѭ���������(l%y{:�H�lΫ���[�t�>�f���Y���z4g��#��Y�����fF;<�10[|a���D٠��@���(1���� ^��ĐK�ʽӷ_q"[sz&h��Ko��f�|)-���@�ܯ<:���a��٥:mj���0��>'7��K)Rѣ+�����?1��-�*�Ħ����X�ɷ�>Ђ<�[F�Cu�;)��.d+z�ܐ�Ib�ʘ���D6S��|{~�90LsX �.0dx���g{nB��o�h�U�F��J��@�FC�)����\�ۃ��WxxI���E<���u06w�Cڳ�����݁��̯F�If��g��J'-NH���(�[���`���R�&�	�Fw\��G��Hʺ�z�U�Õ>E������vSзp	��t�fhƠ��2;�)�*I�N�����l���ll�o �8YW�w�b�z�Ӑ[j_�Q5�5��<��3V%@t%���8�LB|s��	�z�z���8�T�2g �Ot��Jj�^b��c��+8��xz�d��fk�B\V10���x,/LɗQ ܣ�=���c�9��` ��� k�{���ɸ:�C��I�S�ʜS���3�5:Iu3n����Sq�QB�,m-�RZ�I&���o�b/�����yd�_�<6˗m�&��<���q�܃�Ԑ�w1�8;3����G���5�#LC T���g�=I{���'8�*��n�]6��IÊ�saM'*��31��e����Vʆ��D��F�3���;�xs\���ab��tyUw3�;����o�!V�XW�,9=��L��Rк~gxu��OE��8�VZ�P���C�YS��\\�Ւ�Fp&|X�?���@����P
������>�Ĉ�����55Ԉe���Ѥq�e�3���X>a/�Pp�N�ԭ�A��U��D����ft7�Ly�Χ���	��l�&�����K%E�l��1� ��A�ʁ��l�\�ek��4�9r�"ݧ}!��Дk���ؼ�&��tz�/����T�������biLs�So>f���e�P�1	-��J�(Ux���"��7���pL�2iҋ���46uF�[`�Z�Do:VQV�IDt�>��U�V:��iYl��wM,��c0"J
�$�~4��5o��Ck/q�B�	<A�\�ȿ�.e�I�䚾j�aM�W�9z"��K�؇�yz��>�X�UJTI���Ԑ�L,O�΄^����Ṷ5�N�Ө({�qR���ryat�o���]�iI��QZ�{9���A��%5��!gu�+���b�R�	ZUQ��I	�7��W���P���X�Z?	����L��^�/e�����z^��� �}@w��.Ąs��S��B�ƻX.�v�!� ���q "��G���{��tK<F��a��~��c�Z�<5����_2�"3+�EfI��ӬH"�_��8�n���������{`����_=�|�#�34ܣٶؙCڙ /A�R�Z�*�V��+X�zgb�d������a�Z���N��G���.F�y��
�<0v��@f:�O$Ϳ��A��I�m��F)tv\�,��s~��%��w����,��ŷ�ץ�Ei�%�����ѿu���WfR)_�/X) u ���"d�]'cI�:��N3:.���
�s��bS?fw����%���<'�����;���E�X���H0�w�T1��~���G��@�K_��Ѵ1���+��=�o�7��e�X��g�e�M�4_^�����q�Rm����<�俊��R��<��B���vO�j���	#�
0�W�	bTZ���g{��r�C-?�w�9�KI��cG��-���uΣ!cyv8I�* I�+�?nB��։�]M��L���aV ��G��eN8��:by��g��d8σ$1<x4�J�-�f���m�w� G1}�������-�e�M����2� ���K�c��*�ͳ;Ѱ\eQ��hp%th�8bp:�6��~I��Z�����Hp(�ۛ���u�$擊�~ԣ���u��"�Y�>�&���<��xq�hk E����U������y!��K�W[j�@h�8g?W�i<� wSD�� ���k�#Ϲ�ơ22RF�a5G /��ז�ZB�H���zt$܈�c����w��T?�P�VU-E�oă�!�bv��SA���?�
Qw
��-/GIG�c=�;���Oz�V�/,|ˣ�l*�ђ�项����F�0�Vd}����7j�H�\��3^r*\|gEӷG�}��n��ձ?PS#�O(oF��mwj	�gr��W�=Ng^�.�Lci����*t�=|ʞ�k�%)�4�a�h�Z�tGf�P��KҒ	��Y�n2"���J����-�lG2������1)�>t!�V��Jp4hk��/��	K�-����f�s�C-]�$d;����L	`Ε��>���Y>=�y|sl�c�7z��o<�犫�?�0�q�!]�n1��|v���
R�����8ZnP�9k
w }YmzsK 1T�nb�����x��%l�'�(B��Gn��d�uѮ�<�҅4^$�@�nчw�2ս�^�$��,'��������X�}aZe��l�/�L]O@��vF�L��rw��C�l�J�"�I�.��t��/|`FͶߔ:^UV0z�mC)�5w�4��6_�g��)w]@"%0�6�x�+�)��V�2ؘ�-d!��ؚJ�-��ηg�j�Í֋o�(#0��ǆ	\L�����	Ι���e��n]�o����,e�w8���L���.k&�fE?�7jk#C7K�V��I�8E���l�w<$ �V�	h|��{����2�=�ˣ�F�b��^�g�5h��O�������g(���i9`8�Ip%�{�x7��XՈV�S��p.k�чl2s�U-�q���JG�dJC�AR���,��#c!����J����c�Q|���P	�c�l��������O���-��I;N�)p�_�6U�ɱU��zC{�x	
K���������"V�� H�S�D��W�@q_Rz �6Z���%L�?�34��y;L�b"+3��7��9����{�s�{���._�/�������W�+~B^ߢ�h��m݃�6o�o�n�`t��ڑ<%w�����s�  M�yucf��p�n)�ޭ�W�{������G�_8c��-�7��e��oe9!\��B�-���H�Q�8����W�! ��n�l���3 E�DO�c�-�1�sC�b��b�i�C���1i�_���%�=ae`�T�=^���N��
�oj�1:-�a�'4�56����P� �/�K)��G�U��K����5F�l}5$�H�&����3
6�Z��X�q�na��C,��Oi�mED���N�f)�	+Ya��]�mF4�����f$3��h��lL��T[�J*�Z�\��ȩ�>�g���*Rz��J�`�0M���AN��Q�Ȕe@�����V/�f3���ľ�"y�M}�ESE�‒f�J�Y�t�Nd���:���H%B�:;s;\^�Ӈ淠�:q�j����ܐ��>+���"�P�h���d4��2��J{+_��۩�H,xn�����Sg�)N́�2ɇ�A6��1C2E��gD;	�\f�`��`3�
�)c�b	�>�څz��9��0j���~j?�/ʥ��Z���S�K/C�U��= 4��c�(�~@s��,Q@p>i�ċ���v���������[n���+�`|;����������R~��rev����2P+�{w�z$tM��!��LI�[�F��z���^�↕�m=5Gj�0�@�^@�!}�6q�
�mH\��WǸ�#��>&ܮ銵8KY�&��G�Y���������<��ƪY��x[�wo����MI͗vEm�L����Y-��C��I97�����h���츶�Ѯղ�3
����>��*�p�_�����9�,���C:��c#�mƶÇ�-i�P�v}m���R�_M�O�,lK[=�D��֣jU4г��@L�KŨ�?妸�T�G�r�!��S|D=�j��
���'�)��Йn���u+���F3���v�t�)��d�:o��p��<��o+5�,/ѥ�����j�t:e�9˅��h����/�
�8�7����W�ఊ�ؙ�[���w�59�#}lӗz���d��r�5����ץP��$<��D'���f:9bR7u��J
��n�F���j%�5��>�V`�^��O4>��Thw��wb�&��@�����]i&��^���I9�ʹ��JQ�pn�{MMl>��j�!��%V/]�w�I�QA/�!�^MF�Q���qq���,\e������U���"yE'^�f�ޑ~mc���y��\�`ŨP�kP����jK@�gGQ^qئ��$Z�J��MbN	�7����*�����8�8Go��>�H��ϝM��X	�ʊ�o�����Gω�=	��{RG� ��a����+�"�C.��f���*�<t~��c͗�ȏ)�[XF*����� u�M�I�����6�@s�s���X��Qp�`�bY���+:�6:�&=hϖ [k��'�`"�/��f��/����i|<��t��&�%��;���l�5O���zi紘Rҷ�����Gzf=4wL��j\k[�-����$ ��j۷���;6�;�.:�������W�m���k}��Ԟ��Io3�8�lS~P(m��f�nyRǹ���yhh�?�b3��\>�B��>o�441�'�;A89}e�'�ܤ�IL���z߁������)֊+�b�p��yu���N�]+��|�M5��ip�����>1=��,�pl��S:���\�٫�|�O�P㛧P��l��ד��cġ���L]3����W˝Rtnk��2����.U�$ep�2:@k�*mE7wzI"�g����"&��k�9�f�B� ��B��Ȍg�tE~��'Y��w w�h2?�%��]�펮��j:������0��2�=rRI[�����z�F��WPw$o���1d�Ş�Y���Y�aڽ�B���!�ֽ.�����犛�B�s�v$����g4�4v��夜�"����(�FU`
<�S��B�l�Y�z�����T̅V&ǎ�d�<>��������ur�Ж�Ie�@�ӯŝ)��dnG�9����v��y'��M'�F�^��bD��-d����
��[a`�)|�|�JM��0�S6pW���,�V���=k�I���q��������2�*l H���C��b?�vi�4�����c�74��C���p�����dr���V
Kڑ&�t�9qѳ�/,�K�E�&�L�ܥ�tG�Zۜy"Pm��q�,��h)]�R��W�����l�g4��ݲ��\��9z���;ݴ��nV����*�T�S�RbEDlN#P��G�#6N������2�.�+�����/�gӈ#m��P��E�O2gj=!��񈘶�(��Q3�^Y8�a��*�}2�p&�Z{��G��tu'�f��\��a�󞸚�T�~�yij�{_�1�X������Ԯ���ƞ�[�D��������>��ܿ-��v�P�.��7���P��l?ɭ�|#ؿ�� V6��$�Ś���o��H��#&�%޺�&�UۂT������e�o k�\�uF?-Dqdמ��2����fTbd�;�.@"=mJ-�j���0o��T�@]X�>�peW%��SS�3�	��͢ȉ ~�or���gdHk����z���ZȂ��ej��'/B<�\��_���'��J���\��1�=O��Ý,Q~
{%ST�J�N�D|�8������+�3ŭ� ([�S媥��u�O;+W�c��ɋ�+Ȧ<Y�n.�. �.�߳`�
9ry6E���j��YT��{ü�H�s>��+�`M�J&c�b�X����q�ة"GY�%-F�-#+e}d���!�T����z�r'ȡ�2OƬ��
1���}�B��-��f�V5I�����'�7=duf�r�ۡ��'oif�P�>�Tm���5��v�T&���U]m3`,̇�;o�K�(b�
�龰�:� ���������hp��<�4��+��!D��%@��N�P	�1f��i.�fPF9t��@"��2]b-n��������W-}ʺ��[%<\���<��G��0ܰ�{��"7���*��*��|~A����,�E�E6�	��}���'sF�T�"�;�ˌ�K��!�����[�iv%HG$y/D]�g�"q�ڡ���|_o��{P���,xxBRP�g_��	���$}BVdn��`��ˇ���2�>;�Y��4���2[��p�]yD�Ő<���7���r�0]V����F8z����oo�� ���Y���ؕ(����2����[7+�h*\�\J��(��T������j��u�'�N�ׁ��`Y�k���z��ޠ=<;yV��!R�-V�T�\�dMaȳC#����������0[j���Na �����ϟ����`K b�"0c͛��bd��u���
�A!��/�O���zPJŇ��
>Q���/�Y�?�YH����NG"�r1&�f=͐$ep+'	H���"%x��k�͡���4��9�����84��Q���[顣��|m#�~����UroG҂����D��|��,��T顅�B�:��ڐٗגh ̿�v�VȰ.t�}����<�A�!�����i�
�!k��>U'�����V|�k�x�����������ܢ"x{��@�`�}�W�u�7s�3 ���#��H$&�G���q����E������;O���O6ڶ�ߒ�����Z���?[1��R�m���_�A=Xn������5ܕA�S->�/�m�C�U�0�?��2�Z�2�1��f��n����;Ig85ar���+\Bo޵ ��O�(��������-��F�JQ�f7���2�K�VݹsL�72�Vp<�.Av`#~m��c�?�p����Ћ�@�iE5:Y6`:Go�[|E7ז�Ln�"� �r0�ݮ'<�|簥��ID��Zi7�:Lk�-K�s��[z9�����=��ACE��I�7��n�̈́�n$9�E.	�` �&�=I����P��׆ �@��H)ک���Cp�5��x���.!<X@yO���I�z��&heY\61�_v�4E�%�z�/ҠԫM*������ί�;���5	Ev��:	�s���q�owӔ�5�m�2�qBB?�#F�s�^bX-覾�TT3aq]�k�ʎ�Z2�G�"���C��`��� A�ĭ�����3�'�����>,M]57t�W��\B�V\�]�WR
�H�K?՝���[�*�^m�9%�p����㑅x�}JƗ��1�h����^Ar�EO[p��nR0k
���x-��=4-SL�V���H���O4{���z��\� ���7.��JP�K�+�;8��[���������h!uR�=9�W�K� ŊzJ���i%�,����"G�p�x�c������З���� N�M������B�ql "��hm����gcq������c�ix��=����W2�D�q�gViP�������N���.��E��[�`i+�aV�4R���̗�'�!c�#D�R�ulgJ��ޙ]�N�KM�.�*e)�񺣽Fv1^��d���o-���-Ud�Ⱦ�^�,�
I�Y�l��y+��P�$/$�|x�U�Z�z���)���/�[���ё�­�
��4���C'�?X ۲m�j_�}o��-'���u�?�L;��D�fvwlL pN)���K2��qd6o�,��������-g��)G4�(X����V#��L�C7����U��)P%�\���_(K��̈���3�?�ч+.v�Ų���Z�.S��U�ݢ����R��#���u�пX��	e�-*(�QU��$�WL����H��W*o�m�C�K"��C#�B���қu�^9ކ��|3< �&����k�H>\.��v�Z-�g�(��0�@1�^�x�(!�g��o�V��@��@ތ��ߴ#H�ku+�����
*S[ł���L/>�8�-)�����&p�;����-������a_J͞��G��ٝ�V�&Š�꧖�d�W�+W���WC����������Ĕ,��4�I����ک�����)�g��)Z�1,R}JS�;��%m���$c��p�\"�_"=6��3S��e`�.���<'��\�4�G�0�m:���]��
M����JD�2�c�!�
k7Гh�B���� �Q4��׃Z�Xz꼈W�2T@g� ����2Y��(?���u���~ڄ}�Q)�r����42��?�����Y��b��m';*Z&^Lg�S�I��z��HK�6l�M^|j�_\�� m&��D���:ԋp'����w����DNq^h����B@7Q�?|���ňS{��]���xm�q7K/��x�V9ڽ�;��;3vŤ��2%֜՟HlQw��$>i�#���G���J���O_��k��@���6�/��	$O%ڢ�3�,�=��c��=�\������<:QK�8���X,���4�:5��|ɚ5��-�Gys��b��k�#�/ԎIȩ�*��?�{�ݤ�*�qd+UnE�����B)���m��?���޹����v]��.�1{Yoֱd��$'��"����g�y-f�����ᾘ�>VA�eo�C�Ѷ��NJ�͚����3R�o	\����2Ko��@��bZ���t��T�S~NE8_v|�k�"D����cm��1�W��y?�:}d���O/Y��SҊ���DJ�h��ń��M�ܝ�=gMi"�z����������u���뻳k�S��0?y��㏷��T�T�TFѤ�|�K9���!4p�������\yl�s;�����'1�ϐ<�Ҷ�4�+?����K�(x'�Ǿ��mC3c'�z=Q!�:8kWj���G�l5�ER�������_b��J����֯Z?ȕs=烈/�[��s���u���k�p�ȣ`��E ��KHFí%yW��C�'/jt�S�D$�_��B���a�Z�w��Hf�L����Ks���\�"��Kfx6�I/ٛu� 9 �v�/�PH�i�.� 1h$n���k�*��%��gY��$զB76�9�G���*z�SI*����S[�D0�%�hR>A��<A�)=@ۼפ�Zk+.�ŝ�oPz���k����k����5}�rd~���x�\R�\B,�͘�#*�i��Iyn#|�P<s_�*M���5���!d�^����)?C��+hQ����_�/�_�O�i=������gd�8�:S������_V��&]W)�df7�'f�2.մVӲ�|�f�Z]�j���2t?��f7*�{@P��\�/� �t8����ψG6�/�F��<Roy�ZVt=R:Ƚ��9��4^H��G����q�*����|\�`ڤI����2|��ŇZb�zg��������{z�K�H_K޿�R5A�y��VsV�Tǝ��f9ToǬ���e��ro��1Sa�ٗ���Q��� '%M�.�b^�DΔ�����l�s'm�^r��9�ҺC���mQ�	��a�F��	�F�&?
ͬ�z<94���*
��Yh������2�ح�K�d`�(ْte�����%2�$Nk��)�H�WsƮ�$�&]1K�����I4^B!ŧcVoG�P
��NV�S�@�T�W͌�����V�����Ov�6����_���N���-q���~?>wt��[7⒲
����3=7��F��"��[-�7b}{G�����B�;�GpPj����:7�ɹ�I�:�ȉ�;~a_LU�B,.w����և���D;�OC��;�8$��t�rd��]�+�eZ�#��$s���ܦ�P�S�EDÈz�#��lY�?�Y�������U(�md���騘�P��X�yؼ�Ũ�h�w銥���%��@�6��$��/i��y��Q����1��]����j����T�}���x��לr���
({�A�f��3�L[�i~�G2k�TO�ؒ%��|�D?��ԭg�2�����^n#f�\:f� ۷(�}2v���\������)Y^3Ѕ<0���QwRS	~�GB�V��`� �r�֐׋���x�P���'r��ͺS�i<���z���6��-�^h� #X��g�,h!^��|k`���./�I�Zl����?��T��= ~�5=����xo��3�<�k�Fc�PEg�tvz�-�O�P@��:��d���� 1M�D�K �^�П�pn4_M�6���I]���W]OĽ~�v:��y�=��ׄi��j���k��xק�F:X�(խ��[��W�a��I�N�D�r��)H���V��Y�'f̾=���Q��w�*~����p��&�1k�$��Y�@{౧]tsg[���!Tw�z��V�/��RT3�ج �c�d�B���w."F��9����g����ܮ��u�7���~̒g�&X$'Y4(篥���ȶ�ٟ�����=��+�)�W'a�S����Ա<�J|���3���ջ���.u
XN<\/�.��vC���j����9�y,s��!���#Ky�U	����t�x^��:��O�%W!���]<���7!2)�����S��А��U��]�5C?s����6�F^�vi��[��*؅�r�{RT�_���E�TY�S�+�0/��U2�*m'Fg���?<�q}�l_�+]V�����A�lTT�RB[j� ��.��i��g��<��9���ҥ��j�,�_�����2����<#�(9�W,7�,r��f,�ל�p�M��W��0߉Z`G�~�!� �6���8J��2��j�\���3�IV��
#W�Fъa��8���G�fK��yg�O! GUX�|vأW��@l�	 ���`8M[����e-����RM�Qi$��-�y�2�}��]�{O�sf j���Y��^҂�S�+u�b����r�W�3z����?!�C����nĲ�&��ޅX�Qy�c�z��е�'�R�)%�	)w�ɕ��ɢ�H �mґ����%��H���X�%�I�&+�H�+Ȍ��@���<��R�C֯��+�렭�B����f ������_���G�;�$dtc���������KN�h��9�� %��c%��s��3�v���V����p �U��x~��2V�%���g8e��
���1x�Aw/�95�tEctƚV��褆w�2����b�W��m ���g[��i�c����?f�t_|)?��ą[��"srT�N4���'����r���
)E�z�_��kKw_��F�Hc�t<���V貧���1���_oU����t�%D�W�tެ�A0���f�\�x�?�Ȝ���I�)K��.���~/��'xf-�&V�;}#G���=�eE�f�ab,���H�B�(�0ի�\�vV��a��{�_��`�b�)ȇ!Y�1�~`DFڹ�<@v�q9j�:�V�!��Y�^�Li���^�[��A��<$��f}�y��l��
�,�)����q�-O��d��Q�>b��&*~��Z�L;�����:+�3��֔��ԝ�s��C2�,���;}~�x�'�H��2�r�&p>^�T�MO���/���3koտ�%pi�MMn ti�%<r���WM4oGX���Hd3����xDu��mo��Y����f��R牨���]R�Z��C���t�!>w��s��ż`T����J�-?c���
0uBzYے�w;���牚Z0h����sN*K��44��q1'�:v$mҏ-9Fa�O���j�}-G���� [�`�7�xU����۰z��RA���*����%�'��~��8��9�|��}w
p���h\�=��� �~ �K�ݗ;�`�v�n4�']u��{� �]!��.t��#km��@��3�����D�8\h��S�n�����}#��J�,Y:ࠡ\ԚI3g��vS���cJ�;�~w0K�e-���>M#���H�cƔP~e�6��~��	=Ǐ[o��	;��}\�W���u�����А�{2��E��dW�
Oӣ9�Hk%�УЂ���~�� ��δ��}.	�n��㛨2��YNc�	��>��h5�c�?���@�@?��6̗�@����mQrX�&8S6&Iz�>�w5�����z^.��&�R��y��!/2��a���t�S�W`���)@� ���9�X�kg�������nd{�=П���1'� �SZ�v71у��tA�!��v�M'�'�=������E)��k�BP;kiܱ��\[֫�g"��T�^o+����/A���X�Wx��gog�w��s�W��Mf�>��{·�In���Bi�!y����\�>�!�޸4P�ɺvm
������ڵ9^D�޲�d~Qo�h�Oa��B�+��5d�FQ/��Ѩli��tp$#=�Rw޶{N�]��؞�v��}=)y?�����2Ͻ�M�KF���}���MF#��Ȩ��Lu@(��țY&�̬$Z�(g2���HUW?��汒�:T�n�˙	7��Ԕ��b�(cb:�g&C�w��.�C軱�Wå��+,I��ۛ
p��zk���GөOj�H�_���6�#�I�&E��c��)"���1<����4��O� V�֪&"��Y��<��i����Jͬ07�����h�j�&"�#����jK���>^�Ĩܐ���s <�4VJ�&�6���t/L� �������s������Em��"l�)��9�������w�q��T���-�.z�R�i%Š�C��燧v����K�"��b�S������P3��E.vQ�}z~^<�9�Y҄���Fb�*�^)��ۈV�� ���d����]��1P\<$���
�7�y_�*d.8�0�e��D7��j����4�"4�8��4ؚ�~U�q(+�����j�ѥ������=oG�h(���z����<�K��5Am��zs�׎ 1����'���\�ܤ^�^��J�����^��^T;�&�\,�
:�\ -��ɂ_�������g���M�]�6��簲5�h�U�b�
�z|�E�k��,! �"0��m��W*�����\N_����Ë��L�%.�<b�����WIP`�Y5���'�F&Wn"��s�k�w�Ȃ���f�ZE�g�/����~zЧ�v����f̮�W�3JG^�����u���8�?���J�0��tQL�IQ����P�>��r���=�;wz�=�u��3�!���` j{�W��v.�t헨�����bf�$�%/N��.Y�B�He�Lo�M��%z=Y1j�Q�8m*C��>���:D@y~��яZy�c��dXuh�g'h��)hv���S��LH���P��K;6�G�k��)h�Է��q@�z<$j�<�&p�	Z�{{�e��"0��M��»g��*g��>�3���|�
]�B ��GzD��pM�%t$tx���]Z�T��r��.��MS&���ɻ�դ��ֻ�ڐ�luw5���%�;pH����k*H�L(^.�č�=6�F-;�v���e�F���ZB�l�:��(m�:\Xz�s�V�q�����p܇��9� ���ި��an���p�6�W=%�N9��e7Y�y���*7�z,,�:�d�ZTZ�V"�1�������#����V��v�%{T����Ԏ��� ^'�Z6��ׂ�	�m1;��ߟT���tEb'�������s��3?�K�	���kw�
+id��A��� 5�u�F���0(IUI:��@��o/���Ĳ��z�k��S^ r_����`����З���߸g�ʹ��L ��wS_[�]nJ��Uh����a�Q'��Ǚ���2�뵕ؼZ���Z��$���.���o}^L��j�A#��)���v`y8"1�LH�5�>/�:`����%�r
� /,N�&�\����j�K����gI\�b����	;5�xv�OǭGC��a��z��m�tjo���7���Ͼ�./1��9'yLT�W�jc�0`Oۛ\	</���Wv �@��8�����F��	�>�d?|�Q��5!)g�����Kw�/�>���|�L��J0O�  �FH����3>M�H��u�������<%�h��#��Ý��$���ܸ��$��EL��Y�;8wa�C�/!^�����O(Oxo/9���N)���N$&g8��]m.�mY,&���e���{�BL@��q�}|hRe]>�rC��͜��З��5�	�wFČ� �0 v����\�_F0g���l�%�E��F�L-�~vn� �Ex%����{� ��̆�K�۹���5ou�~����r���L�?*��rH�0������Ψ��'Q�~�0��3��.��%��*������i�4Й�&jPK�sB]6��p�P�����o�����A`Q ������B�=U}ь������}���W�O��۾�%�o)��E�@���nj۩n��Cj7�R�s&�����f�W��~R�g��T�|E�v~�'���\�7kÉ��[� 7Ȼ5�J���8�D��Km>���Si�NJ]~�_�@���`fO��A'�M���.KN���Qe�*i:ܮ�^C��g�j(��O?�*�Wk�f����AgM��Ln,4NM�9XKh��I$$|0*����(�rm�������qa�����|����E�M-8d��������9�����	���=7����_���&L����9����D���X��	;��*�%��=k$�$��8ő`.���1��ǋ�'BL|&�Qm��X6��Y�������}.PX���fx4KV���?���¶٠}vH����gߘ���K�6΄W� ��������r��gձ�m���m�~��܄v�Cb�ֶ޹����M��ڶE@��2�H�hde����U}�|XD`2]�^
���\��Њ�����A��ՀM���#�E�)x�q�&!~�g�tO�Ӊ���,-�4�m�u�A�E�b�<M@��l���x�=/�
QO_��I�Yi���L0@��0Qy�%2���rk�C�k}j&�8%�p^r��pD�1p��P�31yE8�	��ߔ>3fذ!Z^�4�d�b��4��;X�F8c��
�{s\A��e��S�b!TJG�)vŽ ���9� R��#i6�JtxF2�� *7�	E�X�N��<ٔk�r�h?����r�k~H�J$7F�Ʊ�%��!���70��V�-�:�=PoMϿ�S>�����sJbJp�� :�G甭�y����,q^�WG�����}�K1{Ђ���(y��=�Jo��?K�0�ߩ��L��]�q,-^f{������>�S��:�M��޾gw&��CNl��������k
�����}�W��t�J#�Rr��������G�gI� �ǝ ] ;(����\ ��X��=/@vp��&0WC��bil>u�Ӳ��+�4�e��YY�+�06�a	����m�֩N����J���0�박C���_�9��CS^r����/��D�t^��������g�F��(��F���G�9��j��Q�P/�hO���l��ɯ�')��'�M����4�/g&���k@���0C��V~�y�F$Ja��fEǎ�9v�g��$̧eԶ��ʘ �T~�.z	YWW�B�6�=zd�(�M�݁�������<���g婈)t��2&x*�I����/"u���.Ը�B���{�['�a&� �X`��aN��WP|�R���W˘��*��Of��"Q)�89F�E�{�j��[����'�{?��ӟ��w���}��녝T�Zf_UꧢK����P�5SU�ND'e�Ky�Ǒ�{K��!w=- ��+\':_ugj.�y��G�uط���S��A��� ��yM`�<�h��ϐ��D,BD���h��$���h;0���J�Q�Z�����ޫ����\��ޖ�k�X����|�@$��O>�ki�Cn.��4�o��E��*�2�O�/�a��K��:^�]��=W����L��</�Y3���劬Tg�L�J�*�AK���>N��J�{���v3�d{�x�iB2��F������V�6�_��%:1�\���O�bzuD��/}�6�Uˮ�� �z���5����xv��F�y	6� 7����*�(A�9�/��W��aҁ}EF����"�!���Eodݟ��/�а ��_�#pW�j[�	�[<�t�ԋ��+���?b3�2�ă<$͸.�ZɧM���,�q�$�3~mC)�m��l�_&^�����܂�:�@;��-6�o�a�VHa_J�_G�)b�_�T�� �ȥ'­�Q~!#�Z$�A�@.�kua/k��Z�jH ����]5�$�LL9Km�Ni�*�8�ٙΗ��	����|�2S=�hH��Y���aCy��>z=jz`ҮM��kW�W�X�sX^�u�|? �3�������Va���t,qj��OF\�O�;�����L!�I�c�9t�NND�B�(�pxCgjw�}3�Ju:��tp��B\'������r���$˙���~�H�����Iu�i��o��nd���xi�W�1>b�a�`�lA^�>y��4D���Z�ܘbS����.L�a���s�����k�N&.� ��1mr��K �������*�݃��9�U ���Q�f�8O-�
6E�-��Y&�ƌ9@B׮���h����)!XbQ-�v0���[���zU���h�/�ߝuzʬ&V�峗\�irJ*ա�JB���{��ԏ��!̃����.�f|������˒C"H��	��J� {��F��_���U�و��Re�>x����|#�D*N[U%�̳���[ �\��G_�%y �x,!#]�
��tU���=��D�FξΏ���3�N�ex#�q��|fz��!z��U�2���uH�&pRd����.~qL�
�r/�:\z��[�˪v0���XTO���5E4�r�6�\�Hl
�
�BI���d����ˊ]o�ͣr��y�W�!�>�)�B�Mc�Ώo�Nz� e]��eO�L��*U��|*f�h�����$����0�&�o#;�t_֢[�a%����D�Nl�%����c^
BI0�3��A(.�፟�׻,.U���Oh��v��8g\?N�ܕ��}���pEHa���AX6�,4�Ͽ*[v�*P����[�<���(�m}>ŶtZ�+��6m�\B!�)+��M̱nm`Z��d��=?���R����tD<e�Okڮ*9] ��r]��L��C֜�{f�E�܌��GXS�t�6�Wj}�i���#��H��K3���+��csu�af��,�����t?$�۫����E$�9P�5�djވDUH3���3�Nam�������m�N7�dk\~r*��2I���ȝF��;�l��>`��������5M��ֶ�����\�'F���]/���_�d�8Yﰥ���!��-���~�S���I���^j�]� ju��u8��g�ƫ��	��UM��X��2��R';1	�.�D�H�z���hF(^��A*�e�����$���8�X6���bT���k +u��
�Ӟ�ė	c��␞�~���ѸJe�|o�is	夊k�$�P�Q宿��T����c�O�:
�r�_�q4�dl�m�c�ޞQu��Tr���ʘ�K	S��W<4���ʶ�Ϧ9ɂ���K�Bi���u�܋����e��B���������������h�濄�_D�k,�����Y2y���C)xUv�ݾWa�iy��(��{�u��+� !��9RxJ�����j����-;O1	����g�M�ڒ���&LRC����>A�:����,&�����7h����מ�(���e4��Q�#o�_�&lPY�rłXJ!<08�XA�������6ڟU�ACTI����F��2x��K�������\��';9uwUEk��5L�N��U�,4�M�U/�:�6�����'�gi���0���1��z删d��j_���ީ[A��v������-�{����z�T̂��x��l��Qg�P����~+�Y�rZ�4�7i�I�PG6&=��t՛8��ݭ���[s7Jo��b1a2ά�}��� b����6}����L2g�$Kh�X-��J� ;*J�؉�뻑U�'�-����Y��G��*�C�n`Ȩa� lp��.&d1�������^S�8�7�gv�b��`΃���gA��p��I�y� ��J���b���?`%��ȕ�c�3�<6G��]�߄MW՘��Z�o�e�����6c���kc��6�E&͇M����O8{z��sY&TC��b-M�J �L�sşT� ������Z�c��wՎǂ�G�Q$�qU�����0�q��x�QB��qFE�@�po���ϖ�,-�m�v�v�PA������������OM�Tu������1Q���BA��a�%F���N��n�o���Y�Cv�%5=���!6�@�5^r�{�`DsI��7�����up?���4��0ǫ�l��&�c[A@DRjŮ����8��7	�����2\��>�k[���Y��w&t��+:�\�C�t���΢��.z���y��S�g@u���7ܐ��2��o�{��A�[����n�ZHXm������
@������=��C3dH c�S��/s�|
ni�X���o}f��09��؝�+yA���E2Cv�  �E����w!��p�_��R���t�C9�p��MF�gjԓ��dg�w��X�?�@h!�ț�KV��Ѧzfr%��I��V�Q�reD�.[�I5�G�9�g�%�=I�%p�:�����ƙ��E�L��Rݺ*ޫ�'��b�ގ�\�9�]���~�V���4�w�mq'���D�t5�dk�xu�N��&"��e�rV�>��ZD��p|s~YmwH���9�?��!%4�����Xl�dV86�|����7��N��T�'~�-���([)}�H������ԉ��������'9�H�m[�2C�:��	�jΐ��á R&��띎ğ�`rwD���jY�K8�N�����#��g0Z'�������+��W���I�����(�n@a�ݲ�a���������+KI?MP���$R��=�s2�j]�:�+��q'��v�xB���-���w:r�w!���O��w�H�f[���}�H����;�X�~A�ث��0� �&�FW��⊬��Hl��<4'm$-�qA&�ڦ�	Eg�[��q�B�� uYM�����#�����p����K�=�9 *����V^�i�srE���--3!�,���J I�l��HƨOA�{��ߕ�S��] zZ꿘XU���Ɏ�n�IJՀ<O/i�ϟ�G����3-H�k�����=N\�!��MS��32���>;ؼ{�/��h%��َ + ">��:��LۑW�%����˝�XkZ�լt�$�_�r���܇��v�f��9^�r�ԭ'�Xg`��g�[3�M8U��q�~�u_�u;>me������e�PC��E]"��Uma�@t�>�Jr����(����a^�o���v#R��&������ݛ����R��a_XĲ���ӟ`/�.&�뽾��H9���o���1
�c�I��.�Ғ�CHټ@'M��i���W��D��ٝ뇿>��nQ	���A���(U�m\��
�'b�Z�satm�H~'+��jV�gy����g�8@�);i�g��ßp~�{X�ɤFMg��:MA�f�� ØD��ƔҶ�+��./2��*� ������z'�P]�k����o�xY��������;� !�c�{5���)�
��{�����[�l���LE-�U˞�*��#g���V���@j<��/�i�-�����997(�s(�ᬄf��q]&�-	3�����nE]#F� Qz-��D�K�[�r�K�#�<��%@k[؝�
WGtk�Bk%����K����#w��֦��qH��s΁�黣^��y$:�n<����a�T9�>�Mx^��+����&s�M�����(p�4��}�Fm��%��tf��UDz����!���vfؤ�a����\1˵N��u��j��e̖��eS�M�U}�/7��4j:�GgE�}T�y���5Vr$ܥTc&\l�5���޴�п�F���!��G:Y+��!��e�L�� ~�h�wz����W�v(,�� ��ɣÎ�r��^v�a�����X�'�.Q��2GWv$�~�q�:�f�ϯ�+�'��b�m�T�C�^ȖX^�+<^�A!ڿ��E<D��<J'y��K��>�(\���e�����ϩ&'��d��^8�g�Gr��pӓ��zI�&�@P�0�<ٮ�V"�E6����*M�jP��_65ό�ZT
 L�)������2��:����Dߋw�E�(/t��-�͒p �C�6%$��u�	��W�v��G_��3"R�P�'�
�<�0>K���m��X�2��$aB�cU H��!VJNĶs�{yaM��~�66���@�Rd=�f�Z�=�$����s-��?���*1�Px����-�@�
����5c�W(sc_��;=l�i<���P��=v֞�q��s�9tf$�\�9�����^��6>]�����^=qF�an�[��\��V� �����u߀.���5��ys̡O:M�t>��~7�:6P�Ԙ��S[�G�r)9��� ��=����݇��5�CBBJWg~�K��*�c����:�,�ۆG�-mr��A,I>�!�X�u��� �t�-�ɦ$_23'�^YP���d �k��P򙭾k.�9�f��H��r��`x�ݜIR( �1�������K�q�ݘ�X!�x�Va���#�}l@8����$�Jv2Ub�?S�|���a�}�����*�b��1��T�@���#������#��?ŷ~_cx�`��AӾU�H��A����IdqɆ؋ج��,�_2Ք��E����B<��z��6V��:_N�w}vs�}MO��È
��1d;C����H����¢��j��r��ǿ�/�ɮN��a@�������ſ�y,EH1	�/����aWų%��T_C���f�or�Ǔzi��{�<	'3_��D�y�����I'i�p�$⋱�ъ3_�\2c֫j1_WҢ��6�}��:V���S����A�w	�^�"A��İNU�ì�/&2Z1�����(}Ü-���Ȍb���?�h4��(�����Ajk��R�j�m�Xz3�� �d�j�V��]����G���0
����/5�����B"��d��|��Trb�t`0K"Q�j���q �T�qy�x��4�	���JJ�00֍��{�;+Ur�[M�go\{��\� i�rBչ��{��h�?�;��w?����k@�����2X�\M����:j~��E�9�u�#��)k��PaU�6k���t9�?y�>��:b�`�0��y�sd�������)[��B  �ҡ�;��_>-H�<D����]��	^�lh�+�5���BhV0.[�:�$��,�4H˪u�K�q[)�N/c	�k�rd��9|VF��˴�oF�qѥ��ƍ>�:�xl1���긡��A�Ep}��7@j܏�����b���%�)ݎ���S缿��:��ƕ��J�õ����N��)��.`�y|a�
�#@\=����9���u���AV�(򑯎�L�����02��a?��X�������	�_�?�]_T��h�o�[�:�6��6l����t�徹�ȪR��k^(�̏�>��e�	p�ϽH�:P[,�����G��؎�Vp��}"1ŕ5�J~�>�4�;����ڮ�ym��9�5�bX�RH|:u��>�k�Sܙ�����,����U�Q���'@K�,���A��2�D:�@߹w�nk9��N�� R���J�M�.U4vb��bF��2�r�?D  l��"�N��� ٨`����k�2�R�i
ҽI�_��*_��QgAڏ6T00���if�w��Է���v�3r]�AU!�y���ҕ�+��Ǽ浜nv)��^��=�[�ĳP��|��-�ؾ�S��o7_��3&���.�FK�s'��^58�禫g�>���ޝij�)�]�l�y�/�dg<_�P*���<��n��Q�lW �'���M�\ꏣ����<�{=A������%٢kf����\)Xr`��`�������hϫ�1!PŸ�2Ҟ����3٪a����U�OF26����}�b'e���7b��x��ԅJ�e5�3�d�{�f�f��;B
n��-��Zp_P��Ķ��6�V'ee��4���R��i>
��h;EŚ�a^*=t]0J���9��?�:��ދȕ!,\�A9kiG�o4r�^/���j�v}1���;��E�"�֮�A,b����X&ر�%9�`��]�I�7^�{"2p*�>��G�w�`��;=.�΂yf�E@T�#��I=ԙ��-�
S�)3e.Ԇ�{;�כP�i*4�| <��3S#��}�۹aFZO�,�7\�T~vˡ;\*8����
���B����Wu;�(TB�Ͳf�AM'��.!�uz��h��R���v�y�[	�, �X�0elgf˟8���-�\W��:v�C��ѽ���ݕ�"���"�v���0UD6�8֊�