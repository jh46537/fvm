��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0�����
����'a���en�,�=y��~{��i�#�sS�Z�àx�WW�Bg������𓇴r�b�ex�Wv�c���V[�4+9o]��\�S�������_���]U��J��]2c���L��<e�@�&���jX�3r|~�SrOa�{NR^����y�R�ΏD�|����m�'�m@�q��S��Ƣ,(�jݎ�4��>X���w�j2�)M��&�wU�=�a�;�k����K���b���ʎ�\������E�\��,D�`�������A\]��J�o�A�����^�.�c�mC5�h�9����N�
�.�C�!�V ˘�٬.#�]�	ޔ.�⏩� j4pTMt��U�uW#�����3��ɐAw����/5���C�اDt�����e���#�h�e�W��QyG	��,ct��{6k-���w�Y&=pK]kS�g7�̝WJ� �
�Y�X�K���L �n��ӡoQU�Iy���r���o2k�aYDx���v~WX������+��xe|F\u�R��0?ked�1G���U��'i��Q8{���=X��c�H����Մ�t>�����T(��k�C���G5�,ɜ���Y�f�qS���X� �f (B:�	Ce�lyB���n�)��Αi���j�c�A_>y�U�s�, T��	C0�4�108��(e�21��&�(�!+L��P�������]]$WI�!m��F`�@�u�9��J������0�p2/���6,-�.�3���Ib�Œ�0�l��^S�������%��a�\ ۘ� "R"l�� y_Đ���KR��u��.�����7��35e��rש3�V�e�B��=j���j䥠�E[�`2�fK�t�����+{��N$,� �d^x�ȅ<��{	��7�{�`��Ʌ�i��zTG��?���E���u�	g�_��"u7\w��DwYƭ�/�-�KF�?ַ�	WI���`��Y�z�k׮�)���2����x�R���C0��M�f3��t�"F�����qu�U�md*&Tx�M��d�k}�A�u>F��X��c!��66����C��[vKI�kFL1KSD�#a,Rm#�;� o��6�)���������iN[>�DZ�1khc0ձ��
�USٺ5��!E��&�01	{8�_���p�1��{_�ju7~s���\��H���e��ϱ��P�y[tb^��Dޣ��q��	�$�v�#��+�����������~��Vkc}N&�5�H�Ѿ� �����׋W���o�_�;����MA����S�jѨ*w�ͧ�;��O���� ��}�����)��  �#
�ن��d9��@�>��0:������?��4��Έ�t������}�z��zdOEM���߳G3E�����2�|�Y
7� �O��%��v�A����g��S[�������S 7�veA��� zS��w���J�P�Jq���������*\&A2h�{O�Uѳ==e��]c�u���@"Gʎ[ګ�_ 隘��� P&Œ�O�E�Y�v��L���!>,�%$OT�u�d�g�-�{�L�\�Z� n��~-$�l��	@���r�#5��:1F�.|��nB/�Þ���oM�>��O�Ƣ��N�ڭ
���ǒ�.h����]��?��r<���\#����6�+�_�X��� �ݺn� HBve0�(H��'�>�y��̈́�VS�Ո+,��R1V�|�њ�'0�L�Lb��,2�bLЈ�Hj���1��4�Ԇ�Q�өo���Նl��U�&�]�z2*��b�4O_5�g�Q�9��)[M���)]���:���2���+)�k�E����sA	��뿒�p����}��:����ned�i_��!Ȝ�ދ ;	�^��3���-�X`��H��mE`�I_h�88gOLWF� ���W3v)'��%� TfO&��k׮��٢dP���~	��y5���l�@���0v�AUp?Dl����šmјݴ�f���up�l�X���_�^1Z�㌏�T0Bʱ�_cL��'��C�ƌ��X;��Ϟ�������*MIs��磛j��Z���}���̰���8W�J��x������kK}td_'�������oN�B�Ӗ�M�3�(?E� D})0gu�LS��Rf*���t����c]DS�@B��Xd�.;��G�1`�y���Z���2�h%������$I古���o@ �]ƴ��/�
z.e�8%��ۡ�U�/�w����N�ۢ�����X~����$�Hi	Yzn����?��b�^	*=w[����@�q��L�N:=Q����_pU�j��h���q�i%D�O�B�K���)����ܚ��Z��	���!���U�*ʺe����L�U;�����%k��2�ȖV�+Z�����h��i��K�>�:޳d<Z��d�^�毶��Y��a��@�[c�I:�13[��>4y��(�B�.���u��l�X5iFNQ{�Z�^2E!]�FyT�>D��[ ���֚W���0v���Ri�&�Q�j�2�<�Z�BV�\{��|��L� �����0�Ym\�OVY�׀ٳ񸲦-��nzTBρ&���rp;��̷��罔�(p��6��8�\հ�?DJnU,M	+��v�yKQ�`�g뾼�F�Z@�v>��|~!p��o�OuZ�!��/[7����oA�@��c��K�Ⱥ�D�g�G������>���101/��j~��(�ϡAA�	HG�5��+�t02����xI�\�|K�G�L��Y��ނ}�H�J$�\)�����Ym�,�%�vĩ�'��6���Qw�w��1�b8\�}8�����mB�����|��t�i��ܘ���+Q��Z���p�G=D[��*����|~�]=���������p��·h��x_�;��N�����i%{7x����b
gC'���V�W�=��/��6����S����ɇ�|�O�2�͍y/BLQ�E�1���A�(vRY�G�E��As�ɑ�F=�V��#�e�o����)�j���ǯ���̎�T���w@��&��d�&^���i�"��ͺN�'��� ��� 3�BRd�QU�r��軽C��w��vv;�l⬈2��mA�'F�T�����<�Is{�] �#�+$c�{h�f��y�a�݋��z
/ζ!,���<4L� �z��&���>u�l�>�b����=���ɾц?@���������f���A��������p����fXe;č���3zU���X��-�w:1��[_�CRL��!c���&W�w���I���^g5�)&4Ot�x6���1�&��N�^�A�FJ���]����9k���4UQ���Lj�Ʈȝ4>é��m#�=�}�y
WJ]%H��J���L�i�Is}�_4�˪��GW�)�%K���_pQ����yG����K�mj ���}{��>F�`-�QT��>~�l��i��1�u���}TF�T�W�O�Y�ڒ?�1Nχ��>������$KR�dF��19����}]{$5���'ba[,��a&+��f1 k��(qT���]tޱ!��0�1�0j)"2e�� �oqf��|�����C2�B�"(%(^�(g��hx���Z���q��쑊�P'�i\�R���g�� a2�A]�J��]5����&���ƍ:3�BJ(�Y��v�$�mۦ�IU������۰����L�1"*%d�פZnX H(jN���Fs;�o����c��k*}�pR��^ �������sQ扣�=z��:B�qi�`IFz�;Hn�8^�+�����f��zل�ĉU6��e��5����=�,��x^&��؟,ظ���`���X���rI�֢��<E��\D�9v?#�l�n���$ ��K��dY�	��NAOkY������ۖ��.�h�ѝn{7�V�����߇�\r#z	�o�������WF���b6� ��E֒b��2�GG,�5���물��+��.f�lU�_.O2��L�#�o�����qFȼ{����8D��"P�0��X�C��V@FM�+ �:��8��^w��ף�Pd=�ݲg�ߍy�o�$P5�Z4�T�{:9�}���>�8S	�}�F˜�ar�E2I|jA,z]yU'ɕ�sq�V����X�$^��VXT���ou>pU@����ҽ��FjǏv(���m���H�aJZ�Q�#d�p����n�x*`���FqF�G��٠�p���5@�R��p���FkB�JE��GgC��6R1l�'i�TMٳ�W���PG'�Չlu�C��O/���2�P�F�*�������VZ�e�t�^	gڐ�z��o��,�w�Ѓ
VW��)������U\_ݨrCY��#��`�.D|g���^�QslT��{H��!7����K!B֔