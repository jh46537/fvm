��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[������0\8�J_R8�C�{B�z��I{iE9�Ъ�+�x	�t�w���V�-L�Ȑ�ۊ�ʭ_�(	��9auo���O������Z-������v���$S���8,��	Y���f�t�d�.�Pu����L�!�c�M?-���	kX��5�n��o����|ӺR�v�-y,��Y2�Uk+�3��d;�ZM��U�c�����ԨWr�ͤ���	����/�L��#|Rhr��(FD�>�,����I�B ;/v�y���;�0�J��qAǝ���!Փt��p �4��:
��Xj�gB�`�k9�޻�|�>�?�Ţ�r%�\�(�����Lc��L��q0о�Z�{���T��oa�Y��?�o����,V�n�1��*��Ў$?1`�ä�OBq��p޹oB(`���~Mc�������y{�/v@`�pIx���t!��o�Q��eƵ��M
��v��ʞ����`�ć�ǵ(���)�A&�\Vn/��~a�ek�^��"�RL�@���#GI��[/U(���?�S��50!�3�#���d���؃���E�	j��!�=oHn����w6)ĩ�3��iUj����e���MG�O d �����`��5�溰�uO���`����-����xPt9åx�D��t��<o�m�c� ��I�����X�W��b̙7�Z�F�3Fߓe��ߋ����&ez�W�4Br4d��R:�x�b�lr;C���-8s��'$����E�b�Դ�ִr�0)q�G2�y
4�њ�9�d�?�y�5��{�>������Y�냲��O���
�$*�㻛��"��#i����>Ú�����G��,���C���s�Q��0��� ��-g@���"d���X�����>kȏY����ʏ��k1�.�h���d>^����4T�,��p�rgaL|����{���ZN�l���%��0LE��iZ�sK8�� ��^oz�[c���ύ�U���8?�y��Ԅ΀8��e!��W�.�m�c�ӲQp[mijy�T�~��^��T�p�hB^ON����*$|��X+��텖3L�pցI8{��
*ڰ�G�f���/��g���i��dX^+&j�u��Kp���su���m>�l�kt��`��S�O�9�TMf��`�E��hx�= �W�L������g�����|��0���Q���M�����댭��zH��;&�_fC� F9�P�̃%�Mc甓�����@zd�CF���Qؠ���H!T 0��k)�����D�&�U+۹����  G����Y�9�`�2�:���Bkˏ�"�Hi� �{��Nu:�S���i%pu�mZ\�	�L;��>�{�[{���?� n7�4D3��#�"v@#����bx�	��(�)�9˞}�#��HE�/�  C�ei�����c��-��D/!�#������aO-�h]Z,�
���|�TH1���O��7G����'�M��7(ႩI��H�?�a�N/Q��U�a:b| ��#�k9L���Ҳ{U0'bp+O.�\�ht8?iuk��PP;	x�&6����*&Ȝ��gC�B���&E����9t=V�Z�����{x���I�%  1�4 �A�_�%�Ǣ�ܫ��q�!V��w�Y�.bt��K�br��N�7��=T�B	����_��LJ�7���m[��o���b�b��JG��O5���˵+7T0:ᬀ�֌�^�	�* E Lp�4�,0����ۥ���訁��>�>;���fDW��rΊ���"���z�D� ��*��[t��i�0ǔ��!����SR)�4qR4H�������bwvp3m����Y�INp	�M��T�R���T�I�k�5l����J�2͖�����*Й��c8���寞�l����O�z\H�#䙬��?ʿXwۢ�����Ꜳ��H��:�T�-� "�@}Q���x��+tJ~�`<�c9�9�Шn��C`3�9sZ��r��8DރE�'�t����4N�ň�~R������i^=6��I�����#��.jv5	�5Ϟ+À�N��v-�PhW�M�R��1̂��ò������FE�ʥ�=t]-�qv4��+<�HRd;�폞*���0LhE{�HVh�L\�8�A��pB(��|�i�o�AB�N1b�	�#`��}�֥W���S�2��6j�D���HsGV�j��ɀ(�X���f\�5,
����Ds�,���b>�cӚ�+��C]�UԒ\g�zj��@hO�%�s?wr�[�̏�a�?��-)E��Cl�Q�!+-���eyX�T֌���i���i*�T]�n%�#��O�i������q��Ч"x%��^��Q5�ᙡ�	J�<��eo���
�K=f�BA�E@6�K�v���9��z"�೼t�����a�B�oܩ��	q�#�K]���愐�W��)?��ׅh�?ǁ/s�7|+g�_'�=��yk�P���,��H���m���4cϖ�.�Fr`��\+0�C3rt��</������O��	�Y�f股l�-��V�O���׈:��UI�F4�Kƅ�u��b�s������0���#���y+�g�kS��FZ-�7��3�Ά�W(ȇ~wg��.XO����(�g��!y�1�WHe��d�i�ZBw��k9{i�g���4.��U�X������*8Jk���ҿSfٲ�}�5Y���~42���O��������@M���JT��3D�촉eϢrh2ȁs������`Pp��.�d�%�M��+<æj�i.�Ft�/����V���{���X�Y f��ͤM�I��ǔ��y�i̟�����+!���P�ܓIlwA?
4���+ֵ��b8͋I;��6�)A�I"��:�4LoC�� @$��g�a��0��1�$�W�R�d_LV��J<�n�'�i����9��6��V�Wo'(B&?B*�Bin7=�����U�R�� Hy�������<�*9������.4s�%���#đQdX�c�%���
/gƷ�'#���P�`����I�����$�}9�r`4&�&]��'����8,ibF�	�]!U��"\dq˜��xgM�Xc����z���@� �+��{d��5L�Dxu5����Ȯ=�c�_n���rk�S*��A�)X��/�_�!��;��s���<���B�w�B��D.c=���'��ǡ�p�z|we���f�����P��z�����QG���81M��7���I׎a-��ₑΆ�S�a+�,f���%z���:�mO��q9����P*�����gʘ��1���h��S���Rl���#�C�ae|˴��{�k�������X�ů9�����e.��n�/s-/AS��o�\�"�ɕ�i8��l0o�>�~o��k��%]ғu�G [IVL�n����33ճ���t����	ݥG��Z���(�"<[�����<�#W�aT��+��H�7����"��hL:V���������s��l{J�����i'8�T��Ρ��;~�ǯ;����c�?ɐ�'y%n1�|0����)q�GIU-S��/&�\W��7RQ���,Bnd�6s �dN��4�33hlRQ����(J�����"���w+�F}hS`���[ab�.��1��UmlW�Ġn�rI~��V�+�	QW\��뱾V��U��BM ��x.��m�HߴU�����m��ZS�A��ilC'����^C=�+^+�䱊��3�>!�23��ǄR���ژ9���Zj	RDL��D�U�n�B��Q�
����TƉ����#0@E����EW�6���Elm�)&�'qov�L0&Ҭ�]˚j�8�~r�ԛ��xE�+��N�q������H��)�&y��P��`l�&&�9�\��*���;j���
\=C`���^%4�l"i�	?Mt�~�v�Ѳ.�r>�v���$q΍ݍ��-~�Y$Вrld���y�鑆@���M�d ��FT �+��.��@q�	��"��qGh[�F@g�Ժ�M���g.}ڀ`�O%Hs$�R>�A�c7L�ʔi�d�~��r{^`�y+ҁ�<�p��W�"�,�5k��Վ�Z��uu�g����茷����K����<����,Ԍ��]�(�V5�1A'�V���w4�_=�F��տ˄���-TF�<�.���o�F���m��r��C"#��� ��\������k�v�\t��߀O0j�=V��l>f{�Q˿Y�S��� h��P�Jp�/f�)��Df񜖣�t��Fՙ�7�3R�ؖtށq�~um�;hd��Y����֢�;�]D��԰��4cf�e]�+⾔��}/U�#m��MX�s�Zj�0\ly�b� �^g�L�"b@j��қWL�'��<�O��~n���u ��4%�O�����0��ӎ<]���~[@��N�A+�L�"�S w���K�b{� ��u�O�������o*�bJ۝|y�o�G
@����+�5)�'I�:�&Τ�w6״{�B�3�CW��<�}"cu�dQ����,�tU2y�3�{D��e����	�G�J�0�D��^*�B��j�q�pI�Fi�%����R�����qO�`Av�!��1(]X	��jr�I�4m�ч�o���KMt4.^~���ԠI�`�c����;X���ƛ���*b�Z�%��ߐ4��N�s�/Vs�1Rۃzr��Ҟ�a��+Pώ"���S��.*��&2{�G>���c�WP �|;N|���5�x����1��w���
��y}u��Y6����BI����U���P�B��ɬ����< �|4�F�X4�i�%����]Y���� B�`A[�m½���%~�&��gJ�����H!N����D�j'�5���J�)��S�G#�Pӄ���vS�V�n� ͊x�Iv�w0v�M\����q��7�����o�V�Q[}�K�x�̈�j�+����IP�%�d;7�PQRs_�1 ň��Ec��3�L���bQu/a榃�H�s�%9�f}��Q5��y�4��o�`&z4g�W2;�
yr�G8g>{6u#|��D`�Ub@�[��,���GUc��>�g�>�*6���-A��v� �99��vߓ-D-�;$^BO3�i��Ȃ�I� [,��>����nn26R�>R����4tL"ÙҴ�e�aK�b�$���kp��\����u?OGu���������-!��oX.Q�9JG�d�~��~Jc��<J�O|9ྜྷ�޲5���ΦFV"�Ҏ��F�y�Ř[i�����.��$ד�T{�9+k5�I����&����)ۓǒ� �	��b�x�^g��'���L#��=)��ȫ����`T�in b8K��Q����beω��\S}IR�p)9�|T���������sD_P��3�TB�l'�\Ur����C�1����UP�$m[2�g�\� |&�pM�M�_��}7 g��dj��5��θ��p1 �$�IA�x��g�Fs��d�C`g<N���	��E�Ћ��?�6��f�Gv�u�� �Oy;���#r�*�9���d|r/o�A:��g��k5��P������l�m�����b}�!��H[���B��]��ٗD8=�~3[�����/@r�X3�w����SV�׶�Eb,@�jV�&�x�;Г���Y��/b�F�Μ䯚��u(y�h�q��I��eQ���0��n�Z����틶�ļ����v��SPQ+9LF��֛I.�n��4��5�Q������c�'��v�� �S�^���l��!Y[im�Z �Gs��G[�k�xn�|����k�~��=�%�A{w|�a�����]�U�ZH�:�>Re�|�j��Hw]\C�AYI�%�fMc2���-e��9�QX�¸�f��ۢf��?S������ߠ}���D��+����u���8 !%���Q<���m�-\q����;>�o|��N�8&K�b��4]�Kc�T�����;f9�5�|;ꟿoF�5!�9MM�SڛFP�%�K�# �{������5�\�wP(·��:0�'����v%�B��q0�����3H��.�]N�ϩ��0}>a���C�*�s ��/�Y�;T���||���3�æ�I�C���*x<�� �J���9P+�%��ǜnzx8x�wuD�M9[݊��$�_�
�A�~��Cݭ�%V �~`��Kmq���g�"������k��U�~滼���C�.�x�RǍ©I ;I�na�$t�M0I�>��aN1-F��@M]�]e���D<���E����W~�.�퓳t���>����83����ܦ`�Qe^)��[�;@�V�k���f��_��(��A�7t��,��@�d��,�e	�X"�M��8>��9�A�* BE4*��;8T������Ef���$l6E����|��J��
�������Ss$-�l�a�*SS�(0I�:w��cLE��Qd��;ݍ�'�Y�G��A�ϲ���%���|zۊ����L8%@ƛ���ï�&���柜��_�f��mINa��n�~�|<�m��^@~r�\���Yo�Ke�	-�̲�S�
��sl�cD|c�~�۷��	QP4[-ώ��[���N��� ��2Ѧvx��"o�a�uEY���O��/��hlb�@a�ؤ'[+"I&�����'�Ni�a� �]F��_�O�����kp�~��\��z���_¬�zRI�5:�˴��'�� }����F�o*̌]��R�m�Ld�_�[ν���r�vb���^3d�W�y�_��������QNN��ZW��:�09_TĆUI���������&[}���AN7x�F��T��9A>_�d���GY��:�W��7���*��VGa�1���潺;�Ũ,F���}ͣ:�]ә����aRG����Fv�Ԕ���� ���DQPL�B̙Q�LK�A�3rfI
�M��gߢh8�.�2y��Y��䇞�i��/���Uv��v���S ����}4��'2��Q�o��k�^�
�!���u4���i��QH���b��K? G�g ��L�L��o��[@q���p���ТqPL���׬p8�i�A�p�ӊ�e�o��pɛ����*�g���R�1k>����d��ᗜ =	x��ך����7�EO�[�J�uY�4�]'}��E���[�dXC���}Ɓy�<����6^�G�a�*ES/��5�U����������:�������PB$���t�z!"�E?9�B4%M:�C���<دC+=��+u�#V_N_y�R°#�DA��2���)&��<dT�r�uY�L����&�&���S����x�kUZ�\_F�� 6��pF���
G��R��i��j����:��˯9���j�+�f���'���@	���R0u9�l �D�1�jno�_�K3,��o�߻!TK6烊��چ�K��`x�3+l��x�U�;g-H�{�'s�=�_m�7ʘ;��$����<��)�H�i�D�n�@�U�F��4�-���߇@ ��M��[�4��NG�z
��"<u7�v��_�9���8F	'�{΄ �����x��u�4'n��1�6>8�~� ^�����sd�]�2^��2Y�Um��.��8ňI\�h0�+�1��˝�AĹ�vG��0i��:�ۜ(ǐ�]vv�d=���܏��*���xoE����%�M�xPq�KG �N3���Sa�3SҘ��p?EuշĀ�m���H�g�3���n慠�/̆���;rں�x:_�p�*B���0;�v�p5e $c��Z �[�F6��g�q�j��x��_J��$�M
;3s�ܱҪ� �&J��sM�#I�Ջ���� �]b��xh����������s�$����T��Qi���/ç��:�o>�E��W	I��7n�K]�&N��m��/L����� yf�gt��L�Wq�4�I����
*O[�	�ez�Q+δ&�pB���u���	���ڍ�]S���.���^��Hp��E}��d���7��9��$s�})l&�G	���<�Z9h��7p��N[[�]X�CGG[R�OVH���H)$om�&7�T��v2�m�[�g�� �ğ�M���*?n���
|�-��� ����Áи�'~:9͞Q-*�hP�y�b�Z(J�iec�t�Ҿ�}�u� � -hI�灧����16+2������c	E�L�vC2������q(�B��;�!�ꩲe����S���Lmy�~�	�\�OO� ����|��7�O2�+=b���[�m�?��t�D�_me"����uw'��>V`5]_b���#	7J	KA���.aF!�����S娦I�gX�L?
����O����Erc��)}m�sf�ɅǛ�sOuC
�%�9�u$n�*�^\P'����-�	�4�������A��E_:���O���{�G�\5 �<��+7n~��%��1%M� n8��+(��Lk1X���L�b)����;j'��P�~j�I��d�t֤�L~�ԁ�f�6�B&��M�\��&��� N��OZ��H���|w#��<��8�8�hӟ`�KUgHԼU7�J��P�s|idO��c^�)l��>�/�d�Q�ݲ��ɉ����S��=���B͑�V�X�6�#u%�Y闬��aT����0&/|�A!����rH�0
��%j[c����;<8(6�f�������~5ꤕ%}�Wj���d��� �K���T��;�JCr��<yH��G+�������ś�2�3��r�9��M�'G�j\!����.C(y������;3o�>=��@E`�7)U���5$�:]r�.��&*Z*,l�a�D��_	��!�  �װ�����Ӱ��9�i�屌�Y�Ҟ
[R�H���%��4 *8���a��ʹ�(%���r�O��\��q�~��^G|�i���b��s��N���Zڄ�|%�Srs�P�h-K��Hb8���~i�l�d��k�M:3��BД	���Ɗv�:����R����M�o2!�,����x\���[2J�IV����al�'��V$�`Op���]�K����'<���2���si��˦�{���*qq`x�Z2��>�c=&T(O�Q��=�Q��C�#�51������&�)�+(1Dh�d�v$�Qֱ}g�Z�V@/)���r	d�o��be䫺����+u=�]��u4�H�wCRlmn%�h©
�`Ky�"V.Z�ʷ�K�i<����ûHTä*�I��s���b����'�>(*W:�������uy�!���h�مE޿$��Yμ�� K�b,Lh|JF���U�aJ���_C^�;�
]L(����C��nl��W8�����n�F��2�t� ��:�o���i���td��j��1�8sce��8^R��e١��aڝY8z��6z1'��a�Q���!GKZ~��j�o�-|@̒�^[:iv��d ��C+�(���2�<Tح��
!�Е�|�@��i �;ٟ&
f����}�%9#�z�K�z*����0����ca���+!䬃Z;#N���+*4�}�q���EC/5�Y��4Vu�����[��0b~�?먲Wl���U/O��n�������`\0�{���q��a��3��C��_�����l�<B���Vd~���0� ���V��梺����v6���w"_�K��ٲM���jl�X ��%���^����1��o�]b����:��:�$:�d�o�s>E�s rg��o�*�f�~d~�m�es��xz��@�P��H�V�嚈�p�p��9��A�m�nJ�zm��NK)�ݫ>~i���sc"�HS�ܲ�a߯��8+��#��˛��\B�IpQ�t�bgc@~��W;P�+H��55w�����>��Gup(�u� �׋�`�}�zHp��d^�Ͼ��2h?9s�x�zO���T�n�h�~ع�j� _��lt5 ��n�_�}�₁T��Z4�ʯ������]\�Ho��`��1���Ԥ_7r��8H��$�A�x1��&��֔
"��a*T�����A�B����՗p�~g�#��wC���ȳ��!GO���%�s|06��NA�]N��$��h��Ύ���]�����n��g��~���ljf����Rђ�=B��	���M�vU����7Ub���|ě�.+7��!�p��,�&�@�y-�Y�z�������0�枈�t� s\�+�>GJ�xFջ�4�ŪS<-����-��cXg4�D���; ���i�����  �x�P��*>�)�H�!���l�;ߓ}=Z�Q��봺ø�#���jf��Z��EvR-��zk�Ԭ�8j}4�|��{�;�iګݐ5S�������.�%��9 k������F�X>�&aM��C�
�":F���~wvR ���BP`��}�M8V�x\7�aߡ��-�O�	A!�����Y��i+Fg�"����
v�Y�=`wz}�)��ue��K�\q�܌�vNK�?"��qX�"r��C:j>����u7�%j�2}O2h�׸1ˠ��-���IՇ�Ƃn���T�(�u�C28��7���&e��r��|�9�����ʄ����z�r��U�u\�)�.~�{����1�V���S���8z�v���E�x�������&���P;����8�i����aV���|��Em�cI�ŕ	�S�K���,F^b6I��-��Z*L�2���?W���:Z�UF�����-zTz�Η��:��KӸ�0Y�qN�����zj��ib��Cg�mS���B3��h���/�P�!�YF�	��J�8	�����Ep���7�k��:k�8Z��\�Fc�QF���7���zE�i6A�����p}/�2J>�0������DCE)�v�~Kd����N��h�7�y}N���2p�79����� .i�
��C��7]y�������P��
Z�&���c�Q��/K�,�z��4�\�t�9;�gf�fD�t�aqD�3v���]�T1<VDj��X�s�')�
�\?W�&�-r��@�)u���q����2J/m�E��J�Q�du�O��h��7i�S��Z�Og?���tzPW˓�� ��D�/`^�<0JJ�٢�u��u��%�4ݬ%���LуH�R�8��T��U"��aO�U[�ͷ�Y6R�0D��T�A���ױ�w�������Y�!��i��I�ƥ3��Q����B�0�Åk��	d�LNkK��wqh��]^
�[�ϳ6yJ����N~EW���/�6�{g0���)�)��C�w+!a{9���� ƫ+8)�y���#|>~5&���v�/�m�E��EcT��@]�1�������mkS v�~k#�Ϭ��mN��w�s�g�rb�Q�u�w͸��+����Ф0��K���ݾ�8�2B;R�gT��L�Ik&A�=����F'Ǔ}.pbt�ȓE�ϮE��E�֤j����i�zt�p
��
U�J����І�F���#1U�_1����*`�n.�Ka���T�HK�q7��Ѡ�'i�w���d�yb{�`�><1ç�JsOY��Zkʇ/�K6�-�^�/L ��w^�|b���_�YhY B�J����T�9�E
">���5��Mp֊�҂|<�q�o� R+0��.���N�1��r��1����kn^�(�$��H'�g$�E�\��O�k�kkz��#n�2�3xT(ՏFL��!'���v4��X�Ĉ"�N�y����p`t�6�����D�6��I��]WW�9�L�P�~�P6�{�/*�ap6���zT����Q�������N �^��Y�ȉl{�֦҇a�9������@,7�5|iL�$����D�H<���k��YӺiҫ��v�L��4��d��j��7�D��&�����<NQ��o��')���R4�.g��-7��u���b!�φ�θ0��).:W�q10<�o�ܔ�I�t�-$\�{�.gi26�*��>��5��ٷlK6�L���r�7���wo�D���.SG�c*�Ak/�S"�����^� �X(z��!�
�Ԛ�Yb��ӃF�r�NoS�B�&[e!�d�^Nx]���)
���RñP�F�UQ;-�<�S�+��#7�&����W���<���.E�DR"��7i�X�������m%_9ӲZ���� I-!h"����|ܸ�ȷ�j�����1�v�z"�������y�T��b�F�a��R��;����U+Wq�L1/��� $�bF}[7�a�$�b^�O}���$�H�^�͏���ҵE�.�Hl�6}�0�[v%�� ����re�e�&��t��ȫ�Z��$�[�?W�I��Mб���/yL:�QD%�x1�� 4m)�r��$ ��sR�E٧�p鑺ŷ���D�R�rg��mJxR��[�C,;�mAM~�9���^���[D�"���S���i��@$b�hs��C̍vq��p���W��a[�"�	M�#���"���aX2�P�˙�J1�V�M�d`iM7�{ ��%��H�%�$�E�ڋu���P!�`����c�A�}���45w$�$%k0�1bVM󪘥�l��s`�h����{?�' ��u�����D��L�0�IO�8�D��e��N�+e��z'�߁��� �rN\j<@��J6Ū�%�qVh��e�G���%�i�dn�!ç��#���LpCx�ӄ���#v����e�N���CK����E[���"��e�W��]�Yے�VtE���'��E/�q:�t�H&?��5hm��/��� ^�����,�G�'?���.�#ݬ�O.f��ݏ������\O��7o�G�FY��>7�׳z[��w)Tn�T�ԃ�E�oz�^���Rz틄����b m�K>X���\L�.�9�D]Os��4 �Jn&�&Q7���א<��dʡe�MY�B$T�e�4t���b��J��Ch��F(<jj8��aB�3��4d<,��Ӵ]}�d4q�sP⟼O�3
ÑE&����%H�jǾ8qͣrw�=R9��j*�%�
:�C��p�D�h����=��LX��ަ,�����ZeB�
V����/����+�I� ����y��I���?�����aF>�	����@��m��=ďzA�<4�	�]O:�Bv���	�"�Ip8lT�2MZ�[_]A���5�x��/@Dlp��e^E����y�n�6�뫓�c�ۛ�)�$��3�^��X:�O�'��$]�>P�&���
�߮}��W�^&�����~% ����YB��V��A��o>	l::C�j
Ol����(5��s��Iq4�S�O��D�̲�p���U�U�_S ��4[	��TcP��4��;���g���ͤe
:���}9����ZE���Jn�Fm�I/�y=�c�ӣ��A���O�Ӌ~�#�*����_��י��~��E�o�IR��8��ц�F�L|Y��zhu|'�c���Xy�'�a�ѐ.{#tu
+��+� ��B��g5�]s��a�#)�%{�v��"��G�; j�Y`x�D;Y(�a���ͬd�cKڨ��7�x�q��oG�0m%Q^L�OD��"٪���Z?ϱQ3�춙��A���M�\�^��n�4@��ڌ�C�/��F��������j�c\�phΥ�f���l��;�q�a����y�S����{w�c�I&��,V������1����Byd;�aҲ����?�ݣ?0VcR��M0kg�k� �;] 	�2Y�U��R��|ڎ��.L��[�W��
�v&�S��dӑJ�*�	�/�*P�91�1m��x���
,O��,@���������4�-��K�5�=���@o�d?i��,e��mYj�[�H�L2�-��eåݰ'����^[��/�ŲG�� �M�@]����2
M��ʩ�8"X��7���!=�#��J~��@�zD�SmT/C�k]��8�8}�� ϵ��NSQ��R'Ԫ�K\��]�36��,��YV�?)�;���n�/�W٨�����Z�%Y�w�Cӯ�Ci��O+�N�yU�HD/7�F�P��5�J��>l\�%>�+!�[2WC���|�F3\�U-�a��?/(n�$���bM��=/�,Pp�f}�%��i�K�-��􅽻c��L6�<Fo��2i�l6��f���{8+����Î��/`�T-9n�*�%}f��C7 �Q�6u��һOV�Ί��x݇nq{���#�I-�����NPڮQ���`C3e \Ԩf4��f����N�QW`��6QB�r�d/:9D��·:}s k�U���ǂiաo�B�RvTG�`iH;-�C�x�!��П��ˉ��Կ��`�U������ܷ5Y}UA�:��K�V6��I*^��I�M:I:�V"7��n[�"�/ lȐ���Y;HtM�v%���+:M��X�J�+Y��G�@��)�f�Dv���Ys��_�ڇ���U��-���Vdn����fL��un��Z~�fP���pתJU��{{h�?�8G�ZD�}>A�����Sd216#Oc��S�N�GK����[�4�G`�����܍tV����h���m��������t[_�%����@`��&�K��������Ru�C����������7<}}}c��#ّLofF���F���~�I� Ѿܞ�2��4�Im�H[�%kW���6���B]��I�pT�4V�[���G�I�~�OT�Ʒ�,�n;����U��K�0���G$�y�z9�e���%0"b?2��},T���q���,vE��̩(�!#T��CR���]~�a���֡-Ғ��{��Dq�u�c��w&�vɦ��c���s�\`��O�8'ڜ�L�̗�%�f|��0����;nzk@5:�`��8G�,X�	�XHF����� ��[��p3��*��$;RN�� r��'e<1�������qf'�f *6��e#�/������_@���T���ee����1�)F��k���?�������J�#<b�S��v3"C\;�zҝP�H�Z��J�{�"��G�^�+�7ޢk ���[ >�dbK�f�a�H���',O�z��5��)��=�v��՜��܊���L��Z�އ�|�D������J�M� �(�$�������5#
��@e�P��C@vU���h�禓�Ӗq�M��l=�����@e�V׌n�ۯ�;��R�\�e���|���3���V�zc���|PB�؇��Ñt������.�^��w�7�Kp_�j1���UA��Ay�e5�-�����T>Pg�#���/?VfpVB�8�3qxak �8��፧����Q���
�}	
�� �vn��[�����-�5��!�HW�$�Й`OA�|)���n�~��"�~�Sx��CE%���̺<�.P�Z��:6�g���H1Rq��9u${c�ev�H��w:в���k0;qgo�ʏJ����,�IN�<��^����'�����Kv�۹���W@�j)��ҠOm�Q���lY�[[=��]����~JQߢgI0"(ju6�����u2sE�)�������b�i��F��j�}{?�`�98WmҤ$$�i+_XW�m1�b\�ҁ86�� �E��26֏�A�P�P5%gBo�R:=ٖ��iL���1����a/8߫<s%/�D/4C�qa�̘S��.��ƓM4^����S�8 G6��}��Zs cta������^��S�m�qSV��O+���ځ~�O����mBmm>+Ե/�Buƚ9��_+�S����J��n�喆��}Q�9�E/m6��&G�+z) �|����2�Fe�"P�x��:��_�N��'}��lgЅCR�y��:1EƒJ-�K�S�ݽ[m,=��-G�p�0׶l�")*@�(Ʃ��Y)`	Ü@��i�?' �b3�-
9�c�j��?G�$�N(�yK�; �8�� �?�@|�����SȪ�d}�����т�U3�=&b���ZK�>O0c�8�f�a԰(,�pQ��⩷�H�FDl�������o#��٤���ˇoC[�	�c�O!;��<�s
�M��}��p�BbmI�{������/Vvk�"L��j6ʬe�k�΅���~�|�f�I̬��l���x�pZm��|{8�<6��~A�1�� �]��u��#��� B���3�7���4M#|1͔�7��4S�57�X�9��
�'^��C���t�і��L�1���
(�ʼ�� ��n*��0����R�I��9o`L�qZ
v3����U5AwRl��TO�ֱU����WC�dnʩ�A�`�R�^���)��3�g����F���LL�K��Gj�B����\�s�g�jݑ�,ڐ��'�����c�5�I��y�rq@�ޓM$-➚!2\���Bf.N�����s�������?TefD~��P'����n��q.�Q؂F��b�en�b:sa���ִ�~t���I��k,���u +�.����pn ��N�9��61�gn�)�6���t�*��)�����7���2p���-n��W������A�ukmQD�t��d�Yj�5|��d���s`G
�8�۲�X ��C� �.�$�;�d��Q��Sm�{wg��,��G�)���Y���+{�Ҳٛ�p8�Z��ۈL(C����9lġ繳����褐mOһ$I���s�S��-���n��*v��˙.u�A%'NS��)؁��FZ`{on.,���_�T��a�<~�i���������M1@9l� �� �
Sh\'�8?��[m�f#l�PJ^�@�|@��Ta��㘛A��iUr��2wKN&j�,�A'��x���D���P�d+��ا��_��1x�)�u����l�s�x��� Xq�3�Q�g���L�����y����/�ӂ��#������'��C�1�T�P8�k\�
���۬S��:���g&�-���]������u	���!�?��p�we	4���m��qǘ���H*	F7�ӫN��F��٥mU6��\�m_;���c�]�>�jQ�t�q��I$�� � 7� ��l��Պ V�y4B��Ad%Vs�߯�Jfp��I<��e�:V�@�/��[B����0��|lAp4:i��0�jtn���-�� ڼ�J��YG�4G&}�����Q�ц_�	:41�Lt%���m��9�+f#sJj�e%�I@
�X����e�i��,��
ŸNZ_4Vφ�W��#Vz[Z$��H|
�{U�?�G�$}��c���R!t�8VKI���ǗM��hI�%<t���F3@��s\�+Sl!2�}d%���r(kǑl%/XT�R�+6#�AXy�.9�.	��e�~D����(��G�ڵ)%X+/�|~�0k�O��v�X;8��)U��z_���^g�&_f���~�(�Νڦr6TB(�t	����n�'�����|o�	���_��3����zE��Afc߅w�Ai�<�c+9l)E��U������(:��p8ec�A�*���ថ3����O�룐���M��8�>���_�`�1*x�r�z�}��6�3^5�,	ms{��5KCC�T�&3
�ó�ǎX�c��ϽWjkW:,�b0�cgh�ƿ��@\���`,~�]�o�\L��&]���X*�5wEv|o��!t�l�S���1Fa'b��2�p/������GJn�����:U�����Z�X�*ޭM{̶�h���O%���3�Y`��&Q˲��hW �-S1` �oN��a�׃��Q�-�(�MP�����!T�n��Y�C��J� ��=�q=��-7. �+��e��|��0Sv�?�F�=���0��ui���.B�[�1�'�4.<��D��a�k�}�vE��B�JO�^*�\v��N[Ñ?_�i�ȓ��j�R�1�ՠ2�[��P��Ԉl$GK��9����45|b9Q�2�0SMe���i��^�}_A��ۜĲ��<۪.�p	�y�*o��Y�$������x�4[��Iw�m;g�����[��O�2���VU�Ҵ�	���TH�׷�M(Fc����-ƚjT�#(��n<������D�r=uN��P˄[��v��=�#^�ěI�
u��"�J��ջT[�djn3oq����ц/X�4"�x��,��NR��^OUg8q���M��M�$����V0���״j�+?N�=1c�q���q=>�Ì%b�zE���&䛓�<�ݓ`�W���R-mp��.�����H���+B�pS���t�3��#y�iE�q���@���c� �3w�`	&�󑦼�Rb؛U<BR����p��\�ρ�Y�t����-���#���%��f�[���艑�+8����Z�uؖ�]�������=������;�q˘�����j�'w[��&w�0�iX���g �CZMX�S��2)�.�� �a�6|�K>�6ȧ����Wݠ $���Gb�-����e��L�/��v�FS�|��_��:�g�ݜ0����r9��ظ�|p�ґ���p��c�.�V%���;h�}'�;a�a���;XA��=-�)�s��[\�[���^����Ւ������������[��/���[�
t�L�A��7h��\6x�YE�x/LT�����tND[�bjSx�]ߗ���OZ��~l��.n��>ܓ���U�&g�mi�:�.I��K���d)f{T@ �<K��I�]í�M�"�s�Ȓ��IX�������\2���M�ױ���L�ͤ����RS�'U��=ࣥ6�ϛm��j����g��k�����G���C��&N�/	yGF�y�޴�]�|��fC^XwD־��O9@�4�BweQ<��ͼ�z�R)���Sk.(w��pb���G�@�=�^7�Ȁ��Z�.����"�o���AP�� �ᒗi��$W Z��&�����)'���DM&�1Tu����B����#>EM��x�Z�'3�\�2��CH�ֺ}���tI��ݸ�#ۓ��(Os���P{��.>�i���^�V���"��{��{�hcX�G�I���{3�p7���ڂr�QqC7��R�l$�V8�<�p�i_�f�i�P&{l��~*�s�He���1����F�K
*���ƙ�t�&Y��^Kd���8�M�xO�D%f�����L=u ��?��Wp]T�E��Ŏ�n
�dG��������Ud��`������m�_̜�j�1?��r
o����?�^Z�=H�x�iE��!E���p�ߘ1�G<�e̝CK7ޠ|m��-B����M(z|\�Q��xn�%�w��߁3%�T���R�O�bm���F*`I�$T>���>/fj�x���֑���16�D�`�R�1-E����]�:q1ǀ���"��r3����������²"�cʧ� ;��z�������	�w���le|z�=�F�Q��v�
���~��t	�𘱈���ۂ-���B��p~{����<���^9ͅ�="�l�'.d�^�j�^�������-YQ�V�������,g,���B��o*��O�-	���	��Jn*�`}rrjf�._�����]h������ZS��Ƚ��.�%�a��p�Y�&Sx�@�aqeh�^�Ş"���J�aVz\���
����kꝌ�^�m+�e-��!V����f$��:��Z�i/9�P}Is\⴨�^�Z�^�v{]����K|���֚U�\�2A��3�ʚ�L �#�Kg���_O�O5�$*t��p��I��i<�cOI�;k35�i�y9�\�]-��V���ِcF�������@�$����v��n�V~0'6�}��![P�C��u��Q�����B�|T���#D�Ҿ��h�P �e����)�,�8�8h��N���^�\�1��:ǂ`)��:�V��e{G�=�o���\�`�s<O&lQ:�Stˆƥ���_�?�1	���`R��qp3O%�ԉ�Y�C�A���LPI��#bO��JM+�v��{e��rͮet�R{�ǟ�e��c�S	BSO�~'���U�H\�蘂S��ň�	�sV�:Ł�N�Ǖj�8�"�?�%��\�B��>9�2��� 4I���+/D��C��`���A-8B�/�K�?|�cKV8lT��6^@��D�Oh�
�W,���
��~����oߜ����,���l��b�ק3z�M�-��g(l�6��E��Lw�qe7*𱜎e���1rǰ}�6B��փ�Ny8��z�
��'�%��3I�U.���tc��6L�o1�}�c/� j�>�EN�ތ$lGZ�-,��5��7��:X��M� ��C�H	~9�?�tI+�f����k�ȣ"���"<2t7�5�%cv�}��3��o�w�P�`I�ɽ�"О|�&"�"��GW���մ-P��bƝ�J`ݫ��A�i���������WXp�LGm�w=+�	c4�U��"Xݹ�'5��vndŔ8�}aϚ�hB`~�H5Ų���}���+��"��0r�Q���p)�������m�K0��2k���T��.�7e��?'
\}d��E�dP�~]�ȱi��5:�B�]#��l����ݹ]�'���R�l�*�;�4��\��n�	aY����>�RDZ�!��J��w��7��� ��Ⱦu��W�G�jm�������ڱ�g�g���/�:����l�_E���Z��6�c\�̬�iO�M��B�1�e�Kc��>?DH��':a�!�$�C���/�<��fW���Ğ7D5��eƛ+<[ǿ�q�f���8-�A���,��@�E��(�QmT�Ǚ<���?�=�Z{�"*d���z�������L]\��Ht��;z�e�H������U�5�W`[6p������������,dI|�?2j)��X�� �U�5 �g��}��|��.��,�o�p^+pW�A����/<�֌Z=�h�\V~@�� ok����s`+O�m�Hl���ICq�V��ڒ7tZ�tѵ��`WNJUF��)���%�	$��MB�S�5Օ`ug�&b�p�]�q3��\�	�M:`:T�j�2��K?2��e�پ�]�\.?,@����<�)��eM�#�x����+�>�ڝX���?�{Ev�H�;�wEH_iB���;酾��8��;�+�.�p���}�1ck[P�RQ�ۡF1q���#xi�SY��?�QC>���a5�7�A�͖X�q\��JO��x
�����P9����;F7���֬���s�<�;�����A,##�@���V
҄J��(�0{�X˔��̼���m�sy���	��Q�2�SH�pb_�7��<�A�!=������#�Hz�@�R���L�l�QC.m�d ���C���#������
ʞ��8^���0-�"�2?u
���66�]��P8�c\��C���?�b:�|�$�
'S&ݎ�g�8Y������z���P�ɱ�S�#Ѷ.�Lơޜ!�������ͺ<�7��ۗJQ[�VV)/.��a����$4=k�sD��y83If+�Mt���j@���{��Ѵɗ��S�c�-��f��_K/��5�]�sy�,�õi>o�2�FfƽU��	�d/d₍��=��c*D�>��U��]�C8J����l[�����n'XmG��b��Ƅɨ be���2�3m��A(������3�ΩD���'G��' c��Ǽop��7�=���|qg����5���������, �Cc7����Ev|�+a������$|ҀǫTDo�(\|���[` ���Bwp1���ʅ�2��)l�	�7���N5=�ad]�ޤT%g:����^��n�����m����4��u�]
��]�+��ҲG�1H>U�����(5�H���1��x�z�zUI�Y���t7:4��LE�jB
Y�)̠KWF5��_�C��ztI��7U����zY1��8�P�m6U.�cfW��x7*fe߿����j:t΄�\�3��I�Q8����Ů�b�^#~���gT�JO[ �Y{p�������TTW�ʍED<S�0�hB�a������=em��糧x|�.�9z��K���?EKZ]�?��	�h��F�E�׷��N�� �Q5Ck�~1���-���2L�ܵ�^|zB�\���I~�B{]�5��~����٠<YxFLF�96s-�"��:/��ÉqN&=�6����
c[t�%���:�~�Į�94�m��I%�������D���	u�Ó��/�L9���Ol{����:�{`�A���+�|��o�`0�&ܝ4�S�l�)�8<O�[BZ�yK������$nCF1��v��Q��y��]��S?̣>PF�:�5|���{�M9��Y޵e�B:�Z����^N���#�D�uʺ��z\61CfKXL�����ۖ���}
I��i��#DG���ݖ���U����	��gۼ�˺t����)ɣ�n��$K�t�61DK��-�%�^R��&�ۘ��7�7�H�t~�<������kB[���_Ь�k�~z�޲:8��+�D;5(�R`�Ԁ�-�4T�{�!I��c\x���)��0�3c��C�.���|����t�Y.��c����&&M�=�.k��sk�x��Ē��}��t�=�0>�R��Xj?��C	FS2mٔ�N��^���5ГY'�,�wL����s<��'\�/�ߨB}��s���I�a��ϺB�K鍃�
�
@�5�l<�
�c���3w#{i��O�\˅��O�y_i�p����t�R��*sΓ������|�e��O�S=��l�u���8eH��Ă������j?Ul?`3"�(�9�t �E�6T� گ�'�6�`_Y70_��d�:���~ܢ0��+][��L��9���.bI��&j��"�A��$ޗ��㩌��j[_�����.�n�ms,���KM�o;Yp?�n�[�F�/�_pp��ot��a`Y8s.�:��2=�&'E�$r����fL�#�xJ�h��{Nd=uPRS)��w����a1�h{Ⲷ��:�%�8�ATmW�>>�Eڄ�8�v�? O��sI�O3M�R��e�2^-�F3���UYRӅ�q䙨��W�T�{xGb��uO�_�;i�24���$��e���#��(��)kz|�CLM,�[w�<��H"|0n�~:�z��h~�F��T%B�8$1O~)�N���$�W7���me��% .36�NPA�oWz�'��'h��M�?�qs1���jz�{.m{3���.k�V��?e!�SD����H�x��{l�	"2�2_�{����W�l?���=�?��D��mA�����(�W�L�f�����:��%��'�D�he0�0�\[���=����	��Խ�<�`��tM\���$�r�$we8Ń���io�q%k�3�k�j����]��]-�ʏU8E;��yL�d9��O��|7dU8]tw�����m���B�T`Q!��}k�˗���h�/�c�a���@G�DJy�ڎHU$��#/�I1E��T*������D�o,�whY��!�7G֡O�J�XP2�x�[�ex�#�X��F\�D�X� r�]Fe9�7�7áw$Vo��5�r�q�����	Y.LPg9�����8���j���V[	��Qt�������e]&�ꜰ�����U�Sݾ�"�p���۲bu�NP�7�V���W"�S�ۘ2ǗX�X��n.bEbP�D������G��S �Y��,����n����]Q��0�/=2�[p���K��B�N�������
ʵ0����H\���Y=Ѭ�wg��NW<�\�"�L�����Ɨ\K��L=�y����|��e��x{��H��T�՘&��d�C8j���C�a�Yp2��\h\ k�Ga�0������Hj���n7E��WC07�BO�����m�j�L˱3���W�%�5��/����ȉ���tt�/�5�Xgk��F�;�2^�Y��(�+L-�R:���;�
T$&�D���g��ASO�L<o�`���v0��W�x�R�?۠5�H�j���H���B�S4$��� �����^�҈oO_��oѡ06��:�}7G5��<r�i����w1�R
k�>����РI{?r�(X���
�U5����$�s���,�K����+
zS����!�������E"���s
�ǹ���J#Gm�W04z&[,���,%�YnM�}�+�JGx;�טH7^�H�ڮ߭����d��L�ف����_�R��͎2L�v�_p�j�x�E@�6���dPB�z]�h����.�O������d����	�ڷ^B�'Yx�>bT�MMIΪ6j/��nWK=����=X˯y�+���G�{Lk�fS)WAc��#	�����w���J��(>����3�>\��Hn��N(�R���ͦqiK�S3i�k��%|��,eSA#�G�o�RW;�%�I�|�Za�?��o��,n�3��>�h>�*���v"F��úh�3���eU��!�� *88 ���D�N�I��T�Fao��B�
��^�lh%�s�8��[V��4h�|\�j��[U��_e���S���Fw���J��ѵ�Fl�7TSeǋ�ul>c��Ej�8�0�U׭��W4����m���{�����_v�U�p�F 폂w�a����M��%�@R�+8X��ZxQ8�0� �^a.����64������(���A%:��+ɱ��zw�r���>MP0>�>�{����J�PmA,s�)���h���
H�hU1Նv�EkTDu�qT��T6�6�OШc��A��g�c9R��k��OL7��6���(K�a��i�lG���/|p���>I�� ����^A���sC�B��Q�kj����!�����H$�.>�|v��ko��t<�t'���`�<�`�AB�f�v~�mw��L�2��>�3$Ԭ�9��r�s��f�9I��tBL�h�[��W�i������,eC8Ɠ�'��ԑ�ӈ��-������|X�?� C��$��H��8�=���_�Qq)�HG]�Z��_�GJ������ĎiH�yP�56�����E����ݯ��h�g�'�đ	ƀ����W���=F_��^F���A>����
��V�Py��[�
��*̹ sT)��ˏEgf%W�h�b����
?�q���vF+�tW<ص�^z��_�+�	$��2@Glg����*�X.���n	����4~02;�c/���bꉃb��c���JY/eY�gbQ��ϕ`�ی���@�V�^7<b�؍F�ǮBg���\q�4���Z�XW�k]l�te�-�V%S�De�e���~W��x�ަ-��t�

�z�&�}O`���)^�"X�6X�:��bϐ��13��:+Y��@��� 1`�h�!I��,��ġ�"c�,��ZX��>Z6��mP���H�D��=#�
aGO�����&`#p�85�p���+4 A 8�@ȠT�+]n;S��;g��|��ز�o�вZ��=�Vd+�7X>�0[�:����^{gմl���tY�IIĬ���QX�@7��a^E�X�-F~����A��B\:�u>�]#�&7"��K�z>n	fD�*a�ҥ Q3�vؿ����3+i��ĩ�B�
+��<�f�+�j\�H�1�rɱ��ly�4�U��\����ԉĲf8le��F��.UNV@�(S:�{$:���{Dn�g}�Z�&�x}�g`��	��3�y�������j�I�����_��G�nc��u&Q���z��G��jc�(�x��i��n��5:�/�[1)M��?� �)�<�I��:��?�cqf�DMak<��|�8��tȭ����:���8n5��(����6�A�I8� |���1�E;�n# �YƳKj��h��jg��8�
ǧM>���8����L�d�&��(�m��H�s݌09��k�!fQ���uP���Tφ{���p�
�4��Z�]&�WH�d7F�����jet�G��CL\���Y��k�m<��J��o[?YIhp�mdWUL1�m�l*G|	�dE� �yu���Ɲ���^$|�Kx�fG�ZM��]qd��HR\�����)�8-&v�\<? �ၸL���KQy��.�~E#�����@1]��&����R���H����y�E�����N
�
q�2a��Ig��B�²羇m,��uv��1ĉ�@]��p	��77F�A6����p1�k����*�l���	��˱�X��W���"j��	�G�̀����U�����B�X#��f���n+�����������g��1�Q�:�k���]�L3E5��!������Ү�-j�:ibv�`yd��j-�B���J)O��D�.��S�Ͻ��|p����	��MOՂ�p�h���g�=BH���ח͜pR��=C���^������2��T`��0��#`"��Lf�k�z��t�bK{S:�yv�0�_� �����E�3φ~�Փ�����^n�S;����Y�p��Qs�H�Z�Kb�nV86�-ul¡��`r^Q�=*7A��p療`�Ǡ�غ��WX��_��l�wɝ=���9��9Hxz��Q�~\�Ͽ��ѿ$I8?�1_4C1�׋�`���>����4x�d�z�H���l-�ʢ�⠱�������cO�����\�F�8�����p�&o�N�Ӟ���ׂ�|>�T_L�G��i�)$Cfb�`	B�%��Ak�V���=���.���ۼl�Yht>���ƀ�
p8I�D$4�o��LFEab3��5AP{[��U>e/ˆ���B��N9I����&
-s���m}�$k��p�$�����I�G]K��9Ґ;�!\ط�s(�6�%��|��:�ɪA'@�B���0C7^�C�ya��3������_I\-��S���#.(��	��F����ng��w@�7���{u�7�E�'M�z�r�� M}>�u*�o��ȮH\���!˸��H�	F�S8�*�¿��oa�VJ���DEh�ٌ��ȉ��q�Ц���<Ч5G\:Wd+T�D�ڔݼx_a� �d�]��-YƤ�]��M St�e��)�]It>
� h=*J�x�ƽ�Y8>�V�%n�2�hhe���#��h�5�f.��{|���c��hx���7�� R}ukO����?������A&��"�4D�$�F!i蚰�oS��@?��m����cAx� �N��[�K�0��}|��zY<C1��W����^	�#�x�
��A�1��-g�)K��;}�ӝ]��$�-XH�d��҆b��J+z(T�N��١zV8Cjt�9�c�V�#5C練����_sd���/;�w�H�Ybv�5�ﲧm�ܿs�������]{ �s>���?�T`�:�Z�ҙ-��"A�SL4�$բb���2��%�aT�[��oic�ˀ��:J�F+��]�#�a����&�5�qʠ����|��%�����>q�!u�a��b.!���A�2̛���Bv1���=�:����#�&�a6���_C�-�]zBs�.��Ϳ�B�Yy���~�҆+��C�ҫ4��7��� M�� h����5�0�΂��]���UI�����_�Bt'��{��n'๨��~�D��������ML��TX�<L�X>�}�|��
�o��O"��~Z�F�$�Fd��\N��d�Y<�#|M:)&e(
�3��|� �]�\m��<�ڠ-��^G�՗�����N�����G�1��_6�J����[>�#5���2�^�����
�9����\��*�p0��z�\��0��7|��e<�M��
�1J"蠔k�NS�g1�I	��0�FL����Q�j ���24 9w�a~�"-ݯ�I�P��� �����~�x#*6J��F�����o9Ԣ���YohL��n���6�֯$��J�Z���!ɗ~�V
yk�2�R"��=�hl��F��rC7���#�g�����sV�