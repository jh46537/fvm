��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)������ɷ,�i#����W���J �~�o	�� dV8�_�>a+����Im��p��}͝��A�z�	��s7ᯠ放�����:9GM�A���ܺ�R�݌��L#Ʋ؜���Y�������
�9*x�&䄣Rm�݁r�oϋ�Z�^�Л��L]�5y
�?!�
h��}��w��)�I�ΙL��'����:-��1!����D��A��#6���5�M�,��u�;�tHP��]�bN�)�R6!0��Jm����/R�����6���ǤI'�L_Ŧo���9x!�vJ�������7��"ڕ�5�Ul�]We���NL�����r����8W���m��_��{5�[b{,:�Vw�b��/�X�H��Z@5I�	�j'��~�9���Vh�/GFw���Mg��68]��:�	c�D��֎��8V���# ��_��9��&@���`c�J&S
� mq7X}����ʠ���� �h n-,͹[���4��QPsl�����MMg���)o���OJ&B`�B$�t�5�z��䓡����<)e7g�#��,bk ���J�!b�X$O���iG���T�j�F����$j�n�w��M�����w$۫����}���J�Ԑ�:�r�h ���m���)؁ƍ�neZ@x��z  ��JK�|�C`.3K����ho+��E���Q&��v6��a�*�i�������m����BU⢏�>xx�p:����5!n�=`M���R*��S��ͱ�:t�l%a��FL��*���}0���I���G8""���+��5��cqlA��*�V��[��NI1J���i6�W���m�M ��z^9Y�U�(��y��Vl(�Y|B���	�]ݬ����?�8���;|�k�j1F��$ aa22+.�<��A�k���|8Ǌx3V}m%aY��\�@�Rs��=��{ހ���˵V�L�b C>OE�t����n6%�l!@Y�����#��@�}:&���-`�7<��p놳��,R)�����vpBى0�=����I���f����y�����T!Ol�&;�<��*���)x_�Hdb�to��O�W�k#�'ڡ�A��3~J*ۣv[��154ˈ�._��(4`ӡ�	ӾEEp<õ���>��78�K$I�h��h��s,yp�������
G���*��6P�h�nX����W���m3�8g�����N���u����a��Ʒ�AK���
#���RB�����I8�ڻ}�e�U��F@���
O9߽z�V��|���	�q��w�ɋ�V��#l�Tp|/��Q���җ����.�Kd�M��D�B}k*'�`֠LU�&~8����B�H��F�FwhI�7b��U��� �$S�ez�ߪ)iO-�� m5�h���`2���!�шhO(�6���d�G�X��������jU��W����M	�\�.�HfՇ&a����|o:=��m��e�,��z~c,B��u�CX��������t^�wBf�(�
��\�i����53�q3&����'�I"�Q���Gh>�>5�T_�_�+�s��1�_���C���ʈ���Np����p�]t�}������D�4�qm�TddjD$�3f��G��h�����-�?�FEd�VV�p)�&�KY��7E���W�4�`ܞ��� ��Si�L��ұ�aS�{@X�U΄�����M=C����.�l��Hv��uG���s��B�k#,�#F��������� ��H�C\Y�
�~X7�#Z�z�:��#�	LS�H�4 2�5|.9���� ��
c���o�6��̫����LS+DU	Z[��rk����ظ�i�ۼV3�0u�������9�*n�dpf�?���}��R���W���1�����͈�?]�$�}��]{(遄���b�.ߨ�ù$+���W�]��҂�����rZ�?9��G�Td��i�Bs}�:�,C���vk�[��7\-Q����&F2c����k˴�q���y��YEP����"�	��(�)?�>�c���y��(p�u�(;�2LBqf��o�Y������d�wҥ��g���ME������;u#���N6{;Sh����zį��',����69�?e�Jx\�례%U  ���Eଣ��$��y�A�z�ʈ�$�2(i<΍�~�����j�[ge��ء6��m�(�{S$��Ǭa�l��B��D�%���s�.s�#���dȎI���4� ���;l ϒPm�fչ�Ц3� Mυ=�����h�XP�Z�ˁ�|Z �#~J��ss�8�X�G�y��v$J�_H�o����ܩ}O�y��WaJ�s��:u������0nB���.:< �բ����㈴�/�Q0��ƹ��:`��6+Ҡ��j�����v},�@� K�!`W����%�{-]���9�^J-}��jw8��~4al+�B�'6`��{a4*T��!��QҬ6}�/�
En����nR�찬�� '>O�!�^�	8��-���C�܆	����EƇeK{_��*��nٵ� ��@��!���M���T�J��աK�6��^e�zgB=D[�����pSGF��\��m�!'�U�=�4\}mDb[�G4С?���i���h�evS��^��˃�!7��]��^ΠpD�蔅E�k�@p��!X��6t��A!uC)�!6�ۓ�"3C�$����M��z"�{ �vzM��=��2�3�?~�r1����<�b�RO�,#q�¯𳺛B;��� V��q��R�Yލ�`����fC�åE[f�����s�ޙg30�^Q�ʪ�٘��;�(�����p���������F�܂�آ����.�xㅊ�Y-��$��[��角��w�m
����o�km��.gz.������1��� /�����}>�5~��8X:��^1ѓ��X�D2�aKY�]vUx��Es43j8
�qҹ�S����G�����Ʉ�o��}"S$��ȭ�/�,U2�kD����{�1FMq��=
K�1<cܲP4q[6�	o�8��1ߩ�O�T����tJ�W 6P�������}���̾3R�Cs��qC���#p?��y�)Vnװnv�@w�H` _Ȼhk��p� ���X��'�����'��	u��h�Sy�,��y�?� "K	�+���7���^���\�!�@>�~*�X��C�P��81AD�� 6G$�f>���B���e`��Iܞ%AsT�b�G����{�u�R�b0�Kz�fr�!�뚍�Dۑ ^����m��]�-��������H!@1�N�;�JR.�� �I��`��Y�`Z�"M��#D�x�>W}��/-l�ɳu5l � XH��G[�-�{���pk̛S
�u����T}��2�
�
~��
s,E~\6���DG�؂d�i��5�{�H Q��?p��8�7�dT	�ٵN�W�89���v=���6�CYUj�d��B���"�GjU:���3�Z�,-`_ш����i�0vw�@�Q�������"8، �1w.��9�EkT(2�&�s��J8�ǺWg*'���S?c�Z�^/�	 U�އ��:��ˡ�ˀ�S�\ߞl�C�(N��5!��=@��P�A6��H���ѷԪm��O��[�I{�L�*	
W�t�;��<B�^�s��i��6h�{n�>�T�4_��P&~��[@�&��� cdO�fC8 ��}���xd����n�,� Vh�f(���%�z�����c�����<��|混f&a���I"֠�LM���轠F���bBԴ�����f�.�� ���>�#��T���&P�-<^[U�
�e��3vT�F�7�BeFJ��tt�.1B�x*�ÉΦI�Ҫ����D��g�f��YqݺO�^�]�O�1(���W�j$Q����&
s'@9�N&���#�	Ʒ�`��\��U��ej�ݍf��	AD}�F�ת����OW}}�3![CЗ*a��kw��9!�O/��y�<k~{��vLu��`�i/�e�WО�ڰ)���P�/�d�S��é�<Ț�"�q�cixԒ�n�0PW
C��_L͏�.��h��_�GW��}M~��7{���6��%��.��p��]�暑msv�SP>f���&�ƾ���`���Ī�������.��M����V��{R�$�D���'0o�)��x`j��`������'Ii�'w�bQ�%S��t�BW�Oh�v��/���]d�?�3.�'Ѹ�VHh�#���v�� u�_|���`�T����:��fS�Ռ%������x�E�GY���"�le���C�.U�փ!���9����ls.9���	Rכ��ms\/�a+�����Ʊc�Vl� i.���:3����;��ۅ�D�%εz�[����i�Z� 0�ê�p�<5-����)Ty}O� fX����
�9�[�)f�O!����@���`��I��rED�Į��;��񵲁�mB��dű�8���������{�H6E}rZ5�0���������ë�A�d��A��w��>��p-(e�dU�%Ϛ�wAS�Zcj,��y�|��qN���������!�R��5�%�/01��*t;:�>]ؑ��,ig&`�jN=�/ ��΋,Ҭ����M��W�Gަܐ7@=K�c��$O"���:?l����8���ٜͩ�MFʻ���%<]��;E�.9Dk)g���y渰�L���uH�UNq�L�]팼�oe����ٵ�@t���?�Iǐ���a��wB��7`�J�2��9a l��o/ ��X	h�^��SӮ8O3�8M0)��!�Ϙ��;sr*�����˴@�X��'^��Z��ŕMF��M�p�$۳Q1���5)��j��ˌL���xu�j���HW??�A�}nZF�\͍הGըe�b�dQϼ�G���O��i��\�F�2pr[��[�����!L���b5��k'B��g6�j�H[��: ;���]��
��3ozD�{rH��܏�3��̬%� Yʻ)@�?�9_;I����,J�"E���١hm���A�΁ Ym��:1C+Æ�ٶ��t�Sk�qohflx%in�2u�%�M�<� ��%}���خT��,��\kr�SB
c3=��� ��o�3��q:������4�?Fht��~	Y��n����PN��[ySf�b�[.+R�-���L0]P83���޲���+���g[��H�X%l;0��m�/�$$����N�H���{��\�pb��~�2_ؔ����-S���:�jkK�n�G(�'ϻ��������E�'@G}����GR��ϕ�.��J�xQX)��:��R���`y]_0�������M_�%!�4j{
bkP�
�梨�;V(^��`x����9�5��_ܖ�϶<�]sk���v*:�3Nj7��

H���;L1��H����&#��T��'bcq�E�2P�<����]��Y���+�P�⌠�Լd��r

���O����{ղ��F�!�>�T{�a$��?�O��Ȝ���B���|��d#����$t�ͺ�6Q�]݃HIS] ��|6F���V�8�6�#�����|����A	�O^�������'[�lS�����W�/��#������$���?�v��ќx6.%�5��T�i���NF�s���~󺽌޳q��@���6�$A;`�Ծ��H{���'��t�KP�!~v���G2���Te�P��s��?�!F8���bcP���̆٪��}s�)���îֆSe_��/�M=~��gԐ� ��N���ۅP�[�*��8��*0��C2�0��빚
����Qc�do�j���_���7��"Z,җ�����J�.���Y�l���d�G������(��Y`k|���Ӿ$�t�\w��Q`SVP�BGQ�%M�,gv��VT�M�%��k6�zw��D�^� B�Ίs+a�4�	�Y7�k�kM$��R��K��:N e��p� �."h�rnH�c~R�oD��ZV��J+l5��p�eL�%t���x��Q�����Wɉ!�*n�����V�K�V�}	�O����-�_�/�f�Jn���~�%�<f�V��I-T�tL��oנ��p�v�ϭϡV���č�C��Nh�$�>���
�I؀��B{�#�FҪ%�m�M	�̂���U�t��^�U��� YM�!^H��CA�����$O�2^&��v���>������lO�f<#�8�w$��W�� kU�M�tWV�F�5�1�ׅ�o'T}B��nlt~�����>B�l.E�_}^�E���O� ���I��w���;t����XI�k��W��l��P���F�:�@�v�_����%փc8�V���[g��s7�ަ�ch��nG� o�X&���ͽ�Ռ�e'#�f���1������7�k�v�D5)�q�>Hڮ�z#gJ7z-��c9ߏ�/��>� �vl�ym���J��s��%�ڿ�M����P�e��i*�u;�b�o��e`(b�o�D6&ڮ��&����Z	���u;�6�'�yi�d�x��{�ҿ$�@rZHFkK%����~�_g;>y��K��J�JF�~��.�T������J�C�W�k�m��&t��]l��O*5��#Y�D�&�Y��<-�-��πcۈ���!vȷ#5ȃ�2F�M�(ϗ�m�E�N�f�����ɬxS�D�j���r���Zo����Z���2`��Ɠ�Y�c?^�=�.��Z���r�L�m��c�ZJ�؄�p�.NZ>���I[P�f�ՠ��/��r�{�-W�E�A�>H��"��B�ζcc>6�ꢸ`1��� ~��L�e�4ɾ�z��[��:7�h���m
3�;��yp��ӈ������.'$��f�s<��H�}�`]?c8���a����G%4՜��aq�z�xT�*d�|DP�A���\�E׳�4��:��e}z7���j�,�5����i�s	:y~4����*�)�KD�)n��8C>C2���,읉�*��4��(��]]�$�?��L����W�:S��j�3�4H{w�c�/i��4f�hf*��Ԫ�`,�� A��՛2�N��4�|�����#[~�v��P�wZ���/U(�	,̫"N��w����r��Y��b*���r�AB�=Ţ^~
}�����/�ȃ�6{��;�����kP�m4��ե ��'��`�۷eH�Q� ��zdDΎv�� E�yu5\te1��jރ�Y�FI����|�4�+0?<��P���iO����Q{9�+�d�������ϔ	�%jߛA�X��7F�e��{���^NᅦP���pḰ�hZ��f�����"�(�<�N�.��Ѿ�3�uOC�t��=����VF�����"{��<��l�e��c&�Fw����;���
��)r4�)�ֶ��*����([N��"�!��~K��:�څ�+K�Y9Q���>�c&kJ�t,$d���$p$�?_9����=�b��I��)�L�::T��ᴱk��M�a_�P*^�`ش��J}W��;"=�.���Y\^<j���a)��%�pG��#�)ŧB5 *P�&~d��1��0�ٖ�'�d��{?��3k�y��.������w���e>��E��SLY%�(���c���b͚���W$��#��x�D��<��1،gq������ x�-MQ#�B�٥��Z�I��=&!��
�h��[���bɗ�P8�V����M"�+���D��g���5&8ۧS�����ʏ�����àS��0�ؾv�ތ�.w��`YuC��a?���ٰ��!gQɨRa1�N2�2�7zua�����l5����D������4�a�{4�~�5R8P�y���#1ʱ�Ffn�Ҝ�����uLJ�N��.���O��>Vn���*ho]�q�x'�A�e��kdA¯[8bS� �[�(D�C$�9���,�����M;'�7F쁠�S� w��O����L�J?[��n�px����EBԐҟ����.�Qv�$}���`KDn�p"Hz�מ~�;UX���ݱ����1OU�,�k�iMJlDT�=�{��r�W?R����p3�E���{H��:H���+��uy~.h��!\��'�G�UǧI׻�'������'�w�{cd.D�غ	,��t���WN.�
[:5�b���J3�5E��h�k��)jCJDÛ��t/��V!*41r�,ap; ®Pu\�W��C�o���k�::�*t@��}���7��|}Ŧ�b=]tztll!3���M���U�8����3��-B���� ��)�q}�K)Ys#]������a ��o�_���������LR��7#J��^��}����%�Q?�ɾI��jܧ|��B�Nsg�gط���������XW��]���uZz�Z�N��Y�lLi� H���lR��>��W�է}2���d�;Q~Y��5W�����6,��71�B��v�N�n/i�Ö��%��p�^Z�F���:7vqM��V���X�$2�z[�_=.�V�佾<�骻��ҏ+e�<-B���9�b�B�ٓ�u3�}�H:3}
����
0�28o�="��&Ɠ��p��u�W����톸��́�R����٧O¯!���$&����,](hz�GҌ���������KH�t�J�����'�PhC��mt��+�l�ǭ� ��!A�Vsi��혵^W����r���9���1�#��h����`g]�$+��V�?R"����N/�kFn�d)~P1 � �\)Hw;ru:kK���s��O͓X�ނ�h���l�_\P��,]$��:Ы��P�"s��Q���jh���y(u'�l��^��� Sq��-)�]��\��\2}�{��u!"|䒭Q����ἦQo��?1�H���g�	b�>eb��u�?�Ȕ8|��ߠ`��2k�m��8#��<[0!0����GU�J���n�R��1l���HV�T":Kɘ��6�(ǟtgP�+��O@B�s�	oV�A�C��a��k6�+Do-Һ6h�9d���z/��<�V����ũ��ʱ�P��P`�r�r���3d2Q�)�I���l���5�Dj�����e�� pW�˰�>��/�*!g�5v��@J:j�Dn#d-��ME^oa% �y��S�QAl�6��C��~�uk��(�ͅT4��e5���Q�
����GBT���6GZk{����gS0�.��ϯ�����H�βj`)�A�+f�d2f��P����˾[8G�e���w���m�!�w_��
P]w㕿M�ԜT�2������ۅ)�2	S볕�?7��ę+�.��ܤ�U-��*Ɯ�w�md���!\2R2�h/F��NprK�Gizi#ͥ�A�8ۭSdD�@�,W�I��Z~ZH��x��/Wqh�7��yKQ��	<\C����A�`�I9O59���	]SM�˪��B$R��p �R�8��-(�t���e��*oķ�Y���k�v����4(3���ڨ�ƴ(A�N&AK����>�􊤂�=���J?xM�%F��|�'!�vw�]YY������=0k�9�S_�����,q$�A�d%G]<��ßL�����I\�-t0po��6���K��^d!�E�V����t�����a���s��M�nH����D����f�F�t���Q�����g{�$eW`��G ���N��@Q~�����s'�m��9s�6ߢX��y�� Is*w��;��|���P^�u�q��kK���y�CT������Ђ�H &`L�
�4�y���:Rٷ=��(����L`�[I�y Y^p_�@o6�!�IT�A��׾��#��R�*��]>�=9	��n eeE�����^od�}ѵ<�w{&� ���=h>|���|��yU1�N����*�g(y����i�J7J�B��`�a��������Y���Xjᆥ ��O�G=�!B<b޿	
~������J8�l��#�a@i�p��,w`���*��ˆE8	�.�걩�h��_3������-�ں[�q���Y��b�<�V��xY)��$d|�w!�V�W������ǉ�z��{32���/$6�}"g]B:U���f�K�Z�æ���Rpf�4�1F��"<+c2g<^Ē����/�Ap�ڋ/�
S[RX����JD&��Z�_B��( ��Gr�[��w�Ӎ"�����ڑ��b�A�|�{M��J�W)��lF;#E|�im,$4{�Vs|�'�j/��,i ��3�ʶ���Ud�
u������aR�b'�-q;d�g�������3N�O��W��Aӯaې�+Z�6��X���aS���U��E'��;��?�$��� ��{�ɞ,��` ��C�2䚲��幽�k�g�2���L���6�� �1��}�b��#��x�!��eXs���̬� ޳�;�鴘��d�$��ށ�8ww����Kx�iG���*`��!�$���hu]��������:�U�z�OA�i$|�'	�WwSW�����;�H�<W��Ĝ	�����)����2R�>��s��}�
F9#�wr����\� (����V�Ű������ϐsI���5��2dU����� �۲"��fJ)��K+�u���	��-<�ʏ�עt1��������#e���F�V��~��V�!M!�Ҹ`0H��&v�T� ^2���^���q�����	������뎑��<�����s�0f�_;'%��'�`ڎݪ��y�*�Q�ޒّ�y6�.PER��RM�CM7+䁕�]�cX�.��h��@������e����a�0	L[�F��lĀ�@>�Lx}�-w�S?�s�C.�u-���("���T
�����0uD�w���P�G���v�%]9�������S�p��14���뷳���H�p�>'��0|��/�kؔ%Ԥ�_7�%ڊ	}g(yK�Nn�nU/l�ig�F��)�&�d[=����xLh�h��eV��M��Ȣ}ݰ��i��Z��Di��Yg^���_@�Xё��nx/�F��D�t�5~���1��葷(�����QA���<����(�m�Q��\��N�x�����a�J�k�Lb!-��\z���Η���#��/�(��|M�ǁ���Zz4��6!���˳Y%�i�����́_�s�����8��K�
�����%�u���8�r{�D�%�QT��hۨŷ[�zQT���=Ɵ�����M���]�8���
UH���>�����k���v��*q-X��ȩ����S��Ə��;qI�F�e�_��^�I���]��d0�����e>�N;��yi׬��W��`��V�)[�T�K!�<5I�j�%Q}��o����@ܹ$(�]p�c
@*�4/�&��]zOXqM�|+��bp��Cҕ�p!!��yV$�a��u,�q
с�$����e[�����m�2����w��"5��#N�d�XJ�-Nφ.���y�Zr�=���R���5'��u,L�O��lÐ��7؂��	i�q"���VUe�v�~�4�b�C�C��9�`��}On?�!@i�v���b���s�|�]��M>�Ֆ��u�U�W4˘�1
��u����;���u,����0�ƒ�[,��c0��WxfU�ZF��ߵo(���hab�OL#��#NO�׸��r+b~��r�M���0SA��Qe��k����8"�v��<������������RG��9ۣ+(!��nr~�"