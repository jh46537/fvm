��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�/�CZ�08Kh�� ry�z����������B��N��VoV�	m��^/EW�ל��!��YF�gC�$�Z�e��d�aEyx��K��T�[#�,<]�\�V��V��a�]k�W���&4K��ho�$2'������	�0̈́6�� �t�_�w
 ���0�-Iȁ�id=v]H�f�/�i�*�ߩ�}�_,BR.� $��h��k`Z��Q�C�$��J�pu>Pg�`�!֯!ҦBW�W�������~��S|~�ꋬ�`4li�~܁��3�>�(]Ͻ�on�yQ�����@l8KEr7�}����{�x�����pCvc�hf&4q�0��z��m(�0BK�G�<�������C��4��G�M�u_FC�F����Z��LV�{k��rƕLvA}|M-M�~������-�-{ӱ��p�t��u0�	]�jrW����'l��l��&�
�����P����^��j	��X�,f��ziU�|���n��8�Ȼ���,ø�r��A�,y����c�Gb:�����>�= 6�u;�O�K,�ؒ�A0u�{aL�j`7�_�f���N��Q�,��<��un�D!#���kf\��l;I��-L�|^�R;�i;���m��b�	c�H���c��=���1>���,�q�B���S��N?-�Hl��3��]o�;G��uR�=;�S	��
�e���D�����R��Hs���j������-���O�$�}��'��
�DW���4�+�K��y���o�)m�Y�fU)�>�A8�,��~N������*p�7A=�%�fB�Y���kLaA��9�XY�_$�4�<f��8~n��6q#��Y� �g�x͋�6󯋭�PP�HG���
N���R���=Xy��b��j�j]OQAtzДc�Ӥ�ÕiA�CSd.�kr�: I��?뇅��Z��;�Y�C;=<��F�L:�w ���'�P�� @�y�|�e�1j�Wio�D�ShxC՞ڏA�

�{�����<v���.�W��i��;�m�P�j�t�(� U?qIT�{ء��?��U'o�%RH��3�K���4=�#�>�*\�<7;O�������	�������~��.&�@����Ov��oxY�
�I�[7ht��f%��Y�j�
�d�[7��r�\�,������U
�����[8������l�2��r >���/���J�cCf��}h�(rX|�����x-xz��2m9���m�lhH�K{8Y������y��o�dmQ3?�u���g{�3fe�.%�b�X���>�R��c���<��w���(N ���][Oc�7��}	���KEH��'���[-Ɩx�R}AmG�h>���!������� ���y�i\���Gܘ8��jX#�(���+���g�@V@R�Dp�@��t錓��̅�<d�I���2�����p&��7C��И�\��L��CZ�X~��I�x(F�k��&�L}n�Je�Ky�E�wB-III�I�~�Y);��ជ�D�	�	�܌_�Ӣ��X^$Y��
2�W����_�TZF8"�\�����s�W��-޾��U`�[,҉��x��3Z3�r|O�pWa�/,��7���3]עl���k�F�|TJh��+ȁĬ��&�+N6:,�a�0-�p��UG�?�����hZ�}V�Y?!/c��<%�؛7��ИQ�[��,�I�X_�#�P�T�ln�z�&�S��g)WyD/��%W�l����v��^x1%�v��h� .�3��t���Ȼ�(�+`zȫ�?>B!,�J'�m�7��t�ٲ����	��]u���
o�;��� b�#A���:�ǈ�_�2�JH-���B�*
C'6���1a��N�lR;p�l�r��̐��ߑ�N=�Q���8-��v'�Yzrí�*�9E
 �=.��aqσ�e��L����|��Wv�5�i���PD~)Z�w�|�q,pե����wR�F�5����{������k�xG�L[�ߏ]Y�?���K�f/;��`��r��E�L���C�ܚ�a�JvW/���c����,٭FOU���r�+@P��v��$��ɝv��{�L�A�5� �nG��.��t��#]Fێ(���T