// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UankhW5XONSEfcLkXirfa6wxwAor0c11PwF6TBjTeF2oyYBOT5mMMF3B/CfTusAt
Pe3WnW6AcIy4dxme6a5cbEj75xHLnhv6L5Gha18x3zbhOPnRrZjsVjpqVJ0UJ+Zv
aqBPn66QPnCe35VYO6FtXfHCWzSAC9T1w63HuAM1tUA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33888)
guAmccqfGBarXBcKbDg7oSLmtxDADFZlQaeOT2TdSOeRXo6eHFDuu1cCNT/36nAK
FBeb3peubOBnvlRamjGVU6DRj2nEXsScOOxevRrvbYwXwUBy8ozcqcU/e4nfSK8+
p/ArmWYhjlG1U2u7fwUTgX4qPM/3ZyS8DhYUdTawPNU95/upnGXdIBuuA+fzbllQ
6+I6C6TfrMWwSg50sYNoFzbrr8orgOnidLm69zVxNDlKpIeZKsXbe6H97A3jMVp2
hKT05tM6T20JIps7bjDaiS8+j+0LtN523P24fJnktJ2YJwmwJDGqQpjQHJz3FWyN
RlwDlxy2C7GDnWwGmHv187nv+17jF7ZanGkBOvLm9AEdLtAR9CLymj9IBl5UhbEP
Jge7pwTLw5ybzjRzr1bQidVSb2Nu2azI1kYZRPCdzdkbe0fFg6UyOyT6mmIs5tkg
ZrVppdM4iRJQeChCpXu8VPVJtQ1Zlg0TsWsqib6EsHsdgXT99HzjYuO9LMhdwI9l
s03AUxNJ961Kh74uezcjh3gQFNjx0gD4UU5U0p48txXnWzbdy++EvcKDGSX9blVE
DVEd6z0BJdXFBuIzRnsZ5vvDC8nyxwDR4noY/C6X0AGJQLOAxngtx+H++7Bvx4yP
o7Fz0mizruxSPpcJYWNdH0kq4tcrcbaFy6HgxroKV9DkeCt3Slw8v8ePn6i+lFmm
mqH5kU4ISBts/h9GfCCMuP6gvEgqmJZoros1IDT+kv9pZj9mV26lKrTpaAJuTcuv
BDyUTpOtGFhToxkack9tsBqvFqk+M6vSvYJuuIR+xorHa7o6T5A1NIIlbv3Y85qB
dK1HAiXXt5ANXFvqzH2qJTc1FLFeHajXZYOVgcSB79AFCeWOCJFW3bVaCpvIFG9o
63NCzTwVRZYr4W/nm1q2oyPHwpNvDHuBTazGbAXtd9NJjjDKIVEmIYkJoKJvyr0q
6t0Q8n9Y3mZX5KeX3upGcDXspWt3KyKNJ5q4x3uhhqBlQgdJ+Fwzl/ivD09WxvUY
YnM/MKX2Rb5QLnFc9/YYB3UZsmhaOpvOmwy1LBypbpo9t+YCMEeUxhst2ESwYVW7
SMlsFjDEEM31kfmtLnHq8rwOZ+MKya16BcpNlPpu+v9TUsQd3IIMceUwbnmmF/+S
5zHeMDzcgFIo0nWAeMxbSrI0Y4UBwQMQgyE4uXXl9M0RNaLWH16CIEWakEMwVZC8
Mwa69Cgc45J6up9jvfePK9eQyKvSbXlCs8I9eb9sgBSWMNWjzBz0QhQ0j5zs3wEP
7EyPlHK2RX5Sd3shcG7Ic9MsxCW5jqMHzD/I366I2tDks8u0n0w/PvkNpSYrCZNM
Z3SeD6d28/nM/IXl0P9hEpkeea9we3FllSGnEvWtv31zBt4wLmzXl2D4djUnggAh
USN66tILOjMNkhsH5219mtCZUiyBJGm33poqqr1lokzcvjxb61QUOY3CTj2nGM2+
YN/uESl+NbFwuF7U03rM/Tx6kDtCIPZ439Yg5uGzqlgH25MA99s+3yCZEDw6vhfL
+tObw4gsiPYiXCdiacttBRXzHuNoDXDmUwnK9/Pi2uT1m7FrdUYn28Y1e1pMt/6f
9B9lRgTGr34WjvOKBS22F+iJr/wnktm324sVmo7NRUuY2BHScrPrFt0fZ5IVfLqF
sHJGLUm6F0a0smM7fNThvEi4fK/zjQYX6Ag477yeJUZMYo1cah41fKPftMjlkYoS
uItZQiWzePj8DNtlq/lYWsEUpO5XSZbJWMNjNNwSIgR7QwqGPGilgqkg8Q5XAo28
0CUSim1mI1478cJb77iD63F9lPe3WMqrc0pExoCweb7PoGVPyjLF2lfFJyIft18E
YPydL7q82hSUqSKTH27xNL3CIE6OP3qzS0rPYRB0K7E+FdTLTBZ/Dng5NQy/y3pL
3QwWQPASnvn+PvIGngT34as/Kfvz3zL4tuKMWAf/Y1UMjsZhzSEEz31WoP+io7my
cMJ53+DLSmV7cd384lQJ2IfNj7qqWAXfkZ51TVrDpKeMEZI1G8CZDyd13aKi89Kg
+SCA5HJSFn2+JyxF/lmMxTxKYm8x4W3KRSnIreGp5KOUccG+ObhA38T+dBQmJ0ep
UnUt/swf7u7leJWzBW7lBHBQCf/ZoiSLlWoY4MINWDl7KLrbMYwBoGQIjNuSoznq
siGk6NqVDD1Zd8eaObyKPRoSkfACW7rFUiGvDccZHaYtC/KRLgjrF049gStieDqY
CFNgtskbhx/Y97clvUeVNdknb2p47Po3RvSvLPuP9mNDen/X9/pCnA8Jj7Xb/KXC
uNSwYd2nr7zCgS+dH/SYgM7TvAGjfjSxAWCsYbD0Fy5K1CNCpRMdO2ejxnauBDCm
36pkYtsvIuKdcDnOi6Zr6jJV8PAlrrxvA5o0RIpTea1aUDgw5XhVIWP32JfJm9Ui
jX58ZmE+YixlVYzhsBtDC7VUS8YavgW4MsR3B1eEo0nw77xP4FS9Ahjez4UujR/i
anwG2bxTAG6Q1I7xwb8HOfj29aDKOTrD2m3LsLSOvlZO3aadDq05ISdO/L2kWFJQ
vgfOl3Upwu9Ee5l5kb56iDD8PrNblKIU8SOI5UcEhmoY+Iw2THe9BNFNZsNrp8Zu
ekVI0i63GPgXxuP1b1rey4miSAn55JXdCMCQ9uhTjD+w2tJoiM4NMCOxZ5HlJ0eG
sR5ztIY3vd44WASYWTswtcHIUe6XF5pof6D+8v/j3Z/i7rXcX6SdaYCrFmBcXD6E
qi1Y3USWt6S6WRbJ/av9LxypaRujmkmyTpZChGfIAWosie+0vun0/DioLSA4Zmh4
T6tlBKSxSHVmSnkAhpd0ZnRJRegJdp+DzDIPSOyoDHbrHtsbYAm+ocwUmoddTE8X
5dq3yJAUn1uoBXw0kkybNWQsiqpJOdAUopui5W5dHv6OKbeay88AnEjUERQJUVPb
vEJqqIIPBa4ifm2CV3HwZMB3DcUdR3340RgFSqJqg57DoKYdpcpwCASEOmSqm1WJ
4gRrzzISP73Y70BYD8Yu7TEQCjgibV8mJHEqPZHNiYUbpN/h8p/RakyOSCz7s98W
PGKlza6BARyZrSZ3m/yf0U7dFR3I6k7WujFDn363Ybwyy8T1NdjL6963x5mn1wSr
iMtEnOdaGA0cDu2P/dJ9EgQnDKGTs216bD+IhcpQLHuiF4l20tXurRSR/boF+PGC
/uJOelpfq+D+pFLwPX2Ql7xtaUHhgDsbuUrlgIIztxmIoNOXz9qLw/Ro7ZjCFkYh
ozNzDsTBQXa6A3NhMP/2Djy6hBo7r/DN1oQOFA3faROZcIbRxLmF9xknR+8aWR2m
8gVOFJZvVTpjbKV9h8AvgXg5i2eYkjWA5dJwAKHWro9a/8c1+6Ct343CzKHtAbfC
Wru3nItSvy8Jp+pNe3XaikIQibVaXLfKiGK/W/e2eVFf/Wx25KaLKvhz5qxWaDzD
S4tUsR2YH+JFLMWGFf7G3q34JcIiUsHi8BnYpOP7Q+CMH9QbZMi5/2aOI7/UjdgJ
CG5v4NGNytj4Ir9QhlsCSNJab4YOn838wp5L2ug0BCWK08xtcCJ8T2dGKSNgSwhQ
XDzJpH8iPPPEyjrqA3pKYxikcSZBwf+kvMRB9iwiWK4bYCRiWV7sZQWjX/rIH0NN
d+GjXvBKNdJIObrhEMPKK6C+84ReZylhVTJGixVmXfyHybQbm95hf6rGgUtD0pqs
6QFlb3ygEyRJNMtoErL23KL0YABaMMSSPNju3hAvBjb/sR1LkpWg2Oj3Py0c952N
ygWZA45q8c+3bMULZDeypRXcwgvtrSTjOcfUSR02NRnl0j6DCGq4dVCkbSAXuSHB
+6qdxTOlueA/9sdyOjDCzC7P2j6bWy2fTBhvT6WbErQoWd+lBGqEmx5eA6bSsVa/
ihvqbd99PMeo5zShnU0lY4MpyTADwrp00ZJPJNjVcIU/fgQQMUU5TfU6n4kr2OyM
d04aLwTe/WPrGMu2gdH3Q9Em9VGi3toY40ws4oviYGc/3kuJ42OHfUk8gmfjXZ3g
64zWBxy1lu38i4p+WBB2G/9qUx95Q578RhBr/zjtF5WcVtFPWCJh0OaTMk3dwj0M
kxG4y5ls05ue+7Adr2zZ3vG0611gYDGDVWbiK7A53z701v4IY2EaV6q99NaEPO/z
+JifJNZ0qIJcOWAU6VafVcWWpCE4rBsFfZz7TGPEni/Eyr8pHP45VrqLORiiknGV
AfXKMxaGn4Emw+daj38GxIUfAM8rH3LkOjm0MMUwq5OurXSUbyU+uXGWOi023Hwa
zX/KI0UpYkPJQbRqpTfTopEbnXg3IHUGhjzAS/HAgDAErYNw+tNO4uEXlKE0FilZ
ANiQeQJZSogKCnMCG4nqVH3LoJwfj+9d4+8Q9CHEocq/iWzav6UsKeaAJd+t+I+7
e3wpAB0pcPSQArWFPdkm88t1oofuInShfvzlgCWhw9s7e0VVNax+wD3fK0WF/Jpq
1kSE6KQ7c2gY1sTcA5EjANzwMjwG4u1NNiopmhSP3DsWqZe8WQ700qXPVD1FGIbH
ie6AeBTwt1NGqRqzbrxtC6FSjdzD+FLANE8wYBpPG4CvBkzOIyKjqe8PUau4+AbT
kh7Ruv+6J91sVB8zuI7GtaAjvF3Apw5bs9SQm3ZqZsKeJvhc218iVtBt64tq2V+B
y0qopKZqU+ekJCmVXHpAIud26n/j4rGXnt50KCxuFks8FE30qqY00KpWE2LsJWiX
fvkNW2cfMlQqaiplIObFflo6aFgpejmdAQQUuBiJKnmN1TKDP3j7RtOQxqlXh4nP
WBgzTv299ERbYPBzlT1LYEs0tliAgzXatd5dY9RpKZLWWKNQRbslXnUCsdcsxyo0
wBXW+myl42Qitm6fNluC/cqmUeFRsV8LWFoECPk9RRT4gx1mm4kcDPf7JS8RQh15
RuZW0V2tc6ysFcoDx1gWC38D38vs8d72HrwdhcUKn7oWYNh/1cOX+Fr8hc2xqalW
aPYhlFOkBaJ34X1nzi8R9UNMYvU9yPPFXQ+e3NA9vmrzWsZIn5LfhBz5MM+oYvqy
k2QblLXJyaHNz6eUqlFwnqCfM+6Jz3v7fVDrC0Zm/N0L/ZE42p0991+6wFRUyZ7t
l5T5XWdyUJzs/w4Husg927fe827tBwwyvWmxhqPr9AXLoMp7TKKTGB5kd5DLPIqc
hC3WXtZOHDbk2Md6eE9pWA49pWJ7UP5zxvnwsDk698EnFtKgvBXz8NDbhcVWJtXt
HA5acFSfak2hPpzG3mqLfNmVefZwrsb8ZOqhbgEQBZ5FbAHh6kDNikEw5MpJJO7N
MUY8O5HrOJN7OUlZriWjfnHyqoRm6vuDwSsj4RJVbBFgIMDBY6qOyYe4t4Sxyr8k
ccGjF/65dg8YuczXSRxy33DQto9knvjmRZvan3Ic66nHcQr89lcDH5Dw2yFaiKww
0wOfTlbpxeUJ5mB8tJ2d+AfxpzHWSD88ev8vcv7ilsf1Q6lDmh3rpW3mJgkMlkyC
98lIwRy7zwUA9Vo57juzLCC+xBHLVKzdTUr6M5fNg6SKwtdx8OQgsl8PxoZ0JjS1
UpRBvMU9e++EKUWHdltN94mfj965oLbuBwGv3Xpqtf331V0oa20dLixhv06FLCby
f83Yw03G1TJ/IS5kT7RvxWoQBfIQH/zapa84Kq2+f5+zTj5gP1MyazrwiXz6h2Gx
kFauReFpGiwEh0cKWOl0Gp4JldOPJKGBTAhSEGrSItU/b0XiH1P9vcU/TYCI8mxR
K7va6sPi9gYSjufA63T9DMAH0OG+IH4tUfmzs9Nc09OcmzpQ8THBxeaKhq8u7lg1
JqDX0ijOiGsFqXgRdpuh/SgYPH7HUxcIPfTlgAF8mAVdZAsflsm6Lv1hexYoHmMw
/boeg3qBjvtOw8sPROGTyBT57NGt0XA5bVJ5SGDy4b97p4QkX9LcnFuIBc3atx+r
3gl89QLLN49DU+xzAAWazGeMnsUlv9xtYg+ijsvKYfF3PlnoTykb4KkWsHDOpYe5
R2/eR7/QGlBIYYre/CwNNtEoTbMm2VQDOgnfq5OawgyJ9t8iaYPTZDhmJZsS3FIj
Eu6Yuv4NeXm9es6UvvUtLWR799AEpYH/P88aVnEA3g/3uWi657lmbu/CJuCzIF2W
DUrPApnIz8PhFqX0xr/JY1kBCWXqtBHG5ZADjMMrahz3NTrjnsqsQirtK5Ik4mvC
+lXslO34JabsK1yDp2sMnebDoGuXW0hVvbtIMoUJ+xsN91uvKxdY+Ws8LABxzMir
z8LYJRoH4Pbnwr2tbXWUgy4SlLgBPVWPntOYJvUGhbROu8zadTziu9y+oa6o514y
KiIgWgAOpTkNQ2GI37+q9VEgUSuj2kePtKsR6DuT1qmu5M5PDuTCIP7azdH3M6Gl
Q2IoULkNYzKApRdHspRpwimLSjWipyV10Ms4ak65ejChFYFaB3jh6fzGSgmZHQdZ
RC1Jy/QVqC2MpkjcfIX8mX8Ms/DFiBNnX/0g235DCT2ez8VzEyyBiPmdoFIugx2Q
DhOlMSwRtbG1OpCpfBJfeTGpyQceSfzOYYtLwhYH2Fhw1eyH7pAN4J9XOvNn83Hz
segk5m2888Wpgc4uF5NubjihqgYnYfjQNMEVxo0BDfadOllAO44+NiJ5+D1D99bd
WWlJvzKN5WaBsfz2gxx8Wmuy+jH6OlTcKeeibt9Ed74o/8mLC6zUGPa8kUl1kIoh
OumarZrqoW+xweph5pltPp5FdwEo4Xprun5knJg4r+B/DH7Lhm8amCVdIiZl/KXA
vcp1IDqonGQcbz2Tqa/fUBJo0xhN6UkYlR56pUQJ3L8tJ02EV0vobEACmtUdH6Pm
Yf3QUEVPngKJnQjdo/l5O97dv+hkSW6g2JcA7dRtUrHgqE6GgEPKzMmtBwrN0HXO
IR33CgtWDxqpkk9+wdQA1emYUiZAm2ae1Udx/L+FNOr4OQdK5M/SJHKrHjyF5tdT
ovlTE0DOVHgd/Ii8SW2vCmuKF/svhrbuIWcWiVQat7CnrSjGEvmcnZUiBRiiS6Rq
TGhrqeKC6AzHuRh+sjeMHMD8JXD+q7qe9339p1V1vJOH45R9jj5h2nnqtAUmCBeU
UqvbornI3sKBuLSwbBs7cvK5ExrjprEs3M/ULo6YAO4HqlVeFULsHtBEIAVyQjsk
PP/kdRyPa94Bo4stTZi2G4+DZjOFJWUQ0ykuX8Z/kkcv1aGyqBppYYb3GUGa4ONN
/T6MSKI9Z2bLKDbu2zHpMv2VuHlIlXzUdlni1GQRxBBQTQg4UEWQCec/tA+IK7Ec
MLzEkbSzwVW4BZ/YIkRC6ZfQUlx4wDCBd+G+IUtK7ZaBo+jpj39a50FJpX1bYbYQ
fkGBmtFE7B/gCGNnu56Xqi8L1qk565BOTrKAQja0vXQ3urtp/k84kdBGth+bdVYO
YXJ8yeMCbgl+KUxJwy10Dmds6I+fACFaNVXLkeMmLrLDwrgUV0OMNtv9pRaarZQH
idd92WLe9JGghzXoUwDZj768A880ZnIEUHHGANbJR8nH/m5n7baUYNZMT/X/OsMV
7QhxMmKxuGtzM7+gqcL3/H2aOeMGTL8+ScCati/5RUf5987ZmWkoX8bC8klzshmw
q200QI0AWr4uqTwOx17UthUKiMgyEJFpydxUsQNj/pwkS0DJu4BqWyhtFaPothD0
evGHARvDnZ1WfXNPvk2UUg9n2DflMnFrRcDhbaxlmYgW0F/RLWsDNmF1XBvf2TUG
qX6hDRGEU9bexgFLh08mNQ9IVJAA1ePNJsIS++uk9pgfHAFAkhzTRW2zqLaa6B8P
goX8/z8mRjKtv7EpZOHh+9OKlVkFbaLW3Lp51Ao/RPdz9oYdbrFPxxMI3fmfjqGy
VWBc5tXxg3m+fDK24vGpr0e82I0OpnOZRMhzkDCIHZIqF4reNs+vP7CatJzoNPnV
jPFF0Nzc1VLYD7dHbLb4ktikvq+QsvNYPxtFTc0HDWJ4JQYMevbXf++PlvmntbsW
+hDtt79+guApAGcvk0V2/on6YzIVY14ZHbktftsRwomKntoA4v2HjfObrvnvY9XZ
IRokl2FR11LZ0MRdb8pGtGrMBq2HX6t7Q7hOu4eMBg2cpJ60LQEaDcyPsUnWzMMN
3Nqv3Dkd/AkJQPmNTvRx6kcDC4NXbcSqxuA6f1NBqCl8cLqRRH4jWtSNVDjtYxm5
29pL1etNJycTMwJAIV5EnWspJecVRY37D7npH4xNnsK7lCiRT5J2jKTeW0VyrAJV
XvdW14qI4t5uRC8ORDREi6OOpWJ0ZAXiRrlGie0NOs/9hu85PBcADyME8RjcgSfW
5zxqGoBpUSAyr2vNBaibPcXZBFv4o6CQ5lgeVy/hJW2M7zwQvGdb34IgKuB8oh0l
KPsSQ2bmlHeU4Si4ee/legHSnT2jWHZ0w5uRz5KHPBpS9mtW+tUAslSjKWgtyrbJ
Dq3W7ke7LyTVnsLCujZ1LG3rRFgE3kmzXP8SqUTaAePXGfe3JyY8g/qCF6wP5AB8
9MFxdpZKXxp/L6SRgbOLql2eChZ+MyLNtPuIdwSdlXqUTnQZ1fYRWHKKl4YIM8C/
NO0ORPwrZWdRIv+1YtrmjSt/CXFVm+A63m/Tm2LVBk3r7B53fXfcYN5hvfeaOMM6
SzxCueEE2NzyLZSnEIfmErVI/RZtlKnldoeGe+jlg7tgqjb0Cs/CpXzPX1O4VUGR
pDixn2bEUT1CkasuAmtZMoW+BBX/B16+vVBWlKmy5MXwTjtHAzPi6Tgbkk4jr07n
vJw+h6xL/1KNcQTVK7ZoD3BQ4XMbuCWkujUEAoJvk+YRJF12/PB1D/8z14mY5h8Z
sGbXO/XvaTDylRAFW4kIbmE6goIepmDTdJU3waOV78e+prntF1ifl11GMq97ncPo
7wS0LUTYUmVbWpAVj+fZUZbe9vEJeJFS6rdQ1MXX3BtCqQSGAp5LuO2GrhKyEkxo
L/U6zQ6wW5+X8yAk9c6//0ZNYmalRU63wMBBle5Zu26uzzYJJQ3EPjwxEfWeMTlk
ExuSkmc+Y6cfDs9TiJgFLRlavV8eJ04mL8ivPB9v2lYh6e5Pq37FQv47EF4UBKsb
0tjR1ElQz9ciPc6kXHJrV10GZNzU/SlQKuohQMHQxzEwjXkbdpmctqGPJObmfYC0
1hFOV9G0AtuJ3ImyUDwjN/lOUENX0c6x9j2250qCJ1YkJpgf/U05drhkv7JvwNKt
PFwJ8Qdge3S33bNi26HLGKG9d+e1awq3Ch6J4l3HHQBmSfLlJxtIFFOv0gspVHkC
zSTjbfZZjU4zECc9H2LYKFnw+/GTUTY9p99tVxi5PBMkQ7KJ+8Xb+kli7rKZvDik
nPtJ4HnbQ6of5xIkbHuQSQs685pad1jdt/ksoYFl9NGzViBfst6lA587zWRqXVsK
bS5fedc5QikfPIksyLzZ+BR/2V3Sutx9srcfJgOp8ZCuE/OteCI89nKO+UfN4Aab
2X/KxeueAzz7Za0IyPFlN70e59tG3ArB4y0bMqOuLe45jjTnKYvXe/oun60ERAEr
DqjXROnyaLpqnfoEWM7vcfjDi5AjD7wuZ0/yZjDKQNBqoxSNs5+ZyaBwRfBW+hIG
jgEC9HASFbR/3cpYQrhPEpTx5l65l2dXTDKt/vv99XVxZrr8shCDYuG6FUcbQRT9
omfHSGSHyua1MOiqeIUNpC9DOcu3VtExWYbJgn7wt9X9E/Wyj8V87c+BCoNA8ZR5
35HW2Fy/MikP78dShc101/LrQoC6aWE+8vwdAF/afZmdzLcXSNF2VM2mKIzbTZVa
yQtdK91aNBzRQkhy82c43391Cb7b/kdqbxHQDdUN/hAMmyyMI1Gx33PmDHO2QLpq
z2Y2UiCq42SAuc16isMA3apgdo9ogNRmYTBEVHMmhvW/3AwLLfZCGCxrzAQrjTzM
nSioPJYEYK6zoVviCAaY/i4/6l23Xfw8TGUJyiP1fGZjpnGkf959i1VUuFld2nhn
N6y4jXJWxAM9sBYSLWwbUZDyKNVAO7dsyIsDIFGQzDr7lRgf9gmkm7mlzDlld+dA
EsR6XgxtbfclT4gUY5f23O9Vb85UcU0ljXhuuIbzp742bezUdf1PHNLS0t2POCxZ
Hd5V9TZadrOBnS3oriyJzqTBlrRYxMbEIiohsAk1H9YPE06NPE1LCE/hoKOasTn1
n6dowr1SQywkTHPKlwn0KTxvrEMzdICp0ILssmo5v+uBlfoUuGOpRFN0ADVxkcwy
YUK7YkHrd+59WDfDVMH+q/2sB/W4S3Jzbgajd13OBsgvbvXLyFI7eXy+jG2Breir
JsNnhT9+PaTvJI8Y0C6xHue/qPz2/hMFoHDpn/+26q5zVVK38My5M7R+mDCx75XK
DJMY3OgtdTPnQQCP11+FTQiADXJmd9gLxieSJnJsfetVPptQPw38+UIGcqIpJtG2
TB+X2WFgRYffFABvBhc3QUpIYF85jb43A9W2yxwYwfwCn2KcpAkvgnoFa9GxsI3Q
kAA9fb3s0sGBJvooKZFL90lZoOvyo7wzA26bP21Wnky17WZzldDvJ4Q2aU7aCEMp
iKccS2wGZTKZ/0j4tWi6jTLOV+sZNfgz3C+G9imgWw+eavHb2+xb2F5/KTYoBp5Z
OOScCGJIG96UfEh8bAtU7Y3xDdqALsHjDm8A8dS89W5HBY3xDBqRVBOA0ba9rHKE
eZg6grcU6UJg998Jb+BVh5/J//fLP/w+KV4K0259dGZQisis4VASAzRTU85deHSO
H4eLD5PoKjxrQr2kHA6nl3MKJxhLMnGk8RYwrg4vpw5wmpGISbbQaxOk/YlxJ4jR
thusVNQNY/aU0opRHyR8Aue0KYjf3Glc9DolWo4FmbR5b5QisiAUcpGvxPw6/ODP
MlmemwlZEo1XWwX+0TxZVooO+ijUj/voGD12yAE6UKPTEimc7uKQ7/+2nkk/okcv
33tb093gLLspjz1Z2NP+ouVkcTLnIW/EAGLMQeP5zarkATiqQ8kMCuaRRCVCbmae
Ms+CPYKmN9uVsI0umEAWvKrXh7q4NKIhE731oImMcUEYEPgAZ6iNnfnnx/rASHTl
Fx8RkvGmBUYkWY0YBbqU36uzAq3V8obv2lIRT1D8EH25ECBfhWIKW8U78obqIzUu
nPzBL/zOGnXghQZywTjJ6v8eaW6WNf0w1dMYWFxDOIUqPUiCk//x4l43hJIbq7aE
IHwrffkMWKtAXkrXtqDbXxbzBOKCOrDIQNiS4+TppQan6hba4I10vaEcPuBSYHjX
wimWguqmHjFGJhUUJElHSTr3BC7N1mA9FSbz2QK9978JTLxdb4Cu/oQ/XY32kgwu
qVjvInzqscUzwkLweeip6SiU9AAyjovMskelL8NCNIMqZCVxeYDnfoG9I9LXW/f+
m0U6ia4V2w0jJSfw3ys38fB5Boetqa3tYr48WamHUlONv91fTtjXFZb1PM8BueL0
viQ+2RGfspWrUDJjX49wNUaQMHAuEF3kFi4SCWvH7yx6dHaIqJjb6SraD88UwcvK
qcYuO4u/1VPuyH+KHwHHvUnvivHR1qM6sTNs0aOl3hccCEIUPyb7gB5Y5ZJMQlHa
W7mRNn11lFlMK9RQ6wgUQ6PxNsjMpFqZHmfQfmPa04Uohi2c1OnspdSGl/sMqVUy
4wrgeDhi82vFhvJVxoJC0uz3rLVg0w8FXTd07zUMWqESBK2dbV3NXnHSxW/ULnMD
wfWMpvRpBi0AeSWbaJjrQbLvs6UWOqRuLUGQ3x6MQiGZI4rwi2kiBxrUZMRH9esV
lU3o4eYIKGBlR3cf34wx0s+BlqIKgp+hgwrWUTatldLH6rXW/i0hQmsQy5PAkrLL
mUUwCF857zHyUBQ+CC1YcoOTDRvaV72Lh1G6VkxUFCvAZy8IwzHeLJMjxohVT3oi
OsTd8SXR/EvpiTjPJ3UEY2gHgkAyd667NcQcJ+s239qiGEmZ/AA+SO2eb1pvjRon
xT/eE9memoVR9ZC+4g83VOmbT/5xgn5MgQCr+UiC/JRJ75ZRRYvNdsWLKUtW1Odf
geGoZA+SX/pxHA8sLDMczMEarYpPo9EUqKvAQUv9KApb3fAhXGdhh8XKfB3gSYXj
qozxsCPX+Bs4yT89VIMgcEqodRlcfdPMRD28X/fBElKUQggQ8p8OYBlRsUzy6zWH
+1an84r898T3decY+RZHPUjWVPSIVMKa+WfHXxn39m1CdURMNnOL2rOUDEhfuzoW
lqukb+sPsavoy8xLGvh7+awBRLChpSNO2ws7amA3fwchIEsU3QQ2/8oka4lUstO8
wWim4juwaZyjBeFPq5kMLtQc8/Bzi3IK8FRS0g2xOw8y/Oxm0jWHvTZC7ADQP3VK
TaAbjDHXUijDmHL0eZoenjTsthlrQJtt06xwp3N8KxxVxiwTBZR80F1S4KzuAaWz
FESBcQJHd+0Hs0s6w9wWXZxxTv557Y/pFTXj9GBLjXFpV1xk0Fp8eKnfSGt2O4CI
p/WkA+itzDOdCHv4ffo0W2tGBp+dS5cKbKWX+7FWigqYT+ff/1NJBsoEExq7Ctsa
i041eOGN8T6QH0vlQ5w3dKGbM54BNjZglRkRxD3SuZytQr+i1G5CLSchkLLj3kGg
+OC/r3Qk1giOLgWvisM0PGStlVYYY0sbcqEpUGFkQS4hPOFzxW7KO9lpCwyf1atp
rUc3w9ZOLAkAb493GVDDkQkPe7SXiqiWnibndTUUWMYAek9JUlX03SEdA+w8qSJJ
5/N95sBMlPdTQRgbQ9iY+nAlOmDuZuyp4pYLHCT39OFmLMfpyAFdaNk+/csajGnI
jFzhwVRDeYp9OMwFOJQXm+ZcU8FiYviYaLqjcASLlYa0XpcsR57dJsXKBbk2WO1E
VjrZp4/DvP6Y8cKNmv9Vg68Drp7v2wUHgr39f4j+5WAq6XdgGKU9++pYjj2JBndE
Jk6lu/TNs3AY0Bp8pzH2pbiImSj9OZxJ4s+36X75ghpwZFXDyh8hMvNp+xV6iJxq
EdN342xJoYEmus7YvohAj7JyIm6Bsd5MAuOsfIQLSD6YoYGY0pjUCh+m8HcZNWfG
Vvu99SII2ebXYRJf9/UhcM/sSrVq+MX3CIV/X+pFTyn/CUN+jg7YBO5k9KYTLd2V
tgAYSsr5XGobv8FACl0WtQyC9fVKEDWcU68bgeohk6EWEGFq3R2ifMUyqa9ajQcz
ZLUpk06YLqhraDQ4tMHsTgITY5fL2XWmOLcrcJxPsVC913OCUmCxPNbkBNCYNEb9
XSvPFfwZVc26uP9PN5OjPenu8/FEiU93wwlKWjrCQEK9iA5eZHLwYRcB/0ZEYnta
XyOi1M46l8L8jtWdaBq1/MjwibPPEMOBEJBOrrvOa2A3GhX3gFsJ5xMnASZ2zQgA
S7sdCs4AFW7PEh+wZMWKadlJYf7VXf9ZW5Fwo9TwlfDztfKqsQ4tRX/fwfYJSo6l
TN6oeCDMVL2QRQ7G5k1OVHX/D5138HrTuzaZgiVcvVu6dAF7jV9BNahYxpgZ0omW
WfIwOz1H5ZyxroRuki1qWbVXj+MPYfT19D8SjkuwoX3ys32QE3Ww5DXpicOj6iSg
Xl34oXPc7gij6F6eth4/Q94JXL0LKc/jHXbmS94qJEVVcvey/eFg9KyWs0HG+hbr
5481i9h/WzgBcwf41a6budBVl80f/OsREZSorKJqRuOoxkYVJLk3UymmFU30kvqG
2mv3HX4WxXV0K/wogYTpUNq4iPJghJ+29Y7fD9NkyyMw+Y75pmD6hpCld1abAgGJ
qtud9q9z2VwGOBdY180hl4NRDiNrLVhPFixQFFleamisqPckqoQnpFcWQSiqpPeD
26gwr2LIDnGvSnVAseHrTAMdDixRV5gt9HqzY6SdXpXn6E0eSKN0p43zpfTgpKPk
QnL+OGzQNq99tadJvZ700K2sGeASiYD/3xJPcYgVXXXfmVc+PurNZbzyE3Xfym5l
2NcwWAzSGNpJ/3JM2fgMnZUPGvEHQcX41vPakefKIVmAfiEAxUyAPjNYuwvsjGm0
mDCODE21561wx9GsJvSFdR0FPQxfxq82U80fFqf8AQmFJsqSx8DBklvamf7F1kwJ
zDsy/G1HY5AnEl8Gdz0NrvHr4i2BNVXyBjQoyhRgXflkmjryKVgSiz32/I9bd7S2
YywFWI29soVfEg4s0yYGf35hkf76VNoMMizWkUUvj4nwK6uNbu8hBi0x333RNxIF
6EhVWRDFm5q2Ewgq5bWrG9+qrc2AyCBwHnPpq84xLghrMfDDrAFMwaGy/CFRylds
aOEvpoIk/TjAOm7ANxGqHJiRoYa6xp6pcsiFi1wqBwSL3TG17/4UUMxNAO/tUwVM
4YBdxoAyZGBxrSgganwrsfXkhKGgXC6p0HOI1cDgKRh9mJJf/WnT5ZfaYiyMqV02
JHqOP4aPdcS0iw+uL+CHbxzVghdPFPJ/FNZIoKfW9DDkcMm2+cGqTO/yIcfy/qIH
lJ1vlRcvoTivsgHdGUgnEBqMluh8MOhHT0EkT7qgztY79eTYmsNAOsQbPQp3n3/I
zuT8T6+a04lWv8lgewlQY5YVXiDCmH22rP1mSBq0RI9Mn/1l9ITz20cpXqc7BP8n
DkANInzlmWxBtsy9gQSalj6Opn7tanj4Sge49f1/4A0l0/vYGL10OziP4+v0Fuex
yesuj2hQpNLFx5SkSRJt5gEHvh5M4Uc0gTzYO3a5ycJN2vB4+ENMv14CEinr6zze
JSDA8izKct48s24jzWIRok7kQ+SrBN7QByOea3h9Q9ADv7whj8axKzi35Tp+aUTz
2fZkjuoJEVGMKb325vG6pMOLkV7HbHRMCCjPMdXKB6KIC57a1hWiv5dPIQaXtEPf
yrRxHR5IahzektHbTK7Lk6z8K41U9CEcHKNHFzLSmZw45Z8y+f4PYFaq1pP0pyJy
CedXnXw9o1yBxCw4KhBxsX7gNgzDNdNvoyluPitd1t3TDUHFQNC6SNrzKM1JSMA7
z5tpjqSghe3MvXlPIuJ2pAOAeBGKMp4d4kREF9uplYPwSbiPZYuI8RoEiIUpnWXg
QTtVgTXP/eBrnV/p6PrdZwf9mfgeCP4sOGfPUPyoeoBh3fuoaWm80Rol4/NBI799
ZIhcm4UuQFpmjSRXhoTiLJpBmpT47r7M3ug5Z5kj6Gc559XLmbkKWrwcPQaak0W7
pcnkassKXy2ctUdoAqYUTBBKbPYWWRVFyrDUdaOJzkbc85QPpIRtEYU5yo68s8Fz
8/np0Uzw+imsY/LvQtY2y83ngXWrIyPNjdPDONSaZGiuUiYOtBsD48smFJNmvo1B
uP9OUb7m+7GmCn4oRbfbjSlirYm/uIeRM4NL8huUd5A8xg1Dpkt5rXgXFjoHcyCV
a2ofDwvNVwSANMYB0Nm9j26yMYFLbG6HFjiUi0fVkdMpp1M14OMFw/iOmqZkb+4m
WdaafQiD9lFhibGHZYZ8jctkGdYzn7YxcnHENQkwXrPZEljvfsvjqGpZDG/eBGbm
al0FIkjSPU2XUySOGZryBN0AkAZ+9Jm+ODS58iHgZiRMcDXEGdFoGe6VDAqQEmHU
DGAUHn8PF1LHKWMm+08m9TPfu7Pm98W76BOJ3Ow/wbAzQSWMzdHYmTfvSsCJRknf
7MLrsXT5vn2CQTW9i+FyYa0LqwbwtM4WCOKhuZULOSAmrpYs1sylo2Za+XZTiRa4
a+be9c7EAYCaHSgvZCZS+4dYryiYmESSJ1owZ4aH2Qqi3McYVvoiOj14o2NwgWd0
LbXw9NlINvFAGdItqh8ClEG9zZsodk/17soNRBE61yKZ8Y66id56tDYVBT729rHI
F7IRRV5+VOSP28GBKOtM9seo/3CWlkcYOQwkyED0azs/VsLIWoiPacF2Z2mCjNaE
IbYk7dAIyXxI1E8gPNgTh3yug0o7oBubT8chnZovElTcH+lU5RMC6eo25m86yiDD
ANH5j8udoehIZTSxb2rrTdQdf6HzH8jHeGjGOSTn96jLkruf4oz3ghd/WdyG4cnv
I28eoHEgZ9kNnTE6x2ZEKBY4/wAsuo9mpnrrmmBkoBRNn+zcQcMNW1uROAGSqdQ4
E4n78NJEY4dcf60TZ764a6sy9e6Y1LPU14kV+2cLh5D6dU7ZsyKToPbgBHHD9Wq1
qOapCco4K6May5n9xtIOpb25ZN5RB6spSihSdJj1MhGkLgrX+Z1T4pettT34mtq6
sYpEUUA1SqYTPm8o6Q9BmeoAs/YjRYqW/aaWU6ZoUDVKYo1qCX9OiqlNMgwVdfIb
aVL4rB1GKdgBd3IcfSQHA2RcKa2RI3jgGS8cZFvnGHUTXmS5kA3cbqRF3LKS2FnH
WuesDSzTjLuG1L8S+czblbH4rUOvqLyMeBx8/DKed2mrFnh1wwCDsBbRh7D+FsTp
RPFpZbBxOnL7uzBzv+AS54AWXNgOcYITsIk0zPvitklWJZbpgEa9tdlaS6EcMXQC
FIHAz13AlCo1ywOhMa+hLEpwywwcdCcB0M4sSYYV+mYEeJJtEfCXS8vQ7CB0YlP8
XwzewtSJ7OEqfo63LEljw9CU8fC4yt+wk+UvAcVcW36hhj4F/5muWq2H0XniLrwt
XlLbph5bGPyGwIMHMfaQlaoEWJWiDUaI8X7d4GxVPav3Wb/cfgc2fjJUybDopefO
5ntGjesJtqfcmlngSgif8t4fRmKufHK1vzc/ugUpXuU3l3kMMMlDRAae7jPdHgtx
T3gL2GVQxEIPzXeorhNhcDMAaN8QuEB8FkZNlNVltHo59zFiJc0GwBEksxGP06ML
PsiP+8G3260ChTcuKgg9XKEhBGT73aql5WEADlSqwPWS2mnL5zscQVqAhaBFu+QH
dG0aLvrg9m32zZg3TnTkICc0AThQMuLJG7ywlOxHm8WfRPA8YvZSggQXa9+F9Xqz
CkI5ILP4JTvwfzDDKiHDTvfVObMrHXRZ0WmSo1ZFdjk5sOpSo+yV683wRXxmYuVK
KPXwrL1P40XW5Dyou3fZQEz9rD3ZQAC81cC7l19ZnnvQ1Sx3MPekY21D58K4xxAc
jkJpayLNk5hsvFl8TNm/ZPjSPi7OEyGvRj5pi7UoUldWKq40ve54r0WJDBCuzHZP
VT0iWnLiPC5+gml38rIP42XZDc5rwTn0bfklJW4t5HXQT2IF4y+X3YOaAKVeFBZ6
+VkvcTEd7pN/t4Wit3wU8zseFLflY4/1NuuRkwu+5sADyNrdOFdTUsCTPqSr3f1/
Dn9T3mm8PQnjgkSLBgclnG2BZ+jV2boRkw1XmlKpLVmawXbJsLUwbHX49ElDoVCP
krfwBkoE1p0Aa6q1TLSYPPjPigZT6HpjzHaEQZMQdditLwLtnJ3HT9MJtV4ORhMI
GW/fNAgjmVAB1NN89HJwsHTc3x6GWMx9/MSDPT6EfPfkmIuvHMxqlqakf1lxK/sJ
uJwhGgIJ82D+2+ewcIVF7rF0wS93BaqZGeHhdu9AkW+sLVxaKQ+zS76b10h+Ugwf
fnQ79p1s8Ys7GPE5MQA5WutHox0yxW1GfSMr84rKSHa59juj6Ngpbr+pt1ITEgTV
4kv10fuCsXYcT9SkofBLawLEsNoKn41yn4tVtvuEWgqqgX1X85IwIrhMHBISRqkS
Ab8hdT9zpYMfVYfVNB5RN4cmbyX0zE5qcxlxPX91twspMxZI4U5pejmTAt7fYKXn
dyQrEKclbOg1Ww1kqDZGbf4cls42+DexmZz6e5nbMb2EL8PMG1Oz7gziUi6o245s
FYJkz+xPr+H/1/ebBRcRVUCCVy3sUx3ij2GX6zgKG2yRG7Ag/Inw5Tm/iLX7Oudo
OEp/VXx6QCzWLMkjzW03MZQ1lrhCFSXLdanoM0V0Z3a30MMzPvV/AyJxir4jTycm
B1zdu4EFJFl8zxvZ/kzL9Ty1Pd9/tggmyTy5C3j7BscHTfuhDgswPqaeKXUaPpeA
M2/BIfyejX373hj/dPmpYldq6OrKYljugG90ILPQKBji+z2SvYIlUQtTgR8tWGEr
Y/ntn1no1XETCYObj3HNPmJR1uMl+GngX5S0Ug8lWZFReytHofZ19z1uJcW58SBz
/WW8xx/e+RV1ol18YBT7+Iot3M1AQpdP+dOnK6Xh3PFVMKEHW8CE6fKgU/cHzHCg
QqhECiJPRdsvwnIRJ7TMlv6k7DTf2/JRnjsELS3FSGG2OrguMaRW5NMf2DkRpIbi
yJpLIa1neQHyCXrXeEBAwiQvcTGRBDfNxrEm3WvcXBqYEEuOqGF8HE/hVLLFWskQ
ATe+TQrRhZj4jHpw2Jee8kBELwmNCnMZVtab6OOaicYsyWLzUdh0WkftX8UxNlwp
K1Cheei/m5ZQ+7tQsNCQCaNog92XarMctQOOhYDz2qdji9+9KAgCPhLtidSbeXwR
qf+JEuPKOsySJXVwtfbjRXRqylDOoiwz91St2tQdI3gAy1hueACzsH7yQ9kZ1PMy
a35yDvY/WgsYOttcXvILs3IxZ6MCEgc+RxsUQSiqdSpf4IHoGCmxuYW+ESMYjsM1
xi9SwtckAwvKSCkqLujJCRXcC6JkN259uZxy4SX1Kf99bJLU6TCaSF4IisbNPgSH
d7KpfWXViXUjMH47ZKQWkUUnI4+5CNP4/13aC+YklYMVdZ+A6H4usaOTpUdy5URe
e+HdtVNFQES+FB3Vgl6FkGtcKfNZTYQBmkEKL9iTxnbm4Hu0IVEmgM280Qpu78A1
paIa9uJvI+QgPopwWcq6EaUOXtyQQipU0Oz2T2gAn37T/0PM69GZajZQhNgJK4ay
FDh/eO9+xU+ZLqfh6sRAIqI2qBZ2kC9d/QRlvaPAQv8hAdWigkjnUVSaA68MBsod
wI92vLNzaPtEjT9D11T3Q6ErZsbxS4ZJQ36zMwbfyCLA72QbDHmZYvnnAktDNCPS
ixlBQloBfnfA/ufiJ9+WWGMX+Fc9PLUNaVMKrKYm9yvp9bqAH2d3N0bixjngLKnr
vGbTG2hQaS54KQw3Ul0oxd3XnuB5qckFqXmtAxaEm2+UzsywFlc2oKrTHxXW69cX
v+/Gnvf/z3BzOtCME6wnItInMMwMPqpfuy8RLVcRnaZIXFIgY+Kcvu1G66852bTX
VyGlKfi6OpYJbRhINtyYhuycMr720mYGpcMvo6wcHDdGPSbMZDGzrRZb59g93PfU
kkFJD4r7725bRfTj5fkp1hav9UuutBb6t0XAiF4pdOV2bM3tYdnPNlAgKFSri+8n
6u4IvGtCq7irPph2/n4agaIoGQdEwXym2lTNl1msvTPFzmczM55KvSFEl/rJuYxA
tkegECpjv6xqZd+c2JQ+ZBq9liAEwjqnWp5pJMmdmFSBPNqJ6JsPBtMcQgYTeRVH
3KpMAJl29/0EVfKE8jD8Tg0/VXLYs662nauL0po7G+1VEF6hRT+OakNrKWN+laGn
WBf5N7oRveGq+cC3lBdKPKzOXrADqQwBCOGcI/1ZOYDD0KgrYr54C9YVPsNF390q
nr+yL9lfvaTCfmfs3ujKVBdudkCXePsaAE/eFGy3R+QatIA6tjMSBeoD9L3jGOvf
T/2Fb0swoXPDGPkJKNynSA4JvyTA+8uv9bAvVum63MJyTgdfdCAke/MDm8xGtUdY
ygbtW1IK1S0w8QolBzJbp0KQeX5yovLJn5StQ++3wvMA28BIH5TGLHTMoT69uWpv
WJp+oB9V1Kqs5fZFKAdRfzwKkwZusFbpX/g6h6Pbhr/pLLchb97gdYiq4iwEkgHX
lrCibLBCTu8GOHK0wz/bXn4/bxNtKkH1F1rlE+1+dGSFWPLjSqX4lueVyzGSQJJA
ToHLLQpJQxSegF5w8QymbsGlZI1jvfv96QEn+R8Q9ucdgCb8Hgt82R354g4A2BnZ
ecz6BO6ao2ELp9FWlKsSK9uFqw2o3K1736kmGnTuiHVIw0x4/nspKZAi5N81Tx/r
m+Fv6mhnDSuQaPWVwcKSSBSXRpqjS+vbczrGfDlcvBUysBtNT0755LyXkPB60QDz
nXVR7Byxcbevg+K7YkStAR4yRE2uXHp/VtjaNeDJQkbb9kqd4RN1Rl7jUmi/Tr4r
N+xYG4e2c6QaK6Is7hVpYRgkkEUPZGbhf0aQKyF3dKmyN9LQCj/PELPRdaGGeXIl
2VLgvV2mIb4D5rHQE2lwJGf5lAsW1ZlcZaU8xr6G+4rECtQKslwVD3GPBg6xtz8I
jiYXymAlbtgWo3LHdGkRtA2f8sTNevlkfrmdFLDnb0Bh8sslbT7dxIcYayB2b3nr
cdXgukUnGcx9b6Pc5MOnKCXNyramX2nUiA3iwWBo6ZmwfZ5iuPvhDmulaY0jctd4
/i4GO3/Ea/ihz5FFWCDRotLywxJz9bMfKlHgsKxjg0X4EdaOBqK9VvYiFtKL4y+1
YDQ03qDvy8SOokKUm8QJ5PlI1wfDoacrGtoEPxfsYPKb7Z+XsjAB71xrNjPJX8P1
j/9TuZv6s7TjADqxsdkCAtkfDdVyEQ7rEuFHAAXSb9wxxoxDxakk2rz1F9SUd+vK
n3eYocsx4cPapLlRVxCZeRWf4EmYEYb7N7rXs9RLRkM4u3YRjGN7E7piUHnjy+ko
ET0LXHid8SiTLz3u638rYPNoqzgpCO46mZ5XunibtB0rHfRnu9Rk+ZXhsLC2g0N/
xzGNqYf2zZPY5kxscWJUfYyqZSAUNsb3Z3jjwWTJa73gZ81xE6Cp/lp499W+PP0O
sHL+lIlzcnD3JnDXrJGazje9sNDmozu70oIS+5fqBlwwKtkr1rSUkUa1q7TBDQXw
XeJbMw5rDfuFfEb0XV/p9eA0v3jyjWpvl2K3w0C49NPuUVy9iU0k2934Oz0aRv9z
EFG2kdKgp1CRhkaBvDU9fqhY5ugdDWNEJcF1D1/rInaVUnQ0KZ44FyW9R5rxDzVq
IGTIG78R2IITwuPu9MEUPyEggJ22vtXt1ddBZFuiAfOfio4Q+sued3r3ZgLhEyQz
aDq4Z6nm/1WGOr8ExQVyktbV1/tDyP4Mdlkx1LhhAnA8JPxWBDs3wnw/N8QJQtuJ
CX3ATepUh3bT8MyCL6GTHlldvSivlVdgG9qVed3NDMavo4SICrsMFnSUk93A2peW
qNfCn6OM7+lWOfqlCFj5fSogclpZzOZqJtv1z7mo3eLnVKJL7IoY0Aq3IZrUvzml
RW9i7Itqe6kWnNNWelMyO1QW4L5sE0BMVH/s8XT62keqFR6q6inhR7+DvrRtmCd2
FfzUTpVKrrlFEX54Zg39O8k78FtsVfn5zzdsBAbfp4lkkMslCDh67ZJUu5kyssRw
pNXK1Wk3szEBruMKWVBq7HnaEooH0hI2NN5zSrJSwUnqU71yBHu+5zn/Owm6rWvw
ujXSaPbwh64rbYIS+YLqbAONN/cVGVTGCDvGScP4Oy2v7inECzw8T3MHOqik4obe
x38POb64ZVzyjSa+LqDYBjJ3a0wUntPw5wjPiK3VCMZd3xM451Q23LYlEdUrK4d8
lcxL/1KghYvEAZK4sK/g8VVA2XnlUVu4SMI5G2l64R2R87Ri2WxKiPvdbJ5fgBaW
vt9lkBrMVZsHo9/Lp6d4Xe8wHuYTdbAT15FoQz+mugKD1fklcRWLnOX4cfmfOA4c
UEXOECY27sQaRJFe2YM5jarP+1RXkJr7W1/tui2fGx4wPavbmnNukQP8udZK2ZD1
HkZzi+0+JtKtJoM6uCG0FOMcs6bMWb2tgeV/ybj0qYjerJWGHK42jyI+DFOFn2Yd
lFVt41SXTpgUdAFVsYt3nQRAzQ5UXVl47EzXs4S9O+NjbdTwkNO+HjUrSTp2uu4E
93M4lzJtgB4bDqp+2uW+Ig4P7rUu29Njrc+hL3zF3t8DD0uz1skLL28VFbmF6GPr
BxJ3yyUnN4IhCPvw1pBxLjdDhkY1U8zJplaTIL7yZEMuQTsH+7NgJKwjW0WYPIx+
NEZQERTA2n5XmRCgr5lGyuPLQh00/2ESi24VTaqb5QQogzGuUEu3gZy8iBqZ8Uca
WXNHteoZOXdN6rCV/8rzPPhELWBJjR+60X0PKmWRdeGpSxGo+n6/ejRiWe2wk4U7
1vy6WCvBXuhDdTQUn8eaAHYLHaermr0rrZe9DVxKZaSS7nO93TPaI20JGQ90zy+W
y1fAZskLY5DOwnASQkF363crs6krZKba9z1qHLrA7IsFUz1cfYMjZVcOjDy1DhfG
TlI/X6327Ap94eE+JBO/DBX+3hAkLTTE0kCv31BqGBmX13V1YFaTSq/+Oa07vuGd
58S8u4JVTrBJy7pY/xt8hcKFKiQRa+WIwEhOFq6AWz52JaRlRIFwOLNpXf4vZQ9s
OMF7LsPS3kqFiwo+ixh6XJLVz7JkBNzzVd8cYUMOfjSkKn1UBF0Bs8aL1V3bjTe2
lfGts+3dmo4mREA+H9dLboxNz+W4wU+0XA1x7GanZjkh71KbMXoR3r14bYbfaK52
fEGO+bsCmzgEzt0vX6tlRVSLNKSxfpCEmVMDCHEoO8mWCFH1GdrxJEqXEGcdxCPO
WO4tZDtVID/7zsyfXlB9EB37JpbGvhWOR+AYVQQsidrGIcOyX0BxUAU12t8agoe8
1DQDzYi7PKEC8KlhXv/kbPFlAWTxgqhFHPZt3ZlxCpT0Oje1vagkKMiOiJj9Wc+L
yNSzEKVawjf+CGuoAWi5KhDjgHuBZh2jC9uEDiQm8wlttqgz986kR6oKltjA8yDj
4Q/lVfdzRoZ1qj5xhKiLVJ3JFDcUFtmfMVoygE22Hy+xagSLhyaqicV6iNSUoaCE
lHWq8e08QSNGA/9rM8UlVwEoPi9rmaYSU2Mk2nZvruBLi1A90/zMeBofHt3IhNnV
W8QVTj+/tm2V4EIyRsmInm5uPUdh7nUS+qtqKQYAWXIVfSHALAZ9jvzOUGbK7H4/
iGKTowbP2bzgw9GWg5+fKuNV6p+X5rEjtiFqIEZKVyc/wBJihO091IyIptWbPuZX
npzScW3zdf5pQTAAnGlYJCWlMni1PakzP4uJuDQ/GRBiWfkebxKc2sdVKhFwN+2Q
qK0D7N2LrrBpSm3oirtg6ZkNHvAKNAZSBova86Ki4ePwBBm4ZMbJQ46LoOPYg7Ur
7bRCS1zStVzByaQjix6Hvyf8BIEkqUrUJSXPhwuh84Z6vkdCOT24OgzWF3H1SW57
QGHqWf14IiQOsinC+5UTSXdAqQSw5SfL6XSOUP+wp9VqMwVTIOuYf7zXmtv/+uk4
vwjtoHmivzWda86++zzQr8BzDHwuPMjLfK1oGKyG6MZDjpFkY2MBo6f+GrQrZEgW
6Md1G7XMtb+xnl0DaKuW6f8zgeVYLD8Drx4CA1q8mJkbH67ZnsUwXrAS6rGrYAtC
gSx35oh2Sj0YuFHeEcwdGwlxo9jI2RfaON4HWFahnaw6M8iojfO1teZGyQ1MyD36
vb9pMz+6ETGGj5fzyptEOFctZTnFregtIuBfrKAJlicjxoLmgx4CW/zkrs5Gb38K
AIDHU4oj/7GJ9BDZTW2KUaTZXS+0q6vRltGaxu78Hhtu9jyDgbPqIQgfzIEf13cg
x7u3FPGFQFTm2HOhSrHgD0tsSBpHy7m2ijRZue0N7p8bOjdinNz/LH80GXaIfSSq
CVblGj4f3l+q3ScahJcP+vsZotcoEU1H0y7ErJI5kCVbjoLcV4pRMrC/rTgudjST
cwTCPGwXaC6x47sCGCnMAi2DrhEiZXA05ep4jOCTapn19zkQTVxTuOeXT/XAeuDt
W7wcmzVXyfQmOEhbl8uXjfY7rJMC2ZRy/rqq26+/h8Qn5aCH0Yti8AnhN3lZnAKX
ei34Mka0bo4cBJ1K8xFvZdwsZxfQR9Gwt7DlCVhIMGm9awj5/eUaUQ8b/FHiCmCO
LXbjvddslpYsS2o9mGHDMUQH3evY+QutGWl8TWKIYxtSAqQ0oNJY3sAL69Y4n713
MvmzEoENKe6jP6U1zlbNLUpAjNP4Ix6eFsvw+O+VyrahyV4oI+Ls7f5vEoKCvVB8
5lyqq2dsVUDKvLfwVEahd/k2uNBzwQ04HZMSmZxOT9YnmqZmWbvF99v84xGRlu1L
sql4XU8mcNXPWP7nxP1Ph/ityKhTvIiGc6IbBzhbGTdq0NzA1XirkKN6gCcHwsQB
EPl/SYCPk9jR3wR6pNL481qwxso/Hd1VmDN49iriAZTU5GtmdGOO0GGjUkBUVAjT
QNRQ2Rn/EY8ivvROFv/kd2lXXIkECnq2XtVRtCfx/cgrUPHcAyCjcPzSlT3A07qc
z2EukA3GMPYT5D+Hft+jn5ZnZhWJgGEjrVWlD5Ry9j2FA7RrXxI1xXZfkZWyRq/7
5iCIQUUhFILQ25BG3eZpmyN2ege3MpU94/VTaeCqn3rpt494jEGsEfh8wRqkx8pH
OloZ6tbZ2IzssANQ3HNlW5UgHtDhMYOHGsCGisd25z18MbnNHJyCfNhjWe220IWC
hX/ayAwxC3SYvJsaF0Ozbf58e88cU13whzi4IHHwgVzGuJLfOSaYiuojuDhZI7by
nLTYOs24vVhVbLfdTM+z/Nuk/Vl4MHEyzYMmPTiX+GRFGm4Pvy6NbcYhU9aPNtZ0
dBmRwVK9uMgzfhNVwxwE/hSZOdVlftXG9/+S6umOYOVi7UUJ+JD70SYYtLgfvjE0
hNytum9jJwscb1vLkRFfnHdmO7L73nurt+jYv20LVu09kllwghPxvKyKi/UdW4mz
qcFxAuww6j/n3qAr7wMKcGRBIHqD3V1AdTRau2/PdFbIdCB92Wi0x3h4VnfEnW3/
wK1JNe6ufU/2IuHoI/BeyUj1xxEVGrFTse91n895ebomqdCBZV+h/oo6w8Kx4rL1
or6xA1F6dC3W8r1/Zt/4c99rwY1hQn+mZz8SAa7lK0NyPkS9SGmn1epvab865SvN
JkTnyHzTm4KXo7rBCnMLVWBlHDMF1CFT3cUYxdNvqxelpEppwcfwduZK1AHbFmps
g2eQwtzV52OHj4EMqNCU92ZLDxr5Eg/gia6sQCjTl43eATomAdN+PxjMRt7oEHhP
Yvt4oHI5QUPnBJNZL6wFR49tAv8tR3ZGwuGPFTGfmlYc+IgxozYhbFy8et4ZZ6Vp
6V0ovmz0ccDdbwtSmdqzTmmDj7hwbZrEH9BxElJWkyga7k6/dL72QZr/ZaNENSJN
6/GMxyQfmcCiVmXZ5V/fM2Sig3TlLNsugnuH/gh53GdJrDPR2DnvltMHpVAr2gJU
TgeOjyTtcIZC94rRg5iFxzW/HJ7RG0/VCNOjL9xpAQ3qG6FnHdtbInQl4RR6MIGr
bNui+nQ2prrjMgG6pA/XlO/6Di6TIpOtk+LJ0OP0Xx4ncDa3wb2qugwlCiAyTAUK
LqWZ7gg8H9nkQk9X1hWfLVY6+OWIwjIatc6k/LgUNI0rFed2gN8X3DMzr2qH3yG1
fyjcCC3BhgFhd3fLXk5q5qiUniMc2VJQCyKKWTkTirxJ09YIqUcmYiIvwA0HjIMI
DeCERFDaTXQUgi/j+1p6qGnOd4Osb6kQOUmSFHtCwmAeCdM7Vu4cpUI0IeX3Ro8I
QVP2FNtJGyP9BjMsxsQaRO/tesl0AUQt8AA4H+2/fTMQT82F/xcBVcJ8KtVMr6FM
mZGIMYnp/ZdwRYUpsSd9vlhofkHP59NIeubMM4s1fVRGJJxZ6OJtlEgt63WDeo5B
uwWQ78W6PV9r2CjnSTW73GP12xVRPoq59pEThIj96+hNpGjgRRQD1o/4hddhuIzb
5mzhNFnsqs2feSjYmaWU9eYPqM1b7ZiaoHAwBLZTiGgzaZa7ftyd52ikf5KfXFa1
tXsq2XI2JR9SeFb+hfkv/gRAF0cHxgb3fXvbV0E2Oc1uZ5QWwGzbBI/YYapmIExF
jgUQV8TJLkjKPv8YUvG02ZaD/85nKFxV70aZ3IIGa2JtFwwWkdO9nZVY/TzYdhro
s7BrhHPpLe7wFHBD541ZMMJCFW+ksnqcXYWgCWZaG+crKE7tZDCYayrIYf1viL0c
o6AWBoc8EJk72jTC+jqrFI1drcjw+1BB84OMZinM4//Z/m5vE33rD06neYArixTg
AwFsGmA2CtJHI7VlYShCxQ77YDzNxas3QdnI83BxZTtVLI7x+EpzEiGDHszzZgUq
qKCfj74QYn9tYhjK3NAruMc4H0aujZgnvS3BaQoNTurDU8GwQrYi3YwgR8EtZDU+
mbUehWzJKgGtZ1LruMHEEsIccTreos1whNshr8VH71zR5z0aY+ef0wWqAgQ3wgGU
gWQT93Ya9YE5D4B2cfK+6LIHuP8P/bq4r+cYs+vWJcpGMwGSWBHrdr9c/3Jt0ygU
aWH8IE0g4egrxV5hxm830FFmXNkbYSPmIi7ZCMSi13tnV1OQYk82GYZqBQUB0Bzl
ZUsOM6odsyVhqEKcvh1WS3HsVD9dEUGEPPFg9ixOz15EtQywXrWIA1Nz9ECrqZQ2
VDFuLPFv6+OLkZd6YArIya+0l4NAx+vX2tjArcdQAsQXML+l6k1dhPmEpbB75D0o
o7rU2TSR5zXq86OazizP0fGj8EuGwDpy+ODO8GYP26i88AAXoNP/5N0npjgXgtL5
vbdCMkcB5zQxB6jFK0ixV/in/EI9/0vB4mKS7l7m1WxQBgcPYBXUetj9Gp3wsnKS
Jm0/DED/B8ZtrHMV9hB3i/HkOc3mXPCX4v1LUi4gxh8DZSkoaFOh+jj2M3BgI4VT
ESM8J8l44RQQQJS88LKNWblJe8anXFdT/QysifnfNNN1OUhnCy0IUrbsDPAbN7pn
NfFeYraa/ord6CkiyyHa/E2gfD+vCUvaltJNB2pAohZLCez98C8XvYeW0/FImzjL
cLXVrU4n1b5F3o5Y1glMXuOFHW2KpZMUBba8xLTnlfm/GNW+ogZl+DaS3hyIFSRd
JyKjwKrSEPRSQrWetknu4gL06H9oS5qEsMhUbNd7CEuBctJd04QenlMX/AjincxI
Pf9E24/0JsYryLBIYH2dl3rC+HCsI2gfBeSLIaezIoOuNpfm/kegyhYfo7pe45v9
m3BVmcVYahWYHRyp9Wjowo5ZkV0oweKI+E+cpH98myfHdoNiWeujpgBI6+RSGDF4
rDB9sRrGEmxpQkk8zIO3VtPPz4WILm85+Zbb4+924SAriXLxAg8ph0mPYxzx9uJ8
4ph/65z5gn0s/b6zIf7jnEVgo04Ozr346YMIbPRnEUcQJRZKz266F/TXa6H+ONV/
wDrw2kzNTZiSc5fa/0YR/mYql6clcnRm5kQ5nguyMHbcyuwqxs77OjWD+er4xcqY
2B0OuA/REu6sfDWDwXpVcQH0yJC8T+zMVbIzHGuomHl+al/4KnJaITvwdomUnoah
yyLOQxby1z6SO0MGjPToOI9E1BppcREHeyTtDYzfyHRMKq5OZwIbNFbjAaldolMi
sjjNfiornvzFwbq2lah88leBlUkAT7nppfwRFMjf5wqI8mD4YuKQ1jvqL8+vF/N6
hwc8jZaRQneF2sPnK4/XmHkICQ9TsHcgjnTe9zH6xfOhEcZeQ/W0NT2kTzVde/rZ
71ddGtOeNFin6IvOqz68qEy9ULAlWIzgRW/SkUKZ2ORW2EPoskKJz8fYnrmxT0LX
2ZcXqd82wMpJA0Kxz4RoVUjpxuSOx0mLlXUQF9SbRhfs4O2PnVpVO8InLnuqUSQy
WVCQsVHqAd7P9d5kA+Qxn6+GHDk83l9/9xfrc1zM41oDmF+zrY1q1CKYgu5HXUI2
/bB2j2ygDVE45yHPIjWzCIgBvcwsaSxg2qtsJ3MA08Hg7yLa7ZQaVJqWGqfYLmCA
Y53egnyCzbEAxHYOhB+97hg+aeHBwopC/zanJVj6s2Sz5X+hUcJ/gjIPC630XOkR
TGpz+EacW/jvTC4ms2OqR9h9FNx2XhIPnKoWnjij8PCeXFkKAYfpvdoaaY32zPLi
gIUi+OpeIB6U5OaiaL6MHTBZm09NxjKdnLxV88o7gbZJgkg3XTMgUTy38lDOJJZP
na3BDKLCaKL4uPp+koSsE/o1XWNb+fOIOWNuYrOrf8oOfu+z53G6jq8IdOuC979E
EaDT5Wcp2TY3allOUEtkPmEz8i8a/GKwN0fSfYFEEpYVFRmwgY/ykjWnR6BHOHgs
4QqRtKcQ8Udt2L14wseZmNvvMXH5qWZrujjIjPzj2AXS6xP9wwcFnos7EI3drQkn
2Yk3pk/rDoFU27YDlemjbyzAH3Wct1vxP86zQb/vozodbIsm6v+aVJgCBRTbX0xO
Ws2mQAT7vkqD+KLzOF1DEaP4GiUmpC4JCI4hfvz3toHVsichMcgUr2axcn+3I/DB
e7Er9h5Rd2yy10z/fGdGl7RmG+nl8F9jIEUTvdQeCSTTkDliAgz3MRQPQ4WN3OX5
JzfHBB5TPSMrFZ6fDpcGdBgdL593YOFkXAMxZSoXvkajmVB9i/GKsw10RGb07pqu
9F5NrClvLRn32/PzQ2T8Dm5UX6huSzZF2PqSXymJDAG9ue+GfjytBjpJ4OZY2kvH
UsbjLcfL2SnY8CeZT9ga01FG/SmjkWbiqAM145DTuavJYKHeycvx/z0kGCxi1tlp
ZjbtDfApIRP7wp3w6kyUCQDw6RVAH2DSZgPGZeKq0+NdQTsx76bAJS8hxpt93MiY
yPXr6WfP42jkIiZ1iuVmCjilC0Bi1ppuzOHk6Wt05zBvbpAHl3sElL4AuRAEc24v
nf6SWo65p2292sqN5EMbEoKOCFedQ5DsNuaqf8fEOjLM3BqW9VZBfXZVxTUvCaUE
W5bY6d1V5twAWbuVK5zClfqdZNg/TPHmZWSiKW7UXWpzPq14xtWHTBGiUEhqBZHY
5N6kvV9RC3PIUC+YOHrd+NtrID0tMkKz+/ds8/wFfMEXsMeW26NgVv03lLIRgEoR
SwKc7jZFabB34owjOS9mN8L8gPvGTb/zVJHWiJqpLHj3Kh+9u+3EgiRtljtxzwV7
uxz2JGCqtlC5iDROkVg3z1sVccVSk3Gx18DBVcdcIcrPFPb91ss2jmk0bKfpNjL5
5KO5YonWL/x9TngrlmWAwmn+XwK+Vz5Bq+uOvZV3o4n45EWorhh6HNyqgcCpMeFU
Pel/jrQt4nnzNIrpdcv3BppsqOf7Ds0EKqyFARSRKtF8iMKsXjy9JJPg6yXRFA5k
8pe6oAISQtv+KTb2HYT+uNcXOT2bb7nHGQ2pEjTqDfYXC9USBLhpjp986pFeVd0x
gcwz0n74BQ9xH35k2+my3jaFxADlzeXv86/3nIIBfrdlyoyY3C8xkbMLnDCuKX6O
2+OjoIY49XEFBGcpDZ0J2/0cesev4O9IxwwzFzzZPKWLElYrJ/9rLYBhvcvwFACQ
+O4Ze2k9gRuuUsQRmgkuOJ6snjildoHxXG5KW5GPjvHf5U1wDD81W8+imiLwtTox
WVcFz+7DxWpmbLx1OAvsBrhtP3nD/L6eIW6FSAzGwtKjBWP0WioZ+vwR6WlqhvWK
fSc8Q0NXC1ZKP7OvSg+ncZAhX+SBssY3P3ZMnio3ltVPTDbmrP81ynCt6YM9vxwM
7E2ez11wffXzwyFMNeF5dAZTvPMcKyjcPDxLmQ5wqO4e713ampTbGT6GALWLJ+lb
rWV2J//vm8KWnVV5Rc2w9uZvwIUI9cG1E+vtIdCWPaMzUpkuJKQVxVTOZT+Oi4nu
A0MEAxq8bSfGYoShtpgR7L7FCwZP+czzqNmLUlualslwiMlCcN6o8rtlFsxkFt20
V8C09JvVaLMV9BNV6fm7WQadlYeQmNsn1r5IA7G84LCBr4pxX3kwKLYyzreNoGd4
FB5DNFAAoCcQKM3NZ7ttfc022BlHOQdIcqyqo6rfNcHn0nMvgCTK8ktl/oUQGBHD
ALCWy/HeEDe+uU6LLtLkxM6e5ZHERNob4UtxiXqS6vksS6EHDUW4De+hwLBzJIf2
dtH8myoQvJL5iRoId7ZevWQR+O4swuLvDrf0cgA0SKBhPucDSs4lelykFgA4nyny
odXrrWY8zQtW7SlIlwEKDD7B3cuSHJEBPIiAnPfX37C6LWYHoxxI7HhdsHR0iu/C
vWdi7nXSkKUautLpv1k/3jWV9ECICtA9NBdmRDYuR8VkeOgsluU77+ikDpTChRCV
5YU0+Rt3Mhnd3U+LFeaIvDCbJScWQVM5kobz2n4SWL9IBvGlGl9fKU0dpsedswD3
vwZk+dbNFgoUx1YNjGiU2r2+UWuvq1ydYIvdFmtMM5WvNDtjQbc2A/3pWO4C2e8g
NtOCz8zt1aeLi/w2erW/kH8SRkGQZWI5WeNNKsywyinevBUnOI82VjFOH1un3SM7
3ANW5dCdqdd66X3fIlMxEbCeiWC8QGcdFyC+9vtAswl+MglyqndF+gFRkguczmX9
t5sY5UIk9FOVhPQfxGi9oKfHtDr4TxIEeDsPH6vgMZZLpuHeIry0VjbJa+r6ns3H
+SEF3Jn2jVzf1MHh0yFL+ET+3EJLpGQhC4fjeT0/xnSgk1/ipDwn0MMk2Bglp6Up
fDswysoRNQUsKEhUMrvlY2KfvnqfRlB8h4TeYEy2gnRWrXaAp5sdcpVgHSsAD1tt
JfTiAoLHmnxHvFMa4b2VgWnrSjd4G7SVRxGfj9fTbdQv7iedmjjpt8PdVAPgakLM
R3RANSLBVJsYIe+xybH+jWGMfbcvxgOVrqdseasXgyfGEqKs7NR1hLjAXRulMyJ6
UNvHZFTlJq8adRcyEHhDvpra6Rqpu2ITmCxAYYBySHnHkGXmv4s7VVStUSHQ1RL+
5YbIS/g3wPFsvzeVrJaGtoUPzXyKK921E+tR3hZQS1tCfVJwAY1lCayqbjfQqkMc
NU6IRtVhGSoFbSbVfqON7obbi34757JiBgLqWVn+GJpQZmlVlxdM/IJ6GBhqoPUz
xTGERNWGUFxWo6FIk1EAPWpYHwtx0Xl3UE2t1uRAPEvhLmO4+7468DHVR+jihkNt
7RoiYcyAxvaXu9ETw9HlgvwjvXOKvmvTwXE5kLDuLQnHeyFJB8KDy197tN1A53wG
LmMfqVFvw1i20ljt8LeCY6XzNEOiUWYuzwcP1xOfOpZIympq2NMZwXL3fHw3cPsz
2dB1IOvQHjGra4ysRJYelbwwR1ma6sfmvgkGMnDGpsE4wMnjhnd+CVdSNVhYXCCN
nlq4lKdqM9DqofaCAxH478Nv3lq4sX6WYfgjygj8YmaBvdaLxxperpXSeH3CaoiT
NrcVI4pvxYtGusXdrcm/c7fcU8ZH9HRtYYp9y5IRWBok6IMW535/gucawyz9c/F9
Wu4qEQfwoZG30XbHIZYQ0nuMlgE9da00KdDpMr1+R3M5XmEm213zqIBc+33WXIpH
UNuZc0IlMoCnyOjg+uDlWnChJiNScWwk6v30vRpafjCaZ1pMyEZMTkmeLjEfMgkO
dtaEwRaM1GY536ceeYC0r7F4dyvJVTWbvKhzbepfcqNgDzimZAQ95VMf9OStSAkL
VA/UimB0FsU7slapkpEPJ+bdoqM1sHg7dZn1sF8n/NRH+mB3tS/ax7akp8AGB6XT
8irNqChL6L4ktNYmk3npqc65vUAONqNSNwRAQz3EfyvAlmSb4LkGj95KxIaZgAU4
7F4nYkInti+ZEzSBUZt038Tt0S0UC7Uv7JZO58fXROW1+3R3RKSDEA7i4+TIBw8y
SXN2H2fBa1SYoALeeCybCH6omGIikH3itlrw3vJyazAXjcl1qRZBfeerlRqtI9zO
zJdeIHo2m/f7rAikXmNNzy1YOWRQIbF6gYZ3JPDX+OVJMVTWn7znzuleOX8LF30Y
NkgFxIVh2GegjzTP6X8xPqadawBoC+W4zzwxrgacBy9qEbuqfiaHkWz2dxYCfWsx
9Ywnr0Ktbi7jeRfJvEVxqkurU+bGeTxzOu5JZEL9jMyoJOvxljqL8WWTLzdHJyu9
jedO7yWkc/U2bznSFd1LAmbI6nFEZuZP8czV6Qeept3pXposa6WP5a2k1yySiuEv
9uF0zFCivFw6InGGBMJO6zBYV5l9Nflcm41u0RZg4hgiHPGqL3gn6GoYu4qV6dEb
9QOItmDu91ai+tbc459MXkBpDqNe4yZmPbBqOHWoh8t7bSXERZYgormzs+LWzBwp
oOMveYidkfdR99va3Y8Xx29824F1damkJlSvJC2mJRMUbieN3OnVwtnx3nl3boiS
AwEfiHJXsmy9jvfhUYS8BqRSMRsR79GkTHY7H7ADZPtezdiORxP4JK39oxQD+RA1
m0MceygU1XzT3BWqLTATtoFprpHNdO1XGoJmMqEMkhLufB4p9lZHMzplDwbtgZWc
/xhWu1jDigfdrn1GVHOv3x3GUocv9HeEEssBXAlBAA2nDCb6uB+J37773O417fqz
SzE0roB/C1UxtiB1Z1nJ+ImRginYDU3maWgLbP6IJCdn4tPCHts3rqt5GgJkGg9a
cEPJP6GCMd/c0xG4Dn1zKgzHSpASiZhbZKtrN3OrO+RvUKB7yDiRCao0Xo0asC5t
YSyEWFYE1OZbQBHN5ukxjhlsMaVaf9s6enmEqZyewE0Bn4FMpfAf2vbp5pHPmebX
YHhsaJ6tjolBY8QqVDE1K8G+lKloRR2uYa2/D9kh9aRy97UsPikiIEgyLq2Blvgs
E469jrrVH1NvC80w0cKQvmvMia9/7NJxUj1gZRXRCM7xp7sJ7HCTegHEX0APqm3R
UI+eiTAeiht9AmexVAhp5mc9WFfvT7laVZWtqR/JbBSGnNHEXdabeGHsvVSN2un6
ePI2l6zXSAOXl+EqI8RNay1d8ocIXHVU35slb5umqczE5uQoPJAifHjIBHlIOC8e
Rxc1nRZFz3YiE+Ry8r1dmfE0QDWkz1eco6U5RQpWOpcyogACws7bLTUFjl4rsYBr
Drx37dg5Z1OB35OgRbhAx8ZQxmWCC0lb5BhLFD5alcfzCX30q1W92YTWyoTb0tf/
3ad/SUBkhHkWqV9PHu5qsKj4cPW4E/OcRFwuiH5gZqD8Po5iO3slHxzhApn/8PXM
go+exV0+rdDWjuHpqGYWxGZLHrd0Sg+PmmZnzZsgaP5hyCzvLCfCdTVqG3I75/Rf
QyEbo/CTNYN2MarLIdtpcbDkv8mmNKk66kgZX+xzMPs8Kg0cRXvFpcjoS4/4ZYbs
5jYpw8jboJ03lqiWgWKnj2HX5zl/XJ2YwqOSGK7cAOG1hoGOET0zRK065jAzwUO6
szap/Qu/bFcC+jSA/fi+O8yTvSbcXAVbgJm16sIBtonbpIA/iadHYIG78gAih4m1
AAffaevWPZxqQu7mGOx/YNnEdk/xQ2N8j0ASMMi7l7mZt5ZfJoMyKV1rVEGSEWAd
nOApdzwlh6pr07ELu1rYWVB837TgEvGrFfJvlECVYWuaNgZ13gUIYLA90t87zZzo
25s0cr59IcRA/VR3Ns3IoyqqSJV5FLmPjl8H0NmsLFmg1RGTvDPgAMK8woD3hPXq
QcDQBCOEVcH+zE03uLjYcVFzXn+r4R9uaRYxnA4Z2gYFNobSD+yZMii1TpkKrKVf
SZeoECYnkc7rdT4peD4ctKtEVt+jx31aUDStD9O0emq+IKsvhj9cmnlrSJSMlKUt
L6+boNnU3MnfGfU7W7VNQdhEeQ+CZVa3ruFEy/SOGVOvYCMojf2q5IB6z271eD+H
I/lLyYgAYm/nmldpBG+t02Yhv2g4KzS66fEugl/Bk1161uWlzSS44f2k2FSPE3tG
AXlyCOxEddkw/lDkh5UTWGOr/FATbh0j1yRjvsphRR70b4sFHrrLfyPFYsfa6799
CUo/4y0+ud5uWAXqK8bqVmf1Wd/ZW0kgkCYPVecbABrwP9VjeBECWFGXTYefmWC6
+VPUhlyYtdelaWeBdj0xQRzqpZEFXbnvHt2WqRJNDHSCX2UHYGOEyXkDxWf36NKF
bQTCL9pgmVdICR+6DLLkoiOBK/X/BHL9cVgEo3WrLs5sQEzzjqFJzJGaPYKb6ojt
muiTuF9paY5jpiTnXqSW8T4zhxWJaFJMYA726inYxfmemg+aNI0oxdVcRejOSC1e
d+JZ7PrS22oSAq4B+qYDxU6tFerNCMDPHNvLY2DgrONqncmN23YJvv8anMkI3b1O
OCSZcwJcKLykhqGPkkZxYOuqDPPgB9MzkYY08sd7T8wH0/UF/Sg5Fp1jVegVI950
jJzImg5TTwlTyNy3Rr989nJhYSHoeHdoW5BIoO3ueC3F3iLanlKkbflgAzeRaArf
4yUfqRg/sQfKqYHfw7mJu/mOMJcaWyzzgbyptauRNvUt6T/jXMxEc8xdlfqInJQG
h4urTr8iC8587xDL37VHgaYiEGZ1PPipUF6W7EtcheOchpDaNXwtzd1RD4que1pa
Etr3mYQ1P40X5gjqUy0hBTFr31IuXuYB7IWFAbo7DJt1fgVkatMu9Cq+cOJ0O9+q
Nvnce41C8ONtmqGdoeePe14LbFVuay2SudAAYnuFY6GoGN0hRgQAgrlyFfeU+TQ0
zODM3ocDTGvhgC1gSmVT44RcyMVEyQBdmEI4KMMPr3E4+NzumR66tHmSITQ2i4lK
fZX8XMMRweBdlEkoZpxH0qPgmWd/3ya9Av09mP8CQmSXEoSKvEZFxEYeoMbPZL65
OuJyXJIcT6fk6H2znbCQ27mGJS7M7UjlewzlFMsp6sva9LoCxPs4e41QFv4hDXC6
eU4nIe1n0tUaY+czKfJbFZaJot+IdYMdSl1uycaDgfIPCRhu2t+hxYKa/f5zeA/X
Bh8hAKEREzj+i5PYJaHixfwQ7FsZpgu+KKcx4YAjsmcYXN7bCIO8yj70cK1GC5ya
S1pwVYUvwho9RYnL0xfnOrQYEsgBcsX1+W4Yb3BSA2IE5Az0QKpldkohpwOnRg8R
9+bcgNzvR4VOMRf/kwnMrHKK5IuSbkYPYPmOlta1g1TQ8F+HkWzA6FxZyol7A4qu
MU9tT8lcp3Jpn4gy7WjNhuIOri0A0RBzZjMyEHUK8RgJzxxjumk/hg8lARE+THnj
MkJZmvdOwBmEG3Rh0IS4MTuwOj/J3DLKro9OS2kG/iAsbgq1QTRJBVmWIsmxk5bG
NOU2HnXR1o6A++VIhRSdDRfg/HtM5cdfvlT7zcK/xJXwEbTZl/XK3n185d1zDARd
z0V+3Dcs+Dhgavg0P/CvE/oiF8vCObpct5OnzoxXdigxLzLAkXJp8iw+iKZhkerc
5N5tuozbKnGd3ZUUahmXnfyt+rOAUQ1Gr3ocuIJ3itkWmVmzFgXCrTSt5TLyDwLB
GLOylpzkx1bzW+3jYzbKx8UdU0lD9dSM/W/yWHon9G5B5f/qBj8nH8swRV3TagQ7
V8rRBU55hpoZu7wlZfGuWJDyGdMJp20x4zjOSmu6ishlnbAfDEOgVh55cZIJrZ31
M/iWYg2658ruFlBgmiKLpDgNdN6Zg93eetJWA4+fA9A/JnWv5bkLh6VSnd4dJttA
jytv1A3hZokR3By8ZKRqAW4hYiBokqzyosy9KNuNX9nVFW49TXl7BJ+57uOyrMsX
NhDusMWGoHzUuuQxy4GIUcywvm0B1J/lWvxaoq40kp0Fc1WdZyi+iui+OkjrJN8D
CtKpdBqu9J7JQR9dlP1J0Zr1p1+/SoNBm+CHg8bnGMyIBS3mNsRWsXOu8xv7dwlk
M7Ctv51P3oIL9H2rTM5QcGjI8hrU/Jf1YsgRH/ghK55sJ3tb9+aywcu5FSpxJzjY
mZZKtx5tidSQQSY2/yUhllQSEsC6H7b9FhHIpeImXgxjLr/Q3bLxRXwwgXrO5rIb
dNONJwvPHRf2DtU5P1JE7yhT7FzP2Br65CJL7ZzwG1uZkCigxtHDAn9MvedxVUO9
vojHTJsBjwEdVCYILsAtRXrKeNFrMj1a0D5lYn2DEc3pIR0Hc5UJuahisaPkvu4c
hIHdnbnAq7dCUZaRcMkPhVV/M27KNlyu0qUVtpPBBbjnf4ovbbdV8AwLif7r1LOD
PwE3aIcZPn9q03IjdkNNqVKCg1w5zVOq2rOTqiQLShmGfByCegnJP7Cj1WXC0k+m
Xn4+1GUJwSLr2L3w/Ob7KbMdOGWEUf2P5jNTWXijZ/UV+xCX+k2VhfeNBlS3NEVc
w6lzLyi5PhqdYhJkxSTa1CuMWt8Rg24reEtCZWW/9kfOt1t46KP+fSyVJMZ2pd7g
n5Jg9VCkhqoLEmmS9Bjp0s1UH9aR8aZT/Bt8hISpo7E0ekFsfjuNyXvLx7S8yFpC
HleZv5RB/1kVPvAm9HmnMLrXg4dHSLlR9WnPGOGxR42rlUdXWQRDUdpFBHOVVwfz
mw5K17hyAkJPNFMHzuMG0I0kgxjytcmWA+dsNBFTCHUqRwkvmm3u5YlRDARTzST3
jvqGfhMhu7EpAOmljiUEA21uGJDTQql+hxjLlQ+nUhDbnZJH1Oza01bUBBQQ4hsh
nTByWoilNasNRY9dqu1+Tfz+DQWCDPlAZlxLhl+gPgzme2tt/XOB+LQTZlYqPpxS
GIp6gV2gygPGbfY2/V4g2xQgl2lPbfhfz6EtLYluBSm57OEXE6As1jJCXbVQad0z
wG+1DgzFJLIGSWYKFrZf4c9GO5QqbS10EnW/2NSAuZD2/ddJeRlAK7MHshYHt9re
H0l3bCQe9G9WbqOX/ec7RXRGUhEQ5cC0AuWAuSLYX5s9QcgRwuSx668qxw34Ua97
9Ch7jkhUmRdyDhHirCJxGFHSJqyeol57THGwiTvEI84kxTyjaGfh1aEhAy/AqhoH
vwLusaL3768PwTvBpBj+lQOpJg+3sP0w57Jo1i6eS0EtBVGB9V7G0bA16MHDi71y
Ep9fHdLRhR0uEVPK6ueVn+lWFQ/g68Orar9jMHq2nAwQla57sRU4aDIdGD/JGeh9
LrcmdEd9r2Fbg1NKSudSNg3Rt0xRFDTw7ienV2GEYIhynXwdRMhSKXOEyhEdy5pW
7rPDmIsLG28RTOiWk+vn8QsL5jV3bZB1AQjkv2FukvjLOD91JyUAlohtuIG7XsAI
x8pKd8yEGXZnz/Pvg0M04yX8v/Q7AxkUgwBa//WPCZEb4jSmwZtm0kbzCqfF7WBy
F9z5aXYfsoWdTsY1rdIK1E9+i84o5/JkoB5FamuZa6Rfq7+32mtlGjlNrUA8lps+
KZbJzcEAAx1fAlpJLZBoBC7jsPyWAAIGk1b8xmzdEEFLksjzKVSjRcQTAqBZGBXa
Ga6wHB5AnUovbWJkVOiK1qCqcG9I3NkXKQce9SRNcvrxM4b5T4fE6OgDSny4eudf
bf/wjk9PEKq4vZRV2GR+SYbg/AE8ggJqsvuy96sNnkdCNBIePwNOg+hTVKGJcSCr
uRDC93yXBt4DXiuH5+r1+Zrxn0sP1aDA5TRrRxzLuuBuV+S3S9rN+c+lTu4cZl3B
ci0rW3VK/GAT/Q5doScrxYlLVaTwnxkG3Y0zEWkft7GNhg6scXMVY6kxJdIPTJ8D
tDp4Csymfa9BficAi/xsRlA+CsZnexga6sR6jx4w0Da+cT9HJevLAlIL2ixWQLL7
AUXMp+KbSozeSLjjVTjk4Yvhm1SXvrowffcB0wMzXvE5+hX7IgKFeL7geh62cQbU
aheurdSxOjMWclJe5lomXRTn/VtF7iFn3nagszDjRVO9eDHjk0g9vMguSbnOY/nD
Hh4tyrYXWDjIMiKQXXbDAJnTTnsY+JOl2gwoSRr0oemQW8DnnQBndsdgVeTMIvUu
LDNqHqFhu0V+osjGBpIAOfvnNyB56dvrcYF01rvXbXtoFh19CezCpdKpHz4tnVjR
b+7ANsJiDP/ZPt9TVsP0OOAGlzI2upaaiRlR0Ng5ogCAFC9WQidTBDBF0ciFFDM3
8pcoYi73PM/6I2CqoOeqFEEFn9yS4TvtND+bfoZoIp9D7wmvqgBLd0W5uPK3OutK
rq7OC4WcAx+5F3ej0MStby8/dhxvfROkJny1w71iHcAziL+fU4u49ervDmY0myPD
ugWg82Tz3VVV5W9mZy59CVQrJ9mjI4XSbrmUFvdX5lj5VWcYVqUN0RX8KtVwHQSh
YDrz/CDnjxKiExytMojq8utwG7R6nXtGnnqprblhJ6R0N2DSTyHMKXxU01Cd3i+j
+dN43zf+pnFkowyXxPF2rTI2NrKNyXj2LP9rbYv4jyxMFIT9fgv52anQ9NpVGyOk
raMJsfOI7s5cMfq2QPxzU7mjmuTQXrM4ARYYHeeo5N97pz5zvm5qDb95Of+xQfNc
HCdEXIjONoYgTkwZ2aENMpZtrS3wHLkWnEc7wEBM5gSwCz+tBpfJM3kxG1TUhYRm
G76ebLyAWsqQAORsj/Dnd5y8wFvwa2Dbc2ICh84mEY7e6gZ3PojCwdfG0zBo6hPm
AuDdz0U0f1IGvAAGFR2KDVjCie7s31141XgqmHs0MiCS1tbrcOCUCvrWwILTST91
XKS1XlULMgIYbQoy1K84y7yYQi1dMFo6jwhsOQ+2jcBt15/ruUr6XCOejhGOSDZc
xRxDDlJa/aYEdrKSqfMXaoSF1eoOh+PLNvESUeoMLqOtcBmnz9pGvA+Iz2ClNQG/
0lxJs48cL+0T2yPBdhxmAl82BhvWKroY3UuE3pExMBh/cF8D+634RwfrxfVUSmdh
Y2vW8M7MgHmgvYMEeDDcT5+BngxMIGSZtdtAIXNaPEiqvFn3J+FW1RxIrLytSTmR
TPs3Tqv7MS5kCANuta2EAzE9QQm7WyjgW2/gTYIa8sCx8FspTVD3FNMnb9xFccfh
h2kLYggLWLYUBx1KLuGGeyMORcqm+Wxtt3f2LDPUWdWdpMOELmIZMj+VRuzaW9Af
HzWUXsRAG7CAF6P9gnKS5erIaMygi0LRrkKubcC4w9L24zT7+IaxBl/2OO0UDmEW
rum1MVCz7sREeX9Q98CdPdFs4iZprUbAim76BTjRJKmOwnFkoZirYac6U4pskkY5
yWlJkCXYVHI1VkBzZBsGxsLFqfwJZ3w292XtDIjnf1tILMIRA79VvkbJm2mazjsB
gIMUYU5K7G4dMMRzfZoXNuFt8J4VSKrJsmPZgSmhfWuS7W7bFvHUqapFWzrW/dDw
ewIoMN0p+UP6OSMnlwXizX92TexNECBk3/oa/bx5lscIvTyzc9kSqjxdWisOIANk
qtKxiLLRjNOD8RE1r4KYMli/Ks5W1FkwADMG/I0j3v1ojuMYLv82PX/a2G5Ry0/e
hujMTBF4IGVcLFdDs+C1r6WxFUNJ7Ml+yCTJRWqdsG+t2XZMbicsuxP+y30AuTu0
29WjCN/fbMNQJWlnMT6tl6aa3mgsmpdb6VjKcTn2i47oUH0p8YVYEkhycTa0hdI1
kyNc9dF5fudFJwuy7UxB6NKmjkvHPExM7ZNqu0vh938Au0b40g8yx9PnUJa1QWBA
ekh8zZ3bY9dvTij/RW5lUMkRirE7m+nVdsVcXNi2RE7Vje7U8IS0mBt+6CDNpNSJ
hOVzRR6oMu0B8VZEoszgyLOCYzFEu5aD3vMJD2HElM/012wvwdXZ+v5atKX5DO/8
7j4lZ9AB+EUSQaV2A7kPeQknKXsHYKSqg7NbRtBsRR8XFMAnfqT50HdsRbKKSwKg
FuV/958ZFuyuCg6TGwK2TQbQTc1Z1dJdiUEzZ6HzW1ob+plLUE/0CpWGIz3UYdGI
KiSyIFe+lxzNLwHk4ur5lA+ixOmjSYc9y8rWLsovmwiKOaIPRP2I10enbmXbF3+J
0dPG6JasW7dcF56osyPGTz8To8Ddf8LPkNrv025uETFhAc0tEKy3g/Q82UTeLWAx
MMGUeREvTMYjwKByA2GLk82a5zAS03ONiOEMwRHIrxSDtUmSIDUcH19yQBcTqz4z
/6pjk021vgXzSJJ56S7ZuO9wSL9XCcF9SiGXRwkP95m2nMR5oFNTRpiHFC/MnI8P
qJDbRgfBul6ysUakIO2q0zZWe7cmyhIlAlR1Bg5/OjAztfjU+c9T1KcWlU1sRra+
enAgKaoSYTIAc3U5QF/iwjW06hjNa5Jd8Nno9F/S1UbZmbdCWcQf9WsKBB1SA6n1
HXOi9aLXIq0c4bQYDfa5SGYotCoGc9Cyg39xinjerLfqwlt8HwbyYuYON+ZrEdaS
ld4zmpESbJlQ89cfX7Da+/3WA5asDduFRlMZ9HCaa3J4enWoE6tDhl9A3f95Bu2G
ySPJHo25gC8uK3TsssgsxjDtnskYu4LaIZ6T2jp+08dmmAKmc37mjZiv+8AMTRjq
IJKJ3Jdd/w89uikZLKMuqaz/D8CagkRCllUPE9xKMrU+GBgd8ScLH+l/Sh+kB1UM
jK9B9JXGKPVDM5f6c6jn2bz8gve0KfTJv13ipj3cSML2Sov3SQiAKbt9iDmzz5dL
csUliFuuCxGT0rXL9po9bSgRuQS1mr9oPMQstCMvBiEvS/l9+vlZkpHlohzhKHOO
B2RohUVddJ7SNneh9Y6kj/bk6DjhToRa1yd9j6Vb7fnDVM/z4hZ7ltu3W0gBT+hz
YhmUP7NXmoppZSQTP9kyL+sB+UVFyzoPTeNVIDbfRzFFTEV8jnj8jk2UXY4Hi2+m
j3g4HTkbTRIkEnEVvByPpZyBq91/eiPl/5XjXHdtFsRpGprALxu2rnqMq6Pgaopn
amOCdqlgXh+HN5OKqwusoMz+B9hv/9yB3N2dh2LXuanDFrNgfe6eebMyz7Gs19J6
9h1OO6fdPqxgNPoXWBGDtrFIl6Sj+tUgSZyvy8qmHxKXvpwdI1AnAP44PwyvQgTa
BE1d74gOsvmohpbQQbh0dZ9jLzhBqyzA3uyI0TkiiDDdukZPDeXl4ViflnK6RmUe
wqJ5PCSIqRN/E3/9ewnc4VC2JIJo1VMbt/xB69r/FtWsNhdSoQlgQ7Yx9EpRutmU
tqoE1/dKfrVsozSK73GDvBWGsytd68/0iz5d6L4OfB9L7LRhZ6douRUY2idB7b99
ZZG2AQZL43niITmQyIwtMSIeaMK3jM15DJ66RaA9WuOgWHw+xZESIaXqsJO1AkOP
pel6rOlqH7rmm6y40rs48D9Fp6/7sMundcufr7/LD36AgbPaxZFTU3DD4p43nsk4
sAF5EBdgIp5hksVo+9z3N+KsX6+wRocqwCOH4+lZNMHWixQhcVI6P1MN9/PCb/bb
FEePE9a1J5ajzeiHnymdU5pu59uJO3G+q9qPU9OHFsnGG5usWmq5Hiij5dcU7Ewx
G73d25M9+LMOmIVjB94S/DchJZvqFqPZ+3nYyhGeRjxG4Qf63kWxBMOTl4ZSPUro
QlEOe19FUgO7J4VQeg+4lUII3asfJ0cdlGNukSoi1JHoH2RxJVDX17z0vsG39UYR
voSIi3hijtpQ7BxEqfz0rtDNNg6+IAbT12V9zaj/HtMCvlJ8kxl4zIcW/NN6vfAn
axhDsuZKOetTnGvhquuUwGUz84+YMaBo3fujsvUNuiCoGFwrqlb86hhMsRvlXuFX
k3l/zEdwdjPHfJjOrSwwHoB09YuPGURmuR71br7ZzQhRaDped4CseHZ7KuENizMh
pLJpmkO3SwqcZwcYfzNB2TJD9l0bf4Xjhd0GjZBKB7WIsARNn9spHhSBqeMjqoVj
Cj5QDtj4DBDG/SeNP7ZfN1InOxzyld2bDkB0kpYJa9AflxWnlXdiRj0Qk32wm+Sz
3tEG1L3rbt0vcIf+r7bNW26fHrs30E1DvokVOLioTpFYFmWm9zMH5tFTYBqIESqP
V+X0RbbllBAz/v0RKuhFJf4wHrqFL9VC4BvSo9elnRp+NjwE/rBvL5MMyt0sjNhT
VuPppKxFwKTsmqdrUKTbVzzQ5lRoGxE4ZXVdStYQErGMNZFcHaXLOvF59x5KYBIV
eHkymWdtvwK+EsV9sfJ5WFfaXMQERWIEzX4mqkbnw9wEev1A0mdVPdb7OfukD65y
TEooOXL72MvnjsR4zRc4QAdBWuBz8xIjWZi+4rHS2M3c5XQFhBF0KvhqeTME1Tbd
uDDvixGI3ESzq5amSe4IvzuDKZMVOKeYKP6NrdKdlOvxCiQuQbJOuQnPOdzlH4aO
J5Vvm1p77IFL46ALQ+FvyHKl+TMo0zflRf+pkXorq+LJqYf9MfALZm71sO4/HHoY
xZloFAFs3fk7DIpBBccM6LmmXn0g8ibw2Izs796/5+GlQTehUwIBB3z+DUjHHilU
ixpAefQjGoiLP06k5AuLHf2W2xgOhvavHfE+h59nUAng5JLkNm/d4eSch+ZIXH/e
DlT61wjDTbv15+2RgA/dYIrkeozTUde3cxuMPn9mpJKMRgt8PLIDFl6S7td77xdL
GxvYnzBkiIFIzOVbf40caqSneRI0kUWuqZZzb3I9aGehgYfhh5H2Smi8RTABGpba
YAgB8j07NfmbK4h91OF4PL093bo7a07fUwbabAiIcwmNRblPqtJmnVH5WOyGp+vV
uMvV/XbAnjruHVHEP10wFt75wkce2tdjJbNXd3vR7UVezRKN/g6muKR2BUSL2+CY
NR9j18RFyQ0o+AlitQ/UsT8JnwgfU0l82X/OhXF42sU1ORA4tfeTOSxKCkEDL1Sd
D2xVdga7oc5mEqP3Y7uVhphPTTfUbNAPnPs835s5+Z35NF7CKhivsbBivj2zhOOS
KuR6JXuuDQpMqK38L3ILtAvyWuYfaerg5tchcSjgiyU/Fp5TX6rSduse/q06NovD
UOHCwOkPHPtrCQTHnEHlDIcSWhiwsvsoPDwBvrGTRIstiLXqAZ6jyqzNJV/1w/rR
p20VeWExQIVcL76x32ebPMwoVzU3v0+inDQ00n7n1uefdX6hfCkDmw7MMiZ4hz3r
OPpZmytD0DBHUn6K57rUnlV1du4iK30JId8x4rfosPyEXAVJ/9WQkDAdwQCiHVEv
mV/nTuqWlPfgv14Va70gDvuZKGUoViNyXoxg0bmNDVchQ1Odr4wRwbtIDvLym8wJ
qv9yYt1LFunVQViED+SXlm6/DaPwu9abpK/HjgHZOa/+T9Shbd3S/wGtp/8PuRHL
rg5UyB4UMj9uFsxTHGm9T3HqO8VugM9NuA2UVraEWiVkw7B0k/eg5R37ijCj/ZJP
3oug+LLKcZoUpiF4Ds3b2RujeGT2lIGPmPO1IUn44ZJTNoP76F108pD9dy722tyS
V1PYjxyN+gEOVbLDdwrgnGlOdcw4kSOKcbSxXosjmMBf8V+6MPr1k6g9zU2VJ7uy
2pS8nneQYYDl2GgpyiyP/9m5OYZL1Ajm3moFyJH6RsN36vctF6qm9USRGBEunWPv
YpUwFmtTK4XNHKbAYvH0rQKpj28Tul+c/YEYjTRGoPm4RfBEN3DPZFeR58JehPU5
uTTFt77JPEp0y2lm2BbUtIotr+GdwF/FHUp7/lyf1zWudQMPFXhSYP/xIoardQr8
55uJX2D2BxzaenS1JPrDk0mhuaS05eVs2xtREaulfFxWQaQa36tW0YQ/GaEInL0p
aTM0Yq+sxDyRuETc8Jf1m0yBdasJUytiWT5U4rLscVRWxYMjhI+jr+iVa4Nj7ssi
laSzzSuNg/aV2PRbHa6t1jxGGQTCJM5aFLRcx0qMEUX/4KRe7Dw6WAP25JW/OS4K
4/cimxVcdaIJ/W4OdxHDadual7cVAtJtZqawMn4Xx9oSk211btCb0T/KTpGqdXBX
Hn54CAlTXbejper+W4x2q08TP8Z/3PlBDNLveFuGQrshuzeNDM2w58+ITzIDnvhu
bHQZIju2asHArpOV3xscvX19MrTdHq8gT1xhzyDhY0Le58Y9lbITndK9fIiz6p7x
2TOPYE40C5NJIA1RQAf5A7M/xAzCAV/rZylY08vX6Wcx3+WR5EYmdb5iDPrLZ3/q
22YhEoBxu+bTLG8QAKhefzZUjnpsnvc8603C2NN7OmrYpPrLHbTtMjKtfZlowHX/
tObkS/UZMqMrdUxIHRa7GpwM4IaPyUhPHkQmNiF/yEdnDkq7leGkLXPLcKFf0Xvn
vhxqMQVk5s+z4azsbplEpe65N9fRk1+jOEuXTfma+wszurKZBJFFkwhPOBg/alKw
XA+biWAN0o5n0nBUUCw2BZbOAuIS1Iuww3AtfW42Mqroc13d/mmS6QTZuFuAnVwn
L+Atm70OcqVJ6NtvsaMDoHpsicpBa6dcHYwajHfI3Iv7kiR6m/O6OG29GTe+Rp/g
UT7xIwmDCz7x9hsa+e5bhg22o0XCeIqIUbOOhgLYrAAmxQzvf2Qzum5sSZwRldzx
SIyaUfRqGgK4QFWDzS47Dx1ZVVf2D7xCXo05U+mtEfgwvOnBW9oZVIDa4/utZEdv
xDF4L8Xita4jJliEpO1c0br4sy9Bc8mKxTpeTOWewrwpu0dDamlcix/JqrQvVpBc
TgaSX/ckd/ze3+4GwEHlcPhzyn5g5MqFYcbJESodYvuIAcfEMiIFD+jhVPEGn1a/
AB42Sd9udU39Grc+NRAGsZ/S/J9b1gXDtxdx/26FN9yY++B94DiOVvfchaCYRLmg
U5bpwpcVb2UiYULHnk4XeUOLlFDymMokSSu9+BuH11YOdkKt9VHK5bW9X8XQDWik
OE7E1d2Mcm8a9sYelnCBGE+bNJy5Z+VjjtGoDy+AxGet8OunDfPkdZbfqH+XBEem
/OeBUh0Jh823MTyjXAy8OEkOG91CRJzYaaEPH/sybmOW/26OjRJPLtvdD0Oujh/u
keoE4YGZu4KS/PUgeF+qWXscY4Qbf0HYPGuomAHLywA2zq4iZJ7MaLe1xR9lVWCE
LuLJ37//jzURJt+HaBeC5QCBLQQequk5Nu/DE6OV491MEuzmEYUybZynFQbSsSLG
qJAZAlIEgf4F7LDpR2Q+u8XqnUf03uo67c4rs2AHf5WxatA2uiKvNJ1N8osGSr4n
I1E0/4DO3ejwtJOL9sA8r/4ZlEiT16Eo7yB8tjq0gf/UHYCcyKnO9DWE7pwZPgnT
Vk+0Ft0lsMI57A0qdnwvfX1bLgbJz4UZMN37K/nRf6vjIG/DOidAKqgkQvC3kP7i
FhjhfRM/X7GRiA7idWW67hkoYzpjFErSOGtJOW7bA5zJugqy2BHtQcsJZwa3jxFd
mR5PowUTtXeodS6zf1HQvuP5TTearm/TaP2c4d21ohDGyz0jVaid6Borkxo2KA2h
ihA1mREbUWrTJanQ7mHI8fqpHB+QJz21ERB1Er4+Etk+Vy2oe26rrkgQjBuu5yCz
6QcFaS1Ij9HveYybqAQGI+CBwZOhJp0ba3K500ws1NpuRT9n0/0gbDj6kvpjBwlq
seB7iCu9QBbZ5NnWIIPt7j846CN3KT72MeGGBA2O62qYJQ950ivYxGAUMXdO3Nq8
N+vyyu/9raANKraOoCyIgVldyUASfEG5VudrUmGBIC+s3jpzkFcthyYXwe5W4XpT
`pragma protect end_protected
