��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�9��.=���es Ɗ��7:8�]��FM�n{��T?��m =?�6bɲ%��!��D��1.�y����� ��*��29=W>.1-�4�!%d�n��m�u�uK.Ѿ�ry�S���N�̇�Z�ৄ�B�T�x���/ck7\D�z!��	tvćh�n��SN:���-5���y|Lވ������fM@��*]�K��A5ቷ��0s��w`m<ř^L<�5�tp�;r���:G^�q��[,B������*��/Plf�a�Z���b���*�)����$_*<�3e���?=ı�A������y#�EH7���A�!e妉ZS؋�
+�������x�<5PtB�k/�[��[I4��R���a����'?�+�B@}ff�<������1Z�=(��I
�OFd��^o]f�S�"�`N��-�;Ӯd^�d��������}�#���uX�8`�f`s���g %��W'|��n�s;���)�:6t�L R`��;�fA7k��\�* ��d���@�1����;�e��#��lAnݻ��ϯ�sww��9��(i1^�P��Y�"w \܇�^�u�����:�>RX��|5��B�e�ˌw����ƶpD�-�v3+�i������ho�2��VWb!OY����D�)�������A��+R'蠥����ܿ,t���P(ګW�R� /^4望��8;���D���<�|�͙�$��0=x�"e�|���vS5PM�Gi($�es�_4��Sg�c���;��w�-����Jő���g��G�:�^��/���t�-.��l(���)]�l�ZE;���S���T�#�t� 堊�Z�
*������Zv$S͊%�H�l�pfW���C�OP7���w�
����H---�""Iu.	B.��æc�g�+g�G��/;�4�#ٺ�-�����g�8�� ]�)����_�B�f�#)�6�M}gR:��t�f�^�����w��`n�A����>��٭%��%^o�>��o�%n��"b�u��%Cz�l[8���ֆ�Ifkr*Ѝ���#�$�ZQ�Tk���0g8ʀ<����Y?�4 �/M��s�P���֊��	���s�평5��rl�P7�=�^�]��=.~�1ם�^�1#����:M�(��m��̗�G,�ݝ<���9򄪋&g@'$��C��6n�#%�h�f��E����8`/��φ����Τ�_=b��.�����ƣC��,�LED��nb+٫�!i��o��Ó���څ$�_��*����-|�|<�b��G�Q��E	�Y-a�n�M�3Q%t��s˹�r!;���l�ߝ��?��q�>�8�]z��t#i7�e�֝�v��ycv�x�i�bD<���F|��7	�٫�W�1�d�N���L����l���,�f�f#&�n�%���l��S����猇u^��<$-�iz�8�ۿ
yCpa�˼�~��
&`,*���a�~�a�_��#�����䮛��F�J�_�˗�� AD�:	�e<s�(�T>h��,?���Օ_ ���0��O��:�JN��I!I�R��y�u!����+�0��Ş���j��O~voI@�g�V�����V*w�
CO��~Z�_���Iz~���F�~��=u5�U�z�n`bu�Wk�7BCo��1�e��坅�L�>���I�i9�w��ۡ� U�v�>U�ҡ�R��D����m?ꃏ��hk�,���a��a����w��k!-�����JU��F�E;s��T��h�X�jfP���21�(hR��|��.�c���:r�Ncg1=��~��|1�^p�(rX�0�E�;>b�Q��[�`�����zyЧ����E.po�2����j�'����}�{�A�q(�$-r���<�9	�޹>��rvua��{���O��mǧ������NW��:�����Y=s��?�S)$c��UXwP�~�]Vn�K�a��oc�\�i���uA���4Z�<5��6��'��]2�����z����*��Y��"!L���K����2�Q�	m�z��N9�3�f����t��v�G,Dr��Ig�0.Z"��m1�E?@�ɉ�B�6����AO��1^�����JF����w����~�u�BW#��#Rԟ� ):iʡ���Y�������p_(�69M0%'��Yh\*^���\�<Gzf���kA@��~�M?Ȅd	j�Fע�w�2f�R�P��.,���`҄��A��u�.[]�;����#������j�	�+*�ѫU��]�&RlI�4�1ʴ�쎔c%�d%�a�V�k��]U���ѫ4hȠ�D�m������1
[V�R�r]@��X�]��$���@�ٿ����b4mEIH�v�FXoSD,���/�~� ����]�u��=�c�ٚ� ��j���'��J�>��.L�g�K���u�D��x�L��MЩ�#�ϭ#�:����|���6�5,1�E*��L�UF[����u����/���#���,]��Fܷ�>�y+�Di'�R�>H�z��2b�F�&�0��{�E��Wn��!���I��դE�[�Yh'#;������7�L�D^��8���/7��5��vӡ�Jε���T��B��l��K�2�Ο��~�UE�������M�J����p��=n�����7ߑK��{�������mE?�<,~{�Z\A{q�#8m��GBvzG�K*�Ĉ"A�c3}O-�����?�o�ձo��쿅b&��(� �X�<���D���\����@F���;�P�*u^^Z�΢��T+ G{�E�P���Cw�,ǐ��$����:k�s�NI�&�b�ܷ � Lh��BL��� 8/7�d��� �r���5��H�+�[̿�?���vF��������>E��6��=�_6�S�o�Y�g�ڽ��hʹd��߲%q[Q0��&j�\�]����NѠ��� �����u�4.ͭa���Yyh���J��2(��6���pq�����#��I����^�mNz��K�+��(+��$q		`�I� =a��[��M��|TW����������F����G9�^ 8����Z��G�nu��e P�|��}�VL����R�Y�f����N;����:j�r_7�0���7h������0A�'�h
,p����c����d�(�ŕ�-N-'V����m�͢� '��Q�-�/+�3����ܦb�:y��z���.1�֋r���F�䣥3�����jw��9�E�Au%��,�/wH�������OMLyGy��$�[���z)���W���N�/���ǿ�