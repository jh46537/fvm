��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��b*]���I��̞m��w^o;�2q��"dS��)����ɿ.�vb���t�WmY{,�#�����C}'-u��d�`N�'�-��

m ��'�3)�f�W���.�-∓��}����Ta��4D�=�����������扊K9WM�i�C�{�7Q+�Tz���)Ŭ��%c�P;�Kֵ��a�6�^�ӻ�r���f\�.�Y���1���xG�}��٦Qp���S˵�^�~Pa�&�=��8`E�JX��;[<�T��^�V(fI_�p�dt���6V��Х.ǲ��@
ք�{)�5=�G�M�lRI!��u�>����y;h?�?�ئ)6P��>4����y��f\&b�\	Sh������MN9[妓�G��i=�ɼ��(�-�%�W��}+��#ء��TT�xZ[e��v孵�jK�Lou��)��ϔ~����X(PD�+X'�h�z�u6R�$�2c�$����-�h�^��׏���p4���&�`|v�m��Ї��g�Y��:��.��}��;�&d�.r�2����fP���_�,�ю�L��1K|�@�#���ytg�o�h�IiyXQ��m
CT1n�7��>���2%U'	@�a��Y���w@/;���\��/���R�X�Q�����\Ow�4A8|����z4�F�2u�D�hn駣zW�%�JOヮٱw�36����F��iw6L-ɲG���9�Kú�?N�	)T�=���昅��Bd5�G��Es��O�Rg���8 e�� U�n��0�"ʀ�U�!ڬt�ѐ�7�Т�~{�92Nݐ|2�sb����iЪ��=jj%vU��M �.溹+C��}׫HZ9v���5m2�,�����-���X\�ؘ+)N�iM��#x�02P�
`!DY!���`���6w��
�VPzWi����1L�տ:��B��;#1f��8��d�t��y�f���2��(�Pdﳲ�m�щe>��.�n���K1Rt|��9}&��R�B?\\��ܺl��#�
��`��8�>�6����&n}$[$V�"���F%&�bJ�r��拌��l�J�oT�ٸ	���ؼ)!�����k��9��3���&���N/f�1a��$M�T�4�$[=Wcs��6��[�&�?E�������6ca�����61G)"�������uz�1
IU�H�/�R��j[�fc����ǋ��;��A�N��v���ϵد�țn�����2Ն^���R��x'[� Ŷ�%	��%4�2�4��o�f)�P�1-�����p	���VY,�!9�B��0�����t�����/�_����w��j;+��5Y5�����G�iE0wC�_ n"�U� 6k��]l'�j�}��cM�-��gC��I��ʌI�ݘN�m���>�:  ���v���M<�~
�S/���D�}�M����F��>��ъD��V��~�t��R�`�g�i�g�3$�ץ���&��?~���"6��XN�N��M<�D��O���@ǎJ|k��:b���ǅW�3���H�r�L����y!!X�h6>�u=�N���B<<���G��ִ�CC.)� Z.i����,�RJ;>��T�sZ&��<���А�B��;�Ԣ	�\�r�HQ��r��k�=�R��7F[�ŤVc��2�!�o�6�`rk}U>����,�T�S�	|�S[� ��w���,�}3��U.�7�a�y�Ѳ����I#	.ti�$��og��կ����n�ڦU��x�4J��~����_[��ܾ��W�o��(�3��ċ�r{l�P1���a����Ւ�{�Q99�p��v���{<:���u��U����k�W�����6&�U��v��c�f/���2o�1ʃ�Tһ�I}=���7��H����;��wpx[N����il�k��2���T`���
8���$M����}wj���WÇ�|;PyO������te�7&�^��J������w�c��3�ZG��siT��0U�|e�o ��� �P�@�#�����?P��c2|-�胏��R�>G:���7v�=cm|��F����|�va]����#.߇<�4���A�S�W%��
	\�3x�5��AVAQ\����o|�vMJ�S�<��N�S�I�����|M��[���������l���ңTe�,\��J��(�Bn�Io���Dd��%v.}�����kn@�&�z��ԯ4:u����l�j����X)��?+��ԟȞ�Yu.���u�S�	��ځ:Y��~3�%�tI�v3ȯg�i(�	�]���R��ɳ5�L:pRQ���oR�!O����/���1��4
C3����ӏ��%�5�N����@��|�.jC<ƫ,��Jsa�f�5>�q&p�R�׃2I���q#�Hy&ΐ�U�;Ø�	r��S�OD�A�F���.GOkTqn*�3�H�jᏋ9�b%�M�N>G��V�(4�س���J�#��ʚ�Z��w���h)��<B��Ђ2����!_AO��Q���<O�F��@ʒeO�&㛡%��<֨���[IS�����T�z�;��W���=�gE_�;����E��k��^�'L8�3@raC��Ǻd�F4�b�)������d"�=��IC��m\�۱��ض<�W�殦!�����f�8�d`AK�jX�ҳ�)�NI�Dr���֓���H��89��b��;r�U�4�Љ��������^0-Ss����/s�h��Ƅ�-o��T�CU��������AXUɎQ��X6{�"a��I.�L"&di&�K8d�ì4i±�Ŵ�Daބ�^/�h45v�y����5.�Q*��$�p<�j�® ��>͠�s��k��3b�*w��$����5�hw�C�X}H};�.*1�:A��ndF�m�mQ��J(��X��w�m����>����:rAFT�fj+��i��	m��Z�0^��`>pS�@YL-}��i�E��&���nH���h���Bn�i�m��mG7�+�G8�5#$���|R���yv
:S�e9K���u�vt���*�G�#c�2P]��6u@��qg4+m �3T���t.�v��^V5�ѽ~����3�}�?X�4��/c�|߾1��(1�X~�fU�6fw��r=]�'�jUC҄�b�`�{:r����i	5.��'C~Av8�UQ.1!D�֗)k�-��uBC��6�w�`�0O��w�e�e�My}+�D�7�G�uڽw��Z��v������k9{�5���OYR����Vlɉ�U#��):]=wB
�皀�~TI�����}}�,bI%=�=E�"�ek��$
~�5�I�� I�P�Q��[��K8G����s��}Y��nq�S�/T�&X��H�Ǻ������Liӯz�����*��I1ݣ��U?y�YC�+\�̻j������e�,�y�Ǹ�%3x�n4| W��4%,��̻/Hn��S���H񳳧Ʊ/��<�g#�ο��1����	�bG��,�z�uq�Q�U�]ҳw4G���b<��ڐ�g�w���Ȑ�w�G��4��]|�V?�LVܙxF �:�����#'fT�S43�V�����~���s5�Y>'�~��0/$�x�/-��<��7(�T�P90��}%��)���L�Q- n%�b��4ʿ��{���:���p&GzJ���v��:/��2|T�K8�\��n.����ɰ#%h.�H�l�q�wO��p${�d�[�A'�Z��g��L��xh0�>c;����H�~VBO��<���=(�c�O���]N�m\��}�_"�_=��D���w�YO�ԅ�ɽ��/O��A�\y<�a�ʳTk��>�S<��f�� ��M����UUP��D/>h�����w������r�l�zg���XBS��sG`6u��YyD&�����hh)�ǀO���|[���[�L�B�>3̷����EDs׃��n�h�/�f�l04�N�պ��į*j��sr�ۖB�'����z������W�;G�a�|���[hw��@��/�?����s�>V�K���aAX�B/NOC�~M�]�Ekh�b�4ێ�r1��>3wX�{i+_�{�p-$c�=\g5s�����zZ�+L�|!8����r#�⋹����>w�hJE�Y�>������~"�f��F�C�u �n�4b���n�����g��H]�Ќ ��?�D1FMT��� �:V�ǄE�#�G�z<(I�»���pq;�?�Rg����������P;�ͮ
��4� �%��U�ǹ_�sD�+)���U��_��l\T��%̂�M������e1@}��&G�@��칡�����Vk���@?Xp�9ö.SrvF]2�U_|R0�e�񗪗�����6m}&�g�r��?Ox��Vs�`��-{ҷ����|m�����ĉ]`TM�P�k�*���UZ�x�zV:�D�!��t%�+V��(��\�l9Y���	�^Q��M4%/�㜀 � =C[BT�-���7�9��ް��w��D�?������I��ǯ}?/�{1����C�L^aS����}�Z�%$���z�&��E�r��Z���J��(I6��+��1��N���
&����TB.o��Р����(h���><��I�u"�=Nl�]��=���vM����5�q�������0 ��.H�~�ckF4�=���7�����uޮ���_ӡ}�R���# ������Kؒ�C˕F�"��j��Ŭ��y����9�O�E���j~������`	:��!r�^-C,~���e38�Պ��T�S��GpË!����Oظ=���ѩ�ɵhLC^<Q)�f�10��"�'�E��Ê���*~�NI�ߜ�
ǈ��^.��tG��D-�B�-�2�,��.#`�@*�L%���E�Q�	�f���U�.�'M���]��B�1�cz�݊�T�u~a����je��.�ϰ�[!ҽ���xY=��c�{�igu]�� �����z�����@\&���8�t��}��}��#����b�S2\���BO�W�Y�-vI�ɐ��E�Dێx��Ȑ�@)���l�Vs}�k���pt}�9Ө-\,�W`Κb&������T;k�����Yő#0g��*�W{�ԥ__����wCĿs�E�m��1�