��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ���>d���G���o���TOZd�A��-��+�A���e�#p݌��S�t�P�1��7I���Sr�742��(�B�'b��q|�6�* D�O��'B�O�L=��y��,
��k��b�@�^��ۿj�$�ftp��/��� ���3'�F�� C�n-�#D��lo�����IHE�z��7��Z��|M��1�<�$"�c��� S'|BLsu���~�O�@{��FW���A�5�Q�=��<a�OL��x�
�r3�)������r}J}ނ�C��v�`a#�	ukѽ���9r�:����9�3>�W vlw/hQ�i������G�a����0�".���b���y(
�+/��.��
+'ҁ����E�������I�;��,ܨ�%\��G�z�!�`�rE�Wϓ�MP����y�u��g���i�^�F����a��ƛ�B�o�H/:�Q!��n��2��Љ���w�����+j����F��"�
�Ӹ:�O>����~���e_D(F_,���AF�i^BEwa=$�Щ^h���i_�T*I}���3\I�A��wv���t���l��\3|=��x�w5]K6�Y!���Uz��!�9>�e���v�;b��L���*�	���]W�ɭ���ܧA��%�-w�Ɵ��X%������S�<̢:�Rl6�����"���?jh܆ �P�D$���ϵB�i��3��ZKu���9�*Ԃw��パ��Cϑ���Gϳ�<��`Mɩ�Jb�[�C��MV�&4i9-��"hM�(���C 1<�8[�'~ҵ�����M|��8l���� Kؓ��r�ƑwlDõ'6K�+��� �V�'��Y`�;O�<�O��R��u�j�z���/B��lk�o� �@S�n�&��&p	w[��|-3.��d��V2���8��5qy������������/��1u!�.:E����~����G!�3�Z�8~6���X��T
�d��M���0j�A˿'+{����KC�7zP�{�a�+�͎��T���N�@���OD��0T0N�3!�HKvq<����>�����	?u+���=�̟�m?�n�n����x�W�A~�o�����l���8�$FɮSy���E_\��-�^�y��/�@���!w^G������\�&G�$ƕM@�bf,h��:���N\���"g�1{�ϕA��UR&UX���ۈ�b�Q��9D��O������R�����}.r^c��L5{OV� f�1��ʳ�g�K�4»L�h�N�;F����2 � �m�"����n�	�(�S����I�Q�g(�J�c6ڴ���g���|o��l���&�`J}+�	L��H
���,�u�6ѻ.L��6�C;Fϕ�q.��rF�Z���,�FN*��,��	�qz]��A���(7���/-�߫p/&?��|ul�{��f1��*���X�'� ���k�N�*@��xA���L��a�3/� �?�ͱƇl]����(o*'��xx�Ŧ��BĈ����)ҋO�$�f�;�d�RP�SKm����a6�����>�Y�Z�hL��/r��q.Q�F�
��76XAv��v�lM~����/�����M1<�����Ӭ�c�{P��"�i���5�Y����k�-����
�Ѵ<q��:����ǥ���C'&�� �\m���6���(�}"��
\����λ0��Y��ʿ��Gp��AG�q���ǘ ������*i�ѸW��c<��
^����Z�Ƹx��[�#���)u2j������y�c(�C��9��1G��R�\i%�̫!�uOI1UDjC�m�1Zܽ�,���6G�O�@ӆ2�� �q ٳ� ��W���LUT�'���s���mﺋOI��f����W�����^����7�y\�#
�]s0$�AK��n���ԁ�%��G�Jf}��k\��;�YI.c�����Ro�A��ۀ]zҶ��I"Q��]Bs���׈��m�(oE#��6�ȡ���T�A�QP�[�!~u�������5>�3��Y��.���	\g�3aZ��Ҡc&�N2�p�0G�����o(�i�Sp��r��v�M��G�Rt�"��=p�5}N(U��F�;ѼX�:�j�=!��=�y���G�2����.is�ͭ3ğ~e6	��Z��+(���΁�֐���v.�R�sW�x�#e��N\�s��qf��tҷ����X(�&�4�ދ���s~}��b&�ԇ�,����?p���FIKs���̃G�;�o�W$2���v5�}&h��Dno�!�b��(aP�[�	U�pG{{�t,ڰ�,I�Y�+�e<�C\��
�����p��o�jN�R��F��Ni��9�~�hSݫ6fy�fq���>�ۯ|��7.�?�Z��cZ@��~���N@�ΕV�W��B��{���&m%2��J���,�!h��#�и�ɨi	I��؉Xy�e�����x���_z��YkpC,?c�h��J�����:ѱ�nG��`�6�%���=I���F�6ӫ|��sa.*
�&�e��|����+Z�����,�'����i.BIy�u��W�Q��[�n�e�){�?<|}[,�����_l��oY9�n��1�m�*?�`�ӎ�$����!�!�Xy�i�-��{Zw<�ȵ�ٷ\s�C��f~� U��U�+O;D�1bņ��nk��lm�:%���z��T�"w�ߵ���q�Qb������.Mx{' �V�Hs��Dw,��F�ꟙ���Y}�ng3i��� F[{mkm2�e,A/!�*3�����H0l?7/SP�����������ۇ�α&�`��0��Ώ����
����o��p�G%8J������0�L+hT�D���[�}j��H����^�Mx�(���x�3�B��jh�Dk�[�3�uʰ�Q/�#U>��N 	�xvZ��g�"(��
9�f����Iq}�#k^mD��Y�V������6��F8�T�����~4�~b��?Ig�c���E�� ��G[;�9�o說�yni70�b�Sw�H�F��ޖ��C�����`Оn�-�>|�F���,c�� ��r�=[¸���@��L�ܛN�H&<6�Vd��o�9�o��`��:QIM��6��3�09�L��H����=�GԂ�bz�c��
bpP����ڇ�c��5�n�b�qjE�2��d^�ڷ�4P�3T
(���7������f���B�ߣ��4_�!��ￄ�9��ڇ�	{�W4�����KzT���a���S=O���dS77�n�!�=�ZI�^ԖƋUE� ����b�T����/��G�oG�+L;T�<w����$qЁ�{!��f��o&�+mO���cc�����0Psrf�e��A�$�':e1H�"���Ǆ���P�5[q��>e�V��H��!@T�n�ZT���@�R'�&���`:����K�R���
���2���i7>t���q�o��;��M츖)c�8���d���Pd_��!X� �-焆���#�U����6Nc��ϧ�ϡ����_�����c��݈F_�^$�|O5��x<.#�*�����E��@}mv#H����RkB��`}-|	y��K-P~�1=��Hb��H����*���-�4 Pp��~j�j�zݴƾI8�إ��:����I=x�� ��sF�&�O+�Il�J2�t�����p �~'4|�ok���	6�6f?����^��*GT��$OU<|AӼ����<�Q1ԅ軋-�����l�Q8�!�PF�8:��l���t�U�O��D-(��q����e�ېدT(�-��Vz��B���`\�懘o���Z�=b�r��-��ae��#-����$��ff�7n�Q+����B���|I���D��>��� t�n"0����W�m���n��F>�ؒʰ���Rpr�*n80�Q�I�S���{ڭ�Eg�G�0�8���!l2}&�b�c��Ĳ�,��
!���Z-d;J���X�N�#�јA����<mt��&�$�	Qq;`Kx}*4��d�XA0&�rOѩ������m�J
�(ÛT5oȆ1Z�),�m���by��a&�kj���ڲ(L�b%�$;���'�yH����`ϛň��X���tE����S�dˎL|�&��n����o�
���G$)��%<F�&6��� �j���w/ҮH�,�6J��(}�یK�"���@�����P�4�@36 �d�	<m�����p?^��iV����Î��Z[�}��_gc�"�b\^��I&1鶣6}*jqn[b��V|�Om�7�����Z���I��|>�D\_�R|h�X�&Jv=,����c�X��gE|�A��?*:TL�OD�>�[�)��x[�Hk� 1>uѱ\&��7<hK|9Rz�����:2j�BJ�&��^�7:�$�\�dF6�����)����4�`�5��5�cl0�q7�X��U�H�j3�6=C|7���S�� ����0T��h*��Oj��_�t�CmT+ߴ��:� O���H��~�P��yFx�<6>�=(t����,~`�94=}�Ѻ�k��/��c��˻/���254_��/LL�?4�)��p��J�=��.Z�����	��-��>>�9RW�=�Ӓ��C����%�E[�M�^��K�NYH���2z���4߷�p����ԒV,P+T�A`B�q2��2c��
�qP���nW��]{�����OV��=K�ftߴqk!c�AD�X���ȫ�k>w0�y�L@�t�$��I�]?/tR#ݲWȻ��}�o����w?��G��Q���z����=���[P��K���s�ʠ�	r�0><F��0��r�;ce2��80f{�a�2eͧK��۹`�Pd�2��K�^��4�.�I�wz�$v�ª��R�_@�(�����g@��_�f��,4m�ڠ��'=b�%��zm�R8n)�O�q\4��������Bf'��|�}�� Ib׌�H�=+�g�����Q��ԇ�t�(�N��tI~���Z��g�@�9�ݺO%`v�z����ھ�RϹ-�Jo�s���!��h�ϣ��>~� ��J-�$-� K�^���������X_�,rlz�ш�_�� S5;��\�Lj�Q{���� lJ�?_EbMм�u|�O^§����볭�����}�N���)oA讫�| v�W����K��^���Bӝc!@@���:�fk.��4��Iy��="�د���E�l;����U<'.)���zɳVw��U\���96!����\? ��s���U��g��iC����i@��h��i��N{Z���[�K��0:#�C��'�����j �#��x� �r��//�#i��� U��h̲�����֑T� �oV�ZIf�h/�n��?$�*�l��'��E�Z�`�< B�c$�����"�����K3����W,�!'�EC�u�/�L�Os7:ăh :I��0qe?�$H�U�i�9 ��2E�{���֍���Z�!C3R�SN+�;˓�;㺹��%&��y�(��)*�{^�H�ȱ�C�;V:p66c8���#m��Fuэ{�����Z0O^VKt~f��_U�e��PZPާrg2������L���&����ٸ��?�݊D�T��N�Z�U�# ��=��p�O;){wT�5,�b�C���`��y|��<�_����)��S4�_�6�j�؜Oc�U��1*aѠ�v��e9���j�����r*O�����#̸���VV˂ŧ�, ӂ�S��Wx(�lz��n���ʷ`���@5Ɇ ��6��bP�w:/��'/V+�n�d����|	�h����>`Y'��!�k���B��4��kw��5�3�TCL���dͩSB�~����6k58L�"��1G�Zc�Nz�m�7|׵L�#�����-Ը8X���FQUe����	����@����$��5_�Dd�Q�`�\������:�v���Å�����b��; �|ʳ�Rl�{���ִ�4�
��?sW:�_LFm�+Ҟ�B�T�I^9�aZ۾_�˟9�p�F8�]�>@>/�����	[tғZ��B�%wA�x���> �V~�������SHս�v�2V��Bp�"T��w�T�ʣK~�B⸎ه��m|��b�8=	CF�o��E��;~H���/|p�xM*�4��S�XA�lɷ������4�ʪ��QH�`���8�ڮ�.F���e���;Gs�\�U�ڙ�`�9�k/`��%U�����0=%ۯ7x�H墭�̹��7w҉<���a��
�0���Oc����mr{��i�Y��-�D�ez}�l(I���.�[09���妇k}�uA'&G�KoY��bG��%�)(e{����^��,A�tp�zP�ӫ	q�%���ੈХ��wU���5����I��R��P�O�y�dQ@�����5�ܥ �V���
��;���A�)Sh?�j��uO0��\�O��Q���!��OM�f��3�m�*���*}� �+e���[����+�����z*K�΃%��nj�V�
��o9�m�ųg�z��Y@��D5x�QA3�hˋ�y��@���M0�/�/�����)jz"	`fq{��W��6h���[<Dܙ>k���5�GU��ل�Q�E8�Kԩ^}2S�lқ��4�Z�~
�/7��@�S���a#O0��Z���RSM t6� z� ��z�H��-�=lʦ��A�������}�N���B^���Nұ������pe�����R�뢉���Y��O
���G�����̐�H^�S�������0��P�E�\0qŇo��,�9��[��,�Z�Xyh��3xFS\�:i�Da[˦&�i���c(��?����#"� 3%?�ρ#����ә����6C����(Q7dg¥�(;���{�c�b\��(N.�Բc�t��m;	5���{O:>t	m��?����C��M�<���]�Mc��R%����"&6`�����V��hB؉���Z������o�\�U�x˧MD������r��z��'!e`	�SJ{�\KWIX��g� �xy#�-��v[ߢ���9�ik�w���.h�24N}���\��������.��r��*>ԃ>��Q\�*c
 >��A���D����(9�j�]�vPl��;��{�ՁU����q�G2����w�k8��N��	��Q����Q&hsLáw����:-	

��]��k�/�2�b�p�Ҵ]�`��b����-��*�ՙDt�H�wƄb|Z�IP� @���y���zv�_�����畨���:�%�$��Hqzt��5�z��:
®�TT2+�:���0�.)�KF]Ă��uh*t��e�*B�p��գ�O�q=��\�b���h��R�ل�{p�rfx��7�I"Y
�p���.[ذG3� 3fNF��y�)��22]C�n*�I|�*�.M�qDs��C͌��}��<P���V�l��Z	1,��d՟���Eڰ�܈�J�M�$��ϵl;p�@)�	V�!�2��(-��/�X��M���`&�H��S�x��Y\+;.�ܗW�
d)�2�j�Q�^N�o�mc��lo������.'?((7�\Z��cv��+�1��(�� |^�ե�r8�M���1nHOȌ殱(��U��՞g������OI�G���N�{���9$�s7����ݔ�v=0��hs^�)�����bLz�cR�y��	�XS�N��O�=o����`�MU��v%��x��`��gϭ�\�:��b�A��B��Vf��L�3<͕f2;�AC��S�6����$B�ޛ��؁��(�l��8�(x�̀�����m}i�4�ے�h3%�|,u�.fcy¨�]l��U��Nk�Tc��2�l��!0�u�N7q���6^zIIѽ/������ r�%�<�k�z�k��D��C�=�m��t��I{y���n���A�W��c���h�d=IHo\��߷y�@����!!km�}po��o��D (���^H���‴}d�l�9�g�F"�z�,o2�/��p�]���F׾�Zt�N��	\�c��[aR�q�R�Q85݊$�0!�9�,���Q6���h�@r��ء��f[Y>gXU��am�[�&L@��ǈ��hr�O`0������1��qa���&���aG��������"��S&���:�@��*"��T�{&A�FjAލ~���$��K�V��qJ+��>
��/i�`:��@[���F�Uԥ�$���55NG�\hm	O)5P3��D�!ŚJ-4��6�hc[*���dB*���Ŋ���K�kr�'3�{
�f��E��3E"��2s�:|�s�a���w�䘐�-Ӡ�[ ,��]�G_@ݼ1�|��E�Z�:��S�1��殥���7 f�UO���Vif��ׯ�(vߚ��$^����st  ���e?+��y���r-�u�7��H�A�|�/�PH��+�G�Cf4pո���2�	�^�?����{]���0"�$�H�\I��G=os��2kD��nOc�]Ηar䖳N�g�\s!m*�d~�nǥ�%)aP@_�d��dd��2Sk:�,CH=�rK++�@|�[>+H�������R7���Ms�n�G��݇�p�|����7�wE'��ϳ�a�+]����94�5ۈ¾���hWg��Q` ��^~�*a8����\$��@���F.���@'RI��`Z�ڹ����C	��5�l��=׶%Y�"u])C�QsY��ݧ';�c�H�Q�	Y�5n��Ӏ�X��*�hѻ\<��	�Z+}�4�m2�dó�v���^C�p}�������F�"�}�*��K�w�j�[�&���*z��~g��g���u���&�ep�Zz/��}���PEO�wI�yDT�(Mu}�D�f�*���IV2=��e�Ό�uyܵ�Kw�.��Y�AÚ\������$,ў{�W��ԗ'`��O�������c��n8,#���c��ɼ��v�_A)k����:j�cC��RJ+�	�<��㛶�w�t���b~�8��c/��q@�m?@f=� :U~z�><�>�$D�#w5��s �7碔�b(XnAU��n�MQ�:���K���\Б��]�_"���H2���������D������� -��f} �aW˷T�� -��t�̍G`�`��n�=^��YУe�2΢y����5O�j<9a5)�m|=�Y�)�����+����W��STIH��9>�'<?�<�o�݉�6�h9�Р"��z�+�7��Ű:�8X���7�;a������AW�Unڃ��?A~������n�"~JBm��x�`Hi$��hj"V�d`}�N�u���F_������5_�˕jfv�p�|T�wE��&����%�$��.[�I�����d30V^���_@c��7ؔ��!lǋQ�@/HIYG�A�B�)�L(�dM�Ѣ�kh��A��t<9��+'�9]�Ѵ�:9��N/�$���֣Ėݝ}m��*���:[�(����� o�	l����/x��q�-w$׮`�+!��Djg?o���M��f����AY�	�{�ZÊ)z��z+�7EL�) �a���3����o���ˠ{WO��Vc�6�	��dh���)�ʝd��z��+����6TD${�Q�|e/�G�<�K��IK��qqHp+ق���\�E�qY\�����'�/�?(�1�:G�Z ,���cZ����g����-t��B"t�u�����\[�;iݯH��<�܈�]�����U�F��0Nw}��;@GFj����l�����/��Qs�ә��E� �(GH����� L�z�ϧ���`�1\$����Մ��yD������U�����Y
#����.s;����~�U]��6�����H!���Cl�7�Y�R�.&U��M���z}�W8�u�dMD0�p�TD��?�	��������ja����/�.�لfO0�bT�q��,��{*����R��$�AcE�h���"�u�M���J�L���`�#�/�p�u