��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"�� $WժOSp: S��B;�V7#\�n=���I�-l��]ɰ�����O�)��& �4~rS�)�iD��3p��'n)��`$I�����>�Um��N���Db���	��$����H�K�k�ӈ� 1+Ez��2���k�}���)TPgM��E��8w0���y�԰1� �+���a4����O�M�?���*E:U?ADcS���yv� ��YaYl4��d�_Gdv�w�-^�|)�mD��
{,y����P=���|��%i��>'�'��W��e�\��1j�)ڼ e�n��d�u��k�nV�v4JwTմ��v��zb7G��𓾏q14���6�j���F��o��V�\�j#w7�C3�9��G~U(��b�K������PH��9$��$���\#U�u��G���KZ�vY�O�n˅��r��kɷ%J#���2T:�Wɒ:��f����T�o�=���]FZi5��h�q5%�^�`��nE���]Y��G�9��KHw��1��_Ɏ�[7L��:Y�)���.��$��re���S����#��!g����`���ae��poC�c�sk����#��3��YYU�ߵJ���l|����J�ޱ�;\2EI�͏e�	
���BD�Hr�f�%�^�%z/�N�h��~�Sd�d�5~�|�ρ�r���m~�����yFy�ә'M��q#yŌ2#L�����+��~���N��y_�.�`�$9�϶^��Y\�L�Q<OHG��ޞg_��=�H뻸sh�W�K`��j�����ؓ�ʙ�ݻ��[��B/��s����R�w炯�7 "=@�׸����6�C)�	vP2��1�#5��o�"� �����p��2��c	�O�T0a�\\d��3���w�~��lӑʪ B��E��\�O�*H\-t�J��-o���&f�[�6�ӷ��8�gv�A)�"�}��F��*�0$�s�����Y�#Rh�E׼��<�T�N|�d��nH�/������i�^̖n��߉>t�ρ����O��N1}~�!�Kɑa#�زʾ��yQ�e�r`tr�:��R� ��@��u�6�VgF��3�d6#)+4�`�Zi�)5��R?�Zځ'�E��70��
 O�w:�g��`-�=EJ�N����MQŘ�k��	 x!�G�7 ��6g!7��C2<�H�6[��h�xW.C̱���pƤUK&;��z�~(-Ԃ�4�78�p�X쐳&3`���:eɊT���_*yaoZ�cO�sqy�9r.�ݽz��ܩ����B �*m�@���bto ����şܡמ����E��m��P�'���hΐ�C��+�>¡���,��Q]�OŤ��pJI�Y�
-#�EP��s������;�u����z�W>l����6�{Ó��J3���|g����T���q9�ˤP��3� 4�ye����dR�43w��;�'!�����9C
č�*�		�P�20�Cz�5L���
N�K&?TF;���[eaw���5���#p�����o1
1���*M��QBkE�x��z|(r���]��}
d�U��pQkpPC��C��