��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbT�L�!�4�ؼ)�Pf�V�p�[�PIO�%�e��
�A� �ǣl�-������[��ȘX$d�u��o᪃Z��a6��y�� ����˻Ci�^U?�O�����u5p�����{��������9Q���]���b���a��FQ��a�}pr1����=w�����^�6e?;S�m�����!*X����Wf�(Aw6Y�.
�|d:߷�w!u�aQ1�Үm�V�[a{Y'�w)uPg�I6�gI��&��@)_�E@��g�,9���G'�y�q�"o5�Fǵ|�O���z'`�X4��xQ%���޳�sP���2i09�d���O��9�\;���1����[[���ަ���,�=�f��)]�0�]��>��#0B����@��*�U��W{Xl�i�$�Pp=�4.�AM�b>��&�6���)�/7�&��K���Ƽ�W+l�]�_K/|tG?�IE���s@�N*�k�=p��T��Swn�ޤ���r��'.d�!J����ջ�w�oaOo(�l��b �g����*����l"���חO�e^��ޕ�W�Ϗh:�h r�����_9�fBװ��e����}C�7�� �}������W��%�L�r���AJ����GaMe D�.y \p��T5����鏎�La<�2a�{���u�o�_�ד�O�#�n�~Q�O�)E�)V��^����iYܠ�S޼���O���:�x�HЈʂB	��<� ���h"%���LvN�:�8���W�36�ͱ� 9���`�H��QIZ�@�w@���D1���0��r�?��p���aZҵ]�|��,3�-�g�x�AT��Q�eq䆊�q3��w�� m4!��? �u_�聾�3�XM�ߊl	�ধ����aW�)��#�=�����I�s��O�Q��2��u&��bY���W1���V���~����v���3��Iީ����U���U�,���������Mk�����s��с���w�`Bg�f�e?Ao�f�ZS>*WBaq�������6�9S���$ῴL��?U�b�$p����WWV�ؽhű�W��*Ѻ(Z�����8��Q�	���nQʓiO>��ojė>��B	�?S��
sys	*@A��-�b ���w��ITU�������������P�ht4��ɻ�۲�\Cl���-�͸(�`���v'>-*��ŵ6�Y(�Vȿ��>8IU�:r��8�{��ۦ�'$�y�o1Z���FA��SA�^����X	j9l)��7�@B5�2a9���a(i8�g,�(Ƙ�-za����LJ�a ����N�]\�zi��'m��<t2�߳�pP�@�(/�pm���}��c����Q)�"� JLۃ����9�Z�Pp1bHSH�ݻz�PW1j�����S��/�uK���Bw���B�D���Y?�o�阪Κ������[���H����y'�(��Ԛ �mI�%�½�W�E�;Y���J�x��,s�9�m�+Nah}�M����'�Z<��$��;���к�ƌ�&( kd�m[~�~���R�:�W�g� %E������եu���uYE Tt�.3){&��ܯ����lf�s����r��_8�8�' C7r�g r�g3��8�5/8Q�E��xI����|e,�!��?׹4a!.?~HC�f���B��iO���-V^;�+�}�p�Eh��|�_�]�Bȉ��)� G�RN�^�{��ʌ��e:���h<T2�)l�<&�(�4:�G(�EO���3oB��l�������z[��QT�a����W�ص���_[>�xu��� �� A�B��Ko���3#�s	���]�=(�㿕�g}r2�r���R3�݆��!�P��:��ukcE�"���V�94[t�%�i�=�%E�,;wI�FE�ȵ���X�n�V���^>�r�&L,)�/�U�K�jGJ�����n�n"<&��ʪ��0����S<x��6"ь��(`�OYj�~���$h�R3S��9�l$�����
�4ϩ�
�!�}��)��І�>]>��{�:������6�E)��Ab��sAn �b��䲽r��T��n���쵰��,q6t��/!�����;�^�0���iNLˁ��,�S�L��i����Xu�pZK?:G�{Xc�*ӒR$��ҦN���0�(h�H.!'.c��z?4�D�9R�Q]+�_���mFF��+��� 8�����
9-��u�0�1t�Ч��d����U�_������Z�3��S�����i`h�r��2U��s��!ޚ\�3��-}n^��8|U,���c��	R-�L^���B.&��K
�w�A�٘cdZ�E�j�n���U�կ�а`�@9�%5��T�*����q��Y�� }��&s��R�_f(4F����\#B�v��n����6/0NR��>�$H<ڸ&��v`�>�/1�rD�*��% ��:!�0rćL��b�̾vl���]W/�
3�)�?f��ۿ,7�]7jk�"`�}_3I�@7�À8��Y�VŘ2�(�5wt��^�_uW{}��e� ���Fޘ�d�$����U�	�@nѶU�`�VWS���LC{kN*B�<W�wNɱ� �U8l��_7��R�J&Y����?z�,X4 �O��q/�f�N�̱9V}�4��vP����<���yl��*%���j�Z{���M�[C	�?*hݥ�~��/��F'.����j\��Fb;'�����Z��֨�IN���u��4�\�1�_$DI�f}z�ـ��R�n��y��KߊV�{��<X�Gػ���o�uV�N~�kHqS�c��0�M�JH����kԐ�ܦ�09�*�a����zK�ڣ��YH�k���ǝ�� 3�Ô�z�g�֞x���xGa��P�.��iͤ�W��U⬟��ٜ�*�J��0n��"F�{$�$�[ϗ3*��,����21����0wa���.`uۄ�����c����c����ǹ6zPf�y�<1xz�3�f������FɅ+��⍴����_����T���'W���M8��0��^��=��F�a�hL;��]�F���u�ф�B���v��o(W�RA�Cb����{��S��[���U�d�W�S��h�����
����.��W�R��)�r0J=�mԷ�rw�����;���@R�$�v�=�&i��F$��>C��:(0t� �RT-���y��5�ߦ��B�g9���u&pn@���(�,鞢
����Q�Λ�J�02��p�m���k �����-X�R7=8�g�ONVZ�=1t<|�ڴs��9���X  t.������
�rn��o|��Suf�~�����ѕ?�G�aXD'�L\����3�kR��m��a����ja(����L��A[9�����1?����U�\c��7k��2�Q
.0t^Uޫ�[�t�UW�8h�$���9�0�gVJ�����>	�G֩�2e�\N/	�̔�AY»#/�{K�K�Oc��|M��̓�cJa0E�/�.H�`�lt?���}ă� ���L+A�K�1�'3�E���7��ɭ(����,���M����Hc٩}Y�"� ��g�?Y�f ;�Φƈ�9�
}�M�%*��BW��U�F��&�t��<�\�A	���2�/䚑�4�3���vy
m���d���ֿ��<)��b8-v1G0)������YȲ}�iY�«������v6~�����ˎ�jH��ʛ��˚�������.�H٨@����qjbs���>vϛ�+v�*=x��أ�}$b�Jd3�1teU��B��ja��$U���G)T>5����Ooթ)4��M^$;aq����ܾ2���Y�������L���
+u+�!#s�0`�����י��Ed�B	�J��9# ��@d���?�7��Pn�������Q�&ek��^O��h����ӟ���n�Yg���S��zk�g�(��^�[����M�? ��5��|�*�)uS��Mt��g�~�����?dr|+�ϭ�ϸ�W<�{�񍈚-�LR�N��i�����T2�	�	�R5&%9\T�z����G���X���K:rn7;>�i	&`�V)7h���;á�Q�{ 8.���	��OQ%!'�p�TRҾ� �w:�^/2E�C���q��)���:kɀAi]=����=�RQ����3�93��W��T^�@�c�W�����+>Э �2�H�u�h� ,T��ӝW��4���5Ͷ������rns[���Д��K�f�r�5g \a��y�p�<B�$����}=�A[�p'�B�F�D<[��j��UIup��0�$�p��YG7���Y�HU�?ъ�\����1`��v}�g�&�7���\�����?	y$��;�_��ɧlQ`��??Z��DvE_�2i@&����W�r���
-��Q�r�JS�җ~�QA�86���J���8k���*�S����4a���u�BG�F���tD��J�k��%���O$���FIP�ߗL�M����w5�LȪ���kyd���]ݠ��.�������p*>�E����	^��2U�И�,�-r��~'uhx��K.䧶1���nս��ީIa�� �He^@>�b�}��].�O�ZT����Á�=ug��ƈKE�e!=�r[6�5���aTww���J���>�,��Y҅@�ｇ�b��U"��D�Q��9�L�ͨ�{YW��+vz��31�	^�eAPG��D5�~?I�b��1���>��3t���ΒP?8݊]y�	����:ä
ހ�}�Y ��"=�W`=(���)�O?�O�O'O~1��՟�������M�F��E�JUPiMq$�D:.��k����(|M�m!����:��3���.��GA��P64� �!��(FGЉҫv4���;�B��+Jd׽�{~6h�c�s�Qp��jc��:�<��2���l��TE�6�����3d�j�L=�%�[���(�.�n��Z���� ��%L��b0I�WԣE�qJ�"�`�~lY\�v���iz%V��+ӵ�,�;�J���ߌ	��_��n�Rw9tf����L>u��a��w�5�Lw�T�J�j�,�f]�����Bf�y�W�0B-}:�-�D?�?n��|����H���t�Y邭n2O7���z0�����`���s;3 �pvWK+��/Ʀ��P��K�
2��`�ʏ&K�EW���4�t���Nը�/��7�Na�ŁDw�����M����(�WvO��<�8g��Z��/�"&$��i_;�����T�J���K}���v%�~r��1z�VEN��aU\�� �W�܇:��ޖ\cd�C������Pј�}-h�y���U�د�D�r��nD]3ŨƺC]�<�x	~�f��`z�����M���/m���mM"�D���Tk��m�������K� pL�{���;'+���( ���/U����R��<�Os3�'���vt����,���Q�ʤ�.��&%�d�v%��L�[2��&φ|��2�=���<?_2K�d��R���Hs���Q���%�j�U�&W�b�V1��r�	��B1R c�Aϻ#��0a.[wj��Fg
�I�6��_"��
U��/�&̑"�"S��?�O���7.������+*J�q����6�HLd���i�vt��W�;Ԇb�C5N�9�)��.{l��~h+�c���;9G�����H�Ju�;�ܴG�/��Nl��騭M5���"�]�Ns�3X�o:�X�*0$'���{Pr��$Y_r��+���Ŭ#��p/ ^��+nY�~�.�%?�_*d�K�]}�d-)�{I�Z�"�$���ʪ@�!XQ3�en�È���0����/�)�:�N]gc'�-(B�
�]��I��Nw�P��w)-b�	.�*pOW/p�څ<�l�U��8e��3f�HN�x���e�%�Q��� %EP�����A��LF7t'�o@E?�X�3&	��*@���1?-�o��k\-)��s-�r�{�P��� �0�/�
��7��H�s����7�'�X�f�b�V�� ���	a�`���[�f8��|�cIg��?�}�-œ�b���'O$�[�7�PW#5g��a��,�����z��Q�;�?�:��rз*�9�u���t�b)�r���&ύ��)!I=��0���W�V=��}��b�/}x1*�$�M��#6���y���?h[���؋�_���vu��]�?NY^̗^瑘�ѿ0�GP�Hm�\z/$�&��>M��N@ݠ���f��٨&N#��H��*2u�����:\��ǤZT��ɛH$[�}8�O�5����
���Ycо#P )[�V*��6��&��^P���f�ֺ�YD�YKQ��+tn9S��f���L�,V�L���B�3qI��F�ٿP�'��S���u�m���Pi��Kf�x��0�x	2��H���:����7P0�Nz.�����gF�����(rZ��|���#kIG�b���q�ןKI�oOo��!������y���g�C��_���+�e@�)ӽ˃ a��%)M&�q�-L��N�5�9K�Å��BULqp���2{��F�������*6��e8�� g��NE�ѥ�F!'Ė����R��H[&�v�"��0�K3`��?�K�ʗa��9:y�/f�г�#Be-Pt!k�
Y�[�Z�+�]YA=R�,y��2v�{��tF��Yu�(}� �1�����a�6d��z_�����!R	P�`q�l�m{�F��:�/���_�Bx]"g���3k����g�u�b��+_���Ԁ���,�x��̲w�m1W7D�Y4Bx�Cv[�� t�?[���)����*6Z#Cns��+v��0[��]gX�O	�_�/�PO���>8߯#��|��	���ؽ���>��c	�p��q��=.����1#��?"ލ��`}�
43*eRL�&���B� 1+�xA��ɶ�p��.�� ����)�=K�2P�ܶb�aO�Is��i���P�X��A�g�O1z�Z����ߞx#YnI��׫���+�� 08#N`����"�;W���v�-c��VI9�+Ch�;�O��!W z��m�3�X��	帿����]�G�&^��$�s;����{>�����;�0Q>��3Mj�m�ĸ��5�<���ߤnk��3��h��S�{���f�*7'�b	^��AN'�W@]����/F���?Cf��4r.ORU��	���8�0�9����B�Y�Dqoc��i�)hÝ1e�X!��0q$������`ˣ���}�CMNd̙Ղ�n�z9�0#��ɴ�qPN�^�m�	�#��E�7pu�^���,���K�ZG�N���x��B,��e�А�E_-}����5���T�*8����tk����P�i0�_�ð�p�t��I_q���h�H>cC�)[���}b	�V�7P�"&���cB�$�xs�5��x3q�g�' ����F��K2�R�O��=�3b�~;�lǿJژDI\vHΤ`�ޟ�BF���Y"�?�¿�k�� ��H˒��TNno^^{�(JD�N,���uȝ9�	��F+K�{��$�i�"uܹP�&����c��Qf��4���G��$�bN{��d��z�:Z��0��jm�0�A�l\��d��;6ڒk>+�/��-�]|	/�šn��t;���TB�)B���mb��x:�l�E����Z.�������������z��:�n����ѺU�/�Lfyq�������)p�-�"�=�YB�E�+Y�����a>�-���6K���:y(��BvI��sh�d�v��@�z�����y�}RI[��I�wJC|�q��%j�y��YHD�\��s��NJ��Ο��z?rs�=W�
��@oH(�*P-��#����� >��L�S��1��`[�������!$�=z��p�7�s����|��W�O��`�>�[�2C����{�!Vg����SM�3��������ͱR�@˯��A�G�Z��q�����qh����^�i@:�p��p4����1����8^~��{���|g�1��!C���LL�_�Vۧ���෵�:����I��jFy�:lu�)y�3��\b��)\D��������
4�֗k�����MS��mȠ�K���dj�A��H�6�e� )$���˄���ڻ`���
�-���n���*�H&S�?�BX���`�*rn�Bi���?�<���w��%o:Y�9���p�llr2�L�e���Iw���B���D���$�7M%�N�R���v��,�F'�Jm�����f���Ӹ�T�~}�4��+����Ĵ8S =q����1�]�,��}xd}����l�e��MQE�W������ӫ2���Xl�`2���k�)a�G��"ͤ�K��R�^� ����bK3�o��S��F'�م4*���]���䇣?�I����M���f��0�����[���g�P��-��bP^�u�E�(dc;=�!�8<Ҍ�p��qx�}�kQo��t��R�8�K3�5|j*�<�
Y�����L��|I���%�=��YC���m��\d��/�G�I�����|`�ņ�UM��Ǥ��%&W>Z��2o��9��_���<)�V���`�	�� UEy�8�(/3j0^�W�h�މ�.��8&���97X�t��Tu}���	�O�
-{Ć�ۤ�&��FΧZEav�g>�-�()}���.��EP��|�t��Lpk?үϻ5u����(:h��Q���a)�.���~���H^3��e �I�7+������K-D�2[��ƹ��������jv3	oSJ
�w��"'C7+�N��~��0eW1�EFh�:f90��y���De�\N���<�$qoF������{��^�)��[Z�L�y*����5��CϼK��Pw�����` ���Λ�W���J�����>���7�� H)��� ��w�s��"Ѣ�S9Ρ~dwn�����6[��o�I!��9'қ=����w�Z���g%��9�����E%��(�5c^jq��<4�叞�p� ����!ކ��rv����L�T���\0��F=�"*J���ň7�]Wq���B����m�4���|�1��ݺ$Vެ�]�#�' k"g?��ڋ
j ������Ϸ�.D��&mz�3q��'g �/�&a�w]I���Z��~��<�[ u_,B��Y\��G8��4y�-�b��>,�N�o^���fW5r\����Vcc!�zJyE�g%�#  )��˚[y������rҒ��i�E���)2w�ll}=J��	���7v��	@���\�s��C������>�i�%�њ����m��+h�X�4d�*5�v��ڐ�����7U�W�=���R�mf�J��vA��K�[�b=!�(�BL�a���Jm�)��.�.uw�GP	�O`}�"0�����;a�)ދ���QҎN��a�#�u�QX)ͯ�:����V�aGT��z��9���l�0[���K�Zz��U�fudz��<ݴ*nf</n=~�6��j��2<!"r
d��O�
�Sc������͸��������A kJ�`�r�3�##���Kdto>�l���DQp�IZ�0n%�.`�]�9܅ꃊ��DJB�(�ϙ-��QY���iѦ��C��V�o���;���r�H�J5���U�]��:���ɟh�̇��]�if�����u��=�߹�t��~�=Gw�4�}攃,ن�T�`f�>NDi�� J���E�Yp�
͕��k4�0���I�r2"J"'ɸ���.:�k+]��J�����c�QM���J%�o`}Wq}w�Y��lopݢ�XN`���Y?R6<�f�>��F���1F$�*VC��q((i7���-�s��睰������We�dy�s?���W���-Λ$��Dl��b��Ҋ�3�6~J��3�\c��՗^h�.Y�����H''�B\����F��5�C��!������y��M�/�q���-��,z�����/]���o zY�D��]���S	��l�a�Jq<|u����a�s_�=��"=���?�];XĻ��.6n��<Ɂ}�ԓ��Bߴ-�@8�L�!i2+���L��u%����l�h*]	��m������/m����K�L'��e�Cܗު]NM�h����|[�B5ڱK$%�LN�� *h�[�#Y��C��p�������7�`�Z_�,n�x�Y�.�z�2	�97X�q�`��\U`����>AǙ: v׼�a�4I� ��^LF1�g��1�ۑ�ψ
��ӱ�wD3=�����R�!'e������Q�K��)��7^���.�"	�������k����	�3w�����A3p`���~��-Ż	��+k螪��߳�i�{ ���^�n73�<���r9}�N}$l��o�D�K_�|�2��k��'
�?��`�4̰<V�&��K󠓸��9��Q�Y�[����w�$ρf�s�ę�1#��kCN��7'��:w�>p���}�����^1�t%�]��?�r���U��dz��N�'�K�7���ms;�9C}6�`������%D�1FK.�_,���c���S�>HD�ؚ�����/n��J�w����[2�,L�nj��P�X�m�?#*�}R,�rl�;�Z̀	?�r�^�`7bHb.�|����F���0j��/sdd�� �����9�%U��s\$.��c`�C�H�R� ���5mCɱ.�ג<�x}Q��Ƙ{�������ߜuޠ`�k0����}Ѯ��e�{:,;�w9�q�"%)���<}�G�n@K�A�$4�1 �/+i�ey_z�����|j��?M�E�Ue��b� �ԯq���4b�]���j�p}e[�Qʴ��lX���E�u��[ٰ�V2���*����t*����[��Р���C�#>��v�����2@�k�x���oڃ9[�Ä:$[n�L*���׈�,���mt�'^Cl�y}�6�X��g��<��+S$��Q��9�A����FB D6�KK��n�Y�)���N�Ս}n�,^�7�|ְ����;�؎����fs��%eD��s�Uk����y@"~�7�O���ܙ-nH/�c'���}��V��ޒ`7�:[:֗�:�ދ��q��>����&�G����?�~�(���r�k��B�p��B���{i}Q��I���M��(��UOݺD'�����̍��c����5w��<�a��i��컸<x�ziJ8��fUV/�=��`�|
|_)m���W��\�}��L�^����jK!B:e��k��:;4���;�}\U2'ߩ�2��l}'����6�{!2}�n{t�Ʒ�U�yN �Y{RE�d/k�J_!|�����1��m�V2��
��6PS"��P��ru@��?���-�$��Ӊ��pc~�Q�S;��@��X�Lb �P��.�k%o7+q<�>�wz���Ҵ�up���o�q=�Y�b��2��:f�_��:��pa�<fm��B�Q� ���ЋYA\�[����?ύjX\������΄,���N�O��O6ϡ�{zG~$�WNH�e����
&�E�X�Z/��}s�\(���F�HU�QXw�5�]J��"cJ�q��Ǫ�V0�ͺ�FxX13ҩJ�j���y_<,8�l~���9(�K�;���3�ي�L*�j���זk���h,�α�q&?4�n�dV�� ��� h��5ܥ�S��c��R2�?�\�BD3p�P
X"��U$��z>�޾��a�]6�>cz0j|x������(��Yϡ��$��^�%S���§�8�ubl�W��<ƻ.Ȁ3�@��3ؤ��gq��`����D7�T(&��ީ]�y��S���5�����hT�Tk�ɗOQjSqE���?�;�����	^,F�c�d��{������J�u�+5�[�v��g�l�#�Y8�O��_�Q�.�RP���7 R��?�!7jA�D�9ր�4�p�ԍ�]u�J����,!��)Ռn���ۏV��WC��ā��5 q��ϐ�ڔ-���W�vX�p�+������+��z6A_ee���GP�V(ܞàe�(rAkp�������Mh���~~�:�=�ћ�s��0�ESUJq'�J�8��]���P�-��M��U�\��i�+؉t�_#`�]~S�>�x��Ih�y0ހ�8 nd��b�nAQ����M���1����gdㆋ1.=_���D(����u&�jCւ��C��i�v/Ѣ��OOn�ͤĦ�Tj;�1F5ň�C�D���M���d.7�^ȌV�*�&��j�X9q��g� r2�İqB}�=�d!��^��g�D�~a��L��B`x׬�=gB,��`���U�]�v;�c�� �B���`� @��KM����!o
����<�vr(����M��X*�D!�n��c��{��*�f���%�ڹ�5�D^d��(HX1�(P"�]�'�sSO��Φ�f��b����%$+/œ�փ�XY���Aoﲵ$��^מ��#�E�`O��b_c	��t��4�_��;�����!A��1tAEh�c�-�@ѓ}hs�kY8pFl%�� H�x׭| %�h����\�iN�|�>ѕ2&�f[o{�f=R��̠�r�W�����}�gbN�΁`sL���]�?�_��r��O���>��	�m�0�/�xӛ -w���U�6c�L���_�h�bFH���`�����n-��-�ڟ?  D}��SI�j	�,�'öj&����ϖ�l�GP��������q�9|U#$4�R�'Dd�	���U6�2��O��-�?��o����Z�	$�?���	�݄���x5XJ}K��B�ms2�0ݗ��=X}��)�tV�HN�;i�+O�|1q�D���AX �"��1-NVUݮ6?�vY�͡��D
��o��
��jͿ�#��֤6S僭�G�B��طRP&Kc9��xً��_�b`H��l���C�R�F�[ʑT�e�{��g�P�_a�叨@cu�%lR4,ԋ�
aُ��W/�CU�����W��U��1e�Ke
�����H�Jz�ɵ���.�S��� �d���..u����Y4m��,CV�-lÌ~ӱDKr)�	�M�8u�Ա�~<��~�x#��~�0>�1�#d���sY�&X���ni���11���"P<��uJ��~�kSI#I9y��_iIK���'&5�?�x&&JO�=�
a�6ԣ�b�yV�dN�KT�V���fBę���@	(���CW��S�D`�AXz��~�.���ӫ��S��ԏ������rW�4�1�3�]�b�=��L6�:��8���~q�|����ʳaE��P3����C ���-�F��)�{�r���x���8	0���P�^���(�c��d+;�EԀD���6�r����XSbu=sv�٘ԏs8���P[[i��mmV��c9�U�aoI<#�i:�'����x0���L�>���1��h��4s�����"�����X����Q旬&�=�W݇��لuu@Wi{;��V�����H�)�H�7�^F�F�S
+n��k둝i�D�AO^aL����f"��OqA�{�{��*� o�n����4�K�	�G���^Uv L���e��:bΌ="d2���vmΧoJ���/��O}׻!9h��9��ͧ�9�G��\|��7��2}���p���$9����p��R�[R���(:�~OT ���7.�В�����"K�R��9�}�)�G���67WI	��3�@e�S�����3���1)dS�ˊ\o��fh�%�v�)�Ǔ{��Jn����Zn�c��Z���Z�48[/�S��ˀ��j�����Ƹڨ/�B2i�{�1� !�귴ZG��|ca�zNL�[:xj�KpXI�'!�u&�<
�S��m��F�pÈ,�K2��ΟZ��cR ?��bA�Wת����Q��4���/T�.���I��L^�Tc.:����C�Ζ4���#��w���]��6oZ� �*�-9O��.�7@4lUY�A���V9Φ8��K�or�v�X��Y�8B��՗���Vi#������w4�*=�D�^w���y���Nd�C�
c�B�f����p95��rMA�S�(bBg���*^�L�'8j�wؖ���@/v�0���jW^)%�p}����	���+���;z�(`��z��߻��U���1�R���q�=)͢��d���kΕ?Ö�(�/�f�/� �/���c��{��"�F�nGP�j��"����;�`=�Y�GxZ�}�]��蠽|;�Oa�)�M��l�� �(@�)g&�]���y*��VI9}�q%\�*\��d��.�H#�u�a���`���_�;���e�:&��ԄVk�}�5t)��ܾCq��������Ȧ#�I��.���!�X�4jJ�ĝ�g�"�&�~�/[�wa�Q��Y��3<�=��`�6�M��� ���2��-�3i}�Q1�L������o|H$��MA����3{�&h�Y���ChzN��H�S��2�o����ȥ���ά�Y߬PN�l�k� �몹Ȱ$��W�D�I�1�#�n����qi�'�k˝l��Í���� \W(ܙ&� �W'�t_4x�qg��yn��|d��2e�l�'�'k��S�#�n�����(��xȫ��l��/��,X�vux�s�Fz����~����S3�����k���p�p1�;��2�]z�[ ����_������kaIe
��R�wG3���-p�'����e�]��[���suce�{͇[�9x�E3�^�U!F� �\��������:$A8�J�#��ݭ���:�HQ�&˝Α}@�����������6g<��I;70G����!-���R��Fֻ��s{���6��{᫦��b�C��ar-A�㡈o�
��Uv����<�-nfͲ��h;4E���q�$�?��p�-S&�����6E,N!@C��v7��qԣ29=Fu�]�mK���mm�癊�I���}N�#vc��[^��.7)1$:����9�39���o�r�����'�z}+��cG��:��;�F���	*+l]���A|Ӭ�c[OJ��A����B�~��Y����sr~x�z�s��?�
I*�LM�XA�*�^��9
�d~�^���m�p�R�Y��]�d�߸��Ջ�I�c�6�?ۮG1,���)h+.�٠s7�F6gMk��8�ixG!1�=$�o_�lW���c�lVG$��૛��!bƂ+h�
�4c	�aԤh7!��W��8]1��,�9REȴ�\��������� �9���#�J��Ӂ����!k\(��#�������+[�F��!�̬[��P%��=� U�����zzjQ&�Yt;8*������I缪�")>M�ES��i-Ď��84+ڮ��0^[��3�Tx��د͕�zB#��#8r5"��Ї������c5�.p2#ϻf�� r����:�`A��Ȓ&���}|KrД��M:*2�!U�1n�Bw��)��q�b�ǹ=�0�v��;S�������9���i#�G?���4r�}�hs�����;���vD��wpo0R�7f͘�ݒ�z���trc>�i��]�L�nԠ,�,��T9��$�!I�T&8��-c�)���s�ܶ ��U��~V�i-M6�X��[�h-]m�c���Ǖ����?G��'9��9(�R2\��T΄�4#����F@^�r�����`o�nZ�]Yʍ����H�d���&[E,���� ��ՉT(pE������%H��Ρ�wo���b��X^�\��j*��յ� $���o��U�������Dr��
�Q�-��8#?���1��:b�,� �,xlM�8���9VD��mR8������0g*����Y��fv?�(C��)��|o�� ��$"F"�4jD|�-�Y\��P'��G��	E
`���0��nR��'�<����L�ȂS��e�2g[��IHB���6CN����+\݂�;�J9�N�r<��ufV�"O8��ٹF�	�w�r�{����C�W�}��B)�i�i�NE�P������z#�sPξ|ي�EC$T3ouR�����J�DU���c[Sr�"snJ������?ȟ���m�"y��%���g�����og�Sr�_�n�'��/T᯶�W}�#i��W���������,�x y\o2D5�9��4�S��G�o�p�~$Ȥ�|�aDq�	��-8�<�d4�M6��D��
R�!�:�����^���X+�N��Z�ܝ΢�]?�eW����51=����܈F��<�� �tn:wQh�]"n��j\�7v	��]�Q%5艺�[̙�J���y
ć=��i	�:�4V���h"��_��٧:�a��Jbʬhs�uO��%���,���p�<���}R0m�a�����"bb8�ώ�nct�N%��qf�G���߄����&a���s�4�Z�W�j�N��%��� �]V�(���})��Y+���"~�5���@���`śѵ�Ɇzt�@1Q����AzJ�]3�G�H~��U���*0�-��T8�迹M)�N'\��\�-��G�y�o��Bi5��e�>���[��|�,�h�r�9y�2
bH�F�ȴ�1 ��d��^�r��v�l�4����=:V��EzE��fj=� �i�.��cmb���1�׬Ƣ=0��&Fǚଈ��a��{}_�?��^��u	J�Z�G�`qo�ȳ�A�?� 
!���۬K��c�6��r
�\$-)BhJ��`�A��A$1Ș)n���s�%��<�,(��k֢���b���x�<	�"�	�W�����'ʾ\���]g{ʖ�<!���"��h
�Ge|�+FP�K�aL`��n���ŏ�yC9�"lA�S�	�q��>��}H�'.FRk��ٿB&���#W���;@�<�W�8v���1Ec�Qo��(�Q��{���u��
cIB� o���7#BO���[e��z�Tv�s:��g�7(-Mf�}b�b��7 �	D1Ĉ�F�N��l'�{V����S�s����x��$g�[VT]���u��E� ���6�"�9�bOt�[E�����@ةQʮڼ��*{A��_]D��PU8��#����<�;��i��i=��q�I;�L�˼�-�HӦ}�0"�y3������0>A�Ge�s����\�֑c�D���rf)5Z=k���:�DzNE����K�Ӄn��tO��}���q���q�Fƌy�����fP5����U�@�Ӡf�g#��=���Z^�����N�.7?�Д�Lt����,��0<%�)V��dրùw�_��$Z'Z�D��䎄��B�i��Ow�~��dʇ��}����u-Es�5�X��%c�T��Z �	@�ggEZ�h�H$�1�[���ي����h�!pj�H��nԕ����<�p[!U�A�?��������rl��u?�N��	5~w�D<PR��@��i�RU���6L�8���u�찲F'�e�6�Վr�����-�*����ڤs��a! �f8o�%Tx��<�>�y�bmYX8$�`1���4qp�-	��5�q��l��)O�cʏ���(buV��H�I2�#;�s��r����>W�Hh"����[�
��["��x,�q�C]��]a5������n&�O�~@��o��� )�h2�����H޲�5R��1Gq�K��̕U�""q�d �r��y���]ͮ���G��N���!���t��Ec0 	T"��� ��\��Y����-�0ʗ|04�
���\�%Sgm���Fs����� <���}�]@��12v� ��Pۿz������W]8��%ڢȯ �%o�9)׬�Т�ٛ�U�"�'�Z#�]�ʑ�sSm��������������g�2;o���k�����N�.q)Fy;��>�Tg^Η�Y4E�csxZo7��*�؇����$dS��+G���@�d��r͎�H�h��M����7�A�TV�}\tk���B������(r`m`Qd-����p@�Ժ���R2fM��ڳ��B��W̓��F����ߋo^'zC	f��{$�5����ϥ�ƞ�յ��A�?��l�A1l-�� ��?�p���UTqi�3��h�1� �����1}T�Dx�����󞏼.�>�mx�V�9<��Y��x�6`�@�X���b5mu����%�V~Hܞ�*f��n�r7H{��q�O4O��"Jaۥ���3*�8�f�/���f�R�f2��T�R��Cx��H�7Ԡ�
Px�LΌB9�Pu=o��x��+t1�"ϔ���
n\kWB7��9?Ϣ4����k>������]\�h�c8������qyŚ��8=���*p��RN��=�Y���TbD�A�t�ʙG������/��9���KU�wlu��g#���V��aS�U,G,���	zY̂vy!𧭌*;�uW�?�j������������⟾��`�F��yc�Ć!�:��I� ��8�5R�����O��L��sȼ�WM�hSU<�b���nʂ)R�ŏ���@�/��<�{F�e���h>���u)�e�Z����-��鄱��/�{�=�5�N{�]�����6P���.>w��%�	��Ъ	=;�c��_���pTE�_Q;�W*�;O��%�zֈ';�*]Zjb��h\�,�����Q>�^�����|4K0�\�-���%Y���\8k�	�x��"�����_ή*%*��R���N�_:�-���Z�2�"���� F,���b���`ԯaN|u�kt@�d2��_/+��>�>��X�M�t~N��{#胖�3�ç=<9-=N)qoOv�T�����3)�Oq�.�SX���I��Mk���s`�Wi3�!`+�4�9��Ib�j�s��0����S�Ys�u�o�K�h�j_2�D>3��}OO�h�����ҪX[�g&��$h ����&�M�Ǭ����om��N��.Ab�A��K<S�����Pf��c���uf�K�Ɔ��w3��}�I�DuTd�vT�G,ٶ�mmﴠ/�Ϫ�#]Mg�f�A q�4�'��m����z�y�����o�=e }���zc��w7	=u6��P_�9������7��ԇ�d����c����]�"���_!΁�>e>�3���E�-��>��̀E�a�IQa0^pK:.��c	':�(�yTf�.�l~�;���ԧ�.V�L�_�l �-�[?i;ˋ�ѳ� a����Ϛ�qZT�m���i����`j$Q�j�=����K�=F"4v�V2`�A����!�a��Hfv&��2L2�.�����Inp��G�T��^��;�T�m,��9�c�?>r�b���Xg�I���� ��z��-���@������?V?��� �{��O�?p��a%��yzu�
��U|.+�a˞9��W�X��8(7+JRj���炋�J��	y� V�y����ͪN�V'����oQZ[I�RX�D��DnZ%�K�v�g��`J��Ϲ>�ul�ȼ�s�Z������}��� �dr���CN�Ӊ]w�	!@!����z��W�O�]J}
���2N��
q�C��r1��$o2�>�����3A�#�G�������=$v�x~���p�Δ��?4g��~������J�U䈶�����n����Wʹ�;1q�W�+����y������.6�\�1�!����is�}"ݒiڅ/?�X�	��a��j�����Q�/@s��Ӡ���\̎F����v�n�.�
�I���ֶ�}q��F	�?�(D�2�M^=q��܆&��>��