��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���tǐ-a�Z��e�l+�H�uW�Љ��Lk�p�@}5�[o�Hݤ|����j�{38��/qlW04\h"��=7P��2.��[��,~�����d���4�o��3%��!�:���&��G�Q5FJ���H�(�m���G	.��I�I�_���]�r(1��k��0��h�&��b��j�����Ǘ�g6Ԥ�f��*��9dS�>}᝟�i�C�C�����Ó�����RǬ�]�BU�����po7(gP�ݴrsе�7�V���~'�u�=��Y��<�(�;?}��Q2_�����-N6�R;SK8�n#1�d��0R*h%]6@�Kp� #�|�S�nj�C���� ,`�T��m7��O볻�ʗ���lUw�{�\�����pL����@��pEkR։��h�����,�Bf}'}'zM��������F�/�ஹ��<1����}��I�j����Q[�uF�"��0.R��ft��f%&k���.C����}���^���*-�a��m�4�I#��zʘ���6��O�S]mQ�o����CH3����V��
A, s��<��h*Dқ�0É_n�(�w���[��=�\D=�SЧ��M����d���x�K'O4S������\�fZТ�Q m'3�#��m�5uTa�-ia6G��>���ŷh���$'���[l.���cƓ�K�O�� �	���Ԟǿ�������qP"5�pY�r�z�$���Ȉ�jղW���k�k�v�������2�?g)�{�**F�~�z�k7� +������(�{�$mDsq'����¸�2�]�\��
���2�`�Ŝ���;�	�%'k�}��g�x9�G����]� MH-�!���\�T��d���Z�3Y�VB�i�rN�'u٭.�Ğ��q�	݋���	zT�"�6P{樎$��V[��ᐐX�¯a��'Z���W?jjI"1F�����v��T.���<���<S��D�Cp���W�v��$��v}t�g�Q���C�'�I�6eq���_xp�z��F�P(��仅rx����A;o�眘�(�*gy\��!��K�8DΜ��^A�Ы8�m<5�G�'�9ڶ����w�������Y��uD�R��B��xB�1l�
���Ô�VeΈA�zǫ��"Q�|W�LquƜ��<�ٯJ��ō߳	���{���0�)��QI_��Q)��X��ҏ%"sV��MC+,��2I����y�Ca!|QU�v�)��ˆ.QC	��U½z�2�3I��7g�k� 4��Yr��{y����~����
ŰS���
�L�x'ӄ�Өm�$βC�����9S`_X��a�m�G}�MD�ө���x��ƯJ}7Z�A�	��Ą�D('Q��p�󌣠��r�U�U�����Ӧ|��\]1L�_�7�2�D�o⋴�ô�T�����e�� D�գ:wL��}�+�Xzŧ��6�ya���ƌFW7��zKd�y���������R<�6�[�B�2��%�H}�=��o���7Ht
��d��I����$�	��w�-��1&7�]ՔŦ��><gN����u̶j:h�0H���Ho�Ô?j�'��z*F�f��ʍ3f��w G�ٝ��;WLE�,�|%n��J�L9Vpi��z�j!��;�4�n��y8���E:��LTAӽ��S+t7*&�PIlS��`^��X��fY����oo�M!��h�3�mwU�Qg��E����̏�,�U2��gΟ�B?�҆�3��nx�~tF�e�����UtBr'�YƊ��FJ��+���.٪���d�v���F9d#*�~Գ�[��sS��(*��8h�|�{���߸�<J�С&T��D�@9urMg8˶�+@t���5ƃ'rB���ʇm�9=���N�����8Gq�����c&1r��+��s8���w&��3�
ӫ����Im�,���'�����tL�
v���B�p �Q�"��D��l�N\��q�������uR�`�-W��Px&E�r��V��K������dB���1ft����赥�:���#�[a~t6��f�ڵ1u6����C߅�׸�>)�J��1D&_-���l��@^yk��ײ����N���^_�e���{��]S��my��)Ә��_�'�6D�F�1���ב(*��Mz
��N�_��):ۢ���� ��DQ��H{eY�,s�z�3��ț��T$f��zN�ڑ�����e唵D����v�>xQ�@�.5^��ۋ/�7�Ý��&&�� C&*Ӣ�QtZqo�RR�!�P��H6��h �pprԬ��!�}+j�)��?�RV�a$ۮ1�*l�rf_��	`����2��Z1�Ěێ�Y!7����HQU��t{*ph~Y�f���� e���M�YO Ӗ���^�	�\��\���p�ξ��"�5[)�z�����g�@����K3�:�9�[���
M�͎��9w��r~ө�]��s��y���Qa�,�5vE��o�Y	��f(U�>�U�{hK����+���pԊS\O�o�KJZJw��T0l@�G�� �]��4�Su�G%�.󨵜S_����,���.�v�����/ ��*KH�_Dp��\��A-�[Km/+$�~�`2��x=E-���[�Lh�����jڅ���^y
�%��`���UL�� �%`#
����8\F��%���Q]:���������fL7�싞�˺��<�"{��
�D��o���ao!3\Y�MO;��f�BM������Jݦ�$��d�y��J�ˡ���M�:�� /ć����$�;7���_�b1��U�#��ZTpw�����ף�'��>��=SMn����͒\wtf\PWyu�]lk	(�{K��Ezw�{Su���ip�cy#��);% ��˼���mx��8D�������͘��sly�-�t�DNf���$�Zh�;v	��c� ���L�ow&Qt^�;�1���Їs�@#�_��蹹>b�.n.,��])\���'�����<wh��
K�#�Hp��<B��j�?�c1q��L��Ԥ�φ��BU1M��f(�w������?G��IK�G[pr�Y@��:�}>���\�$a%��k�D�QH�9�S����.�z�E�F�8�j ��M1��C�G��v�%#�R7|9�����%f��"ʈ�CD�?G��)��z�V$�(Q�#�F�g����D�E_
����v����5���{��bg��8�4AEOS���u�lv(Cڄ�s��5P�n͙�I����s�-J.?ax��rv"83Х��w�\������9�X����Gh���l�Ve�쎈s�D��(�8��~��#0�\��r�f$��)��?EUǃ���v���7[?�op/m��	��=W��W7@�|��U�@���^�XaRE3����VJ�����Ӽ�*�υ#О�4#��_@�a����TLd���wO�١mH)��^����s����?����|�W�2��b��5-�]x������>P�: ��i5"�e�@�Sz��T����(�Zh��ho M�_��<6��� ��k��/2��`��3M���?�vU�("q���L��6S»�6�FUi�N?�?��OֵKj�x�	�u�����o9V�[R����K�� Bpq�7����&8�vQ��_��,'���ڬ*^�}�\2���.&:
���ԧ���AĞ��������5��_�"�b�d<�=�U��͝�@[��D{���q��K�����������VX�m�����q8'����hh��UCI߂����(��?����+�t@��*��qQ5�`+,�V���|��3"��rݪ����Ĺ��f���Ծf�"|�߃4[|˷��X��NX�]�\ޥ�������ZJ=�k�T�k�A��-������&���qI��s���܃�օ�@_O�{��a�i���6; ��yɰ�w=�]����'��1$�c��V���e�gG���|9��v��[=�y(ZOQ��+�pN]���i �+�W�
�#���Z���Z�if�W*U�ܱ�d�`��6�����X��Z���ٱaE-��#���sN.A[�ެ+n���=]R9N7M���0� F`����!�����y��'��ޜ��L��a���SԬ�����3�7U9MtI� P%�+��X�)�'���g(����>?�f	�M5�۴3^͌K'��PQ��s'�=lr�w��葈��Y�}1���Da�^�ګ�v����|����[��G>d.)�$�un�-�u׎�6��Y��$	҈;���a�Z��8��u��-)����ۅyϬs��0jf�|K#>��|vI?GF�v��cC�U��o��-��9��@��r�����}�����O�W�Y1���M��_{���������p��z4�����t�"/�1J���
1j��Q��=J����.t�_Q�������qǹCd�D�o1���i娺vٞ�' PD�Ij��oT����F�ײ��<o�T��{~��R1�W9b{t�;*๺��Cqb칁�+��0A]\l�O)��
�p1���#�;-Q���K�u�AY���1$��{�*�o��,>tK�#�v?K3='���~��yst�K]�xiy��t6?2q�!Ԙ���4S�|8�8?8�`����Q���w���Y��d�
�℗����o����-���
B`W��7�ь�OX��b^s�7��a�^sO-%�Z�ޕ�R�G�t H�EkSl��2�NHY Ԝ�̯w���5`��
�B��3�&�δl���k0Ք�<��C��u9U�,�K9���B�]�N�B_TW$���r�����2$SW x+a���W ��fn�ܩ)��[g�	J��؉[�j�s�eiV�*L P6|��K�ahOl`���8���������aJ#2m��6�1S�}~i%|�"'�y/���m��R�%�p��l3>4h�+��a��;U`��B�4b���\KZ�ީ�Z�)u�����#� e�3�
\w㬪��*�/�V�֦}���o?���6L�]	���?�P=��vۑ�l?�(�$J���Td*a�8�YBD���KdQ9�����]��8T�L�'�Ή:�m�,ޭ�Vf�K�wO/R
T	�+�Y��T������JYj�|�~�[{�+@�KY�p�Oo��K�l����1����G����k���8�:��LQ��Rdݱx�𛾅�{�O'�0��a���K�],s.�����1����G��q�p�*����_���$���I��i%@���E��ɿ��O��0/��#�Y���c` P��K�t0�S���aT"�����h[ա�͔�>�KnѦT��'I�����t��Z�F�k^Z����_���k�^���� ���
������[e�^1�-SC
�|����O�z,\����^�f#��K�	�92EQ��x�g	���3󥷐}[�%��X�L�����$��z��e���U2�?�҉n���A���(��@>m�R����_����?t�*ݶ�B<q��I�}ʆ�m9	Vf�y�h�H�$��NV��Aj�'�O	,�k]' 8	��a���泞�tG�J�@�;�����F��8<��X��D4�qЀ��|����ʼ�������冹a�=�R�2���TB$�r�K*�3]X��Z��.+��1 ��3���muÒ��%�ɀ��F���!k�.�s���f\%��}Ì��n��i��A�����OO���2�[�	�=4��'D��׺a��N���:q��Ą&!��R�U�\9Oإ���������r�S~v���!����m�f���;���-��;�X���9���"���\7���!2��*Z=ۮ�o]WB���0���:(������/ށ���3�!�e�wqk�U�Q���S��s2�2�	��3��G{��I�T�7�Y��ڡ�����r0z��mR��.�sd���� ���Z���f�{�N��3��~��ǮC%��C6G���YS��*��h/$ʓ������u��q�������yJ�94���l1��Â���:/��ΪG/ �U�1冀��&�4���^C3�1�']ʚ�P��V$`�Mg%�����孧sVo�6c��-RmL�x;m9j !��L�+����ORӎ��(p)ե���kf�Ϳ�ֶ>@���C�|Ӓ�qWؿb~�[}'�7�KX�4O�H���g�b�PAc����>l?�.�����X�� ��*֧:��a��O��TZ��y��Y�_���W�����{�]{R�s��S�ejh��J^�{��U�Mmne��y5�O[�׉{;KRQn)!y�o>��6�^$���¿��m���#p�>�Ü��O�C�d�v������y�z��.Zn{T�d^�T���2��d�{����H��Oȥ�?sA��$6;Y��vV�y��=�"t�h>�T��8c����pC{@L=�|�]M68B
w�����{I�Fy���j�~�޻������#nca�g� ����{���P&�+