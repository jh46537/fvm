��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb��N�9��8�
`J�t�+K}=Y��-��.�1bSA/�\�1��Qr5>ڇ�	�3l䑔�5A�󜾘:qG��)ۧ�O����s7庘�<u�
���/��O���j�Qi޿S��JQ������3U`tS|�G�����udB��<hB�#��.�$섵DX� ]��I�ɽ�621Ś�c��|��e�������������L�XV�  �$�P X�=0�!}�S7��e�S���8��p?�U-ZBa4 ��Z��Ҭ��$Ǳ���U^��(����#G��=��hi�;��\�Z��=����7����x�Q�o��v(�S��Xb�c�$�3���`:�V����8���1��*�.]s� �`'��L�=PJ��;D��$5���K��&2��}s�rf N�m貋_ �� �(E��s���{�}���x�U�5/_�"WZ���fR�w�.X�˩���!�*�6d��p 5��%a�1m%n������ႊ��QO��:n�<�̾=	��y}�#2�ba���w�ku�'�J2h:U�!�д����ޭQGF�+K��	�Dpm���~�;��qb�|�X�oG�w��ӄ�M�(�D�k\��[#�Ŋ����X�O`*��E�hGH�5H�.�u�O�z�VY�F�Pb�hSY�]'H��eIi1-�=��]H)�lc���3N�_�2�Ϫ{Z�2���=u����)��d����_Z�!W~�0|�����YV�C�pO�8#!��z����*�}��5�mol�DN��FnZۓw�����>r��ĉ�U�)���!��1KcvDL'��ҿmٗ����T��@�6�u�{���=�ECR����~�p�0Y3f1��8Z	c]ө4z�u�I��_��^��}�b�i�m�S5d��C�.LUk쯾-+�q�"Ш!1@�o�O�{��l�  ES��t3I��A5?Sk�`�+�{�4�&�N�D��k#�g
�mD��t�u%%p����Z6��Z�39��$\񃰉NV}�ɫ��Q��Y��H׋#tl��r��m�� -��MTze ߷M���3�/��.�J�b6S�z�M�i�"��K䗐�����Q_��=i�!�x��:Vw)����6<���N�G%yTؔO����!����|ytP���� T�J��A
(�W��& �?�}WuA\��$�z,F?�
���ba�Z�����.}�j�6�����F��'�,xXb��pRi:{�,Լ�ʉ7����*�k͕ �BE D�&^ҵ9�����J���U��'���)MB8g�T�������`�7�!���:�?��*发�.{�y���M���I5O�b��^EØ�3f�Ͱ-I��up|��#�
�X�6�w�MXɞ����"`V9�I�P���Em�%㸝譝���1" ��O[��ϒ02��7f�
��b7T7	1��ċI��Hgn4m�p�(�n��ӐB�{U��ysW�C��7����0�Y�a>��E\d�Jg<`��+d)O�Q��xTt�R��_��yh��6�L�~G���1I�j���4I��l�,ݻ�V��I��	�G�%�Zb@W4���jӥ�N�y������F��g�5綂��d��}r
o�m����Y&�q���y�jW1]$ge���B$p�|���H`11�YTZ/ �<�Q�X���y�<��.�CB����x���27���g����o^���O�+vm%��mJJ��?�YpV|6���.��+'��Z�ӂ����{�*�B
|�
�m�Cc^�@s'3W� ���0 -8��3�ߐ�a�yumW� ��7���.�7#�$&_��*�6{�1HFd_��u"�ޅ<-V���� �� ��*�$JԇE���j��'�A�_$wR�8�1} ���'�t51�\�r	�`QWNyK�mB�w	�:���J��+�'�r �T?oΠ� /LL����u��E���}\�&�TNH]����x'�(r�oH�l������^;��_a�Va,?])��5C�"���P�T��h�+��`l����S� $�&Q}R|&}m`"��  �M��V��`�����=@�A�Z�EM���ْ��$�Mů��:�^+~X��q�K�,��~^0�`�7�+�⡗�M�M�%��f\B;YW�V�~"�����-vj
 �����ڡC�������9���	��&�?�T�9-��Q�tuu\�ݏ���{��O���v�T�S�k/t�7W���R���EX^�%2�{�c�}UK1���/���r=/R�g�U�TC�f[�zJe���5U�(d�s���K3�Xk��P7apN����8��x颼YM�2bMN�E�?y����5
J�Qe�}yx� ����N��7c5�>���Y�����FU�}6R}U�F���sk#н�T��M�|���X�-�Q��M�X6�G<k36��#��m�|�����h�b	�ZS�JU�M����gO;[���q��M��_C��CuyXv�^M���6��K[>���U*cwU�r����o���S�
%Q���^.`9��o���U��XEJۿtV	/������������~QV��V�]+� F�01��01��{�"�����h{EG�&R�r󫡇W�C#0�A_��o*³ʅ.�����<惀(`�^e��x����Q�lLcS97�\�تQ&v>�č�PU�~�{������N�8QA�:��s��u�c��Ђȥ���
"ׯUaQ�ے	����Q���>kP��%5�'jaL�!��G4f�L�V����qN��򡓗7�œ-��XH��L��$�	2i�=e��i���?7G;V)ݴܾm�q��?��'C�̂�E-�b�x�%U^�a�����U���I7Y¯�=�޷T4��R(v~xSO����d�{~R�r���{��T���2ݚ�7��ٮ�\ğ1����$�("��� X�A�?.6�#狕�x�ؑ��O�H%���TR�=��k����g����7�b���.̇�����a1v��b�b��i4v����\,x< ���:��&��)3S�q9��KLA��Q���S���+>>#"�$%$Ņ���E�5V>0��r�IV7F���@	F �U����]�:�[|��x`�J7��u��N��M?)�ᔹ�f$F���JG'�]#���V�u/bb��yW��DĬ9�G*�{�f<��^�V#�8��W;do��o!��~���*���e����ubBIe�֎q2&8�	���*��>�%�9���&��DE��~��ܲ���w*��>n�n�ݷ6�@؁`D2��jҜ�T�W����~� P?p)W��< ���4ΰH���B�|�(�Ռ U	a�>��~��%���D�2s�)�7����/��4��7^Й��hGr��?;/@tѭ�z�~b�A�U�����`'�.�&o4�׫���Z�|���Ϙc����0��IU�����N����L❷|1[�#4���k��R�pE��c���5���r�3�BA!�?8�����a�²^bi�e�k�ف�ޛ/��A�>(���)VO�LzQ���^K�d�f=�$<�3S�W��3��`�4:��*$�oB?�ϝdO�.�Ȝ�m^�_PM4w��2k�H|���-�;T-o�"��`(q$\Gr�ʬL���u��WFo�K�&*NXf���������$��E@����h���d-�,L$���� oX�e5��΄6�,騦�k�v�H�>�g���Z4<@�DN<���Z�Z���O�w���"�qV��q4�X)���F�f�סۥ]�,����i�1GS��x9,Duf&hRx7����w�v�{��zU���^u���O���o:��?�\	�y���>���gn�����D	��W��7�Ikh�������g�h2v���I�z��r�Y᭡��QK��}�/� N=}�)V2�άg//Q�>E��2y�oP�j��H���-IZ�k����:�oA�Ѡ�
XC�*��d�n�Ozd\��e�[�����G��}":Pc�)�8���� ;�����!ep���"��N�zj˥O����S+}�r%�9։
�EU�ʐ ��xJ�r��>��8p֞[�O,"q��݊{��_���
v3Қ��~,y.5��X>�͠���D�{Y1� ���y��N�V��B���.��/o�X�������;�j������2�o�Ks^ES�i��j̵o�p�� ����Hc�/d�ց�<n
�G���7��oO�09XTL�������N+�8ϓ�����wm� :0�4�V�\"ō�v��w�=W���~	�̋���������W�0|���X����[�����\�;��Û�������^]ح���/ɋ���/U\_¾Q�_���56}��"��o�&��'�.C_Z�2�t;����L���p���CE��ȵ��rT����nF�/fL7�ޞ��ٸ��w���������ѹ��;#��L��Z�Ț4�D0����[��Mm:�0dX�% g���[��A�De���è������ 3��J.K���Y�c�^�)��V�}}�}٪q#G %���(Aq�&O�X��Ə������g�C���ギ���7����ڏ/L$p�:\�~�c@�:)G��7�}��qb�Z�1�R[庫� J#x�� j���>jg��1�_{D{����e�C��#M�0]f����2���4�[RP�ͫ��rCJr�'G0��o�SL��p_r�����聧��l���Β���3#��c�3C�%�c�Lz�c���igl� ���n���*��:��,<S�MY�����n��s�IO��Ce�Ɲ]�A,n\���A�ӭ���~�j�s�rؕUT���P������ 	p�J�)v+!rL���h��W�S�:�B'��	<e!�z�_��~��0�Y2m��5(S� �a���[�.5;�eC��h�GoSO�h��:z�Ђ��q� 8}4�M0�y����h�q7Ø��7�(��x��,���.�W6y/a�Qv	R�=)�k۟���1�����db���=���v���<_�cօp����Q�:L=@�;�h��ro���Ň(�;�6�=�N.=H$��B9�D�mJ&� C���ִM�T�(�-y���,bwD[�b����f�$�.��jW�:�Ȟ�����i�*���|B����tGe�S��Y#��ڞ(Z8ۖ�q� ��Ql�R����_���uZ	���������΅׫��d$4A@
�2��47�+)�f�	t�q��5��W>v�?4����4^:�O�Dpm���&xg�K��d��KK�� �{��lx�9 R���8jN�n;�����!`knw��y��_d_�����xƹ[�-��>�vQ/�N�������)�S@�m<{��e��:B O�����bwbmL�C0-�����h�+V�n��Sܶ���v�s:�=�^��^x#�|}���݄�nS�w�fڍ�b���,�� I}�{��H���p����/�G�PF�课�a3�_٤�c�nh�zAܖ��7�-�\
Qg�T����zBd��GE�&�l��vO�#���d`���z�'�@g��Փ��P�@G�=��H�ڼ�u[�tD-��	t�#�b��}�I�ϼr��Xb�)��E��4��p��BII�P���%뛆��R�������ߐH�;[Ð�'+�	%�ѳfK��G�XabH�Kng�q׶�T�!?^	�OMc��uo�}7J��0��ȏ%W�b�UB�XSM�1��v�a��|�]Z�TSi@X�r�����,L{q��O�տ����=�Ւ�g{�:����q_pT�lO͏�u�êA%py�#�q�3f�u�])b�t��B�qD��n���v�^J�1�Y֘`����%ǒy��tT8�ɉ����� ��WiP�Z�B�3��f������$/໦��������!~`o����<��Jԙa,������͝��(fe��D�=�VA�.�v��$y�F��9ٖw�(՘j�'�B4�̳��}�/�,:%$�)ȻB�@�q���/�d����:�Wi��b��%�L~�~��<-��=j��,?u�l_��ٟc��ؙ�δ{����A��C�9�gr�<����4/w#����K�U���, ���2x���Be)~�xwI8��З%N���N�B������
i6y�Z�S'y1<�[J'�d���:��'���w����ţ`8��-����/��%����o*�aj�N;2�)1�(�ߘ��
��|��J�Ǹ�64�~���'g� R~V_ߟ6������>�c�< ���B\��f
��Lt3�g��e�}��Cm�m\2�I�Y_B5�Wq�Νk���H�3,�"��ԟ"�����bXv�S1�z� 8P��1`�c#�	��Y)���Cئ�#��&u�u_Ĉ��m;-�p?�jW��a��������"�g����-8���k!NjD�U۟D�P^& �t.��O�x��~><"�-�cuFՖ��#Gq��x����'��{$QD�U�%��>�Z�\E���A�x�����EBX�G�l@_����簿I�0�0��Nb!�܀�]et��$�0�tw�R�nM:���/9P����R�r�D�� ��;���_�Ʃg*D���n�o���'9�d�^d1���H��*I�O�a��� 2�i/��e؉x}�M�+��n�m� �r����0���ij�Jf�!Gc�h�ɠ�X:\k�4��#̻K�@�*5A\H �0�5�a:�Z[��!�|;������*s��U/(͒B<����ϕo�o�33zw���$X�Q���y��qO���N�H&�xq~�r�#���f�b���� �;1�`>M��(�6ʐ%��p:�� h�%���D��`R��(�E�쫨zK�l�h��W`�$���U���l�1�L&MsC�:�G���*IU��y���͚B�V� ;6
�:���c����3��x���H��LG	��ݮv�>pa�;��iG#��1�����z�d�'� ��H|f7�F�V�e�Qk�5�����%�9j�O�̜����-����#�����������_��k��a;{�;�X�QPK�J�o��靎�=�PRVPUX;>Ek��L�`��hZ�4z2��[�?Z�D' ���ܴj2Ԥ��j��wJ	�e]k���4������8) �b?şoL2eX�|\�B�+�a��Y��-�u\T/����&��;��Ip+��ԠGc,ңoFH��&���s����nl��7�)k��m&���&��(��㺢~	A�;/+�e����fvL�Eq�p�9L�TPvH��;�f������W��_4��!/9�`5�k��Y@~��a��H�Y&��b�,�zD�.�}����#Fp�R�u��X��ZFzl�i��)O( k�g&)����Q���
H��+A�+_L�>L
9�%��C:R�wD��(Z��3�����-Hg*U8��&ϼ��*�&�u�o �Z6*W��8�՚�:�
Rx��{����4�Rh��:=��\xX�. ��8T�Q�+�np���TNkm�����Z����p�m�7i-Z��"�+�`
�e|��D�����z��P֪��14C���ۮ�����P�jt�3&�_�Wƺ�XPY6Ą@z��Ph�b<�B}�}�A*`��D�N!�no"��Ғc�_����VԊ��;��e�'���>�� �!ꕄ@��\�wG�7m�ct���)
�zz|{��(E�&M$\%8�%�L�������Q{�iW��;+�*{�Z�)-�P��iV3�P�T���*�#6�a�Eَ��q�s̺-_�	�$�lB�#����f{�x���<��l`ڡ'��x��	���BQ��:�Oud��=(�bܻ1�$�����?���=|޳��տ�_=�-ɮ��{��Hk�wW�%�=��T�;@�F�o�/�H���1�mn�<Z�D$��V�RV>F�~^,��Ӽ��(���R1��zJ��~yi�����4Sz�X�/��}x��/�.�e�C��\(fp�il93�o��d�ł�KS%�w�xNٿR��n���j���鐃t��[z.�+F�4(T�%������reE{����-��o5�2b����%N�:�?�w��=P�Ӂ����������Y��r{�u�߽�X���Ol
G�Ɖv��d��jɇ�WK�`P̞��� �g#�)k_z=P@#o렵�(��}G漗�G�������s���<ezY����z���!K��!��xՀJ�Y&D���e	�י�f��48��12)�:�'�	ג�3�d+�����y""��#�G����4N�Qމ��>��@������X�hwo�$Z.����VS2T��7��P�t�l���ٷ����Xz"�)���˃3�?���g�7r`����ի ы��-bP�Q��1��M��	�E��#�ۆe-}���~�(��y^`�
O���Dw�ш��k�e�����9^�D��ZR�d�K�)���-���zZ�s>>��~��
�/N��G|���#mw.��y%4��+�L�g"��E>��R�2d��%����Q�h�-���G��)b(ay�]��&s�F�Q�F�#`�o�� 4/Ѹ'��W����$��Lģ�;뜒0�6`w��*]�ExahM�������l���YԂq�ťG�=�D'�����7�n�e �)�Xw[�Qd���-�$�@A����d����AB�W�`�!s,V)�����Զ>�a�o�)"ϢifM�=�M�����,[���!h�o�Q4M�-ԑ�l*��J��!{
W�*k��n���jhM���a�p��	���Ĝ��f�@@6�T��"Q�?eGY}��KW7A�����|����,h��vL�����צ������W�H�i
�)��w�q�ѧ��}O�o�D�Y����ˁBp=̀L��	�7�1�*�Z�zK!!�9tu3&�u�_��%�4{S���MR�fG��[�@�
� R�N�?I��s�d���v&R��|
t��q�T	�K��'U��������Dc$I��
/�\�d�n$.s߀:P�	��U��\9�I	XN�D�i�N����������j-S+��{fŤ�lPnv���'ɡ��Zh0��z�E�݁����=mZ��RE��b]d�� ����7�������	0J���#dp}<(�����]��7�@���S?���.��(�3֜a�N���(��lBT�~�g'պg
cj��Mx�F��+A�_$	��%�?�OX"�T�$���v��J?��GbE����A	%�=s�k;��Ev�z�D��Suf:a� �xw[�2O"`�.��^i�h>a��:|7F-BD�w�lǏZ�~�J�?�8%������R���l�o�3�QZLŒ����ٍ��p�,�aA!o�kW�k�ǂ�#=񃪋u�y��1���y�
�V1�|���.f��Y
ߌpG��Fp9b~f)l]f_��a�Rdt}�	�����2�O_$�/-��O��CD%�#�wF�Bu͸����/�1B�R�,1�\����&�y��1��ns\)-#Uo�Ô�O�c$pW?m
ʜ�<>i�K8�|+b2	��f����^IF\�I��rk��E�hPe�М����n�������lW��(������8�Ԁbz������j,2��L�{�T�
�^��u�����K�3S��51by��
���OB�?1&�.+�������]yyn��m���(b�.��#��NXUK�W�)W�����/�fn������\�3n��G�*�!�HCIp���(~Zl����?����Ȑ�3��)+ҳJ���2�Q��9��O�'M����b��)�)K��	I�A���Gx۱~楃�XH3$d�y��B������xż����z�U~
K��|�{���@����~�[�����]��"�-j����.�ZSvp��7ި4�t�N������R�m�ɱ����a�[F�o������W�Dg��7h8F���˔Y�@� _WoS�T�,�^�J`W��;`*�O��.ၺ���H��F1�X��G��>�<DH��~����+D���$xҲ��Q�"\U����%|Vg������$O$(*A�ʂ��>�fx��a�Vo;��� ��g&b��}F~H��� �C2'R�jP�N����n�jn�Uְ��
��Z^s ,-<5�W�\�lUJ`ޘ���4)�|��o#йM�~�<���~m����s9�4~���fOP�]�����Y�����"J'�E��:��IgJ�,H��KJ�e���t@et)i'ӧh�{���rJ֜8�<\ �tl�V�f�E���EX>��5�N��<��Qq�tn9�I��t��{RѾ}`#�5qY���;.Ӈ��8���(ή�;��:�����8d��G9����˹�7�*�9�0�#G[N��	v�����z{5Sl�d��#��Yu�w�8��P� �i��T�y�$7l$��AH&:"�"�K�vW�:����A���e�]���]���������
c%�D���F�<bJI�l�{�˿oB9q�U�{��ㆲ��L��+} �Xt;�@D�Ƨ6��K����Y3�Dv"�r[�,K�ւ�OR��3�K�%9��W1��i� AX,),>'%�H8��f�elU�56��@%7�T@�k���~�s�bELL�R?�[�Y��T�&��).�:����V��է_�ʹ~	�',޼��|��U�4X:AN(Ut4B'T�,�*V���7���CT�>������홝i]��AzXA3I��J�M<�ۃ��뵉��G�V�၇�a�(w��-��H����~> ��35+/�4����J��vb� UF�EӪ� �S5�Ͼ�[����c	妇F�Q��Z���ɢ���8ʤv��u�#ȇhQ��̞�o����Ra5����b�����*�ڥ�Qb Ѳ�1q�N��{dT�Ǡ����Q#4���hLL# f!�o�y�{-�]39֠�VYGyo�:)K!�I�co�PsR����9Q>��SqNߺ��
����Si�6�u2���5�݋q	T��$ژ�	9�����R�x�dMH�Cq;�X�;o[&��(��4uR��8+�1�/���<0}�tt����vo�Z��?3��W�e�M`aoЄ����|�xc�����2�Z
! ���-E�����������hC�0ͺm�8��o��D��Q��>�,{Ŏ%�3'�e�`2��S�4d��au��(�Q�^���/D~�&�J�Ơk�Q��Z�[���=u+�y%TC`����-!
���A�.�d��F���
��XU�5�_CM��q�]q��t�-:�����l �7滸ޫiO��׶���1��%�M�.3�R��8�33T��;E=�����<溎�}�3�L�Ր��U�f�D�a �m�g��2�i�^�
c���H~�N]��s�ok���K�M��,Y��:�ǁ(}Q%��X��($\R-��H�N�������ȦI����m�q��?V�wFGC��-��h����� ��eƓ�v�Lx��Fk�ɥ��HO7�M�t�jrע��$�?k�LI�3���j��/�"i�^!�}�$
u���.��O��{m�=���N��%7���1����P�s �S)�M	�M��P�����F��8�%8��+��_+��۾�|F��{�ӈk�=�u����eC�d�n��(cLu%�>a6�B��eJx�q�G9E�o��ʧdP�ՁT� $��T	�@I�S���x��1���i��E!����j"~��8PO���	����uk��gf�<��@��n�M��S��������Ζ+D��#�bh�9l|��.�drA�i�,��a\��/��o#@�D����D�Z~��J~�����v�{頺��iP��~����*����®ݠ�mL2q�5��y{j��`v.��OS�7��&P�ED.8M�I�М�iMp��}Js�x���I���M�h�޳��T 4KJ�|K��M%�~�p���z��`��n��9��{��������5�~�=���٤~L#�(D��p�&RŶ���"M��W�ٜ��g��]@�G�US8Q{5	g���w/� |������`�"�!m2)hc�"���6$|߼��< /�H�����;�DP+b�0�U���F���G4;�#��)�Vs�����j+��۴
,�Z�q#i�O�Ep�]���`�O��ǭD���0��\��3 �bR��l���s�0/���w�+��/�X�ރ���nм7fu��pz�����Ϩ����gkt����	�u�{�����@���@
�߱_�R��!�I�]TDE��C���y�(&@T]\d�����n5��/
L�{B��;�?N����]Ν\�׫?I�i-�.ٯ���Ǳ-�>ֶ�ƞg\ �o�j"2ߚ���q�%��m)��^� 7�\4v�+����Gk�KW6��~j��-��M��a`�/،�]�r��VPZ gCW����oV��$�W`zN6-t�44�X��!��,si��a?��L���;�2
�m����f�r}|,��XC������w\ڕ��H�BH[�������k�$���0��EjD/e!~�j�.�.s�
$*����5�w��NB�<�V�-}O$^�5գ��9��VQ^q�����Ӆ�H�����/SNQ���Y�����Og�������0�q9Ⱦ�������3�F��,�R��T���܂<��;���<�O�l�>�M���>(�
j����b�!y��s/�$uͤ�~��9˼M��P-�':c t������^��-�'���.݇͌E��s�$�j\�:���qk�e[/��3-&-N��n�4T<_E�m���sa:��O<��W%V�i�M���F��C�^�M�G=e��M��u��㧾]�?h��ͳm�Ω6<�㨠k@>��D���l�1�mJa�>GiC��):��UY�@gW���h�	j��a���i��;�i�_���[^4��@� ���	�$���ř���U���K���S�lMQGMm�}��#n��h�!�9�����ZI�
����0Xwi ��������} �풾��%����֥̃�m���yTLq�qͽ��:��V�ӱ�tj�;�B�M�i%6�3g�IA�����r��R#���
Y�*IK������D����@dB����7o��\!�ŒF������ع��TU�^ �Q�TA*�<Ð�95]�Df� ��y����r�,J�^��}�zS�'_�hT)$<��,M�����!���~A��`鳲�1 t�^�}��pՠYy�}m�?«�Z'��{���@��eY,I���]�(�����
�8K���Dq��t�Ԇ�(#�2C���}>���e��sf�!�D|@i�)�D�� �E��ˇ%8�_��)�T�(�Kݘ�?++F���s& ��yXz�E"a:�����y5 ��B�7�ʎ�<>��r!���s�E
�RJV� �=.�Z?���Ͼ���D��p�DT���5��osl2P�Q�����Q'�ʆdS���2�� S�,IUlź�@Ud�2eG��n�,�/ts�la�.#$�Z��C�%�9:r鍮�e��B��*2C��սȆb�="4�|}�&��u�A�6�%���{ptև��o�]���˾�{�<衜��<��.-�\[�L�P�;+Fq�H��;�x�`�Z�uE�b5�m?����q�zN�l_��`�ʛ��})�/�df8V7����+���@���pT���& ��^9�#3�=H}�M�ԭb�i2���P��BUs������"1�ʔ�
7��چ>J-�����(���%#����] 䤓Px|�%�+`�ـ�ɾ�k�v	R\��(JtoJ�_ُG]�����������)M�f��^*�����3���B� ��M�LnX�ޤ8!���Ġ��y���cY1"m�er���"����=j��P�!45vr���N��k�����6eR)b	���.�`c�M����~��Wg�es
��!�V�1����q����RA�#,<.;����Ѯ+�mq��ԄU�%��wm�]��Ó�؃Ɋ!�#Z�(M�@�����v�,���*�L׮�Ua��WMor� ��H�昴lU�3��Ҧ��P8^\��~_��iD ^Ty�	����"N@<���EC�1(��t)��#�j`���0A"�-a��]I���MP�H���[�ך��@�J���~3,��;!	��7��ה�ۓub��Ā���C��O�k �X�w��M�I�Օ-�֬z��>�$�HK��gj�g�?��|�ht[�2z_�b`�#�Q��	%��H[�� �yĕ�`e��`��T�V���.6��z��h�,�`j���3w���w_��#��Bx?�gB�Ԃ�m?���sp=�p~���{x������Ȩ���/�pH|����$禝 ��;�Jqf�����{���]�uS���$�1�êHC��̿�9�]��ȅLw)�ڎ���*6(m��{B��_�lج<2�r�	��>i���mu���i���̊�w��n�ð��G�f/�ԡ?̀�$���7o��k	�,o�B~��tV�i���� tP��i4�'�P#���� �50�c�H�Z��֫���D^�k��ߑS��w9&R--LI]�}��S�:����<ܞZ�6��)Pd��Y�$�X"����<�Š\�{ZB@�%�6�Ry(#���O|*�`�͠oߝ�y��d�˝M��kK�>)�ώp�C2��/N��\Ee��{�-����i�BL_7B<��T��G=�%� 8�\��%���a7=�%C#��2s;����6�i,�8Vj��Cf��o����j�?8�bQ�\g$��<lvB ޱqLt�?�'`__
WDl#_Rx;i�"RA�RL��fd� '��J�'35�uA�����t,���O��J�Ϝ��`���$��׉?��s�˗����jU��5�E�W#]�Ps�?��ךAr9ٓ����\�7T ��������D�.Į���>x��?�ӂwq���5N�X[[|w�'��=�0�x��z(�NyB.�Gq�z����O9�fp\�DhyO"��,2�J�)�

��R���U��8�!@d�)m����T��){��&N�����w���N�tuA-�b4�-H����B��5lԻD�h����kٽ���\����̌��b�"��bش-C���b8����|i�EAE�,�V����>��ؑ��_`!���M��N��戆-��X-����"}9�ߡ����a�Ɏ9�?�!�Hk|�Lݯ�oc����OG�s�y�N#�[
��� ���<�ݺ�)M�.��Q��9[�w�H7V8��<9��Gؙ4�����zC��m���i�D�{�7Cg&����*p��z�������7�b{
@@��}�6�B}�������X�G���{@�jn>�a�Ŗ�#�>���-uE���Ө����|(��6d#�CtQ2��Pղ�.����{N+>b�fk�@�HxUO%�7fm��j�/OЪ>w��4����M�[��[�O����/"݁�_�\^�Eu�|��Uo��y�܌a�o��%�m�4�/d�C�Ttt'?󠵨~�Ѣ�p�"k�N��og���ĸVt���>�8�U�+K q�D_o ��$�&�*��w|h��ף���S;�e#�C&~��oo�G�Z�9N	Ж,[$FOE�^7�?��"�_�~!=_EBK?��v��r_�\��S͙�6�*��|������g,h�o!�R{gσ~*!��*
&{�qx��Jf�hx"�Ǿ$д�0�@�V��A��7�'�E)��g!�r�*�<��2<hg?���Ec�28:@PAd�.V{ηu�{%$��#%C<��*q�Z$N5�"�yj.R���j�fU�9�:L�Yo.�M~N'�<z�y��eXC�l���u/�"�2���
ڿ�4�	�ϩ�-��U�*F�!�
̆os#��QPޓ�N��� >�Ir���1P�l���d,��p���CU�nO�v4;r���t�����Q���~��Gp�r�V���e�t-��qw9����Q:���9�H�=���w���6`-��lж
�_�m�!P7x����$p;!5M5����A��>�{��߫躯"�-\ʙRN5�����)�@XJ����#2��H��O�F�I�4��=|;�Hgkִ��roop��%Q�)�oRX�O����wp�����y���`$]��I�8ȽZȏ�%[�k&S�
�G+��Ip۽E�J�W��@��QR��aGwI���U���|�)|QoV7�D}2�gw�#s��[w���M�31|���GI��d�s�)��Q����=�[qF�䚿�9;��9��O�<$u�]��;9�ˑ�5>P.�y��o1TZ\��c^Ć�ԙ� I��^�A�d�M-�������ʎd�H�֭J"�R�g��|����δ��2���ԓ��̢LS��<��iR��j�<j����l:�3lW��OH�ݞ�?�Lڗ�yŊ�u(0���ټA��߁=B�>���f>��[c�Ґjd����P��vn�J�9�Ǝ�/�-O�}���||脪P����suCP(FE���Fo���!8RZ0aҤ�arÉ��y"�r[��=x�ԋG��ӷQW���ػޥ2����� �������[�ʰE{՗m�7ө��L$)9V�(�!\�<����+-F
���($�lI���9m����C~�ng|�t%px��,ס.�����`��8�����O�͔�J�'A{�����U�&���4hZ/�ߠ�>�j�*23q�dy*�9����;�g�\���\�8Y��sy��綔�*�m�uUm�c5o��NGE����4�tS�4��̯����i� ����8�?�\1�0I�LT�W5n��A8��4�;M�.�!49�A���}d�:���'3���h]��ZҞ���T��$��1�z0�I\j�w�(�b@A���)Y����د�1��[5�zی'��`5�`��03���Q9�A�����@�~��[�P�D;/C�q�y�_���(�ip� E��ޣ�a�0DJ_��\��ќ�����یQ9S
l��Tj,!v�T�c��@9P.���.6c�� 4�� %L(���A	��b��G0߇}��IW7]�:�4s
��^V��%�m�� ���э�ĳ?��U6�;/@~��uc���³v������ 0U�d��2t|-ѹ�%����::*�Z���$�BM�������e&�K�6S5���f��s��������.�4�bk��! u����b2@���$��0�A�v�X��������)����N����ʕ�E
7yb~D~����/�վ��iL�X����{Y��F�*կ(G����,���n)���Ar�����W��W���B6�����~+�7�jL�����V���ǃN����l�B�գ���Un�(s`E�~���77�K�i�8`�Y5v�X/��rEA.9ml�;~{N��>��:#��f]�6owb��t�d��Bwt)7hd��ڭ�EA;嘸���r�b��!�ԥ��	"
�aulr��/$6[���P��M;>������C�;3�^@����S����d��ŵ��x&���K��x5Z}b��rvܲ�R�0� �wz��	�=B ���o��B�D����2�?�jJ�:G���C=� �Q� �S.^Ս�H���7�~��A�j��	�n��%��������_s���hݚl��S|*�y�ʍ>�ɖ����W*���6k�x �P�؀�a�9w���;����+�o���Y��XL]mľ�����6�JkҘ��^p��|7''L�*��,\n�̣� PxB����u0�f+YI�&�{��M�f�B�G4-� �<�Uz~���i��C�U9���48�ՌA�lox�\gר��Y!�<2�C�OM�q�Z7h}ߍ�X�ٞ*�r	sr�ڠO�ڑ��sG��if[۴��O��B����q����Oܗ���<`|L~��HN[u���Q�}�m�ց�+��9���DZ�ReK�,�gkW0�~'D%14����v}�Zہ��$>�+���j��~(��^�_e]��Z��CF��g���X�^{���X���=�:�3�f413�=7ʝ�L76G�0Ik��:q�M"��$�l�E�<�"�&�� IH�8j��^'B.t�_�`K��=��^�U��s��6�~Sc�����}Ƴ�%�w�6AUZR�ީ<�h��c���ξ��V�s���UN���Qu�ZCi�}���XNm����Ŗ��q��(@��Y�S}��Ս%ֳ�x��bR�<��'���,�m�ZE�V0#17Vܪ,�x�^O	�&����C��~�,�E��k.e��VH@�� XO�niB�Mx��� �_��B��`�7k�nx6O����g�ǶG2�j ��1�0k��ﴴQd��u��|����z��g(��ags	��_�*jkf���tƩ�~j��tۇG��~I�Vp+�@�®>����O�r����s����9r�����PBe��x�6����r��K��V�g�[�y�ѓ�2�0hV��Q�':��C4�X�8����O>ڝ?��N��j���M�d\�o��� �+M��9��2���Aʂm���:��RD�GF�?;��$�I��/!AG���'q�7�X�(�D��tᦝ�|o�2l�PV.����(��B�o?����O���<��[�ypZ��˶���GB�l��q�m��+~U� ���k��*����d7���s�B�������
�%#/�1�O����Q��2�6�:�|�5b��1W	͌���O@�'ƹ����h�W�6��S��s5G���ʥ��@�hL��{PT�8�R�N�"0aڬt��,�YdD������8vŹ-&SC�<�1�+�[X��Ɵr��I5��c������f����U7L8x�FЮ�G���*O`�{L�f�7��|�8�!�`�/̗G��Bnu����(�:��!�Z�o��[]����K�_尐�p�	���;;ی����Z�B�'���ͬdx��sJ�T������?j�	�S�
R&.�G�y_2�^c���L�H����=��|�'�B˯='kuR��vF�\��X�e�(�{WbLv��fV6.�ь�c��Y��Yzc�́*�;M(��s[�?�Z^�pk܏{=N��:�N�z�w�fg��X=W~�=Z{WL�SR��n⽏��>r똋.CÚy'吿��U��7�ceè;�Lox��*��Gc����'�ħ�y0q�����}��~X��?��L�U�P��m������M%=Z�2�B �����>f��\�(0;�w�B���F�Ԥ�)�(=	��(��ciXq
�P�ϵSr����X��:�C{z+I���.��: ȴɿ��`��#�������*j]Wd���>!C�PJ�	�RE�4ڵ�7e�2e�a���|
�-�%��**�[K���R�B%E����LA��~u���"лU��:ZLӻ����e^ƚ�O)�p6���.z_�	�aV�7?̹�c�s}�?������ ˤ.��n�J�ý��c'1��d��t��-6�#^L�D��-i�Ǹ�:{��|
G-D�P���j�Z��w��6�E�%�J��j9������׵��cD
�Qن0��"
�th�7Up(�l`��\!��X�ohj�2�
�>A�j���Q*j �nd�A��2�V'�X*��)��e�Nߔ0���2��޼ΗP���B=�%��a�xP�<:�����(bu��y��� /�.>����ӂ��T��E������·r�Y����?�/���Ҧ�	t�I=V��5L����e��]W�:��S�H��g�����`8�06 �����M(x�L
goi��'�A�ɢ�B�5���z5ܽ�q�#e(4z�+�H7�6K�)8�7��h�_	�l���r�����*���éEH��������	� ���7���Z�WQfQ� �kw�?%�9O'w}_2�87PJ3�(݄ub4��z�E鬣��`����ﶃ��
�ڪ��)�o�:��Z�� hp�����-�[2BC�e��X�mܨ�s�ѱ1���ga,q��X֢@�ʝ�<�n5M����#��,́���y���1������f�Uk����>IHru�҆MT�Ht5��5�ڠO��?�R��� �7�M�o�����a�uN�
��/����p4+�cWE#�1�&Xny*Ŏ�huMliSf������yP�X������v�G���(���[)� ����U-�
�Z^ւ��u*)�n��*M�����xE[�O�;H}L6�،�R=�ìE�=g���Ǌ���8)	tÓ&��WS()ب���R��2�H^W�ߩ<��2� �g����>?2����&��L U��D��l6_�: V2�1�'G[�kz�x�*[����͓�����ΟN��:�Y~Y��N)6��?G4n�0����nF�)��y&C9�a=�	%/��P�}�N�oj�Hd�`gT�ժV���M)!/>H�N�7qJA�Q�HMZ���o�p䅶ZtP�Z8�H�7�͚B̞xß/��\����}�����W�>��^�IS�ӿJ`\�$��w)dL՚��;N8v��N(L��&����
�D��"�g[�����t������+eF�7�8n��Y���~��V�S{+K�F��^Mgi���P�#�+0�x{�I���NB�=>�p�.���U��'�2�k�CpL�^3���'U�o��4��J�+Q��$������#�ƶk����<N؃1��v��X;8���^��Z�˨,���<ɻ ��F�U'�M��k�Y�:�z��`�G�jo�eu�{����(1��b���B	v������;�����2��B�y̎��ˡ�,��qp��>�u������"��^E҂Z�=p�¦B�Ƃ�W��)ϳwu����ߝ�,�3z�ȟ���h��=S�p�ZE�F	�@N�tI,mL�%h:1X�^�ԧ:J���Z0{����P�_2 �ė���k ���F�j�HV��HW���M��� �󁥆���	�(�T�9QnU�)& �L슍�c�w�q�̋������L��ϟ蔽5��;@)I�`Z#�%f7A�P���ʎ���9����7_HEQ�\�p2@.ئ�	���#���gf}�D�9 �I��
IR^}���=�}� g�=j'u#|f B� _}�[
�b[g��E�4o������(=Zn|�]�.��X�@�X�7);H1�D�@���W�zf0�;j�����yH���^��	�F�![��*8�,��29�<�\���N���́F�"	x��s�(0���}�Wj�9s���]�al\��A�_\+�*2���T:N�.1H��� ������тð�s�%����ݑ[߁��H�.�]���̱g���Z�ӵ�3vRJ�E�@�������|©��H��틗U����M,�"�怓���N]�PZ�쯗�[*����++�ƴ�Er��n���OX�7��{G�C��#�?eA��>a?�4����#����.4l���Xj3Z�Q��7"�n��O���;O'I�TLEt�W0yҕ\6�����{�!4�V��Y,�鳊��/r�]�\6���(���V�I�Xӟ���>�|�Gc�EL�Ek��9 �53;�Ne�(Za!�e-8Ly �����]L�q�O'{�W���q��S��,�$4[�Q��\���S%��`cz�Fƒ>�����[����ޞt/�����Q^��-|b�PB�ټC9�N������y֨��@]�٩,R!l6'���A�0<�xyB�ur�5�;<�$�ZmI��4�L�C�9$݋_�;(�>�0W���}�9���&��Wy�>3p��"��M�|Dn�����l7ښY�v�`U�{kyسRk*p��=�Z���r㌽I��0����po�)6��H,r��n)G
R3�/�'���jmP,d-5������g�՚��]��v(��c�v��j��d�0�f���{��U$����l�'gD^M��h\�kW��Ӄ�'��G	��,��f��c��h7�t�7��j�z	rkcN	܂"��6)�H&м�˯颜�CR8?t����p8�\O�N⎛���֯�����Qy����RW<��]Z�j�ڊ$�i����42�+@}���6::��̓�W�<c�c���8�f�����ܧW�����N�,�-���tՊk��pz0r�ü̃9������M@<?�I�Z�m?~�?+B�(�<E9X�0�UF�����)���>j�D)�zU~�y��·�l�rE�Ø�R`��G�FS�	��&#M�T��VowJ�!6715��He���j�(��M�gZ�%�tE]A���J�yh?��<7���7��E[�8�0�4�;�����*��Tby:#<�{϶��b�co�A!{ƕa����h�B���t���>T*Ĉ�0�3bM?Pd��J��IHG�H��F�"v��k��zx`1�#ɷ�m/��9z�;�����W��f�~�R��	4���:h�QV�?b?N�y��X�!�_��y&�����]��:�S���3Y��O����u����ހRQ���.s��En�Ȝ�O��S2�uR>��\�W�������a�g�m��\�	����u
m�7<�CQ$,]7Hؠu���d�:�@4��������d�C�{O0���k�6iOy��Q�"�v&���:���6��c���1.	�����͂��/M�ly�t^�y��'3��_��CS"�����=N1AE����ɬ>׷�V4f�S�Q�}Y��{Vy������>3���JdN}ȋ]#�P_/�M]��'3�)j��/��� ����1'�RL-�?���n�~6����0����5!�ja�Sizò�U=?�@���
w���EA���V�T���9�ܗ���� �B�KR`�x�����+Q�4�i�P=&4M����]?��ok�	M�UZL+@2ǥA���#`Oz�D֠�f��"tW
�J��+QD{�75��2�"\v=b)cN+2bpâ@�C6��6�
�f��$lrP��u<��C�`���A���N���hmb�)��F���ۛs�Q��a����3�;����:��{Z�qu �n96Y�Z�ٙ���H�5.�	��ۍ;���5I
��.��2؊���ȼ���ĥt�� ��P4��S�w��I����j�4�73{-!L+���nߴ����3���=�����]Sa �w��a*�7t�ȼ�q:�~�PШ����N��ӵsKh݇�}�.0_��{�Һ;�����#�>Ʌ�C��4W�I�9��&�~N��9\-!z����Ų���W��qR��I����/&2Q
.��O��Ƒ��V��Z�~�W
��T��ɠWǚ�'n����S��s�a�d�ɼɭWʤ:����٠��L�5|�]�!�L�^��<��lK�}�JE��{���J7�wCȸf ��C�rӥ�	w�V�s?���P7������o��M�SW�H�٣�D����Q ����e<ID�g]B�G�>D��IY��{���N+����jy�XIRv�C��+]��V����a��/PV�����'U�������zR�!�@t���q���wE�SC��9Ε����PAWy�n� u;T�1����Sp���!�
���Z~��3�������g��f1�����+�0��Z�=I��Q+f��-�����r�#�w�L㌌