��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O� �R�d��/=���H�/�~6R��2q["�2�*�\'`�y��To���N����"}Ԩ�-Y����Z�Y&%cA�'k���C�>�=].x�>~�ONU�4�,PI�ѓ���~ѕ�Z���rZ�DG3���}�+�}��{���޺H\�H�Ɣ6�2)�y?���'�n�A@��8�<�y:X������]h4�G�9
�����Ƽo���.ά�-x����m��ϛ耖c�Q#�/��O��{�7��(��n��WzT%")Lq&���L��?�{�A�/��|��l�Vm?ޘC7f�U��~VƊ���f����߃�GS��,y�<��yɹY(	��~��h%[�䙗d���_�����:�ر9ӎ�kGȘ����׮"�gun��)���g�͹#��k��Q���2��������S4�%H��F%T�MJ�=q
U��p��?2a�M���X�&y�[Qy=�\n�D�9�L0U���Ᏽ��1���"�r���sX�gO��Ϩ��~R��Q���L��h��.��֧.���>=�I�r�d/�-3Q��dY7�9{�����@���0�=F�?Gx�~��@�p@U}	��g�3K�N��.M ��n��E	�.��WY4�=�.-��isw�	/ۢSI��h ~���gi�b�,�<�b����!#f*���I�}۟8��7%.=��f�~��Nw�$PС8>4L�����x,V]�+�|��b��vn�S,��x��"�V���L-P�xz̪ٝ�XCz� ��TF�4^0�L]um�Fk��,t@��>��E��� "���))�� M��kI\�h�Bw�\��Y��ۥ�Q�T����.:]
Q�=�ĝH�Ԍ�"�3��A)�
5�$��Qee�H��/K����^� c��$��a��~ǩ�{'"��av�{=�P+��:�yy�<�� �/�e��H�� &�!��<H�p���h!���R{��qB�qnI��x!���������_����Tek�^�"��A��f���2�A�����|a�z���X8�FS3�\)q�	�`�?��_�K���v[ȥU�������H���I�_�!����o�)�ՠ}��/G�}�-&�q����^0�j7U��iW0�����LI���X^�;�L�i�(5��)�p�(�v�x���l�oJe^d3�� �K�� ���R���F�:���?p��z�J9��?0�������6�!�U&�úRv�\�H]0�,R�T��	Z�l�{~���?�i9��&�s�XV��6G�qՑ?E#�)���7�����I>����?h����_�2]�3v�e��ϣ�%�[~u*��ɶ�y@o�5�T��/(���&�	z�����S�L���0�s�
��S�@�!곁 �Ϡs�B�
�7�b�R�ԧ�Qe(�]�f%��n ~��2մ��/��R�_k)fi��®$9���ի5�?�}�U����},��ݷ�����'�d���o�h)�����=�� ���C�vy�h�o�y�ȹ��A��7��w
�f��p�NT4��V���1�/����$��4��3;�uD识�5��ٞ�+	��]P���33�G+��ܾ"�c�E/X�ӹ�.�s��̈́�y����%��\Y�km�վPκ|��{�l��)+�.�ٖs9ͭ(�
������&�#*���9�N'��I�ey2x�=��d�$
6��f��%������P]��o��fr�R�b����Oq�#J�f{�`
�J�+�ꅠw����T��������E�t�2G4z;K� ���}��#6��!���7Kj ���<�,(O��,9���0D���oU�tT���@����P�.��AV}c19�Щ0v��!����5�(�#��~�%c��ќZS�0�O�/��}1`|�_���Ð��߉A'�?�A���BJ�.��4�ܣu��^gie��^`��=����$A�J��O���tU:��iz6 kxD�۰�9����3�6���|<��qt�,m5[��g�P6
�&Bc��f�31&g,�;$����s�&Vo�Y�X�z�k��XU����KװB��29��a vv��u7����Z�>XSuw1�%]�c�K�E,ZV��$x'�k�j�}&f\�ZU����Y�/j0r��h'<�N#�c�[��~��Zt���i�IԵ2;j���=�%���4�p���^�<�5�fIY�؈wP�@cF��#�b�������Ղv���Z9/������C#M���e�G�Ү�[��!	e� A�����g�C�F���k|��p�Z5��K5���e��c�֙�.�9��߱"�{�k��*�մ����IAH���L�s�m�C>Q�\� 99ż�ͥ�����Cź\J�|�@���LF2���`��ҝ($Q	!�)�d�A<�>�� JbV�D�B}����"��E)�'�x.��7�TK�+�{�}�FT�z��Ek�L�٦��
&����Tj��I^u*��o!V27)�'�	�"ET���q8��.��Ֆ+x�Y��WO�Yߚ�"E��i�ǘ9֪UE��qT�{�y�$[d�CMW%������>֌c:���V�cnz�$���2 8�����.W�z������j6�;nS�C[�6,<!���d�-�o���� ��-*$(�ql?+��in�0g���Q��),v�km?�R���Vzׂ�谠��υPY��H�67��X�����]�5����(w�j4�p��};-��d�,�H�n?1�V�8�f�s٪]uB�)8a�2;Q>�0LG�kc�V%?����-����:�_�,�kL@��5��-�8�* �ؓ���	����OZ5��f�L���|�͹���m4ŴZ��5(py�YV���u�6z�d<��	��!�}y�@ k��	�\�;��
+���1�Ke����Zz쪘T���z��w�Ϝ�ͽP{��gH��W���}�_;NI�𱃑8H)���1�hkDFӫe!�r�WL�#�:Ε>ݡ��(cW�56E���n�
2��P|�-�@��{�ĳ-��`��3��苠�_'���0�Tݻ���uu�
~1E�K�����$�q���@j-���KB�mE&�9a�>��6x�Ir]�[�N;�w��읟�J�9�NF!$�?����Ǒ;fL��h���.T:(e�G䳧��Ev����I6������X��w�<�w����c~H�-��i�
6Q6��mnd�ˀ%Rl9/���Nւ�Ss^�W]��f2���oC5�08HkČ��ɢ�ⵕ�@�'4��Ҥɯg�(L��͠��҆Or��a`�M�y��D���pFrjF�Ѓ�O��H���+�8����WY�
�k���H���
�'�R ޚ<{�ېD�+L�m���6�&��'j����_5Jxd$���P����Ty��z�b�h7UvT�O5�HHR#����F�-��p��?ٻI[��&ъ�O�7:h�H� �̷p�Ȝ���P���O���f��K�]:�>I��/����������V�ј�Z��T5���ݡMq�K	�cIg����pl6�|#|����� ��:U�lC34:�����S�0l�Bw�7���C]aP5�{o:�\�����"s�����f�K��p6w��<�;e!�o�Ƴ'���+�_�~~�8B���`�D]@v-�x,���Rm�6��L�N(�7��[��˷01�:i��l�Qk�j�z"$z����l�p%�v��<�jRp/�JJ[9���]���?�G�݆�oW��vچ>������O��m�!"�]�lla�g�\�L}d�\�����q!�w許ԧ{A�@e��H{±�K���R	�bv��PC�����XTH�&@�o���X�:�0;(~Z�����{��'tM8b��T���hV�.,G��5�@��QR���H�sT����nP�����;��z��ˋޡ�>��<��6_j[�G�ٱ�徒��$��;5����z���0B�����b(GK��Z����k�ƺ���8�>tמPtnᝂ�x�`T���v�q���'�ۭ�,uZ�{2��q������I�Gpq"�yu׻`��nr�� �nG��<��]�TH�"��&�$���?��.fD���U�Mf�}ۨ�����ʮ��p�]���ܷi�̘]7�W��@�M*��WKn;�h�jC����|���ѵ���(��w�n�����fֻ��N���q�����p�|B�������9us\m1B�%A/^z��ih�
 �@��_�ͭg��̒	�.�#3j�,�'�oD��$��fs,�ݖ����Q
�[V��0w��b��-�<���J��D#��,�}h}��$��$��Jn6#�C,oV�,�"<���ۺ���t�"X%���$���'e.� v`�qS�Z�ꙹ6�� ��ׅ���I/Պ��N��6�E�O#G�W��X	%(_k�M4��X6�(�f�g7N&HGVxK�/�������Nۑ��*w�F��n�=H����pA!;N�O�|�jh��ȇ�)�lT$�	/�j�Y������]|���%�ڴ����8���t�$J�"�!O�x�R5��=q��(�m�a���_8�?�N�j|0+�L�u���]v�Ȫ�<�3���<d2=X ����53�uD��ƭa�N��|��~���Z�(���6t���� �p��E�T���	V;�G�sy�&��7<?F� �~H ����:ה�F9ǀ���kS���LeǮ��<�-;�ʡŦ�)?$;(�����p�ՓfP��� <��D���f��z�U`��pV6͙�a�9Z�n���)��[��Q�#��I�b^knt�X�|@uoe6��6l��Ln���`J�ơ%.�ȟ@q�&�0�`�e�N9�o��e �W�eF��:i�a\s�nL��OI���B�4���y{�Y��Ŀ󡉶���|>�q�U`u���5N�P@Jr�3�C�2)�И,ܩ�:�I�n���=��/Du������͋�.ڃ�=D�h���7M?��ogI�O,g�ֻ�:��"]ģ���\��?XH�P	��F�7���R��[�c�<�s��e3���pܟՕ7#���1�&삂DCnr1��RG;@�2������qiןf��\��n䯢弎��2di-�J�n缒��;�ZS�!uN/�{o"N��\�8����6u�P����e����P����*x�v��Z�����"N8�Vh�pgE�F�@��1裮R�g�{�zT7D��A��m�8�s��b`D_�y0p��ZSF�N9������ߕ��vR2���G�D��,iRU  ��F���q�f2;D�g ��ł1m�i��&�����x@�V�3zy`��d=��9D
��*�ə..�y��[�]��e���J�$�+>��/�JW�3�S~H��(�u�E��R�����>��	�W��{vXE7�ė1�t��r)@���}��X��-����R�Y�A|�˰0���в��7���]ni���P�*|����W�o)��FU��]�59��<���$G�sn��h��]E�.�:þ�d�K�:�8��Eb.�O����F;EܐE���p��S�T��, )?�lߟ�`���d���mP�K����]��0�'��K8��2V�Z��bL)�r�l���r�v���L[��H��i�XHw�7�S׮a-��ڡep�@9��U�l�!8(� L�]�5$&J�?1z�θ��X�O����^�՞�۽&/c�!N��Y������Z>�B.E�9H0!qbz�+a��^.=2����Eu��1��<�c&8�8��PO4���٧w_� �G��l���bOg�֑�%&����Hl U����r�Q��Ӱ���_�5b��ew��rM^�A��e��ǌ	�k��s`�k�?k��$�W{C�)"Q�Qڪ��g<��X��V+x:���|-������Ǝ4w���=Q��ک��:2�	r�|nr��P�����`�!m�ey[%�����8��J�|\�G���FD�Бz���;���Uq{wX���H�oZDX�Q�)��Q�a���&�>����C l�� P��K[3��K�1IM#$WGw�Nꌹ.-���%�E�K����]���X0J�x�Ol]���t�xa��q~��^� N_�d���ɯ���}���˧r�,,�s��^�T���9��$�\z	ܬh��K�eɑ���g��f���s�Ϸ@3��Q� �>Z�ٍ���#%�X�0��P���ԝ�٘�77jL��5�EW�C��eBr�v�O�����$޸m��P	0�O8��V({<S�l��!Ι年U�w����4-��Kc Uƴ�l#È��'��?!j�������_��Np�z͉u�r��$���2�
�q�M�4�g�U}߅[�`�hSf�2��I��n��F�
�Oo�Rj�:3����Z0
{$4U";+�!N��O �H�U��]>��yM��n�
��b�z�̟�}���0�~�3*�}���Sݯ��y�_��@`��\���Cu�L�n��_�t*���"��#�*/�n�Q�L��S���\���C�'��1Y?aEQNNfb�u���KiV`��9*TivLXʉѐ[<�����sA/�.f-�@��o�?�G�"l]�?4�/�lMv������ж��>�%��6)�<�1�+F4�t�`��G� ��w�*�
�P�p�Z7	��k �`�v�Nx�Pn�M��'�rc���h���(<C>k�"�W�V���QuF6�+����1��8��؝��ݪ�u�6(U����H��cn�iJ4�^�}?�^��^e2�������F�]oY�/g�ɎNF60�o/���-QA;c�I/�	�K�qlg_����>�V�v��[�m3�	u�nm���v/y[���Kb�8����z%X�xk��_�H␹��L�GK�-�{"�>�#��������� e1C穆�@�fq���,vc��$�T0pB!^o�x�j�n��Ih�*�9�~h���=�fm4�1���I#v?+�^���i� �l5�$M��-b�܌EB��)
�1���Ї����dĖ8����?�D��zNm�Sn�L�t������4�x��)�"�a��U`�!��YN�%q���g�V���&�I����\�@�2����`��Z�	��99%q���%A?�V������b$Xb���쯟�q��e�IbH�L| w�X��Q!�t=#=��x7��'z�𶞱y�ADhȤq^��~C?%�͕i��^8^c��e0B�w�lNp���~��^F��5N��Уxi��k�?T�6�6���Ӿ��M��.��"Xj'�s���'l�ЖMD���F0�G��Y������w|�	���(��H��Լ�U�P@{ґ�t�c?$�_�pJ:���j�_�BS�M����WS�2�Q�3��2��?w��ꦛ��t����h�I�����#��3�bC7��g�b���Ey;�Xʼ�v�v8�x{JdzB�PJ��y�>�
 _�iUW0	�h5"hU7�4����%� �B��'�n��ݾm�R��U�+S�j8v����	�Z5�  -��蚽G��eV��(���"��gW�R3�6F���S�N$O�Z�9�Z��!%��5c����Q�М.�&L���J��<�V7X4d��RWț�S1��p�v_��S��E޳yg�>���j\���D.ʯv�h��ՙ�(���'b�O�O�%{���8�!W�'o�ǘ�3J�)���g���ﳏ�իv��y~�"1\���ni=���|����Q�p�D9���,��k\�s|Y{�|<wT�u�uK!�����?J����@��JT5ӥ:�F���=V~��1@Zh}2='�h�E�|�`r�UK���u�����Z$���;}�=��U%\�pfU�=:֖甙��
��bt8������e�����T����j��Sk:vE��/xV�E��~����4"[r�A0��%n}�����w�K�l
|�\�j����4��/n��PC�h�M?�A_/l9E�G�\Tsq��]i� l����[�&��HdI屨��7�y��I��e_�t������UM@�59ϫ�cuK�:��N�~$/`��V��
e%��_s<�j���;�a�b�%���L>���y�RhK�p4]'	~#���ƴ��y�I�Ҿx}���Ɣj��9��Z[�V�~ℶ��%|I��U�J_��<`��l+|_�&OtUL]t3ۇ�,�	�R5`�(ʣn�xv��.z�r��P�ŷ��yhSh����t�J�ø�XR�z>�x�s�g�ݷ�8�{I�UA;���_]ˌ�W���b��
2��f���U���8лl&.�}���4(�6�b�E�=����ْM׸̒{�TB��Y�I�5N���T wr�T�|!��(�!�]�D�b�����P���jD�\^s$�S�|l8�M��.V騔��8�xO��&������, g���B(�	�L���rq
7�7j�>�~a�|*�_aa���v���4���zb\�i�5����o�1�o�{����EB��:���G9y4M���AL�����=����/;�l�<m�W��2=|�-�2���m�`�uy��-����߆��#��.�!�ڏ��P2�!}N�ܽ���k���S	��^��u����K���l��d� �V_�PK�z��o5fo�����CX��F�Od��y�� <)Ă�
���5w�خ�k�}�v�҃A�6x��˫�p���C�?���5���A�׷;�j-���f�㘩's3��P��{�ȣF9V�^C�It����o���3υ�`�)K�<��ȷ4au��D���%^���g5��;/o9ʍֿh�5�cJ���(B�YgH�?�C}�G��ռ#a��k����A�����8�����W-	�	�c������P�5}&xE�)�@�e�k+&3�&�~��+p3D����d���JP<���rFA(~qĠ�mE�[����A��� ��:��AȕJ��_����ӻƨG&K��o��[�!J7n��h��*C��5���@�
�e�0�L�>D��Y)Z�DI�d��`���T��ۑ�\�i��1ur���l��o��p���t3cV<�	�d>��ۊ��$�wѮ���Z~��&2�~�T�d7�͘���z;�|��y�1�������!1�ɴ�.r���q��P
��k�{��n�F��.�E�A����H7%H� �Fh���W-a���_�%�Gl��)y��	'��wq�qQɀ�d���l��p���Q%��e��鳂�-�0)m}a���d�������V��v�E$x'��k4����4!�^L���ծя;����z��Y��_��%v"j�H捹pu��Ǒ��X�~/���q�	�1�|p��4�X1����g�yC@���١[]j��.x&��Gp0����Gvdh8��U�B�\��">Y\s�X�_q�w�l7��b۞�
���ڈ!~���m0V�õ�<Qo�������F�ظ/O���Wy���ݖ����X���ȵ����~S�s���tV�c��*�w�}}����3&5�epN�LG�8Xj_ oU�:�tFE�������I�4q�J|����[:RZ�oi'.�OŎ���N%�L4;���&"Qc ͒%�|m�(Ụp�l�>`nf�ɕ���.WB��Gk@,����F�(ni?U\0�0����Qh%5b�< r
�OQr0 �|z��5}?���~���] �{S�6�8�W��pGzi�L: @^�8iV�s���@��¹Q�-rl������
YA��^3${�(����ѯ��DvE#ɕ=�bq�1�`>�\z�g{<���(�8�5;`�r`��k�;����PS���8&d��a�3U�������F�DP�P%��D��q��_h��u)g��~��%(<K::�I�� M����w4�u>{�ө�Ä1(r��Jt�I�s��$��)]ނ�j�Y��������<x���ĆP�m� 3O�*�Ru���h�~�}4�D��'o��k�8��du��e*����#�S.p�x��
m�{�^V�$d^�_!I)恣t�S��-�ji;!v/�p��"9Z�R��B��Zcş���u�qY�����R��j�j}��A'��e�	N�j��Ct*���b��֙*��xA��ݢ�ǿ�;�$z��h�O8T��׷��<^\������q��4#V g�&|�m!�G~+��)ѱ�SMo��t�1�R�w+碘��B�"�`9�
�����J���ڞ
��0wߘ��ó"�&2�VQ\-��6�3\��O��W��5@g7����S2�?��/E�"-rs�snO��C�N��������Zf�M�R���"8�PHN[��;* ��aS���P������_=R��ҺZ ��[��`?I�f���`�t-(�Jf���IZ@,��� �C�H�_���6�'�hKg�G#�#���{�'�r�b<�0~����.�e�C[�ժ��P[��`�
���*���N*�P��Pm�-�L$��Qc��w���\��UPf���uV|���!,�X�`�xa s|�mq_��d��0�>����S�O,��"�2'خ(���~�m�������$���l���PM�Ǒ�}��w��*&QV	��fk��E�q�1َ ƙ� N:>p���g�	55��JQ.����k+F4����&a�Q��Z��Bow���|I�\�C�0r0/=�c%7A��r�f}�0o&⬛�'��+��n������3%?Y��>g�h��s��,s�yA��#�=7���|�7Ɔp
�,����xW=8_��Djq:��j � ܬ��DlƣԄ!�<F�_�v��^3%*~� �K�U�(	���
q9\��
��N �R��W�n�����K%�ᳶ�n���b����}�p�H"���ڲ��;��R3R'�ڟ�K�����w$�褈+\�1
���!Q���_�:o���Wۋ�t��Le�l+�E�8s�Z����%'ǝ�r��I#�2zͩ/F�����:C�3&����PW�AX�� F�"����Q7��P���N�4�:c���6VbF�,�\�4 HQ	t��{Ķĳ�u�PH
ŏ_u٦6�>jF��������Z(ˣ`O ���J�	�4b��pP64��.�p��
��<Pq��hf��L�Nǟ�%7�QъF-b�L`.�N���*����Zޡ�A�RT2���\9���[�+�=�O��vم���x�u�4T\���D�Ho)V���z`'��ؖ�H�`�<\�Ǻ4�P�4�u;�+�5�'*򡿇�˓�g� ���ާ��ԕ�PaR� ��:z�ۤ	��J���̒��ۣ״�t+h�[����E����OC-2	���i�s/g�&��B;L�Nd?��8'��,�A��r��e|쫩�Vo�m:c:��-y�j�|ŧ(t��'D�U���
����N%���Ъ�
c�᫐}��
��JPk�WO��Gu4Ոl���P_�7�g�%H��jO����j[/`�l�V��M��2��5��=�����tBq�X�i�qw�{�T_���tL
��x��2p��*�9�*M'�P����R���V=�28���H�r�n�5�W&v�iG(�밲����@�-$��};$�ܓ�hS�8��0)��*�//���;�-R^��ki���?�J+J)d&�]"�h2�R�I�-9<b�Ix��	,�$��]�`�@[��.���[Ob���|䛵�������J8�_	�L�8�!@��2a���ߏ��hD6�X�nM�=�7=��55
���U�B;L��reh�7�w��Y���ߠo�Ɗ����GA�Xig-�=v�HPZ`��T�m7 >{_��}��f2n���x�$��'hRR��<F~�N���kuz�3��+�6"��7�h񔣤*ÿ�О#P"=ؤљE�(_P���t}���e��C!r�F��,aT\}��MC�}Y�}��zu��V�~�Ҷ}��"�-L� �Z3u )��4R��_X5�QU�g����ϟ?��v����m��8E�����k/��B�a	�m��-���Y9n����q�ok���U�,����U+uf��nC@	FV̥�}Bj�D�3��+���v���N�t{@p��Jw3���%kB婦����h�#�y?�&~���ɍyW�x3Q�B��YJ慓'�y	 #.��~�7�:v/l9׼���"����&�|�Z�b'���t���Ba�J��Z��P�v��e\��8�J�Q~}�9[&OJ���%y<�ʾ�F�VIV�w<��OG��8BI*u�f���$�>on<K�so!�_]�!O�x$�Ļo��cX��g��(v
AU��T[���$ϡ{�O/3~�/�=��<fB�l�7�o!?}o�e�%��������B `��$�2O��[j��׬��^R
tC��?���.�1AW��6�Y�-3��w�w��� �[�@<)V���C��!խqe�hB���)�V��W�%�>JݪۼT��#�&�V�#�GT�є��tb�wfyjD�:K0�����̺7��x��:�[ih���[G9��:�L�5�%���]�t��U�/�K�hz[��}�}h���Ge|�>�v����ڇfR���θ?3fS��Ѯߪ ��?x ��t�/V <�A��W!��-:��;�$dli�nH:ZG�	I9P�1(ڣ�	޾��kA]&���?kc!�l6��5Z����[�$����9W���4�e?ӏВ���F��[(���a�Ȅ�}��pP�p�z�K�$5��L�Zב/�qb�z1�	��ڡ�����X�t�1sm&� �Tz�T��[��o{y��Oټ�G��Ë�s�#s~ ���*����}z�����;=��0q%]��%���4�.�ؚ:U�8�7���F޳�  �x����n�n�o4��)�N���m����m��aޚH���)}����1��yŹtz��tr0R�,)���k��AX��u䌑x�Y��F���`=~��L��s�7/bė����C3-t>�%ö��v�y���h����+v��p���z�,p=�a6>��xxB��{�q_�^I��ΜNf-�&��F�!pz)�!VZ�[�Ў�,y�&#tvO��������{����k���d�8v�1ܓ��2��&	#Jbҗ����j��R|�aW�+��.�r/�N�:͡��b�`C�ٌ���kc�:lK�0�Yx�!�11�,9�vP���9�21<V�S�+���zaԇ�	��(�H	�ϋ%E��+�Ee!L��C��ݦ�M0%���2��TE��h����&S*`Bb�-�Tg ]��,���{��S�G�IS"&1N�`!^*��nBCg7�rp�2<k�u���
�P� S8X��wv��H���\��c�b��`bm�0쭑� 8[S��qE*�/H�&
"��9�
F��y�o�1бY#�?a���ڔOw�h���Q���o���\9g�DL\v'L�o,v��4Հj�V�����&��9�i�]��W�e5g�G��_J0�,R�����!=M�7vB��_�A���k��[���Z>87"�^[~(p�"8��G$B��"��q�J<����� Qe�l�+JIQg�ɗ���.E�����v���Ò���͑k�.S�n��9�I�Q
�f�{5�AA�- ��h�#�B;�&L���Id���F��U�� V5 S�p}�V��5�8�TUކ��9��j7X��܊�u��?�,��۔Z��V]�SX�*���Mw�E������V��5"�$sH6,�� ���.�@��#H�A�N��\��P�O+�ORQ'-�?0����"u|
��aA�8zG����w���� ��Z��b���5����eeH r�.�H�,u�Is;�j!�-����4^���P+9��?���J�cpvo
"�íW,�|I���h��C$�IC�m�R���Y��d���ĳ�bG.�X���Z��#�_��n�%�~3"a��^̫�:��8���LE�W?é�Id�!L���{,A���Ebg8�b-������q����W���ƃ^��^�2Md^�Bo�SBf�˴q�*y�{Y n�_�H�&��]ל�?�RTs�&+������:3f��u�� I����vPO_���{�����&���"%�mq��19Ηk�{29��K+�T���O�;5�y[�{�޴J�?;�G�I��G9uw�x,��#Ϡz��$X��ũ�^��9�a�ާ�4r[�W%��m>y|��y|��.}�����#�`���}'Md��ކ�0_đ�:�Z��վԃ�J{��8���.H�w�X�	�K��[9#o�,��w�r�i���S�5~v����AU��h���)�W��1�ҥ�{��tծ�8�4nEM�Q�cg�$Z���v��'k�ǅI�pJh��Z��XkW,1�-��3�:���;E�PHt�V,�%�s;����4�˶�Z�����z��w�r����P=�*�'�(�[sG��_o�޶+6�V2(���	7����Y�-޻s�΃�h���5l�&w�>��A�cұ8�f��z:���,F �V}_C��y�/�v6{k{F��w���0;[�6�<�t�T(лz�T�c\�m�U2h�#��j�yZy�N�����J.N���zt#>�� YBAX Y!ʾndn��b���Qhz�.����뜘L�EOƴ�I�8G~4P�to&���j�`��(b�Q��[|b��@4��D�?L:��pUk�B���%O�ɸ���0�ȿ)�k��жgI��xG]Ɨ�l�dV�����@�jŬ��> �$��������L V��\zQ���	�w�?.��נo��+LM�1sǃ.��� �k\��̫M��:O�	\ٱ���ncuV�2uo�Ms���@U��h���A��)yj"�aк~�v|�>�p�pc'�%��zT�P.�3�V�̬['�RI8���?�}�m& ���$�0W�%k"�F�ߊ5�ʁ�`�N��~�3
dyqM��k��c�z�}���nJ��f;Qܺf1̏�P	�`o����
9�H��q@׺R�5��&�󢊩>68&ܛT�^wU,	�* �%;7k��p� ͎f/Ļ��n��(���������v�G�*/�+�+.������
���>g	���TA��x�?��s����r�h4ZM�����-ry��p� �9{���H�v�U��4�Äb{Je^�l�b�C��	��� �c���qTmߐ��f߫�(S��e�0oZ2q��Ҙ�+��`�H{�V��Kx\�3{3rT ��sϐu wG����ؼ1�S�=�@���sw�7=�]��2��ylB}�K(��k�*GN�|�>�)�����8���I{M2�k�e�M5���(�L1.���Ǟ�����|]᭕�v��]}n�����<9NU�r*]`\���G��r6F��t<��@�gW�>H��ޝ����2L{J�M����(��jN�m{*p4��1@`��w�������\�3.�|�+��P�D�$�j���kR~,�v^%8�M�[�4I�of*ٕ%�m]���;�L�^e�\�T��:�j���S��%B�e^�� �B'=�ɫ7����\���x����,A�aQ��Z8��%��G��ù��M��72�H�r��`в�I'��%��fk�w���x�C!� �=����l��D�d�a�jW���Q�b�SpM7z�M�9<9_h��SUͣ������$U.�FT�b�O�y��5+�4��t�*���q����g������^Vaf�7�������/`��D��투����D�/5�YW�q������W��`J���4��]A�3e!�c5L���F#��]��MXe�y�~��qa��O�aE�#g%KE�������.�iu��>�����z��h"n4�ܳ@8 X8���]J.��
X���x���D��@<�U>�d�릠U�XH�?���n�$f��7�=w�:�G�|�ȩ
�CNT��p&��oI�3��d�)�4��2ho���7
p�oozɞ��3!��)�h�Rf�
�ks �R%��`�rpsP6 g}P�^򖨽����(�Lq?���>f���
Q�����Y����mS��Ծ��R�E����T�r$�o�
�6v�z���%
߅����H�^Zo�c�h۱y���3��LL�tX ��:Վg������A�;"a��l	���{-����>��9%�̑��t
YE�����A�����`�ؗU� X��{�t��Ck;�i�Bp^����p�
�Pl{/����f�f��G�;ӧ�K$�D�#N�ԍ���!(�b�G���VE�äf>��wdPn�����@�'\��$�X�� �Y�Q�M.��uU��v)�"tc6/E��)5� �q�Iaֲ-���.�c���l���E�5�-<�h\�Zfj;m;������EʎC�l
x�z�����t^����*oxJ���sR�B��a�1���[�$�����Ok��q�Xv���G�N�5�瓐��n1i��/8���F���$�R ���*��Kd��"~�~�dxXk�F��Ʌ������o擫�H�Y���_��Ŵ��矊REE�@	���b�[ܙ�t�����h���84��G�	�c���_F�}��l��
ҫ�sr���^�LI+�� S�]����#"�d3��h�◳ԍ�Q㷛�,T��e���N�����+�sO_�P5.�9�v�s��J����Is��o�A���v��Ba�_*�v��Ҧ9�㝀�%l�&2����,�����;#o�X�*��!�Ū�f?��w������3���cPH�4�37�.�R�בkWV��O��
�=fbn�F�ţH��l1��n���_��n�њ2$uf��O7.�i/�I8Yx��-w����MII�ᾙ5%�pYg�uC�rY����U:2�ٗxV����N����15_����sw���%���>�_�)/�h�,A�˜�B*������J��cq���Z�+�� A&��SI��(��<���Zc�3�5�:��r��6v��i����LVo@��֗uKI8l��3���K�6��*�X�LOv�'-��˓CD�+C����2�}.�cJ�++lnm��%C2�5@ߝ0"`�[F��9�C�-������p��<>QHK����b	:�v�H���dzхM~�V�-ћ��O�c[�;�	�����j�t�:��$>�����3N��������wO�������"D2H�J�������bL��O��=��^x=��"�\�l�VO>J�:y�jV����g�JHi�M�~��LY*�	uMH�T�1�I+l�.�A�N��/yCյ���vw�@ʴ��HE8��?+lγ6:�&/�Qr�7�cA6�
r`��;���v?s�5��@0�n�Q-��Saby�w��m�'��o�/��vbj���L2g�?�[TY����
�BQ�a0��z�$끆HeG��*�3�~h��Q�y�K/~���G�ժ��*�2�����.���8p7ZeJ��?����R��j'�çϋ#b��(<��+X�KI�c`%�;x�:j�:QH��	/p�1���%
S�鑆WEjC��.��H��{�)#���pP�5WW�*�45�[˹�>6dQ�^0��fqO]Be�t��ِ[���|�3���dK�߈�Y�ۇ�����My��ڥ�⮮򁼺�F6�����]%����{֑��J�b�d����ڄ(�U&
ڋ 
�V~��.�{�%#���$�H �U�j��/�4/����*X,�P��K�9	;|!9G�d;��I��9�ֆu�1N�F�\���4���&R��C�2����ߋ�]��}r��\"5.7��\N�ǥ�p#��]\~}s=� [�!6�m�� j<��#8K�]U�EV��X�dt�g��|�g�h;R��w�V�9w{G�h�l��W����^׊�Ʀ��[ԚX�E����Y�Z����~i��|ݫF��'���)���ڸ�m���\*wq�*)�q�gpk�
��a��+�oRn%D-洠'ع�^�5�9؜�c�׿߲�j7U�I�w�lD\�9�`��	#̤�OõvO5���sF�Wf�Pu�؅Q��K�?����5_�.ç&g�
udښr�����hj5ֲt����o+���DD=�RZT�"�#m�)�qܮ�_�+��� !f� =1'�ݣ
zgqv&�˹�*�n�4A}',Q�:�