��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{T#�5~O%�0���tko�^P�fzp���d�MK�)�R,0��B�&9�ҮV�f5�݂R	4�D����} ���D�����o+�h͍t�urQQSy�/�9s}cp� �N���T���H7^��7:_ݻ�ƶC��1B��œDk�*;�*{ozQ��倻Fu�s;2�o��0#���A�ی���9V�h'i��|%�dZq�tW�ViI�P�Tٵm�K�E���~d�'�z�C�0��,
JV��m\4���x&e���vP�e� ��1��e�^)�A�<e;�O���H��k�Z�y<T��@,X��-��Bb�^�f�5b��{�1s����f��BE'��1��l�++�i�Å2ƕ���}#+�҆�l��+����J%�$`f��2]�oQ�q������0�SQ~D	9��?)�<#:6�2:�K��'��u�|Ӈ�Ua0�̾;�d8cB�-������8G#�0�����G�7r�@h�{>�6k�+͹g�U�4�� �K�bC��>9�'z�Ws�Z��-�������_j��]�Z�fT�5����e�xo����Mہ/����B"V�7MZ"@C.�1�f�*km��s����Я������ku��/8��f����]��غ�]�O�Š�۳%����A7([��.	�} W�A����� }�+Ȃ�#�/L�4�O;�y����+��ͳ=�8��q^�$����O�Z92�B�O�ͯg��>�p�������n�j4��+;��e1z���A53�5 ���;�Po���e��w�4������ M�������=e|��h�	����\�B���-��9o�}� 9Y~�29�t�f�Hr3�� ���x|3�uO0iǴ��"�{�뺔#A�l�G?�GV�j���A����}ɺ�]��"�r��Ӽ] �&&��
dj�d���@h��	��đ�p}��;���f�'�hdp���*B2LӃ�Ъ �%������^�D����8�^?J�БImF��eB�Pf0�|�;7��J#��ȡDB���m,Lܕ'�J5�p8�%NLFQ�U�P���m;?}�j 6�B�9Gԋa���T^��m9%�PA$O~����J��J�'q���J;��'��A:;�j�|L����!�s�t2�.��UT���ʆ�� �V���5��B�L�]Qg����R���1��U�;�O�r'*d ������\.PO�֑,���F4�%��>� �p�|��|������ێ |�%�,i�bS�tL�II+ׇ�4C���<I24����KM���[U0<$�T��1ƍ��R�U����&�b�@S��|���(��{
���޷HƯR�A��G�#����{�$��z��ۥ��DPTU��q�O��gR�bO� Z�
h��F+��iޅ��(o"_%��'k
��&�v��z���\0��׬�l���:���خ��iq�-?�Q��mh�ͮH���+����=<�g��@�Ѯ�{�դd=U���Ȁ*�J#7���;y{�9i��Sy?5,��(�32t�ŧ���Y��g�úo�	��z�2�\�q�@(�JJ��>Z�.m�i�+v�����\t*L��[I%Ju��t�]��j�iYx��8;Vw��p�?��$��M��y���E2x��HH���uj��j����3�+4�[�"O8���V���B�1ĸ���g�&�P�k��Ѵ�@��,�z�z]z�ta�?۠"��{�+���(�/�Y_���ȶ�+�u&c��}���g+��H�nN �XؼPy9#�q�B
��W-1C���iN9�ܭ����S�Q5Y�������P��i�sw�-���*�a����:��f��jL�gAf\��_rjec�a��57�٫!@�Ln(�151{�_��h�a^C�]�`���o0���t�����^�n���5����Y��x�x���H���y��p��yQfݹچQ�!��)�E���H|�Q��,|���MX�(��n���G���vw���5#'��0J�,ç�W�u7�j�(��e�~W�ƾ����8�/��OSQ���|X_�P�.���Vj�g��RT�s��1|�8r/M
ep�o(v<�ӱ!�s�(NG���D��kڴ/@���	��9��($N��������d+Jh�����2�9M�>Laś�Z	\An'hv����YDb+,=������U+]l��p�->�����(&�I�&q���FoVN	��b&оo"�wto���r:���Ru�̰ۭ7:*��(�#���Ǯ$�އ��a�kz/�^L�g[ �p*G��x)������׳��j�%,�.���.��
B�����:��Uɨ���z�u!ZsW=W��|!��Gf�=��@5�1���ǥ���f�i�Xq!]���g�"�W��cc��ĿR��� �ē�87SĈ~l�<����=�kB �v?����u��Z�;�WJ}����Rp����QN$����B^�:1��;䧧[xx�4,q�$��|�A�osQ���������E!I�(-�{����)]�4�4�Í:ֳ568@H<~W�h7��"�"WM�����4���	$V�Z
-׽�Q�P�P���^�Xa�<���"W/�/�I������K�*n^���vV�ϻ���@�d�fHY:x�t̓L�/g*O��5�^�Gw�>�5�bD�*���w�s�o��x"�W�PCj}xi��,��=