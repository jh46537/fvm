��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�k*b���f^��g�{uZ�����DJl��NCVs��T�]��"��u��\��UQA
1�TSJ��g���ߵ,Q���b��������W�"���8���tP?����ܮ�=�EJI���M�*���C�_��v7TR�d���!���WW<��m&CI�2G�>f�};/X��[�������s��Z���Edݹ��y�� �'a���}2=�4��:T	�-���Pr�d8�
�
���ؔ0;_*���GOj�ՖƓ�&���d�kz{=1�D`�˨��%G�#-J�Wq����U=����Rn��o<Q��r�O͓�T:�C�;��N	4(�寀$ca��d�z���;x��E6�4(4�#H������؊ n���:�����Ah�w�p��H�i'�N�K�xb�_�L�R�3���:�Vj��R�7g�`���__q�궏�Q��m��2x ��V�1����^<�VEavo5
�ޔp`��u�qXM�"���:6��8q�XW��5�G��h�V���P}8r��;-l�{8��A/�:�g!����
+�
"l//�O
R��G,�|v�ؽiڟ+�}	c$�.l��{�!ث���x��y�U�d���]�N�Ld[���g�y�kR���%&j^~=�^��NZ� �p��s���h�,2u�����rdYY��
�Y�0�=<�/)��pup#��
��gS
�Z=P� 	Lq�q����&WrE�c�0c������Ī6��1�O����0�+�S�k&$��|���l�#Ƭ�m5�D��W��U�㴘�
-����>o#C_.<*y��0��c�nqH�5�h�(�,��|S�p��s[��νQ�Δ롘����H�U` ��t���d��_(���җ��O�,q�2�~[�ӗP��C>f�	�Q?�8�Ӧ�(����s��e���zk=��ҔF�����y��$���т�H*A�fxo#̃"�# W]��_�/1��?�e�H�a���}-�®��۶6x?�'�CpP�V�ŬLm�֪f�]������[��[��*]��.�u/|+�d�ü����!��k8$!�?�vx"R��U�ZC��q~A����k��	J�>\5�c����'L��^F�Yv� WjٳC�Pd�Tңq��>��܂��-��4`}V�Dv2��)�
�n���B�"����Ϫ���kF�ܒ��S��~U�j�O-b�r�1힙;Қ'��{��.5�x����8�*'���=���է�d��6}5zmSG��!�^t��63$z��Ʌ(��Mù$�^Q�(�>�N;;2�*������l�b��{"|q��L��ʔ�1�
!�_��®zc�v��/�[vn�3h�˪YO�Y��`W_�@���%��I�P��3��na���&rb�y�@��p"M�k2���}c:�Q�+),�3Q���aU�Ҟ�@8b����am3��+�d�7QQ�=��"��i, �� lEJ����G�ijӒ��c�!"�G�,�ʘ�V��th�̚�Q'Na|��-}v���8<�%��,�\�9sǶ�p<�\Ku��Mb>�4�ߺ��cz���=�Ї67�X��l���9���]����f/��pF��t�
,����ƀ����T\�DV�3�@A��Qb�(y;!���=���e%RZVuN�.��������7g�^g�T:���ܝIan���"��_�R�?��2�2�y͖���E��>��{��tEڏs�\�Ry�ww�Xz�����p�&��Y0riy�چ����$�B4����gK+����W��5%Na;�J��Yv6�<�$fCۭ��qC�4Ҳ/S�S�r��6�z��- ȃ�?�4�(\@��&��3Opş	_�K�z��8��}���2� z~SH8-��;M*�0dުAQ��̐'��!�>�]_�.�v�+I$ �=�:V"x��}��w}M��+��$Y�C,�y��안�
�{��$UuҔx��!<؉����$��n!���jM�����OS�����<�+Z�h�c�ߕ���ܨ�2�ᩦV�[�Xt̋�������}�6穰�:�J�/����U*z�?��MC�xH�����EŤ�/��GpT�9����ޔ��Z�{��-�74�ɵ�.P��"���r�ؽ�ZBU���5�ܙ7��Ǉس�߯�@H�FA��\���E?��?4-��LF����  #r��GM�ӊy�lu��#�3Jʄ�2dr������ ���tܿ�7��W3xyme�E���N���T$����.yJ�e�͟_�E8�+�E�R��ڶ��vfoE?"������,���ho��/No�@�I@�C춆�}�6��߶����,�ݒ2p�ML�D���5~�O^`�	����r1%fb�9�ҴK��}�K��^D:�ڌqK�p(E�9��0�êRw�o��;�����(�J;�+�~M��pQI4�w�+j.�q�|�eP�53v��^�&��C�\)�e�71���1)s�/�ޮɸ|�> �܀�t�@����q�w���F��9��(�J�4�y�w��`��U�<��V�e��V;�B�;���}���g�./�@<v�K?}����5[g4�����-��ZJ2Pq䷿�>=3�3�nJ���}r�iz����Qrj/����%~oH���6�D(�p�x�(@�YW��N��Is��`lkbi-=�ܧ���\�V��mF��T���~@�Y������Fm��'x�j�%�D�\�����Y�������f��Z���y)���"�]���v�7���z1���q���2UC4��*��Wq�?�����u��_��ϗ:ӕ�y|M�֩�P�7�,(�)���>�	���Hy��HN52��i�m���T�Np�u��O�ݟ#i�����;���q��L��L����׺h�ū�Zf��~u~Ȉ�>zF>	��JZ:'d[�8����a�~���k@P'�@|��9kP*Rc]�اj ���x�u��N*�E�j���� 7.˯63/��N(�F�l��Bƴ��kq�G��
�9�����~��A�<�'�Y���ڰ��1�*LY�O+���֋�����2��r�G(�1AJl���3��ɗ���&!̯۩"Ÿ�wO�Q'I����:�E1���0R- n5��:�+�E�=��͜�5�0�3�*e�&�(ȹ��J��!�a%�|���
�ȫ7�w���f����@s�Jc��D��u�J`�������lek�J["��')�y�Xt�T�ޮY��5������sb�ݗ�\�7�}4� m�	����Gs�3��>x����3�(��9�"�y5ea����5��<ߊ#]���1��ޔ`85(���,sHT9�潐]�x�e�<��D��1Q�k����iO�T������6�$� 7u�a��M-ǟ�_i^�v���䃨nN����)�縉f��҅��`�x�V£��_�e�)SL�kk�)	��U�CA���-1:�j�JI^�8E
Q�m��h���]&��!�]2�ï�ʙ���yu��0��$��IӃ�0����? 4����z��?�6�|�c\;.e�L=�$T���yeo\�L!� 
��X�BMBO��q���2�i��&������ތz�%��\���/H�52����gw�sK��Ͼ90�0�>Pv���#�*�����q����C��� +�P�n�������Ʌ��8��IoL򲷜��Hj˯-�iS��G0�5�K�[BPRp0}E�E��[aƶ��DD�z�!&��3�BR�@ތ!�m͢q����!�܈*!^�"����`�+�T>#i�*�d�V���ˏ���R�2�����/Bt�;����6����=L��۠)fa)�_3�|�e4�g=�y�;��K�kG���2�B�����ӎ�Z���` lw��wI�M}��<�f1�Y=��-���GQ�b��rZu�g����Z:��X�
e�l��|��&��uH��"#�0k��,�ߤQ֜�ͮ��8^���0J�i�f�p.�\v����w�䱣"�F���d�5��-sp�{~z��3zp|	ĻR� ���34����R]C��Y��L(�Bi:"(H�{��u��Zo�@�Gġ�\Ä鐾$̥�l�5�wd��c�d@�5�Kg�-����T7,;�)�.���>�]�X��ʌ���j�sK���qJhP�ؗ����5xQ���j�I:�|=1��r�omE�[QL���\}Ld/���7�j�6`Mn��d�Wq��u��>s�����o������7��Z|�?�t�0ۊ�A�7��S�K<�;��~�PEB�0⳼�<Y�U�����_�喍��B�۹�)}JӍ�XKt7����B]���#E�Ύ$�J����6�0뿃Ĵ���R�y֭�Q�5;�������J.L�-Q�F�>5!��ĢK��Çh��H��Q��!=�y��J	dmLNer���)�/D�Se0���/Q�<����a�k4��ҖՀxv�I�؍�R�{5��_3RA�5G�������%� �@d��R���%��g�̗8-��]|�:�0�����|��G$�1������Ë.��'	9J�֢o&�#Z�6����Rv�bj_����sM�8YQ�R�H����_G���q�\m6z���R��"����}H����ާK��׊����{Ȭ�Vz���%�#a��')t|Gv1�7�N�C��D�-¸���&���4�s���>�oM�����F({��Y�ER�+0��煬{-H'ԵC˂a�Eˢ�:>"�ݞ�B6��R�rU\|��_�]obv��g���]���Jp���ft᧶]�ϑ�+^��9&����S*<P������%�9�{�m����^��%��ұą5h<�TH�+>��k'9�O�4�\�]��N��[�n�O��q���?`�tQ�En;��y�-�V��aENy�)�L8O�@�v(ȭ˩6�g������`�W���I�$^�ʿ�ZI��(�
*v�v/Z0~��^$����dx*�F����X�u0E�=EX������Qf�J��E�l�RΨ�+��/��sO̓�x�]L� �@�����2�O>�r\4d0d�L4f�|T6���^b�������N� �i�i7��ه��������LHK �һ;;D�B�i�u�C7�N���^Uaɮ~�˃�{+��N�H���:���!aɕk�6XB��ϸ�e[aG���iNȑ�	�삯z�u"m��t��ׯ�&S�[�qQ�j-��>��	�V����1�L��G�J�ףZ�Ije�3P����`Ҡ��"P��>�
C<.sq���D&94g?^Ȉ��v&
M��u�E��X�T����TX2���)Q�[�2aA�`W*̏���0/����6�T��(p!�U��?�z{-�--���|(ɛ�,�;����ٚT��nl\@�1�N>q	&��k����{�J&T����շ�Y%�N�KB{d5��Nb�lĤB���"��r��&�TP-��!i��V*ɝ��b������9���r섇�I�d\�*��J��d���3� �aPb�PZ7q�=�[�H�0��gC��Ӧr$�+�`�#$A�lCK�7s�c���ͨ�f+H�y��6c�lt�-m߉P�'XkP�S!��u�o�9�Ƌ~!a����;�F���E��a�ŷ�R_�~�Ϋ
9�Es%����x~���տTf�Vu��,�>�u;8r�.�_�q�h�5�Gi����.t��=�9�׃�,S\�2��z�i» ��һ|�>2We2�xU�j�����̄<�v@�92=k�Ed�c#�Rܽ�#�+Z,�~1q�$,��Iq�O2)j~g����4���]:Jf�+�p��-��YF�+s��k����Y�m���K���B(� ��[m��	f��D��������vVf�"'+���ٟi�j<��l�3_٢,o�xqi�ʠ|F�^C�L�4?��O�n�	��*��ګs�ׂ���D]I��>yE��/��k���z�(1Ϥ���q.�!ڇ�4<
t�뾡q��l�Dym�$�y0I<�%�t�0�k��f�R������_�N�8�γqu�r4�\���˶�HM^j��<��[<P��V�N�a����=�?��h
��pR��I�;=S����͗Q��$q�Y%�����t�-/�:�T�C��T��L����̵h�r��LAiKe	�l \����N5O�`=b��0V�LGTc�P��\p� Vm�C��x���q����^���G�� t�*���
�2\{��!���C��F;T�#�l��N�#��?x��2�'u��:��k��3\d87����pJ��Z�^����
��R�'��b���e|$d f@�)�~����I�,$�vA�3�̑��Q�����Х�p�.�~��O�?����/���K��Z�K�_���.F8 ]��y���s��R��e�Ę�㽲jy���b�GY��#��m�á�-u�ގ;ٙ�֐/�Ăk��xn�F~�� }]��'Zn�9�l�6�k��~�[�3HQq���9����[;ot��H؃���(����V�/q�`9i��C,/
�gd���M��C0�E�W�JR0E�zQ�=�����d����[rW�N�1'�"������>1X�g}G��i�O��7��Y�q �jy�M����$_�`ln�?�z�`�!�FcTX��X��?���K[״_����%����`����q�z���rg�ƽ�M*3����i;y��֍�~[<x�r�f.%(Kg埞N�?yQ�%��:{һ6�N]�Z���b�h����>#��!��D���6�Ʀ�ݡF́,b�0�<����!�����#��9�Y��!K��L��"�S�yՄȲ*Ø��Y߂W�.M�!Ə+Uv���D�fC���L��G��3�ii�����V@LX�u�Xm.�*��Ӿ�@�B��W=��8�[�ɇ1��-��(��n߇�o}<q�o��0')#��eT�}�N�v�Ε0��fof��e��O�@�!� �Ro?�!����hI�d��8{A��w��-�XAa&���Q�)��Pux�� ����~�x=�x��Q������%�9�Y��MI ��!B@����dy��i�6��n�k�J�c���Fb�ǽł(C�ڝ�k��X��$�a�,�-���H����yԫ� GSB�F���.;����%��y��ϟ>�ȀU�~��@XW�L̓�m�]ML.Z1���m�T �?�JZ!� �ẙܚ�d0���=w�����j��衷}N�؅+@aV�����J��J����G�nrV3�W�,%0�y��X�۶��W�p=��^�r��F���ͯ���k�?�5�#�
j�G(sckf����;�৚�~_���P|�G=�q���F�NLCS[�nb� $�i4����Q�n�ӛ�~��] B����S1l�zH�+�/����[؄��	'h�巻�����$A�ayx��Y��n��_� F\5��p/|Mw��,�OB���l���ޥ�'��N9K<'�Mu�����E/�A߼_����ǎ
�\8W�F��y���co0+�:W�K_�>�I��l���&ph��e��'U,Y/�(���:�N��Z�i�<Д�F�j#�鈺�gM�G#�4^�^aĴv;@X��& �Q2��i�q����ZcI|�l�O:Xy�.�;Oqn����Q���R�=�C����ا�1�e�X� �����*�s��:y-�FB��\�7��C>K�qix��y��M�2?� mح�9&�8��h�7�Y�׀Y��X,��7��Q'��%v��}v�rC�۠t����Er��g�K��L��J�V9�cĞp��/�3w`���G�(it'y���H�c7���� ���٣�{
�'��r�;� ��M�
H����"N?>U�*�����^]3��OE���ԃs	��7G-g����\q�W� �G���8ڐ�p��a}�	�]�b���7�a�8��$ݦ�{�Ũ.߳#�˞Zٿ��xݍ���x��	���;�3Inn���2(f�0�9^'��a���r��n���Ě�m)�>��{�b��t]O�5Ҭ3��jF@��Ⱦ`���S%w��Q�q_��F�ݨ+�q��Kf�a8m�33���ӑj ��xՙD��X�)O� �kؖ��oC��Ġd��,s񠷩�㞇ʹ��ě�ih~'@�و����s�����:3=.��l�� 
㤚t����۹W��2	7t��>��S�E��;�r_{��[#Rl���@/�KN�Wx,C�7�<��X�:X\��0v��H���q�R4Ep�H,w�0���ʍ _8�����.9|�44.�
2*��B��m�J�,R��r���
ևmΒ�g��˒�Fo:��f� �2�/Y�ߕ����6���ɽ�	*m�+}�hq3 H�I��+�y�!Ir��~g�����S|�Kۧ����E�j��?�,	�Ǻ=�Y��`(��x����y�],��������ъ����[�{�;%�PM�5��ݭ��ԥz_��x��Ӷ�� i�̂�e ��7�f��R�C�(�����j���&�r�5��=t��
�3�� X�2&������Iv��g2~��'��9�k��֥���n(���E�+W߻����)��6�T�)&����qrk
3�G#���w|[t?\%�d�6K=0��?n��9�'cӱ-ވ��sj�1���ͼ��s��h�s<�;�P$1ɓ��Q��Q�1ڥ����B�x�yF�g��:��0���]u7'�R ?'j$4�:�&a]Y���
�uГ�j$rO{���W���L���_�^�d��K:V�����@�1���۷(��d��/|��7�;MIj!:_�^���Z~���(�ڦD�Ge�Hg�駮^\��"�j�<�bq�K�>N�"�ٔ&a��nW�a+:7}b���/���Ŵ�x9r �<�ß^,�� lϮ�h����%�4��4��zL�b��M�G���ޙ�ex��	�ƽ;�b��f��9��4\ .\��j�h=�Lm��� 5!\`^ ,��Д#`ر�QZR��n�+��[��sR� �o�}��r�� ��Ө��mJx{�<�v�q�*3	K��|Sh?:�:!A%L�}q�� Mc�H���%�	��0!��v��v�T�@A
��*J�K���3�f@*lA�3}�Zk���lٌ�)֞�"�E4v�N�S.Wog�<��&�Z�D�]Z�'3TD;G�G�"O�*�<9�p6�/�y�*O�+���n&�R��5Z�E�����9�K"VU$�F�v.k�վf����ؼ��d�4.s%8�%�{y�4��8Q�,W�o�ɶw��H�xc��P*��y\]��~���:���{��[�с�ߟ" ���L�v���]]Tǘ��xx��̄�>�����E?�v5���U���dTA�&>>�mW�Ę��	ء�?���il��)S���~��>��
)"K-��������'��R�189L���y��[��tu/aN�X^��J[�'!,�>HN�wʂ(ӎ{���- pȈ%w�8p�zs���+���Vj���{[���A��*`1�I�9���F�����2}���~�<�]R�_���\E��/��~���Xt�#���?9��7K7d���#�o��|���!ދ��P�r�P>�{_(��F�n��:[,!Y�{���������9%�7м���%tJI��5�f%p��b&���&m�y�"v�-�tSdl*x��T�󗁢���	v��oYy�m�j�1�Vo�S��be�uڋpE� ��+e���]'�[`=]�_�7��;�������HGY�`�s�tʧ�/�n
`���eƁ|���q���(�}30�O�V��vo�<{��u��J�!9bFd˷������3.a"��^���]!�����;��0���
=�������mN�Y�$��kk�S�֧�X�n�Pjީ�J�}���"�B+��N2�O���Af:�~Y��X$�(�]'S�C�N�댑7���'ZƛM��SXA�Y�)�� �x�N%_�9V���n�%zȳa��q)����}�*Օ����] K_a�8:/�����o�3zE��h�{1 ��0<��,IA~�?�jl��G���-�腊���+NS����m��P�T����=%m�o<�Q��JV�߉������dl�D��il�Z�	Y�����K�_(�+__�/��nF�l�Zo- ����k��4y����\D#�fg��F��K	O�ʉ)G[����q^���͠Bo�k���5�A����Cv������Y�O�[���3���|V��y���XR�̦.�7,��K��6�P+j��ƛӔY
\H����t��p��.;�*�j9���4c��q/���?����s��� �m�,�� �F�2�����45q�s!��>�i"�,�]����*��_H؛'�#�v*x�m��X=�
�UѺD�������*��X�k��p�4��)Aa\ͳ�>xX��e���2@u�����gV���]��x�i���vm�_σ5�	i#�n�=1�O���-R=�o�,�b�b�� ��?�^ �.��B�#��F	��7b���Fi5�'r[��X���G���<k�����k�#G�Ӊ�p�/�\w6�s��O�or
����AfO�d�#6��#Z�gmov���	?R?����ܾax��h��#:m� ��m��(�r�%�rO����E�nb�@aR���4�o���Z�e���3����pG[#����k����)�}t��蓞�7ï�T�BI��G��� ��8n���8�;蜐1~���9�pVkf;M��.h32��cZ��gɦ�e���d3�ak�L[Ső�1B�N���jwx��Cݭ��dl�ąJ���[����͌gv(��	�$��/�y{NǨ��� G����O�فv�Z,�c>����cԜS���#�D�ɯb�f.V(�>��,r�;���$�2���{��bu��������������|�����<��n

�'�(E0x�N- \�p����G� �T��&�`7ϕ0E%{t���v�'�^6��Wڮ���D"7��Os%�	�]��&;�6g;Xrg��'���#춤�>��	_�9Rl	-�D�