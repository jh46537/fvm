��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm����질�95J{۠�_74~�*���i�&��/jx���������ޛ���WBYW���'��R��OL����>�]�
Z��]�/qۮA���4_K�>n���t�f8 =�<Uc7�/��XS��y\r)�������g��)��R���qhho�M�{0�sC���TV!�[�������K��縼>�����OU/�Y�i���托�����bZ�S��r����to���i]8�El87���-=jH��r�Ɛh'���k^�]��[R����+����!��H�6/xq��|��V|��ɚp�1[�<��8�:Qb>h���ȟ�%������j�� ���:�����M�Di(�0{%��so���iW-cO��E�U@�)���H���f�נ��B�Yݘ���U%�W9����\��e�h}p�M��U�s�$�h�]���m��\����ѿ��n{�6ޙ����m�6�9���V���g�c���V@m�7�ٗ��Fk�p��(���'גt$:����}���w��T]'7���-�.��jv���+nG+�H/��᭽���*& 5&���C�|����E���ZF���$��?4*NQ�\�4q�pi�6%�=�qU^wYT���Tf3S���fჂ�]�a�|�y��yպ���h'@�e�v6+W��F�C��}��m�ʉe`��j��԰�c!��~,���-/�ɯ��ô8CI�їm�S�r�X1ʲ�"��f2�1��	�@�U_(z��P�M���N(O��/����\Y��pӋ=2oG��lzNC%��l���۩Y���fD\2�cdB���/�N��g�ִ���i�1��d(g��1Z�xӸb^�ε ��� [��hǮ��Yz=$��!V�����^�//_({�W�5ôHYmUb�m}�3�&��37�;Be�q&�����>
N{u�O�$��/���(����i��\dp��5e�6������$�j�v��W3h��Y���`'z+��}���f���+	���ſf����V��cYsMYW	O9���;�K��|�Һ��:<�	T�$���u�z�\�R�GC�(`�r�ܺ�H\E=B0CH���{ȱc�9�g����" %�ׅ3�ޯ��
�?��U�{�Ꙭd�����4��I�{�LqJC��/�����-�O�d���}���d�&a��e9{�P�s���q� n����;2=����ε���,�7�v�=
�Dw�\��#Y*���_Vv[u`��.�����l���ʋ_/�F�3�MT��,��L1P��_q'�����@X&�>0�FٳJ�?���PV�xb6R�[���W�鋓��ʈ���s�2F)e(�;�b��ɢ�{�zM�誁S��g����E���r�i{�c�Z*�ڮ��l��B���a���*�˓����K��!�k5�c�?���U���J y��Oh��hf2{K�*`T�jr�ʙ���W���"�S>�kZп�h�״K�rj�Ɔ�Q7�,�.�0���"n�׈<�2g���l��բ&���W��Kx��T��K��?N�b����#kW/HP�!��F�r5w��0�gu6� ���k��39���YU�mT�E� �W��eހ��F ܽ_v��b6�[����ٰ�%�)��r
���Kԅ��!9�0�i�������\��P"V��B;�_A v�A�h����o�yARya�1:�p.�]�� |�9o)�9�+�c�{�v� ��25Ҫa����M�&9���s�������:�b��bV��Ԗ ���fS��o0jR�ҫ�	G�������Ȳ�J�	�B��_����)e6��д>)A+<>�d�Wnc*�w~(�[��IӴ��돇\U�FV[	ϕ	�4��4�,[sr�Ă ��x�9\���Y@FDL�>��
���5vi@,ˠt�*��r'���h�ǹ�<}��E]x��╠K�*L4���\�6_Zl[-��=���;��n�wI��]���E��G�D�[����Fl�=�Gy�
�6����$q�i|O<�I�j��O�&�R���pύ�s�2^O�wN���3K&��[��ܢ�Z����h��	�c�ȵ1�P_�s����a��eC��3XU0`[�m�J�������!�պQD���{|�S��#�:���KH�"���XFV�́V)��9�)�#�x�/m���1˨�%��*�K�'���$���
���d!�e V`�)���8VY�zYK��ym�����{���k��b��h�nx�RR���H���}�����.׈zw6�e=�ћ�ģ��Q/�f[�R�J�:���DM�K����L& u�5�y`h�-�3�5a�I&�
��Q��bM��Ihj�@�M�<����Uݶ/��(�u�:��v��;�Ms7λ4�����Jn���YL	�Hc�,�S�@D5k��i =�E&zX@��j�n\�R� F���+�Y���/�uI��X-m9PB�ϝ.������e��^�?Dhz��P�e�������YH7(cRp�v
m�]�0ћ��	?	�4��/��Rhn���T�DT��<{W.m��9I�8�L{�<�:�-���o,�-1 "h�~��t+>9�Ot�;�M24��mm?�7����u�K�����D:�_ �T�����'>�� H�z���Ъ#\d� ���Pt�1���D�1�7��ixЪ�>��:;�a�����3:�Wj�MnK�M�C8J�5�4􂅯��%����϶t�Y�+s�o��࿭[�H�ůy�)@B����|�\�u	�ՠ�<|H|,��ý���qg.��<��H��0i�\�]�xW��n2�O�FW'���+O��$g{9R��v��k�O�V[�C��ۄpRα��o�`�s��Z�m��v���q�������,�=�*�T�e �8NN�V�iT���$��^=�^�ځbͳV��J_ V���#�ZH����3�H�
l���`�Ț��R�?�s��Ʈ+@�̸dR;D����=�w|(ŭ�ù%gk1e�=�5�)�(��Yy#�^�\�#��G��H�v�c�̔�s�w������7z��e���)bX>'u�����xb�,�ji��8n�]��۩�V z��fG���L���7��C�|�N\�$	v��W�%�B�+)TJ��#q��n �D��~��0�+����F�L9�s��Q��
�R���S��Hz!щH3��T������g�Lf�}��"lz��b!��ԯ�?��8R���*���@s?�}v�3�vW)iAJ, edǑ�)P6���Z��{!���Cs3��b��3�)I`�K�˄3�k]���̥x+ւ^�������j�Dޘݙ����1�L?�O�Hjq>�eD��/S�6Hυϣ���Ŗ��M���y6ը(.T\r�0��qp�F	k�ϸ,!>ԙ.r���g�K>ԝ$�a�S7�YD1ph2�Au�<�<�W��&�n5a�:�� �
A��v>��Uz�6l��0-��C����cָ�D�Mb#�qP�)J����r��;��}�<�j����l}��	q���q�8���=ӑ�����VeKM��w���y9q��8t1���&��5kL��N�sPHI����rw�,�$o���4L <�e�c�)5_�0;+I%�!Op%)"h���F���6i��t���1��R9��˕AG-:�.����]��)��a ˃qL%�P [�|�hE�Z��(s �iX�^.�q��;��E�G��Zɭ?�]��.Ѱ���,]��������or)5_!Z���)�e���f� ��Z�j���<{�qޮ�Ԯ�C�gP�d\:��P;��.^
��O�t��"��1���f�||$�?vƽ�s�[�/��,wi������M��4������.уy��T�ė������1>��֛x����H>���\x_�H'D�����F����������ǐۜ���m����f�\P�?�~/�5��ӒO��ۯ��3t� ��k�M,م�KX�C���\Z[�m�K M��?�����>x}�b��fT���8�E����g��o��q��i�P��	HJ�P���P���(����J�X�_|�D0�XF#����<��i�����B�)-0��_�"d�r��Vw�	�� �i����"e��H�վl_/D����Ct��<�
1.�7&�� �~HK�2���N3��Pa�R���%iU+�t�`�dYl�fO�y�����kی��4��	VO���Ը�CzZ�!�ؙfAKU�;��y	7���i�9S�x9G�@�8�ҝ�ݼ	h��Ɯ�b�vu.��b|���5�N��{��GTB�R���8o\���WS�����zI{]Xyt�;d�p)�bp��#O�,���� Bbd�	�9-:-�-9�JM�'y?�\Q�#��"�ބ\����!{�ĺ��G4�H&�f v;p}7��*tH���~�<3��N`���&#e���I��UP��x3�X��uӀWf�*[~��p#�֩[-��4_�Q�,F�@�V��!i�)��-Cॉ����n㋐�����������c�'X,᫨m��j�ˈ������݃R�w�>"�6.�~�_D��V���{2���Uf&�%
W�=A��p���F�!������1"���8|G�#����w��t[L�ᥱf߮���Z*.��aR1�ƨo�\6�y�Fc�����f�F�9)�|#�G�n��U\���.4�tt<�����q2�����}���ݙu�J{�8eqe��(Q��`��#_��(�����t����,=K�U�:v�,��f�d=�3%Ϟ�u�CV���V��n��hf}�]�����fo=�DBI�B��'u�F�w�-M4~���%�J�s.ߛ6���>mO߉�����6i���-�|��4`����dJ��ӬRM�i��+a�$ Xe�sl�3(��b�VPm5�!�e�H�a���cG����k�U��*?�)1��c���B�ء�������5�e�����p�nu��������}=ެ�s�G*������w�(ք�J�SS��ů�R&4�~�i��y���H���~�0}���a�9�z�nx%3ԕbǀ���λ�>>+�F[�*b�	�b���� mc+�$�0�<�XA�������X��)y�oG���~��4Q���Q���.�f�{�ී�i����cM��^�����01�Z*:;֑&�Q�*���i�+2�B�	�8]$nY2���t��g�Lݐ ����kV��>�o�C�;�D\5��.��:./O�Nv��Um� 5��!h<�#V7�����`N���a��{ʂ����X�w֗<sA�!y��8g%b+
�󯓫��M�o�ե��f<��yƁp���HHjԽ�i<�w� �~?ˋ�z�^<��rO;?�cC��ON��v�'�[_8��"�z�}ՎEg�ß�K��䢉�|�>Bl`-����ֈ����0��LQ���U��d;�{��b�UxC�=e�O��q���OZ�q�C�aV����ʳ��I�$�ŋ�|�ag��|�"��b��l��X8��s�!� ��=v��f2�#�����;�3 ��P#�i+hw��B�o����REՏ� W&�Q>N� ���6�1J ���6w�,_�>%�]��w�1MU�0GQ_��7\�+�˽�+��,��A���"Vj��� }��)�L��ݓ��l�F����ۉ7��;A�O��>\���V7�o�R3o����,�Y�݃����:��Nh�	�
���+C����7�&�I4,@�HQ6�5�3%M�4�RzWk�Vc��B#_������h��|����x��5�:��;~Q|�p�X����J�4��G���z��.�-7��Bh!���pَZ��b�P���X4���nA�Y�(^��^��(&�kwOD9�-N�.-J��Y��A���bm{�~bk�5]���=��׃���msXv�d4�2�"�S�G|wk� yʺ��ྨg&��		��mp8���âp��.I	b�g��٪+���;�w	��0<ᨗ��p��Q��|K��WԲ�u�js ��*�O�"O�T�B���$�������Y��-�l+r�� ���m��P��֌	��ħ���_�ƂMm�t���oK�d�_������L7��7�b�\��=�6�88q�Ts�?� �ߚf:��4� _}��|�]�+����u������'��|^ �gA��Yd> �9�u9N�� 2&$����q�k髯�sB��0�\]�it�]��m�J%�Z��!�)[h�]�J�I�}���r���|���hF�:��:>�*w�T@c�U{��KY��[���6�R=�<�u8Bo1Y�t�=���h�KO���Li��x"����a�װ6!�j�^��~��չ�i�wT
V�.F!�1R���"��o�DT�m�fiq�//��:����o�S��s� ;yi�ʈ3Z&����Uz-﯒�[�\JB�^�7R�DmF����`�Q�����
EZ;)t����r�0t������E����"9]�C5�]�"�g�eZl�dŰ�Cʙ�nb�z���ѓ}��!s��X�#��j�/�.1�ǈ�S4�Ϛ�V�������֤��,@�T=\�[T]l����Uy���#q�l�mp�k����j�Y���&`N�4��'֟D���W>]�פ�.[��
s=K���HE�R�~ǅ��0{?L<-&�ѯcֽ�S�:�A�:(} a�t�/���`
�!�$~���B��Ώ*��ud�ܳt���O�â���Ϋ�}�	x�P� e	fV�?T�����Fю]���N�15ܙ$U�k�)�
���:�F�hWm��y��N��^[���	��������q��Z�(־�؆Q+)�h���<4KVRP�)�s�Gj3a�O�k�Ytm?:��	��Ỏ,_�
rrR��%vnr(ަ}p�7'鞯
�y����*O�J\M�n�Ҷ�������<�)�֚����� ���ĩ�1?���n�Ф�<����Q�&s�V45�K'M�&9WT�W�h:}g�G�eOi�֣e��:�Q�1*���o�ՃE	�Qx%r`{,����EP[.���^uC�r.��%~�k !�n۴����.��-�8�؝wS�<�b�D�6č,Mk%R��O�f�����������084% ������b� �*5�!�͵Х	�fzd�H�0���g<����
����K#��	��ٕx*�n�
~�,}<��<v���Ĵ��R�y���U��)�u��E!J���:��ת�#�RT��_i���Tq��S�i�o8���x�փ�*���A�$(��v��`�� 0v塣��}��)��=Qǐ�P� �o�hJ��R���������[O�1\z:���4u�y���V��8�|�����ľ>ܪq�0�� 3��~�d�]PfBH�xP�v�xp�"z�� EF&-A4P����e�ҵ~Yg�9WԧF���s�*���Z�ʬ���%�[d���?w_2��0��|T�(�e"�t�4�}�9N�?>Y�e0Rx��ڨ��r�]kA?����9QdUH�X��� cዔ�24��O6K���tS`�N��R�@[��­�pi݅��ƋP�/P�=�
�y_O��1�M����:�=�ֵ3��Ӕ9���LCGۏjY�eJ�_�?mlǑjvn7F�-�����$؍��햄 t��ѻn%`�FiL��Y����i�ÆNI%d�*>I�>�i1I4�� Cy]��t��lZT���pxi9L�����]h���0|�~�
�m��K��uQo����]�%͋����퓦F��&���U�I@t��x�?J�@�0�2�?�2u�D�����S�$�	��+�
檝�C�ڌ�"��h&CT�r��B����s�N���%L�2!�a����z��ؕ�\F[qZ�.� ��#yߕ)��j��� <����������s�1��a���Z !�l���.���C+�����Y�[��1a"�%E��"[pV}{�o8ٗ�;��7�G]�8 O��?l=g�~Q�F����`?�7�v5̊�������B��R����ӥ���P S?�:�Y%+�F���Գ,��S��W�đ�̲^-ш
X�� Ӯ��\��^����+�gQ|Rtk*�^a��MFV擝���H�o�@�A�C�.�p�?�<ԫ�̇}�<�n%˭��*��kI�-�e�Q����+��\%N���
��]�R,�
�a�#�)�
k��͓~?�Z��ϏI���a����ڎ{������
*�W=J��{Y��=�-�G��`�=kj�SsE��U�0[��5��A�]8�a��o_�vKe"|n9�S�T�r;Y���F3����ѲN�q2��Ь&3�����f�l��P�O���#��(d�?�꡶�B���eW%�I�q��:���,���XE�K��v�;;5�A �k1�4.;ld��j���3�1z+�ï��Ȁ�yy�]Tvʸ�*�N���M�N�*
��tK�ǂ>�!�j�b;�7�mB��kkD�to� �Bk|����G�b2�����~��@��E�d�6��3�(���mtD�%���ƮK������=*Q��&Շ[��|�R��Ӹ�v�(�B�IU���z��N����>��;�˵�眨/�A|M$Tf���N�`��|�,t,7lB�dݺ1��2�ETx�(z���u�O{R�G��t��D� �4�J�G�ȋdWG���V�Ժ���˅xME�,�3�C���_� b��r\L4(��ݪ+͈��z��q��v��^D�z����WҥpC.9�T3�^����I~���(�%Y��v��(��I�r"���_n�.b������3:C�|��<�pw�h�V'��
���G��a��V65������]����%Y_6�ʐv.o��<|]H0�Eb	�ѡ7�0���LŕHˌ�^��L"JɝD��;GO���n"M�	hX�Ǯg��֘&9@�am�MԢ�J�A�a?5��b�Ko|%K���Ņ��&�o���� ���y�tI#�K��x�q[���!�쓾���w��aW�4q�*�;������ؿ�#QV\�=���|�#ɊAP��;�@�D�_����w�|.j@:=�x߈ZB,2w��l�C)�\�b��ߛ��;7���l��Lx�hM-��"���d�^�I0 Q4����Ͼ�f�9���θ�>���6������,og*��X��dj=�`���-�O�<�i=�]����gY^�hEi����x�+t�R�?�f��`�q
��h����=o�H�SD=,s��XmQ�lӘ3�__�<�H�MՄ�b��&ѷ������Z��H��re}a����lau����WM�4M���������m7������q�\+�Ğ��Fci2����������_�Zc��5�����*��$?݆��jD�����sQ��� )(���#����b.5��B�%Nl�̖���yÌy\� �E|}�{k��2���E2Z\�G�u#S���:  �*C�<��nw[@gT����M�%����uv�y-%�I���7�sXL�]!걇
8��m����b ���T���y0�X�J��-=�W�<*O�qyFq�3�!vR���;�:���Yl,��ϧ-���uI&�_�[jx���a<�!=`�u�[�26�~�l�Z�p������M8�Q�#$L9�+0�:G0��;�d�̟],#<��>�G��x�g�Cn--ݎ�Su�B���X����$~ɍ�⪘��e[N_/z'{�i���3�K���Q���G!��ӡÚ��71���Ȯ�/Q*)3����EV��1B�ߚ�/j�g���L{�;8Q����{'6���^�O#��2�'�Y�_��1ԁq>L�}if�B��3!�ʛ Q�R��Txb8�KhgkXs`ݎ\&�u��,I�=j9��L5'�߅ R����#��V���f�P�������b9�Bs�N)X��-�%�	J��Vo�b�/u4!$�� �2U��������d.= �\�3��Wjj�	 b�B����n]Mp�j��]Җ���}`�[)�Q`����q���*L,�{3iO�X���XY6��z����"�=[��C'�0!&
�緽����g���im,Y�=~�����$)<���|��r�D����T'�ťJ�/3�p��<I��<��BL����%q��I�K�e�5GxH	��fw{��� ���q�׿/��'���7�J�PAW4���0��b`�*:��%A���bϩ�/PA:�r���d�x�<L&D/�_l�SGA^9������ GZ��ے�^�r��ga�d�21X�T,<�>lhξb�:@gg�������f�֯�1�;~�]�Ӭ4�����e�����YS��b)l�2�'��;�[|��w,f}Yƿ0JA��ظ��#��sZ��$Ar���>�˧�B|��@���
�"<�jI��/S�$�Q^�r�:��*����������.����Юg�����	IK��q�z
[�K�L!6ւc�i�!=�Ј
;UƠ�u�z@L� +����A���V�"��7�T��>���^�Q��F`S4<ܨi	�%#l.w�}P}�Y�Ɵ
�e��%5'׏
��@�w���Gmc#�:gY�^���'T�5zS�Y>�>V�{�Ah��v�oQ�~p��z>�@�����c���S��;�%��"���s�VQ%����ɍ��iN�X�T��
Lǟ X�@�EӾ
�a�TW �=nuLoGnp���g�nyP�"h����h*R1����,O-���j\?0L���6�(8T�eo�fљ�OwXZ*�s�k��t��]�o���׵��E�SefH	�������9�¶j�T��-^�ޙ�H-I4I�z��B���F>�mՀ�珇�B|�$��˷� �� �l�����]�8A�"u!���ʪC_蹅���($��!^���
K��0+ƒ�9�b<ì����$��]9�c��p�)g��I}�3�_�LR^0V>��	]�I3�G�g��f��ܿ��w�.��'�҂�0/J�3�)A\�؁���/�3�ю�h���� ~�͆��)��P�?��M��WDV�Z�F�6:�&q*=��fX�N�6��Wф���#}����ثD�lG7��!��ȂL����'�<q 9��i�l>Xu߼!�Ĳ��Qu� �l�������T���q�ˑ=��h_��V�[�,>�G^��elb�K��TGw[4�E�=�KX`n����܀�ΖG�;m4F�]�,�4���#��s�s�$B�U�@�0��z�Tݩ������)�ٕ�?�f�t�����>�
����3kz��3鞕��eW��d$�"�ڙR{���]��o�6�1f�c#��^��K$����g2��=[g&�9�a��jiX8�LB=A�DB�^/7����|i��ם'������5w$YwaQJ�g�'�<��(���|�+>>I�~؟��iCRū7[q�-�K���� Ǔ�O2��x�j���[A9��;N2�K8���v���wk��뛦�6�Gy��nBz���^�wD�±	Lt�G�!�|���o�߻Y
��o�c�Iϡ���H���Mi[� �ķmey�s��>Xj5�_�?\�ŉ��%c�-BB>�ޤ�!�PU_0�?��p.]�:[_��p\�}J��)Ie�����Y��u�`s۪8��'n�����Y��P��Ƴ�hfpEC�*t�PX����6�?{���Q��wJ�#MR0z�0h���ɀ��Kb��b�*�V��ۃ��pA�PY�M���],�>02;��ˤ��E����!O ��{��1���L,k�W,.�[|�v����>@3H%�{���AW�W5F���tH�"ף�7�d����M�R̖Y6@~��:��q��az�,�� yK�<�u�dmh2���͠=['s�~�39]�Vߔ7�W�RP�>��/�)Ya�|A��fx�6QC�ϧ?fN�(�<Df-�44A1�2����ov��'�*��^+�%*i�ŧu�,��D���_H���rR��$I/��D��L�@���}U���ζB���m.��;L� S��y���mf��2a��gd���&n��ml��F���m=n��K��u������̖xC�+�������_o��9��{�"Kt��
�h�(CYKӄ�H����mط��0^����2�n��rfy�MoXUx�&b|���E`�Ъݪ�rn%��SGG�������׎�A3c����rP��'�<)��ePZ���kʂ�VA�
VyHrpF�2�5���Lu�����y�;QX	Է�pYS%���,�.���B���m�,�4��^���I���rZ�l��^�������6?(��*Y�:\�.�u��<:�Hh(w�Hz��;U.��F�<'w=�4�#_���zϗLg��"��mȆJބ�m�~�@X��yۚ�f�R|ԕ��d�ح(c�n�'Aۊ��y r]n���	#T��a��cԒ3�ݝu+�h���z�ҵ�@�^�<�I6*���Pɵq<���:���� �0f��q��?	���"�7٢9�5p�y�%�TtqSa��V�N:m����Ɇ��qv�5�)�����S<�`z`_V��0����\PS�,�hN��/��A��n��C�U��ǔ��ux�yʀ߅N���ɿ��KwE"��AC�Q �U�"��*�oI��9v٤1)�ū@�H	�.xL&�d!�?�7���Ls���;)�(g��[L������#�5<Gow�Dx�3�N]ǿ�|�?��`�,�g�����P�B�\#���).�;Ϭg��j��M.�T���N��Y����u  }T�@/���e�K@�ևu%ͷR�3ϼ}�$ܧ?4��P�I�pH��bt���w2Q3=}Y�C;�^p�M[�Q��5��o.`g��',��p��OƮYȽ��h4����o���P#uW���nlbS�3O�~<���ANK��7����6�ٰ͇$��[� 7zs�$H3�Uf�d<a�$�b�rG�����z�k�"��cF~0`Ew�q�4^���`�U�ʢ��u�6�T�Z�������Y/�-��:��-)o�l��>���@��.�F��`ޤ!<;�H�	��z �
�5�"ρ�L¡�p9(9�=����,��K�9+�gݧ��O�"�"��o4<�Վ�HZ3ڰ�TFmu�fB�j��5) 0��Ia�e��4�r�@�+�&xgC��Z_����$F�r�M_��4NQ�Z,�����o�o�.�����]�+5E7/nw�owo�%�:G�7�K���0]���>�,�Cۑ �8Џ��bU�˱����D^Mm(v�rL�%�ɓ�5�'�!|jm2q��F'���Ǥ��	��Jl�?4�bDnR��;XDU7Rz�\zj��3ȒNe�%`���Kq�#ՙ��	��If���Rx4:씱�i�����0�g�5��&�}]����]i��CJP��Q	�F�8o�b��$�3�E��GS!��i��
���؝A {Qr��w�b4�w��W/���7k�Y�p�e��z�	�;r8�4�G�c�,�S%��T�i��	�
����T3_I	̽ ��;�t��o�!�K����������m�UY�����&:�!�Y+�����I�y�������|Rx��K��W��"��R�NlV�S� �#�s5�U:��M�Fft�:;�s;v�>'�u}�O,�%���U�����Ab !�����u�~�%�lo�B�CD��M��V�n���?2���&����$�F���ً��C,A��sn�N��b8W���'�����N�� �E�ԯ�����ռ�v��۵P�����+g.�8�M;�՜l(��7Et�j��*���,�k���Ϊ��%ۻC3s~U�;�;��GRzG Z�"��Wj.ҿ��M��8,z�BݡO�H�� -�~3�Ϡ�%�G�B�ӷw���P�V�_��f͕�KxO"�Q|8�4�,�W*�I�a�g>k�s}=�[�@S��)���If1�\�&_��?�\�Zf�
�4��i��&dl�w�.>n����
��y��l����%u�˱,��p
75Wk��։_x�e�4\�!�f�N�u$�$4�`qEQ��)��O�^�@�z̳T�`~���)��1��Q����.`�A�4��∛���Ķ"�1'�B���e��l)���	
%�W�|��.<��Y_HQ~a�(�Sh9��'ڑ'%Y;����v��m+�P�G�,��0C��C��3�e��*�,cs5j���q"�4�s�����\���R�(��I��آ�Mk)ގ��Ck���QtUs
��t����p(���k���dHr@�=��OјHDa{�����],)��#�c^�wFY�ۓ��z>��J�'>���L4@r�
����E�������b1�Ff]k��}U�1DX<IA��:3#=:t�<��e�@����;KSH���V�{�
��G��%v�XO���i�:�X`R7�ʯ���P/��;}�����2�:��ſC��*�!�,%��ZW�f�9��O���x�d�Ř��3j��@���L��	���55��f����ח�z/A�����/ c�j�W3�!�-���"����@�&�n�:�)�A�$-���9�g�e��(Z����'4˪�[䅫\D*�*��
��B}H�lS3O�K"��S��/��?D�G�0N��Mh��gkZ��v7� Vb�<�p!�H��2�p�l�u�?�� �1v6 ��"毜�웮qS�>_�L�c�7����	
����b� #��v^!4�V���rt�7D Aa�k|#���eA�P�?�P�����\>��^�cc��<8k��z��
��Z�A^8�,F��oX��|�h�x�2���.$*hʤ��z�K���ev?2�)�f�.���%������[$�ι�����C��y,݇�;�ل��᧕z o��敔۸�D\2������"��^��#E�����W��������<V̠%�_󬊪���\�~/�B
Oun�� �ia6	�>Mc��(eٲaG�&'�_K������(��M	�HP�������d�|�3��Y�?4��?�}�96}W�<ɩ���d�5:�uق�����V�������r� H6H�	T za��l�U�1z�f4���d�Mz����}�՞��� P�:��1��Bྖ!6� �Ƌ�@*����1B>2�����)Qg��c�I�����Qq��r7�C$��tZ�KH˥j20���E�mk鏶S�螯
�A�˾|Ђ���X��5����!gVYXRu��0=cD��yX��鰑/�a������D�wm��}i֜I~#Sz�Q��9z��i^�W�v8�g��C ��=`S�)�#�嶹G��ćzwG��-����Y��i�`7{J��T�� /��ˁ�W�Bb#�U��gUR@#��g�0��W��g��Q�'�ǯ��_�oqǿ$�Lu������D#���yh�p�_��1�͂!������Dj5���+}�qU�4�q�����<�fJ
%���299��Ѹ��Tbx��yX;�fj���)��J�M��CГ��<T�r>�;4��qϵr0����r�������Q��U|�� �b���z5 �r�I�3�0MM�NN����T4�����KEPP�� ���]�(Me�������O E�i���1��i�B������>��f�[�l���ʶ@'9�Eo���-n/ze̼���%s� ����L-�j��Dưh�30��(K���2�I1��)o�3N�G�'>��:h�-��AE1b ~K����CHO^����p	#l �_���*�"PF � k-���1���^l(��]�h���B�o�P���������L8l��=-�a���UD��F��Y���ah�Rv�?r�,[��]ƁԔ����]P �[\F��ȂQ�st�������	�|�͸�x����	 ��kŇ;	w(Fq��m�c�L�6��厍�q6���u����Km;��t��c�"��I-C�t������|���c�ۢj|-�g�H��2#jo���7cױsFk�ۗ˕c�?De_����F��!�B�*p6?#��d� ��tG=d��hm��K�0v�{4Ł;������mVt�)�2���gL��;u�MFU��x����M��$�\D%?}�Xg�,"K���I��J��6�#�$�Z����iˣ�Ds�T���cN/���<X�����t	]�����T�F�`b�}��<�Ѳ=�}��G��� *�/�����1�F���6���l���qו��u[[Yp��:~�W-$W�|Y}ݣj@!�7�L.��u�����SF�9x�pxs.�Al�Zms�)Q�l�{Ё7X��Ŀ|����ŭK�7T�u�N�!u,�-$M�|�����8&q�a�}�L2�VKuSX,ǌjg��58s��p࠲tN�-���S�4���y����n��!�4�p����n�YڭS���uP�c�K�R�Ev}����@�Z����Ўc���y�W1U�:�(�kU���+7�J���o8`�(��!#�"��r��ڈ:5a��M���M��i�65wn�8�vW�Kπ�����2f߇�W�*�i��L_>/��U�Ŗ5M���f����p����}���\=Yy��n�3�%wG��b�+]x��s�&�u!4� ��{������ q���~����l���R�tn�J3�ܾ���G�!ԏ��v�X&�����_�N��7�$*��D�
r�S�Ɵ�j���8� �w�#�U���!� �8X��#��\�sQ�##�G��<���<EVzUj��7o�	m�2���lS��l 2��M�&�ae��^ᷛ�Nُ昛.�7!d�㟷���<�����ƳA=��Y5�A~��+���|D8Y��śA�����ȱ��"���Z��hk9�kl�y�$���=�
jM�_θ���1�2z��H�Z>S��yn Kher�>���p%�˴��w"0߳�B� w"��b��t��&\Mjmi��wI��Ǥ}�7�4e#6g| 	ωT���ߜc��GUܡ�\��;#LOy>_6B�[��
\h����7���@~��w��lt�K棠���4�m��Z���zm"���Ⱦ"5pr_��n��(����I �+��G�§{����1]�+Z�����W<��s��g�+�jC��9($�I-� M�B�ٿ"C+"�Д�c!�ԫ1�c U�!Df&�K?ϭ+�?�b���/r"���۠a�1��B��B���&�U�6f30`�Y�"�@�yR�~�j4�E���h�A��tnɘ��pWx��ֳH��N��Ƃ&}7�ĨS�TI[J���g�*���e���5�� >d#��J�N%�l-��G�/au\صwS��ʅ!���k�ėM���y�9�}z�8P��VgNBb� ���/A�05�$r�o�N�����;�x6PL7��X.�"�ɛ�Z��/0���=z8C�� =���;��M��]�WW㊾|:�S���ϖ�����Qso��gb8� �=+Jp���uA6�TƷS���A���y�'+� ?�
�?<8�r7|HqA���v>9��?Z���iti�C�a�������e������2�g��?ҥ�,s�S@���|�_�YZ�sI�J���3lͤ���$�f_�䖯��Z�I�@�I��ڝ`�SH��)Ӯ/�ټg*���GC%�iWxBwxɯ-��u��$�����"є��W��v�L�����g����Å�G9��1�fk�$@7>r��AE2�Ο��|;�G��Z۽T�n}Ž�8����tOr>h}��ԠZ�9�������|7���앁�U&�	�a �6j/�� d���n�:S��D@�3�,����S �]#��5�S�������ڡ��+3�x�ءl�*�U�GH�̻�0�Yo�VC�>���n���ڟ�W����f*�u�,SC����%��R�BkT_��z�_G��t�\u&����`�fA-٨˵uҶ���*BT�Ћu���>�E��Uy��\1��#��7c��A1���\��>�xz���a����ߤ�ն��)=����Mıw!)i.C���&`�gF���~[�̕���`��H�����?P��\pDLz�iD)TZF���2�W9��5�e�U�k�n�#Nr��������:�]�f��ń/-H��G݊"Xm9@o�'�q�9�C�{��tc���d��O��}��t���0�Ϻ����l_;^M�[�p��8)��n�D��>�L��Jf�r2����)��)���}�fT~���՘��I���=֔T�ᾓ�c>(��ڰ\���B��Nw�����u9�/���p��b�8��J�"<�#j��w�ЍNo�q��y�WL�zu����N*�F 0T�7F;� ��ʹ΄dْ;L�p2��0U��8$���>vb��jS0}�_��M����n�]��Z�n�L����Z��c�<ޒ���ѬX�/��&������𻆖�D�S�UP�G�
��.���8^� �C#Pa��n�cL�زF�+��ʢ�������ʡ�qF� )z�t���8����P,� ID�g*��S�So�]?�+A����"3t��]��u������֗&��bZ=�ڡ&j`�R�c�4��bFp�\���YՑ�K��Ç����<n��Ԑ�N���ϩJC�����8t"�J��)�;��r�q���c�p�!�X>[��Tۺ�C���+/�B��;�P��k�:�>�\���=�r"@�B����;W��Lv�D���=�D�Q�^�}E�|*�C����t���pu5�n�o�j�P�VX&��{�&C�Tgi'�V^^��Y�42T(z�V��Qݡ���W��� ��nI���O)L��R[�$��d�OA�+��C�5�Ĭ���#���ũ�2Āa��
%�aB�Xz�Y���Q(Zk��
=��>E�(�S{\=�%�&�h(�%��Z���;'��l�3 �(f��^��P��¾�S�67�"X�W>����_���m�(
C����Y���҉�H�1��c��F��㨱|
=SBJ!8|��9�x�7�$G\��! W�y��Va���9�v�,��	aOM�|H���J�]��W��A~��J��7#_�����Cm�S�|�iq�~��y��UI�;7 )�=�ʱ����i�R@U|�[�;{�$�$c� �.A�ꂙJ�׏ꥎ	L�O��V���׮�wD�V�M�z8A�KK�����|�O�{�[ �Sf����gS� �A~*�%>����.���~���SO��:�c�J?�9\ka5��T妋�/ru�D�����4���'�:��l~����yBtu�ni�����U�rU�2!G�}��C|�+��	��� ��f�޿\��i��䯖]&�Rڢj0�<��NUc�w�IωvT��5Cq��2�50d1�i@�a�j��M�]������K��%aƶ�U��V�y��x@����Hf�,��R+�/Z���#�!u=͑�A|�n/�>r�T���Xu8�gh�{���̉i�IFu�
6��YC��n~��,�ێ^Z`$��%f���� t�*�cƟK;f:��캖4r|���� ��3;�~&%�˄��}����#ɟ��'��y���3,)��'�Qrdd`�}�ڍ��	�Rϑ�չ�އJ�{�o�#�2Vr$a���+�S]�֏*�!����4�VA)��D�����u �f��<��_�\vȶP�� ��@��n#��t�O�r�r�~���{f�?��iJY�u�_GgpE�μ.r���ٖ0^�>�5�?��$p/7b���ѝ�v���n#~f?����["���i_ oz��Ź�Ud��^�0�O�怌�(�����ޮX�����?��\�% )�.�uH6%�[A�Z���]���o�6Z�k�,M��#o>��ab���TU�}�WI����XJc��k|��eNbq�&���9������%r+t��L��[�%ټ���G�<7F�t�R3��H~��b�uc��X9Z����:�S��K�J�U0��#�n��t~y.�9��x)/O�:�v�y`r�{qԾf�/�Dk��p�bWt�A��N(�A�[��U}����gA8��� ��1����Weia���[��c��+!��<��w_%��Xc��W����E2�G��mįd���I�_�ڂ��@�@۠�Ɉ�%�6w�m 
���]�0��?����Zc��x�$����n�D�'uX[6]r�� r�@4�����i]Ѽ�R-8�A�M�p:2�����Ǿ�Z=@�D�
�uGm�;��)��ȵ��n�������M����P�Wf���d}%��fl���d����wPt�(�K?���v?t����Q���Μ�ݦ%5?:��g��m[(J�U�}�Δ�[Kץ��3e��h4�c(2��C ��:�l����GY���0�">_��fc3vf*�����cr�Z�����C��F�^Ӻ�V������̼�Z�3�N�Qg�.�D��m2cS��I�>��u��=yİ�n3�*��5q�N���i�g0��/��cO⍢n�'5���z��kY��IA�S�\�c<�+$M��k�[cAB�7�μEc�<�f@��#h��l����[gX�dV�6¿���5P�Y�\V���9i�C}J�����0��oI#c�4--�\��#�Z��*BM����V�d(�I�컨ɪ���KS�[\Ex	���IE8X�N����G�jڭ�.h.2�b�)+A1�J3�g��)�$.%�q�.lJ���B����G�{��k�֗�������Y\K���h�0��E?0�@`�oẏ�-d���\.�9�W���NW�C9�^R���>2�6�Y�؜@/�@�( nM�7�J.��N�J��U*O�~�dٰ�qF	����-v����=1�����¢�S�e#Γ�r���5�2ے|��Y��[����?.ْh�k�fc�!�ءL͎N2�=Q|������^���Z�sM+��s�j���W��ɍ�g��?- �1I�MS���*r*;	@�bީ�R��'��n/�9�~.�(죲R�jZ5E����rA���l /�	1��38�'��r���� [�ۜ؁��#Eu;���f�z�؟p� ���Q�OU)G��5�����B{Ij�Gy�4b8P�V8����%��,+M-t��샤��[�\��9X:1���Bu�n4<}��\)��tf�2������T�c8��;��>�-�h�Q.Dz��ĚY����� �'��*���T�6.ͭQ�QP^?��X�ׂ(�1�Y�8!񋔁���\�6�vb9�i�I!�9`�_V�K���kf	^� ����e,��|�
��;��0�D
�\�K�"�_�m��3`���3Ǆm��b#�p^����&/%F�j�d�,�l3.��ˤ�E���S�����sT�l���ȃ0m&���XlFoJ���c��7 �=+?�/��7�_/�<<��Dq����|��~��	hԗ^Qk�XA���(�R��>��z�Fh��G},L�i�#.2�g��Z|�61mq��Z���|BT�B�{�܀��*j�Ӫx$��sב�@��#a���C�(&|�	��q*�A4*Ql۠H��L�Sr\>nѧABy>�I�[x8��;��Ӟ��YQ����&��7�>.�=���,:���ZB���.�>s��ߘ_x�3���(�߯wQ����_B����D�z@�EPj!UD1!����ݢ�������2od(����Y*� k&	��6<%�$T�_��	�E����eB/i�VR?� ,]|�n�_��C�shr	�N�_{"Zl��m����M*�39�#A������4�@�2��#*F1�V��}:x�x���ӵ`9��׍A�a�7�2Y��a,�t�rK�E7f	�[�Gə�����>��tDy����-l8s�5j�i�r�#��B�J�Wvn���6M3m���%>"4�5�b����5����/�
�u��k2�@�Ֆ�k,���%$�W�]�ĆJ�U�ʘ�S��I]��V�_�R�0�=�����`��'�Sx�X��t�z�s��+�"�f�T��+\ y8�\�.���N���������RǗ�1h���+�o2:�3{��R���$��������ƨw�I�g��#�}p�nL�UJ�c�r�tQ�͹E<iմ�$Xu����Z)����-z�4=e�l� ��e�^HW���3נ�os�<ؠ
JR�v�ɿ����6����!����� ��Z3�|��"��Mh6d�jr7���K����;�txZ]�^���~��p‷t��|s��/�eۜ���dXd�~=��^R����V��%g􋎝������)�[4�mT�O0�Q����@�<�!�z�#����3f�[/{#�ʱ������'I�F,E��˷��)������Fv��&8mom�i%@���(��9B�C���1��n�}n�R[շ��%�����/��٣$mi�f��պ��G��'!�i�T �����+Aa�U��GQǱ�?�b��肘l�s,���%����Z~<����a��t$�*Ҙ��nz�:x�ﲦk��j�Jn?��
z��)LZ��.&�¯bM,k��-�e��}a�Ա�L'���|@�3xCvH9��� ���,r�#gk�ؠe����KYɏ��ɘA?a��,��erR��/z�n��	v�b�����U����}k�%�#��5U
���;E�q_`���Yȴ��J�S��+x��JH���`��f��Mm?��8�i�����/_9ܬ������D�ʿ���=�엊��B��^V����WA�f���XT�g��o����&�zъ\9fg�N�wJuP{ L7���<�����-	��q�B�N�O��Zy1�թ��h�0Ж�M��h���G4wj��!*&?�{M�4�¶/I�
O�+�tG�%kO�8ޑ�i�-�@X\�r��4j�v��Ǒ��}_K���#�<r�vˌt<���:���@(&�o�ܚ�nX��w��<K�q�`�Y������jA:, ��*�L.K:e�7C�,�t��yGm"��^G	2�Ί�o��j$�s�P�U�Վ�K� h��է��f��33�~v�.ek�n�;^�J����>Ҳ3.bOG$���hWL��X�*��֭d<��tu*���f�6$2Nb�$���e��mW�nd][>>��x��UhxGc��̗�q���pܼ�[�Ew^�ףH1}�J�]������)�8A3#�6k;�2��><�L�Gc�1��N�3���8���m�������w�v�"U�8��](��
�s�h�'����ՠ`7o���abG%|���޲ɠ9f��2?)ʤH�o+9�\��Rj�6|x�ګg�q����q�s�)�ݱ��~�^�ǩ�ž��+&;���c>J�JaK4�SG@��9#�}�����XS�Q�<��oD�t��퀪~ŗ�n�x&q��h�3�{?X��J�6�|����Qy�A/[h�(��T���k��k����>�#���û��G`�`>P��O��K����5����O:�"v��,sbG��c�u*9t�N�r�k?8�<x_���4�U ��V��^�	��z��-�ۍ4ΊK��!���l�O��Ob�V��Fv�ϵt�rN����b���ޢ���
'C�/�Q�W�wD��b1Q\;��Ǧ`��y"&��A@ ����zQ+��4Ι��(��t{���<�R������)�HOc�aC�i��d����~���n���w�jʳ��S���:���U�A������G'�P�(�)vj��2o'��w����P!-��k�|u�痷u[�qW��)؜$�׋�Ks {(<P�1��q�1��S��;�9/�<eJ����1m�0��Z<�Եs9o��",��|O����M�9�]eb��E��G��}�H$}�N��h|��|�]��K�;�o�P�"�Z-�̆'b��4���߳���*�S_`2|��������{�_�1�2��Ɩ�_�譲�#�@��ۂ�6�-(����O��<f$�4x:�'�S�����1��K, �����9�Ð7�����A��+e��j>F^a�������}4�]��=lW�Sq9�,t��0N[�J!Ü
�z��LhȠ�{�A�biq��fX}�� P�;/"fSo�\(��C1�9*�ʬ\�ER����
l�U���)ϩ���hQ��"	kH9Jhe>�.�R�����,}��������Ϙob�#`F�d���CUW�y�B�Y���2̽���r���<��ߵ"�axm$5c��x��a�)��:�7x�K8�:���m5�����)��K��O��-?p2GF�֑#�Y�����0��uBj ��c�������q�x�? l�>�3��ĵ�P��p(�C��cW���$*�Ѡ�iJ�����3h�ǒ��/9#3��Fu�*�d��F�z����'fM�"��9�歠 
=A}��<����J�<���-a�����<�<���k��}��d��X:? 8���v�ŧş�p���:�*ɤ$�rEn1x�g��Q��^���m�l�(�sߠ<�"�W�Xp�G"�6NE��Z|��f P޷���>�5����(t `P�V?	��ES5\_�Ή~k	Pm�C�����ѭ����ɻH�n��t,�hj����eށ;�?�x��fNrM��ZA���v�����J,���W6�Qk�f����y������8T��)�1�ϫ�8�nvls������&�r���
�/>�s�6�:-��h�]����S YE�&�4��?�'�2-�]��nMwN�GIţ��$�3`�LI6��w�ܚu!Q1i��ؘ{�h�0n��0xG%@i��ϟ�o��/mr�H.Qzr����WF�ʆV[��m��Q�uc�r�����+`��O�e�1���X$։=������O�����*�M�\��$r��KzO���ɜ��"�������nYۙ���'��r	"G�=��S� |y;Zm�{IE�)t�h�X�	��+jC_�;V�bm�_dL�H&�T䔅��'Q�e�&~Z����M�'݂E�4T�F�dO�J�g?��zR�t�Ѽf����mn��N� tc5�[�k6���!2=I��|%v�ʫ?Xk�1=�Bqq��x<S�,�_�n�^�'3�6_�~yc�7v�5vI;(`�|2Ѻ�m��X��̽#xF3Z�~�0O���5��3���ȼ�X,Ę�h$�i�����ʩO��%{����:�͔8M�z�L�ĉ����|h��0��z��4�W�������vb"ʷu�a���!��p�]gi�1��U��9��,�3�Y����#0�p�7�ey[Fl���B�2xAeN��,L���]��4��3�F�����8��	E暄��0�-g�q;lD���dn���j�cj��^�a��p0���,y8Cx�z٣HcK�C���e��B��*�u��d\����RzW������-}z�cYs��+�6��������ds��}�+`��bm��l[��25�=K��b�=P���\��Й����î����ځ	y�D�oMU b�>�&nS�$9ə�[W[����J3�0�6�nB6�b�mCO�d�6�B�~�i���Ȯ�9Ȥ�~�a4^�=oL>�>�7+�AjI�?%��G��I!Qfd�y>S�u��k���a���D5���Y2{#;�:�R�i�K�R-ƜQ�?��в���_�{My���	`܏�e��CR�2}�Dơ®y?���q���h�{ϒ��v8a�\��]W�B഍Qm��U0 ,�m� � �_<}(j)�-u�0?�`�>-0��TaQ�R�IE`���/���:c�����G��������ݕ�T!\��{�9/���ta������]x�D�k������Mt!S6�}��ܓE����j�,��"#���ZL R-�6�{qH�<�_���uEw(Iw�&���i�y���{ҥ3�9Lkd`�����叆��F���8Hl4ȸ9��� O1����!^��cs�r;�����;�?�N���^�u���$e�ء�RԆ�T��txuܞ籂̄����B�Q�Jc���\7o����˯�g;Ж=�$�<y�@F�Td���sI�a]2?���I���YK k�v
���2��ρ���Ra�%���c7��[�/��։X�k�7����e�,yG����J�L���ؗ}p�Ey����yɠ�N5����}8U�������!fZ�S��K���D��8��9��hH���0�O"7ԬbX�(>q����74��H*���y�D�$�u���%1�' �j ������ |*��X��3pY8��S�B���[��P(��'���==�kh	���M$m#0��8>�|MG;]HD�ᚔ(��-�M�"����rRY��?1�Dv�/��Ʒg?�h?����}[r������7�sL1i�B�][|�t����N���u*F'҄s�l_X#�}�9�Q��Be&Bʼ����KC�����=x+߻ ��1����5���H������D �'Xk>A4����_"u��L|��E���&_�Q�:�k�Glj�j5JA%O�V*��k +�ߨ3i9�C#Lw������x(��W*G(�5xgcء��w'�l0���?I����¦�g<Bؖ
..X�O6��_mH���U��,>h3cCR*f�A?��1��ɥS`��P݃(�����Z��m�I�YԔ�5-���L�y���-���q�B�Կ�JܦW\���t��ﶯ���8��@�`�!�u�s�-��n��5M�.����%f�lVz����2=_;�#e�R�L��}��'kܯ��iE2�?���Ak�����芖��T��zz���;�1�-��GN:�~-t��������j)�f�E�4�O���I#��>�Bt_	g��Ţ"ͩY`~KGq��$�R8�����ȗ*�����eL�&hy�UX�Z$�*ܥ�1�H��+E��
��`�:Q79�,9X��C[6-#��-�[�˺dP
y��qnЧ1�$t�]�S�Ş���T�	L�Q%3-~p!(UDS�>��	Gk�0��V��k�h�X�FL�2��wJ-I�v�󸬠����Fo8���X���o�X����D@�����	�(��P��7��7~�l����9J��t����3�h��Zb��K񽐮��8�/W|�t�f���A�N���ɿt2V���q���]��)�"�a~T=�n5Qㇷ�1Y+�k�q�Ϋ" ��A;�<���''%e]��>_���LE9�����d�|�})�V��=�20lKp2��Fg5��8��܌����ጵ��r�yMx8�3��C�_�_��k�R2,B�b�{lC��&�#�e>تz�!ٜ��ƌ���D�j
r���֓���Ο���oA�XZY@��)RM����9\��0%��P]{���H��v1h(��[�F��V�F����[���M�k�%C� Jio�h�"�R�p+��ѣ)�V+�}�W�v\��2ɻ���{�L�X�2���&�t���YG����o�.�v���| �P���x�Aa�ߙ@P��r�]-�;4Z 3r�{���o��+#��^m�dܰ��r^���RT'>���}X�C)�w���$z� W�=Uk}�BI��!�9�.��mڏ:'��1��������4����B�#��_@],0�zW��U��U�[O�j&@��B,��{P����Q��x�*M�+��Ad�$h��g�S�ј̓8W&DI��������αn=�,�B��#jh�L7��z��!�`U��^ڍ�P��8d�N
�^ĩ@p��>?@����q��/�����g�E�
�N���Z��eR�c|���o��:L�D��~��d���Z�$��Y�W�=�T�0�0���WK��0���s�9eև#m�Ɛ�c-J��ˡ���U��(N��C�*M�e~�b��I��ߣI�����sݓeau//�1�]>����m�6?�������@f�d�J�w"G��ʔ��;"�w���ڴW����+�M�B���j��õg�^yq��ha:M���Gd�"䪖�;i�"z=ljļR��[�ֵ�s��&�u�|I
9r>�l�Հ�Ņ�u�{3��������_��E<��%�?���s����6*�D�rud�`M�����WxA_�Ptb�'���m�B:^W^�����f��?�yt�ԝ�����׋y��`���5�]vg����8��9��A<�u������nU*��'y1����7�ܑ7�u�[�}�53`d���r�I���x��@�dTY� l�݅����-Z���̠�+��5e��.N���{�_�K`8B,@o4��#�*7J`�B��hLi�R�	�!�J_�G���$��ߨax���g��%4��i��7}�����<Kf��e��I����H����/��a<#��E�[��Ҩ68��E��V#���{��߀�}�'4"~�v��;�4L���_�ǔݖ���ϴ3�ʂ��G�ܢ���j&7)*�	)jQd���A�b��g�eg��|\��^w�8��8=w�m
��^x<���n���h����j@�8��d³����b�����9M�>�rL66jNL��,`�d~cR�W�܃��$�y�a	+���]�`HhJ�.m(j�+*�qu���"��8�B>�ۖ�cFF(�
�A,'�"n:4�E�sUd5��̾���cȟ/� �|$���-d�\E�����ǒ.ҎSѥ�6�[�r�X_��X���fŬ�PFcs��#�t�����C�1�E��͖���H�	����,C�ރi�tgh�}g�?nd)��"�
�,g Jk%\ H���ͨ&t�w�2,�I���2�X=���L3d��"1����&�ʧ}�զܬ��P�j���E�i���\w�e��r$YܖN+
��2<�D8	H�!�G��QP(�6��)��G|�S�p	��b��&�ݢ�����z��� ��D
:�U�������ESy�h���{�5���z��H�Y�`�U�KJ�4+���4Ӑ{9���Y�O���pE�Ac���y�����.޷�3����bgpW��
����Gg�S�l���h+��{v����u W*�셽%�6z���UȄ�c�l����+5�3n[�k�*F�v7V&��g�ִ�;[5Ef�����mŖֺeI�&�q��T�=�,i��ҋ�lq&p׿��cb����G���[6-���b"��;`_3˩�"$�'�a$Ӣ9�GK�=��ER&�ٽ���Ԍ55��[���ޕ5�����f��*��!�����ӛL���p�&��v"`�ߟM�%����^:�=�e8�<wt��uE��r�Z�J%��6���t%�L�Ӟ�?�J���!l�ψ�\�rJ��ig�0��N;��Fpƥ�n^B�N��C�l�F�N1
;����^H]�C������>����
�?Oa���%i���+f��F��,+�g��wrѓzX�������3K|���z�gLE���Ķ���$$<�Gq�s���|��?�e�&ŧ̓e�X��1�g�~��+��
hS��Zhe׍�`���?�7����D�ۓb���c!G{�`�	��%Lc E�#�U�K���:e���-"�k��c3��n4�ٓ�GN���!�[�a"o�P~c���w���m�{�ߖ�0���&;V�t)uD�qˤ�߈x�{�qg�P��
��k�^�j`�U�Q{TM_M�N�[��s�A���4���.(�|$yU`�[1,w��/�oY��Xc���VH.y�u�~��XA~q��!~V��On*�Zl��~kg��X:FDᙶ�J��5/��ly�v�� ̳��@��=�:X8?F:0�Ⱦ���$�j�Ë�Bm��=��w�_ͻ�$(��*yv^�˗3Sު��%�����q��
,t�L�fe*��1�?�}��)W
�#��|+����a��8y��2��.��|"�D6O�l�c�]m��y#�p�7q����2��}���ճ��D6Ts�1Oo6Y������q{xP�ԃ�nvΔl-�c�I�o`pEҮ��@q_�OI%F����v[õ��Ą�]b!%��Jr�G�ޙ�Fl�N�H�����6ࢧHI�_��]�~���U+�&�r��4�Q���5�a���Ԭh�/�C�ӼAg3�f^ݺ� ������9����i���*�v�ob(�
)�ڏ/��BT�'�{
�.NG���F��+��pp=��R�\6[%�s�a]�\��T�p�y�(݊��i�f{ ��xBʖ�ޡ�3���#����b߶�-�t��k��Jv��-JDa�Ag4az�>x '���T����E��ʯ1B)�����V/$�F�ܘ7��b�c����3=�̡�0Y�TX����_�0�K=���]º�a|ɠ�,1���oF@�� 15����y�	(�l޸�z�	#a9�{���{��k�W�,OL|��2��D4��S��82��������}'��|�xVtgjw�WU�Ʊ�E��ُ|$>O�W��J�R?�üg�D���S�_<��yꓸ�m��/��U����iޟ.��U�Ov(���Ã!����k�ORX��
B���x�:��dRDC_����!�lT�e��Z�:>e��A��-��oZ<�)�]\�:�b;��a��ȇ��%U�6,̈́��[��J�L��\��ዷ�=2�������s��(��m���۲ŋm��=b<a�z@ⴇ����\��牠 ���:��rޅ%eO��P\Ӵ���oV5aZ�L �[���Յ�ﰷi1�2�t���ߚ>���f��n�u���Čl�3~(��X�\�i�M(v�Y��ڃ��
,��S�mJ�/a%N��&ir ��l�����aWJ�}%C�{q�S��qlk�=קȐ��2;pI��DV*4��+���<�H�5w�����n��S��E¥ k15>�©b<�5*|��QF5|����Z	/��ue!� 4��r���c���:M�����^�is�wl��wA}�yN��&h˅ǿ���xM3g�Ey8��:\���"��§�}jM�Oap��'�����&`�G���1��&�3Y�}g6�݅;��O��?�%A�7��'
6�`�34� H���f��ڱl�`�T)T��Nq뼟��N'ƥ���]1��O�j�ȲZ��.[�\�&�E�/��=_��t�v,��tȳו&����yk��_�E^��:��̐��$p�E���"�5ʂ���iAr���c�m��ú�c<[&=����22Y�e�3��`�ST����[���
	wӔ2V��f��P�&)2=����;�6�k����A���}vNF ���(�~��Q���F,;�>�LxrTp��O��-ՙٜ΁O69�7�A��̥�o\�E�"�K!��>�G(k_�T�0}�5XM�B��u���e�H�����_��@�.O_!d;�P���@�J�l;S��L�!��N�>�,���Q|���=�I��6�[1���u�_yߒ�B̺�-�Q�Eop����$��K߆���]!EY\.ע���en�I�FzMj%�4@��o*G�����ds~8�*���������V�kD��o)2-ws���͟F�xC�E�%�q0ۂE� �e�2����ʓ5N)�٨���_����ME��yn����������UU�h��`E<�#ی��ڲ�9�Z�S��%똇��:m�2}x�Y��#Uw"b�U��v��'3 S<��b���/,��,i���iޝ.���&=Mr���,&}����=��;{�c�޴����0kh0�7��ajt��ml2z��ٽ��ܮ�p;H1�;������@�C[�etU�D�ceOa�+�4B�X��l�0���7�>%��M�G.�%�r��Xj��~ ��sq��Э��S(ph�K����s�*�����A]\�|V$ܓ�����CBd�2B(����>"Z� S��֍�35�ș�L�C��Ϡ��5�mE>f�-$V��pE��A�3��<�8U�tX�	[~ё�&d����k+�,1�&���mn���-r��Z�;�A�\�B�|h(�r�t?L ������L4pˡ_�lEc�<g'rںc��|G*Ľל��I���������#$���;]�x����h��/��@˶��M%��֖���5}K��=�4'yش���o�!���Wze�,9찹���_�3�AG��p�mg�&)���#���d{P8�B���d=�� �*��E������,��X��U���֬������8�� �H��z�@�Lӯ��2ѽ��9���W�`�ÑR�hB'���Rky�#���>A5�tW6�#�y^;�(��P[*$���(�Q�5���TS�����d�.)��ą��ܞ��+d6���x��O*A�����g�at��k��z�Ԉt:����O}s� ����j�~�,&���)�T��L X�VO�g�4%�򏢙M|���{�$�f��>�%&V5�t�R�:epb⣈��Z��_M�9�Jۃ{I���e#�"�� D�ܛ��wB6��.�mm�\����?%�H�zlTk����t^��aB��0��	e�����d1����j-O����.mo�R�v���.�b�&I���,#��'Q�թ9A
#o���/��gE��O@�����'�R���Ǫt�q����]�S���V1�<Z{�T�������IZrgV�ʩڠɒ+G�cͨy�\�{�|D9Ѭ�p*mК2�eQ��o��3��=��5��N�sC��� B(��Y���ॐ�8=��rD�
�����C��"���з��oj��| ���~��0��'ٹ����C}�.�O��*�I�~����s�.�5�6��W��c�Vﲨ|��:�T���$�����e<@����DDD�xw��k�ꎙ����'o�^���{��G���kJC�����BҎ@w�\r�5�5H#>?M��,B�&O�OjW��	�����	)�!��
��E0� QL���&���u��t�q�q%��1���We�K�x-|��L�:��������,���Y�ў���z:f��s3#������Io�lz���l*�T�>�����q�����/a��JϋH�ALsw�!sc�L9ϣw>�=����@=%왽�����8gy�����*��D���e3:��E�x�z���Vp��j?
������h��\�o��~ݳ�3�4!g�>�� Y׊��/�ѳZs\��џ�a_lP���V���"�x!��䶦���0⛍١>�W�[�_%�	R'�b���)����һ��X���q"k���D�'�����#��$��J�'�!�[(KADU�\��0:��=�gٶF����n�y�׽����SO���n��G�s~?�������p���.&`�)7�@{���h��@����\��	��7"����?i4eIލؽZ:��F{���	3�'>5�� �4.�'�w"�*S������g�[��\>9����5*ȷ&�zH���'֦�wO�O���
K{ǽ�T⁤_T��6p�K��x4´~�ݢ E���@��@��(̰8�}��V�1崶`2/&I�f�ǈQ<�@�>C�*��Y���\O�'�3��u�������H��ٸ\!���H�b��v��&�5pU��
g���-��S�c:�����F���u|���y�����ɭ���Y�П)3���@�dik���8٬<u~���#��?l�4�ё����j��(<���q"�/;P�n=K�2���Z;��jiaoT�oFV���d������a��1�!E̓$x(��i�N9eb�+B]K�$�AAן*,Z/�rI��{}Jr[��W3�f/vH�\�<��f)������{� �[��p��^o�e��'�(�k��;�Lli��+���|�
x�T�L���F�A�'�U��;�:������i�jC���������ߕ���Op:)����Z�.}ܐ�)�`�:��ο��EeJ��K�}��Hm�0�4���<^���m%\O�)3o@vvԊDc[!��HU~�J�^�������W��
�ɵ�u��9��՞�u���Cv1vfu��`B��_�ZUt%�P4Y�i y�d��h�+�	UҾ�.�1�M����O�� ��{���g���4�6����O= �}�a$|q�I��H��޼o�ɿ���*�2�u����`N����U䧤�Zb#�c�'���`D�c`_N�:f�ћ��.��J�����:�j5!Gob"��H_�̊`�� �gw5�kP�9�y�Z��R���3J�Œ�|��L!fKcւ��`>C��Ck�n#c�$��3��|�������q���q�-��E���(�H��\ �f4y�nU��A��������$�;u(Җ�g�κD�dt[��2S���I��0ƨ�10G��f�>B:u鮓L������m�Q�p�\Z���J@ܗ㮨��=���w�hB��9�l�RZSV�5
���v���0:ٱ4��;Yu;�ZEg;���賴r��.?�Mm��@]�#$�*��<�oee�_�.-�U^܀�Y�޴�U'π�jQ��lSyv(B]����Vn�[&�e�M���Pi&ہ,���s�o��l͝Z]�A�4�]6�1�A�X��*�{�����ٍ�1X����~»�Q�
0����G��H�T��CB�8�b�ؐ	9e|8	cv�TJSz��_	@s@ �;?]�oa)�o77�2
�0���]��q��el��_S�MW���ܨ��:���U#��;KaQ�ZI�qb����
S���K�!Ι Us�֚_3=��.�\�)�@x��\��)����