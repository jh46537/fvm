��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħa�gU�]@)},����ע�>S�H����O��QK�\�� � ���ݡ\�t5"��£]�x����b�����{������� t���g/�%Vz��'%麂�����`�t�!���|�Ɍ+D�i��Hȝ���<�h!׹���̨�S����u r �N�G?�v�~U�0�*?AfOtQoweΈ��;��Z�K��Q3u HE�wٖ6=i}^�u�%-�d��T.����I�MBM� Y��W ����;�����a7�,S���cIْ;yP��.B�R��!���R�f�痢��BlZh�w�ƾ�ݾ��iV�}ꝏ�cc��c+G��?'[r2���w�4P�*�lO�>����&`U��p`���-�8���I�{�s[p�(��<*kf��^=�}P*����j���ÙiU���.	�H^��:���b�U�v�[�/�N�0��}��Ŭ�$�78׍���+�L���W-a<�T ��Z#�W��c^v�p˨��z���b&(B:Ja�"�Ȱ5`$�5��NУ�%���=�:g�k�އ�����P�3��@N��1�z�?�����X�4�V�8�Α�AW�����':~qie��uio�F/��u<N]��g�����*�Eh��Yǆ��3�bӏ�I1���Ë��,c�F6�b�8�#�������"�d���h��BC�����;.=�O��rvl_��*1Ę'Ay������๲U��I�"�1ֽBtX��r������H&��U��.�ZLGN{�R�%/?���� D��6�8{[�׹%��A�z����b�T%���,���J��j�aA���fZ�l��/,�ɰz��^Z��{$����nq��RR*��O��@.�r4��ч�B9�"$]���f��	<���vtU �֎c�i��j�AF�8	�fSZ�&�Mg���f�[a�~8g�:ɇ�= 4\�'r��_�D}t�]j��x*�y�=�>�aJ2#hg��ꅭ(uo��-:��j ���l(l������Hz��+�O��/���F
RQvv
�*�M����+F� ���u��ɻ�U�BBev��Fͫ��9#i�̌��V��A�d�_֣�>hf� ��_�g����3�s���	�ӿP#n�k�h�8����7������z�^�����Alq�a~��� �?drt�o�V��H3��v�/�X���r>�>^Ԥ���BJd�����<�����@@��Q������#8�E�2J�9����ͭ���A*���&� �,K/ȅ��>�J�$O����-3��75�m�|�������"lR�T�uhGp�B�: N�$l�2e���:���Ԯ��>�Kyb���+}Sc&~w{��e\^�\(��F��˭�6��k`P ��j1��u�̜���UEw�<�����t�[\2*9 ������n��=�O�`��*��7��:�u��c!��"��bZ-> �����0�f��&wi��ߎ�g�:BP���p�u�2D��5�����u{��aD�dN�]0����ޒ����zG�GI5�=@A)�=2�s���0 _�)�rP+��V�A�\��l��dm8�s�B������@����B�@ Oϔ��_Ԁ�E�P�����A���rb�ͫ���a������H��{fd���l!e ��9M�]/r��.yce��Z����"�P�$��}����s�ؑ��"��E����iz��� �4xqk�;iˠŹ�f�t����3�� ]7�ܠ�/�+�ڴ���+�:]G+$�؏����	x&W�6s�r&�<s9��1|t�=��NK�Fj�7s�Z.+X�X��=%W�H��;xo��E@����!��I�cc\��۹Fb�5L�ڢ�=У^N�;�Z���|��!��Tv[��=�l(�p՟	�8�(�����/���ߌI�X)\��?9��?���X�8��@w��	�F�\�߈�0$�NW��p'�/u1����=C%Wǜ=���O���>�1�,���f�]1��)D�;�h.�{�� ���j;��c��}����H�D����lj3�Z��Y�}�v�.	u�i��qlZ�+<Dc��6����i2��r���	�z*8NJ�֡g��-�YB��]�-�c����C1srW5�U?4��fT٠��i����
�AЈ�a��=&�e� ���rL����4s�؄;v�"��	6�uZ��_�}��4��E'���������lgڤ�&Y��r�Շ�=�q6ù�]�q#�6�N��n��zVME��i(�M0��=ne����7{G��eKZ�7��M�5[�D
�c�� �q��mc��]� ���C%�X}���2���̸L��-������Z+���CL�3HͶ�2�H�%!���yȵOC{����૴� �������U쐒c!-"�@�Y��f��x�f�6�P�߇���\%�Uu4a�Ê�=��t�a�b
�x�dn\9��$�$)ޤ�՚;fDRwt���� 駋���3/a��*'��(&h.֥�j����Y�s;q`�N�F��N߯=B���q
����pʱ��r���Z�i{`�#�s�����tF !8�bBKe���bq3��!t�ټ&��h�>�hW����(�U���pU�����v�Q�Z5��&��vl�Z�*h�oU}U��^d�/����@�c��*FeB@,a�ՐS�c�H1����7�Y���6����K���%�Š-~�B�Y,�`r���ҒQC�|@�qkG�H�E��5S��Qk�2h��Lk�������KkXX�j��~�GT��U��5*=��c�ޥd�1�!�H�U��,e��R�Hd���KD¹B��±�e|j{m����XUt��AP���I�<��yø�����[�i��9H��Y�ۉkzy<O̝_�#���
��ql�jH�S�ˀ]?7S��^֨�<ξ�q��V�LZ��-`��ٔ=�CI��a��b�6X���Bsf�7
�9���?�n��T�7;��e�h�N��K��f�{��a�� F���ɕZ���y�wȫt���z�h�G��������ƶ��c_k@�^��$��5�<�_� חu��E��D�"��G� ���-X�����l�?b�&-�!�4����F�$����^���]׽NT�|�z ������p�c"%1*kn����f\\ds`�K,C�-��V��� ���m�h9�$#0�݅���n �n����+8ro��J��p��j4ߑ���ɥ�E(?��΄F�:ܹ�e�j��W���1�=I�x%�{���/@B��̓��)�eZ-M�2Þ������5s�z����0�u߯�;x�}���m]���;	+�]Y��)wJ���Io���s�L������W�U�����C�W�,�h�&k��R��jwB�7R��F�x���\CTS[/�/w��m^�`��+J�~���R�i�\�%}���e�b05p�-����e��8Q�M�p�~5A���h��z�����(R��Z�-�`H�!�^N6Q��?-�Ή���e����`}�!�N;�UzP"�s��ֆ0-o��# ��2طΑ�չl�N�Sͣ���ZЏ�:['>�Fԟ�QlK��k����
�*Q&A�xx��d��*�0t �����#���t�0?(o������jDY�Fe�
�H��t0��?�w����W�*�����yݫT��S���*I�z�<	�MS|�W[�9����%�t܏��Z��Xa{5��fY���w�`L�:�® @�{�.w�#>%#�X$��K�:in�L'q�����<��	�Lz����z�y�X�������Ύ�ʂF�>]#�v�b̬��طy��dޜ۽����:��T��;�|�4�fE*Ey��g����$��\r�\���0�FTguy�bZA?3�AE@��Qys�	B���ҫ&��-nϭ�o�y�-`�:*~<�U��|�	UfJ��c|��r�Q�8��0;�њ���_>j�V�4^�`\���]��P�{��O��%M��u�5��ܻ�^�+�)1x7�<�l�S�e�e����w	�W�̋ͨ��D���9�Vr�_�wvѽ�s�mf�+��<a��T\�۠W�^ZSG�Y带�ٯA��O�}�8��f8�#�q�@bc��vW���<�!����	�{)j�&r+��OcGט8�Eס4����3 ��"��(#昞��=�K1(O|Ә_Kc�K��4O%^��.%�af BG���1�٠�ʽ���gm���M�K�N(�J�s��(�Z���	�ـv!3[�C���v���j���Aڮ����@ �vR��̈3����_9f\wH���R'i�;�y�y���ѝ�c�˯z�*�r�~����aF��X���+�1=&5���%��+���C����u�4~�@��3RF����/��>�h��}t�`��V��?��U`}V2 ���Y�Y�H`P4�zn��ڝ��,���v8�(d͆o]l�w�$��ܽw_X��h(�*�s��jG�����ɤ�kG/L��Aw�:U���K��T��Ġ����Aa1�Np8����ץ���eݖ��;��A���X�K�v0~���X���((���R���X�t*f�YO	�1�\t�5��p����Zi������6��|��[����Y�oR8�W<)��.�4�h�}'N�]@48ѭ�Dj)�l�1+��݊���-�P�~��w0��AT� ��D٫�Df��rw2:���I@��k�n����/�I��-��x�c�0�cy7����}4��ڨ&;����q�P��'���~׳��BN�5l�}w���|�nDH�<䱶q>��y��7k5{R��&��Xì����(�IWD�6����`���d���=[�ͯ�ߌK*.����)0�;�l{�r�'��+
�K=0���8l�.X��?P	��ܥ#U��AVL�b��#�
[Euz����Q���Π�0A����vG%2�%�����Qd���5�dzg`�$��GL��g����w���B��0[eM}�5j��S���jm&��rURˊ��������6�u`���Q�b�L�����1�4�f�4^
�j
�0�/���	���Ͼ���x�\<�Z�+Gqku�	
�#T2���(�z�M\1������͝��C��t��U�y�*%��f�	u��2��>��͚4�2 �2�lkm��~�f�s1�t��@���?�)}�uy�Q��Yy����9ese�* �����(L���,'z�_�a�����;B��A��r�W��i��n��j~����59���Y	nx�== ��s��vN��N��Rِ���v�T�!�]E��v3T�%R�w�QH$���)5��N/	��&�q����ގ��K�
��#���	a(��b>G�����]�HFdUܩ��^$W��4.%���1�N1V�
X�*�(�+1�%�d_��"���1Z�_�X��^�h7@T��~��`��%��H&o)�ZH��
C�e#Ǻ��N�d9��_rpY�=$].VV�w��30�{��>���Ͳ�W�)�N v�S��;U��29^T8yjL�"���VN����v��+)��N����$��(	�� ���'H��	�J��=w���K�$yAx#��J?�x A��&�)�I�S�'�2�Δ15�g��Sj/����/�ʅ3��_t�u�?�B�`\<\Ɯs�;���\���L�E��F����W�g.�?��.�+P�;�.T$���E�b���5V��[c����tL;��GA��Y�;�Ǩ:�?C����H���Ը��n���?��Hm�C���jw��`-b
BaJ��L/,��A��`й9��d{'���ew[[�w�,8^��o���J�8@9�]�#�Fղ���w��,�B�Lm R��E�`!���y"gҕ��X�Ȝ�*j�CQ*��I���'��8F
��^�\*����wU(g�"��S~2,RՕ��������'�3.'�\h��h����B�:Oۭ�9u�@�:3|��n��1|�  �]g����@I�k���.K���p��z�)�����V�1��z��hzʰj��d�f�{�;)�J��p��4�.ii��d��������m�u�a_:�=b"`/5:���mdZ�u��h�(���*�#�.j��DO�m�4<G��t�L[�LRu��i�q���,_�hC����P��+U�1~ɪ�ߡV��ҿz7�����"��<#��1U$�b�ik��ч��@�;&��5�;������@�H�n���p�Z�!d,�U�w���S�ߟ�|;�f� ^j?^�+"85��s���Ew����V�y��`� �i1����M�ח{)�{��9���գ�ǯ�/���g�3�K�a�����t�кf/�|3	�։��	T>���h�. ^V�D���ӄ�ٴ.�1���CU����X� �n��������>��9`�DmK�3h��'l���k��I��0{�q��%�n8����Ř��UɄY�����8�5h�����+q>6�3�ߍ��cy����ʎ:��I�u���y��֫>�Q1A�t�yOR��`�#m2Eo��V4�1�/�ߞcm^b�=5gd|9�ᝅ�� ��c�_���,tž03����)�_������%�{/�@Rϻ�gyu#7�s����M��^�;M�!T;_��y�jh��F0(��]S��5E �&������ӦN
�Gǽf�o��.{��m:�$aTf>��jG���1o�n�~[�H����_'�9�S�>��~��կ�l���m��<5�&gz"��-�B��uٻ�e��O�~$.���o#�X���=��h���6M��WJ�O� �#9Q��4N�@K�B�gqT����7y�Cz�9������w��,!SE�_29�����a�ݍ�޸x����K��)v�R��U!��O����^
\�*�X;O��v¬sm��Sh]��=���=c�]�	4�����P���w?��D�ʐ'�w�(ܨ��fe~��S��Ѩ	[E�����m��ko�BB��z����qa���sU{�����l�û�]�D�D�L��P�=���>�QsҸ�޵�w2�Ɏ����gq�O��[y+t*��-V���O0��5G�<�r��'�4��)-��k�WS"�:�ѠI���K�m 
/><�xA]x��f!�Zp���qD�'�i��ȸ���6�RM�������x��eHN=�x�H���}CS\Ne�����
��O��x�q�bsn4M����o�j���N+m��j��r�V��<<��%_	��\eO؛�g���I�DgE@ʈM�>�>��o^���@�
5���w�,�v@��6S93&"�9�PbD6����D��+�߹��!!<���J`ʩ��(S|���X�3�+�2&�C���k�]pτ9$��J�T_�>�89�#I����:���#A�ا��S�X��?KqF�a0Ϝꁺi�rU/�Sa��Il���q)�;�����x>�e @0���¡��xch,h-ݪ@������M �*~d}Qu�S���~���?�Z=e��u�����VN�o*����q�>j�	�{�/Ȣ����__�;����~5Y��[׭����L���H1�1C�ĥL�!K��'����{�����w�CpoC��Qn5�������F���6�ཐ;����A'�F����s\x�n�5�Iwg��i��5�,mpu��Z
\B;���oDLDF�U�����lwXɯn5ˡ�m��^����p�ˢ��U�jQF��-U��_���ĴK_��N���o�㍹:�F��4���@�	L���ܤ�8��$��+j��Y^� :̷��ż �c���x�k�z�޻���ߟ�t~�,�����N�L��Ŝ! ���sah�dG�}����:+�0���O�}����m s�V,��Ls0� H�7�+}��$w:�a�;�F��PH�Cfk�y2��Xj·w���ebY]�|r+��=H<nj���miL����q^�����6��@)&B�LD��UO��;"�3�cJ�'Z�� ^��Dr�HJn�0
%�c�?[LBh�]�t��\z���G�0���Km*���~&�b%�a>�� 
,���o����qC�~�G�x�hbX���E>4���c�-T� �/��M*I�'�u���	��'�/�6d!�x���l���F��k{�^H��)OI����zM��%k���9��Y7N칸��UsR��đuM�ni9�?�d0�,S+)�_r)>����P�AY��fM���glF�
�[�Y�ڸP�+�	�q�^&\7?J�E ��C�Ҙ�]fo4��<M��&N��F#���[�J����z�+R�젛��L��&M�~�1�;6�5���pwTf�w�Km)���J;��J�su N�	+/熤�C���|���;aO�ӣ'Gd%���\��)�J���M�W�Y�a��Kܳ~S�'3Uʂ�:+@\VVH%��/�)Ԗ�^�lj�>���q=��Ơ��D��3�qb�T5�F��Ԫ��ϴ �/a'���V�����
B�ǡTb)���K��\��� �|���$��I����ϫ�Ss��m\�m<$��(雮dG���T/Z�����bJ���x`��?A���O&H��0�m䁢,o��Fn�~#�e�`���V8�E=E�/���jG
��;��KyV }�p��t����s9@au��*݇;a��V�qe${������ޯh�q�?<^>CJ�G#�k�'h��-�ZY����H��`[��)�[viI��?%�3񌅽K���j�̬�V��k{�4�Ǫ3�x~:�Y$����.�_�_	������jC���F�W�2���Ϭ@�;d��#��v
��&ډ����c���뿈�*�z!E��5�v�4e��嫳�lu�86���/_/]ŏ�������r�y�.��&�-�������Б?���Æ�A�r0��➂���YP����_��m�D8�o~�j���d{\:VT�xu�o�/>HΏ��3�q�����9�R��}V)"�	����k��BV�,m���=�YQ��k���.M$n��z��7�+|M+* �� ۺ��-�ed�/=%����8"��FŚ@:����m�AU��
W�A��V�W~�{k	�|���kID��tY�F�����%0M�z���Z�ˌ���4�ֻ���eɏ�k�(�q�-KyO���-��q��Ղ���?n�Qv^��i�r���ޔ,� ��xZ?��OE�ߦ���GQ~�"78}�+_m,�'����P�u|����Y�:���E�X���2��F�Lk�I�R��̙h��]������:W�a��J�~f-��d6t��5Ο��t�_t⎇���K�	e���1�,��5����Uf�Ps��*���`S��P�-13�2���G:�h�r�������O��6�:x�Ub�:�a�5G��˹Ov�l0g� r Z�2(Lӎˁ���m ޻����F7��C����9�E7}�sY��|��+���l�1Sa�O��M��������H�����$8���}��ƭx-��}�2ВL}u����p��n*�<OL�Μ�������m���'�i�4]Zt�,���@R���<-��q�D��`x4�7R�_�}A4��� ���
���=*^d�4G��^�[��ஸ�t�T���Š�
���E���x�Y0�Ö/,ՀFu>�d�W����ho0�ɨ4C ���D��:�V� �\�q�J\�ȤG�:B��P`��rh<טC�zBA�ʵ&����Q^�	N�'
@뾂dn�+�֝o�47�6�9
Dy���ųA�M;�i��B%��^-�;��R�!��U_���gyC����h�4��j���x�Y�X�
�������¡ްqȢ�}���O���<tT��s&���� ÐPO�\Z��G^�^�����*T-G�VM�� qB���姘Ić�>�r�O��m�_���As��\�����3���2w�����V'��l<�O��Q���ˣ��U�
/ÿ�C?��͋�K�U�x�9�<w�1�!��
�/~�b5�Č�F'��d���=K�r���,�U_`j��y��a�������lN$�V�:O8���ry$G=T;�gU��h8q���<��!�[t#�}J�����'ǂׁi����O6�2�������Q(\+�{����������N��r�f�Zu��"�}{�ӉR�D�\��G,� ��H䗼Su��2~�b�w���&����F'/:���5X�T�5�ݡI��h��F-�lf�å�[�1&��=X5]�ٻ�r�e�uv����$�-A	����@�@&