��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>����R�JS�d��h�uj;����Y�\9���̠�#_�^U�?�*�L�H^�I���q√��vM�
�f`%*��7"Ї�kW/�Yɝn2�.@/��1&h`�H������۲l���0����7����F����mu;��|O1����o�E;�������0�3k�>�Ra�GȮF����T�yW�(痡"�����^��`�*��h���v���$���y�h����ơI>���cW����F)���wG)Gތ{0Y�r��~�E��u �a�����r�-"�z��=���+l���F�]��U��(�v�b�j����1X1k��.�@���[���b�
3��OW��V4��|4ZR�M�OoCW@���L�#��DL��Fj��Q�`_�u薞p����s6�d��Ta*1���$M�-���{aE_W��t�#ՀMb�#�qؼe��c��1�7�,��p����
Ѹh�pĻ��8���Gz��O�m���-�X�n�WA.�|�_�:Aw$���]z��GH��힦	E���I�Ǎ�Z��z�@o��P��P�yz/��sd�L�ġ��n=�N�ݯ���QT�ţ�U�GB�J��P�;3L縟W~�w�M3*Ui�c���-���@f0H�$F͢^�.���k�cH�
�TӜ~�]�j��a9���_Vŭ���$��&�MĖ�*��j����/�_
�qm���{�d��-3��xO�j�&\��BRTT��0&�0�]Pe��&���QѤ)}6j׾�M�������D-���m2�z�V"��&�Jc�:|�h'^�C��n
��xJ<zʽQ��mG��uY��ՁΆY�J�l���0Pc�}~s���;��%�U����{� u������=���zW N ��.Q�4�K�P�����Z���ݼ�!��W7��Qimvag�������lt�	m�㋖�/=���[J鬁aD6��&&����r
��!�&Y�N�l��'��q!Q�䌹WA�S��=��h��~w�Y�1���_�#
�S�mŀ�����������}�:
y��c�����H5=KM�f�4=g$�Y�'5Nl�{B��	8x�?�4u���r�t���P�@|FU�:�r��������G��Fxt�G����|��Tȕ<@�~v}\6+
��:�J)%���l_�[��MO5i�G�0��"u�(�m�@��؇W�J�|�t�����B����݄p���sQ)�rF��H���B�)d�P!�H��NU*'{�N~1�WĤ���Kh4aS�W����f�d�P�͂vd�PS��Eˡ;�أA��G�c�W������E��-rM(ȓ5�M2f�f^�a���Ph>xSb7x���:�xl���S_G�H�z�#�ջ�b����%��B�'%G�U�|�jC��$A�;A�v����z��O���B�+����E�J[:�M9Qbg+Է/Rv�~��nt��	�`(�G���e�#ͯ�X��H�9R���)�?q�)�6#�,�-^��x#T��ǣ�S"�+H��0���d���%�S�hh+W���곃���#��|�Q\�2�ȥ,��t��_�9Z�B㊵aNwI���c�σ�Sl�->�skVD={͊��L��'�Z'w��bq|Z���%��8
��0� ى:��o%����$� 
�\�������HFԶ=�D>�m���&�+����N�C�	p S���~�uX7�1X< �Ɉ�Y�u]ŝ���B	fΙg�00S�[���+8j]_\z`���!�.f���|���횂����i�����!"����8�z�ၣF�T���|�e�#��v�c\8�Bc�À�"�鋔o�KQ-0�I���cŀ;	�:��躭Rlz1�"� �B�̌�e|���%���!�ż8H���u�Y�h��o8G(��+�~L�F��E4ka\�IA]�g<�NTF���4�￙�b���l�\�L��(�s�[�� $o	l��W��J�(������qg,j7|��A�H�j�\ϵc���`��O8*k�'a��u"��8t�K�F\����N�2�0��#<�|d���vn��荁�7Ʀ�ߠS�)3�6~�	�Ȗ��F�?jU[��sm�\�6~����{ѧQ��n�ІZ��bw.\�_!0�V� ��ۀ/bd�@�~��f�uPnK?$9Z����X͚��4�L-���	�/�d�$=���8>�3��P�v���$6�}�0.�,���)����ӣ�>�Ʒ-�8aQAG����HHՠ��뫄�O�>LF/�]�m�pکf��1�p=!v����ED�9A�R�u0�̚��r�Q3l�.�^$���9l�!uƳy�х�Xpm'=��/���)��X��c�a��ze��,f��7�I�8s�"�v����U>tn���eg
t]A��sƇ��[t��I�!¬�o_��yȄ^�A��[	S��&���glSӁY}�&x����d�m���z
g����L��r8�Sؖ2 "co�Ų�� N���cX�fbͻ(D!{�*Β��hg�!����2.�t1S\:A�Q;&O7-�_��L	-�~������42bc	rdr��Y�M#2�hm:M�ӟ�y���Jإ�T����J0a+5f)&��G�_!��k~�y`�L���*�c$q-22�
��e���a����,|N1kI�>�!v�cP}7����p�!s�Ͷ���Gk��������&*�>1jч�fkx/J86=�J{�����q��u�a��ݞ�&��vƌģ��C�1��8\Z����z�5�	}�����A�.��b�WqC�f=�V� �,@ҋ�lIx������Mh߹�O�U��������H�
�,��gU�3Z�˷,�Ƴ����){)(E������%��p�)5œ� "�:^���j����p���H��i��aa�6�v��e!;yY���\WK� �P(]�i�K��u��ݣyY����|�`O"��+r鲕�D+1/2�+&n�J��E�g)�L}��e�����G۸�(1`9��:b���P��2mVm�=̰J?~�:�l��ps���E�	�#G&�� �2�v�~�Q���Liɏ�a`2td�r�� �����|)�w�=ʚ�o�G&�QZ�L��o��{����dahieZ�+���7p�;�&����������Y�����eN��<�0�_;����'��*���by|��DD��\�>B[����3)����K}�Z�����P:#�S{� ��7yZ6�lL�z"�Tۄ�h)T�����؝�at���h�
��=.>z���>Q(֮7c���ߍdU�ι=�0����+�����;��)>S����Ĺ��H�J5�t�;$-gб�������5%�#�|�d�@m|$�p�L޼
b-��_�|��y01U�q�ܞGy�U�@];ZЬJ�cy��[KQҫ���v�u!J�|_2�ũ��r�/�y���p�S�q�ú�0���0Z�W'X��R�D�j�8�?�7Z	-��=*j����0l�cc��lFu1>��1'�̙K���M�����^o��9r'��IՁ�HE���S����>p��d�IQ���3���_�<R�,ZN���ց�C�#�L���Y�t�_y��z����TviM�/gh��S�P_�X�ٌ.�Knތ��QP��P�2.�Hu#W.�1��'j�ǖ��䡫��%�k;q :�cֈ6s��x��_"T�w���O�ľ���/�m,����O,h��h�H$�'�x򔐈/��V�ì��/�J̴����w]^q�077��t���y�:�������(A� c����W��sD���Ë��෾��'��BL.��q� 2�95�d������B(�H�;��FJ�C����i\����`��p��P���b�$�?���
#�x�4�� lr�O|	E٫1�eN�Og���k "����}�^�4�.5kH%�R̹
:Q�9uZ�>�>��YL�5�D��b���*�7�+�N�l�Z�\w��p+�ju~)�fҨ%�5�7��V]��i��� �ƪ&�Z�g�9���)������*�5�"�n�.�L��hl���#����J�u���Nڷ���1m��<�=/|�%o�-���J|\�p�ڜa�(i`���Y�e^G�֨��&r�Jd�߲֮�*v}�}��	��Fǁ�n_/����5�eQ	���W�1�ƭ*�W{=_H	C��ѭ�:)�oD�DU��DK1�[���H�	�D[��!�̋��(L��IY�	�Pz� v��a3|�v��͌@?c��t� V ���q 4�c<;�e�T�c^pT�>\��(����ڦ�� �H��1�@��˘���Xdi��f`�����?+C�ϛ���wg+n1�ȆŜ�;W��
�����d������[��y��j؂� �eWd9�'�bֹ���.vfl�L�:� �l���!����Je�����ɭ��3��FX����Y��q|�^!VA+�:����IV|�̕�����3+���������0����]����}u�FrFq�^���^X��\-̱���:�?v1@\��'��f�h$��'��r��K��[H&G�2k��t�A�z4|����Nc���CR{��\��	��S�27G��q�D
\�lj�{��uX�!�����N�W�U/�v
���"\3�CE�Ŵj?@Z�Ɓ̙=�Ž-��O�R��6�E�Hb�y��=/ح���x����Br��v���q���b0��Aܚ��ǍKg�L���Z":�.;�&}�x�,߿]�����N��:T�`��C��%x]ｚ�~*k�*�Z�4eJ��5��1[�yŰӮ��A�?\Y_l3�r�t��n�5}��,R�Qwn��zw�V2�z�u�H�u85��^��+{�EY�X�r�Gt"r��%v�+2;÷o�K՛����*���&m�k��q+:SQ��j�u�#�D�]OaẆ<6���ޝ�
���m♞p�	��Xv߆�GԿ7����Ev3���C�\^��V������v���y�S��W�j/A�-��
��n����Ɍ �Jw})%�a,23}&ϝ�#k-�g`YKa;��J��l_���#�]H�x/����chfLH�`Wp08�0'QՐ����%��Ɨӥ�H���R@��{�m��/,r�yƍ��$���]�^>RC��]��޽@C2����}*�J��80��/��P��8k���ľ�	�v�<��4n�aY|�脇skbL�/y%���P�%��"E�ߦ���y��:N�'�(��`���t�4m�0��
���Kqg�]tk��R���T��D����zp$?c��0Z'|h7�*xs,�r6�@lߙ�G����� �ؓ�����3�<{���D/��Tei���z���ݺ��M�+ ML�e���l"��NK���o(8H��x�R��t�z�I`���F�'���i�`N��'&�1�=~�*�4k�P���|Y�Wa�����K�Yц/��ȉ��$�Y0=ګv�&�q]��oT��x����AU6�EE��<'YŧO�yu�q���y��g��|��zb,Ѫ��poF��'���Pd(.Ă�eX�Ғ��]c�^F����O`����`�O�FƊ~reil���8�!�[��W͈�{$3�∮�Oq��<Q?z�U�wO%��w��K�c(T�����&�l��kO����j4�x�-�x�SbAD*;ݳ<��bٚYK����tf$Y�H �J�L�x¢M7;  �gh&��*Ƙ���m�6
;NShE�+=\)�������~��C�Wl�$:Y��m[A�<��0R�܄��1��n���D���
^C
_��Y&��m�_�Y����4i'J��7o��xYϦ��O���{~;���v���k��1_��������J�a�7����Չ�-�:�5��$cg�[q��k{T7�ɶ(��n5O���UhS/V�f��uY�����a��Sn/R'�[RZ�]��ȼA�b[��S�@��e��� ��:�
�>�E����b1�X�_:��Ko,��c
.-�d����+�Y��_1oGi�al՜:m�� ���¤,�J�lԞ# �ieߵF�)�Ց�A�5;~=ب����U l�k�����ΰ�~�[��n�����= Zh�ͺ�3ceu��T�P���F�^y�Obs�P����������ل6l�k8�W�.c����-z<@�Z���B������V�'x�B���u��-�gb�\� 6���;:���+��ƀ�Ӳ�����G��}X�(�ڒ�o��/-�Gz�M�l�,@�+�ߣ���p:�*N6wk:�d��>����Pf� z����F=��U�J�6V0Gr�Ȗ�+�1�&�%��w'��a냈\��@I��"�����?��Su(͆�����*�>��VR�i��k�
E)�b�ࢅ�QCl��_O�S��$���2�q:����#p]E���w�ML�/���[�� 7������3��k���R^Ŝת��Wt@���w���	e�73���ikUY�g��OQՃ�9��)�1�ĩ=#�,�]fhÛ�*�ס�;o(�L�R�xr����^�4y�����-�ΐ.�:A�HJ��
�׽�2t����u�at=#��2ŧ�f�@t{���Ēu��4�k�0�eܸuɇ���(�77&�kk=�KT� imQU��ϵ��8�l_�Z��ޠ|�qIb�-�T���
�d�.?߬/E���~�7�gr��U���B}�N����J.W����v�k�|������<�����`�^��YF߬��'52�z��H/n�/��=�/�%�zj�i�-h�| ��
OK�L/7<�xdq�f8`/5W8k�0KIr�#� ~{��Y�M��h#��gf�ȔY#�*U��}j�u�R@ԫ�r?�Oϙ0�n�����
T�w���`=�/�W�^�c��\��e�s�Q�S�����3�w�=+�D����|+8���q+�����<�PP���IS�K�j|�+�����D�%�~����t�W�(�˖��`�"5w�������dp0���\�Q�Fr?R'%q�G��Rר7��V�n�P}Q�D���b���.{��_^a3nve'.)�I��l�[���l����2�d�
81n�_ C�A�&�4�Ub��7#�����Ҥ9||��$���Pbkps6��ŋYГk����Ou��1=�ű�������r����ŉ�e1d��de��=�������S�F��3e�;g�#��e�Aьc>�B��K0~�a����4�ɓo3�ƬS��̴i̓����ќ��M�A<U��@X�g��H�ős0݆�Ȋm�����l��ˇ3&�Ơ��^�PK�T�j(��25u��������^�`J"��P�ރ*�E��}u��E�rT̥�BGl��;<P�@��I1�U��e!��\��� H�$OE��],m��%�����k�ä�`�;O͙��]l��|C$�K$�-������n���V)�F�8.��ϙ�����q�a���b�.0{�����pW�eZ+���V���b�8A���	U�9�ym�xm?��n�I���$�FϘ��Ƕ�`�+ ��^_�x�k�3�A��\�8^ǠӖ (��E�	�.��4�b���u	-��Y�WD>$�<�H�� |�F5����R����P����KGAv��DU8�����5���*��7�����O��ȿN��^��g 7�b����g�YaM<�5ۜg��/��:=����K�� ��t�t���CJv3�S5����XR{��y˵"Tg�itX�&�+������4��J��?���yl�����+Г����	�h{HF���w�gmP��]q��%8BqM��NeZ��2	�u��eqy�dZM*���n���=~��F��ܢ�*��Q�<�^&'s�.�V�O�gCL�\`�`m}������^lJ��`�������"��@��6�~Y��%طԭ�r��(�>޾�������z�,�����	�4ܜ�z52��XM*ܚ�$ �W������q�y����Hc���#w�D�ID��rH�1������ �� ddA���jρN뚽#舍����.懬�R����|���2YA�}s���A�;k�[éZh�!U�H�@�\i��D���N�Np���wň0����̹l�P'�j��^^���5��G�kH�!�/a�7�P{["�"�G� ����V�'S�2�-ɮniQ�Lf.0j�%�/y����:��+��Q8�;�!� ���Q�v��o��+�v��9� ��~� �r��?h�?=�o���S�{�2�i�h&��n܏����8��GG�q����i/R��j��3�RV
��1}4ip��)������EAEJ�τ2.,l�[�c�� F�TQM�iS	��g?)�^��[�G���_z�x5Z��0P����1� ����mF��@9}�|fúwX4Sʍ�Tk�
9�t� ^�'��i=��}�Q���s�uy?���N���l������\c�X���dY��c�2�����[�Ũo׊wTk!=٤b�$���$d��p�b���7ڊ�Z�(�X�n�7���HP��l���6�/f$8Y�g}���L�P���ߧ{��h����0|b*�:"��
gI>�9�1�<l�IJ�<�"X���c��rx�we�ɇ5f��0ר���)m����탞�o�	3l�!,��� ���UA�[��A)�@���oַ'���B�����Kv�&�ʻ�8fo��o���W*aO&)�2)��@5�d�3&Í��>�S�:�A_)���e���bΔ�����0t���H6�[V��1�m��	��;�"޼���yq���㍱:l�ɴh���m�E���b6I�
 �͢�O����'��M��Ol�q���n"H�Ȟˎ�v��s=f�k �a�rz�㠗���Yc�/甐iC[ӱS�c�[���Z���e���dYm(��2v
B[����>%�_g:�cQEv���+��h��@5�if���K�tž��j-m�\u0��6˵��$�q�����م�2I�`����ayq��,K����ZI�͍E��J˝�k.M��ק����=�B4�����d0�]�O��"]wj����>����e���j0���b</�e��*4�HAK5=�ӟ͵�)�8��E��/�Dc��@`u��-;�i7lXtIo���w u��f0�ub�`y_=�d�C�b �q+�%(��G��3=�q�X��U�B�@e����p]Л4�ck&+Ṽ\�0S���d��#W��W���ֱ�����+�3�Lq�[���8[���t����I|}�6�?��/~�!_��Ko�^�ڗ6�H5'i0q!t\��/��̚�=n7�r;vC�)��J_�\~�� :-/�;p4�v�a��ژ���ʐ�k։\�㤨#��ȥ=U�U��y�#}�������|LP���U��O�ZǶ�ac�8c�A�A��5�Ji�FI�	<Eh�m�Ք�E�z����N3(�d}�}R\.p�f�Y��6��"��\2��|B��t�<�V=4��J�4����Te�x��I|���Ĭ`Qh�m��оx)QP��}C�-��/�����p�[(4U��ԒLlt ����{�i:���`#������O��~�WN�q��g��9��;EF��gbӏ2�����"�g�*zh�7>\�oh�z��_�G>���/�ػab�k��G���M��1.b߮s�6��#�-r�H�X�}cWD̆��2���� $2�)'L���z�#+l,��z�=BJ B� ���n���� ��F#�|��}g7���i���yW(zU�y�~X��������(��i��Mh$�~�b�y.l�I�[4�q;,����1�И���$T�Z���T;,�gxEp�O?f��R�a]�d��K�q�=Gj����D���UF��1�>`�6��"0?B�p|�v����k�,ĭv��=�#=���9X��E����-5,��O+��Q��5���6�Xq[{\���Ϡ��s�c�խ���������[	"��~\������t�`Ӧ�OFs�o��}:��Y�<�:�7@�6O��P5)����D1�~p!*���YbL�d�&��5�������
�?������}�������Z��^��3U0fn�4��1��
�_�܆�An��|�E�U���U�fNy�TPa^���|Aj�FCm�8��'�1��d���x���h��X�,��C��Yd�t@f�b����1���O�Lscد���}#�مWVqA�UI3�}�y-�!���V��G��������u o!J�a��H�V����t[�a��z���B%�h�p΅IO����T�/���e*)��#�?<�Wg\?v4�6=L��u^j%,�g'�����&e�9$r+N�Ƿ�c��?�
��ƪ�n~ͱ
T�[�������!��, ���k6)��s�y�ۤg�7ݻ`;�Egs-)���Ŵ�'��T<Bb��~F�rQ���:~��,�K �Ъq�4dH�o��Qo�2���Z���Q��[Y��;����&��-U�
?���<���[���Y ����`��/c�����%+�,z��&\��^�*�#l���c��<^���)ry�'Gl��o#��q�V�]$��)�9-�p{ڧ�|�e�\�;-���{u)��pW⁢S:$��'��u����Uq���46�g㾯�u��0Xy@Ξ�KX�G���vy]�]�ϽBE�6�{�]�(d���f]{:���Z~:��[[&��%.H-��:�
]|�l�T���狀��f
��#Ћp~�}CcyA_�KE��ق/\�T%V�{��u�Q1{�1�e�%-��ͥW�I\�y��.hOV��X�?��Y��$�˵$�4@Z�{�|���a�o����/s����I�B-=~A@�M����a͍�:��`jc ��y.�S�<��Ka�\�C���FX� iP�( �MY^yQk�ի��d�0%z������K�~�����e.�#��lb��������UX���v(�	�P��q&\�U��f���k� �%'f�h`��\bbN7-�Ne����4©���� ��q���I�W̿�ʳV���)��^��d��V�0vkf�UH�0rD�%�%5�c�m5���x��Q��=��Os�j��Z&k�6�d��S)-5�E����y�pŋ"��y�\n�!�g�	�^�6����O�S+Ii5�)�:�0<�'���0=�G�����5A��P�B!HP!��!�@��f��;����S2�;Mw�/��c	�gW��vI"�40�0�̌�˳�gD��E^,�>�qS��]ъʹ�P}?�lWf����iUw���u匋���nM�h6^����R5���r��"���L4�6�lX�� i#�á	�3RF�da�!����A:\j#`ck(U"�I��/��/�aO��D����o>Y>z��?6�J1��$�����ݯ<Q�;o:����1�,~"�\�t>̑�HZH�q4ʢ�r����.hNb���2|սZ�����󅻖�6�Â���_0�U�U��W������ǰh���T��W���ޔ���� ��Y0A���~���k�����G��E�����,,&a�9O8�y�U̚�K���X�A?�f��̓�l���ֱ!��f!��ѡ�H��MK���Uѯ�@�'�ȗS'�3u����w*k�H��ͤْD��}~�����WI�r�E���b���s
�ef,�E��p�I2�y���}��=�ÉNv�G���ʻ`4y퀘���h�߁f;Db1�����P_f������R��W5O"ا�-��|󴙯����M�ع.[��H|;q�P���'��z���z	� ��h��I0���j��ɦ������:m�H˽1�<3-��� "i8��!O�GӜ��K�U�ߌ���;r����h��;x9���Ҭ_�f�ݨo �������K.b����$Ш�x�/�9ErR=��)=�Kܑ���B�k��f	�< C�	�������2�Z��J�h���{3��Ζ���*p4�D~5���YЁ��������K���#����t��]5@��>9,J#קּ�A���+Pi�@1�ǉ�`;׋�&�?/�f�Y�A�'�X;t��7Y��߸��J4����jT�����Ӧ^ʪt�y[up��
y{�|ЍBX\9`i�����o�R��Y�1~n:�����Kq�Q��x_S��K�T�����Su3����W�_X~(Wg��scU(��<�L)� �x�6t�^�y�y�߭�Nm���Kx�O�x�w�EW������ڔ#��}W��ӛ?W4���jYd�e��Z��sg�b�����K��)��
�\���rH�ֱ�a�E����I�8�4w�5�h8\g�Q�m+�mN�m�W��	/�������Q`�	��r�0��.��I	vQqs�O/�
�.>w�L
����2�G"�����kF��s�:�C!����ɖ�������ʛ�yMN`"��#R0pMгor�`���#��P�f�k>���V��O5�x爹L	�-�oQ sG6C[3���G��Y� l���{��R7��p�QO�t;EX]q����W@FC'��|1��2ǎ�X����5F8��2����s��g}��V�����a��d��}�e�]ʵt��	�O�Co|�B�� "@�a��m1�F�����=�s�;����1���
�prgCS�#x�s2��2QN�m`�86� ��k��� ���;�S��8_�̯�N3��*�❼���?I�Cݺ"�Fh�8�����5��
�I ��l�^��z�2��O�pN��=Ԉ&"�͗�(�B��u��O�-A,�E���ߺ+��<^�����D�p&�VW�_$&��W	�h��3�������6x�=j��n��)z��c�ޝ���{H���Nɕ4�}�k�kd�!��Oh��NC�b@_`�;�o�w��Ag�I&s��8f��M@Gc%|��,��.�r���p��	��ʋG�r�A��P�v�۝�R?g�Ӓ7*�NZ1����q�'�E����9��e����Xm�(A�.��)Kw�<�W�\���]Y��[�f6��#��J��Gx^i�Qg0먐���9��fZ�<�n�Yu<�㤼����9�,no
��E����s���kH�Ai��ɏ��y�ŝyt�� w�&|����8�ނ�
%��V�4�J���3(���/���m�J���}8�H�_瀕ӸAX���:�,���W�lI��k�Y.nobȩ�~	i�/�r[�j���������ޠ�<./+�gR��y�1��1���#���[���J�X�a_�q(D�V�~\)��� �@��0�<A��Q/W�tW���j'j�[^�Ƴ�Y)lB�*#�*�ne�#���:��Ʒ�Cs�*�=QD�����+�m��G�n�鴒�cD��j�w>R�>�fk��ep�1� ��M�0��c�m�l6�E{a�V�w�_�|k����$�[Y����w����v	W�m�K.�c�B���1�<�l4Ȗc�ٖ��gt�<RBLi�7�$����]��'Șo+�G2E���&,Rcq��q��s����}k�USN>�̿�Mb��|��%�z��ZI��޶F'�U���G�g乁+���yn�8?'�5�=��5�I�RhL���+0��X���(����L�(��i�ve�j�L>*���:����ɶ,��k0v�@��^��}"k�gNL�����|��[䄿��t�O�T�a���F��o�mp���A؅�q�������'M/*��t��L� G�-y����u����. ,�A�C���T�5�Ձ��mP6����N����{`#+��\�#�]( �'pM��
���v���ܯ&�P�>�߄��4���Ý��Z��ܤ5o����G8VG?u)�t��W�7��@l�=m;����6HI��@4y
^"����l?�ej�+\[ ��:�m~��K�S=�y�y�(g��M�]����S��� ;zC��X�Z��+~�O�aR:֙��ԯ����-��5�PH�d,D�E]����V�"Eo�L���<��,V�y�A��n{ w��������`����5f6�����w@����Q��7׿!���# ����@�X�#b�/<�������[7p�i[�%��ka:0]Hi�7 �3��~A�?�0�=a�ȋE�7�=s��aUHNȢ��<ȗ���C��}����K�dޡ2b�*z4т�نR��pVףM��c��� ܆����� � ��Q�j��>m���c�2;�2�R���y}\W�|UnB���a� I��J��ţ֋#�T�jj=I<�=܃#L�F�7�cĶ?���$\2�)�/p�М	��J&Z񒽊�Il�	���۸w��8�PN�ygM���0�������)_���$~�}�_y��hG��$ ��N;��͟�I{3����
���S�*%�<�T����b��!z��Y�ߵx��I�W*y�e�����=z|l�ۿ���#��RhQ�N�[2fM�����.�DތC��H�4��A�v�@����vѱW�~1?�M�[��8��!n}kw3	�Q��� �03���I������Y�\�|�Z�\{5��^�V p`��aZ2��hQal|�YRh�tM��_X��p۞/�p���-=`u�K"�nकuaP͟[��� Kz%�L�v6w���O��|r{db�) F�>Xψ��o��u�zi�En�ѰXH%;X��9�9���;U��ý��}&�<u!ͪ{?��[�T�����=���G,��X^��6#�8�X�k����|�άȁ��p)nT�D�`vlY�fha��Sl�Z2�NA�t����i�J(������ ���C�����IZ��U|oO�(��"�;�o9���T�<��������/@���q)�aFBi��sH]��o�~@��[�f��ֵ�t2+~�[�3�v�(����^�������x�Qɳy����H��?���΋,��m�@��8�;���.�s�z� �!��є��U�<P�#ӝ�/��	����![��詆ȍ�O4/I1���#\�6���{��e7�沱�B����ΐ�˷v49� ��h�M���]�X��zeD��U2b��G۷Z߻M���F+��Nʹz}�'�V��G��́o���o�b��5�tG��SsL gV㎧��V]6��A�Y��*�[�2r@P�qp�O�$Mp��o��ƍ��%�o���y} j�r����Yv�vF!¡�ۥ_��Ubo�c��mz1ʈ�8��][��#ps�-q���[!`�Oܧ�/�f�~�B@�"d\TϮ���\lU�G�mNR���k���j<۽T^�[�'N6��c���:L��������`������1�Ґ���~7��#�K[����3s#�;[L�N�P��B��Sh���M�j�zVƌG�ߪiB4s$3�k��"E�^���XE<��T>&�*�+�_ma�f@h|����}DJk�"	��}��� �K�� 7���ع�� ��+�I������}V�q!Ǐv͔(){��̜�{�lx4���e\��UB
�9{4Rq9R��Aa��gk�!|Ч�S����B�^?����d�I�iY��.���J���l�0$l�0W#���)�=��Ը��Wg2��Aދ�f���De8����fN�̶4��x����O�*���� (?�T����7I�q�%�/&Y�<ǀ�AS'�'(u��斅�z8�wja����+�w!����P��M�p�m@������Z����P$�D�u*N�x=�Er*�������+�.�N��������Y}��w�
���_u��G�/�#�od��B0�Md�R^�/ 5���V���@�y`R�p:��)���
�gO'�s2«?k�?)=�u�VW��ǅmK<�!@����'�!�����{��(*"�v�=���5�!8+t�l�E��ĈA��5(�0�v�4�r�2�
��6��y�7�y�,�}2��D������O�J8�g_�yA��tuwo�k �l���{��m��R��@5͸�:���3|�E��ź�Kf)=�,�R��_l�ډGίZ�s|�-?yY�%��Fͻ�&/,0�Y�S��a��Fd?��m���S�@��9p<���p>p�A�69�T�_d*0F��/�:�Ȍi�]7��ԙ����C��:|k����V�&v�Z�"t�$ߨ��)�)ޖBe40}%B�ی_�?���}�� ���R�t�rMyL��,��/���v�|��*�C8�D\Ge�=J��2q��4��\���	%zX���_����ҘXZ���*-�/A�C)Y��<���ծ�6�e�����$~3�r,ɟ�`�(/WJ
��ig�h�a�[�Q��ʦü��}a�>>/";D��k�CE��e�0uѥO\8}y���\�SLO�s�	e�m��jQ�5|��Ə)�``�&^,��kWC��]c�P������T���QW���^�:��I���_�.J-
95�qJ�e��]��G�&	��1��Ԁ���Niʮ�#����������.*dG޷n���@�.���"����V�ѵ{O�;`���~�7��{jz�,�bTό���zk��L�)y~ͮ�b�
�.Rȗ|�HV�*������N��W�;Ж"�~W��^��/S��(���>F5^�+'J�^+O���u	]ultI�:�<�J
^��/��a̧c��
�������YR�V��h�?��WD�ui%�w2�wW���eB�ay�%��l �56�;�����>�}�5��<E����K�A>Կ-gNYms��w3�&7N_�m(/��w�%-�7���>������	/'��?�K�4j��xI	��V���@�"��dg�(rڈ�
�Ⅳ~=�#N�����=����7�������p�oR.)��.d����i�� �����ɚO�e@N`�`��Z":r��]4�ݙ�j���"(>��,��4\J'���������ݴ���pY��`5&q����"+qW0���ʣy��[]A	^�-Oe�!(L��= K��l>-��%3����<7>�ӆ�K?98���0&l���_p���.:3h�Y��!͞���A=��s�vl_1����*l��	s�\����_�r�OD���I� �R�:dȞ��|2E���Yf�Y硏\yE���r�RaM��S�|L�e#�LwB����k�T^��Q�><��}���@#�yl���E[ȥm�ԋ�A�x�@�$�l#]a��L{�$@�NE��Qy��а�R+
������>w��kA�+��b*�#5B�\�sEj��;^��ǣ }n~���BGp��[�o�o_���.�,� �p�9F��ϛɻ}7w�Ƕ�F�Ԇ:&�k0�����N:� u�W��BU��&ɛm
��lF1���g�"��l~P��uԵ�`x��)X4�Xe��R��j��M��o0Ϫhw��K'����^!�%VI1�+��"BCD�P��ԀyMg�iE#�zW�T��#%��hYú����.�w�Aݼ���tb'M�T��J�ᣔ0�H,��}H
���gGD��C�KX�^���z��SIUa�ҁdq 4��g��tAi(�H�e�&ߤB�z�Pap�E2�����R�Ø9���L��s��Vj�ٟ2U� 6�{�(��Z8p�G��&�W���鿏�S�lI��=���~%��:�%�̧N�
ϖ�r �S=u\}E'�ӚnQ`7'-_�+��R_kb�U`�G���e�h�<o����P��3H��[b�ٟ�����A�.K��w.��)���Q!T=z�<���%(${��d�AoaQ�Z�M#?�s��!"f�Ƙ�|E��䂾ciwX�g?(���âg]�w�:�S��(�'rG�Sc���$#`��H�3�@�6�s��RK�ECgs��S(� d&(ܟ�(�Ɵ�CsI��ڌ��&�� �������o���A��@�[�s��u�{�
!�yC=9��ɯͱ��ׁNf�+"
���ʧz��Ӱ�����˻.G[;t�čV �ˈ��w�K�ї.@���I�>�XAo��k��v5Y^�[/8��6l8��ASm�O@�����2=F��(#������X�[��ϼ�c�_L7�!����p����A�����K���(uI��]���M����xw�7BL%�^L��K����Ĵ�p��Fs1d����T��D���L��b���U_p�*�W�	��^�U�T�!�g������+�3K�=`��=�K���'mg�w�J�yqv���dT6+VS���Q¾GU�̬L�}��Ggbx
R��zmS�O>Jz֫z����z�gp�'�u@�2��뷹ѧJ:YX�O�;��t7���8�����	�LK�y��<M?Q����6u����/���s/�XqW��暅R�)1��x���!�?�������g��(F=ي�t�4��u���sܜ��\�h/5K�,�F'�4�#r^Z����E"F8Ph!W{�PǮ*��N�U7���A8��A�=�s�%��P�{9�����YK��In�΄´� V�BuNX�	�_�ՙDf��s�`!��%4���݋��X`j�qg�ǭ������2�M3U�#�o�7ǅp��d�����a.b�b>M���]L��}cp�k��Y�RhPU���)����`����Ql���`�Fg7&ٸdd&�@����2��(�ΧX��3B�D�Ex����>�+� �� 3��8ʎ���pXH�/���Z<�T���3W%<��j�>�T�$�$E�P�B�3@5�W�Sh#��,��"M��$�UR�f�H���BuxrQ��ZC!���h�����M^<�6��p�Z���!}�V�࿾

�D�"b"BO��K�˱F;�,��F)���?��^[��̡Iܩj��z����q���9��]�> ƽB3U��M����"]�����ưi�D4�,�����a�xDF��xO���1B �ph��(e��7��g��p%h�_a���d�%��f��U��&���r���ε�����Y���9V�R{�哈	�,�JyЕC��`gr��A ��� Tb8���䇫�6���*t�z킯����-���d&m΍=���2��,\s��@^��M�I�RK�3M[�|�g�e��	�T�b<@�`�ig�]#�����O�
[�JH��Y��ME䪸i�̿ZG�j��f%��5�x��r��Na�@�]-���v��%���|D�5$,��W��X��������y�{ݖ6ɳӳ2�Om	DVQ��=����Y��̝K ��[�L������e��Z3 �N&�}1i�gq�bb���4Da�Kɲ#]��X��=�d
��k�'�2��c	�䶧�"Z�<A�톄`���2j�y��{��'h�+�M�4w�Ǭ��H~��Х<y�F�v��q��k��.a�ۃ�A눝�����0���cj!K�v�:�Q��$�8�|��A�[� �Z�ce��3e�O��r�4��[��U�f�Ud4w�C���%�*��If=�A����킴]A�%��\�#���/�������.��J�lG%�*���.̔�"u�l�!����5�@
Y���&��w�"����=E��ә����E/������Uph�����2_@�Fㆳ��v�:��Di���M��2�#���uژ�`���ٞ%(�?`�:�M6��A�s*$�^�qo�R|Z������ñ����	e�����:�F�~�㨬�v^�8è�F�����$꼕�P��YE9~Md\����
_��ʩ�(tmZy
*G�J��n�7�Y�.o����Z>���3���w�1^{_q4x�ď�����DOƜI�/�&A�k��n��B3�k^���J��9!�仛�~O�	g����Yθ���Y"j�fg��(2�&n�&~m'�k��}�|<gT��ڐ��e
ݮ����uL!;t����o��J��O��d
.��y'{�o6�y�E��AI��ט0�'�˂�S��uO%�Ϲ������|����Q�9�l�����2֘<{���І�2>�t��y�# ;�����V�^7���	�D����΁>��bA�G!	���
��R�'w�c{s8w��g���tB'҆<Y+]�`�YG)R�OQ��S��A&GVVdDB�Zd�;��6"�Ҏ�Y�zN>SC�����<��2%�+�]�,���%>+^��8"��FZ ���'s�[�n�*;���5���q�./���]��6�`�͊�U@P���\x�*�*�a���W��E���
,�-���)*�׭�S���p�Ì�e�N��H4�i�R|�+��{�o�w�fa��H���h<���,�L�x+�b��m]v�)����ԓwsn/�ݤwoGl'����+��?P�覓ZdҦ���V}��Y�7ӹ	<<���(���چ�Jf�:����R����pf��:d�ݓ-X�y�*���1;"	w���i�!��@,��!�����2	L��]���b��Q�tk�C�y�b�Ԓ�~�������v�D��7����>w�+�
�u-�;r��OQ�7��i�Y?�� �
C�3�;Ԟ�a��_W[/޸����j��?�k�>q���c絼���r$4tE�r���+-�6�����۟�b���^\m.����#>��5T g�FF-�md�D��g�uz@�*Y� ǹA�/�u�;)�Ï\���m�m7�� ��W�R.k1bB�榽���S�|;���d���NF�x��4P��I�G�ǲ�K^��9_8A|�ˬ`�0{��J��i���y��3@M���޿V��;8�Fx�y��"���l�{`�z���Laѻ�/2Y���J�LГ�0��4D�C>=
��yc'(c!���ݨP�������j���,�����M�l ��!��h!f�zR�nu#�5�Q9\�
p�H_�ԇ����������Й�
�Q�}�p��/TC������6r(���r�*�3��ԝٖ��X(��^�JKD��Vw,�,BK`��P	A�����E��#��nP*.�+�{o/�����uŶB_e
��Hx@#�<F�q�Qtq�A֙�B�I"yݴ��O�)�t��n�����*�dɛkߝ�G�3���zkc�L�x��=�Lp�XZ_���ů���a�ŋ����������j,7y��b��=�08�T�ê���=����sS��M���"� ��{F��;�0z⛧5|��"͟i���M�t?�-�k� h��k6D?Q?"M�6<xf�y5��r��zc��x�A�TV��.}6Y��N�֦�懟���|n���}�R�3��/W3�؜I=���5���Zy����p�E�m�L�&ĸݪ�:��JKI�+�� ������w�<L�(�y��9����P'^�0��[6ž��tgD���G)`���LN/1N����ڻ3���z�F���]��.�m��d8b@��Sa��2,qJ�����j<�W� � B�S�'{9TϺ�ɍ2����c��ʥ���1#��&~��tp�B����&Z;����ƙ	P����\�w��@��V$�]�򪃟�+o	��s�����{c��@�:AV��n�Ft���"�t����H����J���%���w�f�U�6��>L�6X�=���>���w�/�r|�#��w%HP�����|��gJ��z�X�\Ti۝�r�(�hk*��W����Ev�;�n{ʾe� ]�p�����g���63� ��)L�.(�$G�����?`��e��C��jVf/1��d��,f�BZ,�;�݇ E��h$���ۺ��*��IE9�C�K���/�A��A�;�N�Ѝ;*��bȓ�j��<H/f H�%K�ԭܳ��u��ͤ�De.��C5:�����aDL��XS���Y�����>�4b�X@��C�t ߹k9�Z�vh� �D��3QSqv:Iv�j)�u!ͨ�a	��Y�I"-�~�E⏱Z_m캑���dU���?
<J甏t�Z�%t&��	z7;�'Իz哝��&.�����F�3�k�����֠|L�N|7�!밠���o��.<�u����Ƚ�>5������o�\��^/��j
�bE�Y;�25���m?Q������b�(
']:��B��=�ǚq�
\���2���3��Y�T0���bl���mH�r��t���ᒃ�)�CV(.��_sL������y�Q������mַKR��}.�-���ן]۬�;2�Y赜�t�\�-xGC��0��u�n߳M�UV[��\�-4�Mt_�V�j���۔���A��?�Wa�s�3-�{�D�3?�q�rI��X��g�Er�t?ؘ�yz"�d�[�bRTѳ��?�pJ��6%�]���)��apx"�ܭr�J֥0Y����<^@� �;��؞|l�R�D1t��HjY��Ժ��a$dq�Z>T�WUŭ�T�ͬm*l�,n_~� ��:����ݘd�ld��UW�	���h�Y�KG"��ƚ'�-,��ɁH�����.p&�z�n/�G��n=��;�`�����nv	7wy��O-h7���X�}j�_h����:��Lrfx%ye:# 9��)I$���"�W��3�M����Z5���
���m^&����l��mX� ��O �;f&�o=��t^6E*+�u�����w��Y������È�H=��c�e������@��R�'���Ѥ�ү�Z�^��_��^�jE����{ŗO�O�^�遤�eBB����U�n_�l�S�h���t����R��S˻E���N�Eo����0q0m�T�JF�dKJ-]ln��A1 [�^D�y�Rp]T �"���V�d��x��B�}�@k��<�!LJ)�81��H��5b�=�dG�L�}C�-��;/4�b^Զ����	���5D�Hq^S/hi*U��w(�X�f�Z�R�I��c��j��T~h��)��q�2Q���,�d[�[˧s�g��N;�����"�2��`N�@���# Hd�ei^���P����2���67KV����rȐc	D:�������ǚT}Hw۱��-{f[1~u=��U釾<ަ����>-�!������m��_����qI0ſr�N�=ם� /̋hQ	�׎�:<�ъS��U3Un�BR��T4�+V�Rj�h!���eC8m��7c�7=�ޅ��`	<�ӅB���!v����fKBmZ��`Sq*�1��'i��Q��;#�bG��ٍ�MrC��Fs���yW�d����}�YxU�v�!� �pd��b1##'��Pf���K�2���4�q���Yģ��Ŵ0���/���6���D�#��XYti�m��X���Ч�����D��\�d�$��c
�J�wm�-_�j�2�FSxo]�z����(�gp':ZG�w�g��le*X���������Qo��X|��ȹ�L����#w�F�h�P���-� �����*�X��|��Jl�DM��ϲf��%(�&a��74 �ޱ��1$w &��QU柴������i�X.�!�����3�;�%>����B���:2č��}G��Y�:D�� w����Jhu����W���`��ך��Sޕ�W����t�y��;j���V��618UT��Aj��L\��{8X�N�o�`7��2V�0 �k��)^����<"¤u�t�������cwB��gj�2#�V�ƣ�G��(uɉ�l��k�!@�r�''?�9�.v��iT�jo���1H����@��12�nXܛ�f0�"��������v&�
��Jˠ�>RU�F �&�e�1�o�A���&8�ii�Kv ����Z�F�B��]��۰��gb����7��e�-���ƳC�G�L���>�Ș��њ1�r��'*&���� +(L���L�$!my��G�U�.�"���V�:uf�R�&����3����>��pV��UJ�^?����yKR ��5�0������GG�{�E7�*�w�C,������/��;Y���d}q�73s��������S��O]H��g�u��ldp-l�D���9�%�=�{�
��_!���E��Tq�*�l���8�Gx��C�z��u���Lc��2g՜@�����x��&)u���]Ţ�U6��w������u���-c��_l��=�ìƁb���QY���s=t� �V��Oq/�ǓRS�]�ưS��Xl�)��-H����z��]a|t'�r���Npʗ��8�g�T��k��)�{��)�0����p��J=�n"�ϣ�n�)F��4~�r;�o'��p4%,bv�-���䍫i$�bJoxCl)m#�~�f�#�
�f��t��g�rѽKy��1�>ͮL��%+-R���9�r
}�) �Gj��ʠ�8�	��&��DʣA	+h O!�|#�)a��2M��ϲ�q<v��I����Ԝ�}��r,���i�����2�`��O�ŭ`��m���AY�v?�A�f�{P�^����Q�HQ�z�:̎
��d�]#R��݁��+)���W��^A�Ű���Z�m�I������nj�ةe�h���s�$����j����p2dX�@�z���n�:�a/*C��s��5&A�c��7���lanO`�+)�I��~I�__q((�@9�-�-'�À�g��,���^1ϲFEb�[��,�R�k�U_H��C�ګ�&c�K���`����� "�����1M[��ՈbM��{!(t�\���-S�5wA��Bej�Aj�y��<�T!����P]�K�&t9�ơ�ϫ=��^΂��=�B>W��Έ-sO�;����e��:2��m6���o<2}����R�c\&�Y��4����|4R��H�ý4w]��1��K���4z!��c��OZ�V"@Y��zϏ��Ԁ��W��c�����Lw4���6�/��4+m8�ݲK{.m��i�b1�5z�Ň:� 7�����i�A\��Ԙ�k$a�07�"*B�@��(@�_����	]zK�7�:_�_:�P�&��d2�;���Xdm ���E�B�_]K58��Mz�U� e��� �2S�<+ �?��4?.\9�b&��!��a0��Y�[���i�{�;E*�c=Sp��1fw�U�m�:y*�\)�?�XyS���N��@��y�+�{��;�m��ˋ�H���{��x���g]��'��5RX��Y�`��"\��\qq��_�N��?�ט�e��LF���-���ۊHg�f��<ᷢ���O���C�2�e��� <�1ϵA�LPN�;�(!_v�:���΃�!3������B����H>��{�]}7��1�ͣ���#�w�X),��c�6h�I07+�
�|�_~p�&Y�3�l۲'L��
��YjZ���4��o�ƣ�
V#���o�ʿ[u�x|��Ф㣍�����so���s�|`5q󮈑�̓������a�w%}*��[	9���;��пO9M����.m�X&�M�-�����q�J��(B[��U����i�l�cb�EQ
GKˁ0y'��Zh�c��w0{�O�}M�k.\�.o�[�j�����L4���%�]��v�(@Ge8WC� ����l�:A�z�*Ts�d�1��+ V4�]Ma�D:Q�ܥ3�J;^�owp�bw�w5��\"0���-�N�ֺj5&=؟'�B���b�+��.h�>�j3b3iK�����%��jE�X�q����R�D|�{��� ��@(�#��H��:Y�
����F?.��\M�?�K�3(cZ�G0�!9�Z�	o}'#��Je'�d��l�I�ع ���V�8j�һ���I	�������𿯈���#�f �'�qqŉ�J-�{��x_�=��V֜�R"a�����ۂ�\�!QT���+��1~P��&mH�����T��\��䪳l(�bp��}4��;�h�|$��5��8H���.&�%ȪO�����Ƹ7G &�4������;7�v��\��g҇�=�F��TK��LQU���(LзkN���
OfH���6M���<�������>A4f?Z!B�d }���ǩ_l
M_����Z�2nt�X�B��^�O��1����Y����_�p �9\ay���O�#�n��O���	�Rm�+u���һS�-��Y��]W+����X'���,��uT*s3�3ϟM�~�2?�;ԅ.���p��[��ӻ����t�Z�\�o��3�����;U�qܭ�ynmc� �]^��RM���u�-9t��)�S}q�5{g��Y:`m������+DC�:	2.9�\�S|���I����C��h���fp�EA����1���5Ύ�j pj�q��É@3�ĜH-�AB8"Y����\v���r�#%���w�RKl0��N��&kO���@X���#�Er�WP4阥��w�L����}�7�t�g 7`���(Y1�����cK���s�h�s���wiLLo�������W���C�����q%�������y��?��>TŴNf"t9*���iz9]#�`�������Y\cY�<���`�,`���>lx#�	�8�%�_?������rV'��a-�B����Wo�����"�&��[�+�.L=�>����-Ig�J�]�T�LV�<ߐ�kۿ<���m@��bC�6��<�|�e���[�c��!S��Vg[��Z�Y\�T�������ya���Ӛ,���~�Ln�o���I!�	q3�����J4)�<��*Zʼ�����ж�c��,��8p�}�NB��1ě�fX�<ߏ�o�����U�B��˺<ǻ�3���1
�2c�����n>һ��i��6*��,��?!i'���k��P��?��� �~���<v�Q��Z�ӊd�&�����TC����@��_������`Y�=��Dl�'�P��#\�˟'�w�m����t������ ��W�^٤��~����<t J_���zP�q�QS'���R����l,KK&G�k�a��p��}`�h<���+e��I/a%�����O�!9��;����9t��lo����}��>Z��%��ڪH,1�"�[4h	'lxޗ��I��;J�=��dJT�[]����6�5��4���?)t����`���,�����:�W	ew6���8��W
��m��)��k�8�V|�G�GFlM��n͇�.
5������x	�yBVD�_e���ꓚ�.�Di��U���2`�����>��4R��Z�������Sg��VM-���Dh]Ad-K��U;̒��|�6W壴��
O��v}U���	�1��_��[�K���4�����F�qw�jȞ�!�[��*"]O�؆ad���"��=�*k��}���Q�p)
�]<䭟�o4�%����y��C�����o�B)����g�}���{L��p�Fޟ�AoI�F0��_��!�b>�/*d�ȟ����P:�74����*	Ƨ.CBV�.	��Y*#3t,���f��^��[Z����N�b'��ho�lq�Z�t����%�8�U�zy�<�P�/�FpN=O�T��o������f�� X3�C��Đ	`��݂�Ȕ���b�����^�/eZ�F�09�u�9��|�a��B= �H��	� ;J�~�jvt<>��F���|"�f@�_n�����=����d�ݪ��˺i.�BY��~s�D��;D��L�kg���-d�uK�Ȃ�c�̣.w��h���NR�lE���6�l�$�%<	�ũ�HQ�_әN	.����׎e�g�/%����hbwV�A�x�\�k�k�}mJ������5��jP�{9���bs�z$��h*���k�d@��տ����1c
���x���ۜ���C�~�99䎩E���H���n�!FǤ��y��X�_�*�qQX]㠡�m|uea��>n�q7���P��9�*4�(o�C#jٻ�qR�ßS4���|�<�F�C����}��m��3QI(��04��x���#�9Ϭܒ�����5sOT�t3��7�s����<���pR��Չ�Z��E�=8(_�!�,���?~_e������B��lҭ����һ:��P��0�F�Pk��E���d#i���B�"�U��մ����W�9������Eػ�8�o�ˁ��*K�Q|�}{x��>��kp�.���<G��#��5�T���7w��v�Pw Ғ
)0^�0���=���#��+��(�m�A��w��.86���MzV�	��F�woF���!�Hc.�5C��s����&���y�O%'v��Z��ه�Y�"�$�p}�ܶ�v�����.��,VB�=$��4�TN&�^J�5W�$��S�B�v@��u�����'��}�j�B4�v'� ��-���X���_ۦE�]�p8�ꮿ�⊒t�_�S��Hݢ���**���Ɲ�!}��n���!'!���;��o��i""�r����:�� U��%43+w���y�w�`a^�rĊQE���8x��&(Ϥ��2��o��h\�_�W�O�`�֢���c^.� ��%�� �S��k�t��k��TP�37�[�>��#�(y[sĈ�E/���2r!�R�{>UB3�}����E�р�rY=U�l�Q̢
!= ��2��wǘ�i�X���f��G�y�A�w�#6�	�"4o��GvV��Ջ��v�u����k���pwkd;˶$���6�QIz� ���y�Ұ�����b��(���p��H�f6�͙.T�B�v�U<�xh�r�{^h��ݹ]CvYv*���q�U���	W,A�f(sG��o��,g�Rn)��G�.����Y�Z�ɩ�cr�{t�n{Tt���+�"���ܪ�J������|�����\��58G��ϭ���\߿�8��}$���AFtʸ#e]�<
��@��#�{�u�Cy+c�G\扚؁�e��s���6���kJ��9Ϩ�I�H��)�v�f���A
�:��n���@�]�s����?�|�"���䄪�!�sR{����%6O�g�"�,W����i&7FR]��4���5��%j�@�#��N-M���Ȑ4���7yFX�5�|h^\���Ja֭�REM�zLI�� ���"�:��%Q�h��Rp�����qLY��/T��jx#M���Hv�V3�~"��Ie����Hk5̤���$ >�olG�b��;-�0��W_�i���v���9��*�X%i(�+𰖒�`��D�_�Ͼ�� ����~�$Tˁb�|V_ˬz����h9{����-���E�^C�r�(��&���n��6`6��Zb�].�GfOfM�w�甬BIb����(v�;�G�:���C���P��r�'�J�Lc�!AsД��؊�$x�tcW��F�f��݋E��g(�ƙ3���ڰ�C����[,�����. �.��C0��u��_VR\�3^=�������5��}t$�HV�	���G�%�dH�x�\�P����w,o��vmQ#��P6f++ٍ�}�f.��P��5X����&��KmP�~p�|n�4��Z��st��W�v1�H�1�bt�A(0����;;�?�g`��;�ܘڻ%W�!��d>˖1"��X��L|9��ޏkל�xG^dy�n��*M�K�F�W�|J��IO��G��b@-'��1����*Rؗ��$_���x��F��C�(D�v]?ڠ!�t�����T���yjDq���h�P�e��J�d{+0xI�������
��	:��pu
 uƫZ��"����$L!���:4_+��l*rԛ=�:��+V�8��kB�j~�&�a��D2�G���tu@�J�E܎��O:`�aƷ7�Ŋ8.��X�~ȭV�Z�~xĉXR0��xDRtJ5�7��W>�᛺ޖ���~T�@?3�@�0�J��^��<pk��i�=׉���?��NU��/Z�kp dM�,�����v��Z�)�n]��%{�ƑǪ��=F��J�������G}�ѥ�P�˧(�7��_�o����H�>��<lh`SBKhzDDp+����ھ�m<��/`^��O�/P��������!��>���b����)a��G*���@��)H��nvw^Tef]���qp�Ui�TdK�XLt_�+�A]�-A���J�۸�]g�#_�H꺞X%p%V�-QyL�o��C-wRWG��y���o�b�K� *��Y�L���;f�j��T��#�Q!Q�G��5j�"�y4�aWv��������p?+`�e�<���%�Λ��jԌ1��YA��\��e�EP?�b�/���i�"����4S�
�n�6Ȝn�gr��e��6�8�U��{�%#��d\̀�|��QҊ�`_����
�z�ڃ�"-ƃD���֢[�N������q
$�#ҹ%�<f�_wWf�'3��� )'e��j,��ri}>�n���#1�=�V�=Q�������QBs�G�e���6��)�G	΁Є�%r�)�Z�w�L�w�n,Wt��y��sɄ���I�;�>{o�wq�}$�}k��S��A���X���H�5�FVZ|7Mf��uR���I��9X��(�4�QPq�o�L��>��a��Ԭ/>;�4�?�	]� ^7��پ�k��ą;�eG����j�e�l�qC"rf�vb��d�j���{��+��m�6�'.|j�@FrIW�
}�ɿ��~��6f8LE*�	�����&ۚ�%<�z��ե����&��\R��&�k�1b>��&ӎ����͇��3�-���v(�Q,$�퉭5z�8-9|����G\�D\��z����,�_�Y�~n��NZ3���c��ozU�"��f�0����M��*^V�_�1|}��7>h�
�x�X%¨�y�.�g����/0��7�q�-,g��LPn�C�}:^���}g-��	�{�=$K��?�q��x�O��ju���-T�12���_�1�`a���DU�r�r/$'?�ԓ��B�R`L�:�{�X��yRJW�U���p�>��S�b�Y��k��{mTr��7��XWsԛC�-��ܽb�7��<8��[������e!���$`d�m���)��������9u:����aY��x�#^�H%����wQ'Z������nΔ��F~mV���$B��0�z��t�!�%F5� ���)eE&�L0��h�+��B~��P7ְ�"Qo:"�uI�tV5A�R���kcWa����=���9%' "F���	�!�_9�l=+ʏu��hs�c7gb���C�Fӵfg���ԧ$��C��- �wY�J���Ν�@�b9�2�Nu��� �;�)�2�O��n��7��/��O��.�]gc�����8�nIjA�l���(���	�s�lO3����'��ҿ�����j-�X���Sr�zA!lO{H�g�d~�������x|f)&��sjL�"�=Y������lynEHc�L��{�r����p��������'�Z�bP�qWHX�1�6����m���Զ�h(B�ɞY亨!U�Sf�^:*�韾^U�p��'�OճR�|R����
"�Op�~�-ݩ�ӹ�/�ZAϮ��g��`\���Lws|�ǋ���]Z}>y.�G������Ҭhu�����t<ĸ7��Q9��~�d���Ol� ��g�
���4sԴVs&�g�T��6���W�=��E���|)�ok���]����q�1�9���cɲԆҟx>eUe���A���-(My���ي�|
29|&��lʆc�Z�c�u%kZ晃��`�?@����?�۾�#֟X\���o����}]ߒF�\���r��E���]0� ���ؼ�Ą��w�$;7�6�Q-_�?r��a�"	a��<��L)ױ8�����B]{ �xзx:9�����B3���{`_��+��ϚJ�Z��9��z2
�}_Ƣ�"ث>	�A&To���Kޭ�j9XQԢ��T>44��Nb4�B1;ų�x�G܄,�s�J�>���:��#�s	��B�=0rƿ�N^�إ�iȎ������mm���	�"�Tj��ޠ� <�j�ml՝�[���F]{RV��o�>x�/�cF�{��Bq�W�9��E�-���<���
^���� ��v��%!�l\����>W/+��6k�9R�RR�x�?�G>�:ہ������fͼ��oUyI��."�x���H�宎�[����E�*6���e�bҿ��
�9�f蔻uv��D&�~���TJyed �%\������ ��l�ϫ_�Q�:�EW<cf��.U*a���7ώe�i0��m���4��iS�fI&�
�.�&��G���l�B�;�f���3"���@��_<�Q�����$}�ؑ+�}A+�hH)�^qy X���O�E���2�l�,�_n�'�f�{!�����ͤ?�!�i����;��՜T��.���m��q��.���I����,x\E�^UB��Lfp��z�==��8�k�����G�d6��i�)ru���ȸc�@T����.� ����o1 ����:�YgykM��0��G#�;�mv-�V�5BZ,p���7>�4��@�q��|!�4|o�6�U��3�s7�vF|7�B�4��/mw�J�l�c|<j�V��W��d8J(gT��eҪ����Ni�G]��Ta_x�^͖�.����"�XU��Nͦ�!��I�s���>ڗr���M޹�{�N,G��ϵ1�����t�\���k�E'm��
V�u���b�����f�&vH�C�C��^caȁ�V^zC���݅ͦH�@��,5����$�;��`�������E�`Wv~wS���Bw���f��ӧ�I/�/ت���Rڇz��~���	�>��a�*��]�+�׏�<4BjPڪ͠Pu#e���D��[�z�˸ogr��vN�;���5�<�	J�W��Y��B@����1v�S��n^c���aKmh��mz��*�tQyZ��� =R��o��Jp�֯��#�D�Ө�HP�p]$��ۆ�2�M�9$h�K�x�TJC����=����oK�� ��<z&ԣU�k͘й��֎������֦On���m0�ʂwx���&�V���X_A� ���5���M���z݇�<s�Uku��V�����V����D�7����ju��p�8�����ƨ����� k8��h��N��M���?�蹠I�=v�+,��B��5�M�bZm<n	/��$lbZ�[��Ű�{�w?��\c��SO���{ږc�Q�( �8�T&�s�m������r�Ƿ�;͑�D3K�9NP��1�9��&]�`|�m�V��E��b�g��c��M:�`D@�����s��ƏW���e'�Y���)�񏜅 �*�����2�\��P���&d�ܪh�|\?yƤ��1\$TMi2B,�y���������T�	*=N,y���5��5`(�V���,�f}ksMr4V��iJ��_&�5��җ`��H-
����r-?Cs%�&�o���k������C�L N_���+�{��Spw�e��k�(�D����G��s|��� �� �Z�K[U�\��Cʺ!�S*���Lf�*C�O<,{(��;
��%�~��ۼɜT�r�T-�Ϳ�u��%�I�wȐGmi�^������]��"
5˗#�)��Hl�?�W�ߧZ�"z�6qqq�ih�,Ḥ����Մ��-���\��z�l���� ����V�j'xD� K)�?v�h�k�����XB1�y"\���+69��k�+[N���DC���U|�ң$�wp�?N��X��@�V˽��m�Fjl��n��q��ˀ��6��a���3�[�D�PJ}�b�=�x�Fޯ 7TH1p%��`�}�;r�';����v,CtA.1U�r�:{���7����'LǊ|H�
�8b��q�� �y��)'����΋���2��� +�aXe�^��K�NP��5�" %�x�����p�p��l|��SϿ�"�qr0�	�ي�S�0pZ��_��t����=hM��_:R��'$ߏ�����!{�1X��d�Q����s~d]?֊E��Eܨ�t9u�}S���JB�T��ػ��
�^�fly�����8��d���C��BMi�Li��D�	!R�6�m��l	�L�9�m�0�V����Z_���TK��)\)�!��(�5�-6	�1Q!'�<��.�o�IQ1���ଃ�,<u���Mj���w睓�&����>���җͳ ���}�;�����]����:�	��.��?Ȇl��hA�3���}\�}
G�ϧ�v7�箈Vh�X���m�:�
�
��[-(���k�q�v9D�J;w5�����ů�u�����N�@~�G:8	��d�k����'��Y��)G�7ʺ�0-�z���r3��L]f��_�e ��&vx�|�wp�=k�1����c,�Y�<,M�m�v���U4��f8�����P��mF�x���� �_�Xz�uC%}c\�T�BrAdW�^H��y��(c�ݕ�m"������<ef��7Z��0�� 뿈���t�eX?d��h�(qu��2���WX�N`��{puHAq����;�'�3^Ќ��8WU�Y�����0jh��ip������.2G>'f�3W��yVT�r���=�Ġg�Q�:������E��{<}PD��T�A�I'��,�mQ.BȎp�L��,|��;�eW�Wt��g ���;,] ��R�|�(��������PS8��)@O�膵�+��ջi�.���S��q��Q��k�5wY$9R�*㮁qR5�ţ��4T4	�&.���.���0 ��1s�X��f&R���S��������; ��l����C�i,��vb�F=�q��d��L�2z~�JOM�X�Q�A@c̈��/�2�X%Ea�M�aB�����Č.B�tU�}�!��SBgצ��JT�m�AA)�Н��.�\Q�� >,���<7
���"�?H1��ȋ �E���xpZ�����6��.ɼ	Q�Ь2�0��8N�J~�4�cj���.`���[�X�cF���g�3�fv�$I�QH��	�7yhY�x����͜�ߎL�zx�Gb�`�s�<*�,:�)�#�,��H�2��aTq���#0�������,��'d���"T��X�.�юEo�t�̽���� �N��X��gS���dtlM/j˧��FǰHtZ�YOtǗ�T�7l���,��܇���@�:�4BV�
g(��*�'��g���U��{��7��!:��B�\�[ؗ�$�"ѱ	�w�5����VդL߂ ��z����t��s����G���)���9�+18�⎏�]%�t{f�zp���	��8B�~̀�PT�D<϶��^��� �H��[ž���J�������U�<��V�7!�$�i��;�߅�"H6���N��3�:�� }��w5��d��C��u�gg�Xv|�R>���e��L\Ӓ��w�S������>��,$#�lg�M���W��vu�N"�|�?� ?&ӧQ}"���"�2�apGD�~^^�qCq<G-X})R�����\��沘�1�AڈɈ\X�Z%FoH�#��湔�{��x���B��)��I��794��K�b����h�W��t�>)���7~�7U������<�y!��|㌑O$���u}Xx+9�|8-�V��lQ�81&���֔��Bvl�x��z,�~<����K���@���Nr�sB�����c��gi��d]S&��39*��D-��\ 20�H�b8u֔��s�'y��<xwc�ug�����dσ��4�u�:Ij��n�� @m�'I?�1A�(M�FejN�civl
��Zp
�� U��F���_����`�s��bj�&E�ɨ�9����9AD�����{�CI�itF��"��Tb�D�� I�r�8y�ⲱaX�(xm���P\� ����M�X~	�U����~+,i �w�����&��q��>�6����
���5م��ICC�����6c���F�3Cy 2��JLpw���oƕֆv�oY3�hy� �)|AHL�
�&����D%;�̲}��f�j�q��#i�	��8�P�Nϼ�p�	A�di��n��������S�3���o����xJngb �ʼKo��뗖��rqj9١��E�|�����C�#Lj�`N0�Y�N�U&q(��^�2hI}? ͘3tF��ҝ#�H֬2���;T��qo'gV�)�C!�������Ɍ�jLǞ_���"�{�؈��	~��l@J����k@}M���Ѭ[��;h�:��X��Ʀ�׮���=��.�/�z�-��u�]��f;-�
��[�B^�� �Q��Q�����]i۝&�����K���3��ҏ��!=�Q��(q,?�_�i��1�;H���ј�t�����k�3m��[�@�V$�������>�7���g?tu�}ې���fQa?+u aljC4�߰�M��>�aw���w�~���˴�mG�0�:�9*�Q
��~rq���AZ>��S������p1Ne�R��Q�����u3E������&�n'z�����v�L���7�����ŭ==4Ӛ����-�-V݄�{�f/w�߁(�ü�����S���&��cz���:���,������H0�z��[�p�H�v���y�R�<D0p��ښ��<�kE��y��l_�Ƽ���h�}0I��*³�K�*c�b���V�}���U� y,4lZ�6C��x�%��ds�eո��#��#dbvE|�ѣ&~���_U�Q��>A��X�x߫��%��v+��f��<�3�'w��m�>�7��1�I�}W`�&ڗ��qިΒ�N��k�h9����Xq<�vޗ�K��|�J,�H D���׳��8�o�C�9����ݓ���"��b��SS�b�DU�߁��.����#��6����x�k�m�ot��jy���@WAM�0���۠����(�M��=�'�G����~Z�s�&��k��{�Le�T�G�{��dA��L"%�%ǋ��1!�����O�Ϙ��5�z�O��R|���pn��g��E�8�~�.���ADK���ƭ*xX�h���e9�EְM!���E���J\��������8]�EC�o�T3�:�����$�3 ���b�� �����>:"Z�yװ�l�K�&�AT�/�FÊQ������J���6�3�̲"SЅ�����:4=��-n
�i����/��$U�'dS����E�N����'�;jD��Tp�q� �oTKDcN #��zU�ЎϹm�J�����ޏ*�>�I.�� ��;����B�w�}?5VKW��Oi�p?��
q&l��y�*��H}ɣ�l�BjE)d���}�ZN�!���<���>X�����<+R��(;���uչK����R.L���#,%{�����*W}�˙�4z�X�@q��q�n�Kn��E7�Q�,�=9>��[�s<l&�2�|b���V��w�����v�T�!�N3�<u�<�QTt�������'�w����O�o�b��^P�'��4M�i��*�A:�;�}��<.���������l���ʐ�/�@�}�u|(FR.��u �2��XF�����$�HiW��'%��`/j��qZ�5��,�8�=�4 @������#%��\)�Dʍ��E������	m������g�=сO��xcҕ��/<��L�'Z�e8���i�
�`��_
�4i!^\O�FER���v��$�U��6��K��Y�KiR�S5����Yp�%���GO<o}+$��0n��y���K4DT#�����^2~��j؎,٠�R}O�@�_�:��w�<3/G�5��ētAv�tK��3��f�k�+��ݼ2�4��!���,���t�e�^3)Ǵ8��a[���#d�F} $��r+���n����hI+��3C`��� ��o� ul�*Z�h��81b(�j�6q�3�0��T�v��R�U�r�~biUE
�9��6j_�Μ]��zlLY���p-RD+�m�X�UPk
k ��$��}!.�;s�|àv�Q�"$` �؀��tS<�E���}���psPg�قX�F�_$u���Do`��@�Y�#b�	0���N[\C�L|�^xX;1�B~Vx<�漐?�B����U6���������!�����D,�w65಍��h���H��ʽ����(߁h��j��������+J.�
�$��N���f��Ӧ�2���.Zd8f3�~��(Iњ�ǋ��i{�G�)Yh<tF����.����:���;w`R�k�_�ο����QÉ�����E]��!c#+X�_3+���;�'��"c�Pڗ3��]����6���d��*]��;rm��]j�į]gl]Ӕ�����3W��C&T�����]�	膦��Ly�H�W��F�C���T�o���-��J^[	��ؼ���<��A[��X ı{�6&g��֝���N�>�d��ޑ>c:�Nʹ_�Y�:8��	b����1�R^E�V�nx�B�A�6�{�dS>�=t	��!��O�jџ9��B���o������x�8�}�	#���7��::g���t�1��fϋo�Vj��"%�;i��U֖�eq���bMj��߫��4YR�+�Y
h�r�3�+y
2%e��e�r�S�4�[��Z� �C��7�q|�8B!1�p��4�e�֝�L.��HG�6�/��1�(�?��_c��ļ�W�z7�_���uܮ�kX2�ԙ�U�@����̉�SW�?\
��#�N��{�`��2JT�/բ��wf đ+��\��F�"�-�_�6ņ?4��;0�Τl�4ݓ�̀����  ��;��"Ӡ��Lޓ����ς$ C��tFz�����ƀ��jv�b+
���^@ǽq�"�Ud'��4�aW�P����ud�@��z�%)��P)�����1�t��y��T������I�9�R["��?�����4I?ҏ2^V� Ѝ��B#� ��h^� �f2����Hl3Td�z��W����4;�#���DɌ��2SH�X��C�D��`g�_~�oK��i|�����ܻy�kΉh���i�G��Ŵ��U����^)�@�eEb'QB�����1�m�lG[��#�;�E�/��J|�FZ�1�J�p�D�
e�G��O@|��&�]��v��e
�{"lH�6q��r9��wr�a���[����$�(��xWɄ mXӼV��8ɛҔ��?t��U�ULb��/�a��2�ZVx���W$�}�$��m[�bJ��$�F�5�dG��ɉ�/�ݷ�����Vc{1��E5f.%�������\1�oA0S��GD�j�4JYe�gTS|����ܾ]l3�o
9�����R.�F	����*���0j~��P�F�iV��)� ߐ�����|�0#���kЏ�%����!豣ZIC���Kw
d���������رDZ<T�S1gDa !��cv�`F�l��/@zW�B_ԝ��UO:�����5h�Av��}�a�ٕ���G?�c�С;���*K�DТZ�rb wz��7����j�~�3U�P��� -�
vZ���t����� ��8Y2���?�����AKʇ�������E�o?o�k��ոT0������c=E>�~�2
YBʯ9f�h�&Gx���A>�W�6B(�5.�;0 (�.(E��n��bQ�����%l�������S|�^�5�8{���=�so���X��Y������}�M34Sd@
v<McтӲu�l�@��	���0��NU()l��s����`N!L���-A��lg�~?�C��<P]�l��Y��!�9^���grо́#�b�����@���j"��~@
�*�	���{yDV%�>��(��C�=v�6��RAE�)�����&�;�fP<n��_Bg���*��H��ח;Kĵ�6�P$�[	��׋�|�&��-�b��ȉWd���sD��ߖ�R  ���HTҾZ����p����������B�*<g��ꌬ��h�!���f+�m����� X[�eY�z�fg>�]r/-H�ˏL~�rʹ�mSx\��K=X[�k��Xn^�NZtѡ��p{�f����7�;>�.1�e2���TRH���[9���AߺK�|C�˾V�4]��w����(g,��9�xhQO����j<�l��0=ĉP��}JB(-i ���B�AT�����==������ x#YlC�H�Dޜ�tb�Vj��AW�F�l�Ť��a\I	,"����j������`��U�e����U�n�K�2���؆b#�9��lR{$���̹]Vjy���>�H�;�g�$4���E�S��掽�F�1
>b������y�b�7x�w'^qN<�͒����k�j�rf�����(��NX��/�ۍy^���0#�Sum����xXv�$�tE!���M�J�o��Pm-�f ��U��I�Í���!��P�N�\��@I\hE���q4� ]=npS��ў���	}{1M���p��D񔃛7��� ��e3 =l
����3xlfA�ay��k�rĵkn\�����,����/������s��/J��:��6`?=I���Q�ඈ�!��� ��̓���e�Ȩ��:�z�+:q�A�*w
o"w���r��0�s�_6,�O+hj���d/�K��Ֆ���a�繮!�* ��i�/� �糂w�Y�R]ZyqO��P_ݻЌЧ̽~��x�_�*�;��3�=��UOGD}Ǖx\��3�_[P�	�P+���i�d9Z���|��V�
G�Y/@�hVۣ{�y`Q9��c�2���HLt([����m/�7��w��j��
;����讒|==6�O��I�Lޗ{���7��r��!��(�x��6+nIJ�Q�Q�gi�t��쳏B�����ylg��Ke)��_�1i̅��F5@�a��V�ʪ�X�?��ز�W��=R��|Ze���'O`��7���J���w�^��`|�w;�<7�[7�Vr��<J>m �8|sK[*�Ee�P��R����ki�ن\��ф9��B�obwg/�}W_�	r��g�q�q�b  lG0�3m�^�"
��1�^Bn<��i��h��^
�ɮ���;=�v�}Ov�T���aubl'q���M�W���?2�ƕ���_|�[%��8�#Y�p®��_
�E�ɛVǺ��Zq���㩷�RV�z��0�H���o�'��5Q��Z
N6*v����6��b�7ml}�F����5����^ak�Os��
�� 1�(e��ߔM!?���m&91��]WA�œJ��1�jd++���iQ��5;5���'t\(�Z�
m�Y ��J�u�9z|-��b�+]�Sl�)U�u7#��!�.3�17�L�PR�)�h�L�Z��Y8�D���v#�3�{٣�W���PQ�8�SQ�uK~�k���'6�1Pߎbl�Jȏ0BM|� b98��K񯞲���=w�5����*;̑�q�u{���sW#$���?���f�1�@\R�&���6��'-�Ty��F5�|u�RBy���4Cp�����c��G�yY�eq�lq���7Od��c|��М]���#�3MƧ�Қ�Ne�t]4F�@!$�#�ɀ'��?d��#�8��a�o�%�������A�*GԛUY�M�!�A��-�{I�e�.�����K��CT�:�؈K乸��=[�!��C��X�x���@[Sտ�����Gw�;G��1����k)�{�v��؟��O��Y��Ck��A)J{h���3�e�x��i]�_1��'�D���V����eD�d-ࡠ��-et���l��h�OTg���ߪM�L��������n��^��st�9�tS�i
���J� �:�gRu��Cc\� ����T7�NP?ӆX!?������̶�w��!�%�J�<mL��W�k���<�Ap��ǥj�xW�Ω��1be|�������ˇ �D\##A9���mn$��L.�2ࠓH� b�#5�2���1����O!�7�jn� ���݉��;��XEz�%,|�4��T���"�ު�<��S/��zL:���#���%�zX��C%����%Nu��j���b���ީ����$��`��zС}����ƫ��K�w>��rX&�����}2cBNk6��&�<�zv�d0h�=7��N �(����k�k%�^r��s
$>]4�h�AɦZן�5J�N��4g����P�,������3�낫��W��6��Js�*^ը�׈��{/�r��ۄD,t�����6FUl��X	�]�����C���p�Hlf<�0i; v.+`!����l�##_�`q�L|������]�L���EY�a$p�ӫ�.�p���%�8+Ǭ�:��M�l#�2�=�����+�e�1�k�`F�ȸ�:�ս��@~nA�Yex^�������u��bZAc�D��Zy��ٞ^�9��.'����~��1	s���R��	>�L�p���'��a�+��&�tc"yܼ�
[�7z'�wGwr���`�J��;q���:�c;o� �z��� �m��an���#��]嘓<>	íe��u�X�=<� 9�G`���y��G�}�d� 	A�a3�?�3)�\b"�����h��8.���
~�zJ�b@�?S���,ʋ9��'�/�ڽ�蘄#�й��d+DAC�Q%���*��f�o],t���D�D��%�FM��иx��WL����a�i��G��J}��
�$���<�ȡ�_��[��M���;Ox�7����J�HI�f]>��f9�K�	��T�%��	\-�m|<��ܔ��*9F�_+hq�ϽTv��J�c	n��̺��{�fw����3ۉ\��Q-ֺ�b� �9��o�fÑzeO���"����v��a���f|S�WYAz q���	 8��_x!�#馲�a��n	�����j`Z.��";�0�09�6�����=��L��N�"<���@%0G���_~�
32Q��Z��U�ʀ�/�V�v��t�К�\U�����ٜ5G�����&a�p*�{���k��ࡦ��d0��.^(�>:�#���ߊ�D��_!z�%
�P{K����dg�/U�y~�3���d�_lD8XAf�2k�~г�w�d�*^i����,g;�H��T�;79��G*B�)�2��O�n~����'[#s��F��[]�-n-���!cP�B��B~{Wx�|�������N;��	)=oΒ��b��a(�j���A��^����>S)�z ��� ,M7��m:dGdTB?����`��+(���n�<6��\��+�\G��VW��)�c��O�	έpe#�(�"��e2����o��v�Ou��d�lBlOJ?Yù�m>�����?��D�!.3+X]+fk=g��ԋ�szlc�t6��v�c��;TCh=EB����0_�뗹=���f������S,�ᰏ)��W�+���&̐��?��ֳƿ<D����U�r$:xK�4(���q'fm+�@�;	��J�+�gt)�^Oi��I�h���C�E#Z ����NN��]1ԏ�ʣ����eVR�^�eT����>�ۙi��c>��u�nDa\�1����+���ܑa��R�ŀ&]4^*`bw�Wd�Զ�6-���.h�[+�AB�Q��w���*7�������ށ&��"ժma"�lL�q;YGo�C�#��O���6��
y�6�=�0�f�">��J<�L*�]�����uY�_C�]�O2a#>��s'�L�r��{kh�ҽN�{�]��ʔiv��A�mZw��a�km�Q���˥����6(Ud~��m�����#��G�Y��/��]��N���:EY���@T�Wgtw�f�f��+^����r�?�\u�dL�\�ǖN�3�1��^HE�62�uп$d�>e�2!�k����T��WK�k�G�Ԋe�.��A���WQ��bK[�x'�p]Fú��%���񥚯�J�M��x�s���,���wx�X��̨ϳ�D9sZ1!t%ڲy,�ݬ�c8���^DN-RPi&��V��~�=U�	�vYKW�(�p����֠��{�&�?@�� ]�袏�V� ��T־i��Ѥ�ie�W
R�qḥ^y�@X����mX��e(O���i�d\L;����=q�8�r�lN5-qV�-E�ZD|�ׁ6��l�r�h7Z=�^��8�bT�~n
uY�{�jE}�D�W�Wۢ�e��/���n���o�_�-866�8MI6\�(:g�E*��0Iл��d\G��"�sY�+5��(K���/�ǚ*���"�b�H'u��t��C�b�Z޴�U�J�PS�� �Na(����˭X�l˔w�X�J�{�np��o����~�!����B����p����|�kFp"~TU��2�c_|��w��)�������_��3��v�A���i�sN6����e�����,]6k�ݳ��J=��q_Z��4�����j�'���7��D�'Q܎��ij�)�/4N=yw���c����?M�h�E�,	�ZV�	_Gz�`gڛus���Gk��)>�|�1R��z{���`�A.TV���nG,]�e�
nwĝ7�}D]E�'�P� ��,T��P��~��tܫ�I�ՙ�N�3;U-���`�z���$g^e�94��-tY?ۉWb _?q���>�S
w�N%�<S�Y�{[ԩ�28�iwUH�}�Yj�r��tpFVg�T�� ��1�UTE�j��U��WJkta�ڷ��?��o�b���Pj�_�
 x�^����W��@;~Ũ�iW2�����W�@�[�n�vI�������`��al�@��*�PI@���v�hԷ���@������q��F�y�nqzQٝȧ��I��2:3�:��"�]������8*��� 'H�|̏1��Ɲ��=��#i�w��|͐������j��"�,!IвW��gx���Z��G>5�;�C����)����\'P�iЉ�yĐ�>IwS�WdY"YF
���!��.�6���Gm�����pʦ^9�n�q�eU�,���m	
؏��ӟ�I����b��Ֆ�'sI�P/cBU��Xh�V��vkz�ML
l�k,����ϓ�]ܺrCÝX��u~����*c'/�Rfl���`;�ڧذ��l�kh4L�	�K��i�ϵa�����6�E^����:e/�@b�&�%�mIz\,#�9l�=� NC^$	"U�G+'���!L���5k�e�K��kP������ϊ�i�k�$�Z���<�K��
�F5�u㌫?_�}���ڪ�f���pME��I`�V�Z뚸�b�(�w�m��%��ώf�{a'�s��\�מR���sm"�ɺ{[l�	8/��~����Jr/[qC��K��m� �q.r b��@���F�
���$y�´��n�֗뛗7����o)�6!�#��X�j@L�g��� �F !�t�B�S+y�֊ c���J�v�&�/.?�a�%7�1���K��Ǵlo�����&5V&�G!1W�@�CfL���B�*�Y'���Zo�h�O�����*{B==��`�����W���J������ ����S#�����%uu2(Hj*�am�[��+����x�d�we#y��cP��Բno��06+��|��o�͎x��i��U����_)�2u��T�ݗi6�c�)E��n�G^-|�Ke�����E���~�)l�Ŷ��R��D��&����b����_h�7F>̊C���"�j�ZB2�c� 1�*K��Է�	�Ͳ�`��E9"0�k/��p���/�2g��1�C��s�;�e�<{�>��3���V,Y���t5�]��a���QC�^&W�Mœ9N^̭KX7�ǉ�]��i�N�c��@��Dga�NMX��ݼ7W�<�������d���R_�u�d�MZ��a�|ɏJ��-��S��a�=r���1���Ga"�Pֻ<���'�I+O.\{���� dv�l6Q\k�}�s�~���0����
�(�a]>��nd��E!�{��E x�0��J6���d�U�u�r��ڦ��}8�?2HmN.�W�K*�e�n-�K��w#��KMC@P�pÊ&� �����5J���*wv�)6��I�TFb/�4PI�{����TKK����E(���V�+w
2vـ(.ƞF��wS�<���o��#�������iԌ�����1�8�%��/��t����7�2��,���iE����]�r��ÑI��ԙ�z��X�'zg��j�R,�%�?�/1�8�BF�ۋf��]%Sqb��;����lo����Z��Z��;��7���C����I�1�bҨ��n�N��~��i�/����|?�.`I�T�3x��!D�a]�)���^~�ŀ��
݈H(5�z�8��u���?�0}��謁#�Z���㬃�/}`M��t۱��K��,w9���f8O9�L�b�����D�B�\���)C��T(��=�z��\�`�W���b`�PL�ʏ�Lo�@�(�N\%w�����'0�}!�0G�湞P�Է�H&`R�8�+��z�0��A �~p����	<� ���7��x;���&/g�.c�����̙���^ߙ	���KsY��3"
4���r�),�<'l��E˸����ט4Z��J3�;Wi?���ǔ�`ϕ'7Vo��e�(-��������sD��_�����F�.zk�
�N%�8G:����6$	��p�*��H��0����i���ZA)� 1j��Ya��*K�[��K�W釕�-d:�8���R�H�w��@a|�mw0 �^&�]g)Ī��{!�tEDp���d4٩܉��%1K�/hO�oh�tɥ좧XON�����MGb��]�
~!P^5�Aw����u�4)OR%NR���Mڅ(KQ��7����)I/��֤O��ϲ���yk�S����R����n�؍	�o����]�^L��7�E���&���z�SN{�׼��j���I��$?��������?����m����t�	9|�uC�
2 �7�HܲP�P���(��.S������)���7o��TaA�ڑ��Dz���z� %��:���υ9J�AT���Ռr�g��o���CG��\j}��Zʒ�%xs�]��Tn��&bQ-��,����tX���SM�}ɹR�Mt��|��_��t@g
Hc��t[�e���ZW���ѼZ*_��ƀ�~u�I��������i��;_;#�� �堈l!fYb�q�*��o�����lY���owJ�b�Ajv�M{�����-
�]�&�2�1�,$�K��p{z����{ule�ॡk�~{����n��	4�,�]�!<F<_>�.��'�
��R������ݾu�X�0C�-0.Gk�,�	����S����iʝL�`�G:��u��{6u�����7:i�Z��6HE�Ϫ���ⲋk!R
o��������Y0�[�@�m;j�4�o�-n��Iҷ��7�r�=�]e+�|)��dKC#:I�sh�W�8��S\�{�:wLI��2�j$��P�{�Wƛ:����<M�3��m}�}�&iw�y��;����a��2�U�w���
��r��̟���=�Ҭ�����8�U���'��^��kn����v,*q����^v��52t�'gS����C�A���7vh����}�T��eܹ�q�`����ѹ (~nɷ������5�%��s쎧\q���v��i��`'���E7C_1[>]�T�e��$����*�z�<�|-�?q6�<>��3`L�� �A`�nA���Z�
���{��O����1=�{�cgCg����z �߾)	�s��NyE��fC�w���a�A\����Mn"���,wK5c��}�/�;}���]�6s;�,G(NL=ֆi��<��;�F�$ŹMh��� aGO�V
X ��?��dx�
���s���r^s�%�%�y���_E'_#����?��+S��[��� �-HN����
�R��FJ��|������`�bU�ϵ���a��ׯ;��2� ^�'�����UɽᩗծH�8�4�<+lD^��VK.��+�!6��K�W�X�J��F�T�� ��7����n�l2������`x�XO;]��.ʪ1�]߬��q/ s�6F����́�R"�X�d�7�#���?�}h�KB��������u(�s+��5�t��MF�a�ɝ�]�S�u�M7��=q.'���Ğ�������r��w��s=�p��OBD?>l�AكrE�/p[Xy��Q8m�E���bĹ�!���I����QVN��T%�ҟ���@;�n`x�P��VR�.u���&Lq�������8����x���s\~��T�����^Vvr�K�"�s��5���_K��ʶ�-N����Le`9��U��,=b/�%���DEk��tkb��k),z2O��5ڒ_. ֤ډ���N�U"t����,JR��c5(
#� ���{�+^��k�c2�͝G���ai�ռ[����r�kh�P��>���<��,��FW�(����Z3�@�k�1�U��D]/�) Rڻ�ܤ�rYu �א���=#u�nZ���S+!@��#�^`
-"8̯�Ԯ~"��r���خ���$����0.�	R��odq�+��I���h%���o�s���_[�*�Ua�>^BP�
�r��k��~���[����>����s�q�˭J6��W�O��U��W\To-(P¤ң��!P���4��\�D+���\���T���Of%�M&=�(D���l�tE�i�yPc�h;碘,��S<�-��gP�����:��BC�V�E`pз�#
�uB6+WRrƍ%��)��~~�7,#�š�����0����+��#\$G��4�����4�+/��R������	�������cF�k�*�:�����4Eb'#3z�}Ŗ£�5>=V���	�dW�d��Ik�ߔԢx��<�\`Ј�	V���V��6J��d�,K�(5y��.�'�o���fK�����i����W8�<��,ZwM,��T�f��-~׺��K`7��Z悔�)���A��/���bܸ���3w�IQ�G@|��.��G��W􏬈Љ I��Xŧ���i7�A��{��� C$���ۓ�u��$��F�SZ�~��k���i7~�σ�Tl����p�3�R��6�ra���1`=�=֨y({O1��N2�Q��L�_���@[�:㤅t*�;[ L�iQ +b���?�s
(5�8y��]#L�y���,U����N��`S��jz������M,��s��d�m)�/ys`�gn����l׽��|h\x��FQ	�\#��7_��i�l�Q}G��@���c����H�#5� �W�x��Y�/�q>����"l\L��z+˞���v�I�*M��l���H�T�9-�c� <�Ƃ|8}�'��d���D+�7A�Ԯn W�^7ݓԨ"wΟ}��,6;C��J�i�J��ȟ�>�>݁�8�V�l"Z�ݪ@;������&�����qdJ��5�(J,/'�^�wDQ ��T �,����lm~Z6���W���]i�9_��v��#���X�^ΉꘘZ�`L>�[<�8��#�Ƈyʃ�1'�鶤|ֱ:�O����_�����c(�w3�w�1Q�i��;�r����k��Q+Ԅ:��|en/�R�C��"�.ب���|����	b&� �xH��(k(/�<�9�Q�i�Xa�h G#�$H�,�w7������#�	���u�j;}Z]��n�&h���7�ϫ:C���5����RE֪YY&pIS�k�@0���2�p4Gs�������>o� �pd0`�	�E-P�R]|cr��mEy����Z�\�O�������#��%&��!I�cX�~oh��|?`���i@���T�5�o����u�O�����_ߑ4�b�����PM�z���ϯ���h�i�-i���<�;c�Y�D�֘�R��i�!)|��;aC�lw;����dO͉��EC}�8��T���I^��RU�͔D�vIh�m�h��+��S867���a�V����o���ĳ�,�BN��u';�*�c�%��ASc��0|`��m)D�z
��b	�|��4T����3.Z4� s踯x;�eW1��c!�,5�ql1Зد�ՖЯ�DN�RZǽ|��#x�$�� �$8=Ą���b��?,d5�AkT���a<���?�G��U��%�)M2�@�}=��~�e���?6�iNէ���۔ч��Ӊ��@6kG��l�>����>vհP�N�?h���kbw�����=u�l�����5t]Zj#��l��>�a���a���{H��Dl��"7�"��0iB��/H=�ݶ��#ޟN��q{��!T^os����ݦ����o��9�
c�qq2��k�c��l;�O�6�w�򷍲kqڿl�� )�ׄ>�@w��k�\̼̾Ǔj�]t�;������'�Hc�	�,�_Q�w6aQ�R;��tl5�â7��12�ڀ��]ڇ����g�mM�ޭ�_D�=�#\��cE���ḻe�����2)�x�5K؏V����VzCF���ZF��*��5a]a��#��r���&���s�D~I�V6_��!@GY���7@�pV��T�����W���9�:Rbo��G�|o�܊��s�o��~�@���Q�V��殢W�:��̤LZW�-h��Q��*DE��p{�Q�z�"�ǂ���5esv�e5��ɾ.ͳǧ�u8J:p��p�*�R�*���RCj�T�P}�>�f$�+��]��Ѧ\Q���<���A�	��wة���[�G��w���P���W�U��?����~�X�f�T����z�.�r:k_vo1�	�XuAԱz[����^���m�meÌ�(���Qrʵ'CBG|5��v�t�<B��(%ς.ۜي0qH6�&���/ȺŌO7r)���f~_����ŉ��ϊɊ�m�={a�?S0n�U���g	N ���o��w*?�Z��[�y��G��90�w�I9̼��jn�-d��=�9��{��l�gj�JT�~��SA�]�egr���ܜ(����?�cR��y~N�� ������ǆM����
.����nƍ�����C�݁�Fo��a�6��26�w/��3�bB�.*J@�%Ӽ�3'%p�%�\�� ��W^U vS;i��'��@dbF�L�h�^�Ry������ a�=��t|�.o�4��Ɏh�BF(��8�����	�ǭ@���@��o�^O���?��i��D�h)��&~V6L��rr�Aϗ��%y�BrB�s�l���'5�'-!�E������W�*W`G09���4�������� ���ė?�r6��N�ꣅ(�Q�2����s�9�����s�\9�	UM��/):b��Vxb�5!�w��7�C����ݟx �֟��Ij��	]���6�Bv������#�棳�Ht�:-ӏs�jhE�/D��n0¥UW�>�'RZo�j��[�``�r׺���!1��1W]������.�=*���0I`��\`i��̈́���c��EM�A���`ʮ��GT �C�G�f3V�?��TÉx�O#�k97n3���e�J��@�G��;���~��=%���H���6�G�?2���N�}S�`�K؂ъb�HŇ�p�kmD�1���a�1ĎMo?��}cD��2�� 4��1��$��Id��ak���1N��>��+,+ћ��S�i����6��NM�_�$�`:�.W�Մ��_S4��Grs��jX���:����=�pF^y�����u��y��E'���&h2��r����uNVm�o$nH�ЬI?ԅ��>V�wq���~-Q��*�Y��ֺ���7��|!� �z�hP����-4)S+3ȿ^9�<�E�}��;��M�]�&Q��L�����lXy�sh���_��a��3�!v��������C�*�/��q��d�i���3�]u�'tt]s��D����m��.Ǹ�����c��F��:V��=}���c��ϳ�ݯ���lɊ�n��d�ں�3�ur���q;��y&n��G�[%]��q�}���H��}��D2._P��t���x��vo�$c��������Tq�����"��P�u�ؔ��q�N͵w(iU�;��6����<z�7*gv�&g@N�x�ڰT'-*9���m�y~�w���w����Q�S�o��*����h��St��̼�r�Y���~�Mkһ�����/f�~���i�~G{�[ۄ��QǺ��$ Ei�q�iX�pd���U�tw�T��(�K����5��7+��A��ǇoՁ􋒃@&�8'����4�B������<���5q��ʍ�_�����g�c["��E�̖�:�T(�.���Gm��AЅ�H�%4l�"~�ԁ��i�YO���s��d�u��7n"kW�o鿱~�8��V"Ű��Bd��4������UMP����ں�U�`�f�!��Xb3 �*Xx�fB��3�?hB�-��,C��m��i}�a���6�G7�<�B$�z߹
�Ͽ�[T{����\Cq���O,)Lp�/J�z��q���ʕ�l�I�?@���n�C��by����ox	w���^]>w�.�>i�|�i���1�?�Yj�V�;e�>
[3�e"'��fð���l�T��k�Ջ~��z@����ĕ���9���a�iږ���K��,a�G�Ϡ�����'��v{��#���:�n',�N,ޠWT�jHn09�v�whꩢ�/����2x�� �J@��}�XR�k�!6Xeo�-� L��t�Fj/��l*���6�����MK2��L��AJ�ْ}
�]s�Q��Q����Z/�:3(��I������JОΏlP�L`0���(����H��M뜨M �)^���D��s~�i���]{93u��U(�����	R٘��>ꧏ��T
ש�`�^��~�GB�S��[����nۈhƫƪۯ�h�6(f��ΰ${�E����g�y�*�"��^OhT
	��%��]M����=�e�F%��hMX,���U�� ���41�O�T�g��+�pS�z��Qv�-,�/��Q��=�c)�{�"�x ��p0����V��'���Q�v2{B񸡞�G;��mu�l���2@0`]��������	��q��:01M���]���;g����@��t�7������P1�T����+�͙�i�I������FK8�jd�&(�-�i�1������/�
�څo�<<����. ����#MÛ�ᤵ��aRs�N"?�	�،�3�4���6���y�������)o[yo9�C�X�M�eؖ�g'�G�c2�=4Y��'ܤ�x�ںe���5�OӸ>�+!�9�e��9�P�glB6�n�x�.;������H��Ĝ:��RL�{�Jhog�/3���ڻ�a�0M����z��(�U�i=r��NΔ���cxo���&��|:����c�2�4!��܉�jʭb�1��Bfo�.>���������r�"��ߟN�	Ĳ�v2��A�u�Ȓ�ebT�E�މվ�7��^/�?5f�!e5���fH6ZGK\�υP;�j��5��a�*��"�|��!2q�Pct�����e6�,��+hdR��
��A�����/�q�:���&$t������j)0�������<.�N\5��=Q>%��H~��^�T�p�F�	^�`���;,��}�;F��^Ϩg�e�@Z�<�[�3a�[�F�L�VFF��.���]`�����KB������Z,zѴ�+���u}���AZ�<�F��G_� ��Z-�d��F6ߌEg���?O�3f�ۙoF;�����cH���lQp���T��;�7t����̼��6v/�KKh�~1K4cA�i�	��b�s-Ŵ���kc��������
Eez�-!8_>��lI
�<K1h�Z�$ֶ����;��-�>�'ѕs��H�VaKo�Eh���6?D�ݒ���qB�B��>�2�~'9ȴ��������W�= r���E���.N"�o�&Њb���(]
'��}gpZ�L�ω�
{�{x�	�ix������I��r��.�Dg�g�8�D��ؤ��s|�r���k���}�-�Pγm��+	gu���k%?d.s���)�d���D$�1x�U�lg.�Vk�V��%͡�05���|@FDc&���+�g����������
r����%ƝS��-�����\�B�{��O���*֑i�۹)���RI����(�	x*����"a�F�����H`I��f��V� )�9�1!	�n�j�e����I��a�R���:�q3S����q4݄0�)c]q�{�C���p��FJ��cѪ�����
-��G��J5�?~�O�p��z��y��PU��p��k�dvk+�"��
��\A���o�����(��ÿ�h#�F	s��h���i[S��YdL8Kv�S?����-�b:�"�&�����[S���2��'��k�����x�ۇ��.Ԓ���4.\z̕��赊`��FK �{��ЍY���e
�������KeU��l�AaK��wTx��m�y,kȷ�"�\[�aݓh���a��|�x�71w�"GD��6�]}�� =��~�����!�m����*�/�#3��R�����{4��<.��˽�l�X�K�th�'KbBH$�����1�U��`H��_�� �C`�w��eS/{z_�gJMm,��s��LCF�� $ �&N0T�����з�"Z�2���
�:��=j��GI3��g��q�eEC63��%���)���6�3'���]��H���8��Z�*�+��G�ۤ_��u$��I+eے�]�fJ�"kyW����TQ(W�+叭6�kX��ve�F%�-O���@F��&�n�^�����z��o��'\�FF��QqE�WP"��Yl-�z��i�wc1!C eU-M�S�~Owꤳ��.�q��Ϣ3qR�3q�HQ���u�����3.�S���h}�q9u/�������m�듙�L6Ol�2bKtP,��,0`���6�>�S/<S�
�(�E��q%ځ2����j�ޱ�́&2���/BdP �?_T�b�G�=�F���m�khl�+��p=��.���I���!��n��!�4Z�.0��X:�
>�P��X�z\�)���܀"z"xD� "I�]��X��&8��k��^��=�;�����KF�R��S�2hٜWþ'��*�2�:�4��!�H�P� �p9�����ɳ��	�%���骱������蹾z}Ș��F����)���僩��I(	H��4�Q��&���+U�����6�;��B8��V⢖w���g*ն�. i�$�d�!"�F�q�"{]w�(8gɜS�] ��
z���pJߺ>�I�ް�)Qև6��<O����-/	�h��Y��˂�`u�*�Xg�I!�����ֱd����J�/�����AR�V&B;K�����f��'/�*1�w�t�-�T}��>����d!����~@�_��gbCd��7����:b�m�z'
<U��j�H5^t6�
�H�q�YW���53�?���vw����㽂򯕕P��C#�O/b�{��(�NmV�4��F�����8_���W�D��I��mI�%�������]�=կj�4�p��ch�w��ke���%e�֛�Q��C�'�X�^8�A�����Ƭ��sB���Mr�՘}(9�����kEM��1��� L	�m�ӉO�:{4�ݻ�n�O��S�ڭ�9��cp�]- W~ً;%NO���[G�|�7��!
1.�Y�'�n�ySځ\^�B�{`�kU�a��?Cl��!�t�$X�)��w,��ˬ�%���S�!��b!�Ŷ��[m�|�_�M�1�+Z����<���x�p�a���sa@��E�� ��2�%�{�@&�-��*�}��	�t�-�Y�#�.6�q��F�$�U�;����y'i��(��7"�}q�&��5�I0���'j�ɩ�8�� �
E���=�ug��)�m2�y��2)�/�� ��g�G��f�7㚺��'&Lo-<�M��f᫥���{q����]?�:VP����QB�E�Y����i�����YV�[���WJ�d��]��}���ϽƠA���B?-���M�\k+�D�w��sɺ*�|���_�:Rִ���ѱ�z"������O:G*b����J��rG�Q{Α���Z�Β�9���l	�z{����Q�[7��N3��c�}��
p*����R@\�����D�/��+F9bN���J��3�ވ�?h�r�m���߃(�Sx����N�)#��;�<\翔I�-����v�A����d�����O�ͺ��,etobYP��y� �*/D�E9(@.�rrr�B@� +������حڊ��?ǖ�L�}ݚ#odj��-�d�H���"	���ƑH-���)�+���s�0�DՔ�s���fe?�����E9�'�)���#����ދΔhK�
�z��!0����E��^����k"䵆���/h4��Y�ۺx�G�Q�e�ɩ��:�N%p;�DO�Qq��c7Qj}%윐	��J��\���&�,���Mb�����]���B�t��CF�c�K���q'�L@`n\<lg�+�w��I)�@jW�_P-8�o>h�;\�'E~Q{�>��L,׬<�6���g��ɋ<bt�K����i����LՃ�i㻟�E;�*�b���B��;0�uW24�#�������ќ�Avo����H��gl�cN�	ӜC�=���̇3A�����~kI'a��m���tw(�EuNAJD� s3JK-�f���2�wql������O�����u���i;i0 {��=�M]{\� ǆ�����\o-�ф�N꠹����M��{I7_<z{����9;��Qg	�/�gV[x�R�N\��D9�
���ݯ{0�5�N�ܷ��� �Yw�[4�W���Ӛw1��k���W��E�y��c��C�����.�s�a�b� x=qSg�H� Ў��� h$�mP�4M�V���y
����-�����Dm����? �?��4&Q�W����B.���\ôѸË���J���z��pL�Rrٖ��4l��p|�gR�����9ŹA�%&5~�!`����f-�[%����0����Uh����֘�~��0]O�Y?�A_�7���*��Ʋetv,�������Mf�-l�t�]�����Ӑyy7�4H�ew��]�]Lݣ���p��Y�V��A�V�i��^_��$�ǈ*p�+�i��݁;����Ν���q2���y�����l��[��KQC�S�NC������`N�^���r�m��Zf�I��gȫ%���E.�v�<�I�A������
SM��8��ƨ1Εi�l�i����o;E�)ViKc5�v�+C���x"[�pn	�t���� �q�t��Ad�|u@�M޳�T�$�
:��R)I���)�ˁ�zG �b��$����(�ҫ���4�@̧K�,Wu.�;��n0\� g��̥ �ו|U����������[_Qʷ�2q��I�0�*���;&�ʔ1���^���2�TOB�.c���٥��a��/J�Ǔ���$-n	��ʾ�5��Q�����|�E������Bz��v[)�u���mx7;��O˵�	9N�aH��xL�� ��0�Kp�H�\�`����RQ�a5�v��T$:�F&�3*�du��C����aLRE��,c�އ�p���X�Fr��E����j��63P�hɽ�2Sa�'������p[������Jkr�}:a(L��t����ܑ_�(�$�{V4�1�Z_���V�4=n����¼��X=������ �|��O�|�ނŚ�F�:�p�$��k��!S(?'�5�B�<���4����k:W?��������{U�?\��A�G���DiT
J�['y��I\��Y�M`��L:J
S�D�r|������p�%�{�[�ъc�����}�,�+}bv���^�z��ml�J��d�,S'w���4h
יS�/
�-9�����~7�"*�0�ڐ��Å�8:Щ>F$A�h�^4��4��%���2�.��� ��S7��ݗq��l�����&i�h�"+w�ձ���,F|CГ�,h7:]x5\B��"�H�g��;4��;��G�_���bc��r�D��4����p�u�^��|������B���F0\:�&��5]�-Q4kZKW���C�*=9&��P���?8<5��)��#��l\���O�.�ĽN��/���%!Z[`���+b�J���v/�D�8��	(��.��4�C�g(Y��v�|�.��PY���}�m��_�Ph�7 ��3�(���!'�9̈ν(�S�=W��6<=jXuYU��ǩ���3Ak�P��i�Q�Wz��`ݞ᪗-�V��Y�`�o�g�g�JT&�����bLJ�����q���O�9�fK�1Xٔw?+�m��(>Q�����҈�	�b%�"Rt�\vދ���O��+�n�BgJ�L���d���=Kg;��������~b_�V�r�>�Z���?�_�e̡���l��(`�h������LgMB�������(D�1��9��ޔ`Yl��p^��(4,��׾��M��.�n�����d�N�a��(��ȪgSB�#��>i��}?�SV�/Jb��2��*8&7�>f�j�'	��j�B��� ~ =N��$)��,]�����i�na�r�c�ٚ�"�"UP����L��[|(i���r��+����4�fg~|������I]�j8d:\x��i@�GG͑\Ž�]�\F���E����7����J빂ՠr��Hp��u�:��<��>.�qR��l��1孍�}���$��2�|�ZS��7�Z��;�Hd�RD��Q�R�c��T���.�,m��c�D��vsZ����n�`B<�{� -s젱�
� ��"����[� <��+�.oD�qx���u�#���$!9��ڶ]�J�ދ�5�(0��ņ������6��D<��C����ѯ�\P���
�"��3��`���ƌ�i\�R��Kx(�]3oo�5j�u�#(�ɍ
��R����{��$F�-e+|^j<�g��^R���		�y�e7DQ��`�VCҋ�>���Ӛ��s}�����佟���&�r�F�*����DQ�|X��	����LH�S�rʐ\"x�M��X-�*C�yr6��M�t&ơ�9�(l��gL@WJ�$yd��_������x��˩���R~~'�E�A+6s{��g�2%O��d6��9\
��߇8���a����9O�2��`>�<��Lc&�rb��eq ��o�������{��7���DU���T��p�{8W��X��gдg:ׄP��j'���HP�	1N�6��a��`hg�"�6�pX��&��8����u�qui�� F�2���W2����,�d����y��Ci��w v궺�ͤ��F�0�bPj:��[�GFDI�-hM�:m�v��>/�H#5¼R�CՐ�~'��'3Z���h����F�È4�U�s��2�xG��LVQʥ5��;XE��A�`�N[בa��D<�R|���������%l�6'��fխ嚥�⍼�1�<�噞��t���_8>���n��(L`�6k�'c8U���9�sv�n8 �K�5�����^#�������	g����>u��0�!i�����UH�?6� bHF��-�G$U���4��u|Q�f��Fy���f��4�Fj�>�qT\~f�Y�9��	b/�Q���2�x]���������7/9��B�|�A'��h�1o���Z$W�� �n�2�&�O
�E4�`G�|l(�c`-<G?>B&�`��TU��������c'�t��R�*��y�p����q��q6�`����x�oS�OZ>�{�k1�9~g��WK�8����Cn�ϵ�8]8}#J�^R{��AyVc�zakp�l�N�O�Z�C���'����|K>��l��{}J:[�py	� �^�h�no�,������)�lI�����g�`X~px� ��]�>&�ښ+�c�L)ͭ�
ؿ���2�±��N�B�N2�{1�|Fs�xy!��`�P"��IvYd�o, �*�J��	t��:�Z�1 ��S�*�ap�;�Qpт(��x�%V�4&(�ЩoF6�yI��X6HJU0e��S�^NO�vL��Ae�'�'YQ�R����Yb�O��%W/�X#�)����:���~��7l��<e���p�I��h�DeT2��/;�.^�{,�R��Ў8K���bִ�m��s_Z���A�*eJ�����`q*��
Ю͹#��.�D��ި����8���t�JF�l@�)��tV�I�޶�1��>�ߪ c��q�����Ƅ����!c4���UY�c�[�_S�}2��~~��	�����|{	�ohu � �o�7T�6�+9R�@�� ץH,���K�
���B��1�09�ӦH�51n�Ċ(H�:d�) -����4tw*�ZZ�R�S,��f� �� ���5��GH�t��F�kπY&��,ya�I_HHZ����9�zVf��Ca�#U����P�RJ5�N"��!������PBW�a���8���I��1��.���gQ�&e� 7�1 �<~Ź5�	1�0��w� ~+2���N��#ܜ`>oR���K��G�a�t9R��w�x�ߩQ���m�>�c����@2��yZ´>�W��.�2�)����w�<��0�J�?5�0��vks��I�C:)v<3�Y,>$�eP5��|�J5�Y偮Bť-˺߱�2���K�U�Mc�|��Dn�Jn"����pF�3�9�ѥ���",S:+ZcY��8[������W��JE@���9Q�U!�j�ش^0M�_�A�Y��O(���5֤Xn���B����:h!͞��uO�:��dÎ�,�O{?S�ѱt�)��f#5�}1���M^5�B|�[A��^=!Ɉ�v��1�.+y�{s~�p��e0�e�<�x��>��ZtJu$%��a��rZ�g�q��@4�Yɂm�4S~�9ˇ���
�t��V�{�|s��2����β���A�) �&��l&��k�U(�E��ԍ �F���͇1yr�X�����IT]��ZG1C�1�糰����Ys�gz�L���~lP0�?\i�ڔb��{N큸�jZ�W��}qy�ű�U�s�>�L�Y�J�c�<����<�$�ٞv��"��E�a��kae�)�O����OA����yuaG�����>��=���A�1�ѹ?q��ΨU�y�|'uy�;�;����.5�Wn
���k�%����:pC7F)�F�QZ���PK�$D�����Ξ4a<��X��m����i��пK����7�A� �g�r�F�d���n6��Px��+���-،�g�kmSt�zu����} k�IN�iR��������(��g�9����W�JW��᣷e���oi�u�C��7	�/��~nפ�A5@�p#C)���J+O�n�A"�ïs��t�V�#��|qza�^�p���<����$���B�
I�C��!#�Y��eaX��Mg*+)R�Ō�/��fmeY�
��w�G|��!�(����B<!\�S�d���)���ҙ��c�0sPe�ӯ�O�?��pр�AvKl�<�ϝ�4��g��b�$�bs�++�Y��^�s��R��<��m�;�Q�!݉�vZ7��t�G٧��_{f