��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�������s�h�qQ Ҵ�pp%�bs�!F1���|W��ٍi�\��չˇ���7Ge�+��9�*m@Mm��A��/f��XT��݌��GP�s��Ɔ4)c��f6�}jwS�����r��j����Īf�t�8J�gmdD����I��h9EWC0^����T�
�we�g 7H�����2�^/����t��PY��Ivs�b�q@>y�%K�~���*0p�w������
��w��{R�8u-C���_f(ZG��|���/zg��P�sIY+�e���<8%���⌚��8gn*rp,����_{���W���J��fM����D�~ۂx�Q|�hCުŶ�_����[�����������=�՞����6�����o��B�#A�����4��5s�32.�^�`�!c菂Q�h�;�wטvm���Jy�#�d�d��_ǫ&؁�	_��8q�,e��e���O���<������э	�gS<�U��� hNH8h��]z�R�| ��1�%��N�G��L�f�e�F�xO�3�]_��	F���� :H
�q�<* 3��j�6ԩt��/�I�?��S���9�Z�p�؜�'�����h����ȫwմ��g�FLs2��r��|G���>��d�ڙ�5���>g�3��ü<c��y�:ʑ��
�pR���+��L&�g�j.~Ǻ�$IR	����4t>�w��46�;rc��[���P��k9�5�I��Iʈ�+ZV_=�$Vj��rx�����>G<C��K�J:B����e5٥Gp+���hJ�Q9�Rc�coF�n��o��̑��3��e�ѱҎ*Q zfc�f|>7���z�`��]���	�d��=S��]tppiO��N��ѵ���_ ����_}����4�`��nA&vȇ� 3��<�XG�/�2��$a6�^�.���=-QR�h !$�GM~ Dw�2u�lc�P�z3Z Α�:H��#	�i,�*�<�κ�{��=#J�00�t5�a׼F���},B�+����$����j:nx'N#ݽ
�Q_ξ����Yw�ޭ�1�E�!�
3�e�,�\��u[�lw��#������1�ӳח.vt�_,.	hk�QƯ3j�AhE��}�=C_�c�K�p����t��>7<�����k29xx�%Ƶ�o�JT�i�0t��4?��� ���v�z��ɦ��k��!8�J=�X�y��/}�ksֹC(���˒�N�@�$K	�ڂ5^��)s���,�bt?�S�ˬ��*I��k��a��\z5��P����[6�z�9�-x�./<�$�X&ǘk�F�u�=�&�Gx�w�+P��-�QV�S*Q��KR���EW��x��ِ�#]����x�M�8(#S�2?�s=j�Ѕ[C��hTB�Ɵ\{��vz#sd�hR-�'�R�0ԅ��5,%Sn);����z!{�>�aiCŐ0��F�7
��3n����_���� #Ä+�nO���;��2�,N�oS=͝��
e�	��@�	�WE����L�~�q�����'¬��T$��S1W���y��;���~)�[��CI����x�+�e��}Z�x�Sh�ag�Zb���Z��!$]�So��#�~-�����~���Fiج��tXeX�ԌAn���y%�7�[�����E��I(��0�Q��eXJ♓k�~D��l�@����W;�����`i ���lE�q�� %N�R8��yz��g9��[5n-s]�L�nJ���3�G5lnhd�M��PK�o��;\ģ+��/���3_�98��ެ��޽Bɮ��5�����;���������>�:D�mfHG{�?���f.�0*`\L�{��A��I��@����eݧ�(Z�Ə(H����� ��Qk:����I���=�6/�D�D�-SF��a�/��Sm`0b-�ظ�4ݵ�[娘g�P��Z�q�t#0
9��!u�]����i;$_�.0gDl(P� )�(�f�¢��6��!G~(0���o;k�p3c<�d� a0�nw��S�1d:�2ϕ?؃��_~Қ��*��n�KobJqi�z1��dԤ�����V!٭:	���8lPh=����ц�HS�Br��AG`��N7�����_���2������JW����mt�1
�7PQ�Wd�&ƈY!���o��4�ϝ渓6�� ���c�ߥQ1�9ꐠ�����NF�Q+gLx��Ui�o�|Lv����|ް���f������Fg�q���B���z)?�27�ɔ�!��*'2�aD�͋k�7O�)����_������g�-Y"A�)C7RG�[���M"1s��/d�d�K��C�>W�� ��;K/5�]����L�0Xp��0nL�$mb�<���:~=���7���á]1��;�u��;�F�?�%p��0I���|;�`��>�j�h�mRoC.�ؼ�t'�a�CZ��+y�C{�{y<̊;���[��L1�Icbe�AۡL�n�<�{8סu���TVJ����{J6�P��-l[�0�e�w�;߁pq����������tFT�7�K��(kF�eK��{f�k�Zz#��)T�i�gO�\��UL�ذZt�w�j��=��-��ݫ	_�F���#�z���)��
�zTѫ�x��� ��!5��a�
��: ���<Ő3�
T�}�^H��h�T�b=��,�Ԃ0��k�T=�1��(9��(�yɢb����5�R����I5:�ȃ��Yh�G��Rs':���{c��}��\��\g!��|��g�i�+z<�l%PE��$�[�*��I�/o�!/�]:�M~���z;�w���T���%޷~/(�p3��MU�!�٨���=��)��ቚ�}�Yg�6��$��]��cTV:=W��n�)+aN!��Z�fg�ƕEӰC��k�����o*._?��o��w�s���wy%�~��Iu(O�J5LU:�t\��f���\^��vp� N΋!�C�B��h$boup��#5+���h���<�U�E���A�t����4��E�b�Eh�"˞M��Mg�"�nd�'d�C�fw�@bg����#8�#������}��0i�o�Ѣ������O>�ʸV``Ҿ�$%����(w;a�V�G��<LH�[FƯrG�m=k�)T�fxe���Wk�l E���T�@cG�N�ɩ����_v���N�i��0�#��M��<Wj҉���j��y	pi�����a��z"\bN^�gaQ�+�>+� ��t.|�JZ�|n�j.�2@�S-Zn�(`�6m�� ���H�A9Q+��#���,-� �ڮ����b��ʹ��o֦]�2�4O������R�=��=�l���~xL��y.~o�OVv���5��{��6>����*�Y/��<ZDn����DA�d��������l��]?CY�Vo�%�] h��2�а���|CV�T4@��4�X��`�&�`P�W�-��H*Xv<���Կd��9cӞ�����0��6M��ؽ%�?D�v�ج��,����Y�Y�`�W@�F�&���F�G��������Y�S��46nd'C�3P}�����k(fV��`j���B��X~$KG�ݔ��P��D���z�XL��.t �yL�f�Ⱥ�������E�ŦK\��+���V�`8�Ƅ����N��e��l���u ��o��t�W�1��ƈ)�3��f\ށJ�x� )X�Q��ޔ@�w���@!e��h���2u�*�E�|%��c|64^_0�� Ɉ6��H�]��R��`��+Z��[�@��ƴ�E����GZPZ���Q��\hO�aI q�¦��e���gP͊�d����=r�r�yXy��+.qX׌�V����I^c��'�id�0z���˄?�R��ޅ/3h�l5��
�En U��$6lB���3jC�k'	��X�)�\]�n� �~>�T'4:o�9h�v޴^��d�d/�?�T?�>�e�f-{g�����Ty��fΟ�bv�͊~#������
R��A>o _c�0Ac����ͦL�/��vydO^[�[8�b�J���S�O5_"�#�)`5�Կ	��^��d�y;*O�w*�����g̮ʔے*"�?���R�73���&VC��Ο�ڛ������-+>�*P�JF�::�,Z��5]�cVb���6�^���IBo�q�(&=�xu"fo�[\���±��.y��9��6�����_��ړ�0��g�>7�8~FʁҌ��s��%�vfǭb�pɃ�p���ݯ.]=� C�9^��hbb�!J�n�>���M�8C'���ZSTtAڜW�:�	��0p��"�գ�������s�UD��4�z�r�GrE��߻q�k�CDCƳ[��6x��Ք���;�K���w;�3�v���D���Dnz;Yw�i(&�P�MP���|e
T0���W�� �G��b�p�s=�M}j.v����
�w�P�R��MA���a��L��YN�i9�gR�P0r<����E�vZ)���^�	+���r]�Kq����Z���z ��I�*O�V���
[�'���ĺ�B��ާ��X�V�h�$�SKu��ɶ�TʰO1jm�*�ǀ�s�O
���j��< RP���Ɨ�\z��V�q�� ]������T�,�v���q�V72��Sp����Y\�i����[(��)��3%�d�=\r"�{����k���._��K�m��<&����&�4#\ӝi*e�{G�M���k�8Ӫy�L�Y����NС�i�;w`��T�0��c�����39Z��.s���d��o�+�]�ކ����L��!�TQB�X����r=����d�Mg��9����1���z�&�����LS���܁���Y���-*U��u8z��P��0k�}57��$���awB��Z�E��^x]�9o.:��@�X#ѣ�6to�:S;x�M%��=�*T����89�@�KPK)d�n�,�J6�H���c|w�!3����z�&�Qv�*o��Ԫ�9f��<�#XQ��w�[�c���B��Ԛ]��6��LD�y�,>����7�+���:��f����Ƣ�a�e�vC�x):R��lf�՛��?�o�``�Y�S�'����cr��AnS~ȣ�n'z���a�l�s�N��gUl�I�k�,־ �s��WJ�악��nxO�d�.	��i7 ��j'�e&.��A2-���!{o��tbkH�JI����I���xs+�7��V/�x:�¨�~���V�����b��߈�H���2\sѯ�o���A��-�U�2�4��`�]�; ���;>�u���y=*]�d��I�����7�[%��]�P{��׀@J�4��D.���Z�kf:���#(��]�+E��x&^[�~���R���NBe|+bi���D����Τo띾���h�(#��l�(�<� �Ӛ[:�\ezR$1��.R��-�Z��^���"Xz� �m�T/՛��E���G��%��Aˠ�LJ��I��(;ō�fj�ۙ���y��y���7l�b����@�)�TJ�dh��:9n��F�-ԖT�%ǜ4}��6���4������!n�� F6�L�(L�d�;��E�YZ]�2��-]����6i���'�T��������CQ����ִ� �-��T�c�@F*�Vѿ_�q�kr5
��$��$�G�ۢ�`�Y.ّ
������^�=��u���a����k�P+�Y�A�g;뒔`�_Vf}wC�l�;��%�)]��hz׿X�H		eM�czi���m�Q�#@���lu�m{�kg'�f�����"&����ւ]=Xu戰홈n�Z证���%���g��z ��}��a[�a��"X�5��D�¿�D�������t����1�M����*�g-E`$�9\�톝ce����J�"T'@k�"�na��D.X��*���g�E����UA>�U��$v6I�E�r0�EL�����RZp�Ы�F bVW�_Z�?W�����¿�FN�����:ȥޔ�V�����9�~�W6�y/0�(��k7~���򠘜�g2�P�B<뢱@"�x���[�b�����V�;qz�)����v^��U�zs:đ	!>���ˎ[�>M�\�r�B������i�:I��'����+��UOYR/CWUV�q��\%޷:%S�[�R�m�Mpn9��� ��{����>+�����7��M���<5`���k0�n�~S�'b'/�j�!��)��<aݫ�B�
<��?b^�Q����2�M0�KI��}wU*����T6&	Bүcň��o�=�]G�%۞�"m�-�M��n��� �m��B�o���ҁ�~65��؁�:x=z���պ'���pm�����7W��8�\�C�2v`��/I�M�"O�DmL\�9�7�B� :�{ƚ���}5���>�Q�S��S���mpg�aj(5���a��,�d�^P�}�D�P�B/ �m��	�����؛6ڳ�V.�.��ų���$��e��安l���C�6��ژ7��Z�c�i��cO �߶A�8�յ_E����FU04��SvA�������K���§���}M���bت|��a���5t���F���8
��#w�QG�nm����O��$qsY���k5�6�.�u�u���t1���-�5�������.2�g�SE�U`���4bV@�}�$ҋ�ɲ9�I.1���0z�<���#zR���W��a&i����p�Abd�e1�%�&�ۑ=�*Q���tj[m�O�}�-�[eޢǗ~�6U��Eh"c+��6kNl݄��I̻�â�ӥ�{�
���J^.^?[��v䘣��_��5��_ �@�hD�t˂艏�Z� �{QDq:���o"�+'bq���G���B�Qh�hHD�C��`���)����;ǿ�I�j�h�S/-�-tFYk�Α� �#H����� :[0	�۴���!�onE�����/U�?m��y��k�K%�mS����m�'ꖏ�_�ʗI����?wgn�^�K��f��^��z�w&*P�J!f��sGft���r��g�9e�	�6̟�-K������YBZ��79*�5#�� .�m䗎/$9D8tO���:5{I"�/6���.�D��}x����X��wk��v�����s ���E��H,�;�����'������=�Ǔt[� MK�s��9o ��ZW�5��B�1���j��G�*j3GHk�B�<�#�J���:�l��V�k��uc�r����թ
ѽe�j-x������3����T���Tq����$�����Tx��mT�Q���oCK��4qG��I��3�m�j�,�|��,��L��yE�7+�\Lr�+��H�9�z�e8��|�oLvJ��ť�`�7�"ƻM��/h�� �\��Җ�p=�7�6��^�j#�a�^ȘdH���|Վqו{��A����5H�Y�}�3x���O)�}YnX��̢�껟;~��N;�e���Z���0�{�`5Ǔ�e��3�#�k}
v�2HQ�0VnZވ|�R�\5��?}`�N��/��NÔa��D%m#C?���F�uc�������-�]�F)����<�
�	}	;0��%��5	��-���mn��h[��F�ٹP����Z: q]�tq�cĀ����T�Y{{���0z��.�T\�V���n��TP/"��1+C�5+SN�8��@-W�}U��h�O�a^�2��A��W�Q��	��\	{o�R����_Y5Қ�Y]�D�?ٔ�ި�F\�F*	UF+��������t=���'("�w��ο��M�1u$��IA�|i>� �;*�T (�Q�(��e�b������L-���*��.p��L<�c&Afe�ΪR\�RIU��Z����zV9���R���:.63y+>�^����"�"�8o[K+��kn^�
�u�6^��}���J+6�(b��^��5�6�R7{�ͥg֯)���?�{Aj�;7a,K�}O,�[|��5�̤�$��:Һ>����
���#���^�*ߊ֒�m���U-��Я�ğ��F=�v_S	���ę���u�2$(�G��a���1�٣W������%��h0�MSM����х�e%�s�.� y�̊�mM+�c��;n��]{���̫����2K3�:�dSZ@r�*��/��+�U:�b	�q?V��[.o'�TGB'�*[E�:��6	�uA>�Y�v-�,��!���J���t����;��[�3��8��6�윿��yΚ�KӀ-�13H��q���k��?����4��%͸�2]:V��t� �傌V��ރ�8B�Q
�4��G�H:'�l��U{���핚��9��N�ѱ��w	�,dnw�Z�\�%��,v��o���<����FS�"�B�SN�j�ۧ�y�c�?.��(�c�)��=x�#}Sv�,�L�W�5S��[=K�1fWN�ya��9�ep�'n7��S�n!�>"	�t��Q�2�Q�Oa�e��P��V/!�}&����f���4��d�/��2"�|��{��9+�	ct�ǒ�0p"�c��ε�B����N"i,K��9&I���j��,�j�!@rqݥ�����{��EP�d
�A� J��j�����a�D����]֭�vˮ�	�%�	E��z��h����e�GO`�ܷ�h��C���8.'ݰ���<��ت�Y�d}����ɍ�Y'�P*E ���w�^I�4���>��*��#a��w����:�؛-��#����'s4�_�?�M�j��V��ۻ��ޟ�ey���j̙�w���pd��p҆ �1Kx&���;\hJpʅz�NKKA��\�����	:TM�i�h'�<����4�����
q�'�I{�gU����|·��֮�A�c���a#֚Ƹr�L6'��b���J.6t����<�����V ��w�x�t�՘غ1�W�^9g���&*��5M} d�I�!��.�p��8�ad�(�K�V���i�-���� O��`7��@�i���|�s�9%>�en��2rD���tpF��U�*�E�t���<7���W"��LK1'S�����tɕ�!�W����j�^��>��&�v����֚iIt�����$���g��w�_)��o�i�}�^B�y���G�t�U������Đ}��O��M`��v�o�X�l��7q�/[���`K�v�u�7�+���1��×�IOrS�K��7�쯁��|������杙�_^��eϙ�<���u9��c�& �$��)�}��_Ix�jn�Gz���.��`��X��Č�J�.$� ]+!�%�q���.K���7-ݑ<�yܿ�'�M�m�̩��6#��*ch`�cIkхN�t���;���{���%�+��|�����kk���g���[�x#G���H��`�JE�z܆)�)C��x��w�E4^c7��'䅭���c��n�8��σrN�fg�N?M���<Z��؍�����`��q����L���ϊ�f,����S�VU��:�(o���֜�&r�j��CQ��N���ݣH�f�b���-��4n�¹1\������n���.[��-Q@J�Z`VZ�0�V��&��9�s�U��ݎ.��T����(��H��g3�:�;S5&��q�}����~�P�2������9�v0�:nghy��B0��z�K�C9�Qp��R�O��4_<e���>�_K��m4\�q���F[`�E����Z���vJ-�2D�t���ܫ�l��G��*R��!�.1tF����b��Tp�w����Mj�=`����7�9@~��ËT�`J�	=�˓?��������h44\��=���M���w2�ۉ�V|�8�_�Rsߠ��H$(��>���b@a$y�=k Q��	�j\������7��ۋ%�����O�۾�X'�ⷫA،�����B���@}b�e$sP{#�-�� ��:�"��p�溆���k:`���$��>�)��4V�%;���30��VZ#;��u�<���	�%+�W���A��d�Y�Z��3 [�G(
 iJ�GG!��dF�-yԯ�B�_���l�n����-,�kV,�F�u����Ȳ ���њ�-�%�˟<�gh�V}��$��)u'%������}�GM�Llu+�o ������P�"ң��q�q�LB���A5���@4iT7 >6��LԐ�?�GG����3 >�	��j b�܋���u��%��a�_���痵΂�xj/��h^<����kD���^y���:>��L�Dl��&��at��j,6"Oj��Ô�o��Ė{g-���s�xf�tkCs��Udu�3��g>�Q��>K�)�(|چ"�����3�^���r�	1p��g�O�s@mI� N���R.�M�z�{l�����f��o�g�P�zSC�ds��/M��)M�M;�����i�`���[o[��h0�O�8p9���;����Ѩ�C)��t"vxnq��F�!����rˋ�C�m_�#R���2�`/�M_���3�������b7\��օ�k�ď���龢��A����򛪌TP�r�ڵTbG�$pP��W��"�2����ěmC�c��:�M���O�'��q�%ٱ�����d�������蹰�o�8�U+��U�w�W�@\��MiR���C�R�=�u��
y��de��* �r��h�vYr�g~"��ɾ��fS�t\���RC����p�Y�=n�dW��%�,��Ps�[�r���A�j�Hz��Nǅ��J��^i��$\9W�ؙ)˺[���en��l��զg�WY��K]?4~K��k�B�T��]܋��w��e�	�,S����&��ko�$������t
\�]�3�A�U�lZ�*��p*���>!�|��J��>C^ķ�m��]"м�C	���jR��"�Qj��n���(/n�o٘�9�qb��QW�z/;���d� �X�ܣDVz�t{͌�益(ؙoozڛ���{����ý�q^������vPwUU��U�:G�(���s*L��� G�ǆhf�����GiO�W+3z�B��|	@�aB�k�9M�r5L"�H=���&�	ՠ]���N���u�1�9��<�Liׁ&�yi -s��Y��i����&����Y����k�8�l)��� ��J&o+�.U��j�x�8X]T����&�Թ����Ԋ��D���+g��-ߩ-2�����Vwq�{W��|��d��B�s�p�z�J��.���6�j���?��ɾπ�t���O��-oп��OC%���Ր�3�~_qJ�O���,�T~�+AO��yfq�sl��]���k�R�.="PQ}�tm|;�]�)y�pU`NI<e��c�G�����=��a�]8�d�k��
�Wd��H�>���?؝�?_�T��m�m�}/fԀ蟎��J��˕�u��k�P!�h�fӸ��uz6dĕ��B� �g�&���x[+~r��Z5_1nk��d~��I�Y/P$!}�=����*z`��61��cR����m��n%| ��FK^��l�6|��5���'��H�v��o45M�� ��uS�/�?�zV���:x���"���g�y����D�Ӽ�6e�"�K�Y�W��#��4����s���z�j�D&_��z��u��+�,��V��7hM�с���'�X��d'�NR��XJf�|M�#����%?��ǧ���,�gZش���wbzz`@ސ+������ʧ3=3��ytv��o�Q��M�ؘ�m4\ʼ�j�%h��-�XU�?b],��1���bԛE�~���$�����9�c��
o*��	X�4���8����"�~5'��@�����@�A��y��`�Rl(=�p����{ �ka��b%�w�m��X)$�Fȣ�tj�:�M�y�ܑV���n#���އ���x��˽�7�I��0��RmB:�M�K�0��@���	h�ۺ"���BP|K[,~I���dك����;��6Gq��vJ�&��+r���L���%�S�8y��dul�!����8��DA��o���Ԯ@t��}��Y���L���A+�a�"2�A�4���^�J'�;�5���&��K���ޱi�c�)�����&�;߿���$�Ja_�ƥ�	��r�g�Ine�<�1�N������ٰ�A� ,n�uU�8�S-p�¨�J�s�B&>�j�C,��tpjSt�^���
��q,�1�e�J�z
��f��
�ʈ+���U";�x)�k�7�������3���1P�KT��% �b7vZ	���[�|��~�~.��n�FC�l�I�W���Vb���H�-��.}�~���пu�ŘT]x����~����vg���9vb���3�T��1�ް�c"�1r��!K���0��r~BMӏ�RS��әJ�89�q�"��k�)�w�X�vKIF��Z��n�����xs��࣐I#��e�AG瘑{�-@G؀��c��<������, z����-�-�5�!�.(tmq಻#M���ئKN��o��cD΂V)��?>US�$��b��I\l��@�Hd\����?�e�n/_G9񗧱�U:lK/��b�J�Ҭ{9�>B�L'g�vTP˵�O4W�`{���k����P՝J^rd��'�LX]�bj�2+mY��
�V�	ޛm	��ؚ�"�yr�pӌ�HD�y����v4�L�wv��1����K<Y3��t����>M>����	��~m�2VL�A?��X�[H��Ϋ���C��qL{2gz�}�r[ �3v���;D��0�"�j���.Xs�G��ُ�$9�}��B�'�u��z[�P� i�k"�9@5TU��JbP�AC�Y��uzL6�8M%N����&�	���N��[G�~s���5���͈�2��0O*0O��������>�J��:3�e\z���T�Jp>f����	🤧c_�u"y�ۼ�W�rTBq<Ծ���r�#B��k��q^�MVa�-�F�����s��(pޅ>�S��;Ӻn;׳����l+��:�}�_� t�y����,b�e�P�^N�ЯC�����l<PI��U��`cq��<��r��J���uy��~/����H{E �=���4�e��ޱ��w�WV�%h�b�\բ�����H3��	'�<D$$8�G�|�b�mwh�D�'�u R�s�T>kGD����J=��+X�3�>�m;��b=�I��Px��	���ˏ
���>m�"=��X��N[�ݡ�mh��L�X
{c��z�� ����TF�m�H�sy�s3��yvz�ʈ��T�YG#�9����6ayy��zq��<_���V�-g<X�UY��5hz;��E��ys���D��"��m.���{q�?���_�
4����r�-{	$$#<�I�wO�=�U=��Z<�L�7�"fnQ���&�(����E�5�_Ba���l�F�R�l/�]��F"� �a��
X?�;��9�G����1�Ua�@
�M�:j�q:�9	���	��-�1�W���s��Hj��[D�8���B��̥��VXsw����a��M�tq�F�u+ji��|�5m����J���?����XV忦n����z�ͧ�|�!��m4z�^��������U�7?�Y�'��ڟƧ������93����vxLA)Cyaj�(�_ILZ���6�.��͘��:i�׵2�}-"�3َ�Q���y:<����Rl�jy�f{���H�_�6�t;TQz	����M�c�,R\���p�l��^�Z�$���5�V"�n:.�|�u�A�^+�<���dp�!���y���U>SFm��+�M�¡E��S=��J�X�G'nJ�9(�t���[�ns_�Hې�U�k�y��?mg��,L�S�
)p�$���	��n���9�$z�v�[�����;l���D�=� �j����K��y�I����҂�;���:�� _K�Ⱥ׎�Q����~�����N�Ly�Zإ	c�T��)%���W�������E�Mh7[�s[���}h$�bQ(-�#_���?!�\U�}��'!zr�9�B;Q��i�q�K]��#mz�/>��sQ�z��فo���KV>Wli�S%�D�_�+��d|l�8�'�S,�8U0;M����m�\�y�׉��nǥk�8`\��5�C�J����H ��S�B�O%�:6-^��
�йf#>2��`e.𻫛ߘ�L�����|}NҸ�Ƒ�3'�HK��]V*��c����O�,�C^�������{-!�	f;�g�P�|�`�݇?��m=���tۧ���/�����sV����]r�Ǖ����J��5��O;�1S�S�f�j���?�]��k�WLI��Lg�r��J�B�z�#I��?5���?�?�١�=Ę��ot-�M��C��K�Pr����
J��c�Ry >`~tM5�01�ٯԣ}G�F��DՃ�cB#[ʸڴ�&q��삮I�7���C�� 9� �s�U`��߽�d�,IX��-�U�����)�Tb�1�����_�9�l����Uu�v��@�r�i_�.`�5r�[�F@���S,�@<u,��K�S�Ǳ�t�� }H=x�ʧ�vBlK��N#s�}	�3g"8�r�����7���-�z�����gǰ��H�.��`�b+��í������ДP��7��4E�f�0X��#�C�_�DS���a�CsJ0�/���w�8��D�0
!�f��>�N�^���8�^Om�HEz�����.�E�udp��z;'�����u���6����@�S�!x�kYc7 e�R��9�VLW�e�6o��q%���o?����CʮB1����̖p٫̯�Gz�$y�);��yV��S,9�!^�b�?y�h�"�z��-Êw�d�!�����*�۹P�}�p������D��r�*��E}2�%i�
�sUy�S�ʞ���pC9$#�k�#G�QB��Y*�t��3�uk����5Zb�G�#!7�؇q	@oϋf�����Q֏��z��$�AY��e�=���£ �	SB�@�Q^]�C���u.��d���l��$��F0�����B�}v0_ #U�y��,WGGg�v�� ��Z�a������;,��~�8��5��ş,�2]-b����o�VXS�-\p�J�s�����w6�n$&z�����O �G������hq3��3.�$����N�Fv��jB�G������
��t��P��7=^�j�
	cQg��	������8���B�H���N�h'j,��Q͆�f�.?`���Z�d��F��Zt�:.��*	���dF��0�6ca�E��І�Y�YW�q�`p4�������@Gtp�p�]Ti~V�+��Uyr4L=��%�5�߁��4�� ��ѳ�����ECQU��G���[y9#�ۥ?���q�L��V=��K�1���<{�`�ؘ�g�aK�6�� � :�gr2���q���ꗈ�iwJ!�浵#�Hy~k�j�2xGv�0�/4��[�1�2K=϶�|��=��?��=_)-�ï SbK��|�5����^+�l�@���ӕh��A������߬P�~�J���mO&��*�Zj,�����[3[j�A�⊿�u(\�� T��~H�@<z��R�0�Q]"���#���++z�whg���s�]V��|4���]m$q(_���so*�S�Ap�A��.s�HR�����s�d��W�\�����I�{�}免{\�>�Z0�|#���ˢ��kv�$Av~'X���0��yL��O����y�21�;�D���EZ�J��Y�Z%��3(���B��+���-��� I���I$.U���3�c�o�Epc�@�,�1���h�|a��\UV�ɋR�6lƯjW��NY&�d�@H�� %{�ZޠOoFj�'¬z�;�o�\y;�BHg������ݪԘ_e�f�>���3�f�+���G��֠�(O�Z�D�^9^_~�Kۨ�+��LG�Ӿ�t�6U�{k�7#x;�5}I'����2�UO*�w� �4�<D�0�4�x�����@ԅ��!��3�.�6��uhʺM(=��b�~��y���ž�#syյ�vh�i{���"~��m}R�$�T�����]~�ؔ��9{�@@�c����t����h��]��-jA�O�]��W�\��b<