��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c$�����Ԁ�R<W�����d��2k�i��T �M��&`(��d&��G����ſ��IDvW�"W$5�=#��*#��)�J]��+��%3���R���uq�����N%i��u�b����G���P��L�n�Z�([sMv5:5}��A����f��;�����-��xN��е4��{0mp�~F@~g��Q�}�,��h�����d�p��kFKN}�{���Ug^�}��:؏~�]�ǽo:�gs���-B[�c5�sP䫷(K� w�SP;p�y�>���$pՃ��g?��gp$_)D��ˊ=�Vt>�-6�
��Z8�M��P��~��}$������ivO@jt�X?
:e�ǻ�p�o���$�=�o�v]�8����v^x��oaE>��� I�T<�Vq�HΗ��D��Cx���kxהS<�f�Ĺ���8�0��0U��!�.�%Xr���]=K��:��$��@��;�5P��_go�f��jƔ���yHܳ��_�d�K���� w`�a��V;�]9ng��� ���|Q�b���,L5i�~���`������Hs�]@r\r2���Ɇ�x�H�����m\`�?���� 2��HnU
��|�Jq��J�<h��>k����t�/���m,m�! "hrv�C�$�����%�L=\M�m!3Y����G[�~��@M
�R�hA��V)+��jW�w�[-˱���LT�d���e9wa��0�G�擵�F���O���v�`�o<��0���`�|��im>�3/��R>���mOV{=bԃ>cQe��e2��:Q�U���Aǜ����yn���ߔ�AI��a�����r�2@:�ܕ(M�f�Q�1�/�
���Ag�p���TV9�J)��59��"�S-H]��(�4L<��AʡwA��!=a�q�0�����.Q�M��@b%��P4�T����;�m�2���edS]����X��jЫ�C��:��{��$̂�4�]��\�Q�d���/��	�Ŵ1e����܊\��)�Nx��ބ]e<DA��E�x�6�6r��'�0�}j�N�����.Lx��΀�f��CJ2��y�X�ǋ�I�G�3��^�ww
�1�O��0��pF���ݛ�Q��?ߢ�	�@C>N��J�b�w4fB]M��B��	'�0��Ƿ*tk�;��j��n EQa��@+d3qCfS�@�0X�p?!�??���	��+:ʃ��m0u��Z�?�(�aOr,c2���@����������gҿ��~B��l���<S�`�2�?�0@�B�F+����1�d^���u'�7��+�6ȷɭeI���J�5c��D�!K���u#���CȚ��2F��5$/w����_�ӎ��[/�F?���:�-m���d,��Ү?m;q��i��y�KQ>D�M�~��N	(�M"��;1<FH}�a-&/�I�!���9Mtm�WW]������Y%����� ��w���U:���|P�JO�ƻЁ'r�q��X�����m��]F4܃��Wy����g��<ą�8�M�l�rt�Ɋ��̮0�O)���a�:��.1!K�����(�8ҫ�}t9��OF��sҮ��(��N���-́���i0m��a�ǽ?�g�!7o��!x���a��'o'�pZZ��^��	b�.�Of��1!+�B�"rP�Qy�
���}:�V��� ��LZ$Ͻ����ˀ�������˻���S���_��d�xU\��'�����(�}N	b�".�y��I=%H��=�����g�?��S��й�Q���s�'L��WA����<����E��.������+ƞ�?p��+�\}�L��5S^���B��}1Wk�7ڌ<b2u�Q���iȀ���L�ﭻ��=��KiӼA���<�.k�Aqk�)R;���RˏT=$u�n��A�\3^�4]�D�" �#�!�z�rʎL�����<jg�Y�m4��I��z33��Iw�4�s�j@OR��.^����D�����bz�ǘ]�'���b��u�&E�\��c�XK?-N��@��X�����^�85����[/BE��������@�n]5�x�$�gz>�m�@.@x��`���fhW 7`p��TH=,2�Ԏ�%��Z=(#q
d���rT:����YZ?�g��SPͩ�L�p�+/��������������;�D��O��:��i�$�ѽ?�)�ޓh��G�=���T
rdOUK�/j1�ղׯ�U�*p~�t��A�[��I������HHG��y�v��v�/��l�Gl�1�`;��>�r��R���iQܯ��)�q��%�ش���]k
�L�T�"vYBS)����`���r�q�&>ښ�c�AB�~�4�&��D��2�CGq�Z�O��� V�r�����d!�]r8o�2�tJ���'�8����2���z�N�5c�����]���X� �HKW�$��#"��V�_оU�ʥ�貏U��av�j]��2��|���j ��Rp�r�g��A�����f\+'!�rI^ ����գ���90�$���S~��|�����Qk��~TT�e�ջ�c��f"�h~E�!�j���k�3�뱊m�GU�t��|x]�mCE	��8kD���lۥ�*�q��Te~�uݧ�}o��OU/��N����/F��C�J��^_���'(qR���4�����7�9Hۉ��~֩���K��]� (
�k��a��ۿ�!Of�X>>mlk�%�J�NdSz
�>�`���jH̶A��D<*cU������^cs*Ic?ϫ���� }ڳE����V�M���e�R��(p��4K�U'�=��o+���}	 �ʛ5�)P����"��~�O���� Qy�~���D~�	Y4�_�C!�� ��8ÚK�X�$����uYRY�^�|� y�ὶ|��GM���#D P�\:��m�Av�ܲo.|�Ҕ���ŉ��I�J�����=N]e�E��q�$��f��;�@-%Q�D����_���ً_ŒS��af\�x�+�9�P�{�����ANgP�����YL���������ub8�Y��/],�S�JW��z�b���A<�9t"L�S�P��-z�˞C��_i�����h���FS{�^	� Ԡ�ݒ��O�*��O"��ݾ`�{���8�df`x���Yh�'V)��ܳ����m(�UI��K��w"9��YM��z�񈀢�h�+�أ��l����H�~	b9Mx�ڳ��e\��{pD�=-�ig����͘�b5=X����ɳ�2���@=;d��S��+���^�$~}�dݧ�$+��}/�ߧ��n٩�ǧ����O�FJŠ-�b��A��.J����fi�a�O�鵹}�bK��$9��6���1�0&���B,���l-�5������Hg-��=uڒ���ҙ7v��e�E�����#��}���'eJ���i��!YP]��p>��{=��yy<p�����M���ޭh���/O<� [	P�"w:n�(��f�H5Y�Ii�kd�fL5���`��w �:�
���Ꮙ���q����k1h$$d�3ES�$
���h�
1��pH*�ޖ�O�)U�Z�J�(hgL3=�a]_�vJP,c#��5պHC�~�/�E� A�[�S]r2c[\������AHʊ�0��A9�Yل�	��I���Y;�A����'�$��v�TNm�r� �H�,|�3�ןY-�={ۙ>�
�KKP=�����ꊹ	 [/Hr��ͱp�����`�]{N�ď������wKD%v$�ZaEįX�Ťl�t=����`3�[{ ���	m<b	���@��8f)��k��s�&�j�(Ԥ�#������z��>`�^��Y	^w��|{6m�˫��Ұ�j����RAKZG�~������ccVI���E��ЍQu���be	)��q�b�-�EF�k( ��ߞ~;�O�����]h����5@�����?7(�[��+ur�w�0����?���E����F���z���^��w�o�P���?���{���h�����,V�H����IlsXx	|S}�>�.C*vq�x-��M��A��:��d��~d9���[�f0��ږm�ګ��LRj�q��\t?Ѹ�D�o���.ċ��Rz�)�ZsW {�n�t�^/���AB1�Ig3ݩ��Ψ�	���`����t]��YJu��|���4(a�����u��D;�z��c�D6�=��u:�ZŬ��\o�KD;���t_��2!���
���
�t-�j��E�c���|FZ�X����u
tê܊U(S��͎X����a�����Ife̙֔ֈS�S	�㔜�r�Ț,tك�Q��>+�}M��rdx��:��Oֵ�Jt� Ҁ͹��\���!��z�Y���1��9Y�lI�0�L`:���g��#w�?���f��q�LN�2��Vw� |�2r��C���N�wC�!�%^���%�Tc�����g��tU0�G3���w��<M®��7C#o�>�DQ/�FSY%�6r�5��<�YpK�� �{�"8���{1'���](�3��\&o�����y�uÆ����ȹ
��l&���l��p��NZό.GNc/�9W>:�m`�1��(�.�1�g>W.X�򃤘�Lۚ�Y�ğauILz���ɿ^���=���L;����W��p�I�w�G39��#^�	>��(q������*kl*��j�̚�v�n��ݲqc|��*�����_����|K��q]!����_-�F�b��ۼɦд�Q����� f^/j�1��2�4��R2�_�������uDc��=N�n^�D`��5�;B&��I��L�N�+��f�&ZQ�-�x�yr�1C�̑��."�c(��.� ��������Q�*�d�뿼��AM J+X0��!X��w
y雹����R��j������>�(E��MN�]T���(Rs_�LtT���<&�#[�B�,�8��