��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&??��vD����j)�g����*V�Z7���[�*H�1�6Ք9��/i�fxL`˾����rF�d�ɘ����&8��'y��Wy��zw3� F3à�:��l����z�n��dr�q���i��<g-X0��\�uy2�����k~��r~�
*�A�>iϒ���]-y������j��PmaO}����s�>��������친����hu°��������/2���7�,���W/��d��-��|�ό�`��~JR3{Hޮ������~>���sOh1�(�D/Mw��	e_�fvn9�(�
R+t����E9�#>S�#od)�>H�່���_@�Sbf����[�"�aNx��c7>T�4��N���!��}#�ݽ=�RG�����e�w��D��m���$������i��_��H��M(=�XASV��&O���fU+���G>��?�尲��䌧���ƽõe�yU�;{Bwm�@�H���?C�!d��e�>B<���^�K��4}��2�K�נʐ�W�h$�5�+:�����3�t���S�W�z�c*�K��M&�[�9��x(h�aI5J�)5,)�|L����(�YȤ�;@�rf0������0�w妩d�*�x*]Bk��Or��oϠ���C���?�]1k��}!��|I����]�K�믕P�_x���T-]�o?4�z|�^	x�>ǩ�Y�B�����)��C�
���̢
���;�v��{�کn2�p����LY�w ��o��ofic4�|J�}6����������+�V��E4���[mv<^;� �â�Z���|{��7(R����?jՅ�4�m& ��"�8�uX�a�>�<���(�_p��>*��]�D�g��!�O�ݠD�c�Xy�3"�5J��I�:���)w<Hڈ �ֶ�ZV���
 e"f����i�[�v�)p�qd$�ߗ]4fU((!�_2��*ZVƍ�=;]��y�Wn�!9ZTa��RRX=�T��m�H]�.��\#6c�$c��:���2y�������	,�������I��2VÈ9I��N�������渂@���U[]{Y�ar��Sw�Ꝥ+Ǫ��Z�M�������.��%0�+P��:��i���%t���߮^�f�2!��ua)�����6W�u�$ӌ��~�����~�<v����Q���=I���bIp�f�I������FVr%T��r[y��4�ޱ�C�0��׷�:���XJV�+�"���d�CS%����2���lgH*�� ���1�#������X�;ERӽ�0�vDz����(-fZ�=��m��c�hF*1�g���z0A�ꠞp�,��ͻ��q�i��l��7�SL���=V��7ϯ����!%��&�R����_�AM�MO�cY��+�.],yF4����G*��]����Йg���Skbg��Zcp3���q�H�0m�`^� Sq[�h]�=T����r�.�C�D�+AN�@�g1��mEpHHVR��rU��^���Y�/�����>m"M�����N�Te�6(K�ێd+w��Z����$}q�����	���:�����^r��D�J��`�o�u��εm�\�a��َa��%�.�/f�����L��A蔶GE�S�ʋuG�W
���j��dY��_�� ��8��B�.=h|�2P�Sm���;w36�b�W�6�k�e_�a-�pǁ�_!0#���<�\x��@
���ۏ/���OI�-�
�[�V=�U��@�����H����(8�a��A84�'����,�QG1�0�Gm&��_~���D�cz}�=}9����(�<B�������PD�Y�Z �֩X!��V�Ԁ����H�DDIͯe ^�Oa?v��<8-%_i�J��$h���й"�i68R�\��[�n���E?԰�,/�7�ġ����2�<z�o���B:��~UO��D����LH��T�a���*�Q��v	:kY
Ei0FF7��Г	R�?�F5�rM�0�<���e�z�� x_RO2�P;T����]{z�,V��X4���HH�Q(xeD���J*��`r�l���*���D竵S�jD�o��To_2mL;�;g��L��v��η;�Ƽ'O��FO6�B���W��M8�TI,����>�.���=b�R����=�����G.�gdv1��{�m��<��t~o4�w9��<?�ՠO8�&�FS� O���5�Q�b@�\��m�( �m�*��k��h��}�.��av����oe��tX��8�e0�×pi�����4��Ĝ|;5�f�KS.���k����7KM��z�y0�;��:��ց|�@j ��mv?b��`�b�������T�m��m^�z�[�*]*�P��n6'Z߼�>���e����mb'zh�9�ݩ��'Ⰵ��ΐ*P��a9d��'rX䧜�DH�dj߻,��Q��G�!.W��t{O���ǵ�~��g�>�IȗI1�#�f��U����5�������kR��0oR���_��^�`�V_����ͥVe��R�R���UP�<�

�(��l�P��\,����c���ys�'>������H+�㾪�pk��UL�G׬��~1�E{����A�PNK��&�4�w1Z)�;�˒�� T���5�U��c�~(�]N{˄��59���sRE�*$���Q�~��+����B��`�����P�l�d��'�A�Ӝ��m����]�7m��zs�xߪ%\�%�3|Ic�A�*���<f~
DGɲ�A���t���=�3��܄��Jv��y!7A�q0��}����(��qE�l".H��u�V�g���R��a���ac�]\:�5܃�:\�-�YH�G�B��\tf�.�7�J�It�F�ٟ�11'�`�\)>~	��#2�-<����!�}}�A>|F��X\�F ��۳��<J���H��*2Sr~bي��-�J��5��=��M�8-퟽WmO��!!��`ɨ�I{b�%)Y{YVq, ��Z�)��3eu���X�b��bC����;;�ya��V�-�{��)�O�N��!����1V�Ҕ�ٰ�2u�棽 ����R/��$WM�hn@�6!Oƣ�8m�W���Ә�n��|��G>z��꣫"7��:(��C�8<����CM������}��c�l%�4S��ٜϘ�fk�t�l�Ko��V�ߊnlΊ�}�V�]�J�6� �q�׹��NN�t=ei�9Ǉ�tl ,�Ij[gI��Հ����+�x�k�D�f����Y���]��T[[�� n,���6m#���$%�Z?e0���ۻq%D���=�	�Դ�p��^\�Uۊ��V�@��y�S�c��̒)ܨ�o�K�_)�"
�/}c�I��Ձ4:ÖE L-�v|�w&��ĵм�ի�p��B���3�Ī]�Hk1i=�"Z���g�g��
�i�BЀ{tz��2Ջin�L؋��\��Y]��Y���W�^���lGP�z�Z(��=yަg��k������~-�	�edJ֫)n��W�@~�6DkX�LΈ){b���N��sg�_��R�%ԑwm�Ng������wU��v�O��޽��1z�((AX�ΗwC�_J��I.��|��J ���~S.R��Ē9�U�[��՟<WP�,����nI.�Dӈ�V��:;M{#A7ܭ�3Yp�wU��=�*��H�]������ZP]�#�+oT�;����5+2�L>��DFid��e��<��[�xY�6(�&���G"+J]O9tϩ��˦g�� ��1g�1v�6�Whr�xI�I[��%�*��d�]�.��g���,/6�A�v�az�>%���U�Ls;=ez\ﲎ�yJ��LȌ)���.��0G�U?�ѿ���g��T5Q~Dݧ(3?�
)"<�a�D����f4���h�[lc�W*ī6���J?'N%[^�៹:�L���6�TuQ8|O���AEx=z�5b�["��Б��7�S�T�E@w�k�w�S>Fml��1JL��������u��S&RY_�k
�]�>ޕ��	��5i��u�����ɜ�[��i��m��/V"�N��d����'8������I��|���Z�'_�Ɲn��*^o&^���l��[7�N���%��vq\<�?����}�n��1�@����q8�ba�2�jK��㴶�`x0�xi�4��Te���IAFΩ*��*.' �R�a��+��5~RsbSƆ�L�����t�Kѿ�g{�mue�O��-mn�lwK���Ư�X����>��|��ki9Ĵ�}uL�$2�� M�d��XM"Q�j��D���ʘ�E��0ͧC�	w��D��ӗ5S:��(�GS�2�����?V�)�73��Ù-�)����t*}�>�����u	�'..`C�(l��8~��Xz��m�Or7<ғ�&�P�oݛ���m���7 �+�Ȥ]j}����,��J͖h&l�s�PBJ#J����Zz���3�[Zz<��N��4�|ӱ����(+�|x���ׯU_���/dJ�l�'��5��zq���
X+���$-`	/j�}�<ʁ+����9M@o1��[�S������%�s����g_�n����R����Һ��,���]�!:/.��b
F]��]���z�]"����.��s��nj���c9��|�s�4Qs�P�؏j��-��;C\�1RBL���8UB��g]M+�h�@����R���n/�a�a
�j-y������ZpZH9,�_^U�ǚ~�T�O���j~(�ʬV�u�pMN$f���४*F>x��J�3�L��I������2f�C�k�>�?'�@�H�G����S!�&c;��m�2n�Ys�7���������=�#~浃��x� ��E���-�ZحL7 O-u��ST}�y�(�'��TS�����s���Ϟ4.-����9��4ęj,����%��}�kR�lTZ��r4L�=2uҟLofճ�����i�����r�|ZϏw���2\�����PF4:���miр����f< >`F��+do�w�-�l(���N�̓�ГW�c���1m�<���pi��Gy�|��:a$W�-�^ �5�xO��D�T�]����%�3L�V�Ae�K��c&,��XǼ-䟺���~�Zѧ�j�<<�����ըn��*��c&H��kڛ��%����Vɏ�]6����`a��֫��N�Ў�ct��q�	i�9��k��������Dp��5��#�1M)b�[���"Bݎa�,oo�[8������Ɛ(��ä��gCK��Al{rP�TB� a��[d���S�}��y"cDm]蟺����%o+�9�.�J�8�P"�����}G�9�_�����D9:
e�1n�-2�vf�o��lH�_mz�t�����bUa%�B��u�Z�����wn����Ai���У�j�?��U2��U�ܒ��A�˒/��HS�x�@��-�'W����rrf� ���-L�-RI�/�6�nN`�5�ۀ�dh5Z��$���o	��Q��u�$�T��j)��r^�@�m5C�uݺM:E�Bhf�0[/1����P�Łd�Ϭ7d��])_�&?⻜��E�ߖ�ګD��Ad	�ܠ��
HQ8���}T�yk-�eIlXm�+�뫩�����kM3T��3��e��J�H8��j5�;�61�+�M+��9,�.6f,��^5�1���Ij ���W�6�*�=��ע	��>�
k��E�jg� ��B����$"��Wu�A��B}s��3�/�wC��Nz��Gh�����I�oH��} �C���� #w�GB�����9<ޅn�w ��o�d	(B��Į��������-+��U�/�-^Y��
o�j�Ld�X�B�V<�r"�q><j������*Iv�,�m�mO*�7�AE����4��}ǨC%��x���L`4�)�ޛ���l�<���)����n�L`>܋^b$���3�6�vv���;��G�r�2��~�]"_��{��MC_۾���֓I�8��]�6O�v^���J�	���W�{$��)�V}n�������X�����m�+ic�7&�cAq�$TZ�=��9K���G����*Uk��V�ͪ+�J쓬�e���⢓ô]g��)�TmԧA�I�y�l�FG��pz�Ĺ�{:��Ѷ�X�	�_��_D*ioa�O'��^h�2�qVz����A�^���(B�خ>kZ�R:� 㬺o��Q�a���O���r� E߲y;]�BED=��^ky�
bO�`���*iam;颿�m���h ������u��C&`g���\��7�-��Т9��0���|��.!dN����<��]FB��n�3 ����Q/�h�랧�i�7~ߡxZ!��T۰���_2�TN��E���n��i:�r�g�� +��ʁ	�ţMԐ��+�{�U���������%��]`�car6����CxG"��� \2zټAi;���~Kz�ga��-N�s��S�#����mߏr�z|]Ӿ"�Ġ�d}<EPj	y/BH���Um7�Vκ�T��`��j�'��s��ߓֿ���J�ǃ�0Hx=��.l9���<��x�	-~Z��q�N]s	�|k�9xb����Ѩ*��v�+^-��(漌>b�gP�����t˂�n�"��f����Ȯ^U��r7�/��ys�M�y%)�%��ߪ�0����uEɊc�0u!q䓄X���$ň4 ��+�YT�8t�w�P���mF�޿��b
̗��"�@�����Ί�! �H隿O��Fw��I]=!��s��*�ط"�/,(cJp�0����!������5����i�[�W�v+!I:�+��AǨ��BҠ�S��ώ�5�3"�~�)a̠F��u�fAP
�0�y.:��5�I"h�>�}�0ej ��]ߺ��<Ϊ):����I��{�E0WLºq:�=���;��T�w����P�̬x{�N��o�Au�<�f>�Ɋ��W^���] Cns��W!oI�����=Z�}D}�O�!� Ɋ�3A0�~El�74#��kpF��������#�j���F��'���Y�X_��S�.}�w�w���<j�&t=K� ��H�H��
Gn��a@ߝ�'(p��j��	�[Ec�%����G)�!�R��y$��-ͻ1�tͫ�3f㦏W�/c<�L����m^>��.��?Cǰ�l�|p
F��Uҋ��?��qm���Bs�5��$�ϯ-+3�b.�����
*z.���%�*�|�-��4�J�L��-�S>�Z1l��G?�L�ԍ�t:aȄNk�����bC�n�.Fù7�2�p�]z�����1%�k�� �����pph�]z�=�Ȕ��O >�`��%N<=�x��d]dr�і:y+��Br�Y�9�P�RJH��3�u5?�Ne[�5�!���Ͽ�-�N'JA����P��j}Y/� C}�B���O9��ǄZ�lj�z?+�*⠀��>A ~ޚ�	��.�p�]�ԕR���8����SE�k]�
�kg�qWT氢u�`so~����c%���ꕎ�kF��-��~\_�*옊�O���dJ�y�P_�8a�����-/aLq!�P��!XE3&k#W���M�kJBB)XJf}����m.�� �MX��e�c���)C׺�P�2q�1E ����T�2bf��*~��O�'���2粇&�2q���;�-B?�vs`��v8R4�@�ƻ�8(�0o�R���񏧾�2nqj0?46�C���V@�[�E����-�ȹ��0n[/�}?p��c�<%�V�]e�7����#]�I��S�%�M�����HYbH:C�-Nc,�!��&@��[�Ek���= �u��V�<U^�齩�
'"!c����|.����]��́2�:���}T��Y_6b[�U6q�������W����v78�s��:h�A(���m�!��ɚ��)!|��= ʅ���؉��8$o�����w��5:�n��%�E֌����GA$e+mxS� V%���6��{�vB�v��X��Q�ҡ<�[�����)Dm��a�$ƪ��^sr{;4�Ѝ���!��ش�VX��;��/�%Ϲd�x��ȥ��:J]m˝*!V�0?KG�]��P&\�QJIJ����VW�k3�E]�
���˂����?��3��*�E�[�cyc!�r��gg:�!oi�T��E���,#pt����N�oo��R���J����A�A�	L~w�y?�ǜ�R�'�
���X�z���� y��G]P�w�ע���'���1�S�	1ƴN�:�=F��?5�k�l$J�X��s�xbB-�����$��11��Uv���)h��#(n��5@ﰢ-����Q,y��L�5�85������.�Ԣ�Ɛ@f���`��jF�%����g5���n} uI7�i �_FT:q�8���,���-��7����_�	z�G� 2�B�=�Q���Eo+�%=l��iZ&��0	���}j��l�#D��-��|�r�����ƎVU�\��q��&9�p��Cz�O3��3��c��oZ�p�w�	�Z���^I��Mv�څx;TV8?����� U������tC@���յ�=��rq�J��a�s����w�@��[ח1���F��1�������1�ݓ؏��	��"�:%�v7���4,�sP�
��KߘR��􍝸1O�����R�����$Y�d/�5�Y���w��>C�4�̢T ��혰ߐi��T��&_q;���cd�O?w&A�ұ;@ ��Ek��ڨ�a��*�{X��r����(T��a1�xג� �f�kcn]�|�ʈ8='Z��@�����MYXn�x��#�dk	��ͳ@u�~k5Q�E����Ǟ�ʪ;���qg2�z����E�����x'��#�p�'�\ڳ�� /^�k8�mf59D�s9r�pP�0B'Ǻ�_i��W�^��)ɴ��\X��V  $�D�/삡I�#����X{f�����q���)и��,����i�5��%L[�xDv�s.�(	�v23��6��p�鉄��"�|��  �q������O�k���2Q@��I��r.<��c�f��ٔ��W�L�7��{�����F�����!Ry<wJ�TB	�k��g~d��2����9{̿��u������~S���/��xV�M�^g�5ю�+ka��,��AQ�%�Sď,�Dd� :�-�M�KZ� ���-<:���)��J�l���'��֒���B�߸q�A��Q�rJ0��xt�f4옕�����"R^�
m�W�7�0�53O{��}�hL��s�`���!$���p�g\��+n{Ճ��a����9{[�T>qN��\�ωύ�s!,J���J3�i�P!A��t�ц �B���M�~��6���-v=G�9QB~���L�����-k�i&v�-�����'�x�3�`�{lژ�۾JA*�=��3�H信�o��qg�~�#��I}6��=�x9�[�q���}
T�D>aG*V�:p��ho��9sl9��
�9��/���q�2��Tj&ܸ�j_�⯖b���a.�����q����Zf��:��u�r1d�m��Ħc�J%nj�hl�^���Y��X픬�i\MDoU����nW+�:x�T���i�3�?����C�L(,u���F��l}Q�c:Q������YV>#!����7JC�Pa`J�~�8��^ƫ�-k,����s���yz��j���L>��dִ}�����Nd�4�Sło��Y	���d�11�d��E�^Lx���.����XC����ݞ�yw1.�(�4��׿}=��WX�M`����0��Jr]׆ܵᢾb�f�@�S{o�-S�WG�D�����.�����I"��ڍ�o��OM���u&v��S;�1G$W�16����f	B��5PݤHҡ��A��ߌ�&���Oz%��H�dџ������zW�/�U�6�o3h`�������[�d���eفI����'FB�R� �fL��C[�C@O���Uį��(P��`L���]���Y�^���n��R��'���U�7zL���YA�J��/Z����Z@�C��n�f���}X��Ⱥ�s8h��S���D�P@G�:&Ȣ�i�{�-��5O��pf�nw�4wC�p�2��v����f~�ZL=��L@�*�C��w],�ݽ<�j��n���j�2���e��n�0ϔ��\Ǚ4&wb��is�>�S��+T��w�Z�	���l�z]ri�[�`>	�ml���z"��׈hGm����͉��o��+�L��f4H��C����<PX������A'-�.,�4�W��?����4"�
_N��D���a�w�ܟ٢w��7�ҦU/�����$�7�dPLqu�
�ā�|�&��� R~�Q�,(2�>�;���UĒ�2b�H�kXlt��+����pz؀ېȹ�+�c���;x�`Jŵ7�,��9S`�#�`�f�#ڌZxA����~Q��vT ��T��u�ޒ�"�g��ǾFV���\a��@4�+��Yq�b��x�d ��N�]�\�A����0wLӮ��kl+g�*�����	t}�T���_"?�7܂eE�>���	��]  l֡̀����nN�@���>R�	7Lu����1�WO"v���f<N%@Tc��#G���Ɗ�V��r�J5�9fTT���nH��e�����kC��U��e9^: ���g�3�W��u#
�����l>�#��l.\������[�Ώ)����ދ�_쑒F��f&��KJ��w�JE�P�ꙥ�a5��ᥓ�`y�%Z���M����ȥ*�h<[�f��\�C�hRe�i�z�����O�C���W�.��hG��iRqg��vװ�4�����O�V�sv��Oh�u�s��,.*���)-�HN8v8L�{�`�+2�y�d�f�eW�A���+��[ay��gW=͔��	R5�e:��v9��
��5[YB�sA��1O''���q�k������K��5)R0 2L�ɧς��ҽ�R��8�lf ����6���H��2�ֹ0/�d���J�Y�()���I���E�e����c{���դ'�hD(	 �')�	�%Y:��4����N�D�y.��F�������ě����%�.H��%C�AgI�I�2m���r�k�JoT6�@�/�fc��F��f�����C�!�Z�{@�K^5s�~��	[�3�@R�l��I�>T�Ѭ4�#@k>�3�@��V�;Ю�Q�wdb���ټ+�ʼ�l�v�2�hH�[<1��=���Bib:h�� �nٲ�V�.m��o�Y�+�Kb�T���j y�M�[��}��~�G^������S��ȸL¸jv����f΂i����O��4��E+���A��a�N�.I5\�B.�^�/�ƛ���{z�I�>ֲ��3�!��ؘ��5\�Ԋ�?��ߺ�*���k�&� cœ/[~��x�Ӯ;T���7|���)�	#���l����ք ˎ��n���2�F0Ӳi_�/���ن�:�K�#�2���V�͊�|�|7��UtO��@)|��{S��X_���(O�o�Đ���`r�����Aun>���W|��<z2�o5�P�*`�KM�T���6/W�I�۫z��D�n��qX�5��|-�y�A���G��������Q�7:v�E�n�K�w��e�O�ys��7����-ϊ�+M����!����汈���H�'���B���l4cl� �� �̑0��|�hy��?UC�<��g7{{�	_	ց=Î*1�a�֍q~�RpB?��>~-�?�LeTC߱G�u�<Lq�$|lhn���D���	�b-���(���$-�{Y��y���u8����v$����V�9�]�x�-ԇ���J�� s~1S�vbz�����`6��:b�H��[ӗzm#��:�v+[��8#SBVq�?�tǆ���3�{���3B�8�W�Syڙ��k�����62�0����O/�����T�K���܀���������""�e8�шh����-�c@J>m�U�_y�6&�M-m�ȩ�2
��4"	��.���:]���d\ �}��iaB֥��q,X�E����֦=Rs_Q ���S��nЯ�Iw��4�z�Ǽ�\�K*^<���s����I<P�t�nd3u��x��3�`�����Gڹfӱ!`�]W�J�=դH�]��cli�����v���Ĥ+�՛�Y�G�d��IO�=�-b��?�1S�������
����n�}��dd�o�:�1��8���/0�;��"Eg�n�g �#�͢3 �4n��Vw��b2&#*�������b����������(�RS@�"c�d?Z��p#
�y-���¬�BזּXGĮ[e7;��Mi|���e��\����Y%�!��Q�����e��C�V�_|>��yA�CM�W�w�z�թv���$���y�j�^�6#���
+ 8�<�����
M�t~f�!Є~_�v��ֈ�/=}��	P5�Uw����2>�r�e��qR��;*��э�����[�q��̻�]&>�?u5��8/L��Fl��ƎyU������y:KEf�\{�h�>6	,NwO�Mt<��S&� ��'�D
��=^�9��^iD� �b�$>����:�s��vJ���e.�p�z���KN5�<�}�\	��R�a���|j֍ȹ�_M��uv��9�3��/� ����6�!,{=tqƘ貿��F+c�T���BS~���]���@�:�n�6�9�]h��B߲Nϵ�>V��,H��C�c�aڕ)~ѓ\w*�(�����ٹ�b�
���h��(I�;'�",y�q�ճkR����ӊ�)6+�Z���°�=�c]4��P��F�u�y̢��/�[�}��n�]���Mr��l�|����{�(�˟� ��*J�:��;��L���c���`��L����U[{L-]`��j��O�3����E��r�Xv�G���L9��G���e�[�c�A�K�N!��~�⒇0O�kA*��}G�ܶ�J�f`w��e;4��.oJ7yL�>L`)����C���ܸ_��{t��P"�e�.���3�?��� �����yb�R#P�ʡ�Gaf�J���0΃\1����r����Q:;p�r�~�.�d�S��h�ņ�'�@(�.[����� ���$��G4��5!,K��0b1�B9>�ȂC� \�,������>��Ү���Ca�%{k���"�8��R&R
èP\��}�y�3�B	o*����u՗n�Ys�n�d:}���T���c�H�L�X�a3O��u6{�(1y
�d%�p?���b�lfQ�9۩^vu�5·k �{�5i�7hqx���YE؝��dk��[��n���=Z�ۺH�(�]�`Y�oa���BD�2MZ?e����/�����6_�Ύőd6K�3�K�������	s��k�#{�vZ������)��t���q�#��<=)
~�������d[�/=�K��bƢ.�Ϻ'xb^��->ҐX0%F�i.\ܱ�W��,�= g�x�=�sX��D��YJ��Zr�Cs�T�/Tˑ�e>M��ӹ)a�l��Y�ARж3qTALcU��a�ƮE}%{����� ��݁@������a泄��.t����>;�Tڔ8�S+/�T�G�?o�&�-.����������9�"(<��^l�n7LD>����8�"�y|���L�ş] &g��j�*y��a��6�F�p,$�1�bd�)>����|.3�?
��S�9{kh_�#gL4��r�jT�L�$��)w���'������ȗ�j�&�Ԏ�WY��z��$l�,R�Sf:&&|
�;ԗ��)�O���JF��԰^�)�J�=%��3�h��l(DQS�S�#�_���ֶK��B�_k�S?�Xg�у]����q�~7N�h��q��?�	W�1���-��ǳx�\k�C���ƺ%��N�AIG%i����i�K��� �@m��b)�W	l��5 ��ĢO�D����T��R����h�ҋ䎶�����M��[VNK��G�:P�Qw5�TQ��b�&}� �c|�R��M�c��v��Ël�j[����4k�����(5�Č�"JKK �9I�5� f����-�-�T�4
�CZU�;.3@3��A꘢!������@��x��=�7M��`���!��m^
�a�.v��Z�f���lk��E1B(@H��z�N��jO�/��˶#~dI �� �F�f�M�¤>gd��������{�P�����dG���<}�x 0���dM�u�$��x�]Pd+�7 �>z��M 2N;ak1y�5�pB��6�'�!�tO�����C�R���39MIKW^|�	�O��G�
�x�w�휳��E�[S��*ib�l�A5$�D�3����J=^��,4�Ʃn�B�\�Є�|��bs���B�.`�J2�S��T2�mq�D$�'�ȢV��I4�[��+�h�4_d���|�V$�]|~�����E��*XRb�Q�i����+��_l���X��M�B荤$L�K�����=�����a!��95/ȉ���W��q0�(F0	�U���K�ݚâ+�]S�:0�Ǵ;IO��!������=���A�I��	��KҌ�͆'/�:�����U`����b��?�l�ͻE���5���� ݈MDp~���N�� $6��iZU���I#f�s�=dw� m����=��f��9��XpY2�fG5��»$�@Bm��vz �xTt�%͢K&*�nM/A�ܨz�É�v��a	�� ���K�r��qq��jJB��xJ�1���e��&�Z�6�HB�=:�;ic�ǍJQ�¹��
7m���??Ăwb=��b��XA���p�Hj�|k`F%��3
͛\��׆q+���4'7�:�q�E�F�E�l�^�owI�@����� !`�����Ś��Mx�%��h�gI�;�4|�s���m�����13x��5�W��U�h�p����F�C��S��7p�;y�C �բ�(��J���7�w�4|��k�� )J���N��
>t��]��U��o�d��e�<�[���k1o��p�㡡Ʃ{ոXu|,^��~���m�ȸ�p�b��sp�`|���o�E�BG�S�Fu=z{���������M���#/S�uW� �����M����o��(g�n�v��A'9��b�+�Sv��JJ6�c�� {P�����@y� �ڼw��YD�aNne���h��a���0X54y��f��{# ��
P��Ϯm:��Pz�̐<x� x�o�Pm��s�N����Jm�CA��TObg��o
�uj��K���!h\����#���'��\b8���4�N�`u^������QQĮY6��V��TA�'�(��E=�Y $x��	�{�O1!$�����9x�y�ר����a�1JI�v��c�Cn��w"F8�	�{�1P��J�c�I�݆NܳW.���ɑ����gD�l�E]��(u/��s�H�r�m6{z�I����i	"�Zl�@?Ğ�a�mq�54�0�����]a�'I$��P�3�TNp|�J�#�o���T�N����\'g��Fk�˖ �@ j�D���3Y��Ѱ��
��ir��|���`�����k΢��e29���E�+Ȅ�wN��04��>~�(62p��Q`4'K�"rM����lM�_@ �Az��+X����B���Ɇ˩�ܦq��@�s��E�11����X�{{��D���d�����`f)0�{95ض��W��F�=���� (8p��[�VӁ�ІRh6���f�Q���`f���5�|ķ�Q�KQQ��P Ƣ	��Cϴ�eg	Y:�]�;S��kn�DGQC��S�5(l��bv�X���7�q=7���L�����J����ʌ������E�y�yF��Z�:�?-�)\7��t��c0��jv���a��oœGm=�cP�:����Q'�r�����@�,'�����s�	˼@U�s� }�#�֐?����ż�4Q�&���+W���٨���;����p�C���g�m�RRo* *d��/G��c�HE�pS7�e`�j� �2�F��x�B+�v�㺍��x����3��l�1���Æp�瑅pz���4�75Y��9_��������O��g�*��$��`5����@�B�3�*
�
��ǔ�`
�'c*r#��9�Z����&u������4�N��{7Hn��a&%�~�J^r��o�=+�F�:�bcb�d�[J����g�[v�|���+�t梿��Ƿ���X(���8N�����YjeR�|�m��y��f��o���<v����n�2}��llK��领����{6��G2ه��	�d�hب�f�<.%u����\:k�&�I�^�m� ������9A}z�8Y�q!�+z�1��d��ik9(_� > S���/sx�ϼ�y�9�teW�N]׊���KW�u��MO�D�S�=���q|&�c�?�.~
>��2�⌅
�N&����Ҕ��ϝ���$�aU�5�I�3S��ڭ�?\'N8��G���*���PV�P���gbT>3h��'{�V�y����3��DCcy�0�9:�����>�Ԅ�)C�H�%�w�	���Kl�����)�txB �B����@4mF�,1`���Pޠ�{�hM�ʝ�K����JO#iC;T�	
��Ȃ��OR"ǲA�d��5�K�M* ��q�.�\��^��,�_��l|3:�gV��2=OA�_n;?�q���w�-��I��UKd~'��}��
p?F�4����W�>(�ǹ�D�e��I��\��K�hE�����
}2��H4ʬ�@߶�K��c���'*;��u�������P����'$Hḧ�Iȡ��\��.D�H@��.��"�����p��[0
N�X@� 9)��[�KV|���e���6�RR�:�oq,�bH�;¼r��b@�����F�;�3�km�*,���WcUc���I�6f���Â3&X���P�t�	���r�7w6�Ƕu�uI�j��N��� ���"mM��HA�~�i��?�rw���S�Euۘqæ}g�)�+�L쎹U��w\��ݻ��k��-V��v�/IGa�d��9��G��Y\����ލ��i&H�7x4L7P�-xn��֨�3b�4'�����Ufk�Ƴ�-�D�ћL�O,��4㨄�J��#�&�ֻd�{G7�،U��d]�C�9`��j���*|�'�uL���p4�K�=^(W?~d���9P�UCu,�VM��c:�"��0�)��c"�"&<���n\L�4S�������8`����L��4�$!{��Y+�]%9��_���U[�J@�i-��񠦹�:�ƹ�h�w��Hm�ƾ,��(=��"�}�&�i|'W�W|ܡ�`S�e\��������NX�
�����x^9d%PK��s��틂��I�ė�rD˧�A�p�Za��6%U� 	���'��#8�<h�[�����PĘ��`U����=�k>���&Cr�IMLOHR�����
b!B���#)S�og��M��:'��tN'�i�5�Gק�@�<�����������V��!A�Sb��C�:$]���������>]��b���*9;MZ�j)���VL�3�q7ڏ���v?ʋ���A*���(Cm@�y�:�����ȡd��l��$ G��7��	Xѕ rf�)T�[I�G�X�_-�ɂ,��{�[H��ч��]XК%��n��� 9��:f�*��.ڷ��"݄��^M/�{�I|�8�"z���`�Z��.��g�Ɋ#١�"���pH-�m/�>ݪ��&��?W<g�Y����gv��Qg���⋣�Q'`񧯹W����bĵ[�V��[Ld�3���|�ɽ�%*�� >'w�#���i�G2l�R[�p��v�{���P
����k����=�jۘ�x���-bbE��<Z �0'�1�푕N�Ȭ�΍�ƀ�(wRj�9�GI-��f���0d��8��_+�C����s�� �耗��ī���X�	r�޾�i/d�u��Y�[�Q$��{��
��2�;0��og��2F��1�j�U7K�O?��n�ty^��R2d�����T��4���0�%�>� ��S]e�G;$�P
��RD��~�:w7H+�]���#+���P=-V�R49�gzG"|Fڊy�N�Q��C�>V�9~����=a� 3�e4�j� �ȧ�0Zf�����',��ǬŦ��h�7��m��G�[�{��cҲK�#ku��������M�笛�I���G��,1��#%�����3v-�qg�n�i�8�m���%�it8G�rWj�ћWg��T+�KXoa_V�L����Mby�Ƙ���A׿j�3�ly�y=M����=�@wH�"��]����nvl{�h��/3ye;�h��X�P�L��~��=C�`�ށV���
�&��_p�&INs{�y����ׯ�8|�[މ3B�-Yo���h���Mar����H�R�ނ�4nf�_�)������)�o�
��K�J >�]f=_�??��)+x-u��*r;��L{�HS�S� ��M���ԓ��Ӻ��_I�	�� R}U^QS�8�j�R��3�U �k�!Q��%��W�q�D��rni![�������iU��	Lt��8�듮Ԁ�Ω�F���u���5D	��<-���x(ajfxU��F�L���(��������Yc��gNF739h�T
�B;[xU����}�Q!�n�Ed��:�Y �B��ݶԚ�j99��7��*#M�M��#�/~���sA�k35�>��D�օqi7)�yMeQX��&'��;jn�7�#�����-d�3�X@&]��T>Ix�\_�n�骷���N/|�S���R�W��fՑѕ�ි��Up՝�
;)�ґ���ʠ������Ǔ#Nֹ}��ɝ�B,�?���u�����LisK�B�'J�^��.<΃�/X�AJ� ���ݾ���B�e����_��趘�"8�C\��-�8���/2���U&m������]�Mv|�?�=?��ꥣ (�C�I��ȳ�{T�m�\Kw�&#?��� �s�o��\r�'5��Q���ߞh���0F���f�����rg��|�srj(�z���|���6���1*�.����(v;ْM��\�rv�й�}�����(�i�̧	�;`�2/ӹ�㭣NC����R�6�#R�TB��V�:X�Z�7�.�"�Yl���:�W7�0b;��{��kA>��5\����G/4�i*N��n)s��=d!����0��a��̬\�.3��Rg�P�CG�M<��D�渫V�Fp>�#��<s�W|�j����'�	�U�}�9|��HUO+Ȏ�]����ɴ��YG�6�4o��k���/,���#s$)�� �ʀ[��=t;�z�ƹ��������3JL�>�5�%e�)�F���(S��vX�J���k����Nv2ma���\>Ŵ��"�$(��t<�Y���Wݙ�
�l�k@�^��J�^ܓɿ���\IH1�&h�Z �zVP�6��Y*, ��c<5'��r���Hݥ�A�6Ue�� �2}��Pe��s��ê�+�'��ٌ\%�.�Vε�lѣFkڑ2��>ʞ��"��2����t�oL�D>�&v`Hu�(I��O�?Q9�-�H#�i�)�����::�9������h��m�9�Sb�B��$1�� �ZwpM�R&��P��z�ӆ����4�@9&@��bՅT,<����^h?h@�,	�V�-j+RI|_��y�K@�6�y�;<���Nڪ�K]Dl��Z�G+X$��a2E�D���i��T��Z�<�Y������Z�Y!�X�S]����8c2Xt��M���y�>�B��PA���M
�:˓�Me�O�	v�;�<�d�wr�vu�n��^nQ��ү�lw��JS=�D �/�������D�K5H��x&����a|Y� {tkX/�V�|���+����",�l6�`���^�`�kl�c�n5�S�o�"��P�[�����_�#��*�=9�U"�Kѐ��u�T���)W� 5�#4�W\���|��+7�	(��k�^��J��Q�~�f%�����gQ޵ރ?Q��&�;���_Z ��#��(�O�ݓ��1�W�$zǭ�WAzݻx�[E�� Y�t^eks,���k{��t��O@�E)��E�;��au�<��K���'�G��S�	l�=�/hH�ELsD]_�ﲡ+dG$��);B��$�(�����o5P��� �U���3��StD����)�ȫa�d���!G����0 Gx�2lZ�Y��r,b�U�������"�Q�~��i�Fzw6 (��-6Um��ϗ�#/��^���9�����<G�V5#�c�ez���K�{	D+�HQ֗QX�c?���J|,��z�Sexд���eb�l�A.cᎃ�j���M3.!Z�t֝=K�%����Q�s�8��z ��xQ�yH��㒲K�����uWg������R1�y��`X�^F���n��.���cZ���q�-+%;�i�NO�yl.<�@-\g�>��g�n��f����5����"��+h� ��v�:�� ��l�Jqk:��M��x��^Cm4�'���T��>ʵ����_����+c۪���I��(�x��#!�m,O�:��fH�4Yle��C����e��'�d%Z�����A��#rx����$/'� T����E&������l���-&�:μB�=�Ӑ�@�S6���^��V>��/�J����mQc%�����6�4��D�f�ki�I��Q�6,�?#�� :���Z�P������'��(Kv=��q��$�:^T�s���.t�}��z��1I�|��V���H�ee�T)��O��`@�K� ���َ��0!nX ��G��Fij�O<O�m5��@~�a&�Wܗ�/�ݎ}�^�;�A�y��V���l>����"8$���"� o L�.�'n�(��_�-f2��H���?UsH��#q/0~��3Sz&�Cሷ�倳"9r`�M�!�"��˶ȩh6�Ju��'������l�!�߭[	v�7�lC��w�%V��`����,�e�t{lY��a&f}ey!��k�T2�ok$# ���c���c?�r[-��.x�v5^o`-u@���X8�68���Z�93�"W�6��:e������Q�|�r�P�q�K�ԍ�J6;iߙ��TR��p��?��W���:�H[�Q��Q(ڧ��y*�uަ �d���~p~tX'p�$N�ûQ�%��H)��m���ʒ�Zڕ�f��
eq��Ơ&��z�7�#�C��u����Q�J���dܙ�A����:|��4|+�d'|�#��\�e@Eڻu'4]����Wd~���V�&P��';�A�����V�� ���Ո��m���3��1b-
��aWO�(���{9KQ��g����N������42���]�]`���-pd@��Q�9_�e$_?�MhD^�ԭ���C�RPsr�Bc���Oil��r.���ЈADu�;^J��o���Gc�Y̰\�����~��ew9��ܦ,P��6u�$W�D�D b9��)�2������ȳݿ���js%��ӼB�q��� I	t���<	�؛�kF�;�րT,��Ʃ�U;s�10-�)�������ՠ��Uo1����z.��rw4�j�F�uGUV����w5^��4�x6t�b<������|7����cf	~��ΏG��k:&���Z�Ƣ�8�?��&����n�9�{�@v`O"!�3���cRq���u�p]��\@x�X$G�.���)����W�5��J&乔6}i�;z.����(�

Բ�J΅E���zB~�?��I�ɕ$���n����uF(�����Bŀ�>�6��I1����-�ѿ>�.c�=�elʸ��d�0� ��=�i�E0;M��YɨzY\E��Xi9&�M[�xo�UBl,��b����"�^g�2M�EV�.ʋ4�%��=����ѱ�h�C��� �pB�!`g;X}n��m�++��:v[ɼ�O
�O)�F������ʲ�]��J"�[�cK��gK�o)FAVN�ߧn�-8�0��1�B��Ϙ�F=�;5z���Q�JE1�
�!��X��$)� V���n�CXi:�p�.��5F�j�Aڌ���p�����U��E�b��{��-��J ��GI�� �rM��Ԇ
N���o�y/�=B�;��0)0�P�	��z~ ^S���J������]$F��������[m����@&�I�7�4=�F���1��tI���tC�"?�2���sw��񩱺j�Ƴ7��T�N���y��%�g���@�a.�6t2�o �i�8J��f�|[���d�����E��jy�9�Ì�Ҥm1���q����X��&����{`b��[_o�Ϝ�����t���Ҹ>�1#Sd!�o�ۚ�I�����Ej����	�a�0{YS:q�4&�ܢ&_K���j�h�x+N����������]YT���8���-��:�&3�(���g�\�V�y��ɐ��U��"�|���9�6"(�4�i����(OP����΀~����3w �m�N��\�߃�0�h2/:	�H�����SU�E���$`վ�^��ь�2�7&f��,���8: ����p���\١ ���?�䅈ޖ���B��цmiҞ�gP7޿���e옃�9Љ8�9�g,	���/��`cI�؅li��"��?8�e?���&�dA�%�?d����ݧP^�r�a�
��.E$�9���ҷJ����^;|ۃ�/Bi>��C��aP��t@��➳�%$������([Hd5��c:���)*X�����xT3҆�hy�繤�(7�ԉW+���c�(�:�T��ˊ�����m�F,�؃�;V��l�;&���7����i��A�@�u�2���~�T����қ�	4�F\E��k�����_���cJ�:�����ߌU��Q3XYd�z��WT�y����]��� ����n �E��b�o3�y9�t%S���1�?A�Zp Wi`@'�^�r#�	�����O&�~(L�w)��>��m5�%V��
��ŁF�[K�R�Pz���]8���-�PY�kxN)���<����{ҩꙃE!qh$�����.L J�K뵋r6J�Y*�+#
�x_і=�9�Γ���2CԮYJε#Ǯ���a@4��ȷ�`d7um�<,��<�j�C�01Q�nB����SY�b�&@������d�Q�>��M���q@C�%Y��m�q�m�*uC�%��9xy�oo��L͙
�O��4_��"����dE"�%��x3�UjyV�]z�x����Z����Sݩ2���$�{d���u�8����F/d򒷦�3q�?;i�ek�\R�\�����$#��{�b@��l�{ᡓ�e��r f��	����w;no(fr��^��-n�X��(�>��}{d�8X1�)�2�B���l�siK6��ffCr|�'�\7ș󜗖��=u�%��7}Yl��P�.3sQ瓛L�6^��C�xn�3|�cn#K���_�KF����1���S��,m�p�iKq_s��<�O^:��m?��,��JRˮ�������I(r��sBhkP��F(^�q��i[��+'�0q�Sz�72�y�P����h�LS�ү�b^^�;�rt^��՜j�
�k)�3�n�D��mpP��a;>t�#Nd�����O�ـ8�q��	����g~�Z>�M0��c���luf���??����h���v0?';4��Vb3���͏OP�<�
����Y�>�]�FW>Y%��؅X�hȨ���m��i�����4�AQ[=t8�|"��;���r�b�L�Me��<\W��Z/^��"��J�`7� ��8Yqg�@Yn ���&G������{�v���å݈�� p����fU�u�0|U��G�~����=��z\?�g�^��%��ɟ����A���-_;���f �s�ܱ"紁����Y�6��M��ܦ�v.��f�'��"�Q��Jǫ�TB�#��Z��byVi�yP�z�t�P�[�̣[��#����B�$�=FN|��������B�#��Ƙ+�,h%&
m������0
���� �<F�Ò"�&�ޙ�K8�@?�/���ʍ4�I/r��C��@���vB��l�`�N�������o��h2�1�""�����T��b2O�Ǣɨu���A{r��صR��3�mfL��D�]��$��@S�%X��� sG4�HfI@To`��S�l?�Vlӆ�2_x�M#�c�j3�w"~ςx���`V��m^B�$��!0��q_S��eB�̈́ᰛ�[_����������g�gy������|m�X}utz����K�_=�6Z"`0
�v�zݮ_A2!
���8F�LB������0�Zfb��w8�A�q��iK�ٸ���^��?��p�j-��/!V4�1��9�F�`�o�uECE�+hN���Fm���P��C�g��ӟR�=��b��%d
�ivZ��+�U�����88��mIܪ��p$�B�����֛q��Ћ�6hm��Xl=��99�r�ĕ��U�p�W'ԓt5�7ۏ�XI�>���W�[ȩ0���8�?��m�?��)F��58���iJ�����Y�׸5��>�j�"%;�-�P��[�^ ?�����e��(�04�+ƾ �SveY���V�c/ZԨ�?�j)���'�:=�p$)Z��K�H$�ha�\Ϛ��1�HN:�L�U��}��F�� R܌�\Ǻv޿ C{P_���k�[��Ɏ/�*���x^|��+�l`�8-=��Ts�Թ��F�C���zu4� ��� !�+x\@1_)����v�`�D��n� Bo\#�XCU��GL�kO���>;+��,=fdJ�EJ� n�M��.ر��M;O�C�W�)ī��gJ���7�]�.{Ej�� f�~��l�x���r7�O���p��*0���Q�[Ryl"��4�Iz��Tp�)�h��1�v-�d8��8�u(��ÿ�׽��6�<3�=��1�a�UA\��{�R���ݍ�J��;각)��=\��l/�78�3�l�_7E��d�:���%J1�AÙO��0h	x�DL��$$[��W��GD\�b�K� &�Љ���-w���О}�7җ�X'�޵qL��~�x�Sus+�ui�r�x��`����eO���V��,<�_�A!`|`z�ƿ�6�I�s���̓ȾDf�"�s(�H���y���'l�Dǣ�o5)��ѐ,̐8�R\��:��ǋ����m����@�'��l/�^ƙK돠R!�|I ����3��k
/�r�^�QL��6{�S��4�DY�"+�<�tLa"��� �y�(1m)K��b��W+�>��
?ť�ڑUb���E˕���|�k�v5EI#o��wB��+��F9ر��$���N�'�ۂ2��<H�����\~�łš���'��b��{-�4���L���c��8��(:������!���'�J�����<�e���2�Yz��N$el瘲guF��X]vM�<s�ɢܬ��-��*+U*�z�,�*X0ȃ�"`D����9(���g�º��'{B���+u��2��4�C0݄y��y�ꥀ��.㟟�-b%�5�S����� ����0���|8KlAGK`��-�*��'����������%n� �+�?|1�N��H`�"���W��C���A��8�g����t>�7T"���Q	��-�~GK����0�o�LvM���^a�r�a-(�h:�-���&4�9�W<X�yI1��
(�(y3�])���{pR(��
�Pݬ�w8�몦�6*�γ����W�k�K��񴌁����T�2�]�P��쩗I��&Tv���/;�Ƹ����������޸lB(|��Չ�FM�'�q�wؠ�߯�1��k��S�1�nЭ���$�*Z�K"��`�x��i����d�t^��q�M���ރ*���5��>P����2?R����������4��Ӹ��O��вR'uؑLp����S�x?!�d��$�HVW���?9z�S�Z�R�ŦsEj�s�9�;��0���/��y��<c�'>�R���,����lq$�`�~�[�k�S�B���o�_W;�ֵi�+_D���9ኹ�_~� ��v�D��j��kG�`��>��q�U�4v�bah���b�P�����0g��I'� Ҋ6�3X��K��]�������;��7f�X�f �?�B)�=aR�Q߇�����/b�����6�[�]Uhk�t=$Qv�����	nYj�O���W��㍁QO�D�`�r�]�|�î-MMT:�>�u� 8!LzO�@�Yd�s)y�gȘn�����"'b9z#�X��� .�F��S��.�Hw�,���8�1/�0���*V�$��X��+U
�m���?����ঞ}���h�9S���7n�� ����ݩ�(W��9U6s�F0�j���	*�)���X���3�Mc@h�2!|b���;��1�-咖h��73͡G��;�a��l�a���j��J���Z���O��|�n�H�]��"!�wlJ�5s'%h���9��]��}-$ߢ��y�jj1����������F�l��>�>�ǪV�?<`H=(�t!)OrN�#泓龄��4E�Z����$�[?�@��QO <1�)<�I��7a��p��6P��ʿ&�9�ű1c�2}��~�C�
��u���O�T�Upxa�Guk�}��ٔY��P�3Ůgζ��a.��e��t�7jbv	:Ҥw6T@�m!x������?���-�x:�'-,�vX,Bξ�adi+}c�����zD�{�%&%du;'�@�=]�d�ʏ��[�0�,C�|_�^��9�t�YX}7ݺg��y�!�n�n�F[�r�S�N^4:Ni2�����;��%NaB"Ȋ�����t$��o�wY\I:��JD��2d"���ߣ�^��˴F����!���0�o)sA�bf��Nn�����(3��޻H��S9�d���r��M��+16�9P"C	��S��F�hx��%�C�Q֚'W����8<}v���䆇��^�֙ �'h�oq[%��ў_���f&�-����f���nj�+:U����T�����V�i�1�ǬK�=��1�C�֟��d�~���/�y���tLI2xӲ���,�BiX-`��1��5�柯.�����˗� qG#��XB9���r������q��X����|�V���)���:��!}�d���o�����0�E��}͋�Ge �|�mY���� �@��Y����Ӄŭ�(`�L��enG��y�w7g�t��-!�պ	.\�ԭ6 �!���4�&��ߟ����ܩ��� �v6p���\v4LFE,E�gp°�)i=�ߢ^�*��Χ)+$�ww�?�K!o�;eE��t���0��!���/��*�U>��&[�`��EXPA���AI*���℄�ҲJ]5���g��Oa	�њ���Dr���y�8�c �6(�ؕW<����j��q��OSL�c��R��Ь��g �>�zY�kX��؜㔸�;�j0�$)r	y��A�evt�	��q��ʗ|X��0��u�1�w[��jU��|i��R�,��G8��m�z�T�E�:���0%	�ׇ���$��}CE��A<T�"�T��}�TE�� a��2Tg�p�r�RC������|;	㠎�oV�lV
u�$d�3[�8q���p�=(� 7Ǽ���0��r��?aѰ�H�S�
���7�!����AF,;�Υ��|tK�-��)�;N�����yo���?�0��xG=h���8����W��$sl#�@�[�ja�/��v1�\���<��o�>z�M�����1=\� �o>�����3�PA8pTx�0�R���t"�����wa2��Y(7WΎ��/l����o��o9].��h5���T0���4,�ˤp��\j�8,����-r�?Z�ƾ�f�3���Hc��&�;�mܪ��#�Ǒmk��k<��w6�n��T��L"������'�9JW����O�f��ȩ��Y/���:Td����:�'�TJ.�����W<nW�'l鴅�eu�6����hV��D[�|6Lf�lqq\5>�@���2�_ͻBl<��U���[��C2��
�~�������tå�`y��@��d��4��5C���h� S��Q�2^�Q�@�m�6Y�
tN�QU��8����<_��0RZ�t��3($�Z�����q?R�M�sqo���p�4���d!0���ly��-��n6��f���9�8L�-;�� �2����s8,xmt3�� 0���L
�Ab�(�x�W��w���$4v����X�_#e�.w���4��� q���=(�T�o�9W�E�ˋ �=�� �XpF ���>X�nV�:�~4�H�H����7w<�F��/�����f��X~Z[�(W��#�%iL�#;�����+3��V�5���d��#<��4_@�8�:7Y
���Zp�����H�?�G�`bb�1��b��]-� �O<f����9N8������1��p�Q�	�(׏4$Vn���eɪ�$�5���bz%��_�[���Zmx(Ђ;�y�p��P�m���-j���qP��w��v�#��~@dF�[f��Rk��������ѱ	�N�[��(�H����&�*�Mف���|���;v���F���b��~�����pF`e��P�Cύ�ٻs��j��f]Y)=Y0�r-�Kwe`2Х�`����!�uzH�F�5�Np�D����)�z�wPi��ɉ�
p��.�]�%�!��<0��C�f�U��RS9��u����и;,1�� �RU��:̓�[��v_Tu���z������)un���s*@�W r�;�J���t��qH-��ůg��&�R� ���
X�x�0��H�ே0�I�����1�x�ӥ;��L��_�uj�x#�B��5�ҳ�笃�������*��l�kV%[����7h��~vH^���=R鍐y���&&�B��������KhIw�&����5zk����X��p������}x�>X[�e�ڐ�=�ݥg���?��n`h8:
Q�V�f�O�s..�B�f�Db�[9�;�
�w�����T��c5����y��P�_]6���LK�C���P����P�A��Q����I��u�