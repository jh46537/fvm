��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK���ʗ̹����#���)��*��:bE@�+��Q����}h���je��UAM혅�5�֬�U���9�� -	�nn�&��!��I���s�O�ӏj�_*���;\-����i�S���p�����h��u�c����kW��<��6�A�`Y����W<%�S�-x0闀�sk�
�_�j-�NIԹ�O�5�حx�Ү�����4�nHG���R�REH$CR�FKg��i�RwL4�>���e�-��;��\v���t�_���>�,��/"�����p��g*x���W�?\�%�&f�>�Ӆa`��:��P��k"F�^@��gk���9q�&?�l�)g 6S�
���l�N��*(p�݉��G3S�VG��3���[2��Թ+�J��]�b:w��6~ӷ���A���&�'"x��jQ�'S �v B���r�OA<�Q�����߽g�fki.��nsz�3�<�_���%='g�j��R�^�R�����E���F�F��h6� ֠�C|W�Al�8�M0����Z Ս��[�	�dɨ+�ݯf�[��ʭ`����S�##�Z�h�5wi��;�� �Z�wF�篣�OV�
Uȗ4����,�m�\i�N�э�#�y
8��[���Ap�юF���� �p�zeu8nm��qt[�pFr�sa9=,ˁ/�kr�t=^�T	��_,#����ىM�����6���X�S�ш�|e�+}ȥօ%
�-AV���kK����}!J�x���UTa�SՒWӤ�����S*��gE#����b�֠_��R}6���׿u?�;��.��+�Y�2�H��7o.(�ꐿ����"�"��\X�=�]}�M0Ư�>Y�&�-:������I#̘�a���^�[_��흇����,�'PB��N3���Rk=������aZ�V<3�c����_~�zIE�dgH���sd-�/�&Z;�j��ȱ-����$Da$�yJ��K�O������	�$_8��O��[JB@���a��R$ ����t�ڝƟzF�-񨻿��8a�oS�h�����X�#���0�)J�|gze+F��m�&���X7�e��fW��e��|���!B����k�S7�!|��dS�_��^�Q�k>p���6�p,�1�n>���KLWٹZ�X������`���D�Oz炃��U^g�����+&���F$'?ky���[spNz����*��o���nB�]��Q-⟵�ȹ�t�4&�Z�8DQ���!���<a��Ž���}٧���muGM�@+���0�mUB�Ya\���S�O�Qm�1Ho1)6#�v���a�5lA#%Gi(V������C�ԍ)�`Y ��J�AE"5�����k�|G8�6�5%ކᑳ�e����)�^��a�����i�ݛ[q}6")K��>Lе�&���-�Q>�*j.���*		��{`�7�<y�r2W�r�V�-�y�l� �%{��Y�|��P�rҎǲ`��9Y]U��FI��l�k�RO��"g^�#½��))��j>oO����m|H�%7O��ٔ�s�Օ�.�O��H�ut�̶��U��%iN-ʿb�Z_j���l�J��`6xs���x��j���ھ9�ެ/�sU�e��m#�c�Q
���&@�&5W��Y�[^Ŏ;m༤7��� h�����&��%>�<�`%E[�'	��.v�~�X0�t��`��D�){�+H�/tY��+p�C�����$��b���5]0��w/	�KL�d�c��>�*�ɚ��3H5f��9x.6Gᦄ��g�T�\���P� ��^Co��R����%ᨧ�X3;�Ι����Hl�<z��,�l{u(�Y��j_|��C�c�Kh�r�3�l�/!�)`����cgm*<���Yᕗ�;��E�9eW�����i��@��+�v��Q.��.���#������ŗ�A��SU�����J���1f�Mx���%,�C���O�B=��غ�C�P|�"Gr�1�?#���Q���9YvrَSDV�X4>���|rWj����L�j���EQ���];���0�ދ�U�Q0H��+��ts6r��9�mc�g��z�_Q,}��4=-���t�������i$�7p!k�Zq���T���6P���!4�82#R������M*꛴�݀���d}���E�/O�r�,VMޞީe�ǭ"A����e�,|�3
H����t3���:��@٢d�_��PJ�a�s4F̬�Z �>t�P�G�3��!��:9W�������=�(����xYK�
��	F^���rG�=�3��g�G�|�0G��Y��<�5Њ}�2F����D:�-yơ��J�y`�*����,��8��:g�9LZ:Υ�x�&w�O�! �LN0_��Sd�kg���2�}WO��7���w�@~�6[:}�2���h2Bqӟbv�I����E��@TV)�v6��6��aT���d�Fn,v|����?
,yFt��]�N�~EaS�c�O���>m���J( 7Zw�LV?I����(6�A��ԿfuSy6�C����:���g��_p
�6�z�&���W��+�V(��6���^��e���!���)�]�m^�K(j�8���y"D�@_I�G� �P-ɷ�g�����u��h�����y���R?r����b�8j���$�B�[`{�|^A4ͅ��dm=Vzif)B�Bw �0���M�!p-���]W�8�[Ȱ�.Y%�4�Y��M	��g�Xw!2�x_ �dH?y�<Jo�-��jI�+u>몛*�7��[�qWAަ�|u�pҶ߳���8��DK~�=!�bg���1ZP������ȴ��<)��' L��n|��#�g_G6����c�X����s�W-���	�֋��U˧|��Ǩf�>ifPK�J��RԹ�ͪ{4ɜ^y��z��2_�"�lI��y��*�IF%�T�K(af���jrٻ�Y�-\0ʬ-��G'GuVd}�w5��j��}Z�i���W�@Vp��J� �uO ���Hu�Na(��{&��U?C,m�X0I&M%���G^,^��_�4P6ѐ�G�Y_u��vC�]qP8�!m�e�;�i�BV��bI�n����B!a�6�@��QiM��Ԩ���x(���C���X��J�T	c{K���R�$�e�K�.� nڲ�cV�Π#�b�ָwD>�����N����]i�~�Ry1��R�U~/E'C���E;Fa�^�Ե#��ün��`!ҕ#XKV�1��~������ �uw�������@����2�&�߄�;]��j��b���F4bA�f�t������h�]Ly2�����X $�]�d� ��|V��n�?"o���#/bX9RF����j�A��"�ei��oT=�]��Hj.�rf����s0R؎nK��Q��K�n�9ɭB��@�fݭ T��*즼�! �\��>HǝL���v<�đJ�
�\Ć�����+��(e��@hb/�q�tr� ��ޚ�z$��!R�1R��X��z�A�𻍫��b�p��9���\B�A2-�=ƴM��8/�$� -�[���o^꠳�g%�|�;����\��@yVK�\e0;mUZ��ns����D��&ǺT���V��T%�$E�r7\��ݿ҇l�LRo�en�0�i����Ž�u�$�$ϻ(cvC.u2�$��5ic��%(�x�Fg�_�;�G��G�ѱ�'`y�(����|�`#��M=�'����|�ScU	W���"6�jwy�qq�B7�������#�b`6���`&S+7���C�:��f)�>�8ʸu4�i���A�p��TM�J�@\!$�V�����N�j������J��1p�<ܼʙ�rgb� ��Y�J�5�����^7�yC<��/�@��F��e�ʢ-:�5�Գ��Ɲ��s|��\
Ƞ��E�1�s��7I �c{�|�'��6����Ԙi��)�R�>�2���U��5�L�rV�)z+��@LT�
"�eZ�mG����ݖci��5 /��X�6ל6���\E��U���<4ʹ�m����4Ć��4�0��7$�nd�K�I% �8���Ȳ��فK�x�D��kĲ��8��7ɦc��;�:ޣ�uKL�R���*[tU~���xz�$��#����@�U�2p����Ǐ4R�,q��B�~*��/4}X�~���ق5���|x�8���n����^��#Ȅ��u���"5����t�U�&U����oYu�MV�l�jbS�C�QWO��'�o<^Q ���W���ǲ��I�����1�2�?�X�
���O��)'i��=�;��mS�Z�g�G�Y�����6�F/��(I<y�t!��8�vIp3W���įx"J;U����g�<#P�E�	^�cY�7h(GLi��*��}���D��8 �-��A<^O���+.#]u`���J�q�jX�=O�s���*�t�S�Fc�N� I���w~q#D�Z�#�qe�S �GS�5d�@|�����9'aįl #�Z���;�-�a�ih�lR�^��B����Ւ��oBBcC���܊G{j��Z���d/���d���{�/V�������Ģ���� *݀[��̸��8�ݮP���w	���4��/��i�Ӯ�M?�x-��%P�)S���KH;���D�j��8F`��8�dx��S�Z �Rܽ�����/9�M�;I�IN����-J��RJo�3���u�iH�pk��ls�o��*�A��B�ߩz{'�k)���&���攢_;��Z����wZ"¾� ��sq�;�l���H~N^f��E<��<�M���t����Pl�4�o=J���/�L}ǡy8h$g�`&cb'MM/u#�c 'X+o�~=�%^T��?2���,b�5Iv��-2�*}y�!pi+�3�o�-B�d_%	�8�-��<i�>����o�q��~R^�Gmxî���M"����%�\���=� �ݞ$��-)�4?��۩Î�p�����Y�UR���?Š�e�Hۓ*����TqgN�-�I)�֞5�B{���#=�L��Ը�Pg�D�~Z��_,�(� ��Qg�V?���M����Q��8]�?�3>�8��h=�]F3�7��|�/�7~�]���g� ͶL\�yc��0�X���`��ߔ�:QvZ�� �&O"�TAo�w���\���d]È��sY;�����ء �a���<Q���'�Az���	'uV�`��U���@KZ�"��o�("	>TFτ@O�[��e���l=�'�U�u�Ud�+�% z}t�㦲N���N.S���Ja�A>$��i��=�b��]xلk�Aok�щSQ��^���W��Ɗ=L�E}$T���{�0�F���ŭ��i�C]N��r��qWÊ���+�7�f0Rsrn"��|���A����t׺����8����y"���x\����S�B��,�+�Y�@a�rц�Ѵ_FC&�Cϳ&Ʉ�F�g�O|�����hI;	tS��c����8��^�� b4�i����{	n��6(���.HK�VrpU5ݫE�D�ɑ s-W�,�Kk�E%��7��7����F���:CLB�1}�Q���2���1��]�8��l��c��0���P��Y��K�4E�3��,���ͬ䑇������%�}�5�4'���Kxj�xu�y(p@_����Yp,CT�Z$�f[|8�fb@Tv���7;qj�=1��p��M��Z�7�s�x!�tr���Q�y��-\�U�F��6��cy�ּ��f���U�ާ�̽RC>t�`�]p�o/+���V�k.l=�>!�/��[�ߛQT��D�B%'�������
FOG��!�	70�2v�%�V!���c��JRz��fa9�Z��̔���ҩ�����������q����-�� ���SY_�Ҳv��EL�`�bV0G�����ԝB�*s�e�a�6HgX�å��~=[�­8�$';y�^1}-��Mt)�Gj���U46�̳��&U�I6�/����
L��pD�\����+���� ��Eg���*�#$�Nh*8{��a��Wq���K��E/t�7�0`o�MMƝ&Q'�aD���TN���ק�4-	8opﵲg��t��E�?e���jl�:��2(%�r))k�MR<.�)���<�Y���m��D\6�m��lN���l9�m��F�k��2���L{��ـ�a�m_��՟p) �RAf���+�B`8����$F�z����|���k�I\���<�@�%�%2�e(��y���ռ�f�r�����y�A6��r����Gm7)��R`o�U<�g�,̣q�r:�M�r�	�����@��B
EM,~j��IM��ϺD67Y�]%���9F��J�;b�C�uZB!�Ư�b��w���� W�I��?��,�~�x���>�w��j��+�SkPZ�������*8�}�º�]h�w_�H�G�K^���I���N$�(%Z��@��Ƞ���|��vlզ�u ĸO�߂��`c���z@>x�%ѱ�S�-��U?�7C�4�~�F݅cs���e�F��Qɽ�R�dUY��2bس	�C�`�9Ag�+߈�g��pܐ��n������}�<ү7���:H����f~sn�K��L���oSĜ�!�u_p�
�C�*�׆��uǸ����ģXm��m�T@~�nF�X���}�U��u���F]����R�hT�� ���g�e 1Rt{����q-`��q�<�.g��"9!���-*�4�F�`�s*|�r� �ƹ�=:[g�xOJѸ�1���S��q���x�+�:=�?�]�啒�g��Ef��V��1z�(�����_J�'��!S�)�;�+�=��2�e�Gׁ����^<�@�'��U��bCn�a@b>^D�%<E�'`�՛��`
���L
~���!�,��_�c��I��6�ϡN�-T�}Z�7g�聖=�M<ޜ��xL����r$��)��Q.�(���m�C��r�h�_D8wϹg�,�����7`!�4E�ɖ�Ǒ�ç� �@�d����t}�����7W�H�׻���)	����~X~��U�ܽ�N��������b�'�J��T���v������8�\��Ʋ�! �i�f�=RZ��S��;	!�_��3�b�Hǵ�f�����*{�x�N��f�p�t	��$]W~D��L�~�bI��2M���$.��I�-`_/y����^����$�֘Fz$�e'�(�@�8IG��)�u�þ�C8�I>*���'��/酑�a�+2���^p�-̐",�T�<�'�f��Rw1"9PC�ȄNxi��E�>Sn�?q2�J~�#����>f�c�e�F_�wk��4"�G48]��=�%o]����P-ؚ\�5��������H ���:d[̔����ǍʩO����ؓ�$XH��Q,I��ȳ��,)�,���<	������n�tS�p����x����gλ~&�-|�b4̈́�
��M�s-ڼ�K� )�g���8"�H&�`=���q��lGK7j�����b����Wt�����k� ���n�'N����|�Gپ�x���ɳ4�z"w��N	���~OZ("����P��q+�z+t�ӻ�N��`�R�@�2��Jw4HBa�.�Ϥ������ˈu�vL���i����M�7�,E�M�w�nu�cwA�|�x	�#a��5���W����]Pb���\�ø�d@�k���I�\�%LY���CEh��N�)�NQ�JP�&�q��~̍~��O���e�1�k׿xך��3!?K=��C�B)ԋ���op��[��-J\/3�"�{���R���V�eIXt�	M�C=�Xh{���$�%��&���$��I�e���7���m�
H�,G	o��qW�y?�4R��������[R�C<���4y[���M9�8�9@+Nӧ�f��������*G�p�_�\�?�49Yw%N�'h�0��ry@���k�+>�_V�L2i|�QxF~޾6 �%"d�1g�M������!��W��۶o)+K�Fm��u���50��G�А�ʥ�OA#�Ҍ�����	iS������O��=��ɩ���1�%z�7E�u(�OZ�~wp���TT���NZ�S(�2J�N`�(�,�~/��^��j<W��FA⟱tm������w����t�7���<�"e!�2��0_/�sNx����˂�	WC;�@�a/����NvN�jB=Vz���r�K�:<�oT	"cM�a�X=3�<6֝���ȅgz)(�-?f)��ϳ3wi�:�В���r�j��b8V����L���umv]��t�	O��TVǬ��h�UK$5M0��6��z2� �7;a�)���܇���s|�b��w{ݵf<�u ����4N8/�-対�:�w������I^�zԱJK����R\C\B��c�&̺Lvq��&�V$�:�AVݷ�sv��,�z����~�}d�(T\[���㶲��Ȥ7�|}�]�^J%�߳��q�X�&�>�ʖ�A���\�c���\�C���m\ �k�O��ԁ�5�PK=N�$�?rH@{mAHo����k��'&y�/Ev��5��J���N���%p�X�
-��&^O;Sș@��6
��~ͽc���a�Y�Q��y��n��R�����ě��f��[`���uĳ�	�m�GV7���v��抪�x!����Z�G�T��l��NX��;H�0�׎
+���_��L^-� J  ��j	��q�*����M�ϞY���Q��ܤy'�)8��[����ѓ/_�A��Cp��Zw�g�cfx��YZ��\ðǉ�a���鋙�Y��|(���{�h3�]�}q�7l����ȴбr�$m�\u����S�(�r�Ƭr�Z���������R˽����v��}���AdTsZ�o���y`hvWEZ���
�z�`���e�э��YX+t	F�B���`{�NpAd	�z�UvNz����M�/�l�2�)@d<�+������I�O6 �t�4|Pz��x��$��^��:j6��_��@���݄&��'i�Q��	AW�a���O����w������>� 6�J�!c>R`�rLo ��A1��Ϊ���*�&��3JȒEBD-�3U��|��j���BN�cn1�F�un���o;�[�N�8�X�M�����J��yu�y�;�,T�Tl��^U��i�:o���tr�7KV樽2��.���9q~P4�H!����A��x���I�O��F����� F�04x�>���\�B�������X%�ң�!��u��B���g��Bu/Bp�����'+]�T���o���}�|��q
X��;��l{�]A��R��d��X�h�m����* X]��(��l��PO�w���,-vN� �j�G�a�(&m�S1����&+Y��1�Q��3�����L�C7�����<CaC��"i�}V���o���4%r����܉�Y�^8�@���7�� ����u�,�*���������t'��n|��XH�z�6��_RH���c�v���6f��,����V>�\����d�b#��P�B���N��/��bgc��9�tD[E�nUĻ֌���3&%���i�Ö�:���tS�0Uy�cQ��e�ݼUH��s��ۧ���W����v\j���ey]���|�������ܮU4E�.�O�Ro�:kXO	9hY���NWs��P�K�<���7R$� �sJ�O�R��l-q9�Ep�3��cO������b��h�<���?QA��l�=]�c�v�$�<�Fd��ndH�W�CV/
rc{����zo���*ε����,��h{�I�|�^6��r-A�P*ْ}辸M��r���r�G]A��6(-�B���d�ُ��|�Y���L������|���K|��+l�����:���:(��@��!�t2��� ^�y���ӪZ�"���׏�E�xBz��l��7��3�
�쯤ds�8�}G��XO�C�0xnϳ)7��(�\��֞.'C �X�fkq-w������[;,Er�k�R\�;�q.�oJ��nR.���M �P�X�]�ೌW� Ca	r���$Na$.��|#Ri=X�旂��Y�?Ҧ�u#�#�?#gvO�i�3�*`1� ��W���q/p�rf*��]/L$�	x�E�]�f���I��1�.>����Q���}��zp��w���5�L��[� �����BMAn۾�z��j�������G��.c�LO���������
P� @a�*8�7�=\�_��o�/�����Zp�F	psYg,�J�#ܷ��ݰ'�
a� ���\���5��)���V�Zڞ����Pu(�k��RK϶��[��/�+1HT{9,S��H����޻^U�)G8Pj��׾����b��*�&�fk�z���]��)b���l�v&1E[��@1��9��� %���+���(v 1��/	�C���k���AO�o���G5��@��;���-s�6 ��p�����.`晙��\�>,���Tժ!Xb��:�b������aN����l�)�@yE�b;�i�#s�<�=:ޟ�g�$�� O���\#�t��A��+�	G@�P� 'r�1�6&+�����c����w�*���T;JJ�/�'�� ñ��iY�h�����N��Gy���C0��a���S.J[�����EJ�E�Xr>�;��t��T����;6��-��V��'��D��P}3�B�&�N�	`B%�G�e�|p���Φ���sࣷd]9�<Q�/H-�-?�h��9ӝC�x���s�`_���N2*]/���}0i�:C�X�L^���,>���/����\���I���(h�{!j�k�Fx��3�׾�>��ܾm�G񺺍�\��ܐ������ѥ�{B��b�O���Sز��E��^9�!���x���� ����y�lp�q�B�һ��L�6�����P>�WBNd�Bʓ4A�����Bk��[]嶢�W=�q�FzLY3C��wk��[y��`z�P���E�B��O72����t���ZSsk�μ'܁��L��X�u�`p/���z��EB�&�2�=P��O�	-�����Ϥ���as@�u��)�1�������j�bܮ/oD0���?�e��В���ٜ�A�_���(7����%�.7Y��Y�(���R�?�Nkl�.������n�;s1֔��t������<KZ^y��4`��|�y��C�2k�GΩPk�覿=_Oa�G���S�U�N�G�-���օ�Xv��z���ܵ)>����ъ������t��RW�j0�d�w��F<��{���~�'7Sr������nG�3�5~m�gX�L�.���;F+�����4��^ Ԡ��DW�����0?��k��%&���c�KÎ9Y^Ɏ$)���*��7��,�)��	 ��L�m�sq���ܡ���ǭ9�^��e구y{\���+����_��ׄ��d��|������_X�e�*8�9�(��N}��~�u#)�fq'���a?gS�6��Ő@<Ӗ�I������2��|��V��CZ~eu�I��Y�������E��LH�H�]�k��`�t��Z�5�������U�a�����.&#�d�i�~űG4�(;C ��`C50FW�K��>����Szm�1p�����x%���:K���v��%kKG��4����� nT�x�'���ӊ�~�B,�z3`�-�Q��P�jv�~RO����`.����) �s���.����O��)_�����SWz-+�3�����K�D�邦i+8����̕(�Z;X��"A�{ĭfZ�OY�΋_����P��O��
���s���.�e)|�쳦[���O7�M/�[�}3~_�WO�̧jn���S�b�C�o��׀%S��K�TJ��^��s�s.ئ~d�O����-���`�%'��m#��)�P�DW��Cw㮊N�W �K0:]��m��!�����/�`��"�d�4��~� ��q�Z���SJ��������7��H�?�܇K�Q���Fa�	���K؆�B�WK���q�	�ɓ瓸_�S�D��}RIIA�YѰ��G��ru��#W�������SE(!|Kn���(�r�Û�����/}�"I���1�;��%�?j˩N���n)� �[�%��K[i^-X�-���gX�a�����_ld�@�u����zC�9Ⱦ��Չ�Y՟��iW'���{�Hs��;ٔ.�%E���Q� 79�� �Ц�m�&{��T��Cu�U��������^�~
�V�G!������y�95�@=����a.g�%` ��7/�Ttr,�L�1�`�:��q.��TE`��x��Lb�������`���g��r�i~�����g��� I�����v��p2�X��kH����U�B��f�#'.�ŷxKDi��q��n����J�ћ �� ޣ������ >��V��'��+\N��W^%q�����P���C�D01��h����F�m?݋�4�Z#�g�tA�/��W�_��]�c��yns^�k^��A|IW�F��xm�.�ٗ2�D�*�һ���C�n���U��a-b=V���<IH/]��c���c����e�s�oi���nt�
�����uބ�BN��(���n��K��|^Jk-{���:#�"G���i�<tp�-'�8Kd|%��M�X�E0���?ڻ�E3�3��^W�ɻ�E�e!4��動�@��绬>�_	b(V�z`�Ǔ�k_GƬ7���[���j:�{�A�i4�O�2T��¤��|4'"�ݺ�ֽ��+s�
���9"�����l`�k��Q2$;�mŞH���<� ��̐5��ܾt�)`9�q%[���_���Ib#�k\8�Ȝ����6�8�
�ώ�T�gxf��DmK��T���|�ɇ��Ș��;QA��ZYI�;�R�R#^�Q��x�d�~ͧ��̲���1�G�+��ӭ�_Y��D�O�`#����dy��OKM�s�X˞���[l��D9"-�ה'q�?��*ps�x~NS�V�m�S���7��h��	�c��)�,ޒ�4�bp~�y��Ш_����Q[�ֲ�(G��,����dq��P�C����<aW��@a�	�^+�+�2��)��0�Zpq�`����|&Ҟ���,hK	�mo�I+C�`����
m�� ��'"j�Hѳ��LM����X��� -`ȔJ	�*a5��I^q��%��q-�Qe�Ё�x�j�f�F7���$�!�F�ݷ�J,�߅�m��,&����h\A�i����S~>�y_	���'T��W�2cS���1���
��Cd^^໣p���tbme�짤W�zki�t�X<U&�:�39�wь�[������#��xoJ�{'-եJ��Ad"�]g���#��>������b3̵a��
%Dul��[�@����o���c��^9A�"=�V����>y��;��3q���I�;U�����R@�w���/�y�z�DO��?3nQ��e�0h��[b�?�<����9��ڜT��{���炤;9���E���ɩq����r�R	��R�펒�>����ŉ�]�s&zlx�#�I�9{��"��,P�"Ī*5]��)h@w(&�7���`���o���C��̔����vo�8���y��9(Ll��!����Z����yf��n������'>�kP��3WfĂ
琕;J�d��R��Y�^{*8�C�''~���u�y΅��QM����TL<ʤ��C�Ȩ
�g�:��
��Aa�N�h{Ȓ�%u����2�x
W�cPP�Нajy�AX��zo1����W�_�A���1X_�Ԓ-y[j�k���f�����4ѐ�w=��>,���O�|1�F�?p=��b�Hc��W|�j�y�Q38+�Ki�����6���Ϝ@\M=3�Cf���F�9&4�ѐ*�T�'T��^cԴ^v�2��CVt��-QƋ?�t]�ث% ��ǧ�X���pޗ���k�/�
|�1V4�A���g�`��Jr��~����R�g����<��E��5ƥ�(|�'��hQ>���^��E�ę��שj�$/�>0�Ho�y�����o��M�lVȄ ��s�7�A�W��z��g�G�&��]9�`X<���_*0�A�3ٮm\�B%A�$K�� B������m�Ũ��+~l���}+�+�\�Y,�Pȟ��5�����.-N7Y�J4I!vΩ�^͕L`-@	�,��:��xFɉ@�;��6���a�M�9���h�p�ܞ�ߴ�U�������hi��NV�
�#1V>g�睹�[@���x��q���Ġ��i�z�WNk�mx�me�����
.� �r�x�	Df�u��j*��"dĶ�}�V�ؽ�}�n���_Z_g�®
�g,Y�~�tU�C�Dx�So�Mcի3�ݷe��DR�|�*o�5&���'�r]]�`���W���:����+�q��;+�,�=|�7x�2s�9�~ *��7�H��MP�-Q�ܬ}�[S�;@�������PN3��Y��]����,�`��}�6[��Yn��V����&�\v{$��rɤ|;UL콚���+�4K'��/�\��|lh+���6I�s�@��O���u�/�ڥ�%\�^�r��2P )j$�p֯��u��O�:1��0u���<��:��0C��)f[��Ä��h	+Diɔ/E�E���/9 �:�I����U���Q�@�MņM���*HxRJ�q����w��B�l��E��
>]�l�y�����5�U)Y��E�1L�=�ҍBr &`IF���o�6p��h�����S�z	����V���S+T�_����]�V�w�?^�K�>d<s��;��*��?�>�r������BU������F��_��xUT�T��
�u�l����
>֞l�lZX΃X�^�4	B�I�/J��T�g~I-��
��=�h�a":��U/�����1���\�["N�Rµ����&%���^�C���L{�W��;'����s�|1T�f��D�'��w�U�˹��{�\��U����v$K��
�b�O�����]�4舦�>�/Q���T@)s�mJ>f
5�.�p/9�y�kS�1�y#�,�8�5�!�~̝�M�N�5i�ⰰ�a�����I�@����P����g�J��Z�*-x��K����Þ����}}�����Q�N��}`�V�2��_�-c��N�����[��/E�/���5_`=s���?��}�I�'�_~���J�5�}ki/\7�ˆ��������{2��-� �D����'9��E� ��Iݲ7N��Q�?���VW�=����L1�0�ba2�SWZΛč��Soќ-c�
�f3(Q �ū(�5�X�ϢG��[[⟋	~[�JN]�ʂT���EA��l-�+%�^�0w���x�W�H3d@H�UPf�2-�g���d�������W��1�s����,VƔ]R�dѪpp,�̡����CPo�p|_�t�IX{�F�}��=/�/K�@��u
�����?y��5���`��c	4��o�x(xÉ�r|������E공bޮ�ؼ{��+�>��Y9
�w�~i�U{< �;騊]�1)|F|XA�M��5�y��Ư�6${�e�pc2�F�Z�ri�{��k�<�;_���W6����������5����r�]%�����Ӆ;�'a'`�5Ԩ`<���[?`&�tR�j{m�N˅�B�_�_�G䖇�8�dؘ����g�>!|.vnc����B��;c��If�u��+�$���e,J冕�� �ܷT}F{i#Ƽ���U�Fgf>հ�L�ɋ��|������h�Pt���������4��'��|����X�$�ҥ��|M�F.����7����{�C�k������d��Ȭt�y����W�	�_+ �%��#Q����/UO�g���]~�7Q��Z�駩�J��MB���QR�qRB����
^�沎)��$�'�_e�^ζ��	L�h	�0Z�G�T��0m0����;V�e��-����2dݒ�z�;ܺ)��ت�����I��ǌ�Ұ�����!!(ָ��cN��)t���ʣ�!b��?[F X�&@;���<�ԕgk�iQf)S��*�X��C>���' JLe��1����ߛ�ؗ���y)�!i} ڪ���|�{����'�Z�<l��w����x
�CTN0��V�t�()�Z�N�ծ59���������x��"}�z�M�k����5��_F���1�	��~`IGh~��+�Ӿ����Ƈ�4����"ty{�%�{��[c��1��Y���e�k?D o��q�>K��Jy�{�;��y��<��\X`��	��Rg�De>�1�6ͧ��g���D)��[���&I��5��xÖM��1����Y���2_ǭ����B��<�m�F2�ߋ6��vl�F�j���dA�Em����GK��'Ȝ�1��S�c���
 Z�����>� �wX�<��X�͘��ζX�����9#�Pӻ���;�Q����f�S��d�fwdV$�5�U#)�� �N��-a��96�/c'��`1r�Z�����kB�c�VF�l��F�|���rN�LaQV�j�$?8��F*�w��5�}����b���Ws�� ���Y&��]U�O�<��M}ڃum�~�3�O��O?�
;�շ�,��mJ��I�1�r(\�N�uP}�%�:�Qàk-R��q/֭�9k��q���pY��ʰ*�z;����V.
5Y�l��0�ȋ=M���������ފ��� +1�����<�� }�a�!h�i��d�z9�a�)�'��O���s9�A�jo�OQ��P�
�r�z�__�,wz'�u��,�\�����#2�Z%?&2ls�g��z�邅��R�]ZH�z�yw����Œl^��hC��~@ ��K�'�j}�~6 *��k�_�-�@R��V�0I8$O	�m�� �a�[��,�e���d!����c�D�g{X�IN'T$z���_&�C���s�I��Y&�ԓ�1n�ח��Y���m�5{� z!��CG��g�1#��EŜщ�E�wLСQ���ߒ�,fT�C�y	U,a�Q,�ޔ��zܵ�n�e�!���6�#��po+
�B���H3R��2Rnڇи<�d��>SM��x�����s�~�����_�BVS�p�*���SN:����_�F�I�x��N�"�;l	m���p2}�[VD��π�pmQ���*�T��:(,�"�RI�/�-ղF�Q�|���1U�Q�o�c�B�o�&TI'K��eS��Z�m����E��
�����@��a)ǎ�Vi�{�|3�6���D��\��(��M<ܫ����'˔�.�Xc�T%�[�WB��OY݄�����d�SIP��s]�`��d�*<�-Uo���k����:�jN-���Q~
w�&9+L��Q����IEB���6�mAZ��%���-E��D���tA��y�|� �����g�~:"�(�=��e���ư������
��eI�l���	|�Y��rM�9w�H������b�s]�E��җ4�{���Į:P�&��QC?�+S���㠁j`�%1;�@������� ��
��=>G5��7;�&����c&�-�p�����gB���(�(]��g�Q��G��;wG�Dٻ�S��9�)yW��_B�4@ 8J ��Q6'�T�2����9s��N� �EБ�E}�b��o�m ������C��ȸL�Y��h�u��\���KӢi��+ 2�-?�gK����Ȯ�>j@X�L%�Z�Ѽ��jDͰT$y˯"���j��|/�Q;mz|��*�x��QXO��Bt�y1c�Rҧ�F�EU�|�@w˔���0˟�G��J, �&_H�gKr:����_�R��t,���s�K�,���v${ds�+�s��#\�������{�kz��m���׍�S�đK�ň���F�tѩ�l����Y/*�yz�J�YJ�i��'�(��� ��H�A��ȑ]��\��A�a|�g�r�:��{ơ^�6��;w��J��@�on����>�h/vl�1SE[��NUU��k���GѾo׻��2�b�[e8P��"M3|uе��SR�������ܯ&+���
0�Թƃx"�p��b�;E���N�rW�b�����W鑦�2�������a��6��\DP��F*��Ht��G=#�kL/ǖM)��Bt4�urr�����3����_6t1�2M�;�#����yd,�z����ʲ
���v]��Bɬޛ*&���-}��E���;_D�-~�	��� 3���BS7O=~Fk#��τ�\2�N��4	�k�����ފ�A��W2�}z!o5(�ע	t����4Z��
k�B�48n误�/˸���T]E�3X��8Y�8�����-��a�Y����`�d,���:n�hRp�k�i"�z�@S��ħ*�^D�L��+&ъݛ�BH����������ZnM�5p�Ţ�#�\���8	� �U�qu�(�>s���V�\O��L�e˦��PKd�bWc"p���ޥoh��q�� ����w������&��ZX�0񪓛z1���W�׌��~s�M�*��"E��<���P�;Ɯ��!2�ˤ'!X�bQ��Dp��ۤ���}�]��	9X�S��sɦ*�@���r,ǲ�@M�Zfqe|����������mNZ��f��Õ� ��p]L�شNy��._Q[�b�T��_&9�B���R�����8tG�pZXas����#��\���5?G��Zhv>a.� m�@<�?bW�,x��_�!��A��	�a��_Bh_� �\ł�|@&�!�	��ٕ����O�T�_��kaS�������,�h��'���>ԥgf;�$��	�k!��^Y��bw&O����V�ۙ����8n=G����*QM!)�"X�ɘ�D���뼰�7!�Dod2?�h�|-f۩��Z0�8�	�{��� �~�^g�Ơ�l��yz���Y-�'侔{uiG����z�k͚�1e��J���l]���<�6�Zϕ���3\,7�/�z�(y�b�
�k~��j���s��S��Ӥ�u��2�Ya�	��ۡ��b��� �� �����0�6�k���)�QL�����k)ƆU�����S:�?d�(���7�Կc~~�?ij��	��Έ�=�(�u6��:_�����$�D߬,�����j���/���2�]r7o@,�j&4tI�0��O]j9�n�D����3�����9��0�0�+j��Rڿ>m���_� �Ln�jy����z�_�*~ɭX[��XHe�ݍ*��\��'��L> n�W�����5o0��S��l�M�<�p��d?Lc��K2���@j˟4�vN��4��[��V9+���w���X��xl�bkx�2u=�^��̀�erZ��V�g��ďT=��|�u6��4D�ܤY­}e���{�̳��T�/�y�T$D����e;�h������\�1�t�-�A�O���3Ś�1d��؞�U��O��A��-w�������]�3�n�g(�����߂�'}���^z�~N�vR �0�ȉHj�O��fq�R�fA�K_O0��r��24����]%���2��vIeh_G���e�����<�>�q��ڛ�9<M�z;�$��s<ܳ|E�ߐ_X�ΰ7�(Fg�MS*��k��
��.Z7E���T Qlq��5�Z���7m'�᳝9�`�h�O��
	��s�B�,e� t��X�	����sà�mD�uܓ�RM=�~4�qo��M��F��?�n��	�"l�v�S���1]sC��揅4H��胎���~�&��[� �& �ϡ,4��q����C,�M���M��]x�":g������>ᄅ�>!��8����T��@u���18�Bb��'�1���O�^f�!��_�҈���ݤ��R@�<��
U<T>U�]�:���7.�=(	e��w����sa>$�Vl ҁ��:���/��.��˃���_3a���n4�b�~���s�Y�8[�F�dsi���o^��ݐ�I�L�:U�#�	�?�a\,�ڤ��k!@N�ɰ�~���xӅ& ����
5��e[�V�67`o�.�꩏�~��9��2�1��`sMoE�c�c=�#B�*��LF�a�<�\GBd=*�Z�V�h�����ۖ'��Q���4�)JC|[ӈna�#ӊjщ���6p:$C{�X`.��;���X�&lv�Y��W�I�˞���0�Z�qXE�(XCT��F���px��G�ڞ��#�n�-����e�&R��&WQ�v�`n A�c'�. i(h�Pr�r�đ�L���Ev���ʙ՘�}l)��~���������
/��hح���Y�	�����i�:]��l�.�6Ne�
[�@͂ʜbn�J�4�a��$>�j��/Dz��˲[��������K!]�`� Q���~Q���+��=H��?�����'}M9�/�^�Ղ7�p�%W�G�\Rg}�=pT�jacW�a��V�L|[G��2/2h�v�?�xf�Sữߴh>^��=bMh$��������2�,,� ����ܓ�醙����K��@��r�s/�d�'ICpw��,v�i�J�da�q-ch~����v,am�{p��[���J�]k��Z��S`�V̦�Ғ�>�i�jJ(N���U���2�����F��6Vk!YZ����kg��q��i>�`�[8)�Y*a;�V%�ۮ�I�Ki��u��8u����Ǵ���\�a��>�m�!9Z?��ew�������h+��v�^��g�pi��-��棡|!yfUp� �Bx�;4�*Y�?�ו�l���)~;Tw�,{	]5�� ��v��'x ��b�ڷ_��S��rfk�<}�<i�B�)ol#�Bݨ��f�<�ǹ
W����M<Uz׋�1|�s\�Xԁ�����I�S�6�Ə���F���*⅋um
���m��#6��d��f��F�����!:����k�I^���^�H9����ևY����9p�J0�;�9*�\ˉ�46 �q����'�c��\�9�"��i�˫�y��eP�"�MI��G�n�W��[-g���{�&��2�o������E������Tp�ފ]j�k��r�֛�	�g�0\��F>!7<�m��W˔����yћ�:����O�!��|C�!0<�p�|�޸�������>h���|�_�ȸ:M�s�nS�)}F�X��a
� �N��r�Yݑu���}�o�^�l��U6�=;zG��ǋۊ���
��}u����5�Q�\ӱ�e���2���ݖ$2�v_qd�@��~1/��@�_R��PQc'[P�<n�J,Qu���;kV�6�$�tRLm1�k����v��&�ؒ�r \�l;��7 �AV>����6��ݐ�2>R2!�kSe\31�'�+d	�hLx�#~~��A4V�1����F�#L��ԚU�>�V%�|��,��L�_YӅ�ָ�do�E#ԯV�q�9���y��U)=�[ޣE��-n����#�4~5��I9�PrnpCsX7�ڳ����H�������[�p͊���uh�,(�/1Pn���N�@������x�3zL#x�iD�ݡ��؀�!�%Ei^`��o�m3�%>��9�~�8C�
���.�<(R��V�+�'"�2�S�=˩&�<�h���ב���˰ ���5��󠐘���E�P�.�ܝ���D� ��*+��*D��Y~��5�h�	uQ��O����Y݂~v��Ln��5��ՙ3
j�Xy��ĉW6g��k>Ɲ�K`�f�
�:
��G�Kg�f��Р9OU�H����� �:�*�.~h�o�}H�^f���sfv��%�<�c��B��@yإ�z�w]�`s@���n)�G:��.���j���k�}��e��<T� t y���0rOGBǠ���!_ɰ;A�:�k����p��
%hH�⚷vML&�g=9�C��f*y8mB���G�H�����I��	�.y
Ň֑T*��(ތw��j{1�0��ͩ����ŀ���lA�;�d(MQE0�'�w���-W��Y����ia��;����]4�;�#z����B镓 �r��*���o(��1��6���y��I
��(i�VyO4����H�C���Fkɞ�)-@?�F�\7ԋ����A��n?28E�{�c�c��ag�#�v��w��tCϞ��L����/{�����<�O3y9$�N�:dB�<�(y�Y���!U֢� +E"���5WU�Z��@.�@1�I�np����T��pg����,�V��9$࿖�CR�t��V����԰lߑ�D�=WT���^��Ժ�M\D� �̀��:��9��8\�R�Xe�스m�
8��n���J��r���"�H�`/{iY�Ɂ�֍�s�\�H���u����H��1:�/��ʩ�K�Wl8���BI�X�<��mt��._�d��b�s|vq��9]�a���/��L��o]u�̀���&O9�ˁ�T���@�y�܌�I�)'����e�w����"�
�4�Pm�X�T�:�;m�!��՘%��$oz	@3���&��u�L~
^P�Z�.���b�:�{E0�m�*�Em�o�sV1�XOg�K?]W����pW�p�f�޵�Q�a�^T�������� YB}[
�:�Jy�΂�����5��ev�)���.���MA�����wJ�v�N��<ϡo.�2Ɂ�DŻmN�9D�pR+1�ʷ&m��}������O����{�w|O%G�SO�#�U7J5����l+Q��u�xB|���Y��[�UQ��0���Ev:ku��Z?�(!E�P3
��7l6��Q��-ş.�	S��"k�B�Ve���;O��ұm�H�R��h���+V=�o�>�i�AO�@�Oߡ�a�k�p�_( �5��|}�7c��C)���!l/��Z�A�AU�	l\���7��u�J�$Z���LInz)i����� mB�t:���4�h�LyJ	�P�x,�
���qm�2 ���h��%���:���%A�ƈ�OK�O
�o�|3�Qw���wt�J.6s\�Ix��ڙ�� m7s5��[]�������@H�a��T�, #��/F����o�,�9�� .�(vk� �
�bt������v��2��B�� y�(���iԲ泸 Su��LtO����Lد2�$#1�[?�'	�_ !I������dd�<�� �I#D�#L�����k����̺*W׀&,��Z��t�;2�oI��K��B�@�L�
�Z�r����DK�SD�+qet��r'Wy$��|GF (�K���ČX�������������.��ab2�d]P�u	4��� �cRے�>_�U���oç����;��_R�Ok聤�`���Ⱥ��gCw�3)�[x5�6���Qym@�|}�5�C�Tv*�X���=����Cq����3�u��a�?��[�7�-F	8}�_q��Ɨ��C��Ϙ��1����4O�li��Z�Ez�xA%'��]L��Hw��w�Q�^�l���U�2������46�`���5�P�`�ək$jh ��ӯ�.0�o�=	9��f��&Ȝ���J�_��D��B��:(�)�F�g2gu�[V�+֥��i^�R���1�V@|2��;�EN��ol�L�/��V���o9c�kb� {u��A\����������8�n�&7�U��j=��48,�����u����X��?�z�d�hw{�o���5��|P��'�J��'�~��շ�IEL�xi�g�RA��f�ז�q��������0 ��ݹwP��}���j�=���؄뱫��%��x�G5��M��Znp}���K��J�#F΃��ܴ�A+F^��n��V��q�[�\VCO�_��4����b�TH��f��e�nf:�3�_G�)���:>9h�bBVZƈz¡���Y��sr6#�~���T�(�j,i
���2��a�R^sD�|�ދ��u�kd�5�R	ͫ����������p������4O�J`����8�F�W�z�ݡ �87�Iƨ&,E}SZ)ٌ��3�e/�j�y�2��V^	+'EO<���T<�Z4,�����z�*��U��r(��gP�"��$��R�Z��ö\��ﴗa0������wX���ȸ�n��6e��@[f�����Ŭ(�9B(�s�לH��L�|�u�f�|��`Xs��t���`!e��.�����P��?Ꝝ��^q�ۙ����@��`�F�p:�Z��&��3���f3T)?�A���5��85N��ɫ�0k���O'����e��w|]��V��A�Ҷ�Xi ��t&F�;�|�iYgmP��p�E%K��e(�w��g�+��0O,�%��-p�..�4�Ʈ�4r\�@x�p��L�BK\�w"������,S�}4D2�$o>��@�K9���G�A ���즩@�i��͐����x���m�+�!x��K���@�t�i{�X�7���h�)�aؕ,8S�1<��\0�UqG�S̗�{;^��$���|������kj槅8�J�V���x�U�̠S�
42��U,���V�&h����G�V�X�}�Cd^�%��3"j�Nw�����?�q�B�;���t�d�4YxC:O�x���o
��A%���OT/.�M����-S���Xd�Stk~0��(<��v�"���:�jC6�lw7|_�""�%ٷEG�v�� 5���(S�$��bq*8������	宿����P���h�Hty �e"/-̒�Њ�b럋����H��֖�!2�AR_�AK��<l�m}�ւ����Z�U�e�F�v��艤;�q�S!=��ìX�S%&j�8���C@;<�pC�^5�B	� ɷ��o�1�7\��4�����
�.LPG��g�p���I���GN���V���a
� 8�넅�K!�
���Mz���K�����i��f*msvw��RGyǨ��j\DI�.�(ԥ :�$��)�_1�������KѺB&�\� �c!4���+ܡ��H!_�dgB�)�
��C"�A�JSW�.,QO�Ap�l�GK�s��"ޡ�Ɏ�w���7�>pH_���?Ǖ�y���0o*�0��pm�j\�-�L�O@QpO�(
|N���Q�r�J�A����;�<?�#R�����;@LU�oڷ�ڹߦG�NgA��ף�
�����p��Wi��VK�w���c-�����ȹ#�����8:����\���Ŝ
c/(�M>x:�e���l��c;���ߜX��*Ӆ��J=I'^��a�����ه�41Q��n	�����q�Z��69)5R(��K�m�R��M}��Zc��9��N۩�����Z5�u���<���a淝\��Oi��f�N\�𕝔�eP��f�IDᎪ�hhP�9"rMMe��V�F���t G���U���-]��\Đ
АlwZ��4��*7��[���／]�?(i`���c���&�h�m��f� I=��Y����5�!��/^G�������U�-t��0��)%���%�O.�c�;�Q�)4y�t����#ߒ��u-�>�r8�<5W���ɺ���Y���#PiQl�;��
I�oC�d��g�2�I�tj5�������=1�W_c�}�x��b*6��t�'?�K	m�3����v^ڳ�O>|]mĜ��r�҃�-����9�VA0�������B�ߴ�p�{ٻ0yFI���k�]f�×�R����x{�[����W�H_�~�^���`/9g&CV��7��hI����:w`)�:�	Z�����RL�1⸖+�=�X�`�x�xygL�	�_��>�`�Y�v�D|�0$��,����$x�MՋQ��sNrojUP�����X7?�r���
���6�t�J͈��z�>�@����h�7z1�0F�Y` @V�|�%ə������#�%V]���3��R{�I��ñN޶{�Y�#Y�KKX����e���.i��í�O�Gj�"V�Wq�U(�����FPv�r�Up S�w�4�o���ġ��V@���$�{Ko�3�m�꠮�fq�)�C:N��=
�P�H���gd�?�2�1dm�� Ȅ�<%P�!��K;���k�j!'��*�&Zw$�}�u2��D��o����6 w�Xv��&���XB�Q�M�>����Ɍ���@O�nS��/_ߜ�@�&�Tȓ9t�/���!���8MR�+�H�o����]Awk$��?xP��6|a��Ӂ�Ժ�|��Ly�	j@k[^Z�4���������#z�F7|�	�h)������,L��+���w�U ?�B��mЃֲ���g*��XfR���k�9h
 *�^����ۯ1�OH�\��2�t�»��l��WQ�L&t	��f8^�ܠ�g��Ξʢ�1@�Ć?(G=�z�HL8�J��c�ORJ(�C7ҤA�L#�R�yZ'���9�;��S������,,�aSi0cԱ�ށA�w\��eE1�ݎ?E��5S)�{l@��&��+��]u%�'��\��U��2��T�n�BJ��2-~���v���X�0�<33�m̿U�HN�5�(7�9{�~J^��H�^K
U�N� 4x�I��[#y����zfs�z9����G6�'���¾��@M���W��l,�֊�'O�Y��Z��	�v�UO��ˢJWʙBq����J��<�7�0�3V;�[i!�jdz�Ԑ����S�/��3%C( hM���4k����Ů
vu]��eu�9k=�AK��A��HJ}J�){�o޾��TG��L��+�d�9����c�}K��#A�0T��2Q���f�A_��p��!":���@��Y�[���^F]^`q���Tfk#7��L#�+Π,.�5k�����hn�]��E���߸����BxF�ItPp�n"~3�b`A2�м��@wx8����٧�C�q�0YA���	��.,�+�ʚ�@��w�,�G9�g�_�T.�����\p�I=�gg��"�#�1BZub,�e�n!�ט/���c~dP�n��Zf���⥷�Id_��y1��R���/AUҢ�[��	%�&��kr�{\���AS@�J�4���v�]���SR,�$�y���h�����g�2��$���q�i�b���+���@ g��Ob�<�7R��i�1��¿���	�c�j<q�A|1��3�[��	�<*� 
s/�mj�u�|8�P����T-��%p9�J�f�������>k�$�X�zIޙ��|���6�e��b]�wiپZ�)����s��~y� Q����%��O��}:�� ���\��p��	C"�`����osA���/�х.��o"8�G*l�W���^�����`�QU\���`(�$�,�e��䁞 9��S�:;�ˑ9��<;D�5@�Mp)�0$l�U���.����drX0�]��*���mk�n0�/ڞ���3�T��pN����ɞ��yl����MB��y���Ҭ�zܗ��y��w���h~�֑Q�8���#��Ի�!ܪl���2Y-�|
}���Wk���ʛ��7�h�Q�<�
0C�G_q���mbB S� �E>?���(�T
�LHm�l��!�J�2�o���	�r�k����1!����/��x�-���Y(S��i��q=�y)l;�RԤ�մ-�cz[����=8��.��#����Tw9�{*1XDT�m�'�C_ps������ĝj��M�������"��jh�� �]=��Gi/�����E�gU;�Ǵ̎[\	�F�l,W�N؉���GfO[	�N����[��jolk]��S�!��@5Q������1��LDn�^m񐨝˨��� �m�BaaسG[a/�<����E�ma
���?�bƔ�l����drV��v�k\��rWX�l�\�Y��e{TMt�h�����оW0�����+���CE���B�j���a��N_�����/�Ǟ�4%G��]���.�ӆ��+	 ����d��B�d�x^J�,*:�Kx�U+VYC���R��v����NbޡTàd�-֞�V���3����J�[��, @.�g���B���W��#�SHk�CD�����Q)��0'v;��`�2����$�	7�zUG�� �GK�4Q82ͳQRb:e�H,���x��y9�!2�o�_�M��#zR����\e��K�LP��4q2�52�1���HAS\O��F�sS�/<�'��}�0=+j8��!�),�L�-�Uǉ)���m/���&מ��6��o��;hS�CS�á2B�J�6�;"��ፐ��������*ɋ��1��p~����K��k���,R�h�v��m�|S�Z��UҲ�?�ܱX�Wq���)]�3dH�����,��i:)��/%^����i��>a��@p#���A��{�R�\��M$?�;	5T�	�[�V۠��� ���y�\0Û$��d��4�T��a��U�xyW2m/@���J0rq�����p�XS�����D��|�'�d�	�;��04�-)])���k�h�Bt��hl�)��ܑD����	��R��ٴ^Xj���|�~��;+��b}�r��Ko�,�7�݊��5h��� _�-�A��0���/;����'��� >Ö����b��,�W�&���U3Z^�����8ى!?������ X]�������j ��~l��={�yZ\92pߚ����}��;�3E�BZ~�������V)�.�'2�{�T�=(G��M�g�mǪ�2��/�R��w׷�1��z�.J)Ү#�o��{|1��>�����֞�d��';�csoMu�:!�H|:%~^��y�ͧ�BdK�+H�>?��*>Pd?q ��]��R��&��
���w%�:�	sW��L�������r(z7�l���8j�s �(�k�E+0�x _��	S�)�Hi9�z�}a���ߤ4�[��H?���S��[��W������g�O(�i�1*)�)�:0v�:])�i��e��o$��]k�K�[o����/'���K�?�1[�֤�1�)�hWQˊc�j�ȕ�RG0{w�3�B(y��T�ͫhb�#g<L��s5���=���kv��̓�i���;`������5��WI	��P"�H'	���Y��Q�Kڤ��v�<',@3d�Ht�w�}��t�5�y8k#m(�۴�xq:<EcZf"P��J�γP�޹8š��l}��)�ǩYI�X[�R�n4i�]����QMHY���5���w�DC\�
���e�m��}��I�j�C��vN@H�0bh� ��rNC�4����ޯ�� 3���}y����Q��,�\��̔��'�����~����#�ƌ	ݐ�sF��`�[q<����~j�4H0C�d���$K"]xt���AM�B����[���\��#㥋�豰��-��R��]͏�ENM�Q��K%���n�2��WLw�����K�AV|���%� /Z��I'������@ɥ	;̴���K3�!0n���v��O�%�QÁ~�f.�h�Q�oZi��Ho�jV﷖�at�����Ŏ9��0qY�����/�� �c�M��Ԃ��o��VtqD>-(#?Pˠ#�ּL����B$w�D�A�5�
Jjtl�ʗ�O��V�}s�d�v�E�t���;"=AM�mșKVET5T��־*��I�]��r��Ln�7���;�Z�"����x,H��Tt@g���}��0�n�ȔWD#�BEv���ҿ��5FaA8�0J':2[���{}����H"	�ف��}/+x������jM����6<����{�}-��<W#k�im�E�!2/��|V�³
�yҸ/u��埬��h�\"bj'���5G�]ee���u���ӝ<��<�K���m4/ƺe�Q"g�x_]T&�@̽$``��t�.���,֚f�yc=-��=�E������=��?8���=T��Wm��n/��6R�g��In�C�TJ�K6�u��^�J~�6�������w�a�T�ٚ�%\�/Y���ajI`	BrƫV��r:	ܦ����)�����a&a7D��W<όh�8��������HZ�h ��d�ЖO��M�i�~��A��C�&.p�vu�Z��%(}Q�9s,60���sI��c�%��6m�N�E�d�K�:�������Y�U�;a�k�iS�-�q͠���!��3EW�&$�w�hnA�9&*���1�1j#8{*3Y�`�A-����	t�ӲGEc�e} V:m�n�*����Xc�z��7�]p���A��v�e��HZ�*�O�7kv^u&)Nh63��\�]���|zG��a��C�����N���I����{�[�w�tY
Jt��E�S؟�p��nŻ����.�j8���I���A����Xъ>�I�����2����T7��������5��'l��h�kS��)Rx��&�	����
Ͱ��G{��6&/M'qh26.�DC��#W�����'�����^
�6�F�������	KXr�ł
�^���&q��Ȉ�X�З�Bc�#0�J�h���()�CwIxC����2e����I9U��l6>L�Q�ZЛ{�ʓN���b�i�^�"�/͡�،���6f�U��'n�Ii������
�����dr$�4�����m�Rf����v�l��9�l9����+�Y]�������@}�{ܟ�P"������zS������٤=A����Bv)�%`�)���@36:�t�O-��MiU�9��M������Q[2�c`F$|���VO�,�JI��Yi�M�[e���@�ậ-HbQc&�0c���Ct�=�����s�'s���������نʔ�[�Cw��,��D������Is��~���d�Jur�,�#UP��өLǥ�G�j���d4A�6���	B{B�h�p�C{k���������$T��@�_���{īDɸ 0�y����|pE.��j����a(��_ȯ�Fܵ��9N3L�I{t�4�ӕ@����/����X�-�I�����4��t�8O�F?��m�JW+��-�XQڵ�Uc�EP���VSo����'l�:~����U׭�)������B�7�vmK��{�uXP,���	z{r�t�������R���tb�h"���;a0M��_�~�� E��������&�ct��=��*�lڄ�!mK��o��8�w�0��+j�@���i��J�ߘ �Ȭ
ހ6Hi��X�#&��iB��80����h�/ʏ:�S�H�<\d@�C��y7R#�[K74iLu*Cux2KB���y�N�˕Jj;��t��H4�����:�<�	��_�6���lu�c��G�t�G
��ыe�*#`|S�,�r����%��������Ŗ�\ύ$ο�J�|��T�b�=jM�����^�p��Ë��s�ٴ�D.4���9����CQ���@	�|��fzG�7Zk���t��Sߖ��]e:�ɮ~��P��gQ�\���:m��K0�,R�n�E@S�5�&ډ	��V}#pD��>��ieo�n�1��J�{&��bI<�����~lc�:�q�Y�7��^�R��5Ζ��p�5cEJ�fi�+��f �6�Ʊ.��F�Z�}�C�|��.��!nO9�5��2�頤��p	��꼬$a83��s���7�^I�4{r:��M=�ē�nQ��.���}1X�+�W���B��Q�8�N���0�4�u^�{�~�H�N��o����
��j�۟�N��Y�]ô^��n`���O��!V�������"��j�g}s-ה���ʲ�PD�&���H���~M�fv'�Ƿɰj�*���r@�R�~+e@��;T��V���y`A#/@��gc�O�d��'~�x7򜇔�$z�^����f�GLy�x�|���}W�#QU]��vȑ��#�R2��M�W�?Ԣf���aF,��m�G����ׯ�O����<Ū�|Z<��ca�/ܳ��&��a�Y�o�o��� -`�N����Q��b߰�ᬅ�r��ip��d�e�Y�{��.FϵUa���Т�c�{з�=� ���R��������!������,i�ӹ�>��㠼�vMԎ�+T��ꇘ��ʌ}��9#,�=7��,	� ��!����L�hN3W?a��ԗ�o�.d�rJw)�d���R`��:�sw 8��d�����BȎ\7��E��LFE�8&^��g��]�~�����l�ɂ�.N�)����Z�+ƍ�� _�����d)-�^��B��mo`_�n���]��<�0��:�ސ�a�l�	�!>���hg��@y1��'k��M��M���(i��Z_�;���@%BFV�X�x�{Ǔ��@9o�ɮƉLP�>W)dW)���G����L�HB�p��5Hί��x'C�k}l��L���g8m�3�����(��܄ݬ����T%c�gc��rPW�A�Rr��+�j��@�p�c��S�T��i�rwI��W!
Q;}ȶc�.������)��6�=gX3���W�b���f�D�
��I����c����NN���k9U�^v)��u;|O���*�|�յ�8�װ��1���MT0>��o�뽓��e��yV@,;S�f;����.�)�n�w��@.	r��e7�{�K)+S�k�F�u�6�n�ܘ*�vǵ��Bz����í�Q��ⳁ}&�!�!K�ϟ���C�g��3xK*SH��ON&Y'�v��z߂�I7�2�y\��Q���7,��}	��n�����Jmjfx(�O��SJ�����WJџ3����q���3�j�ϳlM�A�=���@Xq*xX��3]�X�C�x��������w��
?��<��x�+�iȍM�{B�����Хw�R�ƌ��h�4d<��9@�.��9���c��V����0ꦍac'��X��\�b;�H�ٌ�����6�4mC�0�pMI4ry��x旤עe3��Q�ui�Q�X���)�r�x�`��cQ�=
�P$����q!�^�m����,�*�x:G<h���`ܐ`����������@̼A|�<7Y�j��@�\]���� r��E���@�4��"`iKp�E��(Xp$�����8�>������&��2hZ�y!�(tE��ai��)�>�t�)iY��_=0����6��R`)MNG��5��{d}�DōkY�Q6e�JO�T
���$��5dhE�N?6g��6q���A$R�8�~IKөI�L��q7w<6i�-Q���(?B�/,ۂy�UTp�h,u�V5���p��7�1��3_Ť]�[����Yиl����i�"�]���8^+��g����!|fԬb��p%�w�V�u�B?H��t!�����jh�㋜��BsĠqxp��Ft�j�L�fkd]�k&g���RZZ��A\>���_̰�s�凵������
���F���r�!������R��[����L����߽M��	e�ʭ'������ٰEF��zb�/q��3o
<Ilc�]Q�S� Xh6��:�dg1���1��@r=۩���C����e��N"O��\��aguF�N�<cf<YV:k�/���?��˄�v\���Z��jYP�B'�-#x�OG��W||��B�Z���	���75���^٧�	Ļ�@ʺ��yf;��u_>3�=֮���la�<�U����0`��~�� )�I�w��5���{-���D�]!5-�H�qi�]?�� /��,H��1�p!CS�=J�<�퍒�E��� ��^�4���4-�)|���������(�D��y��N�pLg�I$���h�sӘ��\ �20W_�kt̽���T��?NA�ލY'T��T*�8!�-Т�X�Z��z��(�c�	'@�`�Џ��i�"�S=� ���O��g.x��J;�lEb'�f��H�K�rT�Q;��+�[7jsƏ�{ـ��/�j�P<��S�OA�/iѠ��ު��>�N���z�-0v�Ŗ�T8�MR@]�g0�S�l�5W����5�oZ9.�I�7�PT �@��u�b �=��|#�Z(a:��q	,�۾�=+8���S/#<�wO���� ^�Y� ����Mg������
ū|�ɓ�\�V��E'�P�4�u�l�<�7ti��/vd�;`��x�*�qNW�>?
�\�m2YP��LF���a�J�xP�R_F�P��>���~�F����6/(\�/\�Ϯ���P*8�5�x����ϸ�VF�sӱuZ(e�^0�=��r -�qX�g3,��K�y���Rqs���"�v��Ooxj�*ǀʒ�U{�}��ć�$�����zF'7�,8��*F�bP�&�ԠJT�j�ƍ4��s*�պ�*h~<��Y���!#��椞��e]f�z����.�%u���4�mL���س���݌��?�g��n���-������V�R����y��7�Q���~�<s� .̅Ɔ�������n� ��XX�(孔��$�q?�L;���D	U|m�F�7��N��f����J헑�뀱e�
�ױ��?8�Fz�a���z���Dg��i�^�f���0�"57�]�+4�OM����	t��4me���ߓ�yP"*��^l��)�OIF�1��M!4���v@W�^�t��ed��ńCM���m���w�@0F���!��6����E�F�rE���&M2���Đ9���C�!,�!F�ä�+��4 �W���~Xا�4Q::KZ�������J��? оI5=���X�B*$���.E��a�
�r�n�ۨ�fI���љ�9��`3��ӂ��i"˺[��X��g
�NG�U��%�sϒ�t~'H:�RT�D,���A�Hl����0���|��Ւ���T�#�F�����)�f��uS[@'x�d@~��	
�._>�qƮI	��9�-��i��9=Z�r��k���s�	fZ��J�|���g9�������8�>�\����hp���͓�'������ļm�1�B-{�$^���XP	�FvD�Yʂ�
�!�/�A���#�??�ID��(O����!���#��zȅb�?���9��06[u��a8�S���ƧR��.�;Q�E���U�m;cb�� 3���`yP-6�U<=�N��SXZe4�K���}`z�$�"V^��>������Rv>�@$Ȫ
U�j�e�A<x��]Y"����t�l�&�Ї1(N��y�I3=kz�Щ��F�'����#�"����z���n®� pj�]{��S���@�k:��m��5�l~�~�RyIEi��ht�[�p���u�,a��'��#x6�ݐ�4C+�	u�ڥ&�(��,` �h���G�N��� ���q�\��@A�����ו��l�!�&\���"J!)Ƥv�(T }�4�:4X��nm���;��Sw�hd}4/�C�	i9e�;���2E]�Δ�l�P������ո.��**a̎ ��^H	��f7�jDr�R0��@��v������߆��3Hl�+}q~M<}Zm�=B����;��N6���a���s�v�����(l�R����%0��5u�1�[|��ʹ��ueMB�ǯ�����1fK�`˅[T`b�:0����qJW�<$#^���`��� �_c�p���0�ϛ�IL�"����w�I��*B<�]	�\��N:+/
M����C�	�.Ι]5��/g���7a�I+��v�]����A��US	����䥮��H���������G7����B|鑼�2^���\�ڄ�C�j�B�s�?�Y�N���{����Gxn��`��ݥ���H(� �Į�7u�"/�������bdM/*Bp?
v�I����.oW��=F�*t���F�|�HV��2o������d�bf<��B�!;�L:���yP#��Q�bW��`r��:���^͒0�E���.�|�N3ٻa�T�Z��Q|g��&�[!�ݱ�;��Qk��h#1v�O�ƌ��!�E�uʅ����A3��w a.�(�$�r��ª��ZoWnB�[J�r���4�QzͶ�X���8�����ڰx�`�#��U�.��Q�\ބ�Q����**+�0
�H�V��@+�z��M$Fޟ3zK�>}V����6�@�������'�����e�@7�-�"GM?�z���Kp�.*\r"�(��Ȇ��sO��h�Ӱ�;�!& *`�S�l70�{�xA�ݎTGɥC�&�,����?�T�s�7b���|���p��cΔY�����r�K�18~x�L���oJ�|~y���c �ϷJ�>*��1���"��?��OyO�9����?�����c��f][!NU�!���DV�E[ �#L����©#��ړ�f=kQ��8u��,�%�E���V�{�VNܧ:ϣX�z�𤸽�����V�֕,�=D׬d�]$m�3���w�رK�����yFy��m�P�T��Y���K�4.M����������5&Dl�$���)U��,�?�j�I�{W�J`Y�t��Y���x����E�AJt��Z�����!e�w�Y���xh�7[������a
����kj�����/g��54�m�/Ւ8�z�㇡��|�����N��nF[(��t���2�4E�M��(���:	n!_+q#E��-�o�w�-%4�$œQD$v&2�א�z )�;+1�7�g�=u���k
�%��T�n�Ԫ�iT#�Ͱ*���$��_�!o�k�`6��@������2�ޡ�2��(��9�21�+g+�g�>"x`��KrQ��Bi,�<#�w
���ڼ
�V�˾�ޢ"�Z�ʁ�{{����~B�d�[������^)�F�L���o���T1��;���M6��\��t�>C:����K��{j�ͩg3�5��,,�DZ��6Nuo9��@8���;����N\�`�~�Qp�L���١qF�͆���5����)���� ,�*�ۉ�P1d	��]�D݀^���(Q<a�^��'��J�Zui?�AdO�"���H��������?rpM	=����?iZ��/��ư�9���s�����b*޸��-zI����XBg��uu�)�I�7Czr�i�kd��}}����\����W��M�jeQD�O��#z�vԝ_�{��Fۅ<���
�b�2)/#�a��u�C@�����.�Q��4�V�d啕�&�@���U�"�S&���_���9l_b�#�[�F=�_tR���j�ZA��%�{CY�7����Ҁ]1C���79�� �`>8��0>^���ڰ�����e�e���3�T~ܛ'��O��w��G��$���ߒ�y_A��
�� ��W�s����MT��QT�f`%]�p��m9��y�p��� $���}���f�q�6��
�J�h��"T�+fX�IƗSn�үI0$� {�KMhq�n��y�A��_dC��҂���gE�8�j�X���{�%p�qEVi�0�Ƣ+���Lq�x����Q�3�	�x-#Pг^�t�ZG�2�5��hx���Z&'Lk�:�J���%��5H�'��;���nn;ҽ�<H�|��# Y����}�1R\��&Di��Ep�A�{w}��ίIT�AS�R��Ç�IBv�_��p(�US��"zg
xL��������s��Ќ}�}��Pf ��;�`8�Y��Ah����0dCĶ�P2�t%;�_���zRJ�F|����
;M ��V8�	̍�(`d��w��J�j�_S*��t��*�I�-2#�n�H�υD���؝�[�h� p~X['^"�Ւ��H�!��BYGސ�=a-{�@�HMN��n�'�2�h�������4��J��~���/����2�JO�g�3��w���=�S�z�*����;e��Qn���f�to�h{B�������a.���3W>��W}�f���(ei��M�+�y&϶�G?�U��ۏe�M	�KѸq�
et{e��[�"��B������_W��5���LbT=��-O\㍽;��>�H���T���R�bb�mbH���p�q��ph:HX�3�wԱCi�*������(���,ܘW� �̓��\nmS��@�#�F育�lY��9c�7Mw煁��ygl� �|ˊ�6"p���(u��k텓�m�^��o�Y�VUW#������Sk� ��٣T���-��������q42���_�&( ^���+�/�|�kX�sJ)#V��t����]���3���WK1!�|.h���Z�f9ul����H��*n!�J�ѥ������u��LR�Sy���|��PY�9���LZ�{dd4� Asҟ�̿diq�X?y�!]a�U��ܩ0��|y�Kh�Jƶַ*���@!�}�`�����}�V;z����<��heSU�%���F���B<�;2�N�C=fry�N���Ŕ6:��E�S��Q*�B�tڪώL�S��x�����мo�A�{�l	H��Ϛ�~#N �j���}�ǣZ��y级�����,@�.�ǎ�6��o��/0ӗv2)֨����5Jg�S�Y��f
�ni����C�X^���o��>��G�"ics[\��/�{fʣ��L���7�Wt�]]�x��,nCC�Y�۩#!pxd���m��V��ez�
�
��8��*�5�E�k-����z�3 ��ށM���ѻ��\����5I5��&&��=���RS��O鹥�[������;?��J���-�T��jz�D�=U��5|���������J=͸�^�(��0��%�'�0���FC��Y�h+e�����cT-�3�"�d���d\k��#n�+bȋzB3c�6�� n�EY����>p����l�{b���'����kHc�3bA������t�f�B����W�_���Tn̸��'��c���p�K�Fs�����#����Ux�b�Eܿ
	͚~>���^B��K��/�8]�o&C��ozp�6i
�3����`(F��s�(�=ܮ?R�j�i�<'N�Rl�N���n���R��qq>�����|����R�v��~�:��{���3��X�ґ�/��v���������2m`�/80'#l��W�4$�Y�K1b���M��Ԗd�Jr��`A��KX^��8%FC� ^~�C���bz��9�*��Ï���4��SuDY�+g��c�����i>���9�t@*5��f�O�[����iidv��#����s��e!U��yN6�q��E��i"���9,V5���U{�6�?��c��vI��C����R#6A�Q.�2pV�����\�S����sٽ�fM���[��+��!9��oZ��A�#F�p��Nǌ�}�ie�$��f�sz�}gBC{�3�d��K��\� ��uoa1*�ʑ���;`�5�x&�F/���9h��"���wC�f�C�?���`���ΒKߚmqN������U���Q�iQ��U7N���
Nz�n��a�H"� ���K>�����������*H#���q����D��֎C�w�O�{�����^'<|D�)ͯ\hJk�&� *��>���d��z�Y�kQmo�G�c;�v��[�UR��ݵ��|�v"d0���`������b�K!�v'��f�i�UE"�?�n�P�>����zGOo�lNr���{�}�����E�L�Cm`շφ\s�*�|��Űֆ$��\���;�b�.����O�����;����?#�w�:vA�kV`��ჿ��u���G�|u`�s�̌8T�g��Ȉ#���@'�K_�f`�k��1K$u���w���(��U�F�w�6F��h��x�'{�(NUl�����N<(w�\��{A�$pǖ��Cr��V����u���)j����2��O��-Nk����덟�yfp\5���+��C�y�&���8�^Tٹ�ldw&e��y�D���*qp���z�4�"��E�i�eA���m$���1���G:W6�,��|�o�p�a�+�
����Zb�\AV�Չ<w%̘���)�A⏹y�^3��#l6e6 �3�~u�~�x��_��n���W���� ����xډW�
� ��Gq�7���bc]X;�L�ߎ�r�p�_F�4����E���C�!̳�U���usRDOIB.��V�2���T�w��}sh.S`�mo%��pT缎>��ʩ�|��	'�o%���'�k&A�O{i�4Ag�`��C�~�悅���p�b���n�Tv*K��fm�#���O�a�iE�p��tCnGQ��������$*;X�%x�S�J9�%��Oܱ�ˆHP�����Q2u��"���)���;ADV�xx)Ar���í��:F�O���a��͜!w^�p���z��DN��.�/�N��@dI~B[M���.�l����@GuI�N,`�RN�d�g�|)�V8ЗaJ�e�� 9�5+�AlS����q>����b�0FY��V+���j���g��������|�y�G�f�e���+(��wAF��M�;C�BÓ�+\b�{��|������#��]�4�@.��7G�/��V���;8K��{��K�!qR�(/Y����{л���n�؝�v����^���h@v��H/��.��3�f@ �QW�d� ���&;�(]� �|m?h�<9����$ Å�2��A�g���-��@`�U�ܓ��,��~�lq��]���8EM�ʂ1c �/2�6�:e�!W��lPx`>8Va�\&�!�i[��9�&ߢ���h�.���Cwk᷒���)��~�V�P\p\��W	p${�}��`m=���*��t����H�A� ����Ξ��kK��)Ƅ��(Z4�9"
�˿i{�(c�ØsL�̠��y
?��k)��v�,�Cy5D��IªOW�Ͱ�,^���Ew͹WI�_Z"�V�/h�$*�`�<���嬂V��W��U�Bm/K��,m�V��P����b��?����O�iT/�9��'Yb0��,8- �
l`vg�)��TUf
P%{��3��,����o�k ;^&(N�\��{?%���eu�P��^+�m���Uejj{�b(wKvw��O���?���	������ڛY!?��x��T�}8�g<c��GaK4 �S-��[I�&���_�w/��2t�́�-�q�+���ڙ)�^���j�A���%G����"$�^m���-٫K
N\[��.hkO��A����ܵ�
{��P�GZ��Y�,���Z�(�,<%Na�e�X�3�,,�L}�a�0����H�`�~l]�oQ�k�m�&�k�ٖ�9,�j*�(uG�zC@�[a�b'��
�:F� jk�w����'���_ʠ�o�K>M{j-���7݂�'*dX���$��GAdʰ�5������U~"�h�׆���3m�\�5��F�?|�6�b���L����}�v��@%Wy[:�*��P�&����n(	�/�$�ɿ9�E��BQ�;v�Xv�g�0�F,ߦT |=�����wtP�8jS[�LCY�#�=��������h���cƱ�b_��>��Qw�{�nd�7Y7
4��.AZ�16�Qc��5y��X%7��k(�w1Нu�P��`,w�i-r�?݀L��W�D8�p73��^��uS�tRJ;.��S]_J J�짱���oq^�_�"�͆hzc0(N���>#��K9�̤��?e��iɕ����e�b��wɖEgu���xF%Dڌ���o��vx������ඝ\����� ���R��޲�jC<�ُл4����j��F�T���bJr�3��ܑ�u;��Tۀ�	�A�����
��~�� F��G�o�Z8���CJ�.���%6�.-n(OM!�I���3���o�U�QJH��, j}�F1��M�H��{� qCpu��n�->��-I�� J��gI%k}J!��%`Zt�'f�%i��H� ��0P�Մ���~�8����-I���9B?ӉX�ny6�ۄ��{�p?,�g���# �|
��e= ���ZKL3��jט$���+�DaQk ���3��4=���L;7��iN�`�_� d�e%�=�R+�����/G�$t�҈�2�ڑms�~�o�1W%zt:��Z����C�djN=K�j3�OD�8��Lm;b]����}ϩ_��rq��w�p�C0�0ͻu�j���ިi�[�g"�%��B��K{���P��K�}��r7J�]r�~�L���]�E�>��ZYw�U��l�r��*�J�w�V�gJ�f��̂xQ-�Į,�/�+!f*@�.U�k��+y6���-�#�ȑǙ`J�(����tn�`�=b���l�H�@��ý��Q��^��D��U�j}��rI�޸�:�8aT��o!+3�9jM]�tx�.�'�$)���^���hC	�����ӑ���ϒ8C�1}����8�)���
#��?KT��|��Р��&�@�����Z�e���X��;���Q>�,*�u�SEg������̞������e^�J�9z_�pvh"�ᒾ���!�+���B��1��`o���ڶz
�f�n�JiP-�1)I,w��6Cy��ʚUh��[α^Lyg����[��9=���hi���msV���Z] ���v�7(�m�Թ!�T�����+�(��w�zk3����ucJ���ҳ����y�"��>�SJ�Z�:���c�S�a�~�G(�	��뵏pͬޭW�T�Ή�V	�o��Ȃ��?@�������b�WR$"�t�C��|��|�V�Ӝ�c�o�e�'x�.Q��@_�Q<�,�Qj	�2��!�nw�Τ��Q�X22t��R
�ګ�ؾb���BaBD�t��0Y��%h���T��+����h�a�3&��-ZNCs��Um���Ǵ
őn@���=�`Wr�E��ܐ<.q�U��R��e3�E�νŃ�C:Gׂ�Tu�k���*�N!3���]^BԪyM�LX��l�����(E�;C"$�)A�ɶ{J�N ɦ�>�c��F�(C�^��5��Z��M��,Q�8�t���w:D�#<Q�0���<��~â�9 ��z���q.-0}���w3pz@i=���x�?,�YIU� ��AJ��0��7�q���+D>b�����@�,6~I�Թ>���[��0 �:ai$|��w�`7K��ղE~h��4�l�Z T'o��lͶ���{�~?j�[KQT@��!�䭂���^�����@�d1�܁4������-��i���j0	��ZӞp΄�ص��	�?��,��W^ќ��l�=�ީ;on�iE��'7x���m��$������p���n�t��P�0�؀;��'��+�{)��:��=�؉�3�0A��sk� )'����iqQ��ķ!~�<r�^1_s�)��͍@�J�I^�$��	�M���vnL	�W�V�w{�M�)��__3��-��Y�Z�>�,Po�T�)�__���	n�0��jzI��/�JG�~!�����Ca�g��>^���d�;7E����ej�� 1K��P�:H�s���/\:�ո���e�� ��>�+�\��C�:6e�-NuQN7��o'P��0����<��>�8/Ӹ����������8Fd5VR6��9��^۔>N�E�;�ѡaR<�L~�L���lC��^��;�3ϡ�3�	�� �[�[n���l�֛k��a �)�f����e���W	��Xq�<^�}~�>'*i�޳Yο���$�K�d:W�W6|^q��Ih��A4�����l��Љ�輿e�o(�J�!��4�f���i���A~�0��*kV�ł������CA���BW1L��2m�BNHG}���)��8���e�8��}���[8+��m��}(�ʂ�^���_t��@z��&*�Ջ�$�,e�2k�O��+ss4`1�4ƸFt�&�ZGb���]t P���X��|�6M��?�FMh��� ��	\�}��59���_t�,k������������¡|A�,yj�#ص|�1���p]�˺��H�א�;���o��~�v��~I�-mk���M_Ϥ��9{v�cN1 dݷ���ݧ��ijm���b`4V�U��+��#� ������b\�H�׎skc>Ժl1�p��������mf(X���a��S��_y�ʩ(��^���I0�F7�AZ�ز[�W�(��V��k������PWB�A=��ya8�|��W�Q���@JHq�F]<�L���9�"m���k���Ş����B N]|2�Kp� �hJ�d�'������s�&��m�
����"{�� �ل8�i��o�D�/�+�L��@��;F;qI����$h`ΰ�XP����A��K��������7��"Jҏ5�?�&���3n]�'�w����/���c�֒k�Q9�L��B��8E��1U�����a"�:s�a��8o��]6�>��0l��4�8�.r�/*���Ra�`Zsa��Ջ_�0�H����ȗ�OD
�%j�6������ljM�}�	�3���t�k>χg�DE\�Jy	������P=@VI���T�Ad��x<�G�@B+C��~ �wN�Q ���5����l��|%�g>����ϾL��UJ�=�h$i|�+��7��u�ϻ
+/�KB	T���]�c`)nEY���q[���pԵ��'=Jw/b�x�/:ڠQ�o\��w��'�dg�ե��\�1M�n*I�/�6�b���a:"�TjbW%j(+��&{�hY*d[��R
H��<���hMmF�v6ص<a�gr��R�Uk�����\HC6f˟�M���E�B#�C���yH��LN9�f�H�tV#��c����YA�8��C����M�#񽄑�~��X&�R'-H��l������}c'V����D4���4"�02�Wi��-^�5ѵf�4���sk�w�:��q�N
jHޛר<��G�((H\�%�o�	z��҅>C�CM�`�+\ГUz-B�.ٞ���;�U�y�U;F��ʳ���8d��]��6�3�A��e4H�](ya0�$��!�l��g�j�uH�Ē�i��X
�ҰO:�b_I��oC�Fq�I�qf�L|U������B��mQ���$3���"���?Î�fܣ{�{4����/�4�W?`Z�/FnP�ԅ<��L+�j܍so3՗Ꭲ� � �Κ�����fm�*8@����+������Ѽ9��8��B���8��m���-��GrUs�BA�	Y)�j� {PvT8���b��%L���WZ��ƾ�0S�7��@9������80B����gK�ո��Ё��v%�xmދ�!2�� sۊK�v ������1A}�3	�peǐ��VaV&<�͢}	fK�^���M��
@�Ej_�@����]�Uʨ�9�c��0�@��}�� �[ZXn�
�5d��l�]��+���Q"�9g(ly|���q�q^��	�����߳�]������@�
JF���bCpN59�~~��$`}��2-b$�'p���d�v��� D�V�>��\��*XH�l���ll~R-��"���Z�Q�m�؇��M�&*�*u���+�cU?_#��!��^�]\�ʔ�#�_�W��m����^�m�����5J��1Bo��`g����O�L֨�s<gT5����WZ|
��%r̅��=���3��YR�\l6���Bx�W!�s���%�jh�}�it\ޞ�}6R�DhqN��"&}��q�����eQ���Ǖ�Q9x��tP�T/rWD#���?~��y�-����75�]��(^�8�e%$	;~����}�C�TxNv�-�&��A:9�:��.%6���n���PF��ɿ�.C��T����2@�ү^�V���ǜ����[�������Ů�=���0�i	�?������t57����e�����i��{2��������cF���%��f�[��)4�`do�a� ��M,TM�����i8�'��h�Q&�(?N��dZSC�7�6��َ.R�]{�=����a���i�v.�~���E�X����N�%���Y������w���9�i��&�L�����ث����O=�����6$�!-��ȼ-8:�|�$��M��7i�Q�OM�r�',��������SX`��C�A��
'_������*Ah��̂�<���9t��v������L��uv�!"�o�@$�U8~Jt��<j�Z�W\�a�vE�P@�a��\D῵�+7A�[Qxv��n�*<��$�Kߋ�O��Ojc�#2�m�NB�배Y�a��.��ɖ��Ӟ��Au��H�T�ϰ	o.>4e_ �c8����&Qz���
�絓�>Yz!.�ω��bS粃	�y�Ms��|�j�)wH^��6@1�`�PM�?�Ʈ	γ�&J�0� �YS]������fI)���χ��E7Q��>�;O�g��|��7K��%ې�HVV�<��j�
&��V74��s�Y��0GJ�EH��~���/7�sj����W���_(�inH��Bo�d�ޞ����nm�A�' �l��E"���<5��L~8�cUJc�΄Ѝ��D�e߆�5~�� ���ڌ�pHLo N�O�p�tYR�{=�Ԅ�����:���9 ��{,��wH�/}
k�z<;���V⥡�<��Gfs��n���WՀۄ�l^X^w�}��hDw_������H��G��&��d$Jn�o�� =V��C'75��<)�,���䑑C�PE�wK���+�-�&���~a�\��B+]5{�ԫ�-�0<��a���T �&*Z>Ǩ��-[p��:�a)y��q�&�����?�(�@&j��٪Ko$���G�`��[~�f�¤\u��!��XQ����"j�C�&O=\rݿD��K� iB�H8Zd���Mn1�O�>E)4�@�_Yf�X��v�Yq������)�,)]Pv�C�K��n'ũ�ׄ�H�vH�W"{/<��@����yZ���̜�k=��j��Q�pe_ Oo�llp�.B��
&Í� ��K��N$L�����s�ki�������{qg��C�k7�����0ߖE�<wb�:L�f-1����Ɩ�	��Z���/��Kj�_�	X!�ɀDp��S�j�z��}�ƴ��b��<��/I�]E-��s��+��6���C��8`������Sc�g�?��s�.�a&���?^s��)���(hN����o��e8���{SB_�]�T֟/Ҩ�&�6��p�~INύ>{ &�y9�5�k�G�u���#�`;�
�+4�-6ӍB'!��m O���x,A�3�P>�@}��w��y>]�t���/�  @�8�
ˀ��O�ZL�m�[X�p�Uhl,� kD��E��B��P���{ ������D[�`f�⚻��J�H���/�Z���'��P�5u;����@n@�AV�8'ۢ�oˠ�X@�^��bl��&6agڇ��g�����9�݅|
Z^�:��|�U�-��b�r�|��*�{�췇�&*�Xuè��썉�A�Z�큣VPTRO��=<�U��\<$���l����Z�l\/vTT�u� u5i�)�x�ZŸ�;�r���5zf)��U�{dW�mQ��@7o���u-���Gw[m|gZ�m����"*{>���'�4�zx+��8�F�j�x�(���$��+��]fo!.^�=P�G�OBcB�]b�^���$�W�(٥��,<`�L$9(��u#�:��*������S�)1c��Z������h�''�g��D�W����|z��:�K�a�"�̶h&QJ
k�b�=R�i�(�y�]" $�}�ͳ�7�]i�p�fӯ�&[���Eك����{��{�H]1�e٪��-���®��ê����ܕ7�W�<���Nn s|x:�L�_/I<�N�z�N"��^1�5�!f�x~�g�=AG�S�̏j��񻚅`�vӃ�5����������Z?l��a����H�jʺ%)o��I;~��I�[3t�
�HB�ڗ�|�:wK�
e���$��;��ڣ�Ho� ���[�a΋3֭>#-g���{�_;QLL'��`�*��j�`81�	�y���p��ࡌ\H�Y�t��T��涅��{, ��&�������mR��������bm��M���r���_��@�43�2�:(~��愇�kF�lP���&L�\��0V��v�06��B�v�FN��X�)�|SZAa�$g5���~�b�%Cꐟ��#�ߓ������*gT���[����s��<U�̖�`�x�꿽	����W���i�su��IN��(<:l�3�F`��'oN��lF�ʮ��y���#D�t5ݓC����E�`��F�-��!�21,/���IV�g��+0���(�r��x�W�	������!��_�G�i��^���̻߫g6�܅oPa��|�;��)���a�e,�K
��z"ywkJ���N�&q$�.����"��^�3��u�D�k���9�Cp��	�i�Q�)�� ���!��BR��,a����^�� �@�@�0��1����ʌ�9�>�S�ռ�O�OB�����S 	�������M��w���Ma�-�G��ZŬ*�6HR1���?XCU�;��U���������y(g�Whe���7�.+-��g���z�@�^���p���@!�e cGU������E�Ʃ��XKe���k-x��B�ˤ�r�������F6�>��W�������7&@���������Ɓ¶�:�n.6�y��cŉ��X�3��$v5%2X��(�-]x9O?��B��;k�d8E�{�p�Z�A �y��3����V����b
H�BAћw�����k���ς��(�m3�* ��,�(M�t���2Ҭ�xS��=���[%?���P,S�w���a��X�G�ܵ��LjX�6���@��J�a�F$m���I��u�
}:�5���Y��C�Cb[�����r!�t�㘆��L}�牭��`�Ҵ�n w(���3����� <9@@;4��B2�-��';�,˹��(bP�-'QK�4x�G*�"G���
�M������D)�Y� �6��F�d���m���|��;F+�[e�g��:�e�,6ȰZ��w�����pHD�z��}�xr�je|�G�-,w	{�}5��B4���< f����,�)7z ���&Эm��}.Γ�M�>�<�̧@DP�?�s3:��ѹ�� ���X�~�W'���r7��T��٘a�7Ҡ_l0� s<M6#wjX���1�=�!�mo��)�'��R*�U�Y�U�|:���0�e�bP:Ai���+^���BC�\��[Մ��ҳ�ՍV��N��)�U��eA9#�Z�sd�q��0mN�l�a(ʛ�_���w�]�-o�Xy��T }�	���9I�J;2x�'��=����4��!�L�Z����|T2���<;�:1��1^qO��Su�[G`�Q
���p�L�83{��<[o�0E���c�T�(�y%bA`:򳶷�l��to�WK�
�/�8���l�텕IՅ��3U`�j״^���𗔊ν5_ʄ��q���?[yٳ7�����/~	6_��A�e������٪Ӌ���buk��ĤpG��F�1�bW(vǏ��)f)7Sj|�Ba;�}N�ݽ�&K��]��|�E������c�: �gx�3��.�}\���'��3=T\�cT9�%a˜f�6k;3��2I�W� Y�U��'�d7�1�	���=��������[�ʯvH9���t�s+r��yg��T��9���ş�������28�l�h�e?��s�9I�W�f�h�wLo�=�W�r0³H;�����l�qx>z�?�~*hԩ��4X�Ǘ$��hre��<`��9����]�3�7_(����L0��i�'Ym"��@Yn�Ⱦ%�����9�Ϛ�.f�9���A�1Z�Ni�M
m��|s��>zi=�\ⱼ����6\�XK��j��FpvX}�g�!a����.��H!�[\�fg�?���f����	�}�����nk�q���/�{jFp�
�����qLq�7��ۅ+;yvou�}����CT.��f�i[���Kԝ���J��q�Y��}��dxG(��%ח�>V�}�53�ᣠ993���,�3Ji*�uw �b�Ư��{<��J�'��-��G��� �P7t��G��IL�Xj���Z�o�^i�u��+ot�(,.P-z�1�#/�
�V����z8l�V��ݐ�� W���,_��pM�q�p��<i�*��G�=*��^ۧ#�<`�L}Z�tftz���u��<5�+`y��m��w���x$b(�Ŏ��@�¦Eχ��� fR��?�hj*`�gأu���ͅ�t�𝧂�Ny��h��-��W��3�1<GlB�fe˼��E�~���̷�������#4ܯ���h����
���{pTx�1 ���=��-��v_����;*.	���;ڬ��=���D5�|�A"�49'\����\�i���8��!�)�c�j��ςѺ������ж� W�j������T�~�r�� ���+Kӈ�b�^���9]%���'��w������fȢ�[q)l�m�+�hY�����&��U|߅��z�6�Bn��(^�ÅEw(���֖���de*:��1�&����/jg&r�GX�v�!��7Q7����{n����Cg��{��43��?��eB�CD�%����"��{��i��:h]}�_�r\L�F=���~���0U��-�V�+�Ž���L�cx2�w���)�Ǔ:�;ZT�|P�_G�Bݝ��;-E|�����P�bx.��0u,0�I�������y��Y��-$�u:��m�;�AoX>����Ó0�g¥y�?J۞��}E�6&K�`C 4��t �.�tny^���̈U�P�w%lN�Qs���/�	�KŊ�-�����p����9%C|4�B��:P�}t,
U˟�܄�-�]�h�Q�� =	��X8��)��!'����赯/L��Ě�r� E>���f6L]u�iS5�D,�'5S�gTl�$`��9�m
4A��!sbh�ei���)K��X��̃�<d}��������r�4��	����o�l��ѐ���9{��r[\BVen�E�t�#�3Cy��ߺ�2`�Wk�a��c�K���4F���b.�qB`)�"�Ncf1��1�ڮ/g.w:�u�h_��"Jq�Z&4|}�Z)Z�o��'	/�B�jQ3Lӽ:��Mn,���	>t�xX��+]L���ޗ��Dr�^�f3࿢H'٭h[��bμ+�4�)ŬS[	_�J���[�y�4�F*c��l����q�p"���о�榨z]�Z�:�@��'�����0�xH���D����G����
~'��K�>vN����c�����|�d�T��
���������V��V�(��hkx�����mZ��8�Ǎ�[Ͷi� �C�A��dҨ���/SN/���wv��Xmn�����4����jꌥ�6��K�������<����7P(��m���Sa�6� }amHLG#>7�UR��{E����~Ÿt�o�D�'�[B�ٖa@ȡ%���)ov)ȇ���@g=�8��Cl�N�/��)������P��/��f`�>(�����WN6�W�!"g�i���$���qA��Ʃ����AFTi�3�<��S>L�B�L��q7�!��~a���%�ε�7�}T��i�>�_~v�3t5E�X�
�_`��O��Ֆr%5\pJ�P{ �8awUvE�Vm��D	�YɪP��T:_ݽ��/"��rQ(�Rl{�-W��Oo�P�~N_g��?���$��)��=F�2	�=��D��g���X,m(t<CX<��K�\|"�^*O�#�� �h�xY8ΐ7�H�A���&�294<�u��l�� ��Lk����>B�˨*H�+�/�ehu\�H<%	/Ų@+����&T��Ɣ����F �j*b�Ȝ�	<��6˂F�?���Ch�Of<H<T����5{wE<&GX���uzwu��V�k$�☔,@l$m���D�kr�̻���n=�?%��_/ܡ~�
���i�`�O3G�&�4ۙ}���+%�n!U 5��A�����:I��ڹVJ�.�K+U�};;oF��f���|,��_�۾�$��s��vŝ�>��3�]e��.���b��i�R~KH�V[8�
�m.Ȏ���tع���"�0ث�4���q/^�ϔ/��]��;{�3��-�����U.���M���J�����X���9�4���!)�X���(��֭m]�kqYWx�=7[�M�����Jd��7�#\�t7(Yy�-�ʱ���u\!���I���Ok�W<���� 6�w<*�N��i!qt;�G�i^����� )�*a�r�qH���tE��X��/m�r��sC�����d�ʫ�j-�;IR��T���}��]�{m��,���������y0is�x�������R��W�"'�����qG�/l'bY�����H��8�Ni̠�G���7>��
��Z8o7嶅�)q�ۍw�`�ç�.��U�vtz)��'9g,(�v'#�W�7�����r/���b$��+aɜ�j^�x�(�
<_hJ��rػ?^ǌX�X�w�yR��2%�C���ɀ<���� >�N���%ģ��Y`���yW*�.Bì��؈!V��l�A(X�sm�����BT�&	����-�n��h�l��r���ʛCp�;�;��S��t��G}�w��h	e
�R�!wK�#�(h�Ɏ�6Fky�,��s)��?�'�e�$@t�VK���B���ې�A$2攒��I�"/B,�����6���mz��ԏg�O���Dd��+s���@9�45JOC��a�-��$o0���/R�Q��I���m��Q��/��Z�^��lx��>�7^�|�%>�],����?s�����C����"'\UNt��>y���퓅��;+ٽ�\�^�}��~��W�`��|F~V�D��N͂fu�F��t�~1��-����C<��z
�	W���g���5&���~�ms�D]��8V����N�N�T��[�Ǽ���j>
�B�僅��2�:Uqr�%�!�c�_�����Oܷ�P�]PN�� ��{b1�Myl#�p�Ђ�Y�U,{�l}�gnBE�t-�bTq������@�!�ҁ{ۊ�+�u7�N�����q�=�h�"-�n:&?p���Q���Ƭo��wYW��ժt�:�u�ߢ��>�`��^�p�3�Ӣ��ض7�O�26�T(O�D�EA�m��2�M�Y�Ua$��L�y8�R�_�����Cx� .��]�%:0�2��r&H�pM��WM�&��xn���k��l�S�q�v kW�?H�JLHE�al5�N��mԟ�,�{�aڹ�9�w9#j�4.SJ�D��gD�N�:��O����ڟ/8�]�Ҥb�f����	'��a 5��	)l�.l{Љn�_�QԑX��騟y �@��z�4Ŏ�`탚%Kz�KhRȓioV�AE���΂������{�5�Ӻ�!��k��b������Uw>1[�;�+�X'� ��X�=����0��,��l#%�Q0c�ƣL����y�������`�}�ᗈINTϻ�-BH���{�.X�;+1?�*��E-3����,xO1�N�~�H,ZI�ߦ΃ȯ�9�<�����G�jEc�t0���LRo 1ơF�y�#C�(�6P���,K��!	(�,�g���t�V4[�]U���taD���_I���t��:F�|��i�8�Ď᥿C��=�&��X���^�e8v�I�3��c�;Z��ւ��R�z�k(KYiڢB�A�qK�J�5��ҥQ�����������ۀ�Ap)�e�A#���	���|��mlD�d��@������S><�:8���R2T?0V�%� �X9��p���he�[M*Kp�}��v4��/�ZyZ1[���X�7�a'"�t%S:%��}!�� '�r+�����f�4x�	z�p��Cͱ&�3w=T��P���ت+dv��0��� I
3�
�me�K`8���B������B�a$fsc�F���+�)o �wG���"�j��p.|�7�
���EW�[v���b���A*xg[ͼT���[��߬��*Jz$ǡj���˶
�"b�>4]�Z��.�R]:�7�U^��- �Tm���E�r���ʩ���R�XJ�f��<J>����Wc�Iع�c�����,�͆:$�
BD�t�4��G��c�UHڠ�8?��*DTx��c�!��=�:(^)9��~�o4|�H��{�݌�����%g�C��*���cF�6{��iz���3X��0�����OL䀱�F26p�/֓,1���F�Ue���+S���]t�Y�!��AF\�۩V �V3�`��Y4��䢻�qs�D>i	a��ʗ'��o�(�26._:�\b�#�ͽU�t<p;J8�Դ�)Ԕ��o�Y����e[:���O�~�w<V-���aJg�fX�.�m,��������+��? �:k���A
�p��.��*�Ll�bI(��u7������C�c�׶��[�N^�BSdɰ��6�v=zqȆ-�8�E͛�� P,x	n�~�g��t�6-	�D 2����{��E������4����K_Ca�G�]c���a�[]F�V�j�!<����'���ڐ��tB��;�P�_���(v�^�K$����r<Y� �w�t>��5O��<K�; [ќ�U��	�����=��cX��g����m7V@��P��&�mu҆��6ڡun�[�[U~���k���1�|���Ռv\v���/s�?�0 �)�qo@@�!���8��۵��۫�{�_����-�܇�S�b�ZP���$e�*�$�.e+�.'d1�a��׳�H഻v\��4��I%�-x� >&Y1����9�=Xk\:���&��4&��S|8��6�/�`�$�R91(�O��N�:�6[[<tS�Nj[*E_9|ۢ��y�R_!C�-��d�~��u�f(�K&�eqЇ^���y.S�ъ�i���r��o׆���z�9�ٰQ����v�?������\��KT��C��5h~�\_�֋��:	K��J��If����R߫�e�����qcbC��A"&���$#V�'�.���L���y�/l�h�T�M�k��a��$��W�K��Pw]�`�	QL�cG���>bJ���ɔ2oa�;G�(+� ?�w�dmW�5�igr�C}����#D���%�/'��=��|�٠)����"�.	��v)N�ܱv�W;>׮�ϑt	���v�7��](�0��o�c
D���1?�G�y�.]<�N_�\I��ᨱl��|�.�蔱 �o���R�6�@�uF��D���Bn*K�Jq"����\�9u��N� 9�Dm�)�0�T"M~|2ԏ��r���G(YP�!�C���Hw�B
��zgc�ɐ��y!k��_�cz*��V}�$>Q��Z��!���_����&��$�՝%�|�l�;�E��-�����h|�v��&�m��W{�oBmr	ZҖ`����YJr*�l�]��������X[����6A��%�����Ì.0�3+�]O2��ZB��R3(sw�D75�A|_�W'�Nl U�|��xA����,��O �AX��:2x�O��YJ���+��]�N�Wx��AE	u��x��{8=���p���EP}��ہ}�
�"�C\�zL��^�5
כ�U+������Æ�r_fk�1]�X�p���E�S�q��~��&�wȵ�cK�ƥ��d;De~������ݡ�;�ͮ;�3��0�ml@H�V�bR?1e��&%_�\X��b��}Q��*@��.v�b܈�uͅ�?)�H�-?Zwf�gP��-������Qs	���0� ?�_��D�l� �tQK5쐞rO�6$T(�$\�zpv�%��N"�w
�:ʴ��[h�OF=���h�l���V�� ��!W�}�+�}��+]dU���N?��B� c���
�l�M��	�~V�y��v�w��l��W��\������r��Ns�Z�qh��919YV~S��� 5v���cTLp �I��8��>۸H�*1V�hw���j'+�a4����E�R�p���3��  ��䩁"�􁄕Ӈ�K��K ���t�Ϙ�p�/�Du��͇�L	�D�њ��ֵLL�_>f�`�&���PND�L�,����b��X;<R��]�wO5� J5��Φ�F�g2Ͷ[�Y�V;��D5ҋ<�Ѐ��,�w��H��"<�
6U�,a��8���-(��<��p���oVu;wU6o��dɺ���ա|�������;�����y��ٮ�j���1�+y�i���XL�"�ݖ#ȺrZ���³�6�D=N5�̟R;1HJo2���A�=���7���K+�LJ�zR֥0۝�������i1U�����EUoV�ny�(���o�
���Ș���̖$��#�%č�r��S��Lv"�����K�4�D��:�z��(z�#����� ��N��)��o0OHʫ�9�;f��i�ߙj�d�O����[�l�����
♸7���p����r�&��?߫��()P�G���Q�>[2��o+��3;S wu���p0�alF��x���(���L}o����jf�0��
z[�Hhn�o��a�=ùf���xojںJx	I����6t1t\�j����x�"��|�hNA��b�p<TR���#�y>v&z��`KVh�׮@9h4Pb���TQ%��F���)�,�q>�!��7��Y�D��M�0�>�@鍁w؛jb�J��X#��.-F�(+e� f{1�ګ#�n�DQ~G����K1���ۗ�ۑ�|%�9�@|�-cb���< �:S��>�� ��N�����oC��lP��`ɝ�J
mj���������U������,��Y��dK�CN��M�3�&��=6;
%�,\�}�_�Oq��?7�{����Zr�rXw���ʽ�:�>&$%3y~C?"8�#_��KB
��D8.N#Ǵz���n�F�����bB���������ǭ�!�{g8��a�1�#����p��y���S�=��
�ܯ���`�
W�;�F�z�9%@H�F� �!����q^וpI�	����+=�Z�8R>e$����9��`_�*�w�w�/_�n Y��4�U�&�=c��y�0�h�.�~�њ'>̤8I^C��7��#����F:������vT����G�^��%�ȃ��`C1���������"�}s&��+~�~���!��� �:�]���(��,1�Bsx����y�m��+d.����\�w-_�.SP��S,�31<�W���U_�c�dTi��s^¦P`XBDH����j&yuWs��ߓ�~E����'��e�xݟ��ic���c^��Wr�~ei�(�9؁*xu5��%�B��C��8�:�����Q{{�T������+�Rϊ��}��ܪ��Q T�Đ?��o����I�8%������v��tm{���q�Y�dX�x	�׊�nnU��<���(K���p��jx#n}��Jǔa�<v��������\�!��#l��l��>�iH�Y"DQ���� 2U�7
���E$p�4���?�"����j�Җk���h @����E��i��#_D*s��J�p�}�L��M*Pgb_��oo/3onФ���d��8�5�q�E�;���Ԭ��z��SH���� P�P���z�O��A���DMvC�_c���JB3��OV��c�U L�
�,�~s����}���S�D��ܣ�"݉�n�����OGm���?6O�<�7�"�SJ�@2�t:�RM`qs<˻OB{�C��w�x)�\���:l�GD�V)�\�T��l8�mt��ƨ����u ۺQ��JY�d���p*��~	v&{L���t���ϫ(?}�#��.��i�-1ژ��ŧ�	�uv9�)�����ۈ�vV
9Ϛ�R�5��VI$	�HJgȉ�>(җv���=�ٔh���D#y劕*!O�p�^�H�t�'�%:�)��wb�K�+���=��rb��ڏ�/������F�����1���ȎĸT�&�5w&�t���q��T��K��K�#\R?#q�kD��m��� �Ӷ�O�p�ų{����'-�磱�f����Z���d�n�;OI)�j�t ET(n�
~�'aG��V4Xe�\PR,�j/��wqթ3���pzj�/J���ṱ_nT�LVI�\��w�gl,cs�z<j��!=�/�呺c�8�ga�����)�HkG@	��xކ�4��1�cO��䀹�<Ķ�:o��K���rWG
���d���u8��"
N_�Hӕ��[����~��W������7��c<H�z*L�n����89*�N�-����Xo�����C��N)�ކwJ%D�^�2ሜ�˨%�׼O��JHa�d$!,b�)(zE�>E'=�6l1�Wd���N�L�bʘx�Hs�|��B�ջ�����5TD�T2��T���C?;���L>�=6Ko�nFF�1� �	����$��K�V���4f�n���im���c����H�ĕDk�<N�V��̵����c5�u3|Tm7�î��F�t��lo�4�3��2�����u|#��-<��k��f�.+�[� �;*fUަJ�i	<§��q�2w����[��RW��8��A��D7�^�gN�d7 q��R�8csz
o�HzK�YC �:��;�#��B�{�ڞ��On���!��U�U��5Zћ��J��N[�:��������KO�5��^�e�'���f�б���(�R�L�c_�)f}�"���Z`  3u�!��������,~�Ȭ�zi�-ީ��
�)ep�g�o�$ $�:3c��g��߷�]A���W��P�� ��_e���/�!$�U���I������O����BzpG,�,��^儰���oE�&A�Ô��6���v[,/�eer}�Į��6��ʩ���TH�jW� ���Jnv�?C�]����K(?�r�[RU����}*�"��\^TAz1�+�����m��3���������4P��Wʣ�X~�u�,k�]���_7D���8��Eu
!T�[g:�O
&	�TqB�](��Ky��B\m�0� �ݾb�m��ޯ0�;�b��d �WtΠ���]\���%�Zd��Ƚ�&~ޞ�܇9��&��0�;3i^�TJ�~<�ސK� �2��}p�%6�N'Ґ�e���ǄG�۝�{����ɞ(�� ������y�(V7�C�>,�h�u;�t�e�$�w(%�+Lq�lS�,���,*%/Ju$t(�Sf($�(��t�r����w�[f���Bd��מ���
�w�*��V�'G��!.�Y>,n��g��~�j��0X8�7��bx��J;��N�h����7�}�P|�N��Շ�=�B��6!�my��-mհ�j)�X��ܒ���s',�~ ��m��l�,��SI�gT�M���T�I��QŪ��Ǯ��z��1�{3N�a�gk�%t8�&�x���q۸t�AӁL���m�y:G�4����r	f�tX�-��t�q.Ӿ�M*��Ji�;��u�<kqޘ����{N4qG��W��0�aJsx�%��8���m������]w�c���c�KD:ٶ7�7'%/� ^3���-���M�t����L)��x��,�Y�u��w��l�+�?�=H"�O� �	�$o�yd��gzP�Ժ'�8P���(�^v�o��������~;a�Fle�'Dk�	�
;���kBPq*��m���m���������`O�,~�i4h�*�ǯ�M�Oj��}��H @�6Zi�9�.Lo��Nל�J�^ ��L�kC�� ��g��Q���T�V.�qI�h�ٷ��Eh�t��.T����s��d#�Jͤ�C��Wϓ0P7U̪���n�ʢ!<��t�q&<�n�E�*j{����)5����t[(��Z���0_�O���{�F\�a�e�l�#����o��ek��'��8/�9ϧ���R��	��ӻ�&74�R��*�=	[���xq�j�Sp2��Z��|^na�4L�jTw�*=�ߤ�0�����1�Mߵ�F"��BR�20Lx�b0�.~��(TJv=Ip��P�K��<(C_dn����\��+]Yj��v���Xy��:ZN���N����l�ֿE�.� |@����M�����Z0���O���.d�Y��t4=����x֌�3Q��֍ƸKs�Bʽ������H�-��'�5���vx,~������'㜘�X�X�<�*�*�b�V��z� �>��I�;�t0t7�1�mIcfL,�� �g�"���^�d"��s� ����I����6ԯS ��ޕƩ3IU�Kx1NeZ?�^|�.� 3T L�ތ�K�Ϙɂ���N/w8�5π��y�8Nv�dR��Xq���211a��#8���>�S�����-D:�,�]�ɪY���\�P"��Fy��=�5�#��C��~�2�TJ�ȿ{�t��&p�\���4�h$ _�:l� yM蜴H%�Zhb� vhj>�[C��,�LqY8�8��8�e��O�?~�7d�$A��u�T�]�}x�b����d��c�"3�le	DMZ���7�����%��� ���2O�K�0������S\��K��;���@ �N����=K�� ^J�Y�p�_"��c�[���]��@��-��nD65�4|�� ��uj�T��YL��d�� 1,Y�ݙ����V0�e���Bqo�򟾛
Ȧ����xj��u���0nX?���5�Ň�S\������Cb�
��*��zg�P�����,H��:�D��r���O���0s��9���z�����u���r��^��z�HWa���a'Л�c>�ȋ���rzU��̂"�2ve�	�P�����gxNф�&u�@e�ڰ�n �C=�����sۇ�m�FI�=o�{ %��hb����W$�w]EBd�Y����U|�=nƻ~i�][���LR�A����D���d��a�hbY_̓g��M]z>���c�%�?��5v����`YKS-�gr�f�x5�kz�L�M�E����M1ٛ�����ٯ�ǳ�����6/��w}���"�m��(Me䧎�r�����<��.��!��r�ϗ4�6���`�c���M4���-)�߂�z�$�PՑ���-�]b�z�ZZ���Pl6��م��([^=uv|>۪�˜ǩO�3>o4��N�&�뚴�<� r���I]��t���*-���[�ǨW%�^�ɯ�L����*RT��?�g��^&Y]0��?I�L�{��ӥq;�����Cg~޺�*>��vX���F�е�eN��>���_j�u�$}�#B�&@�4⎪K�Il��Z��6�Qn��0��Ī���+S�x4+e�> �M�h���>�̭����{��B�JN��������JˍV!�ZG�q�5kEA�-������PM#����w2�/�9�<���i�?*��`�9,�`b�+ނ*����̡k��;9������Ĉ(3�m�EK#+��bk�S�-��vw[7��,~���bw����]��r�	�I-�?U�>�B���Hhh�e�+�����}j�M��lV�Y��h��c�/�P�۟�0�Trƒ�V�Bs�<{I.��(�ww?�&�� J(:�����ߓ#i�4x���mY��7$Y$�5�[BhFH��-~�Eo�W�Ҵi���H���x��hBi�q����!���������ܲ����+<���u �6��%�;�;'��oJ�#�Ok8�F�u�'{�#v������HoD�~�t���Sv��r�t�.�y��}g��8�p՜V]��	��=˅�Gݿ�0t^�;��b��wm8��+cRH�a[)Q���/�$��W��f��v ;w[���$�*hV�����2����`��Ac.S��h�b�&{����4���9C���M���!���	�Y^�������U�[�db;e�X��d��ɏ ��e����?H��"� [8�����\%5�H[,�@�V�x�ʿ��sڅ��ͼ2���:�B��bu1_�ynL>l���b�k�-�S�˨\	{*��@�"�r�3S6��16�����T��𱬭�x%).:3*�ӉuV��';kf�Z=�����Lۂ\cr�Ϊ#I��F�{z�lp	:Z�^/��]wX[�$g�bO�w*�>M�{U'���EY��س�l(ؼ�8��R]�F[]ĞVg8!396�U|՘6?��
{`��ȡ���	Ow�!+�vTZU�y�t`+��ӎ��!m�Y��0��
2"��pi���)�����ۢ�F�{cB���PХ �L܏n�=YwY�41{������Yαg�|����sH�ow�愹�������d�Zx�C�켽�7�m��Zq�l���_�	f�-Aܒ*놂+^��_�
���)��.J�m"l	
	�f�՜R���̬qd�7/'�A��J���W-��02�'�׆~n�6C�y4H)��/�P��\�� ���2�c"sV�	:p^K<,d2�7m�<�Q��bRu^*}�Y8���%('c*�[n��h��x���y9��="#_G���o��8��/�[r޵��/��쬨���.��]����:��7��|^S25{�~��!�qEZL�ћ$�!�e}���j�,j앰�+ܔ��Q
��답�'6��6����P�O����G�N�Í��u��r�:%@n_�<t
L��	`K�R���4��ol]f�p�f$"Wf�J$�0�Ƥ9�D;g�QR�<B����f |�E����6o� <*���ף��
���D$�[r[b�D2�T��ǒy�k��M����Q��a��o��X!S���Y6_�|q_ه��.�k�_�Ϥ
��YY�PnN�R�7Ā2p�ȕ�[c"=v�@a��|����&#�&hh��������M&�!0������P F���]�*n%���v��fL�a���8����xzPY��*,^�,\�p�M�BX�<	�v���!Ol��"��]�%]==���w��T��Zоf��|����(h�ts�zԐڸu�>��q�C�
@���eȼ���I�b�q2j����������T2�4Q�IV>J��Z��#�A��?Wp��c���:X-�|_t�����A2.Ϟ�:��L�����#����{�9,׆�-��s�2�&7��=��s��\�
`��v�Q(��]�U�O�|c�����k����G�3r:0���+�B�e!�)f)�V-�R���Q�>�<I�i	���?bL����@�`�3'���^����U��+A�wU��s�����(�����t
[s�gq�ܾQ��#�Aj��6d�qB ����*#��U	���r��H�9Y�7�ng��P���#��׮��� x#���,T	Mf��,��bL�mw�$h��Y��z6ִ��_+ܽ�^���\�{\K����r���g�^�r��i��*C�j>9������a�V&/�e�n$�t�ŕ?��28���:�Tѓ�F��N��
�c�	�l�MH�����@1�״L�vI�S�:tf9���Աt�4�w�F���RO��Pi�43���� �(W��s�9H�ijb��L��m�%5Ȋ�Uv�s�����2�1t�����n �N*��>e��'�	*֔��{|#�+l'�RQ�RV�,KH+��
���:�qS�@^9?l�GR���т��Y��n�`%�[��T,פ�Y��#��5����a�׭�Ǟ�w���9V@���X����hg5~���Dt�M�8n��Si���#?v���ټ����a�j�LH�t�?A��E�� Ԁ�=�By�k�b9�W�<
1ү���%��r�
��6����	�I�{?Їc� g+�����DA<�Z$��0��,���f����T"���)�9���5ʗ%X
h"��g*�����U=��S��Q`v�������E�D>Q�c�<�@у������\1�JF�X��� �Nc��8&r�_\���Rc9i�l3k�N�t�K�7��Q���ɫq�J����+�žQ���ڭ>�0��=<�9�A˱�����{p�#�d�g��;3v+��tF�� �I��{��X&���t\��P�L嗉1�48�u�� UW�Ա�!vrь 
8�6u곚���Aw�1m�D�\U���@��Œ5�Ng;8n�B�������!�:��'N,�?ghJ���~*ߋ�5�$�����aA�Ga���F1�&��M���X����&^�.�z��J��r���u�:(�0�`����X#"ğݘGs��h����W;%zN\#t��e0;/�.qȬ�X�$) � J���|�@6u�%h�\:�f��~7W�`�E�\� ��[�@����r��
��P^�����1g�3��r%���E^���&��Q�kx�e�%X��WA)^y�ֶz�	�3�j�/�"[��>,�� c\������z��%s�Y��`�������!GkP�F�?pd��Ov������Zh�5a��#��V�qH�}����=eS�;a-ɼR�WdĄ}뛁��~EA����/�"���sb�=�o��G���=Kuѷ'��rԲ^���"@�@t�
Y�bu�h�p�z�l�᥀��:��$����Kc�����Ǝ>ir��e�Q���&Y��T`�K���	�}?$�m�Aչ'�em��<��Z�y��������dG��M��m�V4��;�Ô �{$��-18
����O K����}���;pB`�T�Z�G����w�I�2����l����)s��q���ȫD�4Ԉ�@�|����G����S�vC<�zJ\���� �o����qr5��R�bq�9b@oP�5L�cXQ^/P���~Ѐ�`ZN��n�~/���伆m��*��I?E7���T���k���(l��h�$tԻ��񡄊$z]�p+�1��ez����؋C���KΜQp}Qo5�k�Qnw&����{:�0�>�7�zY�R��!@H�c������^��J��+N�h1|��w�&�W���)�,�Y�G2��_өy=<kz�~�~�~"9�B��JsR�/pS��,u/�b���N�o6A�!�aE8v����s9h��H	A.���Z�$C������Θ����p�p� ZU����y���xX��H*ˏo������l=�{���_�b��ep�	�Tz�>S��������#�vv�/?�c�E�9��QGY&��4y���V9nNܘ���
�/��&��W�S�
��&X�.2H���'5ۼ�6s!G�8���EҔ���Tڂ`o�����,�%D�(D�tNŨ'�j��N�=�]'���~Y�g��<��WpXIZ��_BA�����w��61�(�_[Q��`��i��#�ա����\ch��a��󞔋d�A/>�FXQ���c+<EE�!�U��*UND��D���q랶�F��U�O�}A�����d���Xs�@5{jL;�1��?f�	�I�U�O�o�H��jn0�LFor!���D&�:�n
���R�\HgĢ%�2���t������*�(N���;�!�჆e +�#ɦg�і��h�S�E��s��R�	-E�!}pc/�V�ҁ�F�z��`��w���o(}�[�4^���^T"j�d���a�W�gT��Fȴ�h���'�G��WY��}�z�?_TZm~_$Y6'�lV�!���l�,�X�I�K82me���;��G%�xh�>��GO{V\��vY��� χ5���\�jm��U�-)��@�j]#��(�eI���J���߈�]�)��'�b_8-lxn�t�j���z�v��l�]�
�V�~�ΜuU҇��#����2UY�bw��F�j�Nؗ$#���v4�����ԭi"�Y�[�<ab��m+%s_�Q��4`׉.�!�0���B�Y�A��B��@�ܥ<����v�@��Գ�TcR��d<ɀ�,[Ǜݮ����-�B�T�d�x�� ` 	E����?r1��h�����Vä|�|�=�`eRM1���C�B�].���bw�k8�C��=��\���D[���� ���b��[�*������\�dd��nF�&6��K� j7��6���q�������~V~V��GV}+�yJ��?��/��AG+�y�|�l5�	�.�f=:��G8�Q���ډ� �6v�d�nk�CM��)�*�1�!W��̿��	��fP���_�t���4�CЂ�T�d�{���X��m���y�G||2�U�Y X&���{�Q�{���2�8rxDY�y�������M�!	WX�Y+^IFcOv�Y��k2A��~Y�c�hSOj���M��j���sE��og`41T5�t�	Z�r(��Etu�r ��vç���.������̓������'��hp�GE���U�>_cje�qΖ�t�oJ�v��y:�Ӿ��dc�jx�E#m��ʢб��\�~�AμD'y�i�[�T݅~�Un|����u�~�T6}S��%B��#����h;א:4,4����jL������_������F
+�/
�+1e��^���!K�U�8\�IC0���,�ό�)�f�0S�O�5"aKm,t�	�u����,�~�n�D{�2z��J���4��h	�`��;m�{I໼k����5-������ɬ�w��`����NO1fPKEg���A3[�k��*�c�͕��D>�`�Mk)�׉�i��PLP9�Ob��� �F.��[�m �U�9�X`6Ж�w��,�V�� q����4���$�~���R�<<�A#Mr���彜'���#��/��)1uJ��j)Q49N�������X�:P��"_�	�k�\d��g����P7��z ��L�	1r������M������K+|vm)q���}��
�-��a�n�F�8���0�������smm��"w*��E��"Hܜ\�0ۜs���ր�oá�Ѹޣk)����8؅-����[�Z��MR0���g����n|�k�)����E?0�0"�7ƫ��@�;�E���pȓ�}�(����f�6�DVMG9^{x��_&���]H��>5-!��=f`�"�o�����4�!N��T�"h��N ���!F�vDr/p�|drh	�M>\B:�d���:F��@6��|Q g�궬>9x-Y��5j�/o�}�Äf���jˀr��F#��-8e�bJh�0�L$��p_��A<�w[��@P�-���)=Gvc:I_�����A�u?�ʝF7f��	6.6����CB�(�(Ta� �DV8�Z�*/&ף���*�qF9��5�2`픙g��٫zg�����XP�O���&8Pn�����q�{��[�8�hX@w���૝c�݁0�>��5sn�����Z
��ͣ��W֤�8��_�=���['8�b����q�z0�$�zH/�5�F���J@����ƭj*|G�՜kI@�
짼}y~b@Y"��_Rn��ysv>��L�,#�#�)(�X���(��q^�M޷�R��{O�h���h(>0<�8���z[�8v�� k��ܕ-�������T.\'�hv�9���OT�m��#^�ș������H"��H$�H'2[�_-S�k��	��#���E�|�_���D��D�|�r���<|J�H+�1�ͪ�H`rM9Gv��\-����y�/ҡ!iԿI�����?Ub�� Y�
ے�ɍ��m�Yٌ���,���z	4��s�V褂����/�s���rr3��L�1������v+��1�}Cq�P�-:���@�~|C��5�W$��W�����կ*I����;?\���X� �jÐ�셺vH�-?-�yCT����w�c����$��P�aZ#��\t�!W]0Ee|�z�%\`��\���@Y���U9�,&�T����LPiZ��iz���Y��>-a��Vw��᥏9�E�7����!~�)=��v
GH�ܗ���Z����qW���2��I�Jg��\ê㪻O�3>��ܴ�`X�F�U�vܼ݆��b9bL��(>�.�w튈j���gؤ�~��A�lE"�Q\Y? ���a�.��ٛc$L��?�>Oĭ�h}q�e�8V�F�W�o'���QD�lz���`�F}���� �wTxq��{�Op�3Ѱ�|R�]b3/k�����8ڊ�[в�PM�H)M��1`tμ�%�&��U#<$�uz��_>��A�Օb�/���&�ޓ���Ux�ЍE%`��`7<�
��[��$���{7T�|5�uO���29Kx��T�s��ɗ�5�A㦪��}�y���b1�B���ߞ��s��kO�|��e׉�����q^��0�n���V&�����@q����re���0��T���!>]ɭZ�P�}�.��N����gd�wD��#̋A��M��}�P�D��t#]���Vɲ"]��y�X��$pj�zY}�.��L!&�,$d���G��.͋��F�q'3�-�ð�����.����rU`����T��1g �ΧX�`���V���J̓��Hg5u�-����*{3z�r?��_�@�kQ���>� ���$��M��̇
���]t
���H�)Z�E�����a�w��i���=�f��3�,�.�r.˞9O���[)�y�{Bcq+N��v2�'�y�:����%I_k)�N�#��=��\Y����r~x�a�������GZ�Y���g�p��uKuҍ������-P=�����1��Q^�g��~p����cF��o���V�J�2��e��F��5.*}�ľ��6$���G���:E�~yvȟ��j��߁i��$��1��1�xhE�w�!+�;���G�\�\��J�a������L����%�yo�?&�$���"8˗+�|VԂ��/�C��+G�V��wꙷ�o�l)6	L׀g����6�v������?zW�q����w�@�V]a��������M����׺S�aw�K�I6It����6������C2�<��B���3x��B��oj��U/7 ��)\X���+W�,`�Ƃ���태��o���ֺse�;�����G��,���� ��d^`1~�m�C�;�H���Q�����}����$�����o���J�[s]Y�G��vH���_#��ZC��E�R8w�$�L�iG�J���V��Nz�5	��w}[ơ��+��icS�:��-[4~�ֿ@G����㜶B+�^�1th��C��|r�7f��!�>�j;�]�20�ñ ]|��8�(S�Jӹ}����rw�t�!a!����h���2S��?[��6���ݖ���k{�7��̲���H����9������qE vЁR=k�+���p�����RTF��&Q�G����	���`mY6ǹ�uaN��8+��f[���1�+�n~j�hR	Ɓ�>�ZK�]��J6v]��y�V�������&"��?#��_��_�]��V�;g�}��ڂ�W�}�[Ŏ@���߿�_����ZZǊ��(��c:����:�Q�.���A
��8�}~)���y�0/�_'�"GV�m0<aF� JYx�lU��ī+hI8�#Zj�z�?�Y�@���|�hk�ć��U�c~>z5֭*��(�ߛ+ygD�'�^u���Ԯ0F�7����� K� U�9v*�N����#�փ?���
��
q5l%P�ba�_*U�x���ܼ!kD��^17�>~I^�N� pϞG��}�}�Q˹�w��3��'��ݬ��i�7����s����&���Ap8?�\k�_�^(��p����c�;������bG,8�.�<w�V��yr��ub	 �>�>��Ax�e��=ߓb�����d�i�ԃ��@�`V:��~��2�U>)P�Y_Bl�~I�*,U,��	S��5xo�[���&R;�HQK�nh�Y.	/��*��PDl]$0a��C�+۵/ O�̢bc͠z��b9�q��NEċ,�(K'	d��׼���x|w���Cx&L�g�)��%��,���ӓE�'��p� Ξ�+tS/��<�Y�����0�P&j�ɴ�=��ň��F�O?�b8���D�S]�Mc�6�d}5��ͧ���þ(Hf| �[��-�৒d|'����"��p�*�t��7�j�șf��2���jO�U��n\�~6���S�9��q`q��\-�K�[ͷ|���zA��m�D��5�A�ӭ�]Rj�9��K4�/�̉�`5�D�	�Vǡ�U�3��ӏ�q���v�!7�{�Z��U֬LC��+��)����^�)���[�X}�n˝��A"%ɡ\~�!�P��b_���E>v �����7�Ze&[�;��VU����IY,2�6�IS�����Lz�����m�dG��]�kh#��b��(�u�Hj�/ڿ�L��c�֯�j�K�?IH8ې�~A�k�l��E�;��4��5�(g�+TJBz"�vT��p8�j��|3i]N8��4/.0w�66╼��o��y$v�5�:���-�2�Q ���$�J]LZ�Z �o�%��� e����A��O D��e[�/3���s��t�PL%���{���/�k�� ���$�
`<�� �B(�4��M9�x�fڳ�;��i9�q)�G*zU�-x��bR����I;�q��U\��uVU�;m�P�(�he�)kt�cgĢN��E�݃'�/�����6/��X���S	��U: �d$�:�0�T�-\�:S�a� ����T��#8�����%��'�4.T��@�c~~oiE<4���u��{QOֶǤ��\Z��t�����$��w�%>ʌ�N03E�|b�˘X�g�w��ؓ�y�TA�d3��_C���w���B�$?1�UL�Q�vMz
ѕ\���T�9����4Ug��*[�?8�dh��#�p�*��f�d�����)���	�/�c�b?pIA����g�s03�I�N5����%�cv-06hcc���&8~]�Z�6ҜCB�3��:Ι�l��69g����z�'Y�{���R�1�uB�|�;��kT�?P�={�Nm�JT���l��S��t)��`,���j	l��K�A#\a�pC���m>k��2��M0B	�2&�+!��Q�*u�M�1���_]X��,Z޶�,�C�m"����c���RI
Mc��[�ڂ�s�Z`Q���ԍ�R6>��_��h�/n�'���"릴�R���J���^�n��2�6=�(�p}cɅ�a}�Ɍ��T�jY.�<ڱF�麑��)B }y-��9��>ö(�瘟��������\���SV����&>!���*�A�4�X�K�ϑ��KG\���wb��˘NL=|�k�&/&�&�<�*����d��h��٨���r�{�	���郔�
�N��f��L;��V�i�.�ղ���2#'QN`$���B����A��i�
���g�,�l�����N�hhlR��*�<L���푝6M���3&^I��)x��~X�����5�q)�&���()hU�Մ�>��D}�4�K��ȫ��-����8�+p�7�]�A|�ڡN���,���/��Ϯ~�P��^%�*i�fcp�H��7�,���1�ؚl�!���#?�l��.��_�v��S3l����c%`��EU�x�%�k:#/^��\����=��uN���[ 敀
�"�/�!Ǆ�8��m��M��}r�� ��]5:ү�L�Zi���<�wq~��V%6��}����v��7,s�2��/U��$l-?���@,szD��C�]��]�H��x�O.Ȯ��\�������	�����4`~G��r���깢�PtV�nS�]`E<OeP�QK�}~+�Mo`Eg[��>O$��J[͂�˖O$�,W_�����p_ˀ�tR��p�ꢗ/�e�PE�Ҧ�v��ڄC��ts��l��b��p�b�j���� ��U2��~WZ9b�ʹ2�&|H�K�6�m_�"A�
E] ���.l�p�p��S����Ц�ϡ��եT���U�p�6�+'�����D@s2F�<'��$����.�#�1���Q��:kG_峹��<�D��M�8o�G����������9��d�d������]��`�UM
ן�G:ɶ�Qwm��]M����me�q`��x���Hr,��V���� )6�i�_躳���T�
w"ǚDV|A7�<]S΃�cqi�CM��R[��B��\�f��=���Ѱ����՚/G����"�"mhj���uRh�������T(͒����+N�Y���+�����T��s�\�њ�!�f�d�Ϟ�5�a�H����)o��2}�;kX�*I����H	�(7�k/p$��lS%���b�8��m���n�<�	f�ߨtߎ~#���u��L�xe�L�:�}n�-�!7ܲedN�Ié������E���3m���z~*ʂ����)�o�ɖԅ�����ԋ�)��lq}�V�m�O/�G8�+�ET;6ᆲ-���xi0:�����cՓ�0%ֵOL�W��Ml8�d�p+����̮���_���1-v������td�1�7��G@�v�3:�M������
�'z�NB�.Tbd���$�x�]��	�U�����6�Fx����y�l�'�7�zd���օX�ysw�Gcw�3�g����ƹP*<���%w�f��p���Ysx�p�s��ml�_��1��D,��RS�)���^Q�e�W!Ɍ.8���a)5?חdQ�V�l�BF3�[���W��},H�	�M8xU[S�U%����Jt�mT����	Þ����	Y&�7�f�khjFa��9�6�<v�+�DD�����,�_�h��!�Y�=N�8�7[���4K#?�Kc�"j1�@�����jaFđ+����h�t��G��3(?5Us@�c(ݙ���9�J��'q����k�x�,��s���0�Y���!�h��c|�ʢ&&4��A��U>��[�����b%={�KoǛY�ߪ���6#I�d7�"�M,Wt$) �D�"����0�͌�PIw`&9n�d�����R���٬��ѥ�?̬J��$��w�qi���lGJ������������x�=�J �.c�E�#Mء�w�0�RjZ��D�>�*ԹyA�|��p�'���蝑��D��%m�fv�62n��b�nʧ-(����x��rv�Iف��
�u�t�:�,P��F&��C������VN�u:+�R(ze4U1b��i�oE,��+������('�X�m�9P��r{4���FRX�����U|�ƒ���@w>�Rr�L�~�Bõ�`�&ӿZ�0�k<&��K�ee�r��2�=�A�%�W�3tVp|��:d|�bY���Rn��7�q^_��j�JԴ7Y<�t[��]�3�A{l�r>�kQ�����?�iZ��U�C�jT2�N��X�� H��ux��m-�)�:�4�YV���T^�ݤeB*b�
B�?\zxo��a�s��,Ťi)w�F���xMX/
q���>����4���y�;��b�Jn���ڼk����,$z|}����J��+�`B���Y�I�X�T�}��MF�����!By��/��a�u-v'�� ��H��<?ftt�U�&1�6���Ku	����`B��`N�����$���@��چ���U�ey�u�7��L��=�I��ԏIlU�0IT���������`�\���cH�ȟ���-�}i�~���k诞wE짯{�FU	��xN���.�8����TK�&�-�����ܸۍzl�Hb8�h|�F)��{��#�%����!�0��-";����aK�o�Ok)�~��?2� M5�}\�@,�]���,E��'(j<���j�+?�jᡟ�����v�H��.�F�u��MT�}���^Z�T���Y�*��y�=�^�3Q�Si�1�*!�Y)�[���Z�}�����Q-�;��W���gI[�$Ү2缰ߑ��|�nL�e��L$+��a���o)�/LI^�@w���%�^[�7��̂ �E�#�J�n��r�w��" �{�D��ypM�;�y�%F�����ڪE�dj�	��5_uu�����zg>|������u;�����N�N{��${Lp��
C\[�0�Ti��P�����P�O��T���ث��
�'{ዯ�Z�.���R���o�#j[&��*h�
���eĊ�ሧ|�B��zV�f*�9|��!��{3=P��r��8�����Zύ�,��ȯˡ>�pk֐.�Z�E\�ҵ����əry��i'��p�9b��{R�/�5cI
+�b2���z77#��n^e��H�x�A��R��E�޵&d�R�و�[�I�^�؝A���@(��ڲ�"�7D�$��)9Ê��IBI�c�3���ګ�V����E�	;�D��s=���ʠ�TWz�`/ۣfVF^��^20��Z5��:��><Jw����w>���+7���;\e�?�+�c�p�DN�\�O���wz ��c4�P�'���jz׍���;A��������:|�<��7�$�J�XTP�L�D�u��,@����Z�^�D��%���4��Dq�9I�#r3,��}�>�����B� ��q����}�\}��ܔ\	�Y����(���yֱ̧"%�D<<���	��3Ͷ8ї� �U{�Nz�;�z�_�+�b���t��b�"�FgW����$]I�z㉪W/�U������[��BY�8:�����,���י
�v���KeL*J���O��l�����l���N��8��_wFy��͂%�6�F��O�P��%�(t&���j׺����NϚ%F��^#�������Xj)q}?�]GeM���j�q�y0Up���J�e�k��Hx��`c�a��Zh��xV�$�}�����EO(o�H�w�ů/\m\F�(���-n��O�vo���N�2�v���8����+��u5K�.�I91�1���os5���-�b�$
4�� ��f�连���d? �iLX���A�Rȅ���@��'��l����6+�zve�I�2�X9 	�q|M�yoV��@����E���0�kub���.�΀�
 �xJ8k���HM鈜��������D�#�ֺ�/�E�%9� �y��[�KW��Onl���{A�Z�����G���ٽ�L��l!��u�:��
}CR��L��[�*� j����%Lx�A@+� ����{������@�>���?l
���ٗw�1 �3�ʛ�ʋ��+�ǁY兩���}�|{fc�#)��?�^�yj	8�|/��;��Ą��[ӗY�|x1Ro��'��p{����uv�03�rAeɝJ��8['p�"���Z��M�xG�v�U0��a
],]x��#P����.��;�"�YP��/���e�p�a��~
�J��쮨Ͼ�/�<��.c��^���7y��o��� !���c�-֔�F�Ř��Ň��*ѷv�����	 ��,c�e��>&���	1�L��:3�㼓_谊�^�sq_^��K��j-�]m�[���u�a��[$�S-t��Y/�!�tMo��3b9�K�*JM;!��dŝןp �LcÂ8Ҏh�}�K(o��d"eU�*�]��8$����:q+&�J�c�Q��*n�$��@��U�K0_1�y���>d���L��g���\�w�y�Mn���<�$8�+��&�5|�M$���D�[#i���X�I݉�܋�Uso!H�W���&�a*�I��W�4���ԇ���A��5�؁��x-�8���p��!�q��7�_�mJň��:�[�l.�ݴ�,��M�i�m�D(o����������o8�`u��q7.5K=UO�g�ʇ����}��V�p[=-`����\�1��2�=��)�p���7Uˡ~na�!;|���0��qhx"M��fɸ//j:Ǻ}p��-�vh�5&i�O�7�ޥ�0�⤾�?�%�D�C�M������P0�4^,�{�Z�Kx�>��
�����W���yD����~-=)K�դ�jμ*�<Xy/{Tv�E2;���h5�ؾcǨ�]��]�m��Ә�������2��FPEtO��oc�@!���H�ޯ�.(Z��5�_s�U؋�������o�~F�f��:?�2T��QNN2m��ۑ��VnB0t��D�4�����A��	�� "�	��yI�2Ԏ�v����b�/f����#�>�,F<�j8M�6���3âoH)��� ��E�]�Cq�F&��8<c���v���H�'�x�R�|����*޾"�x- {I,w��aE�h�	!#�"��h8�n����+a�j,��]X��B��y�e}o:�1�v�P��ț,,pRi���E*\��z;S�[f�$d��u�9�E	5��#G�$k`l]p��>K����4,1�G��Ͻ=Zx�QF�Yc,b��H#pnQ�Q���X�y���U�,^���š;@p%E��F�C�z_#��O�Ղ3}��D�'�wǫ�E�@��O�}�U�ʳ3p9��康XM��<.$|P׍�a�単~��x�V�WJ����hS�D�*�¸D��C�W(���1��l�7�����_�#��E]�I�12r2���nXw��h%�[��\��
r��Y1�!��:|�N1۝�}�����޴ÀG�)tE����EZ=^v#-Ѭ՛���]�@4_j���aIG��nD�ӻ[��ӕ�_��L��
q��R���0J�j�N�y^Če���5]�)��p�^a,��\F^�`��ںc !�I;��)�h����+�Le���.��y3��f��&)T�D���z�ka38<X��G����a�+_�ct�ȫ�' Kh�<�����ӭ�'E\F���M�Q�]W���
*)7�V��y������:7#�䎘��1��낵=��eΨ���륋��`���QG�-�3T�Н�R��J؝r�
��x��7�2%<�� Psޓ�	��8���T��ğ�:�M�q�D�U�Y�{o���d�,��,����3β_ kg�d��L�%/���
)�A�(�F6*�b�o�n��Zݥ���઺t���X<�t��n�O�<sci�r��N_����b\|��+��% �q���$��[����	���<wQy�� !�Zk�EL��κ1��<�gs�d����Ch��u�O����X���n�@"���wQ��ːU��x'�y!a��9��̽,#�|��[d����/�59�j�n?��u�����~�XػnE�P4��c!�ӕ4V���RLM��ז�{�����T:8��Q�v�G�� ��{�#�ʖ�G:�
��r_�йe�q w��U�P�A��v�`&�
�[e�}����N6:qZ>��֓M�}%��;�x<4��p3����*��H�U׻�o��P�߰Z�_?!_\H9������u�C���%7�!ѓ�o�U���l�&#�C�*O|~u+��%>�:���Qw�񇭹�Ƴ�֨ͨ���;��N�vC�X��>��Ύ>;�}Ir����D���z����O^�y*W9<�K��t�=	�G,YF��qݮv��3��(>�z��|��V�FV����67xY B�@�懲��#lLԸ��-�v��9���[ܹ=�W�\�K���ʑ�$f� �?�c�q� Qu� �8��g��Ԃr���׭s?�R����ȶc�Yٵ�B��~W$E�[22R1�������nXkYrF�R;%��R��x,�\��ԙ;��@�X�P�SU�&p�A�ݐ�f}〗K�_���!������P{q� �',[�,&�Ӑϋ�%�k���ơ���6��p��ƣ~��R�n�����|���(%�a�p�C�g�Q�h��#������]JI���m02@8�KUg�3��3��7ƈc��{��n���f�{��3o`W�� �$�oR4v/@C@���c �+��@�%狰t&ϲ���M�����5�����_o7]�{x͔=�-r鰼��Eg+9�N9'1}�<�J��]�%|ʫ���eˑ���:���F^߻!.Y�@�����*��@ވq
V�����׳g���g�Á��K�S`1��z
�G��{�G,Z��V{��k���1os�l��]�Ϛ��t����4u�-�$ϐl,Y!�!��Ma~��s��L!�5x;yz*�4EM� 1'/�s�S�C����j�L�>$�u�&��xt��;_c�R�omU����4;���?���D}��|�;6��b�^���@�뭛y`u��ٲ�,�^��7���k���߱�A\G�2z=#�B�G<ȁ1�L__�3�#e��qH�"*{�5?��1����Q2������;��N��S��9��K����$-��r�'W��U���0�ɳ�)��q���Ԉju�ܦV%T�s�Ʒ��'�ƺG�"��(]���.Ͻ��H��ʴ&��B]�?fA��Vr�v2�M
M�ب�`	GgAÖ���ᾊ�{h���^������k��;��4ǡ�;1(i56�ݖ_�dLڅ-*�Mk��+*��{��V��H�E��W-[���﫡�3 ����{r�W�2��g�	[�#핒`&����q:�p� e�����"��%��F
�7Du��~�dn]���/5\�3p� q H�.
���[UU[%b�Xw֥m��HY|��:�95)�R�4:]�&���էګ�r�I��2�S�n�l%��>DLbJ�8�mY�@�#��l�^�Zm�6�7�i�Z���~�D�?�g�*�����+˘�tь���{�^Pf�|�Ԇ`�o.����n0h3T�q	�n<��$�������й�5+�#�5Nƕ���=<z���6(���'6�22K7Ў6��d�}��N-��Z�H)3�R��Z4�$pUމ�2ȭc����O�|��t�ύ���'s��S�9$���*��t���\ ��bMH�DիMt;�P
n�)Wޝ�o^R;��M���)Ol~�'+��aw��a�6P�=������W��V���%*c)�����@`��w���`������:	�
+I�좰���6G�I���N)�ǰl흓�־J"83��F�(�����_c</圵]�����¶k�߻�[�&�0��5�Lzʊs_��I�Z*$�� �c�T��K��B�tM}�sH��Z��,5z���|B�DM���s+٠��K�J)�*�s-�m����b������-�@��@*<�=�DU#��NG]T�T�2ϲ�v�z��>n�X$!�)�FԷ�y�IN8h���n��~�Gq�M9/
gO&��wA����W�$�w���zЙU%��+߶���/}k�>O $'���JhFh�E}�a�h�p�������Co���_����x�.���kK;o���r톊�d�y�.���k�2��b��A��w�2Y	����e`cޱ�G����&I=H���8�{��dӳ5�GQ�H�l.�gF��h�jNv��K%s��v�zV����L'�@$�s͠K4!���B_�m,<{�Y�ޖI�T�vM�/9ɭ��d1\���V��T1��O�;E����{�D��[s�5��v�7q���V��^����&U���E�A�xz�y'P?\a �ޭ�
�zFfY��)�Ia����u�Q��R%PpFf�v!vbJ��~E�=]������å���}��;�ռ��9@-�<8j�P��rJ2�ن���-�C����2Ӵ� �5s�:h�k�=�h�%�����v��=�'�g�2MP�-
�W�o�s�+<R졣KV���V�*Υ�0JA�&�ތ�/��Jt�ݶ��e��h׿_��kO��v��y�-h���~k�rN(X�z~ͩ���=1j�����NB�>3)GC�:i��K-��R��IC*���Z�0���1g�V����;jL\b�X$T��fgCY�W%M~��2o4�����z]�f� 5�g9����uOu����F�,����Ω�($WS�d�Y��JA�d`���m�G�1.ԥp��@Is�GhOf��xG'wQ�:��&�~6Ї�_s�����U��X22	�F"�F8��Ϩ��$t�?w�>�����Ue�^�Q�����tJN	��#Q��{H�z�B��~�f�z�Zt}�qx�]Q�Ơv���K\X�-N#�5����'.�2��A1X:�� ������A��{++XTs⎀�g.�z:�����݋���߯ͧo�L�I�Ͷ'"��\�p��B�<(P5�Ѓm<"Bwt~�2��_׍��el�;��ɼ7��]=� Kx�y�\'6e��|���xr����@L(' ��уC|�;�ƓZ���
��j��#ӳ���,Tdל�:~Cj����qND��c�-4���V��-x�|'��;< �ѧ `<�+�UN�m�]q�"�z��ҍ/r��O�|$]�_��
��!ڠ��;��oL�[6�9��W�s8I�sU�{�I鹤�c'���ӡ�(�y|o�7Ę1�$�o�'	����'�ZL����#��Ob���}�S�����n����o��sBX���'JD/].����x:�+T8��re�r����g�׫_I�b�~���Hc�'c� l�)�V>�\�|*�|c����𸀾 ֆ�	��AU#�٭���@A��6�k�6�쥎������G��i���~� ����0DQ���L(R
i�E��B3H"�s`�9�����������We=�h�XB�yw����)��vF�#+ ,C���S�A�H%�v(LB�ٍ��-F����oI+��l�?E�m�v�F �!�	n�Y-�:���a� Sۂ�  �B�	6_�����{u�_~��j(�P]�AɎ�f��~�RY�NNK��y4���"̹ۻvחwދ䊊�*�'�c�� 8��ߟ�;"�|��4��i���0�Qb�Wi�[[b���]B�Ih8���]�E��/��#Y�.N��3�kp��ũiԔt�ZP�88z���`��zɏ#��= �-vj�������ٿ����)�N�4Ù��h�i��������aX2�O���^����]�yt��LG:\���"{ڥ���G����ѺK�S3q��J�H$sOh~��������	�e�(� �5�ڰ�l�$6'x7\� ҼX����X3T��T���������>��L�"*&�р_:����J��嫨+r�~�#�?ߘ͢M��B>��h�P?��&v�R����I8�x�tK׼��-|Yw�RËܩ�f�%<���iK04jS-�ن��m�
�`��y�6uuۃq����E�d-�8��5r
VZ5�<d���}�b�[v�"j�.{�C�yE����8sy��k�L;I?:���oON"B���V�I�nUZ�L��tޖZ1�<K>p�]݄ul5:r�ȴ 	��-�fx�\���Z��&��Lo|�b(�.�j��?k>���^����!������r��]�dO;v�UU�/�m�:�q��J�e:c�P��i5��(J��{�[����r͊/�S��U��$�(=����bJ�/k�o�3�^������H����!��I"���"��|�
�*��c6Q�PZ��Ah(��]/�.�p���m8���vm��PA��d���ǹ�6-s���QH9f�h��}q��3���!Y�BE�W�����YM�o b��R�eP�.�)IW���X~�ā=��MF�ݓ��ݼ�I��JUR�.	����.��&h)��N�2�o��5�fy��1�AJJn1�*hL2�����x���#� 7��:i���@}��T��ă2��7I�s��hHo	 ���N1��
���4��E��&f�KS̗��㫠��r0��\YL���N��n3г,�������		��sT��6���>7&�[{�B[���7F����!m2��(��Zs!���$,�mGv��P)v�m����m�:r�ߝKj2��ҩB�)x�,�!A'���cى�׈s�t8{.��(�8�t��@4P�cp�,i�q{W�N�W��Dc�qiJ�IZ`Gf�Umt]��A5� lю��R�gî  �Ł���P2w�p���S�,��G���@X������s��WR204�Wi1ۊ�����R�7/c�`�w�O$ץ9����%�I�J��ձ�Cj� �U���-0�?ffD���,��:@��U��B���Z��>f?���+ʻz��GU�Ce��~I,���m���2���W�C���
�s�%#�|wW��ab���t͙��c��aLL5^�$�{Z,ֲ��­��(�����A��L!�7��Mv�,�g��22S~���i���Y�p�#��
��i��È����^C8ٍ�Q�.!�)���H0O!5<���7�#W�	'�ʀ�������dbW}����y���Ƴ��ȓ?��5�D@yѳ��L��ȧ���m����Vxz��� d�B	OВ��b���U݆_3s���-�;9V6v[c�\�E��f�jt��p���f����~v�ۍ�b��6��8Nn[p쬈�����/�ݵ��8��Gv�s�N�2E�B�~Ԕ�),+�U��M�|۝^.�`��ҹL�k���4F�i�����PI޸C7���1�ls�>@�-A�@��5��JU�6-y�ОSGLrʱ>l�4bm�W,�!�b�L�l��C��6�����fJ~Tl<̗�*YZ���GR"�W팦��8�|5��I�	�q<�C����'�,l)��/�9T-������0�n1�������I:b�!��Vp�Gѵހ5�pޗ�lf6�&8�jb/�6?b_����W7��x�ݪ"�a�ͩ��-��-���7���],����4"kz���zI�-��l���qAl�B��F#/�������uU�h_�� t_��쾳��Y� .k>*�+���$��m��aq
��-�A2S��"�h��|�v{�lsM��
$J-;r��kc�_�}�5wňiI���IGfś��U�y�X���"�pD���=3�rxv�+� �~j�2"�Aq@���g�~1F��������?C]���h�	����yf��i�5�M��ݱ':;'����� 30ls��⑃~}��4�gz-�Nq�o�^�ɰ�&u��3�kL�+]:O-�3u+% ��3EfD�ʘ�s4^��87P?j^���k��g��� ׮�W����&4����&�0���N���?Ӆ*�=���m �̖�z�bVrZ�ٌ��}���uSO��f����Pp�렢7��9������a�X�r[h��3h*$�����BX��v��
�/��j��h��2�����G��a�<~�B@m�t�5#�Q�1�\q�(2'ER�˲10��'���9��Zj�S� �)���R�	9M����R��_��ڍ��S52��m͐��1��KAP��3V�C��E��к�}bR$ع���<�-�q���F
��D���0�m�1��3޸g 
a��<][9
�Y"b,�y�!���1X��~�����d�1B W����IQI�)lvBZ�E�&Ji�yT�G�7�b�-˗���:X����
B�&q/�]=2^tL��'����z�6��֜h����&8��q4�(�s9����ѝ}'][�Er:����/�\mň������b1�(�"l�3=Z��q`q���1V
��V%���~,�%&�
��
�E�H頦�LX()ch��WZ��ŷ�$Á����Շ-jȃw��f�� ^+{m�Φ!f/��N.߈z�N&eƣK/sYa	ĻH,95�Deȗ.��{�����9þ��~g� I�PD���l�)�P���/�I-��}��屲�l�b	�L�z!8׬h�}p(\/�6��O'�Wh3T��V@a_R`%kPy��-.+�A�hw=2d�T&�[i�MJ��N�e� _*%+������� ������D_J�	����kQq�G�3C픵�>���쭕�	����r�\`>1�;�+æ�h�F���Ip���4=ߣW��_K$��v^{���750~��Q�`��?i�C 	��W�C4�1�zt�/Rv�����
�!|<E�JY3.�j�����#n�\)Wf���#=�ŧ�a#��[�Q�u�4�=�����Tř��P)�%X���֩����}s�.w	�mbs�)��5���lreC�*hO�����|���#ގ[��y,ī��i��x�m���=��i��X����Ja���eH�Ka�T�-�{gc���w]� �ʅ�'�{3�e���	�4��#$&A�j�٬MԿp%�� ����^�p�\Ru�UvAI����-�r�;����(�|��Ҫ6��b�z�W�v�������~�n�|���Xy8p�J�hy���c��ڃ��v�23O�]��&_ƒ�vC�bd���>��Q�g�q����%���ras�,$#����~x���#��\HM�=��K4�`�Y�x6+���,��y�w%ނ���Ζ��g�Ў�ւ�3��%�A��n�߬�Ged��R��;��6~��^���̰�|E���
['����^uh�C2}���tݏ�^A��|��dag�w�3>�K�=fz\Q�2��7dQ����Ƽ���5��vQ�z���+.0A�}���u�Ę.gҦZ�������W:�-�6�V��|�&5ʟ��3�Ĝo���#!侉C������ۦ��.�L�rTu�.tR�pq��L(k��٢����a0����}��듥��kȔ�h�TԜ#���,0l����ߥvHY�e�6آ�%��w���d/�7�ѲiK����v<X�2��L�x�#�*���ع���F5Դ�e;��®��E�F�e���
�1�
�	A#��׍څ8�a�q+��jC)�?8(TN#^#Y����F��D�y�%M
�p�H���<���+y�#
��K��~��۬p�ybՎ��B����9xŽ�1�(Y>���	K]���n���JG�$E�-HN�dҪ��T<U�9�[�׏^�U(ۿ��_�lUq��q�g�Y��a�2kk�mS����c^��_I֡����\��N=��B���jZ�t[y���s�hz�v���V�9�4��{����4���mzD��o��k"�&�	�k9֐��Nh����|�S��*���e��� �?�k�j�O� z����*�_`�\�l��,ܜ���F�k�{���O�J&]����8���]-�0��4귢˴���B���\x1���_���gRZ�=Xr����o8�#��`�����ؿv��i8��<������.�����Y<�$`�m
V�k�Lia�-�C(,<�F������z�9���3)�5�`���B��,Cѫb�H(�4a�c��E�����s��m�,Z�.p�s\�e|���`�O���[/e\��Û~H'���=�Y���]�Fp�Lh��t�	C���r,S�2X��ӳt��v�K��ݨ�A��M�9�4��8v�(�L5?V�{M���8�MK�x&3>��ha�C�8{a� _<�m�G(��%��M*ފ��.�/�u/�/3�a�����.I�k};	���pD�e������? (^n��/�X��`@���>�C��\>Z��A#	Ĳb� )���u���92���$RsiMup�Ms3��`G�0C�	7s?)�oxq�JG���RO �������ŕ�64�u��\�%pa��܂�կY�1�j'�!�n�n'�Lf��$S�*�#���H�8�o���/@J ��>�b��{�?aK;�2�H�����\������4$eÇ-��a$�׭�c�__����䚌G�̒��AKwFnm�󥠒�r�p47FS��vi���\'�}>��/j��W��E��<�r���l҆�	~��&jt���,�/!8�-�p�0�q!��mOwu�i�9�C�dA��B�YWK��`�yY"��t/s+L��`M"~hKx$��J=�������sJ_#B3%��(�zYC��S�+�#k�+�%>��/hJ�� [��Z(3�ײ��K�M��!ol+�wU~�j��dv�We����S��5�b���z���Χ�+��qP?��pq��f�5d>��?^�[H�JA1��8�ރ1�Y�'�{�5�$��d+i��t1����kC5jH��G���_�
o�*��68�(<�Y�ǃ��a=,2���/��+*�E벜?t%�`�t�(�K�Q��=G��w|������z�?&���U�fP����ߏ"��?����k�n�r��w����4�-E.��򻙂fJϒI�7�3#��@u��pbt�7���/�3����%:&<�"���lOb|�GM�=��#��3�K���7���~�����Wo��O�I��M=������I����	%�~+���'���d��Ag�<|�;�<�>�� K_6�7c����<�J12��%w�G��TB��h1A�� *��Qe#�?\]z���j��!�lxR2`�O��/x�g�a��ᾓ��}3���i$4�WW�]nb�.�w����Dꞥ ��O4D�gܵƔU>H��	MF�������"�{P&�>5:�����>Ώ/�
$�T(*����z*���ƙfEL�̋e��Lw�@����q�!�W���5m?�UK��k�
Ry-:K`�Y��q�96
�>�Zo��$��#]A����No"�vm3E�3M^����tl��Ք�� Xv3�����;K�Aj/y�l�@� 0*n�s\Z����K����e���J�x�Y�?��O�w��wM���*��N$��|}k� w��v���?na�,*�M�����G:�V�ΥQ�����ꢃ�,�/y߫G5�x%�=oq�D%*d�L���7���ZMkK��ƞQc�Ծ$�k��6VInM����L�!m�	�f��&1�)aClP>u��ٞ���#/S^�g�F��z�|�����s+4�t�h��/�k�[�X��Gl:���5{�(�)F��� H�skk�jS�m��5
V�ѽ���[�Ь��`�+OMwS�_�%67�5�s4�D����^�`�r�$���2C>��7f�h��9��C�R�~�C]��IeIA�6Wu.� � �r��D���'3��q+i��L�@�?M��rӃj�Cң �����>��ښ@wX���/�眦#�r���j�z��?U��������5��؂m���6HY� zH'5�"�$��?BMm)���Sr�z���FzܹC��~���!���k]?C��~�̇G�'��a�o��G� ��AQz0ܺN�  ��&(�������pA=��3,��$�?���G��qlG�oUg�b�N���Y<Y9=<a�	!C ���,����-͹x�GC�I;�v+�Tu�`�t�p��j,u0 ���,�P��J�w�p(����������ߣ��TM_�SJ���dazh��D�|F���-�@��`��{W)���7>^	�|SC�� 
q>�l��u[��sK�5��3�F��C�]f=�ݑs*���]O���}���֖��i}���六P%��P��*����hxX���QԺ����;��o���^�[aA�5���W�	���f��FC;Q��gbmS��Ό+�$)@�Ҥ׿��!UHn��I��Y���h'�~�ʕ`�8s�h��e�0��`�bF���%Ձ2�kWҘ&s�-��J�V�|�l��.qM[��a��Z5X��!�Ih�T�ø���z��1!�b}��b�1�1���"�������ƍ�.f��z���DX�x��σ�!,���.�zxpzT6�@���o�t����@�O5�Ä���եW�w�JۧLh��s�鵷�Ŭ�n|I�A)TOC�4���_�u��ٯ�U���Ip(`Ѣc���d3��B[q�E}�߹�������*��h�+���*�0��Gʉ����N��u��^�Ԏ��^z�a��^K�h�&��^���kz�(��zsI9D��؅3��_��z�Y�u t0�g�2�Nx�ZD�r�k��CWw��G�gKk��Ug;���}���88�����Y!FׄR�.�>���6�_j���˖�M�q�����,q&˪�0��RJ{L���JS�u"�i�_���qJ�捿���y '$\�yТ��)�ešof"y���7w���|�ߘ��&-��t!�g�|m]�h� ;�-��֪�$S����dR�L����d��v-��U("�ä(ߘ��]�L��}�l'"�� �9�xM����K.�]��Jay�孪������pW|nq����ĪY�����7�+a�t��48|���~��Q�B��A࿘��L^g�n}&��#�ҹT�2!�<�6G� 4)Ŵ9f�E����)�A)�������Ctj1N���x�n4�h$�lH��>޼	p��)�!Z�Ǣ��m��{+�	�m�3��	_��乐�8F�qHo1~�
��~�����޼���ti�7[e������CC���{�r���@~B��;�xG��%fݍTw�l��Yh�Deyȹ>miL��VG��&�6�r�G�X��>�`~�Tq!(��ĕ\��<H=K�P�}���	���-�὎bd��J�v��`�4R��{�4_���2�̰�v�=c�2�����R�+d�g��t5���1�ӬOf�9�l���=]-������e!F�ބ���g����m�i�JwpiO�$'(?{�|�T=�6�q�:ٽ6� _1�o�ZB�Y��Ӿ���i�C,���*�����(��ߢ��w̬W_[l��}HM��U�|�]����Y��`q;��v9�Ee&-~�d�#�x/F7��j�]�����FW:gT~�Mk"A��T"��|+����lIθʞ��/g�e[��,�,��$ù�U���E���S�N���J]['�>\�̢y#L�%8�v���Z�d^lRH�� Ay��UE�J\�`���(�e�E�3��]J��Ebҥ�n�f^?L [qB�K����jvXNr
��vJ�G�Ck6Ш�R�5�YLʝ�$7��`E�GŮ�[�����j��̂0O��Bo�9l�v��B��c۾��ĊN-�Vq�ܞ�Ipv}@-�u�*���wk#������+"�"q���kM��4���E-�+'7�DP��Gn���u����
���X����$1b<��@�u<�a��˷TB��LI������L�yw���Y��b�^bw	�xQ���l�I�3����Z-��9��v��I7���~ �?ZYȵ�f�;��f�����E�9V�h�0��r�4&�v�D"c����K4��妨�%2V�*R*��K�\�u;���C���"�����]� ��]�6����Xv��3��]t�f���z�xX[��_+ ������ܶ����l~�1`�V�6����.��,%�>�ٴ���W�<`�ӗ���~fӪިA��L�ZFc,FT��j� 5��7.����:6?�V�䷷�+��D��:|�l_�+H�qO?>��z��)#(a��8g"�f9��e�ϡ��\��z�a;�������J�pI�K;u��|)�N��J�?���/����;��/�n������)������\�V��㼈H'똼��fZ�Jj|2��PO|��W!�5��W��%Ώ��Y�8K�I���R�~p�ط�-���q;��Re���D<���SI.�2S�������c���.e�`�MAy'+|����/PAٞW��y��4)4<�ȗi�Ա��w���G��T�� 2�Y:�J���m3�D��y�����7>�]?b���;�.�!�giJ��y?��Mڣ�
x��<����t�E��*g nyG�
:XZ��ޑ�a�|��i�h�J�l�b�>����f�]X���K/W��8JOzE��;�T�cK�Mp����4(��C�(T�ك�/,V��.�h��UM�47KX?�:/Q����3�h��6���*��d��{W'�ڷCb��+����3�d��tS�갽q8ͧ��Nd>�́3l]�^�A a���n��D�t�Ȭ�pV~z�p�����A#p�>�S�7u��se>_MnZ<`Ѧ�l�T)L�j2S�����ݧ��{Y��r������~��H���������O�[ا!(i*��MܯӪ�r�t���k�x���C�E��C>�nd/��B�ū]s<�5	IT�^�)�lq6�T�hgx4�uy�t�E�M�'�6�>�^W�#��sbP����\l�c\�,�H%T ��IȂ���٭}DZwg	��R�1���ɖi��h�@����_��[�Ǘ�5^�����A���of��#�=d/�c�K	��;�g�x��"Y;����\5��	%�*���t�v�=�.�yq�[��= �����+񇗈�'j��]���^�"�jsCCշ�<u�Y�L2.�k�_�8����HŶ׼I�K`�b� ��׮�~i�K�t�EdJvSH������3���/*�����0�W3�zy%e���&ԗPFg3uĸ�j`���Q���x��Jn>�d{��z�3�ap�8G&[�tk���6
ܯ����ZWpEU�l�W40'b>�1Ȱ"�%_� ��a(�^b�3L�$̺��ķ@s
�L�iD{A#�zdϷ��)@�
���ሹ�HP`��_�"L���P�:/��:j��R����Y~�ѕ)>-'��ݻ�>�q�޻���}�Un4��F�(ȁ]�7�w�y�&W�;�f�IG��3ɛ�f�4`�.N��tη��u2�����4MF�O����!��5 81E�/��r͋��h�Xew;%/�Z3�t��Kg#��2��cK��=�P��g
�tl�ݤO.{���+��<q�ޡ��!�����3Fn 2(�Kb����"��t)��d�q�<�TSZ�����^0Do�Yb;����(�"�)��PCd�c�����p#HNZ��2�=��Nj}|����%O��}��E��N��#pu�ˡ�o��@�ƃ��vƧ�T��B_Rg�DG;*(�2c�2AC
�s永I��L�����M���P�k�v1
�je��7�S���uU�/Nx#R����}��n��� �U���p���D����KfקE��]N��n8�,��0�0D��� �.�G54��
;Y����J�����⃎=���Gn�vg��[.s��"�d<��9E~�=,ȟ*U�Z&
H���0xj���)hU��þ�?��^}x�B틲+���`DT� v�!�M�o[�.GaCiRi���d�_h���o���� ".��:��q%�!��Q��H3<�+���Pf�Hgo={��ȱS�D=ՙ�I�@�����><�j#�\%a��V����pa"��s�*p��B2b��� tQ�oŻI٠�Z�j�`ܝvl�3�x7-�o^T
e�t�#��W� k0|*7��Q,L�Z UV�=:a�Er6�=�Z�ԉR�V�X�肦�sh���m�1�.��(����]�`�L�s�R#��wT���RI:V����Cs�
^����]���#����
<��J8Z�VX�c�����$�Zn�OSJ�,��<IK��5���Y��9ye�S����&�D*܉�爲p�A��H���1n��ߊ��Q��۰��7�*nk���~�5� N\y�"aҶt����-I�bU`]�)����d6T�ߢ�B��xD��e����N��T�\8P��VQh���<�yPX�A��ˏ�a�f)x�7�$�Pw���n�U�"
��vl�M�P�݅��ݔiP��@,J:"JMeXd ����Y}ן��\� �*��_,B1?:<��O�K��/���|o�_�@��p���*��O�����K3������9��3]@�>�(�*K���m ����cIx��r����~�I�2V������8}D�M�-=-���mzC�|�%]��a�tl�H���j�����E�m[-�R(�2$�)�R�x��Q3�;��-(҃�_Pw�G/��G��O�_'b�Qa�qc�,���cP��N�!8��G-�a�GK3��uU'�)�ø�f4��]4��z*�<�sN��
^��2�J)���~+�B��x��S�5�	�&���<�okR9	�]�}�g��̤�g,�IA�4�>�#����A��!�8�nJvO<�w�
��������J�OR0.� jp��0>j��5̏
k���N�Oƿ��S形e�WBj-���䏾��F�[���亂@�	�n��n�Z�%d���);	nO�T�(�p����[��$q�l�>l�z��~�&E}1�~3#�ra�$��=C�����)�=���Uk �5�{�	��K%�	���S5q�3���}����ӥ ���ͣ+0��&Y1xB�F���^k�����L����V�#ާ{��{\��M�"��m>�@�$&��O=��,x�n��8�X����&�Q���J�+��p���Jy���}y���O�3���5 ������7�F(e~�����Lſ������:b%��|=��+k�-�Ι|�>sz� �fg�R����
�-�+�֗M�R��ͥ6�,�{���hS�~�#�����Tc:˓�����S6��2��h�
�f�J��N\�.�����	Y�v�'����Hk������v:T��3�/�+�ؤ^���U=��GD�WZ8hqd��	���Oǽ��?^nI�7
��c�~tX�iZV0�A�����VN�=��>t�xKr�	���J]���,�� Rj�rHZ�@�(T�F����+�@�����"��"ɕ��^���9	���NT�^�A����=S2���+ȜT�A UngL�FŘ��UQ�'�	w�F�fܖ���l��b�,��ȱ�g?��U�T�h	rA���ѕՉU)F@��=��T��fX�C�����$��v��⫞�P�w��qs3]���Q��}2�锎��wtBJD���l_���pOZJ�F��M�}�7ؿ���G�"��.
���F9�Q���ՏVx�J�0���Rcl��Xi�D�~rM�O"�_X�\1F4����[����L��Y���o��vw�h6Bò_ϯR���ͤdVNo��A��2��x-��G,5��F�T��r��?�od�Q�����*�PIs��Bj��˜��r������p傞�^�{���9 ˄�cQ/a�pX���8F~�oDE�xu �qw��Z1b��?|d��ma�թ0��9�����aw�fckg��%�qw��d�%�k<|��
��,����p�|�`9��
���_�����,`�TFR�V���ۀ3E��j�쯭ܸ�j�8�:���Z��Z�vh��j�Fj1�ɲ�K���4���Cm�u���DOo����W�n�����Ê�1u8{�&�C����D�}�	z78��hgP^�q�`��Dc��Pl�K��U˻ک��rcM�B���m��2�Q�*�9���d����q��+!���ީ��k<}&ѝ��Za&�E�oML\*�xv�E���: %�Էi�M�ɞ��L�أ<�$C�6�B��irR-�
�#�l�"�Z����#��r2��F�"��1~��G�M�)�6y��2ځ�j[�,��t���ٸ�c�;��@\n�k=s�O�G��Ã�V
��'�/\A�ɚ�SO)�{���U@��MM�0RSs6��f�@z��q��]V�������(�;'�BZ��JyT����CՉ�j�S��ۈ��fB�����bk�٦b�@���J{�_y}Wb�j2�8��N�%� *Luvw-@�����m�8�#,m�l�W���n�H��fJ�E��/��a��I�� ����^�U�J��9���O�5�텨<�Ȏ)�� ��V4�������� _&\����l����*��5��c �E1���h_��AǠ�R5�A\}y�T�ǘ�tv�Y��@Y�Z���I}��"@|� 9K��9��/4�%x�|Y�1g4ߟ^x���,��M��OYW�@�y�AǓ�Y�Ow^���n���i.l�X�1g��;�uRtS5�uJ��Z��>ܸ�!M��� �Z��	���\�S0؏C�ڠ8*�Sz����I�Yl�h�+N���pԧ�������gS�&#�5- ���OU�\I
OQ8��9�=��v?��da�����䈊eY!��\z^����G|�0,�-�G)��_��G'(8�m�ҽ�2��{�)]�mm��濉W;-U���flz���8�=�90��mX7SD%��x�*��� �OnD]�:&��=���2�������e[��$}銎��ț���>����
5�r�8�?ws҅˭d��p�N�?���tTc+?8��$ {�x|D<	}EM��!�Д�����' 8�� ��LQ�0X~�
��hC�0��,gI��kl�tm.ݬ����R^�����p�	'�kN��,Ṡ�B���������=?���M�'Ij9���� �2�o�Y�0&/2vm-�^�]kB0 ��Ɩ�slu���5��1�=�p/l����0�59�`�'�ϒ�z�R����R�蘫��{��T�)�1i/:�:ڌ^��:?i�k��ǇN��������D�1oJ޹v�r�D�;mX�b�p��2���؄�y����@�>��=��8#HE�s���x�D�VJ��/0��C�'�{(�E%5�{S6/ �8�?�܊R*O�hYXO�a�~������\�Z�a
���s��s1>w�G�a�u�m���*f���E�)bqrK�D��Y`8��U�o��S-�k��wuȭ��^���I���&i� �����=7�mD8X�w��+$$u��)�}��s��S�Ca� bG������q��y��nutEވ���r���������B��W��M7C����*��q��

����{h DN�/����hS�u�l�C4;_�0cx�*4s����m�=�(�4�
(�ÏE%`<���h;6�d���%��%&�����FK�ʟK�9�,��7η�9\R�Nل`��w����Z��P|uZ�aH��j/�̹1�p�����̕�׌�'�7�w>|����?���Z�߆��Y��s�<'"Bhr(1b�t)���=G߷"�� ����)Zz�^>�C���!�a'[=e���K��L�RV����x�K������St��w��1֭�jR�8b�D++��'_�Y���4�U�H=�������ܙ(��N(,����	uz^��.X ��������AeLh��h��I�0��d����Z�X/���(��Л��u��S����r���yq3r]�E�?��ߖ�
�B2��#u���(P�5q�1���L�ty`��?�Sh`�-U]�����'�O����Hl��S��֊��8h�|6�����y-ߣ���}H��H�Et	9�uGo�]�|9<��z;!`[P�KP�7���ǔ�Z��.������ڤ��J�2P��Y�v)lv�W���U,���C�q� �$��.�h;�� I���	|x�y��znY.u�)���"�23S������'�f�1��M�-�t���\������N6���,��u	#�HGV��"�4'09����.��7h8]_U�'�5;�Lw�9���*��RG�>OLn����K��80Ь�7A�9��y�9����K[W�E5G����!�?5�]y�����eT��'aV2E=E��	�--?�k_�Y��X������G�X�8m�(D��/O�Pͳ��?\�[�ܯ�Yv��Y�T&F{����7�n����t*F��ʱ��w;@a�: O[�͟A�ռM�0�*PT�5�|?��^z�`c��L���y�X�7����{j��[��
�u�E�V��btz>�:���oS8���T��.3�ݲx語 �Sq3�gz�����}����?������uziI�gCev��鈩|��8��a�PY�.�i�]ad�������P�����W˰�Z�J�rl߽�<v�7��#�8q@M���M����������:�S�C�b�vW�n|C@B{�tW����"H"��5[xS8�Ǫ�XWp�p�+�C�-o�b]O������-cvp��]�2ّܩW�[u;��8;�J�/C_N��<�P��-��\�������o݁�/���L��m>dV���%��2́�#��+��G�� ����߸��($��8#K,�
�A��RR�OsțS�d��K��{����ى�.>�>�:he�ݝ:���$b9
���s@�_h���A�����|=ǔ�e�,��Qƫ7</��K<��L�z�~�lR�xW7�����R��#���rH*aਜ਼�=BTo,U��=H�\
���
	ٗ#o�X3��o��� X��ᦸ��~����2��)r�س-��v�-7rH�3�B�Ũ�9Tɧ�R��4.p#[���Q-�3�1)�G8�W㪋���<f�i��š���s�����8���ii2ـ燶W2�nG�[�\���/�G�vA�7�I�NWD�34#��tq;�����A��+P噡n�%��.W����ێ�n���p�/��}U'S��3��dTj����~��@����s��.*kǿ��U��qiFg��m\�~>)��VI��D����\a>]K����!X*�N����A�N���=O���|�&�Xʥ����U��aͽ�v݃?�C{��°	��<��]����7eN�
���0���GΓG��Y�B!��'�,B��H��R�]��$�xN%���Z䛘ϲ�Z���������~��ʚ�U����w�lm�h�;a��7?�+S�|�?�=�W>�YY�b��<,~�8�/�JZzȠ���}/.I�2nfĴM��*���a�@uuW���P�܇p6�w���|j�ȭC����ps���m�ќ�d��1j��F(����5"�z��OG��)�v-�2�Ki�^o@Fj�S@"N����%��Lا2kqWP�řj��5��y#���OC��cUg�6
�y��%��R|�i% �rcIn�G���
��>c�ˠE�|5-����ڥ*_6�*2����P#6��G�C��Е��m��^ևj����l���~���X�G1��U.�<<��J�2���Qhj��AX�� !�� �@5���Y�Ц��i�"�[�QK���	��F߾h�Y��kмhX���yJ9�h��*r*�yD1b *E��{@|O5�p��B����R�VS	�Y'A���
���L�М�KE�O���Q���H.������i�]n�$8��!�m�ƓM �d��%�t�|S������d���d!�P�l8X��pcv�m+ ��V�w�V��m�g�e7�@�>��i����6�ʕ�� j��J��?6�Țd�e��W��RЩ� ���Ұ�mtE�H1�T���=sA
	
���sIb�av�@�����~a�����XL습�ݷ�hTp�~o{�$��m ���j2J
��d���f��D�ȴN�ܩ����%Q�h���2��]�~3��N�������62YW�.b���]��M���sۙHǰ���TG��NW.��������!҇��ĺi4��|� �q�����-�q{M�[6��2@��{���q4,���\�2+Myl<7pT�����}'�怽
ΥS{ś�i9�����}`�������0ds�(��59k�����bz�#S���[�.n�F�!�N ��ǐ������QĻ]��o���R�:�M´���Ok���lB8*������ǳ} c,l�B�Zh����[V�K{�2�p�Y+��+��Wf�A��a0^q���!��S���1|�L��JlW�V�ٖ�L��s�؝�$�%2�9v'ސ��z�[�mO�e=��/ߴ�HM��|�j���e��C���$�ؙ;@��P8��ӊ��Q�9���a �U�PK�5V���@���$����Әss�M�c<D�yQ��ݷVl�\Z�Ӈ�uS15f2�����mDg�� �4��[7p:I��FR�����e���}�l�O��AO�4s�1&" �d� �������y�����yl�@��T�sr�jx^6�D�I~����ݕ���J�3�O.0�؂=q~���q=n�ڙ�#���1w퐡!d.����#�+��K�]Շ����R�����Zw�z�f�z����e�G(��f �ϝ}F́$��ïA��K��}�C���p��|<��v�B_��	=ެ
�Fn��w����
���� ��� ��U8ٞ)��,��y�Iןk�X<_gzC�������rA����"���B#����	�z.o%��w�ЀCjBʱp��I���&ݜ@/����K��A%t��_^���Jn��Ne����$�XL��۸~�8�p�S{�t��t�� e��v�wL�Y1#�@g��AL�6�K%�D����ρ�z���&,qԸ�g�qmR���6q�\7�FI�&`�Ԙ%�ߞ����ij	����C]����9�3���] ��6��y��u3|��s��9�kX�g>�?E�{������n�ŕ�^�-E�X�|���2���:�uC�X,�����a��,чMQ�C��vs��I~=<w�`%��R��;����?��A	�ݒr�'� ��6㯗��	�@l�)�axZ����fo�&��Pl��޿op��%Y$�^�ɵj���%MU6�;�a����ِ�C�A.�J��y)�@L
���J܆�]ȃ�_x�U�>\5-!�����1�t�E�M�,����	J���j��9��z��)�8��n�jѫ��U.�(��k24��e�"��JV��ύZ�q���s��&}��ʲ����@Hi>��A�������n�7�SZ֢�Ov�����zF�X���qHC�շj���w��Fl7�TRL��nJ�Q� �Τ_��EZ��C�YP�bX0!.�*����JZG�m?�Ó��a�;�ԘP�C�l�S52l�G��d:�I�� |}t����)����7�2���� =�*p�і���}Q`���zd  Vˉ�uhjt*�aBr;��և��Fs$ ��C67L5#��,Yl�y����H��3�@�␧]�ҥu���WJ T\�Q�{p�jM���u!�.ⳢK�5�/�H�H.�п���;K�-c>�b�����@pRӐ�E��'�Y͢�&�����͖Sι`���/������7?�Y� ��yᛂ{1�?H!�I����.ПABH�ȇ:�<ָ�e�ˆe�?��k�]�9.�����Qq��!�mue4��>鐓�e
��抦����cx������Q�
-W^�&d�M�(��e�Rշ#QND��#E� ��Y��|�T�m쵸��|�
g4̸�]@'�&Ǭ_�;�qV� ��x�(3�2�X�EZ�;'��x�0a���w�N^��b(���� �x��Gs�d+��j���0c�Kߍv�U����鰩�LUu��������j����?(׬�=:M+�_�l�����+�� ��㙘$�ꎥ-�<�g �|����3�˯t�;��2(EW����EV%�5�����"�_�m�t��s��_|���#�,'�\����M�0ı�����u�<�M{���7���.<N�sd��,R�s�cO��I4��qZ���?;t�]]}�� +S�C�|A>ȟ0v�Ct�ɃA���"��R:��W��G$P��f>ܺ���>Z�)��\9g5�%�x-��(�����Vҝ���hP��U\�6���<i�x�?�Cj5��x��^���ɔ�=>0���!J���3�|��Ѹ��\�����ی����Ϣb�gØk4��(]��+'NM�$!��}��,D-_�,G�o�z�4D�8��G,�5��^:(rPiD�.����ф�V1���`=G�}�0܂]���m�r�6[3��j�vcذ�'���/˹s$�A�0JX�[ȱ��㪠F�����������Ql.��=�\��=�Ӿ����������l��$k�+��a8Cbg]�R���+���F��<���CAlx�d����4H�~�0ti�dk�~���ݖ� U[�k����b70"*9�+�c��@��"/$��5�!�y��7�s+�̓e���l�©)s��>&�4]�*#*Bpx8F�m}8:�+�p�H'�㯩R�t#�.������ǈ�fx�zA�e\�٭����dy��`�?]�}��q���]�v�I4|Y��1��+��ҍR8B55(�� cY7�͗_R��+!H�嘘ݽ�M����/t]a�a��B�����FJ#�۳.��g:B��c/@X�%���F���<��x	�� u^(%�Ғ`#�xL[Q0�Ԯ\��:⌨����̫r���W2(r �ҷ�O�JzD����x��^	�;����Y�+�Zɚ�I}h�s86��/kĐo��*��.�v�H��h�8��Oʢ�<��r�C�o.��4�T��7�lp��4�<­�����`u���� ��؞�/�j��'<��=�H[��¸ʄ�a$��|��jgd�JŮa��B�_�_�m�z�B/�ՐL�W� s�oaf�2"h�����4./e-��2"6�끬f"���~��l�;f���g%�����^E���/6H�J���wE݅��	��g�n�j<���NE5����h�O�`� �l˲KL3�G��|	�;���E�=��2���n�>9\s����КiAX6��t��,��3	o��O�-��VN�h����s���iL���=c�n�*]`Fv���v`��Nz�h~�| 	�2Ȇl'�+}�I0�|Gu���Vۖt`�YU����͘3��6*���C�
�z������tJ]�4 ���h�Tˏ��e//~���PY�d�d�U���O	��L�$o`1G_��� ��_�RK��6�3X$�)QV���cL�b��g!ߊ�Gyv�0K��������L���ˊ��?X/?���L����_�"�L��b���IirE��ɸ��zu\�zVg�5��6(�/e)7MEA��P���iޡ��|��/(�<��H��� �����|���9��Oz�⹁����N��<q��f�d�!�a��>�>�j7�)8�DR�%P�2�.C�P�$U��=���픯+��q��]7�Zq@���g�A1Rh�u��@��V?Im�n���Ԥ�u��o�D�P�^?*[���y	�@|3D#��Hh���R��
���n����rM��s��]'�{�m[�D�C	�`��R%0o]Ew�:�x��Ԯ�����}�p�
UPnU�KLܖP��/�)}8�Ə<#ckݥ5qs�ܭ-�l�}i��*�}Q�.>�%������X����$�!��k����W�Nį�Wş FtK��>%A�PW�Jt)wu�2��+ �B�e���?�r��D͎��@��kg3����rp�|�9��Ei-�j��EH`���1/w����	���#�^ZoY�P�.^>TEI�lщYd\�11�]ߗDp����)��Wɕ�`QR<	������XўZ�rk?c�u��N[��;�JT��r�]Q���^�a�pK�(b8��p��x�kvC+zWx��]�����v�NG;�Y�=Q�<x�)D��I�`$�Υ�[�ē�d�NN���`�A��5_�'�w��.���)L�	����%�����y{��C9`�c���Y��+�o1�@~��A��u��!��X�ʾ	kv�[�����[\�.�p�+�k4��$��Qz�.6��C�{,�?�4�z
oQט��)����$:V��J��_
6�+��[@�-AE�Sl0��� ��FS�_ ���i+3�yɽP<*����^�f�\���'�amA��\&��gب�µp���V�N�;�܁Po��[�t�(�y�ǽƄ"�w���ѽ�G}/g���|�n0�h�i� �e���$�#�7�A�>���/ľ_X�b��R{a&�[���}Ÿ�g����w`�tlJ�Q��F�c��.�?k�ﶝ�!w� `�܃���{(Pr���IM�X�v�'���������[���Ǵ���������,���`y1O���� ��^���dO1��T|�g���h�^Sί�z
$�c���6�Ԣ����͛'�)��!$L�L��]��%Z�U�qDj�C������А�o��5���f{�g�x6���~��S���+.r��v/�q�ES_M&4'�]�>|'�8�ĒB�+[$#l�^�6��X��ZA�Lvź|����#�bF���#���1���:�4އ��hN
e�h1�|{9<7c�)�0"
e���,��?rU�e�\Y�6���)�e���{,������;�%h &Q�"�ŰŴ�8���4v��Dߨ�%tlQ��LX�ǐI�Z�,�Gs��[G`-�d.�v����'��NO��$���_XA����N4���b�t)�X8ظR縛��l�;���S4r�..�)LI���k�Ս���B�/3\�񲸺���5��3�S�|A�ҮP������#��tT%����;~.^[ѹZ���r���`Ӱ���DX���E��z�/�q�x׆.��h>^ �D�v����x]xW���-�,B��S�Y�T_Y� ��~������7���Jcg�w�X(�q�&"S��]�|b�d���
/����E2�hO���D�kR��|�R�g��d��A3{�Zq�0�w�?Ǌ4q��I~�!!��g�C���b0��&�<1o1�����/ȍ��.��ǃ;�� '����ZI���=}&��,��oiR��v�=�s�:���Ј�x�ˠM�����m W�a��1��u5�F����=�bW�,�l��5�d>��e�@�Q2��n��z)��EL��!��U$
���jo��D�\5b~$��Hh�e�!��� (��~v8j�Q�#c�1>#���N�Iq)%R��&J���0tK����r�� P,o�%D	�}a`l-,��ئ<�X�
�+Mb�&�4wm'C�߹Q���c���3�,_�n���a�B��B�Â��q����ꌻ�;��u�������q���ctϽΦ�W�uɘ}�/U�m���R�Mr�Y_��n��*����g~Xl�O��6��ʮ6�!��4~�738��ЗJ��8�^x+��������x�$,��6zv�Ta�:�T㏴>1�gTV�:9��W��D��2؛hwg��S}:���k�� �C1
�
�t?����|�i4�z��OE0'��A��n]4���QӪ�l�ꈌ*�uv��_�+d=S�|ry�i%�%�#𲷒x�V�o�Qj.�g��aE6��#	`E>��'�_��k�x�
K�*�46���>��Y��%���w��Ko�j��pxs���F����8�08���q�!���r�iiZ8����'Y>:\�p��Ph8�v�%U׽M��B�=s��Dj(�i{E��%��a�OP}�<ٝ)�5��*�GZa(̢(g�rN㪶��aS��Ӂ��q�w�m~�H�� �
�!�AK�ʫ��n[��D��;khX�H�N �_��]E7\�}�4�׭���gƝ�Q�"�X�0SI���钟.ď6o�Ñp�EZYx��J��{�T/ �?-{�R��'�������ư���I�����ҔS���oZ��8�p���Յ�xV�y�Ek���B
FR(-��s��Ưr՚���_��
10��l��ĶW��k{8��x�̯Bkk��˔�֐�I���Q+��O(��{ǂ�QD$�K�A�a���P7��r��������E�5k
��/me�|DGw���t�bZ�N�y�C��T
�[Ua�fV)�8�Kd��,=4�IQ*z�bf�H(�/�WR�Vf����q����]����*����L���ѣ��\��fKߴ2
�<�&�����S��+�D�	�BU�I��5�l����'�%h�iOT+��s�`FrF�	"�r�o��/����@�,��'�}-���m�Y$�i�!Ľ��/g�p��R�!9�����"�������*{h����O��:|��eSh2[��p���f[�3�g�b�$p��M_�h��b�8Xe��x�Qtp�w���߰kȌY[7�<��ƵU�\Q����Eim�D��ɏ
���C���}&�������D�T#C�0�عM��f��g�O�,��_B��9�S�\�Њ; |�Z~��pW�)Ɖ���PE�JO:�標�z�jj�B
���HP�S��r��akY1?�@/��� �2,ɉ�ZN��t+k��<�=��H����xE�����v��Q�ﺢ�vu��:7z��_g��g=�J|�aWm{T�����W:��ǳ�9���	���3Ey1@��k4�b9�I�ɚJK�h晀@�ώ�$�$D�'ե�@@�qQ5��|��w�<��(�N�ې�a�pBM�'Yw�������@����ue�	���R{���z¸�u���L��Ⱥ� �@8쥷�v���a4x�K�I�U��x�.X�g�	�s���'|�mH��~��CxV��on1� �x���L��'��3C��pRer�5՚6|���J��E4�=_�8ɛ&F�����い�>a�9�bTx�#(v���%���4$�\�����ZRm��*���D��� �:�#ұ�e��#3k���06��X��!KGxa#"���dMZ��X@'�L/b)^�u��@6]�po�kᰊ�2���?�H��:�5!���h�yk���y�B�<M��k�L&��r<gG{^2�p���� �U��{%��%T6���
$Drc[N]$D&���>'� �4�`�K-�c�>���ҤN̻��6n��k�z&;���A�����eo�X��K�����.��ѢW� �)$)Յ�y)�E���v��k��A����b�%ND$��S�wU��:ちS�-w��=(t��)f~���)��Š�����l*�^�y`���(D(�Ψ޹�H)5�h�6�c��z�y�d���OɥN�-W�K��&t�0*׿���Hy}��/n�ޡ6���0�HB�`#,�_��d�DfؽĿ���A�:�B`���wI�j0���g ����q>:x{Qu�g�N�[&߾#�$0�_U��0�W֒77��Ĳ��"�i���N<#���NE4�G��B�y4���¥d��@�!�q>�'ɳr�j��_P�/dAWT�Q� ��a��8���)�uү ��z������4���`�U��hI"{2�"��5�_����A�$i#VNb	JNzzT8�4��$x����v�nl�.Y=,��-VX  ��f�EN^rd�V6^'4o+��"� �j�ݓv4'|�4��9�"	X��c)�R���ʉ��'�B��K��?���*�WwS0����I�����3����v;j)iTdM�����+�&[�h��CYKo=l�9²7̸[�m�,��'+�o+3BkJ��Ā]]��|'>�ރz+�����?�t�q�+��h�A�������%�pu��r��ڗu[�0Iy���
�=�u+�"�5�M����^N�����4�l҃d@�b���|�S�_6�T�b�t$PX�M��zAŠ5j��S�ɸ��(��ix�N�Ig��S̊7%Y��ʞ;�Z�� {t��BK��>�V��L@)��8�؍��$����$�k2��DV�B�����|:��&E�Z�(�#g�p'%�	�\��j;�pjSx�l�Vb��/<
osH�ȞEW��@��M�QK��0#�4�j�ifv�~!W��<�������@d	F4����40J���PE�^�Y��_=B�K̾6|n��TP͜�e0ɼ�z
�S��<x:&���y�q3�NJ��c��1�A�6.��ʚ����/Vkh(E�m�k��Ey=��ݿ��؏32i�#�V%��y�;��~�$��DXn�ĸlB?]CU������
D�o��F|d�|�Q6���U\�r��X���R[ٰ(�
u�o��2Lj�&�}G/P�ѕfj����f�j�m�"e�O;!x���]Հ��	��f��_55B�eуG����D9x)�������"�Rtr�-#�A�`�E����Vʃ58Ho��a���wY�_��m&'�02�4���3${��ٚ����8�)��Fx֞�Ȟ?<ޯn��0U[|G��Z��"��sCD��j�m�@�5��Z��v'q!��HO�1�P-��C� (�2ޡƶ[ ��Q5��8��M����� Z,0���2xe�O���еbƫBfP���w,�(� F���N!ڨH����TVB=Q�>y�[�(���Z����e�-�$e���#7�Mm1uϋ�}K��7E0|D���e9Dz�zæ�xf���3���H� ��e�ee_��Y��������R_�g{�N���/�ӳ���s6��V�(�N
^�bL������V)l�W<��"`�>N�r i�t
������.�+�zQ�G`F���E��q�~+rrtT�6�2��:�Fe�DtJ�̈́&ָ;C�X�*���F����ԓl����G�B~o��,]Ss���p~�|�;da��7]��������ݹ8F�|9!�2r�6��'x�%��J|x�)�[Y>���2����d�-Rn�@+0�Y55��g2�Cۑ����Μ�S��@j���n��w�|r<g�5_��0�������T�}�"(-��z�}	Iɬ�3���[�ؐ_��%�	�U�l֒��D��r�	�2q�'	�X�"���כv�C�o��r��Ue.��j��4��! �S���6ES�B-��{�k�����`��V.�P��oDZ����v��� �S��l��l���D��!4$F>�/Ц����wP׎��m�� ��d \� S�5|-�e*2������b�
�
0�!ˍO��exR�M�̈́䦰!t���=Lq.��4U|������Y�6��zP������d����baW�Y��wm�-�4�mك\����Z�r]��0��Aɟ����Gu_SJ�����~|C~�»�J��v*]�{�MULc3<$���{ɬԡ����F�u4存o�K�oh̙�RR�����ـ���%
>ˮ���(�t��[���ꪠ�~DMD��
�`0Ԥd�	��<d��3㋑KG���X~���LCP���|G�� B��u_��7N�<�E���Ep�z��H[J&X1��:�~?:;9��\֨i5���k�̨	C�&W�6x�|ۊh��3�]�qC���Ƈp����+w���|�IT�Ӎ�V�_r��\�1�LykR���u����Q�6�-u^��@���b�`�њ<Rf���Ol�Ó���V��#㧷/��k!���(UE�� �E^ηy�R��O�ཡU�m,ڝ���f$������a)֣��^
͘Z�O2Β���7x5U�����4V@0l��*!3��8��D�d>�䣷Uʷ(g��!K/����,��[�b�W��wǯ�ۿR��@dU��c����(8樂	Z>���x�����
h�{����sg�\J9w�n��h���a�z�h^
�� q�D���?��qS���,�2�(�
�n��W��ڀ�����1���*.�ۮ���fP����p(��k��v`�U���u9�Wۼh��h+��p�ߛ�6T�< p����q�1�*�W��]�'"�,�hj�R���9���z��`Ԫ����c�/�Ė�6���۹����<�uY�����4G�G�ħpv8Z�2����*QeWP�o��$�Q�ʏN!9K16��1��sc�R�?alC�
V�����@��Y-{�VR]�����BLZ���l��?Fq�_��q�S`]g��%�j�)� �⮢Z"��5}���5�登zF~�5	�4{n��R��nxPn���ཷT0k���mb+��H�y:sK��f�;��;��V��j��P�>��C_u�]
��m>��������s�q��Z�^�l���
#۱ش\����1�[�D��;+�"�?W�6�	s
=~=&�R��0b�H}fo�<,�\}t$�<w��7	�'�'xke�$�=N�SP�E�[�5�]�{�6���\s.��������,�4W�'��1�2+9��R���6dh�&��<&�HɤU��|����"'/B���`"x^�|���!�"��� ?���
�;�^ϯ�3�7z��$G�e�'���ߥ�ۋc&U�3i/�ǐ+�Pj����)�I������qzd1�z$�{�Lo=��厉U���~�U�j�D�=jօ�5��lZ�(���ѱ�����-2|P�Jv��=�����-^�I��#I�������*����vC�%��y�E��x!'��u�r���4A�
p�st1�n�_�pd���iC�X'₴��4��	�g0E���pz/x�S�$I2ʻ��ƤyX�f���y�ٝ���0���2�ḝ�|2�/�k�OY���*׷-V:i��m�o��Ɉ��!�������H6�����ds�"�w
��g��n��m������b��<t�Y���b!AA�vd��,��}^OCl��3Z�F��#ak�̆g�X�"��|4c�{e��pR��u@۔qd��3�݂:���m6�o ˤA��-���U ��Vit3�7�1h�X�w�}���[�K|�X����N���AVΦzR�z��iv�g%�� �Չ�ޕ�{��J�t��!���X(�iҿ�k.)Ǟ������ؒ)Bh�8ľ�q$��^] �(v�`,8��#,FnZ� �L^��ױixj1���=6�Mx���:�J�C�L�E�(?'a�Cp�GKMoP�������Sc.2���f �Vu ��l��q���V���T��ņ��ރz�O�xf>��Q�����ޫ;k��&�¾�Q��|�O���C9���>���K"��F�C���v듰t�HW�"��vu:+�ihH�g";���a�5�!�I�X�)�V �q��yt!��J .��l�*��p{��3N���ׄd;�*U�`&���;d���פ���O�Y4ǝ�ϭ��m�j�c�%4��O`gNr��62�F~����qC����9?˸��渂�������e��}����:��\tKS�l� �t#�KkB6��	��ek�7��"��K���&�c��M/�鲋G���e=�˰R��#�Ā���d�t,�s�h{�`��� v�<�%���f���\����u8��ϝt|a��ȥ�A�M��c����E��.�h�2�w��kV%I������<b_*e0.���q��z 9�ԢF��(�t�I3�.ۈ�u٭��@��ܕW�7$j����{���X&/�e�mȘ����w*n���Grb��֓n15�?������8���^�Cet���lCI˷øj�H�
�E&�#�hyLY�����#�O�:g�L�����h�ȫ�� �`x���t�sD%�^��b������u|�һ0!�Fy�`R�~�t�˯��g�!��rA@u]I��\w���1Ie������(m���D�f�7�1޹vWq�Ҽ-Y d���+�E�m���:;�YĿ�������6��h#��w��6/�������vFu��r���fm��@��u~���UX�R�K�]�����W�yLHCOn��.�?�Zdh�����IR� 0��jgI�J#�ѐ^�D��1�	D\�*~�u_���):7���9���YLBȊ���Jb���h\�Z,8אj�"�ߎһ��)�@}�����<���A�p6�2�;K��AD�E��S.1�m���^���hx�Hʜ�v6x����@�R.�|�*�%�=F���ӓ�7A�|֖f%,j�=�x�R�ݛg�v|HX��b4��ɚ��v�h�.q��"�\\��y�0�*E0x�-,����'�ҫ�N��"Ҋ�#�n#6�c^&��؊�ȕ m�%*�d�R[��'=�g����ƍ#d�&�]���ruU��ڸ�:P�Z�X0z�����#+�I�b] �#0�C7M;���NIE>��S�]�>ǹ�m�C��B�QoY⤺�8Ln!"�Y99U��]X�"tp!?V��|`�5��Љ�ް������u@���[!ۛ��֣|VJ�z��d�"��(�,M��a�G���Ͱbi��՞"�᠘�`b�m��eiy����I����NM !;���� ��˱��4�k�Ba���n���H�R��	���6��X,����q�XI����1)J|�
Ub?`��c{XL_��G��RT�3_��o[wY�+)���k�2ev�j��u9���o�8?����M���q"~JI���a�֝�J+��v�^�z��ߒV�Y㍲B���p�"�i���_�Tl��Ś��i�E��v�a�F��ā�,��Y�]���N_��e����s�n��@�����pP� X3�[��3�=��@y|R��L�{�*�zn�y��m�/t����^_C\�ƥH�g�[�s�"�)��j����]+-#>�>Et��Б���K�~JST4X����S����݌`����$��Y��!���A�V����K��X�U�˹ж�P�Y[�H��U��o:9�,3$<�՜�L(���m⥙���Q�1H������U���H9�� %��|乫yG�$����A���>a�2��FBk���oQ��G}u�S<J��U[���Yc5�o��l��}�ܜ,��|n��;ݴj;���oY�=�~;�Ԍ�n_bll�k�[�(:��1FE�.����	fW��"�I6�HR�°��Aa7����f'�HX+�7q���"�Q,Ε�.�������<�Q�=�)[-"铲W� Z��+-B~��E:�Z�p��>SzQ���1�ׯ��R�z�"��(>cGޕ��]`�i��4V�{JsD���ϝ]E�gUݖ�B@rn�\�n�������'D���H௏BĎ.�K�P�	�5�*����W�4���X�������K ��@����L�ȫ����5�λ��k�m���/ӆ��O0�7�@}J���_�����}������YNZ����"4�V L�M��$r��0v)�e��N�uß�"�y�sc���K����zkoCnQE%ɜ�h�����V�������]�q��+ag��z� �c2����dY|�<�p���[�GM�N�~ų<�S����9H�b`k�Z0�S^�d�m黫�tQ�)�R��m. .�M7��b�{����'S�1�}r�f�N�:�)9�(X�(�^jjY�;�]"̜?ũ��6�]�0�9'zļl��U3I|��㻖T_��C`#��Xa��Y���@W�dṁ�Y5�`+���L�-?,W��BdǶ3��c��t̉Ϣ!�.E�Lv��wP��f�w�n�(��|� ���fܠS�M�t�|#_����|�#�Y�5�4���& *��(�)Y�T�iC�<r]]C9�����3gā�����Y/;:ΘB5��P���Xd+n�.�y�\�Ct�:;��>�Y1���nHn���*u��4T+3���t�}�����(	ɶr�I�@��\�ԧ8�	2Jv6a�"�<WXGx���Y�d���8�Wc�L$%D���܌���D����%ĸ��<�,��7뮕xB�?z�Q������[��n���m���1���:��Ⳣ<�ֽ$0GC���И�(+��`�L�~�����o�n��1 '�h�b���6�T"�-'�8;.�O8%W�i�����{��q���B��g�1��du���S�����/�H����ІYv)Łl��>'�;T�C���;�f�}�H���LƎ���4���&��u>ZGVl�U���3Q!�|�#4�p]�Rg� %�݃i�+PP��l��b9QI������&7 :���m�zIY��\��8��i�1��B�H6���r㍏�Q5���Xi��9�zl0�Uz��bݭ �i�E ����-5*�a�ܧnSc��jfk,@�����Ҡ���/�5�c�Ĥd<S����0��/�X�>�U���+�*�
}�	�lQ&Qg��~���� �g���>ɓ�a�ڒ��y�j��!�0S	���U*���/����eDy"��0J��Ibo%?������<�Q�t���Ɉ
�6���'�g�@>W䔘-���`�b͕�`�$�-|�?VRkm^{��-.]�p�Z ��u��roĵ��q�1�����0��Z	��׳�-�o $�o} ��S�]�k��
�9�3�����`C�Y�<�W��
��/ΧGY�(�8=��:Y>J�n�sc�)�ā�1&�$�a��z?G�^L��[��-pE��j���M�����sgv@Q��+����B����J�?�\�b��2�S����Y�.���{�O��s��-��JTS_TZr�5�Y��u�ʲqn&F�L�ܹ��X�(������%�?���6�b�nK��Y����'N��!����xsV�ց�c��pҒSp�Z����b�����B����U:ȼ;=�'�,f�fv���H ��Zc��)�#��פ����n���q�;r��pz��ٔf�I+��<��a�f�(A�kٓC�	cڊ ��q`��k��� �d�� ��;J���P�0���,V�\�v5���6�����e�8��M�n,90���gxg&q�بv��r��������r��R��qH��;�k]�G��]�=Ar4X���S� ��1!giQ
���l:�#��B�ݭ�(K�9̭2����F�gE��^�`yaW�Gz  ίŤ���I��!d&w�K$����K��ķ�Q�"J�U)��xִJ��Y�~Y�j�	 �0����8�uw��i��&�(Gռ	ܖ��P�k/�L��jHl����O�F]��x�I��S��ⅼw4��ˋ�-�.�>E��/C��/�>����U��z���u�q�_hc��t�)9��cT��z1 w�L�c�a�����2��tl�띮�_��ɡ#HӺ"[%ץa���b5p.�&�r�m%�P#�t�\�tt
(2�tjGyX_vR���5��q�>��Q�
�sd��1�J����Uot����]�v?�6)V�����nh��ܳ�}6�u�uB":�&ڮ��%y����:��{ZB�T˵y�!:�H�>Ou�A�0F]:�h�����	��y&�!{3��Db
*��<����]��gF0���1w�0��<��,�o#����6�xc�mD�щ�f��Y9���^`#�/]X�c+�{�Xݙ���g���! Ͳ}K�IXRs(�&E�U{PVa����
�$pa��p�J��:?�����w�����?|��ڸ&��iN��f�m�l�ğǤB�j��屳�v���ǋ[��}��j���D��JBz������5�Y��#J��b���Sq7��È�%_�3ʛtdllq2�ٮ�l2'�t~w�贈F�����r�
�1,^ӓ�C�,_s��pO��E��q&��:�S%�˞K�Z�L��#�7���6˭ftC�qr~i��\:���+됸ʍ�!(�����l�J�-À��B�*�Rbl	�����?b�n"n˞��CxYw��� ��A��S6�??�o�cn/��۹Ͼ$#d�E%8F����3���%�yH@�]��균�񍙩_ 2�W�����S.��p.�jW�Z�)�"���t�Վ��$6�ԉE(/�9�7,��*�.M/1��t8#�)��)�j��^�5z7 �_�� ���qeˉ��Rb���Ӥ"}���s�E���.ui�<��yY�z��<GF��p��>ʧ�$����^�I�6��h�u= G ����@J��;K�3��3w�2�s�b�G?P���d�����X�	)�>'�&Ѳ�c$��w��9�^�8�C0u:V����r����*8�ֈ"0�i5?�KSO�TJK�Ms�
�#��,�o�`K"�0O����@�v�d���?�,cWu(��9T!Wk���d�_�Η��a�Y�BS����Ӱր9�	K����I,h�').I��@��w4h��5�uD-M9W�]��!�v�}�.��$��"�9�e�%�7p�)[MP���:���*��0S��E2z ?�lW���1����q��(��IhI7�{6� ֵ�j�No��bh����	h1��«
�S4BO��[�r���0���I(4��x�#̈���V�^I}��X�>e;��������p�JS����(N�/h������+\X���s�a��u�$˦�J�j���B�ݤk�%��d�����z�?tÈ�H�#���,���F"�K@����/�|�4Q���n�5y�o
ݾ��^����4^A9r��3:au�8`6��4@�N��4&P�]���&Ƅ]2��⟊��E�[����h�]_J�.(��ZZ�ևՅm�pi���wC:Ͼ�%�,�d�\�ݷfm;!]K=C޷�2@(�
mI��O�A[r�P�bq��.[���Wk�N?�JC�H��TO�3��	�����Զ�����a&Qq������w�n>�	Қ�(�a�Eż�l���o������'���[����qyޔMQ����o�:a��x�9�����F�
�R�����) )1n�������94�<���Ⱦ�,�Ԓłə�6[������>��yI�4����3)(zy�*g L#�&�#L�r�pnRqV��+�� /^W�8�W�O����_��f:��$�3w%�r
�T�����tkq@ո*Q���;s����^w�2���<�~�T@�;�Z������oi�ly��o8*YȒ����r�e�Kh�����o�76$�4L���h��ѧ��Rs�	�,P��E�I��Lrk.l���., �"	\H�٤,������-��m,�8q�J,vFM���py�i�t��9�tͥ�b�t���լfӗ#>U3���V޷P���8w�h�+Y��nǤ9GX��U��Zd���+]���F��.�6j��Jշ�U�J��B��^�|�F�^
�`����3�Z-&3�l���������4��}'$�P�»}��0��%e��9�3��Mr�ɧHj�m倛�=��^%�se*��c�õ�����k�u�M��"&����C�N�xE�9w���V�ձ\Z;�+�Mz�q��Ζ�v�9��C��T���mi��>���ն�mEd�j���x/��)R��2~�4�ߒɲ!��I0�!�wc��;M���jT�C l��h�䀶[P�yQi-���̨��i�B^V�CI�u��ഒ�L�|�h�'
$�W�SOG����:�d�m�wI�����%1��J��ր�y�N��Լ)cO�s* HzZxA�N4g!�@M���C��<���g?���ag�����f��9�ʦ�3������~碔*J �K��` �H\��[��3����OL�«��&����Ԃ@���&�f��[��%tw��9ҏ���{S���pN0gmm6���fV,+|�.����c`
5u<^V��\?��w��4f|��zώF�Ҍ=%�Q���ZmM+֦�m��b�ߦN.n$��EN��I��_��ufJ�Rl�C3���	h8"��FA8r��?��%���>�����6�\����q,b5�Y6��E�S�!��(L8@wH4I⭣�"����m;'�k}Aà4n�<"�t���V���#����ǧHU���I�%r�O�?��ש��y��HW��{;Y<a*G�7����ۆ$X�z7դ]~�����[W!����2#��|y8��l Go=4����]�u�
"�g��	�$�k�h�޸��;�8��lԔY��Ѷ�I�[�W�@�==��L��~{j~��u�.��g��D��j�
��*/��=	���E��@L�GF�/�Lf��k�<�rH��
s��k?�]����*	�8�:+��\�� �e�㷷k{�j:�Ql5��!�u�!8exw�'S8̏/Id$ �m���^$�@�-�X�n���.%��2�9g˓�Zn�"lܳw�0#S��~o��Xk��y�H
�K�����M�D���-q����%���|�`���')\�+��`;`���$~J�u}��(�ySX���^s'��8޾��i>��b�Qu�֓}���ߝ�A������Xc�QdnGV�O9���W�@�U�Ft�]�-��CfA1�;+��F��]��U Qr7)�D�b���`:'����Y���v4�i���S��R@rZҗ�>���h[�泌�����J1o{�kD�/� krU��_vTR�TC���P2�����_��&�b�hW��TO�ѵX����,�1��N����	��l]v�@/3Ӻ#ȐΜ9�y�D��>[S�}ܭյ{�g2�?Ha�p����{�B���Vje����{o�6bW
�A�6X*�̧_o��C4� �n�#����������l<n;̳x�k��R���3���*��F�EV �X�����$�T���4��+�_�u�1w�ɟ3�Jct��B,��D������oJ*T�°<A�b<r'KO6�W�<�L�m!C6�8p�����	�Y+�j�Ɇ�E����g;j�.�p�������l1���8�RIXPQ�y������3K�U��U?so��$���<�vl�l�"��F�yT۬,�D�������C��@bL�.��N�z9��31����y����j���0�O./y<ߣF�F%[t#~Ͻ¬\�w��h��\���?���=�z�e$A��UY�!�#�원���/��%/���]N%��u�bvxB�Heo{�;�ϕt�WF�{_P���>�(�j������&h�uB��q���#/��W�b*���m���a&-�Dʹ߉�x4i��ʡ����٢�ҙ���	E�� kհ���"����v�/��N�	��{���<��+��}���&c_��U1�V�ǡ#Y���L��E�o���� /&O_b7�8���T2`A p�^�2#�8�D��}�G��Ӏ\�G �����~ϔ���^� �h�f�#?���<�3r8Ig
l2L˞G�M�Fl
C\��O24s黈��tz>�$W�]`�݋�N��JY�o������-^h�B�5];�w�q��M���>����B������O��PN���_�5��_�|/� ��1�&�����k=�=dX��.8�?>tւ5��s�!���t��]yn8��cΐ��r��d��d�5=4��愾a�d�����u9_�o�CmE��t`8�Q�`Yp��QG\�u�r~�m�0$,;��}�W�W~�Z��e	]�ѕ���w6�D,t��r�(�~��H��Ό�pG��NB&��vO�H����p�W�c�uj#��c /%��M����@G�հ��;�����eP+^*[�y2��
���bKI��W��:hPV[���?#i�3k2��Y��-J|���K�v%�����5����w������b ���6�DX�z�6x�2�V����\^�P"�;�2Z�Qܓ�ꝼ�G �t��䝹v.����PuxAv��Ired�+��dRE�Lq;��d��8L�@
�ؒ:��J�M�I}�	q�0L��	���6�D��kC��-�v��ۃU��YŃmtV�`�
�* =���C�?��G��	�-�[S�)1PU*��P�N>��&�bQ>?��l9�����Q_����#3#�jiy��@Iø3��*ٙ��40���˄`���E��H��%J�n�Ƃmg�s��n��d����C^�d(fZ�����n���%��r�V�
����e��V3��$�O�	Ӽ!YP8#��On�6ڔ$����`���1Ch�Dv��i�u�X����-*����P���*ک���'Mu�sh?W�]�c�r�um�O��H��U\B�]��(�������b�pLqJz��l����z����,��l�m\ʈ��B�Ż�)�k�����:]�a��rNVq�����v�U�s�G����}7��q3e��EF�� �S$F�*o�i1pY���:�bA2�����?�O �?/<,��(��0�l���4ّ�`!{����&�?�pVQrR<��3�����d�	�w��b���6y�W�WZ�}[׵,Z.t�5<��=n�E�&nE
�Y�Rz��Y��;.$ۯ�����U��pm�LL�:�N#=w���}�I�i�1:��ӳz�s�I��$�� 
H
-
N�76!c�t����gu�sG���&��@q��|��K�Ia4��V��DQ����eu��`����h鬮�W�)�� U�Q��Y�|�*�Q����KT�rww]hWg`1[S�}-� !�ml��F+��������2�Ebl-b���
��r��h�la��������0ȗ@w>��f�H��o}�J�j0��i�SS��c֣�¾%�Ǧ�����Ѭ��Ʌn�M����cV�2��N-�m(zݪx�qo��y~��U0`5��B��OC���'��XF.ɫI�����{A����<h7!��}ѨLsۣ�:ᇓ���H��:*��!x;u7����*U��E��/����|��䤅Y9��?GÈ'Emi��?����J���K�9�ܷ�hv�Ჲ�'�&Ą}
9$ħ׳��B@Fv�]J"�����.*������ u��>#�"Y����Fq�_��v��j,�h%�al��pPu)�h�FH�tu��N��`��-�-�P6���0h����h!�Ke�'s��[���@=��&���/>M?�j_=�����&QD|z�!*Ԩί�C]�Aj�N�@�46n����95�0����e&����,��Jڈ��O��H�T�+�~3�@?�\Ez��7]��c�1֎_E.��7��	+G��s��{Ko3km���*�Ԋ�%�>2� �Z<z��� �a��}�i$�e-��Jx_��ls�aU���SC7�|�^"���oؓGh*d����AŎ
�N��*R�H
�?�X��)�9�����®��3z��6d������8#�k,��^���CX���`�J����߰
,N(��"��7�uI�W�U�,�,�켏OyyM�[����7�G[n7�Yr���/j>K;�����CJ*|,$�/΅�i�5���)X���0N5�Cw:�X����V&�`0����l���d/�g>�]�)���u��I���w'��/>(�-��Jf�Im&� d�@�`^"[��Wo��]T��P�ON���b	����R�b��u҆�n��J��Ȇ��i4�޻�oz��mm�����G�ӌ`���v�PSZ ٿ�(����2 �j�Z�xf�\e�uN�/к��y������I�3���O^%-�/`�"� ����>h��D@��, @�|�zA�L�i���r��x�&��^�	\��q��:�5qD!g��1A�̲O�<V�&���|��j�#�v��;Y��{�yE� ���ͤM����g1V@�-	R���*�g�n2�Z��v�a��ǘ֡�7U���/jK��)�Xj��z��"��~���G���y���Z0��W����W0KBf�R�/g�	6�WU0��^3��˃�e��
q1�C'_I��>�i�`�o	���2���r�OM�V)��)�c��c�uq bd����)ftN�pspj�������w�/_������}�>�
n���؂��1����ۤ���ܟ�]�9:�7�B�6*<6U8�<�]�A%�~n�e��7p\���FRTj�4���;)�\'=q�\h�����6���F%z�9��Te�O�!B٬ǎE�h/1HtA���6f�^�{�~���aE�La����q��1�X��hԎRF����sѦ��Q�?Tnn�=�.��W�ZP%��zl��
�����S����Z���7Y�Jb��ֱz���`�s_���kᲃ�7l���:�vM��?���3��{9�9�g�� FBi�X[�u�}�g�. ������6�;����43��y��ą��q6)k+:�gXI�:6�����ǣ�DH8�Ȗ�������J�6�t��A�����:���}��T��ϴ��ƨ?We�Lv0�A
3�S���rD����<b`���	�`��ߠ�]_ ����F��xֻ^@(?RA��d�¶ hAt��6���`ӆ�[�D���K?C�����[�d�4�D������� �_�y��(In$e�[K��'-߮�2�~!؅c���"
���2ث}2��(�@,���kA>yj�o߽� �1m���(�!�'��7ilY Ra���SL)#����>�??�"I��%�} ��k(Ot4 ��X�>6��5��Q�;���7��FЊ��q_85�⮣��N��w�0^Z�����="�� Ne��^1�����`xm�NS�O��z�z&�+�(e�2&��8M���Jm�}�/�E��O��;~�C�fe�%�����L�*C��4��fO1b_JBup&,�S��Ԥ&�;M�wz��x|�B-����@�%z����C��^����QF_.!1}n��d����3�C���+�I	�Ś�U|����j�8�>	L�����tH��V�B3�D�`6�e��wve��!�_�/���s�/�@'m�D�dj��X 5H��-���ޠ y0w�fxv�	I�͡�ֽ���P�棋�yv�Pw�AO �5���1>Jk�aD٘2U�\� �[���79O��M���4��w���Δ��t�{��pe��M�<a�t����Q+��ŧ�bV3v���{�s{��j��C�]�}y��6�FU�?�@�u#/Փ& *0d�s
�U�Z���	Z8#�-�uDe�0�׽����{<9HW-���X����K0+	r���h��Jh��!\G���-],*v�W����ن����+f�q:�x$a��Wc`�6:�C�o��!�����Q�\�C3�Ic�����̎�xcIZ�iDm�]�ۊ����)l�z�lgkFW<�いy`�x �}pSd�:�NP3���Y�y�/ΉK1�H#��O�h2��W������`y[�s��W�ޭ=�~8��,�Pz�
�PS�+0ʠ��s�6��9�b��pJ3��C{��.��?BK�s�Ha�:�;Ka�|B�)�nQ��(������FA�𲦫�_G{oq��y\��������9��p��p�t �ӷ�8���zqRp��˾rV��1+���hoխ.]��V�؞�JL�Ӈ�����ݴ$������z�}�h���P9��k8��o�g%�.�&�.�7ކ�aJ�՝Y>�.{�M�@z��8f*��5u�K�E�c�y�2�7�ϋ�-|Ŭ�Ű�:��n̘Sņ��'���8	�s�������Qrm�Q�ݏ���h
m��>��d�"��0E����lx ��`Hl��'�Nsf,����H�����ma��[��k,�����T
7@���j�##ؔ��d�Eރ��8a.��OGRC+Y����� !b���o�!���ϑ�����O��j|t]IS΄#���/wUv~U���f�(��[��]�t��Z��_/���x�iTWxbc��v�c��8ۂ��~P�SRH90��oV�9�s�{�����gP�c�բ�k�d(�U�HD�FJP�����T��o��n�މ�.�֬�N(i����J�67�um��%�'� Mt�\������%�y�=tL2\&ZF�T����t���ݨx`4F�&���Dc���_��`�I����	^��*����+OV��v�o �*D�Le�q2y/k��r������)�kx�^�G� ��9�/�7@����)�Ly} iG8�u��M則�/B-?Fe�7�?l$��#Gx�@����|���!���"�Ѥ��x5�%.!���R�Y�L�gy�fa��"�s}��-"7�]a�E�cF{�YL�0l�� �K���r��Y��"2�}�a;P�3
c*?��!Ǹ�29���T9�5��4�w�j[\�Rt����K:Q4��+Esd���u�<k�}���v�� �g	۔efzB���>bՙSC�uO���6�H/��h�6�Y���ڠ�@EU��t����UNBh�_�z>�n�D�&v�H���k�Q��$���]�g�H9P�@!⫭<��B�j;��7�#4>i�˕郥{�tA+u������L�l�e&�V�Z$��n�&��x��-r��♶�_�N֘v��^��!�8�u;?N������81G�,�fQ/h�:�+I9i�e�V��	��f&�����OW��MNQ@��| T�,�gnzbs�y���a&��%��0fC��^1�M�g�v6<�&|6�L�՗�T�$-�GBG�V�1�����h$��8�n3'>a/#%�쉲�(3��ÝS	����t�n��k�ṕ㑢,�=-I�ęA�6R��Y�z�t`Q��y1��Wn_�a�+ii�ˍS{�$P����?z��QW�?\uu:��k1��ۺ9�~���5�k!5І,&��f���	�+�h�Jj��(�Wȿ�mV�+�U�8v���EE����¾�u�c�;]{}�I�>��w()IԯV��p�>��S%Q8P=P����m�Be"��
b��ʴU�t�؇%�l?�:j<�����s�1c���ͫe�ϪGͯ0F�e84���dO�%���5����4k���DJ�nM�p涿|O�#���T|� !��9�4jץ����;YG�h�0���=�8�P滥:M����U��ƹ�,����e�h���S:����7zy��q��vn�W������`�F5���b;Q�'�t�Ue�ɇ��� n���3�g�x�t��"ٺ]�s��0;x��Up�I�8�����`>�xr|��J��̡=�6��"0N�E�iD4��rԕ�����TX�T �Ç����ʺi��!���}8Ԫ�L]F	�J[�&�d*'�調�b��Jnꈂd�#��!�I���6�� ��/�RR��M'�������5'�۱?t¦맳�8B���1y��CF���ZW%�ew�� �����2'7�|��Q�ޝ��qL�1�l�/��:�4��w`%�I+�k�RYo�b�Ѱ��n�*7p&��BT$i�2pY�j�R��+�)�Ķ�N\�}$N;=�l������څ���G+�o���<ۨn��co\����F����H�����y���Mz�#�/�3;mı4�<`A�DA4`���!���&�k�׊��ІV[�x�b��f�`�.[u�Tt��G/r�L%*[Rl����I��{�c�z�~�a��v�J"�cA�w�ZT+?���E!���'�w �4Cl�_�Bhg���RjCY�@*��?ZIW}c7�pE#.Wh_E��1(��J\�0��j��p���s�El�����;(�&�~���}{5q�AD���KC�D^.���ϗ���Ie	�È����q����0�l��6��4�J���u�UY��HE$�-�ҝ����^�'ж����'�[��}�t*l �d��v����}�i�����a-�4ܴ��� 4�~�t��Υnm}	�oK�@�&�����Z��Tp--���1l3 �j`h���s���.G�l��"_-��Nw�=���IdC���ִ�Q �T5'�5!WU��������1�I@��@�q��`]h��]�n�)'E�d�d?5ʓ��X�zg��i����U��>��o��r��^�jY?C��;Z�\�q5�E#=2�� g�������K�o`ƴ�]���Li�m�o�Sn=o>e��C����f��<Vo"���
�l�鳽D��� �
w �)����f4�P���*g�dfv]�7W"�_TZ	*�i��{`�S^���!P�w'��5�������lD��J���%� b��R�<E�le�x��NO��<7ۧ?�,\�k,-s ��|z�V�"LZ�]UN��=PY��BA�u!i*����.Ͷ9�����m��B�7�!�:�?�����z�����b2��7�?�y���8e7�Q�SPz���eVY�w]�?�UP�L�H����Q��\�`X�[몯dF5c.�/��ӄ����!�U�PU�u�!8è����ǏUϔ��m�A�P�F�9�*S��Р53O�A`9���T]rR�����.2�{��<��%�����$��
y����Z��T|���E���'���YO����[��ɔS���~z�
�WS���>xH�lq���#�)Mq�f{�+ZS��V1�s�.�LX(hW��~L鹇�l�N�z��Y��3�Th,~/���+�O���1��q��}�vQ������rK΃\�S��4�1M����h�|1u��׍�"��.<wn�#�Xf}�p�\޽�*�p��w�?�;a@c��z��ƈ����8�d�g���\��nX���ͬ�/��6�f��N����~Y��[ "<���s*iV|7�M~e�������ʶ���4����^de	٬m�w�-X����ю�[ζ �(���aŬy���ЉvŎD�� A������	��eT���{�Z��H�T�Z&�oLr���ڔh
�E��R"�D�<KlPM�Z�b�t� ��Յ��@��w�t{�(,�hO�\}Ξau۶�e�3����ʄ���5�:i������d$A]Y����_?�ޒp�V�.~0q������]��;�����b��Q����+�P��GVox<����>h(��;A.c��Y�6tcČ�/��{q�1D�G�AA'T��3�bC��U�<d��Y�*���B���0�hB����VU/�Ҕ<�=
��z$Ȃ�m.���M,�G�j�4J�����אa� ٵE���C��wOz����r"�Ul� -@M�ڻ��ȕŀ��צ�霄�����Ŝ�ſ-��<+}C�"��tg~�G���Y�"n��w ���N�h*z��ѫdt�d�y�-���4	>�犹�F�9 �-�I��wqC�oeƸ7��mc��>��BѼmW-�{{^I9�XLac�6�%�e���3��(�$���Kdю� �2NP��Ah`�k=����r�Ə��f��N�=�����<��w@A�G��RS���f;1�/
3Ο�M�� �ۇ�K���Y��f/������GVl�b����V٫�n�Ͼ��p���8��$�5�5���scnH��3��)��~4l`4�F��<���,Së���hIK��ΡIe�f&+�����WFsb�����x�F�r�ݧ�6?��x�~s�'��Ey!��d���֚d�BZ��*�y�A���3T��eƧ&�*�����kEP1�?��	�m5������W/��n��Vx%��h �ӕ�<�pPUX�6�f��7#k��@�����D}�y]��K�1�~��+7h(�C��l�:��fᙱ� �l�07c����ri^�ht�ּC�u�ԅ��]b<˕�H����d�� ���ɗ�k
��H7��;�8��t� q���-?�Ѫ�l�JR�@���d9�8JF�o[(cǠշXT݃�PoT�+�Zě�(�S
�ޡ�����)_�o���	%Zu���^�5��t�[��~!K�:�p}"�ck'�>�R� ���N��Ƴ߃.m-"�uw^y�ޱ�c� �T�M!���+�պYgI���Վ�o>O���{F�b���+4� -��vt�����|�n�"�aV�*0�%P@K�t�� ���1�8�v����'�h�6��'�@���L+��R�=�=���0�ߎV���9��껖���m� �//r�i�W�a��q^�ԍ��d�B��٦������~'�p~�5;_��o�Da�x$�T�V�I���[����/=�2V�7�c��|����1���6u�� w��NPk4+l�'��X@"��<�$.��R��+�l�HK٫CbE�ND0�;c�i ��ةy�Ѽ\	����
~	�E'��u���Ι�X�\���?qw/D)
ZN[�.�Nڍ�Βʎ&� �H$���N�a�����\2`�zg��o�$��Q��x2�rm&���v�9|��cEW[7�ِ}P*�ݶS�Qu{�(�72�}C��XyY�aRtTyڕB������P�}��=4P�H�mğ��v�l�;?�i�O����AQ���Y<]UB��`q![��|ܷ]�r�	����7�L�"M���wk�)�=o����6���]`��ޢ�?�Ӿ���;�	����?U��� �����]�W��*����+����F�B咭�
����.�����VN��D]dk�����x��J
{fI.�*�YҲ��[����x��H�C]z^4����S�*��ci�=�g�bq�#|��J�}�V4�ޱS��$n���8H�����0��� ���N)��g��a�gH�3�i�֟��Z��d�p��AX�ƄF���k��H��7@P�CCes�{���͔S�E܏{mz�j���k�{q/6�4=�>�{��v�g���6���}SUR�PsaX֘��b���gb���vE�o�0��O��c���
�c�Lo}��6Q%"�!��*4e6�[iRXz�^HݭC�X��L]N@�JxM�&?	R2�G�;�|�K3��}������e��1�s("��1Y�?�C0������ˈ(%l�d�q�\�'ބOעdڑ�7=lD��j��z~�����O�$1KH��y�����;ߌm�e�O)I&y3��'1��fJ:߮�ƣ'�zo��&�_C@��>SP*KsF.�	���ګ��d�P��L��{љ=M�6��ۜ#o� %��!�>H�|���_4iQ��t��h����T�x�;7�V�Mb��۸��U����@@�c`A�SUc�ͮCqY֢��.��O1l�?�cA��s���k�p�^�A�(�����zс�����4�zv�UU�B|<_�f�%��e>�T�_ZQXW󫼿|P�s7�R�+�y_o����_ջ�	�J���y;؀��N����X�]��XD��Yt�(n���ozBiul_�~��l\��qh2EHL�G�k���Y����m-۩{ȧ�^����̠E��>��8��k}�{�c�����"����.��k�>��@'U,�Z�M.3��i����}.Cb�r�a_\z�����4o���#��:mCY:Im�`Y������*�)�T����pyB�~|hg�7dmK���v�g�8�[�m�X�$8y��tR�)�5NeeI��s����wO�È2`ҁ�k5�`�vڿ���I�P�~]��m7!Z������Y��/X�v~z�R�P �y��mJ�Vs�r�"r�e!&QA�}1���!�n��=�M�՝%�O���m�D��s	�J�* ���Ɇ�Wt�3k��m�g7�Q��rd�[8tS^@�k��~(�%x�T�:�H)�W�i'5���^�Uۧz��6%@b�֘O(�R��=T.�}H�����ߡK6{p #D%�������RI�HW#;�?��z�֥J����n�E]i�2�!CG�k����x�v`�G$�����6�F�~d����%<���ȁ��%�I�8=b[K
��ݍ^��jb����B�T"���ѳ[�N���X�|���2v�gx��r���y�,�'K����"�[��d�-���}��p��'l^ƛ|/��r�� �j�#j��_��d�E�K�#F+����#�P�ҵ�/�ٟ�ykq��Wc?��*����Y	u�L�@�Z�-��}V��#�wQu��t^P�tU�:��1ʎ�n����.�I#[��axΒk��Yg͌�@�������Q��Β[��,�G۹��s��H�PA2�+�兌@��p�]-@�H�,#����3[��V�����#���>��Tm�*�YY�G�� _��"�y#���W��7e�+}7���l(�	��=0�1vܗد����|yp��(����F�SdO�^�Y?}om�M��UI��B@�5Ch�����U�<x�\e/�)����n}�Qh��(��o��vK\�'�w�,6���-�?��L]�*,�<�l�0��/ጆ�a��?V��	�$�yp�yo�����\�8���)d��'��G�*؁��m���%"��
���g�T��u�%@Y�o>��CƆ�:�@r7���!iS��w�sP�e�����R���S�Bi|a@��=%�'��-�U��x�� pH�}	���ޖ�AcrqL8�|��&y��p%_�����`���n�,��0F���ǮaDmCHb�jy)�	���d'G�R���pIݩ��8T��5'�E@�;�q��`���N٣5��cA��c�ò�����FăaWʿjb�d1S�t]�i���=�H���(d^��g�ė|� �V�A=x2����dh@=&��~*{5v���M-��}�9�V}Gޭ-�{������,Q��R���,�Y��h��W�}E��7�3����
�����F�T�0�6�"j���Q����4�	S����{��\ �QG�x�<���,\-��hx����J4:����	CϤ�"!��s`�����t0rz����P���kY�;�gW|!#���6\ջ����T~�r�Ɗ��|2����1�LW�n��&�c��[$KF^]���H/j��M�Di(~*)�V�������R�x0�E's_lwlN�A��~��n X�V4�
�"h�l��u�>ռV X[K��	��o�A��u��R�̌LG�}8;�D*�Ǚ��1+�h����U}/�@}ھ˪�=n�C�z�T\������(g:�`�����������)��i7E5uU������x�� ��כĭ��s1�B�g�B�Xj��S�t��ǯR8+���ܩ�a�;a&�I�y��rړ�j�j���TG���4�D��ܔ�^G
2�*��һ7�����3�v�����P�(��<Mxx_zz�TUsK���H��[!��!{�]1�����?6�/ݺ9H����gˀ�t����9��Z�$�r	?`�V���^��y$1����0Ԗ��[��#�(+��sg"\;�e(��f36��Ƈz��G��|���DE5JI� YiA�#�#�w���q������'��l�JŜVJk��u����ۃb/6�*Cp�&�k�?'CGZ��1v�(w�%�Ds��i���#��MyyMT�Ú�����h��˓l��`X��\|��m�M�%���^�pK3b=�~����^#�6�Ļ� ����i/m���A�.�ف3C�n#׈%4�c�Ӿz@�E��M�M����C{��'�Dp&'��`�N�a4��S��]�=�o�2LCy��Z� ��z��_ԕ�pAN�+u�Jd[��)5R��pߜ=K�n�JQو-(-�W�j��7�K�9�~�9�P��E�Ӊu���ʸ����Ț�
�7墒5���^݊M��~�}^��	k�V�C0�����ԼA�c8G�!x�]��G�gm������E��+�6^6�Gʽr��w"����p���
'Җ��!�?�'���jވ+jbW�Z�z�By��A���66����R�Yl� �dG3�c�7��n���fC�"�d���O�3�r��=c@U�W@�/�-�P�Q3#|�����QsR�A��!�
�+rABd�u����
f��,=���x&�:0�R��M7�NwT9)/��㫀3ҍޥ.����ߨõ�)���E��>8�<��VB�v��>c�����u)ZcWGhg��!���
�^��wW��wy���p�n��p�}��1��վ~�F�P��zlT���0���#�؁����b;�,"W,d� ��j��lH�
.w<2������H�	y)����� ��� 7{�[��x�3\w+J�iAҴ��|phTC�eX��/�GSϷh�@s���+6�fu�������R�Z�8���P*��%���ZFW�R[�$<"��9�1�ק@���P�D]������	�=�Q�cZL�/�a�n<�4��sdx!F�L;T�|���G�."�v?��L�N���T+v����_6���ô~ �e� ^X/�VoB�ʈ�m�Le~�Q�+@��zdr�"=���܎���R��J��Wج�Iq�wS����T�&4�p`�)��!��*����D���"��'4O( �W����n06��n�����u���n���аz%��A��� �ط���PW3i��3�|��s�(����A�u�q	��rة���3z���I�s�Kt�1���$�a�N@��Q��n�3�<L^�A�` ֔N$��(��ǐ�z�� E�7����!�49#Bn�ߌ�d��R~��"WIL[N�9��7��8#�1����9�ׂ:��	8�aVZ۸dhxѧf˟�U�O�H}:�"�0����B�|��4�����K��0�pK���0u�s�|������On���^�c������`K�F��S�+N�u���$�*n��b������)�m�����.{��b�*6���p�g�@�K�f�};_|k9��yji\t���<�*1�ﮥO+'(8z�?��:ĸXˮ/�����o���,K�����}�d0��`���c�~���{'I:���v}'H6��
�M<��0��W�ؑr�N�g=��Zs�>c�b�'��{<�ׯX	��ی����V(x�"}�,��������=>�0����$��@v!ڿ~)���<�Ěw����t��W���^��JB��~��d㧇���?yv��d1"減I7�M��(������S=�Jm�h>��k��>&�P��Xw{0�g�g��P%���ܤ޴�^�S<�D�7.b������p�w�O�UAl)��E���]��x/k��j�,Ό�	ǜ즊�B��Ed�se[gL�4jqP�tu�]�^�%Bb��;+̒5ן[Ta.dM��g�w��n�£YP�_��r70�+e��+�n̐- ҃�ϠoU@]�v|�/
ԝ@�I��9�;!�2��b
�}����+J"0����~i�z4��G��T�e�NV q�G���ӽ�k�\z��"� JS���������Zd>
u�l�"G?��1����6�|E��~\�#�.G�bώ,�uƑ����c+�_kY��WM�������O�np�h�Яk���x�z*�7� I�
:�| �$qԅZ�S6� �N�FGM~��)�T���XO�b�^<n5�m��L��A���=＆b*�=�p殹�u��1�ܣLx F��X=���Z7#�ls�E��sԞ�)����1�]e��Ԡˆ��vkda��!����4��հ}m)@1}���N3E���k���!�|�2�A���-�ǻ!�'6�86@,����R�0!�6��($Y؄�<�z�ڢ��m @ʄ�N?��m5���E�T�XKE���x��`]c8����i�� _�(]mc�����0w���P�����1�]H����>�K��iV����z�aO�x��"�*D!P�e�y ���7U}�QL7@����Lu%A�@�!���Jc���-?Hs��H�
����a�y����5ѻb���r�~0�~�22��m�k���]CշfM:=v#e�����I=i��S�MA���.ˁ�7NlDk�A��U'��k`���ĵ�*F�SW��Wi���P��>=�B�!��bH'���!ɂ�%�)�%�	V������3H�Q��-w[��ae5K%������년��!��S����l#� �e"b��n��v�O��)K��4.>����(���	�B��������с5 	Ki�4��%���E��{&<i�]�n@���Dh�m3� ��HD` �$�Ȏ�2U�Ą͎Lo9X��}���`�B��<��%Ҙ�4�d��;��lߺ�����
��iM�w�!���b�v�}��ϩy�Up�1���c���mL)�;?4�Un*��m��>�H���q�T�(*��QR�L<n��~��� ��k����wHCCH����J%��*�65��Vq�E�:�g�\��OS.�}��;�B�oݗ�M_n �-ܐN�ZĄ;�((�b���T�.��v���?;���ϗ�g7OE����^��ԡc�s�[鞊��P= S3��WV��n���B�v}�.����;ꖬy%���ݎD�r1�P�U�����f���2�#���iI���T���t��_h�8�vC��p�!�
V,|\�c�Ǎ��&��Q��S��R�/>�p�~����K��=?u�TTX�o��[��j����#8,�ɢr�	��	����q�e��Ԝ#8 �$͐���PQ`�
�p�4=?�N���2O\S<���+�F��M��V��~��nm��g�&�T�槝�C,+9�z�獵��d��S�\� ���G��P94/((-&�u��&�K��h��Ǵ��ٱM�Sf�EY��2؟q2�!X<�L�m`���"&���-��8@<֫u;�b22�4��:�:a�P
"q��c�䄉��B���v8�GT�N�!��Bk�|����@�-s�تS$bWe���?�ڣ�ѹ�o�k����9k0��uJ��j��Aj��Mw����i�(=}�����;[�>�tb�ϯ }	p��10����sp��~zE$�^&����]�,D��ݍ?��f���8��k�M�u��`��Jߋ���(�����Y �T��V���`E{G�z�{l�
�O-�7WGV��m� ��o��Jf�����>��h�%�o���})�����*�����6vG���V�z���7���J&�e-D�w�܀�CS3w%���&�ԍ�������'��(	��2eB^hP�w��{֎�"�ԕ���X�=3�2|��;GJ?|�i�o\�axh�Y1��^���s�rVӡrq"57��k�O�!T�I'Y@���ծf&Q=sk�)`�])��z������I.��%(�b���������n��D�0B8n�5�x�-E8T�k��T���8Ch�^4�pI�>��li$����@�M��M��h~�կ�r ���>R@ X�\��f��`�����G��A���n�d���ʘ��ī���Mc�<�Wb�	��}<>Cd)4�}��#ߍ�Jr�ޫ�k+/�9�H'����U ��4����߇�
�!�jT+v�ْ���� >	Gu*�Ǥ?���y���^�U��k�9��9�����Kv���H�9O��#̇\}_��;��� 4+ 櫩p�u+��NY��b��ԙ��ϽH
e���G�~t0�y𤁸�nW��~,+L��S=��x,K��!�5�U9ࠒ��ͽrYw�qVy��q�!�Nj�79Ӷ�حc�2p�&U���_RL�JST�UΨ������h��s]�WP�0έ�O�A�K�q�1OG�Q%�R3R(���q{���Ѡz�C�RU�� ���p��e���:��ԍ��q����܋75J����5���>q�n�/'���R-�CL���C��qM˓��N�dėad���b�+!x�P!�$7�ez��>[m{| G�е���h��^z���)�Z��١�+6�_�6 4w;ʳ%��͜K}���������X˷��w3n ����/N,�Jxpݥ�����:�j[H�'���N�@,Ӎ/oq����*H�0HD���~�r5�.�\��P��Ts�:�Cˉ��x��b�~Q�C}南W��2k|
�U��ǿ1G �K� ��s�n����H�εv�G4]9�8[\G}���{'�ʌ(U�O!jv|�qc�5�� ˚�"-�#��K�T,l۷Y��*/�Ģփ`#�9Y��lߍh�$�.P[�e�=v���q������j�1����I˴�K�%dr4S��cT_�X<��3t�i�Ɉ�rN��y����;�?\�:4=��9�L������3�� {}��澬|�"����es�{����@ꥺ
	.������[ŵi�$|��7�m&��JF$^6,�i�%��ʢ;{|%h��A��Z ��V�>��?�����|,f��$G \ǾN%i�"@DRD�x�L�3 �xq?鄤~�؄�������|�2���zs��L��f�-T�l��i(���b�M3�#*~��ͧ��Tӣ<V��y���4.�&�����Z�O7OZ��<滙����b��0�I`RqcAϑ�7�KJ�9�V����Ǔ��A:TiXX�6*N4He��'�_0�d<�R�0�j}�.�LO^!)��t{�m��!Z�u4G
6T�R������;
�h��ל���/q���j���g����U}g�1m���hǡ��<���8sWA�z�+D�}�!��yt����nkt���t�/dk����'�����,�srZ
��]��:�,�s�&m��@/2cM�+�YV�?'���/������틍g����n��ǣxo�gC���b�-�8p�R��݀���Ƃ����v\6w���t������i�i�u<N�ِ�/=�w`���QZ���".q��bt���������-�U�=&�@�1a@�XJW4W>����?�ɐ��PF����^�%���l��� ~������&s��"�5���a�%�$o�6�1BEyQ�{�
v�|ҷ\���d�EOkJ䭹j����M"�����h���a�����P�||x��5�>��5���f�ЬT���w�X�P>�ݝN��7E���#A�����/��r�|�baJmb�j5��c�>�u�|X~z��7���-�_���8��0<�x��z�h�*j=-�|[��`�?���4��tS����H�^�O}�CC������L^����t[5v"g~W��r#Kπ酜SՀ`����[��T?�L����Ob�Z~9�^�����e��K�t��{r��UMlM�%/����9v+E������)�����w%��Ϋ#0]��@y���uqk)/K���S�T�(W��"����7�`�lw��0b팼
�e��>p��_�T��#��{EI|i��'`��l4:^�X����~�G#(b�+x�{7��f��a��i�[�s|��V>���P�<�2x+�8M㲜�Եyb���X�D��6�U4�D��2�@T
�w:HhK�R�ˈϏ���9�=��v��!��/@;�7�`1F�n3/�0P�N�W�_��5�Ri]�;,a��1���PEx�*�U�Y�vU�׿�X�V��K�7�1~$=�
�ug�R��OJ��׊��6�<��'��	tAw�}��"� ��3_`X$�M`�>�ȝ�y���<���ɼ��))�,�$l�O������0��+@�D{��V�MZ�HR[Ф$6�M�!x$����7I��(�/A�4���B������?Z@��!���(k��Jj�]�Z�B��Ǥ��>�.p,�zL����"��!b2pf���>�_�lN�����xC�1u����D��qB����:(�=N��[X&�q;A~�`xw~Grwv�l83�c���]�\`y}B�Tpb���؉t���o"qˍ�����ge��&Q���V�JY٤RG��f��D?�p}nfT����U�#���?;�b����r0��w��
�&���ۯ�h������d�.�N�.�$��/6�C_e;�e�So縑#��D^����6v^�03{}�1:��n��/X�XM/q�2���Ce*�`QZޞ�J�N�G�BFk$z�@�t���kRq>�}�&}2r5�:;���]y���f�[��?�����6�#w]kꆚ�<!lp�'g�O�<�>��a��	���u׫���A�����k�A0�qd��m�by�����V��,�RR��he��?�n���$�у//dU��96 q�� ��p��P���6�T��גt���ŰƋd�j�����a��f5P���b��l/�[���+�o+F�,Cp��'�tu�qyc 5�-B�=���.�fv��Թu�u�й\����8tD~o�Dݙ����!&��pE{3�ج �W]k�W�"7��U��LN�S/PT0.i�mM̢�8�Xh⭒�Β4{c��$�v��J��͌쥭}yB���H�Z�xu�1S��1����h��
;5�ml����@Ri%H_�)�1��YK���`�̤��ʠHO�4g�9��V�rr�yZ>��ϓ�����I���V@��`�\?x�R�jK�b��%`�R��O��~��	w�����p� ݡ@��b4����#|![s���*�> �t��X��6����G�d�j��+�'��?ņ5M�^o�:^�T���Ch��X9�kw�X�pP�8DP�/M����}2j���[/\~��8?���o���oȤ�z3m��[�P����Ҏ�eC��mIa�ڱ����I쾱7:t���
�|3?Gf����rk ɮ��
����CPd�����7U=Yљ�_�I8�H� zz(����|��(��R�q
*�!��N�x���iݕ�όe�]��t������-�4�%t��51<�T�*�����^\Ϩ5�X:Fi�|Cn��Ƀ7�H��|1|l�*m�o�P�Z���Y�п�'�[{�& ����O��u�;}� e�^��I�X�,�w��Z'p�J煨�	 .V	)SL�"���^>ߘ�3�¿�	A���N:-z|��#��9g�;��5��\W�*r2<�t���_^����]^yd�eMV=�(x�ThILÐ�V�Яƣ�\ԞjR���]~Fj��Kڕw��az��1֮9�m�M��;�%�������O�CMB���Bo�ѳ��,l�de�g�e )�6{�樵1h�6R+/�v�G镦�C1i7��$�	<�ʉ{ uH!_��p��L��-)fepIt5��z�Ӊ2d�4f3{�!���{^zOc���أ���P-�ĞF��z��&���>�+i�� f^P�H�o�$*I�-�~��H�� *D_Sq}��.6$] )C;e�^Cm��������^A%�-���%�����*��@?�F��P�}�s��"yV��z=���2*J��{3�����`g�[��g���<�z�8��W�������1X�@�Cׇ��ę%2$��$��(��!G�'6����Hq�1�*�ѩ�� � 3��Y�b���Dd��uo��(�R�KP8��
�y��Q�m)>�܁ϵK�.�G-��n^����L�{�$~����xl~��Zt�䭵r%}�,�j��������+6�ck�$A,���ȕ�p|:@��� �wl�DѢ�#^yv~�%������g{��E����ea�s/5g�)KiIlG=��D��	�R�4@	��������K�I[���td��7-V����p��A����|��9+��N�)��5���T�<�9'���n�4��uO���a�9��v6"'&�������q�xIi��.`n��i��66<͹_S[U�7^����E�i�]-������֟"�_1mk��c�Ҕx�7gh��欉��-����}+gƜ�藳��.�����z��y�}��V<�W�&�&l������S]�f��ͯ�?m���ϫ�4Pc�O��%b��U2{0�%��L\u�;F�-.vxc�O�&R�����b_�Q1���Rr��_!�����j-YQZ��,X�m�j#��:�XX�Wlq
��`��3jefJ��o�BUQB��o�NS�Y�q^�J��k�<�|��2`�S��9�������T�("x��t@|D�3�e�����{N�d������
`���9lGJ���Ỳ�
ª���W�"�����C|�tZ$M��|O:zX�x��N$����@
��04�:P;���1��Z;�L ���M��Zi��	�J��ƒ,�7nbz=W3��]�ٔ$z�՝ ��B'1㶏��6R,Wܭ��V向�����j�צ��=Xt�¡b �SKw�ț�*�^ �}�3d2�eUl8�����Ks5���b>�ƾt���/�� e��(.�6ց��`�W '���]}K)'������!£7�B���άk���o�M��:�u���z��<Z�)�>����b(f.ؑ��_��;��b1����l����xw�lX�R��L�K�2����΃��Z�}����p=߀��A �NX��CJ�Ty�̦���a��J�ήDMr-z4{v]��mAE ?���ް�"D�=����H�ՁΓ�Y���Xs�n5��;]�ES��M�ئ
iK�h�M�E�p�Lc�;I������W
��Pܖ��,D�th���� ^:��mx��v�\Rj�0:	��,l��'H! 5ՕA��qE=��L&*��h�J���Ẳ`c��gVW=��
�p��6/��9�0`j��n�8-�is(G`��7-E��T�=z˃&�F-���ڱv���p�@����k�*�Y=i�
�|s1����<�:4��m�֛=ʸ4vXV;TI{�kJ"��e��,�X�}����{����@y�J�uQ�e��p�Q���}*�56ˢ�?�s�;wL��@��)r/���{>YNg�Kr�rK*��c5ɇ3�Z	D�;8��b1虒}�`����g⹫){����Dש����c�S~5ƈ����%)v��R���-+hV^�m�ڇ���y��#�/0�~�Q��. ��"&��� cP�_����������x��v�h@j=���}`��R�}�F��$�\��P0a�B��弇�J�[g�7�d8M�2P�7�_ʓz
��=V����(���>z}�]�0,��mA�?/o��Ĕ�!�w诙v��uG�1��F�!-�9v]��'���:����Bc�r!��*�Cb;'����F~_��44s�ʼl��4��݅v�O�5a">��y�1F]�y��˺כ3�������H�oE_��c�b�w��e�aR�Bv���G6��&���Q^��� :�Ǿ�FR����ĸ%B޻�Zl�6�d�=؂�D�+-��˗�n�=����a��C��l��X�O��f�0k��6O�J!Z��̢�hY=���Η�(�6Q0˔:�\���A��xF��GYu
�=]إ2'�¦P�[
ںD�g9�����P��#���`��LK����g�N��s�۴{J~�����<�p�`�,��u���KK]7d�[A'�x�T]ַ�Ɣ�w?Q��/�qC��k��"=�^݌�ќ�On[���e��s�>��֊��f|���J��;�f9�*����u	����{��tM������&��	��^�aWb2�V��W߿��!�&4�&� ��\�KI�q��BEl�ǉQ"ܮ��-U�IE�8֑�L�����먨J�$�$�V�$ӆ0|��pdؿo�,_0��e����[������$r�\� �'�F��Y�'L�*[�mKG�Bʰr��l���<E���,�5(��K@����:KA���hp��&����ĝ\��I�_%m+�w,2-����Y�����d���2��O�D:
�����x�Z�bٸ��F�g����ZΟTQMG������qTƯ�~I|T� 8xn���V���2 8I��~W>_��D���uڿ0ڿ�M�/Lc�l0kP�^C
��I�͠DuF�U����c� �F�������Y���
��VS���/�4R'�<�<����v�)�r��i���JLU����l�S�EE��K�qq���
K���/����;Y��sb�����ER#0`��qoå����yjJw�cq�E�A�C��x���vX�X�gx�+��2s�>R|~���^��o�b����3��w:�{�+Uh���w�_����<��S۟;�>
�^�Z.+���6��yE;Q�x����#��m� �,�a�-�Z��\�@�@v*Ř�����3�Z�5����"N��TGv�(����7=���,�tb��9}�Ud.K�����9���ok���/���~���4q�q��b>W#l����5y���Ʈ>?{1S@��T[�*��:�l.�b��@�ŢR�f�K��B�\�,J��:6zo�]&W��J5����G/�l��|+h��Z�C@��i���_��Sxפ���|��%b�濤���L����S�о7AbАQ�i�rjz��z-�_q�q��+�H�п��9�>�.uZnGn��O�r�f�Wlr�\��|�u���ۅ ��d�V11L��FGj;?�{g r��2*������0�c喷�����Շ�F5�(�;��X��Q���'�H�H��aL��o62F����g�R���e���~���g���P��։���DrN��CVh�\�
p��m�\l(-�yS��F)HL� ��p�b,��gXy����
�1���"�8馾+B����~ �j:r�[6�Ѧr4��\��-���j�u��蝋Q��H��?��.=�jd�D���*����V�Jf�>�5{I�x�J��8 &[���t��`�6{2Ty�����w!�2EZF��y���φ,��/�>oʳ�
U׈��$8<?�w�b�1�a�����saߒM��٫z1�ӎc]�;��x�tݭ���>C'�ζؼ:)Y~#��Cǰ|�	zZ#�rS��4�4gK
/$��!2��S#Z�[/Fm���T�V��/5�<�e�����TR�o&s� u⿙q�|m���#��Sc����������&��6[�C�b���;�L#>�oe>Q�~�q����ď&-Nt4	b�]��(կ�@���<ˠm��9�q��.X�B��%R��~�4S钄�
@IV4�,d��6�G�}y���>-�Fۆ�9Z��:��3��u/���K�6~t`^�{�-O�^T���h���r�2�3J*�?:����
��2��#�{Y�N�-���Bt�Ew���@�����`��G��<�,r0��b�U)����>��;F*�����"������xa�>�Ɖ[H�������%��7�9Q��=-�Np�Z�7˫�(���ćT������f'��v���n��]���|`8�xmi�<��H�(�~;i|��~�@u����E��B���m��w�:*��Ǯ#j-���#��#��=N�m󮍇��9s��Ӛ�� ������Y0j�o/3�З��Sp;L���5䚰ޤ�a�HR��\Ԧ��;��4�5wϋf�$P�*ő�^ů��`ӕ��5�V��+x�1�Ô���4p@�1/�Y��a�y�u�v��~��F_Mq��=mRpl��ۅ��f`��-����7c����ðuy8r��>���;Q�[���MQ�e�������g���az��9����%Bt�i[���r�e���u΀M;uݜ�"	F�]�+>�.�B������&��iK~�-b�&�A����4���9ƐK�Hy��;�q'�T��5�ɫDP���ف2��W!\�;"�t��?�2�(��~�l���\n1���'���^fO5��}v�_�u��k,x9���3�T:���ݮ��Ȁ1'��v�5VO��ﭜ5~\���*��d� �����itdu�@�>��lCd�+�ٜ�6E<mk����J�4�� 7�/��;��@_�3��7�,��<��7n"1��J���Ek����`u/j��}v��ǫY@<1xcA����FS��2���4�^�1 D�����Q�V���ُB	
K��Y�NBAr�>xMR��e�X�\�t0�Hg��s�h��w=��;Q�r���p��ل��⮘
@��w�d�?�_��G���p&��0�N1^k�"��"^����4ߝU�� �8>響��X��Xn��PJ�T�F�I�R�̉�����M���p�D���9|O;�k�d�9/�����Αm~���� ��F,�	o#8���̈v>vzC2~��t�|u���XF�|�^��Q�tk�pנ�&M�C�~	�V��:l�����j���%.�_��Z���̝y�A��R��5ӷ�����".��t� �=�ق`�l��4�pb��'m����@���$'�=>1�B�q �Mq����e8�p|�T��sp�����"S� Vi>p�ʥ\J��^@S�-���'ٶq�RZ����Z�
<��x����^����i��0��$��D򾣗d��6J]���}*9b�g��-�!@��ʈ(5�<��Kkɮ��j^�^���Q��Jбssa'GhiQ�����~��{�]���t{GP�I`o�ѫE3���HZ��R5`�Z�s���R��]�Ǭ�kFg�Q[������� -^�ǔlFa��2�8�*Vl/C�8�xq.'�>�d�1�Q�:i�]�*Rɂ���A���1�u}[�'�'|��p����a���e���-;��"-�
Z2�sk��qߨ�8��C���[	1!��#|w����qBU�u�� �K?��Qj���\��EZa�Q<�⼫��>��{U�h ɝ���5�d��Wv�-TXC�n�m�خߔ����	���G� T�aGAcbr#qZ���]fzG�Q|��c��pf�M�1�`K)�)@��J|�c���/Z��,��V���d}a��!j�5V�KDgVm�G�CU�u�����u�I��OU�)eYj�0]W˝�W�ʔ����#�U������@���\$#ސ�� ,#��$�I�e�!H)v�����۰��y�<�ًO��ŭE�����|�o��@y�`����K�����쵭[�ͮur-��埈iϷ�(�A���o�̙[����	:�t	�&�9�#�J�K��կn��Q�M2b���@�Ɍ�wk�Vo�-���t}�H 2�u���5�?�ˋ	Un>5{/��nJW�dˋV)vK�����ǖ��]2o#����
7�]�|�L��l�8��cE;b<HR^�����>�r>�H_����g��X�*�[V�XW��)?�""������4�H�	��J ����qĨ���n��F �ڑ�(
lɷ��F�7/�#[��K�)r�<�`���r�طI�4slt63u�yy����{p�qā���7br_N�9jft0�ы^��Zdt��I��>��4�j)�z�����	��eŞ��R��J����,D��r���_m �`���{ֆ�&;�d���K���Kn���h����Z0���P�,���}��͟�B����_�X��$�d�9�[��!��̞yu~hb��u���,I9elL7�E�E\,Gӑ���j����E����)a##W�l��4\��g&U�qE�F><��C��!�����n)��M�K���Һ��Q����Zѝ��&ֵ�@�O�q����C+�a�7���(�+����0����H����f�2(B�$�Đ۩��e�t�tzE�y�>ڸǘ��R����Zw���M��?�*�8�C۴ ;+�8zMG����}]���"������Eˇ'a��
�(ц�wj��3Hڨ�ı#$	$�rn�f[�K�6�\�L��8e��\ա�)��z;݇�o*(W�!�<G��u8���z��H�
��Ūa�����8%U�ņ.X~�z��;����y�0]dA��9�
�p�9�Kf�_�?H��z]�g	|��=E����<>�'�)��K��i�#�R�������>�����UIW�)4N�̋F����Q�A�I��i���$��6ަZͮ�#�.�(pޕ�����(]�P�q�5����Ӭ�Xt?6�ޯs0��/��<L+5G�iM���׆d�?� ql�C���l�D�wPя��A}����Ԭ�!�0y��W�j�1��:�d( ���(�3�t��Q5�p;����ym3��~lU�/l�t-?��/WbAzyy%�Y��.�Ƃ�������� A�@�s���������5�,��t�� ?<�7��t�R$Z^�3��L�7�믃m�3�{��������e�2��w��ψ�i�_��\hO�
����`̤wR�5,^�(�M(P�ٱ�/�l��l��U������Fy��+}�V9�Ǡ��p�a'��0��7�3�w=aPM��2b��f����Vz�b�'�h��	̐���PER�r-,V��X��2�7R�h5?�A��,��j(z���O?�n����v��p�>����;�!�;C�ur2)�*���lxN�@n8}*���.�h�#���w����k�P�p��S�p̬JT���YX4�vn(�"/��f�du��W�Xt�¾�ln%r��?���Y8�d�+�p��׭�6�1i�)*��s X�nT���0�a���iaۘyW��o��?�y=��KJ�0�i�n���~���d�
!#���:V]���"Hr�ji�BG;=-z� �!W.6D��ei��a��c�Rz�/=+��6��$���h��8��K�[�����j�DŇ�R��X����jn�!V A e�O+&Q�$�c��VZ>�۝�� �ʪ�&��[�Om�%Qi3��=�E�bE`)Pax�Qd��P*�9,pͬܜPg<��3Q�
�ՑR��6do�Rd����6{�[W�3�<S�pD���f�q��ze���9��`��k��ܬ��Aa�ָ�F���a.��6�����ݖ����T]Lq�����1_~Y�ᾉ��4f�`�yn���˕`,�Ù��zk�ߺJ��!y�SʲU�bԺ��H�6U��tΐXV�Y4U�Mkd�E{|I����
��(B!�[��4dw>A�H76d�R��S�Q��U��Hh$�f�%�0��f��բ�<�|޽T�_����X�z�(��r����ˌ��������LV߷aƥRx����;���h���Y�'�:hp��s�&�����M@�T���r}��`�i����G��Q�ɀ���x:�)`S�_	T�Z� ���5���ɟeⰎ��1����zdC-��\�*��	��~y�m,@pE)�hݐ#a����n_�����Vv'�q'5J���30u>`9�/��K=����<�|���jra_���r[D���v�]��Qj�s/�l�h%�a��	}\���~+
?.�\%P�S2�\[�dӹ�F�Rᜡ����T�� ���5҂�d_�PY-<X����j�L�^n���#,�Ԣ~xζ�0q�b���3q(�-�V�r�6T�;v�>v�$��<0���؏k��]�O)�b��}��ۖ_+Y���M
mp�6A<��3@�A��źh��ue����1��QB���3
�߬t��m�cv������[�p��*��n/�=c���!�
��v��@� g�<?IX�0A��Z,Pm�=^՚!Y��G0�N�`�b	Tv��6?8��(�#�� ����繘ߒ���E�,;MFm�9ѭ:d��m��/+ş�<�䵓 ��;NE������C��,�z�#��<�jhw �	�TFMX��Q��3q04挷[sR�<	 O�9������,J��e��<�L�87��[�/�ß�@D���S8�����l�C#t�����].w�@��L_�V˿[Dށ�C�y���-?ֈ1�����],]����*:t��:��8紝q�Dj ?��U�J@�H�<������?��D��5�T��"�iT��ZF��%�u5Ib �h��GIN?���؟���[o�vF�q{Ԃ�� T�۴|��Id]�� H��Nkj=̏�YF��͵��?����#�[���$�QE���^��/����A\���t�Og�ŭ54�7L�x�:��5�|�+;%/�XxR/*A�b��Ͽ�
$�3�o!�Y$PV>c���<n�)n���.���q�0��r�c�`�ǻqq���kk6 �4L�������o�����6(h�Q�S��Z���y, n �v�������A��K�rޓR���O�t;cv��L����TԸ��1G��*s�+�ߣZ�������#C����.7�x�t�$�O��{��`	z�f��aR�5�&������Ke�Z?�_�p�&�,������V�oT��h�j�v8«"~�W;�NoYw$R����y��.��X�wj��A�r}Ks�=/#�f���6�b��K�9��X����B*�]	<�7��N=�]��K4���es�W~Y8sj��r>]��R�:-�mU��+��Eo�9*d| (��Q�}����l����=�
Y+rB�R��9z��WjJM��p��Q��|3L>dX��'.��{(xn~eڪ���C^}�{�;�W���	�jZ���nNR�e8�,�z����a��?�� GF���N�4�
��TX��w����3�2`w �4𙸍b�>]���t:c�����5�F��Π��}�E�t|�	��=zK�YƈŪ�ф���졥#V�%~�V��Ɠ� d{E}�A>o�E�5��I������j��]W)�L��TCp��z�����	j�c#������h�q�W�0$���O7VN}V-�F�D����ʤf���xx�j�8�f}M|�0	�W>xk�)��$%K������$2\����wj)N��ę6(����8oP�C�9�(�z�e��6��7r��ž~U� �\ջ�ݕ�!��J$�����a���Ų�,���TД�3��v<�}w]Q�:�<��Q(�G�V�UgB�	Ŷhyd��B:~9��{�G�I��x"e��.i�=7�:.��N�0j!�8Y(���B�/^,���Y�g������d@䯱�L�/�Uo��q_q5��!i�\�f'r�T/b�Hж�F�!�c�*����u��
�tg�(�5Q���5h"$/|z��/���%��_*U�,ac`Be� ��\N��y������)-e�(p���<oX�bT���Pԥ.���"��\a���}��5�(��32�sZ����J%RX���6h+@2u��9��,�U	�m1�1z��,	"��c��DG�!�?5P��`�`����Oc�¨ݿN�Gj����ڱ|*���Mzr�F��el�db�s�EVP�JE��9����Z���T���ĽEѿ�s��o<��i��"�b1�$��k3��;m�����%�@3rݸ�"<duN��&��p���г��p����g���Ɩğ9��0I��Ṫ��4��l�����C*l�����$VEbRF�r���zW!N�v���'vl�o�����KÌ����{Uqe��D��~�^*U�[%4#��猝L]����u�©I4ֻ�[��6�2���H��(�PÔ�z+qԇ��V	�AS)�:'����c �'Ĺz���έ�t錣��{� �g����s4�gk�y�w�j�r�s���JY�[�O��`��<�x~�R�t?�K�� A�ʻ��a_��N�aC�-q�+W>���+�&��ω5��+_��n�WY�;���a@�+8Ks�!�fՉJ�*�)�$�d����B5��x�1qԊ�ͤ���.;��[�8��M��|Oemm�)� �yW�>��6nt8�Uo��4�����7�*Ɉ�/Iŕ.�<��:xS��7��%NW�"	�[9'{5q�2/��EdG�L�����\�����^�B3#�]ʛ(J/i�}4@�F%�pB]�R�F�P7����)k��;�,�4�����]i��b��CQ7:,��;�S6�dq��� �t�
�j�BL��3u��/}���3f��l��A�*6�"���#�����dVS7�V:���f%�mcX��p6�z�y�暓J����:�l��b̷�X�\��p8���5+�8��i�P�X&n����Q]S�?2&�YɆ�+�Aw�y��Ӂ8�&S�Z���v�A��wq��*;�z��e�3���4b?��N��ީ�������縡`52M��<�������g��>���5�z�L=�|ѐ�����I�J�`��gQ�������%Gn�"]~�-~ �Td�������/av��W������c�F	8ƫ��+ѝbwݬtg~��ұ��,}*��ys�H	qt������������v�����+�MI\?��t���;���6��n̔�ߕ�����ne&\�4ʌ%E1;�[
:��bZ���*~�EΚ_
�{!�w8�<1���.�A�����e�����,@*1B�����S�k���d1�>Y�x�9L����g��7 �4���DY��:�#�0灊`��&v%��S�$�(c�XSꈛ����|���3��ܖy���K�r ݝsO�����㵧�r��:��`"g�����t��A��Z����Z�mXX�VM��Q�w
G��o��X�G�ST*d�Oz�LiTx^� �Kl��ā@fs��MwL����7��K㚝��^�:�0i�_�)��Չ���T�Y�(T������押�1�>,���`ݭ޻=�-�����p&)�J�o��Z�0�^7��RA\�Kv7��x�'n)뱮�5�Ȯ�ԗ�_��CO���d�n���{�PE$t
ᔱyY�QD�D���bf�j��?o�jײ�~*I������s�C�P�����W��Wv�Ҋc�-�z�z��[�s�);?,ᐠ�mu�x������u1/�/W�zW���Q���b�O
64j�M�5�C�Ii�dQ����|�6̡YO���O+�z� V�i��N_w^}bYC�����@��๙�O���e���Ƙ�*&��M5*�aذ�H,u^��=�s���(�e��;���s�.Y�+�%*)Ns�����jm߫�-d�v��� ௓2:�%��J� �j���Ƅn\��V�?�׏*��&>!��^q�hs�Kt�3j=�|x-�}�M���T� �\�ӽ��OO�HgW*�||����:�qYE���-��i��niA�Й�h��P5�;<�x:�R��y��k��~�2��Z!�Z���+�ġ�Y�>^*���xњn�}$kh�_� m�2��`��/�����|����������ܘɍ�d4�!4Ac#�����|����2���@f�����|O$@0b�Agl"f@��6z�xov1
�$	��	�c����^X�#�w�s�w���vF���ϭ�9�/��e˝�}�?r͋�_;i|欵�a"{�!�Zx��b�z��/{Xjz\My~]���g�7�y�,Hrk�Kd�:ҋ�v���X����)h1�\��Q�d���܀��,�:�C�"�+����Z���A�[���ɇ���d o0_Zd܇�g�(9��<��"/k1-3��ت?O#����v��r�W�R/j�������-y���� /�jj����ʲS��.y�s�Fc.P��H�He��m�1�9�������@���W��i��m$ퟁ���ю({�\;��\]Ln��1d�DO�rQ�R���O�bJ��2�m!�G��B8�����dm���U��EӼ�+�|u��Ȉ$�e��y�U�˟ܔ���]F9���KM#	 1b�V�!��*��7�<�gA�16.�hb��K㓶�y�ь^X�Ҏ���.g��]�.��pwfOO=�o����0|��m��%/��cZc�m&C�g��TX�ɍ�p��~�A5��U=Ad�*��,�����`�[����vY!���V=Z�
/j�	�$�<��V��@�$t2�F��J�lf�EWh�g�.[��Hoط�s��@_Au�B`�De2Ԥ��]�l-&��wZ�����3XǦ�s���m�=��Ox��B�����g���%�q�҃��{��*?��k����� W�Њ&�B�;�MC���T�ڏ5���I�d�w�'� ��߅���z/�?���[�T�u����U�����A����^.�g	?X}1y$r�I|f������Ğ\�3�L�����'���~�f�¤&��~ۦ_�K:nkZ�e�W�����D��P�}�⣷�˼��5��mi[��{f���,e%��-	�dF�y*mDA�k��Z��Q=�d�n�{[H����]��^�a�	���۔�ﰍ���l>�b�`�7��G�=�p!R��P�oj��0,�g`��U���v�2DZ)p�~"��Aǁ	�����x�+��E��bw����ԃ"Q�B
�d��t�2۟�����F#��s�>������K\�ۧ����ҷ�ѕ��H+���G�ټ�h�^v���%�綕[j`��n�4�I|�F���������y�*�r[25��v�,~n���LX�Z�J��{������+�aF;fY����sr�*��Y�W��2�~�V��F*��w��{�~#�'�o�	���6F��rD�	~�,�H��Z\(��!k"��c5&J�L8�Ί�i̧P�U-�V:^��^`b����^��Hs��[-;ܯ�p��#��hR�zR�nk���Qd%Vj=!{� �)1NL�7�W�����B&�����+�N���R�K�{�Q->��V��[=�$X�ߪ0�w:&�����KJ:p��&�ϵ!(u�'?�VF�V*��g82o'Omɯ��nCVSo������FA�G:F���d�2c;f�Z����F�������'2�N4A"�5h��#M�n%���6a��P�0=���+�Ģ������Ө���'nP�D<ɷ��B���nd�I�;���N�ah?\� �������$�*�іNQae�*������H���^ugq���������̢;T�<Z��5x�/y�[\V��e^��o���E�v��Z	��q�WVs�w¿R��F���c[����������)'��������2�y���F?X~����U�s��'�ȠEj}�'.��[{lJ%���X�T>����|RHk�� -f����}W֑�)#	ۍNP�j\	 (|��9��5(�U�����S�kPjl�}Fc�zǜ+�������0S���܌��M|�Ig9t�Y��_|�������U��/��|����E�.M��W	�Mg�'ڐ1v��J��-nV�j_[bfR7d��D���R4F���䇱�,��[��oKk�<V��Q7$��X@��z:ƙQ	� G�0^cp"�T��_.�G��ό���£	=���F+��!l�+����C�r6��2����usDu���f�=��#0���-�9E�9�L��J�{��"�^��.�>�s�ם���FK
.&/8I=\�X #/��g3�@#����0�FA���' �z���L5�����c���X��	����͚�u�U�d2(�j��&y�3�*ZW�Ksk)�J�RqYS��̽�����j���O��[k����T�mtr�=����F��q��v�:?���j^��5ؾ\�Wg��s��"��q����x�P2��֟-?�2�ˉ:3\rW+�Qd�Oԁ�h���V
�
 }����*M����t8��e=神���l�!��˷<F�};���?2K�m���k��<�3�O[AɻB��5��>	�|Oq�Nu��=!��Y����-g�:�r	o,6��`����)�OI�,:��뢗%[��C��֕9_���<�*Z��,��Y;� ��SQ�X�0vI:6�5�I�e��P�����,�H���,�I��&���kt�����4,��ɡ��=p�g�֊�H���b	n���&�R��/�-z߶���K �#��ZM�^��4?_��k]�$&�� �N����o���2��JQ�%�8SW��nir����N#5,���_�0)94�,��:� ��O��(.����!�]N��1�w���+d�/����ᛒI-���W,RB�>����YuJ�Ei���i>�+�F$8��ZpT���늓j��2��M����B/B���M��Z8NX�|Qf\H������x&h��m~7���E7L�%���?�Y%� ��Ϭ*�x�D��Q\�(u����1׫uv��@fy�ә���2Ī}�!�i����IjU��
�T'ê���/E�<�dN���7� Û�Đ{����Hzv�L�aH��`�*��̦�u*�I��=.r�ƅ�Q�,U�W]��ΰ���A�#��U�LO����ؽ`!k-�q�<Pc�5�B�識WY�VovSbk����4���� ̀#��Pv�J]z���`�<!�\eN�i@����*Dt5S#�E8�f� )������홤��Z� �U4��"��1�GQ��Y��KV%��x�M�q/
'vM��~�~�F�C�R�7P٤�.����s�Wz&�t݁�	ݑ�����v-�a����ȧ�� ����%��B���\�+�@�I�BZs��?�f���������nw�����֪����A ���+�A�[���J,A�5Σ�y������g��S�u��?�8Ucb��,��{5q�gf������1�QA��o�Ђ$�N˜��a�����xS6Ҳ@|�ڜ��<�OTϡo�}�>96z���,�3/����-ʮ4��3��:����G����s�*Cj�X���}���}�@�M���T�-���_ښ�����X=����H�������[ma��L6m��j��g/A O�����=��:�^�2��4=�M�ϮeZ>4l���0�g�1=�&5=z��� {�g�3	�Γ��
�
��F ­���k�����XIP���@�A~��Q�To���⢈Ŝ�vG��Hv�j�9�m��9��1��-Vcu$����4�\�Ao���b�#m��Ҋ�,�$�r���_rb���퓅]�l��6gAD�󤖨 }��lϐ�3Y*koq�k�Bw٬(�ҝƥ\D��p������	��dp��Hw��T4�U�{�3�wn�Ѵ��}3\vDP�d�S4>W�ۓ��H4Zl|�+X�2�E��$� g8
�*�ە�J1�	ӨW0�:�o�:N�hnư�!��o�(tXi��~zrp�[�9ې*i�(�ih��I��,e�vp�T�Mb�Y%ZD+B�Q��-��ː��h߇H�l�1�e�Vk�����@���v�L�\_�kB�W��&>��f�8 ���%�=����#�d��I �:^�lI�9�<X&��$�8B�|S�Y�*������	�@�0��^���Ŋ"B0¡~n�������Hw���ϓ}�Є�cF�rи�o�#[��>k���2a�1+&h7�:�t��\c��v�hY~����7���"a�#���&����n�9�[�+�bb����!W�x����f��vIV����w{hs
��X1V��1�$H��a��.���h��9�>C;,��N����͒?x �Jf)�ސc��u��.X:L��|�:�u���+7�P�u�FakC�Ո��;wL��"zZ�9��*KM�0kQ�Ti�k�$��E#�ظ�E��* �ܥ�$�����U��Óg��9WX��K�p���'��.�̽u8�+�����r��~OU¿LK'��ZI�Ub�Dud���>�E`�Q���r1��CO�ب��#G�l�\+l����5�ݝ�A��9�wln��v ���	m�>R.t�	R}��&�6ԂG#�U��ܗ���(x�ީ�"���%�@o�ȅl���ӈ9q{0?��s"�*��|z.�{�{���{K>��$u>�>y��"���9��jH"^a,%��aԎ@Ҋ�Q�|Ã��/��{!X\�B��X����q������%6�R�tĺ�Q-���@��)(����*-"�3[����X��4�2*g{?r�w5UЎ{!�7����t�5m� �����e^��7��B�;��3����ZtT�r����N�[|�>�S��l���Cp0�D"�c�ɡ��C���Pav��Zf�x�y�Q���#��mٗ�y<��$�ƅ5.�4�����c�[�pq���aԺe6G�Χ�
�;���b��v����)[X���\��	���K�em�A�:NÂ[�0�zL�Sz�����	�I�"��p��#8S�p��\��<��_?{����!�=�魉���$ը�&$�����
HY�y�1�a�_5,��#�iJ�+�A��ri���f�)�b�LY>�����xb`���)����{(��5"ig(O��:���ެ�-pD�@w���I��ЗD��	:^�����m��-�*�	�lL�&b���J`ˍf����A�L
>��pj�m/��T�X30�@:l��b�Q�r���P�b�d���ZO�bخ��M�;�4F�>��ZCmr�+I(���ܮ�7Z�-t���ȅ�D�/ <��bkm�rf�I�)5鶔�Ǻ�O�-\/���dqI�Z| �ū����W
��o�����O#0�@��B���[^'�F1I��/s�[5��_$�m�d�� 7c_��Z�&`�n��u�Nvw�g!5�1�0F�������<�ҔKC��Ӯ��;��,[�.�3i��]1�q� �=���׃#��[��0ӗ_C�I䛇�w�/g�PQ�.��wAT�~V��h͖ΦyRs���Fҕ֦�\ejk�`-[�XIǣ��B�����K���&q�A��Iʞ���)�h<[A^�ŜlΒ��?��Z�_�֢+�
A��vy�,B�|"�\��V�;n���f��͓����8��Go����-қ�yAq=�\!M(�HprN~뭄�a5�ۜ%N)�=Z�������kڰ�i.ȅ����H�h+'�;�͎�@$U-�$�[w��A֦Z�hVa:[��G�e�F���{�Nɯ�Itp������c�D9~�t,|*3�\ t�}q|��rD�f�~!2�����KoE��N*p�&��;�)f���R������ف�smF���p���S�nW��y[���"ǮySX`�M14�M�l�g���b29��n�%�q*�m@����6#�����I�B�q(��8��
������U�u�K���r�y�3P�	Z�M�_���&��.r<���x��)�Kt�G��a8":	��wp� %�cf��4��/��^y�	-1��}�˃�j�ӂs;�M�Xy$�&�I��7�V�;�bGM�> C�T�Ql������P�,�)Cc3.�Cn�0G�������/N�����aq �b�.��[:ܼ*�J;n9�]X	�Ѫ�2�.���t�C�\���Qp��O]ݻsBL?�
r�������?*bm��myȖ��;h����\a�x^�@4�]/����'�;"�;�������@iQۉ˧�l���m�'�_gw��S��tF\�*����y� �����Z��B��#02`��H���l��F��B-�
���¡nRa0��U�Z1$7Ω�Byb{ܓ8��{���z4��i�K�-��HJ�J����k�Df�%��q�6�?�VZ(�o�~h=c�����述s�|fڼ�3i��qw����>B�D$�`��W�<VZ#u�����/���/o� ����e�<u0�<w�%l�����P���\cn6'=**���g�l�u��)�&���M��q����}-�d'�Ko�&�oaP������[M�tW�B�r@�۰3<WuӸ���ރ���T�#��d�g>�_�]��;ZB��E&=��j�X%�
I��	���c��\lŊ�Y�%�$�\����KA	D �A^A��C��\�y�"�������{�U�V��f�rI�-�?���}�#+h@�S
�i��퍆��?t��߮זY*�A����@c�E�����)>&�{5+wTԙ��	X0�~n|�;�/H������!�?4Y�ϕ��i�6�#��k���7d�������Se�{��y�Z��r]�����H])�[b����
m-n ����ۣ�`_3��,_+v����	��/[[�_k�eލ��[�Y�@H]Kl�DCT`z4� )�u�4^k" ���#�nu�Xq��o�r��?�6�Q�d�͓Yx	�)N�1�������+�6��>��r�I�՟J���6Q�<n���-�q5�k�ElVf��C�,2�mֽN��ĸ\�:���_�G� ���|%�N�5�?TLf���R��k�Ho��;3���V�����OY%�AA�8�'�� �ȁ�l�@X.�/�������x����b�hep,��e��W�*�"(2
ħw#��1W��ZF��B�J���!��:t}u5t$�"���`T�5M.
��!Q�����B!�m�����Sa��{Wp
�5󕏂Oe2��9�����$�l%M���U�:�9����ھl�����Y�k<'�#���M�*�}�Xי�I�����)���wX���;�\�0�X�������ǣ�G�)W��p���L��	��U���"���u������{�*�_6g����u����ް�J�fԖ��2�*k����jp���(��C�9}�^��m��"���M�	�/A�Mx^��1��S��HƬ4�(�$v��M~H���ln���?�{�f��qH�k����_�;e�g��^3N�1B�ťt;~�jeU�ݖ���{����� ?���5��eKP��R�����9�l�\tG侱\�d��5/��t���Ĉ��(��:��}4�X�@�J��.�N�J�u�Ow�ͺ#H�˪᫒�If?��ƤyV*��A@�ҵ�\nʰ���G��3�:z4�,����q�m�?C�c$բ8̨U���)���2@�r�`�R3;!���,r��=Q�KC�	�|�����81р紆�y�0d&o]�QH�e,/֢��s�f�ުٝʽ�=��h��<����{�D%��@؜R�M_���pc��V�E�ʣ*����So>D5�A������Z� ��[>�����&0�p��]5��7t�[���z��@� ��S�A�AهF!��8y�n3T����W'�^2�W��:�l}�w�,���S�N�����~�S���ܐg!�IL4��v�,g4��d�����·L��(�tB}�[�v� � �ɾ��������Z:z��HH��)3F'�5Ŏ�jj���>-~����)jߚ��i�xY�.%^\.k���9��ȓ��q5��d�����p��K��ϑ$#lx�(��C�t��pPJ�1����ܫR�����s���-)X;a��t���o�
6K�#1b�2f��o�͟���݁�U�v�g���8b����D�2�|L1|�cud����6��de��X+r�K���l�"CP#�g�X���i�yW����X�]4^��ܲ�$����d��C<�J�H(�+��c/\�%DĦ��[�SB9}�2�]�L�D�E����j�X�aFS-E�|��XǶH�Pǃ��9��.D^���d��.7��&>o�9.{����w򬚡���.�ǲl�?����M��hS�:�uV������^���o���M�6��8qi�Q-��S��L��͒���!��n
��|ie.��^<o� �֣����b��~p�~k>L�?ymc꧖�1'jg����t��ȁB/�5��P��F�4��[@�3忨�Kϙ���"�p�������n
^^�������itlL>Ex}_�@1;�5]��Ǎ�b��j�W�TKt#<-�W���e��$U@��-��T�����}+?�ʒl����X�Z��md�$V�ߎ&CM1ò����R�Ĵ��_��C�bt�ro
.�Ӿ͙�
p�����q)}�B�AyK�=B���0M����Kl�~�p͡~�?�^$�0Л/i��g�2S���"D�:S������W[�\$K��L<�� i�ԻY�J�pM��1����κ/�r�����W�sM�0>fش$�7��U�:洗=���r2^1�i���T^���r���n��w:{c���'�z�ǌ~�_�1���T+?l/����)�����-�&�����m����=C�a|��yDz{Ժ�a�'�56�瘾��{I���c���'f��[l2S�n��(�a�|cJd� K�����xk� A��6oa�Z���3�&�"���q�w�`
�M��8�$�B�{���
(���Xy�P��iW��@iΥtے��~:'��-ȗE�;�&�2�q�|!��O��겴��΍��(;�y���ګ�'�@�����Tij�m��
;��l���k���0"4�+d���ۖsF��+a��;��2��}P��P�)E4j�il�M���Y�ܫ�x�|5��ca�qsN����Ѯ����9+e����tK� ��C��5g�R5sq'�����;�z�Y�>)���&��v���0�q+�7�hDLQe�" ;pW�-dT���z,�L�c4��l�S��_�gQ�3}��}v7Ǟk�u��'��z�G-�)Sh�v�g��� �̄K�Z敜�{T+���p���,
?��WҰԭ<P{I�r`sd�ܛao����i��2��Wzq���]�3f.��7v�@K���&�@�j��o�Ϭ*?�[Q[�5�+��ڈ��b2EaM�$�1F�[����x�����������J�$nx@�J��QZj���c���l�x|�޽��ج��`�,���n���x��y�GhB�{QSmu�é�W���.����w�oO�3/�o�:�$��Z(0q7�T���� ���L�5Y��k~��U�t����\���v���e@S�7:�X�;��j�`�!���~��8��}<V��=H�{u���x�تGc`�y LL�y�3�S�$۸�_�Š�ـ�c�]��wG֏[�3$v�fɳ�x�*qL��F�4$	� ��79�S�ַ�¬Fr�D���6��b���?j���Aɨ���1�e�J�{�@,į7�я#a���N��� ;�3���)���k*7���ט�jN ��s��؏	'3�O�"�m/�?G���x��ы5�
\:��u�w��kq�Go��;r[O�(I��!��>ޫ3� �'h�[����F�ڹ�� Uĺ�bx.�`�1���w|^Ϛ�,�{����e�H� ��+���{CE[F�Q���I�2�^���Ǣ��~eF�͑-��P����x�GZ��}a�@O�U{դ�o�b r��~�q4�C��Ȗ��z#��w���d0�&A>apj	L���D�bl�~�X$���T�t[(~��lЂfn��N�lT�N��!Ԋ>G"0���h|#W���J�YN���r8Wo:m�B�i����m8v3܌��@p�/�C�kP�{o���<eg5p��	U�Ͼ��g>rk��@�j8�� Z9�7��e�s�ٝcYoLS��3��??�����������\?\^�2�^�'u
�>�yq?�
�'Z�h��v��k"��	��TWp�MO�eNH���
�ب%┒Cޢ�3Ɨ���O��0�L̅sҴ[���R:@%��A�ߊo)������ �����3�R�o��p���Y��|8�XH��Y-�p<@V]T�'�cV6
�yn�̆�����<	�bcXGa����b���-8������=���9Qh�ri�jx��>%Q�s�+��[܃�rC��A!�)7e�Gꃱ���Y�u�Y}�
�Ӯ���A���T�A�	���B�ݼ�G�C�)j@�|�`�D�{��A޸Jڭ�GO�!��]&��ڮ�:=F���Ç<݋a��D/<�I��@��`��Ҽ	+�i(���U[���\Y�=��״7��#,.���k9���|G���=��j'+�X��Ȧ|���k���zs�+��F~GY����v0N�T)
"��1_Z0V~��N�*����_��+͠�n�+l%�z�r��$��|W�g2�E����4�e�;�:��� �-�� �\��+��0�LN�}�0ȅ|���i^��S�0�կe1z��H��MC4x��WJ�v����!��g��v(D�Q�Y��S�E���1>�D��/5"���u�8Dm��5L=g �>6���N%ܹ.桞򃾙����A�=���F+�X�#�5q��˄��࿹��1NvR�t���]���e�=�
%H���?���c�^k�2����"�U&�)���U�;���eG2����"�cC���fqy`q*�v�����'��j�U�t_�h��88������H�-\�ƉH�PrT�ڱ;�Ϸ�jؘN�|��=�5Y9��l߫��ȀZ�����]�>�D�K�(�]=�w�1 �	w�=�_Lo_'A$V�
����!=�٩��g�$i�Ky}2�9�F�P~Ufzm$��7O����>w��T�.�����8W25 r0��=���N���{~5=�eH�
��	?r�iH�	ܟg@��̼��W�����m7��\��Q��{|����V2�6c�
������M�[q;�W!z���%�݋��a��:�?����8�rJ��q�CH�}��� �Ca?�m�8\'���ڐC�O6��P�����f�4&���v]\��7�S$P0��'������R�|+�)�^��;ٺw�r����ѹ4�~���y9��B���]�j�F��H"@�Volp��B鰊�rI��KY�N*w?\�U���[o5��3�7G�3�zh	e�Z�US-�QSC�9�zأ�����&@���½�]����=pvK��P�X�3^�~fJ$0~H�/�/�<5d�.^l�����UR�^�����ϓ?�J�7u<}�"z�鰙������v� �K���>����@u��-\7=�Q�Q,�g�QV�!&^�����Pǖͮ�����E��H�30?�4K����lN?y���F�[3����� ���h֪̒��$�N�p���\1�kԼ>���њ�Q5}�)��$���1���Zk-���*�����)+�v=��~6��\����:���	���m�� �G�3�B�.M�o�`��RB)���+�d�t��I��@vOؗ9�ps�Ώ�����$��r�x�?�G�*�v(�\�%ͺ��7�T#w�N�K�9PW,U��p�L��J?�!h�>OK8���h����T�K�5oн��ٵaXR#Nۊ̦*g)TWI�� drO3��uQu*�H���4�V��I�|B��Ip�����Q���TFm�Mvbs�P;���2���"YD�:s_1;���b=U��r��-���W�2� ��T��"WX�:�i���B���*� Z�'5��3�c��6'<7�z�Dk�U�A7k:�=L3�}N e�Yռ��ŊN��x.9�P�<�Ҙ.����<a���`�"�̮*3���q��`/����N[����%k)C�%i��y����<u.s��T��=�Z&�\��Q_E�[�(R�S�O�ן�֡N~�̽���͌�,Fܪ���z4}��9��J����ߘvŝ#5������D����
k�|�S~P_fjX8�r��O�/�$��˧��o�dn�w_	�A�hK4�Qg =x��Cx���O��z���Ӓl��`���W2�����'����e���<f���s
sJ��Vg�{񎢉H�y��Ck��WFUs(���B�':'��X�,nSIa.���t�}�I�=;E�b����d���X���]�WBc.�J�M�KD�e�
4�"�,g��.���w�"�
�,!��Z��1��5���f��g2�����yM�t���2�YIle���.W��{�n���(Hڌ�����E�����K�*��F/#�CVc *t�S�V:xف:��ۋ�H�M2�C�4A%�&��.��8���N7����f���߉u8��( N4�ã"�K�\-���g�E���zW��Gw%��}v�������<�����h ����5���I	4�-Q��ݖ��!�?U�*}�gv�:��6!ю�?ۉ�yC��lᣓ�d�޹��;�;��C}��N���Yh�����K�x��?z/�b����@Lj`�\z\\=%���I�G�@��G�y5 ��[�/.\�nK�98q�3K�͏�$��3�w9������`�+���x�D;��!!I�0�=�ƀ*��u�I�;�������T�����<�I�$[�Zb�VP����ڻ���o��;y��i���?)M;��.����ME�h������;���&J�o�=�2wS�i�B��{NfW~���x�ݯ܎T�n|@�����.y��>��>�#u6�'�^D��Mf֎���&ɯ�z@ο���}q��W�FhO����E�(�4��G�̗@�0��=�g�fsS�� �y�f����gO앸H����wm�+�7���q!j=F�T�����[�Z�	�4�z�+ft�>�u����L����a�/��qMDHpCj"2�%�fC��IٲR2VgA|d�S��h��7(�*�L+7���Qp����˞�y̫����M�_*�����q��6D���P�`��d�C��2�;*L����+B3�do��3@j��&8�$�s<���=��E�n�ܩ��~,�^)��T�;�2�,S9�t[N�RӚE�{�{�[`ߟS��#�N�1��/�~�ܸG�Wb�V�	Ɏ�Y�1�B�3����U�4�?��StF� ������+)����妮b�N_��N�>Q��\��#�C���Ќ0��f
����Ц��֋Y$r`;"*pۡAJɥXː><��¨c���h��b�&�2�� `�>�&�,Ȗ���J��S�8޷E�$v��pU�n�u+�Th)����a.mi�����S��ܒ�'b��a[�K+���
I#`(��#mv��҃��Qe-� ���̻O���u~[T{bѠ.Y7w�ҶOP�q�n�1�%��=�+�]�����2���ĵx�ᯓ��?Ӯ��S��	"�p��3�3����K<��A����nNg���E׽��@Xc��>W;={o5��8���()�
�:�L�Y���� �o����7O>ص���_�v9۹)�����MƧ 
��J \�l��,���3�;\ѝ$$�/�{c�pR�IX��R�Ϥ�=2?1~���/Hٱ�昈��Y�QX��D|Y�����3�*�m?AG˦;��`�$��׈E���A�B!WI��;�Ƣ��4�% ��OX�59:���w��K�$� ��CAB:� �:��b���)� �����Ҝ��Q��xNըߟ���"qvJp�>�)*cb.Y���և��H�ʎ��X'�>:��\���4�˰�&�"+W��<jLa�Sl�|~k����� }K��O��c�uvr�J�
ND��[�gh�:�
r��W�}s�e��[<%�a�������]QR+Qk��jg�f����T&�ժA�-��L���r	ӬG��M��"�xG��suE����t�E�Y{�]_�ܟ��65F\���:k����;u��8��M��7�$�#��8A9��H,��-�(�N�I%�փO�YUw}OC�Wr\Rj���`���"�"�r���i�+64�_�#W��aW�6����⹍<q�z��E<'��?�i9k��Z���F5�,�J�N{�ET�#�ՆЮѬ�i��,[�w���.\���gݸ@�4mÞ�T��L�OFӝ�s�(�A��{; �I � �z���S����0� ۉ�na��P�
d��"��s�rOi�mx%��K�� |���mϿ�&�ǅ�P	���Nl�6�eX�1�*�H4���ߨ{}�v
�];Vq��)���ᦩ��:i>��9D�Y��݆ΰ�MqD���`l�*�2�[3O�XP������H<4@5�p*�	��s���� `E{��G��a�q?v�vD�8�d�t<�0I�nd��m���n���A`u�6+�O�[`@v���
����_�8w���K��l�e���銑5Z8�p�U��J�����_M�D"�<��<���C���>pN��3�J�O��@�GĖF �y���',#�<}(�Ǆ
ƌ�l�9_  3�~�Ff6�=����CQ`�Ա���cX2k���h��
�)��p��a}S?�dЎ�����	��u%�(ĺ�C��qjaIjv�d�)
�V_Pʬ���{(��۷���9�%Ti.\��fk&�Ǽ`ɩvCY��<V�T��cH�cH���JE)�vA����OU���K�u�F9�&_��(xf԰6���{&3!��kOd�ʞB�����E����<�ܬѲ���t~��kt�g�q�����o�i����]��&ZLp9�Z3_J�F��i14���V������}�]��nW�����y�>,ހJmK��j�B�N�s��E��ʘ��J�Oip@X-�,Q��g��h�sw�.n�jΝ0��7g���r�.���)"���������"����� S���H�e���X����=�C$���)#�n�j"���P�[U����Y]�Ko���H�C������6z�1|�Ga]�[���S��/�~{��g���;#�
G/?z?�+7]RD 1A�#��L��8cL�!�4F�v���8b�y�^yK�#�t;����Hs@�`�%	�ŎQ����^�7��> eKP�Se��\��7J�7��2�XCQ��L����.]V��mB����<��(������_��ɘ�t֛��l�V6 �VP/������?��J������]	��-����������rxURX�l�#�>Ha_��&j{�ِijI��9��ӌGpn�D9���?q�4����n����}oJ��2����Z�kh�wto��9r5�"n7��_b(,�e LC���׹zL�k�R瘼cyyu� �����T�/��=��Q�L�2H�#�ZO;{�lR�_��	�^uQR�j1��4	�3!R��e�>�I���u��SI��[�s�t�?8v*C38ZLA��ѡ�n��ښ�n��;Ix�1#dMnj����6h�(�h���{A�k���_���{8x[��º��|�5���Λv� ��?P�G
�|!{Y'y�Q����b'�����lq�q��ͮ��u��f;Ξc<��#6n:4�A'����@�k٪�$��k&��R��֝z%h`xs��ah����훂d���񝥃;�x	�h\������p����E�;��k�g�'��h���l.2�U�X	ǜ6�\�&��_v��Y�&4\��&]6^�݋��D���5B9�֤��m�H�C6�c�>���?�%���U[�;ɶ��/Q��a��5@ .�á��}�L(PU*;�(:���}	N�N�6�#k �kɚ������]m��d	�D�!!�㙃��D�����"�*����8��.��O5�Z^G�9,�贠S����b���@�����P�"3ya	�, f��g�HH� ���^S7�W�x� ~[�!�[w�4?��{I»�LR���WȆ��$W���F��cv�+�M�[٧�"�Fm�l_�Ж'c(�TÜ���ذm ������j*ܮ0鲜���n�����T;3J��}�E	x�-x�{�� P��?3��"'�Ӗ��M��ނHnˉX&Cd����[o�)��P( ���{�!wp�%��o�7I�S�� ����߅+�E2Y�-�;�ӯ�е�c��9&��|���x/����tm���k�y����2�]6��e��0`o0h3�pI&H�f�t��� �Ի��C�ߗ�;u@JB��b�2��SMQ�J/� �biķ�$S�4�:�m�`&�V
{�V��{5�3�A�ƈ�JʀR�]"�XDb��0��Da�8�B�1<B�'��x��PR)l��4n��<�
.S=)PЏ���C\�/S���So�$�N���ń���F�m3�h���p%c_�l�pY!yW �\����R��P�[��!�U���T�������-<a3;�l���q%�u����8����8���d������C����LX��&<g�Cf�R�8��w:��x�h�6��)ܔWI��'�9 �$�L蘽_L���F��g%uq��V���8�U5���>M��鬿�Da��<�#�������
��I��8�*�R�W��8������e�����~K�=�娌W�?{]��l�žkG�����-8)�1Z9]@O��K��(�D��(��r��R��|�g�J1-����E��c�4㧒����B*Ҕ��+nJ���s|'��,�fk=�/T� ţ���F���.�c���[d9�H1����_p�c��3x�6�içV�ߙQU�$2rv_
�G7�r�����i��Tf�*�&<h�)0������S�� �_�Ǔd�Lm���-�]G}��j�1�lz�n�>��Eɀäf��5*9��� Ul�Z>#g�r��o2�.�p-�j����)�1��O�}�T �<Xv���-������@)�&�J��]N)�����Z���H#���!��B�Y~>]:)=8z<�Ry�q
�(���&-�F���m�����gZ4<
�'Y�?�?��kƎX};�h��\O�+���T�/{����*C ����ܬ ����S��i�U|j�w� ��9�����[��Ԉ��)<�y8��vt�)s�ؘ�`��������2"��,�w�V�G��c�Iz��j�x�ϼ���p�
.;�\��Q�����č�dIϒ_EE���m�s���C�� !��$_���R�'�rG�	�z��}�>g��&$�<�"�}g7Up�LQy>.�m����m�!򱽻5���n�+�&=��a3��&c�].�e
{m6��lv�������D
 ��u��G��ŉ��a��,P��IIG�6���0\c*D�q4g`�ϥUF���h����h�o�dP*Qe�/7Y
���
D ��Mb�L��N�L�,^\����'T�<�{�EZ��7���8K-j}�=M�Zb�3��>�ʹL�9������J���tU�bs�}���N��$q`�������BQ��<4��mZ�CV��lD.!Z��+�~z���?uܢ�+FY?��^���L|�h���n��̖B#d��`^����T�ۨ@�4��/_��&ggkY$pB(�f+`�J��h�������p�a�'N�w�Iy�6���S��+�"���g���dSr��z��Ģ��w���g#����{� 2fk��^Ȯ��W_�*w��=�Ų����xG)�$����ڛȕZ)%x�V���d���8G��,��s��CjV�9�a[˲���O#��D��3|k���m٭�#�E�@Z:�_ե�s���%��X���V���c{g�l�y�����v*�3���̌�Dm����vϰ��7�r�Q��MJ��_uUp��HA�}�� |��&*N��-l'7Z�?���C[�R}��I����חh"8��#���w�w{`�����m��ﮠ10�y� �鰍y���Ç��������+W�Mly�
?l&w7��\�]���T�7��`��� �&d�.�"?ˠ��I�=�Q5�sX�|�ki�3��|=�~��ZF��2����0�)��eĴ�P/>Q���'n�z��N�JH��F��zo�kμ/�HI���qTw0�#M��U���}�%���Q��Ke�XD�����*����/+\1�W��~;��/>j%�	��e��2��89�b��� �ME��6voV��� @�����`w���@���3G g/JE78�d���,���:�g���l�Fu%��ҾP>���!l�	t�,OQ䮉c	�x�aO{�4(�2��eֆ�bQ����]p��xz.ĕ���L/�w��w�s�;���mM��j�ѾQ�0gb�nCgv�Z�}�[������~R��D�O��8���V�k���o90�f���X��0@Ci�g�i�jn�oZI�
��nǡ�v; + w��"������Gら�8jyr�\WK���I��(�S=�"�R�p�ͤ�s�bd�)q^�r��Nu8��T����{��_�n��㫤�����Ot�b�{�O�Ƿ��M'I{ ���}��d*��ռ)�I��}X��#-�/㥂.�Y+��hQ�i�L�M��7ه�V�(|��P�� ������:�E�'8���M.h��~�<�PӢG��>>�O���X���eKUի�]n�)��J��ɍ�1Y4�N)��`y�qjZ�wIJ�z^�H���'�@_ت��t�_�Q͕��[^�����b����eu��V>��T�5�}�A��"��ٯOO���Q�$�~��9R��g�E�Wź���6Qza�;:C��a��)�{�����vN�������p�h�S'���a�+���ԉ�os�JgAh�D�$���E��؏7A���E<ƾ焅:
C��)�!�b�i׷ZM�w�L}�q��_A*���K�����?;U�^�ѣ�,1�"�"�6����Zm�mw���e�peFa�NZ9�q��1
NK%�;����;�� �P�T��i�X"�C��${�ד�݇��{���{|�'b*�W��0wʁa`֙���a�������+�|Y���D}e"՛կ��L3%��"�2*�cծ<��5���
)�R��E���Qܑ>$(c�t]�*o�_J�sܒ��_�t��TD&�ˢ�j)x����\� ���{�7��gFՏ*K�!�,
�P�L��R�"TGwӀ�H-[M(O�g�b�" sf�A�o"�l��+b>I_�$v�F*"e���L;p��ʤ�:��L���d��q�;�X�OL�~r9���2�M��%8Q9�/zC�7�ϻ[Z�
��<��C�k[�%w�m��H�� ;�C�r��]�TLѵ������e��9r�`�}�}IS8@���T��<���| }�[�E�c%	=EJP.�3״�Y���5E���U��I����Ix���_B� #�ܯ7��S�R.�Q�yxb��J��h�xa~��wb8w�� �9!��)�u�ףXҪ�t:�.����|&�g�r��&M���yK���\8�H*�V�,z9��n'��P�BuU�ؖg�-G�#s�C)t7��~C�1�e�f����?]/:IP���'���J��9�ͮ
���(�'����?�:Y�*����d��zⱔ����iu�ti�A�b1	����ߟ�k^G���Q� �rL�i�ď���c":�'�,����$'�+������^����%�k�u�?f�/1�tV�i?+�1;���Y��-+'Z���[U�A�?5б���q�5m1{�£��tF_Wr�E����5����Ṕ�h����ɫD W%�4M	��\pE����֍��S�4%�:�9< ��3��$3��Β$����������X�hM|����鳏q�?�=��\yAȨ�?�`W�4��]���p�i����M���A����`✿V	UZ�͚-���ՠ$���I�,s�\ s�Yh��e���ưHJk1��Ƕ��"�$��ǰ��W*�Zng~+u·Y�N��q-��sy��n�W?�|M2�%�ߟ����03���F�o �!�<�-w�_�frI��`\�#6���	�:N �/�u�
�K��m�r���גOn�zV��̏�k|ÄC��=�Y�-�h�Iy$[}�~JlS2���i�.�E[�Vr�(�
<9ص�����٪��OM�����'KB4_�K�ȇ����J���)�@��������vC]��,�ep�P�]�hd���!��~����x^�"��~�sVߚP�r��ȭQ���[]�ؽ� ���`�&u�N���ݑ�}��s�0NL�?4�}�?S��e��5�gU�dEܺBE5�Y�h����{z`#	�ԗ�J/\�v�d��I�`;��G��Z����7��xE�F�=HF��B�r�y�e�����a��o�WNR��ɾ�����Z����
kϑLf�?�q|�����R�J/gb��i��s�:�u��	��Y�!��SI�wX!W�	䟝e�7�vǄscWQ�$xԝH�B���z����>��:`�jfw�[���G�čr;�1��a MO4!О(���Ѫ���	��Vi]�v�K����KԮ�M$�K�����T��4��;�bv���h������pxHas�%����}\9�e|mr
=܎[�y�T��8z�fM�U5l�^���v���Wv�oPLo��c>��%���J�ه��!�j��Z���j�;�3K��dzoN��)�*Y��3��5��g	����n'>�,I0�UoЏ���j�f�s�F����:}�#F^�I�VK������2IVPT��z������)�B�����4�q�4����x��������Ɩ�Mk�����G�47�虷QE(��K�Uf:c�X`;0��R���)Y��W�U����~�e{qߨ3�ga��i���`�8\d��~�cw; =s�!�=�������w�aC������̌S���h���]W.�s�A5�P0�5V
/�������d�r��0=�&qMG��.O��pK0�R /T*���!��p�3��v�_�ܠ����8�����w�v��$� <`P�p��N���I,�#R��xs`��v��-7�G���=�m-�x��C���� �8\2����%1p�7&v����mx��nq�Q��� ����{mq���Gk��� ��CЬ0!N�3�Oԉ.��>���K�ܝDZ�b0��wr���\x��2�t[A�X���B;�Qt<$iT> �]9����2Fr���Nю�۩q�H#ҵ�P��ݵ����q����*�)���`nYý��!��5�f��lO�{.�b�^�D�[ #�G <F�Ʌ��~�*��p��2rG����Q$�S����'��Fſ��_�2A CL �SJ�{�?.�G�n[T� ���@��+ZGΎëτ���L'��������H�{r'6�Ru�o_D��Uz&����>O}KH�:I�~�z�>t���3����"K����CR0G��"*�2
u#	&.#�.���dm�u�|V���$�U.��\�.�W���[�ӳ�\�,Ce��}�P0븚�<B���Zn���U�X��>�ވr��Ϥ~n���Y��Æ��#*�zw1�b��s�@���}8�_����� (�%`f�`Ts���~�K�����N�L��ry;�!�?o�at���2�V$�^��c�f
^ʓ�`d����]_5�c)��|U��ٯt�]�7ɳ�|�O��b���3�hh`�wD=PsBQ�� �:
H׍��7'�jg ��¡7c��2�-���c��zb�į�#���Ъ,�M��0�M��3^�D���V �+�AĎG؆����ː~�W�*O?N����=ô���P�ǳ�H�,_��&�ߵ��"=8,�wF})��K�����+��S���CD�׬��@L��T}��[`�}���=��;Q�pLc����(��6�J���[ٮ�>F��P-ZB��'�;����RЉ�fg�.;7���/!���n0�NfhŪ,q�e2z��×w�٬,փ��E���"f��s~��":eI��c��-@\����� ��@�ݤH�]sτ���ikY�o��a�;_l) ��6Ν��V�<����%��o.�9N_ܾ�>&>�X@ok8��9@}�C�m!�'��ͬ���G�y�m�4�K��U�6m�'儻j���5/J�F?���x�� 9��^��??��)Jb�����Znϱ �/f9N-�d	ۏ"�ҳ��K�ЁY{k@8�L����Ll��\�17�&�K�$Yb+&��F21qq1>
��1���L�����4��c܄�~1����d^�B��N�OB,�9��;�ZV6U�������s�zK�=v~�����`���B6M0JM�o���|��^��D\��d��5�2_xYY��^̭G6ѝTy��\���x�=��^��3�x���w];ZwY��w�6S!Ts.���<&q�O-�Q�;�.�dZ!�Xm�q�ҁ�~��U�#!�c�y��/@ &B�b���K��с!��)j��`��.�ApwD��W��/'ch�P�T����-��ew�~<��SYiۙx�h'�ۂW��*u+.�ve��bXˡD�)�aK(�����'YێWb��ɜw/����(]Q>gd�kD�>Ţ/~U=B��><g�fC���gTb�bɓ�l�g�.��$�D
��	�ta��1�[=%x���U�Q,�S!�+7�}q/��J��^�k+X����k�gvZ���۵� �r�!Z�5Ey6��֬-�b/�s��c+��x��w^	8W"?Z�<�F�'�}!�~"k P֜{r6hǵ#|���BI!U��c
v�JpJ�ܥ�o�~E�Xዓ$��PN�H�^��+���C�/�R�\�L�������)ߕ#tSyI��v�$����ŖG�XJ��I�y,���n¼� ���Y\*�9��}t׆y�l�*�[F�c���&�a��ޗO_6�{����-��ٺ�~����]��N`�r�%�/F���௡�H\�8L�0A���~A�Y"t�	k�-�ӡ�fb���VЄ�D�ߏ�&PdŠ�a̗��pC�>��p�h<OϿ_E���_�O�6���!CsH�`/Z�x<�0O� ���ɬU�؜�wC��+0~6�a�Ll�뛐-��~|P޿X���o�B�_��8���#q�:����^Ѡ%�<�yEV�Oc�Z�3��uӣc�Z�Rm�=�/}���S|T��p�DGA��qEB=jq��s��Q�P�����[�Ì��U�)�'�];=K/V�� r��6��.ؗ� DG��L,�C����v�#?�~���ʌC�[�D��GB:|��_�.��lbИ�*�kug�m2@��sO�$�)a�&��l ��C�k�d����F]�;�̳(�C����Q�E����*~Ox�
	�����ɧaj�]����ݕ�Z��"9��k�`*X�x]���,C��y��2�a
t�\��~�)L�^Ԓ�	\P�^��s�',J���t������oW!q��5�%3T��$n�M�8�v��gB�B�d��̥���s�j
���'WI���]�J%�6D*s��̥�<�g�c���H�tH��WÝ��p�~�C?#,������T!�J�+:%�g�g�ᵸԕ�u$s�HOa�3��b�z�ƈ��f��c�#�;N��>Aq��!�{�;r1�يH��f����f�^�ꑁ/��k�F(�5��|�zj�?�1Ԑ!������K�Jױ^�lJ�>.~n�� �)� ���$~e�B3���_���`�3���q{$�Rv}�r�Q�9fѺ�jq&�g�\ݴ�MZ�O��"�DrQ�+�荆��� xs���n�MwPJP�}�L�+ƠR��ZЗ����i����K(l�_�a�t��52k����V�U���Dz�k�b�|�z�c׊�O��1;��l �J/��B��r���os ��(����o�a��2��,RNW���p��'�Ͽqaiv��Ԕz�'�M������Ҥ���m�cï.y�0���>7/u�I���:y����$�j�Hڈ�tk8InqE�ʸ#�_�4_�]�b�Dw�V
P���%��3am��jm��n	�� �'
?k�)���I�6P�.Fc_q�-��������/���R:8D�;��7t��N�4v�G�
 fԔ�(�����ȯ��g$+��_1��}�=�K���&�6��n��嫢� 6�m�lP��	@��"�k�w�P�d�5`��^,���Oj?�s^�=�F*PԢ	Q��T���K ��FOIy!]�)@�Oex�]��K9;(pw(�>�:�P��nK����GՊG�xb���	����.�����:q�� X>�� )Y���Cd�:���2(� GfD��'��X����0}���5�i<�K9��>��n?�s�l�+⪐&����uL���%W㡫�#��Zt[�Ppj���i ��g�'-U
5WD}�@n�[R�uM|f�)�s��̩��9FC�rvWk��#P��I�ˡ��jX��(�B� ���K�^�M�l�����K�w��}q�%\l��C#+;DC~��j�>%��̓��`��i4a&Y���bb�UT,��1�xe/�*B�9��?WS���&�l8����ĉ
8�%���~�mV��I��w����$t�_~����E|���o.��Er�:�]LNc$�Lj4�Qx\�]]������>sa ><rxG`�R�l\>0�K�e���)Ec7�&��2QD������s6ov�	���85ezv�����z��\�D�t0.1k;�(�R����
��O�+����%��&؍0�.w<�?t�1�����_��0���W�*e���E����i��5���鮤����;4�܀���CQ�_"������ʋ'�x�n+O���U�Ԏ�Xт�ݟ��)L#Y�4o����;�"�0���gּ�88���x���6P�7i�5T]����'����j\th��k*)��|4�z��)�[f�rp���s��OH��G�!g�B�ᯩ�&nbl[��U��)B֔]
�Ų�o	��r��j�I�P�o�n�6�3�N�� �0A�{�A��.|�wqr�P���5�0�E��o�E�OUgf�BdP�#�\ٶH�iB�ѯFTk���<�@�>�k��!�A��i��2��|]��	?%	C�T�IS�ý����]������I�=IǂC& �O@�����&�'�#������^����	,���
��`���	;BL���O���1�A�B�����(�����~�+r���|��&f�Iһ���z�)� b��ȕ����h���ӚU�Y�
C�_@��D���~:�H��� O�ٜ��PĬ�Ӵ���~ܪ`�Lu)���K��41�U8��Êu)�HF_�,LVD��K�t���4f�<����c���z�{3.�s:.�MY�QQ/��U�y!	�'�s�@/�
�r���Fñ؍�x���0��0Go�_�c_�wwy&f[}w)��(�S������/I���^�_X��-e;Mͯ���:�.��?�X���CQZ��% 󰲂�Y'��weI�-V��I�E	,�/����t�#���u�TPi����������y��K�Ï��X����1Wr{f��rw	۔X��N���V�#V��H��+=Qo���J�0��B��u����q��@�����O1ˀ@!�R2&�`��\Z��Vo8�~Ǿ��l��������O��b���tg�m��j�K���P��Ӳ!Â@��-����!�i�&��e�s����Ny�|��]���1�)\�I�Y�����)�-��^=�	U+�L�i٩Ĵ�~�a�����7���%<���o�CudUt=�<�J�D�ɍ��c���?�^��>����^����y\��88���X���/�v�O�S$��:�]E�g��X.��Ù�?k�l�$�o6���ѫ��O��^(���op+����.B�Q��G-�����Qa,4x�F�;�j���,pa�L�yz�o�k.	Ni��8;]�B}�c���"�Kp��o���e}D�Ϊ���	JU ��g�Űu���۽n��ި�2y��ł���i �(b}:�c���R������ i�'o@
NU^�-�K8�L@Z�B�!}Ii撞`a�|a����D�/��z�7��v�]�JVQF���%S�)��-2=�d_��I1�T�!�u��h����;$��ߙ8��e�%3_���(���h/�T��}S3�.�NK��qYwH*p^��K�(�b���ǐ��T���a�E�G�8���t��\��M���s��X1���n��p&�0���<�#��A��N���ܞhe��(CH���a���2ܿBf9T:�rgN. c�L��OS���� E�<
_u`$(m����Ǎ�[�Ȧ�E@>��	��]���	� �͌�<?=MM';�߯�,�3��uL�q�@2���eB�~��s��ob���M����X:�!,C����R������߆�I�D��1b��z�zN�L���`/�6�=W����V�=$�x\Ì�o1�}�۫�]8�
H���l}Ʉ���.iKo*���Yx��o�վ������!r��a@W�w�z��]�u�qw��������?m���q�ow�HX���Q�9|`���2qW-Q�uS�3�]n�ߘ�6�#��J��BDg����_s�!8(�O+`�/��591p@����X�|?��(�9�:?�RE#Rr̻�$!RM�Y�Ox�Y�0nq��sϧoW�&Fb�D�ǧuw��D1���̅@Ց\5*�@&I�\����[P�1�{��b?��]��Zk�o`��S�1Rn��v��V�`�H�)B�։57���y���+6�U��ߑ:);m�y�\F1�~v��A@�Tg3[
O!0ĺ<#�T����8S��'��z7~[��p�9�g�N2��Α�▏$J�7�\�4s�u�V��n��yϏ��W�M5��]�H)D1ZL�:�z,͕����ME�/v�MZ�s�o>-D�;�
���������kh*ʅ��x�w�籀�*���Ƹ�~��E��ŀ�m��Y"Q1�c�ΤY�F ����>>/4h�!-&x�����fX`4>�D����F�.����Wu�{�}��l>�N��qr�w8ҋ�N�k����
[D����rVCp�:�Š�t�e�?<s�V�!aQ /�*����_�$�G/�؊F	�G� [݅��'Π���U(ة��S�{�ҝ샨�jm'8hr���`�6R��y��3^��7_�����{�e���ɖ3	Q��΁`��A�A�A=���K b�Оȇ�e������_��*�٩�7_���N�XxFJ�/���@9h�p��x��j��i�K��'C2�A�/�j-��c��knl�g���L�O��_K��
��A���!�^XQ�"��X��$>@"����ɱ-���ϓ��d��[`F��&�;zwp�e�V���o�ι\�KM���� ;�I�|J^�<�,�M��%$�+�Tj��2i��HN�+��}�+Yh�湰=�UJ��<M���O��κ�Ɂ ;���ߨ`*�JEN�&�}����.*6ǜ�_������/����qSȅ�_�<\V~>o�z\�M@b��9���T�Ä��v�S�	BY���0����êX�I4�"$Gh��*�ب��e�Y:X�M=�$� )�z�:�Y�+�D�1k��\�9?��gG;W>F2���\�r�EB��.
oS�Iou��<m�I8pm`����d+�\�'s��W!�@����@Pǲ�@�8o6毉��'A�������x�y,-�kHKd'��N"�2���l���ʐ1��SR�A<^��C;��4���z�l#e3�vbD}��,!@�Ucm�]�.Q�P+�Ҍ��	���* F�Ӗb:���n|�YE}�z��~ds≫�Y~����}���֭����mY�sYOm�^9�F�������%ٍ(E��]߆��{�r_���]a�.�Iy�ڐ��2�t[�ڪ�FL������۬�]�2/~�w_A�
X}���	��`z�T����Ѯ��'�-iYQ�M��*�Qa��J��-ۙ��b�X��N�$R�@�ˈ�+���
�5�p�۩F��F������$꯭a۟�2P��`�[JKنf��g�g�'������L�7�!�G���.j��)�N�WuC�~|T��>*1��q�|�
���{	�f�ys� �ؠ�[�����}�/{H���"�7T���w���
�0��G�P��u�����e!s�AO��	w�K1�/Z���/�	�M��m.���|56{��֒��}��7F�*�\{M�a����e���yn����sW,
����~����_@Be��sG%Web�N\	��2�0��G<�K�љ���>�j���Fq �;>�8�q!��B��+���6��n�-#�S ƹ������^������է�h�x.�jJ6�2�!ִ�I�����fއ�q�[�W��=خJ>�w^�ˊ�o	+Z"��6ü������e���r�&Zz�Y���!�W:5~?��.��>�F�n�2z U�۶}# oڀv����S+x��0�d&�3#(h��S	0M|dWZ���j�Yu�b|�P�Q������mo�����6<x$��\_B-&x�_TJ���bvǪ1��o���JE��Jq1���io�Xx[�K��)b�Sw��Q������jf�ְ ����T�R��O���o�fw48����<P"�}�� ���kج�R�F����n�^�iil6�Ưs
46<�M��jH�IZ�K�Z�`�H&�L���+�?Brh���ZN?����l�V5ո�: ֋���/[���p��3���t_���{��_Ȫ	Ƹ�&Gn��[u:Q�ȑ�$�eTw
�-�zojZ�7�%�*��{�g�%����#����ZJϐ:^����L��)P�`��s"d`!��Q���B2IP�X��.�*1��s��U���I��4��5Y~g�je���Zl��!�(t�wUr_����~�*�]n�|w���< ����\xPMޝ�o5罍����J��Z4�e�C�{�(�%?���p�bԈ��c�4�5F`0A�H���&`����S�5쀘	����p&{�Y>�j��uY�tKb���.�$�H.��$)�`��j��·'�S�*�>��g)A��
Q�(ܡ,~�N���	���Y,�#�B���w����0�BWS��:��pݶn��F�sd+�MPaL5��=Ko�g����D����/LC��5j۾�/,͟V��8ː�]�z��X]˰�[���m�T�a~˒��-qHȊ!����_����,�06ΌG�<,w��\���w6�WM��Y��W���wQmu�뒎p��ڜ�44�z�!;�ٸ�o���|�n���-0��1�xM�����W_)M�vI�cg�	�$��zK���f"1���e$فR��DeE�ʹW"�fѼN���3Й1��Ƈ�;=�!��9�@4#�w�sZ��a_���֍�7����]K9T���	��vK����Ω�ȱ�aغLl_g�|�X�+���u�C�
Ozc�ɪ��4Q���������f#��z�B'�S�c�nzD�ܞ��"0�[q�*���懑4� m��@�|N���t���vS\ԥ�dOֹ9�C���X�4/GK�Z j���I@d�)�w=�+J��V�nm�(72v�Tc��U��b.tY��X��E>}�J�0 =�"����L[%Q�8���-��:V��+̓`�V�J.�۲ʩ	� _�E�!"��W?�������ӄ�7�i�s׀}iؖ����G+0�dTir4�^���$�U��6�'�F&�З��f��+�H�Iy������_̮�,�F��I�L����E9��y�l�v_�-ء[#v�&�˜Vu4<}V�۠�$�{�E�O_y� Pl�`:�3��d���ztVC���.��:�4f�B���w����ۈ�i��*I�����ǡ���X�)����s��G�nxT$��yYT����(�����)�H����8�#�"�X7U9$���8?j�@��:�kHxP�A�>���g�g�̨����B�
y��glȥ�b�L��o��$K��$���c�|Sg�կI�K�����������g"�hF;�ה ?&��pܐ7��:��|Æ��'B��T����C9�c�=!�	�[����vo�8�A%�)-�ع�'�Ո�d��m�Mn�9̂۬��x~1�L�~�h���p��j@��D�����ȫ�9��nM�ɭ>����Y.P�T���%U�`�<ٺ.�f�~56��RB�i"��y�q�2���c	a�_l�f���V�E����n��'���+4�$�M8�Z��c93�`��L�0h�PQ%M]To��L��+�2�8�.�m*_��c8F����ر�K����\W�?m�q�5G�z�?��v�I�C���g�{����"rQ\��Y��f��L�ܖ�-�-!EJ:�@�5+�;#c����^5��I�L��,�2�q��L� #4�,��"��1��V������t�r�)�qJ�&�����mQf���ݪr,���UqfD��.2t��7o�/n]�������]GX�3�!�i�l]����:}���ϛ�P
�J���.]cb����i�+��:6E�u��P;)�T/7DkU�)�s��۴.B�&%ci���׾�i(#W�>�s�-�+z���m�&S��>�w�����C��_�q����_��G.��M�#���(�<�fó5O���P�}[�H�k�_�&*f$�e�M�CX=�`n��U]����#uǏo�-�a/�����]�T�':A(Hr%m�2xb��N�߃ۿh�MZ �Q��C3E��P%�\+��ş@[\��yi��6�+�0����{� {Gކu��{���]�M�w��Vʥl���̤3���k}�o�m��GB�M�q1����5:�{^�:���5$�CI���eo��n�01�W��6�Ehb,�o���6~���������U�4�텱���xh���
uS�1>�sy��P\��U���mA{ 7oy�͉<���it�xFn;�R��&U���<�W%�?6��g<r�v�_�y9X�4�2?a�_\��è>�.�k��(���>�m����l��Ȁ)��ؼDB���Q��#�s^��d�Y2���=&�o��)�zEK��Y�bNZj��X&�Gmd������o���%���
A3��$��uu�@s'Tߕp)!/��r{���Zl���$�^�f,��� ��7��F���8o��J� 鹠��A/Gp��םɛ�il����G��]R=
��j�J�J��Y�ۃ�w���I�`[e�g�mM�u�U�P�SbJ�W�(��O�'��9��j�{@��nwM�:�����-�{A�#�*�
̺�"-.�2{�y�W����nE �LFt��*@ߖ6�����<ev뵜>w������*ޣ*�]q1Pf/t����C���D7���f�Z�NmW��EN)HTm��{����>�2���Xa�2��&��)�u�������!���4y��w̦��Ŕ�5����H�;���Yy*�*�<��X_��@�;��%���u0X)n�{�����ך�Hk��Ζq�7@=M̒-��;0�x
6�b2F����
8�ex`~�^Y^�J|�k�ь�E:�e��`�8��(4�^�^&�B5�N�Lh�L���-�[EPEۢ2�-�Ca��M
��/�˪�ߡ$�$鍺o�m0�G2��_:��lC<�!B�/���n{4v�-�,�\REE��B�>LD��}o�ɕ ���/��K�Q�����g�YIƸ=�����6Y���X�̾�P(+RiA芟��>Z4}�h@^��s�p����6i!%�b���*Aѯ6*���$�ӓ����BOʑen�a��"c nU����b�-���3��z	�OY�� �[�9��B����?F&ͭm���q�h�����Rɑ˻��/S�c�0��\��N����q>���]>!s��(-I碥���j���,�����6PM��<5?��4�ńke$��p|�b��[i�����&��$���0T:��* �`�B�xR����ͬ���>�����8��<>�%�]�{�F�LֳN�K�E�"x�a�_�h���0��~�D��iR�;�sΰ�`���e�\'��3���һ�WiB~}4q��@=>:f�V����#�����Y+s�m6P����I
���cg$z��i�hHf(]g��`o)$�ѿĺr�4����)wѺ�z4[�a�6@����]�j��I<�a�}�4�[�d6I�r����lS��BL�z�U@ṽ�vFL;�+���`��,
��1Ck����=G��B�p/�0)J�1�V��d'.�Uy��	 ���砻����ti� FAmgɵ|����K�\CX�v���+w#m��j���殃�����x� �4����)h�oѽ�;��a�E���M�4�¶Op�eQN�A{}�7J����c�ϞPD��d-�Q\�����YZ�F���Q")T�/���'��"zp��r��9PDA��n晐���>h��Y�3�Cj����m����7*�/�;>�m旒t+�:L��tr�	�0�Ć�K��~�3����娡����Җ�R�S��8�d��-�#i�*�����GX�tvy�2*T��^N��u�~.�n��_�][�ݹ��DW�zo��ٔ} �mq�� �6A���%�wj5���ǧ�n32� �<H�P�H<-.��LGUX��Z�^=!*{�	���V�=���#�.WKx��e4{��Dֈ���>�� t���ǩ(6�g��9j�kWđ�H���w뀰ü��� V|��r��8��l�e��'�3���R%j���y�@fD� ��J�b ����J�r�����M����^���qCc}W"�O�Q@$07yKsϟ3B����#�}�o����(��]M�?3
-<�L�,��V��?�~���gkrO�gb47Un9�����mTC�.A4�پi�MZ�>*tκ�$�L��㪿=���dS��a���ֶ2�/����b�0�Q��W�S���y"�Q?�p��+:�������� �	E����F����~��$����ќC�(u�`D�g�$�8��������]�怇�i�)��� {^���j���0L��I�x�y~��䇺k��tۯ��d	���Ä0���N��U�P�4�:gvXlF;a{����g���{y����/B2�5K�"x��!�R�fZ$�8[,P�0/TNM;���>!�|��Lŀ�>�̳	3^�3�R"�ט@O�c��C�j�~Q�x; �e���"
�3^7<8�%�]��ͺ-����@{!6��}+�^X��	�t�$��U�o.e_*�UT��'yD���p�3�ɩ^�@�:v���$�X���eQ9د���*z����-;!\>�Jk��1y/870y�1o���w���}Q���;@�+�E�t��J�����k���3pZ�pλo
k#�*oΜ�o���5�X�w���z��'�'+Y`��HW0��9��u2�84����(�Y�%�=e��(�=� p��9�@ܯ5I�#\��]���𳕢��m{�Q~�静Tr�ta�g�D��R��1/}N��iO+r�;���?�7�^��?����MGs$�e%�!kd�Sυ�JJ�/m�m�a1g@4c�ģ�6azj��:�W(0=�`�OW���T���lUR�f�CN�����:q���H֦C.�ȇ�q�G//��k��`i:T%�c,�� l:��|tL~�nE��f��-�}<������{<E��쯂��C�U��u�����f���7�o�e�/������O����{�΁���<����%g�p�U��p�
�?����V���]j��`/Q���M���4�'�	�a���?x�7%�MTo���/����A�^/a�=�&x��M ��C��
��X�f��r╠�=�*c���M���X���=j�c#u?��cs�_��@0�G�ī�Hq���[��_�[M>R݆��Ŵ����/��{ZR�c��6�}̟�t�s�z4A�x%�jP�G�� K���4E���=8�f��A��*��v��tJ��ۇu��bY�E��o(�
Y��Y\���^nȥLn$n>=�&��T��v�ބo��F���C�~{v��[��E\!�V��ޗI�ә��r�j���o�[K����1�U��E��(.��_���7�'����&=���ú(� �)a��#��v���7���`���H�*L����)Z� �Q��nB��n�D�	��(��gZ���-�J8Z+�ᤨ�t���UJ�4�h�
�q�x`ϟf�L��E�k(
��4�[�~�I%�~�>�\,�&���fyF�Q�W��j�J�����@�7�b��Aj�Ʊ�+�m�o�5l� ���3�!����[x컸�M�׽�]A�Ӱ��L�Td�Ž�.?��6��EL-�1�j<�N�u����ĸn��i-�@[7��I'~�ԤO=oo�>�`��a4ul�&^9��6�m ��[F^x=j�65q�ؓ�^`s���i���*����B�>�I�Q��X�i=��^�Fܨ��C��<�hs$��֖�S�IYI`��=m���4�9@W�$���WU3��ܼ	�fbi��"�~3]bh�S[��4�d���g�Q�0+0�*��l$@k���d�OQ����үE��d8��s�����=�x�\"���9r�Ma�X�uv�������z=�5�7�q~d	i\�∗�2/�c�E�� ,Q�>�zZ�!�VQL�ʧ.��u�{ɾ�pw�E�H/-�aWh�&AV���m���(ya�'���7w�@�̘�(�Ih�Us�h
�����q��A��Fv�x��_|d�K5[�h�L���6��Wl���|X����֨�p� �ؙl �X���w?��p�d�l��*-�p��sĈa�el]��=ǱF�4�|,�B�����IQ�h��Z�4�Tv��@wYĥ�>��� ����0�̝�-�b���Ш7�=:���sB[���N�V擤U�!��
X��0��ȳ�-��f9I-�f�gT%�`u��rkg}�V��F똋"q1�3����Q�ߖnvK�؀��8�U�|A��U��н��]�,BW��C��l~&u�)Tƒ`��j��E�.O���/<���0�Y��;ܳXE1nQ�:F�Ӗ����|�-
>�mK��:�4�0|�� g�jU�2����=b��-���P�I�2T9D�v��̆��h�d��ku�� �CE޾���L/�2�b�@26cE������?��2�G�I������:q4�����X��j ��F��w�ނ;��C�P��>̕��h������ԕ ��z������>M�$F����[Z<ԖtA����Qfwp�.b}��s�������)�O��8&�"�g:��X�|u'��Z�6ߒ�'a�)|3�����������+���c��R�^y��dđ�a���_�o�Hq������/�,l~j�����֨�$���R��z�����9�U[aʧ<>'�� �
:�������M������-����J�d���&�U��ߏ,�����X��v�_�;�iue�j��#�f����l���< ��ɛ*.���Z���l�m��Ї��u�@�e.䥱�H@Jj�������~@��ĳ��%R��!����Ic[�D��H|��tm�J�߰bY7T�x+IeO���	�,Z*�رތ�A6t�/X���� ��"���VE%.st|��	�_��w[T��=G2��L�,B���������5��k=��"ts����{�Z[i��D
n�t%�q*�dX]��\�.�^FD=ZE�7���C�=�����t�JGt��4͗A�Ψ{M�x�1 �xr�#+s�F��׊���$��X�̰���@�wu��.��յ� ��gU��AV9Ϥ�^A䔰V�8Ϙ�� �Ċ ��- 7�'}UO6���=2	Ą5U�����T*��*��}�roF��K���7D��A��BR�f!e�^M�쌥���"�UVE��Z�����t�M~�n��To����r`�>�#)��k�^�)s,�*Mb���'�k֞r��բ7ӯ�;�!(T�xhsf����Feθ1��\S��ǅ��kT���;2�l�P��)@���r�D M���Uq�n�t��³^��!:9ym55��������D�|��"����X�-�^��]�M,�Н�N����лK��^N��1�FIr)x�u�)����������.¯�.�u�S����ޑ�;rx��]�P�j>C�A
8�����@��0�帧t�e��[�Lc����V7���@�寀N3v�N�ނ	��X����5��5	��<���b�Dr���|:�5��{5�N?vk�i����6¦��M��ّ/����GlF���TId3�h��$�U�[αVK1��bu���/���� �,�`���x��1�d�DFR��i[����b�*�_lwI��y� rH�$�R���pͷ]�ū�pL�̜�]\�SRBфG���	��GU}{%̰�)�M�c�LCOq���j��ئ��� �����#AOd8��32
`H��#b��U�j�4PK&�*�5�R���b!�������C�A
-�_U��,�N\ n��4�XM���k^�d�;S�G7R��ۤL(VC{]*(	����A�w��6�ߵ=���Q�*f�T�c�ru�P��f֊1�M�v��n��P6�N��Y�$�L�)�t�<�M��2`Ku�
���d�_T���5o��/�X�H�ж�lGV	�ǜ��E'�曵ߋLEu6�u����w�����O�W�8��ɰ�v���I��e�ou�:j��Ɏ��'��ۺ)+ȡ
R���'ڠǢ:E�m��v��>�'�8�AR�"Ѐ�I~Ԯ�e8�*��sH������H6��g��������i��&�Ϡ�L�'���n��*�߶ZGT�. N%rY���(�����D����jV��a�i�;��,˵��l5$�2�aiخL��sp�u�~����}-lpF����|E��d�;�RI�Ś�x�2x��\<��
Jh��B����G����	��L+?�qk[�,Ĥ�!Kst�},�>c��E�>���Ep�0|���b�"c')Ta�s{�2c��M�Ã.2+i� a�5�^^k.�3��vS�P��H��g��Sq)��������Dn�S,�Y��7 ����]v �zu��gn����X����0�W��ÎR�T�������P���y̇�_�]�3�p�cv�_W od�.����t}�*#��S�'hD����I�����L���'����A�hk��]|�ky n�� �>D+�*2$��6x'�A��G�	�J�G(���6(-�����e��79)��E�*U6��u̻�4�r���-����l�<m���ͪ������և<:ϐ�M��	�M���(^��9_��/I��NmS�j���_][1�\-��!s�-?g����"ʘ3O�V���L���H�������-No�ԽD]?d(�f<�zT8��R/k�J��t'Jn��o��4��͜z�TQx�ۡ���dkPb~O�e�����h��c����u�I��C}��a�_D0��pw_/w�C���K?R��7�u	O�7����l�$-JF��3m�[<�����)�&���woN�,X�Ѹ��>SrR`'xu�(�W_����d�@d�Z
�����,����d-���C�R��8�C��ny	 �;]�h���N�؀P�E����,�l�F��~��꣆�[���z6iy�����i���T�i�� ��\��n$7ԲX_�ߵ��cK��w��+2jz�";)�vw��<�ғ��d�Ej��������q�E�3�� �D�l6�^+�L��vz�p� *�\��d<�>-?�R���Ui����_qD�=���Q�\�2�����6�+p)+�D�� =b�h��y�7�|�����`-
�6�h�(�k�D��|� W�	��QyUQP���br��;���[�+�$�?�c�ڍ��>�a������h������U�O������ڐ�6�'�E<G�T	���RK̏bO��I�&_�a��Q��wqܐ�Ϭ�!��,���"�#_}u�����i���`���5B�|��4}���䯅z���y�1[���VѲ�Y�|���-��cw�w�� Թf�k���).���v�L	c��P��~X�0=V����N1�g��࿋���L�s:�igo��3�����9�7���B�|�Ǐ ��!�(sa�U�����>������`���-�="����;��!2�� ����Ě��3�aa��1�#D�C"-T{��x��	?�b�T�d�<z�]a�@��Xm5hC�����?��Y�W�zpXL���X�H[-�*E�����$���(v �?@�ڱH�2��4+P������2�ӏ��8�nǌ�����SF���Ė�����TႧF0Pn�ǻd�{6N�	�U J�2@78K"��Bt�?a9,Lo*�{B�����Pgc1n�2{�'6GK�w����r'nV9g���|.g)ܸT�Iy�
��[��7z������N[1 �J挴x( �e6����Op"�A_k����1pM�1��0Wm���ԔhUˎ̜J�q�L<r~�>��%|��Ʌb��B�Ct�֜0]B[^��J�@ʅ���Ɛ1��n�*.w<��鲽Q`�3.���>?�����c��nq��>H�P;�i�f��<W��*�l�ܤ}��_D�yY0��[bD�VO���o�,�n�0��C�>����26�xfwL�T��1��W�����^V��]6s�ͭ���jv?:mm��`��$�PB�����J���X0�2IU�n�.,d���w�3���/GFK�P�Ħ2F��A�+���o[wA�u�,�0�X0 �R{ \�b���l� {-���q���5��C�#a�
�j���Cx�|���'f�+%�1�=���-�T�&H�B��B����Wx9,�_�����\��޾��.IC?C�%ÐCC_�ѴS���`Ta����1�+݁�pSacz�#�W�Ůe����ex79��Ĩ�$�R/s�W�o��q�pW<S����Q#(N�ߒ���c�w�n��߷A���qf�m�W�'$j4�v�`T�?9U���]Ʌz	���f�����G��D�u��֐��������K�б�`��6d,I����X?<����`��x��Ͳ��)�Χ��	�6;=�5���)�<�����0E5@��0���
��K
n�E&�w�#� ���o��[���׆hFdH3�َ�o� e�!�O�ސ�"���U��q�V{���W�׫=���	ܧN�Q�~�{�����܎��V'����B>�Ҍ:2!�N\�� ����ulpܪ4ևgXܪV�[�d�UanFuj�$���÷�D 0:rK��{�!���~O����p
�$1����u�v�Z����z�HfC�I>ѥ3 ���{�v�:W��(�Z��=UX�i��7@�L��f.L�DG�ՙLr)I�p�q��.�Zc�D��5� `�.�;��>��C/�m��I�&h܌�<_�i���َnA��<G���J��Қ`os$Յny�թ)DO���tjH:f�^�X�[��TRL�	:��4�x�W��ʹL@U���e�Z�zFxǓp�NG�A#+��e٫-�$j3J�b�*�mc���x�ܺ��8�Qk׸4���|g���%������K�h7�UT*rV&�Q��	x�ȯY#YY�]�u���6t���8�OD���#��s��DY����"��M���}�c9�
��-�,�>��{�	�c��+��73�IAͭ�@�G���u>���r�Y]r�'���ʓ_S���W�
����:�Po�g"�cR�^i�MYO���n��mwej�R�Gp�
]}Hg�i'��lD�i�LxG��f�҂W�ON���h�п��x�x�_*�R8;��ﵚ���7�y"�%��]��8�$?�u���W�HF����>$�YY�脣]�^.� 0��{��Y�kt!�p�-�����7�����k8g��E��6���<��(��AַLO�3�9}ڇ��\P�������4ik�%�����ɥ��d��s����5�蜄�����	;��f���>�v�L�/7�IL⶛Ee�C��}͗���M�X���xH�1��Mr��!K�ϘވLg��yv�Xo�U�{�#�g����n����t�$��+!%؝�m}P��B}ɓuO Kps����)<�m��,�ȏ��Z1(D���[Ae0Q:c��<Ȭ�ѷd�똂(��O��7;��TfW��[$��
"Z��=0>5�� e(��ixН�:�����ɽG���a���<�2ю**�۬�g���Ă��|gт��l�&9�:;j�Oh�~k$�xKkz�򋮋��ME�kdW�P���j_3��2�jÅl�SHy�i�>P[�/1D�,p�P�A+�K��!LgD��P�O٢c�a�1�@��F+���4-�0��M�o"��0�\I�_u�� z����?0�c ?ף,E*P��,$��b��։���+�q6�L����煟Ao�eĂ��E3T
X s�ְ���`{BJ�E|[L_��ɠk��:l��J����^>�|>vi������Z;uu�[D�^�Ϧ�\��8��<��.2�+%�N�k�D������O�4�p��4Nqt�Y�����d��3��Q~XA�O��Ѻ�Kd��_% �z���6] )a~b��ONz������y
ocLq�(�ot��[�]�'.�6R���Kq��l�;���}��2wK�e}-K�]Y�=���w��U�~q}E���2܇@���
���z��TT�J�g�E+pL�xS(��]0�f�/*�����:���XǗj�$���ҕ����&�:v����2���?'�%�Ѐ&��/(}d.�ћk�!)��0���|p�+���C�w=D�ֵ��z^b҄�/FV\�y��K1�^5�ꋶ)d���b@ ~H	�&�����0����d��9�k�8����З�E�����=+D�e�O=�7Yg̦��O��(��aI��l�,����r�;�Y�MG �����|�l&��^�"�� 	� �|輪�דa>l���t�m7u;뾆��U�7����Z�~��/�`�#�,�C�0HW7��1<f��;��g�􂜧T�R���e�iJ>���הb$�k��o�=����C���Cf@�ք�K�{�G�ko1�h�Z�_S���� �����?�\�M#�h�5����<ST���,{N��/f}x���CV�����?8}��!@v3W ]^u߻��Ӥy�r[�.�R���1��ǅY��T,�>�z����3Ƒ]��7����8�v�|~thW��vW�{7|��6zL���[z�ݴU?�I	��P��n�ԈS�:}��N�i�~�W�X*�R[+Zn��,;3���蕟�B3����������Lԣ��[e��:�&T&u����IDRH�ԼR.�{�+�bG5��Xsϳ��t��#m��ǔ��ۼ�t�8��{�Y��=���&
X�pN/0Fek�I}���l^L!�$�V�d�M�3'���d�$Ƶ!k�����b �,�:g�$�$So�Bǣߴ��v���a������u:�xG <�nD^SC^��]�H�?`�<��M��[�KFZR{�ݠ�4��B�˵Iu"k��\�U�.�?�
he"��0+yS�AȌ�ǥbC�ӲJ�1)(�%c���f�j_j�y�rM�]G��?�&s8�"LO� ��U��o;�)����G��7�O>l�AW�/r�]85�^h���\�V[���\�5A0]u�.ʿ��£]�i��XĂ�=|I!�ڎ��27u�C%����UCT����e�>�n<�γ6�)��D�,�o1x�_�Cɺ�h�W�)�����j�$��#�r��(�L�l�a�n�d���:"io�
��a�7c����N�jOzZC�()��k,�A�G���cWι�Tq�����M�H6����n;@�탃�tA�)���޸��fD�������2y���O����H^/70bS0k��}iFW��N�5�W�u��U���Ӫ��.
R�o���]�@�7iW��W���D>��I��� W3��ǆ<X+Qxgm�I�Rޫ��h�z�v?l���Z�؝�1����U����2z�_���ۓV���2��]"r�,��>} �QZWZ���[�I���%�ʧ��i��ET��9{_�.a�}��8�!���P�%��ie���
��&��&1��@���zL�p�Z�ց�7������jM�@�>]��l�V��B�'��'0z��J�j�5HB�� w��]�@��
D��<�����Q�d5�v��h�/쇌�n\�6ݷ��3�ڡD
RN�"Nmy�(�0'&�д�>��aZ��[xr pIc�!���KlN۴��zMO�L��
�;�E���?�;5Fh�h}��0eO�������0���í�e��|����x�Ԯ��b��WƄ���Լ��W��Ԭ��D��E�X�To�{-;;;�a悅TrϞ��C{�oA��ie|�]����1#��a��oMK������}�$ݙS ��qd^~����s��b�_���w�l�c��*�l�,�U����g��p�E,�SL���7�O|'ײ ���{NZ�7�A���5����d���5΂6-̢.�x�葉�~�\��T�'�:>&��OB�x̳%V��=�?���H���U����"� !��Ӑ��i�%8�(ns�ՍT�ȍ��PE�� �|�z��g�ǅ,d�M��R�ӹ�����ӹ�{���O)�ɇQkp3�bX��� �O:|C�J����<�m���DCF�܄R�7�N *6Ԭ_%�|�X]����7��@�!~?R�J�'�����,�����ζ��HDԳ�+^8��.m@ݩS,@��P�9t�����k�Z�~����Y�d�KrD�u�v���n1	V��������������S���'Y�j�X����'�3�~��{Gۉ�D;��&�\"uN&u�'�K�8s�l��]�ՅP��w��̍��U0������ �$�t��������D�r5v [�rA粈��Ȇ��.{�/$K��oN<��X���d��gΥ|l��S��`䋢1��T�O-6Gk������(;���(�a?
.�P��I�gx!��yw�XPӐ�4�WCe�s��dňV�sy��/2��B�s�'ѓ���	�N2"9�k^���^=���)� �IpE�`L��ۅ���E�<'yD�ҷ�<Ҫ�uz�ӌ��&I/;�j)�/��3��k"l6 i+�/�8�!�\�U��J��=/��؝5��6�Y=]k��:���0�dF>æ��8�����eŤI�GLʧ��k��Ň�B_'c���A�!�q6��{Z_J!���V�ō���KTri^F���X�~�p�ˢgOg����4�Q�D�� Ltt�`q{�-\ےVo�g?=Im�?���:�ļX97�\|���J�T�F/o�|�b���~b��GrG8�l�
�
sY6�. �^z�Vz]1yu���ۻh��=L~:O&�����P3���ȳ��_D0~D�!���k�����g�j��\�I��hwҹ��}��5��;�^|i�X}�^���X�~D؉�0Ƥ}ap��{���ҷL;Y_�s����9T��J��7�0p�F��]�?�ة1�`�bϵ�[�w��D��c+:l��͙h�S��T2��,� )W�q@�]�QW����]���_o�(��'k��w�ѳ;Z�fC-�v�����_zF5\����=[M=}K�gKb�ݪ3�����<*�,���x<I�P>�2�9s�Dn�x�����dsH�(c	�x��j��Dm2�
����ޠ� ��!]P�
�)�֎��G����_\@�C���i�Q��XtUt�GF�7��I5;����ty���b�5���O!���!��R�w�5ے�T �H�c�y�U����kca�o1�l|�H0X�����~�@i�L�EK���?���J�����e��n衘Y��p�1B�s8��=(��	0�&��|`�,#�p``���@�{���h��&O�k?/�v������0v"�����_��1�Y�/�7?U*��)*�?q�=q�b^2o�І�`j����q��~cK�ݱ�!"/�ǀvC&��\��[�X{ ���W%VX�9:AN��oI79���nj/(�� ۨ�s�tS�>����R����1�0�&.h�X<&p���
�����<�0�}����8x�L���vJ p��l[�L�U Afh"i��^W#�~ޱ�������&Xbv��~�؎kNM�����ۓ��p)��(L���`5�y�����1�z�-hӅ`�N����8taD��Vu�f���M��.�C��S	�J]3�Cs�n�;
�V5E�� �^���<�H����<U@ج@m`��f�HC��&�
���2`e�}G�F�#d�.g佌҇n
z��r1�}#|#��=�1F�ͶU�6�ܫ_�w�!XL�xTb�^�8����7��6��5 �"�Y?�w�����W^�.+O}8D��ųC��:
E�ڽ]��0��HL�*���e�)l���aK-���Pn�"���#�T߰9�Q��'q�`�;%\)Y_j_�˗0�Qߖ���p3�k*��:�>��WP묬� H:�3�a�~o&7��)8���p�M�g���r͌����(�]��"�*�.@���� �C:�6)��A*6g�	e�u��b�^�ǎ �I���2/�Q������w�0WnB�-�XaA�wK������VP�RR�/�C�p�w�v�ӺPEb�h^�
e��ڶٵ�U����ssH4��G��B���VW�(�O�y*O��\����HR��W������.]mT��w�=�*�y����N��m���y�ֶr���WY�)��J'�Ƴ΋d��.6�s��`f�ִ���b�
�[D]��QHY6W'E!;U][v�N�U�Z����'�]P�tA����e��ᾴ!$HF��T�:�P?	��9�����0��߽����<-H������
"�ԧvה�s͂����o׾a��H�lk�R�F���5t$�@��9	��(_n��mT>��5���AUt�!;U 8��<bxƷڝ�UҌzŠ!�߷�2���t�	��,��6 KTx���3�ȯJʱׁ2ZR=.Wc��͟�e�<<�9[i�ŕWv���'�`�<�Z�'��U>��v��l���!��"��6+�;3���Eh�ӎh�Dm�!�����_/���-Ϻ��X��F&�sQz��Wa
5�����t���eI~fd"(�s�+
�牀�C\��"�w�?$�H=t���\Ȩ����T^$;\sf�;'HL�|n+Y(W����|Q��___�6��� �����jƚg�ęb���Ar���uq�ů�z�N�s��j<�VU�n�\�av��uiA�+����fs���${
/<��zj"VQ�χȬ�U������ʍk^	{���p�����9�7�����5D#3�x�f�=�Ov�G_�GA��p� ����7��Q�B�h��<�~-ԁnxo{L���j�7̉OOr��)���7"��=�9�4,)h1���eD�⧄r�'�PO��·��;޸�M�j��`8ױ��~}{��ɭ`��% �!�m�F���4Q��g��U�2�o$f�	��Zy9�ܞT��P���w!Y��E-J�W o{'Ե��.#8ө7c�dDZ1�#�d�3�U���֘@b�Ok�?�-�`�RV�7<��m����gS��z��	A�h�>2�k��BwU�.c�	#���w��Ga��J�}������g�)�,K>�i���޲套
	����7���e���C��� �:R�orM�e��w�
ʻC�%�����޹���#E8�ql�0m	er�ގd��fM�N�� �u9��K�c'XD�����N�+���G-���T3�����i�	<|���e��7��nS4l��.�W�A����_#�l.-�κ�~�l���bn\�/����/�-4�X
�"P����֦a��a	�Hf_�~��O�q�vl@��jH��q��y'߰{CY=��ns9�qr��(������št�QX�}A���
�l�l�����P�&�K�ѓ�S������R�?=�$ͩ^��s�y��	��_�"��l���P���a]`|��*�{�����e�\��G�>��LSi0g�]/��~�
-�|mG,O����,ӹ8�vL}n�bB�CIP�i���g"��À$͕� >H芼�{|мZ�	�K�=;~�9��+���	T�0 (���׀ǀΎ��i�e��o6�����ZN/28(�OJ��#K��Q�q� *j���NILX����.�����yb�pm�^U��1a9��U��~��1�]yU5��3m$a%�8@�o��<��BɆ�1�	d!$�-�/
����W�Y�ڃ�;?��9�#KM�|�|"B*;��/��B�a�I]��Ec�S�;��
&�����Kօ=�Qr"�������+n?�JjH��;�|�,�4�WyD��76>�m��򹾬v����Ș�~^�r�o\�od�l�����@�&9"|�>ਐ��aH�1b�n�,��	�j[����wT���Ϟ�b� �L0m�|V'-��4�îiZ`d�ډ�R�R�(�l 8-�����ߠ�/&�|��e$���ḀcWdI����´�J[j�&e�W#��j�)�E�4]��;��|.���]J*DI��,�jȭ��s��9py�C��_���mE'�� 5��|�m6	���L�U&U΂\�<�	���10 I�X�>�Hu�[WsP�Uo��g}U��_�Bxr-���e�?")}�����E�b�{��m);�^v�m��F�]p=N�ly�UE�1��q���N}����U�͠�{�i���g�YI�#��X�G��ё͒�Iʸ��`[�Iw������$��l��-tz������-}�6��f�	ӑ�!�ӃK0���~/��2����4�`��.z�U�*�/�m͞�zz�FY�����4D���	'Fe�
�Qz&��eS�_=��U}���m�kt�z9���M��(Te'� ���.�('�?�p�$��'���e�4h�>v�98r]� ��ه�E�"ب3]$��uo~��b՘̽�~x�G�r�x}?�Y��L,W��l���W���Jۣ�J Q9�d��@�ڄ��j���?!��w��7��ވL5y�D��-���+�z�!���?���Ϲ��^��K�f�� ��
�^D�t�����e���<����G�.V=Ee���S�JV���/�����x��Ȗ��R'�?n�.�8��jB1�ø�����x��٫�QK�0�6�XCw�j��+{	�'`�	��6@,���;#W��_�m�q��ZԔ��;�� ɱT�2�
�̥+�ܧ��-�nSCzo[�U>��!w*������B���RqeQЬ�FX�y�,�	�ը$/��GI��gw}4�%b������j|��Ka?6��Q�A��U�}cwZ�S�ZU�lP���F�"�&z$�!�`f�l�Olz�+�Hz�s�+&��2�|\�6q����5�.䊵Q�r��`8��]E�ށ �����$��1C���N8.5\���*�]�B��?����Q�i�I �63ګ��ML:��Υ9U�>����-wSno,�L��e7{��h����
`�ΗY����n��`A�RG�ukuV^ڵ%��u��������b�s��/�\8?��7;
�n��#�V�Q�-,��3�E�E�T�����W5V	�^ymk葥�ƅ��m*s��m崶D�B�@�����Z�<��Ԃ>Y��7�GJ�Iv l%M��Z �a��s	�#�{���
j`�A4�O`�ߖ�؃��h6q8��%��"� $�5���(	p�lj�=ӄKu�o��?+�'!�L�;GZ�A�h�!kv`��zL@$�P$�Y-��.��d]�O��yb����
�L�[z��f�8)�U�7�����k�)�9	ٲ'�[����ض��sLP�l�;���8�t�Kj��%e�ة��=�x��a�ѩ��4�)FG�g�(Wԋ#���4_{��WU-��Z����]YUj|�7�;�ӇZ�tg�G�K��uo-�܉�ͼzҰo�*��x���Nk�!���P��'f�w�
�斒�)�v���a�����#=
��U��әl�J��2z;���ܶ�[����@zz�薒Z� ��1y)��H��R�~�}�I#��A���F���̬��	~�\x	�Eo���z������٨�[�@c���dVT�^��A��Ѐ��:���iB��>����,�7��� �y�8�����i�@M���(�������k���?�	z�|�sFX38�go��S�aUh@���d^�Э�T�ϊ:g� ������o�z�mR���`�D���2�V����<��H۪A^�h�x��b����$���x&�=�V�[�F�FNQ��w���qX*
�5V�����5�ǐ��
/:|(�0�͛ N�I�K9����ƷA���,�ɖa�a�!Q����U�X��ba B�u�k�޷�'�+��F��9��c�Jkh<����� 
%#�b�O Holz��oy��W��Ѹ�s�y�k�ч"��ͽ�3ñ�v��UZuQN�c͖���o��c�_&l�F�HMi9Z&]�!���V���
;�~���3�P�q0F��m�y��B�ĳ#��~Շ�85�������b���yo�~�۠��Zn j�	�\�V��GI$$��k�_tP�Z]ZFx�n�(�7���Z��=b�i^�$�K����Ҍp�Ն�O��X-��֖��vT���(�Mca���'����۴�8^��QD]pn�}�-h%�L�J�WC���dAD	�u�c[�Ti��hǫfv�B�}饝�m��������`$!� s�$"��5X��ϕ>8���9��(Q��E�DY�����bA	�A�@�T�3��*#bn���f���H�st�~ᲅ�D�`"}ԏV�� s�a��`�jw��t��0vq�w��F������1^�W��:��P�B��*@��2Z�t�����q�*�B�Fc���ۀ��V�	ŗ�x���Ft�NN?7�L�p��s���H��P�C�k!Ⱥ�#ě���dI�!��>3�KW�z��,@X�A|tQd.��|��Ov!5Ϲ����C��x�D�t.�����Ӵ��ҍ��ٴ��+Ù09��]���o�Ց�W�y*�o4�)UG��,Yu�4�
(WwB�r��2���R�3�{�K\�UK�R����P �R��ϩUCQf�����5��*�=�W��^���-���OV��#�
Crΐ�=��^��â�}+�~��`�[�Z����[8^i��Gt����wu��f��G {�t�$^��v5r�$�췂��
�ﴚa�J��;���ɃE��;��]W���}�hʭ(� ������WW6�s��":�.�0�9K�k�A�s��pvp9�X�8�"�y=�Pz�-����#V5�ɷ�O���O��{��L�������A����WT5�!�_�o�4�f<�s �kP�]��}��*N��@�c n~b����K��� z�!za��+�ý%3{�{�'F2��i�,Џ�ɔ�,���������&���1�~�{|�Z���A^��D}N��2���ߴ�,��f�>���FpYx�?B>�3?�R�� U^>�=-�V�}$7@^���Z�|�����0d�T֎�¢�M�Pc�F5F�.#F��8�b�e�l~K6 /�L5�j�}ZG�S�a���
:���Q�Q���Mh���;-��:�HD�� ��^4�U��(3�[�|Zϭ�yT$Oy^ʸ��<M��h�LX����.=K2qs�n �D�;Ej~hkQ��Q5d`����v���V�[�ԋt��#Rp@���n6�n�xȷݒY�)Hr�6�1e��~�i���sg���I<Ġv�/�A�����0qw�@�bRB��h� �-���E��s!��&DB�ɸ����5��v����!�4��v�S�vi�/�9�9�>M�s-���}l��f�=`��s1��wD�@���)����*�VC��ȝȦ�,��C)��Z��c��di�>�z#�m�nn,+�]2�Y�6��뵤���R�?lu^�7�����%�Ѷ�5?@V>� ��C�y&9�T��]��\�Hg����o	[�y����sDj
{�yՓՌ_�CΪ�n�K�m����Hqm�p��3̦G��m)������iPCQ���ݓ�fz%Q��ݠla����+đn��Z�=��ϣ��t'xA���	��cA+���"��Ɲ�]�2�W��=����Ur��7�����kə�4)���C�ݨp�7�I�GTK>��g�}F�p(ǡ\���y�nռ��~z.y�!��SG�(i�;P��*�eQb�J�e���B���b��><pÕ��.=�̠h���m�Pq��p�ot���o��]7h(w��-��9��A,���w�)ɉ�W=n��9[�yR�WX��X���>
���#�4��!)�k����k����o�R�����Ыk�����l@�h�>�0�L�B�U'�t��h;Ʀ�!����������{6J�/��tF���C�V��w"�)�cs3��./�8{�������>�尙͸b\3*��N�|���h���.��h�]AE��<�_3�
�.�SSq�����-��A���j�,�s-=�����_W7'��{�[o���H��:~8<��{^}7��{���rɁng�!"�m�I�r?���Kw_D��E��y��(��s��#����^��(���������0�?�4
Ŷ�'�.5<!\��|׍e�]9(7#�B�H� ��ڭg:�K���"Cc�ƏTE��4��܆�c��S7�OR�#nnW��-*�G)�:10�3�7��Q�$���(*��8ʶ�M���;a��"[�,i̡�z�F�>�2�ʂ��Mu����xu���%Ml6�;9�4����Uz��~�A���r�A�`��h�d�M�r�[}C�K����B��-~~�F�y�-��ȟ�[ڻ
��L>N�f���Ȯ\������;z��1��)��x�-�r�����Y��	���]��t�L⟼OӨ)=Аy�̈��?��mg�˒�]*�g�nS��!�^|0��=�o�E���=M�lS3I1�?����`��*k��KM�aĺ[9�sb�����#r8��j\���JEE�Ҋ���t��'�Y�p����z�fd�̞ӌ�1��o����y�lR<�P����`B_�Uğ\�N�B2���@U#���ؖ1�о�2>f������;xb���T%=��ϘVVb�]O�0FT9����]�+�E�F=8mk��<X�P)tv@�*�FX�����'�����!�B�Ώ��#�X�>�j���9*KDi���f"z�!s�T�g6�=C@B� =ۂ&wI������&º^��h�	ށ��H�� 2�r_��Χ� \!B���i������;10Ҫ��^yY������ΰt�Ux���B+�,�Q�<�6\h����?��+���I7���+�������n�(��y�7d%4)3�<*{�j��_A���=�Y���'�?��7�ß�l`-�g�.O�vӷF\��y[δ:		^������*��O���	m��\���s�;!V9���4:�����I�M�&a����9��)��o����<���L����b]�,����P���z[[M�`e]�/��o����򝷧e�eg�m���gU�k=��9�ӘO��z��;J�vRP�^J�	�I:Vӈ���T#���vE�y�0�@�'d���U�J�N�V���G~����I��/�F+�-�+��\���4Q?��YLQ䰤T�z"$$�Ǟv���Q��*����B��(u���<ߪ��}{���������L'����U��1�^���@�W��ގ��B����R�}�+/�	)�E2�1 �}N'�C� �A�Ç��#N��z>l�%���!8<�d#ųH'T��9	��O���α�y��uݡ`����u}=�L}d�����}X����us���3:�:]���R(C�6����Oŵ��k���t6��Rѧ�0�BQ��]*�𳾲��A���{�i��QZ�jClG�?Mn�Y*_Z`��z��.���MW�c�l���Fi��{�+�I�9_���.^j�Ы^1P���f�CU�"T��4$6U����k'W��w��1n��S2 ??1@��&�W�ͅ��kL�O��A��j:�#��uS�dRā03���/�nW���Z�I*�{��9Zn���ʌػD�i�wvl��m�����v�X�{��&��J��Okz�y��}�#%d϶���f���D�B� 	�8��c��G	���Y�b{��{1�m�vYR����lN����M�:}.�f�/d�g�F���A�dY��|ɻ�b&<�ӄd�����hK+p�D�Kug�9�Ȧ��TfF�2�#;�F��M��ߑ ��@d���Zd!�2.K�}���z�0���w�҇!���J�<��������{�Dki��?��Yr�s��~n�Os�ǝ��[�V�����<���g'}RKa�\��YS�llϟV'!	Y&�L o˻��^����:�M��^;��f�>ҏ�>�>�:�Rd8>��-��@�ڭ|��`G�����vb����C����рli���]������H9)5o>�T��S�d���h�C8���q6���l
}id''r���h�S���t���>�C+-�.E����.�=\x��S���/G|іУdw���l8 ��'�K�1���9�����.q&�Ie�:�ؐ�h ��
�������6`������c�l���O�M��
6o�})|U]Xl��M��=�X�P�K�uP��#�:졄�[���2��h��S��Ə)�/^�/0Ϝ���z��īBiȏ�8� �.�z1����0[Vd3��[
򽬩���>��Y)#�H�_�&��̋{��I��2 [@L]փUTDE�l����E�SN�p��@�0����[I.n��*=��	�5'���6_l�t��@]Q^J,�QѤ���Am�z�[nq�G�T$ەU�tou���\��Ӌが/(V�H!N:T%�;Bv�n]��{��d��b�W�h���qS� �e���ښJ���G ɝ��`��F(o^�(#]\=�fF�	  5�ZɜX�~~���%�*�H� 9����1_��������EW|h!�j	�n5�r�"�-
l���v�`k�,�F�,*�4IԵ�h�y����SsJ�E��/��]�3g�i�O�\����= ݀W
�u߷�([Og5d���O����*]��+����g+�*P��xh=n@��H�^A���i��:r>j{����t��8�� ��y�3��*�W2?��h���1RMG\�'�4��Nl���y�))� y�t7a�S��M���g��Nc~��5�1��e�< �X0�Ә�]�����}�sup>L��|�&yXl��*
5�>�
	%زI���wط�n�j6)�@jɹ���,s�?�����CM��T�V�#>��av�#8O���}�U�%�ݎѮ	����U�6������[Q�g�5l�d�`�[�u���_tNC�2N�UX<�0B�'&����"����K�"�����d�v�m���i�J����#6@���OT̓QQ~P�N�W��x��%7g4��w��#i����>�!5P����[�Dj�`s@���G7��Wec������)���ˌ&����ti��pbhל��+�Xj<!�b!f/<�u�����O�R��G*�$�ݞ$��Si^[s�$�����������\z��&u��`1�ZH��9�AV�4�֑���K/�/2x�`L�EI��ɿ���U��e�#�~u�~t�s�:v#mLWLȖ��{���G2�`�ӹ���=C�����>�Y����[$�c��V�����TI�3�+l]P>y�B���Ojbix8��a�W41�?�[$����M0�=7�ר��a>�c��D;@z��_���lx\Ŕs*q����&O��VȘT��7�tn�^�g��Ja�GF���_�ݷ/[�6�ʅ���y� ռԢ�M�w�q� <��(��]�i^���P��C���VW�.�_%�N��� ��{�j�5C��.98�u��Qw	vI9N/����$>}{{U^�U|UKIт5O@i�>��F����BL)3]f���y�j+u���w�9ї_Ԑ��$��,�H�9�?X�� �Bݾ�`�;ɺ��s�.@�vaZ���E�C�l��sb�})��Fw]��G
S����Y��~�֫
W0�������߬�7���)L���)�a#�(�|��Irl������jI����q�_�sǖ:і+������_�8�hD�H�H����6sR+k�Aen	�{<�՞?2�����V*I�����^��Mm"�//X�p�4gk����/����8\���l�\^��ZQP�1��=	����ϫP�3"8U������h������ҥ췔ֶܼ� ����ˀ{̈��]B���A����I����,��T��[Q�"2�X�^�l�������� ���n�5�b���t`E	�y~���̦`�Ƿ	����%�Rk��nv��( h�Kj���ڇ���Y�e��4�g�f��3�Ǘ�L��y7�c$��oؒ{��w������A�� �J[��I2ӭ��Hb�	z+m�fI�矐�Uc��H	���	h��Q��vc��ð*�QI7K�Ɖ��8\�? =�u%q+�ϝ'������z�,�!�������F&��8�pL�خt�"�{(On�������:� ז]��+8�G�ݫQ��1r)������G;]"๽ՙƪ��Od���UL7��&��&7�Ƕ�/�Y�'yy�]�'��7��.��+��[�XӪ��]{j �{X4�M�v��s�-Q�u��L�f�欂�1���B0y�8�	J�n����e��e��59�l��f-o�\��ތ��NB(���'>M%��7��Ok���ƪ�;�|+&_���˿$d#�HL���'k�a���BM�+T�����iԺ�D�m�J�)M��S*�(�"����	�j�k������~�c�݇R��i �n�%����7�dػ��?bԡ��ǃ�}�<&�2
�uvi됁IjUr��Rv ��K4�^���Xgv쥛m�1N�*��i�:�Z.�S�(0q6��Cjr��t;~b ܻ� 鱻àbS�����^Ue)��JUZ$pA2�����$0A�������-���y)t:exׅSb�{�x����T�-1�!a�_���S�����j�hKFl޲��|�|N+��L?�B<t꫏6V.�Ш2F��Y������n��l"w>im+�+��=�s��ĸ�e�5-�b3DK/�A��_��Tപ.+W�$8e-ߏ8,)Wua��_��'&���C]Ц�W�XЧ��圉��T쪋[/��p��D+��f���6PwG�A]���X��O�������S����T�[$��﹡FD(��hr���d�[��1�j�"0 �OR�v���ڋ�'�uk�XVw+O���U��G�B�X�xo������.���.X�r.��^��sJ��S��YA'�nӰW��.�Es������Q��ܷ͵�kāt�₻,����$����2�E�����Br��/k��_��8�.ҵ5"��C%����a���kd��j\#
b�Y�>@Y�e�EF�$�K,i���Z��"�φ�Y�+�m�� ����HbY�EQ��E�(�]�&��mh`(Uy|E>��
�3J��A� �B����	�q�y�|�r�ސ^�F�j'kd��!يD�?5)v�y� >nඬ;r�����~KB"��&A�.^�S���<�@��YZV��<<�lG�a_*ڿ��=F��rйy��b�(邻��
�cG���|�'��[�~�F6E��ťxET����Q\���2;���Bd��5]z�2���oA�C�O��{�g�h�Wc�G�F�׾�D�L2�m-0ղ���O�� o�|�2PW�,��џ�q�A���������9v2 ��I�9t��N�%���m���_�BK��׊" �V�����<�	1��������=9�@��� j���,��*)�Tc�Hr�y��s��.q��t�nm��M�>t1x�Z 
Us��5w=�o)T����"
'�/�[*��bi���@�c"�o��a��{q$j|*ڪÚ/�{1 �/����0{��To�|Η�<昮�p��v��(2Gc?>+�$�,{s���$˩�,����O_�)0�{#���Dm�	hH����2��'waK����/�r4�O�0�@_=���Z��=�r��G�zl�Q�'�{�z/^�E�'+��Ֆ5ᾚ����j/�n��A��L�@��s�Z���橹&m��E{�gv�ga�IbG?�[�EA�m�嶈%��#S����Jb�<FWJd
p���%S��w"�~�
h8�D!-l�'����AO��\��q4R�qQ7��>�y{��h s�^*V�����>���8��?���V�v7^����L֌�|�� 9e��t����%Z-����v�e�l����x*���E�����po������J����pHށ�X}����\?��=�ŵf�l���Q��^�F�:��:����(����v�K�g�3F�_`5Qz�T�n�o��
�n�����B���|�i��@&;)��>�ک~�`��BH8�K�x�O����q�V�%�kƧ�nv��Um���0o�f�W��$�僆^����N�h��YCL��&UĆ�N��:\�%&��{1��܁/߰v�3�{�O�2!2�n{!�&����I]���\)���p�M#YjbD�����؏Kى uR֨�&y�;�Х��7�J`aW]DH��|c�ݦ���.�z�!c�A�y)�d�a�{�M*�ڷ�,�G&�	��_���Q]��Y�V[�9���k�0��%������]��C�d�����I8���+������_c��s��~*#����)�u4 �64��\֑h`!u`Z���f[��t���w�B��,�V�-��X#�c�$�,
]�<c8�
�������1r��AP�Dz���_b� �$�EYcz��o(� �%�#���B{�;n�#Fn�hc@�Ua��Z��?� �CS[C��~*cm���f0�+��QDN�1 �K���F�iմew��-z���0��ws���2F�ϕ^�ެN<�r���&��뀃���L�8h��F4��(��Or�(��q�L}�,c�.,ƾݍ���HS����=�-
j�@��~|a�5��tO8#v�M��%r�2����O�
��*'���b����{5�?��#�R�H����]�A҉OC��e\����+�[��4Q���iVX���(n�]ޭ�V^�-A�;�j>�+�=u9�������>�)n`܁�kAbO��bD{�Z�Rj�/̓ल$�5pSE�xƻ'�@�~G����I����� @j���S|ƄQ���[�Y9˻]8�VA��!?k?�{�ʰϜ�$4��<���r��S 3�E�ߍ"�ܚ�	���ي?���6:+�`C`;	����*�Ԇw+���'sQh�l���Q�<�l���T�^^���J�]c��*��(t	aV��7��'j�y�-� �cM<�T��_F�˜xO�Bf�ӃMO ���5H��&B��c:� �&�B�'+�B��p�T�d�ϸ��dtP���u$�Cu��e`N�\q��F���M�� +���e��1 ��u�@��^\�a^���X��4�#qH�`�H<'�б4��4��K�?(�����"7� d`����h�Q���9��O�!О��|��x:���I���ϧ��S7rd�t�Yz�ϯk.܅	ɌZ�ut����)�I������dR�YJs}����*�h7V�Gp�M��q����,Ag��MЈ�ݱPĽ���e��M���w}~=��I8t�͎T��L5v���֞�kѪE�[�:a��Fw�J�������7u���/&�$��b��["J2G�v'V-F��S�R2��̮}��Z�	*r��D��u|sW=ҡ�&�W4� B�HI������w� @�g��&��p
&W@È;�d����[��e:���Ȃ�U��# (�dn�L� Q��O�,Z�p	����S���i\�r\���t~+��d�?���q� �W�9̡(/1P#�^v���k$�o�:C�V��
�O�R(����|�������i9	���MX1����z�d�2A%{9d1��*b�2�+v����C2���o�)h��n���i?H��"�I*A��K�R�����ȕ���:�7����D��X�����]=�]q-_Lv�aB���,�8m6�9|�>TT�vМ�Vμ�>���d|O.�u[Mq#i=:��(�z���>��矺�&	��~���'`��D�L�~��n/�5��t���ϓ�����O��5�5��"=��=�bK� ��u�`� �p��X�6�P�uW�I�N�&�B[Ԗ�����s�%��׬��@õA��K����ǯ���A%o9�ݑ��I�+��r����l9�(N&����j_�$Q�����0X
�I) �5Ұ&��&��m�r
� �\-����_��/GfF:��{�\3t����@�t��q.c�R�U1�0�B� 3��P�Y]�-��M~yK t�� �N���>�{� 2�9�����?Mq6��wt	��QT�4�;؞Zk#}e�m��Sgr
�����xo-Z��&[��X�Dnh�	��w�Įhp�������ڷ5�g(��z=�ݼ���$Z��e�v:^����U����+�C9�w����L��L;����y�jn�S(�%����>e�S�!�)Y+?SY������ļ�=���ľ	����/�[�&1����i;���8�έ���|ǄO�P ��P~��ئ��9��ȪWO��� ���m�0��ðg������������"x g���P;�o%�����U���-��5��Eg��"�Σ�n�m��چ���^�6�[`���UJ��Ap\4I2��]fq�FlJ7��A��/��.�4���$�`��F���)��9x�	�/w_$)���0(g�Y�
��N�6(l�.��)w�	w�j�s���Sω�EC_�:#�[�_�� >}�/�[3!ײ�Է(��u�@�J�r<�o��q#݌}����exY_���H���%6~<�j��2�R<��ʡ�$��m5{�S��m(��@�;e�H����Z���!�%^ƣhAF4Y�eZ��Q�I�4�D���/Lcb�^$/�J�R�$�m)�9Ї�
��Ғsw�o�˃�)���G�b���<\�JV�-�?x�p)�x93`����ͱ5 ]��C@h\��'�����e�l�x����0����w)6 x&=�����S��Y��9t��R� EG�p���?3"h�HO����k}��ƃ�́Í�/����Ba1X����q�.��C�̌4*�g�8iu0I��J�t>
d+�e)x8����0�����n�x..�����cq���v5}�3�;��	�nD8*���J�>'Ыn%�>�,��tB�p�V�-R�"���V�[�Y-�-ly;F�^���J�?mJ�	�ိ��4�%��[0d�+�WV�0�!X�ږ����o]����; 8�M�a�Lo�x��I����)�X���Z����	��&���4l/�ql��9�ߋ|���� -~f��t�cQ:6}gg�0g�^��r����.b<o����~!nʑ_�����@~u���M#X^�>:/!�_�&pT�z�Z�DX���#B� �����D����A-'���i�:�5%8�0�#�]ÛW���9�2�N��ɩI��cFzb&MD��=Z��l�}pҚ���D/,�}�4���6�륊�K���K��UX���sH�M�m��DCL�`�k���.�3)��"WO��4�^��Z���'�+��9�6X��h{^؊�����\���m�m�[9T�s�J$[��q�����^���篲���u�F�yBYk-
 �ęީm��K�j�~�����p�Xͦ��d�=8:�����4Ֆ��Z1ݠ,-�Cq+iB8?-ez)ʩO�������\����gO����UE�r:^�k����&����-4���cn���"���3�:ڹ���T�m��8�����+ܩ|k�>�WGVv�t�Ǫ_� A�!����+����Ă�31���� ��+5d�|S?�C�LιfL�o-���[�'.G��nH�}p��ƹ"3�*J>��y��(J���	b��3.>�b6�/����ZF��.�(`��,R���J�C���P�bg����,�v���X��F�]��s.�ј�/��L��M߻s#����9�{2�?Co��Qa��a����k�*���;�CRl�	�@���ң��*����s"FH��+V��d��w��E�j�L����,J�)G�T���v	d�!l�i��_(�IL��V_Tm�Q�d;6�Ô;N3�,U!u���Ƣ����n$�<��$�����]���af��F�z%�r>\�����!��R���#�03�+kʳ&�s���[%��>	��V��;D8�S���Ņ�M�v?i���������	7'������
������p#�x��%?�|��A	ƘO�z9Z�gr�(p�,G��VSӦp����~U/|$�W��6}Y.�e�'���(��a������5w�܋b��G� �7��{V���+�ÆV��&L��t�Kx()<�X���m�H�[:��6��B��_��։�Rω*�n�]葼���i+�%���<#-��4�V�����c�,U��g&�(I��Ҿy�Z���9��1�Eⱎ<�����ѝ(�ýT�FO��TĴ�2��'0�,-��}�;�%�'z	��'��^�?��T��*�VRV��a�`j��M�l�Q��L�0�A���z����?��ܬ��߀�6����j��9�=�ԓ/�ӣ6Nr^iB�7���)CV��'!^��p�s@/�88mZ�S~�$���&⎑��׎��a�6Y���M$�y`��$�?���+�	Uy��-H�Sƀc�d���`Չ>},�K]��?�H����qdO������8i��x�oo�`�*��#y�˅hWzSˀ�~�/R����%ƢD^�2����,��!酣��-Z����t��a�4;��'��GfI��4۞{G�8�W��L�%z���Y�������a,(>�}���8�،�¬�A&����F�|q�:p�l[�2�N��M��[��JS�����3�&���pTy��>	S6^:��,�VS�L��.�D�.l�N1^��/�9p#qM�-��`��s�r���vw��!���cQ}�R�i|�� �!��8���=�>�L9E�V"&�~pܕ�O;����H��z�%8�7ô5k��Z���}�}�?$��o���>`~�\���߁�WI�W�^_��3�=����p�8��&mrG�3�L�m���&�;�?X�e}X������e9���,�.��f��4��M`?J��nx���8��i~��;/���$A ���hx���Z*w����В��J�R;�*4X �]}�jI!�G]r�`J}(���������m�uMB�g���HeN��pM���E��A��&_���� ��/�P�
k,:B�����d�C���=+��Μ�oW;!��.�&���h6s��0��'^_<���!�����u8�/ �������`V�`��e�ކe�� ���d�0��V�-yI^��}�R�P/$���;��MPa!�$�LHj���O`�Ê�#���J��W�8/,���������o\�6�j���'��Jw����3���M��U~P��;���La����'�g$�!���1�K@���`sl�]CM��N�FRʍȲ��aE�y"U�%$��TĚ�e�R搼�LJ���?h
X�"_A�ҝ��l��k�9	�g�u���X�v���^_�Wilj�9􇠿�� ��O�[��ݰ?�c���z�ٯ���]�['3e��
2�X;�P���A]+�����A��o\���������{�d4����-;M)��(� 7@q�K0Ki	DRvV�,��H�:���8-K�t��T��+
?�h(����L�ZM�N2k�=������>aί���h7���8FbMA��j�^�k��7V�TW�HQՑ�QQ=�cf���,�G���4B&q9�ĕ��8�Ӕ=�����m�+�mN$��D�>���������9�+���T�i ��۾#|���V��,Ӭ	`��>cL�J!W�S�ѣ����z�ś�8 �eOBn^SPwq^�=a�|��M���J�VR�:��yП�O��g��a'�ߨ)��;�t���J�����Rj&Rl!��M���"�������'��������f�A�|:����B~����r>�(YY���S��(�Pr�/�u#��Ĭi�{�"Q	A�F欘7g�
$���~~`]z0����f[T�)Ie��}��#3���;�"Vvk��y��Z�0̻��>��:�L��IW�b�/$�4K�I`�z~�b��Ɋ-�}f�O��˼J���4l��F�<�o�|�S�W2FS�4x`����4vc�|#.>�_�O"�\j��N�8~��?�*��3��d^��8x����W�x��� Q��˾�Bo�K�G���<dk��e5_���ѹ��� 0_�Dp�?�=���M�Us����� �����8�[���t��k�'��T~z�Y�!T���"�\o����O?��ѫ�	����9��S*W��;�|�L��'oQ��5Y��A$�v"�p\]5�]��	���0��s�kG ޼w��@`����Ļ�n��3 �~��(�q�%��8����q����96��E��@>��l��� n.I�O�Y�K � ��:s�m��U�q*Tq?{��1EZ����i�V @Ȝ����-�:�j���k��b� ���O�i��$�20�s����m�օ���_ ��Oj���(�y���fTErGT�颓���o@5,#K�{h �1���E��Į��*>�R�Q�M�Y�#cF1���F�`�yÆ�+y��Q�wԎ����D�H>�Ós�@�����,�K�����8KcV�=Z�nNla�Be, W�C��]-q�
��ūa�!7�ꅹ}�.��M�R�=X���; n���a����~�����-�"*v��cK��T��)�Q����j��~�I�P��'�AM7��+X���`jc��IX���>H༉�nj�"ަޡM�'�ʃ2�@|��ܐ<h7����c�o��.�/�r�d&L+��p{�v��u~h�.w�Iq�����9��W�G��ӈx:`T�u sġ���>p��,"�e:��J 5/
~/E��&��!���I�)����?'έ�[�0�"9�3�' �_~��@q�r_��HΆ��`����"g��-��a�/>;�	�-0~��V_�fE\�:��2�!]!��WLf���Gi����sd*d��}�R�+%�"�/�5_|X�W��}	s�Q�ڹ���'~7�bj�I��-���bP��ƕ\�4�#	o�x�|�r�l`:gЊM��D���b6�m�#���o0���-��p	[�z�~�AvN��5��w�n7+��01Z�H*���Uպ�b(3aE3^���&�n�R�%� m���D��0�A��`�r�8�+���z`or?�n�}4�����5�Fq4�9�7���,�ۍ�'_������u��p�㼁�;j&��4ѕU.1
�ϑ����e �؛[�%}�W�W�h~ߔTI���� �m���( 
�w-�Ȩ����ө'1�J�7�g�͠��Q9y�{�)R*�Q(��0�B�?s[y�u$s0���u��9s�>�ȯ���h������a)[lý��t���X��t.K�y����E�����Mk�ޜ���M�rm�愬��Kx{� 2�N�k����C�7ʘ襶�;��;
����Y�2l&��[�Is�wT�1���$*{E�F��yޝ�~�=60�?�^���(1��nǤ����Vwy��}K��e�? �ܗ�?�*�!��j�~�Ղ���:�����N0��C���ז�Tr�ݤ��-efa����+�:��mz�d�G}��}g�U�\���R�y����Cȓ�LK ��7Tb���Z��yӬM��<�
�
��C���������1X��r�MsIaSޚ;���
#YjB�mB��Oq��l��K�
_rY�<��+�P*vѫ6x�*� �a�;���xOD�>�T��҂Nnh}E�����S��؁E�B��B���p0�J�h��oO� AZ���C1W���^C�0L����E��������Y��@�Y��MA�ƛ�	�f�0�\o6Ǡq�+ ]���|�����$���"��
:�'�X���(�c�F=����D�]/��Z7�8TP6��p�K'�Pjx)������h��ʿ��~�=��P���.$�!���K����zW�i�?��#����su�τ	!��J��g���-��]6���� ��1�Y`���5=}��g��J������_v'��n�7I�"��c�>R�@O0�36X�����k�)�^i4�<�@�c�|��T._������ܘ,�g��[���?sc��D@�0�'ix�	�gT��{Y�>��ƁT*b��<4����J'Jw�%'�ۂ|����?�W�߮�sa�^E�N)�OI�i�Ĵ�jc�@���K��s(�l�����!9������+��в2m���j\c�*9���E�'�ל.��-@K(�G��V�9�Z�5ߏ2���;S2��^���r���]�?�L�)��nGa���8�������AQ� `#�º5�h��J����L��Y�8�p+mg�qy"�M�4և��g� ��2Ǡ�j9 >���P��o���;	� ��?��eD�;2w?�;P�]{]bޙ���~W˦�eEi��O��*�^~�m	�P ��`�lЧ΃��,��uj��G1Qr�D�	R��f�d�;�6Z	ͥ��."�;C��|n4�r�Nq�K�y9β�~I���	h����"��H*�
Y�E�-c�&Wj�F����� Y��`����R@ I��t�Rna�A�+x�K�D�V"x��{�0
0����f�v�z�	n�����9�!��=g.!j;S g��A�����l؆�@�=�,p]��IY���w":V��8i�/�U1I��ʅ��g;�i�� 7Yڃ˚'��|��ذhbG\��o��|� 1#d�S=a����E�V�\N�YZI1��t�_�)n�دA��УS�u�Y��<s��$=�P!%y�����r{�ӯ-����gpp{��XAHC6iS�Y�C�B1[�N6!��)�Z�ng����Z�#olo��a;Q��|�滏QY�pC��0�V��W�����+�G3��E�� !�4��1T#;����Ip�V������h��*$�����[�1�d�S@��vA���_yI�>�@��R���{�R���O%��*��~4YYA阅����6�ߗJ�Z�U��`ɴ������n\<�_q�e�R��}�@�'p����Ṋ�	���R����fF9�۰N���O�s^].���Gg��^�{�as
=2��EbT	\Oa��_�-,�]טc�W#��x2`ǅv�Sd��^��r�crM��)�iu��*L},5`l�r��DL2+�>֧�ٻL���͝,�B�+�8��6���=��	��a"�?�htĦ0�C�,[�d.�5�z��9��@N9��^ŧ�S��[�����'>i�����$PT�%@��Y���{t�2P��Է�X�z0��R�������?�b�N��+�N�ŷ����P17��VI_��('��VB����y"� D����g"�$T7Z��󷳓sVw����e���j���i`���/�p��v4���<�;�_���_�6�TJjd#(Z8���Q,-;�U$�x%�`K��&e���+��IBc7�����<%#~+���X���>�V��id��, 	����aO�S8��������MJ�}��_G�0�U����@�]�=_��[_+~u�)p`����qt~�#ԑ1�Ҧ�d�i�6���{��_���sE��|E�t�Ԩ�r�/3t��!�h��A�bS��w��5!/U��ԉީ-�ݎ���N�hza$I;W�\���|p@~�9���f�q�Y��A:i$���&�.߻w�x�2��x�&�����!|)��O�Sm{i!q�QΨ5��g&P찮��NJ�ĺ�qg.P"Q����uef_���q}z����Q�7�Xo����1�������L1��AF�u����J@�7�V���B17�b=��0t%	��8��l����!�����Fh#ܚcl��I(XOBˁ�}�u;ּ�D�M�k�%p��o��� ��P����e�_���xK�6F�k%���B ��.>�",�+��̷��PB\҈�L��s���⮄��&�a,�~��<�K瀆��x�լ�a���W��N<�ߕ��h�W&�	FKWj�)�j=�l0J{�	��P��K�s�^�lsO�y޸��R"��-`0����Ч'B^&0<\�����9����6���Un�Z���w���S������X�ݗ� Y?�d]{k-���7U�}�R�Uʪʧ�BE��=���p�q�X����7-���������V���*R:˰��r��_sN��'7�1?Ȭ�ڂ�AxJK���r�6��*�|���m�^<v�Z��Kr��D�j�%��J�ٽ�+��@�	���O�y>>EZH;fW H�WN�+��v��m�F�hOY�M��	b�q�E&;ƣ��0l��������f'�8`�"�.��i��a�x6�<��gֲ���]��M/�|0�ѼL�ϴQ���1������]���^��q̙�����3} �#⌷����F�J��� �;��?�ԑ�K���[�*�m����5[#I%B>-�ދ�!��e*� ������s��i�|�d�,ɁM���h�����}q"ޏ'�9�;��ew㲣�2�Fz��`���\�,��m��sl�,��x� �����	m��2�ЗY� �çR��1�ˬ��ٓ������wYO��<�>���Prh�iX>������(�}/}�&���V�K� �l������~Bs�b=
W��EA��Law��!Pl���l���^
�*⭁�_6���Kj�N5s �g*Y�I#���h>F��H��f�o�����@�r���{��Q��_�o;��_W�W��2��Ƌ<�ˤ^๠�Qy	��$�Qa�%Aʪ0i�CH��hBiL��>UԢ�� =�i�$�¹�'�]"�/ϭ���Io��@��W5�w�z�����;8`����Y�XK#'�6}$em�"%��k}�,u�ݰ���Z�n�W�p��nȚm9�_���pk�8�����Z�	=���x�k�V�����l�9d�+j���XQ~	�O��6�����Q����{d�)�
Tć5����⿾�7�͵(��zUD<�9�R���N��圂���ͫ�9��2��G���K�2 ��\��z<�^�7Q �W��x��M!l�쥢��j�I!Z����ňM�q1�=�'ZIf/�̰���X{�NG�,`��ʵ4�ʧc�R���g[�H�`oQ �?�{�?����Js�$W�!q�2�|������=ts/S��TLv���+��sR&���/����o�:.��J�5�r�;�<q�u����u����*�:8|V��ΊKF�k���E*2*�L#p��o����1��=_cQ<4�.g�R��Z�:�XQ������?�ʌ�U���w��?f�n� ����0�u����h�7���Q.̼ǗD��.���̠�sO+
�,xq<0�~����@t2�)�p�3�
�Z��xwC�i�@��qZ�C�+HG0x��m��ޑ�>�Lv���������ЕFX��L�� �M�&[<�z��}�M¼:���
M�ED��3/&�˥1����쾇 }�֏��cJ �.T��N�����r"�:��Z���A��T_*���'�`G(2��q� ��?��bG�<X�c��2��oZr���埙9Sx���i��2}�zn�H��~W��1;q�^!�)jB/g+u��}�QZ���lT���K�9���_+X�z~�(j�GH+��k�R�����!�;��H�]�b8�u�z��檵q6���"���]��6Y�ͨ���	e[���0���;����9@���S1�=O(T�+��K�;�HbV��_�[9�é��S0�T�BD;֛@
�������`�B��h2��i>�C;-8�����O�����(j6���v�/����8g�����x�Qv��n/2��=3� 6�Oڄ*�{�7�i��5��)V�����K��Rr8X!fĔ7<�<��#� ya b< g�{`ʨ.��|
�����T�eM�U��d2�����������k`r?���	:+��Z�$��(���~�)L.x����	� 5L�*��,-k/�X�fޭ;\���˒�+<��1zXwȾ�.���Y":q�c��&X�꿀�6}�����4�m%�eQd��\dsb]�j�3�vy6sPʽ,�!��<d2�)��\,�"�;=��N��-̽	� }Z��ލ|���R�H^#��$c�OJ�M)��}�&$��������~z��^�K�tRd�DR��$s*�æ��K	�'������_��X��j�K��ܘ7�O�*j���)��k ϚIzފ�F`�p�u{���ƋГ��Û��O�D%�֓S/r�L.�.�rx��&4�����擆u�Q$�Jv�]oSX�G�a�Ơu}[z�7�C��ib^Wi�_
'���Ӆm�FS���5�+ y\]�M�|3;DT�iS�_=�d=��z��	���d�\�=!K���{����7�������1|�-�2h
��5ȐnTc
c,$2���F��߸c���k�,�f]P�W�1s�X����v}�s��ƺ��OwM#6j�q�N�K�S]*�Ǌ�L���P��=Vmkwm�0��mhLo�7
Ɩ.�e�*�4�!�b��8�~��A��w=�#���օ�򝰟]�8r��M\go ���EW����pKf�ѩ�3`D�,=�4C%\Ky?.��_�_Y��o�@�=��P��3��n�Q�:�:+�5�����1�����������և��^�3E��k���'�y\��]�}��#R�C\�J�ԃ�Sj�DѨ5Y��Z9��r<SD_���x�n	��mjRu�OK��ϲh���؃W~^��u|б�pj�Cw�� �_���B~�Q:�n3
몖���
�����£3r��b�\#,uD����4��W^���s�PyJ�s(�ss��K��#z.���Հ��н]u�[Ң��P�u�y�ݭ�ل��6hJ�ĥ��WJ^�q6���?��Q[Q �F�@��������p�pb��qgDQzat�.��5W�?W���es���c,I8
�)Eoc5:N����M( �r"�D9���Aw��r ����z\b�I`��]�Ēqڻ�����Oݘ��&�4�$jM]>�B*plRݾKdb#	GG���8H�׽��_�eۘ�J����^����9i���z�/���H/n���VN4;P�ih�S��09F�K)�Gz�nq�\e
f*|���k[����K_[��|V��Ե7S��������o�	:���7��M��ڐ~�_v�9�V�ފaN*�w����`���h8n��A��.��"Ry�e�L�l�%k�y�\�Q�ﳛ�!��/k߫�z+���r��<A;��랥w�i妯t5o�6E5w�f	{MBU���J2,7�"1�G��b�|^u��ڰh�=p����V����m�h6{��II�7j p^��5R���	��,���s�m�$� �礹�T\��RJ�aiS����&���O�TȄ���k!��

,d,��6� ���	@�.�hꣵ��"�h�j2��zp�zA\,Ҋ��췔l�}WO���\<Q�1��%ynna�R�O���A������X�C�����Y��.���h�������]����d�8�^���!f��K�1a�)RA2��-����9�K6#�c�!�2q�"��d�����gSh�����B6w�)yzب?;���v9.؇j����� �H�-�%�IY�������ї��*�h��
�Z�n�I��͏��?ɺ��b�a~�y�W���Ğ�PCȖB�ZL��Jl����o�m��zM��4�q�!���kuB��E�}tek�?�$�� � �r=��F�؅�e��6�8�ԃ��v	+���y)Q!S)�4�uv��ߘ�))T��놃��E���f���,�&y�i�4g�Q
yC�$K��1��9�$�JxB�n�n�b?����g䱷�
R#�gQ#���S��{��ߗ�"?��������0�|ܩmۂ|��t]Ss������'p���zR���ɼ!�a���ر�&���ů�mOe�1��i����/��)�gۆ�R|>(���[��VR/Ak����Z��l�0��sn�l_�����v@G�&�)sT�0n��u�!�zE����z�.��M=|-d]�N�R��y�9��q���1_0��� �hz}h �R�RK���+���{W*�fsU��Gf��\��q	h K
+_A�f[��K�������ÀM���� +��|B�E�lNB�_���b���vB����%w��m�k�����2�33`��̠�}�|9�Z��u�f��׺V����E�a��gވ�7^iU�1]>��ͱ�f��?D%q��e�A��{<�F�6���z�Z9�-57q�/M�Ake��tW5,H�aXզ�լ�ɫ̏ڳ��Cb���R�j��b�ٸ �C�Jz*�4`���YF3��v�P�PR����!`�i�H�8��n�AN$/��������D�[����K�qc�\�
J`��<Z��v��_O��e��v��Yn	n�Yc�=�����c����!�x)��b!�$M&j, V�L,��x�R9s�-+,
=�����y\�����W���)�"��/`�<V�N�(���$!Ƥ�������H�e��zEwͅ�ۗ	�HVz��*oCDUQ[� 9]'hY�}7� kD����(|��E7n������E���`ফ6���5��%24ߕ�}&l��������?!~�v�m@0��$��ߩ�ߏ-�%����Q?�����s�̺��mL3�3�}�S���n�>R��n�RO�ωoC�xB��yO-6bf)�+8���1^d����f�dr��~Q4_^�����C������ͬ����U;�<Yf��Jg��`�L%�i� ��K�p��^�'�3!��-`%Y�W_L�i��w2s��ZX��/-����wˆ���oX�P8����P�H���\�v�]�
��wM���'��@{/�i!��lK�}1����\t,S(�����9�Z:��0�d��6Ŷj��\5R���MZ�S+5(LMb�]����"�C�}M;c��������;n	=��ui�zQ��[����\�Lj��~��������
��ئ���#�G�B�+^���y^�����<
?��7*�����/�y�
�B�6�+OШSG����/���K� �h6)1|�X~��S"a��Y���!7������������(�]��y3u���c �3
[���?������u��g�#��y<��V���}�G.R�]�=����|���2��������.i;J8K�����M�xQ�c6�����Mt�"
֮��-�RY����6�&�u�4ã��q[�O�(��G����/}BF��;��a�4��Ш�nl�
�?��+JU��v;mj�;@�w�Zvķw�W��
z;q�I��^p���E �/�oX�د����}���h���Ѭ�|�2ۀl�� �
BkQ���]��U5(�hS���YPSR6`k�R��K����f8�Z�,�����R&ߍPW�d�:�����1��x�M���E`7�G�FmyW�YY�v˙�*b>�|5ϐYYS�ؾ&@S/,$�ms�l�H�݃ԟ9�&����|����N�� Sv�s��z�Xe���2�|P��j|�uv�	õTQ��\ 
Foj'��1����s0岶�J�7>2�3�*	:�a9nf���"�#.ò�uեг�XG��[)$	�Bڸ=%�h�I��T+�W��z�iYۙ���x���i#�ʨ�6�x���cy���\����M��?/��٣s�_	~Y��M`���O%������n%�>�2׭���_�*t�(��5s�RԚ�ZټHW�Yn<�e����5�-���}�c]�W�F!^u�"�,�gJ+6�������w�n��u����n�ꯧ8�U�Vmz�4�>Uc�7ڑe�d5�K����¾T5�2M�>�&���%!���	��	闔�[�*ϸ�֕�w$�����6O����J�%�9z?-�Ʈ�Ty�:zé�`8�s�H,��w��>�s2�f<��@xm�f�xcy̖�a��;�EI[�Xe�� �ϕ�8;1�!��ǭC?x�:+���v��R��H�åטu�܆��/}�E�n���E�4�a�cv��8��:+J��,%��m� �%��I�2�s���yu���c�sX��N�mQn�ؗS�C�q�H�7-��u��.�>С������1�Wmv������t��+J]};����hl��ƻ�= ��+Px\�-Κ�|�jӓ�elw��|{�-��&�ە3�n6���~�(��@{H�3��I@��+5�,�m$r_¢ق��O��GgA���	�hl��s�	r�S�q:Ni�K�knJ��t��cjR)����QX��.�W���#�)ؖf��d���ɦ4F�؝�p6�(�W��x��AǮ$�"�&�W�փ�u���g���K����?�!Հ��:e]?��s�BZ�o���� /�c�|̼f.i�� XO�/�-Т�����'_U�)�q1�!߬��h��3tM�,zm涐%���M�Ib�:�08J����ֽ^3�!㏅�-��_?!�Oy��u}��:�N�����:)�M�9�BL�%Ǜ!ܻ%}��/��U�sR<T�l�C��0���S� ��	������XM�b$K�����!�XL��Fq벜l����E\�vL������Hd���n�oձ�g�h�1�ZFmm�� }*���A�G�٤V����E����#'���>�O@��/]�N�h����X$���|8����{�>W�J�x��fL�UZ"�!�mb���F�s�[.�H��~jHG8M������	2#�����svŗ�b�>e?��8��1,%	���g�r�M��l�OݤM�"�r�;��hK���ZU�+��~VoA�i���땭���d�>3��E2�c�����}~�]��{�#һ�Od�'���ۉ�$d�ϝyW'�����>�����5B���a��@�����(�]`ך葯4A"¶�$_^� ՠ��C2V��Z؎��\9��V��;f��,��;���"��?�b!0_���p������^�f�ѷv�B����-��T�ڮ/H 6�(:�)�����y�X�4�e�䅗�\�v���z�\Ж��=h�j��N�xM�&��u�x@*L��$��-�&x����?��ĵ�������;�k\d���{��4T��&AiR�2��4uǓ���ay�+P����Ė<J�<`�y���*6�q]�:e?���W*�0�]"�((W�o��?�H%���.�K"���������M,m��LA>�I3W�/	���@�l�}"�^�'�d8�N����
��9�'j�� ��(]�w�]�Y(��W�!�\�Ao	�؛�{䌉�';�	?�|�BԤE�WY����ò
��Y5�]p�ld�F�WW��&�����:���>דH���k�B� ~����(�p�����<�'�Ţ�w
8�RX��9v�Q{q��T��u�j�B��٣������V�����*i��,��E��Zr��p�;�-A���ԃ2��y.��2�[�5ac�Na�e�����n����)S6c��dor��4���:�	����6nU����U��-e�H'���XY�!K^��-��d����zS����ԗ�'2��� �g��lG���i��	L ����,�v�1��/9��='��(^��l�#[��InI���)rfd��N�?���D)'���X�K�
��!����X�l@d��]�!��G�$C�,�K�%ڍ�1��4$r�D��v�j"��g��(��O<g9(vh�H>��°�e�>�]��+��`)�}rx3�q">��Q��s��tj�,-��C�s�� �܍�V��H'��yc�0=<y��쪧){�G���ϐ��
4E>J�>Ě�Nv�i{!:b�1���K�-�%DZ$�7������*��uh�4�%F-��<^Y�ǎ�� �Z�^^T��,s^�}9�:�o9����?;z�J�;�z�/S���5e9����iR�Fq�x�hLD�m�����'��[��u>{�q����@�_LE#{��4.~�۔�-Yz�j���b)��/w��O�;�A&0v2�m���QS����?�	k0���u�0�$�Y;��T~����4^�8,� 1b�O;d�c�0�%d���^>�>BF~�P'�F�F V�19�?�U�`���1l�*|h��Dn�U�qtw�У�cw`Ӫ�R�!��rC�c�:!���+
�FD��x�{��B(��zVNwO�Qn���%S�� ���<�4��'I'\h/����gd�u�e��&P�,p�~1�%G�Y 𕈞����0a�˦W|)���?�[GW���ȷ��[���������	�cj�5�;�ʶed�Q�o m���3���Gj��~�M������6f�" l��-��
��.#���B��5���N�l�e!�����"M�Dq�O���w���]D��1SS���	����7U#9�P]$�ٳmjYXX�n�	L2ËI�?Й���J��)ov+�艜�>hI�"{��nE|��O|��-A�1^n ��0&�S��;r��n���p���)�o��1����"b �_��wK
�i%�!��O��q�0s�cO�'�R�Dv��ͪ��ū.�%�o������)�����㐑ѧ�$��N�� oiW}�XtG�9�ճ���h3f�1������G����jx�6F�hC$[w�����IY�C%�Ro��с�+��Z+6t�O��d��2������(8�
Q�P�{N�
�d���˶>�H|VRh��xUH��yQ��HV�/6�:*<�U~�U���z$V#�'s-ٞ��غ�Q�H��1�Xq�!=a	<�+�OO�T&��L�꒑xZ���o�âƧ�ǣ�ɿv�9��wz;/�᭄��!T��&�k�O�n�@D�}����7h���>��ũŃ���r�Fe�.�������OS�� ���n��J�K�8�2&��t@��q�[4E��@?ꉺ�$C���4��/�JE*c������k�1��l��?ҧ��T蔽����o�|l�z�<�5�L��:�*������3(}::�j�,a�R�]��)��Ooq�̱�������L�����ƕY�:S��t���)-rO�g����%�SU��}F���fј���I��vaG8{�`и��:�K��ق2])�]��P���8��x�{�G�شG��w�e���C��%�R�bM�Y��8J���i��z�O^}�i���Z7�w��M,�~^���v��8�����&dī�@Y�G3����)��57!,`yWۑ�t~�uZP��8ǂ�X� 	u�l:�k��MX����S��E��\��K��J�e��}�	��v8��(�;o�"4�������4��Ɇ	�Uh[6���L��]UzV���ֻ�ZU�y� k1gb��*�+��f�#������Z�I�
pg��P&e��-���j��1k#\�y3.�����)m�$�[����'6z����?F��>5QM�?�I��+Lo���L�|�(�9H농��2[R�x�CHf�Ow�̥t�I�<)(�G�B�;�N�%X��`���ݑx6�3Js�_����%�H*X���`�ap���G��!*��#�-O�dUt�t�x|ёi<�����c�"rJL�Y�Ogנ��
�j��-iz\B2���arc�Wj�S�"��0�̑ʹ.�!l|��� �KkX��88��J�����J��}&��
�����GqP9	b�'[~U;S?�u�>�3�l�B��|�悖c���"O��9��@-q�{�h��1���J�1s>�x�7w�N-��c�F����^<�3�p�B���a�BEm���Ͽ�=�8�a��ws(}��:�o��a��U;ifP ��	|Uԋ���J#�1JP�9��*��@B�Lf���b�B�Vm�@��lOH-��0HR�"�h�W�(���¼��e�l�4&��[�B�r�>]w�RP������ucÊ�*8�xE|�~6�vyOỈ44p�Lr517�pߒF��.���b�Ϲ.�6����.� �`HP7���'2�#�-��Z?z's����+&9�X�(�b(��d����.�Ó���v\�E/ί��/R�iAl�'��Ql߲9Hbw5��Q����**��<I}�T�((~R��Xa{��ҐpU�a�<��6�#�
y#�����ƙ�������Wӆ]�$��hK��c��{�BjQ�`��݄ �j��>d�g�[��ͣe�{��E��Ce��%���	HP�Eh�ŲLy��X"�`y�t4bԀ���R�gST���c���)��.��1���f�����)�����5<`Xā�%�"�����YJz`���o{�����.�!�@������ݽT������]U��I���i�Lƴ�6`[0e=2l����C��@Ӄ���d�V��E�ZLk7��U��UԸ��soFe×�e�˽���"c78hDXC�� C��`N�G�!���QVnA�+����H"�U�/�b�:��X�A�������c_����l�R�N	�#[���[=�\�[�C��0���$Z<��;�\	c*0}��j��7�\�m��L_���G�ӗʽ෥�T%����}���#D,��H��7:�+DP�.�ôn48���HV�����ޤ��"��q��L�Ź�tuL�W5X�����L���UުN����	s4���+��@[,�ͯ\q��j��\9V8qJ�9Q�c�������:�6C<�����E/�Um�=���4��:m�4szn`��l&����lg�1�M�)p�D�l?�2�K�},<�s���n��wE�!���4d ����L�D������a��o�7(�Ř��O�����`��{�kR~Y��isp��_#_<�hy��<���E��o73{O�(�y�e�Ni�e�!�nP3��V������v��3t�w�i�u�B��@�Jg��f;x5$Ȯ �%���#p�?�û�ҳ��Z��`�k��: �{��K.��$x� Kf�ݾ���xCR�N���nU��]���X��i&�χ�xc�Hp�,��c��5�-�+�`�M�5�`F����ȅ �Z��+𙤀#(��I):\����>󻝢�e9萁2�T���1�w^��¤���z� �Ϟ�H�K�6wv곮�ve��P�P+�_����pH(�ͮt��z��q<a6:��� �Z�#��u��-�!@����a
h3ȴ"�����S��Cf*ƪ�/�����g���Ծ�@�c����l4��5��|��I�1�L����][t��VI��n� ��=�
d.	��PR&�*D�����m`O�Jzb��1�ȫv��C�g%�)��<��}�U</�bG����M4�m����sI1�|Z��ijq�0�V`��0���y8��2�,wFy�$}����k2���XM/9JT&��W(�0:�
���f���8p��"�,�2-%^n���g1�`'N���}���I� ]\�Vך��q&x��t�^�~�%KGD�"8MQ�����u@p)�D��m~pY� ^�*L����(�L`cv�	�N������ғ�OP�Ka�Ӛh3��ȃ�|\�`�#��ј�.aIu��Y��&!p�d���!�F+�P.�`��J�Z9;����&W~���=��Yz��&����Ѡv��h.r��#��{@�Wz�K� �k(���!���l����՛|l�s���s.SΣ��VO}GF�d<Uő����7�1ת�VU@W΋�E�X~6���H譖1��8��֎���1�O���0)� ����͹P���d�k�5����W�Ю��7��Wo����(�&ma�p����_��'���A����*�z��M��F�r
Or�#��<0���,�e��$��`�&��e��~�=���͏ 2gԗ~�R�}ZQ��N�xK�*oh���3E�*���1�0�&b�$��8r%n~�
u���^t�&^-pz���t�f9N	.&�������a�H:�����J�=���5�	,ￖ�S��T����r+LYfuY*�����~/NጠPe��h��{ؾ�v__� ���v���O})�p��$��Ar��< r�<��H��w c�߭�,M;���L�W_hwB.�yQ�"�Apl�E�|�����7�7�e�-d��&٘�7��w��E%����c��������ε�A�6�^���$˶"�$���)��R��\ք�	�Vj}J����2_��Q$qí������h��0X'K��Dv��aU�6:��v�%��ŕů�/��U�|�����Z1J٢��F��g�!(m[vF5���`Ĝ[7��|��{z��kX����l��Nhui�	6���K�N�����G9$ ���.��⪨}ɇ���T�:b�ڔ���xal�.MAW��A�}rq��d�Wg�#�z__l����rD�rG��q��<�%��
����Qbެ�����Q�C|�����u-�H݄�kJs��u��P=_�o����  ��#������H�}�3��Lp>�����Mv���`7�q��jYn ���r���`�*��Y�}7�/³�g.-�`������ڝ������F��U��{�1���+Wھ,˘BھɈ�=�У����v('���d1f�Ng7	Ni�'	�IY�K�Rx�sut� о~�a�"s�!��~O�i���:�'�z*G�q���T������W��g'VZ����Q8f:��D�$�j��c[ewV[�S���`�>H9��d\���0})�$�[�#�/���'۴#[	��j�@�Wy5'@\V�2���Q�*q�-��?sOx&_�]��r���Ll��'�u�,8Z���-]FJkyBw��
�N@���0���~��	��Md+������&㯭��Z����f�x��{� 6e���ɽA��[���GW[�"�j��Ě:���\���s(��a�#�ٿ<&̯5�	J�M��'�g�(k����z��r�����$���2�x.}���v�B�.$bu���gN8Å��2�5�*�4�$e�$e�N�Ơ!N��P����}e�&'�:����%Ħ�L�Mn�rjk>/7�4On��݂*�#ү
���<4���O�?�[�*����"�� ��f�B	��fy�v�W0ۣgV�Au��uٝ�|D[�����d��tB��8�L$�&�`��g{6}��unz��w��\c���ɑ���;F�@��K�ۊ���d�,[Jm���,57<Ʒ2��l��XVx�����2��E��3h���m��wȔ�L�0��R:s����2jk�&ԉ���6\�
�6�d��L��}�G{Z7�yɡ�T��w�5��}ZɃ��`��)/�^γ��W���%ƨ����<\:��w��Q�Q�G�o���7���x\�Pg���(g�*����!�$N
2墹����9��Õ%�s����o�Ʊ��B�f�����\������zQ�P*}A�JV��h��ۺE�aCǶʷ,����n*�w��f|�oz�E��.���PK���H���A�	�B|�Wt����� �z.E�;����mƆ?N+ߙ��u{Z�-d�W5��U��w�S�E~:N���٧�z����I�,�2�Z(b�'�ɉu��0glcg���P�����щm��D���i�T�^�
wZ���7�&��?h��ﰉ$��xSC�N�O��[)���_1�[���Hp6��(Vk�xjO��Sݛ�
67rd�'���h���O,BO�\}0��_|i+f	Du���ؙ4⋘��5�N2~]��9iH�2J�>p2yL��'Þ���:�X�D-)�T�(K7@"Ŧc	1PS����암�Ipk"o�1M��w6�\)2��)l����;�iP;����!��{���A�gh|� )�����'����M�t?F����\��$W�/>�A]Y��[(�`���`"�Q�����I�w�GJ5����U�q��gC�p��C�m�c_&$�n:�s$���"��k-�,D��TQPf6u��}V���i�sx�H�ꃼ��VE'��n������â��,�KE}SQa��9�ؔ[{6�0���Z+R����Λ�����j�a3��1F��K�-����e.Ɩ�Z(� ����Q��ckDb��$r�T3MA7?(�,?�%�d���Z���,��(�آ�yS����3�µn�i,9�	Jb�4I�S�Is<��8�ݗ ��)�*�d ����M#S�D=�Krד_� �)㯹����3�R��^կ��wK�T��4���p��3��O_����������?+Wђ�!��j�Y)kLTVݴʵ�ar��� ��TM�j��q��#{��K�^��4� X�Q�<b���R���V�z{�h*��ci��ĥV��hCr���S�L"}^�>q�ٲ�k��&U��8�|I�%c!�9�l��$[�F�@����H��}�����D�)�p1By���=A�?��L)`k�:I!�Fj@]�
���[��<���n��y�_C˒$+�@Ҭ�0ٶr��Ol}i�O0J���j�v?g��ֽo���1Ì>g T-
a�t���͟!������\�g�a$�BJ�I���,�#��Z�u&�O�aK{:�[w X%?�-$�(�yɨ����e�9�o���$�A̕ ����͘�����J�!Ұoy����鿻���M���~u}�B�E ��k&$
����V4)k��0�|��@��u��cG9LM@����k�}�#��;յҴ�$�7��̕Jp��y��OM�^�LA���$D:K�_KA�1;Ɯ�;�!��w5%U��x�z���|?��|V��a�_�xN���,_+1��On0�TF��D���Z��
<L�BA�E����+����Z��9 N�!ñ��Tx[%� i���
Ęp�]q�RI"�}/�M��hz�{����9~��:J��%')D7q�
�D)����du�[t��i���*a���'X@+X�H�����1IЊç�1C��������ڑXx܇�� ˷�I*\�w�״D��~Y�(7άl��=�L������$�N�a����T/�fk��6��uƒ��2�i"�"����d�z.l��>���� �@�O� 23���y<H %M�丹y���T|B�)��)#_|j��s�o�5t$̣%a���S���a��.�d�n�J4
+(��J������[����o���[������9�Ʉ�!"wIb���g��R���m-�	�VȻ���ퟙ�H�Č��2!����$xv�|�f���y[�H4&���$<����)�.��e]��[����Z�v��|���"�=�]}�[L�j�Y���/�v�v�~�L�ω��5̈́��x�qv����q��v'�<_\�/4s!1/aX��3a����غ�{4)n��ܵp�λ�\'��{�f��*�6�Ȱ\d^�g�]�ۻ��=��#��<d��$$2���lD2�C�M��"�Z�1�r;��_��������̨#e�؁ǎ��,����16]ɏ��~HS3ݲ��ū�7ZGx�>��T&g[�>*������B�.8$[H���e'*Z��bE�����\��ou�v�K}�yT�[���d�3,�Yt�����k$�4��P}W�?��j7L���ê��+g��|��D2�5NvQ�p��!��;��^rŶ���-e����G��:���?-����	���^[�o����l�H>��T���U�w� h�!��$�y���)�ٙ-v�o:5���ɞ&҆��pa�[�:P�+����a�l1�"����{�K�4mK1�5%>9u\���Gm������[b�aI���~뎼~�u���?ކC��ʞ�g[���O|���	k=�P�dYA�%�k����&J�����Y�S��� шd�`�=vg]�=Tg�SO�w��	�E���¡��a����	#�
	�n�+�P-�QU��3	a�)���+�q.-Di��m�U����*��y���c04��?5�ĳ��0���#�v�38΁�g9ٝ$s#����~8ܚ�a6vS�i`������a�F6o�������^�h=�)��]񲏈J(��kY��{�Ն��Q�29gH�?����>��9�*����m���p�'�it%�8� �On�1ߗ��om띊��@��I/b͢t	�c ��اd��=8=!�G/�MbXC�F=Ɛ���#�x'�7�)���{L�����z�������)cLHXC�kQ���'�N�h�ѻv�rrbi�炸���g���B�?S��%ҿ��
-ٯ.0�5�^zQ@�P\j�"ES����t��}S�{)�|��W~"��B=>~yU#��9HsE6f���v����"�v��Q�����MV�h�հ4�Q����
��a�ުgX�ZD�ۥ�g�t��'֏�.��e�CU�'0�'h�, �<G�JK��!ǰRۛ�H�OB���g�����$�+)#���-��ڏf��>��S��wUt|�]���n���o�����!�7��`��!��� ,]}�8��>�����9_�"U!e	,�EƝ-�$�kw���2w����J���$�G9�Mp9͓(�ó��-�}jqx��1q~���ė�<�Rʩ±��gy|
�'mR�g'^��5�,'4���2��w�Ȉs���ŀI�\��e���L��}|��:t׶��=�VSf����ӎ>���<���X�B�&��l.��쭃�N���>�3�߷v>�f�@:A�Fae�]��r^|�4�/�u��;5B`dėK�y9�I%������ ��_"3=>�c~�g�z���§��P����K�S�G�F+��F5�`��JۦI4X�C��Ջ�����8"SS#s�	�mO��:�5��dQ>���d6����X��>5]�f�k���5+j�)^$�o�رȂ&�.&� �Kp�d��yB����|�:���Ț�!
�r�G?�P8Yh �e������8"}pWZ�LL���p��>ȸ�e��4�	:z�$q�u�w X�)	�Ͱ�QGF]�����TK��j-*T�@�h�Ñs�(����t4��j���Y�v۫N�N��1f#r/�8u���|t����E��N[LW�0|mz߽���P�>�v$y�ٴ{�]�o¦.`aNM��X��r��锠֬I%��Е�����]Н �$r�`b�V�~xubJ {��O�.^7(�O�X�A�&.RC�=����f�v�a;!-�$+��~]����z�SD�0#��s�X�W������I�]�?��R�nwH�1���&��j�g�(�D�w�|����y��t1��@�:�m�Qx:��H�g�EL��)�a��6u�y����:-&	�5�.R��ݡA�w4R��u6ir�G4�҉`i1Hp�aĹφIͧ��+�$KH��T+�t/�3��BQ����b��:�zck����7�����u<�,���9��ݵ�A�ϊ��KL�A(~�F�|��Z��A�d�k�Jw�&V%�E�f�YX�%���Y�~'jFw�~��7�r�Є���V� N.��]��"X���o���b?!�]���E6KjP��PU'�����t�w��I�0H��pf�j�HՁ�RnF�p�TD�Y>���w���bw�Q�Bc�@A��`Z�s���O�����t��3v&Nv�����S�R^J�}\�i������VDn���V|Ի���O�)��S�%�T�C�g��;+��_g�O	�ˆ`�a�<짽�cm���P�F�����]03�ǫ&P�_n��"9D�u�����ɣ#Q����G� LO 9_�]���C%��Z�Zü|*�Tg2p�5��S���Uq�N�䞲�`o��xh mų�D�He&�uR�#g�kh�x;u�s�%8��Ǜ`�42���ep�k��z��HsA���qX#��5<��'j�,p��yHH#�v.�n�����i�x���^iX�b%�q�#�[&����D�s)�s�i�밍�%j}9��}#k}�`=b;�:b�{8����)��e�i.g�P�<X���9�+`���N~�]���l9�1M?PW7���&�X�--�B�������@ѽ��i+^�}a�'�{������.S��Cf�m.�Қ�)E��^������[%��������Q!�o��%�����ΙTC1�����T�Z_��u���ص���(��sM��9��m�g��e��^ә��,Ē,�gaQ3����Ю���I�!� `����r�-0��z�mr�QxwJ�M�\c~�(���vLL�����4��%���8������{ջ�Fu�8�{����78A�a�&��M��J,G�ߎ^O�0�E;�PPxw�����g���ӄE+�Ֆ��2���y0�ة����`&���uQ��Ƙ�u.��)�9мW�A/p+2��:M�^��FU/l*��,BTf8����l�Y\�0��	U�+ ����~<�(%��(8�k���d:�3>i����ǘY�0�>]'';��H�ڑ�jTbw���-�N<���Ȗ�>>�h`�[��ʌn������|ͦ���L��Tt�Cz68�hLp����Q�Ac�k`40LZ�vEj��	�El��s��L7Rn�y;��]��aÜ��˦E�t�S
%��m�g"}�
�#�Y@Kw��-�kw�zm(�-KL�Y�p
�������x��9���ﰉ��ܦ�	�K�뎅_&|_��4-�VZ�؁K�,l�Vĭ�s�Nz$3�cآ�;,�9e���zC�V��!5���F��!�����n��To  ��u%%(���7�H�e�0+�^>���Q�Tv�S�������S���/����e�t�;�]=O���nM���"��F�J�5�ˊ�){���C_Ѣ�+1\��^{�/�ؔ<އ/�^/5��7��`^�x�ؐ�^Y.���	����Q��#�-��#�n�Y��Q�W�`�71��m k.T+�Aߙg^�O����ˇ��h4���.,�F2h@n���k��H/Se"�	���B����}�G+$�V��m���z������m!������_�P	hď��J�K��� �(o 
�s��Mk`��GX��+��������K�F8y#�[y��[E�%��3�Ĝ%k��*�я`U�6��7XY]54����N�A��1�<r��C8�7z�{x�vӖ��l���2dyl5+~����w�����������$��E����_1�<K1aV�e(�§�̭�h*-ʴ&����ܤJ;դ�z~KXܖ���2l�X-��,6���� �a�@S���Jv�˃68& �{9T������)��^��B8V�.��\��Ԣ⧰*�r_��^�w��[�@W��bC]_�cؔ�V��Z��d\4�p.��5m���axH�:0\���+���<�a	x����b�G����_�q�*������uv&�oHo�w_�9��`�5]�m��^�נȊ?}}:��,����m��x��^s{�����I:�E���wz����c{}$D���iұ��F�\��a�R�e�K�K�B*�[ea@�bj���oJz��VoGU��w��64�H�,����N7�ޙ�����к=u�mt+}�R9�T�!�f��񿳻iQlje;"SYUR�X�I[��6#m]����1)Ѓ5^yy�jb����p��-��ρ���w�}̲���B�UP�a�*oBע��oe���Qn�9%GI�<� �W@��z�ۚ�_��e��=�NǱ���E����:���ǵ肕��]��?nc_�hw����2��ۡC�� PIz�F�;��A�ҹ��v69�M�5�|QA��V{k�%s��6>�7[h�rAu�h�c'�T[�̴�XR�;U�
���R
���V����zZ��(J�nx�y�f2��6�W���)��Y���K�"ʊ�.���g���h��X$'O�<$ޒX�b_}�� ��K�9��&������J�I��R�(F��|-�g��y�z�4�i�sk�|@]�3U�g�J|��eO�	oUZ�1�������P����+�'�/���j�V�(R��՛��̋����>(�6�#M�~t�"��_EK�}��Q�"9���e�G�ƙ���n�=)��!��^X��;rfҗ���
{��*d�~����S!��� sX����q�z�o��Y'z�Km�Lܣv�; /F�� j+A�f��#E�߉^�ϗ�R��6�u�7�W<3�'����*V��y�h��V0����~�Hz����څ��N�y#�"�DB�B~'��m���P;�/�w�A���
��FfP��t8��L*sX�E��O����G�z��z���N�?�߬�ô?����C�C�d�(�E\��.5AFX�?>��8�;r/�اpH�I|�i��o��+<��h��=��Ip���L�~��B�������؄��.�O�Ewʥ&�zY�!�6TH��D����϶�HN�*�{fIF`ΉLD{&4��`��̻��!�5�6Lr����(�K�/y]�z���":��ix~~.S�|�v��ӌ�iQ��	"�'dA2���A�H0�F�����h[�Zi�+ɊO9=�g���K{jÖ+?L���'��x�7��]�a��C܌��Z�0eޗ)�j+A {5��á[���?�"*���e�T^�0bPb�tA���
�u-��\�R�nԊ=S/���<����ԙ���� ��D#Q��J�q>�l�n��ŨH���J���R����U���K���:���<��}����!yB�Q�]%��^{��U�tLR�$�$MP|̪����2T���ˤ����[exzۻ�P� ��%�!a-�e�������寖�����,y�w[��0�\�M���� �ȿ��G�����F!��	:�}l�V&���2�&��E����fE�S�r�Y_}r����g��UB�A�]��#�_vE��)Y�1޼�'�A/�z��}��Z5�rT�Y	]�x��N��3�����������P�˟8�ldygQ�8�[^��8�^����t~[�]cz�����Dҝ4Ў����D5m}��\��-�섉�6n�*��v�s�}�_G����g �1���b't�06��q�-X�A����f�����3�Ij��)z�c`�f[�ޮq���xM�@
X%��.�tݥ���-���F+LG艙��a��Pr�Ś�-{�3R\ZZA;~H�4Ο��IU��H'[��&v�����29�����	BN�TѢ�
�'����/���+�=6��+.G�J��U�G `���ae���p�9
��7=�?��� ��ۍ��u��I��U��v(�h���v!ڑ��c$e@!aa�������T��@i<@}٪O�o�@��yӫ�������]��|(�Av:̩��TѪZSڭ�hB��M*���y���k�T�V;б>zo�bxK�iK.,�P\,�<�);2)T|y�SJƂ�T�z^
b�6��A������,�]�y8�'kW���8m'�m�K���'�m���S��#�-�Cb�=�зy��u~����]!�V&.{� ��t7�?JO��q�9p�:T�����	U�u׽{+�e�eΪ��O�O�:���E�4�x$n>���|�e�R����6y��m֤j2�$Y��N���S�A���vv�`���/���Z����䦕�2}�
��<�<��[h�5'��ZҾ���B����y���YK�n?:)��"Ro� ��c�����\T�Äv�-�|r�<{�x�R����\�h���`�MƗ#�C8��#Tk�K�@��Xi��߈�m4�(cf�¨x�X��K]�p�ൡ�.)}h��wT3�l,ӕ>~=AgF$�x����[F�H0,�!(ݦ~)r�AF/���;��:� ހ�p�T��`�l�B�Bț���į���c3y��܇Tc�!�9�!���[1<X

�x��D�܌-`Xj@r��dQ�Z=2^*kQ:<{ٞ<��n�\��l�e]b�5�fR��p�P��w�J_�W�J��T֊�$�����1����K	.���2B+
��c�,���%*0�x}f|w�����k�Sai�1�B/�&+>���aSpHc�2Q56Č�kξ��&S��_�2u9��s�W�<C�۝�^�6K�&tP����/_��i:�v���kH�AT虫6�f�by>j�E�u�'�m���>��b��H���S�ch������	�&Ӛ���I���E��X��y�wf~������$����G�g��E ����r���	�mn��ݻj�q�20,m�t�[Ҵp���czT�݆�3��M6_}��� m2��TYd�R �b2L��0��ɇ��^-tF7:�!�0��h�o%����-�(�0�x��`-aV��:aH���[�Q����l����16և���ڡ4+��#뫱���`{N��ʺۥR���V��V��H`d������϶caQ�;��K�a�O��hC�Θl��/t0� ǔ��QHH��7�m��Ù��V�O"�O>go�hQ��' j�	f�wɻ����,(��*<��.P oϋLrB��$]���Nuu�����l7��mMtz���sR[<J��E,�?ߥ)��H��pN֋�������\�I)�S�e��u�i5�j�e�z��K��#��)�[��i�N
Ct�>�1u����ևi�<|*WȂr�lM���4��*��LHӕ����7����=n�ˮS�hj$������!��Ѵ �Oq�|���bLd��h+E5[�~�ll�#�s�8��?�w�R.���M��+.%B���E��Ԍ�G���#=�ύ�QkL9��)k	���Oo}+�Rj�;�$�aCq����u�����9O�V-7kV�J��F�|-W�.1>m<�����ԋ� ����Mh����v�n�27�3���%�ZIn@V�%�S蛷�����火C{fS�c�559�X#���z��iW�A64zq8�Q릥
I\�9�m)L��>�(/�f��i����	~Kh�dx� '-'�%XIt5�;�5���Q�yf�����j�Xmλ���?�]�$.(2���cE�魠��
�RM�:��}N�l�d�Ąb��W� ����'(���fv^���3��̜σk����y���f�ʇ�p3߷Y�I�x�T��\�QN#�qn7��2d���+�5~x�q��)�6<�o.�Q�C4����*���� >a�7'u	���R�"v�O:��"|�XR�m���F�6(�ηR�,�)�l��&�-����i��K�;8���!\N26?�*/����T��9[TPdBa~1��3��d�����E���Ͱl�(�<F�.P���Z��ԧKB��_�2�9,�S�~ۼwl��gG�y:m��cm��hk;�>�\��b>�T��:v��Hҵ`�A�����
M�i%{�>����P�2v0^�'�er� L��	*�q���T]"0p�t�t�um�R�K��l=��(�q)�O�9*�/F�Yf�b��A�$��B�#�*�6��������d%�����͹Smn�|D*���w� !�<7��-�8�k݂���Ʌ�31�2Ԉ<a9��	�L��J�wx[�[�5�������Lb0�R�i�U엓t��1�)�a�ǒ�}Z�Υ�M� �΅��AWEi/��G�k+�B<���s ��f��vWY��±���75'��գ�.+�JJ�u��uO�OT���u$����I���K�S�o~x�'��d�'7g��e��M��:?�6���~�Z�_��a�C#dj�x��>c�,C�R�+���lY��m��.��M�e9]�E����Cϰ;GB*D�|G�U�aSⱧ"Q?��m�����Ǖd
�J.�:�V CQSO��"�j�lJ��t�Pڷ	��-��o�Q+1h+b�[ֻ�2��\T��e�3���UL!+���P�TX1�&�w��u�
���Z��3�R��u]� �W�m���e�����fSnC߶�>�ܝ�]8��uoh	8U�f�����;Բz�_+��j��]�)jL�s<�C�8T��"�8V��4����R����7�����x�C��Ɵ|/�j��.��e�Ǽ_��ة3�Xkk��	�K�c
�"����ŦY�!�$z�y �{t֊���(x�m�54���KOD8��r>��W˯J�%���#s��vU�o����^�gc��p�N0L���:�:�Y�����WX���0�G���5����Z#$�����5ڡ0�\�
$��2��
r�~���S���"T ?-8	�Կ${A�9]�]���4���.�l4AE�p�>}�k`��[�B���sY��"dqܩcTl�}D��}?#����G��E��j��Ű������iC'E���=gIFڿ�:w
BǤ��Z�mĥ~ۂu�P]C<��`�y� 4p
����=���^�g���c�=7���5��[���s�Y�uG�W:�ڰ��U� Vd㌛��%�l�;�+%�8��������u���\N��bl�=��6V<$�>�c)����}a�a��ݝS�"mi	�X �s-�l��d�ϝ�|�M���c�w-kg�
?x��~E�9�u����4�2`R4����v]�t{\1ےt#J�'ި����NSV������G@c}����rV��88��kB��TlK�� �*vl��n������&�N  }k��U9\�=a�Cر{$��� L�+}��I�z��Do�B��n�f ���s��,���yO�pt|Lhy����rMθ7��@�nS�"y�y0��#?#�h�8�ANlT��g;k� \B���VN�81����}�>���'�k=�߬Y�w1�~\��\������j�r�Z�l���_�07�$�5}��y�������q�%����Xn;@���*���*î}�e�w;�g�U�N����7�4�5N���5��2�q��lR�u�Č�8" �1!�uA�#ۢ�F�?Ppa��V@/�&�j�?1dx�$�X�ZU�ʛ$t3j�f!弼&��\��p�U��.\H9js�Sw���.�WX�$)�|�̓�#�J)��R�Q�>�m`���d�������,˭�W*�ɢ�`Յ4 ����3�D,�b��kِ�|������gje[����[,F�r̆�T��ƉLf��'vVq%^���[���>p�e)p���⬩��PG�t�,���(�B�k�'�I��n^Woi0�ʀ�D�%z#�n�<N���� I�K�xR\���ԣ�A,J�y��T�'���s���FfR���ϣ_%QX�3���%p45�. �ޮ)pP���mݝ:j�nh3Y0�.vq#v���^!0e���8���PЗ^�/64����Ǣ�	�[V3�r���K�c��P/Mv�:oc��	�&�$�Q~��En9��t�+)�Ҟ牥�>G�U�ՉY�����N��^���v����c�a�B��9�� o$�� �J9��=�f�mqMvT�ub�K�[ڣ�`�����1�-W_{/`na��x��چU$�w�vdL���;/�iUĺ�
v����<�w
�3��ރ�3���n�ܨ�=�N�� ���X-�w�:�s2p[��o��)o�"�T��+���a@��yQ̹�SZ�T^�qvy��?��4����C<��+*�8�f�������`��ՙu��<�%��7�ƎLㆩσ��"]Hp6Y�㳿_������V�U�m7��Q�6�QCPN�f�)��r�S����Q������r|a�aC(�ݢy�+�$�@�R�
���>$�E(Hn�<儨塗u`�٩-q���/��ŵq=T��޹LJ�4X�nX�#!���[�a~(����"hH�D�/��/iU��u�`���gӲX�7��y�upB��$�I��?����y��Y������.(Vm�K_<�Jױ?����s�7W��;��_[lz�&K������oqP�h�q$���<<��UI��J���w>s7�0e+�8숦�<��0�`����V����pB&5�j^����ҧ����.,2����\<h?�g�n��ܞ���V��ļ�h�4����ZF��X������-�a�lv� *�&UA7�w��st�n�m�����8�i�x:vs��S�ԫ{e�����Ŝ���G�r�h�0O���爄�/*М�i,��P�F�|vKVZ�!�xK.Q���JVB�%bGyy��X���k:���H��s��FN�l�z���;Fa[:�8x�*��9h�7=��QΞ�� 'AAR׊¡���?C
g���Ra�	�aPR�Ǌ�j|����$�ꊊGPQ��[ŒOseY�r��4�ׄ�ڙh��
>׬J��jr�4��xf�")��j��t��n2�aTu�h�i� B��O�Q��_?O��a�1�	��@>'�M��A
�-8��i&���d:v}��$�^�n��d�S;LI��@2pa}�z�ӏ���7���v��*���1�G��Y@V�b�!GT�Ss��cQ��^�B}�OP�2�]���牱�7�� �;p^Tej����ठ:[��UO�uvPQ�pK(o�#�s�(�6�2��rl�`v����1PF����=I��?���C��aB �_f`�4/���;.L~^ţ�af�+���\����lp��C5l<<B7����K�\ϹY�K�<��.f
3k�+�ϵu�wwa�+�4n�+�b�{���*���F�h�����]�ǟ/C�W�?�gQ���Y����M�T���2�b��3�����D�Ϩߠ�
���T��I�Rt��e2���9�F���1����ճ���0� ܪ,N%�oL�����\�c���
nT��!���֖g���O�3J?��Yd�TG�o��������o�r�[=r��^��ALJwb��.��e�_���˚�x�L��ߙ�?m�!Ӛ�%E��a�����Uy8��ͣ�jy�����/�'6�4��n��9i�,�*B���<Xa�{�$^���� ���Q��I	�~�p]c ư����Ѩ@�,L?(9l�����`_k chX���+�~�6�S�CP9�ׅh�SQQ�׫�<��l���7���*4��E���I��#U��#��*������Ƹ��Y��7/����?ojM����q}�/�;���L��[Q�&�%A�m�9�x���0P���ɬ,(�GN` ,�;i�Io�0�-9#���S�t�����Ӹ��q�al(\��6�ؤSC���z9l_��AŌ�ɜ���X֑a�6?���Ǝ�@���O����v�UW�u� �{� ���H�B��N�/�C����&J �i�}�k�ds2T���<��`�Y/N�ԗ�������<h[9�Ȇo�#�7kJ���"���Z�����Z�8݅mIw�@)w=2�J�$M�#%p$u���X������3�[��j	���^���b�$W�x)�,�3��b#p�x�@��B%rPZ�ϼI�yr�j��#���t	��|�ʩ�ϯޗn�����?��,���U��>�H����P�ʥZ��!�n�aFi����
��D�׌{ځ����E5Nɂ �Z�4�7���L6�8Vǹә0��)m�ϵ��[�z{ٷ;X��x*Hg�0�|�#f�a�gmQH,O��S��E�F�P�� >���*��z�c�!ÐY�,F"�A�769�m�
��Ed�"��*��6�6`��$�"�* �^AL,����I%�� v��z���ԯ�~�/�CC�&�F_gI���{�E\7�HV%��p�A�\�8}WY@ @�&;�il�⣉�Z��:��*b�Z@���q�����-=y6i�wJ���_�ڼ�;k
eA�T126�g=2�7ϯj�z/U��sF6�Z�i�$�M@ ��P2YD�3sk�<N3�Q�]/�}D6��܋,�w~p��i��a��}��.*�Ɉ�@!����}wf�pU��g��@�[��/��B4G�j@(؄ǋ&v��h��Qk ���3*<'5�"�`�!f��:�����X��b~�FgU�;�\�5 �#,gk�>)��,k,�H����Єc�����d\A�� f30%GJL�I����y)W����v��MJL��p����%�S�Q�m��I�p�_���S�N ������{L,��S;����V���t�m��9]>	�br{�e�;�AŒ��_�j=G��f�IUˬa5Yw\����X��z~���,�!���t����	{�1H�(B��B~2��4�!}������=~G���J���/��g6�*߲gWzi}xF���0�2��5C/���M���v���3��nR����'8륮����(e�o�(��ϴ"ݯ�Qͺ��"��=�E�R�n�������s>�i	�L����I����:{F�˛B@�{�y7s!��j�h!ۢ���#e"��f�
\H�(�'t�Ѿ�j�9�纊5����ɖm�쩘����0�
��4��)����V`�y����m���CD��}���]��g�)���R�E|N���w��������,�Y���=�`�F�����c��Rt�+7?2)��Ɣ�;��1|�l��j[�B�瓲��`LG�mC։���q��`F`.��4a!$�"#� �Ё�sʐ�S��]�!0ل��j�BMIr�m��'4�e �+ +ܝDX��n��҈-���u�\�S4{R�1�O�bj>��<m}��kU����\�%��HeI�d���UeR���ĕ�d}��"!�Ɠ+v��撣tDe����?��l�фA�����D�{LSƖ�+��3gW]p��Y~ӓf�V��~�[�1�n��3����9�)a��b3`�jy�L�#;BX�z`o}y�<Br>X�7.�T��`��$A����/%8�bp�a��}��=��r��1<`�wo��,*�cA+i�2�1M7�e��%�J�,C����C#�8`����F'��Z+=�C�x��'�u	(��\4�� �VZ,�~�
)�i3�jm>�Z������O�{�^U������:��������MZ�M�C#��~qM�m`�D���x��A�7�K�
�7v��W�$̿�>{�"ic�4�9uw����L�ү\	)��w>H)^�CZ/*o�z�R�{	`+��}�\���ʿ�K����?d�S_�������l���k����ڄ���\(�v��a�~��ؠ�o2�<���S�$�сT��8'�֜Ձ4��]E��8Է��H�@!���O2�:l�GѨ�˅a��d_{��\�����z���^�nWgR�]�ݩzG&��!�HB�ej'�+�j�_�= 	O�co����0������;e�&B�|��*������( {�_y~M�*�� �=���TS�Q���+qY�������������ݸ�yr�m[��+��@�ж7���UnJNE
l���❹�������U��/L�a����9c�gv< ���l���;�\��U�QM�!�A'���h�r�1�kf߮Ez��^��נy��/ �����Lf|;�MU!9�z�$	O�W���Q)��)T.)��'���W>���M"�"��7ZQ�ӜH�T����p��쯀-����8vzd����c	_���	:��?�&�7F�����h��v�r}1�O�g�-'A���1Y����e�5����)[s���J7ÿS��<]����;'�}0��0L�A/�i��Xr�@w�%!�lT��'%�i�@��-Bmp���W"�eS��QPbe��|&$�Gj.W���\�M���r織-�@�@!����߬��~��Ӏy�3���bR�#T�p�mMK0�w�۟9\}�����
V,x�O��lekvx'F�I}/��Xݻ/��+�gP_C��Y_��o��q��M��X2�!�5�ְe�ơ����� �,uP1h͇!�}����3�@Uo��I�
�T��9��b0l�1�d�;l0J��F�`fk'?��O���
o���Y����/����鞳���8������,�mmQF{�a2^���L�,ۦ`ܴp�,����O_F��2X9D=�x�1/�f�`l�5�|�"b����Q����m�y@��H�.�e�!sb��*�u�QZ�6(��8��fOG;<�@�>�q�F+���D7�HhMm��w�7[��V�@Δ���M�|թ�!dJ���3ҕ<w��N�y����Z�k�A�Z���S�'�%��x�O�U0pk`y;�Yt�H���� ����S��{g�@t���^�Io�;���u%�}�m8��伮�sb�ǒK�
b�B�?[u|F�R"珲b�	�Ӣ��_Yo�sr�I{"r{�q�-�2�pw�#�)ǹ(�l��kb�ߞ�<��4ҽ����  ��� 	u�x.���t�`C�����)�xy���\t:�fJ�*
�z�	&иߥ�f��Ip�$Έ���E�T�A�l1l�4��j%7��	7������J�bpy{���*U�qeַ�J�(���x��e��r�H����bu����:+���#(7�������U&Ḱ��?κX}��k���d�F՞v���m��_ʴ��dHx2b��M�^޾���9�A|��M�2�;}W-�N�׍����wbv�R�L �e�W�^b]�-�(��|�ؖ���,UK��8�IJh����
��#���ޚ��V\kl�N�9]Q�71, ���cv��G/�=�Li[��w)�,�)le����h�X��Ĭ�7j(L�����*r��m�
:d/��Г ���|�B#/9h]2���"[:�mld�m7?L���MY$��/��}
f��h��n��ϛ;�g�1�%����\&#3F~�"{v��$�行�C��rGlG�7�������0�̜�5�v������3	�d����������m��0�������[��������v�x^��l���}��[�l��Қj�W���i �I����ٚX���1	&_2��JF$A�<���.f��s�G��w2�^t��ZC�)n��edGtA��bB|�����(�̟i'��E����{�P����͍�E[�r�ݿs]��w2Ӣk�ii�<'@ ������P�М�'2�~~)�J�ѭ���b�a��?ƈ���"9�������b�7��P��*k���Ԩ�^��r1�3�K�H�A��Jf#f�h�����zϋ�:!���e \�&�5d�_�\�	�M�ߦ+�fN��H�Et�rt/b*ل����:T���d��cM; �Ԫ�z%
���H�iӅ��i�p�Fe3)3`=�����[Nz�/ຶ� yG~=rL�A�'u��4l�P��$Xk�����/<s��!��U�LJ�V���˒)��l���=�7i���C+�A"3�<�=�\�Eԣ%�@�a���x��rÀ�5x���|/IV�KoY'�(,5l�GOQ`�o�E��IԔ���8�P��"Zٓ����:�ǜ�'xh�����uABG���A����am �2>^,��:p�2�F�C�JDEШ���B7a�G��v"�=�W�4-!*6;(`����Աt0j�� �g�S�����@�� ���y��U�pi�;���[y�O\ҷ�����=?�w���������N��h��ux�[;,jt�m+����j�t.к&�e��M�o�l3��v��͸C��s�̓�U����I9{(�fI����^$U��9rx=�UAc���#��9�����v�zAl"�>5 �6j꽱!b"�}��fԧ�4�y�1�O�cT2d?Sn$������i�P5X�|��v�<FX���6B(�1��:�z��3���߆�cV��8W0�P���YI�'�R���I�uɿ՜�Y2�,�BT�0���\i�e��P	WC��d���çc����Ȇ| ^?o*��!��~���a.�Y{T�Ry�%=��ܷ��gX\JzO�G;#Y�p�C�Z���L�kS�F���ٮ3#	P~�^š���H����=q��h�Y���=��!��+	�⹛�ØA�D�ف".���h��eauĚ����Q�,�5 �|��t �3[O��5�2����:��k�&L"]��u7���d��y�EQ�IV��iC��Y���^TZ7gz����m4Z�������I�AW@���A�#HQ9���N��a�IX���ބY!蔍T��D�];��o�~���;�t2��؉x!�锗�,�8r>7�q@�|b�9!��$���8��z唪������^S�m�$D.IXa�S�"4�4�jR8	��DCԺ�9���
�p�}d�|����tA��Ѷ�~/�{H�L�m��iD��r�B�4��r�Y�\��"���Ti9��"Uo��5E����_���9�4Q��[��E@�I��kH�Q���FJ�(��-�U�A	
@�j�������͵���7�����g��g�	[D�^L7Ԃ�d-�ETxZ�����V��&&���@�ZI':����c�)&�с�)EĮ$�ܢ�������B43��o<�aǚ�3eA͓~6= �Y4�Εء�7��^<L��#�-�C�w�)�0,��Н�f1�h7
+,�#%ۡfЭ�MuDE�i���(��ml���Gp���$��G[Će��r evl���9b^����,:�1�0H�
f���eU��XU9x��T��B�ɰ�e�f��|e����'}��#f�����JN��6�͖䬵�Yt���Z�,�c����� ��Ǐ7�˝[
磳��c�䁑z0i��t���
5�2�?)Y��n+1%8�d<ƉD�����~qU
خ��	 �"V	�ͧP�7��J�D]i	��n]����!��]�`��`����A��g]��f+l'S���
������s���!�j`��4㪳�C�)"okeⲀ�v�!~�������ņv=`,Th���Mt���TN��t̄���&PK,N4�x+j(�)m����Ԃ0a��&�9h��
 e��q ������{�>�aܥ�̎����-�S�4�\k���VN�p����#��mX�>�����r���J�g7��s��$?5��!���2����0��dv_�
�D	=8���(8�I�AH;�[E�D����ۭf��2�����B��؏ �B�G���#*�Tz�%�x�O��N��TQ��R�d���Y\��$��ꂽ��ʅ�Y�R��n,�OB\�~�P�7�o�s�ة�Z�D�C�W��#�����6�z#��� a��VC^� 3jZ�09A^�Zt
z�m&A�zx�{ʙJ�'�8�s4�'���2At9�v�b��ih����������u�Oq�^Q�~#����2�9J�1J�� W��w�* ��o��K|���[W5(M��f� �H��[���{4�q=UQ._m��gd��%Jü<�Ϋ�����A�ym|��l�kQ�׵�ns�ja�e�\��x�MI�\��������Y��>n�ƒ��7hW�pA(̻�Գu/��zm��!�؟�J�5��G�DY��gj��V�	����*�=x#��k�s�]��BC��SO>ze���&��}.�V'��r�2����"TP�#0��fQ��ٱs�I����m^�p&A�RG�K��� ��mT�v���y�`�1�kFP�F�}�)�������5ļ�[�e�� �(Y���tw�;�.?'~���<9��0,�H9>�GȎ��~�
/υG�ř�\Ye_G�uA�����0HH,Q��2�¬cl�H|�!����:'��fI���lY�k��T����a[����n~TC�9E��E�4��5�H0Z]�vg���)�i=���q7�ei�vj(<;�2����1�ٰ;�p�d53�R�q��^x�FU�����y�[G8\{��E�6�&{fe배m�����Q�	̉&��0��t��\���u(��I�S��r�e��������ʝ�ߙ�����#�3�$����,�~&��3�H�W���f��a�>Q�9�6Lw���wt������3#�`J���.	��߅�#���A�W;���7K�WG�o>�
	�2�{s���^o'�������)'E����KYBn㳞5�US��!A�Y����.��l�y�aE����N�̟0O��1ZAJk�əi���<8����	|U��<kh�[f�W2Ph��V[E}�_Ⱦ o�"�Y���UP��n��.l� \u��$�n���m�CHR��JF^h;J�`���߇Q��厖V��>=ei�Gp鿴i��YҀ-I
��a�e��B��y�=K3�*�5����s�ޡۯ͒ox���i�`���
鱁����KI- �H��ZA9\��)(�� #��6��9��,n����5��Pg��õ�NXz9Xf񬐥�.x�]�ĈkpO�O��|'�����=>�%#j��}=���8����:�1_ˈ$.�'A󣔊s?��:�i28�B�J�$@���yA�z�B����U�o�D{�MT�q��e� ��*HI|�ß�(׉������i��Πe��4���^�D��K�����q�5� ܺ+_K��5K��c*��y�Z.m[ρ��v�K��ٗ���%HE��(�r4�϶%;��O.C�`��}ȫ2����v����DĪ�M�a=K������+����i�k���N�����_^	B���K�S3X[ʺT@�q緣���(_M>H���$N�8���+�0x�3��	IJ-�$�uh�Y]�� ]�$v2ޗ%�L��û%����bZ┈o�M�5�ߚ��a�7�k96Q�0��~4|(�*c�Dj�cI��X��^]�su�!b���)�������*.��=Iܘ���~��iki�%e.H��ւަ�;�H��ۘ�>D�hQGl�ǃ��JmV�MmOkIߏ���#��S��c��?�1�0í�Or��뜝���iZ�1�eH4�4���mz�	�'�ԋ�6��Fv6�WC(�-��'�̳��سq��q��=M�]b����G�K��:��ָ��r�w�B � ƈ�i��l?�r�ȹn�[O��s��)������>�S4���05������~�B.k(�
��SO�+��0��R�:�9�Xy^���J�o�������l�HݟĮj'=��K8���d���	��Q����s휿�j �ӅMj���T����Ό=7���{�ԋ��T��':kg�g�6��(9��	U�f��	c��x�l���0o;uw����u�$+��V�Ŋ�_���L X�Õ�ݖ�nn9>s�ñOD��.�;��As,�xD�)�]ZK�zՊʚ�j�Zg�Bqi�aE5�B�]��HGHs�j�#�|��?�2��>���1;�ǧ�� N������_Zi��2��N;6VKPQ3���:�"����*�y�9��>p�0��e޸��g�*�!q��@�N=z7�����	�\ݘ�b�,�:�T�.h�$0s�8 � �e�jU�	(�;_�s��X���{a�1�ڸH���y����/ �䜜�y[��Bc�t�B���0K4�%+�ן��D�2��.�?�j���#�y<�:�}7O��bL>��n�s��a��C����ibC}E��CM��f���a�@�]�)7���R�����a��+prӿ���F�oך�;O����p^urr):d�ެ1�Dr��ղ�!8}��{bjKŹ�C=5�ĳ@&;8�M3�~Ҕd�t�	HD�����̸�O5ۙ�lHc��5�L3�V�C	�(�
 ���?S���u�y;�[�$	��Kw��F=p��}�[)g{�� �U�Ы&N��J��c'��^�q�q��%�����1�˖,5`=�?pSw/�cÑ�3Ӗx��;,��ô[���iůl�Z*��W�n9���K�z�A���aL��[��K���ܞ�y���c����r��A���{��+��ؐ���8#�8�������==�k"
�)w!�`$���vb
1��w�Я���g�W�*/`+5�Z-ţ�_jb10� ��_�YQxm���d��"�y�fVñӷ�7�(�DQ{������P��^�J��X����%��$H�����4��-���AJ[�G*��������S�<Vክ
��l�2�B:1���S���*�q6[��$�=�R56�K)��������:.҈�=�؏�{��?f��>��t�R-��(�]�;:�3[]��mx����ip9c{�2��k)��)��ѥ�QJ6K'�װ�N����}�� �#�v��nZ8"��@n2�w/v���YnN��<Zx�p��}�l����	��Wp7L}L���b��ΥY�Oe�	t�m���%�(K��������dO���[����

Z>^�ϸ��7�!	�}�KĘ� _��� � ����*/�o-���$�h0��ks�4*���#_2wDV�r\^CCØe��}I��ea�4���ox�%����5y�z��j��Zyᑒv/�^ �y�l��w�=#� N}o��#rr�o֬(ߒ�)������̝���%zǌ�'r��Lc����F�4B����.�F���见��R\C�'g��e\c�!	��ʊ�\��Un ��:Ҥ��s�v�,�� zb�c��1Wj��/��)W���R2A��R]Y*��vga��賐u��:�'�� �������)��f��|�*ܲ�$�w%�������F�9��u"���u������GL�:�Ho�E@"�Ky�8Й6¸��HUF��.?��_{�2T�i�5�S���(��2RH��_���-)��]Q��Ċ�:�J�j������:��LZ7T������ٶ��\�l�J���+Q����"���['���M�6�1�3�v!���H_r/G��/m��.��N*�pJf �sܛs,�=mF��\t:�z�6�>z�zW�j�q�(��2��Q/~�93���k�Q�#�3#{�J-����I����-���w�uֈ���̪��Q_\���*u�
r���' Po���M}��O����`��p�/rK �hש�5���"G|��b[�6��Z��C�A'Y'�C��u�,�i8��8+�i���ׁ_w�Ӭ9@�4�H����@�ʮ�	��t��{��bO���j��u��g�����s�h��E|�M36�b���t\�����.:��N�+�%)$� 4��f2��� {��$�3FF�T��m������k����?[GO"�fb���!!$dDۂh*�QI����h<�^��V�T�S_B�1��6�J^N?��%��F`Bm�5�8rm��Ȫ� ��L^��q/��e׋���}�x�}�WƓ�- �˰��^H�Ԕ�{[UIT͋�ν/M"���Y�94�J��@�0qE~��L��A�O�C�O]a7�!� 
p�%��ƚ�6.74�!!�H�;���̊@�Zy�"�&�aq-ܵa�(ʛ���������__::��j}h�A_�$���"��z�s�؀C�?���40����zV%�tP^����o�b64�-!�N��oU��Z��/Q+J�DaJ����#X�d�Q&N�o>���\h�5���ǘ��#Y��	�7��=L�+�E��{���^�-V��ѼSx�|��A}u�#��N�j:��8^+�f��iP�5Z��𿃊����w���f�8���]s�,�,>�a�{��E8��ִr�E�Ъ��T��}e�8���8�A7a��t4�C�W��>t� �{���!�h���y�YZ�h�h5�菜@�T���b���>^@�2o����Hn��XCq�
p$.$D)�x$��\�kv�n��&��K���D���pLʥX}&��T�JQbh��j�#����Czws�e3R�&�J����Y5}n��N��0�
MG��c����:"�ZC��R�Z�wKBw^˕�[a\d�z`�5]9��JLs�+�J��0��>������#��"I� X`wŧ��Џ��(�@��X\�N��n��^f4F2�7��j諈��8�ҟ���'[�:�|��Ӌ�Y�8�:�U(V؄�O�Qƒ�f��h�.TRhY\�"�KX�6b��NT����q��Z��`������O@|�f�L�|D��Lz�"��.8=R:{q��;׺�%4vF�^�0��w��Q�̵>�'_b*'�wS�ѱ�k��!�m{��7�/�:7¬4`k6��c S��w��	0���\���;`���Kd;�r��+�]��?��������zA�[mU�(*6�'ݛ�ę!l�C�/�/?��V�vF��-? 1��e��L�f����9���e��gˬ�԰�Y�H�C}�ˆ���B���_��!�	L�N|�5!T�?�E�rs}����v�̓�� ����n�{n\��NԆ���)(���F����_ ��R���5=��Yp���xb,�vm��ˆi�� ��j�+c|�#~���NdQ
��%���G:�1%c� �c}����ͤP�.ho��˟yK0�lGZXUY�#՞QJ!e��X$Ҡ�s��y}�
)�Ĩ6E�0U�񙳁{�z���}�R��ٲ=��}�W����L���lh���A�f�p����߇EFW�P��d�ٝi�|�s��ַ�d*l*����vn�r���u�8:r�#ꞣ��P���v/{=��pz��Qj,n����������d�y�mgS�A¹�Γ-��]�c���<�܇�O|4���D��:��#���c\���a���m�1��>z�RV�9"�#��D+���K��h�8�@�@tv��M���b��cL(ش��VVI�/���FԢ����Ѭs��3�<&�m��	f+���i��t�m�6�N6 �@,�����@�8{��9��8�3����ɪ��V���(�H����k��u6Wc����b)�S�X#��J���чQv$���3	�v[o�qN�U��0��Z�+,��9\�Ȟ�niQĂjiJv��&�r�D����8Ӌ��z����X,ID�Xp]Os�Q�G�LAJ #�!j�@#�0���S�N$��1>.C��G����ٶ��e���N�[���k�ͯ��X0��/���.�h4@�K��dN/:a,���/R��"�E���;��n�T����_�λ`1���S�1+͈�P���z���/j���B�E�вuFzhV/�vOXpT�������Nv�3�-�Χ���;�J;��k���P˫
oY�K�4���E���m �Qu� l��Q�oS|SH�d���}*��g:����0���8H�a������0q�/g�@a*�g���W����9S���T�$'.����O3o�.�Ր��~�B˪1d��r�z����$6��o>H�5qKZ� c�8r����&�*��f���#�+ ~xt@��c��b�\RK�	���4mi�3���~�.�Lׄ*�ao492�{qy0�M��O+uL���Rm�<��z̽�n�������Br�,��3ס_-�WP����Ͱ�.��+�$��zf�ͪˮ��wW�Q�m ���x�O^/ԂX���'D��r��T�oi@��hS�#�ߚun���?q�W��pY �/�&���ST�0�!�!g�^^ \���8��3\�8}^S��'�����@<��ޟ�!H�L����:B�f��~��������h�<Vb������ÍY1(!
4#Ϡ�KR�,�I)x��'�Ġ��f?��իdxYׅk,�s���U?�܏�ʺ�zah$����E��˔���xs#�@ A���Ub��(��3zk����U2<�}\;J:�~�>".m��+x_et�lP ��Z��'Pm�=��c�;�60���e�G�>I����RY���TB��6��0�j��"n��o�;B�Axމ�0��H�rbE�L�?�{X�D�a෾����r��)׷I_���g_kM�)��/f,�aʴ٩2t�~2\H�C�R�*[u��q�Y�h�F�����/8s�p�o��]s����ڿ��l��C��J��c��W�*�R�2�
w"�5�s-��ì۵��^	����o��Mp̜�9��g���):��Z��!:����⍯WK{�f�d����D�zфN���W����
B������6�J� �}&���Ԕ{Q���|C	 =����(Q�4���a�.
hKKӄ�|ZM���d2��� ���j�����۟�Bs-�f��mm�x�,R��
�=�2Y�{9�"���R��2�u�xj�k"�ʻ�r0"T��o�J�A�u�nQ)�DF(�fN�!o���P{�i�iI8U�s3�=D|�Q,�	�j:~�q�V�t����
W��)�vSfP0(WW��L����7�|F`%a`�П�w�~5��Xq��'���n�r�P�p&*����߁C��N��;J��5�R��w���4tV'~�hk��f���f3��X6^�������Cw�a����[;�I<��0���O��������4�7�yka��;�#؛�c0�"���D�� K;�,-w�C?Ԇ���,�yX���l$F�E�]����(�i�.'1gFt|�أ�0�g�,���b�l@2j�`���خ�ߪ��� �ogU>�$v�Q-a���DmGw���B3+2�c�]����5�0+�o����wn���/��_�P��g��)�!HTW噵89!��/d�虳�d�o:�f����'��J����ݭUL,l�*�	E>N���E��E�Z�v��6(�S���9��Q��s?.�P���F�C��&�n<	z�ͼ�BM��ic瓺�.-��9��ƑI����W��G���h���A�]!�g��h��s��t��+�T�Z ������@�{���cO�y� t���bq�h���(��-�|���
K��U��a����m1�Ѻ�D��	���.�l�4�7_/�^XbV����"}���K0*�:�m嫿��R�b�o���0n��8ϑ��;*#��ԣ��q5�nׄ�?ҥ"�v���/��V�OA�C�s��b�݊�T$s�d�	� &2x駅XE�N� ,�,ȃX�nLЪZ@�b���ڷ_p�N�iy�'��Z��j���W��{Ȫ �O�Y�Yo2g��ZE?HN&���M��� y6�����ہnڪF4��U��;J(�֍t���r�c)�)zڨ�w�0	���n��ZDo[�up,��"���^�^g�ja(,MՋV\z@"����Fw�p!u��@���f�ґ�Y�����XI�z����OѠm��Vo����tZ�����?(��+.�\��q��J�F�����+x��tYr����{ʉ4�s����?�`�10�"M�?�7Z���\E�Q���^��"$N/$L�������&h�!d#o��#�I���1e�6�����q�(���o"��&���I�$��N�1�|d�ekϾf��w�� �5�!h�����pj��<a=���ɱ/V��A�u0��]:!֞��Z_k��AMN��ΰmcr�9hk;aR��p[-a��]ibM-�;4�K�3~Y@�4^��Y2>�DQ��5G�p����!�[�D�XE��/�}t�uɩn�� ���w�����r�����n��raN��0�G��_d>G��N	M�p����F�T���}��7ė�Mt�w�xg�;a�J�����+���|X��h���Z����[hb�£�)M��W�9co�9̲��|��zhgyK'�!w�N��i!7bn�ZY@1Fs�u�/ڻ��l�G%q�{��D0#��t������2-��z���b�f�D,jY��a�̫~m�����FA{=5�u4�aP@Ɋ0E��)�e�̀�	9Ԕ���]K�<Sɱ
�_�<K�Q�x>�H7S�Bݡ.X���0�c;���� !�|��ײ�7:Nh�O������Q_���N�d�!(�6_��ruPX�\b��K��Iv��pv&��$tB�PQ~��^S1}ϳV��c�3睱�V�?��ۅ��0�
��@M�H'2hb��v%<��i��5���5��!�<�����tί������)n�3ɸ��WV������
���?Ey���]��yW�u�.b�;�Xx6�!,L�%{�넏p)m�� �?��u	NR��&��QZ8�F�y,)ϳ���#���竝�\�4�)���p�U0������i?6��E�W��~��[TOm��`���
h�G}"��)���������Ќv݇�.���
�ܩ���\Ȑ�O,���0��=ܳ1�5J���u1ԓF#g̽|�2l��ploˢY�]�T��1�L��[��}��{a�dyKC�T�̪�O�$�Υ�lWB&b5��e<R5��?S�)��#JW��th��w���#�n�%��M�Da	Ĵ�l�r~�0�Ǣ��w߿���\
PQ���u��ا"��
�>��G��r���#���[�	SK:(�|ٛw�?沺�Õ�>~����q�z�ЕD1������V���Xq�8���s�ʮX[���B?`�!{Ӻ9Q4ZY��w;
�3L����"��mBPl���p�E7�wJ�=m��-k����mH��8z�!�o��J�jJ��X�؋Z�z�Mz��u�|1z
��6�	i������r����9�%�����p��E�-�5�޸�6�U����pxe�����S�.rx{ϕ�nw �ǜz�xQ�Q��$l� ��;P3e6n�*��qЫ�L��6]])������!x_�υ�s��r]ލ���N2�q߯$��jkV�$����������c<� cp��x��=��f�K���%X�?�bf��`�ޤ
�N�A�Y���0�4�+��4�c$�J��':C*Ǉ�Q|Z�*���c������qT)+u*�#F@�$�b�Y4�����&�lM��5�1�x��Pz�����E৾�������k��ed[dPw9_ ��(-[`aviʴā7LCT0S�q�O	{5H�4@`Z�؉�3��=ؓ�H*j���P�@���>vE]��)k�t5<,Ɔǲ�o6����X .���Gѹ�:%z�����Hn����{��A�����~�;ˊ��5�rxa"�A1�_��g_�G��xDTT�ʽ��'3�e8��B6'^�h]���l�#���݆ 2�s�iS�^C+��:��G�S�~S�In�db$}�%ˬ��풽
BO!K�~�XW�Տ��"�6�&s��#��b�~[>��=��Rt��wή��覆M�z j� ���Ŝ�q<�2�Wy֘�J/�z�o��($K������6�I����EZ��%M�)�"�X�.��lLE�I�ι�T��p7'�{j��I-�#�$ �o��NT���P�9�º���2�N��q�_).����Qбͷh�� ���,��C��6��87��v���,���у��s���Vc\�d��2�N��D�������XH�����̅��lڡ��lR�2Q� �D��߇r��Veqe�r�!����l!f���3��+�ҋ��u�t'_��d�$�H�V�v����euӜvkF�,��ۊ�O/	H,x��@&�O,u�:H��w�-
E��"
kŉ�CF��Y�X��{�4w����SM��p	�lGw����1����r��R��{Q)zan��;2�B��Ɋg�	So�[bk���v1z@�g�˩�ޑ�@|`����V0��M1vK�Rq��<i����`~I�iX����"`�.5��ʑ�ώ(�M�H8\u�F���'L�³�K�E)s dB[2�L�A���f:)�RqUA�?���ʥV~.Q��c4Q�B ��<C�m�Zi��C����AP��&�E����9�%�sJ�=�x�3����n��U֏&��lIn��?�������_�Xh��Cp�[�C�0	R�#��Z�	�����?"��U� �Z��<F)����AC��&%���Ǩ8a,;�s��0�7����F�˞0Db�wu�l���5���n^�!]P�U��a�%��9��2����M�_��Ïz5گL��5�����v�oh4ڧb���%ej�5S!�}8gl�4��b���4,�U��\���~U'��n/R�ﻧ�|3�ZO��=ԟ��2GU'NF�[Qr"i�KNn�EU�9��i�x��|S����Z��GRC�V���"́�H�+|�O�"#_,��h��m��,��9A��'���C��Z��K.B�+E�v��}�x���cR�tU��ϫ��خM^���kdm�� ��&ߒ)L��R��+�3-ð��ht�K���@�qa���G=y}8��ѧɍg9�M8�fq���6�6L�:�`ub�|G�6Z�f�s� �����BM�)L<�7.h�����-�%9eE5�iר}�y��X(b��~]<�f�-�(�В��ߝ�w�8�#��ECx�H:g�XPi���m�[�2�.����X��弇��!�P��uҹ]��y�`�ￒyV-\����V�iS�-�=�P35L��5$H;�Z�q��M��Ӊc��>�u��N���h_� s%9!x~u|o-�z����~�s5��X��&�\��'����"��
9�.cW��2�q
�B^��KK�����F�T� �'ɳO�s�8��c�	J��]�A
�hR�=��<_��(SY��=��?طHJT�5
�Y�HAtJV��AWM���wy��?'�,�v+��q�
�w���)3�����X�y�p0�N�*ׂ��zj+�.P��X��a�G��W��Da�������bX����]M���Qv��A��lM,2��EZ%� ˨�H���g_�VLZ��)�6iBoR�g&���	��m
�8���q�#zMHP�T��Z��?醃D��QC�rGEы�`N���L��ĝ��=p1�n&�s��b�7|:���#o�'((ӛ�Ɵ��ohw㴼O�r.�Y����h�5ɴ�J$��� ���򂃡�.���k��UfT�`c�VX0	1��
���FwuW��ů<r9�����&i��XG���P��R�i����3���?%���m��1gF/1�Ɓ厪����]3^�6��dX�@�L0�+��ΚKԷ���[P����ܚ�"e��
!&�7]4I@t�W��^Ca�r��n���f��>s�����pX�\'Y������!�|l[����T٭�dPD�>D�$,X8<����nթ:�s���,'k*w7�+Tb�m���+B�&�"�<���;{��z���g;���]j� >s$��_��A�\$���Q��1��#��{K'�Qq�#�5�~=����+��T���P7v�����o�Hp=V-�� �@�IѝzQ�8�s:�=��$"���O��i�jU1(�4�\��n}��5��m�^Bw�߯6'���:ޗB�Ke�{��'�N�4B63\KU��g5{is��c�O����c ,�V0��A�P¿[�o��c�^J� ��MD|�9}&k�c�0�М(Rl_�����I�'x,�w8��@�3��7�x�}�������! �:�5�w-]U�W��z�`�{<4�>�z����J�-)ȄO 2�d1F���*r�%��D�L�Q��Iȸa�BW��	�o��ݼ�N���S�ޥV�]9	���C�
���u��r<���'�f �P����D��T9�� �#�	)y�8���>9�G�+ob��@Edu�O�ӛ�U_w�b�O�B|�c�Qԍ!�D�<5ǖ�ϟ�u+uG�A�j����k������e�_5���o������2��Q(�̾'Ȋ�{J�Y׋��0�g<l=,j-�}���� #�*R�	�"�؏U��Jn�? �	��P���S����UϘo�z�6�,�XƑ���d�ߝ��ٯ<˨}�%%�����\O0K��F����.�i#�M�x�"�b�[|7[�1^���N�(� cu��&�$�~zA?����`�O&lY�Z�Z��\�Άoy�bx��IS^Q�qw��~Fn��	r�&���l���PC�G&�M�����CW�o���{��N��-��<ϟ�(
RcŻ�X),a�@�������"AX�"�/�6���;�OK��#�~�f�E|�bW���E�1���<��0��@q���M?���� ن�Qi"T`��UI`(�i�A�e�TN��Qs�`T��zF����|���G���`[Q�����8#p=4I��7����Y~�$X�eU'h� ܕ�����zr4�(;��ga]B�Q�C,Ɇ�k���)XM
J���&��X;eXX~�SƗe+>rZ��%��dC�t�����F��+N�O�*������U��;,�6��k�%�r8�TWn�,��}��'��B���M��v�7~���.��R�k0Ժ��$�y�x�>5�#G!��"�f�����ĉ���6�yH+(�Qnrغ�w���.
��k.׮Lc�
8?�9�Ũ��6��$���p�4NHF���Ŝ����2u���!f)���xf����.6�����
���-Q�w ٫������+�ias�h5H��쥅a�H�L$�\m����j�L/�����^�
��_���Ps�dd\bK{����[��D��$x�ֳ�����)�����s����ˎ���T��&�{!����Ư��,����H��	J�����p>����Zy���W�{�a�b^�|m�BRQ:?�4Z|ge��UڦRc���>n��y��<��P�0�!�5[�lz������0��k�9��hU�`����`�{e�H����3<�,�X�z��)#5DU$6kwUC��C�u�x���I��A3>w~��_�kD�(�5؆`��4��Kv76 .��]�%����*Tir�&dLi��(��)���y���2��§���	UX����D���� �G��B$�NM!L�ήHY\����Vj��S�$��~ O�@��pBv@�&>���s�v�>�8!�D���qXW�c��?�y6$[�q�l�q��ӹNY�6D۔�AL]y�6��ӻ3��[\�G�F���}��w-^�����!E'N[
��Rm�[.,Q���P�輰���R�Aɗ�4�=&6�����`����U+u�n�H� w.���Ml�g�������� R~�n�KL=���������V��S/��W��i���N��	��n����2�2��t�m'=�~�N�V�X!�?�>e;�l������L����o�!�˙����U��H��	h߷��_�f�_�9����^��̴������%i&�WLQ4�:C�({�'ϔD�}}N7ڼtF��Tc����E�2ݵ3*�`/y=�E�B�ѕ��6ٺ0���ZP]��t6�M<���OE0WT�%�� 	��%���8T]6�N��~_m*+�LZ}mO�v���l����_]�� b9�)50}wC[�Irl�xѰE��u��2	��:��z1[�@7�Q�Q�$��DdZz#���Ѣ[X4"��2|\�s�|�-�?��K�y��θ�Y�E������G�)� ]t���Æ��� N_�!���Ӽ�*E�5'.C�^��[�ki�jW%�nU�N3��;�g!h^g��.6ת��ߊnxȖ�]uLGE�%���g�P�P�pzݚÁ�m}�.�*�}�0Ҍ��� �w���x�졤�M"�s�Fb?;���E,j�&���q�ӌ���GEip���\���f*͵�� >��YE\����H���تsO��g,�����n�V��&�I��J�b�U�}��=���TG
�L��7p�sL/9w,ML�6��Nc�U�_Ua���y�� 8T �ԝ1!���ME�sj�&km���pM���R�g_:���LF��?���Ց�}V���k�j��8�7��|7�����tͮ�c�4�D{����1��v��kl��: ��@Y�*F�V�{T/7�=��$x	ЂƓ��ŭ�\��������"�MG�?�r�3�p-ɎS0��ܷ� ��MD�k��
���*��`�)#cZ����{w��T��A��A���e)@�K�J��.&�Ҋ�)yhJE}�)s��a���V���y�����Ktߥ�Cו��P�C�O���$��Kr�B��o�D����Q7:,�=ŷ�����U�D([�}�5c.���Y3�.��n�&��S��-�X�߸��$#kF�����;��Iؤ��.�����ì�rTa�miJC����Ƽ�F*��N��1�R�߭�	l�}۶ACo�0��dD�0h�YŻu��Ǟ!��8�^���t�%9�#0Pɫ�u�1Ǧ��$&|�s9?� gp�I�܊�*��A� ӏ��|��+�7�{�o��S71�[�Ͷ�~?��{��U����\a�Cm�W|��b?f�L�,��m7{�1�u�wA�aja��_��]�}r/v�RI����j�}2+,�]%���E��d4�]<#���1??���6����Y\7%H;�����s^�/
�Y���"�a�![��f/�/��@?G3/�����ⱥ�������ǜsWT��1m�2:ܮL�d\$j�P4�n�W��.�:�_8�A���h㣐��`�fKkA;��M[�'9�i����t��`�s�kń~&�,?��+��7[����X��<�6��	H)���<��	$3�U�Y�/VK�$��(�1��9��+��/��^Y�({��S?��<!L�`���|�� :���)+I����ӈ/N��y'WA2)�VuŖ���496�I͈�G�q����g�]�^�����d�n˯A�K���%�M � p�>��J�s!���{�}���l(R�.Fi�?i�o�>H,
rT����y~���N#x�N ��"K�wHq��s�K������j�t�h;�� �b���9����bDX:Y�T:b�qWu^"N��iA)ߔn����G�Ō��K����ɲ�C�-H4X���^��췋�����F��^kd����r����q���BVT��z�i�X�k�7���vntwEft;�S�J��K�$B2F��1���n~�V��s���]��XRE:��s��$]���l���a�\��Vķ$4��C�����NEɺ�3|�=8X�P��hQ��-:��˩ZJ����ƅ8~�ІI[Q������ai7�4��T���-��	U�ٱQ��,��Mt`��1̯Y�R����1�5r���t"���̡�[h
�-Jc�y���'$�+�P�N���th3[z���0��L�sO)L��{2=&yl�)��+�A��"Ub�b>�[���`U�쑚Q~+]`h����{{S0Z�XΏQU�Oy�M ��˨g��u��A�,8#��L�ӫ8?i���đ|��J���5e���S<��)c_aB-w�P�[��.���ܦ�f�u�qG�:�S�n�W�6���Nz#�� 
J�U ��*��ѴBP�*F�	���zh�pk�ý�ǘ<�����9��85��ݣ�ϱ�w�Le춢Ab��y�U�/�n��C�ޡ�I�����ZFT������/mF�|��e�j��6�W�=��_s;tF��ujz��lФ��"A@w��#� $m�ډ��+����3��?�S=F��\RO�v����Q	��{�n��Õ��Z�8���}}Frd��*�� Ex��+��M�ΑQ�"�oƹ�9I��V%��'�2Y��O�݉����L��6$�)6��a����*��I���;7sdA���D�������)kμǟ�L� Z8bhM�$��6��n���嵹	|�"����XѦ>�#`D2�����ˍ����W{U�?(�ý�$����� �w�}p=fP�A��Tm�1��A�]z����+� �-Vş�;-�-4���\[lx���舉���]��٣��;އ��������*ͯ0�MR�VͥӅU[��f�2���} �Q����M����8@�8�]���B:��DD�̑�|�u!�>����?����f�8���Hk�M#X�mS�������o~�a[7�"ޠyr�]*��Q�մ%v��)O �����H�>`������a�B%=ፆ6h(�ϋk�Ƣά���^mμ�黊�ne �ͅ�-S	�5+������IZ�o܀�.����p�%���:��_XQ�!\�q��a�.�5d]e��/�4�]���	��0�m'1'8�s�(��Gf�*j���X���c�l�Clx6�>+N��[fO)�HT`����'K��{��{�3D�%�N�Je� X����t�`BGG��9�@u�| �7s��*��Ӟ�q!ݥ�nd��v��%��g�����%JZ��"��6��h�fQ�݋��?�nFN�<e�Q�����&9ަ���Z�E���j,�8���� �t��K)��Z�u8��y���F!��V�dw�q���~���N?}Y9��5������%P^zT�V���6�s�4ߡE@u�����u�' �RT4��<�66��}w8�b�Hh`����{�E՚�rM�=&��jß��MC�mه�O��]�t!�v$���ev���	��=г�~@��tB�?V8���K
%��<���[�l��N�|M�I&��:����u3S�cV��2�tr �����dG��W��#��ry};J.j��?��H8������f/s�eŧ6�[s���r�h�py�q�6��q�n�#;��"�}׹w���k~�
���4�c@�$�ӥm�'��� �zC�l�����B�y`#~B�N�+���:�B�Y_yئ��,�%���YsI&�c�q���,j��=���mN�& �RV����+��p��3)V);�G��9Z�c��8oWg�����ĝ�ry������ޱ�/��hx*��˃��������0II+��Y`�2M�v���k���8c�4�k�lr�8�'���,��An��Ŏz^�e�.՝��@\d����cZ!,�f�ޙ3����g����r��ƏTBI��l���⪶�k(�a����b���7)L;�>9	��S}OjNX��@�t���(s�W�J�~�W�$y��ȳ��]MKq<�Uj����R�	N6|����V�#���݄A_7rD����oh���{%���G�@��̸M�s�	����:���d[����D�z�TǓ�[��>m�̀|�+�@�p���.� 8,~�2(a�oTi�������CE���)캀����1�;���e\;�vv{�ɀ+k$(����?�����(x�w��ϓ�3���@���,C
8��e��]�׶��� �[瑍S��	�v�BMK��AX�(N8�f/�5W��~�k�9�w�]�!����bQ�-����`Z�X1�w'�VY;��bu:^�R����;��eg�8�F��d#ͻ�Z����A��Ј�Ydk�@*��+��E����J��Ac2;F�l���Y����"l�9s9�������4E�^�A��,�i��}^`(2��B�Y6X͓��؊XA�}�u֝�R͛樉��=�� �`o����>=����K��h2z��s<�z��w��%�P"�RGj4�+ZR�@6��h�eȰ��I>1U��@��<�f:�U�`q���V ��6�D��b�8�`���Ȳ֘	~�h/\�K��y����!9�C�$�4�"�;9���Գs;��}F3�tx0�F,��v=�(�
�	������÷2rrd�K)�P}�i�DL�51��Y�@5�ۄJ{���<`���p~9�(�7Sv��ǎ���n���~i��n�c�1������o'��wy:��2{V8�j!�P��"`ec='�j:#�J���$Y�2�oT�"��cZ ��cr���%-ԩ��GCz/z^�++=�i��'�\>1�����d�5��I �G��� �1�1![��@�s��6�W���<����q�/O�L��u��XyA��m%�T�����!h/Maʍ�3�=u�{,��;g��o�!��Pg�ج`X<8��J_~/\G��E�a�%B���?TcR���d�Q�j>^��Hz��ϑ褓�OI�&��r4ꁙ{O�C������K:���i���(L$�m�ʛRy��=�U+�n��6��7�|ވx��`nY���L*E��=%�������ͥ����꾤Oݑ#%t��6��7�(��c.-;9�Qc]m%Th�s3B�{�N��7t���yZ��.�~�g�d���l>R�����j�}� �F�����э�eW��xL���ϫ��⻞bI^Ev[ ����c�C�ew���_'h.f��b�ȋ�&���I�J4n��������~�#���bfy���v������ȚG���PHp�|��������=(za�C�t	�1��و�G}��:�Ψ)G@0�*�ã4�sV�b]T/�9Q�s�e#{�Y��.?Ut�5p��w�?E�bE	��C��nk��s�k#��T���׮�)I�P;eH�*�z�|ny�6TN2p4��O�`X<����͔$���D�ּș�Dλ�j4��+��p��v���r��ڤ�%P��u�X�v�K�"�c2�M��E.9�(c���&�����~�\�~� ��zxI��yǋNw0dP�R����J�,�z�Y��(;��E
^� yu���q�ܑ&)�x�Ô`��Ǝ6���P��������_���{��)��l��0�3m�S]���]I.z�� Oɇ<̟�;A�x[���|�=��!$o,\�ؐRy3�q:3+�I���D����}9m}��p��Z�C���~?z݀cZ:6�q�()��u�;H�gZ;�@d�*!1�͘H�٨���%\��6vA�w����<�v>Xe]�v�c�ܼx��	$�~gQc.�!#�$0��N�F��2��zJ�|)b����¥Y�S ����P���6L9���p�V�3ۍ�7�#��^´>��84��76!W�WE���#Z3�~l2��pDc"���.i�����k����x2��&��yXGk�S��3�J{��oN!�t�iﲼe��r� ~���=̀�E�c�[Y�	�uj<�C*�����6S��T���q���.��kH���m��E�������h�S��_�klg�9[~�n{��Q�rʨV8f�Rg�Yi�R����J.�7�rz�v{����� �n/�]�zX#Q`�'j�\ۜZ����N����
�@EӅ�P;�kn������'��U ���Sd��C$as�3h�u���� @)![5�òl�t�=�tLD.� _q>Z��)<P��J���.KrT)�'�<M�w�U:%wAoL����xL�!f��z%-s���^��������l!�r����n2\��}y�X]+	�f�+�'�z�/�����h�D�<w�o@[��(@ �ўԸ~�"��0.S>��?*��?Ƃ�0'�V�IF�J�h5HE��
i�z��6�o,��?�e��h#�:W��Y��pKG+���$�l[�)�t$��u5�g�7"w5��ۥj�Q"�� ���珷:n0����
 ��ٌI_:�o�
� �b.DM�j�U���u�'ǖ9��|�,�Zt�(8�.[핓��T�2~���� )��ѩ��X��$҆��ci�B�C����>L��t��i�y�uŽ�W.�����3��f��V�V<Zo� y�$�m�l,�:AyG����3t��pѵ��JCU��j%|~��s2=��d�C^�����5�gi�YSv��%�3c�s=���k0R�)��g`d2�k!*t���N�d7��d�-��)� �J�O[�B��»`&�C������%f�5�/���4�<��������[9������ �n��ʅCUl�ig������SԦ�o��+�b�ĀL�6	vqmX���g@7����%�&Ys�6�����YaU��XL��L$��(*e!Z�ku)]f�>1��Cov���G�,����E�G�IԂ� �2�Zr��وK�>��ۖ�7c Q��pì+�h�~ү|��zIG
�\��tޣ��2�\x�@>��!&���ř/X��~�)�U2�8��#«�'�>�`�>s�8BKs"����M�xǔM��е`�ѫ�^��bOg����ɞ���ƾ*��Y��	�zn!�/��>֣?�;^Dc�c�A��5W��خ�����" b�dGd�5��x1�VaT�\�'`?�'h�m�Ss���E��d�qF���ɥb~��?2�6��1<�g������0o"�-J~Z�/�5��cq�������QsV$�V�����Cp)f6��R��^p� }���\�J��,��.�M�+w�ޚls:��&�bl�B�|!����{�����6z5��y�����#׶H�*��[zP)����oזW�R��b���uc�d��4@�]_�A� �u�5_DV~ݦ��%�1=gL/���zw(��'y7�q��(����G�k6�s�6������1`%)��`����y� /.��5��\ҋrkv=y�|Ь�5��Mc���Ej�g���zb� xG�fF��]�'��\$��>��]�����L[+�G5U��Mv����/��87tRթT���KQUx1���z�<���B�Ľ��#8�wh�C%^I7�u.1;҉����Q���� �-$3P�����[V��(S&�9GBc�ܝ�θ��w®W5�`�`���^(�ϡf��x�t�����x�]�k^�#N���?&��B����?5Ә�F��!|�O�u���Y)�����9Ƚ{#�]�L�����Hcn\�T�G�<.CsN���}��v��w8lkf
�0d�p����Z��?�3>�կ���li��qCs� ���l���P�Z����U��vz��)��h��ɴ���4�!e��;�#�.�QÇ��0}}��g��nN4�א0��'��YV����:�3����5����}︖h�t\�P�*%�jWl��1��l��	��.����c��`�~���QeKC����`���K���e�������!�ve�/Js��֞�h�k�r�fL��������z�ٵV!�jb(;3{F^�2����_i���QX�8��hr$!�66I�[���	�V�kINDܦ/{O�UZ�� R�X2�f�Vy�
���;w�6K�S¢ұ"��3��06P5˰�Hl�ga1�L�8^돵��Nz�~��a ��Xe�^D�dmO��L�D�@e�L(P�G%3�h�+@MU�ܿ����'
�T�AEC*��{q5��"�����z�M�Kz���jL��S�6N�U]�����i��n�P�x�O��*{�4�������S�EP@��\re��K��tp_v#N����;�%�k��wI��r���L���Bds��Q��D��iuk����Cq�{�\&�ڐ*s�^[���S��g�#����2'�o�l�x�B+�R�ǚ΍�	8�T��8�l�����ٜJ6���f8JnG�)�,�#���	�x	�%��}a���CJFgz��?Y����Q��m����e�W����倐{�b�>P?J��&=�r�Sb���B7w�󰻩�5�~8��l��;�]�pڅr��`5<n�Kz���%&<0��^*�����Ct�ܱ3B>�>��it���)@V�$FlN��?��g!��\���=
�Ua��K�Eje���ƗNz�&XL$>��$���:���$�l�׌UA$�<�y��g�9��oO2����b���/z�'�S��ҔTעbVV��30|�?)��G/�v��%�/�[V#<���9[�~g�ZM&�w�/΋�0�(�#8��D'���pkT�Φg6;ބ�$����������t��/�&�ǆĴ�ÇȚ.��Fɖ5�PV�l��#R�,���uZ�F�^�)�}T���]��C�{�?�[s��p=�%�����o�0r�ޞ�P�m��ѭ��E'J�u�}�'����V�F@�B��6{���
@=`��۳i=��-� �|��0�m��@�R�q�P:����X�_��"��.���e����s�p���"�JZ��HO���l���Z+�����1��D.�(1�-�t�*$��χ�f�m�H�<��Pc�i�-hR�I.ʅ���^�u������K�Z�a�� �O׸�y�k�
|��;�!c��.��X�"}/d-Wz��&��~�J]y�u.%}����(���?k���e���7����=�F-���| �OZ`��(h�ɿpQ���x�l�3�������<7!�<��@�;�ƁZ M g_�%���}2s"7��¦�.��H5' ����	�<˜e6�_W�6p�Y���CP�
���K��f6�|;�1e#	5B��܏�K!�z!�&��A�rN=ﴳ.0�dD�ִX�A���z�eZ$+��<nR�$�wF1�Ƿw��i}^� ��Y���wP�Í��Se�f������
[͆�BA�c�r1���F���>ʋ���@"Xp�^D2���T�J#��T�5�	�S�3�.�3˜	ᐁ���l��� |��|���ºǝ�}��W.vI�<h�{ތ�H��`�������G�9(rM�h���Z��R��M��B2ƈ���[�'��=Җ*����Ԛ�.���{jG@#
c�K�� X*D�+���*�z���F���l�6�O׆�r�7� |�,��X�����	�� ��T]p؜	��R��z�@�L�^�0�Ùܦ�����>>m�v�Ҕ�;�B�[�([�c��{�!�����r��U��/::W��B~����fyg\�<��={�Byj��I6$/���H{	Q�P�S��ĉs�e�i�[H�ELo3���K� K�Bή,#?��1���n��#��N+mwI�2P E�U	o&�9@��&�)��M+��VK��FF�t4CvP,��H��V��T Ա��!@rraC����؉�R��!��e��Mznr�Ӕ��u���+w����6�6Þ���6�6o�x��B5ow8�F-|P%��z�otj�W2�)=+E��h�p�ur)�k��rs7L�W]ޅh��a��������z�B>��$�Ⱥf�� ]3���ȟ���o3@���%�V&x��;g�Vs��6G[�m}�� �b����Id��>��I[Ҳ$_�����2r��T��P�X�4��@N�r�����m��Q�,v3h}�kH 3l��ݷ����( �h-���!�D�wq;��=D)4��$�۷SG��c�H�&*��i����/U���V��z0�D���#,eK�Ѱ^Z=i�r�����bo~�_7M���#(\JL=�|9�%�GAB���ʗ0h�z�R��
�{�ojY�8-��d���M�~̝c��#��x�E�#L�{���5� ��n��㡖)��U���k�v��@-rEΘ�DI�H�6���2У�HId+c�[ʐ�Γ#�(�*=9700��.��iG�����+R�� TMt>z��9�B�I���d�[�W���\�����iݰ���&�tѸ�Y�Gx� 	*1F�_XR�硕��9�pS��z�N�U�pf�V�AX�墣�0���>�dE*�2��m����ۘU/�)�0�~� K�waÓ}�	�o1=�m�����&���k��������,4���.����N���2��R+vH�n�~�B���� E�G���`�ͷr]���N�M����Г�d����
Tt��+�Nkw�E��[���G�����ב�	����A�&�
�\�n���W[l�-O�s^��Jt�ag�g[�n���<�L�8_��u�K�7U��Y�če�gs����$6hÒ��FW%�+��.X����ϥz��M�$�{Ep��_ ��~�XJ�<ãF�5�ty
8�dJc�4��ţ�	��B
�ɭ�Cv͑�_(^ [�P�kh����)~X�F�z�Lf�����Zۋ�Tk�na����2��� �L����=H� �g���5���II����AD�e�'�v	cg��u��Vz�-��������0�=e!	߸(A��CU�ۺ�������kN�<�ԪTz���*#dJaDlCuX��~�X���/�3
�����`����bU�2�R����M����y#�&}��[
��z���[A��-��64?��@�Q�1��>��e��R� y�`J"s�ro��E;Ì�9^c23L�$��	s&��mSxO�e�^!�]6ܼ�h�#ҋ)�1����,)o�h|�%�Y�z�=%�\C����{��/dOG���v��_H��[�'�k�v��`�%Kkt���e�)a$O"���@�=o�k�q�M�2-̯j�y�[�M�*�3@�������wNg���9������Kweɞ��0V���5E=ˣ�9!5|EI��Ui�3|��8�o+.�sr�1����! �?�<J�ц�c��bڗ&r,���m�0XFTJ�|��`�*�A>'��?�'M`&6�r��>�ynE�5�g7:�mC����sG���(U���e�B>n��5%B����!���>D��˅��Wb���
h���&qX�w�S=-�J������֜��9#B�UI�/�v�.\��A���	���+sY�(��6Ƨ1�!u! �a76�Ua�>���\���ˀ3���X�6fjK��0ًǚ&�?+%�x��P�����m�fM^X�i���>O^�p^�8���GZ(�<�N���S�>���oN��݆��+݆���I��r3�b@��8��
/я�j�Jz|8ꁞ�M�C���Cf���R-On3�L~���'M��tM}j��sn1���R_��o&�<ꈣxM24b�,�Ŧ�a�wD���;$u�ysE�X�RP��_F�㡷9���KE5q��ء$XA�yr�?m��d���a����5���]�i�G�jS!�ũh���7�	��ߋ �?����&U�r���� ��{���ܴH�pq�A�Q��=R��m�#�44��A���f�	�1�����b�W�� |6iI���[L��_���y��rM�󇲂o����}�՛"P��?d��*�t��b���*MDC�L�xUJ/u����a�앆O-j	����F��h���]�<=�Jݎ	���R0M�߫��;%�o�����"f�z�q��ܚ�����C�/�kyNlׅ�O��`�gە:��ϒT@�_^x��\V����M���|�FP7X�U�q�t�I[mM�4��y�z6W<�W	��d�|��u���l3�w��T~$��~�� 8Z#Zt������Z���=ӢW�l��)-������ӯ����n�׈�l��YJ�
UDʥO�d:��w��(��J]_��b�,�H�gR�5'0���
����s\�dT=_X��o�ceD�^#����B�l�5)��Ph� �!U;�7�}���yP3L C��<�͗P�9Q��Ѕ�$s�O�+?�F�io��� q��g�ѩ�g��#ԅ$Ys��!$a[C-���h1�'g����%?�2��.h0�0�,�����},���ˏC�Y<R=8���0 �w�  ]���HI���������L���>%2����0M�i~7cr��7Y\�b<39���}&��x�����#g�g}.:qgs�t/fI\����X�p���	�\`$��Mx���\I9$_Ek{�a[�P�3j�|������@��de}�؂5���笵1�Z���?	@���p���ϓ-k|Ф9*��Ê���ennBf���YX��EB!Υ6
�뛝uD`��8���ɸ+��O��v�=LY�%���0�
��؝���VR�a�b�W�y�Z��'Vq�~��D*�2r�����&��4����,>���2M�|y�d�J�1��s����c"�,�ap���=�>M�ձ�=+�d��&�ԏ�ݚ$��*D����˘�=E���
׼�S|����
�m�EC~�c뼆���s5-g���Ã���B����^#1��*%����9r�>6*j��MW�����.F��� ��-������&�Zo����D0�R�G2�,7�L<g�# ���t�Ҙ^�s���Ʒ"�4��?꾶g�?���\�zޢ��A�֗�9u) $1��ʰiq� �^/�b`KS[��[�g�謕60A���6e]�gR���/����,Е���Y¯Z��j�C�2u�S��2�ɺ%����2�g5�ΕH_<�7��5Ż1�ꔰ�C����T3����P�R�	0��I�8^��7
�g���'�"5������7�s����Z�dT�IF�"����{*��m�Q��S���*�V����s�aqi����hz�Z�������6EƤ��LF<��#K?��;�
��}Gi���l]Q�(ʶ&����bEȆi�8�N�P�K��F[��<*[{�/��G��YN�߃����0��Ľ���$D�lΡ܈c��➊���gsC�X�[h5�a�L�ޯ�nr{���Vʱlw���a�
�p��*�iN�������$�bn��y��^��(�7o�~�i�~oH�e���*�I(L�{��3G�����S�*�q������Β�qsB�9�����#.��V_�X�Z�m��م����$��N/���$:���մB�)�k�-d��L�}>}B��8к�%����>�V���:���g��+t�.�'�LV���+3b�ݕ6��4�u�6_'��x��.Rjoq��ps
�c��(P�d��~�gld%4��o�ޟVZ��Q��:��c��a� MX5B��� �?"N!��f[�hs�'��(7J}6OfW
~�O��fǯ~c�wj�/TV���(�H����)��A�{J&���������<� ���}ь�%�����	@�o~կ,:h@>N�bϖ�l���~�_�l�� ֚�*�sI��D@��^`c{��M��Ǘ?c������Éb����{��]y ��,�z�����0T$��pN8��R$�	�(�D��#]���i0\<P�4���<�
�1�-c�
0�R"~̝�XK��H�2���CԻ�y�2ƆC NM[�)=4�*��J��z������>�A|�jt�0���6Ġ��(|�G��Y��[fO*�L��@)O�E���N�V�>N~o�I��X1��h���E���h�"|��Z���6�Lc�� �C���k�9?*kbss&Ͳ_.�����n������;�J�D
�>�jC��]bq�$55e��V�'���*7?��2g(C�f�lp_c� �������^pyq��$�#x}}h��ᘕ�f���;Cv��Ny{_Z��O�o
"�3��|Hm��4R
����O*8����D��I� ��\��u�r3���Aу��h��q_R\��jmq��:�-��1�N��'��
\̺KE��諕�7�����W<{��%ԟ��t��T0�q�g�~]�a7��m��D���A���������ң�H��`�s�ǔ1������k���+f�7���������pl����USls�"uEI�"ft=$��"�B�w@�W�Re_*]ڠ,@1�MA)d�����)�P�$U�s]�P�	y��fc��	7�_R���W��g��o�����jI�a�s��D��F��n��V��.���1�;���.W��B���� �@�!an��>&%�:�\/jnZ�[sO�`l+:����pT��.�8��K�D�Y8!�v�޷z#3z�$�$
��a�@Y:?�[uA�%�V�⭙�FT��L�'~��~�A:���F�T�W`ق2(�����.�ld��[�8;:����E�~��sOi:�7��xE����o^¬f���!a��ދ��1^�.��]�I�FЌ�I�U�z16�S0��!�N$q�B����q�4d=x�wrb&�Dl��zR���G�5q~HSJ����݅`�����NI�Wd-ڪ%�ͪ����� �*�L�X'����������!4I�gv�� �7|�l���;���ҹ2�%�ތ��Τ�qh�B�G����|"i����\@0��T������΁�=%d�{)d`CT�'�ݎaM�~�;TeF�#YjC������:�΋������y��OE|Cx�5�j���Ry�|\uʗ�|<���GP�i�E,Kb�-��o-���S�g	u����b)b48�"H3|4� ����l!����gl�&�x��D���+����y[y\䟼|���*pa�S�h�2��H� Cs�nP���â��ݚ�mߨ����\��^s:�J2z-<�I�����X0�Z����L����>)7k������VX�Z�j��%_,�U�E��}�ixTwT�&�I��H������]z��Y���0d�i|H3
��/�w��؁�8L��Zr���i��j��,dm��C��?��I$?�"F��^�a.I�J3��6�r���w�0	��2#|��ؖ�|�E���Z�@��BeB@2�������c���ݦ.W����^ŉ�4����ie
�3Jd�4��F�h�L<Hz��(6���֔�&�DJd�2P�� �&�~>�3j���O���D|?7�b\�)��LA`�+n�8�.CڮR�Z0�4cq����9�"��t��8�.��aB��qǶ�
����$���61đ7VV�F�j�>�	���	������{�Z�����K�WoQPŚ���V���IFS%3)�j2&��!*0c�8�u��F�^Ӳ��u��/�4����!�����-�ý�9�+�Kq0�e��#W ���T��jTZ{�G/�!��"v�I?�1����s�t��&�c]s�T�q�[��`rL������@�#`���Od����^l�)��⢯���v8e_��2�H�10oԵ%����3�f5�� ����&�~V8]f�oǋf��V�U�G����M��篟��Aڶ"� ؤ̒z���e�C&�f4>�
��3��|��L�gٶ`�^�]E{�+��%��%��c5��VQA|2�[�i��e]t�"��v��6�|�μֶ$+�?��[��4#���o����Yo�<�ͷ6G��� ���(,��Ԇ�ƨ�w�	ڧ=��w3ib<�|/�� ��֓>_�gm�N>'��xaGGA��4�x�ct�R���(c2�Y����Ӽ�Ǖ�I��N�
~��0�Y���/G9�;�����u��}��A�#��
LS�*|��4�;@�[�R��#�և��V��m�r����!+�h-@��5=!щ"�����n���?�^��e�����RR&.��}$�kc��ƹ�R�����L/<�Á���F�7_�n��ſUk�S��&��2����s�iV��&�eI[	�S3�:G� �Nz���4`���a��E解��\~�,�dn��`���l}�Z	���n���w���s�l�-$%�%���z%��lb͙��8A������R���/��ĸ�]�&���4"}�I���bE�t7���1�:k����*��a��4
�d*��-��zP'q�-�uW��g���zh!�U�:����w���z���Xy
���V�h�/,����37���$�k�26��v��;���� ��D��]Ç�j�Jh*%s�(�/5m*=W�,NG����F��� R��5@�j[k#L��k�M<�w���i��}{��Ha�8w�T�F��g���CEXk0o�>�K�Y��7I�S�W�>�ȌcB\��y��1t�Tӷ!�K���` x�&=���
;F3G~/j��ß^R�g�K5v?eN�o"�3�������[�1$0�r8�/�\_?f�
T1A�M���Jw�Ӕ�9,X�O3!�>=�����Ɍ��W�O��A52�!��A�Ep��<龌��,�t��?�ۂ��0�7��S�?qN��-���������3��,��6���fL����q�gZQ�0�.L �&�{�3#���8����9~�
��S�B�jEtv_��̀qA�A<19ZAܗiPX��On�����9zC	���c�J��������ԓeu0̀q���Y��@��W{/MLRtr������dQ+o�"�\u,*��ח�؟��Y�n���m@\p�ѻ�[���|��Y�ck0���H<wL�c]g��/�7LE ���VY�%,M����}�Q���-Y��f�R�ڱY�x-�h��1�݋C������ɗW|��\1���h�
�?�>�T�³E�人N�S�]���/�
 ��a�� �(��)ζ}E�5��o��Ձ�d�pfI��[ıM��b�!��On߉�$mܱ��ǩW���]3�T����5N�k��m�H�G</$�FɲMM�+��07r��֌xϏa���5����,8$����7탘+��8�k}
{��#�O�ċX��:�s@�W��"�	v)7R�Z� �������03w��w��
��Cs{���{?�1p�"Hv�sc3	?�	����w��J7XA71�Mw�_�C�-(��O?4N�r�ԭ�k�/�)��>P�K$<[f���:a��ϵ���+�T�*��P���A{�b�M�r�>rZ2H r��;���/��љ���=OB�r�󤷼��9�'پ��P.�W�v- �=�`�z>vR��k�*��piO��N���z�ZK���
�謖tj��6�mgA������Z0�����DEr������W��:���C�)
M��z�x0wN��c�K�0tH�a�}+��7����̇'侂���lr��`��y|��*�Y�-H��/_I+ϝ+�/k3�����T]ۓ���VD�Ps�͵����3�JW��8PV�#�Tw��_�&<t��0LX6z���si/(7t������I�C�_�1`A���+eW��jF���tF������l��fR��*p��c�z��FR��i1׮TdP���W����(u��U�ouI����I�B���<*Yʋ����ܶ5B�?���I�+pϿ��G�߲�;}�^��:��5>g�f�x�햡(��6��J�/�[�����<:� �|ڤ;��%�Q%b��_�	Cv�16��1�}�������]�o� ɻ���F;��]<�:j�!�ǐ�8�L1y����`��m�A����7Ǳx�X��w}�ÊUpݟ�g��u��|0}��g��`��
hE*l��(_+��3�5 ���(��bL8'�IX�����(�����]���y�]
�yr�Q�X�5ݱ|Գގ�DJ6� 5�)����R�t"⦋��ݩ?�%��95�ޠ���nz6$�V�u�w�K����3kX8� b5�x�^����=L��	 $*�%�t,�#Y8t�[L�v�|`��J��+�I����ђ��|��R�I6�Q����'}�W��1�k�o�~;Oj�]�Z���%3}1�J�����"ճ�j���0=��Uy�(s>U�E��4�n��`�b�M�d���CF>������L]3���9R݋G��EKA�)RCY��cO^�!ӻ{N�%Ֆ��hS~��ʋ6���dņ�O��O�jT��>5E�x�m5����sH�dދ|~�y��*}Ko
�}�R��AД�S�a��.�#�q���5�!O ۆ��/K����бn�$���$d"İ�WD�sȋ�Hg�b�!�W�������>�u�6 �Vn��uJ�f��>=8��k>��w��3��d�5w��5����/o܄IL�W�������ȎG��!�䡰�XS_g��鴧��Af^׳��Y�S!���~߬C_}En4�y��J%�� s.�Q��o�t�.^ ����P�r�9P0~���{$���CuS�([q�S���0�O�!P/�7�^xk#��i�2N깉)���z��Fם>�}1���&�&���P�v���Cu�<Yle���ףkZ3�ν����1j�t�v��(Nv��hK!O�[k��2p{�7���r\��<@`�|����n�v �*@��/�f��ko/�G+[Q�F��bgnj6Z��;Z���"�z�?�/�����.���l��/
Q'�.	w�܎�_�v� 2j"�t�i�ޟ��)���XD�����'��f�!�x@�hV16��9�W/���L�p�ˬ��G�7�����v�I�ڍ�<=&CY�
�P|����C'a!NȪ_�˶�:���	�˄*��U|�2HB�S���i|j2�Q2����1iV'����^�q��
�U��.�h[��m�l���#��ȏc�N��C�EտmC���4K
�@֨�rv4��5��Q�|#��}����' I�O~[$�lhltS���Ũm"Q�7a^�?.��ƈ�zc^�'`�'�~��H�r�#�ߥ�9�YH�r�˹��mW]t&�
�10G�-��\��ڊ}g�w�TD���-#�̾8p����K�I1�0i-�6���*����-��g��+@��P���s��⤛�5��?� ��мH�GO$~ez�M	R����$OREt�>�vw�1'L��QQ����AG�sh㬨�F�*N�?R�7��s�p	��L��E+�^�c�.C358���Q<>>��RD鼅+���t���/p}D4���t�|���RtF��G'�M���~�h|UJ"�]��k~���^A&�<T?��'��E�ܫ���"��/�/*P��><h^<wNDa@\�����z�R��9Wt��:"��S$R�dw\�o�5nB�S_���\k���J��^ n�j��Si�@819�ؽ|�Ҍ�I:j�m���a���a'��E�ě�����?~r�%���e�rQXx�h���M�6ZԺ�(�S8�w��-н)B~��o\E����F��NA��r?���H��$)����/��g��L9ή�����}܍+�w�X)���F�������7XD�?y�3f��{5�iNE"K�NA���ţm>u( �"h��/��X�DZ�-k6�5��a�^jˌσʂ�;B�0��UT?����s��X���Ar��HSUx�ŉ��[��θ�Ӎ(�z����4E�� d���Ɔ)1{:��+�z�jYv)$��N�m%4vk����D���� R�T��P����Ĳ���|s�ʞ�z,Ё�"����ķzc��E��?��4� |��A�w�u��X�c���Y��XgY/�:
����4T��IHF=�X,�˦b�d���c,v�Ps�
�F���*�鳅��2{>��n,Θ��/T�D���d �bP*,vm~�{k��x��T{�^�z���r�Xm 96p�!�˓��~�Uz�(o�\!,�7�/!����V�K٧�
�bG�"����y�$�xw�n��	Z��]y,�`���kZ �%r%-_9�&�P(�R�'�$ wHe.�� ����ˑ6�+ri�/^�?ٹ�v��	u
#���w1w�-ֳ]�Ҷ)��q����nx��\< Y�ɾ��A�d�S�;�� �s7�7�����R�����X��Ms� ��"��W�X�0&僴��#i,�{2V���&���o�g�4*7K#�=4�j��V��C�k��Ǿ�����;�����k�	�(w�$j[l4l���'����p�u��k+��%N�r���������;o7F����	��0ez);[2�1A���Z���(�M�O���ǞΧ�G�E���%Umd��N��D�07�)\MYϭ���*�Ԣ�h��Ԡf�,)�\��D��x�^�[K�ַ���}6qq�<�h.C^�4�NZ��X�<Ϝ�qg�&a��F�Vq��y�Y�w�Y S����3�e9t������v����r�Fִ��3��H.E�;���Q5�4�dHk��B�����1 ������H�RN��ȝ�h�SI�7bX�3���e��u-�������l���pzd#��*a�O0)ढ़� 4�Fۯ}z��A��>�'8�iy�������F������?��͒��e��Ww-�8��B�(�y[�ғ��pw
���d�tl1�6�| �G�na��8�'��6�4��`�����2�Əxy0�ݝ�����W6��{�o⺸��Ò.��,i�F�$�ݓ�R+���=J�T��caH
��1[��@8��e��a_�>6�@<S,�N����U"n�i�~N֪=f5ԜmsQ�����S�р��w��GS���k�վ{^���BA�]���2�}=aGN��e<hum�I�q���AY�����	s�5�s\xus EX�u��w�W'[�Mz��4���fQ:�ȇޒb߶ֈ��_Z���W.���&e&����~�`�8�E�z�vw�1sY�����UzW��3��\�N�L�Opș�qf�q���-�����Ҧ1����>-�cc�i�a�����ky'Q�@���/l�Hsb�iv/*o'���Z�(z�խ� F�l�7c�eX��8���Ӎ�Ĕ5TA�/�/O�S7
һ����z[̭�<7�[9
�G����a��Y,�a�H���3l��do����ȏY0p��.�'}䀬׺�ݺ�۬�ziV�]ed��ѱE�z]\"bSF���\�T��~�:��_�lT�o�_��`�:��ة3��s�">��s\��^�ԧIű�؄��3WK
!�s$��ګ�Q�䂸�N(w��B|,�5Y�v�p+��Nq� �&�&vsr�3�������A���!읪�:|��������^�y�c��ڦ�i�v��_*$��8yZ��"���5�fg���=O�P8����W�Pr�.�y�Ưw����?�C��E��/�(��I0�Qu]Ba|�8�w�qB\�m���:YI\B��د�ȣ���)D[A���8V�C_���
e:`4�C9��@z�q�r)�?��Hֈ|����z�D�"���~(f�i$-��-j�Z<�#l�Ϳ_��ǟ	 swk��I����EN^<4��]B��A�ڍ��ڗ��m.T2g�<�h���:��� g��q_͗���6�,ՓM?.�	�l;QO��G���(�!!
�����1�¶��B�A�.o���x$�P��G�q�L��-� r����q�Yt�Il�f�9i� Y(D0I����1��lmb�3=����Ig��Փ�{��<�xD�Q�Æ*O�ڑ+�z�����1���rS�M[$hE��}��t�Gj�s������"��t<ƈ�jvJf��U�����8���D�7m�֡�Š,%��;�^�W�'Z^ ���~�����o0B�W��pQ�u��Ƅϐ�V~��f��z�0�SS�A3٥�F��-���k� ��IY�ِ�ܖ���VQ\KяA�a��`���T����������ړ8��o��~�˶�a8�(̕�?�=#<�?~%N;s��&��Ҝ�pz�F�?md��IƵ���뒍�O,����Vǘ���O��|��A��z(�ב�ꓯ���&G7���G:�I�f�Lf/N|\�9MB����p;e����r�Z���L4�� �[wv#�t����)*.!Q��l����R"C4��^t f�q)��h5�Z���� �P?���/5����tl�f N���+��D�X�C����4Bwwu��G�:��=�ۜ��x�9��
W�B� ͵��NUމ㠱:(�ks���4 ��8�A��j���9W������e.:�����s"�g�mݨ3��%j[�����K�"QQ�%��5q=#� ��G.�g�b���e���}��n�F�M	,����d�B��Z�ƭ���+�Lt-cU�#������.���7���jb�M�b�S����C��
h}��T���WCs�5�L���̦�l��%6�"��s�$��m}�MxuBm]3�?oW�2�/|��s�K��\Nj1��R��[����2���9�l�/�qKtj=
�������}Sx�4�� �>^���'вz�
6�!0p�Mi~�e,b���lL'��(��ӎ��r�W�������.�j���4�jأ�R��z��b�d�Mp�!�؛Y�2��U�;�}C7�&^y��S�L�=�*D�c�p[8'It�E_����}������V��D�f=����5Mn���"9�СJ��[!��pVK�Q<jH��w.�Z,��[ K�V��چ(���x�h� �T�2�p[��
�%��j�}h��dovN{]YG٫�i�E�7%���[i9����q\}��诮z:�v]mfW�#�(�S��)+f|���e��߄p����ZH�)_q��L{ڧ�#%�^�d@�;��%��B�{�y�P��m�Dx|r�����Q�O��+T�ŇD����g:�0�˯7�{��(4^]�L�����`ZrQ�?g�f*�&~��iD@׭h�4�]���Ǉ��X���#�a�
b��O�R}#?�
���M�%G���ũ"�����F^6�Ʊƻq�
�74�3�BvT�2�tA�_�:K��r�(�G����B��=��*�4_���8󜦺���2��p�]�@�N䢶� �3�k�'ɮ��#����:����Ao���6���I��<�á4��ݷ��:8�C)=��]˭�0Bb�Ȉ���r)^}�d_�phe�?�-�:�/�3��D@�_Y 1�(��L4	_}X8�L{t>v��V˗�,�n�*PJSۙ�M��6n��f�A�ꖯ%l���C�iE�m�K�"��ka������_�erO�H��e��0LtW��%�
�p�9*�&m�P��;yB���Ww�a��l�̟��yNL���$����ܷ:��ޯB����SG����S��t�M�6/ic��,�tq�ZVg_/{+��D�Tiǰw���.;s��d���؍�*���hT�.t�U�jί�N�fDCO؊'}Aė{��锛��8���}�/r�.}ԉ��V锤G�	t8���aL��ؤ��~�0�7}���J.@�Mv���H�	����z�UH�5�O*bN���lUٶԪ����_n�Awn����z�``����j6$�cbq�?��0Pͷ�s�Y����s��ގ���e��A~kٯ��X�� �H�[�+u�����C��n�R~��#��L�x̎Dt������e��fs�Ɯ�0�����gz���t��?��ػy�
��d�N#C�2����Oa���I�t�m(�2 D*���I_��gd���2���Ays+&wDS��^$�B�M�άa#�t�3����5Q���R��!s��#8pl�S/�F}�I+ICE�t�26,��6�M���'�=��(WS&�V�n��݁*��Nzڞ�O��O��&�+��<�L���	u'q����X/�b/�K�Ru�^
g텄��G��x����F�Y�S�u=}ΉS�(�3�;Y�"gm��&�̸6}����M��l75ե~t�UA�!���7������)[ŷ��j9�[���#��|�c+��G�-�����sl�ޯ��������Jvw8˄���Mn��-�À���`e�= �.HRI�V��FLH� ��Iӛ�
?�50VX*������V��p@�Ѭx���{�	�^�O�8�ɍm�p^xN*<m������d<K�^�6�M���Д��?w~��}�r�u��EФ%�ٚ������񡴼�#{��G6��F���Q�!fd��*jkdÿ?&_������&;Zц0��N_�(�z,�צ�Q)b���|���7��Hen�dl�����҃���.'k�z;WH}5���sm���X~�@��+���qÕ�������t�G[5������B'���\��"t+^yN�����k��s@>�or�dd;��k�m�F�pk��:�	`�U�����F�i^���M���^zܯ�7Fp�i��3�-� �:�MKATiv�HB�-r���U��>>���7���8(K�޺�I>��h�h���죯g�7��w�إ���}���֙����]��7��l�M�U�D)����ä��"/Z���^fń�<#p=7~'[�+ ��EY{)=J���meTʥ�����[1�f~8IW���7_�bpg$���V���ʙS�'���/��~���J|SV�G���B���r�=�\��NU����4���u��
�l1
=*��R�+ݚ��w`��Gq!"��-n#S�/S_"����AO���E�?�C�cǈޚ�oȀ�~V֋�E�l<����z4���ku��Ə�s���P:��.���=������\;�Í�al$��24����.�7�����s�y�LXqο;bn�;*�7�s#�����>y�x: ��J�-��S_���B�˻�(��6i0F�0 %�2��[����4���?�ڷ�E���S�����iC��lwn�7E�30uBU��*n
��q3���OBgŊU"���<�!͑@EXX�~ 
u-%~-��&	�����m��D�����s�a"b��q���l�*`#��b�׵��C	�g/�˷��"�!R�]��)�ކb�b��D�H��;��'8�[�x�1�F[OA.��O�K�ȴ��$�UN�H��)���=9��i���0K�I�7���ۍ�G���bq����8Щ��!�����Cŗ0I2W$�U)�������s��K1j?���i�ԥ�lUÆ_��=��l�o����F���G&��i�������9g���Ф��[�EͬC�����A�c�9J�7�ĴP�uoS�=�5�B����"���� 4т�h�/xY,c8QS��g��|��-�9�'e�Wv�#�c=4[J�K],WCO�vip�D��h�!����O��n�gr�Z�H12���w�#���s@f�Q��3[��NT����y��l��!��.V�c
n?���L��20��<�t��]c�SA��
�2�>{�Q�Ͻ[�U���>�Q,�o)r���n�e�ٯ�\Ϟ��7i[@x��&W1;�Vk(�8�Osw�r���F����݃  n��/��&�0�V��b�� �k��7NM��x��Պ�m��5m��M�B��SɣD�(� �i))�"����fz ������4�'A�K�q����m  ym�y��0C�7&���,Y�QcKę��/.��p*e�{�o٦6���Z����F��~eY���/y��)!��{����&�K	%��ٲ� ��9w��.���(Z���~�G�)Z�8�l�Γ�D��/u�q$9�e8��Z���/���2&8Q�ʭ�cf���0�!d��9�7XX�Q�Fh��qSٸ��P�C	!%10;a�6�fi��GSA�▿;u�+���]Ѽ�l�f��Ԫ�/Ꟍjk�Ǣ\#Ϟ�+I-o�dg�C��׸�>SA��h\]:�Q�������M� ��c��0U�_�Nh�:0J��0����.$U�S��)�v���_GW�]T^���!�	�u��o��H�m�+�ⷊ<�~�~�'tf9#� �����y{
<nO15��ߤN4��H<t��b�b�Fy�MY,/�kG�.�W'^���P�'Ɩ-�ǜP�@Obr�pQ�:$_5�F=��-9��%B���@�� e|""��Gre	�a8v{�vv�yV0��� �P�,y����H��_6����d7	��)ݞ��R�����6fI�fU"��'���08�N��\��������/Y��f��WY�.M%�e�عz㣜]:�R[����P���]Z:?�lS����*�N�'x�g��/�Xx)
U|��3�Uݖ���4^cY����N�{��~1�<�۱���(R�p�DJ֫[�@h+�'�,�!��^�D��^<@����������?�	���>+��H�Ô]W�q8N��x�#6%B�n\{HҦ�) �b�S�G��~Iv�4�9;<�b�� G�iR ��2 t��k3k'�k�%�����)�5��\�ڞ�m+ac�e�b���؍�������a�ZUJ��9���s���s���'ڂ;�렡��p����G3�TY�-޾$3sb=�=�?Ƿ��E���&�aG��(9�o8J �fQ����l�h�k��	Ò$K����*EՇi��.��W�P�|�_����)'׿�}v6Y�Rb�G�hۃ ��z]��[�>	>f��t�c��JIJ�ܧ%"n ��J~I�����:�D8�O�T��|t�$��ӒB��Ν(�W����{��y���G,ɾiv��vx�vu`��O���t�y���2�i�����$�_�����ӽ����Ar�Tjh^�Ea�P��W�����Π���P&�Wx��ϱt@vm,�Ԥ�4:)B�㚯��#EOR��F�T:�ip4�,�o�{l ������`���=m�k ���;=YN?�4m{#l��	�3YM?�q����r�q��\dY�������l�?�94. ����2�ۂ���2�����Jx�8�O����V��Q���R �dvY��H�!\���Z��>x�Mn�ӛM�9$P������o8y����l�T��134�[c����0�I+R�'[�#���'N@ژ��ďt�������wM �X�^�{��Dt�!�����SHGXG�`�����p�W�]�-<k�F����
�N�N<2.�OA���K(��ˏ��4v_�x*|>#&p<(u��6G@ҙ��?��SZ�0��X��c'#�\c�_�� RKE�/��]�P���	٦����)X��uDS~��H�����<�r}�T5N�!70�����&S�N�����ǠWA�d����}�U� ^�'C���0�����(x-�f�EE)��K~�3{���bD�v�ȲT��4��R�GA��׺�R�]+&u��x�2ٚQ>ם>�h�	��F>=���vS�{2��X\%t�4�G6Y��\ŕ?C"$8�Ci�c|�g��/�ҝ��u�sR,��RM7U�q���ˣ:c���VmX)+�L/"I`�G���*��M�r�����C׳�����H����)�jF�1ݲ��Ւ���n|������d�?���x��9�R K�����/���+^����}���l����4�	�10��DMv�挂����c�2g֊L@�	�Fa7h2�#۝��K�/�I-ߘ��&�I�HQ�����M��tE�?g����O:�d9R0�T6hA0�'x�O�g�.Zs����(��_}i�8_n(�;¥��N�ٕ3E��H�}׀Z���J>�u�tgN��;T��@aqu��HZ�ZP��j��q��I��]���+U]�X"��/!;=T�;Z[6�r�{���`#w(�&KZ�	Y����1�JI�q�Cl�-6D���#������`�A�m+��c�~:����њ�a�TLV��l��X��{�H����l�
�|��^�*���N_&ֻ ���u��$A�$@��)MgJ%�I}�ң���q>(ō��ؼ�g����ۘW�e>�!���H��?�}��t�9}���J4�C~O�������Ԙ��6�y;ɫz`L��oS���56j9����g�ؠ۳G�c�@�6�S/XO\E���Ua5Y�/祜�yk#<��|�������a�l�z>�4��sk��>!֫��3��;�) �H�݁ڵx8��q_#a<�A7��K�Q��9�9E�8J�>'�d ���ނ&�C�M���k���X��^��-��*�НH!_Y�Y�h�(��X�9�<���xFK�4�Rª]\:>�,	wx��an�KY�+;Z����	���h���_�9�E��B$u�iV�IaS����	���|֊��"����0�̓��k2޹�?8ǻ.�jM�Li���֗���
]j�0� �c�ƪ��X΋7����,��x�k�
ܷan܌Ԑ��Bve�s`�����G@�����k(����d�́u����R!��)�L,���0�V��g��GVxDj��'�+c�L�$ Y�Ż��=,�{V��PGX�~��y�B�ޡ�]��Y���
U�錝X��m����{ѯ���m�n��u#��w�d'���>�(N{�@sr.���@���=�?��ͨ�mCh)�v����o���U���.�Ba+�uJ��v�;Źb\r^m�&V�U�J�9�����w���pC� �sB���!�P�Z��bZ�r���X�8�}0.��9k�O��{E>7{��^�)�,s��ח׋ߞZ��ö.�a��V�*�<��ܜn\c�����:g��l�v�l]��-�ҭ����FNdx�B;.���wN����"���9j|ҫ�����w�r���9��o5P��?�-�z�d�
 ��z!��raa9I/Ӿ�g���|���J�@�l:�eL�����)E:���Y��L2[`&�\�#wE���GmW�����1�9|�K-H�����
��g{���4�u�����a��K�═g���c'S�=S�[�[�D�'�V)L*re,�%�3ST������1ہ ����gI�T*� {NO���o�K���!\j�i�an��j�|�=s�g������Qjtt���sna����&<.�%S��!�p�.�X�8N�M�NE����\}��{O������SM�7�����Lz|�VkO�07�$�<��F��1˧�M�3�F��d̍d��Ɔ9,��e#7�z�n��c���?���\:
	�0ɽ2�+'���w�g�%�A\j��y��ɰ�Y] d����L�r6�앞�굫\���6 �K��7˘)8��K�.���f=��8�8`^��ַz iy��x� w�k��c��x���d��΃��5ޘ7"�M$����Β΋>J��mrｍK�U:��}�w稺G��:~~��5${؋�]Nz�BU��6�ы��҆�p�m#����/�B�J���༻�d�݂C����[T��52:�Cg�>��q^�u������"��]���� �����'j^_���S�C��d�Z����p��㋨ K���|����=i+@����C�'�Nt���h��"*55n��9��!��y��B��HW�����TA������9\Ӂ\Ng��ؔ�0�ŀJ�31�UIV(�-Vk�smE2�)�����kS�M#]�[M��{�=4Sv�;��ku���#صȌX�Vnlj��i (�4���e�]A�h93$g^��pa<Jv�ȥ��<��wO�|d�mgy'�]a�y���E�&��/�����@t ��߭�z�.F�~��$¼�T��Ӕ�l�1ݽ_������X��wy��b=�q��7@fO��k��+w�~�LJ����)_��Q����������s��~N2��69j��V�,x�]�-�Ar�����ݞ8X��rì�y�)� �i� �T������GD��I�E���g�?F��oL��eWȶ�5��Ζ=.�"���".����I�fA���(~��b2�c����m��1RO��Ϫ�O��x�����OB�j�PK�g!O���:�K\����G���WG���V��H�wT��*%��g�ۿ�wm�bHb�+�e�M�S��p�]NX���ޭ��������T�_.O�5�T<E)�-���$����Kv�ہN�
������ {L?)+ǩ,"`20<��v�W�jr����l�:��:�c]J��&7a��IP���"�x�Y�����l:j_޻�P�Y"Z�Z�����4�#���1��!�UIu?�gU��>u���X��[�0;ŤH��sL�����WF��.	�1�R6�-g�Pg�����nv�?Z0Lj�����l냢�biIR��8�w�*�R���)%��Q(�����|d~�]�B�<�>���J��=�lƱ�K݀�j$2~A}�`�k���Q�:�J�c��z�t���U��	�]�i�`J�_6��6*$sf��8���\_[��fzس'T��'��,�"?��2�Q5��dކg�&0�{}La%	��su����T�ͷ���رd�&M�r�z���}�m�u�D��g4�	�s�K��W ����V�ܙ�>ȉ�b��I��Ts�}�l���)�\Y�<�V��).��r�z~��,+��o��Ux!\���=�jm�ܐ��T�8��@PDF<�j͟�66@�3iM�r���F�59�<�wkt���^M��NRӥ���g*ws�V��8��4���w�=,Т�7�џ���?:����a��-dP��2u����+��8na(BA�E<���ґs_F�c�D�����E-7(��+��v,Oy�rzu�>��#�Z.����b25 镗���يM�XAd�zj��߮Q��++���A�����
A�A�;���|��#���΢9y�8��'����t�(�_�����gʑ-�}1N���xM�(T~��̱�.���|�̄��;M�H�ٓ����!W�^]'�Z��O�ķ_p,�d��4�?�&�$:<P�Q�Q��B�D�� |�T�%~ߛв\�R���cP��� (�d��aZo�5uQ�s^2�
l������P�A��%7�A뇷�N3k$7�:��u1�WQ-�+�N��&Z��98;�PT�Y�$�H�+����?MGw�輯�R�ȶ�>ؗ�[6��?��fr�|p��B�z��[����	z�́a��}2TnB&��lЂ�rD�]�1�*k+V{�-Zp����+�*����/�q�� �T��ɬG9�|�6����p�^	�5�&l�F�U�E��� ���ԜZ�g-]XŢO�In�T�:����}\'�-�����N��J�L �2B�6��xK�f�����`n�D2�,���.)r/���$��fҊn�$N]E�P�� ��}|�0t�j!:I��3A�4	�6�@-j1M��c&zsס֫�z���7�>��4���4:��f��o�Z7�,X@z�ݽ3�"ހc�Z-����E'�id(��N��{!@�4��R�d�qQH#$�nA���;�#�\y<��׷�����Wp����k�"����X�B8/4��,\#�I蜶��kϰ��+�,�����<�B�U&Ām�( ��1����������&�Ο�h�bV���GZ�Ͽ6_�Ǝ0�E!j"ţ�H�O�W�G����AX�B�/��l�Q��Q���^�?G:�׬C��|
�����w�٬&i�'u4��e�I�
 �c�W�����X��jeri1��������e:��]�>	txŶB7ĵ[�u��o�%����\�!8��G���}
˖�;�n �w�
�h��<S�Ne�9�ʱ��#'�ԛ?�u+���(^ߐ�+B����X��B���Q�@|J�dK?J#��̸���ѽ�#i7���M9���׭�D-�t��(�+Q꾍ͭ���ȧ�B�4��ɯ��U����sO5�v�ΉD+1�t��� ,p���K^ ��Wő� ��6D�����ͪc\���4�pi�5�8b�E	]6��a�'Ȓr�%�@��H��ɑxֱ	��i�K��=�'�v�b�����nV.����lf������g*�X�W���,����8��1��ļ(
�2�ՍO�նn���Tng3&dE���TK��0`s�[��;Kh,k�h5�2
b>�i�nS���xH��Wu�g��|wm�o�H�����N8�UZ ��d�{�ڧ@ʽD���~���'S}Sn�pR(���;��dp�F�_Y��!p�.�+�*��cz�G�%�^�W�t��M����&��򛡵��1V����Y�Y!��Oqg��yƈ���E���Pn�|ч��?�O��G%ll�͎*_�x��=�*`X�<��o��&H$��dSͿ�E��vn��뎶�Q�: �s�5�k��_V�H��O��t����/r��f��y�=i�/Yqc~M�¦��V_T�vN�rۑ�	=B�j�\+˴;�=�[�=D�V�߻�1J��yk��N1/�)�����S�aLS�GqK��W@��B؞�/O�S�8�q��x����!
�y���W|���젂�l���y�ߣV�;ȎޘhN������ǹ��s0S�օIf[[��N3� ��ȃ�E���^"��g�5І[�p�㕙���}�����R%J*���P�����*)Q����\?���sP5��S�c��k ��Y��C� �z �`M
>q�^��4��TA�n|�����_�۾Y���8������×/i�����"��fGS@]{���U�H}`b^�s����N�����s"�Dأ#)~!�z{�ߗ]!%�a������Ni�A�fO���(��P�e�V��E���kYz��:��)ŏlY;I��7���lI#�E���d���H���2�
�_f=8�{��.��u?Nμ��=�E�9����¸lb/��S�v�Y�~¸�t#�F�8�,}#ǃ�����O�N�j9
�3C��e���7Y ��'_5)�����w�d}�{s���@KPM��jpl�c�ɗz�u��n��<!��\���@͏ؽoC�|�?�{�ՠד�6�<��ANJ��Op{\�{}o�r��E��\���5�:���)����>�L�WP�hUT�����9��57X����G�pK��KZ̐��ޅ��V�9��諟���o�FG�7�VB��U����m�1���F��?h�֬�dq]q�R?�5^���� �-JQWLȝg؉a��=�S'm�tha��� ���L���W!U����o��%-��GN�V����w�(#��q��� 8C�+��i>[���I�U�D�c\�g��M�<�!���a�	*���yU�m��b�Jk��3�
�1�{��iCƞ��`m���٫�h����P|�9�l��"�}��٧}C�+�Y�����l')�]�[�}�+n-nZ�P�5��i�����f�^3�3ˏy�[���&�-���;(�X�p=�WA�K��ĀS����k�U�W�0ݔS�8�0�O4`F�V��u�b�N�e�G�s�Cq����l#��K?L�=�����)��؏9hau�MH8 ��F��*��9:�z�����:l���G��KS�V���\��.�7	�Dc�١��Є�-�� �N�Β?ܨX�(�Sm�?��W)���!R�/�-��'uX{���2H��<���V��6��F��m���x�W��-+�������<�_�]L/
x��T�t�ML�@m��R�G� ���(!%v�t��0b*,�o'��S���±+�a�1�ӳ�0x�Φ"ܑ'y��vl3����.�)�)�fS/�C��=<*�����/`�h��E�Md�����"6�^&��x��ԍ����8\�)�~�(�Q�?Bl���r?Z�/��#��v���x'W�,����v(.�#�Dqdd�P�nJ�T�@7�N@�:}���O8�?2�|��~�a���_�H5���D�&��D��;�ڪ�1B�K5N�Ԛ/�['�|�1mc�ޮw�����g�ntQElU\x��̒�?����#�-f%���{;+�c�c�9������ K'�С����)1�I�y��w�uO-C�H�1�0ji�LI�6p������cO������Ax��7?�MP�ky�7���	{���S��o�8�% ��`�kb_��u~��E�Yn����%5h�HU�i����Q���rkh�|k��S��|��O�,=b���&Y�����2h+!B�'���B�����"�`���[�Ia�*�|��鲠ޢ��1h�`oU�h!c]x���5�(�&Z�q���n�r�\yP�\5E��uZ����G�W�O�jl����qi;k&T�u��6��^��e����ZP~Cy��!�P�
&};�<8W��u)d�����?wC�E��;7<��H(�� ^�w)����FhJ���nX��G��;gb-4��<��*b�͑#��p'��w/F�g��ϯ�X[���}]�Ű��d7/ɟ�mJb����TӔ�A��Я~\��&���tY�kw�g���=�\x<򨵸��܃�(�b��SÒ��bޮT��;;�q5b�P��ڒ����X�3sP���ڐd�=���u]����,��v:��Œ�yE(q�<�๨����;@�G��/n�ɵ���3�6V��?CP��*��O �)�[�f�K:��Hw#���a�7-L�3K��͆i44d	�i���;c�9���wOp}�fΓU���Y��W(�jĽ�J(hSF����UT�t�`1���s	�J8��q�T:��*��2�6��8::W���IZw�s��q�6;W�s[��L��� Mמ�{�Oȉ[�U{�ֲ�@9�1Ӎ���R�,��s&�
�n��_���f!	�g%��X�.6�9���/�|I,�L����
7��N��b�v�s�:u�nӟ9�e�QHwh㔼г��y��U�b�hä٬��5����(�=9\M>kWsD��b��M�`Q�ֽ���?\�e�`�4|8W�7�����!r�~XB���ø��*�6�`�=7��i�nbP	C"��E��Π�@��&��!��[*�9Y�᰼@<��X[����5!#���X�4_Z,@��zp)�ʕ�@!��sJ�
k5��$�����άH�z�qǼDޡc�����V��%-��i5&�� +�i�������k��H����:t���8Q1�`��z.��=VS�q_��f� �>aoP��K�5��Pbk���]
v� ŝ��kcV��Ƀ�"��`�]�܂+�54�p�B��A��)�����/���a���X�
���/���h�Di���n>YM1��N̐;/�4j�����+��fno2c����kc.�q��#x��бZ�ω�в�Ԇ�9�j~�_b4�,��[��$jO@�������Ԭ#_��x���N�a����*�[�X��"TW� !W��4��J�86��g�Q0���I�*�<�K��4�-���j�p%$��qY��C��߰N�*�udZ}L����_}GYL�ۯ#��㜀�#C�1�)WQ6(� ����(;�^�j�oѤr& ��Lb���*�J�Q��?df���
Y�_d��#�N�!a�x#t��q���#�+<���r4]��i��.��P鞽��@dF���E���c��W����8U!n��H31В�]���u^�g��cU�0FeM���YOƤ	0�c�q �u�3�D�1�.{څ��9�T��m���r�cEfSD\��
�B�&�D�}&�l>["{���f9��Ҵc�P�%S�@R;�3�T)/y�=s�P1s��'H�E4ܱ�T���g`3���@��Z�ؙ~����9��m��m�R|Ǩ����~Z^��>I?Q��T.���З�L��*�wޯ��N��ѡ8�p�����_��5��%n�-����}a�)))��yP4lW!(=dN�1-���8�3���ݠ)o�5MQvܬ\���@��⟫$���`�� ?�U��7��1c�[��l�(bFB f������'���3$n<��ly�l��ߧ���a0�Q~�����[�5��IG��?�~ֳN8vc��fķQ��;g|�9�������$�£U��[��:�6.Oo�Q���֞C�D]c�ɾ����#��Lo놦y ^#��z?�Ob��~Z�7�8x�Ia|]��ֿ�yغ}�;@ ������0�59���]d��SR�v%E	��x<,T�}nS�(�6�c�a��j��7j��
}���KGRj�5
��y���ǰ�"Wi=��7�C1�\E����=.j9[�u��l2�h`�C=�{�~��֕:
�E��5�	���Gb�8�U��)�5�*��Q����1��m��|>���"Dr����R�*s�-��;2�B}|�yZ搼@��KP- <\�mN��"��3�r� �>(��M�o�qIA�ݠ3�q��'���{���M��3J�L��[$�B�q�5-�@uE��J�\��He�{b��#b�|���p������੍�"��\�]�2�t��uC���\��9g����`��A6�w�_�-Rg���r��_�+���"X�#[��
 �ȩ�\�1Q�J���9�&L��*^��zmJo&g�8�B-Z>���7�#�n��zMu)i��jcn����m�b�)�� z��������R{7�1��<�kD[����>j߫���\�����3 ���d����<��t��7Q��?��$��"3@<�6K(eX^�}��--�a��vX�^z�@=�L$�d��5�1*��߼������B֪~ �(���w�C�f���V��W�{�&s\�3��7V�ED<�p��4�8��n�
�J�m���솸��q� �����A��h�#1�+`�z8����E����;Ym������V�B��B�Å�\J��p3�%7�V$1/Mh�[�^5�> ��r����nN���Z���D����	q�p0X^qӰYġ����N������I<�mK<�O.[H�=�F�R�y;�L����d\�s�ʿYhK���v�l
���,��jS�G_�e�� �����} �k���}�@ y_�q��Ӓ�n�_��T�RZ��eo�v�j:77۬L��ޠ5B��Lѱ�B�|�i���@�"��<P��GG=��ɹ���|�k��P��J;* �I�1v,��p:5�*O,�ad�o�sn+H��kS��`$�k!�M�3���;��}yW��\��i�9�L0�X���Ї)��QQ%�rv-�b���IcA����8/A�`�``'��fl}'\O,ҩg���G`7�Ứ�y�ik^�#�jdN6폘�hؼW��w�4,��ǧb�*(g�����^�(���g��g��u�������D���%�,50����$|#�����u����<���䩪F�����"ͱ�9���L	�j�M�J�\R�C_�2�|��D{R�7<>{'��3�.��%�A��w�Ζ��W���Z�4�����������aK�R��]Zt���Itf����o4؎k���1ܢT��%�]����m��͋a�m��#����[��fQ*����6C,ۈ\�oEQc���Nk4���pƺ��P�-�>ƊD�/���v�$�)^�j�{)Vm?��=-����RMEz��f�M��eOGI�w`�f#��o2���-�h�kWb� mϮ|u���t�p�U�Ɨ~}�I��'�\Z�F?�лvC8V�� �_�EO�);	���u��%�H�=����L$���1�ي�u��M�L�=�s<��5x���{�+�e;�F�lGz:�~�B�N�]3�������}i��v������i���S'��{%�ܖ����9/���f��i��y��z�4rnCB3[f���KE&�BK��K��C�q�Mȁ����Λ���yþ�́�04���O+0�La)�jh�ύQ��	���*�$�Kf�-g"8������|�,��h�YL)�+�\�੺�C]'�		/�K6���Ɋ�_�����#r��
3N�Aȷ�3����|�f��p�O<��U��?'�����"��?��
���5�^��f�>2�I��M'��[=���,���L	��no5j�����!^Xm�PFy��3y��P�~������"�!r�2ѻD(\E�T�d4�"nr��RJCK����:��5yɑG;*s�x���eޑ�IE�(쥅�8,}��bW<��y�d2�.�
dzj�׉��5��y���}t�VU}�J���,Ia{+���������1�QG)�p^JnMe���|�OYDplObgj���Du�	�o�gE���Y��V����"U ��2=ʏ�B�\�,%h�1le�w���`g7���7�_i��cÓ͗U`b�os�Y��ڱ�k��*�D��~J5bUȢ���*r�i�p��o��\qdWA���`^%F�ֹ, �T�g�ԇ��Xf����pG£J�Y��f��vN����o.9�lH�W*m֌��_�Hs�"�Wӗ1�ȼ�-��z��\}2�i��>���6�qX��!v���W���ʾ�����֖�9� 4�����/�f��ݥ��KǇ^���j�Y�:��3B�=��9���B�!ո������W��]�(��$��YJ�Ck �:k,F\�����-�g�����T��#�Y��@$*�H�Ju��jZ�S�:�'�֌�(���X9V�׾5me#�¨dI��Ǵͷ��e�~*v�������_h���Ǳ��&��lMG�Gf�rR�Ԫ��i�}�a�SUfԧ3�,7�塤Q$��A1 �l�bK%��U�gm�g���V�����<����ll���6(�N���=�K���\�,$P�^�?�|�#Z�	��R_	��0I�F__R�� ��۰o.�T�� :٪�3pc��Z.�I͛#���ȗ����Xy]��QF��9�2dk���5�S.��}����r��,����oXBz��@:=Le��o��q����{#���q���Uv�mDP�V�~1�`EW��E��d�v�I�7��X*���(́f`�S|N=-�ұ��M�]91#uL;[@W���|����"�*�ȴ���cI��d�x{�p��|��G�vC���/��J7�4I)�4�Co,m�I�8�BR��S��a��E#�*Vmi��d� ���U�+1�8@Id'�"�$�>�.�=�q�(�KZ�M�Q*!H5���T�6��;�P��%U`��V���k��Qu~�\4>x����S�����E<����:X,x�0}ꢶrJ;���ƒ<�+�a)��5�Qv����S`wt�e�Ii���J���ڜ:s��ݭ��,��N�bs�yw>ܜaV��؉���k{��E����q�q���'?����rT��!\bhكZ�BQ�)�e��]-��;���\�e�y�CV5(Kc��v{�0J�=������ԣ
灭�>��^�>:&�����>+rq�.�m u��d���[*�ֿ�`������gi��W��;_)f�n��B��k$}��d�A�V��B�%��H�$�&J���md��h��>�Q��ig{C�e�3��#o��~J�n��4J�s��i)�J�,u���8��LP��NK�F�Pp�LA�}��E?-��ӿF�1��tdg���9�n�n�MJ�7{r�H�P��2-0��6 o|���P���}@e��OL������MiH����/�eC��#Z5|*]������ì��.,y3(\�p3�tK�jbl��,����e��M�^���zO�q�9�M�	yK�ko|�k��n�M/ʧm����)|����S��WȺO�u� �����gf��I�ڊ8�X��e�Jzl�R�.}�fJY$K���0�;����=�#�{Nٵ���Vj���J��)d��P���`�ڦL8Jܴ�&~q�VXLt'C� �ij�#�b�M,e.)�ꌂ
v�:�Pg K���ᩦ\>{�r�K���U�Zp�v������3�x�k�\�ݮo��m@�[t�-RQύ�2�, YVeRπ[���_�=.��)��qlS�}ä�V��7����Jw��}��+�{��ޚc�ď�a�Xҥ�
O#
�i���w�)����/)��Q��o嬯;+`<�q�:-���:�A�;�V>�}5�urU�k�Ɉ���!<�M?�q/F$?�%�և��^�5Dʹ������@yq�U�<���J�(�%�ĄB&�$�'���Eo5�u�RO�	��C���TT���Ka��>}e�D�;6��ϗ=4��ed��w񨢛\��C����@a��p���}��R�e�a��<y�PO�Ғ�ͤ0� f�F���`}��n��Ё�rۭ葰�HΆx F0�!���(F���v�O^��A�b�r��^��Ő���@�w�6j2[�Wd�c>D%K��t�Ȏ���)�P������u�s�o
y�z�dy�B��P�p�n��w��H«��y�d�!�&+���Z �_sz��y
6Ӽ��K��fN)Ɓ�t/�"2�lԻ��HF?J�#��7���i:�����L�nSz�(H?�@��L����q�@?y(9Ii�J�ַ/�|s�E!�����ԛ24ϊ�kb������9��|3�}"���Ec�eg��)��ph�����W��ٌ�#5]�gy����u��o2�h���W+�bC����o_p���DiP�ާ[հ6Mֱ���3��q�Q�D!$6���GS�b��/�
��H�m*D���C}}ty�f�p���(åV���Dp(b0-N *�g�ʪ�}����!�h��'���6v���N�Ǘ
�Ug쯒�0�l�Ќ��*�3td!S\���#�hy���pV�EOM��++"����Sk���dC�̳$8ۖdrhh���]�Y*�2^0G� ��Ļ����D�x�Ѩ"UmR��n��l,2y
�"��N޵8��>�X�e���)�8�}�}�b�.ly�~�e��_v�q��S|�����[���Ff*IA�/��m�2���ġo�IB_E��6��L�b8UB?roE_�����	۸v?����*io �8�^%��aF�-�j���x���]�f���.���	�������|�(��J�#�;����W�j��e� yo�� }�{��;1p�:�6D���֧��Q����@�`P0��A�/�44�x1�˽:�tP<$y"�9#�OZ�N��bƚM���V�\��U��o��Z��1�|,�T��sb�����y���[v;E=4���no�F��!̱������g� o:/;zT@<�I:Ex��y��:���H^����[G\�ˮ�^�ie��m�60W5xN��>5�ċ����'��|�;I2��+n%>[�a9T�QR���iX	����K�3f����4��$�p�n�J��x���V����\h[HD[�ߘ»�_���WJR�]�Ō�)R�m��a�=�"V��ҡ�!��s3�1�I]rU1��ߪ�O�N�F�v@�G�Y=�.=���z�D{�s�yh�G�$����lJ��O(��ކ��`��p�h8���R��q�<�w�p/����'�F�ķ�u�V��[�9�(2�*t(�蔊�r��˝��-Y{a�b�{���sî4��F����Mܫۙx��\���A�Z�d��?�=�a:԰�_޴��g�8�x�&��&���߇4��ԯ`���↘��F��
�E}8xxX���R"�U��p%��n�9$m4m�r�V��H ��������t�-<�=&�BV�皭;�2f���,P12�{� �͈C��������U"�E{b
�� ��s���ڧZ�_� �Zt�_�n=��'0�V�Y�D-��)-���Rg p����R@�;P{p��}��6)��R��q5�[Ϳk�)��DW�(�&�����8"��̆q��#`�|7#�73���?�=�7�6��(�:�)"�f�s��:��8?l��|���]?f)xĶ}[O:4yZ$�w&�ۙ��|-~�Y�CE�o���J1Ga5��ʏ��%MP(q��.�2Tv�"[rꭞM�b:��`]1�BPgmOH��>'TMB'X���Mw�[�g-+c�O&��O��7������z0P��1�S���%xK&ռil#N��%�I��m��n �9�:�h1�-���n�'��[��!C-�%�礀���Q��%u(�h�%D&�8"ޛڃ��>A�9������D���&�Ew��`V�Ɔ���W��=R&�^Ǹ��t���Ӧ�1d�`p�Ks�#o���&��|�n�DH�|%�ZϗA��hn�'�w͓r86���,y/	�ʌh����-��[F��u�.>���^��3��x����L%��+��!pz���`h�K��ɱʌ���B���� ��������˖͟�E�â��x��H��m#�=GY���wT!����l�ͧ�}-3�&>�a̿�'؀�-3
���zF�Z��&%�=R��^�ٷ�:��>�c�1Uً�](�r7��<c��cyl�d��b��B�����(CH�<�Dg���?:A�	�=��+�D�$����B��[:�̄���m��b¨�%��0:h�Iz��Dl1��=���E���f�"sh�I��~'M{9��)�>�3Z2�w��&8��Q:	7�{cn�x�Ii߼�j��w�i����Ы(���=̊��ʙB� h}=v�K=;	���u�h��Ϟ���0��ƒ��Z2�K4qV��k]D��:3eqD���!������󟨢$�fR��~��"���#�QzWm��ݻ�Vk�2�R2���6�A���ga�z#/���G��d �Ҭf�܁��׌î��#ƫ�L�[�k@���yJRc|�p`�b�ՆsE�]nv�g�+���1O���rT�g���7+�>��k��ÿ��ؔ��.M�	Q�6�"g�Q��Xna�Ő�J�O �P�)ݯ���~_�:M�ڣ;r�v���8�<�ł��Xq]�Q�]h�{3ɺ)�H2�x�$alm|]<*���'H�����I�3��[��6 ��f�
]jd�vϗ��#��zx�p��&��L�Ů�]o��J:�<���`�g��`a���?��"ϒzf��5/�e��Z���/I���R:x�Xu/ֵ�	�C}������Ű�ŞS)�9�;[��[�3`n����ޘX���,2��b
�2��02����e#�����d�	���6���E���t�R���ʵ����D����F��m���6�r�wg����.���w���zxl��KaL�ǲi��u�ϟ����������¥�h��ERS��%_u��hu;�ܦ�Pk>mf,r��r��M$�dW�GS���K��v��8o\�r��H+�9�/���}�F����2[�E������d�XٖJm�ۗƆ��-j;F\]K^X�p�?hW_ �)���r��l %�V8�p7%. c�Xs�ƍˍ���_��d�:o��� ��.ά�&�˭Q�y�NR�Ȩ�����]2mc�i�X�+B���S<�?�}�;��� é�p�){,X�����s���Tw�)�Bp}8�r�2�Ș�Ts}:,��n �Ȫ)˻�� u�]��B ƛ@�r�a�䌸2�*2��Q��4U)�#�c�*a0�Z%�rEz�-�Z�ɥ���v�B*�� ���p��e|7�?�ʦ�֊�Q�e�*D�nN�+y�~%5TD������A�?F�(ǖ�O`Ȗ�f���M���SY �����B<{K�J���#��X��D�'h�x�rd�Nd�߷��@����Z+�[򐛬� j�����w[�c���9X%}�(�r��p[Kd����B3�lt�-S�صy�=�eX��Q3�H9Ap�a�j��!��fn�Fw+�T:����&��[*�M����]k;��[��b�p՛����_�����VO�(�=�9���7JZ�+z�m�<mTj�����;����~8��B��c@P���J�ۘ�[h\;�7�Ç"���'CA�V*�V�ߴ\xT<T�^���M<t}��6�|V�W�T�"��c*=���+��X�M�Yf�R��CSO��O]Cے���ƃC�7��@Qކ�Z�5ʕ���?*9n�3t0���2���y0�ܦS1SN��g`r��Z�T�%%l1۵�>�.5�k��4��M����	�Ts�
�:��A5�0h�#�.@���F)��DK�nJ�2�hyN�!�m~�7�=:�
܅Lz��G�#�)�m�+#^n�šW[~��K���s|ru���tA�ȵ�-��������V���k�;��.��;�!7�})U;)�&=����5���]��2U����lJ�qz'"բ���w�L'p"���p(��D�}��7Q��-�0�u��ViAV X�W�,!w�S>�F�ւ33��Yy/r�L_ٜ�O��G�Agma�]$Ȗ���%���cy�S:'措�߃���*��lk��D�m��3���pO�^P�����
�R܏֧����M�@#��+�`@����(��6��!q��GQ�"z8-�V����2萎�W�譴�&mF:Dm=CG����HT����isu�غ�{;}��5 ���.���7^�!����^���e���3t��G'SK���/Ɍ�/-	��*�)�}Jv{�跒�����P�
#���ܩ]c���<�L��d�_ߚ�{b?�B�N�L����x#p�8�Z��E}0РMa�
T��т��z1�\�p�	�o��MuҀ~�)���d5�;��=e����V�d�$q��u����A&>?0��K�Yqm�7�C���T��$X�W?Oͤ���s	��P�(��H6�`EF�ކg��w�;��é�ƛU{i��h��O-dٳ�[�a�6���wY�T3���~�K!D��P�UC~P�H~�ͅG[�]з�MG�!�!�s��Z�f�b�&��
�u��6���fSZ&k&���e8C��<U�@�s`Z���L�lhFw�B&�{;��~�"�@�(v.���K[�
���\���s��$'>*�Y�����O־I��H����[�b���3\3�8Җ�^��D���x48H��K��}d?;�b��@����MgM5DT�Gb� ��L%����#e�zHV�B�r�۽M[|"<�C,�/�i��w=f2����P��l|̥�ck��h�nr�NO1�t��B�IJg��(���;[)��yf#�q�کJ%����?T����&��G�X��	�M�z�~9Y�n��pS�|�KieN�O���f�y��!t���#mdH�gY��3e�
и��G��xD�Pևv����.�'I͈�z�M�|���� B%�/�i1�;�u�QcJ�	`^&\��� �+���d�(�b��J)]�H����b<�m���~�� �\Ď��n<����������	"�N!P�;��#jr/�1h^�=vNTŚ`٬��ƚRKKYz��=�$v��g޴ob7WB�x�3��>���u�E��2��2\���oN�\�e��2�W�|��d�
ng��oШEp�.9�|�'���\��G��w	���-��V}��Ù��4O���Q��(�ueȝ�&��a�� �1���Xv�f����N:��]�#ꅹG�R��H-p�/vkz�Zjf��화"ְ[I��]�ΏKF�y���cD���XpwH<�Q�Hc.���ř��^����B�@�6�r.�������-�2G�����ǒ��f�ǀ$�����j�T���������?�fʲZ���(�=%��Y��ΩS{pPG�w��8�'o&EU�ߌ�1���5�t���W�xu}8|��; ��Y>�>09�� #��Rrrvn ��qL�>H��dM��K{=n��jX�!y��C��W�DtՆ`8(���(N6�6X����͒h��&T��I㽞9���޺3�2�V�[.ӌ -Rֈ6���w��g����(���d�3V�8^�����'�A���݌LgE��*%&C�<3��Jݣ ���6�����PƄ�_���7���c�P�tL�q=�J�44��}7?�0}��:q��~C��P?�hr���2G���G�$;�&�ͺZ�*�pC��ez(�l�H��v�T�e��s�wh{B�*u55�+�m{��x���4�/o�h�۪��+��F��R��㇐��ȫ�HGa���(����g(�6������b��y�}����/�]��]YZi�ӥʞ�UI���lѲ��:i�7�N�x+RM���SR�tAl���~秢��-a-�M8v�mq���L�I:�jC����n���KF��A�L&�P��_�+�4X�qs�T��3�o�[L�$�j�]cs���R��2��}|��x��0Iʒ%��\�]]{�U���J��.�+}1��I�;��lPĴ��g{��>t����~�Œ��!Uj�0�~)�]xm&Q���7K����N��Qf������ʚ��`���J��Ț����q�X�����:M���jk˼	N�d�qo�����a�՛�Va@��?q������&�]Y�`��}�Q"?s�J���|.�ќ�ݩ���^K��J���.�uu�XË��2����4�\ a}]D��5LKMB�Ώ%#�O��x!�{�}����ET՝:Jמ㺮nr�"�xMU��1��8����k.��n��&>�Ǧ��u���ݺ¨P�uM��>T���퐆�6V��u�ܢ!��a������	��+1��w#�st?M0z�S��ݒ�/�$A�r�1������P�[{O���s!K�O�h������$Ƌ�|v S=8��N�ws����������wl���z�1�4�r�k/�8W>�ƚ�ž���:��l�5��x��l�d���8�7��'�v뱭�-���M�nn$'1]��X���p�ԙ�a��7�{A���f)ivQ�4���-��M*�����4��#�ݿ�4V���l�b��E��r�	����-��L4S6�#'n��R�e̢?�t�v_.f�F���p�{׀�����, ���$�0��r�Uy4���P�ė�y/t�^��� ��)nձN^����L,�C&� �{�e�����޹d�	�.]=z�яh�Hmr�=�t�yF<CH����Q�_rv�|8g`t�����U�����,�X��̈́�����R3�<�{ە�.�,�3�1^s�~D�ز9�|xC���lr��P�j���",ס*-"r8���eio�M[�n�T_���D�򧎷��0�>̳�mJ���&���#�I ~�E�~q��W��Oա0>6Dߘm�^��EW�R3񡓵g��3���>��:���Р�-���4g�8���{aK�Fk�����=���W �H<��]���*%V�]Y��:����_����7�_,uq R���E��@VS��e�}2�O�J#P�&�x����:+�fO�;�K��6���R�8���x�1�O	�A`8�Qc͗؅dCR�!{]�S%<�n������}�]u�%fJ��:���fx��4F�d��x���򍠓�W2�.�J-�g4�"�-������U(q�ɻ�B��:�i�m������+�����~H�`P��Ug ?�Dm��3C���	��\�|9��X�:���a�ߨ�gy.f���%��jr#Q�`�$� y�B��Tcx3P�dnr,�;�@��Χ�Q�A�����mc!����	��b�߻�w���}��B�6�9��?2t$.�w����{3����t�,#��V�_�^a�o�icA_�
�b�+��ҝ<�$���h~D���ۓDbdCpT!�Ĩ��7�{xx���%4>�M4�E`�S{N��O�����F>����h�7����ת��0;���D:Jj<�s$&ʵX�t�b���3Ta�����?:C}-z.�q��Փ�i�Z�G���R����,T�UN�-�E�����1M��C����<���-�r�ȩ1��lVL�����Por����.
�XWx�(�����J�E�6v9��$or��o�J��(1�Z���4�o�g�٬�p�]����:�}Qǋ& �{0^F��i;h��g����99z<<Z�dqZ$1��s��hG^vy�F���m<�M���x�~��X7G�X}Q�������E�W���6G�D�}���W��?��y�H]�W�)ކo��E��'�-ݱe���n6;=�>ݻ+*��gn-saj�o�]��p�{���{�����M-_3��cnW-GZ'o�;ΛBTrd�h�T�t�{�s�P�J�{���|$ω{��~ۦiZ�T���\��c��P:	���GQf+Ű���K�L�d+`��n�ڛ��=eK�8Mw��r]o�Z@�M��Un��QsKP�W���ge��Z/9b�H~�օC�!%�S~�uC���[e=>6��w%U"�V�L*���;��ɢ�y�eA@{�.�>&D·zUP�&��]��>��# �wi���Xw�\	Z�߃�O/�Y9/"7���H ��xq�h{�&�3X���.?���M����P�&5��