// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:30 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ogf7IszXTek2mcStBmPuqDGGKPO8hr4d++G3MlRTeRhuTnBKAZiTOyiqr8W8099e
+mENIBWcBWvj/qPEZHVhOK1csmFQ9PUALWKEM7bDi8MV6ra8bogMGbnODAw/K8aN
cyK4oBCG5uzK6kmXzl5hXcAuDtUEbdGJwKCQJqT5lYU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5248)
SOhQ1doLxWtgaFz0h50m02vLhxGG0eUYezktT5zpJnumE+kB4Tl6QvS9GUJ6plyJ
KTnmm3NYGNBa5Cx98fPs2FVKYO6hI8R5UiynnfoMPlpBRCzXRZ5SEuWoxzercjzM
YufIRViJXdPwYyK0WkpwCxsV8qd2bt1up86PjwL9Aoyrjy4sqxZaZEXQfllyka3p
TF8k59NC/XC+Vu951roLaXykatsI/mPTV42J3DsVKpbXzSHJsn23E46HVgF7PPJM
qK+C/XsY7yFOYE4tfrjRjYMJA8BS55EgZhZqEOU22dGVfkLfE43vYWJrkpKTfUm1
7wu+rf8yv18JwHtp8cWvfemuq8E5RjPwVtDoZkMTSeI8f21WPl4k2gvIj708yBzl
D1OEKTDOmQ2E1Tgmvg7BiWneJJxHi8aRYe7xfh+tZ1yLG8UXV30ga/luPkK4VYn+
CWhjcViWjdSi1Uv8Z9iSsIZDjNLlDCcVG4bnGvTTLXbHrjIPl0y2dFqUE60YHhu4
hlWzwJjtXuCbScey3S+/h0sH4UNR8DbBmuT1WdbUEytcnQzTa4sgMvcLFhAUJZgR
y73eXglMxOOjRRJ/YYAZDtIV8MHKuLBy3ze6Qnygh4+iOPitVceXP0n6zED5jq53
bKa8dsaIl0AsOYh2QfSU2b5HegDtbbNL29BQp6zwgbfZczbkosu/BGwcrVms9C/w
5mNPIS1QNf+TF16EECdaQGma2XfcnX8n1VhPCGlq32kasOITbNN1ul3/zKLEHZEn
hJi2EgzIAmWcB5sZlg8dbYGuxCZYexnRv+aH42fedB5FSODUXvNPSYqf82CCPAJ6
IwLh7tAjzLgCnJRlZmW2e7Z7tDl+PBiibs7uSxtzNqjvX+rVGraSPRSJ6NBdyckB
jj/eGo2R7f/vK+pO3EF8F1LU5phEyhyMJui/urXxV7/qMdWq7CSzMigIq9QW5tNQ
80K5X31kAiX46nLPdWlMMBXPma+c0dnDzWVsfWngk2dQO9eWMZ8e5TSzyOxgLxTo
jZonL/brTTKE1/GRN6R3aEZeiHbBjj89dVFjkx+URwyyKRCNvg0cvwKmlGUg17ln
0KQhnzOmP0MCE16eLCR38Pi7DonGgcyQ5yzHLHicqJUS5UIo/CrFR4TsA6izMbZ8
+puUuiAdGgbK7pgM88u05JW98B6coa0c1tsczcwwhcF9xgrP4zJdRtDJOB7Lv+tL
o+9lukPJA8xvT6ao88QIUvoP8Hgxh8tTnm2Nvk0B/11iPVFhzgUE7yi7Wpm8sgBn
GaR6+p43d8te49KF8s57KwSx2xK+Q5MVO6mje5n61t0HirQW/0Vvmz/yRijLvTOB
pHk+SDbR7pJDVobogYuF21M3tL1XHn8g1Xngx0ElNGMds0XiYqZV8TjKk+QWb+xM
g9IPTa7Ac6Di7h9HaHSSiXzgDHOD9aBmeZG+VLTO8+f0XzkrXmGnN+/+LR3eHIYd
/Fm+D/SJBiVrSTPrGHoJKNPZBwnDIV5ROg3vv+1shs8y4OSB858ce36JdOTC+WsW
Wa41rNwS9gm2AUbFs4L/I0bc/AzddAtONCMaGwaOtSIgY1ub+d20Ql5YpqECLZrE
vCJF+ms7xRRHtyAGPLZlscvWWrHCa3KfB+0fYn6rm++qc+ASTmOEDjtM1sZHX2VZ
csovL0Vk6Wn88f8/+lEa00RLjEb9XW5dwM6ruf52YxJwBu4oFEBCiVXGS4RIimi5
xe9crOhAsgD4qnh8fjaOK/92EACykFzXMkLbN0wS3Lum98bajvgT+DOKfMjm6nQP
v/rOHf706PHZfopj4ZIIe5h8xLvudesdIidGZGdDWaFQOqBlA0/mfySyUSXThWeo
4FyX9QqYjTz94OpwEaqlfF8TN+sEiYV3vWbqGJ52Qd25yeY5NapgnY1qR6wUJaC3
yVaKX6FRGZIF6StZx1CeZ54lpPgu/yugjG12s50aoXieHYfW/NDCxpOEih5xN4Du
+cIBhMtPGznSzBX+bSVRQaOFv2wDch6AmbkDlrf15+C8eZvg30ZBHNrgp8bNtML3
f73WUDGKo0Kh/IbCiwo901fMDiiNMK5OBiikW+i5hJUVxgYCGvn9HWqpsUogIgNL
0OqnfUfP1bYA9OgYQtxw36Noa34YCbPFdm4c3jsbfGOliFW6+cfsGcx6b2LYqN68
ems14u+FtD1BRVL+FZ61mGJl3Pe9aJzPHpz8BHSqjjXvzc2Sma6BTOC9XrGNpLby
/1WjA5LGfYK+3Q+gEzhpMQNlb8zDRa5+C+ve023LB6rPbSkjZ85z3+yooTCIjTry
rIZer8ZoNi+PdB1zuQs486xFho9gYvRd7FGA4dCeiki2JIWGL0Cp/3bNcCKeke53
dD9GCcigIysTTAo7kJuQ+o4L3arKUe0bcr7HQ9u4XFj3U4/r6UDwmrpqZU9T1lMs
+Sd3Wxjs3FJNMH4En+iIxUZYrqg7pYsTQWqL0DmKLpS3cb9v8UffRHidnSkpfkmu
IM3OZYcvBLJI9KyCpfSon+jP+nr4kJTK01/A+bvikIxJlfrwNGqk7ILvBvHIVYPp
nUKLBQXtthpJvlxy2viBFBZ6WE2nBZ0oBkeXymMLt7hD+6BJIpJo4jyoDNOFyQNn
ibLBVJd6QgXI7jE51xE+zKgLPicLHWU2IJi6fTqRmqV3w5y7JmWvsV45+rPPYjlh
6H0eqJ2zifrxyqYPZ+Zuhlg2BrZFPm+cTElCiTiT5jcwblka13vV9h+40Io72ncq
dR4LeFRMCQnwDTrfqLJmuKh6O6efe3QhL7MZOYVngC6MmT4IC/ruGv5X0VAZopiY
Lvuvp6fRDoHoKJvnOeyeQCjvKCE3yAoM1vR9CZJZPZogaAm1EPYpF1LE59J8qMDg
4SJOy8VQmI/t8a5YkKHyrysnqAZFhf3cacMbfVPMFxYVzAJGjDgsyqNVXLEowF1b
eTJIbqELLUyX46owfVqXFagsHQ203SqZf1ph7XYC0+d60OwU/qSqtJXJKw10LVI7
ckGG74gaHUdDY7WG9KyPuMIpSdBO0GE2FoE41U93mzr+a6alFTWSzq/+4N6aTmCg
5YniTJ8wJ9qIVN7PlrWlB/Bgxfy33ku4SWUsOC0lShp6TyhT8WFG3idk2KvTrw4Y
iWDfyzprXwr4UdMhO7pVrzxtRdEd8v/uTqxwPgXDkwO3MWjKfEsgc7djEckusGPB
7L4C62af/xg88Hv0YNwvH0EXGQZhMFG8yKApUAMkcvFnMyKBOMlYsjh0TEJEenoY
2nfodQFF7dILCgviZFgFOA/WUnxWOmY1nTe3ktbqkP4wxvcHKG/vC5eCJ7uPZf93
aldabU1FehgtosnyPakGFAtRqk+opdJWmjWM8W/kse8887H1Z/10Ca6mKr8VR/oM
kOkSB8OvGcTuihRF/GUIoeodd4HjJ2MR9qDRbssgj/xIYKcJ0t4aLMeWJw6DBGo+
3uHUTdMJMbIWcIBdqAbJU59NO8ksWBlNO2h17uCUJHlZFl+uN/K1e2WeDxtr7qnb
TjCZPPBjk5EM9W+U4QDs9egy6dzllMVj7WksTH6ZqqnnVu/f0T1A0BqgMjW9aNpK
+uW49UkZ3bTqgFgALmcuBXusu7vJYuT79QM1DsFS/6D/TK19ubKv/VIDPayR5Z6z
NI+GFuQweCjgj4O5OQPT4V9uhqZw+drxww3FJeVV9bJ0/0+XfRwZSxuQPHmi3OJm
buox8TXAHj5WGibZBjbiXjBTppx6kof7UkWeFyBbgoJDT7loRv4sELAHcH2I0The
kgl88jb9Bivcld3jC7ASKFzst5ZpSALBuIqfnKChx+Bg0DQDkYD/BAQNbL93FLJx
pqnEb9cIqiCyN4EHODjUShp3/J6DnVIwKJmttroMcf0o2UTQqeJyYvBSmqh99C+2
pI5w9QNWEaygobKaWOjEQJgvEYLRFnclZ28loV5qMJLf0+DI/HG5Gi5ERr41jqEz
tvvBEGUeQiR2KZX5X897xIbtcpo1r/y5honstRwIam16KERPCxA3io66Zg5xW5k+
V0IxEDAVDACpgKdau34QcJAH5m2D3CmKeKJr+XQ+LKFaMrfBy9mO2vP+y/889yAB
ZJH5G4WgBtvYVdfXqh6dWmXvh8y17JYaPci3uoFScszsNDL1Pn8g0NVEaers8aY3
cwOrnL7LN+jUW6JHGWCscwznt7xwDr2YtVYTGz8Wk9JvNQg1Y7Sfr51LCkP6e0Lt
HDMe57M/y74eoVt/rBO0UxDACVG2UZJcuxGq2auU+Xh9HM56Bxj5XbXRSASDKZQ0
tOqdbw8SWEdQLGQTjTZfnjOT2TT/72HeWvYnHWI+z350lp5Nm84X+9flvcIEmkyZ
W0aNb/xMf/waAxoODomxPoWqmpl1a64PGKKnoAA5CnuLxXCVEOEqBc6eAw2oG7MQ
VJ9d/5Cx1Nr/ILzuiUwPdn33TvVVcGBmyQiZ90HcZn+6XI/KLM5H7ZzwxvX3Pnb0
6eyi8qW6F3mEjvFB/qfAEw9M9YIz8WdE7DQW3y2XrsAmEtFTlUbap9OUV8iTIDgA
BRMbDFB2vgayAA+R3Aw7fPrSdytGecHYYO6LWSbKXN3r7NW6dgDa3L/voW+LwuLM
PNkh3Zo3mInnAYDuEboNoRBpTxvt5i0xuQ4IrhWr9KDOzEcMHg//hBCf8hH+mf+S
JpdjZFm1IJZo7OYX/u0BJzaCflzMZIIUeve4m2+LlG6KeMKy8aeJOokoQozjDfvm
FQxLkWVIrPhxuG5E1rtltY1Yl4I+Dn3H+qpLS5vMzZi8vniCX7ybwqL4Lj0DCzju
xD8Xmp0GgGb3NtDslQ97ThrFY7fbWsRo5Zy02ViVHdL+liuw/4zJdRtY/LxXeL5B
+VqI58DT8sHYKW5h1WN0ieIV/l2B6+fUKdsIMP1lFl+hmBBTba6sNMNpnF/cXKY9
vATe+4R/loQmFqbQbUhV1/MHjuXO75L4q/kgURXboIZDOIct1fyA1vWZ3eQoeO3t
PehBe9qRhnYvaTOMcTDJ05WyRHQiJk32jzoRltsyBlk2MikHIzrihqLLukrDcdtw
42YfVAbtd/WtJtv/f/tjTck7QZJXWFIQbqNNS9vVAPBtayryNUL7AEK+pZMoI7X7
6g9FY04rh5ytmp/FPaomngTUIqtKPkyB9irrx8eNSBElIQ0SIEW/APr8YlwFafRC
WGcyBV8uy0GEHVyhXbb0xld29xOnBDozsJFbG9JBqEpz3i+21wwQ7T56uvHrNvL3
MgPJ6vlwHuwCqLsduaVdMG90sHiDY2jr13SCUlJOtiRtaeB6Tm5iuTZ8gOLhbp4L
gyxY0cbulUGscvHNCrUEEz6F2ba1nAxNUdL791BFJQO7/HhyalRZr7LAsCRCC63E
wLLLLnXuyAJ5cUwss7Lc7XWzJax8Sxj2j1uZT+IVaSc6X2UzzEjJhk9wr5BpcSe5
miL54sgDLcKydcmgfZe5wJ8Eg5sJhXnRZyvVPwAVyPteEFfWWwDnRionpEh4Y4QI
2wKjsJHrrcD78tBVpKiYwVZTj1HhhWTi537yK+OfoYdW44QAGJx+Sl3acKrfDRWV
LFxnQM+45lxIkTplyfXYg5KtXSGHGamZS0WXee1sflNbRseq+CtRAcV5lZje++Xj
skVxhSLObk4WqMnzs319iJ9guJ0utxjrx6ezKHvLM9hkBQ05GNC1zP3BiZMnK8Lq
EYkAbGPkKKRqFPMPhNuK7pioEuJmV3OL4cJRk7Vu7Pm8f2sH4A1+ZNwEh0YYe8Gn
B1fVGItkivAZyJl7j00P3ck9yZTb8fos01Hfnu4vVfne3tzBllVUY171E28raNhb
6CbkupCJ9MV4/CC0iW4Ta8VO1zVYMRVnichQBSCoxWK7uDk02jd3oLhC64vqh9Yr
WbFDnL1v0zhMM4Tv4EB+SbUyGjZaUCS/aL2vzSjAo6TWV5DJ9sndgAfwZwjdiyJh
xP0tzEW9x3Qk0P9D+miQdOCXiz/2U9Av6lHws7DtrNci6IOznRlV5ZkkYTmMcIez
5pZ9y19fb3yonK2/nls7xfMwVQ5y79LxNnKSzaIPrPIJdzvXYy2UJXN214Tf9CUP
+80cF4vo1YuHCTeJBlLD2wBg9SmdRdzNe6HOo9trp/3frcvNX88DZ4UAFxeZc72c
wdsdV/XF7Fg/W1LDJwrIZQJ9qJ7u7vDWCEMid0qPnX0VWfqQzbZLITa3eErrq3uj
0qsNFZcDWnAGjQnCGcgrcVpmUh5D0Gvj2I1wYth0MPqCpLsEGgjwG5W6A7k9JsRo
vw2UGLoBp7LBcFFQaQZ6ZtkQexUbQh1LQyJNjABzHraKJHb4cvoPApvASG6yQLbG
tMgZOyxvPy7AFeoOUrQiNQnoaoQCnEdKtIsNVSurbg14r9NSVS6IPqHueZop2pb2
sjLy3oz/cnD4jEvDAg3Kg6w0AIE96RcUsWvS8vVBWJmUpd7c+BHxO3XqtCgOEZP8
IkwWqyIgARRXxB/KjrcmLYkIPg3xOtD8v+mVBVtufdwLhEdw+Yu4qNfRj5RZSC2C
ejVMPxDEXDDXoTlDx9lt6XpGSpOvoAyTjKK8Q4V3QhtGajZ2YnSGCeye70xfv2y6
UbI7jtRHDoO/RiR3pLQ+2aoFJ1+EGzWhDowY6oaDduEgwM+o3HRIKGqz0CspK8AU
l0WYbI2QLwAL6dql3ucpEYVCxTXi7xigkyIEx48DWhp1G/jsELhjN0VUTk9zSzST
oOwVVYqIQ3PTURurWcnVBYc+FEklMu78HEZZgC4SpNZ6qbx3qa8b6KLK/A6k4ZsW
q2LQFdwOTKpLw1iOpeZMkeTv8Tom1msk9GI/3dx6YmbN3Lc9X7xRNFX4EPZNaKXH
mhRCUMUMMSswbRdBg2S8kMQ8sqI+1OmQrja3M2QFquubfrrk7h7rCASVbrme6iqs
VJeiRy5PoEMTOpycShOO+0tIafe4Z9AI4c+702r5ORP1ihawQzO5Sz2VJKruaNRr
iP3pNZpbnX4jazIweHZzkw==
`pragma protect end_protected
