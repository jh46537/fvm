��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<����d3��i��:��@:$���;��U��zV>���=c��Pz�zaz�pwU�8��CiA��d1����T�
-7?�.Q=/9��[�k��E����kax[O�}�&���\k%~����DԮ�A��8;ݎ�����\q�}�q�(�dP�u��.9L7��}�x �p�������1^��,�*����r;�^�%&��Ӑ���T�t�B�ۤi��
��\X����M�H�r������ד`AG��ޓ�o�W��)x$�a��rM�Q���p1���#�,��r�Mg�
��G���?�O��f��9SH���1�KHbbpg��c�� ��?�A������p�b��pE�X��%���I	Fz(�sX����3e>g'��Xl��I�Hn��d�N��|x������[���e�(cܝȰ����עʧR^k&�;��9�����`�HTۋ��0��jjL#������[��ɥx��3�T��G�4�e���US�D��q���AC@�]B-���v���x���bE�~�/����p�_�*�%V iJ�[�s�?���!͹Y,��@\�6�Y��w �[���9׹¼/}6y�@<�v!��T�ӷ�=*Xbf�����^(�1�Ä��"�3��3ϸ�N%�릢�{��S~t��q�q�/d$�:f��z��IA��}��a8����֥O&�h�����3¿ܪ��^��w�2ܛ�ɼ�uA��6;)�#�(���xI��xrH�.Ʉ���.��y��{L�2+��7�T��F~k`/�J۟�������v�{Y���+V�)Tv.HhJ=�9����t�
")ج@�%�$�ɏ�c�)��dZQ>@�t��4��[�K�� 4�55������0��N��r������=�gDk��X���ס�M�o�&J�Ϯ׺���nj0�Y���ڑ��S�xM�T�N鸡8Ôp��|d�>��5�(b���զ�y�қ���~ω�^>�4�$9x��K���n�����\SWJ_�n�!��`u�G�f�a�!�����ǩ��̖d�!c�`5�M�^۝�4�U����Q!F��f�R�6a��#��Ցݨc���B��e����:�_��+=?�F>TqVA������զӍ7���.(Ώ�r�z��<��;�ҝ�vc��Y���݈��'�����������ぷ9|~�H��隹8;�b`���{�J�y����l� a�!4���h�M�2ms@FңK���j�����t��=��HV"f+�񻏨�ӻ<�)*��Arx�����Ϙ\4�����א��5�yRJ�����;�fQ�gq��o��䛰c�$� C��Rr?�P��7�"�n��,����H.=�ə�;zc��0؅�1���쫻�#�p����je6s�o�)�݋���&���g��᫂��:�W����&������Y�V":����5�	^,ω_9�fV�#���e9�Nr��@Y�ժ�w8y�{��%u_K����π��m�9��V-Clg�`�<1BR\���'q�ט�L��H[HY��=����l[9������R���H�:�i53F.�u�R5���Z7]@�2´��-�/��0�V���%.��I�@]Z5�F�Y�s6��D7E����Y4 G�������N3���ǵ��/��6��t�d`��SH3�"艫v�p�as��+��4{�����I�H6�-�3{���,v{�SΏ���+��L^J��\�}�w&,lE�8zh���瀴���\���b�n�,�XPAN~��t�Iw(�Ť%���O��D�{s���J`U�����ī3�L=��2���u7�M��<��r0#��]!���m�5�����~4�ws�3�1�6��`��̭W��i^=Uhc�����ݻ_@�Y٘�6��Hh�o�����\	��L!�l�5ޏ��$��H~�QqQ���M�[��#�xO������*�'�<��*��؄�KM���_��"���D� otZ�O��x<�VO���CT:ܷ��YJA0$Z�ͭ3����l�oe��/71+��-�ŏu��m��,�8�9�����jdԽ�-�h9�4j��ϡ�q}vw�,	)���3�#j��]��%ǫ(Ԑc��.v�5]vDg��r5�gg�h�!��X2�U��p�M���W���'?D��!���z6Cr�IB
��5�(��X�!X����Bt�k�� DV�P7g�v.��H&r4Zc�,�9Ӑ�>��5t�>�,�#�k|�܄8zo�c#�|���X	c`#CSY%\5�W���SU�N�*0P��9ҭRS��-�4*���#�}N%+qH]U]Cύ �BEf�,#<:�cF���M���Q�s
N+<�o/U'����t�E�3�6T��0A9�~���0b	.�U���x-%&�muY�+|���q8�gDW;�5�o�dEY�[�%B���AS�?)Q� �?1�$�Sh0"직n�v�x�q��b�Yv��FN��Ī�\Vk��Cօ�7L�P@H�KĘ�@w���‰[r/�*p�xqhA$p�z9d���] �aف-���@+������4�[�n�3��q���=�s�,�k���l�@�q�_FΧ=*=����P
�Wz�r�b��.I�:3� ���z�İH^f�A��i����d����Nĸ�\���n]���b��˦)�%B�M��z,5�'���3�^*��h�g��S�Ȗ�Ŏ?� H����%Оz��X,<F����2^Y���-gMEWc|��dR������F�Cs7@K��e�L�%�It����t�]} ��LK6;�/8��جud\���%�sDP�M�к�����I��D���0�?��D5�~k;�%p���d��0ٮ�>�Hx����v�.2�+}��]u5�-|[v�ǲϕ6�A'bg�1&r��q,��g��gN�}1ܓ@����r����Ǧ�9�"�~��fU���>�	�8<p�/S�Yu&�H�����Pr�^(!!%�U͈_2�Dn�I�0�[�W���hХgT�f�Atl��Rvm��
	濇�%�����Xt���V�JV7�b�\]�n����Ux�Ѐ=��HZF,P����8wuŰk_n�?:�&8ƫc{TrV�Gw�@��y����l�i�C�=o��S���_ٱ�Zx*`c�>}O�Mճ��tt]��+��+���*N����&�}H=���.+��sG/�b�-����$�j��m�b��@{�mF���x��T�v�)G� Bo'��W����{c
DKʞ��R��m�	�BR�`G�4�3��Y���'as�,C�(Xu	���Zh0R)V);��ՖrH]�*��T������+�*�ז����k�Rv]R�����d�V������.x����ԡ�j�,����qL�앃K͝7��֚����_�'��̸�.�6��r�i���^�87���ճ*p�?h�)m�4{��`o�F�]�e�+�}�:�m-}}͉:9 U�����:�5��r�آ$mq������8��J��|� �^i �����)n����&h��V���1Ǘ>�n��J]g����D{q��ly3�
Gi�i;̏�&I*n��x"�b�H�ڲe�}.����stO�[���R4�o���0z.��~U��+�9�A�c������_^�J�C}�b]mgD�L?&(��0�q�8k���F�7����F��@��2*�`b�i����K�e5��ݐ���DH���}>�gUg�=�)ݜ�u�B�w���D�2�S�1%$��Sk	"|���w��뇙����g�>o� �US:�R���YAqXU�s�i�ʻ*�K�0�Ih�CBI?C���A�`�j$�5¿<[��,�^'|�?��:�dusN���t�dN#3���_�يC,q� {���WvB�,puy�g�H���j��Ԍop�����cU$ Ǵyi�Es�4�+�Og�=(�=�g�e���uÉAx�M,�s˧r?0&�;>;^]a�ɗv4������\j2�:s&��;&���>�q/��S�a8[t��ku% ��;���$���`2ַ儂�
�W�G{S�4i�Q���k�(A"q�]��'BS��9I�ǔ�6}�Vwo�4�!A��;e�fa��y��h�ttN�j*k���(�f˜�H�(���T�9Z*��^j�Ș�=�G�	�)�0B�͠Lֿ��΃֕�@�o�������T{����[�/���#u�ܐF�Ểx�k`��!eӕ�c�(����Rҹf!�,��+�,<tQ��8bz�t�����:%:�U��٩�(�#�[Cpn��r$�
U�!���D	,4� ���M�5���p��  �x��,�s3�K�@�KxF�%����Q�.� P�NRCD$��Ī�ev�w�f`g̵����8�y_�z��N��7C�x�AL#v�x,ץFݙ��L�)q����+� =x]�6|����[���4`�����/�^}�.˥]�5r��@�D�"�_%j��g�]�
��Syp�f���e�tW�l�K�F��H�/׷�Y�Z5�-�w6�.�=�%,QĀ�=b ���.�"��x�N�ݺs1��ON��x�&�Ӌ��\����I�5�23� ����^Xf��)*�� ����
�I��/�j{�PS4h'��Ō�ܺyJ��W����I+�s���g����d��nT|�W&!�>��z&���ke֩_�+Ǉ�]�o���5�ې���b��R���?�[�֑	��2]}#��z)�'���j؁���p�"����;[5���ׄiܻ�7=|w�.����P=/Po-��fe((���n�W��*/��8�iᅮ�[��4��iJ��5�)�1�^��VU j�g��L����.�*�IHǇ�����r�$�d��2��~��u�A@���29]h�q�߀\i��#�~>dX�%O����f&Y�P��{;L;7�wof��q�9�*װ�Խ�=��׳AL�����W����
�;�(@v�o�<�0|�>e�O�Y�7��M��VBg�Af��(���hbi��Ek�E��W�����K���2+0�=i�%3ׁȀآŐ�%d�)�ڦ* ���_�ˊGF�ܤx����=&��w��e/T�q�Ux��������)��-�2JA�M�p��3����g�$}�q�؛�T>�yܦ,�1���`��tEF����h�yC���6)��?�j0��2��E�P��q�q3�W�r�(�=�\eg/>я ���3�II2�d��|�ˮ?�M=[�< �$/���#1ҏǫ!��=��H�2�q��4<�3����jH�D�Q�ȞtB+Y�G�[�3��ZA���v:�v�
�n����(�p����	9�a�"�u�]��Ȑ��M�m�OR����A��������
Y�]=A9P��8���U�s��1�4�r9��������%�#8�0d�� �L]�_׼/U	W%��K�(*�X�%{hPB\_l��}��D�	���@a/J�$M.L�����˰2�(�8�����ܞ��	pO��Dސ��K6)2�w~��\L{�17� &����Z���w���0���qjh�"r+E���+M��
 ���i�z�,Q0�l��N�2
gL>�l'p���,=��Ƕm%��칀0�[����ګ\#�ު�Μ����)�����}0N��1Q�M�>M1��Q�[wj��Fd2ܗ�hH!P"�.�hNm�bz���A>�B�>ܐ�n�O޳I'�@�'oD��� Qj���D���DD/�����}��G�-�=��	{��:�I�#��z��3�����r��π�l%���eԩ𒾡��%�jRU����������/ٶޚE�ߖN���Ahm%�3���]����o;b�n�Lp��������a�|Tt�gw�C4������| Yv1��_wy��|��2�Ơ�����nI/�
���ԙ�K������M��EIƃq��K��JW�NCD��}/)iW|x�Gz��;R�Vۺ`�+0g���4���ZP����v'x�G��ZK��=�;�~sA"��ҀQh�:�ɑ����W���M/�p�����r���4�x�����"�X���T>l�38����?�+W]wA��N�'Ii�$�Qؔ����q�P�k`Q�:�Um�����8���5��}8bt�j�S�Ͻ� v�n�=�L�:E�h.w���Z�.��˶�������#����<�8ʀ�Ǚ�s�{:p�5�b���8Jf�xy�`��d��}�
�*6�Q���.|��e�5�%��x�)nk9��b���F�E����=T��Zw1��,�Z�erv�+
Zh�n��D����$�
	#io�U����%�͆��D*OsI�B�`�B#�{�����7.Cs}kb��ef���N�e�1O?��r(&ZK/X��,���8�1�P=o~#>��;S�Z��̞������zq!W��>'՗�b����Sa�-h���8�y>��u�TێOQ#7�*'�1w>Z�ݲ"��u�k�6����N�x��n��;'�lF���<D�o�� ����Ol)��v��&�]�G���E�u��`xP���(cAK�8R�K�3��Ҋ-��A�Oe����)�ղx�G��(#{������j�ܧ#>�7Tqhߩe��La����UK�v���j�K
��q����砃.��|�.t�sLެ2����Kg�,*>4����_�]-.�3w�\��f�f`}7}�����bmU���J9�R�T�K)��;���W���.d�f1��\u�D� q�~��q��N���n�?�!�'��6B�FTp�xl���z�	媨6��sR���LC������x3�g��B��_���{��f|qwa/T.΁�j�{������:��$����@@�*�909���W���&��n���-s�@U��/�}kbÔWI0}�:�M4Y��^~�?g�})�G<�P&���\����C���Z��<�A�tJ�ŪL�9��jc�%�ʿ������Թ�$���r�*�q�|�$n���V�Np+N�)B�� %�L�6H�`�l,
�3��Ng|�k����-p���S2D�J|�"F��ٸ��b�=��VdsH*���>�>��TkǪ��ҙCfҚ�[�(���婖��E��R�Dd����xG�����7w��cb:*��+��-�_=�'F�l�[:�d� �
(�����}��\/�����a�4�b�Yw>_as��ӎ�e҂��h�ѰLª`�[,mL=���ˮ �mn�b�̛7M��J�
@"�]��[�z��j�`d�?�t��L���&2�/3*<���X<v�����:���@a����r���K�2����L^��q��bP�G
�qhbw��M��g�+�%vm��J���v'�2�H�w���!��S�pX�t�ho_����̿0Hk���ה�+�u��K!Y�N<��9O(7�����D���.X�;p
��l�h�q�6��ww�v"��7���^:���:n<�,���$+D.&-���ۑۋ�d?�{e���������sM+? r�����֜���w`�%�؟u��Ł���=�ٽ1� �P�h��[�}�R�À��SMK������7�x�=�9f/!�ay�xz(p��}H�]�ݸ�W[�]$R�I.4�q��b��]&��Gi��:�����${���Ȇ���L���Y��/����"�Ǆ��q�27�m��M��Q[�m�������