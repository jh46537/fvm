��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�����:��=3�J�r	=�� M@Q �:���!+��?kC6U�T/���&��	�bK����V��D�Db������V��yfʀIG�D�Cs㠆�.�`OI"��\��L'1dA_���%��:��c���'P���G��4BS�_VW�#�6����ZT�v�O�! Q1�fX�<o��3���x4��̢�!i}���IZ���C} ���ӣ��L�l�,��Z���#)GO2��ׁ0 ���_y��7�����m��n��tGo$�=x:�U���������3�YX�"}�ۋF1�0� �-3��{^Yt_-����W1�>_��M�-�����������&9�^�?�ʄ�BϦ�s�V�gW��ĉ�Y@B��9`wg������t�I���Y�<���A�T�L�Z5p�C3Y���D��N<�;�n6��y��S�s�ok����h[��������A�{ZΜ�_6�^��l�T0�`:�SUbD�o�u�,T|�,�|���hD؂9r�����ou{����>�G����5Υi�p#�^<
?F����ȕD�`��	]f��B�r{9��wOM��=v�ٴHt�.`}&E���x��Q����en�f����=3�"�^p_[����B��&#����l_<:/l3��H 8�}$�vq
�_�� ���h����f�8ɰ�� f���c:�=�a!�LAŦ���<�`�C�4��t����?r���52K�؜2�o�>��}v�.ER��v-�?UmS�)Yu�t�e;�F�]|���H���:)�> ��WCqu��˵8������.}+V�>���-kΩb�����_�c`� :h���*�WFBk<{��&�)/}�����	���Pu�Ր[����e��tD�/�2?��e��h� ���ޅn�V�2��-��vM���P������P�p����wg`��2*�(f����5c[������<w�˵n`~
l>d�� ����=���d��T�����T"��#H�w��f_,��#�69�ھ���B��R���17��)�u��,4���Ɏ����s�©��J�7�IU�8���~���?� �����u�½���+�@"	>�6�� D�G�4���2|j�V&5O�+>%���m<�}�]��vƓ�f$=���F�m�H.��V�Ze2|%�e�7�F������"�*4�;���0�?�S�+j��#���(;��H
TwDD ��/��<u>�n�@��� �����~�g���O�&�a���g���gb�=�Ͷ�T_�\�.�Hc3�gE`�$.h��F�7��:GaOw�����z|n3/��M턞�	x�HID��8�ٸ�H�{�d]H?�I�x��,"��a��MQ
ɷ�8�@{C���S�9-��.�,�Kn�)ll�&Q@e�:��e���+��9�W)��9/i����P��%�q���D)����ľ�5�Sr�D`�U�b���~�U1� �gI�e��]���
i��Zw�|��ȑH�z��Uf���]�� b�ɰ=Y��gY�.1&L�ae�E)�خ�v�$���#��>���Pi^\=�5b�v1��{����Pa�y k0B�
���^��Q���%q]+���U���t��CR�0�G�YߒEvSp���Q<�Q);M/A����䗾��������t!�����#R9P� �ݻ��V�!檶 s�	�J���� 8��ە��zL��W�nt&n��ѻ���䣮 ̜Gy�̆�i��7OI�m
�]��A����,�7�j���pR�Wf��/��Ld]N��N��[[04Vp9eJ�4{���a�Lns��lqe����dBT���x�ĜϚ�Z ��7��z�����D&�w<��b����L?K����2�*���x�����L@M�1Or�Q�+PLI���d�&�.t6�������F��c��E'�`+s1>�_)���)���3
_~�L��N|����?�\O��l	����X����?w�~���M�\x�i(��wd�1|�K��)R�>�2����-�b�wEI�CF��8eI�Y-�r��(\��k����017�_x�����RF>8����vx��t5v��&�b�r������?���;��n��~���ޭZq�Q��Q6��3�\u���{-���v`.��{���l�V\���G�9	��Q��
$��xKBWXy<�)�D�YcY���#����5�<U��N�&J��R�QEZ��|$�a ��*�F��j��Q�����l\ճ|�a�U�7��d�/K�6lb��[�/��Ӡ]aJ��՗�a�"W��m{�z�b5k�#�y����z����<K-�����i�r{gˉ���޴�c"H�Gk�>�{�[v� �{e,��6��\�߂����
�c��&��B/ʫᐶ�� o}�,`�[�"��f Է����MrA��xs��U�j��?��u�����h���O�V3/����
5���d43�N�;VwB����Z3�l�$=մ�͔��q��p���ǶfK�������Mn����tٟO�W{� |*�۴-D�N)ג�B��J^��3�y-*�:��,8���,�
m�)���Ob}I�jB�Ō�^%�i �uC�?W%��bG0u�#��5cs{J�o�#r���K�g�q��0�c���,�ɐ�;��2Ȯ���yΏ�x:3���}�m�T�Ý9wcP����B���ٱu��0X�xf��������_x)�&:=K�"�, �d�ㅢ7ޑT"*@b�:���`�C�MS����ݔ�Z�a��X���|%�(2�)�����G�\B�e�5�C[T*j�CbJ�%+�?g����FT=1�R�6lx�B[�ٙ+`t��č�6g�*LWCN��jm�$Z�׭Waů�Pa���\�(^@���{�dJ-ju42��D�&���t"��Hc�&�'�f�I��}���%q�@>���TI���*@�y^���d�w��ߨ�Bi_���c,c�v���'�w'�H��ͅ�Q����]a��S�aѪ����Ja�eU�Q���p'���'R�����1|^b̚+(�7j4˝��ܕ-��:���t���n]K�������)ۅCՖ�H@6��g|x�ǽkj׍Ƚ �>�.S�ds��0|�^h���7J������!Zv�٦*���v�bK��F K�Oz�ys�z)�A�%����i��L�1をSBNѠ�ƁB,�9x\��%O�ԇ\��� U�8�C����u�歱~ra��!�nwW�W(�9�!�фϼ���Pc��"�Cl�]�0�9���u}S7�1�-�46!t�=��a��s�,��ᕇAn]!2`9��d-p�t�ʚ�@[[
��ch�� �dp�,�oD%d
�r᎛:YNI_]�\�	�NF.!�5���F�!ך$6oFIۺ _4���7Gȗ�@ph�l��xێC'�K��Q5ur1�V�~T&�,�I:�??���u�"�)@L �0Wml�/D��!f'��
!��HQ�<}�  {3 d���P�7�ݼ��2��Z����m$Pn��\�l�Gk�����k�ˤ����12|����̦�����^ю\������6���>`�K��>j���B4�Y�'iG�/PSee�a�N�]C�t�MD��|၍Q��3��)����GxE$�ِ΢}��")����v�v���%U�|4��d�ի�����H�K��!�<ޣ��0� �&�ޏ�䍧7��:�+���Km�:�3m���\2���4#�u̒��.���d�7�&����H��+KP�FsW��B�z�;��k������(��06cn��Mғ,M���j`Fwy���:w�Ch�QU��M��t���
�8�E�-��~]X�+�1d�`l�&�l��2�a�h��G(�M�e�'a��`.%lH֧��E�Zl��"	��-���P�Ա�>N��X��L����}�a�\I� (ZI�6.��T�
��t(ϥuz� ��o�`��W{v>t�X�1*c�G,_V9���l-��j�e��
~�$f�ܦ"|�&�S�V;o��yۙ<����"?�%>�ő��^�H��2�a�6���{�aб�3�L-0+ e��GO�t�$d�OU��H3��Zw��S�������C$o�/<E�m*.���!��K����K���#E��3�}�z��Z�o'q��R���z���=M}�u{�&�y� �&�9�_۰}'���+'N�3
�~��o�!�-�_�2�UpK�k5���т�n��ҷ1���Y!��}=uB���@���{]�
k�2���#mM1Ό��d^�\ןJ-�<:	��0+:LgwF��c�a2K)�t5��KӔ<��x��$m:	��it��'v��B/�=�����
D�A�b_X�lO�l:J*	B�����r����?��^�`�����
�wub������3�tM��/	�#�}�4����2.7H��}��H�Nr ��q?I1�1��v�i���������@W��3��?A2����]~�A��[��)��9����u/L�s��%pyn��Pƫ�aC,3������o�rC���(�q�;TN�l��ᇤ�^��)d8/��q��r��g��'�t/6f���tu���ҤC7�-\�=f���=�E���[�M�cS�]J1͈��T�S�Y�pw$�`�c�K���h������sk��p�U�����Fא��[��#ӕ�*�G���<zE-`�l�Xg!�N1	�Q o]a�D�8/�}el��JIH����gpb9K�������F�+�}��`ǎ�I�	�C}P�s�j�
M������ףt���<;�S=9^����Ri� �5xB�����z[��.$�h�����JQ�;s��t|��њ��G� �Ck%��y������D���F�g�"٤��d���;�l��%��3���U�B��b��&���]�w���h %:�Ԥ6sFĹx��pw�](�R��<�&��L� �o�-)	�Ś9UW�N�+�L����E�w<h��h(��i�Gb�&a]�\8��H�?5z���Ʊ�o{]�%�ۏ��sNʃ*��P{m��,���7eT59l�u
��p���^��.
T��Q�C��H�>�����2=�>�������pFl��}.�#���W�J�o����:AKvp��~q��G<'Ƞ~7jᨆ��d��:�w��*�_K�hi��|x���+څd����KBW�c��\q�L^�"��2܍S ��boL��q��/V"2}����m6�^���σ����q�Ȣwq�<�I��3�D���X��o�>O{u�'qh�L���C���''J�/ꂿ�8��Qh�c�fnR2��'u dװ��HOj ���(lQ$���oU}���GO)'��X�#�4������;���M=x����*����9hѳ�'�Sڛ7�:�q�ey�j����(?��N���� �_�LV�G-�]"J����@��EZ����30h��w��o�Z�N� ) ��m��|�#��k�>M)P��ŭ�,ro�v���W�7KG�P4�z����{�9]~2s��U \��&�z���TL�%6�>�L��+���zD��P ��	o��FD}�m̖Y
�f��?kE����'������{��ue*J�O}�w�g�N�u$�_�,'l�~���`��Dq�E�ǵ����!���vD�"���������o��jnO��P8&�v�/"uC�}:؀���p*�e^+��u_����,�8��z��A�!|�h��X2^�~����4��S���]Jp�}�|3���e�פo}�^np<6���)GT�q��I�r֋9�{���֮����I	H���٭�
�B�����c������Ϧ�e?j�Rl�.�R3���:[:���/0)V:{;ok�]��|�\�Wh>�tn��EvM�S�TM�`�����Hu����䨲�F�K�J����b�79/�cۄ�Y�Z��J��y1(��jǸ��*�Лc��]�ɰ��UњN����?�B[C�}���Cj��g�*�%9E�A�w���&ٯp5�ms��D�s����Ѵ�����2��%"8�9s��(���E�R��*�%��MN�������W@Y$�Y���*�v7d��ڮ��p �$�;4�VK��2���󋁅�z�n��A�&�\iq��[Y�@퓻��Jѿ	fH�u�Q=V�K�бEU��+gQ�~����)�V�̌}����h�/h|���yq���Z݈le�څP�mn[TZ�U'��p1�ZO�i�)�5W���k�
Xx~&��8|�0����y�����v�8G1�M�
E>��SOi /Ψvs	E�=��-i�#N���#w4
��V����uPB6��0V�7��#��3��\Tg��i쐺i����	+�R՚��Un��s�e�`Aq��;z��6��6ȳ�	}�ic���]�0/�e�����V�!� !i�C��܇��q�m=!y��V�A+e_�6);&���Ч�K}Ȣ�]�s��A�5� K��OgN�4<�{Q�_�����X��U�u�-�7i�m&eR������p��o�s�ItN���B��튅��+���l�$0�i����� 2_���9�D`�3+S���%>`�K���M���8�}���g�˹�3נ�3��G'�Yg�+�\���ƇC^��1=�9Q#���i�֬��0C<���U�w��d�)W�u�����A�#\��ݠ�3�۟�vw�8l�2�2BH#9N�"��Oin�#�O4O�&ֹTL
}vC���ӪUߟ������c*-��e���(�y9���C���w�A�k! �.i@�󛆯?!�������#P���?�T͖��w�`�3�2l�'��}8{� T�y�P�#l�r�߂h��S �X_���+�k˪G���@����o�x�̋�.��&[�O���h�5��J�y�@���9~|hdc]�i�ǐyr9��?��8>�ˑw��O��j����h������J�j��L}M��Z{PNM*��be�13|18����-���_�.�g��L_��<Ԅڕ��ԋ�A�����vW�ԗy���ᯋ�1�i`��Hkg�)����o��&l6ܘs��Y�d�6��tY�{�^\���o�y@ ˋ���K��9�|�&�����"t[�s���h����[��7	IAt��}���FV7��`Rz����֝��GY���{��&|^U4����TP��Q\&�?�6�@�(����ՍpF��
�p)��O�$��=�O*Ȕ����޴j�>̄����H�ig=c��t�"���qY�cZu�<�y��K�F< �V#�̵����T�N����ϸ�J�+"UD���P�RW�8s�z�_&��a,�<�WI'�\J#V5�$����|,`9�?#NC�葥��{ Y�RƛI����F��5o�>(|��t����n�o��y�3tX��"G 5#�:����J�F��I}5��FvP�nRD���C��*����1���f��419:�Ft��^
�K��ʺr`���&�5�������D+?T��C�����O�\Θ�Z��R�(�ٜ�<ۍUVb�n�v2y��:����c��4�b}�U�I��y�v�m�7{�oV�$=	��f��Â��,޽1��	!�ވYв-�(�*�8_���Ҷ�T�VH.ǹ�����.�@],<dU���;��*rԎ�� n �Q�X�(=Zr����8�#< �Q]���t*p	,���S��]L�3�F��;��¹�p>�S�k��0y၎�X�����K䖸�p7�O�8�,�:�R.WTe������[��6N�_�kN��U@��sA��k=�<g-T(�$����G@Y��qVy�]MqnN��[��R���QL�J��n�ǽ�0|v���AA�I���/A	b(�W�T�^f�� �4�1e�+U�� i:K`m�� u�o$�o3bO��I� Vc.���I���:0}K����c�^�rr���Ŕ�Śz��VQ�ڍz����LIY�br��iJ�֐��f;�����V>z�t^���BA��w���wu+���0�SW;u�QKb�c��u^�����S0��5�(!�+�~���Ґ��u�l�'��:|�+���_&��[,�8�����	G2u�f��>�
��Ƀ8�W#7��U�AD�����Xs��ȑ?�#ޖh�I�z��{9�LO��ѤN��e�d	��l*�[h�+f|t�4���]|�wl~��|���DK25U��=�Ɣ=̗��	R���������f��M�p{���a�7���v��J��6��3��}�%��B��S�����Z@D�����x����!*�`|*!G?xj�,�D9��o��qY����t!*b�r�#O(_��n���͛7���S�;MC4��ƙ�=��R����?�ט�@�?�������m��:w�c�����^񣅵*�i�Sz�fLo9��t7#h=Lqx�`l�}FŖ�!|� ���I43M.���da�pڶ�b��XA��k����!��Za�s���ϧs$u= �P�u�X�]YT=L�^��GX� +�8��#����7��,���m�'N�Vѽ���*�#@i���_���\�1x�TD�����|��6C�|	�
�'������ᙪ�i�$LXdZ�G�G��fkm�&����F����#�Ŀ�䬾�-~M��[$ܵ�	!���X p������qŶ�����Џ�����i�a�]Ә���V���������0=iB7x(�/�^���yBб�Q����>9/�9Vd���֌���E��@/_ü;W3	�e/>��O���Z���n�!�Ca�����S��݆�����M�vL��e�i�b��`�?�ry���LZ�7s�\T�']��iu&	����e���$�uz��� ��@���Պ1ZN���E!�	������"|M6�D���;����Ifۙ3X��,Һtw_:�{P��jf�P��p�n���`6�˵�b�S8���\��$$(����)�������Td0Z$���5�����2�����)��~E��Hx��kQ�<C�2B� ���tA���q���?�/4���{�L7p�Z^�?�	Y	YO��r�_�)�Nk���y3r�(sd��E2��Æ�Ӟv�-�ze>��1.�7x���C�t��J�~	�T}��`��3�R�ҬW��:�@������!�Z��v�g�lV�^PJ�����𷪰Ҷ���#��b��OWF�J��e{���v��1����%��Vp���@��J�{���K�ݵ'���!���*�q�]U14w/���Xq�j�AVK���g�F��ĒMrx���_�[V�I��!��vߦ�;s��n����m\�%�&P��V�����NGuu&=�V���p��ҹ]Ԛ�'QN9zݧ۹cS�C-�0ui�$I�[�����@���l�f{��L �k<F<��j5Y�4�1�~U�˥9�>�\�
F��0����w��CV��'��o��'��D�"��� ��c����-�.g�DŲn��w�痖J�І�|�*%	�S�{���	׷:��qvĮ\�SuopJ�.]-��4����Ӎ�/�l�ӌ����\��C�n�лxԐ�	e���O�(�Ÿ��q�������ZWAEpN�u����ya�{�A1�+ȇݙ���J=��ܱ6u�htQҝ�94�+�d�m?H�KdE���,řmC|�Cp�t�wi g�M���u��F��Ϻ}����4,1��_b�]8�zp����D-��G'�)�V�͓�vdhB}�	�]�VR�J[��@��J�v��46*��1��5�2�җ�r��I�:jַA&w��3�T�Z��I
hI�f���2I
���j���*]�ϕ���}K+ƀӆoiP����w��.)��U�i"�ƟrB�-�no��B��D��S��ɨ9Ϊ�,�'JO�{wc���c�'��5P���0^t� ��D��|��e E®�N޶���HUT�L[���bzv�����^6є�W*�R�vܗ
P�Zm�`6�S7IT�5�*�2����V��ڞ�^Y۔�8���:��^kh�ȦC:��� ���+u�I��G>�X7�q�j�e������j�&a�J����� T��~*�?��M��#p�k㩽�mH�(�bT�o)���b�j���8O��{��	e4���rc�3�(��cM�&W7���Q����=��L��'��)Ap�Uf봖��,��ݠ�dò{˝�R(?��]���s�Pyl+��N;JrdB����X����p�������KC �� -��d ��
�@o8���Ƅ�u"���Zی,/6�gF���(�	�0k��`[`���Nѓ7��c�� 5��9��;����OwA���X΄Nb^��n�}����rp� �1Ƕ�|[p�+��7[�x�)oW ����<�+���8-�ZgV�[}ib	���ַe�}᷆#0�Br �Ʒ�>5�A�ޱ_����IS�Oţ'b\ݧ�&_|}։HHP�c'A�o k�Kp���=�E�D�-ڼ�<���l��4l�n-EE]!)榰�ݰ��"!2𓝟�kb5M�e֞��U]��}Y�n���Ⱥ.]��ST;FoV����$���*8b����2�gE���邠��g���E[��g'�������/S�h�"�^s׳e1C��=t�.�܆��0���H��n�����	�"v6�(���X���X�h�]3mM&�m
L�e�,���̟�N��"l���F#�ϯ;x���Xէu��f��)�g܍�+����,�|{�'P��/�?���O�p��dP�
G�� X�&`l�i�J�Eg��%���!ܛ�=W�	�:U�^��6
�{k�28ƀ�C,EL�c5Ol%��3��尔��a��4�Ӏ�]�T*X�y�n4jn�� 5?��4'�N��z���U�\��|���0'=�mfΫ���1�Q�u*�l�?y;��#��+jR��r�@�I���<���Dg�Ŵ�<֖o[��.�#���17��c*�|�O�g<Հ`�e�sk7</ڐ7��W�XIJ�A�3T��`���L��=e@����orɋT5�,.�D�S?d��0���rb�u+!����=�gJ���^¹[��g�``_��_�,V2���1�g�����c�?o�R�!.�r��co�h4t��H9@̲+E���sM�%���pCW�(b�qx�R�x&)��a��i��cyw���*u���:����[��k-C��x�e���[�R�c@ݍ�&��Qp$�z$^���s>��(49�L��I�q�6l�8��V��{4��朆�S�/���u_�|��u5�M�
���y�و!�sV|�-[����19}�`*�2}��=�;v��P73�d������	qt����2Q@4��ĝ$�z��뚫��#��L�A��D�n
����,G�����ߠU��lނ+���x���{;�� 0-�w�Mk���¸��`�r�f��W�E}T�E���� ˹��T�RwF�2Զi���]�p-�*�JO)ξ_�'F��+�<O���V؝�;��:���$T�d�#�'&�t�2�R�1:V{ ���A+���6�͟�k+��/X��H��{�y��ax��v�}Z�IÉ���/�q�+]���J!������҇�'�p�D�мg��%��Y��	B��s'Px�����S��jږ�cj��(�!��	��Dҁj��,P��e�Żzk�!F��m�{{j�6܁23Pp�:<�9����D�������'�r�r�:��s"U�j����f���3�<������E%w�R,�5�[kE�� ǒ�u�H��q<@<8����
99�@03'j����-��Zɓ��N���Q2������b�����|ś{@�y��>�Yo��%�5���&U�dL4^Aʹ/z[�k�����^�G)R�����7�gRzU�gWc�6ɕQ�>(1��|g������t�a��Qk�<�\��ផ��;3�2�+X6����t�0ZO� |o�ۀ>$w%3�˸�s�C�<��S�I�	�Ѓ�&��čb�B�q��gk#��'sH�/VǇ�n-4 ��RPc���N����8��NS�=/%�L���n��ʻ�.P|�(����ز-����!8�=�c��m��t2�2��j֠n��=<9�\�]Ɠ6F�4�\���@�N���@��)��8�&"��$���E���@Q��Z�;�S��U�΢��]3�zh�;	0F��Wo�k���`֗���%�]@^i@����+��Ϙ]��X"d"+z_�lw��pKKk�3R%�k>u�h'����]��N:z^�1ȭW�ws���Dk�	W����L-:e;7�JC�&&�3�K����> �0э&A�QS$�Kվ�����t�̤�!b�;O,��8]�zC�P��� ��u�NiMN������*?2����~z�m}xry��B�W;A�n7�`��<ܮR�:sj�q1RмZ<x^b��N6�I��f�b�4.(90��'Ԣ�P�% �U�F�XݔЊ�]*9Ћt̉�p�8����er��J`�\|}l/�홻6:v_'	xx�S��c�-�K>w��-7��������촊R&h<���o�I� ���s��e�`�T[x��m�H�	��5C�iܚCj���V"��pxAL�d�ҸeL���e���M��[+o�AmO�#y� � ��;��|鿿A_�_����0�/x�&�0��Fz(%��PJ��' `���q��E��,���͎�*���-�0����9oY�Z���g����