��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�r�A�\xnc�"� �z�g�B Ԝ�:���ɴ�^����-�p[]tx9XHޅ��)��5��� i��]�jq}�5�Y�?W���������%��ѓ����<��o���Y�gխ����O3�/�)[vb�ޙ>U��xdb��`�R\�Y��2���e;)�	k.�3�X?+"�A>�����(�r�2��ӆ`uvSc��Ho�wu�%J=i�d�K"q/��<s���L�;6
�
����!Yx���;�ڟ���k�bM�и�U�c��ߙ/A'�C`y�i/��r?��l�m�e�j2Aԯ9��Ia(ǋS�=�#z���Sjݓg�l�3�G�d��p�B~��w��*H�����"7;��4�����kN{���Y:{2�/[ �cI_җ@���.(� ��K\����Ư�z��"�ٯ��L/�^�� E�Y2߆S.�䁔<Q���(��{��@0&�8��Xu���IWar�~�I�W��A�a�����do� ��G�p�E�
Y���Y}�V��c����^ ���lw���[�9��k��1E�,����uak_�yx����}w$ ���8`�SId��������4g߃}��<���\��8]��P�:��I�{e�Wjto	��@ͩ���B��]�
�P��f�;�R���@`0FY��V�ۺ9O.L����|���IB�Fi�?Y1�o,ú
͵�P�Tom�w�>�Wƙ���[Xb�Z��fX
�颱+ߏ��}Ø:i8W`F�(�*����ڈ�}�W�7�D*w�ɕ��h�����g纜h����Dߍ#�-�!�#��ή�؜�����#�&I/1`*�|�}��񝦛��_rU�ʞ4�����r�(R:��ݪy�ى��BOp�G�$�n�F̌9�;�Jh/�*{K���I�`��ó���(�y���ͲQ`�h$� QCB�rHA�� ��\�f3��o����A�bgQ֦�O�a�1�^�� ���ڜ���t�N-��9�ϸ&̠�pg��
d��<cV��8�/���3�/bq���Xz�n9{�=��`J�P9�iR	S�=�m��|L}�����V���?6*Ü��A��YR�2~��4"fz2;�`�8G���Ȟ�i����)�Hm ]�����5�X0e?>[�P1��֜R����b/젽�f�x#�2�0G�Y�C�Ov]���c鹷�b�މ�P]gO���6]��\�q�#��y�J|��ÿ���z�U{��uy����C�ҵ�V�Ŀ*^�  ��RC�̑_�(i:��w���H�G�y�;��x���8|�K3Z�?��檓��AB�	@�[Z�M���U�6�E�_LX���/��#7e]��%�*&��춤]���L>����=B� ���]h�H�z!�J��BQ�"Qé�Ft��@��u�m��/Z�����@c9�ˀ��t^4V����	�W��Fi�r��s��et��Z�,a�Q'*����~~�5^c�q�ڥYe)�L��\X�K�Mx�{�h�����ܔs�+o����8��{�N���sM]"(�6������I��w.6U0�˕��3��(T�{�b�Bk
]�����y��� �0!D%&z�����Z;��<).s�u�h�0����$��V�hOX^q��i'�xT��3�:H��O������^>4,i�|,���������|f�\��/�i�u�%-�DN�Jt��l���W�^#�Y�<՞�{.V�At�u�8�g���s�+Vީ�_BLϵfunK��:r�%'ho�%\�6�Z*����nM�xT�v��	`Y���ň��Pk�躬�:Ux�
+ᜄ�b};-�>�=�lF��:/ɇgo"`�$���U]�K��t�}cl��[��D5ʠ�����ƺ����"`���/V"�-0�Q^����W��/Ch�$��c���	i]]�4�\�8o��DZ��������w�T�bڶ䁒>W���<zﮱ�����7e�nQm�
�_%��@,J��t�I@E�8�U��B��%$;��܋g�5D��C�s�?�xFWs\2	��_�nn��p���`�ur�F������)}9��Ǧv��:�\�V{ha�k���>h�0��l�R�y(��4܅��Uˈ��LX�Qַ�x�	�M���l�w��S�x��z�"�E��w-1�Go�o�N����������Y����=���e�=�*���,\qS��A!�k��B��ß5"����	<�_?�$��:;X���� �U���ŵ?B��P�=$M-�6��}��Z�8������ǉoLj6���n�(m��>�P=�::x}t|�7�M���Vu�TiTH�η���:��������:����[|n9 �V�;VDEg�IiW���F�����;مQGj*wd��Z>��3��~#�a
��l����bM�� 3��O��=��b��I�́X+��^�`h�2��2��I��ʴ˗��m�����ޏ�/���?��r��}�o�.�+�3��oQ�2�\r}\,U�+P�*�E����g��߶))o9߭zǝ�:=8�vF6�������bfz\����u)�A�W�LfO<
+c�rXo4!��y �v�C��b��\�/)I��.�lJs��팑�2,�M&�/����ծG�l��/]�Q:Ș)�U�[��1���9uOP ��^�]�pG�����]��@�����6���^q2Q{5^�۳�ذ�.�_��Y�z�̗
w@��/�5Y=nBzT�L�?��O*mL�"�Ꚋf����D�(yLi�� �C��U_���� �hP��Ő����[�uK:|��!��"�|Awd��C�C��[ː(XOJ����P>E:�!�^�2�a{�Ի�g5m/�<������O�������H�6����Ĝﲺv�*��Y�4�R�<�����`�6Vw~𳷰���*X��������O����<�nl�y`���q'�s����ϭ褙f�B'F�E3�[^Ru�����Jn�h�*��<��]��W�Y��y�����7�|��N�աB ��� ��$�� C�s�S�[�X'x��,XK�z1����%A�waMG(ϛ��4|���o�f�T��L;�M#���1uk9x#�b�8?8c7�g294~x�I���XQ�(Yꉴ�Y��fl�v�~l���W�z�_��&�e�Ik)�q�\_����_�^rӈt��+�5bh����?E�7�W��7tGDz�?#�Yl���q)��{ч���������ż�
'�:jxS���6�]IZ�
=��׵n���|�}a ��ns?5Ë��'������m��a#���3@h��˯����vЉ�h)��y�A�F�y����vyY��Ԅ]�N;:6�i�B^5�Y��W4NTFܾq�5ƍ��%�
�d��lw#��f��m�5%4Ʉ�x�W���e_�Q�s9���1��!52pN��`����)��6I�N��߆��67W�w�2ʰ��#��j�� �=�I�^�L�|9��(��	�{đ�c��M� ]�".�����H����vb�A+���p-=RQ�w���LV�lY�HV*��w�� @&�nHMUp�hkBrh���bE";�u��\:�g��$�F][+7�@�g�\�� L(sp-	r��=�̕$>��Mw�U�Q��m�z��h��S����ȳ�~��h۹��]L��`�pD���m�k�8��Fg�+�q�t�� P�ɚ���{�� �^�'���̝�n�˚]Mտ����9�u�BD�u`z$�P�v y����C�	?�������"� I#>�/*�L�s>+�	��+t��7���W��N�K��WN����5�"q�%b�m ���
Oi��_Fv���Ϩ�+E �i\H���[�p�}���f-ц���DBbc�N���L����� ��N�$�7}����O����.�2&^w���1�y�[����� �{t����?��$�?���7���jY��Y��,*��@�RcO:i3������֚m���( V;^@�LOLf/E�̆K�}X����0¢�'\�Q����G5.���i��7�Z��$�xJ�1�)J�都]�S\.����/�	�IE�?5�
c�v�4cP��wuU��t5c)!���37�¥2U��`RO�/4A�D�ՖRy���o��vu��^T��z�#�6�\f5��v���ړ��`bz6��V�UOnᣁ�ƥa7�R�j��_���݆'Zp�~07_��E�<�HѕKeg����Dx���3�٣���'Fjǳ�i��LÂ���|ɏ��P\\�C�h��6��1��i��I���3��eb?'�k���B�_�*;L��$�����q��Սҟ�0��z띮A�9-���I-��%�:F�nv����������6#�8���i��2� �f�'��;��y�71�'�wd�a��
Zm��ƕ��j�x5��ST��`�u���A�f�C�VDdS�e�2���m�mP���9S�� M����"#ַ�i�9�E!_��G}`v#�6����`��_.ؑ|Re|>���
��x��lq��\��ĊĆ���~.k�*��y�����E�Aj��?�><��3,&�|.-� �q:����x/�f�s�q,$��&W.,m�ID�Q��L[+9�Q��G'��}�\�e�Ur��n(u#��oL���#g+��՛>�&E�9��Z� %e�u-���G�{� �{夑�?^8
��H|�O��רU�#��g%+���L�G����_��</u�U$�f�u�Ӻ������G�S� �������j��/�~W�8u��NC���#3d��{����]�D�~�v�^�6�xu���v׬}���# �Ԙ��<�|L�YΝ6���l�i5-C��?vT#^=������`*���6�ӷx�iG�w����E�BC��9�	=�n�.��L1j��n�1ӋQ�S{C�۫��~�;�� ��`T%���&N�ޭ��&D�/\}����x#����~eb�k���{zo��ɨ��ۅEu��07���d9�D��.�������?�҉e@ݕ� ^��pRX��7�fkOy���Ҿ��u�҆����E�3k��h;	���L�!�?k�2�=q�`��Wi̃lp6>QZ�1��c��`�E�����r�N�D(T�3�����M��p�Ux`˔N�cGbU�����^x3]�����+^_"�v�k�UrAPOjI@���N�ljǆ�����^E��Yc��M�<s���Ϯ�S�&\S2�S�8��޵K��ZǦ��a˪fOؤ`-�519�t�Yv���#�W��?�w@d�H�����	������+3\�ׂ�0E��)�7�b��yd�� 9��S�K�M�#�? ����Ǡ"Δxg����b<�O	E���S�d�McR��3]�<u���{ry��r�O�2]�@&��d!_��,�K��O���-Aѯp�C��!O`�2u�/+K4��{erA��A0ut%5��J(�w�SÐ�U�uM"4�3�3ӤErϧA��p�^_;�x��lۄ����C�b[��kJ����qS�����r��A��P%��o�|�"�5p�EX����.����N���)K�8W�DO亅[Bo�����l"[�O����#�IG�6YA'7	Ŗ�j)bǗ��O�H�:���
ys�)��]3�	��\�ت\|%�����N��sӞ+���3+�
��t�H�P���������U=���V��:z�d��Tۇ�׭L���^��$͐'�*�b�!e����Jkl_К�a�R�͆tR�LX��� �	��
\��nd�݃u�݋��mǬ'\�u����,L�����̌��Rư	�~�2�W��o9�ؘT8
F�����u5Ԯ,���XW�:�hx^��c���P�� �ā8ڇ`��4�d{��8�<�3����r�\�r�DP0�����P����zҝv��	�g���س	�Q��[�Ъ� �g 꼝�����?mV�cZ�F^�:e�֐�7��B�A��U��;m�E�={�3���r�#B;;���`W�_ԯ3�
M�4�Dޏh�ϋʃ������{/�f�B7�����*_1 ډNy�@����7�̉�ë}h����,H��We�'�hRH�Ď�Şh����.픖z_!1��Jt�jY�TUb�ڨ_�z��j��?&_l�}��A��3%Ч3qSK?��3�d�����m����$\�)����S�M�!
��N��b���F����(du��6W��A��J�=-�O��T2������4
]쒕^)$KTɨ�-5�b'���0/�d�+܎-��$��&�1�9�hr��;�J�Ph3��~�G'�i�a�gi�5��T�9Kn��`��O�5�r�q�W7X�=�ej|���M�O�}
�9i�\̋�Z�����Z>���ڟA5��c˺�����3Ex�F]��,Jc	҅Ȏ���iA����Q�5:��Q5�{��)���,f��sO��y�/8o���c.�����蒸�7�il[U�����&��X��$9w�\�>������ng�AsK�c5�56w?̗ox�&Fj���x��<�H�Ag�ev�K����o��������A�9-�w���p��$�ʵ{yŶ%��b���ӕ�5�gF2����<`�IZ�������M9�w�p�"��zB�h�M`$�o�A��k���H�=���E%ů�o�����8�j����8$�Flf9~2-R ��ՔaϢ��g���Ro�N ���\T�lx	���&���� ��B1f��!ec	R���H�!����]�O�m������8vw#p��9OBD������Ax��"���2�kH?m%������7��u����=��O�2]�j�\��^y���=��?�_4�� �-���ײ>�$�3�5o����U_}�?��O	J̞5"�0?�ǋ���+�~���R�����,�70����504C���C��>Z҄�7Y1 Mq@${��fn����ѮfX���~u
�á�~/7�@,?B��[I���)6��U������4� u�߉����/48��Ձ�4�=�������[
�U)�*p�-���خny;�m��??���|Y��څ䆧��Ԕf1'��x�TI0���hќ��A�7�(��s:��*����ةw������ l�`�ծ����J�T����]��;����O�ll�s�����q)��ke���j��}*�W6����N#ɼ0Y�B�t��
6��~�[��G����jJj2���wp]ck(8�e���<_ r�~-,�=S21�QGi� �jP�3	v����"А8��)�ȤU�/���h�0M������^�u�ہc��d�a͙`+�����
�㜍��]aQ]1��.ړ��W5�`�T%=bV�񁔙6{�#Ѥ�=�Q]tn�T���g����|� LX:��U�\c��P�Q`�����Y�������*�p[�ڪ���q�)lc�a�!�?0N���ᨀ޺�1w�I8�f�6OY�B}�ꁪ&�I�39b�y��))�r�^6�ɉc�N�}M瀷��@u���Ah?�����]�4T�;C��MBLb���>5(�z=�L]/Cսŉ�,p� �Ր��
c�\�/����#��Qp���;Ԍ*$c�Dp��@2�����܁��=�	�����L�P�?۴ߘ���T�֬Y��AFs"�d��o�W�����4�g�M����	����7��f���j�M4��җ�/��.��
y���޶���lJo5o��W��̧�uU>�LI�PH�Gu_[�d�Qk��e��1�$� �/�!�wz��;<�e�,ڎ�RVe����d�Qt~+��a}$8�N� �X���y�S\eR�J&��JH�!�Ț���=�/bu)��}�����<vQM��`��Ҵ�@��ݱ�S��HD����j��7���P���9V�O�����ATW�'���i��t��h���%�3m���p�R�HK+��5�9�	%�]A��Տ��ڲٜj�f���`�a񕱪��.Z
�x�B���Z�o����9,U������Zɰ����H�Ŗ�@�O���u�&�T�
���	��[�8èihK�%�{[/�pe�۪�b�0n�&�y[Q$�8b�Ȏ�A:��u�������6L��a�t�^i��sM�S־�U��; H�-D�9�O�n-虏'b+Q�����6Fp1L��є���֭��/�c�M��4OT�{%xOe���#5�U�b��p>3���b�%ɠR�TF�}Jky\(F&c��2�@L����K>듉�I��\�dJy���n��?E��o�� ;v��� �i���"��Z�tJͯ+r5�h��]�ʍG�2�*�<����CV����8����;�jڑ�����A���8RN8�.��A�+­���h�~�k>iI�rԦ�b��9y�/}��kˢ�Y��e���*�o��z�i�81�F#@�QN��ttр��f��9k�?	�5^�������M�;�`5e��u���:E� �o#�3��(�C|7��s"�/AHe���A�#U,��缙�����?Oc!+�0�u��43��DE	�r%�g:_�/6t� `X+�OF�R�������t
OOc�N���Z�d �&Q�S��U;��]�PW�@9%qM6�T�#?�a6&���K`2�.�l��7j�^��)A�#��~����3kNWn2��Ug)��d|���:Eޝ�J���ř~�:�Hm���"\�p|��Ba�������*	O�`n�TC%|u�r�6�^+)5�ǹۖ�d��WP���s�N}�:���~��_���b4�C�>k?a��me�^3�אc�5T�^S����)��������;�����ѧ|�X2����K��&aO�h;Zd�铝�LQ�"��D��٥��U�q�p�X =�!,��4�$-#�n�
���cZ~n'������!,H�`�D�����(��^��άyvnם�l�=B!��sY��pl�Qz��Md���@F��	~��ż��tN}�v{z��:J�|�S ؉ �����b{x>>{��n�'K�����w��]+��q��٪�	���[��(?m�7^�	���Y�8����a׿=�ץ��!�~�P\�Ih%J%oM�݂*�����d	��g��0��87���W�e�
6?V����c�&dՍ�ͯ�XdC-|
��J߬�$[ �4��>����F�k~5?����]��� r��\���,����k9:A\�Q�m�E��
҃�EO	KU��,_ht��F�V7O���I��eP��o�ޥeP�H�3r�v��Fmg4gt���q XZ�/h�k�k�V	G�5����:��8%:)���i:���{nAZ�u�� a3 ���sh��x�N:S�v���[#Z���D)�	;�W7T�w� ɼ����s��Rsl)���f�m�?n$����}�/���5����kx��;	>�C���#�A�n@���O�˙�w:����K�y�(* l숪��Q�{噪�7 DVk!RCEؕ��J�~�? ����N�6t��]3\F�N���`��؊
���&���˰bA1j������1�x+��9�@�^T��m�R)"�&8��$�[p5Q��'�t\�a�F8�/�ϑ{�m�P�|X�~�/�!��CN�E�f��!���	�p�kC�����cVe	����O��L���x/�h�b˺�v�Vs_Ll4�����yʼ�*Ȓ���<?&�as/��zw�~ x�O3�,�Gt:���Ѓ�l�l�Yn���zFw�up�$(�d��1�H��dy5���B��n��W%$M�R[5(ӝѝrR�z[ �A_X�DOs��x��W)]s;Dq�H�:� P��
�)϶��$!��oI��8I�.[���?��m �Ìi-����GRoeb��
��L�訧Y��Z.��oRQTA�����Њ��Z�r����x7]S���ny7N'�
5A$�������mm�7���b�^��wz�s����f�����.ZM�� Ei(^s�7ӊ�?�H�)���N�0�*15u��̢?X�Wi���9�n�bN�!�S3���r�,k�;�vIT�t�R�8!�v-������B�� fX-x�AP��㘎�����}�Z�����^! �Y�kϻ��g����F�@��)ۮf��TN�/'ϳ>o'��x���R�������U�0RQ�8[��M�A�[n+���7�Qj���c����!��9iVܑB]և5���9%�~�k����W�����d 	��r�u7v��b՗��\���F
]�s���N+�$p�h"�b��5n0�
4�Jg\��8ڰ�Z��ǜ`�gc��X&�j7���� ��2O�%��j���5��.B:�i+N���;uP���
H��4Z��R�h\p�Op�B��2"�����eR��:H'#��kx[Ih�y��{0�5������ݞ.�����/���.[~{�Ӓ�d�!T�ٺgZ�[�����o�g��'96�����LO�Z}Љ�d��q��` ��g�x[P��=]�lqҚ�G�ٻu@�Eh:4q0_��Mh���ʚ�?�%��¡I��!Hd,A~r�5�S
��2�����7�_�2����$`U��5!��c��6��/P΋�|�̓
ps��.��Q�܂is���vm~�e,���a���M�M��LB��ױ�1��d�i���1��Ύ��8�SC���RῶCR���/�ς�3�;E\b��}�'�2D��H�Ä�~0��Z�F��j��Y�����(�Q�`VH����n��T2��:�Vr�k7[�*k4Tm ۫�i��.\ĩ����+���bG���ߗ��i�WV�P$c��g��>�}��"{�6��8���lL�� �CĖ�H��̏VKۚ_͔m�c
7�^�|/��m��`��_�Y���|dF�W�~���̊?uҞ�h=���f�y� ������k]� s��_ �~�Wm9�r���(��GSݸ�(��W�ꊻS'��KC>J�R�0	����Oٗ��Dx��BL1�J��$+R}��X�
��,�C�g��g���?ɹ]#~�m��G�0��\��Tǚ�cغ���E�k��s+�_�[�=o�fX��ø�g�� ��hW�O!����X�dx`:�=E���~��#���g;� �㷦��Tb�m�W���ے�4�X��o����u�v?���n�K���H�1(�H�������)]%W�`��QT���ê��:'��	H�+Ft�I��s'R�np�恫����	*m���
}��/���s�A(I�]�cE��,���%u]rݎ3���^B�R`��%/fc�/K���T޼%;K��X�i?��a�BRG��W������&�@D�Rp�ʵ�� J�}f���-�܄@U�#e���d��+(����}�U�����=�3-q��;I��aR��ٖ4|�S���'�z�5�P��5/Mɀl7Ro#{�H{ᜨ� ^�|�I�I�ɜ��c��� ����:Z�+%`;����4�8�kD�0ӳ���2tˣӍ\�|�(k1��C���dS>!��d9�#9�η)D���;��"�aq�o\��M��O�>��F%.�u���kG)qTR���QsH5r�?%����V��FJР��Ztf���\)-�\v���t ��V뚲Ky�Yr*q<���� ��R�)I���@�+�����3{:��^������p�Mc�z&�L��������e��!��N�^�n����֒�9R>l�j���7��>����u���P�NHÉ�C��f7Iٗ6���ٓp�)8�49U��\�O��aOL|��ʂQlJU O�nzأ�!4W����"�E�� ��CNd,^Pu*C����n 7�
�eD�$A�C�y`�07��.������Y�+� jHB�#M�0vM.���xG���U9����:ǒ b<^��4�� `t3��+�2����)��FJ�������@Gn*��>�쯸�I;Eʁ�tɠ�	���p9lN�2Q7z:pW��*�}�h��8;�%���l`v��&f<�L�S�y�/�"ƭ�0G��#]I�����L�q��L���fZЎW�7�8y�W��4ܐ�@���8�`���901��%�+D�1��(ЂN��Ĉ̅�c.�����m(����N�<ߊ1�\`�;0$���e��Ip��޽QZ8�s�	��jo%�B���tf탗���vވ�owHo-PY/
���¥��vȐc����p>{�Ѭ��է��i�o_<��M�ܝ�+�S�~c͌�?����'|�0$_�5�K;� ��(Pݻ�I�ҷUr؞�2��O������Pte���;���ЃL�^��hb0�n�����ң^�0z6�C@Y�+0��ƚ:��Ɛʞ;�킵�{S���x2FS<�½�K�Y����䛋	�x%ꢐ	�5+�����*�X�42X��]^�9�+�i6����x"\��"�y}���$3���7�6w�VԎh�p��{iG��+�j���H������܃=]ox���׹�%Z���T��D�]s��^g�>�ϳi���L*�E㔘�%�p�b��(�÷��|�L���3�_�]w�6�p��m,��P Owo�b��7Ó���� )��")��w������C��{9�\+�?VO��x'����+Η���̾$�C�Í�2�w��c��U��ظv2\�5���y��Pk�Es��&�M�eq�CA\T IiC��.�,G��l��{�9�<����A/�,N�j��+�Ί<◴c�}]�r@�;����Z@'�{Uje�Z�d�՜���j�>sMA�j���
2J��$�N��UVt4��,x��yB�]$�á���$&�Br��X�d7[��g}l��[T�>�l��'���P˵O�]\~P��T�{VL�?���Ws`>ֵ�x�;eOķ�tG;x�F�$��75��h�4F�=��G�Ym����a��f$�O������ЯyM����#�Z�QB�7^��1���� T�h[М�f����+*=0�D�~&P�ձ�6�e@��}��F���8�����Q�~��N�h+��z?�iVC�0�3ӕh؄�i���^�b�3��XE�9�
ƻ�)3I����3-s�U�ҍf��XQO�{�J��kLl���	JC�~�����ǠAX��3�W5̀�]l�E!�^���A��d<k������:si��{l��G���?�i��� �C�'�I3v^&�/8Tg��X�8�"Ze��!0�JH�U�#��@�r+���6��'��k�8!��=;�L&�.�|�;�Su�ح�Wj�[��&���X|��$�Jx�4ؗ޼��h�xp���`�EF�4�I!Ne�	%�,�]Щ����+9����E#^���m���Va��,�aj[�/���*p�AF�ͭ"d<���d�]��,�W���}Ui�F��ѕ%�����\���m!-���P�.��{��f,�t_��n��{	��%[�����oJ1�
?��<B_R0��Xٝ�#Iލ�2f�3:�yl��b�T�,�ޅg�#S�;X�� g��}��,K�Vtu!3v'���$����s�$?���0}�,'���vބ�h�t�)�qa�

�՘�X5t�X�>ʊMw�q_�S��_	�I�*"bz-�����N�	��WN�z
>����%~Ϙ?��P^����˸R���4�z�Wyl����_kwuб�j/@� `�a��Y ��p�ԅ,E
K{ֽŧ����e�׭�=]V���?��ov� %��i����|�����$|����i�1�S\vy�x�:H!N6>�����k�3����x�Fݑ\vy���3ِ��_a�_��j)��z��>_]�KሌG�!_)���j+��X�H�=D5�h�����F(?a��v�3��g�
&G�_�S�#F����&A����$&u{d�|�|M�#.B�&+�l�YE����D�**�<sV�"*Om�h����L�\��ܪ����{�~ 
.8x�{^
�}5Q
b�73�l7�
�`�>T��JZҏ��>Sa��=�X�-A���r�h�GU;�Z�����F��:�:�uk�z�Z�����f�S�m^��w�.$05�a0k��,�4<�����p�����K����S?�庭}to@r:��s�7��Ȼ�f_���$�z[�X�݃����� )�1����NQ4��O����$�o�}e�b)?�Ư2#"f�����0FJm�m�[餪��Τ�� /�͢L����2n�����(��sSN����+��P�t��):��%�Ds
���l0��$�ӥ%�����1 �Pu�I��@Q57� �x!�\NؠU'IVc��ǆ ����e��%��2lR�ʕ���a�(�E�Í��$��t~���Rb�����-���$�{^�	���a6���	�E���LL��ڕ��'��>Sz"�y�rdk�o�c���$S89]�n�� [�#Dhr{��w!�
�=6��6����yM���N�Z��K,�OBw���[Z�.B�䃔He����7��ޓE�q��ZM�aV�x�?:�ʕ��:@�Ξ����
H`�E&�a&��'F8-�`Y�2?�3gyh�������pR��B2�!��"\��������Bnaa-�nC�±px×�j���eC+�X���cTzKZ�$U�*)�׊�+M�&ױ>,�b����i$�~���{�C�����(�4��H���H��@�|��:���{�W���Ciϱ��[FC,_��n��2���҆9ɔ�����(�T[�=,c���_�_�[y_���,��3�vRǼww�������׽�.���Xd�N�x�Zeab��w�^q. 	X�{ė�<f���3�u��eG�1��e:�*�=U��Lb3��5ã��X�9�[Jk����(OqP&����f��Z�\s����l8i&U&�uSո{�~�v�j�0��8H�i}Mt�j �Y�!�`�+�c¨���A{�ƃ
BŰ/�������G����t�����+G7��B��}�t�	"��+����2Ҟ��@��5lO������y#~%�qX�!~,Q0m�����^�8��T�l�1�p��0L������}8w����cq眱���S%�ʼ8e?{Qٷ��eq�-�^��xq�׊��l���J�Q\���#��%̷�w�[٘�Q9{��Z�+��Q�������y)ي/[<E}���)����kC�G�W�u���]�(R[�Av���U��A�"]��}��?c.A�������ИA��r���&���J�E��	.|�=E���_Ț1��Q���z�nnX���G�	+:K�.T_�d��K,h�q�>�R����U���4�Ȃ�^��q/�hu����WV0;�����#���
�Ī��Պ���S��{R�B��=��bg���
r�6����\}q^B���H��t��N(�=j;�,B���C5g�U�z�(�'�g�.~�8��k���	Wn��o�u[Λձ��d�O�)ε &+?Yr�	X(�J���#<�E�*ˇ8�
���:��^F�
j|�ZΥ�w]�N�}��!q��*#�ո�� N�jҧx����0���i`����CUUA�.���8�9�L�X��&�����&�5����4h�jl��������9��/,�^� F����-д�!�TA;�c�i��*�#-�#��a��_mC6��L'�|�Wqq���k�cbN�!#k��k)������������M��8$��$����x�	k�[&��d�h���M�֮��D4����!3�3�>n���֙��f;���6�qBU�xb*�м��{�vǏ��x�R��Z�)�Gtb��JG��X�������&�[��]�ψ�Mc=���τ�,�)�M�f�T!� �?��^� 1�1�+��0�τ:Ō.A�4��uT5�]�/	��T�n�d0��:U{[!ѯm�p��N�n��������J��H�S������!D��T�Dp�']
�r�KF6cHFV2S�n���������~���&�U���TL�KI�3t]���Q�qb>�\�4�˽�"�w?��� �x�:��W��+�Ņ���@���MJ�Xn�8B�,�VjȌ����Ƽ���|�&.iv�]��%z��q��Wꖘܺ��gpB�$�6Or��R�SZP��eY#�I7�^�Xvv֝�eJ$k�st��qǢE�w�� �4�`8= �P�p����c�$;]�3�ڵ���^'g@\��U����hB̙Ԇmb��r�f��F��Z��E���=T�{�TV4X9j��/��������{i��]�lY �h������,�KkQ��j�?����-��f:v�5�4��r<c�����NM�Uf�$����b��awe�zȀ���4���T0t�(O�{�I���OH�4�9I4��-&�F��n.pcP��f��9#2q�Ok��������돥_s>�*��ʍ����.r=��G��3����GS@�쇛e��]�>�(�&�� �ʰ�)��Z�Y(+����'�
����'_�C	ӧ}����1-�j�0,$��8I��Q��+&����r��>�X��u�����"���AOA�>ְ�������/�������+`���FP��v4�0{( ������3ZY�
����P���2�3p����4.MG��N��/�0�f�/�!��0��/�����J�뫐��QI������]��F"��Z44�1���&�<a�ct�=�1�+��ꯨY<h'b�\����]�^^�F�!��()�֯r�۱7
����v^�v���������
4��X	=B�K=�c(8y�Q�V��O]|��&1U F����P�jQ�{�)�6��<��"`-��F�z�|F@�x=����R5[��ìa� l�4�Q��*K+� &v���|ۘ���g#:lOP�A6i�u�;�κ�BZF9�c�%�$��B���:ֳ�F�#���?�7��Y8a	�����W\ձ�Ptbd�"�܉h�a
��(�ߨTLu9%$�
���k{g�u[�u�J��$F��#�U��a����e���n� ����,S�S�����X=�aPaN�D�錕�Ȍ�����ę�Onb�^^%�1sy%B���T��EX�1٨�mW���+۞�Yr���w ���ţ��+MUd*�O��,ԋ᪐��K���A��E�u��W�%�L�1�m+.�M�9Ei��x4�7�pqN)AW�Z}ߚ��>i�nB}�]G�9���f�n�/�v�e^K��]�I�-ꇻ��($���ڡ��8�V�f���OV��,�9����r�Z-ͻ����s�^|Y��������A�/`v,9^��{n�$�đ�rκ�1nCܒw2j���f}防�i&UH���뻣�4)H{ټ����͸�����
`��ɧO��Z�/��;3/5mq8��H���sVޚ�F��0��|>M�x`X���D2ك4��D�����u��|�=(����o����S��^���g'U�\�X"�8}�}k���%[��[O+���S��3M:�D�V�K�XEw<VZ����녀ѷx:9��Pp�yd�J���m��,-1�bo�f��jYd �Ϭ(��4��u34�i�M�}C�6��'�$h���M� :ǒ^^���F�m�W#��Ց�n����)�Q�\�meX2��A��"���%��u���I��n�N��}����*v��ꡇ/I#��w�'��}��zכ_�3�"��tӻY6�5taiW�R���Lc��J�6���Q?�T?n��4���P�"�Hh�������D��j�Sh�,{��ؒ���զM����[�(Վq;u#�������:{pcaMWR�����rvѪ���m���S���ʬJ2�
����y��ÿ��Sg~�>�y1�)Ѭ�%6�U���R�T%��UiA�v�Q���Tq6Zĩ�)���
Gs%Ǧ)���G7��Q)-���].�WT��˕��/j��v�ύq��=v�rgm�)�����A`�4rN@���j�5>�ϡn Q���|�D��p-�O��y��#�y��r������u!������ؠr�|��$��+Z\�@�>�2��^r!�ņn���#���2z�O�h�uőħ5r�h����`��e�1;@�?�#�ѱm��}g"��/�b���Tk`E��+����	���@�
U�l~!tGȁfP͕zh����=4�B�{8�2ݓ:�/�5- ��!��.8�țf�ww�EW_��bX�4���@66-h��|y���v�'w62��F?D[��Ii:�|f��GT��Mn0fC�"��
2G릎s�JDeH*��k��oD �����ٹaP��A��#gaS{��I���Y9�RmeY{�h.�Ni����� ����L@Fg}!b�(Y��FD"��I��2/I�U��ͷU7 j"LW�?W��]RwK	��ɦG�=<庒q�"ń܄��f�C��8�Ez�+�%���`�m�cC*Ǎ�/��'�o�(�%m��.E9�j�R[�<(��9�����y���8\���+�6
�Y�~���NCI��m��XἻ���W�Uz/4��o:k�,�R���Q�5D�y%����%Ԣn21�1�jߺ��D��"�W{&�s���qp<�뜇�N��t)anB�r=��g 0�Hf}A����
n���^�:
i\�=p�}�:Ew���z�G.M.���ld�	?�7�}!=��đ	�fC�Fj݊&���S�e��0+��2 a�5R��F�
�O%�K�Fl���v �`��n�&(�n�H�ۇ*j}��  �T�32CIV�)Gz9�H��|�}=�<�C����,�ގ�lʧ9�^F���>���b���]=��R���Ƒ(�ȭ@�
x����P�+.�i�>��f�w��ɬ���G14_#�3�ĵ�r�wV����c�Qs�J-��ʂ��H BΓ�w�"��-ܛ*6Y����'�ʭ�z���j쏧�j���ݾ_i~�_|+HW�ފ�or?���"�\��}��ݡ���]�����m~,�Z�x^+ٗ|KS5��n���[p6p�Q&�1��/�ܛY���Jon���-̃�#� ��g�6�}U��� �UX��a��i�Nˀ�~%!�	s����V�[�;�&�.Kj�@�Fe�7,]��w����~���Q�<L��}-�F{;�'��%��G_�ރ��4ti�U>++ ��U
Y� &})>r*�5SőJ&���X�4�A;��bLv7�}��EҎ�2R�cl:��W^�"�L�4K��v/Ĳ�k������XJ�p�5I�?`dJ|ڐI
F�*�C�A2m�~�v
�$���&50��a a�$�Y.�z��~v�10�}�@>�od��yO9���'>կ!�A�5��E~k	b�'���Gi�l�'ߙ�cJ-�+m��wݴ��a1�d�����n��>��Z9f�)̊t,�N��!`�GG=��|���Q&��m쬪A��Ui[��'����W�D�c\�?1W">n�z���E�8Of�r.x� x��z5�E���M/�\<��l4��E_�x�S�|O"STO��qu�t'���Ў���Q���M��=Yf��kC^����V�m�H��p^i�c�w�����֬%_�3�$���#�92���]���l��+][����Q�Zp��e��|LB�$���N�O�����������S%K��U
��('	%h�����G�?yC-��b��\rgc6���b��x( s�Jg�}������q�� )�ǻ�6�'�+P��b�@V�[(�(_
Rfu2�}�堆�c��J���at
w#j��*�^��s��筠����y�nl:N����N%'�f�^�6��p0k��nI*��
�� ��D.S�<�#R�T����Ĥ~o#����X��{>�E� ��W �F�*��]N��~��
tO.��E�=�FFC�V�R�G��z��R�� ��8�W�a��A�j�5+r�	:���}.|���r<������6&�[Fn����D��O�8�n]ٗJ"?k�{�����%���Ln{\-������,�*�T��
u9"[�#p����P"*�7f��0�x2���]��SZq�_�s�︇�(�$j�*!��W���$��+`Hܻk�a�,�BQF�6ji)L��)�L�E9��A@��O[�y5(|J��*kR��s'�za��U�8?�&ְ	x����s&N�H���v	���6�� �%�d:\�B�$����@°�J���F��'߫iǂ;o �*L�4~���F���q����mdѺ�Pi�h�qT�n�R�ܯa�����W��I?.�wͧ��8}+g�a)$��ʃ�	"�`�`���H���`��4��������,��]�=-�oH`ޔ�*�)��v׍��Z��Io�٩"�6�]�2����킫a�Ӹ�H���R�{X.&����+��ק����.,<�N87�)X:>xo^w͜�}��1����M���۸g�-��m%5F��s�n�2ɩ�Qy0�oXn�k�!8g۹��2��
����r���`�'�u�%�H�1���e�[�,��U�p6` n�u�c����8�QU^�V�,�X�0j#k/$�e*[�QB���:�Q�i�o���љ!D�oR%uO@��,�Q-�W7]�0���0G�VQ(��Õ�U��g1����]j���q+Xm|�q��T��a�e�($��#��h��ތ�{��f��� q+��;���eLE��e�9K�q�K�É�_�dc�����*��^���(��5 ������7���x]���<n�x�(�'@x8�ŖMpt��=Q�@u�ٴ�F�{��M� ULFڶ��L�J�И���PwGF�A�f� X�|��"i�FG�C��*ΰ����Zg����z�`��u�����*�׿
�����Z�Z+E�`�X�S?�j&�oƌ�)�竤L�;�$�Q^�4]Ύ��[v��S��5�����Sw��+����7�z��[3X�
;���}Y^�w�D��� ��*V���9�m8P�<���2lg�Bgpx����-�����(�~���Q>�05m��0���2' �F��l{+pB��K&*��u����^����fg���p`��!�-�I���(w�2ݟ�E%�*詃~	�H�Xk�)$�x�1D_�%z�^��Ni�T_K����J���I�&͝���UxQ{l�{.��1�����yeM�����0	���	Ό|(�HZ@�Mb����Uٔ�������H|����/�U��#"߄�hK�^9ޝ�\0��܎ăӝ |�X����!R��gBE����i��F^���|��X�'�^��ߴ^���!��_�(_0_���
UQ�8K7����_O�������36��O1��]������ׯ��"RH�Sq��5�A���r������jZ��_�i��Įb���Rm�sK�I��y)Ȍ�&��BJq��e��oh#�$���k�G�Zr����|8��Qͻ5I��ة@�Lɳ��N�ӝ�Z�X�j9��4�,�XOV�T� �+ᇳ��ZS-ų�Zu"����a(��S.�V.�:�����o�BL{z�ȤG�B=L6���y�Q7d7�8�i<t�b��2���D8r7 s�#��	[��0��4�?!�.�.�x�:K:��wS��58�/g���o�b�\�&.�D���I�ׁSF�_��M�Ou��p�1�a�YP"��H���l��K��T��+'�*�/��N7���7�j��H��7C�.|"'��j�<�Y����p��Q(0��h!p���6�V��@�>A�ufL��=/G����d�i3��n�E� �A_2�x}�!P[ύWʦ�RNc���Nq����Ơ��fӖ�O��Ǐ(�i��VU������ˇluU!W�&ha~ډ�|�?���6�����x���A�_�1o�-�i�$�2
 ��M$�E��J�iCM�}��O��f��T�衮�W�S�m1ƃL�:��y�ɵῇʽҠͯv	��/1��uLRQ3�ܼ+���âXl��{C�ݖ~(��D^�Ij��+� |2Ød�k�ߴ�B�^V,��0�=���;��?��i[��E/�}�50LJ�ZI�g��C��<������C�kC����臚�=�u�\ˀb T�B�N�������g��k���zP�.Yҕ�ʆOjۄ��(�x��b�Әd���Lk�Sdƪb�M�]�}3�_[�?C5�ϟff�	ǋ��`4u�wJA2-�~���ow�R6?hq�� f��7d�&�aڟOB���~#��ep���;}k�A[~b�
�B�s��^^d�'h�����#ooY�hK��	Cg�T�ݫ��9�����̀��|���f��Ix�).vI���M 1�h�]�h��i��@F�X�I ����ِ7O�Xag��EGگN��2��ᨳ4��>�S��7#��&o��=���h�8�;D��(".	P���IK��<��t=WVE3�tٞ�](�W�Y*�P�{��C8 ��<ڰ������Tw���@Ѽ�̍���4Z�?;�ˇ�)�0�/x�Ԏ�n0��O�S�-�����㧡��v]ޖ�U�MK�Պ۴y������L��Ú/�~GI	����Y�LJ��gc�5�� �c�,���CAF�����<u�%)\�C	���K� ���M$-�F��@1�׹klz�֩rY��u��k5�h3и���~�ߔ0݂� ���2zŕ"g:�m��z���f�?���^�1-Ǽ)i�/��w����8�eK��ϕ0�D�a7�YJO��іaAz��4d9 �*�k��x^9�� �XI�)p���Cӗ�Sƾ����v�^�B��	@	�޹Y�.\M�XZ����D�!�ͨ�H�U�i�ݦ�u��՝�V�������(��W��ŭ�*�nڃ�7�;��U	�������@��j����אT8�=I~���I���H^����w�f)Zb�������3��0x@��{�0�y�!�,W�;G���t�6�h~��k1k��@�_�Ry��v���6k�ڧ;��!��ق�w��DWpG:^V��o��hS����h�?m��e\�g?{��6���G/�B��Y�d���sd��s�췱��s�C3/�!*��a7��[���!�������Z90��=+���M��EՅ>�H&Nt�kui0�ML�r�|�ͣ.�	�TO0��|7�{������z�p0{�����r�lmH���<9�Qn�>��U��B|�	�
R����x��y�\x�[���0/G�~̥[�Ir�W�/��.୬Y�-]�����&��9P9�Oͳ��|{Z�H-w	��gx���m+o�� ���#�%_��kҔ��"��S*��Ѱ;�D���8V+{�}2�g����l�FF�G�$�?`}�.~;�^�@�@-��>�~rV�D���C#) ��eCc�ʴ�#d����ێlb$5}��`��3,���#���~F�X��h0���{O��,�\�a�{vh���i0@���B�d�/#�E K���
����"
��e-Gnڡ�~���S��6��o�������~q�b�}ѧ+Ģޝ	}���������'?Ǳ,��(�V��j�@�ަ�,�ۤ|�;�q�KB�i�E�=�#Ǹ�{��m�֜=���*ʂ��2�Tַ(�͓�܏�+�V�r��?�Z�7�A��W���# ,L�����*	`}J֖���[}P�[��	 �xc4��勘� �\�Nה��h�f�88t�@�@��}�O�m���'4U�qN�TL^>��C�R�dD