��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]N���!�XR���դ��oL^�8���m����T�&���t�Tj5�Q��W�Jߢ��A��XYbDD��B��v;�9����`�%�� I_9�2��Q��p���J�{��U4��v����6��6�ؾ*����h�\է����q�>��V�F#��֫ ��ґ�V+�7�s߬N���2>�4���۝��a��TxbkU��k����~d� Q�n�.�K�-Eֺ.�U*l�[�zv��Dt@'����/�`���)�"�T��K�`hR�jC��}���$�m=�x�/\���5n ��f�Vj" _3��%�e����P�sB�����,'n���T�J�RHz#c����M���+���5��B8��C�8����e�81�ms�u����+e�b#����T2ի.~�q��� ��a3X#�?�E_ML�4+���C%R�����V&�p�=.�Lo�&TׁH�`�i�Tg�iz�r��C�
�R[�N�� ���q3$��]���_^�2�~B���uR�\�ʓE��=��|J���>ռ`�9ʽ�E.�'�Y�ѡ�Nj�-B�ݩ<V�`���Lp���ӵ��{�p�v�`�OՁ�:r�\�r���v�E�o�3�Wi�ب�H!�/�� �|��n穯S���׵�wa��Q� �ܶ1_$�mH���ةZ��"��)6͡�Jٓ.V2��UgO��a�RrT�U��a��ƅ��0��!��p��(�&��V{�����4?�OK��{vKD��)�$�!�v ���ǳ�k��A�Wy届g�H�Akw6^�P��i�
�� �hn�ؤ���N�''��|cFȼ��$��;�Nc����u�z�/�5:L�',���#�%v��lg�"�,�k�PE��/u�t��Ը�����t�������C�dߢ]����_��jo#WS�+�ׯP�������R�oӁa���8��ƎK�"U�nЬ�b�]ᓟ��Y�$ܞ���3��"0u� I()�S� ;r���I�p�L��';#��VV*m[#A���MI%�"4�Y�s�H��cO �H�q���w%����}6	$���hv�w����I�DP4.�����B��2�i���*���~U���/'z����?Cޕ�s<?��O�7�n?w�� �r�����
�s�����6*�'���C�+o;ye7�>�Op"��uR�������Ma=e�zc�Q����Ϡ	˦I��D��匸�c��u*�aCx������}�8�n.܉���6_����G�bNj(�[biޚv���D�7D��!Ʃ�֞�7��(k��y�9r�ī��U5W����R2�����E|Ġ�案��u��͘a�)~�쏽���Qȱ:�*Ϥ�j�)��� �{���{ц��d��Hj��S��>�P�D^Q��Df���s'��2�L��m�ۮ���В�N�	1���m��L9d�ƥ(U/�-��"i+���a�bʐ�jH�/H%uZl[Ԣ~»�x�U�a����K��i���2�T�w�Kt6u���,jĩ����)�@��[7&}�6�q[��[%�r|s�Bg����C���w��-�W�Зf�A[�ڑ���#h�,Ee��bzw_ב�]�64u.^�iV��&Of@��},jht�ϊ�Z��V�w�WV��5k`�X�l��p҉B����N�����&{�w8��ǚ�����.}ň��=9�0�,��K�.��%��I�7�|�A#�<SKK������r>6�"�*�݌-6f�?��(�4m� 9��&'��P��ہ�mR�X!J�
�o�4���l�~�[�/����L�Tw7�f�W<1B;"4�~�����t~6Er)Ts(��?p
#c]��>+�y'�O�ʗ�g�i��R.�����q~���9�Э}Z��ɏ)�'�r'�:u3�1��\�$��A��a��wr�7M
�f?���zj�X�5D+^-tj�h��Ѓ)�̅w���[����{kU��:0I�K4 ��@e��x�)��s��`�B'�&5�7��>0 L~؁�0YZ�2�E�_^� j���޲�M	�G�'w�&�aڭ�7��'-���N&1���-����~��K�ǐ�%�>�!��0�g�
k��d'�YqR�.idB�N�5�ӧ�S��;_S�jN'�)I��������7^w0�q�D����t�g��k
 �%?����Q	O�ī|���e��8�],K#�:�ħ�S筺�/���`���Q�����[T�F�^��l�z���3�#V�o����;��j,�I�����>{���׀�������u`qp����X��$t%t[��%(���v q��\eJoڎ͎�O��g�����U��sx˯�G��a2�x� [P�Z>XkCOȈdB�E.I4o�9�<q��^$\&�k��7��f��i���Y��t�y���-"a�Ml�����[uŘu�["kJ��b��Y���,��btx6c[$�&	�N�[(����4���:�\����6�o���e�́г9%m�B
 YW�*���&�i��X֝�pV��q�T�#�*e%��vY�t^X�&n��<	�˖ߋ��y�|�$�̎x!�C�s2�Y]�a>���=��
{P�L����/9�,�Αۖc\ЕU�S���x ŧ?HЌ����=M>��&9\�;d�1씈����fZ�g��<��  y���:��|mO�g�J��L�
t�#���aq����:��o�._&~�FT��`���܅>��9@�$1���8E(�9�8�����C!�گd��u]�8��L5c��Z۬IU���q��H�O.c�������Ϊ40W#�����];�$�l򓁌_�
��>;���At�"f��-8�{(�pQg]�Eac�5�
=�Ǝ�e��)�d�ϴ�"̶ߗg$lU��(F�ư�01�B)'�Q��|��L���\
W��V9�g�Ջ�\�AT����fDU{+c�h���<g,ӻ�����M���j�/1mYԇ
`�����y�>f<�~��X�h&4B��Jmu���nCn�_k5D�s��h���t+���2GyI*�����9TO�1�n��R�̈́�h�d�������8l���%�����
����#m�Zb�_�S_���ر�/K�����zB��n�1/��\{��Ub��!�N鼇����#�Ү(5�`�w���2�8����H�=%���oBS1��pl�a['\�r���?|QGPI/1Y������*U�-R�geA*��0��43���H�1q";Mc�ϵ�P*%�T+�) *Je��1�s��W�%�0ĥ�~gcNT��"��,�#�A�����zge�5�ވ���DH�qO6�nK~�R��M1�F��SQ�~�+L�L�S����E�O��CW���撮�Y1���0�Y�c�ߐ���o@��dH�EE5E� -��Փ��/�\��fsx��F�lW��u�{
\S$?D�iKWF��+�EUX��������/dn2�9�eg��Ⅷ9/Vbb�}�t'�nQ����9��i��F�0���@���E����:wo�Z�eI��;S�Uo����F0�dU��(���\��d��W"���m��$	��x�����p�|��{��Ķ��ŃVK�-���56�6��V��0}��]�W"3|�?��zW'*���1c8oS�Y�{V�O�����G ����`X2"��ê��/�	#g���E�p[�/|����7i���D�n�OP��c��'�c[i�kj�@�1�ɤQ�<��;*2�i`�
P�S�ѐ���J���+�]��9�����9yO��gϟ���ҁu��5a�/e=5�B	[`Uq����s��[���ՄaQ��4'�Ar���i;�ǒ"*�h��M�H���p�Lv桘3tk�2 ��d<������K|�:	�H���{ew�Hm�G��ٹ�5L���!5�fڞ���^�_��R��U\r̠�2ZSF���Ĵf���b&��9���tLG��.��V-��H�}�F�I��d~ܰ_��^xJ@�`9�8��@,���-J�6��7��L�(���sbǽ[B�Q��5q=��s��!7������SJt�-�*�77N�mڏ^L�x��yՒ�j�s(k��_b�%>EJ�F��n9H��Lz��#�~L�<>K�J-�<�༘~i�	&$��R-�!*P��f�ny@7���"���+F.�w���<e��c���٠ڄe�{�zH�p�?�:��Нƛ����;&�|�v\���iE��I��Gjj�0sWW�(�W�g���x�Z�H�ڱ֎�Q=?w�J��v���s	�P��榨3k^v�#:��rُ��v�%,�>���~�[���cf�w?Mx.hQyj�v)�:O�L�1_,�0�V�)��1C����%����;��ҵ���+Lm���� !U�K�-XPC�,�te{����n����Y���k����������O�Y��]�w������-�xM(����T�� 1��**��Ǝ�Ĩ��(��,���dm��aڼ��Q��[�SڗO�hn��ʖ��E�j[~�q��?�=�	~��u�e';�0���
V9zNL}Q����V"��ߘ�6@#��R;�	��Ł����I%K��Z�SL{}�s��kl�3��d�ܧ��H���8�/�,E?�d�nWvX�Β�i�o	��dN�=��B:"������O�:\�����YXF��x�Q�]�f��Vu*8-���1�+^ߧ��'��4��ݾ�DrZ(\on�,{|�m�-��x�O�&^�z�0eY���=��{C��b�I�V����_����n���>��ԃd2���nU**AA����.�Ы)fwM^z�V}Io��\ۢA�C��:���̓w��T��ka*��?��=�\�hx��Y�o7����SI��OM膮���sa�B���8/S�����c@�@��ֻ���ݥLPXt}�n_#_b�Àl8q��9v̅s��Oi
kݨ���BAS@�� �냢��S�&�aM�7;(�J*q��)S�.�ڴ1+��X����v��/�"i5d��'�l��+?amI��c{x3b�d���|�.��7I@�l���!m>g�.�4��M��s>��y�+�Q�
�)�X/�s�4�}�u+>e%$.�)��E�0��1AЄ���5
�'������V�]��\j�O�ah�3�^wt����3����ޫ��1�z�sL*�OF��̑�Q����Ľ���j���V$ސm�x�b�#���e޸s
���l���,u�:X��d�ӌb�;��ڤ����U	qPZ���O�.7���ւ>knt0'J�j�-Ofnޏ�՟i<���ʹ��φW&_2&���	~@�R���QY@�2�w�I/1��3��z	�Ȣ
�s�]F�)V�M�\����;��[�f�6'7#/_ۼ�t ���(��\�����"�Y
��)йX��MZ�x �>%��N�ʽ��.��GE�Y�6���<tƩH*˷<��g�q�
NV�4����x�u`8?�`J ���5N�Wt͏�����%Nn��ylv�A�5�*�������΄V��"�7Fy_�s��u�Md%Q2Q���u��$/;@ P=�-~��<��:^��k�p�P3�"��o%�� ����e��XX�`tsϐ;̪������������x���g*�eK�Ǒ�]��W�f|���i�A�*�T��uYr�ʐ1�צ]A�����z��͜���c��7�*D֕�j@h<��?���p�	Cs��$n��F�d���O~n�v`^u3@ ��`�⦉2���QⶈE�3���YZ�X�	`�����ϝ]��������%��S�M� �.�O��m��
���/ ��3��W¾%e���"�����ӑ���I�5���o�ϊ'c~�G��ҢbOIA��p�7M҄G��B�������R������>8.W�!�zJ>0���K�x�����9(f�����˴��̎�x7�#�ɭ*F���SO��,�Vn������Hdg淧��{w��|�л��u�9ȈI�|sh�Ԟ�c��=�ti�1�m�E�c6<�s��vݲO�����򑐱��<��c�&r��5Nȃm�<��Z1�o���<xkf��l �U�m�ݢ�[��@�}������.���w��x|�QnA^A0\pZs���y+�ݒ��x�3�|��X:[r;�y�/<�XL9gD��F�v�Jv͢yY�k�-1����#���I����f&e~��,ʻ.]���H�-fn��̝���63�(Qc����b�/��0�sY�-�u�1)��N�Sf0�*�9)7���n�*��U�� ���)~�$v��6jՌ�����Ӗ oY���<ٴ)�}<���bP)�^��ή����j�-Ǻ���1>���'���������hM�z*��č�t��I	Ǳܝ<�f7s� ��J��i�Ɍ3�u�F�b<�Xٟ�ge���`V1zk�m6#��J(��JX
!��)���TCԖW܊��h����H���I:�A�jCxz�-"	������y�죋�saa�9rSd!#�� 8O}�K/��e4�K`{~4(�u�"��p�}� ��`� ������n����Z�_��ƭ����D�K�j�����pz�-u�naR��6T��J�����~Y�A�{V��������%y�+��-\Z�;m��G�kaV<7U���MqH50b|�.��(�+���O�5|X+(�^҅�lC�kl�C�uW�M�����3�Q4�|���������Z��n�aU̽V6q0Qv����߂�C�	=�VO{I�**,=����	a���� �����P ���Hu�%;s�"�6��1)zY�|8��4�$��0 ��9/_V������p���M�ls�[�/�O��pB��T%�m�ZC��s�^D��d���ńA[�0���%�x�P"s�ɽ��B�R����6J����e�x�7p9.��uA䨟q&��o6�w��:����$��L	��S/��Ⱥ��|��H%�3�1���UFQ�d���)��C,Y���pX?"�U�N�q��-*/�t�F�0�:��jv�@"�0?�S_�)x0�NL	�]�Ԩ��s*o�Ee���r�L�>��S#����RST쀿1M3�!s��:d�' ��t�����l����,Ҍ4�X��{�5$� �<O�>%/������wH=~ �%�Ï�͋sĜ�ۤ�ʢx�R�ҟ�$�HL��`H�a�m���z�/x�9D��a˙�	E��S��ڲ�\H<�-r�n���w��I�c�Z^1���W�$Cw����a=�x{�����UgU?�ɺA���̝�a�'Y��b���Ҋ(��P��A�|�eNӟk�_��ṱ1wƾ�й�w�ҕ3xx���M�vBk�Q�9I<֟�˴x`����!E_�OU��m����s�-�/�L?mED�7>�v�9�~S�ݖv������.@H��yG�ep�a�OX^�Q�}~x�h@�.�3�K��}_E.lO��"~<��	�zC���|��0bB��t�*1�Ƌ��h�pY�TJwf�'�����N�����0�b������/h�M��fm�d�Y=�/�;�*b���~"PԐ �7�Z���7����SK�}ܸ פ�U��w`�&N^�ꫯ��;�J�Vk(���6a�p�&����	Z	W0��H�E^�O��|b)x��k�������u�������OwS���_
#�`�[�?^��-��lY����y�*�9� ��*jK�M��-��"�>��To�;-��(0\vTg�q�����R�3�熔+>�,a��G�/�I�~�X�.ݤѝ��P��_�������0�I��)�y x��N.������́��s�~6c&G��q���S�H*�N����p��)է�v�ݬ�u���zĂs#��u�p7U(JmQ|�Wt�P�?D6�ik}�#�V
�!�N�N(��8��s-8�3�=�������Ӄ,0�II�{L^&79�:6m@���~��r,c�U�`{��������4^q���Gt�%m�6i׌Ϧ���^jcϹ�dAb��'�~V,�yq�	��_��l�R�'*V�^���� 4C�.!6��9����WW�U�I��`У�#���ۈ���1x,v"���Q��g��UW��1N�0��T�7-yf��ƪ��h����c�|��u�ˤ_�)�����(s�n��"�{s���
�r�:_���2):׌�x��b�2�䜨��x��x�x��_�����s�ЏG3�*�����TU�Heoc)���Cp�����E�Y�-�胏��e���k*�m���xl�P
\~Vv�
K��I_��J邃�@�W�&�B&��~���7j,��דcG߈� �{Ln��HFj���l\�w��}0�4�@�-|�=L,��m�c�m���E��i�p��Q�!�w
��{Uo�i��s�g5#�z��hp���T�m#-?��&�� 	u���sb��K+��a(p���[M���&v>3r`p�vO��%I'�r����W��<���d�\�ԫ+$ĞP�v:cT�� G���/h�MҚ�7����-y�J�����Ԇ�����)���6�AF�����"� ��6���64���@`Y���G�*5֐�d�~�p�$�ʺ�WA�*Nj�.�J����$K��YaH#E����X�@�}��ET�c#Q,���H�
踛K��|6v5���S�fb����Q����[�Z��(6�	K?A`S~8�Y��n�thUJ<��me�Pld�0t�
v�.(�4@I��ȯ��	'�H#O�������-����]��4�����4%ˎ��u^��ӫ��|�ng\�| �pV=�/�Q�������j	jp�!�/����8F{G]!<�⇻�җ�A�[���fX��������.����A{H�H}$K(��1�)X��t�uy�0�-U ?���]�c� J��H;����q�u���Wn����5_�����"
o�U��9�U�p����'3��^B?uX���x�� *��d����y*i�������L�X�52��2��uq3��s�:�$^�ǬbU!��(E��Ń|	��<�
jt Q �k�e!7�^`�\�����Sh��,{�L*�uN��ɧHx��ni#�0/|��U�˻��41����^�hq�js��Y����XE0,������)��:����j2�	�a?�`�t����](��O����+��IR�ʽR�i�1\�#X��v��M����`
�>H�,�	�-���j�������iu�e<�V�`�*7��)� ��ۋ��@��l���B���w�O�Z���|�̌͞
�k*��&U���>�J���(8���!g�bg�x?9�[W[�
Q|�V`H�c�⸠����Z�$9�2��{��i�ɸ$"�ȃe45И��]b�{F��==@`�%��� �uZظ_�D����!�J�V<�ω%�tC��L� |�R�p��\�|��;q�@��εw��˻���/�?���I%��{\=8�m(�	���FP�Q��l�'�"s��T[�����Kv�	�%�x�^��C>���Vw2.!�F X��h����<5��5ڕy�pc���[��I�_9��gC��"�xA���?-�0����YH!�l�&��Q��C���d�&Pe����!�mC5�Sp�7�S%m�3�)�6�ߥ'śGC��W�e��2�_h���.kʙ�L%K��sd��ҋG2E��d��a�U���*Y�J�J=w$=*�7�k�l�o���y׊��C[�Yo��?�b�EcW�&s$#��ف;�_��.Ɗ�+�o���~%�]F�&IR|���<7ƾN�x�C'�9�z���m{HъK��=�N���X���z��������B�PٿX1R,�
�,Z�J�	�:�s�C���]�g;	V&-t�]�P�g��О5/Q\ ��Y�d��N��[�z��+
�u�!-0�l)���cV��mpJ�����2�_�LbH}]�-�j/ۺ��e��x���^�,�A[���e�P���lnA���p�ꛊ 嵳��LlKn�ͧ�I�cqӄ␢϶��.��ڈn�\�''ؿ�=�'6�&�B��|˧W���z��	��!Uċ�[7�-k­�~��Dץc߄���A��$|X����<��G��Y��(#v��X��X	�b�9��Jc�ڎ��yAֈ�m�A����J��fN��$�lz�nGa����i�m��Խ������j���ZX��0K4:��Y��V��b������zǛ./�tB\ގ `����e}a�"�ب��W��b�����pẉ�Z����Z5-2Ȕ�m���%������������8�JSv�R)-�hc�/�!��3�{�ɠ�k�{������{�g6㵳��F�J�H���%���σ�K_~>�Cɂq��he�bB��pE^���m�-����7hT�l�1�V�{ad�8S15���[j�-7{Ng�N�.��]qa�S��l��xl0t���
4l���+��8�o���ܘA"�{�:��;X�՚���yp��8�[�����|�7o����tq8h��Ui�F[�C]!��`h�U�#(i���#/���'������Z�K+�~����]¼�M��P�מ�R�d�D�O�;(m:d�Z`vST���3�G��L.�C���x��� 'P��hɣ00��[�(`���p�-��];W'ž�$�#���E��d��C�,�k.�z�w9�/�AW��5��@�Jܦ��O�[�i��B�-/ր����1 ��/�J�1`���닲�t���a�v�,D�a_OG(\��b�t�fL����㲳���-i�Fy��	�`ȷ�!�Yo#���]mceQp��
�JA��y,	�r��Ƕ�G"��V�H��z͌cm��(zD��%j��b#�������V8��7���pPR_�� `D.�1�E}I ?#�_Yə���Û�V#/�r��lҕXR���a�A��L8H�3K�@�F��,�/���	.$i���F�b[�ȋ���O�S��Z���H=	9RE��^3���hՅ�L����Mp��ε0�d�����2�)��ᾷ�d���\!z^+�|�Q,���O���/�m��?��E����|�Ysh	����ǎ��b�]�'��mfJi�� ��Nl��K��O�"V D�î�r��\��sv��0���oy�����O��jS����Qz����xi2�N�f�/�8�����!�c1\G��	��G"&�vßr}N�Oܓ��y�h�M�����.�8=(I.NWY�� ������bG-�%�2����ށ�
�s�14}�S�t�I5�W���-�	7G�MC�v�2���g�MJ�ɗkBvp�lݎ��o�D�9c��܎���¾<f��Ȧ�أk�Zc�]|�-���m�f2��#O{����`w��{jRm��O��y�_��^�v|�Y�^?��ymSQ�]r��e�/�>Y��8�G�Zh���32��p�BH��MA��oQ�,mf��(u���o��		֛oi4�J�����xQM� u�3#�J:����Y�-��A��|;[!إ��|���`'T���U�(�<
O��f����Z�]�`43kIU^��W<��*��f��`����iSs�]R��E��[���Q������*���ua�N��������9.MZ��0qQ|��0��n=%1ݭ�"N�S$�jc�94C�Q��#��ut�Au�4Y�T�;�M�:%������9~��,���U��^[t��� �������؄��-��ݨN���������Cd+�
ĵ������p����0%/���rMO�C}B0��=���Q��T�Fׁi�Opv�0t@���s�!�U��;.R��b��"�k~��AO��xn��8�� ��ҟvD��A/@�O�p���T����l�!˺(Ϣ�XEi��̉(_;��r�us���]�x��l�g����ʷ��[j������_��V�H��+��-I����ȳh�i%������-�/!!��&ۯy�?�s�rs��iJ^Zܽ��i�S�>���m�p�ɇ>��S�
Vr��Y�l���'�{�t3�Ci
��vq�S�A�\]�˙�q���s��!-�i��i['5H��钟�(���&A},���-sشB]k�9�ab���c4G{��5ڟm��o\g��a7!�z���lbw�p����� d_z!?c�[#�+U����yˌ��-f�h�*]�6ؒ펵��N!���h�>���ʘƹuz��Ϭl_/=; �������x�x���Qt*n�ѩYnuާz�s���F���lM���g�z�M�,8ɏ��Ӟ�y���*]`��iĨ	�bp%1u�3�Jӌ���u���O�b>tjC�Lx�r���Z��\j���./��EƟj� �$W��ܪ}�xf������"�y_tGW�b��$ѧ�B2�7qu\�S�D��ަEW�;�He
��س�+�Ղ�#Q�N���G�6݇��U���x��["������;�fi�f�K�[����j��l\.Ud��_��M�u@�U�s�9�׶��h��^c�g�=���}AV^����H/�FP��8�z]�Ã��V�7��!,m.�Yޅ��O
2�G����G��y��>0�kFm��B�����s<�	Q8�З�Vt�����7ha������	l۱~���F	��XiIq�+;}#��ؾԿ��@Z`�xo�����5$㠁 �R�#���a�6cH��S��஝�6r�:9C�}�U�+BŖ �i��R˙�=6ޜ����ʀ����;!���'���3�E�����W9}ܾ����d�ɾ~��Q��C�ׁ�\�N�?O�[?��lEܻZ�nq�/e�/Əġ7k?��gJL/�{�p�).J ��b�H�Fs-�M�!X�pv�L4��7�2��Yv�[z	k[@��FM��wy�Yy�Q6���0�FW�Y!)ô��	З��`~Q������!;\�%�����^����\�!�nu޶6��W`]O9y�l�Ş;U�k�/��IGͪX�E�p�p6o��ͤ���ll��v�jA��5�Օ�,FZ���D���R�y$��]5$���r%$#Xм�����~��;� ���v�I%DΙ:��-F��$"�2ذZ-S� 7e����H 5�5�A�m�_�K�W�������̏݇q��*��*B�cx�G;Ҕ�o�v��7+S���U	1���Z�/�c������i�}|S�	z�]e�s+lO0�=�i��+{��;��}�v&�[���!��=E�� ��*��R�Y�������2p"�:�U���ۯ;�X��;�4�fç�$:g\�4�
��9L�&z~+Kq`cM��^%�mNWꢟ��P�O���˷_2�z��$�-�T��(��k������x�R�h��|��tG�6(8`�~�i���˶�f!=�	9N�H[ώN�]�$&J��9��/��O+f�Q�?�G'h1�xhF�ulB���xW@��e\����A�c�aքSP���A�V��f�\v��A�=��(�.\i�>�)��o�Ä$�9#<�I�o����%y���)U���K�\0L�{m�Ev�Ps�]ur!��Sz���m�!�\�^N�~��<gcgǐ0�S��S�S���/;؈�/%��ò��s���m�|�K�ŨvO�P,�/�R�^��,hJ��
�"�~eā�!	�
G]�!A��L9��#U�cћ���N𼹘	��P���y�ƀ���-��n�O�>�R�wW�;��4�gM��}OBۅ��T8*Շ����N�RʋڥXQ�����	=F��f���E�L��G�@�Vy�������,zT?o}{�U������{C�~:��=7B�Rȭ5��Ƣ��c�����a�����^������^��ڱ��V;0$�	key�o�kr#h8-L[j���]��x]y��>1�74O�cj�Pk<��?�� �,��|R��%�f��=j��Ys�xY:Dod��݊$6�K���j�S�"�y����6ţ�	�:��7Pe�&�n2;�������>�aߜ�^>��	�w�kx��#��~e97�����D���*1�}���p���ƺ�f"�cH�N(6�1��Eo��"&6I�[��r�!��?�5|�A�9�[���㴷��k��&?���o���$ɛ��*�Rm�K��7x��[��n�ؕ\��&C0gf����� ;:�mu�������늏D�� ���j����2B�ok,Z��8eq�%������5��$lw��6��=@L��*!Lc]T����;/����:x���|�M�V�����$$#�f��8B[3S}��]\�Xf����ځ`�7��ʱ�\��xsuе�D�M%xS����k�%�Q���6~�� f��D|�C����{�3���1�!4+���@��G=�5�L ���𧲶R��itR�r�ǅ��v�}g�*!\`�ы_�|^i��)�H��1�����§��Bt���Y��L-�X%*��u�:lhc��`Ct�!`C��5�Q��r;t��B Ϲ���?F�+�	t���M���w��+������NX�>*������qT�����`�V
��Ra��aAyq��}�!��(�y��F��!,B=�M2�{�7�n&�c(M�EqV�#+�wjȯ˗4�T��v�s'�М�{�=mS'��}ȡU�qER1�����$=An�Ԝ��0�a�	���s�T~�đF�a1\��ϩ`�0�����B��h�P��v�m���Z�f�?�ͅ��:��%������!�A}K7I��b���ż�,3Ƚaa�s˪ή��L�=���~�ڑz�~o������Y�^хe���^_W�-�U�j��Ec �˕�o�,�v���]B���H-,i�±�L�����R�R��J���S5�C�)�w×{�����D���R瀷��fX=���҇��]U/ �z���
4�Ý��x�g�Ql�OT�I�,���q(���c�~����)�Y)S��w�D�//��f��USc
�LQ]��H�����r�0b��`2o�0ˍ� UMW�z�R��=�����L���LQ_���R���M^F�!����9��sad����=�[`�V9�ˊ�f?���Pz�y��Q�%���3��Ŵ��a�1F0d�~�窍jKa]�K��5�WG�[tpn��Sy��s3C~W-�����x	a��[�ӿCOP�,=ELȳG��-�D
=�a��#@'��/�^Z����Y�$�=����Ŋ���2Rh1`STf([��u�M���1�+���b���g���A���w�&d^��։�~��z�	����"��z?���!g�o�7��"��M��Y3���M~�H���,D*�S�*.i��D���h�
띮(#8��
��z�q����Ɩ��w��\�zH���o�4�����%���>^V�3:o�A�������c�ޓ@
���FY�m�k�p��\ZL���M1�~w.�'��Ox���B�qkV��ש��U���Y�VP
��i�a����7I�o[@Re;����eΝ���刪��_�;V���	�N\7>�ne�?z˱8�Ӱ~�k�x "/L�������/�Q2������Ye8���G}��*�Ф�Y �	C��Y�C����uyW�u]��&���Dgɺ�����ms��Poi����W���q�