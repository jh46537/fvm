��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i��e�EHM�O�ｱ	v��V��a�"��l
<<b��~L�v�S�l��J�b�`$n�	���u�'B�:?2��� /������k\�4�H-�Ϊ�ԝ*o�ռ|:�1�]9l�������P�q�x?��~Ij�ukS��O���ף���ל�����<��?�,�#��ʫ�o�f}������b�)��3��zx�'0�b�L����_u��R*��}z�`�9NR�o#�/x�kK�Mg��sST��p�<��8�ܠ�M���cl��+;��V 9;�<��u�^�gV&�|Wγ�g��/���vB�C�����+���� Vځ��I�_ ��~�["5�>�bol~ˆ�
��A$�ʐ���`�!�R|IVQ�7��� �>�k�9|< <�i<A�,�C� �V��)KA6���؁&}��ee�Z�$�i��L\Tn]�u>�N���?��*e��VYL�_��Kֳ�/�Z.�ѵ`� 	K��&�֨Z#��B�s�����Zj���c�!�²��s���i�ԥ���a�Ɣ����?�yw���>�_�%.�j��t�@73r
il��/[ 4� WQ
"�s�V9�{��\���؍a��_�{h5�/6�t���;�i7J��6���҈k�� '�����*EE�>��z?�^��� f+L�I�x1?����9�ڿ]sN6�$ڭ�ۧ�=��&�fO���$�Ȧ��`b�I*fS��� i��%k��yH8PBi�4�o�\�vj����n�
��궂lѢ�M�pfN�7�����ϱέ�׽��_U3*%�n<�*�E�zuU�n7;p�]�:�{�h�g������UX�\UY�L��v�d��6P�/*[[$FW^i�g|����w �~�ѹ<�)��'�%h�0��4���>�E����˼�^��{�aB�.�>�a�>�L��W��W:7Nw�����ya�f�k��;�0��DgpJױ���rz���Zt�̄>����� #��@�P���_�� ���Y��s�����=��L'��_���L3 ��c٘����q��!l.[àRv�{���l�|��(��{4�a���	 ma,.n���o�)����坰~M����ރ)�)ۑ�� O0�G �@�7nf�<�����(�o�룗q劐��,���>u�s/���0������z�S%�:Rp50Y5>^�TQ"��n�si����R��J�iՍ�LD��E}[��{��Y����r�x��媴�F��K����"��������̄��C��ȣ�&<�����{��ޫ-����	�>аG�d����3�� j+���d·�^^ݳ�ȷ���!�[���m��gC�gQw"r-E���R��?E����﹈}D�I)�g�y	�;r�����K��$������h�v�?����׎P�z:���rY�l�2����������!.Z8����Y�'t@a���6�xJ>YH�0�z�0z{{Y@�����~�#����(=��������]o��*֍���n���o�����I�VҸ�bVX���#%Ů��<����۝\!���&�7\��ok����wxk�l�:
�oԮ\��NdT8Y�W(N���&�:/̥��]�[�y�T�?�> �z�e��,�К��4ddoa#۸׊� �ENb��*��
/�"w_��#��*䜇sN���dHL�}�kM��&�
��渏0��EX z��^��X&���y�� f#k�p �Ԑ��D�7�����:�"*W.�yf����A-�	�����ň��90>���g��M����I�#�h�n5m®������mU�����	Zj��4?���T\�h������3}��/^���
�%m�F`�f�rQ&�u�D$��ה>����>��������%��o�m��x���+�>]��)%��NΥ�5�'1$�"�~���l�����`Xվ��d4��6.K3�f��t�1E��f�����8�$��>�2'������ɺW��X�b�����8Ɂ�N��c��ReV&���ȇ��c�#�e��2ۏz���i!�-��������O=	�mפ�F��^�{9O��<���l}gd�-"h���=O,���Nu�Y�&^>��Ё�O0����T�����7�l�N�U���Y>�G�C`z�3[W(y@9��K�(㖲h�u���X�`V-�nr�����q#ݾ�׽�|���Fj��"���6s���dJ������ҿ{G����w>��a�VhLY1�����a?rX����W���0�^ef�:�����Z���ܭt�iA�@w�&B<	�c�,���;Wܛh���_��Q�P)Zov���y�rZ������DŋQ�<�ų�� �`��K�"{��z��T��aطx\Y���}b[�b/s���U�꾻�o�/H�$�N����38}���0� �ϼ��K*ؾp���� [��F��h��Z0�B>��Ff��o�f!e��̀��N*]��'����	��/j��ۑ�wX���֣�3v����-���L){Έ|��p��ە^NW��a ��M���-Kڥ���������`\Xp�ORov�'��#�%
��G
�j�;�d���[�4ǿ���bEد��(%w�"��a�d3|�3�}@��m]׾�!Γ2���rwي̬Lc[�Z��*���s%Q[��/�^pGv��1L����Ƀ-x��+��s7����hZ�R���:����<���u���+@8Y������ʲ��'9�!mj�2��e�>!dޕ8<��^0��_�q�>�y���N�u- �	q���,����~���RjL&��È��B�,�����y}�7Ʉ#n�w
������UhW�IP���P겪�}q9jC���X����s?���-Lж;!�,<ߩ��"[�Qas��
'>��=�s�Q��h~E�����Y8���"y��� �ub���Br�`[��ib	�h�۠fx
�����`%8)���&yMeHB##'��2����E���!�R����0��������|hD��D���ĺ,ܑ棾��G����6��ߞu1����(y{�x������'Te����<�ǅ�끺�AL���笒���n�ܲ�J�j"b��� NHgJ�GŻ&J�x3o䡫r�s��C�F��`H�Ue��{�#pK�F!N,V���FϿ�:���6���s��X��9��E��@~�Ƀ�ՙ_����2Gvvd��� ��;��'n�����Je��4`�uA���6?#2��L����m%8)��Õ��d�hC�$:,��A%^��ijHu�~�~^J6�r�@ z�aqӺ{6`���
�z)�&Q�z�qh���;p����J��R����C+���yb^"�r�y��(*k�h~Qd� \�c�
��q�Au����X�;��l#ŘHw�^iq��T׬�Z6��&O��֋�O�?�Ӹ�$�6��Nh��/�S��6�M��9�@�`�]�36�"I���!����Lb�@5�0g업v��l�ٍe(��e*ك˩����}�3������UvMj������f��w����n�a稩�"�e�#Y�l1����G���w����9���.8#�ziP��K��5�f��=ӌJ:�8��z�X=W�u�>��!�I�����i�o��T��� d���LWH���g���Ҹ3�E�(���>�-�hs��篣�dO���G�`A]�
��n#1����Y�')8�ޑ�i�X;D�_�i��<#�ثIʽ<�����c��9�Z�h�g������E-I�S����ĚQb��	�.�$z(��"���:�&��՘Yd)�t�R���z��R�1��h��X;_�'�����&�����?Y�{��0V��!�/��kip��碕�[w[̸�{RS�Ht�U��"��UH��g�Dݸ�d�y��-HJ�2�dV���V�I j6>��U�����	���i����I���GJ^=:�}��M�Q֢�)w�$�Z��+�,}��"�$%ȵ߃W-� ڨ���$( �75��:�����r���1��N��6wO7�$�j���<�;A��b�a~�[Hei�E7��f��B�����e�~ǿ��S� �eo����a5Ř�[���5U��f
�Ѡ�s�S�ƈ�p�Y'�n>:y;ծ�h/B�疴J�b�/�*LiT��辈>y����,,�,;�����g,�h����=�/�)q;��S�G�t��]^WV�I E�G�hP�~�ף��1?�i�",���D��iW�G�8�������>��n~v�Esd����Ö+QA幫�K��AA�w���vP��0q��?Ed��e��!�҃�Qr����i�pI��xI9�/���lA�pr��������&H�a�CÍ����A�"��U2=y�m&-�_���g'�,���!VA&8�I�����؜��.t�$$�@h�[���\���ك/~�Fψ�������>%}��獑�J1u���Ыٛp��if�=vv��Rm����^7j�	�_�	�s�F-��\��P�7�WD3��ݦK��l�e�Z3�e��J>���i��¶���/Vq˵�X�vr��}c �7DBg����T� #!-`��y��#�7֜�&H0��>	���Ojoe��j��(�k���0�u��n�cKB0x휹i<�����]�� �-�Z
+�; �i��j���3�~��箂�K��yjLiw����8�khû倛���c^j�_��ww&^���^][}��(�ޜ�9�VQ��y������B�!�f
�T��-���~�����1S�W�^�?b*��ؾ� 4d�:v�U]`]i.�	�Bh�K���� �hn�:1�a�����h���Y�B���%��ce+h˒/�1�H�����Xb
���.\�~�p�ubf+��A�b���L�Q���ࡴ3ϧ'�0^�_��'bv+����wd(T�e�z�����n� 5�C�-�鷠�MG��)�}E�0D �i��<��G)O߷��������R��F�3'H�N~�gS�pn�څXpV�kT�聛�������nK7�c��*%��uȩp�<{E�)G+�^DA��e%�ڽY
Z��G@&0��"��9Y�m\���)K��f�A���L�k3$?�v^OBYt.�	~��O�����`,�3��^ �3G���X��a��(����輱��a)���kKb�cB�3GH�'2T͏�u��r�#ٶ>��-BMhzy�� d�=*S�A��<HĞ�!�OR�m�8px���Ư�x�������\> r����H���K���͊�r���L�ŉB�@qs��涛��rcy49�Di=�6���Ή4�JBF�.um��0���-n�J�-x�w
륝j���Q!~X���/f���L�f�_��Z�����NW$��V�(5�n�1���-m׈�E�������`&]�-�D�p6o&4A0�C����er�o�	�n�����3(ĭ�X�o+�=~?�ބ��;B��]��Шߕ�rل�
���b������3������Z��R���E�n	g�n{u�f^�g�9�S6xƴS�pD��*�?N3쑑�_?A5[�@j��A>�[�Hw��;���鯍�8i��Ron&N���!Y0>�P�C�(�l|�HO*5�K)���<���1��vG�x�0�i�FY�	O�#��#��S���S�%���t���Xv�^�����f=�A�F�J�k�3X�K���c1q�=��|�P�h�K�	���\�HѠrK�  '#��(���WKĿ�*~n�����ތ���&�x��<����y/�����FsE�[�̐P�s�~b��,L��I,{��v�8��O52`�B�����aR���mh*�&��-�͂G�-����4 �-V��w����[��T�m_����ԏ�Uk��m>VzZ��q���Wo}<��J�*�������Q؀A�Wb>:�M�/��}����}L٤�a�@8��E������"��Hh���h;YZ߰�(
�9�#3hI���e���݇� ��geN^f)������Y_PzOu��Mb4¯�� x�P9}B�8���/������I�Zԟ
�c��b�X�,2�I`�Kr����G������� ����?T(���@�dx���v��ۦK�q�g�X��S��f���كAo��&�j���l]�QЕ^�p�T��;�������a�۴�fË�Ĳz���8�����k�U�pG��}t�e�a���ӛ��ߤ^��O�f5~�Nd��4ao�B�݊���MG�M
Дj����r�B7�jM����,����� S#�8.��M���0z�����Ƕ_�(5��~LG(�1�_����9u���\>-��O�5Ϯ]��d ��{(Z��@��t�RRr�;�9�/WԼJ1�[!��t��-#}��ga|�}f���Fݜ���P�L��R���s�ˊ��S8|Jq�9)�n.�9ψ#�Gd!6a�K��:\���ƚ�J�����;P�d1"ͬ���9�����k�i����F�����&H�+ �>���33=W�]뒀�X���s�A���JwѴ�)��!HQ��pU ۀES�s\&�Ĭ����a��j'��!��cY)	L�O�q
�3�x���t3���V2g�G�8?%�Op;: wLL��la�\tй��'����أ�㊚��W��嘋�H�lg��qV����u(����M$�q-���fܫ��>��p���f�Dg�np�Dg�0��Ρ�(�&^�.{�K�8�i�/�Y�i�Z�FP�aQ?ۜ@B	�zU�?$L�BLע�Zd5d�]^�v�:9R�t�0?��3��i=*�QT�/����c��i!OZg睍.���k��Kc1&M��c^.PY�!�H��&8\���T�]9�2�I���_'P��b.�C_Z�sv/�3���5��PA�s6{3���(�"<k�G̈���h�xm�q��Ϝi�}'0�?<�=�nF;)�Kb�����:���-Q�=� ]|h7=	it�р믢��ks�>nu>,@�c�U�P�.aX後��	=v��t���l/�_�CuS�z��tulxk��Lߡ,B�8>*7�U�d�v�	�pJ��/���4j�E�e.j�W�(��s��M�b�=����ފY��Y�|�]h���1�`֬�+��/���L��H���5��P�H�DtR[��A����������A�
�����oRi�L�E5?R��U�h�l�Āٚ|�
�10��ۍ=ś�c�@�41]ܟt b�,��+�Z�i��������4˗ds{:#�
̩�N��J�<�Y+8���G>��9�i;���L�*�����ݍ�aeӉ鐤�����ǵn�#gki��`)�O�s+�1f�~J�<��o��
��r8S2���Ur�9����f��v Cmy��M��R��{�I�P�)�`s�l-�_~Ê�B,�n��W�>v����C��<�jU�Fc%�@��T�R����t���4���!��".Kh���#���[�f 4=��hwr��u��-kY��;d������*�����T6�|R=�k�i�5ղ!�]�"�Qt��&О+�q+3:]�ժvAQ��c9<ȝ��ϭ��ϵ^�4tnu��@�{M.��t�O*F��U����/�T{���s��ד���:=؜�Ҭx��u-
Cv8�G��I�5@G�rUmѝCe{�J��t�H�{�(V'�@�xϒ�.U�J�����xJ�9w���x
�X�Y�L�)�ୃ���5k�V�r�[;J@|�y���U�����D�}��9eT9'}��O�l[���[ࠨAW]�����QǞz��G����˭'�kW��N@����1it\�'}�S��9i�5�䎖�9��}ؒ�<�w[�m������e)����Ⱥ��D�fiԀ�O. j6�w	a�5]������>ZRg)��+�^s��:D��r��In˅�@�Ny�|
U���^yj���[�k�\Af�L:��LӖe�Z��Q�*坂Pv0�����P�c8�uXuPE���Fy�޷���8�u�p��������=D����GxꈊjnQ�8�3U�����"�}�Q�(6P��U�����C8.�`@�5tK�1"��3�G6��*��޴�P����+�w -��WU��6'�x���t:�Т�c�Cŗ!�R�L�fh��ʥv��M3	=<}0�:����>��eF��S��~?��Lp# V^D�JaHc���Oh��X��]�̔e	j��'��+vH�-$5�}���H�@��z�$l��;@�V/��S��n v�	��$�ee�Ip�*|� �9��5�˳���x"��e�W������ECw����P�u�A������`ГY	���OW� �K��|�OS��g�y�I�.MZ��
��f�M���)��E8�:1+�*T�4J@yw�8x��~�J��0�X������SMbp^��5��:]���:<��JImt�h�Z��5AJ��H҅AcW��$�J�8�bM�0��)m��!���^شy�[�u"���Y�*;Ay������ Cs��9��˘J�k�2��G��j�tt�Q���밟�t���]۸�@C�Z,��f0�%Mҭ͖$t��Z�Z �
�w�	4���*�{�%Ӣ!K���h@tXcRM�e�P�}'�0?�h;Cs!E���^�{_l�kB�fr2�e )��k�����|ɛ#�����<&��旲�oK]C)��� ���rܣ�Ց#.���E-�gSR9�:f�3>��~�H�P����9R�s��
�S�F�N��Ʋ>��kH�P�Ph�2S��y��Y��Y��)���i����=6��8�p��;�㓹23��zće�)�!j��A.����`���B����94�N<����
��/,�Ɖ��U�mM���융��c�t,�Ἀ,t��⦞��t��JSq�Iɂ�yPX���>��|=KZ�y
�Q������Qc�}�O����_�Ǥ�ݮ�C��Z�X��|���d���ÅE�O�B\tQP@��j��R>�+5�B|�#E'���ИqX8�>����c��a
4�mJ�Ӗ�o�:㪖1Cy|�ݘ+���l7�r��A�A�^x�.�> <�#S:�2W/����IyP+��QX ��Cs$��|�t�H��� ��r���<ˌ�x7�r#.��+oX�%�'T�(�%�=9ʺ����L��%mX�ٸ�~@�����:֊V����s�92X�VK�]�r�j�� h��_D��)CԇР�	Ƈp�qƭ٭����P�F�D �t��&��7��N�y��`^����	�>�0t��ը���}�1��_�T&���W����}?7�_���/mRN<C�6�#K�sr��?����t �|jfsKrt� �����GSϨ�:m�njE�ͯ&����ѷJo��ٛ�u���ި�,|�k�^7?e�6)���6�;<��(	cкF�}M����������Q(�>�bȔ<]�ܟ��pLc��{�&t�����ղae�W,�k����ftZ��j�����LIe3�yS�P�U�7�����R��@��}�g;���GB���}H3�����q+�j���MF�5�i�9E�b	h�k��eT��[�Dpa5�ZND�E�T��m$�@�4kP�l��⒤�dvr�%�X�8N;�b�\!����[���g��2�i�)a.M�;�V�H��1خF�c���K	ӏ�+�=�#����}�#`��q�a|(l���;�5J�=��<���K_9G����w��S������`�wN��y۰��%"�U_�Z��%Q�KU�"�ɳ(�2D��ո�3/�dd�+��� rg3PM �o�T��X2�=m*f�a� �//��a�^��W+�M�C��|���y!:�숞�3�����	>b�徳`������)�b�sR���DPE��u^�n���W����H]�UC\͜B�Y��I��A��X�>��+��h���TB�T�O#J,��?��sC��E�B�+��L�eڷ��Ҍ������q*9l� �y�ou��L�D�b$��$d���J�[��s_�{��	��ֈ�F�l|am׌`~D���7�xo������j�6��B|2�)�P7��N�q�{]�S�c�I E��R\m%��Y�y�)���w-�/�
����?d\�C�tCP��o�-�K�����U��V�������EP��c�%��	:���ze���ui%�y�-
�"|"��'`������������}%��ۉ�P�U T臮� |�^I q����7��
��	��_N�ꩼ-4�Og��cE۩���w� �T��VE�����D�?��)W�A��M0c�R���Ϙ�E���/>
gcSۑ�ۘ�|W/YR[�E�ǠM۠Tƶ�7����%o�/�`��u�;��f�35�=CS����`��Fg=h	�-�3'�Qd݇���}�UE�2`��zj�F ���6N�@�/(�'�̌z+/���P q����oS��=�S��k�ic���f�%��Z�'HrTZ�˦��}p�X7ט~�rD���϶[�<hUT҆�v�[<d�j��䞔[)=~���������ȒX�ؤ��-��W:�$9|�ׁ��h�ړ$T�XV'ֵ��V��4-��9Χ��D�h��'��Ù�p�6���{����@
��vīM`��ҥf]�[	e�^uJI&����i:F��Dm�P����xĘ(3�	����L�r��7-`���������w��^��v�5���m)�FNc� /~�~�+⻳| ̳<L9*y�>3 |[��CFiO�+s�4&�֩��,��L8�w�cM��������	�YB�=/�
$=���%@�4�?1E�[��bgJk��A}�d�"J�����C&_{d���+��q��CޛB W�V����-�4��B�G��fM�������b��J ��R�NY�s?J�H_"���C��=e2r�
��d�3G�(�y�EiE�R$�YR���H�7��&���ZJy��#�ԯKlB�4=v�H2O�ܢ�`�@
ـ%~"ß�%+ %����'َ�C�-?[�c�o���e��m�u�cm�_���}����Ik�_Ms���rl�cL�fO���G���J���?�W���v���:h,ڜ8�u[��I6dh�U�I��� H��O*(2��Xad��py��M�w^��'�냻�0�a*\��� ����1���^�[�>f�jڣ~Y*�&���E`L5���x�D���bu���@�j%����
:!̏u���¿F�{X�~w�f'尬3��;�v�L����p����?�\U6���JFa3&��	H�5!_HM&� 0$ފ�V,V�>�x�M{���Bp�Ң�����Eu"*��^	_��qZ�I���:Y�hLt��b�έ5�Z�/�qYy05n�wuM6��O�=��(��[�ub��~��V|8�{_ ��Jg�ŌN��y��',�ǐ���4�tj�r�Ľ2��X /Y��UV-g��Cip���'�Bp�T��b�.9�o"|���)㴸MͻE�5}.選���Ǥ�[��+�<x�D�a���d�k�֤�e���V����^&���d����ʦː�Q���s���_�Z�@����Њ~S5�2|��
�Cl[�g�-26��m7i;To��/�I#�Sd���X����g6�!�mjv�%(M�!�<��a����J��2w����ܫ�L�^[��^��z��%� ���D����Yc5�R8���p��Q̡Ύ3}�]ԖI�ĝؚ��$�����&a�	��/�H����W3��<:"H{p?��IF3���!.�Y/��p��x����Y����$x�Ѷ)�u�M�S�h+����-�`�f�7F�=��Yxh�ˣ��8�5���*&�u��rЈ��,��S�g� n^X��a�K��ɗ��Ad���_p�{�2�t�Zn9��yz�~�uZ_�IO�7���CX7B0�n�Iem �h��C��f�`,�7?s��Z�����]��s5v��6*
��Q����}��j�/�K�B���e^� ����""�S�⛔�I�l ���.��Y^��"ܒ:�9؀87&���*a�E"p�G-��y�)U�{Ft�+�a�1����Uv}�~�<�ؽ��*#")�5�-���"�pC��tW]5A�)c�A'%V[�n���a�m`S�b9�_F���x�e'����37mƧ3��bO����X�nѨҴr�������E-���U��<��۽n�!J��O��F�I�9RƦ(�������+���[E�(xŬ�lU�����a �F��$=<d�Y�4B��X�_-�Օ�����'��#>�� ��Sd2b͊��2#!l=Z.�?�瞇Dߏ�{-߁g�w�
詠q��i�#^��1��p��1�BT�50#NoN��]��;�U;�
�,'N	���R hD�o�f_�.���j����>j��A�I�9|envdTtzG�����{d
���?�2M���`�b���"��uo���~�|4�6!�4O?�`.RT��S��֞ډ�J l�����70+�6���nn��a/V׫�@$�����4$�^k��󱗇w'���F�N??5���CW�@�UC�҆���wI��;��h'�[c%Y4ł^%w�mH.t��oA7@g��?.�Z��h�,<č���i}Wy`��St�!m�w3�i3��%z��E��۲ZZ��J�M��l�J�/)	wY(�]�y�@q� �}vn�rIw��P@s��/?Ao��!rC�K��l�������i8�O5��V���ҡ*���MǞ�-�!V���A�Z.
�!�]H�yg�G����%��<�}��8���+\3��:�n�������q����R1�3ҷE�EfL���H_��b�@��t�waȉd ��M�v�m{�5�K8�!�H �,e��	P�:�>�۞�}~Ȕ�[��VE��k3�����K�a��6��$����TǾ_���v7��q��ǫ}^הWs_U��ߺ�<�3����vO�	{yg��o��W̎�D3�7 ��E�m���;��ɠ<s:g��`�O��v���{����ܔH[���#�
i���%.h�VT��4�)�V������^�U�"�����0�(�r�Q��ֺ�����$OY�`qC����e��������~z���x��K�(9ڹu��f������o �D�6�<w��YN0m|CaJ���P�F �ͼfj�kbcq�\)�Sm�l���Eh꫑S�2!���*4X�و�I.��ģ�����B:g���� �"����2ɇ~����=�6���0mflP�Ԡ8�F�e�w����x�G��{�F��y���A�����y����PG�@�۾��ۋ��e�@�|����-s�J���5_��v�8^���=C�ŀ��P,��<=������m�8�.Z�����T�l����h��%^,������WL4����J=?,OI,������泦�9����?{)de��Ρ0���������q϶�=	Nˋ��)�ܞ� ��gy�� ���Ix261F�B\�`zD2�`�黆A쩠��bc�F:�H~d���l����o�o>[���Vy��qR��y�Fy�4,^b�C!w[�E��Ze���a�BxtW��s�ԏ�2�M��i(���I��,F�P-Z��H�} zR�*���+m5�T!z+�cc�B��~�"E�$O��dB�5�º9-

�ui���3��k�'���5D���Y��烠���a��,kD8��75�AvJϱ٩�{<��6�0Wȑ:~��*��2��t�
���J_k�-L���i�s��<f���nU������"[4����PV����p�Q��e�
�݈XVc�pUv]�x�
A�7��8t��/MQ��gau1#|��M`*ށ�B�W����r�������&[[����zʰ����_-���..��?�(s�\�/Z����l�ZZ��'9����͌_	/������} .�)�\G/���λ���#F�l�h�]eD-��F�߱��s�!у�G>�v�>8���L0�)�5,��� v����v�&([��[�7��݅/ꌢ�jIz�R��T]%��<$��H� ����^3�N�:��Ӧ�7ؒ�� ���d�Q\l)2j/�`����L}ٓ �c���9Ǹ��������m����{�N���acR���J�A��P��u���&&�d�-m<��aa�i�-	����f?eV�8����,�B.����J ����uXj��N7����+�dq���*�+��G����}`��m[�O+KM�1��x��$�/k�D]�P�#�Q���u�,}?KĒY;�p�U����+~3N�
�$W6=�2\�u}��阻��nu��
��33x���u�q��z������L�C�� C��-�bx����Z "ÄS�y�ꖙ���u�C���#�̰����!]w[�88����'!c��t ��50L�8�e�w�w�9tJE��Z�G&�+���ʝ|�S?���\6��t�T?��RS�/;��4�ۿS��)���Eu�@59+�u���6���i�L�.K��a�ޏ�`�	s����./�uq�����%��˩�$����!6��>�����!�3�)�caV���T
n+�t�U�l�5*�َ$PoٴHՋu� |�4.kݙ�)N���2�SuJ����񏬏�3= |�)M����T������G˺p)߁7�`vF��Ҏu�5��-���3��<e���� ��d���inF� �p7H�-�XW2"�p�㎻�EqBj��p��\�#燊B�~f��Q��Êu�����H�N�A2�'�Vy�զ�ݗ��i�g��&vΨ4�$�?��=�H`�#�QK�"+~�Ϊ2le�AW�`�Q�ChV���\v���)�
�*H�i�U��*}�$�O�]j�V�m�s���Q���E?��~��{t���0�gk{���a��S��(���`W�K멠L7aɴ�H�?��'�&��\�]U��5�(O<T��L��h���P�z���;	�2|3�ߔ�j���)�pq˓TxE�ޱ�H�K�m��l��x�X`	�;蜂������FS��Nj�(��(j�Z=
�#�ܘcS�#����ڗO��md:Q������\�W�HE�����n=<#��B+o�6>���Ps����luA :.�P�f�p�M�PyTu3&л�B�/��R��0�"E1?<j��N˲lթ}���V�x5���ք�����9b��QrE1����}��{�O��E��q.'���7
�?Ҕ7�~e��	Z9�a�{�<qc~#[8"�}�GNt�V�����^p�6'S��G���ݙ/��BآC��p�>R"I��0�}�]?��2zBI�e0|8y{32I�J�֨W�:ᎆ�'�;��m�XuII�V�x��)[�����މg2�l���SZE�����Y�ea^�k�xM�	mX����΅�('���bi&��r���[S:Y�� Q���{����5p��hT%8�n�djT��#P��������Ƙ�r����υ�bb������-�H:N���+Z��]O2 �h�^3��h@�.=$���h1��53y4������F[�J�y�h�M�X�M���J}�D+�OCC1z���y?�K9!�N+�s:ï=�nLx�]��#������ьKt����z[C��B����߂��W���Mà"l��e�,ɭ�#��i�Hv= ��52(�b�i�A�^�82J�P��G��G
|�����Ch�͍�����X��ICF*4Vq]��1�>KhG����~*�@]֙�yG��4�5����U��KՋ��k�`�����S�cEy9V�!k�Z�[�M���/�a2�&���sQ(��郕���q3������uJ(�����E�|�Lwi<��7�$��L>.�͠ќĐw���/����Vj6g�$��˛�L�DY��~|�H���^�Rԣ>��^pպn���S�Mr�~K����s>��1f���9.�zpS�F�m�1�L�!;M���g�~�l9�Bo_Tv��gi�V��da���,���5X�#2� @��[��T�I9�Χ+�{�`h&+-�5��|����Q?�HTt]Z8^U�P���N͜[���S��?tx�r.+1�(F��=V�ꭡ���8$
E%� �9#R�]��?���R���.4p�%��[�Fi��~9��o���x%�𣫂�oS�B�����t�:a
��D+cD+���;�n!5m��,���>̩Yi!�J~� 2&{���X^&��r�W-\��\/��|� ����;qF��uV����挩�XT����~��(_wE��YV0�<m�� �B��	Mꦴ���WR"���%.@0W�yQw}�y .#�>%�$<���N-f{��8���Oc�*�y[�c����s+�Gܣ�,��^�8�&ab���*�<�s��VW�5r:�hk���WdA5���B�cHN�x/d�d�B6��k�ɓ��Q�&.���\׽��"��SȪHX��m�s�BL�������xU;M��x�V嚿�M��C��2<�k0��dao?�� �ۍ�2�Ċ����$�&�H�O��+���֪7o�)��/�!�!��/�_���~�"�j	(�+t�]��k�#z~�W���z
�HdO�J�&�9#�}����ns	ZD����mb02�����}�t�S۔�c,Y��Qv�선��E۾�?8�Ϫ\F⏜0��C�T1o;�V������Gt�6���G�$ۡ�����^A]k4S�#em䞡�U,T8�T��7�1����	J��a�Q�-�:�2�b�鴽!H�1P���Dkn�񅏠y�KެTM �7<�:�ƫP�i�Ak����w��Q��b{��4�Q��âJ#����e�cPL_���_��&HE�^�_��K����}6Q�	�[� ��/�Ͱ"�X�ӛz'�nV3]�H?���F�����`\�J��A�ͬ�T?�O���E�R��J��T1�EH������
�u�t�@x�3����g*�X;�r��o���S���	�;���e9�Q�s��O����Z�ń��uF|fqІjf�47=b���ù=�Λ~�ƙ�|[v O�"��f}��s�z�d�L�d�RӆS b����䝝�5n��yĳ�Ü�oP�,��~q,/+��f����
H8�57�-�*,��y�ԭ�о@�YŷC�������,�<⒨�l.�e��r�ܡ����w,��S�s-��f�� k�yx�mS�F�g�8X��w`y�H����U��xB2�?vp���V�8N����m=��c�`�gm^�-ըNHb�Mڻf�*t|�</�G�T����8�������WP�}ܽ80��L��Kq]%�m�;�hN����'���7fc�[�̖�3��
�o�8{&9h��w`1�z�(am0琰>G�_A�ֽA'���.�!�4��Lt�\y���ۭd>��!o��K���/е���Km�3* �t�`��sWH9ڲϊ�t8-�
�p�)(��D�8�g��,]���^CL�6/њ�t�+>�Q�Y"5����9)4"kPv�lS�Z~]����>Ư�>) �����5�$Wl�=�"dD�Z#�Ϋ?����c��
rGfc�1��_ #
4;5���)-EXè���9����i��eHg7���:mPK�Y�|&�������X�����y!��A	�%$�<'�bĀ~6/nD���h�q��BȠ��c��ɟ�J�������Ta���@�Ĉ��:���
��1�kᙇeNa�Tްؔ@�ٌ�g�^p�K5�ڷ[�k���B�����s�!��` `��?m�!˕����]${�v݌�=��8x1��L�:�PTt�I��l��me��b>_����h|��U�J�0��ܷ���N�mD���>5^_�c�?��s���y3c��J�5ƪ(#q.1�B-�!���v�X��޿�YFX9�,cyl�{2�^�\�Cm�䊇�\�kɄ�
�e�����)vJ���'�.���,��|�8�'UeO���ʦ2)j�F9?̞����*1����u�y�>c��InPkj88�F��-:ŵ�C��_h����%��ޚ��&P�s?��rӞ�R�uධ���ސf���|���7�p�~~�ƶ��@|&chW��o_m�9·C�67.;�{��ـ}KNd�k�r�0��"��cA��vM������lK'ܤG9�(��Y�>����_���P�I8"�h��vKr������V�������i���x�Hp�9�iY�7����OL#����K�?�Ҏ�a���hw��Ql���ҀO��f�T�#�4Q�,z�$�@m���4�<S�B�Dh��.'�b�w�S� Q�+j��a��X�dD�*����s���ub�y[ܚ�3{�������6$:���]n"=;��3M�g� ��O��i�2k���)ql��٢
�q ���X�sj|�œ/��%yC\>�Ւn��/��*FH��V;Ä�.vs&�}lʲsEv@s�i�S��Xb��0c�3l睰�͘���m���<�.g��X*q�%'H�)��Z0R�����'0���خ�K�k�l�����+RĊ��F��:��	Yb���1f�����`~�{
�9���EsTO�!� �wJc*c�4#���'d-����1t"����LM�d������-a�ǥl���r$�F0l:Uw�6�)/L�uo��V�W��mJW%�vw����ȖϿ� >��hʛL�������s�BV=�"���`ɻZ����gg��q��� �Q�d�Zq����'�0�}�4���5�Ws^}�M9�Hq�d,��H��������p��FE�*�0k�
s-7ؕ��d_����/"%�w$���������}Y�!��Y�F\b�pe�ӆ��*�ï�%h���Iê��3�����
��у�E靿��L�>���$��O�\�N!
��ѓ��2��O��e����T�x
�8^>F�������[���T����ʽ�T�*|sc.���y�fJ��+@_Яر��
 �g�(����7"I�^��b\�!�XZ� �uLc��E�s�N����X�0i筏{�8�l��Rfy�Z����*O<q]a���-��hN�f��	
����ڈ�T�P�m_m�O��H�@���#�zO �`뫆�.�����jϻ��A��M��[�B�7��q.�dm`Kؒ��r�gti9v�.�M���d>q��my)>b�`>�+wb�+��N\�7���a����~��K� �y
�t��beX*kVP�w����ܼ^��| "��r������&��k�z7s�g�MV~ֳ�s��F�(d��9�sV�՟4�.����$���|���p+�C�Z�����ԕA>�Z�t��?�7e�ô�@Nlr1l�p�q��3�B�,�R1����՝���P
���K� <�>�y��wah\e�*�Q,^mT`7�����M�!|�ڈ�ճ����Y���G�C�ǅ�08|$=�k�+��/�ލ5��剤!��	C�����pn�� >KQS�;{��'��Ó܊�g�m/ҔS��k���V�=�Ⱥ�W�i �OO�&��;2	a��I��7�x'>?Oچ��J0�B\oNr���>�e���g�w*w?ป ��������^"":ʮ��p���� ŀ��;�۸1eՊ(���%b^�`��͙5��
������t�������;WI�����څ)�¬��6��D	rt��sns��o�N��$G:������f���Lk]&t��)�AЛ:u�,@�8��-	!S���ck �J���-!��=1;�hp�zhg�ճܕx6���y~rғ=��qkg�@����7-d���:��܌�U�����Z1��m 	��錛?"!2yJ��'��Nw���hsԏ���ҙ��p��i�]�Fe�Cv��<J��Yh%}AZ�|H@�)�3�W��\է�p��8�/E:��4�a��ĺ�������[G�I
|`���ۨR��R"#�H��gn��f$��7��M��[��V�en �駤�?��zв�ʗ�$��\�9���Z��="�w"�ey7�;�т�X�0�$���2�����B,^�*���vu��RǼ�\a��N�x@:@U�S~3�s��>$rz�f.!>��F|������0&��~�����}�� ՟FreVEs+)v�`�/��Q�8[V�^W�b��@�������\��{�^�_�?�m�W���`�NL��R�%~���\h#�S����i��O����Yg]��+�YCR7�J�SWM�L�c��ͱߤ�E�z[y���9S�0�\ϟ��ϛ_/���
�S�g���lt��������(�v������\�6JD׭A<Լ-.��.3-�"����ɏ��"R�1v I57c�o�"����n$�˝w��[1���ts%�	~��ە�ͼ�5u�]۸(�SG��B-�\�S����0��ts�M@��Б��vL���(�M�i+^\�m��Hr9M3�(iH��H�J)�:ykl�Y�$/:�T����Q�Jd��z8�܃��r��)�ߥhnHL0~�����Þcց���	�l�|�D���t���!�?=�I�j�r�x��q_�tg[P���?�z�9Ԩ	��K�%#f5�Y��@*�,2�ü��{��X��c�qGC������9F~���$�8��v�K��³~?��B��21�~��ӭ��<�5�bz�ǋ�I�� =Pxi4���s��"���ϊ���
�K����<��dl!`����N��7>�N�_�ԲcV8e-�x��=3xc+}�����+7�X�k
c�*O_�@��BO&�F��6nv�d��I�n��A2 ��P��[��ѡqT���씛]�c%N�N�L�н���3�0�ܛmG�0���V�H�Ͻ�����v��4�'�
�!T�RL�= ;���\F�������{ɔ����0�?7����9��
il��q����3�	��`W��ܦI�v熛}�Ѝ3}���� ,k��t��v᠎`��%�p���D�tYk�[�\�nld��ل���c�I��5k�_N�Ds�D�Z�\_RUO��c�~c�dBE[j�]h��Vn�l�}�͒���ބMZy����Ʋ�7�������ݍG����{'�s�o����;�2b�pE��s\3L�$�k���QJ� �i6��{�wr�&LT�}3�V�L�xCB�l��?��	�V��ϴ���c�|��F�G��H�w��Y��8]G-󽈝�8�e4�ޠ�w��梎�~Ĺ߿2i��HӀ�����x��
vW01v5�b�b����C����e�����e�v��yX���f1�S��YS��:ʧ|%'�Qtw���L҆��&��m��n�s~'��v%/�1�|�������ă�ˮL�v�7���]�C��k���=z�oذWg��
�]D`�3'�v��Os9���L7�;�<��p�<�ڥ>	(�D��~�(2<��"�:D\�ǣ+e庍�`+�����4�_(�z�?��Zd��P�R�
��8��x�Մ/�𝡓+�:��3� $���oCg�	F_1��7�OH3n�/?�{ZBbQ=� ����i1ȼpr�yj��u��9S�2�-��^�/G��\=#�`�fǑYs� �{v�����rW	a���OZ1�K$����j�_yR��`N�AQ����+�Bf�\+L�׋.�ܝ�es�\���Ό{M~��ZO�}�ߋ2����{"��I<���.���0�B����];����5�K.y��[D��wL�~�����6����Ģ��*$���>٫���̝۪�������B<<�v�ϵ1ۈ*�\5����0 O���5�
���!ΥV�t:Ȁ	h�Ɖz?�:2�npͽiFhܫ�`���$����؉"*e�Ŏ�*�����#�ʧ
:Q��i����i��84'�C>��tm����[�����v��ɀ_e�@����+Z�,i�m����m�¢�R
��V��n F����r�����2���T�M��>,y^ҙ�m@�Zd�ē��?~G���Gb7�7��/j+pK3|��H
�m�A���=��4���灇�7� QIgx�����|����\�v|f�ê=��z5R����R�s��/�G���o�c����/g������j���_�b�`��HJsў��䐕uL�!�v��&�(�~S��C6�eM��zh�� x�l�������Ϝ�J��	��r�eI�iQk� �o$�.��X��Ea��b����.s߽[Vǃ-Pis���pG�[*�w]sC��׎�|�9#�����fUU�O� �x��^�����4za�2��V+A��q-�ƾ���vR]a)I��t6.N��~	93�1�hN�~�*���0dtT1�h��/��T�P���]
�y����f��o`z�~��*;T8�a�w�� �Ono	e��훼U�9�ER:�>AY������0n�:lE@C�k+��<��=Ț�d #b�"��~[t:�y~���<�z�S���	��4�P�7���~e���^�y�+������E�l�Um}y�z@����?�k�l�$�(�����x��1ꮏ�e@���i-�5
�z2��z�����b���3D��Plt�/Fu�S�yF��Q�Ě�v���-z�;,e+HE&��֣䓉��5-Sy9����N���8�	�-� � ��q��;�@�uR�ۺ���fvs�
�c\�9�VL���qʆ�a�T�V�v�$��Ͻm ��}JNr���tq�/p4�m?�@�Z$][K���dX+�\��0~u}���q��6�1���1QV+)�R�3]��j���`���e������ipMUw -E~	(�6�:��v��2Q�5��d//d��d�|�$S��!�(]��Df�4��.����tJ�&�L�|����1��lswe(�kB٭�~�V����D��V�)�С���9�F�}.b�M2+͵B��MRL�N%��6��W+vޥ�����&K�
�5X.]~|4���:h.�	�yoP��&�}�h�,��M���R�Tfmy�?/.�}��.������f2 �Ǐ�����9��$���Ҳ9�~M Z�  Kj���1K���ֿ����� �(��8�P��,^[RE,1h�t_%�{�e��цIL�lW�z���_���p�v�=>$�uѣ���.A����W��8`�ŧwO@¶y
�a�=8���5�������CAic:�N0k~u�E�F�\�b�$5^ʹ�~p	�p���ٸs�j��л������눎l�o����s��h������C��L˜�_ҌCB"�/2�������,PF��h�뤔+��QB���c�]�0����(둌�m'�3n֒i�EMv�l�W�&�Sٝ��C36@S[�.XW�\)q���樝>T�G�K�4�8U#�_C��#�dQlv���!�<��+,}���Wx����o�Z�:�*�gM��IJ��R��n�*�.�G�x��̱��jCrS+���
S��	ޅ�_�YS��z�{�p��oӄ)�wiQ/0jɝ�&���m�h-}�4��%܍��y�D�����Ҕ��6G�;#H��@�-�2fQ�n22�����U)Wt�<'j�k?��t�� �е/ǝ]4!�����~vm����ln�W G�������z)�M��a�:&p��� y�����5dy'���o�@#�K^؁*!c�}��0� =Oa�"]���\P$$�A��@igN�k�CY"q��- ��n��IE��p(��(�$e2�.�E>����::~O�D7q.B�����0k%>�<��	F�����5�t���cv�A�<��ΧB�E>�r�w�Qvg6_Uehg
^w�릤�Β~m��-���7�2���X�M�B�z|@�5�!w���9#�NXR�e�
��Y�˳ZZ#��lkY�Ԙ*��d�Ym�yK���Ok�5;��M���8�T��')�d���<�s��⩤Ø"<��)����N]�B\;�k�N09�xF��M�IU��jd9B���&��ui���k�m�%B$�2�#����3�􅿱{�y~��k����y(7eN�p���6�C�#�u#���D�Ń����о@2J���).�2�r\pĆ���@z*��?}ѵ�|v�,3ĸ����O8�Z����C�:��n+�-C�����M�i��"Cw��|~�6T�&��
I7-��!���s�x�J<)|l��l���#��$8ky������=:�P��h�t��<$1�Z���pU�L���� �b�J��h���XT��Z��������3��7�ӑ<����T[ج�5׈` g�>אSM_X��6�~��
BxL<��Jk@���{Mc>de�3a�:��K���������O���L�\I�xLǜ��qI�pq�z0���>�Ҍ� �#q����$�(xOʢ��hz�lU�ca�͆�:��7�{���)C�C�iz휒�S��!qw(�d�O����rHc�r��.�}R'�5��"�DFZn9V����&�7�g2"*<]BJ����y:7���	U����O���i@ �g�Be���PP��QqaL(��N�ߥ�V�������k�⺮Q@�+y�1�4�ȘU��	��,+�f	 `���c:u�E��ַګ>3�c�C��T.!Ib-�ԓ�����,+���� p�*�H��$#m����J��Vj�.<;���*t �G�ջ�+T�䦩��gԑEp܏�E�E��q��[��.�UQ��ƷZ�+q5<����v�fR)�����g�"�k׵��0�Ae�OιA��K���A��t��s*�W!%ĘψǍ|k��ZV֭qbNxO��n�qx%|�Yc��mg�{�Ɲ��i�U����܋I^�5�S��koB�	�iѺ�˞3[Q�]]F����4��������?���y��;�i`^�l^���t7�S�@֖��u|4�~ �-.�t�/#`�۲�<:at �2���%�~�٦5�� k�U�\l�<�ַ�=)�� ��������B1�|U<��������iqQ'�6I�7z��짒�p��l�^�{����}z������@Ƌ%C��i+NP||����C3�4�h�fރ;�%��\w�}�W;������(�o�Ә%��2��\6�E�vZ��شO�QB�B��T��C�/�!�</����� ��͂��a�d%��q�Ӂ������׋�Z�(N,)��[�s��2��i,8cO�-1�A�m�*��ʎm͜N��Yڂe��sx�SG	��T���z�#��,'�iF���E���(�O� �@�1��e5 Ɏe�l�X[�l��ŕz+i����#�j���7�Cw�q ��m��`�����c�ڲF��IPk��}ny��{�r��>%�	F��'�2��r�M���kTb��Vi�N���;<|�L���ũ�揔"ax���������
���W�s��"鮾	�ےm�_3Ǭ�h/�@�q
��	��3)� ��4�=!o���t*�<�Vf�i�M����/8���ҧ��V���~&�� l �i�r����ƖŶ�o��kN�4�du�L`x�@�Y�O8&��k���+����K�nTh��ݐ�ܱ�u�P�/���]�:��&���ߚ�4PL�xJN�+L�VƎE�?��l2&��J<Y	?v����Pv�r�2�v�r}렴eH��<�R�fd$�f���}t�h���J}ƛ����5��
� �V}���;eN.<7h"�k�t��C��5m:'��/���%����J�b�-�����U��55�5\���%�`��tI�?�����/Qe����D���5��kի�9ŗ��Y��D����\V�D�t=���%C��*ޒ��� ��x
Jpgh4+*�[�T\�TW�vT��W5��10�$X	۵rwc�PF���M,�P�, Z�qw�q��)G퀁県Z����0������@���&�f0��%f %oZ�����1�3�wy`��gpl���G��ʰߡ��UK�\�b^����;�Dϱƾp>Ŧ�ڕ�3zr�}��1�$y/�9��U^��0��]��[���QQ�����9��S�(�}�I�@��ok �7K"�����.�8���V��n<�*���<i86��~�d�i}$�O&�՛�<�b�{�~�R�L�ȶ������e�М	?cc��&�:�X�ΜD�dJ�\���m��e�.����wQ����V��㭷b��k�ι�:��܃�� �z���;���^�0����f��F�:���IWJ�� }W��i<)˜ ;�6X΃�U :��Y���*f2��1P�,X�}�TU��֜2<�8]�؂��7���G&�,y�eH��͘��� �j5@�ŏ��[ƊBPO� 8� A~��D�.fK.r��������AdY1bl��b��`�y�������7��r����y��}�<?jt���n�Z�jJ�r$��rH�}�������z"}Z�%"��i˦=���?z�o�X�΅A�f±��2y�h-lĩ=��V!bƥ�����/�jꦄ/\,�o��ز6���_�^`����4�C���v���:�`~�h���4x��ç��ܦ�Sw��Kǔ�����q���.{6�F6�#M�w�-������V�u�t.6�ǻ#|Bj��;������$��f�F羃�C%�H6��L0�}m�㕲T%�1�Q��~�å��9�[��k�`|�uw��W'��ϰ9�B���#�����ڗ�\v��4�6��IA���M
*n4�[��Ho\�(Zi���x_K�n��Z�ہe�6��`Z�u&��軞[�^f�	]Q?��-L�`T_'�EC)��}� ����F���?�(��k.?|3��#*~Y��ݢ���ֲ�P��$�#���M���'�f���j���F������)�hL�#Px��&Z����%]��{\�5 9L띧4�)�&��aI� �(�Y��G@�F���`rg�Hi�pK*��S�X�����	�H	���F����RY6���*��Э��Z��α�bVT�_ݽ���p8��P���X�E�"��]�&��]`���\��Ac�^�F@68YШ���S��)IVך��'�z&��p�'~��r�"�Z���Ws�KF�(��`��iw��c���O9M3�.��ϋ�am�LS���R�iɋ��j������EQv�Δ���N9��MP5q-�l�ɭ/y�0"*��U��R&��e���n�Z�I|Q�O��������e�w�̞�~���B$�
$��nF�(Ĉe+PwEӊv�%Z"Á.֤�r����y�e.�@n!�<��5Rɛ�I�фE��KlƢ}ɠ����D:�M?��mߓ�������ot��<g���h_�h����2�E;�M!��O H~K����Il��:�4�C�E��ދKN���b�;8��V��+ש �������	���N:�[Kj�ݐ����������㮽�'#j������� �V>{I��sX�v�#�l���re���(�gĲ�YY�R؆�l�0��~rn�K@Z�f�\��J��s1+u��|�C�}%͕ުmo\�j���6� � ��f���Mc��<kj�N�j`0��ڎ���'�g�)4�?���݃�,�i+GSZ��N�����Q���Sm!i�*# eh��j�C������z�<y{=0ؙ��g�t]�����X�ϐCs�*M�_���7d߱�ߍ���<^���\���lo/"�r����Y�MEh^@4�(hc�A��R��<L�	�C�Ɲ,����ئ�b���Oɡ%[���08��B����:��7WݾFuΜ�qxS:�e���3��ZN(�r^:��Ց	��;���"��s��ȟ�-��͓���p��O<$#Y�$w�u�Y#x44���2��8�ot�m��Y��!�L��CMizIQ�T}�|�E'x&ADu��F:Ǽ)g+~wd[��Q���:�[��7N���$��]�q��P�T��_����0��(���L���Z$��%|ƕ��*+ӏ��F��E���0�8,^[�����,G��4 ���j���i�0Ye�|*L>��:�E�*f�
'h�\�[A�#��
�?{��}}��ӌEN��JvT��0kܡ�&��(��8�Fv�}s�K�G��c�"H����%�7��\�ԩ��GU�S8╭�� `Ky���=y�VԒ�윅�ݽi�*���eSX�q��3�	��%�\5���8���!Hq6.��9��� \����]0Z�� ��{I�׬�	�V�A9���V��+��P�H1������8�ɢ��\�e��l�z��� ����Yܨ��~���.�#@ܹ�A*ܡ�i�f�A�Rf$n���ִ�G!�2\q;�\��r`Q�o�{�e�i�ҬM��m)�8�{��C O��Ah��	�hIޘu����CJ?�����c�ܠ?�L���L��ޘD��vB���*K�^|ϧ��g�g��J�9���|<ڒ����e�%à��58>�n���8�/f�	 ��z#�KDt�a�G�Wz��@�>���u�}��Z���q3  �2�x>�n�֥��|;�=�x���n�Y{�G�Rb���W'Iu�*j���ر�:��tZz���tzY�J����"|���G��!�<ˏ�E̢���O��܅�Ý��Dx)B5.�D���-hৡ
�DIÔ
@�T�h��c��g�C���<[�6�&s�*���?�*+	����>7���*��o�&�r����&�$��3s����2��"���2�"X>2�\:x���y�����I���EM_�������P��#��r�A�6�H�;��{�.���/~d�)���|D�,5�_O�z��Z��sp�
Չ��<�>�^�	�'����?��^[�X��j�����wkn��=+�2qY�^���� ����)��|�|d,�^X�/-4%o�Oq {ź��YJ7�R��蝰V�X��L��KǙRN��C���ť4���r�y���;�O�+�W��S�0�;�������z��@��У�?m���e_����.�K�Al��Tn�rCYX�V�8K�#�/��U���c�Y��Ņ���Ƚq�;�A���5A��q��*ತ����I�.Ӌ@W�(��\EW��In��;p��{۱}b&���im�	��D���v٬��ߔ���f��$'XԒ@C�'G��]K�s>�*A�1]�b��B*7kJ�1�zuD�8H�?%�+�k]��ƜP�c����A���"��
��q����wFN9a50+ê^UפոՃfUlH[��i\���B��M�y5����lҡ����0�@����i����%A�(�oz��7+3|�|�?�:�*N]�� r5 v��>㐸�Vk�dR�����'C}	2<t#����q��xa�P��7{K)>���諭�h,��ϢX�7\�A}\�8�c�%��Z /}G��'K���$�t���Y�ۃ������*�ϳ�$iCW�sƇ�T������1<�/��
���!��p+��]���Z"�
�S�|���77�Zi�%�iɗs���D@���@*�<ô��w���9�@����s�ͣ 1����h�\���ow{1�K�P1h>�n�t�� c@p$�;(5^���;^�,b�sϹ������x ��v ��N��K�F��� t�z��0�HL�2&n�;�a���ZVsR�fNA�*h��If���W�^�DfN$f�Y�:�����9���|���n �OB��>�S9HC��?Ÿ��,ށ�<�H��_�b�X�R(�VL���^Q^�H�nK��L 2%F�����
�ˢ��d���Wxy��ya�˃ӳa�P�x����u��A�QM�~��
�V��NgÈ����T���A�m��bE���ݼ�L�s���� bs�G��/+���
�P�.� �8g�m��ܷ�՗h)�eD!چ/�o��u3m������{�_퐨\�ǬϚ�+g��K=}�/�kT'6�`A?w��ZR�cyu���S�0�F�(�hVcg*�pQ�4�Y�1-�R����M�
}.��񔔞�RM�œ:�5¾���ˊ�<�8� �k&x�Qf.�c� �Ob�B��})�R�lcW�Y��l�T�x�� >U�R4�US:^�ӻ��%�
ğH��1 ɛ��ER[�v��, ����^���w���i_02����7h]0���*�2�a׏5���C�%�D�p��e�����G�P�s�ȳ-l�P	����#x��B�a�S�x�f�x�X����@K �_�bq[A� }k=����*V�f.?4�S��Z-��ݕm�oq��K����U�aW2
WH����I��ľ���&�9޼�)����P��0m$FMK.i�� 51�XF.�Q���U�r��K� ��S��L�kS�m���
�$�o�+&�c?|�fj��D&���,$��,Z�Eɶ�-U|��I݃q.�؊sm/5��9�}�q��8�'��>nЎ���C4~J���o\_CY�W��uݴ���F��t\U/�L�/�q�XUTq�ұ�p�O�"����Ѽ�1/�W~��m��jU*�v~�J�O�Pd��lo���|(�,1�@T�?@,w+K
�}��pm\r��2w��=}�!�	ԋ�s���.i�,Eߌ� 7��Z��:5b�+_��2��A��ܠ̭աX!{͂'���<9�ߔ��L�����z�*���"E��O�(����e3>q�l�����j � ����ĺ����%��������vm��fK�y�W�������+B�A�C"E���g�>38w��?��	z��_���r[oJO�`wGَ̐;��?P�WrEk��D��a֚2�;��:k���St��Aee1!�W�R�p�~�u��|��*�P�=$����NNS��

���YPs�	}��s��֮�.�jH�V�Y)�� �������Gp�&Ҡ�j��(� ���v����6y	Gr�R���2Q  ,�/���5��t�jܚ3�yB�&��{NϠ��L�Ւo�j�NN#k5���㋡�S@���02`k��6-��}��vn�L�gc&2`w�{k��;���us�?B�]k�t,�NM�y��um	_V{�g���Ü(\j��~*;���f�T\��cR�������A��FH�7�����8��e�*��A蠥���0���>�`�!��m�����}����2iu5����	��£T
Zi=T��N�LG�kM{��A��,�.��C��_��Q�*���������0"�`�i���U�P��D�W~�L`��D���;�J��#�M@ei����K0!Y)�z�V�Y@�݉��B��E��rNq�����Y-�9����p���M�a������yC�.�嫭JÁl��TB�Vfz�� 1�4�C����J��9�R����t�ynŔ�h �c�� g5=�L�n�������n%��f���exN���{
��jg�w��uI�36��p-�U;�o}��z�&Q�(�Oۗ��r�-��ޣ1n��� �wAl���G�B���~�k �}ݛ��>�1�o%'����5-�Ad
3!Zʽ]����v��-��ü���y*��Qlzƾ���m��4����ݴ1f��J3��c���@�hd#A�,d��i�%��81,#�5b�W�������"h��L��{B[�a^Y�x��r�fN7_�-&ԅܯ�)�t?�C%,�
�Ê �.꡹@Oǈ�רi�j�]��Q����N�?�~ ��'��� ٬7������`܏��?��\IYy�i^v��.a���5�Q��,���>�J�^]�K� �/��^H�!e~������X,�5	�dL]�斄35�6R�0��[
x[�g3�UP����j����k(��s��8��2X���^/���25?#e��X�uQ�s��
�	*f��;�G��s|��9 v% �0\K�	$�2��3L���͛�ȄV`Ez͞?	�+e��Z1p- Vȏ_��Oӟ�AR�on����n��-t���W�~wIm3-X�W��_!n=�\�>�nAw�Zc��)�B��Q��Ъ
d�~��T�l��gR̃�稨y�����N6#�l0��Id�R�c���.$#�ϫ�CFcu~4tY�Fd�*���WY�@�i�����tH���%9,0�ԓi<؏Ҏ�AOi��@�ȮZ6���1��F�Z�3����#"�%U�䜋�{���&�oXQ���\.{�ɃK�5\��P� �u��*^�^�XU�<�����wMK� ���P�σ1��� %��'��oŎ����������0�[GV|�7���'/�V��%�i��-���M��������:����������D�B=cf��/�/���qU}9���}~lR��UF= X�Y��4=�3����x)��oc�ai�~��Ǥ%���t� 4@*��>\���"��aל sU��[��9zA�w#�k�Eͩ�,��=l���^�N -zd���q��|�y���8-��Ω��>>�]~f9��$T��î8�&�`�S��^��y(�_��h_��h����3~��s̡fl��.�R��↫j�р�{E�
�o��.��"TӖe��v�^���3�`p�LA55a��'�ҥ�%SM�;�	:%��Q�Q�$(�֙�෣A���~�� ���uX�&�m����Q�"���0)���_�d=N}S�v�R�t"� �h�����-\~��/0#���<�y���܍RvV��_Ӷ��͍���p�&�43e��6�$���{jOl����~�~��4b1q��R��*�)cK�t�Q��5�h��c�,�j5)9�^���da��*;5�A��5y]t4#�l�C��L^�h.;��Dz�r�,(Ya�*'�t`�F[��g�sd��g	����`)�!�>�⭐��5����.�40�ibQ�g@�5Kv��bY�$����g�;��ޙ��S~���b@��a�=)��*f��+�1A��X�9ǉaT(��=Y�l�� �$a�$`0Z�]/Z��Kb�~�Q���$Cڣ딡����G�&rG�Z.�&�#M�����ı�*Y�?kS��a2q���<�Ӱ���K��@�Ҵ�M�%��gT��J�K1���A:25
��1U&6�^zs�PwGf��5ʂ̚:���S�/�=K0�ʍ��r�i^2����^���UK�x�����9;2�3zL��뭦���&2�$�u�C��u��s�tm?3жG�E����rR�Z���4Ů+���%vLy%�h;(�C�g�FʰGE}�#7����[��3_0E��Wٜ����v�kи;TU@*[�(���zo��k�+��'�NIj���,�A����^x����-�eW?U=L�fI�jڀ '��!;�|m],����R�KxeBg�J���=|!8('�N���kql٘�=,{Q��M'�
�����==�5��ݕXWu,�jN�"�ڐ]��!�j���_���L��\���T�������4})�Ϊ�1�R �~�^n[!,2����v�񝬱�*�/QE�e0�#��3�Nc�#2�b�T�mE���q���M��q~���K>|����kVc�t���Z�S��� �ꡏ���i��ζ������ߌYpJ����|Lx��Z�?��%�+l��'��ӵpxi�ǻ�2xz�դ��t~�f��x<V�|S{<gt�*4ৢ�~�x��3n��X[; l <g�iO+�,?F�Ё@>�:X�J5:��0��Q�;EY��rX�]�E�ӳӅ���f��M]�8��Am\<������|&��M{~�,����1�⠕��1�o�1��P#�c��h�p�h�Jc����@��������	�@o��²�~��(ї.;�S�7���1{o͖�bU{F��R��jcO9�9�Y\��g�`]�x���<�~��U�a��߈��O������y��o��UB9O����
HEע�u�%p8���Y#�n[�n���J�ĳl�!;[ǩex�����d��6��
2D|�w4D���5%U����I�v����R����A��Aei�Ǔ��]��)��R)����  Y�g�h��o�:�%��e���)HB�e��^q6͎�R!�~l(�C����嶻�MP8e��iZP����>�R^8�p���\���A�_�!h<�1�m��N����O�3��eg(;A��J�>AS���$f���"�kc�	R��Ȩ�<�xiT�)w�i<���t� �v߽vеD┌�W`'�����L�	Н�V�2��y�+�7�.8Wak�3	��n\pK�@6��2X�D�v�+k�y�݌%sT��s+���S>�W0�R3�`�~A2��3��O����n]:T!���5>�}�m�S@����21��K�/�
6�VEL%JvZD~�$:2]�3�n��k�ԭ�i�t��|�\o ���W~�{9��z`c:&�Lz0��'�	��'��d3�����n�����J8�L�h�{�Ϣ���m�s�@�uk7��"���7G!ZmG����}Q$N�����Q�J�C�a��!�-��Jt�j�I��"̢��e׹��E]Yo��5,��\fL�jS�A(���A�
u��J��(�c��QHmi��°x'4��|��m��-���p2[��2��v�����q,U����/9�_!�Ț�����d�}�7���J0�*�3��wm) {i_n�S���eN�&�ҧE'���=ƓaА�Gߐ7�k��{ܫR��K�X`җڝO<�$�D���W�g� �#!4,ַ��(�\��^e�=g�D�GE1�o)��mZ������}�J�+�/��9��`�)d�41g�3+v-�f��+�K�}�@�^�?�Y.�郱z@}��q]d����4˔i���U��E��F�2���*^ВwK�;'y�����[U��MJ_��^<��r�����݅�<e� �S���M�WF})���+Kӣxw��}0��hLŞ[��zx��ihͳ��׫�d#bF|�Fvxҕ��H3����EU�b�ܭ͹HMd���P���Kd�&s���6���lbq��3|��-�MI!|�>I_>��e0����'Eߦ�y���gb/���3����&T�W<}	ۡ�}m���"؟�b�J&ys��g�sǅ��r�
t���|��x= �`����Z�YQ}��A^�Jh�i��`	�<� �� ����8��V[��p��A�xl�@�<o@��}���&x�T �����!�.h�Td�96c�E�<���ȢO�nO��lq�T_u���T>���M$�ާ�L.V�hlwz��O@����g����\�qc�9M�u��It�
ҙ�h5��j-&��L��[����`=4:�'�c�F�t$
�wA������G"-c�R����t��h|��y�-wP��{1�O��77�� �9��{@\�IR��9�v ;6 y�T�S5�˩�s�
�ϩ�6ɾ����� ,�^��S3 �|L�`ސH9���P�Fu�P��6���x�嗨����| �G��$��}9���R~��t	�^a���ƙ�,�ѫj��z��F�Yʞr�<Z��6<�)�g���,��������Н3��g�f�ExcN�/ר_��ɹ��<�����c�0�w�u����V/A�Sk�q/�vʬ&�ęOA��a�j��S$P@sw�|��(U��$����[r�I������ϧY=��ˣz_��5b�y��{I�<��T�P,���(f����ȭ�Nb�e����/˒��}��F�>)2{S�{du{˼��'BT	wB�����hp�O0�w5�R�j*J�g1�5?n�0y�� ��T9^9�nW2{Lgy4��Յ�Q�~�8��$�	��9�y�"�&0���'�ы-� �)�ß�M�O���a�[���o�e���x7^wd3u7��_j"��P�E
 �T	��)������V���l�W�n�$R���K�8�ur�;�}����w����媬��T�k�,��A��*j���D�e�&ϙFh٤�)K�L�f�1I�HV�Q���1G��l�������˿��w���ҘQ\�U�E�9�!� ���Bk�!"��&��CC@5��DJV�u̒=u��Q�pӰ���I�����-��}5����\�2.t��?D�)4��A��RŅ�d�q`��� ���q��2�i����*�@R:�,]O#
eg-�Q*���<4<)��i�C�%���R�Gp�G�S�N�/�xa���������r��J�	��$������e`VFBxM�,��*Bh��Ɵ-�n��(h�dEX�����S!�%�T�4rB�MMguui���CIf`MB��ONx-� ��65�������[�-�w�.R���_��A��BｆC���tLzI�Fè{fH��QW�G���?�f�����.�x����M�$�)�ph4��Y����i�ơ`m�W�s� &O���f4�*��"-ڢB�%�#���L�^���-�CV'>Vw�?��5T�r��4(p�cQ!��ۀ���Ǝ�Q�XK()c�_P���_�V ����S��%���~M��@����>��זA�^(��ca��M�����B�!�����/�$'s���Rd޼���_������%CM�i?��R�N�F]�ɫ���e%��T�����Zƪ�;m�(8s�+�>h�y�w'A�Lg�v�M3-�ME��G�|�J:F���OXFS77�?��޳��d�o�j���˻_1��|��P���1���h�:�d��n���_5i�7��Ǌ���w� /x����mU��*?�����iXp�u��W0�BGxOm���0�򖸪ٙ�����.��"�D
��&�zP1�eQ6�q�M��܎?G��\D�q�����$��^;S������t.�������*�t;�UV��q�3D�'���;+� M�Y���Ԟ�g�d�X�c�3���D�ɹº��E�?wŝ�o�<�t�+[8
�j;����o��P����A�Z��:�0Z`��1����G�G*wٍ|:t@i�	���S�5vW���'שX��|�`�ꀜG!5�g�ϱ��u�ȍ���I�<��C�\�����\	Z�>�{�[�1�Z<쳩�!и8K��?�}4I�q7��p����V��$��Y�wi�ov�ӫWbo�5UN��jnny��eY��΃�%���ۇ/���8�Z�]�0!�ə��c�����Ӟ�0���p��PMtw�`w�mSj�N2o8E~˙jk=aQ$1�E�^�O0�k�:C��L={��&H�R���ȺU���?����١��蹋l���8.脌p̮������ChR!H�	���!ϯ��(o:�MO-��������?���X3�S�Y�i�7��7%͗) e ��'P�MA���3����}��m�l2��Z�4|-���+5���:f?���Öu"čg~�*4{�N�偙?Q�i^v���I���d͞��|{�hG�6l$Uyɏx�ENq�X����k@���*�����]�ߞ׉�!����~_��S)�.���f��5�g�0a�\�[��젣��P�@%�����&!yE�q��
T4��O���R|�p���+tsm���3O�����^5\@Gh�t\b se�3��>$1�����������m��{��T��$��ee�P��/h9� D���K�U�^bW�}B��Y>B�C���p�n�*��a��RY�|P���;N��Es���& �Zh�V�Q	CUBc+��EL�8!�JҊ�h>����_����[��ȣ	b�'tTl���������P�Ck˖�6[r��+�j�]���1��o�Ә?i)���ȍ�4uj� Ӡ\�q�^7�%$�R�1?�R�oV5��a0�>i�a �pސ��5�-��X ��Z{��-�+�Cfw4�$��*8m	�&��t�+�B0�ErD ��q���dY�����B?��M�������֑=!�f�4��[��X]�1�2!��Y�J��W/0�Q**Pt�oGwq(�� ��<[���w��퇉rv�hr�L��x՝�YM�ҳ�B@���p�Tf��B�ez7�9�F���a�\*q*75ŅT,�"�����D�Rj��秌BMI(؍�^X�Y��E{��S����h`F��|±,.-G�e\�g%M봝0 �[`�q�@�ԯS�����*R��
����CJ?��ܮ�C�,S�d�
BHh�8��Is��)&K�����&C����#MM�1����r�r#�_����0 �<�Fںi��1�V��e�I��'��f�צ��"�\������vΗc:�xU�O����^O@�`/M́p�KV���c2��g���� ������01M�&|�K��Jպ�_K H�Cpk�7�MAC�rj�:TE4C?�üjA7�h�1�;P	�������:��G��TE��'1��c�=�G�YT�WA52��[,�Ik�?W�{^J��w��
�����@m0c_$;"H���.�'U��`���q� ����3�C��F�\�z4�.�S���n͊"����-	͐+�o̬`�嶾x��,`�	{taǻ�?3�?�l�UO�Ja��$����l#Wk�Q_�3K�eb��X�O�ŀL���C�|�1�X��S/���FEE�ȳD�s�Ѧ��=��`��1w�t��_�>_��I����_"$�4�w�kwa@M$��ހ��ז�&�p?{��zxW����7��mCt�%�%:�����x��R�=��юa�:�\�I�o�����ܟ����
�Z�k����.V���|M��3����7������9�UR��2�3֥�Һ��W��׍��`BL�Vs������*��1��w =H��ə�- Pߋ"b��ب2{s�=��ݟ\X��ע5����q�����z�����>�p����&uJ�$�4�7�� <�m�+�C.ֶ����$�6"ĪXQ �4���!����͕a�.���^w.O�ڧ� [�Ր�{�b^�z�x�o6�C�u��a�~�ªN�"@H{<>H�)�fWC��q�}-ys#�5gk_�q��H��{���{��Ae��DZ_�7ߛ�juҶ��;����/@fk��!'�!\ �Aȉw�x��E54�Y9z�/̒���ʶTaᔩX�M�LY��u崈DV��p�,M���.��v�w�?Q�8��ݿ���=�F�q�m �t�A������8�n(pv�NI�ֆ_Y\e^���=9�&�/[����"6`|�`�ס����DD_��ydy^!+K?�g�o�2�!a-�����I{RJҜ��%>��1K���qb����0��hol��NA����I�+W�m}&rq3m*ʍk�U�9�3�+N��+�/sB)Nr����Ert�z�-4�N��k���c��gy ���mO|G�3���8��ɔ�C}�Y%�g�f�[`������q��g��n�.��_����#lM�e'�X��������%E
�qS�6l�bBi5M�P�bB#�`u����ґ������x?GGZ�Ӊx��<M+�y���(Mr3oT ��*��*����ȓ�l�*U�l\G<�Mʝ���fR<�(�ꬖEtZjF��v���z��ja3��yG��T�>ÍEt����U��=�r�.���CͼmDȖ�vP�磆�8��9m^��-T�E:~�;����h���s�"�J���_%O4؇n��(Y�(��&��&w�+x�EYyXn
���u�c�Jc̕gh�u쒈���rt���kD02��ݎ.��ue�|�N@��D��{���YH��ԵG���Y 0V�f��7|ܝ�<�s�?9�i�B,��_VE�����@ݾ�����<�ZzA?/H^�u�w�ɪNu��e�b\�T}4�9g�T�@���Bˡ�Lǌ����9��@����n���j���=n�5,��E눞,v0�ʁ0���|�?b�R���(�l��|T>���T�o���Dq��0��@k����O�B�%ƪt#��D(8�������	ѻ"��鉃��C��]d���={�i�鄌�:�FG�j���5%�@�i�e�ZwF#�G?�d?���Q	<J�t�b��ݢ��f��3H��(m�"V
~��(/ F�ǈ�ڙ�&�N�!h�m��JF���z��9\���PmB�b��H�"ֱ�K<���U����w蟍3=oܻP���_$Kq{�[�����{8_����U�X8�w,@U�O��p�[9���}���f�#�"I0$�����C�I}�~�
���}�.D���9������Ç�u�kk���ЭfM�F
��q���8�C<b��`��)T�9�+Gk��ꗾ��}��6���9.Z@�[T_�i�n�ud�ݸ�VV|!o���w9��rh��Z;���ql��m3���Ł���ЮW�.Z��1��i���xM�&��/�=A�[@�S[�~�vam�ʵi�9O�A��q��� g�1 U1W����9/����3�\����Ic���+���C�e���cx%�>�b��A
;F�C�y���iݡ�gw0�>�F��A�wĊ��[���g =��r��-F:_��'�sݸ�+\��l@�}�sn"R����ܔo8��ߍ�oY¯�Zg�4g23"ac���-�h9"�^�顷	�T{��v؅���P��s��3�4�����?Ʃ��_$ԟ�T"�i���i��G����OVK�1S�&�������W�O�ĳ''ZŎR���:��%n�)��חS��=mrO_w9g�2VKxS�@'��%�\>b���U�|c��4>���+�K��ÆI� �W�t��h'\���m�����ը��f�2��kz�\���2��t�9�t=b2-wK�@��m���� *:d��,�6�j|����;i���{a@�J}�xIػ}��b�م��u�u
��! ����m��ޏUOmn��?�^k���G+Ճ+.��g�1r��iT~
b�vn9����^������;��5���"nG��R����0!b�&5��U��c�!�Ck/��ȁ;�D"�,-�w�S�Il��;y��tf�Cy��5��uB�m�o����:Ƅ=*�H�	�L�T0�<M�o�B����E#X���툆�����>�1���OOr��Ԍ9��
FĈ)Z��t�^N��'���������촩4Z;�Wy�8n��>c`��f#�Ï�S#�4�o�>�˓� �i��{siѺ$�R�?Ҥ璚M�n��X�'������9O?��N�^�PM%V��I٩|J�?���ۆ\)����G�Ͳ��ӷ*�Y��K:��D��G���M8لI�8�#�H�z[�Qיf�U{�6dN��;�`E9����f4�Ņ8�sJI���Y��H����f\�Lh�B���$)�V��P-����_3���zN�����<ܘ�%�b�?���^-@�X�o��Ȯؔ�?Yy���ͷY�fA��j���H���Z�$�D*P�i���)�.>�q���%���5�7�Č��j^�c�<1����Qăhd��kF��غ�����DR]��q���2���]wP�H"����@�Ўe��d�kUa��.��Ny��,T��Q=e�z�ʽ�Z8��E)nZ� �لX���d1���3�\�\(fG�����Q��Z67�YH�E��R6��<��=����
9���2�L,��q8�ι�/de�Ur6�z�ʓb�A P] _+��hF��2�S�Tp�B$M������2�{��pT{�u�.�� �l6P���3���;�1��X���)��^��r�55�</dGM����x�k�:�JLu��؞5(d����nK�/�V��W�Sǋ�#ƚ�<˝��������8��}������Q�n�H)#�U�����[BQ�lǛU�F�9��K�!����5T-;"�f����n)[�aQHx$1�"�E�3"an_�[���p$�u �ƿ�rmZ����%SN��\�l'�ۃ�YO�1IT~"��#�Dlz ��Q�DT��^C+X7��%�d��Y�V�d0�k��ҁ\k�	�}�3��U`���J0�
��G�<��n�����S���LR���:y^����(���hMv�|ja��)Z
iyậ�@,�bd�~�vͤ���:`�4,���&��E�9`G���ڃ9�O`T��&���Fc,:���-��7Ю�~j6{ܤ6�]}�� �S�ȓaT�jH���#� S�C7'�`L�������nB"~�!-��T.AҏM�| Kh��6�'*��+�F�5LO�������}xW�^�(tӶB�wS0��au	0�N�L�O��6�PY����u��")b��*)c��XQ����[W$7v��2�EE�Z��݈�T`)�7���ɧ�6N��<�.*T6���7b#Ic���%'�L���?WP)�~6��"����h`^�M��0X��>u��IY �H�%���~�[�&hw��^ū1� ^�5�&�q8���y�b��췙7ڷ ���B|�u�N��%��a�8�����U?ǟfۑ�P�y��._���3���0ܩ�8�-�g�bf�f�j�n��I������Q�L�~���K����g��? P@<@�nb��������e��M%e~�,��tـo[�D��K�)x|3��V;�\iJ�������B�J�����t�`�z^�i������$ٚ��.(_߷q��H���Q�Sl�o"Fr���"	��S�(����T�o�4&��h�S��d�>�Z�{H�k �x��e��dGǉ��σ64�a��Cu<�h~t.0�g.{a����(�M��!ws�d5Y��p2^>� m�e`T"��,f�G�g\���,�@p�&�b�k�W|:P���^{~K�H��P�X!�׌��a�Ot3�a��Y/ii�03��@�w����:��n`������p�0����3<���{K��ʶ���o_2a���3�}��2)�T� 	}� ���}�%��A2�:Id�)�P<�~_���5|��~
�e������]@zF��O<nvf��m�)�_�+	�]���N@�A4�������ǟc+�E#C�JǋR��Qr/\85b~a��RF�U�l�W(��kbނ�'��T�Y�ȼ��Ƴx�E�n;���Hl)�܀��+?la^B}�l�.��hU07mq�\���j;N�Ľ�	X�jsCF>!K�� 8�m��O�,����2�&P��(v�<V�`}��*���������
ӱU xa�V�g��!����2����� �?z�4��qk	�vf*B��I��З�5z�&
�NƆ����J�\(R!���S�~��~U���;�~������DR���f�`�ta8ڜ���a=�`�`]b�����XMԖ0��#K���g������-Y��d�����aO�iݵl��t#V�د�Y�b��ɨ^ޏ.�.O&�xV$�|7���<��D�O�nM\~��-��~PI�H�f�{>�Ŝ�%__�lne��{ʜ��x�x*]=�b?��q`$�Y �L� ������=S��?	�������}g���/Bo}��	?�=/LT/��޵�C�XÄ���ػ�$�Qj����w�s�a �����`����Ŝ����p���Jy�8b��]�C�{ʫ�HeM�d���Z6���TÛ<�υ���d�ÃmMT҃0�ۄ�x??��/驂��}���t����z{s�(�]0��~���7�8:���#��Ț��T�ʇc�!Q����W����}��V��o�Y��|�Gs��3�x�����ү�W�n�{���� �C�栃E�<����HO�3�M�����{��t�3��[��щ�i3*�z$#�OK�P�A.PUN�;�w8�ݰOhV�\kˤ�Ł�Tź�%ΰ��'�C?T3,>?��{Ӭn3ć׾+��{% %]�S�3��0�2�D�$�UY�|�2���~�rd��n�_�Ð�@�$�y�o�EU�M�iH���	w)'��p�3���ԕ_�M��9�` !�hj0��J�%��R| ���e�u�"�4ʋ���1�����ɻ�= *��q�o,����P��!��%�!Ǩׅ��#��{Dz����J�:rB��L���L|���ӌ	�	��<�K� c��4��c��s�W!�4索���`u�s�i���vT�t�M�S�S]KM�cAw��yF�Y{��s��K��;#~�p��Q~�ݺs`��TRLň�Eff�%���]L��Lc燮`���Lr7\#�r�t���5��ȏ�}�92?�8K�gYu:r�{K���`Us"ˊ,'�I���&�����#�yOG-��7�E�����i���)�_�oSpn?�K�����[<A���H �Q3Mnk���R��9p��5K�s������ڍ@�}$S:�@5|vDY��L������^��9�2�y�"_3wq|�� Ç���Z�zP��Q���a��]kX�Z�����/�S��Q�G��k��EӱJQ���
$��0�W����{�]X��XWaE��ƨ�la#%PD���k�`0j�3>�͕n���70h0��fE38{��Q�����ܜ���>��n��V/��\��Ոs�J���y�"�1
�` ��O@A��kٖ����!M$������w���Pn���c��w����Y��		
1���.���Q;'��O!Ɖa��C|Հ�� Ͱ�W��X�b�u��n&�/o�z�,.���~��X���D�q�-OܻJ`�������%����g�����Ή�]�J��7��uW����W~� I>��(�����b����s�*�Rk�>왿�S��}��	�=�:A�t��&�>�Q��{��5���!RK%��@^��O�tt�̩g;�=֞c4iw?�ʪ"��P9j�2��n�[�Y��#��D0=��U2����%�tx��o9��=esE/Bn���?2gx��τ�[�O��_*���QU�&�M����f�C�N�xy�z���1$�{��o7�'�;�l�|����Ne�&���@x9��8���v��T/����'z|��n���ֱ�,��G0��]zJ�
�ؼ+��K�	��s�}�$��Jֆ�(YZdf����4��zed䂖�Z����I-��-�&�lt�Nz���`�"��r�<���[�Ƒ����H�#�{�f������x�&o��J�rP͢�#r]|���`�:����>q=��i*��C�S�F{V�F+��y���Z׆บ)C1). U\j���5d�?�PBB1���~�B3��\�5���JK�*!���hFsA��{�.ܲH�����pt�8�&�M�9?�QەC��/��zb�� N�J݁|�����ʛKર��V�mWR�~.1IO]y'HL[b|)�����D�8�7vѪ�,�H���F4����aK0)V�PHY��!5��֥���Ѭ����D�m�����<�V��Iߟ�3�g:�1�4{㹾��'�'����}�s�lڐ�(&���_��y~8�Q��${��.�*0�=jv�3,�L)Seo��<f!��\*�|��e���[��jVp)���5V8��^�w/F�п��DH�Y�I;�R��Z����d!�z��|#��������*��_�!i��S187t,���Y)�P��4(�r�,��ױ��Fj�#ҥJJ�7��!��+]<Jc���g�C����rj���Q{s]�9҈Ҋ�	�2�2f�O��n�R �BԦ��NJ�ь��^�A�
�X���H��%��G2���Ѱ.��V?���4�
\���P{̋����;cg^ZXD䮘2MP�աM,��g�3��z�0뮪��R�|H�a���U�=�H�c"B AL�L�KS�URڻ���]�d��	\�R����s�s����K�rt|x'J�m<�Sw��%Pj����BJ�=9��)����S뗢A@]�q��v�C)b>�a�+	M+yg�|��D�yz�(M�9�f�pl�����l;��u��,�Ul�pg���+��IНIĢh�Q1�
s����|@����niZ��p����_s��Z��g9C��hp$^藷8�Fg�?�0w�D�ͨ���:*n��x�5���cF���@��qM��f�@{��zѠ�S���J1���! ݅"Sx.%����Ho36���P�a�c�s��I��Y<ٜ�����%�h"��̽n9;}���.��e�����ud(�(�#&�����@%�,�ƌ[9`�*"�A��uz�MCb�����	�,��N���y�̛>ȳ@,��m_�Wd��Q ��Q�p��[C�bä(����O�2o�i�X�7q^Jg����Ffy�F�2=�;�_s:��n�b_ǜ��$���g��7���F�����r?��?�5IR���Gr�[�2���k��ؙ���}\O�q��o��xJ�m��k.�4?��8M�Ӟ��ڊ;uy-�bqk0N	9�,��FA5,ι�L`�j�Ϛ������eO�a��D�>"�}��M߽3��7q����e���2wm�R�*�s�ǯ�sP?n�I��&6ϯ�O�ho<_ۜ�Jef�q͕�֟����si����;Ƒ0a�/���]�^r���nY��i
�,�q�'�s~��3�d�U���z������8�6]f*�����
p�#;p��8L��QR=}����X�GYp�i�=�,1�W�a��6��)�a��΀����\C�|�#���E�i6��0�a��"�
J��R�$���) u�8\����Q�|9�;%��Ċ����(��$}���KC$.��sJ ��Ɲ���wP�����]`�F����ЩX�T{��٭�3K�i��u_
�ʷ�khj���ѻ缟�� �������TB��
-4����/���Z� ��E�r��|�{ͼ<�,�*��V���2V��BlE�>?��7���9S���]���3�H�� �d���dc�����mf�-�v���Ȍ��4��
/#�����'�HJf2����ɼ!�[_��<�C��}�L��z�`�3h�RQ