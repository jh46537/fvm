��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�Y֢�08)�	�SX����%�4���l����E٩\�C��?V[,��Wꤦ�}�f���[�V.�Co+��"�Ar�/e�O��\X��kN��>=�(1���?b���v.�4��RΥ��3����n�MvB�^C�`*Bp:Y����E�K�?���n�G��4��7��S]rq�L۶t�D� ��`��!�������t֪^G�o{CH$HM�t(�Vh'TY>6��ن\,��:j��Cެ��A���4�(�7ܨ�i}��Ċ��978(l�e)wqH�H/O<Z��,���PR�(����)�ދ�*
��*���*��,��fowQ�;�?�o��XH�krzW�IF�M��~'�/]hT~�N��6�8��7��3��)mS&ُ���*���N��f($a�\��$�����t������`Tr�X�'��� DK��Nܜx����� �������=ˑ;e�YuLT/�p!��R)�OA$�J��O�_�F�w]9�>U�^��s��ƺ�g�N�?X�M��g��%{f~][iA�z���f2x{���?n/�yw>��3�Bbz�B*^],�»�6�k�Y�qI�4p
�b�1|�	5�J)�0��#�;�3��/��̓��#z,�ǻ�\P";�[�٠J�˒�K��3�x�z����u�J�w.r��p3X��R����65i���H�dE9�u盽(K�п�݅����e���tI�r������[�Q�ib�M��q�[
�'����+���Kw�[�1ѝ7�T �$���&J
��&�:'��[9��*_v��Z�������0xe��%6�B�Rz��k]�K�O�ⵔ��q0�TZ=�1������R�`�R�_��s��9+6@���D��׍��|Qү���֍�пtO������4*W/���0�s�yE@�k Ҍ�|�.|�}���y��!�S2[%cji�� $f��G|7"�@�1�W��lԭ�Gi��ͫX�����G�� �r�`ð;��7v(�(�L�*P�iN��ڕ'4�kr���_f�<�;(l����q��ɳs�T��Q"5RlXR���hS��`sK0@R����_嘹�g�7�\X��h�p�B�f���a"�(�y.�L�Vز�� ��Jz(���R�)h
�n;4�q��WF��"*�X���Ǔ�Z;9,K��7.�8���p	0�z�e�/�{�����6�[�#��g��Uz4�%8�x��M�5�H�A�=C�ց!�%��P#�o���&!{���-��^j)��Y�?F!@0�.����i5��,��JM��k[�<.+����D�~_B���5��V���=�L]�苃��`H��y	����l �̀E?�7S�a�3+S��Wi��RV��ZY_��F��9�;�y^[�tN@cfI#�ּ�m�)���=���a���K�f&����-�߯CH�[rL�p���*!�Wd957ԕ��)L9����\�@;2�yh4_�Zl΀�sI�#|b)��a��|�-�_x���w�S��������-|95��N]��GS��_��pv$�����b�Y�����-}q�#ذ7�|��y�!��b�K}9���ǚ�.�Zp�&���W�5����R�U��=99�T�W+���/S�&�=B$W�H�F��1��C:K�!���V�����4�XQ���Ş/��7o���͹��B_nA�"F�>��t[P�^�'�A�Aw��!~��X����N��Ƌ�C��K�"�wU��A����F�>s�r��[�ކx ��Z�����G^�y�B"G-3�y��$�a�M����tS��Xӥ�j���6R�*I��o�HV���hQ�)�?���]�Lx��9Ѡ+91B�ˈ2^K�I@�%�'��/�t�O��x
��ΚU�d���W���ژ�Cѱ6�Lc1)M+�6}d�n>_H4�H-� :��4�r3���,���f,�*��V�@��?H�@��ۚzTT��P����~��n5g��{�9ظ�a>`������X��|7��J d����+Xm���Y�,i��v����J��>���gN�)$��[s�ڬ��(���}�b]��f;ҭ����G�%Jb�t�e�s6I�Djb8b�Y|U��osItr��_.:��y*U��9}c�F��2���8b<YSd��O}!

�6�c:�f�Ơ>����dF ��8��F�U�k�ڝ��(CO�6�ɹ{�)r�E��X���E�������lVD7~��/����&�>�������?�n�2�V2��g�{��I���x�ͣ���u�$��q^�,�(����mNK�gT4ǘ�$r m���Tt3��E˹9���c�$iy�����GD��Pe� ڒ������a��5�tm�6X k�.��2c#�V���:��\oٳ%�	4��E�M!���t#�_<(�g�0��8�9L��+�h���OV�\Ѵ��;�B�`����Q�*���/�1mc^3���cS�O��u��St0m���:�F$9Qؠ�[�̓�s�=̙Nʼ��;I�d�*`�3F���f�������5̏�F_��C�j�!�r&8b�S^Ŭ�chY�t ��΂zY3ul�W'���<�v=�/��AsGw3\[���u0 ���Ҁ��������bX��JM�W��L�)��5��`�S�qW����H��s�!H�d>���:��дxuT�6u�O����gp�	 �)�8vw�Mm�}d*E�ca�#��A��o C[�L5�Ԡ0��A�2�l���sK�h&)-�Xp��yx�P>��Ȧ���N��6������ɉ!G<�x�i._�S�y�Ѐ�x�6��Ѱ'0��=�Z��Y/����9��~�U�9.e������)"�'�,?)�D��`���A�<�z�z� ��l$R/�%��Pg���2��zH}��~>OC3��r��E�;VJ��o���9�cY�c����8���S�8W��!`�-�z-�����Yd$V�{�)�IF��`�JI��\gi�ܝv,�>Ρ_�uV�|ٷ�iu��� ����1��.r�V��>r^xM�}Q������:��P0}	n�Vt�ʙ:�L6vWG��<��)ow�������D�@t���O6@�7zz�ȳJ��T>�$&� ��g�V��r9�:�������d�$Ӿ�i\�b�R�������>,��� ���^x�Q'����_�*YZ��ms�Mn����q��Vd�I��Ԡ�r6R�lU�:t$��W5i#k)��1���t�jpY�_�:й7�2߫s�ķ�R�LB�S�<ZW�g�Rc�y�ܚ�x�h^[Aw��J�⢚�6�zK�nw��1���2���
������w	-��
m�t얀5��Ύe�;o_�%~V��Nv`��T����Bz�|.5Oa&��V�|�PaE�>\R�h*!&:�	ۨ {����	R|�,j`_�b[òC��K������a�3s:���_À���I�^��r	���4��8��nXa}h-���Ƅk�m�_ef�σ�7�Ӆ���%*�>8W����#���ɦ�5�e��*�B�Pe��W�C���Q����E�	�%.�-�,�E� ��^"� �\E;�>da�r����TN[����QWW�)u��.<q\�L�\�T�ߝa%�Bc����L����.�����h���d��LjO�o��[���s-��0�Jċ�9dp�1f����'։L��?hh��7׷?����/�s��xtػR�8�z��4I�.T��g�`+��&x�'��=���<B����J�-<���T-@<�Ʒf	^�-1�*�U�+m5[�|����C���G�so�[krc�9!*�����t�ޣH>n� ��gy�rw���� ��ۦ����m7��2���V���ڈ�t0�v"�ר�
�n��p�L��r�m�yS:�$�8�M(~���s���_�Q-���|L�}��<�֤l�d���I\�w��H�C��$�
��bٷ��-�3�ܟ�`�N4ͧ��/����[�GR�6d+�E��ߖ/l}Xs��Z�����L@c��^A�?C�U'���Y�d�qB���٩�Gft��ǁ
M_1���4韝/��<FM#e������=�lql�hB>�@D.b�^�G��*���bd�b1K[���{D��?�tu��`Lft� �����A��X-Uq����ds,��C����w��SfA�*��HkC�;�m��z2I�j`�M�Hr�^� ��L�9B�1�V�LBt���f���i����K���r�.wl9$-(vp�7����$�}~kyXXbG�����Y���`�
 ��̺����A��z��>�s�8kHNF{�X6:#��t�o�hq�ao����K�J�w�F���Z�B*�.-q���oZ�Ejݡ�2	b��[�s�'-�		��t32&�2��md�1�s�q6[��GܕP|;���t	I�X2��k%�Eĝl�gQ�d��=����*'$��u�3�7�{��c��H��~�� cr�rZ�W��P�W��,�������=ab�
 ����!��;ii��
+G���d�����y�&]����Y��$02�_`��/�(���l#{aa�w�,��x턍*7��Q�����}� �dy>�{�X��emRq�<9���`ʇ2��@Z3�R�����
^�SM��.i�O��[�H�Ђb��N'�S��q^�
��->8|��*���uk�X#k�����+�0���c�'8�p�B��2|Ud�,�,Օz��/(����W��Q��J�~�{x`�)I��,b�2�������@�"&����Wv[�i�n��W�L�s���k +�+$�^F���X�T�:�'<��%7�#���q��[������b�Zj-�/�/�v�0p���
`ŋs ①��!�,�q@bU̦��W����k~�����1�3����Z�؟|,ɍ��fa� 
��D��mѶ�eU;���sis�%)�cw�g�����;ľ-+���(~��\