// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZoQNCBFvXhwWAo/CBpnAvA7QkTCPzcIE5sMu+B/N+X+H3oY5T8GS9n9HB3t+Yft8
s71zw76xvUGMUdwCxglFDkDtc7o4FKqDhK3+kknj3t1rETyJNmJhzNNtqQhL6fOl
SqaUfAMkshYRT88N2r2I7ur5WLTBrx2Vxqd3ycJFd00=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8896)
6KCQo7i4w1iuEaaD2R3P3iN5C2M8sZF1Vm+RJpcdLyRF518E9RvFR6ydANdnZDvH
g72XR5R81Chl+LpTnUey3IwBuEg/+UE7KxkLERc163ljRnw5T5PADazXTn6qZjVH
cdY+XDHYuwPbQehuIsWmb8sk+o8HHoJ0f6dXLYj6QVq63Z4o2bnLfw034zJfhzyb
Mpol5qVqFHEf8+83v7qxkJKCrusBU6pHImIKCHUHqZoSVI9RcaNR+HAma454qPaO
kOclEbdpSgZ3UgJ9BcAwUzTaJm/Q+V/Miqk7NLyJ0/FLjcYBasK6T7Uuv3CRMsLa
hNU6tZJS1LBDfbIEBykJHJUnjsxVMvCHDTioaqZBMWVZq2aBlrKcYaz24s20qnHC
b35EmdtVc/ZL+ohNZdDzAI/l8o4U8lwdU68ylwwT6FFgDJWcsdkqFBbPQQwzVyhN
KXE5pBzvOztUEMOFOjq2psQrM1ruc7BTtAMypm7WFyFull8N4847Y0mb/e3V9mUS
vJgstvuANFeCpte6ynj1K7h3QB0Ds+6azxz0sEh4qu82F5damJlzYu011dU28AnF
kkOcWUuHtMqQ+jFNAysSOdwKFA5rHjK9ySt4Q5WKTixxwmWR9dW8n3MGRSeYNKMK
pS3gVnxH3Ifnd+i+dDcIzxSX5VQy+eLiXWrRB6oMRQwYWHycKzQH27xnBifDpFQC
Uz9maYvBZY3qG+PFihIFJECAdskikvwI68BufjtmjqjtecWDZAQT0Cd+94CDhhIT
4qgw6mIvDq9fESX5QXkfoyKBY8ppafeH8Ryu4QtfBkw8l3jEwtP7DQTlc39aGpu8
CpattateXLVQLD+1cPfiBssGg8b/N9rFiGm9tmYUbm2Oset47W6hv9jvuhTI0H38
Q4eGW1yDbaxPM/LT0PmB7t6ucUWCtXMJ660+Y/zXRKrrk8lGNRCIkEiUPMgSADAo
AGt0ecHOXsvtp0I1/YWkOJj22QH5HVyCaRszW8W69/J9s0HlSMkqSCmSa71C9Cgn
6+4RxyDewyRHS2L0PcodXwyvtbSvMOsM3lI9spd2i+GZbpsQQA5BXoi5v2NwApxH
7c5klaf3med6+LHPa3DBxMOwVbDqOrzqz1Y5bMRs0kCVilNy3xxeVwKOMx+9AEuk
ESbZnDv3bwGGxWK2ffwH+ccNM1t/nWy+/w/z6QutZQsONwggtPUGcw6gp5tEO2EK
k2gkPs0Vgz7M7VSSLk1sA+B3wnaMVpKVvvDZAJcJa7Se2VQOv0RCsAppswrKFX8E
IdNj+mNgafaMgUAGWxhb3smNAQr9Hqmj171R6Q5BZNgR+zXVJJeK3AvER20EiSNw
TxEag63fNRY8uWIhnRdfiwf4G9l4ZLdOBcEDCwuFbgO+qlNFjGIi7WHvDyb26z9j
mwIa3eIOZHeK2avbYM2Pdx4TnBELU6CJktC2mu9EMLN/gnl83vd+cwc6t9w14CJB
sbUT3H+v6Fs4VSYvImcB1vhq57H0l6jCRgg+pag8VDcWoLVtKZ75qOcCZKFYmWQQ
tF6KPLNn0MEcaOCgJYIHME+nl0300c86WOSAn3ByG+D7TSwZjeG3iQjxrotwa9o+
Xju0Ne/kRgfI6TTCMxsKOzC1vzGHruPAOa4PHadrZ+P/dyDXnVk+Ok2r8geXulyb
0cukDSDyWY/akVnBMubt5Lk//KiQnr2IvZ2bmwEu7hWVWEWsTtbk92U4X2C7BHEj
CfqvcBB2/QazroW/pO7s5Hy4EiHHsZVQ4F2Y7DJA3r6j0GAFRIpV+OKff/mZk38G
txsWQRFfRSFOPCBRoO2waIpG2+35hpptDKSgvoQy+hXc8eqf+1Tz48cGl+t2wSGS
4ZVPFiNcT3yCXRMMa/DX2lWG+DtU0suy7LuHWz1gQOtqxbnAxmeaiJ7/Ye7DWKqK
KtYlrru/7xG6PYxV3GOjg8QGDUQ3lOGSpWJouiWSTqeiZ/t3DpfDAXgf5BchT3Nn
j/AiyitICBmPXvBvdgQUswRemjw6rMXD2MKMLURVG8VoIUCseYH48lG6mEr/UQCG
H4lTFcGsesWpycOW30djJE2w8G7ksBPsQ4g49R57Xaz+DeNuFuvi3JI5dWeXoVH6
uzpNeGg5v3UBFs8X7MrX18hw9RqI/Jh8N4OwdRZCuiu5HFijvBGKhSjTBynZh2C1
1LtGqYOE6wlzJTH64SBqQ+URNaS6grUtWpIiDfMrCB8s2H6kENYiCjrfIWRsWPV0
TA66xRDg0WzQHGLrT/uQQbD2SSOhO7+Sv8tQEpJqk0qhlJpllcV/1o0Jr/fup7mR
skd+lNJbUFoke6oxHbdf9tXis0UhTkZEgbtr9GW4zN17wAoJpOF+WOck5wcdZzkx
TjHdG1HUUTbLOtBEpM5JzFiyG0ndCTocMB3uhnxEC2T+Kywz9CtPOoM0YwngAaek
qbU8g/bNWfUK421lfUZd8RyO2c7upxl+fbLUuzSTDWyNy7U8Qfwl0xU+o8i/l09p
UAsZ1/HKSqknFZOOAMzsSrvXjOp6gLbNHIRwICvPNAO5bFEh92bSzKo1H2C/H8dd
/QFEjCCFtIOfacr7XYLHw4xwcP1wqYGnygMF4G7FtYjRmsPukojgUVZsU0uvGh4H
lFc+4iZV0Sxv23wDjgSPEEYpN5xYreDYW0Lt5CksPc9FTzKMlS6TtBHkFuFQH01v
fBbdja0gQa1Kz57jJUzXHeyXcCaziULRg7ILsgGxqrddv04Ctms58UFYuZvgxetz
//WCrENazOGZr3pBRqT9mBjtSHWyVbG6pf30UcMfObKQXBtA7UMvyTE+ASF6YhWd
TO2nInVm0t/qKfvlb3p2sOiZFNCcfJ8Wl1zbOLRY86iOQAgxNwZaMjhOvqQaljVT
g/TN3rKb3G/etsQwUoSK5TKRAk12kfNxop5NAkYODVwRgUEEyJTMPCAtfH/OJDsJ
1wpB8C+OT9Gg659FqoWKXWFpthwe45N04jXLLKnRLI0gb1iyBlEYztlg0VKxpqjQ
UtfhTqTD6HYAQmf8T2yJN1Ot4diU/aGhoaf2GpwiPOvAMtkRyGE1AXlkfbj/oks5
QZAOC5eKNxx/wEXK9/hBPBSskFj8Rh+nvgIms6fMOkmM6ekafESClfpm/BZVJuZP
ZnIpEl955DuOlznGkqNTg9itknpbNJZkt9WcnTdWz6b+6khe2ne3hNngr950TrYh
JkXKvcNl4vzFqVjfHYIMCjNU+imY3+ASQDyc/UoD2m+p14M7xKSYBRaAGOI9G5Gc
4/v8+nC0S4IFGNQAASG0g6PV2KAYZIaEZCun/QShdwrIuzOvNvRuTJQ1i8IPa0ko
iesGg9W1RZQDv4CQat/RFPoaBkU4n5KG24EZkyQm602ZMtjuFP9CpZlfUgSwckoU
SeNpWsdxv/yk9X6KqHBcgQrkgGEUQS17zlyYSFtEU0+B37GHKnX/xCtDdKLFP0Xb
qAhpBDKfIti5ZXD77iKxamm1bKzlNSsTfprYUqegJbLulJ2Ht7o88P0IkX1eDRTF
WZk0MirR0jKz527BdljGK1FAgLhnvXCUb+RZDpsHwRNR778s9TvRQq1PmupNMjUn
1NCE0W81O+2YC369S1PluJ84Q3rcPsWccFk3UQz6oSnuya72DxoOOr8aKxq20amq
uJE1AXkC+iBm40T24h60n4kfhaBXIayhPW+scbW6lcwZYMCS7ZGzLE6aVUOssGGe
IH8ipt/18lI9lb0rkAD2bDKDX9WangK3tvvv7mzl5Wc1mLc2vxW5SSdIkB0ot/5m
5iZhQnwSs3aDEUJB+RwfCBykTjGy4KyZ20BfDexNvbJmP7333dbe42D3uqfms43r
m1B/0fO0uWvqQArP8JEXB1PNJ0MU3pCz4dwX6zVGM6SdtmVcnVIdqOrPhsWnm9kC
nwtQTUfJP/g79lDjO8FXpLrHFRnT/zwOiR0drEQLPLBg3IvUMvSop2UrNXeM3+ZT
tvia2tjOqCVw03/Le3Yepx3v4Y8eqYxoGy7cw5VkKW5DxkFyEtd/hmdUZUNTjdoc
DI6U+nXuxFgwQnMfs6P6IT1gZpPXnfpdl/HCdzbCoX4m6cSGeSNruzsZUiHVHCrc
Af9T0m47kPAmjIn9G3TzqDH/MfdXzHWAhzfOtY0wbH7/JYivgSez8LMZp/kgRf0g
D72fvMzXdZX8pcPehHyPDOiouuB3lgW9fsm0zLv8Q6x6udedOypEXcpbsLMBxB1F
OntA8eYx0oQqJCl7Acc+olNUG7yjHCc/74z8B88dGhEUFuj5sTa/ISnFpk5kf4NV
AurV/qNPIJGobcZo9h/TVqms+DV6p4YKiQV0K0XBpADVFwmLPN3Cd/gBU0YYp0wF
9NEypT4TyYQoEItPUnGkOZ7NKlJ164TPsEXWnNc+ltRKJcipJXXaDGEM5+v/vXfj
8kH//gVEni4S6ljobE/CTqe49GcHwxMO0euPYrZSydhXBhXF10hETbDrbAJRprSt
81yQ4SeVXbZRt8qPPQ6fJIkt5Q1V1or5zKqDfu0kJJ/Lvvs4awx0q22iwF1K9vP0
gM9ERJ7Ai/ZzPaHxLUVLvAWrgwSuXcgjEvA8zEThUMlhfmCJ+DKaSfTD0yvIZkgX
nLvpi93KYeZSShc8OyWeSfGe+soaKaO3CvXuBtFvV+IX4/xRm9g4so1+kUJmCcRV
zGxCozFVbZJe5jZjjZH9JwZjKlz8y5ua+7fDZeRhIY8zVHpk31/JECywi6o+lbGY
KmywRhTcbyxPEfFDiQBfO/k0g6mAqmzxtUbyNUZGjbWPn/ohxE0DzXAbMVjZENAD
M7mkFOD7z+DJL2puqCs83PUrxVAmmpkHAOAkuwTaoelqiuortruNufXmk73/dG9N
wMv5Iwdw4/t54PlV8u+DaCXne1J59FZzlZeHsozHlPWwkBXMQvzCzy2GkVzLh9L4
hVlYxKn7LT+yZa6bUGtMyD7kgu5/cs3BJhAnsKcG+Pf81HwjfB9u7UxBgro03ny8
l5cwnr11RwFF6KaufK6lJQE79mhh8RYCPlV+DpHWKuuwL7R6T9bf9KsaUaxwZAtC
XsG1uq09gujCR1oQPEFvmm4zWaxqKgmuQBkM49N9rIivL9xd7gprCHYRJFLcojNj
kNrAn5l4y+VC+XSpgvy1rtn0IUVXTjWwQMA1exeAMfCu1ggIOBAq8IvOGtO8LuyZ
c953mynhMWMruzMno6xJfb9p1xEjLupDg2JHpW3TXnpAxLxi/5yXQ/AutGeiocmI
aRUilO6s18Rc3JpUkoA1Fklu0LakdimknxuP1AfKt/xYlOori9yvz9tJXjaWF0h+
bok9sHcWCHqMFuNcbIzA6RSPo4cEKkfd+ExMCeCSDv85GciBgDcvU3rbGzgGCC3W
iOy8Zh7CWZX4BDkUJEDkW6C4TDHokPQjhjBLxW/pIKby+4iEnACFaFhb1k/fMgyM
pFgW7X464Pxl6YEoubXWllpVsQL0WywGTpYfu8iY5aYDhU4ITRicsW/SAYojfAnX
61BtfAwlXmCayUVqjGjoRrYwQdGjJ/hLtub7oCG7K61XaPKCLZPwVmu3XBmQCoTx
mK3SR8ROSOs6YPYCgp0hja+NX75qRSk1aw3/zM6Y9tw0NHG0snjnehTkhzTvIK92
zist/9CAyBUU5b0j88Q3mNPP4zqyP+uDJiA/2KUQdgZucUFa61yzMzG1M3AV8o52
MgGIwrkiKnAxFnBOj5S3/zjVLIGbopIZbtI0M3Zpv+0kmj7KwxLPQkB7fCyy9h08
fNX1TSTUdiKcwi1N5LtsCH3eBD+dzlY+WD02IV6DMkorrIEqvWbsvD1humdEfyQe
auDrj2NwSha9tEiRq4xkwD1WdVm9xLMB88J/pJbv346N+V3m9pMy0Dm7fp5Uizv7
RJvaytGgNFlAQlYXi+vIxz6NTcf6LsfYRBjT43yQu3uCuodVMcWic587YLx4w5Hk
noKs0q2W+qtcvIidEFUTTxIdqQC3gI3RKpx0OR+GW3us+P4TAUiZSrf2ix1ny2yf
XTvu7EzAZaWcox7TDTAa7gVr+uKQTH7AeIc3pB3V4TzdvQy5voJAdxAxdwgPfyOj
OAb3L6MMQleP2nkD4l3kZoiZUM4ISFfj7TAmPVbDwqNMsB62WlAhuVkyzX3m5IT0
LF61ArbmA3gUToS+TNnHUv5bwK0YPe4b47AYo/+lFdV4KCz75XEpFIe2tTBqHRSJ
DcWbraHpRcTzkna83wODUzKBWNobokiAud/Tma5giqFgI+afNNGfAOx//U/Zt6Fp
M68jkRl+bCapypiunowOeeoEC6QusSv/YDEvDfB5tqxlduYCrgsOLjbMtQtC82ot
3Y64expguR9ht79NLUG8KCpovWfQ4vubNxDa/A3KJE831yiRjdtXrG/tL0pIaTQ/
sNNPFns4vxdAmnxRGEr4H6lrKRcPtCGevUkJ6cEuzB2Zyc6HML4yVRRBVwg9tU2e
Nq9cHBalxWay1U6AKjZFze6lMx2F1LOWw5txXESi8H/9VLd/9mEETFH+0gbfpfky
tfafLTxSJY3D+asbYanIYMjVYnaaTFwynj54BlguvkyhkEXq0CwjsS58BqbgDApL
jAuJR9KDklShxzNNPOXqHeMqytjjxH5hTKN/ndMBa1zDYUHNCmpL0/ORip7S5dfY
MilrYN68W9qkjaEl9X0KQQSldCAPqPQNBOiMoQvjWU8tDArPn+/9cKT0G0y/2Ngl
xZF42jesrIKPPofEarJFYnycqz4b+G2kIUVqzAdnLq2nBtYJjvz+v5Grajo753H6
NwRw/yaUIO6UILltPQe+iNDGP/rtPV55EcuH6T7oBj6/I241NwXvW1rwZRviqP8k
vDqIuxahvux8DQl8c8NLhaZcgpuigkND1qQRQ1vJNa+NbdRsyIfU/igoPoeI88wj
mHcYz2FO7dUjdlURUPtuV7IntCHwmKH0ld+LyAA811sa4NOpRyPGnUa0+9HaYvOV
eFHW+k+ioJobkx0aea6/Xhp5MGmoqX5iTAoSwhp/3/0CW1FrCkYb3WZy6XYNN+l1
IV0aJpm+3zA2h2caJU1zJ5DDUSV6ykDqIPLeWRg7AF+kB2e/Wb3Z9NVPPsFeUVm9
mYJ8+iYIpUqijpGD3cQi30jcAHMRUrSplfiT50IkxoyCRgBi9Y3wYVQrEeouhITD
K5AA8upc9NO7WRn/mzVdYyV1Bc9C2zr7eQitacmHK1SHy20y1Mh/DW/T7L0SVFJk
HeSDwJAOnDOgrC2JWpIs0gLXXSHAz4ZJIpeRGOKKok8nyaq3sg0jJDU9NBBIcX/R
tmy7PZ4dZ5oiqomX8TTayDpXGQlN+j3FFCpBkXLSWy4T0tTVF/sQ2ZMJAV9UNs3N
c4kFWGJpPz16hWBCAzULUF1568+DziTZYo1cUId9Tsd0cgilnvGABmTyI/g1696Z
2EhfSdMXdRkmVFfi7VCl9Tm/oDqFGH3xi7ToycerJ5b78suo+ZI782SIUDcm0K2n
a+lEwQ9cwC2SrUDXDYqPUfJUR+RGHWj3oFKS2tpWkXGj8SwipULmFqlF+k3kLdJr
PrdCKnPrE+RzkTzPzENzmRT2GL2N6cVaUC5m1zEtBT8eMPB6+Wg4KJCvIHoVaLXP
8/sXqQbScNJottFETIX1oT5AA1fx9PnORCF0hTiHA+cmimpig5ccQkLRbL4XpxVv
oY4fSZxVW7ItESWeaAvx8oloYs9wGrMu8eyPe5kAobO4Xv1S0bpJvg3A2f/GJvDz
dfY2ljECkH0GE3dXhyh19yQobmwf7AEFQplKi+M+1HPznrlWpNXABwJm5j7sql/Y
XZoqlalXyi0iFEhed2MqvJYYRGZXWGqxxfO0E4IhNU5QZljds6kF6cqfHCF3sIdg
/shjUumRjME6SU/Tvj7kNnx533kK7hFNP2h6xMzQLLdVF80py/3lkx20QceTwjs4
k75IYqfQA9txo7/u1Cisa4r7lbw4VWHhsg8ITebTLM5zTHY9xSqmTMjMglb6RfvE
uGJ4WLuq2iLGbKwIFdy8D+ld4+IW1iqQnwDDZYZGra076SCaVVybrMZItGs3N0lZ
YIIW0V9CwZU/RhONOfocfNskoYxrtPAXklVe4c7tFfuieIxCPVZ3jx89sWuLest+
WUILIRGDMoRYSWgWcTPqH83ofsOCbDK0j4RJlSsQFxtncy7B4rp55YzoqNp9MT4L
r7CCGY5g+DLnvcRZ8BhUrVI9zK+c53ZTNhANV1CvhCKI6mq8goahSr2EY4MT1uCR
0ZpEtgqXlbZ8K8sC1ZJ2v+BiduAnKYCUeiC1qxjlh5zGaPYcfWX4UdQROuIwlcON
HSazMab5UkGVxZxgi3wAPncI90YHI/w1Kv1HyGNfoyj9ky7x48p9RdE1lu9mbg7r
8EQ1+DkPhXLJIj96H+Tj6ftTZ/CivSnb/CQvRVH2R4IRzf5uAVqvVaJXh31ZSkh5
+DVuJo6PqWNPEtho7jG6faVHModw+HARrh85IWm2Jluxr/QIahElrvHAMmV3jxGm
I/mOdoImQGLO/3FL4Mi4LXxrCjzmCdWGN3gVKekXQQ4yoyBNkXLggHsElzPO/PZP
deCHwoOQ2MT+BLDfL2cF1Df6Gp0aTwpoic9fI9W3wcJQtrXl/x1eRy0jl6zOFy8M
2RjJ9qTl7UxtUh1S48QbNZzopA8aJe6yGqLo71DC02VrvtxeFRbFFUzMhIkQMEzz
oAoKv50YbpNhvGfJqWfyygiR7WssUgGoMpO1tJ/5rTDkkBPrbH6lmio3UFB37q02
szVkAQn05quVte9CvHhN2uIx3oPZn/aWdozmh6J3LwWO+NcdzEAdB1npGd9s+/nK
fpyJCI5T1KSdQzVWHIrahHC/jvXe7EqElHYwdWyq0WdAGXI7VaUM+H0iM2fPLoTz
UpN5oOYSAuoThRQhIBXRJQrjPClL9ptw8gzGRdKzW2lLd5cbfx62Qn2foKFKqUor
yYJpWOZ+tjv5On/cIU4lTWpV9+Fyl6WpuwiwVU1bECiTr6yuuHf5V/HfLmpE7mlE
m/q02KvW+9YyLBxZzYDXrnT+I3aEd5gYqmEr86m3LpRCkCRAzjaDltd8iE0yYEW5
Nl6x7pr7ecdfGfDdsPlQOPbQeLDYMLzQnITaIpXdXFbyLmM5LGGOpyNnJZ7YhT4K
JW3w8OWxCDr3bkkw5+LtDDkbpfLH20Hp8vtTVsvdXFm+JmcsLpo8Lf+Ka+NK5HeR
pp+7OCPLughPxSUFpo4TCbCpBMa/wc+mGwbrWJk8zDFaLB0kg/E1lAsEeuexZV5V
lskpIAaFzyNmamzhE30CSRPOD9X5+51K+YOUOt0eC4r9dMZ5xgBL6lfQ8IOkEYHW
wm8RhBrnb3rEau7LzAxTjGsbO3thrS0VUew5WAN3nkc4NtTD8a/Qjj+vcYMgq4yS
7sB5xNX1Rp6KOO8F+0DugNtcxulHhdh6SEwot13P/mC25liGihxD5yeiZ5pFLA6a
z5Kf7OL4sA3gbql67talZoAdepLEtkOi+QtqCxMXBnY5VFpdVdF7XSYvQpPir0i7
tRCRQu6j/AqFDAxUGeZOkBKZnE28UpJPIddjL8r6chUQIMgRDAwpkUJKtG6YMInG
gIbafy4GGKklgwPmUlAT4HE12lMkrq98gab1XR8N+mnhRWrkPE/+FBINJ/dS+6mm
KlSqyr5rfEkr6m+lEFZn7M3wPZZqUv8+SsP/CTPin2V9XAMYD7nIAe3XSNJ2+Qvf
v/5PfvdMbM92zmuqFbEWXsbVtZhhNwp6sF7ZbIwMQq5abLKH5Wjn9uHcnvjRaW2k
NG6epEvCOgAuzPG94VwLrLjuqfVSipDWNV81DCuIcBa8yYtvmcNGG8Jp2watYieG
GHqgNAcqyAqn6VRKnsKAvGB1fC48q7nH8C4nZ50KwiS8tZ1SKlVJRcZciZvNqoe/
AnTU99Cw1FSTFaSkfasytfTHLz/6XTBx7gg60OzjzKHy3aKY4GDjRaLC+eVJWR7B
CFWTdOAmg9oNQKjWRcLb5/qjHIk5l0i28eBVFJ4fvcesWydV3aNfQvmoSn6xQlQw
xn2kJmKwpXHpAOrvk8kn82k3oq0Q3okyA3jVkkbs0NhFdQ3/5olQt1S8sPavqE3F
w+DUKDWa3Vyqc1YhzJI9IsAedmO3nXuHJ2gftNm/2sjMyEcNj7YqsD5AdzB0uQbg
gEcFYCkycnhQncVY67wx3/5iTkcVEBuRcq4ToDIk/9BmXNqqLbNpOaAK67/wFGCY
c+TAkXmDPA9BS4S4+pCewL8UoZRjc4Vy/YTlVAsZ1do8/cME645RIwSoYKD9XhB0
23m9QoC3rUZbsPQdZ9ZyqFZu0Cyjr/69WkG0XfijqBHwCrhq/70u0sKEIo36hOjX
501G8FJHAvHTB0Mifp9zWliN8+gJFsm0KC9X/wZbAj73wgDPVKVHAF0QptW5jAKq
ZdX5Kmc7823iH3ZVgIIWvTxTeIboQu0JBXL9TCQO2C+K9D2zOv8J00H6D5R/mdyU
QeLflduxZhlteivAP8BttL2bygADgCTqr27JLn5j9s8TBZ5o6NMWbFFfqsiCMsSZ
PyJufGyJaH7Pba72ClWVPDZvDandrZUJwFLsx3+uwV8DTkjkD8qMtv3wQd+LgiYf
0DBlJt7PXUWIUrknu3g7KpYG7cQ1/Sc2PhaQmZR8f97WVt4UflHFUT2G5eIZwaD6
ANGT5OXEI+trDLMfmf7YEn3c5IAZdlmlzS4ZEmmEFwGCstsupRDv71wYqxgd9rPR
uhXkHhBOrTk1ME+HEIUr/4YACGJ5t19lNFWLjpDnrrNCqwibu8ixIVdvFbCN1217
GFuYcx5HZ6ib+blnV0Zd1adqDkrQZ6B1eBvzaflN2yYnr0W2I0uMCXvqqdhPJkH8
60YKs2oK3E8JLV8Dc4ujjJdvb5qFOA8f6Gnmj9arlul5sqpCrMuvqftYmGC9Of3E
z2otnMSFbt6ZYx5rF7f3FJMphAWJQIcHybgyVT+I4+3gw7MU7cWzuqsA/c6nQ4X/
XLJzi76QjQKOz59L3l5DiMUu3pkEtYM3Zb823Zzls61kfoTXb1YQBsFt+vDEwDYk
MCRmyklu2kM4xO8vBLzh1psYWBN6OBb4Wi2husmdhelRu16T776jAySfZr+E/S0P
fKeZ2flr53EYEtmCNzRmiJm16RQcewrYASHaTHJSTicpEulZZ2JH/pH409z7PneX
4oXIoWdG9Ceu4quFiROo5Blt/4wvNeoorjyaVc0XdB0VtMWHhcd4+YHmwLHJrYnx
Kz+6ivJqNBHTecisgTYO/m9+aGLouKRCACb0wXShq7tawAYxcpOP1k9vysy9pAWd
5wjnpCmDmkB0XqEBPKDlwa43c4etQ9nqdFhk+f5Itw2Tc0so/FgtsoIwwa37WUQb
VK0T5F/yQBU5J3pZaJIxaCJ0eQip3Ns2XPf8Rzo9YCPh8o9eovFm9X2R133C8MSj
4nN5rKM1/hXHtbX+AlZS2nwwzcU+5ieVp2xBmKnKjARaID4x5+R+J7kR8MP4nkRS
BYp+kxtNnfiEQMX6crzx0D4k5sBWUjeTlygOnfUIEFLvGVJdNPrRJZ7WY6Gp+wRK
l/kwTl2hlsWNdGglh7rMAvtTi7P+MIq0pK9Ru5UBhxbWe9jz2PuSuTX3OxIc0iZg
qxWO5640DYoSg3yeQQdTlsV94ZbppP7tK+s2OvlxH0X8X4kLRjeVjRK6Ev+Cgd5/
8a2jtFJ4wCspp3UKqO9gaj1zaazmzsfiHs5n3LWPTaWQ+ZrNHVTg0dRF7yhknGFt
CD6T3RG9Y2N/fPr/mK3fqXNiffN+PQ9cnfs950yg7fxjCEeQkwAtYbacHa0hX1Kg
XSyFGU/amK3ekg84Ckf+XA==
`pragma protect end_protected
