// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QJxuMpYiJlSwt00PUCvngAfmtLmEqXDayR0Zy+fA8difAAv4Aq3n14hCniDMI6DP
qAYQeP94uzvnvSTylzZqE8y2lwi5mj+mh5A6+vjGq1ym6uxPDuG/tN3x082Hq/zP
g3PBhU/AN1CYrOMi3xMMKMjJ0qfH+UPqq0aiEY2T+Is=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30544)
bS69qgX2juJ9YZU4H9KXTMKe/VxfZjB20nCsLDvJjU+F8mB7NTRVbcmuzjTYOeoO
NHfznpGZQUCPaOFLcUzMZkRbEWXgYZN/LCTGtn/geO2fdzOJwCqQkLesypk08SoU
i589T+vu62u+hG1f5bKuGtAiIyNinVc/gyny2lJCfPCOWvoAJxTIfIHrTJoeA096
I/9JAsYSsKtYk5/GtLYOgdYN2hPvmnVJKLmzVFEqZfAs7qKmsrjakdj5LRl1CBL9
WaHtncMkJoRxADuvGoP45TWV2LfJGWy3B5Vjxn1p4jFa9/6yi841/pFm5e2l6Hvf
EMqfMZgUZS2po6tO6qFtJbEU9wJ1GKVTsxhn2LzJN61CDZHx0bD3mNoh7it8HIki
otA+6rH8ZewTqt8kxDaO3PIAfbK8bHC3T6fo94/gDC+d3xNkpTCMv4i36ACDmBu8
nuGWEkErvjNgp1aSuzLFs6owy00ReFgp7NDBsigt2Lvma+pt/wa+ItAjcLCJCb55
TEed+RK1BGDznoqkWbqCp55FHkqIYh51mGTXMT7rBxB22n7/vwM7JBieabHkKH+9
PwpOWyGWFkC90750bTHfg3S+a0X1O8QAtKQqKbdD6WKimGKzuIeqRbZYPhZshlTH
m08g7ER5jCTXbpev+nfF40N0CVZo3/5brIwNhDtxoGOHlL/Wk5kRDsHBhw47EH/H
OqR5BIkSpAOcO05+yXBdzk+rY/wLd19DWSaPvB8kxp82Gj1TEovmaccCeTbSz3Ij
cjTIvvrepDGZinkRaOot6ZKOetqA81PekU/3UEsQzTQTAzqC/CjamdkfHgbf2XBx
5CFhnW6fQjC9eUHWkSJM/8b/MdpVXImM8sYBWWaFkMB/hnv2Kl/CG2iwDJ+FxFEq
W9VqpwnSFh2Cp0MRxi3wVQ+AeNzGPH/4remuIPPI2U+pKUq+XPtSomqrK4/0wy67
FWTqSvlEH269VdmFzKyMg4Y6S8GW/kDumL2P7jxIGam8Yn98KCiFts7vxPUSe8Dm
68GclQIejAnvDQDENkmKaP13e9fdUCiBZTHB5JlKFzAyQmpl2o0AsygLpDmmt39D
t46VeqlA/2edrKnp/QbnRwpkID8jiplO1NZyexywMv7nOQmGB6s7fZ3Wn4dialqV
LcNhbKJYGKm+eq4PiVmIPrHXkpiCLcAInC1qO8jWTviFl0eqlMIa64uG9VyBEt3j
OCJS3i6bbRQhRm/PplYM4EMsQDkpCS2ZCvMvPFqB8Xwiqdv3C2MoltgizzXvCMF/
EXzyGSVJoQHRuwlyWni+WHqA2LpxuLFmj/JXyZHrd+sXn5lY3p3TtznftBvUP3aU
T4Vvq7s3oeCfbwGv5ZS2r+FtyA/xBOrmxp0eVgXM0UHfhjSxs82+zG6i8KZEUhmk
1QP01rgqeQlsJ0Odp4hWthmtMWiVJt/+QGJEgJ+RmdgIoTzoBAfJxjuOX11K95xr
BUi/FTKraClhN0mzoRcDkRq4XY0ccg5+5NyZR6TsMgk1nrk2NUfZjS0CtR5FkepU
N7brBIoT3xFjsZBJtLHEK6sfn/rFo2U1DnLk8kYAbXHI2vUT193OIETm74u5B3Fn
JGEl+R3zzgNKPSEQMDLEI5TJMpJsyEU3SZmK7FSzdThUWEtiBK+1d8KD3HzePLzW
w8KIMgmdEbqhlbCLiBrk8kmfPfiW4sxO/V4AsSDEwPe/FW7qOQTrqMPkAJFx5WKQ
Bx3c8je9zuOFEtN9S/7oFjFz0dR2JAT4Xvk2U9UyQazOx8TkNgwiRPgIsGg05O+6
RwmqoGr/WRmzxlWNPaEE+/Z6P8a2gsAnm9zZCdql2QEK582zMQzOlqFtepDuCCBw
FIjT3r7sMpfKhhz+yN3mPtZzAVmOrdi7RUmaV0jZs4KKBXYCHFEsDl10S6AvPBHa
2yoXAEIcqBBL4+G4erBbA7e47qWv4jTVIBDEXIgX/49MqI2LqBEpjaRSad3VabAj
f8JZb4kRo6FWa2f+2kQt0mK50BPAW4BGMR5dCySUxyh+0ivE0ygZVd3j+kjgvBkU
P/0LSW9kBL7BC1zZ44ZBUaekdUoOUtjpFOR0NtLU1EcseCtLrkyfmu0cvS3/HWKY
FWJQLo8aEtq9fv+FhFSTSrRd5s03IlphngCRhjgbiHvwwxTJrTURhK1Wki3124dP
+2aYafFerGHpnn/zLs4hXHlTx8O2n0FqR4vNiPfXPFZbH8ZaFCaE8YInDzJXxEaq
L+JTvB0dwdKwoIZk5iX6P1xrqEYkl2iHccC1lO5d68lc86TONSp4rTYy5ZTDz9oc
nLOX2Twv0CLNYYor0vy/uILsKRT7Ckz3Fu7RNMpLVEzDqC8FGyCaizmI1Evq5IGQ
oJWM22ZqZqdX3LKcSmY7PJXHJ9kUYe8yc8cW+Po2FZss1jvvdjo5nmqvpZZ2TMW+
F7BeGdMs7R+DD8dZfgkcsFGhULzAPf75V+pfje49CTX3jZvoY54sas5yH0zDTzhy
0HvDEQ9H9hd1PBoK4VV57IWTGB/44/bh2/L+FfN7JwBAmWz+jPb60oV1F4bl4Grr
Iwn/Jpt9nzjkMI8/D5fZhQa+H4gc+vXDOmUqFWVmKcpTD99+2zpZVzzER/zNkSFd
l0WQuwR2pLZQO9ENk5SjGZFZq7I5eZ9woHUATTJNeve8YI0IlEf1JEAwFULUdh7+
lJ4D9QN3+vmUoLMjEbOkJnmZAJrS1whHz78WLarMOHt6FJQwtTOie9BPdmrVO4WW
2EZapJ+gC37PGm9AwbcFwFcF45QS8s3fdsRsMhl9wnEOglwdMiOfnFOlEIC2Yewe
2FXZw+ajGIL2+UV4bK4QtX9L6WxtbA3dUU0h2iPsPYaqnZ0t1AHgkiD0479n92FI
/ITNlyJXm3rEpV6wgxA7j7yLWtwTiqGthAWzwkZ0Zm5XJo3fzMsuf2eu/tAPpwaB
lJ+YA2OFpQqmBaeWSnTeHiFQfVtY8ZW+5p7DCnyKKZmnkMXWzWnRilPEKy21AK8z
JluPe6SaAeTOpvaFdg3lqsTneHT3GmmWpGU6YecMDEx2642vS/07cua2BhIyLVga
A4MDQag00gIOhZktZkGZJLten4xV0bX7BU4tx3pFf67T80QQw5vj8xe54kOrhptc
RWXySyJzWYLlBp9lVEPMih2d19SQadE32si6byIduJIMNIWqERKtwy5Rn8zLdsqG
Q3beX6yM5SZ4GboFKfXgwI58g82wFXmOAWNUjjDj+i4MHtZNfC2kXbqRdHK7Khxn
oaR80zBsXk/fgByubtXA+WuhYqjijpCc5S3s9m/H6pd9jrONcAeIE709h9BbLDN+
rNkuYELAnh00EY0jdB1CjJBtToEZEeGnqGnjT9/YzOoQZRKCyH6tqN8IgZAP2UWR
Fe2r6a+Z469Fg6vGUyWAaNWPXrGAnx9GSHuzGKDbQyPtSskmkg9SUN1pnkKOu1Bh
sfRGbngC7R96DZ5QWiXbyGjAI4XBsOSupgl5KJzMjfPBqg4i68yOBiEe21VLq/D5
ekjGcGU5i6ubBmYaQW8f8uH6oNSTnznYiJj2AavMWn4e9XqomcPx8VRBAf+DUZyL
d4YkmNvX3rv8NZfsGEm8ENTPTfqnYlbDhXzv6yzMaFD4fHZvJqyFmpcprKhyMawF
o5TTnQK/Y1o8Y8im31zgvQ45qUNxpSB/p3f3ussl0BYa8/w3ezXj4EZDOLafmseY
MFIfAHeWk8HBIaooyZIIxYRCpnvIBdyIQyG+3O6wezOpm+Czdj3aJrhk5ckWPwF+
Pg8CFkA12k75C964XH3m250myqU2pUPvwe3C86Yh5vjKxIaqVRQvCT4Gum/WJ29v
hRDkNbf/KcWVZ/C0ySCuiGdRDjiP2vYTXGJyl20wbl/SdlbSqTW/BkvXK2E0dswr
tNP72lVMTXtAuG0MBo00fyB4EOwisby/28jPd3a3mq4TpZmhSRScXdZPWev7lCYz
IcHuNt1dttidG+9EV0ugBncPAYcsWczkJhEDKEJuqr8fIT48o3TRxEIfLkMrRoak
z1fTJmOqgifh3ENhKUfWPwyHcXyKs5MXyjRPxqn23HMeQghcvoqVlaOPuQXj29C2
IcMg1FxA6cGwglf1efnC6De/39zJgU8y34yMAFQo08hTQdWgjAEjBCX+R2tuFcUI
1FRACpu44yR8LmAsQ+0xuQDWmh8WMtSQI/jCMPUA77obMyz6Ib2zq81ZtVrBb7kQ
P7R+x/PEHYCeYw1w8ihs7ZWEAHMG+EKCWfoNEibwJpG8mc4C1gk7K9g1ngKNkjzB
SHC3jYHLQWKmDQrC3RohQeSrglgxaqvSlRK6Xwhjd+GKU5deC0oluR+VJVSaZG2Z
ebz+iPsqN4QqGLiig27ixmVhW1qH+64hUx75pOvL2VFrjAxjP/G1P52Xlip0M0Le
6+j9tBPTVIaAtpYpyTUA8L/bgHhhM2pz5k6H4hIpJSAoCz/nebOWP2lzJNBbH4b7
1uFkZpdrfu+JsjXIopzOWb/nX1FzKPagDyu1UR8LOuR7meu+9syiinNXu3ydbICc
6j6sOrDTH9viQZGJSPpWeT0uNONiUzej4MfHrILvZgGbr0YvgVYvH1WCSlZAxW1j
gtUm/pSHoMYcuKS6hbbgIFPGrVE2sqTzVvDqkA0yYKoKlB1B65tvR7wLbN0dBtPi
C863Z5oI/jfCbVCaqQmpNFZY489ZO1+BFnJRUW1WD+uxgqstpO+SsQ7IjbaUxF4q
8+4UGaslyGkyiaENKub1OUNEFiYxPvuygplBk6LDYSRaWUF2ht0v7aLYEKAfjh9F
raGk/7OGHJQXBYPWVpX++yCbvZOphdUHGSL7ueaxuHZtIi0/2WrRuqnO/A5Tsmem
1bcbGw1OU7qmCVL7RV3/vkG8b5oF9PjfCmckF5yNcPK5wRCwIjgiooVTMIwl2rvQ
O3KKgcMv74eV+/sbwEvyBA8XsLKSv9r47zXA5woKGXcgq7H8zrp9glpxDvry6gAo
2qGL9Gglbth9xkeVARra6TZVpV2pIoTK+wl7VWh7l8YBcrgKUHkcnng0Apfkdqqc
LzbnbzgdmqBeHyGr6Z5LMb5VhcY/kTSWxP+txfVmao3eGtzG8PbeDti3CokHfTdj
8/SfD0V4kcegmEqNNNumUHKT2SBGuDFBjtaFNvQmLSOTFUp0ehCF33eV7SILsA7B
N/L94xiLlQRUOXwmG3RGAE5jpzH0ofZbkrQOtIzNKhP0CTcvLMrP48FQAJQuJF/b
X/ax2L90UbBiNA0jWIzzqodv1pn9pP1y+3MmMhk1J/SyuA02QZaC+2jQ9gr/VNPK
UQ75k8OoDnrypntzfmP0MBOHBuu2kfBZ3lt3ovCKYswLssOJZm5nyJxR5vajHxR+
X7eVEeeDWVbbmR+6kXKllR3+NAsO0mOraDONghBfTtVD/oZ/+IkLy3OJyDy1wkDj
3RvCSiy14UuqCjhUX7IXQ4Kq3m6C5mUvHzRNMl7YNx4sGaet0n+rnHSEJOMJBrdK
KdIArcMBaZw3Gm5qT7wCTK0PP1sawRGZ1kqqnzXqWEqqthld+ZQABoF2PK0JOIrg
TvGya6bCYHy0m1MYqkMgyA9raHr8yzgGh/guWFfHPdlm7t++ioW2DkGhIq05ZG4Y
19pSzk3/zhIMlkl9eXbBPQ3kWNe2o5kO5lRVPgKuJi/q5hGLyla6Cb4ub6OPk92e
r/rE1LEoCySKroKV90RBK51zB+3IcYo04jd97EeiKCk29fJpJOFneiP9nNAiLDrS
vRyZkfXiu3BbvZnnZv7GzrVu4g6tJ6MnXIb30Zw88zmiJIhGQCXpTSvDcMDtJU7Y
P49QeIUaGO3lKusZaR+rss8j+tXHVP+g++pJUjc5/sMz0yfcQg2t6A++ObjLN3e+
J0cL2w5cL2brxbIgzUoWrPepafpYimFYPoj8FkaUi3XcHIBBdTmPTh4a3N0huIC9
AVpQ9DNdQKmy7MEOZzodW0lquw6WRZ7yLJC6l6zl3INA4tEIcmSzF7CqW4fj/O6E
2Fzbe25V/EMWX+3mZOJEgTLx9S101fT9Yhu0Khw8OpKXjqVwlYVJI4cOE1QsMHm2
Wv7vlBK4wZSaffQfshQLGzDiSHrdQyY4VWk31T8iqADRGWfoad2yAbTGCjUHMKwP
C+yDH5Ed11naNbTFvFHpCEc9FLHro3MEpGKABHtAikiSisDIjQuO+TtVTd1rHghJ
w/oMXo5gSxk2bHw35sLfmsP/Lp7PH3VnB+03asw1/ooMaXAgx41ppaSlQMFIMVE2
MpcY6hE/T4ePoTsFXLEAkXrrehegJZEWUXpb/zl2DkCXR+RllxZKU65JL1tRlDQj
RAQz10Ka9+WdQtOcYaWqpj+I+Ske985inbsC8mf+uWzoiUV3dzLXURdTHjYkBkke
yN2u7tyfBMvibTk/wvzEi0x78icRXyt2gp7bV7UY3KyGh9taAW8MJG8PNP/UEF14
wLTdit4xbSTfrcvSmYPUS9afyPr0mtUmdqb51sY9wTZiXKUvsozaey+nhfMPz9gb
YbIlWY5kzQgW42Bvouh+4HmcczEdd/m+mFAywl5drhEA1eJrw6KrBnzUHIQ3ih8x
Scj2ewCWvKzaYX7b46hfI6xQob+FWM7fTia1BSY4f6Rcx6y7xWGfpahqB6+xyool
ZlZwfb/q60o2sdem8WBP64CzfgD5tuZNwJMAv03sS9+GpV2GTKeZxhuH2TqOYfXt
QS9YiB+tXLlDRSA7tOmxxDt0uogfx60s/nrVmt+MrSHyXNYgkJ94ZmfO9q5cOg5E
m7RQ2ynC58hSN2MoIh3NdSDHoVDrqVT3RaDaUa+BVexdZDwNWBqwd1gZTT5SxPYz
KUsgNiIjE7Q45x+jdA0C3HwKV4/w+YIwFOivYinPRJnIai+jacbcvi3kETlxqlq7
G3rZcicGI3OIdPE9i/4CMIdS0COtv0/Zx5odNLc7WmSauOsNNpqrGGmRoywXgeRA
Z2wASoEUUEm2gkfgCa+WYGjPvJuu6rhB960sudQw1RKQVn6OIZjJcImtu5/naCMX
aXOkkp3jIjUzvvL9dutsHPW/eessyhL2HxywfEAPv61zetkEZmKtbAZxh+/MVZdu
j7Kgdeka0iu934HoGK7Q9nkpC2cAPlqAHqPDfuwCWuHbp22MW4yII5dz3LXR3MX0
Z4ty5+febolYHjrwm8aUSVm/W2tsA/NuIWN9FPTQuu32pqhUq1ZOTMr5Ws2DQJhG
0lrtgO+KayEagGroYo4ghgEfQ2sceOuoRq0P1m/zfiijcMNTHuoOVilEQGszR//f
nl4mWU52JEOn6dpH7Qac/31cSOAw+mUUiOvZCZh9ffC8VY0n1V4YB3N9dXQgBkEw
LXdW+8IgSmmydjdQJ/P832SCZUigUl7IDa88uMqACUbZHsRdpjIMx1d5yc8XNLHJ
qZZ1b3kRrjmYFy8gsDc+WWDL6FSrcKvkBXChNfA6a7m+7yZsYne3Rs8tM7t/KZkD
MGAjpTnSf3XZilkeHxmEXQ8wpz6s0SsIUHv6z9tqz6sqGZ3k4dd9muXTxAUq2plY
7cYmjlrtIzYcZxR0G4L0kIzKF70k5V6y7huFm882URIMTvFMupjexO8EkR6SXFLq
iXqycUOaiyK0jUYthJ4Ugyv4oXcPuWCA34maRvi/gf/uuXP7rfEkcWFtcFNOm5ps
eiVIsU3w3HOX55HF15v/bDnR6o1Ypm2m/qmkvwGfJf9H+7ud41M+l5xah3ovB394
a9nvHG1FPiJKNfgTOYmDN6fAgEvmBRd/T/Mh0o4mE/VWTT8Qr5TcYt3TNf/qb305
MxG8S81f+s4GRVmiv19khfSOwuWWv1CvIel23Eqsp2h2t6RkhkAHdxiUsmPmD/rA
ktJ5mBEg6bYpIdVa0xmRdeiMmZmolZO9s710ds7mv25xrVTbX5EksK1NPAWvysed
7dDRVpRYd4o+8v2FNoWGW3QkCEoNdVbHGK7BfV/g9IkU2CmWpZPrFy8vb+yQD525
txjYHCbfQRSY1f7MMQPoSnIEVOjBjiu7rajdRbONMf6sU2xYi6FYfKxWq5GjQvkD
bSm4ES8muA8DkgLpGHBgpvlAilaXz2H5hIXhFcKTlxPtHzW8QTHPcD214kqn1s9e
Lv5WrO0jJatotFGMHREd2yjShPm65JNnQdpcIo5qYv4r+P8IXBaicCpBkfK/KNRs
IRe3Bs/S0GRd/srWhfooEZG1hxpAxmCWCpYfewILmX9mTgJyR9U/Ro181Ljl9a49
5/MdDLA0zovOsk162PZ78ah5vPG2FoJpHyzBIr2WJWsic9c2EYfq78snxnHnOq+s
iHescUyeIwTsA82oRwgZG62ccyoSDF6Z5Gu4vyKmrqT+8MFbFNCkCmrC5TR0nZMy
xUYEs7YbHZ1MwJk7Pil2nCJIK+7m6wUycZUTi6kVUwi/egKz56WD4nN/3+XwII1q
uMNmWpnfVHcyVGL0HM6XXWPIFDjphBx4rLOBI1wu0N4zkn6dn/gqZMml7iiCr2Gj
3Klq5hNHsSpm7q/XpSRn/7vyIR8U3fh1R3W3vtC6FpARQk7XM8d4BV6f4B35MlvW
3fZ5OSKLEE8GPNG7kQnK9LAD6S11GYAfknG4jh1VTLVFY37sxGe3/vzmIg+N4V1i
42nuakPWtv5VM8rud4wHHub/pppO/q6Q8xq6eMqQuXK3wVgEBLsB2ky5uxEo6uWC
s08zUU1rzPUh7MGEl5LW1h+sZBVsmLBsn5XTTjZ3F27nXG4oPcb4eGP96SG25nI3
Q0vi5vhO8psAGHqw7eudGi8TfsAq0B/SMks8AUg0DfMGZFqWhWH0WIsCH5Uv3/aP
5JXdZVBZOrYXW9tfIX4wSrjZ7oGmELzCzU/ns8T59jQybexEDNgs6eZ+282eK+Fw
K5ThslUqEZFrVll3ozNBkD8FwoLaLCIdgkpiTxluLpc6WOEIihTmS+LtLSsEFtMi
vuzGIJWI2xlL9DmlQGEpoBDFdNFt0UzNDJj6dfzBqzoRKR7BzlDMsk44iV4kg4hI
vFxxSjQ8lDvViXJ3zqUB1jtaHfwCwpyX73Zn4fdo8Pc8SuKsMsvZGc3R6viaU4fH
joEcu9C6Fp1pGDuyNx1K6i8MMneW+dmlHAplq2GNZvYEzVT1BG8M0Q7sOPf8d2W7
CM7b/8Fhx4SypUlQrzhZdu1RSli6SFIpcTaiwjciH+UN49v8YIlCcGX0lPM5NYZd
Ipz2FT0mA0QrY7PFnaQy5XP7/v37mntkeTVmBnZtb8W8GzdCIiWXTppK/KhKMKq1
GRY2aaY2HzMOpIKerFrOpY9wccykzo8Vh9GSe4UTaL4KQHEZhHupHN6Gafz9a2zT
y8QN5uGM8b/P/BGUHuTyJFysZUWAqYJ1XiFlqqxVnlwF1JB6drKM7QFbFKLPGKz8
L60sNqs8L7mHQ+XhA1jnKb6eiAfiCGu44Yax2KukRqlv8QZxEEM6CsUSeKDD5dN2
LLyqItjjS9ptA5H9IfypNePJBB02chwaTr2P9b3h+vgXPKHGP8LVlIwHsm3zz5d8
MMiVB41cHFH5co4rQK46+dWsN1jRzpwjvrPbQ1N/SD0AtxdRkrdaRQSv9Xknltqa
N8F8SNY2X46qUFRwiwQfudY2sm6vLPe4VledR2lcmgdI5FeEtWJW4mwpiWhCFJQD
Y2hzpytCo/LqImZzRjKrL0eLwAbyXza9RINajdC+Svps7+3FbkPoPFm1ZnXMRjh5
1/nHBF7FBchKkIxYACK9XesEE7GaczO8fwPf8ie4ecnowTTJszvVCLlqzAXA+D/A
tNW3oqG16gpa3f9ZqYV0yzidsbV/Z8ODLUOoKQDOHTMHlgozHyA+H5xNTTu/4lTQ
tZoV8hNnwuX3RgaB8mHjk3izEEFSOsCl1sxhPr7K4GohbpspTpZZdnpooXDJrmh+
WFwuxAf08rUvG/lc2W+DTBAzgru8wTNyKCntEndtt5EARenlsRgVQCnL+LA3Lgye
LqBWAccsKEUiqQEjNZKZPjJJMOS6UC4TuPNChYExWgrqiAx3UIV9iSrg1e5yDwcd
TBP0+KxapMt4wPUfpvy+uOqF6ZBipEoSj5zQPsTujkeRTEc1P3d5XI8oIisigU2n
3vloU+ixas3aPX65/f+3YWnU8TPbwFj0X9Zz0nTp2cWtAFgz0fR8f5chk1XL2fQU
bJzQV7D2TgQJJB7KPhoHMqGRLZyT+o6MenujXEgxOclxS5FZN6hWF5SSXZdTBSx1
RIlXvr23dlq0Lv7UV1GLg8zOXWuOYEAIUEHwkTjeihqGSbS4rDK4nurWDQJjn4Ee
QthbJmkYRaOssEnQxKsWcEX5ravRIYJ4AgOsaT0ehtJOgFn9Mq3wkxJanW7g1GY+
MeTTqOeRqZ55/4aNraM/3+qFRkcEvz+VE2Mr4Djz8acNootpMvOt0L8qMIYr6K0f
bK475eUjlm3jwq4NBHKGHdGqhkLgTfgVnkxJgUi+VRS+/4/B/dQTVNOqmPzO3obV
0v5icLdG6pkr2mY+HLyjzJKijAHUvpTm+oGQWhUdf9cmhs4ZjQBOdzoRRAdbgK5w
PikYwtEX9YIdILuV+pnf9Pk9weg/KW+4bAcB1LSYzpBV3TSLQXXzxi1dnln/UrQh
70oNKXVJR9nNDMIapUZCAxnQv3xkXQtnsKOfIyleTup4lbHM0SkSWOiLi+R7+DnG
aCkmMvZGq+tH+DA/kf9sYo78Iaf+i5EE9sIebJ+brLKuTabpJX1XjqlcVIN2undO
uCuCOA6XOE7/X3TKftCHlqrfNlCItwO0T2e3UpsfUO1MshgrbO1EcpIT9wCStbNa
c5wf6Xl9YsaZnAOkeGuwC/NqFOUxF84HLPCm4QgZjuO38tdOrtfLtslSGHAhPK/C
DizrYaW3/beLEewn/pHvkjM8Sq0qRXwGitm5W6guhjCvotA2XAurDjSFZDXe0Nkb
Ncn6Hx0sfDS6nruGi4+aUiZilk1k5228xJ7XYsjiYlBgBXq7nmn/A0jLZxkg+VZJ
y10oaYggauhLphDWhLTn5PCYChGZqX3qaCXJo9oQQuRd3sCt9IPW23RnbLrFLiQP
r3KMH9DbtWmO7/DIJps9+qqOqUUpu6lHwMNLl8EPIin5Q+9kypzgxZu6B484gcTN
AR/TO3xcdhcBS/OkE01ioeDyW7kLgUn+iDeFSqG5z7XcPd0BxmMVGs8saAUuf0zU
8oI6mnAqI0Q3sfJU9YpcTkkFSmb8OOAxW2IMQd/zI8JA4088KE8qK5sMGj1njyIT
FcjB9nqmQ7Y7lpsxTPc5lSEgg+cV+aSVIajjV/PXScJFdLmhlNg6ubgbI4WvVhda
n9O10ZjuoyzgciNnzXVYTYqvk1Wr+VDYRGemn3tmeOnVeELaL9O9DVA+wvyYGfm3
FqL0j59/JG58acGOsPySxxs8YvJgiueNyBnLYs2iW6KtvwLpxgFw65gneFH0dyA4
M8eyJ3LZU27m2/xWdZXmhrh/vKwyMOlqkgj7Etycirdrn1APNtoWB65LIc2yP50v
z4MH7P7omTA1wpoysI6b0nh4SIen/590aW830/iNlY7lMQbl6Cby4C8JrGtO4Xeb
xWULbzYKuFqphRgCPWNmq2p1PtqC3BA2n2FSgfSH/dsUhQ2+0/AhdLhN+wHBO/RQ
cNHtVpD+SyMxrqkomPnVXjLNnvfiNFFEpCWORc8t88wasqbOyfCG8/VzpDnJchPd
E87BWcHU+PwYw3SW7FvHZ25ahDWZ4IfrjfWiD7Zbz+AMkCNeXCaW3rysmUgo1ufX
L72G0pEiTUgrwr4+11khOKnvDdxLANmvaIbVcMXy4cLt2P9DXJcs3JhRWdUmwKlE
s2sfSHuSTDXWq+/0S5bOrHtSxMhpDT6Vcy5cnyuCrdXmWoWNs1Ul//4AtRRAO9rx
8On95o3mwLYloa/rjxA/e9KaTgcW2/3s+d82DZlx3d1rsaL/5vtRFt2MDYkxqrNk
33nehMpTZHFWAHNMK04Tk+koJmp3LeKhVze3Jd5bdhqakmkvrjKJnhEvNwxeQGrC
UdIzp7nVc4WtaOkZgx2kmzShLw+AuQFLYNEK13x8XOTeSzWQgxbowlw6gwDTvuee
oHHMlvaNUOZlMSKYZhP88Dg3F+URFzjBcRsPaNAOhEJ889WJyZSlfLXdG93SV0Co
VChKzq1RewlFsiY6TwPTh0QfrDnk7KQGFkSnUZQgIbY0qP8qJL+jWSfmJB1n5EHh
Bqf3h+5Z/ck71PaKfOGSarEaCpqK6CfjKVlxt/tWlQEZ0sApVKxtHkJGLBn4A2G8
dkrDskv6sc/+eMivvjKwBGZBP+p/q4xMEwa+mWoJyVcPj7pjNoE19CFrw9Ediw4G
+iblfGs3lAHXGVN55hCvJGKB+I9b9p/F5UHKXyEMqxtalevtc9m0SlXDbl+FgZIe
TZyoNnarB+xklwrlv4C9k7z0QZVMzkA5UI8beTJ1hEczqyzizpb/OtnnuFT7liXx
1z3gIHsIJ75qB0O0gvPpyo6+fcmTK3FiwyzUnY6BSxwTRatwVZEfH+/S/hmdzgLr
i1c0OvrrDXWF8xnPH9R3vdIVCQWNVcXUeCfxBmx3JheeLv4Sm+I5XACxr8Z7Adbc
SBY/qghzWpwxbQ0ctcIXd8A7DZ/QplJvkGUIfB/sPvGYloJvuz1NsC/Cl53s6r0c
ZRi4brF+EVuGd7UYGbULT+5OISTlqhIj00hBgah5RtQ9K7hbtVCltVylFcL3TKer
uerQ+0G0NeyGkQKEIQUDedU+VxsI/y3ioPQ8e4u6qUVKsiBKiFvglPN6BVQgNfsa
hVw9/jOJkSFDQ1/6rG00M7S/KmZlO3oVo9FO7ClJWYyu2/QpBlF1yZSRYX30tdSu
v1tonu3blh//V0n5vfCe2nhGb2CMoz4mEeTta+Ad8mhFRTrixZK387GH8Ij5K1Gp
7TxuY4J+BA4GUnqjxvmwF0EsdhVu3AVMgJso6/JKOHmUGPWAcCCBAKUFZkCS4MWe
s76cs6+sTixm/YaIpo5TugjW4EAqhjicjLW7HMCoEsT4kl6Wnqve3aSY054VDbdw
50bZ3FoJrqxh7x2a3rtOD+XY/BbkMy+rBhiF6x2Rz6Bb6JPTocpswvEqQ5mN0z3G
8QKYHgTHpiWii7KpXWv8a2R9EWutYZOyylcNiw8eOxRaewtSsYnbylU6FJAxagHG
PNSrlQbxApPlZiebadAV4tFPRxJ6dhsbrtuYDG7M66o3cBArDkT/nDdsIATy7RN6
cnICgKtoVgdlP3zVG7SeGLHTw92TK15eQeQx/eYCb8He9RhF6rhaelWN+YTfBvEg
loTUAhi53rQElLn9WwGFYxy/rzHe3G8SA/OPy4PocMrr4CjclCt2aXyCfodC/zoQ
BvpLEZGhWVwnJ2QalOQlB2yyEudGPZLSGDxdEMres7POOGmF0unhkq6xzEoa+/Js
JlON7Z1L1ZQrdFQFeYwcSwp3JDDTcR2Hbu6/FHX8zmivNJnM2dHrO0AT7L0W3e3k
sV33iq1GDv9my2G3+GwqKda+70QRg2JEDGbNuQ4AN5ob2euBEf2sGZiiu4qSbp8W
4m8koFyzj3ngvl5TfAymevsI87iYpndLG4x/y+ytiQ/FE8HpT/rD0RxJptiVLFEp
d7heAZglVApcS/6Eql6ik5OFgF51SmwcrEJjfKW/4/q6GW2qHJkdYyTaeAY025Vv
Ct6DFFuNTF4bAv0U3DJzM1nDNJpJ8uajvwc0odO6zwDOIrSaBIZLyOdgXXvlKucn
m57plw4Z9LOsqfEoPVg/Pl94u58yyYLX7SaN+eIh8/DAGW66rItpNAQh0hQlUva1
SLSKxdiMVo5+FaPkHwu73sZtE7gBddd7osO3tSmYVAOEJYEHIel5pRMkPk+ZHYFD
DvLEOqzNrNWxk2wxU7KnvmqexKowCVp1PCzYe23zG7xQp77/FSZv4xfDaaxagxKS
HlWwyDzPUL9VFhDLWUs9N3PpxaRYnsW9Q+Ge0lZNMCdkaXO1gQ5AI0llarmbLixS
kfBPqq1JUo27wR2FUoNivuMSXw7KY4kJHU9abCwCBhMoqQosMCvNyoa2gOhIdvqd
/Tfz2fL3zyfJM3SZrOvt/EPhjKgW1JtH98913i3/AHEn3B/qXez8L7FMvB5HcOC0
t0HifH8I32lmd5VnZ//FXbNVsSYmTCpGxXnPYHkuOQ8Qy6IwYavuvlXnhLGac4z5
MS0PqniVKtnaJHBw+YUwzKiHRNRv3e43spyYPwt4JdFN4fIKvBkD4WuFRocndwsn
PlrdUwGkTxCEvXCydFzyHtnGTNKn/WK3XjAOw+yW2L7vtp/nyOeRVVmNxEmKS4/T
9/ljWqaP4czO86VusEIINnIC8ki/Zv6gMi9mNAJh1PNRJFstPyTNaJnKKxQPem4D
Dx41fhKVxc+qbpgFNHzf8cn624ZMjBrn54taIPZ3LhNm04Mr6suNcUCYnq1Ow+ad
I8yIdY0db9OoloOEIUkNwZxE3SmLztcR304+iEpc9INlhPhox7dXscJKT+7Q/OIL
R2h0d5ccTXnEgJzsCqFAwzwoES8zVHK1Fxgigk3OE6l7BSdfKEFpdCBwA+sHLArr
xNFZdeNA8+JfNJpr7qB2Nn+ReCfaxR0KMdKSojvT8ViK/Z4FvSGPMWTpE7EETZJN
IWQrYp7JTmJHKjFjZns1Qc8kP5UUJGH8s9l4T+CJeJ+3VpJlHt03EFQQjltS4Xv7
bVQtC980Rb5NjzoEA+WkjIfsWubGAC/ean9jDTm23hvHsZMsksYLUqs+lP8V7LF1
0PR74TBBvEbV6xeqFfEQq5imU7DFvLnNDMZPF+KN/wzU9CAGAsdkhMDQVO6rANy/
+wzcQbbBDhECN8tEkBWrtmlxRlLFmxNt1Ja+usrFzFGasdY8VVWN1lefNrMvvmOl
D2d5rrEcabiJu8W36Dp9YaCh02ZRmNvYBcgvKDPntVDLZWRvmS0wq4+0cHam//eh
X4EB+URnMNVJjx/10P5LT54LU4IDowhazn1OoGccEcgmUxhiK2irqObTcvt3YA7j
+QmHvlYUA2asGo6w9dymwHpULGNk7WemLwRSWAcECEyD9V4L91yllzjLUy+5QwRp
Ch7/73MHD49jNodf0/P0vuTRNhWfr0KcE5MYfm6cnhWbAeSqVtUVgOl+ZTy6Z5JA
FXa5iuUzjjrzysm01i1yL0bTnHxRbWElWS6nUn+hFSJ5S4K2oqs4xdIKeCUZ1hYV
vvPteOnFxBUDt3juZrklX8ZdIgU7NGM/HKNWHdoYEvOtBcj4SYMI3Fafq3sTjCBq
y1zTBowuQB7U4YSW1Di3PRgDlCq5ELGfvhHg/1WNhccR3nyBYGiI5CxoMl0J2hXw
3NN2pzskTMqLDox9Y/Zvz50gSpYYHFGfgGCKFa6j65AKKHeHIndNclcgf3Yq6MfP
MRH91dTjPucXYX4QVGuKEtvswNnl0iCz7X9T3jz+zRuMTYDJOAfGrEXcpdBhPr7P
0a1Px4t/mvSfN0SCURF9FHAhCUbKdrit+kk8+17ywPsx4k+CZ2caJz+L1jKrGYGo
wlA6UteN7mjrCm6Q/TUI8Nz61iyFm1Rv47WBZuOeuEHtQX6xaMg0ng6WV5nZbNvW
iBYHolfOo922AdKN7subdTewUQzktK7eVU/4PpN9YW7sdLhEjQNVC9ZEFBpXcnxW
zsxY8fU1h9Hq2Dj+B3Gm0QSLcevkxDKAXUiFoT6UAtEyTSNIpNTYcZpuj2w96De9
OTvWzM+rMP02wlhyK7AG2pweGpZtcVjuqaPdH3cg5jyCKnk31wCXGASxbwjHXI13
uJB1ZqCZWSbMLQecWKgR0gVJEkY+TbKD3ppGIuu0yE++k8rTEy6WithQayajL6hu
BIfB1P6CCH/eLKyDt/PH7z7D7fUU5nm10Ff5U4V0I6Mb0iZ2J8Zsxbd6X+PA3jLk
ZUmYG0yiba2kU1i9E3qMtNa6J6HidlIKCOKEPu8qCHxdA6RypQaUU4W+kS2/ZY+K
wPevU1Evc0qiIgM8DBM6QIzqrLtmAjREnmetAzL76P9F0VcL+TAd9GmCeZBSlHcI
3D0Pcyed2ge2bvmOPFfbzWtfaMKdv7B6EzuTQbux0CkJDt19NhprqHJyI25VTFPb
oI4Ih7Ra9g86EytGeR7IyAbl8xU0c1IUlNW2DqDUYjiOAKr5bDfDTKX8HvQX9qOV
S/4D595qB9kBu5UnRdxA4+DyRJb3MIio5vJiIa7C2nLCkz2fm/C+i3p2gRRpJCqp
cKqVfLVssb+SAG8WXTMWPixl8sG0iEFiWqnA0eq6F0ullj3cyiNxXsJDXXtDkZhK
9Fig0mNHk6x/pgPQE3LXCbD65yaZMnFs6lGwbUiZXg/2NiTJksybmn8IWzMLqYlI
+QkZVEsdQYAouNxMoHvLb4XyHze/oqNTQRVouaGc/cRoRDflSj8gz9Z/KEFYJd/e
Suy8cOJZwMlihcsh4AHI/bdVKMrvFPsKSjUx5fCLDy0rKxbZL7Rnwj0p5HZ2G7PU
jcw4lyExHdbijGvPp9WBHi5aOyZq7geNKN0bJ37yrKn+wYl+lnYNpbx4ovMlwEJ0
t/YbHE+zmhdZLW2O0+Bhgbn7J+ffIMNN/cwp382Rn5M74fXLmKGAzQnhSeiJrKl/
EX3fCLUwFdkJ7HUqZCK4QweeX1pVe8LyxlvR7U5eY8dfh7ugvYV0zMtlegJipUPD
6ikMTk/yW8gvN3AWA6u1UT1b2Wj/9sbx76U1VhXXe9KhTO5z4d3/VeL8XbaQS+XC
GYGaabfCp7CGIjCEJFRYqEqXbuWO3zhIOhB+7YYH14c03A6cjd+L7nsG7G+Dnj63
tQTwCUe2pqs97QAgCw0FTsEI5/I3i+CbCjwl5Tb7+hrhrIrkvJDU1njN4qBAm9Xz
Rr4qkEpjJAtr9imc8cP7RSRRBTTV3sHl7U8yik/cXM/ZpNdjY9RRsQHB8UG3PZU8
GthSCksTkiUr1q5LKIL6valJKSnodTYM9ALVTrImBo97opsnkXH6hNsOz4wyN0Jf
1Foz9OyMzIEcOiVh76IBaKoCvLMozyBRvo8PBw7EQHvH4FskpxCtSRM3CCD1zfFc
2lY0c72FL51bLRFZvo0A8sIdc7P5cSoh6vksXsp+nMm4oReSHUgoc6qNEzt34LrV
EL3vMU+S2QIkVSxI24APZDochFfL4dd+udcSftDdGQWsg92NMFq/QiCom9Qah1Nm
VG0dADf/n/NKNhZfjbM/ju8rxgaoD3XMCtG2I19J8kfMX4vx1jhPhB8r4CCUhXtG
yJ7n1x2YeO0X9vVv+IxpGv4Gm0gHdpd5aZuA93FZfhS+mbA2k4gKP7yiJw5fI4dk
Y3TEG2SKfgGoF4zEi4NQuwo6bxfkWaENHH5keA6Wu9PXGcyBnfEJYRFFeaNv15tF
pj+nJJw9PpYFmeC2efEB2UpVUzhH3lyg0BwlBbe6cp3oIFHLBQ/VMtEEJAzJlzo7
NA43r3usZbdcFmZQKMvoASq1dhDsw5r5P8BfWpG4isjHJLRYwMWxKSRW19HGcY/9
P8qDkORqZPWL7f1DBR7u1Sqxio+4KlTDKB4hjwUDhotg6d6bGlZReun8+dtFeYHx
GykuwuHonORpGjfYYfs7z4gV2h/+KKs8iYvcN7e07xr7lTfQQYH/0273h/fK1iR1
A0y9Q313IJO2YsEbw/sGqbQYSo7DbiF6a98F2stg3WU0HhtBf0kGiS5NpxhcgO2h
JYUgjs60YgT4+jKskqkNEKY7Xi0IZUfp4WDA22bT5rf4xwed9sWZVyCEbjkb99KE
M+ii+5q9hMfw7pOESB5jCBr9tsmjDa5VhwLGxPUnWBXh6lPnzi3/x0y+wwvJ3PkJ
5nsa33R0ROea2A/Ozyc1oWSBhRSSuugzbmEWazeDsVZg/Dl6qyHNDq4g7TWcmwWd
a33lzmD4gl3W562SwRDV941/N0h7JR/AiJqnjBj+/H2+aVUFbfUz5C0Y977VqqRz
1axdY9UJd1BEIEfCtRztrCq8V346gG8mga7uPX2SQP3ks8KaiNIWodun+3KXytvM
jYaOY9wAP69Ns4nHSS2I3ugyDHu7ORrmzn3EEpCAm+n0Ho7VDxse413fESjg5q3q
2PlOPgNTGZIH/A17G2ZuR/29FBL4j1TTZJFD28fRU1suI4AATJiQ6sZjmwO17Ze8
q0OwRKf1Tzgln6JKSZtiUrKidcWt2H2n7E2kMYcj8UlzzwhTkkdBQ6BWHsSyxkQP
Da2Y7eUGOspJhJUeJEED5tKwVVEWA7+B8xU6cg4/5wxPN+KQ/3KohCCM7G+4lx+h
hY8Th3PfvZqx2yB5MLCoUGcinowij1e/+5ZPalCil3oSruvLAiIGBfspk+JsGHCQ
g+4i0L3TAQ2ywmUoe31jeYZHtClOAI5HYR1DMlloNiLZXbc0M9AAreQsCEaKYLHi
dZP4E0P7heacZ47XpfL1tjrJ9wOnCKQ5vtXxr/rf7vIKzWuI896T4jSNXSR0ZhTq
8Bvo+vjUbfgw49WEwzCH5Fl2n78TjTHLrqlh4UvWy+vyh8YkNiBFkVtQc005UgEe
uq/t7VkMD1y8Cf8UVJj/9U9hao/x1OcOgeG4o3J2J4t4nIm1v3Wtz61WzfCGSChf
uB1VTFpD/PZm/HW6medvLWG5EMXyVmhNycJLO0DrtKCbCIW19eSMd0YuWbApbZaj
wQGEOSlnXMfXG8TNVyInAQc16vpijDad1si9YUp7/OEN1VFcbi6VtbLVMjM7FDSk
hpFERpb7kojGEbJW7BRuEIebqasx7jmOqHIhc5MCOUdXzp/CW0796Ik7LelhVxtk
COqAhnQA2AQPva5VVNxmitNClbagjOYGSqUnEBmWTXtnuU23CviLQ4moFlb479lc
+7snsvyLUcXD06t1O+lsUqlx9niIUmL8OWn0wT2J6g90YvkptsP+p/McuPS/9Z+M
txOdeLri9SOTG2YMeTghZos5dQ4yq4e0uiZQjObY8o0aDKRsHl63wsyF9om25QaV
SXBqCNMnFnFEaJtPpyfxT2v17zrRozPARRPL9Br3ML1NDWRfp9NNmMG0GcCLAT+s
Zq4SYPolN2JcF7Lmzusq3Nt9HKJP/4bCpBI+U9RoSYjMUNEP+D69XNMiMBozagGW
Ettxl5ejZrAxXZvFmkkeN8MZr9c0CFHCFTf+5vv+7jnJw1E7iQ+ztcWWik1nO73V
t27QPlY8ZzupSi+bxwDMWMij+Biwunfj3q9uWVgkNgrAbzFN4dZ8UgiYTKe9tDqp
f43euipBnzCNJbJD5yTf00wz6WHM7l0Xt2XrJ2KYCMsqHBhMw0Bwm8N6eDHAn9HN
VOxSd/z+DsD1W7jOQRYc6L+VC07CV/U6OHYpX2VgE0IAkAN7myta2cHPsxpJUznr
2TWOdqslBw+CLqRPDV6YOENWKf2446ySyJ40Ecv77sWns3dcZJs5iU1dJ3MPDZWZ
EGMzHU12P4JxOL+wn5bqITb7+MTjCeda5F7gS5Io8RuJGSiTFKJ/lO/JjSVP3BVI
R2K+vy1wMfBjO4sU/098+hbj9Lp5X65BEzLO5xOcLciAF6SguPEiE7golLbHTSW/
gctwByrLjHa3OKmUPRNi7GQrx4XmwZFfqfk/9HUy4+VI5qNPePOhdg8LiREANfjY
I3KDHW1JEDmpFKIEUL7hahjJXxhG5OlPTJGYEr1huBe+goVZZesEBMgd82Hr31u4
MsRhMI3mxaF1BF7XJ0zMHui6cxBmYURas9OswczzydsQDF/NRYFjoliNA7im/xfN
2AtRJkLtZjsu8u0JxVUjqRV8+FM5GumQbNo48mwgZZK3ij+dT7zPhRghGYpK20wN
ZWeUIl/TuULcIHc8sV27F4bESXNQ/pDPhJHIObJPejPJlEHtD9xaMfa9CBlF1Ywt
8vsp8nF13ck7zsouAzD1WRC9N9fFfWJAwtkpuyroSNWffgNSVYT1phEjvBh4yJxi
yyUlRYUakjZoiEg1xDPJ/WW65ro2jz43LcZ1aipPIZy2l6qKhK8EQ4uBTGbtfvrM
coJTncBj8AusXmOX/Z3Cash3NHMnbJxOaGOyYRhUlo4/aZRjaXe3h0F26NFPkAnD
Gc2fFVepj4rY2hbVvLiW73dWoCe1n9ZyfYho5eGCxVQ9aeYf5qD0rNiJD1PmN6lc
CFn8Yad6RfB1rIVL4vFjNrSiNA0dl+BklwlpGGYjZhe3lqn/CHmN84JqNEL8wk3f
IWAOSdN+ow22vcoWZDbPEi1kzCvdWWboQh1iWbC3LTeZiE0fd+wSIAY3AB/nLXU4
nJDg3Dcp2dHXa47h/cJKmGeDLkuLQgC99WBNzFWva7j0YSMC6iJbAaEYllVhYTgA
kXJCnxAQu2aEvyqJts4xSG/yut7qOfupyWI7z6yjVzlK3QJplR/U/v2mh4fDeN7y
pS8hMdLJg3bljU0seEuKVeJcCUA+HnRBiT1/NHWZx3Nlr7EcAD0C3MqT3BLQTHU+
Xk9mvCY4VkNZT4IhsGayw06BVDczc4SUzLqFwRHsUpiy1lF1ltjGutf3h1+gpj3P
sJYQcwhGwXiekkQ/lOVr86EUSFhed1sspgu5nnsnhq7raK8sXJeazhEtZJp6WvWI
zvi8Of77OM224OtPTjDVREvLTwQs7lU5LI24I11IZZyPdg8XgEuJ1Gpip4/x7byf
jOZj3BEliOjK8lpPoGr8eJHkfYGdiEgvdRRPgPtuDDibuY7cuFlQkDxTYZh/nuFC
CvIUOJqT+iYVlqIhOIcqrOd7q0qzqGlsyoZQCIM8gSPRN6o47bFD1qfi6Y0xd1pG
Dn2ULNj/Dl/lchKtoczLqkymKRAhxtZZF3joBzU2di8ylYOLDnkQUxKu80fyVj0W
EvydB/napiU3n0V6glndowzt4Jzjc9jvUBFcC1CbWqDy+FkUw+8V9y2kfum7xkrj
61kHiY60UPWKrdKcZFVZPXz6+AXrpzj1VKpDXIr9l+6K9tXP7AzVD+AZP5AH4RSB
Bd+yFJrVMbLzpgHBXUqeVw4K/lFQIQkw9avH5zJrrAc4WTXnP0uIoS3gH8c644Do
gk2JWQ7yzMTdWZdsEFgR4vU00N0s6u4wOeC6//Zm/Utak2lAcd8IWdIBjIjFJPfx
fMuL1XCE3TFRrjxEZIKVxSstALUfud7mHePR1ltQpOiZEmZUU2mdGnltcxcu/6VY
LdltxXVkcmK28Ssoa9qK8jXldoEfkBuv2pgwZ/IFIv31QAxwsvZkpi/qu6e0nWFI
KhtTcDVi8hEzLCm80xBsgVmXn0eeoGIqQKx2BRVE6UPfLSGF+r+6YPedS1QUvGjU
S3uZu3nu8LBvH5BZHqR3ZSw+O6s3ZQytKPO1d4B2KvfE7cvi4fvhzH5Nz2n2/DtK
o6kAW2Pok3xe+aiVLQFrneW0jghKhZUFLOicva48uL/RukDE7e427Q/p/VyMk+X/
sxRyxZmTFr3YrfpzDDTsQ6V9cln09B5rxTyjT0QPTNcCCjuIur+LBaN5Yek/eGbU
0dPAWt0PMPTOzHCSZNOPX4pAuE57XmxjT2XOQS5dkVhLTkDeM2fAlyNh0M5BKjL6
oMKuGz2/CgDQ4HG+hhfFM+FSJJc31GrOIKGubYX6gKaLgpWm7DXX2K14PUTn9Dyq
6URcrPgYIKJ/TlaUUauYhSoG1SMt5TXT8NdSXvvEPOUfkxH1cp18yUBxynqM3Qmp
h3WA1jQ4Fkvh5dKfxaBBnSs+JiMVF3ET/qQhKxvBI1qdIWQCj4qrckGkXJ8ZT+MA
Aw6e46Bdr5iH9NBKAJs+wH3/az/buBH10ow2rAZ2TgwPzZuecQwSRTBuOHszpWic
ffHq30zuGcxAuNQybXEdoNdzQboASC8gHDaF5hNPzjijwhYrxw8meBpnoXxOF3z+
QxnlRlrxZiBXV5saNZZJGIubFGi+5FHKSj30DcboBqI1un885h1IFEOwynl/pDUJ
sU9pW/dJkbWslYk0sPkX+04390cbXkuUBEwiiZVqWu3XjL7soGhyrrYRBrb2abJb
dzUXwlQpOKW2RNbWVI3JZuk1NT3paEbG5TL3XoC49qSEgtYF4xfAuFmPPDTEW00J
2F9Hl9fMpCXalUqtj3HmHnCTEntGcmmEt4Bd5tdMqL5DpdaENjLfdfRz+rLLV32G
Nn27KVHO6GLgvwJ1Cw+oiWs4utgYfe4CE/lCA+8srZIFr/vRBsxZgr2ebkksriCT
r4tg65XQ3G/MIMqclMbuzs7axbctdkHI7YeVCcZmKZRy/Dl723HQc8EZSbKUI2tR
qmKsJSpO5ImY2+zoF6B+m5j648B2BnOs1RvO53lJ7YmbSVDiKjUpwQO/r11jYZvp
gbhLz+BhCweFvZdNBZCm/ZZ7aLMB3Id0dVUYb6LKuAcmoKvZsDM0ZFPw/zXIoVBo
9Y6vsTaBTqgCgORrjHJthP1H9zHT6BowimKGY7s9Yn5UkNsB1lQgg3axdkBFKLlp
df1j+5qXtA13jyt+tqrKNMMBariFkJPSZs3AzFrejUuxYY+ZL4Fr8FZebtnsw1Zx
I3HgMbLupImMAF0SdiFe7csSSLUWibBhbuvbP7b1PRN7k2592YECF0Tv4HlXiOM+
Y9JIa4X1vJfzILDaJVJ35Qzs9d3EZmueM+4Abn86vsEkD/fSRIyAJkMPYj0q7vjf
jiRnIolY1vizD4d0IJvcEeiegIe3Jq/AmYg9tbHSjlbOpy+tHL3EcrgH/PslFIOB
z1nSLc071cm4jR/7l3SvCoPyBAvyp9niqnsz/BpqnEojAjQDaWOvC60zEyLVdU7D
vh71lhOzetwMGYLOfEhNnYo8gFItW/muuWAnqpO3SLxBLDx98w7RVVKCFMjKNUyr
s5HMG0zHe6CaLTQFPYd6XM5LGfjSzjny9g7VF4rPiuARaMNsra0o2CKsgpOij2Et
0Q9C2abGYfUomtDnr/mR+oaSJRYOSRpg/N6imcIWO1yTsOqCV7XZMoKUKg5+QRWv
C3EI0Jz7z4aguE3bnw5CcnRErFX67MmnwYyRPBtS0NqX35RNnb4a+Dz3IMOHUOGq
UlH5sKh8W4OAWbuwbhpdh5gnGB/N82EjjtLniTV4Q8PfuaKUpQQ5ueOk3No33YIp
Aa7URPXh41f2xMLx94Z7Uz/3lc96I2n4B1KzeW9hOVIInC3mF+J9WXGtKxt/ua4v
6QCWlXyR2o7zT1ts9TdexFeB/O5qpGN9xbOrMFMwPsUFwAPtj8xwE6MugeSH6e9C
v/1ZuMYa/TLD+6qylMug/8bMmDDUCdGp5bPS0bUQK3OreG2axbSdp792Z8FCRZit
m16byYdN5lw8Wk2sHVvaMXXA0QaBsLcG7X0LOlYm+6072la3bJOrGNkrwFjcMlKn
qumJVqFiIp42Pre67GfKYMzZ8xJOrXOajUyoJBPPrQ/dgO1ElEgKlzGqKbm+goPf
6TgAlULZxN9iIatD87+hsQZBW4pS7paF2ea1QI3fswy6ew17LhzVGNLhWcOgaAMF
7eq4mgJCypvM/qRJKwyLdHs5U7NI0aQtP1UwOgfsKihiZ1+woAIOyvZRfq69OR4z
tqaVWDwzt+OOWplPP/NryZMNcfqDOahXrLpnzKbgFoTnoEoXV12KbACTrvUj+gLc
KxTXmFqAoGRO86m0l6WQ/c3+t7P0uqWukqrDiyvKwBMrJodVk/pbsEqiozqMdjmW
o2j1r7Zfv3hpFEDnst8mXIJJcQcDruL2UrkKa3LlvQiMELPaHmoiN/l219Q+twAD
VuCbfOKwTACE4e1IBLrKbJxzKc64ZsLABaa4YNCysQ9A0VSzfr+RYUl5wZSWTSn5
pTqdIAXKCUiwfpd2nnNNjogVmjrk16FG+Gq/1HZqOCb+FCHesUGD1sZTWGripWNR
EfJxHRVnVJiogvBq9I2NUlpfNLXaOnlqqTnwK9WADKxsCWmXtDF1UL+hFkhVkSEU
OEWpUS3xQ1JoEd8JjAhGstHjH40VaYBVFxMoeS+4yJsllPdLb7ptwwJ7l/xss/F+
H5/BbQWMg0ghpaE2cxHM40YibIy6R8oLmfoL58ppXbOX6iDVhcGn9DnUGb6rMuer
ZdlUWTMKXmx1IWEHPR7uLBhY5Yek4wQv7y3WCMzcB/IRzSRfW79rIZPHeQu+VDyV
/K5kqsuhjlkDBSdwZCdYYr1r6FEXjXN5smo4OqA3pdyJZZdL6fOZMCJg6Yk0F5mu
5EUIQC38xaTu/EhfOJYZ9T8n4lJuKqbxT0VuMNTaYqZ5QOIA98WwZVqiZ98crOQO
zqbHdp4SJwV+JBUmVRCDu95V5Uu/UVIozndDiJCa7bXXjwq7tP5VGN6k1+EWj7//
Hqh08r6iW7Rw0aDiheqRkfwRqO2TRnCy0AYK8Qy4m6Ld4fdwf1RklQfBkufRdyN8
wXWwoTmrN0utDBUoYA/ntXbucrxixEt9CFv3N9PMILky8Y9HjctLbwliHWuC6oQa
yw+hP2EITjLidpYJmx6Qs+gJaAtrpmLnK9rZssA1NKWdkV1FlBuAY8oTnol9vlhO
O+JdbLfwW5fLRiDzv+8TUHJKWCSWiNGNxQC54B+mBEmF5+yWmUGim+rePhMGwz12
4EusYOjDFa2h8+gywNHJcApOtPrEhRVl8pWHW98+xlkxBqgyvDfMDJyORW2vFtho
1hxGe1wQd88aY2C/W3oDwDWOWpwcHdx3CkJkTFLlwRy7524A0Kw2j5IlZ4tE3ZaJ
RK2ahBT5ezu0wqaFD+UH2ybIRpncpHLjMhg442RHkMAQ8Q66YRJ6GykPUHWySwHx
k07V+WkTJSUUHFUAeITzH/1XerH314d0J+dc50WA4KLuhbvzQIZwkTaCLVfUphi+
mHWQMubR0GyjFWoUr8qhCWMjf+bty7Zx8FY+3VuijX4g74Q1VS9PvEB6t561M1it
Z9UIaTslyDP8j2rWIfjbqlB8I+0aoMsZmpVcgU8XYMIqaFefLfgHYhkrvOBXssAp
UlU3cZerRYg3SyqrzjRHMW93/2KVXy9Z1KjVv3WmdznXO84w/e7heszWWY9a7elV
l65tMEJzbKx7pz8HVivBmaIk4E2IBnlopwOoHzTPUiItZgcpY6sgixZjeqC7yd4y
7yUFsz6fqsBTb1HldwO6XXmI/b0I9G00D/m3J0RVuEscUj0lc97LWh3+E3sNLt+p
SCv4NQaerUb5t/q55AXRWtDsNNmmrG2R9F3TwuJNvWvVnoW5h1olEd55d+YJe494
4PLRzwWfGxAJDzMEpDDRLM2trqUmtitM7VU6HL/ws1T81Qx+IdW+I41qektTwhRD
WQ4wDzyIeX7AN71iKd1xX2zYZCrO+X6Ag3XeJucO6VUYJ6B3ic4AGcXRxORmPby9
hu7vS08udbF71NP4zMmGaFGVXfJuug3+zlJBTS4Rdd4BmoXxgNuHgzCAA91ennlI
8+zw4iOCNpskJ3+L7MJ199j7tu0o/X7Qq+YjyJACesUfyki3D2PCXlWWRNU5lG5Y
g7hcs/i2i/QD6Vb8x9j5aBCwhjp8VtAD1slNKZAXd7XkifK+okhX9dj8DnRvKFp9
5em355UXDexHybiWzkE5N7xqjU8RwHuX3xjCoEBiXmpetcs192i6/r8koRClmSjj
EJZ11ixdb3RW9Rye7m6pfpaK3O4c01vaMTaTxeCGqbeNS0EVBRR9iiDsbxBtdr7T
kEcMpVC5zTX/FoRQHzW5pT8V4zr3HnKZ0AzS5SuNJOmKIr6OzznbzqBAOAOcUXFH
3JfMffvuPcO2RMMNPaVKhPTg1f4xYNUJ4toVlZcpF0z5P5EtoHIRzsdgfIGCz+k/
pqWowBm1TxtsuUCuf1croGK4kV2wdxiJFVN+jlmbQoajiuA+feIduTQMPNq1YYCC
YFHjGfQBfPF6cc9j572nl1iAFHed7T5KxyUk7BPnZNtf/NdS2flu8l7bvPKuVe3z
vWIzhjesRr834MfyP8T4VGIWq0ialzy4ZjcfCx9oPhlG/opcPSVVKBhR+nk+In0m
RVYB6jRQePcqE3bBxG/KDMf2h7+K5E10yOR++SGhWojo7+rl+2rggW/j6B2C2uht
1H5je8R4RyQhmV0HOZ7XfLwBuzyZXOFkUlhYHbR7qwPEAUWVw2VJ6/EAnnc8LDI5
J94rwUh4MZwCt8CMfkSH44NuSBiihPIrPKRAtF77Qj5Jg875O2tdZqliiuHod5dK
jJbJfkkI8NbyEcpM3viR/h38wJi3N+jXS3o0sSEYgSeIcTjmWY27pQ/GYyD6qa+Z
9Uj/W4XUfeQyv8fUC6docXpqPC9ltDe640WyIW04DItkkPYvpqVQ8evfVwunOQht
AnzgVO9roknm7fJvQ3umO8Zex7pLwA3rV3TtKyQuhXSnL8tCGxs89h3ncKx1srLs
SKYQCsP6GCDh64Lkkdtvq3DL4b6UwqAoLtkCRMD7msuMLRskCefYyHSDAuCHBt3s
Ew8aSTWtAnJL5LlvwaF1f5QL3qzCDfQLmxY8sJie8qGJv82zvWA0T/fh7sRN19Ir
cCSRloCEvSkU/9fOVwR4p6iefzIujg/KRJK5kYzlAD6msYLZT7ZvVpJMQ70cQ9a3
SphapD3JM9p7wSyIGLDOAz+OJ9Vo6zYyQLvzmoy7MVZvE/XzgVR9JUD7O57uGq7p
wcyaadhhAvJ7guD5Ib4oirlJ1e0GfKDGsKkQnB/PP4r9xZgGjepCPSodIGvNpTeN
VylQVt4LBunhX+06yRomQo/O50rzgHZPrw/Fy2y75y4Y7NsNecvLADG/b6SPIa3y
Hj5HEwFkT2RVCyeeovrAhTw6iqtZRtc4eyRxhAv3qNaBVdkgBXhMRE7r9T39cyyn
w2mcFnjCxO7qcCCx3U8FYGl61eH5cN4CFZAXe2lMXREPKTL+uWEET2QZJKngqNX8
yKV6Gml9dpc7IT6qkyFl9MHUT5Go0t9NxiiYknCP4WI6Gd49DntiofNRzY0LIQg4
hCq3SeOHIwyp7XV5Ul2c2sTD6f6GjHLfKDPqgSg4M3iLFS1fp7XU9c3QKc2I0ezS
OG+tWAPLtlmUm9TkoV5jEnmocPtEbtrnwXbqJhpMH4IQcNck4jmfFuIV/DN3m2dJ
b8wTtHw3dabxaeNOjsOZvtTl0Ab5y9w33COW0BAtu0BJhiJxDPRTwjVnx5MOePny
FXk199hItQI+EQsvtOHbUie3gr2Z1+tWQ+2iNjm+OkmnL3FjslugsDBVnAHDsjTi
NdadCYLc/Ypq4kRboUMJRddgnSiOogcG+m7AVEtalkvd6MSJKySzdQLsR3kCD8it
5PVZB5Pxrt5V4PmQZrqTtOqGd62GjxaYca2Ukso3if8Aq1odi3MO9+ylg9T//w/H
D5iihYRlJMjC8AG5Uef0T1wN2FMnoBDyr4av6qbVr/yxdUtcwnQYAkZiQEebnjnv
KyLeznem7s4mkZY9h6HqMu/CbLJlm5J0nqM4RwTvSm631gCRTngALD9QdC0a5/dD
EoMYSatrR8r2TgrPEZlBnpqxMP9o4pQCd3fdT0aseyrLCi2M+VfiMycPIbApkQbW
niOqPDFsrG0wSvpWeMec/NeJ5Lj8/ZTMYoQYiOv4kuqsFiM1HSaPnVEzJu+GVMuO
hDmB+vi3xVUDsMBQJMWZ8zn/gngt3kiLj4XX4U+zATUzD1Z2VlQnhoHVtJXyPtbU
ZysxlxCCc0vIszqEkvmJTSJ+8PF5UvwCjLeKK3+F1+7QwxG1D8d7Wg1nMbVb6U0q
OkmxUJgxIlM70PRk1+EPQ2cq/w3W9rTEHJXHsQ+2utgz2bKjDhcCKeBXPtf+Otxa
4upuADuaCG4/ZkZd50fscfLnnZ6t3Ov/i8Q09kwrVJ2X3q74hD3XSV0O7w+JLbgi
V0UN6qDAbEPG+1VUlpmi5S4t7Yiuuc/gwkG3f+AK1CLlUaA8J9A+vhZeSVpehG5B
uN4LnCYTIgWvc1RkMhVQBpavxdz8sh0sHzsUNFA/s6kmV3TAoMJtRl7OlZ6sUqLu
oqS5QqXgGkuFFF7JNbyMXz3/n8LUjk38FXMxLKqTKsUBSXA30ECyTZBcZuITzXz2
6WUw7XGt+yyAxPFHW5vLEz8CwRMLpAqErfOeUqttWFc244w6UFhQzL7OMvHJBXsg
621sW7vvhtlWRm77M5L+6eAPdSlfz0xP9ByoxhjJd9J+pzOgiKrCtzbjCgfdAlo6
MDn21rY1TNUDvaKEcy1qEsbumdBuj9SDkbsj8PQyw7MyY5onUa+3dGinA1tar17M
logRZjz+0tH/pFeFnQblERgQtVpaQpydTnG8OZAX8ucYYKnwjCA8Ne7BtCHXeTit
WU2voRh6UdnGP1Q+cCTW/AJHoCJuTIrq1dzkHfP1/2Zqq3wK7m8bt1J7QJ5BlDuY
3kodJpZhs9s58oaOq4jK2uVZTt2O+gP0UpER5qTUxTM3gF0Eo0hn0cfyBVRtf61a
DJSj7eddCAEMIvciUWLqd87yIUt8Eubw1jVbowTQeYGE/7T1QH8Qq4rksjXw/qPn
F8bGRgFb8SM6tDolSEHTbI51Pla3pO0XjHQkknth9E/xoX/IJ1/iQGSvEvwNuQg+
hRT/AQkb1VK6X5RnQqZMLZI3Yg95xoPSNmWOwjD3DTt2jMyuyQ2ZgP81GIBFMzw1
OAxSPy6DlP6y11AZD1G7fvu6EmGyz+LTY2qu0oK+bzazds0NCAR9fkP50oWzkcPk
eey0JjjC+24baza/X6cqiDz0Ui9EInfXqm5D/Yc+SLo4+KnFdvgJKtXQ5K5sib0J
POuLFfpjMRqf9EuvgpiCAo21SAWsCURA49ONuNtxhJt72ThF3I57oCnreqKNyyp6
YIdMS4oJCS8zP2BMDDcE/rbIqkWXWUeYLk/aUYqlb0LLxP9gkynCtsrpwGivfXLX
uevaO5jDxbuyQoauxH/RhW0a2589aE2p5PPmcNqWPs3AK1k+KY6kpqvxuLnS7Khe
EfP4wmi/Egu+04RLmQF7Q/FSgh6NsiWhIgQf5xXl+GrSqR8XaXyVcTq88PZLxKPp
d/RsqHf8KRZz/WmfWb6GmfvhP0fr8duKENQj4cEBoVXFnBnWncyM5tirs7BCokib
kZqDpqWx3eVWubowDV6BPcfC5hUdDpcsKgBHGltwMOn1zyzCOVyEbPQLaHgJwvA4
WhzLQVAk4tKErwJZZaQOQKeDenxWfmvVCIqlyMX0Z+45m4anFtsoh77nNj7wxvmT
9ioNMr4AyoPpL74XNV+JB6HjxnHw3rodd9+0Dmp3PYoK5QIZNN4EOF+8TscFgkUk
iRkQB2ao24oG0fPr1D1YPsSANcvgKzaSG2z+Sol11fFB6JVbhQ9//mYi8usxKR8+
qgIzCFVbnyCOzuLMFJvvmEk9hHOB7GWaXA8Roye6Jz7ebuvzkZFSTGg073ZLcs6Q
Ed/291C+XBoc3VsvEWeJCqnaa+yvKyjBYPAw9IqEVY+gJYm7IC1+qDzN/4Loq2Cu
0YJs+IeTgwwE4BzW7fMFAN/PAUbhlvtUTUhqmpjY9H3OrKM1DAizwaubvlw5d+BK
PqzYphXx/YXO6m9e+S6ESvzjLEQPcT0a8SSU9V0r/kRp6Bi42bTlPXRA8u/C59Av
OZ1fPyJ5vhv/teCtJaf4Waw/Dj94DB3diB8c6C6ePuGVR/Ky6tN67ywAM6KaVhLP
pdjD8Fnb/nLVZT2f3QmyR5zP0p+vcApVYVU+Qv53LzOOmtiRyE4UteTPRqPgpCyk
npcOnsS6UObmECwxsWvl5QfuYbdKenNjM2Pd00rE5CLV5tNQ75aGAT8fhDz2AcQz
41VUh1z227N2exZtoaRL11e8D8nxEfgVYBvHxplGoNw3EwPa970c3g+hyLCIBk4p
BUsijS0dqhGG3kHOKepxbIJbCrD+JvLpMJcn27w5jbjoGKVN2UntcTjJOZv1uMPD
xjm9G3GlPXZi4F5yxUa6dsUSScGxYnnHyq5mpI37ZtwrWJkLYOX9i5JaPq2N7opa
mLcLHJvaeYdnZeIwTTyEYQ1sdc7CD4X5G4iYDau4/a8r6ZmNg91+P+a9141/NBgX
3ouTZl02Ecr2pNNs608Lx78JKJDOk7FjZmbbW3ohmcaHPIsS405gASQ0X8M0A8wl
Oo8y82jVyFtvV/NP/VTGRJ72CUtEYKANPMuayl4qX13c2QEQ+KvobixpNtrxtoqW
RNFXYBqWVTfvvmzrdG5JjK438gZwgh+41Roy/YFE8BQ4m9rUeLvxbnEQ8FuTOEOK
qnDZ1/05WqZBWxEwwtUZmc3K+VzArk0yFrvAZkiMBECDL9AIAMTV5LX2qoDodqcG
lZtyqZRgNsAjImqNixp6oRojsJB1kR/tZmRB0v7GERoTPd7lUc+BqPDOn2IyKhQB
gjdOTsFQxcvGFOJoC7GzlC627Txht/rwAMfSKHsncJamDmRGsa1PceDqEcqbSfWD
3W7SQFPhtcM5PzBGu9nVcewo+rL0NbtBOJNDQdxI0ahfCQSk6Xq6HuUH/4JzG1jG
zpKsAxbtJOoRFfMGjtu/mnm0LfanKvgPVHgXju4K7PhjeFQAKPuDTWFPEFTw5NSJ
kp/UTEcvCaLbivdtpYl+ztQL+MB7/iZzow01MNOMo4uaJdVTsPiAgBcZsxnuMJ2g
JfGxxXqHHmYxA07LD21jw2Hym6Z/JG3RtsUVyARYb+r0Hpd5CTu1f6zkxRiGEK98
T7ccKdJBugvYIDR0+y5EY89GSBHyD/yxjOIp0xvaBLxIXnFgizNqY31j3okQ1ZlP
sim0+zgD8Sw+L32FbvKvSpCtMqS7yGx8GjV/2+0BzbsIyzCHKLwhbEuwjb5sjABY
AbUiJ5BIZdZf38s7xvNcLpzkmiyJ0sN9G4KcHNZukA1ec6biTIIFXJsPZH0zvQBr
riCYJMueZxTtLTLBGpJHoXOmhGvntEBf2NWMMGNGAv4NTNYhBjkqOV1t41ZJHxF2
If0Sd+35+OkvoOX+EKlqRO7JIbeEoZ/AX5C/CSLv0kX8pwYb4TUiUN4frFAxp6+8
d6W+5yUNA72XZn4vbuJl+36w20kHrNMWOfFKhtxidAjqHx1UvkJe6Owxl9N/XMUm
qtELfkqyFp80hifnjx7gYiqOm3DrawUXMcRMDVXwu3ZBhgLGtzhMkHMn4STLpRHV
9qE+kgpQuPLffjEaNoFt8JL15U/M2HVEnh+YrargDTb2ALZnVMKDj+1xmAnhUGcT
05MthF1RuvF0LEZiC/yHtIxnA09FjHcT1o+YnpLvIVybUD7lVBTwT4O4302SNoES
DhmH51tMdQymBnqUkbu3X6rlsxSdre25XOVSSBvnGB+6ea8QXd3pN0qiwUyXmi/J
KLuSNYKK0UVrs2dZDumF4NFtM4ig6Dlb7a/qCnn1/EP/vleqQP++j/trAm0ig4Bx
LRr8+OXXXDNNzPXEJu9/SbRBzJqlXrgr7pV3+UAPJdwuv8zBl6QCMP6KFuyfezaT
1SAk1AD3h5ADT/9DLHqyAGlyK2yJS18fjbTfK3Dk2jlW+fO7H4Fg/wywPpKj6dl+
ywO53lfYtemzGVRwuDQJN3fmeSZ+D+maJfNUi0CC6miNYgZDNdWmDhJivPyQut0q
JrDeVSo6jnsycl3UBRxwcL6FAu85L0OS4ljd8Behgm9YIINavEliRP5qBVWL+pEf
dJuIdM+P6JKO1Y7+PmDF7bn9x6eSTmqMFFNB93jT2s9CwGeyvWsyKyZqMNUSj2iY
bbezaDXWPEVKcYhT+SVsn3pcNf4pXWuBcU7pMgVK6Ceuc7t6j/O2KHfnrst0Jml4
LBevKunb+M7rrJek0tGv9IexmTrg65TJ5IIt3ajCkPWIfP9jsPxI/It0m2ay2hwF
xthOCIeXoGqCjwyau8tevDZXjOCkcAeGPEtUZWSF+YKAEtSIz9n9UFdriihlx4gq
cTF/5B0xfNpLdon2iJZlDItB0enQGAaRWrPJ6d5NkoWIdb1gFRnShxIiV/ySrf1S
t2a94UY5OESVV0WP25DRQ161zUEn0up7Py0lsWTT1cLcQaj+hJkruJE8+IcKVbYB
+6L524qP1d+ICDnTPl7pnPzMTQaFCGAsch3kx+gUHxoM2JkMlRiyKaw1pk3wRRT8
2Xqvb8fucG3vSRz0sMfK5aU6HLuMznSnOQZKIta4ix195bm/Cx3e+7uKATgnKsrx
4Ov0HsjCiOlhVXJc3a7l66i8qnI5DyY0mdxslVpUhPv61PMLG9l05PchW+2ug5bj
3QZiroq+pQupDpVBwqmmsB4oHxbeewqeOLD8JPL1qe7v6aUq/3nboz81m3J2q+Wo
TRhLRnrdVIrvZNFYgnVdaxV/1Wrd78f2ublY/gfuG+PVDhcWMtWEGXFZN6VVq1EJ
D09zTAWxPZO4T/aq29iPY9N8Yt2+3Nq8eY3iiSKI6+KOU2h1LNodk2EErUYwCjRD
Q5PpMMoyoWfxLlQHir0QE9U+H/6GLC6qWBl1Kq7zIOI2ivDGGwdGMRbyZmT8Po5U
Kg1ayloZUHs6BQ3UKDH1LGtTzdWz/9uAQ8ecKZhZP/G7QJJBgrdmRd3yY+AzcCQM
Wz7ml3J06Ya53gw7XKfUI14MRjjOBX82VAAuCXxhGVjZ9uv0N/179wTckfUKVykW
4vy0Z3+hS4DwH4L2y3858dKHW7SRyUPHkNBkI3m9a3hY9x4ALrcBwnl2Jz2JAZjo
plVoSL30WWvfs0RIKY3qnkqwayjL96U5+9fpVJoLhvHTfUNVE68U0ucN2KaEAZOv
pUryvQvnTk1/bTvieOAR8ztbfPVWnmDS1kflrHbM//Ccq7g3wRra6Z8Jv1XyaoWu
ntJMQQAPReqobUsUy+YLzDwuhjqEVqHj/71hDPJyELXjUdkTPQ2Qt4WoOjEghNoq
Yj4IpMBHKdcV+oJuI2In74U50/hCMN+nFQ4bC/V0c9t4jev3KNTNG04Y/LSPcsrk
2cuQNz8CLbHh+71TEXBNFqCaPRzrLHPh2xZoSmgNhx5J5yKiQgUMeBS8LSvdbzf4
g6zlH+pn4k7Y5Ir9DfILEmaMmWkR6Tzli6DTV59A/GRK1JoPupbB7RakxBrQjqps
cnCYjCe4PdRSRUQT4m8r8mHmenv3vO+tJ4hULDGJVcNPryhkH5okJLmaDA+hXqkr
HLFHULn1fTvreCN9oEdcGcuxpAX8EDtZpBuKjVkKeHTIvt+jjQQG6fcxz5FmzDYG
Xp6KXjobzB7Jt84e8bayfNVqNeWL4FTAkr4vhR+mXQG2sJW40HqBz5+nhNAcbCCF
f3WKnvsLSUuDplQW7UBvr0CiMnguiD2qwBJW6vO8F0LGBKkK20ia2Dn4Vn/ejpg3
N9PDIqVv6byFdXqzH8eLdD16uCJN0OOCWzvmhj15bmVJBZ7afR4wkWB//w7Zjhhd
kx7q33+s15fPbnobC0GpWr6zvUu88rODgtUX4nTPtKFfgIgBWuLYhBAAUaVzuCvl
CIOzhZuhVITiy7GJu0zE7BhzJ+u+roXH/TJDPK4gFXhAsmr0XwsIC8IlcNYhcyKx
7kjwvivvkeUTO/+4E2aXY6b+W+IdvPHxRnCL5N55ry2iIhBLweFMdWURqGoruk8j
ibHvE2go0VJ+RGnzvuwndaIRw+84Z2VT4EHODdaNk7yYwXNAwe1XeoZlFxzhU5Ka
viCJwj/BaG7emU2GY0zpBoIyClhK9JaRViXbuIXrpz0detYZH1RCKPlypPe+IDp2
gB5JscDuHXgOvE1AXzyzE8+mvvOBVed8s/DDNye7+beY1wLP3es+C+xB/DU05D4c
TMoKLggK8WyF00msnVdmQ7QmMY6lCiqhZDt7UrEGrH+fDgoVn4t0fegyxFaRo0jZ
qbphfUglznFWVktXN1fwt5b59SsHau6ecPkFG2q0OZ7Tc25CE6ucBLvBoYXKQ55R
x5nREPmlcNwmxptO/oCaJEt/5m1QbBgClOYBKV+MYQjcoUPoJBKcD89Jgg/b++7A
F8BsFcdcY7XemDbpTnTKyyoCx0xbJ4C6D3g2RcDSpxMPsdutFH8fc+TrxDGvpKTt
4o4bzt01/Xa8OURGBkl7Ai/XJuqV65ceJRcJPcriaMZRWkjb+g7qyvexzstE9X3+
NlQqh8iTS9nFotpHEN7m22Q7cD+vgLW0Ek0AOKu6SoilwWwyDYZsXRDaI9QoQsaI
355mXM1PehFdIJl/FoGxxgAWbpaVtFA1T7xrucvdKFK+Cq+iN3/nR9+w+z4wofY4
BzfYCQr+FfG9AQVe4/5ZScZLppm55i+lgY2Av/E/WJdIUWOfF/pZqF/3sZjuo1VJ
tOPnJC/6W13qLIqkosdvS0II8znV/iYH18vCiujEdSh4IaFI32mL5IMkShRH0M50
Qh5DMl+dsohfvZ/Zl5AM7IOk7QWmeMUVKhuIqN/VwuIBa9huo37s3Tp0TtsbXRlz
vbCLkv7kQA2sf+2QawET9I9S6vMOcV098G/LKtaTZuUCXsdQpHO7Ebe7/xUcYHX9
GuZFI7SZoOussRaDKzbxT6sUTuDE1KwkMCvD/5VflbpqJKvIjxphjfBtFa92RF9B
nR29tff9oEsXFEfaHK87XdQh9HdxJfASEgaEMVtcCF4BfRZURqpP/3FjVQCwKpxZ
C77MJh8pAFL3vCgpzJZwbpxqHtjTs+vZ3Y4Ldcbnnfoj2k6QZ7Ba05cEQTBu7Qkz
zOlaO/uRC9gGrrfp5jNOKvBBCgys15O8viym6xkKLGXqWSY0X4gqHIuW+kGIAJ8P
q/kgur3XWBQ68JIiVjr1wSWwIcOMgxItBpuHU1cfCZ5Kg6gt84t+q7VS6u2MKtBm
i2sXNggtqRUXW2T1SDwKAVh6OMz5HYXKx2C/EPiNW0tmjOjb1F/A0QTqI8IghU+1
BSO8V6syan/2fp5gWYEDzI6/Wj31rsfXoP8Yn53wzY132AwkdSmje34a8yMbypAm
LQLVph9NWVX7mMeDxgascn8ym71dRz7hBIgt6LJwE1s/IH+C7S5OX20aIHID4wiX
rXiqRkHQ3srPppsjputVWi1DdL3B0uOxb5OoOckTPUrTPcewuz2mXwRH2OskAGmh
R8akhZavRFnTmuLPdV/RYZ8YWXi85Iil/DaDk1FbYGprrbC8AagCUkCNvtjcUDwy
ag/xsEFJ2QGQZakoNGx6td36kVToZvaYK33ay02AV8mvKyAKGoeNQ9LGDntWqHjb
mo8GmemDuTMOzRN1oqxsJHKAdx9zzPt9uTLDxHlCKkLW/VeaReoGFJtDfFeN0rv+
3kM7cWe63kknw+0pYPUBjr/SKCG5o3EpWx2ooy7Xa+dHifsy4A28dXvNRJNiaOPE
toGNOTE+aFQaN87zejfrh70XeesDl0rdBX9NuMZLEyF2mpiP+IhWeUS2s8/qVhxW
TZOIH9EpwrgTHLdtPNSsWEaNcyM7rJdQoNkIy1DXNKqAxJ2e3GCsPaT+OVBlenEM
H52QPE8wxSOkXbUnxFoSZNmkjca08ZAf4kcV1JmMJ/bgwLHCmXLoh8+IwYkwN6pP
y1Z4KW3eialf4LVWIciw34oZXAblblxsRaYsgIrdZevHnDcxTJ7E7gyt3DkdwoEY
UPYR0bEphYj3DzrLvtyHJi084xTJzJgFzCRwZjQx3u+cM8OOaswbUaFwKrIMMq9f
fTmNc1XLt+CVYLRwlw+HN9VUfOno1w1bmxSznHyVJDDACjlZ1FRAsT8uC54iL7qf
3gxOnaMZCCyETfrGX9NxXNVMwWOs8ec8HNqxRjxr16z+mH/BFkW6NqC+3XutyHNG
XjV7QYwWe6y5Phqq0qHheU1HIVXc7lDCJ31ms7EkMnmDqlH6M0rTDKZ9THRKlgDp
Q3P5AhIPe2Sk9+n9v/hCR7wa12DEfklllVvn0+NUdJVhJ+T/d5z8iQucoBrUNh5g
4q+0alKZJVyjKRdBxR5yzT/t4yLvuhLd5DSPtKXJ6BN3H5IrytQfKbCPavZQk8zg
/f3U79Ob5zCUxlJEIXxd8rybjTyQZzaT04Xss/NQG5lVb3oXahgIv7qhsG4TlTju
9O+vPX5ptNSDaeIUV/WhDRp0cZqfi6PLbfbjR71EKylEIy8NG7yIVlXrbGxWvCsr
uMi1VJKxyy8E+px1Lvu8JNTeogyXUQwDH+wxsvGuPf8fJSiYGKCW3SPDsMUhVPZ2
iQxWOm5IBK5R4/am6F/ne1tXeR/AFSKEgrgprazn0kLV2cD4kTPOrVZsFhqXsvau
hB/yVZ4RDCYbpn23vQk0Io68R6rlzjDDw5Lm+Wro45TFGEsFyd9G3Yo7qrs/VbSO
77sOMePs9nj7r0FwTcIGYXPZtKKoGadlaPSPTN81gY2h6mPhVMGA9JI6n2zc1M8b
lTBrPv27dAURGVChB6oHneR+lef4usKGwXfAJMtMrWfgPSWMOGZwP/H9DG39fNZh
TtNrIgm0cU3UjNe//5kpxkgo62J7wArFHFhBVLP+41d7fpo3x8cfwU4ptcBZpB72
ie8Djtz598bklwF07hxbqqeMPmh8mn79HLdwvpYOcrSqzVz5aM5+vpHPKHQ6CHX9
pBhXaS3G05K6IokAMdhoCAouDUwL8cz9u9mp5doDllcLGEVUAtBjtNW1araH3kh5
syQXbxXzwYBhceKAaEaJax+2BYnyuPOdHib7MEdOvPhpAIUHiqp7j4ivewSz77aR
Ymur/gmntekMnzpTrOYeH8NlX+ir3izC6qCKoCvEYBaHk3HQQfykYfEVH6ZH2dBn
biZcRmt2Mz42kkKczQnTmabdSi1EXUAP7Z2bT+n5a+buPo5fdAFmarhiBlSOwD9i
+V5prHHxQQCRXvhEtGzUxJZTechz7fTvXc7tC31BOZKUlbr4aW2xaWmRq+fEVzud
YLomgP1G/g0zGMPlV0kPnRCE4j/yzCltaxqzJCX1lHHmdISwqqgHR3p82NbR/DVi
K21m4QN799HjbhbOtR1m2Ay34Pm9XDHNOzgmqPiXOS0StQbWr3Xxle00Tn56pd+r
+XqkaG6ufqoIgeORRkFFXexOV3/pLruXFDKl4u4nrZ7RJqTMMy7Ng71EX6KR+sNI
X8k5JjepU8O0wvpfyjebiBiGwLLx0Z/vSmBu3Z2ifquQ5LUxrTgJL/usxq5FaCEm
9X26LbK17dEYwMP72ryjR5vZL02jJnZ+IGh2JFGqFPIbJCAQGXyNP0lHfI+2p/ZX
bnlsBbvXyjlQ0Hvv9xATw6WjhY3+YYSapAqI4xSlXy7IgXDoJTejbUbYBHIprLRt
zbVCkM+dEuj5MjzmTgrD4Cjg9eO2MRkLSwxw9J2XSq7HABbrUwBu2B8SFLlm38cB
bpemMM334eL+cnJ96RmQes62nHU8EDSaRmBgSRxM2ZeHgKYP0wnZ1YZ6NGe/ezn2
Hf6QJZyz5B4wuFLPuEid3IG/EineNIq5HwkgWyZ7cpKYjWIhAFgCizDDPjgkYjmh
9ePBHB5bnsbahG3SUjBe/irbKkscWoXaB4iEx6KvsomzDAMXtGC8FJW+WH+PbbpW
/jy8nZp8jVFAyYXMmyZduRR+0sBAed0TfBLuZOZYJmN8DpePYioqVjDMjExYoiX6
L+qR+PRT7R7VAqHLIqu1fhQ2DIO6X5TwT4VUZELgQUEaofO/T0bU0BdA6VEVSnuQ
sM61DDJ2zpwQPratXAOuMxEqFUdTL9LVvOVGH1HO700znRVpzzC2SSX1GNnm52Ou
QqWtMNlb/sfbZ6WqaYHfovV7avSs9+CE1F51jjNvB64VcC32Nol64u02HOT3af0f
uRDbNBxXr7egrip6ZPVc0+pG4098ZTON0tcbt0jd/itPkbyE9Fp/hSq0I7xlf/II
Wb2Mz3RT5VEvzFrs4SOCJBFQ5hu0T6ejbXRbM1vyhmAq/hfvcJgNAs0Z+QU2e3ak
QOsEIzpSRG2pM1FuGKoMoJB2brOq9cckmCtZNxho7MUR/UwUe47jYpqpsqmQTe0f
yEIU8BDOTFG9tDms10Wuh5mVfSvKzIJdWQN+47EP/RHkyeamJctTmlpudMgu0STO
/uzbKqdwnbSIC4TM4NrLx3W6ny1xvgRyIRSAl+JfCMoyt9vo+aZijlWWS11Z9MC+
C9IhvxE9qKcMtaXhVicH6JT9Cdc7umtXTlff4NucHROBISykLF0rbE4hTUX8AAAq
VIrpcwsWnVA45JdjVmSf3D3UCfKWw8gYzRVkl97Ep1rMxzb+uU0ATNYDy/Fm2PVQ
0fa0lSMkVY/I/QczuuTiQu6jcDBWiAFRLNSjqmwKAas1013YFHerUun1b0dPk1Ny
pCYxyIMUE6PfeGy5JUK42hbFNCCp53xt34yUSCs0K/zwzxa+7N4rdwxbRQNUDTdw
ZvvRj7ZFu5KKqNE+CQCDFswXkw0fJLMnHvzbYbUr5BmWhGNVwYX3TCBnkIgUgOu7
RsmRbaQl0tcl6aMHb2cLREaD/DYQaKI2Zbkz10h3Rg1qhChghUpIuw4Bi2TGsZu+
oqtgxK88AWZYlN/EvJcvaMLpp7ueXoZKUrDWSUTCDPVXUjp9pJzq6nWHt/kgDQTW
I66+gbBnhVNsvgY2gVgxrJtUwn7IM3/pvL6rXWbS3hibyRjLoZjoX5Bh+505ZqJA
zBVXaikE8mN928XmE0Gd4/WYbcl/gxCU5j3l4yx373bkiDB8ODNxfVkn7ECDhPaW
eovQh9Cx6O3VrTXxeDi2iJvAwBDyIOetOLBcNabktM/NYxkxoy6h9HK2cYnSkh4+
5ub+beQ6g50IGjtxQtILfQiNABdhn6G5tQxA4Emmc1keMXhkB4Ki1QGoyEGAS+O9
Xo83s8MBNKL41XizinZrBTXcN3lTSjwy41dg+vfgDXMNRT2jnc0N074kHjVNrjyb
AUXf8xv8tegr3Ik+cpwCNclY+2Qe2uNI4XT3fdsdoIbf4gIlyedX4Y94FMz77rA9
bJtvA5jVgw74qRtVO2Z0fH4UBJXuACFmho8+aIBw8npvyfsLEvJDJA+IaOSYtbsN
x564hl2gJF0QeFb+PCYXD/ZRoL2FX4jUWx5IGONiqBO76ldKjKPDHLjSj48dJjpQ
o/ne2Bl6/z2vscolnneRgVcW+XGOcGD2OQZDSlaFSQHNorf8bRbQtNcEC8vKC9ZP
UhHhQMoCvMKcP6cbHCR8drT7artfPQayxtIQrOJzVFSM2h150llFrCiPIeb0hIrZ
WE5kyMEaB1Jg+JDat7UMWlwsNTbSy5PPqhC3/jfn+BLD26AbMCALbgOFsQ8AV9rp
oqo89yClh01iUwVo+Li3X1muXinWa7zvNZ2gt+gCZ7B5Np30EfWoAvR5p3JKoYJj
nG8RggCxQjNJnH68KcvNQd/MiQESOs74WL9IVBbT2EuzNj9oNY2U7aYvtE/jXVFX
F+gX17rQugQqXslxNaa4+uhunP6HCQM0bracmTQPgMT96SrhVc1OizLG4tsr0iSv
TB/+35slNCp+PTqDsHYQ3Ao65EaM4Sq7tgyjyIhAlQaVsF+h68SYSCxVXSjLZcXu
psDSLSq1BswCOFnY3n458C7SecMYnRfFozqUkhW7ahzOSbOuYBN32cIP4EbVGt8g
msGTjUXdgJpg0bCUzZScNfUtVylTw8v/V82Kw5OIULH/jEKdwhnukYZsrsg26RdD
OiB1VD/BCzHOHz8uMAiKzrzROdrQV7MbBZpaj3QsLjKoH91Aww8TZm9kdx19NSRz
oL10llnj2ie6FufFyHb18USzgYHs0GhKDBi3cpaB9644bH7caRHDpXYSivls4ZRQ
DPy7q3KyH9CzTbcctxqXJSK/+X9Mw1xeigAfcDdfo5Ud13ZDMqCCep3Hf8Ir7OhK
Mpjqo02RaWXQkb7B11EEz5Coe2/d7Qet+dWiowOL/LxZynIfhcvy+1id9VbPSsME
LZZoTh0ReV2TzzY0gpaXWKNpJHtFnTF/8XeC2oMJnsO/w4I1oS/PHft5P+5IXeIR
yjs0XNozgS4dSBGRI0s3+7xJZ8kmPmGQouSDI3vBTgAaRDo8MaefzFGImWB2YQfV
4oy6vHM3B19oxwoaHlRP1omxF6v805COgYF1kCKC48+nNltlcny5fc7Dwfnvsj5z
QItG0GPwPXJYnNlNlKH05BJzh6e/TH5wGGZ/yUXhkH1xo5YjObz8XDRaaP9DkYi1
bDUZKsIWBN2t3IoaPb+5YrYkPHfE78Sde199aNkBW9mTadALNt37Pj5XSSxIoeGU
FV8XPJr4gZL4wKZinpuctFcj8q366nEC1PHkwvicE0xj8B30iLeWQeCD06medhQG
3xLHe4VPYsO42c+j7FMN/3W+6WekytWVm1TLzeWH8j5+yFR9+TutlI/OHu6pF9iL
tcNxLgBMDrm3eEupV1pg0qSxiSD7Avrd6WyUMCeaGeDTIMUcNlRj6dwV/fRhUFUx
lGK3nUJzptBxUWneYoVO1R/d9F72WWD9uq2Fc3FSJykpnisGXB1qvRKMQjDFzhC1
a+k6SMngDtL91wYih/lSD5h04OWrqhyMNUrqdj/J2vMDnFLFrrIG39URDHPBYknD
j+lLbroATvHtLgIq/Tqu8sC6qXX8CQPWR3wvA7noPcaSL/T+bRhZG9+fQYODWqaW
qX14UtyKMZtiiUjXeJjokwYlLleTb//mo6XisU2oktGYXBKlWol8T4bbU2R6hbT3
/r7TCfKWRaoOaloM9zCJnuG2WkVqwmv7bvhII9wjGH43vgidmn4avsAzdNL0p/YO
f3SEEV45Kujicy+FUuEX1NFi7hMJHZP+lw8T2dEuGk+xhK/szD9buHe0k3ITwfTF
iAyM3RVjgjq+aa2S60FGhQ==
`pragma protect end_protected
