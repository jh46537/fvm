��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ5,��kF��#��o`�Ylw�ve�ѹ�}��'�?�|+@��D&�l���]
�>��ݖga�ec:��A	��gG��T��j)�����R͒Wpq:-E�e�g�vd.C"��?C���-C���V��]��6�>H��nj
��1�|p��j^��@��#d��.`�^%@���*#�'d#�Z|%�,G�5z61�^�r��Ap����XxK?�c9nȏ�Y�4��
dW�8��u�8�ud�*�������.^���(�)Iqv���h��q�y��'hVv���%���i��K�U�&-2����٧�?s�P\m/x-e��\)���b��k��ׁ�D�GT&H�ԉ}�:(�B��C譂b�k��&������h
����Y��!�1�E�FL
���x��*h�^�� �^��u�� ���D�* �߲��܁2q���{~!����10+Ɏ�7��h����b�e�{Gݜ�XmK���$ ;���@ `Ԕ9]�ț��E`
Al�o,�n�u��$��,8F���Ȇ�I� �@�Ј��g���ш&�j�s���A�����V-��3k'D�����^���W��Eу=Z��,:�l6%K�jm|uUKU�;c�y��y��/�5��q	�1͸ۏ�P�����\�Ul���A�1�B4o���, ORԘ��o�]�6���Vj������mTLwDУL	y=S"���̩���~BѺ}�v/��%����O��hcr�Ē�C�cxn �5����g��� �c�`ʧ|ˡ�C`��U`��bT�f��}�?Y|F������nq�X�F��1�B+>��b�L�!��k�g����ևF�	�+N��1���K1����8z�W�	��E�Ir��r�
�jd�P}-,� O��'#6S�����U�j���=yy@Hs���T��k��Y��4�T�et�#4��A&�t�8lY��k�Fo�>��~!����(UNC����|��h�A�~ЪN[���G��z Y��1Hh3	*rX����|vڎ��ܶ�$�O��y��s�f����{uY��JuA9̓z83��I;�6�U�L���*Z=r&W���0b�k�q�{��]!��	�n���_CP�����@Z���E��l/�����R���\��Y�R����C�u��cp��=��&�o��o��J=̰:��4�)���
�,��~���0���IO�_���B�p��;����]���]xX����d�C�3�M(��+�~��X:rCxws�"&̾�1
81�S����`M���l,>.��	�}�0��\3Հ�w5D	L���0q����F�
>{X)�hD����z�;2Ԟ	N�����u_�3�3��� ϫg�fς�J��o�DY���X5W��*���-	��V�U�N	��W�����%��x�l����ז��^Hjv�����9�f(��
����E?봌� / ���6���Ee􌋮52|rҎZ���{j^ZA�y��#��o }6��7����8M��iŋ��C���2��n%�J#oj�G.��x�ѧe]��G���nFA�sK�k�Q;�Tl�O��Y��$',�����!���w�J�N�Q���nM�7&Y�(�s��%$~��_��X������@W=�4�-�&QQTAպꫯ�;˹��ڧD�gh zY���Hj�*|#O��!.�CN�
�W-+ㅚ�̲�"��<ۘ Z齮	u���q����R"	��LD\0$�@������c���� D�'߹��6��@|��Nװ�����c+������������3���;�s�)�|l�3�u��ȱ���G	>�S2�uʊ>lB]���s����[>�k���ǩ!��lo������燏�q�!�`M� kz�/$�m'!��e�=]U|F���6U~\)�`_52h���N�C!��m-�!���e?ua�G\0�i.N�^J_>A��fCI�����姭l&�+=��a`��9wY:���!f^VX����w{� �ã<������2a�I\��B��lD����F2����q�B����b��v`��/w�����V��1�6�o�� .+y֐��6�g!ou֜^�ovޕ�D�L�s&=NWe)����6]t2�^.�������#�bНO+�icZ�&���h:��ȥ'6-�`x��5��V��D#��	�`�B��Vs�/�ʴ�Zt���d?��t-N�o�����ҙG���aCS���9�^-|QOeJ}�hw�{p���ǚ��|�.@��Ho��r�n����|�2�#��e�� 
�gD�J숤��D_�Ψ���>��烴�s����"W���^V���:>D����0�a:w�}�X;�W&��4R�υh�m|���Bk޿x���]#�U�L;^*�3�n�1Њ4ɣܧ�~�Ul�]��-�B�u�U7���DmB�.����Dİ+��3q��^h*��8��0'��X��ys(���������R�� ��ۨ-�����b!l	|��G�w��uF.��yOS�R�F)0&� ߃�<0�� �K(��q�V9�j�1j٭)F/�m�D��6�ع2T�K�1��Tz�oڛ�o&��R���m �ܰ�z c/�����nP}��,�I���]7�U�y�� �{(,�Ռ�z�(3��ɋ��Ÿ(z6�����=��s罏�nwت��A��S�ʌ�i�ra0Lt̨�E�o�f��,z������d+Y��')��-�X=8�U"���qɆPȢFY�R�R"�Q��=Qnֶ�#�c/F�@G��Jߌ:��}u�w�W������3i��g��/iJ3mE���-c5:yZ1p�-��%E�Q�;7*|E�e��l���-�i���1��h�u�Ȓ�P�Wl���
��ZXc�M��풖�X�O=8����ɴџ7vz�^���彍WA�g�8�հF��w1T�C���~VfέK_h��lI�����IO�l�!CG�HA	!%��.̖�ه. �'Q�lhF��!�r=%tN]�Y��]�0�� 0!��O��S���
��*ٔ�fHp&��o�	��?Q�ۧrǋn���XD���E���Nן����p%.=Q�gx,�l�:I��~Rx��|�[��S��wֳ��B_���`���!������ĳz黃����N!�eȽ�����V��d�� �W�{.���PU�?3R#�0���n���`x�t�������UY;��`���j~GDH���_��ɒ��+��>Iq�m�����˛�����:�!Dj�[�R��]��$��E8�ߖ���s�In(��s���Z�ȯ*l�����e5�߉;�;Y|\�����+�S\���������?@d�#]C�z�)H:�m�
l�>���$���3B�E�ͻ�VHB(7��@hoB|P�|pj����HB�@+��-�#޴�	��t���EV{�����l��ۉ�ͮo��RKUm�9Q�*�kǦfX���߇	"�Ru��s�Q%��&��J����q�ǅ�U��@.��%;�����v�;'�3�����HO�'�g���)��y!M���
�=�K���T;�x�q}�I��2�5��ê}�#zРU]���y9��W�,��Ƅ��1�iu!V/��r����h�<�d����<8��A���ڈ�k�d��Ɉ8ף���������r�[?�Z���G�}�]ה��ʀ5����eQ��!����l��F<h�*�w��wC��2jJ�(58?L�� �e��j�O ��5r3�ĭA�Ƨ?l�Mz4n�of=A���a�63�7-��h���.
o���b�bE� X� ��I6�ʝ{�,2���������Z�j�b�z��FW<�k0o��n���<�'�$y9�/1? ��S�዇��4V�x��M+zh��U֢U.�U+�Ҥ��n��A)�e5(��AT����u�d q8�"��Ib��4i"��֊�j�OX����� �A��f�K5�>q�	N�%�4 (G��f��zsV(Xa���(��5x<V��:sK��M���m�Ri*�Ղ(eTZq`�M�$������=z4-]�!�CW�h�X��[K��x�8ȉ91T�� ��j���(�G��QEew#�A���'�<lމ�oV�'B �H#�xL����VfǦ��
���fD(iЃH�=:.5VB��۟`l9�Al[����M�|��Q��2��(/w�c��T��g�%*7N4UԂ ^=��8�K�:��'��}�(��[��G��*��_�U���aO��$0��#A���]� m���Y����~n�Ѝ���0�m���?z�t��
��n v��nSq)��1=�O�1��J�/���.�E��I�T|�M�*L�D%��N T����-)Si�5�Ȓ>���K�#{&$0پX��0x�K�LX���Av����L�P��:]5�No&8�!@��A�Cl����X}�ܒTc�4�Y��E��N�]���x�U7 ���ϣ�k�}�V�MjŠ��P�O*�9��1ݮ�2��d X<nO�I�A��Ԏ���Ԏ���K߼��&�e��� |�ݕ�Iٕ�-��i:���OOQ|��ނL��	�ɺ�<���S�0��!�ߝ�p���8�S1v������a��~�H��\����8�j��M�Oc�9�43��Q`[$��i�B�������^��j΢������^ڽ0 ��26ļ�fs=�Sh�*܂I{˵��%��	�t'`J(�/����Ww��L�x#h�$&Fgb���/<�P#�߯h���W	+��M+�L|�u��=��w�"X�[��M1	��R��^����7F����q�.�!�͕M\[��M�h �
��7'ɛ��9�b����`��yʷ��O�ǔ����sp!_��IB�ᩖa���"c+�z-OƗ($8r��0fZ��l�̓5h���H����7�ihF��^l�6v�<)ǭ����ߧ��^��f�qZɳ["~�A�:��)���I�pZ���dW�l:1��V�TC5%���([����V-��`Mg�e���M��y��t�I���e��b�R��DH��[lFh�QP�STDCq��b�$�0�h��m3�S�m�=Z:�9|��V:�Ǎ����B�mM@�R��6o�� ӐF<�n�>~�x?��V�}m�dM>j w��N|#u��ΰp>��b�3���[L?�n��wI@� V �đU�!Z0�ҏ~�Cbk�ظ�n8AHl�9�J|4��������U���ߍ(�MH,�#��W�'5��/�0ۇ��	�p�j�y[RZ�tx+��r6,�>�7�__2Bp��I\�9h��H͹S�fE(@=��P�9��A�B�5,&L5�ԡ'��Q��ៜ<��;]s���Or���y0���t�4�����qz.����%�a%�y�
}~(��9`�>B�S��
��6;/�����jWCP�.z��c[o3��D��]o�Ch�w1�x�]�O�9A�k�EL
�"(��nQ?�\V��E������5!�����F��\���1��@̿)�:Uҿ�^�����Le ������zKM^w=�>���R�(�QǭMA��[��c,>�]R��fP�V����g/�;�^�^Sr��oWG�I$6�m2��z�N�]�����(��Dtf��O��wVZ ��F$�l`�_��������_�A=��"h]��m���� f��{(��K6�q*��z�M�(@�}op�3�0���
�`,����|Ӥè�Rx����������4��x�!�ifZ�1*;e���.�(1�q�V:w=O��}P����"o��˔�ˣZ9CJ��t��e����O�;�k�9���0������������^�B�yz��<� �� ��YO�W����1��D)i)ѫe����[6W=q�;=B�TXԘ��5�Ha�O�=�W�Q��EW���Ԗ{���7�-��
�NrB{�.�I(d�E�c�a��*�Xx�2=�*v�JS�ވ�하��41�o��?�ڀ���f_Z����#�)���x�'Y2�n�BH�5v�����1�iD 1n�E��nE2�s���e8�U����#&�'��}�;�Em0��W�&�4��F'"~ÛH�?�P�2��B�7�񢥄3mp���R�ۢ	�!���vTs�ɐ�-�'�ΐ�#���#��z9:�r��U���
�����L*����⧳mwvo�V�h���$}=RXZ_��=0��ZbZ�m���	?��5\#@���ۼIK���)x�Vx��Z����`��F�	��fy#�V.�*��*+�.�k���s�"l��9��JeO�����!x[>ޯe� Q��K��n�'(��׼�ҍ}�U
�q`���A<[�	���9e���'�1�?p�8\�'L�b O�5��AA� ���I�!��-Gbs�y��ȸ�%k�����Y
�%�Md/�*m�yo�rlZ�"b�,Pm!Q��Z+��Nj06�~,���*+	?�T���y� z��M�/��
�Iۗ���O���� ��;�^xU\�w2�<y"cM���>ԥe"|s�XQӘ2����R�۔��|����S��c�df�Ę`����\mMh����iG�퉪6�헌9�CN�r@��j$=����F:K��d���nT&V�d�{'�Ke�9�BZ�0���.�	(ZP_*���t,��f�����*PK!�5/���ڲr��ک��Au�DIQ_��50�ũm]�ı��f���=_tzur�/fK6z�H����:����
iu���6c��>HR����fc��)�����+�^mw���8��e�)�B%��*Ǚ�	Z�ڿ؝#�����׷D�hl�Q�^�����zƊMRL�	�����J�~��6�iܾ�R�$V����]�#�h�.ƺ�_tT�x%�\��. ���j�t�-6�_�	ˋ
��7���o��}�zcT&�-��@�0�͍@7����=�b��2I�nd[Ll�D"'�=|�"��d7/�����'$״���ϗ��Ќ8�֌J<Ϻ�F�)#�Հ�g	Q{�57X�����r�2c�%�r���fg׭pk�,x��ؚ̻^
�l:]���{���|�ʀ~G�s菢D����V��:�)�@m�}e�?�u���H��$b��6�LtF|��]r<+��W�)g�y��P���L�)��}������é�N������O���Z�����M�T�����^j~L�ik���S����&��0֎�Ђ�%,����$(����}D�}"��[�L�N����8��Zg//�2Lވ�Ӣ�l7\�3"�h{a��� ���������k;�"b�L�k�5i�B���i&&82��n�M*(��U��:?��Km�|(�cay���`��.O�����9�B�����`���RFZ�Akťr"s�W"�A(�X�(#���8�X;��MV8�7MvϭĦ�	VԘ�X��]��%�+��H��ǟ���J]b���ȏ�������fx����>��׉X����
y���be1��!�ʣ+Y��AdˠV���=��&`SØ�t�j�~���C�n���1|�������#k��n������J�d"A�7e��x�T�D��!y꧎G����L�[s��$�˚�@��\9�3�H�e��}±�7�7���ɾ[/�6.��L�������'b��F���o�[P���PQ@
�"��~���ORW����3J��uR���}I������s�)av�
�oY3ß�M�weh:�6�8�U9z�.ըӡZ#"TH�%秧�9w q�Z8^��^��>N�[�Q�V\7�e�g(� ���M�[b}-�+
7v'?���ЋxW�(��+�q%,�r�u}"������Oʈ�|��M�:"���t���l=d���̭�>ݫ.��T\�`[�'����7��O&%D��!��	O�@��-~,��{��}LN���嫑ѧ�kh����uY5@b�u}SG�H�cWc�s��6�6��Z�Ȯ0$�o���~���������Y������6m�}h:b0v�'�l�>�GM:��{I���:'�L�J�-��<�^��]�	t4+r|/J~�G%�_���#�!+p��g���C��c����Q~F���%�*{����%��-m9"O~b6���<�?��EZZA�8c�LsuXr��-�3�$<�@#�r��V����:j��gJ�z4��1��ܯ���=�I�|W�܌Ґ��)%�rl���Uv��p��2���7K��}Op�S�9�L�ӗ��
Wx� Epz�*= B(�\z��u/�d+��e��"���������^�b�S �v������t:FkC��F~*6�i�F��E5�'eЮ�����p�F���`�.�#
YN�qG��X��g����1�i��	��­�Ӓذ���(i:_�"�k��B�P�y�Ŏ�G�#��BA'h".��p�,/���q��SL�ԭP^8�R�X�;��ɂ��_)���%���`.0ݺM�1���~���@�=�<}��ń
�m�(?�DC��$_ɺ��w��6�/�?(�����`�bv,��4�� �e�jC �>��F��x-�EЧH1��AIZ� ����7tX�!�>|��$23\�TH�G�&5eW��B v�ƪ��C��a����C�+-)�����	EO�X�+�+���&f�<:��;\n�^N3aX���Op:�{�W�3����k�G�R�Fx�,�Zɼ���l��<��l�>�(mY���Ge��l��\�A��H4��歒qǅQ�G���V�/�o�8�z�9���*}�����W�tg��k<3; �.:����R�x��M�ˎ&�33m!/�8�1s!AKo����n�z���7k��d7e�&�������x3)`��e�%�N����ba{�e��A�#DB�m���]1{���S��~��$��i�����I�%��L����P;��`����[&6g�q�k���.�u�����6�Z���]��f2�����hoW剴/�����&A(`s���;%Y����G�Ȕ72�Ē0,Ԕ/?S�D��?��x��u�}�Ѡ�z��g�R&�m�d��.kFJ��>.Z�:���͜*��O�;�!�M���T[x!0⫫!������=>7t�&M��Y��Sa�i(� 5�Q�ūJK7"������g.�>��؇���K���r����*�{�.9�/�|x��$�q��s�uH�OV?��텎aT�0����.p7ZJ%�Q-��cogi����҂X���w ����*�m	�� ��ޙ��x1)�.�?q�2T[����kjQS�z��7>��꜏7���-���J�ގl ś�-ʓ���T�_q�;������d`��b�l�*��t�)�`H ���nR���b�?��Q"�g�Q��hy;��q�
*hs5!HkDl_��y����.
0lI�,�څ|�&�Ri��D�|p�w����^� ��z�O�v����ݵ�u艊^�OR��!���f�WU��r	ER����u�������L�cch��Q7}z���E4_���5�8��Ȗ?<�C{3Tl�(�<���p#ȥ���_���ۑ�����1�r^�ZvIS���o�`^��`��(ކ�b,�j��.q?������	y�����#�{����ѱ�G9�?˚j4M���W�xz�B��(�(J�.�s ˆ����j=�3/��,#�|,iC�:���^�|_�=Q�}Dc�;-�}��ţJ%-�k�ꔩ.�WC(�E=�Ҍf ��Y'7F��D�dT�n�1EC�U�Ŷ��D@�?�;@c�)�j�XҋeX��.�����{[����>��tP�my,�	��i�q�"E:�����e��C��5�r�4�vMB#Mo �;ؙD�\�J��|	�N`�o����)��D*�-x�@v�y�{μ�K8���<�0��!��������;�o��!�
Z�JG�x*�n�f�P0��O�Mo�w���E4;I@�H7�[��9x�@���(n%���2�.0h���,t0��X"�%�r� 2h��@f$xy0���i%�Ó�v4^�IB���^PB�9l
>J����#3*]oNzM����/�2���@=X����w�wS�I�ΚT�)���V�hp�>PJ�*|����F� 4�v_��͒-��ۊL;�<ŮK�!a��o3菶�3�Ї_o	�"w��ͤ#Va�ݍ=��b��A��`�ϜOi3�QR�z�yz�/��/�}�4�*��}ޕ�Cb�~�rph/Z&:W��$�B�9��]�^I�\#�j}��|-�-�(�:�)x��Mr���pe�-�V$X"�rf��Y^�c�&d���.�����1�\�����?���5�Ƹ ]xZ11�rݲ����M�d+E�du$'>��o����	E�-3�DC��`�^�4���<��
���W�H��w�4�?�r��-l}�����CHKEg�$a���%��pPS?���M�7�X�瘭D�DZ�Rp�l�14,)#<���*��]p�RKW��8ָ �_�`��F(��!����	�vG�����a鍏�WLF�&���Fg
�K��]d�Q<���q�ʱـ�A��-+O�Q�1E,��߹�D��y�{��^HZ�$٠n�O������'��F���@dÙ�P���C�g��p�;�J�K#�g�X}J�9Ϧ���z���*G�����>/[�#�-*���{״���1���I�.�X�ߎ�፰,�M���;�n-�=�1 �3�I.z���wn��%��
��U��V���H]��Dy��!�Z��Bd�.8�X�ً�/4�S��Z~�a��*%ug�{�`3y�W�̢�N�����iD��&�s��C4&r�HJ>��dM�]W��L)!�Z��ێ�j���6��Z�U�w1 �M�M�$�/�Ď�o^w�->Ue�䪋rk�n:��8!?�����\�?є7��s^n��!��h�� ����u~�C�Y�x8\e���'.����+��>����cq<?X���S"��WZ�"Ov0�L�̚k�]�emi���Iu}�~1縀 [y)wQXӄ?Nl��U�Ӕ��bxa���|(�7X���|H�q9|E'(��S������N��	��[*@Y��,/ud�J���d�6�^Eo�[����\�=uS݅�>Vti��A�mj|��