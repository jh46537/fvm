��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���ጨ��KN�`��[��h����z\��Q�ɼ.`i6��f�c���t?^"��Q��Ŏ]�D�-h���N��ߤq	�#�F��U[�T�d�4��s��`ԗαPB�� SE ��i����G�KdRG��N��Ks�Y^�@�
�K��n.�mG��\>S#[��� T=G1���T�/����u��zѣq��s��?*	3�̘T��{xh�E�Ĳ6��w�A�ײ��b����V�f�N��umya�2ܲE����@�݅��X�<���WT��/�����̶���,(Rg�?�Uig;h���4�Ubf@b'�N��-@V���g��m��[��9juhn�NM���$�EY-��N������ty�CMbD�~�JT�͔��ԡ+��t����C<J�;�ud�L�2��1":FP�I��Iq����i7jL �٪��tJ�#�q:!.�8W�-p.f�I������h�|�~�;���i G@�D��l�Gb���a(!�A>I+���z�k,����r_`����DI
������SX���C<��#z��P�z����5yr*�-Cf� �t����2��ʼ`��7���V;R������YZ�*2���N�hےQv��z��KH����"Aq��.k�Ꮯ���p��++�'�Т}o�V&qJ�O�<쳌��ϰV�=ھ�g��������ѡN������M�8��t/��D�	[�oE=i�͈�4\m��i?0K*�_���Ey_��T��&~�q�J}�J}@N��td�}[+��\� �1��ؗm���������#29�s��z�}��t��f��ٝrt�a��Yx䃴����[�����Z�`��aW��I�K�e+f�&;��: ����Bf#'�ӯ3J��P����oD�T�zJ�nɬDo�B6QMmk�Y�����@���+A�����r��X��~�V��!���/>�yޜ�P`P|hEBr%�[Y"����lO㗑���Y�%*۬|a�e	�D�/o f640�]��,%�lT����u�������ȗ�u��R4�5�|��?�p�i!��^^r�;G����-��X�U���&9�ɫ�s�IK�3:�@��r:c0}����6���2��εV�k��;[�6̔�7I�`��M�	"��_��s�+�'JBL�0�A����S�X�	
3��Sg�c���3���3�	;NՉ������$���z�݄�.������n�����H�,��T���u�Y��~����2��� p��?����1��|�4 Fq��r`o!�l�}�1������Gj0��|���!����(X��=#�z�'�k����|N^��T`}��b ��������b��2�d�X�x��lP����쬳+�P� #U���!��M/P��.���z0%]RF��ضx�=����r�&���&A��}�[R-[l��h;���~b�9�I����s����NJ^zlV48|� �G��
#�Ob�����Q=A��U��4��"N��I�Յԏ@�*5m�l��A�t>�����u��G�	�ѿ׉	�^KJu�xh�<�"�#4M ��Vp�F?y���zh�R�d��L�VGz�'^s. �Mo�S����f��*��~FFS u\�����f�L,X��q\���.�ۢ���޾r���T$a�+��1��J�zf =�e#�Q�CC���!��[�8qtD�o�R�<J5Nҏ�}�j��ZX/!a�o��)
�@�{G�b�4 Adh+�0O�{	�sh0>�ۄȋ@\j�֏�2�jڊ/�9R���/�}�P��	qi"�F6�z0� �(\�t��Wd�w����["A�m0,Ηʘ��v���`c`v'j�V���<)T � ^�B	{5��j�[�M��5��w�f}������sN�|n�-�S�eg���U��O���5��j�:ձ �3U=����O��)_�ڦh�����"�V�
�N�bH��˿�[�uͷ�@K0N�-1Pl���G�J�;e���o�ZN�pѥ�L	��\��_h+A�>�7rw(���=���Z�-ֵ_!�G�r�.aK3�Sة�j��I��Ý��+�b,m��f�Sڷ��^�m��	2�;�?����RH����[�^����(b����Ʊ]-g�_���{^��b���1�����~��dy�k�b�y�+�]�����H�oX��K3��Y�x&ʥ�1մH?�(��֭���Eg����(ʇ���5����ŵ"N�*a�.��e�a�a�`�^M)�/�{���^�@U^�'��}9��$J�x�{��#�]��p�ԅ���a\<�s1�f�:!�MX~: ��Av�X�Z&�)����͕_'
n?%� �3�o
�b����q]�(p?|K1���ڤO߭k�� [ؙ
^@1=�Փ7�0w���c�@{��%�2[���qŎ/����zg�Հ=j�!�I<fw�?��x�'��i��W�&qdwGT�$���p�_x@�_X����Ef̡�b)�̡c�CO��Ћ^b5�+��v��q�!Hqi�x���S�}�'#��$�3n�� ${:�	hW�.B�<���w��]�eY��]X���濩ݻ�m2����@'�����u�W�7��;x~��ƃ0Q	��=����g�;H�Bs�'a� $#�-�qq�� �k]x��ܺ�"(�e�?=�[���{��$��O����S|�6��d]'���v����n//�|�`O���k���@4����;ďkݽW�9�i�������V��"����'=���� <�"uXr|�i��w��ћu�j@�;B�����X9���}}u�W"m�.=py.2f=���0U �\���'�<�Ԑm�{��h��B� ��8�ã^HM�B����e�)��O�����ڭ�>��Z�Ȗ���	�Ȗ�c�����m@6w���,��A0���g,��݁�\Z�U�n� ׄY�c�'M�CS��v���^;�,�z:�w�ˉW���3�JE��w�����Qu��JP�$�
�v䥣9��(ᔎ�mȍ<W�Z(�����? �T}i����T�� Y�$�1��=O"�d�?%��#���`�E�F�܂�kCo�!����ٚy�+kї+Y�O�,-C���S+O��6W;�O�r����d�X�p*�t�m�������7|;΢�<�߭s+��>F��[Uےzҫ1&�sE�"9���iM}� /�vN䔝E����r��>�bO|�wDx��93�d�i"���Aԯ���� R@l^v�去S��[	���.�j�ᴗ��#P%z�g�<�#��0�@b�3�t�m��n5�QȪ�-ϙsö���^e�,��c��/�e��>Y*/{��.h�ӭĞ��3V�Uſ^�O�q/3�e�Qni������wﵝ'8Q.�5K;���f�h��#8�����	R 	�S�����P� �1%�X�A��ed�S�c���e���V}cJ�2"
�23�!֓��,�-�R��������k�+��Q�8�Jar�vZw���,u}���#h��x�I=f�#���P}ֺp�4K@3
g�ܥ@p+��v�z��2����dX�8�'��\ �.��Lm䆀r�D��7ޥ|]�D�ę��?��$�
rmckm�֨�+��"��B=:�W*	1Ɠ���pN,��p�-�'�[�х��)��������b�{=�c����s���v�$�o��t�ر"�'[t�-�B�,H�$^� �����L�����A����=�0��ŋOI~X����=.�8�W_�1*�4�'�9rX\�q�Lr��)\��CC�P~���CB�v����~Nv�*RJ*�$��|؝�{�]"f���t��#:/D�_�����7{#�1��|Z�i�|B81���ɰf�t������t5�C�(�wGm��Sa�j73W��HZM�HT���0��f��y�Q�:��&0 ��������
�G�N���t$��D���Qm�ׄ���Z��`݁QnP��2~�P��Pz�0K5RE���/31/Lu�U�&�����q;�w�y��`�1�S�}�59�W�lh@�V�ѶP;Ƙ�F���j
}},t�ь�o+�	Wo(0d��h���TKe*MU5sV>��\$�{�H�o	�6��S�K��� 9e�Y�`�|���^�B5�U����Қ�H/�@�RH<A%���������Z|2D���/���LDð��'���;������l��̽=��$���l
��gm��R��D����X��P�6:�
��t�*n�:ȟz���=���S%�����]"���d}y+�7�m�}�\H q�u��]Es�N�Y���Oƹ�v�X\[8���E)����0����1:ec9�Z�X9%�����~
U�@�#�1�ޱm�)?b`������Oz9X?�,v�1�������^�l��q��gi�0<���}��i��,�L.��R�y�[��b�[�׃������|1J�d�>���EN*��_T��b�i����
-(Y99{6��,w��Pl1�4Ǌ��/�_��}G��ZQ�|0�NgB�ㅑ��K���E�Ì�� �Kʖ*X{���P�����/㭂���(��")��Ҫ�������x$�p�gGxX�-Z�@���}q����fl�1�xE_��T/�U��Z�|�ѯb��n��_���r	� E8�,�-P��2�Y���J"�crL��2'��1�8������5�ල�~ ʤX���g�4�i��a,��"�J����� �-�c�"b��E�:�'���s9��e�Q��mH��}�#Zt�<�v^pQ��K�3����+����z�Z�Tă�I��v�nQ�6T�M����+�}�����Lm۵@�H�Wü���'�jk�Y��BSS�]V������O
�
F�1M!�_�8b��m�#Y��O�����_�J��A���-PL��n%�6)��ɡ�|V�S�F��H�Ӳ	��|{���+��`�Q=n�%M�d�� IG
tA�@�m��͕nq-��Jw%dD+���������n˟�~�*)!}���n��ʉ�D�.0��Y[9a�R=,����RY�F�s.+�>8��"s2(����w����+�yrD�T{t<<�:�ϵ#�5h�`���I��P�j5=�F+R�������D�ş}O���@{$���?�,'��a�+(<����ڋ�����k�D�K)ǯ>4gZ3�IEe�o����&z �:"�+�V��̹'N�����K/�U�y�H��b�`X'#�B���!���=V�8K��kTl-�,e�5p�.R���K��6EGq�L�	2'��ؘ)B�~o�z���D�2龷PUr���[5��<�f^�N��������M.�ߟeg��5
?­��ο4Q��J�A����9����c�8���qiHZ�j��zU�)᎒�R�gX�S�SڣA�Kc�fb�\A?teh�߭&2[D�� �"`�[јA"�ٕj�w�h;
��cS��w��c�l���C,As�H�#by�lOx��2\�9��+B�����e�����d6ߺ�OQ~�= �+H�94ܲ���CtR�������\�6�;��gz���<ɋQ�8���̳/�6������¦Ů�v*���cg����()��c�H7G����\�A��s��3��ʚw.x��6���h���2��k�ܜrh�����qܺGЩq����*P)RS�W�[?W���@�չ��ot=�` �w�T���<��<l���C���;�1S�pG1� ��,*#��	Z_wN;���#D����O��.�E.��])����yĽvM�bd�����*����[9~^u�Y�E�X�I�ί�o���x&\g���yO8�ŢT��w[�\煜5/����Q�Ihs�:��g��%�5����I3�����!`��q�fN�W�C�����djV��H����*?�*}�ͷ���Z-�y��5�iC��������R���)v�������{�?��fES�p����	���?D#��$�I�K�d"��P�}[ߑc(� ��:��~��ww	��Q����!�������^��6(H������=�,��(Z����ns�c�n&o�A����?��yX��Q�_�N!e�Hԫ�z������(���