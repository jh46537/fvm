��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���9�{RԱ[ж�8�����������/a��:��#Շrb�,��Y�)n��M��Ӡ�5H�������w�� �Gx� �Vg~�r�5�t���5�Ш>@�t���57�s�f}U�������2'�k�l�E�g�ܒL�������(B`#�%��ǩ��b�y�ّ��o�ka�0��4�~u���͸c"�x���3_�XlB���J\f��E�W����	�]��8� HI{�s�zq ���s,=�G�:F�V����Y�e>�V4e�i��_�F`�mg�_}j��&���\���B�꼗5�%_����^��Q��q�o
|�zyFB	�9{i������ag�rʲ5Fe��Eó?T6��}��K����JN>Cgc��Ӛ�cH�`��(B�� �l��j�*���gjdų���\fٙG�%���$�����tXS)�N�����f�td���kt��*ؽ3��t�����-w��^XY���L��K@�Y<&��F���F7=��g���=�p41�z�Y~��%dh~��5���$/_,���\d���b�J�Jc�i)vs�L��]�U�Z4~,��7E,�~�<�bЄ��
c�B�(/��kЇ�6+���?'��X-%��,*Cd\�H�QJw��Y��)�>d*5Jy/�����֌��%�G(�^`��R0hL�U����v�A�k�3uNh��V�3SIK9�X2D+�����ٟ�`3ѝ�6&�
*��G�ӗBLc ��0n���m�:Ҵ|�Srv��?�Ь��P�[-�?��MW>!Oq�#���gXݤ���i�����K���h��^4�;C�p!��z�3���&1��И`iS�j=�%ݸ�T	�@���z' �O��ތ��R�֦���;Ӫ1���o�����Q�D����]�sgk����'����~�D��Q�؋����tm&��N�Yd�ROY�ϗ/���K�)��{xB��|��(�0�����Yfۓ\����Dg�� �%�{��tvǐ�y�v�#@`��U�1>&"��^�Y�UFU�/X��R��6E(�7��؟�o��r��{��~��L]鈗�[;��킢�y*��*m:{N5�3�_Q	��}����do�f�l�X;�=���?�;J��4/�VEo��$�Fj��)�����}B}�y��zbY=��۞e�!rGV�}�:Q��U��?�?������S�eS��[{G��)�n6Ƃ{؄X������K4Dا��;<��C��X7zs*i�.a�ߌ�i��?
Nu�`�i*h���C�-�Wi��KKMM�<{���~AD&�o�W⾋��1G��rE;��Bj�T�)wE��+�K竹��@�v;�S��x�~*GtN�ӕ���1\�w��!�/hj�Au";C�2��g������4�ʭd^�g���q7ҿSOjB�f���M��H�!\�qs����z��?ϥl��Ê�Qu#�+n��,��k�^F��\A�;�Fn�+|����#9Y��b����*� Dۀ����O឴`*T�զoJ`���8obH���ՠ��z)��Gj�0��s9�RD
� �xAa��B���U�V�!�+m�V�\.1bO��#���jN _Z�I�h���S﫥Bq�>u��F[�uvL!s@^�B���R��\y�)y���b��`!p����͖P�%摮���:t�W��t�na��#�I��bnŪ/['! 5�����I]��3�8b#�HFã�K2��zD�v��o�
�L%�e����O���ԩ�0r�*��I��Y-���dՆ��� �4�%�G���оh=�����WA��.��{����+�Oy��~)��Լ�B݈
�L�o���S��� �é'������v	~�%~�3=��ukMv�����Y�,�Mڂ�"�o"�l�Q���O�9�iRƾ@h��݊��K�X��+�_����e%R�}½�B����.�$�8d=�V!k:,����.A�Y�6^Tf^��J^+.�x}�i[��y�V@d0h�a:�\A�;��l�t]�&�)��pOd����;�>枖Di���k�#���z��k%EO������|n�#�愧ߧ����M�X�Z�J�:_`�WW����:�u��,��<��Q-l�Ne|�R�X["}�W���7�$РR��/4������>?A1,	~FZL\]�Y�Z��4��ρ+��3��n �+`{p5�͖Q�w���%Y��
���Ӧ�m�-��@7��"(�\���^u�L�}�s{� 6H���ø���%�S�I/c�׵����?��F���	��4��-���3��A���ֲN���s,�4 �^{�����O��և�ZC\(�°_���/ca�p�իJ<�x�4��6��-!:��>�mɠ���׸��~�h,�n��I/���s�b˴hv��@�%"�Td|�X�KQRj����̙���/����O�I��*���5a���y�z�z�3�9D$��2H��q�'��>S��0]c �pǴy��Nʶ�	M��%cU0��t��5t����'�}��?�:	��� 7K,_���ML�)l�����8�a�g���ny��
_6�q��7��(�_0#�+�����h��0��-@�8�\�����WO������>��#����sW���,�rp��.T2s����op_f�Ȏ��[N��)&��	��Drw0R�Oє�l�(����P6Mdɛ��p�� ����q��W�)Y���<-).F�MO��3�4�uZ����m�C��=�8�U	��a�_Tж8Ɔ�۰f��Vq�oFU��̿�U�V̷������Y[ ��M<�G�(V���p�Zg8����o��i檓��-��Nj//�l����EeZl"Ǒ �.H|��m�`�o8O�O��+�=��A�I�c�PTLY�n�\�GpPd��O��k��6Q�Es}�{�0]�g[^��+��4#���:��4��������n)� ��:[���i)of �,����D�-e7V���q� ���oVt�SgI�N��^�9�ģ�g6��hC4;%ZR*��h@��ܔ�v��0���*
�p��;�r��f��yZ$<�1b�<U�m�᲻�K�R2����<L���l
��6���2i�
~��(b��G�� 
�R�|� -����yj
l x��؃Am�8�ؿy��%}��9������v#��!�:�`-��U|6�e���Xr�G�Sb끞���?�VƤ�h����� �D��L�	1Jn�+?�׹dE��j~��U���k\�y:E���C�L�������� �߹X��H1x���)؞�
���.�x�I���1�h���R�;��B!_,rR�C��G���U2�%+�\�?�������k�ʢ��Xj
��|g�#
*���8���(e#���pHv�U��GC�K�?�sG��ʐc�8E2X��(O��yp�q���P�N�[0����\^]�s�O$�9;X�o��x�`s�'�I4j;(n,�T��"�l��@�"�]�/#עI%���z�
�� ��ב��v��&8���mT�8xBe�7pv�6�k��ol	P#c��T"b/��s^c�������nD��4xJ:��3�'�8�&����_E��ǩ}s9�\���@q��]q%TD�yĿl�kS����\����#o�	��_K��}��Z��a�Mn}�h�NF v��`=���#����U
mEn�b'��o��=�)M'w�.`�����Lճ吃�m�+����B��%���r�?�s���C��]6k{A�c�6~���Z�KC�ȭ�����©���qHD��,z�wLߍ?�A�"�6�	T��4q�6��{���'�	)h�n�T���V�1�Iؚ�n6	��N�g1\�\�#?�*�HQB��	+F�Ʋ
���z�|�R�BVm���>�xM�9��Y6���N�SEr��,t����]=��1VX@o�0�a5�l�F}���0_rO�k&Zؑ�>vM�ITy=�9@Bz���r;gvI��V��F}�(PT��]�	T�A�;,H�DY��ֶ�xϏ8v�3H�J~us�;uz	W��,[©0���X n��� �AYsY�"Θ����ך��l�ft���-�O�d��
rl-nC���X��@K�ߌ�u�j\J��/Y��)�A��.s�����\�)�=l���E��w����W�aҾ��P�4��$��4���3�h*���g��0 �V��k�l�s����;�|�}%�(x�S��Od�$Tn��@W�IU���%(��4A�A��X�+��N@B`?A����#�L'^L�ӈ��I������4�B�1��nVJ0�>�(�5A���i?��h��ql�2h���m��qf~l%.S%�Ƅ��$�ue�.���A�䁬�|C��V�;u$�g!h�`�B�.P�1-��ѝ�v���u�6�ZO��,vN��<5
8��)�1�'���8+���X����X��kY|)�U�i�r�+�
�*,E������um��G5�Q��cS�0�_�k�f0�8�K��I���	��Fޜ������zG]�|�Ne��V����'�-b>�ȸ��(;=�<�_·+���&t��"���W�ҵX��v��u��AC̓Bk�Ո�����'�S��^����w�hW4�zOүp�z��ioBN���<$H��T�T�
絺[�Q(�~s����s�v���?}���J�N�۬�.�N��%��\��9\3aL�����}mx{�b~8�!��2mG�en�`�p�.��m�6S7���j�3��:�ީ,��1jN�sW]P*Ņ8�07k����W��@.v��:�h�Ώ_�	{�i��G���ū� ;Ga���m�b��!�d�Q�
��/ݎ��}��UL<$���W���?s������8����?+9�
!�YQ8����;@(�ZII���7O����y5�&���.�ga*�̀Z�5D��_���&��"`����G1�y�=$C/�ҡT�.X�m$� ��^n,��l2�̧���ik%����y�(�G4���(L�)�����t��Q���=�#pP��]���7xRsf�
l�<��P'`�Aͼw%@TջbϹR�6t�o{�I6��U�l�j�]+��W��U�o	��e��K4��*��`�8�"�Ɉ�"EwXV��@��;8^M�QC�gX.2��C/?+c�=�?A�6W5�ꔅ��E�ζ�.پ0r��s��S���T��!RV��Ân� '�N��hR���<׊�x�!���T��{��v�FʌbBݮ�Z:x�,qsu�;���oȤ�+�W����m�Ϝ6%0��i	�R@4�{<q�d۪��=�h������X�ݖ��K�w���]����S���<��{�<]����R�4-��~����E[�Ƙ8�ٗ8��`5ny*AԱux�|<�Yx�ڪ�-�ڑU�V�&y�*� ��7܋���2���G�B�W���c#٬���k`��:FT0i����]�o(+?�H(��aϋ�#
�pҪa��Ë��pF�g*�r��c,����CG%��j�5��I�U�t��C��#��J�j��wg����A�J��R���|Q�>�*�L}��^�%�Eo܂[dʒ�^[�n������~P�	�5������rՆ��X�@i���k#Ii�@�I����l.�Br����&�]R5Ѻr6a�~��~>�hHwV�O/��m�	7�N`]�p#�<�N_l����Z~@?�
|9��kG��ܐ*c����\�]0�B�'�!m����u�I_��S�q�.pT>��pT����<o�u��J��>H\�>P��W��S�65Z�������Өэ���n]��z遉���i���"^��IX�`��tǜ4����=(����4<8��,b�i�:c��tH\*X��2��W��Ww���!���s�."3o;�d���tz��^�>j�Ѐi��V���~0b���9�����qM�i����s���F�]�w'�ܢ.��1���7�ò=���æwX�e��0��,l3��J��tz��אrmy�{K��i�{��U�_�>��K*�tT�<��28ٞ"p��;=Sd��F����������ωpddQ��n4��~n6��B��_��5=T@q����?X4$��,�xc�Ra(K��2� ����][{+4�&�Q�&HU�q�4���+��c���S>�X�����H6��x���&x��D5��:5�<(b�!�p�x)�
(�j�#�݅��^E�"�m��5���TOɩUW�D*�	�s�f�.ޙ����0j�aYL)��;��l�����6���Gl]+W~�&7��G0�vo�
y/��߿�2ܗ�����u4���ٷb`N9SGF���*�Q?S-�lO͢e�u�E;��L��i�n5�g�-:Q(�C��;RP�\���8��A�v����'�r=c'xa���~c��%z�;4���Uf:vo��!�@�#*c�Y�
��Z82;�[��+pwIDŵպ��c/���c�d���.i�"�M��>��0́�T�d��H�8�~Gn�%:=tӱ4��	7PU[�)��Eڐ���,��MP]��i���3Cu2U�vg|ιpQ���9t+4�~i�kp������O�l<Bݾ�qF��B��w�F���8����x���"���1rZ0�t����Ce��\FpI����7@��
Z
fV%��K��9x�Ey�c~u�Ǝ��ޟ�7-GI�r�x���+�%X�h��W�}�����ըF���-�N�ǉ,��}ް��$\����B��fn��G�- ����Q§x*�z����eτR�z�k���㷮�*����ص�xP���9���v%an�WQ�@Eb_>{�������N��n���V���x'F���ƙ��ռ:&�;�.��h@p%��{�FXxQ�ER�[b��Pz�T"�[`D֐�i�h�i<6ۙ_��N�S�J� Ϋ�X�����m����vry��]�m6��R=�>w?z�,fk���\O��qT�f���7�:&v���W3���qV��.t������<Z��bW	�L�c7`�a�8��:��}�|3�>�]�u�L���8*�5����,^Iˌ�[-z��K��Ą�OO�������z���[�3���+�jtK��� �C�1{�z0H��{��T��g��՞��kؤ4G�Ef�2��N��S4?��Ɠ�̐C�f�8e��hy���M��̼ ����#�3����L�z������jyMC8'|�̠�x��BE��1�w�����b�(h�Q�l���'�����Et�Ư�<'p����?:���DL�v���!</I3>+�O� {�?G=�>=ᕲc���CJŗ�	tj�� .o���-�������<\޸L�숕�0��,l��Z}�9�j��N��W���b�I�����E�6TυM_�˧	v�J
��ܙ���=Vڅ�6� �u�f4���eܷ2R���AK.����M�꣝织V�.��;��Tbր?�" ���0��P<��A�q9nv4w��bH���U�'�x�w�E�h2r�^�z����o�#��/
]�d}o��rmB���3v���C|��fX�9�n��e:��|����=�ăz�g�_#�)���O�ή���wۊš���g`!�	��u�y�vGT��x#� A����Lpv ���ǳ�;�]�)�â�Yy6�@,>pօ��b��BB�Pa���
���m��TG9� ��[b����C˱a�;5f0��B����2� M��d�k��z|C����{X��6E�G�ڲ�0h�CZ�*�"�C�P�Pߔ䢖 άHn�<]ko�$8��IbO]$r�9$�y�<���è�����7:���v���˱��Of��e��8�+e�ۆ�>���c�r��-�������@K�y#Ym�|�:5�_��hb�����X��#դSnΆ��	z�YeG�$���U�z�/�b��.�xjQ�����eo�t2KM��9!��e�ԓ:�~m���;��W����[����O�>�#��R�1b�ظ��m��t1�i}6�IZ�4\�B�rg��Ac�f���
�����3��̟�g;d}��}o���nd�Mw�=x���C�14l&�z@\�.�R"[- w�v�V�tZ�b!�L>�����3��񈍻e����ch����Z�H�'YG}�u�� 6�+�Aa%_��*�cĽ��]v�3|7�Y6���D��p���B\2�s�Q���~��j���M��g���"cm4=E�g4Dl9�|*���M�_��m���Y�ID�`R>�O�LhB����C�"d����T nU�l�M#~��RH�HBGX���b{��'����c�P7��]��D*�4/��4����Pe���!�����$�O/��(=o�e�d!��C����ڊ�δ����y���1� U��@��G� ��O�>�jg�
2 5�����L�[@_��8�����XF+�{�[i���������V&S� u��2D����PWb�E�Or���'x&pc�b������N��V@�����ea�)��'���/�u�A������`�*D�������.|U�к���~>�޾B]�܎����y��5 �nSr���:]A֔�8�1����iS ���l�����<W�?	ic��_��w�h��H�a�#~9�zG��	aEHvs���=,ˬ|��Wo)��>��������/���	����JBʶ�f�S�Y��zT�86m	siΓ�-�Uu|մY��}�����l�����2��ؕQـ�r����%������r�w2�R���iQ�,@�&�,r7��P�F�T��V��;��ګ{�^��GK#ʦ�s��V &}��=��������fs蕡������u�F:��z?R%!I�~@����M��9�T���s_��󜶛W�pt�Ō,������Lq�`n!l��&�����h( !�)�s�� �H'=�
rg�ߋ�E��al4�D`�6��ҶI$m�����qת��C�uom�����H��d��H��b����Õ�%����9+c��&Tj�����{�̱���>w��.����k��k!<��ŉ�66$��K�]s]�����Ĥ5yl=� �qb��J:��L'���y���n��JV@ �'�=�` ������������"p_��@���OS>��5\c���^z� S����I]�(�#��섖�o�{i+�y�A�c���ZV	&^�{������Gǽ�6�@��d�}���(X᫇c8��4�˸j���m�4H���'8͵�?�M\��E-uփ��7�o#3�	��������Z5��~��VJGP�2�S�Չ�P��b����D��atU7z��A4o!�ġXd��ڈ����^ {�rJ��=X��q���_-}�e�[en�4��N�P�춥�G��%�^_W����8M���/,A~�Z�Y�7nF��K���-����>!�\a_^q	출�x��@��G^V}���z+���\�=�DT5�(�,�+Q0�lqV�������0��D
�Ҭy����MN��ع=L�HӂY�y�+�a�L��I9�B��XdS� ���
(��M8�id,���~�FG�]a��s� �% �X�	�Ծo@8�����S��sN����C$��Re�5�O�L�,�y�>�f��dϷ�ܐ�T��R�ۅ�1��k�ؕ@( �>�I��G!F 7���EB�Aĸ�+5�~�-�P�v��:����iuB�n>��ߡ�	'k�|�er�f��?a��mPJs�WN4�ej+0�+�m-�?�.s��4L74֖��f���A����m�{��f0Y&�U��+��iE!|=���_Io�9g/��zl��q��Á���p�	>�K8�D[���vX`�m}Jt�)�a�) ���1������ ��u��q�v�h�Z6'�*0��C�e��[��d�4�J�T2�?���}Lĳ͍=�ܸ!�sa��Mj�d{���쥙2?7��s<Dj3���o�h�H��p4����*��}�:n�e,�����z���B��;w���e2:��e��E�S�9��uLBo��=3M��A8)2G{���0{�}8�IdT�4/� �-���h~���4��ysG\&��ۍzw��qf�<Ӂ�������8��K�ե�%���8Ⱥ�&�C����s5�����N�i6�����*�A�ӱXD �*7�T��>2��g?��SZ�HA���n�H���+9,t�PU����*��e4 �41�D��S~�H%U�<(�	K��x�9�%��8��kJ��Z�j�D
��i>%l��d���\�J[��u���spfUpb�"��NMh��Gw�5'�]��C��\� 7��;�P8��i�6߂�K=j�2v��d��A�����C���Nq 	���8̷ $�$D� ��z^�kZ��V���1Q��d!����N7�V�{}��q���`������b�N�����7���O��T�g�@�]z|P:��9�uF�d��1���}!OT.��I��y�`@�[tK��{	�gd�e#�N9�?�U�)����l�N7+Ѵ��cX)��^��2���̆f�ܤ�Bum���QoWa|ʪ�q�k9�~�{���ܡ�x�������H�g�[��)�*�>�8�)���h�9���c��"+~B��_�S�K���(0x�^ì�ೇi�,�&�p��Lx�R-NVE�D&�D���A�FK����D��sw��no�!�yGpf�x} ��0܂��/�1�a0��d��oV�
���.����QsOuc5��rMKqW��':h&\Q���D ����C���b捛�� ���aA���G�;zA�n�xn!DX���?��Z�w�p*����6V>5�/�Lc
�;�2��[����4�N���s��H�9��0kH-�{�����'Ŧ��\�?�ָ1�ɮJ"WH�7���P��3�+	W2�ݺCf���{�����ۦm�fSY�=�!.v�4�:�=ր�s�P��߁�u���/���n2!-cLw�����<۱��$鴰M��W���\�O��+�fvc���Od��Km&2�����+?�t�Zƅo�u�mJ"1	(t�Mk��5�S�_�����њ"���_?���gc��)��Ў��{O����Th�v���i�;�Z�}/���}�m#"�Ke�M�\>D��G3�jC�ՙ%�f�T����9@�� .� ��7JH������Z�g���c��M'�)]��`,�}y�s΃��+fq�X�Pۺ�6}y�H�\�E]���E��m�}㿾��?�`�J��ӄy��x�C����؂V����ٱF�� 6:�k� yI���Nj�c�p�~<���W�B��{3��ҝ��?�֊��)mk�`�W��\�4\=.�Uz�U8�<�	1ed&�km,3W���%B�8#���Aډ���S2�:���T��
t:����k��r2�򱢳lrV��?mU#�))�Yʢ�]qD��>���]��:sj�7de�g]��4ҽJ��~a��`���(�x���
��6�ܯZJ��](p���΅5b1��|;��'}��-�W!�ip�����((�a����E�xY�Ĥ&���o@E��=�|�%�����e��X��6|��4�!���p���������A|���R���\a��&ת\��M���p��^o�����q[;g%K�J|�[�s��i�iO�(����B�[|	����ux�{�7��q yj(����>�>F5�|O�R��Y-�Y�YW���7~[!�vt��aGn��&UlT��K�D���Ԣ�7"i<���q�M�>{��g�Y���ݜn��c2��%��Un�\�����A������N��NHa�G���h�J
��)sgoB5�	��i��y��Ƕ�/�� ��� 8�4"^��>�G�bCL�hW��ۗ���y*?B �)3IP�(�ϒ���ے��a�줯@48ن ���ъ��⭝M�T,hҏ�f�+Z��YHXU��oZ�%>�ɑ�F*�-���A0��F)�,�L���-�Z��^u�3﷟,�nl�ͼ֜OJE����/4Ggg1��PG��0à�p,AͶR�Bt�"��>�z�:;� �4�93	�=x�о쌁�>}�9ή�_6:���>YH�a��r0V�w�����Z��0s����w�������<�#j��B�1 ���*�dK⏇����Wu����Y��(4P6��/�H/��#��*���n��PF$�җ���9_8ݕ�!�&U�V ��|�t�B�\tN�_d�}/82��v� � ��m礥���{�X,��o�gtq�t Yntk.2K�jV�����G|#r�%�x��aSlRi�=�n'�5d�|Եhq��Ih�n��Z�{�4���l%��O�������������6�Z�.D�d�x���Q���Vc��.�|�õg���Q���]�wK�z��`튗|�>�p�t���2#��ٚsV��	25�g�����9+���I�ru�N�609'�
?���#���)܏���`ATA�z2�oo�6�HB����qi�^����u�G7_B6� �Af�$��k�4���*t�S�<��wT8��� �b�����<��ᕪ���k�v��a�Vxɫ]���IͰ��ɵK�93�E8W>Nq꾌=	���A�%�l	Z)AN��GV�����vf/?TlAN���8�F�ű��-�7?���ގ�B�W��,Ң]��u0l��'<q'����b�t�~P�^��Mn�8�і����皶�f�ꞿS���s�%���h����mf�n�\���2�/��6�q�T�#o����H�'�_"[����+[K�W1p������Gz#,5�s�77�Qc��pF���N�ߍ�$��<�ce\�g��A�D� �g��\Pgt����ާ�Q�}��~;��l'�Ȭ����3*���s5�k�[{��~{�ɲ����|s�-��:
ͅl��ar�#B�Hah�Ȭ`jT�����#i�Г:^WśwO��m�C�����T�r�E�X�`j��P�<����w:�UEɭw�Y�
��Ld˯�gm;�+8�R+<��<-9	�pa�)I��GV�ҀL|�4ueU�ی�-��C)�L��Ӯ����/'}��&i	�;��P=�t�sM6�$�e�+3����*�]-M�1�����@���;Ԥ�ΡE�m+O8^��%��V�e6V �����T��]ƻ��&�?��$w�$�/
2��Ň�����$T(�?�����!`!�ՓꏴJ&� K@�щ�I��H[-O�#�����8�D88�n�y���o���E
�!Dױ�U��ϓ0�В���T�給����\��Ű|�1��z�P��/�k^��5�����p��A�6t��m�c&�A`���gTj�UW����/E�S�7��d�$��Q-�-&T�$�e��o��[$��濄��ۑ�UR�_������p��F�hӎxD�9<#��E��"R)�a��^��\K�DRlVD��WǗᬉB�����F�J�s�S��q�7���>I;]�wu��C9�]���@ j]��m������9b�X�Ք�!�2��Ȕ�ߌH���$:��/���'��e@}��U�Z
��XJ��6�6����nB�O����ɪ~�����.���r�A��%�%z�;�z`��yPн�w�Y.y2��r7�)ʆ�ۻk#�����-��� 9!J� x~瞣b���4��A�����(ed�r-��Pog�L��*��ѫ��ä���z�$h�`�o�b�_`��4��HP%��a����9G.�X��{��g�(�2���R�03iNo^u���x�����r(	E��TKP<���I{i�x�Qg���1
�)�
�|���^�9�g����@O�6���m��jO����dt'Y�v�=��uݗ���x���k���#���"x%�e���./�2m_��ǸPgiϩ�&���	�C���+1���7���8$�0W0�5�ɴ�m�?L B��F�j���XR8{F(�#���&��p�bJN��9':@���S�IL�;�;
S;�]�-� ��_�a.I��5�Zܑ_�R���7�<����+0acH-JJ�9�T�����wP`��jl��_kN�AqE":�Ѓ�ҽ#}��r��n�`����Ov����ݚ���oݏ�{�i��co��Po�
E,�p���i�2b���th���.�R�=����(g~a!����~�jTց�Y�e�#�E�O����|�r��7~���_OuĠg���k髪
5q��t� z'�������$�����+z��^��F|-),����[8��3�{�*�Ђ���\���/'�Y�^ �_����+�V�~l�$� b���o��G'E�$�`gr��S-﷚�#ԟ�P#24���+���㌻Q��rH1���b٢������ֹXx��s�kJ�c�UZ�[&��%N��֓]J$�M4�Ɏ&�	A���;q�M7a�3��oa�I�����!�	\ ^���ƃ�ZԒ*6������;���ER���:deBEWr�N'��xgԡ�D������Q�h�k��Uv��iﯙuk���WK����VM�r���\wG���X=�q`6�1�J��U�:���:Q�A�����{#,lz��>�� z��o��ȃ#�����>��~.�}�'O�o�-cm!	��_J+���68�$���U��-84����$)|o'��}���d�T������="�+�CX��:���q@�J�S�C����3h��M9���I5�SdLV��Ha������+6��hk9E���z5��H�.	�*P ��d׉���j�6LƮ'���N�d���y�F6��ĺ2݋��}� ��(���F��k\@._:���-{�2��p�	��#Z�Z��.����;��{	_�������� 2����"ZV	�T��t'���đ8�����*�Ts^��0 ߘ%)��8���D05N �zv����� X���Wg��ۓ1>N��V;	�Fjޡ%I/�'lq�P�s�n%�#O����S��i��Q�WU��ʘdֈ���L"�p��}>���"0�g1'�AN�Ÿ*��4�"��Ă�X26�c�E�Q�O�`���k!����k�b��(h)k&;�LkaǍ�P��g%Eh�J������P�ڑ���آ�a��CC�L��vf
�^��3�]C��
AU��P%B(/����b�^0�e�W�=�����r([/�#��7#��:���(��q���
H�{�(��v�λwm��F��s��������m&f����zE��q�XcJ�p��'�9O�^�k)��=�v�p#i��7�m@A�_��d[?� ���5����7��/<�)�`�tl�A��r����}oR�)[2�7�뜚#��F�Pa��*��Y��V�*7��fۮI���0y�zfȽ��O � V�a<=S��D��	���~*]��7�)u�t���~u����h��K�j�؁P��.�p34K��|G)`�@��5�$�.+xg~���NY�-@�7�[}~�)An���j
@�S��1�����K1�¬�vM�O�(d���l�|e?w=Byi����cƒ/x	߾����i��:uC��P��&�yVsw���i�.�3�����5��C��;'sP+A����K#���S�� �䧄��̬ԫ=BF0�xr<�7s �ϧ<Z���ɵ�~�B�2k��K|���(�������Uk��A*�#m���Z�� |�@��IF�`�R�Qh�Pͻ�|����42����<~ʏ7�a���Re#|B�+��yW�]�5k��K	�T9�2]]�?,Ñ��	��v!�u�_�:�lUD�ֶǉ �U�:�mTV�!1/����
)� b(��)N$4]�F0�>�
 ��`~��Չ�8��}"A�c���T�yM��=E�#���A�r�+g��ؑ���.�s�R�Ne|�>O�K�(�˚*��v��兕X���Im��8��l)�/��+Ǝ2���\oҶ������ZRa��2�։/0
l^�T������wf�f�y�ᚴ��v/6�&�u� ���!Q�D2�5�~k̲��r��6����1VD���̓���T�K����IF)��ߖh1�$D���(0V�aP+o�Ƣj�O�"�$�!�;J"��+}@�<n�ߕ��X�zf��_n�W�kw�y|�OW�ht^B�w�����������ljXv���amqRb