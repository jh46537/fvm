��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���M���Z����;��b��=��98������<U�o��&5����O��ƭF��ы���m�t<�� �WSs�������()�M,6<������z�ȤSb$�dRw8^�0��?.׬|����I.����$�`�kU���(� �F`Q�	��A"���C�[5O���L�PX�5)!A�d���i�C�L&-0�벖�� �͓��غ�y�PQ "��8���S��<ĉm��g9I�ּ6��#@��� ��I>*�E��_�T��b+�S�7��6E���^1���񹂨�;?��t�A������6/+?}�ʱ4^��P��p�Gv:��8+P��ռ}H�WIiGI�=��l�u�z�d�?"�+]X��>�^�O�hU�^Z�w����.u��o���R}�g�$��lr��ϸ����Br\2�RT�����b�2F��,$ۆuڳޛ#�φn�1[@�����K1���c(!L?>dб�j ��'#�߳?>�H�N^^�y�i�Y��=ٷ�� ���K�MƖq�	�4NE�[]}G��h��	��z�K�_A)̧r���ݽ����l'_D�|�E��`�UC\ֺ�]F)���EI#��7[���xef��|3���{������w!N=����䥂�UP���X_ zBG~�j�e
!I�><��;`H�Y+��|4������H���݆��l�C�^���đ	(��#��B�+�.3zkR�/5�<��w�=�N�""�'��c�J��]�	!�Ǜ�A�����N�g�op���i�}���ۙ�lQ=�A���uK���ڔ��o��t�ٚyR ��S
����%���k��+����2���[#|Cm���0XRК-V�DMꎡX��+��r:�I�"����mQi�SA^�Um��� ��z�Jdt�c������LxrA�1��O�ЦQ�i�#��M%�!��o.��%ot�<46����z�Ƽ�PZj�Ǯ��0�-"�n�>!�C�j���+==��?'����Ls�vF��~5�4�܋��n��ua��[��rϘ�j�+�J��Q(�l��OP�u����̒Q�R�&	/��de4X!|g�	-�����L�F��z�BO�v��6��7�x�J�p+l	�}I���'f����Z��h�Y',�x�g���l���|I�{}�?��^*6��n�z�hT��W���)���f�9J9�BA�|W���&2��ǅ)����`\��{��}-Y��^x�A����W�r�b��m���y���Szx��9vq5`(pd�d"���� Y��E�X�q�1�"P���Q�*�J]�7��D�H���s�ƭRyoLF�W㭇��>)+�tS	5�L��<��9�p��ھ�<	�Z��m�|O
O�5F/_qy�}7�9sQ�ɸ
_���5J�#��)�E9=3�f��y�6��Ox��nj��A֊�H2%j��$��Tn�FG�<+ë�ÚV��A?�h�w@C���sv{$�e<�|�(�C�ȭ��MZ������n�������6�"�p�Uj�}v��߼Q��hnx�X��E�:5q�.��&�*�]�>�K����1Q[E�D��=��2|�:`�xV�D�
�����Ĳ(N��l�9?\c��!�H���5I�l��4Mx��p^���l��
��&�4Aއ����@���IA��D
��T׮[N۹����uw?h�j���50, Q����8�G��^����P��q��A{��8L��!�&����T�����w�ȸ�s���&�+�Mjm�&�9!���f��=�#k	���U���9nǵn/#E�0 �odf?��G���(�0�Nιnۗ	]�s�Zn���lP,�]׈_���pt^y��R܊�F���^�a4��VG,O��Ĕ@M4��l�nj�y �&Y�72L�`�n��&�7�/���Z�;�:z5���wM&�T}=���F��ޝ8
��\!��D/�c]�Y.�J��<��O��7�[���O�1꿃e��{���D��k�N��:w��6��DvCҍ�3�h��{u�Z�A��\�������h^h�ȕp�9��I�����pE;V�@&#�n�s��S��������T������/��g��\��ǜ�3�ۆ�:�k>�h�Z+�*�/�2�9a���$���>7�l1��Z@l�s$tk��:{J+�iR�Zyøbn���©#j��+�H=�bL�϶�����s�@� Ay�x��-�&-��&����Q�}o ��q ��I�z�6��!~��VKX/�H.	��
�IoAlQ���y�2��d�"b��
htX��\#������䍆�� %���ﴰ��w�9�.��/�z�Z:�nӅ��o>�v����nl�f���3]��X�UO�E>�]�o��H<|t;������/��Oe��N>�~���r��w dl�)D2�8\w�Џ���\�[�^ϮW.����e<��I�1�<&�w��gi�dIj���2��B����8`��>x���=X20�'�sp��O���#s.,�`��u��.:�Eb�z�z�]ql��yJ"F����{%g���%�a��0�/p~��a�9��-,������a���<JJ�/	kQjݯ�e��p�u1�L�,s35��r�V��x�%^�:Q��]{/��󈵌�a舦[ǝoo>��s
>�h_��8�a�b��;�I��ԟ�&�=Aq�:���D�=:�2�U\b˟o��-�'��]�ʁ��i��N{���.��q��	�w�k�,$�[�?5��{|�F���u��M�A�oOq�
7��,�f��t_VH.�aP��Ӂ�-n%l