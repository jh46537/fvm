��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��b*]���I��̞m��w^o;�2q�Ŭ���O%�.7{�n�|���Ob�Tx����q�1�	J�p-֝�ԬHP���"��%s�"bD�K���_��tݟ 9Y{�(������gf���x+;S�	6���/�؝��/C��hb����CC��:�<�s����ZƓ[�>��^U�m�(�1_h~<ژ�G��;�����J�����K�#1f.)V
�� �� �OKr��1� �cO� '����%��agy+��!nS����8Q�ˎ�\Ic^���^��i�\(d��7��������M�~���R�at�q���|��^p矵�W��b5�>�)[�B�����{L�N��!W�y` $�P����m��'�ѓz&��vyJ���8��]tP��W��*�<c�d�S�������2��RUW��`�����X<�D	���W�`�
��ensl	�����#�E�[MϦa��ߪ�~�����`�S[��g��^��l���PϨ���Wu���|۲̋tB?ဏ G��ﻀ%Ϋ;8��Ҹ���ށ�	/�����L�9q
v�����Fk��5��J�z�A`��-fp�:� �$( T��&"٢��w8h. ���s���*t 1AuD�DF�#q��_h������%����y�� �ņ�H?ķF��%�WM� ��a\Q�����K�
ۏO�c�Ƥ�Dl�x��%>����[����h�zXZB�l9ȫX�B ����2i63%�;��w:<��u�5w�YC5��ʷ��t��|O'݁�~�ƍ0XP��B�sKT��	��T�����θV�g���Pn�q�@�6I�uX�B䎼4*�]��n ���ǓXX�	O�G� �n�r��'e�I�*�ǚp`*{N[rnF��j�I�Z|-:UQ���2��� �#	��}5�!X0H�����=�V[?�(o`�����XZ�����D�o�2�;;��}�'�!���ŮэaX�dm¨������2_��O�{|�����%��zW����>^pL������4�	1�4�sW��g�N��b����dd<
g�u�=��r�dd������&��EM$����)*��w*ѻ��|�?�XJ!�J���iꎴ�l�OЭ����?��z��*���lg�{�l
/\�>U1<��~��%'$F)18t�'��~j|r�
�������g,1kL�q�3� SLY�~!��ӡ��W-�F��d���x�
�����{��m7+�)שaD5K����ko��:^�T�.�sm*����y� 06$�ɚ���3n�'�u��M��"ݼR2���5�`;@�y5�aZ�8˓RY��X�RZ��������-[�� �P�q�Y��Ͼ���J��Zq),g��t�{�dh�;f����ew���'NC�7A�f�0+�*��v��'$޳��zLy��h'j�[��TӀ�'���:h`V�-��qU�\[�I�.i�1�?ș�<w�y�]�1����W%H��CL0��TpZW�5�����Z���34+�o'U �zT���#����(���/�vl���[\FgFl���W׆<�%��X���.|�?��Q�����O�"�sL���1�����g�FõN�m���������X��m䶕�+�C��-�������	Ñ�>�e�"�r�[
�{��n{O�M��;2�x�#�b �a��:���7��w���?~Ɩ�R��	�-�ـ�H[QO�V��`ş 5T�Ж�x
��(��=iv�e,�7�G���1���Ɔ���E��
��k4EX�d�m���m�g0g��D�TR&qh�pm�!>��ηY�0[�p���m��8�'�N��)���DxY�C2ķL��ީ��q'��e _�8gD��QL��	zz���b�1)����W�k	�nF����Н��}�\D�-^:h�W�4�&�c��*aau�������K�qkP&��jR���[�4Hޑ�g�����hO^'��Ă�/o� k��su��M� 
L
u,ZK>�`�gwYu
����x3����a�1�f���c�%c��v|עU�Pi���Fh�vMs��}�ij����4��@� \9U~ζ�*�RuS���u�a���?�mߓ�D���I�*��P��4��y7Ry+�=NDڟ��$b�Y�(�h�2R��9��t���z
T#�����A�����N��
 �QAO�G�u'��F<w������R��g'{�$�`�vP�Qb���d%�����鱍171� ˸�^��tn�)^�i8�ūR��9�xSnw	R'w��su�Z��"�[��~���o>���3+�C,�㷫���`͵�� ��kc��F�`Q鳆�vc��e�9���/�gv��)ޠ`j'����]��̀~���h;*��{��M ����L�BL���BĘ@���H���a�e;�"���.VQi*�+ޞ]��o�$';æL��r#�(�Ƶ���^�Gp��� ��δ�̌Z�#A��KF�c��we�.�s�I�+��@&kp4�RQ�a��$C����@�Ӱ��1�"�����j��-h�S=:�'b��3�v���ȍ���N(m2�? ��F�E��8��0@���1�Z��~�gg}���y'��ȅ�����������Ď���x�P)��ͱ���I���1�5�<v�פv�N�[3�m��Z���s���#�J�;A�1��b@���zg��u ,LJ�(s����A: 9u�+���)���`��.�������I�?k���,��C�=����[lݺ����%'T'8�ؿw��*������szu��I���X�R'�}9��v����]�?�h������F����MW�e�Ll�	�	��ӈJ�
�i�&JV���搉� �N�|o̙o!dz���h;�3�":AL����^�kL^����+=�󫰏E�1jV*�r˧+��S����Fi10�t��)�|3�ؐheb��[<T�xQG,�BL`3�]�q��7&�
)RSͱ�43*`�C�p����vשlg/;Sj?"�%3��Xzq�����췷8N�{D�D��W.���bP��4���
���U�VUM������
5HidTP"�˙������׮#���_%�m�3�~�h5ŷ�Җ<��ҿ�s�ڎ�El���!���a��oC�f�
�Ӝ��*m�O�������0����e�k&��1	�uq��;�^@�hA��G&�8ؽ}r�8b��ɊRSФ����n��%�Uǫ�,��˦�،&�y�����(�6w+�\6)*�";�����'HL9�LDpt�����޶X\gR[ۉd��������u�l�6��j�V�i ���� 5(��A��+z�D!��y��5�xDeXw�hQ���?�r#oa�������]l����]XcC �s��.��lv  �x���2FS�M���v�?�$uRB�e��lp���$�<~�H��j��Nw�#1���X���z��ӱa�:_�`g\O}[w��9��;�$�����sWPO��u�����_�C��	x�1u�)�����Q�WS�9�:A#f�/�) �d�ǘ�++��Ӈ�G���U���A�B��8l�W9�tr@�L�U��(��`�X��~�%1"W��u9�z,3�T8�*~��{mZ�(�#t�9+��rxm-���z���t�)׻���Pg<���a�1�����ev-IN�������[E߭�h��0�3�U�jJ�����HZ -w���Ppͼk����'5���r��y�prż���� ,�}�h��Tp���n���N4B�a 3���
<\�%���B���-�f�_/,̬�
Z���bQ�^�noe�e4���!,���c�۶/q @į�ǔ���q����0u-+H�B�,�9�HZ�Q�X	P� 㩞��ӻtNL��O��(��	h�@�7w��"�@�r�1�ƿa/m��h�����杸��U��A�}Q�/�.�&�۔�
�c���8/���D�11+T<��U���،(͍�Qo�o�4��� `�"� c��Bot��F�5�	L��ɉE	�D�@F/"y�f��=�o����-i���L��h��Jt`��5��W�or�µyC��B�
�d(d0by�b�S��w�UҘ�s/Y���@ҳ�7-��'8�a_�1y�R��]W���b�3V��1�(T���wnm_Q\��Q�G9��D�Q�8��-͒��h,���?,����������׸�T,�ww8�:D���{��}�P0��KvM����WQ�9jV��?c�,ΒofN�_�4:��7�%��М��z%�#����V�$w��FN��`ڼ2���z���=Ч��F2��2T�`�]?�
Ȯ9VF����c����
7��@�1iw�M*�h��e=m�Vq�خC�d��I�s�ZPe����	RA��"[D���M��4/p2�8��	g�T��7���y�����&��A��D��lZڊ�GԻ�e��W���/5wo�!G~3M��E}Pjk+�ܸ���we:�$�l�]�_,��'�1�u���J��(� �"��k�y�4��)��%m��'���<��l�dr�|���+qPg����z��G"�ҍrѣ�}B���!?�J||i7jh9�n������Z�i�Qj&KW������0*a�`�u�׿�-���7<q��|ɹ׊�횧��h�_��)�8��z�|s��8p���=#�� M١/Kf�Ϩ����}��A7�Հ��i	ܠ^�A�F�_x4�qꠣYn�� עV�9-��e�"Ec�]+��T�r�M|2�B���r���37��K�C��8�������n
�&2���h�Z��e?�&.��� An�!�s��~܁e8U�;h��xs������R6JI����
�y�(�{�}!Ӫߪ���ut�SV�Eu�0��%�����jSU���T6��S�����25��)��� ����S-�F���4e�{�C�Ub<,�$�A�� ,�P0rj��w�PyN2��k�����v�O���j��J{�*n]>��x��>�B�QT&�t�W	�
i�m�Op 
ʃ���b��O�<S�3�ȩHb䧧#���c�\�Z����X�hi�HڟR�B��F1�^C�Ip��h%��d�����)x�chpܨ.!�R����ch�x1:��