// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K+nB9pWcP1+S+p7rIssLU0ykOZaArR8A1uaPjZl0s+T8/uwvS6GMzi36A1XxlcoT
xPbyXp9jy+sU6YAanoKdKqLDRKw6nUBv8EmNyiBy6DoYy/IGjW1fPZ4tfKNuM1jo
1MJoPAL/9lhFnDnhg1fB7w2gbKKQh1SxxWFgu01bkPA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6048)
rLWIfwZYf95ulhi7tZpU+gfv3aJbKe1Zj63OCQOhgKgJJPI/fU8GwnOxxaHJ9PkO
/GQVF6NBCus/kFFrkVkgUPXR7B92R1RPbIz9ISnv0/OLhPNkYL57CpOWzRHaPE5p
X2IC0UG4Bkdmtq8OXE2IH6K+krKtrbTO331rwC1Bj0TAe84a3NyCRtJY3o/OIR2R
XQ46NBfpojDznJEnCeDmCYS6CR3DfMJ+WLzqJbNS9MuiDXE8aW/9mmczsBoc8486
1QkXvBF2hoB/NzIj8YjcdadOfXCP/aawDJr086RtGvfXlGl63HYfnCi9vg84mpxk
du74akORJ8ULd9F9RSwxeykUyLQS/8bpjU5RbQEB7FXkOt+kQNQ3YSvUPWiHYkuS
JI41/14Tki4Rv/VaK6bhRUxMhueA4ss2DkCah4Dn0xGPC99pLaQ/+xvxGhkuu6OM
Frq0hNu8e+ArpMl38rItWXWgdybx3MmtieJp1ZKmBX36slXJwLybRhwWGZEuo0be
7trA49kBjxkUDS6p4iw8fT2esV58ybFaOFV26gqDBU7K3iMxinzdXTEtbzyn6HvN
8skEMhQRw8rhJr6dw2LNG03xlKXtVlKhg2j1gDfB3XCD/W4+dBvGLrmNFR4kQp+S
jzhk65A3Xaw3/BNQdogD2J18NDU/jiRrwzqAaynkuNWwSWbdzoyr6BR2XkOBdpQb
/sOk8fqsfnhrIdGtOxGgR5AcgIMR7iJ9HBzgsC1iiyBbOvyqZXLFb8+iqBfCPTVE
Mezc0ptASsP2vRMKrhecyHdUqTVUGYbv6loTiYn2ksU1mgr9C24fb5DPKJk6iwib
rSZvFQfA2bX7eRRi/vEcymyi2lCbzxS7GX5H3Fk3Z+Qwx/Ss+8b/T0QuvbHbR8aL
qXgmEQ4Hdn4vR1RyKzPnDZtRqQY292Tsw3i0dcS2ff/o5gsmoer5f2gGmMRnVJrY
42+vayCthGiP1EpQakHFbEWee5S12Md9d0Mj6lLJjYYOle58P9u1OsoGzJNYZ2zP
F0hdVIRqH1Xxgjr1M+1PdE716LGTcGYRt7FHHeKSA3UktmjLtGXtAD0GnkNmui2e
WADg0jOU5P1y7nNniUSz74XPRw61Gd8X3U8g7qj3ICY2Nz95MB7bwJIvNgHU4YQH
zS85KGYj1oDav0JFhmkGJS2T5AWbk3MOGhoefmy0iMHpQlxVCCMCGgWpc5PmBnlA
FkDyOiOtF2qD9SRVxfSe0mvK4tx/RBbUofF867uR+8Ii0yM0EHXq5zWznE2pvg4M
/833CkvPJVh3IKEW0hyIM5bffU8T2Mb5bEMizM8jWrDZt9lksM2pofeaan61IWot
4M9GaX//AY+epFeYcYxB4nsq6E4DFzXVY3//lsRfRELmS2KLCC3JDa1EyfE1hxdg
uNrch/5edCekyXxJ19kr93ZongnA3SH3/cDe8hzNkrZtb1aRTT3NAlw+B/2aZ27A
kcW98WP6+92K4skSM1f4ZiZo89tmLuAZ6hOPK/DSh32TrHhBHHDSfrY8Y8f73gms
PAVOsKdZKstYkF5lFB7N2aYQjszBDaOip0ZjbBycpHJh8OHh/+hS1d7eBzDLBdgS
3jOf8LA+GIpwufQEBRaf6tXpisy+8tjIIgsscji/k8hmBiF26TRFoRnjUGQyHzb2
OeAX0Ms4is22KtaTY79dwmIdBHmO/dodVIUCAEm+8f6zm1u61McmDT2zZCBDz81T
ut8eQb9N+C5cHg8osaROPg7cTzgo8CaqW29v1REe+prRtzyxqWE2plBPH4OlFn4m
TNtYS8flGAbAO0r9kxTcbsvo3DhWLtq1eyWXuEXUOujRbnGQwVzBM6zS7iMcTM6w
QECufbL49n4XraWTnHTsnxOCnvfvJ8V8q+l5fYNt8j4wdXKE0oOYeI0KIJmzPm71
s7KYrB6e7CkmLKbMhFAPLKCQ3Yn1fBGiU3+eckw9jAy8bxP9VN4qnm50uxJuQEAA
I2YM8Px3u9ZxawDcJUmamIB6Um9ZEm8IPDmExofmGTXKBwwhNFykj2E++QOEU4ss
4qGQzpHx6YXMR+FxoUR9wHAirQD0U3r/9r1RcYWzI4cT+ms5zWugzsSW7ZzyVM6N
rg1gU3mnA7+byfgz8GO+TLUP5o4kOVEcT73kr6VjTGjWfuu8kKg66CN7VvvtkE9o
/P7Wnpl0kDcrpMLQepg8O1zATip3XZO8HAqRvhwWzeTrN/M3jpmV/FvwzTf88jzs
VBhHl1G83UnZcS457jZoiS99g1+v9O+hNBdVzFluQ+mbu3LhZrgmrEIvscY0lL9d
doLExVOMiDhb1NEXFlNXtYClnwTEC78QgzQljsVBdRoekhjKW1j2EzYE4Q2xJ9rU
1VvELl3XypAjAYiYdZlQ+xUiYKnNBukyRQ7iE0IrFP7V//2D6N44euhkK9z0a2pA
TyM0f1pwsrU04TVlsraQ/arbmU1/veXcJ6la315FWe5cgG+wDFWTnl6y72066tEp
DmJMmUk+uF1X+e7TIFBMHLHje5I3G5ReBmkpZ02yegCDVeL/OXnwjGMn5S1SC/SV
3fB9kxDP5r1d6HGCgSCeWitlq2/vzAZDNbLMP/FMn3qDJYBXE/Pg7jgo79LMLpdA
eQfWDMYBy81z/J/yvGoAApLm2ejWrL3S5wih9HYYs2NpMuBBaZlAceEeQE4RJkvH
javJjy7eu/3G6Tx/n1KRQ39PrB9R0MmsXOE03cTiloMFVOO+sGWJVYJTrJWGWQ8N
PHkUzZDqFrDRTIBtHkdLnz0SPoL8xgvVOIzUJ4ZGKP3B3cWECKIuMRkf7uxfJj0U
CNFQQdXXrdOma0ip3bIHvI9vym96mPkcup+LLre1E8dwer3c1cGMI0jnY55TTKKe
Mh09y3fT8Mc6p8Wmhw2q/SsjZHP0xrWDQIRH5EGOBQoW8FJLd2W4TN4ndEAYDPz3
8Z9zhAyrWE12swa2LyCDUT5x8NSVpXUJbX2ydGUve2HKldzA5xhZr9ZuSLelP1Bj
rUAjK6SvKQA5DSxDjSiCS0IdNJuDCY07YDER2wSsHHFbFvbvefCYMnzfpHneVEV2
FszRNgqOoSzCvUhtwnEgdmkK3zf7m0yabo+FM3b/ZioOKQWwk+MVdQHSC0xIGPXE
AS4Ea5/mvmSzHHEHmioTKYbgDLUt2C/7ynaECmVYHckkrRU8HgFNsk0xc0adegNJ
3wdgkNjbKeOi0MdF8cR+oj3BhRTW/j6XuUDXEFpC2QGkashSAkxZyERH794atmq6
99SFpi6yoQ085zDfOrnrQu+oZcfjutjYmQ0xx4xHlCVSv14yGHNlA+svhOEeaBBf
FW8033pAou8MGwK5+sH7pm3GVKHK628smP+V2goaHfnSeaspT25j1gAYhEAtn15i
53xEAQGYENkNxCvi0XqMFpDCWH/KK+xCnPGxIsPPnxlXDHJdoTO9KQOQhuy1hytj
gLzQvnJxiMfhiI/dMmAdgyflBNdCXRj/6k460nN2hrBtcT49e33qGIFxd2BCLaZY
tfdpiv0W/POEku/oX4WVXfSmm94wtqHd+aau0n4Gr4hpGgyy1T75xs8fDNZKt3o9
jrllsaLAaomZLcj+UG43mm7qiaOuhIxuyjU7cB6ywcM77/kcHe4J9wqEK8K09gmk
u6nuAvsWHLcTOR83aVz6kXyZ6OCIwlV3HrNpjUG0UON53B2/M0/1a4GpXQa8C6jV
YinJgMcG1BpmTQFjHL06OLuTj2gnE7jcdRg8cfiT8dkoTJnt9iFSk0hhwqQFrJXe
mbYuE5HcHkZXai0lZ2jkPgx7gQ4tsrG+uh19w7E71qzFlH4bEszn7BQW9A541Vio
GgKiD72B52w8Uot8HqXXZ2Susv9FF2QO5MWW6UNgRDF5ugOHs4Y9NcnzIiQpAFpk
ruGiIXUng0O1HH2DpL5JKjpxkot7atSq9TwiHlXiT3QZ1jmIdJlgHEouo8lAIQVp
YCMXilGZYreHp6BLvx1WltJgG/9mpV2XT0jArTZI2KerEhFWC5dX0wKttFxN6Rie
9/63OIWZfwEgBfDFcYsYQSEZ6THfUdJpkg3KPd0p/4RpesD1xNUrMESRmYFLAHnb
kDIbnEZBWuFemIYRRVVO3KefW9gWNTXj/LaalTxnhbwb0UuSDG6pU63TRJBoMqlp
21G+CEZoU1JxituQaNyeDJx5A2R3MPmHXnjSlWbPLvszPs7fEbqCOmzASRo4hbNk
+TMIi/mzp6Tan5rKB2rbv2Gb+PcYKMUVlYoaknRkxV8PRcQ4Znkqa78/xuzaVjvo
Kt3QrNwDl7ZQgfAUSuIOziKZltpPERlIEP/zNaZh2yK1HK/fqKrGtwjGeUIbWmzW
M6lm0c5bIEKDoMo16LeP7EtXQa5C0i4cwgtTGU31+sQKmtJaJ122k8aqI4B2Hqws
XHVp/siKY7zYRvbAt9wXYwofFoVQ0jnCN3R4Nm2glebau6Ks5VOI0vJYPzX4cPM5
pwHyyUdStjrel1FHB8EZHgzcwPFDkQKzZzKPR6QgTvrs+tPp/VuL0Xa6A52oVn1I
4PqrxWM2tz9OP1BdCOBVOxAMvtF1g9eWdQepBFrI98+70ckqSf59gK/TMm6QfbRf
I4pfyJtXnqG1yVQ9e845/Y8rd+61k5oTzhMDHMNiOT1rBFx7dv22VGHgSYIZmiiR
Q24Rx0Xa/u/dsN9fIAUBfiKePpvatuZYgO2g+ZtDU4jYNaHhYGJZV85547ITiwgb
l0zMM2VTw70kpJRFA9h9/H+mbqK42efdBhw9vyKXh6CkWIM5iZz07LqQQxGNEanx
m1JrAJG69w8nZ1aF1L/0DelRBVJmPJJ1dZbNb/7m+H00SrlphIBsv2VRbaCzjb5I
tpPNtB56EBJG8yhhF1UJiqa4qDGZsDsYdg/B3PKF4v2FwOb436IbGSj96pMDem0V
uaGBnUwLWmuYY92qntG+Jf3BbhDd2CK+KEPikyNUQqBOEUwkAPLGr8LfJtBeeBzC
mFUVRQEBLtA6AVVa7doq1MrPAQeC5a4U150E3EdOrrJQK4To01yfLZ4Xrfr4cTAN
IxXjknZwNeFnTtAziNlGZ/lOuTwx827wBpib4gfyJ02jsee+wAhfLJ6kbvAi8ZXB
tfrdmwBbhldPu3ZYRg8yoPf5w5J4QZVKPTwcIBz/VPhyPIRSAhym9C7F0OtPrPZp
uqzV2yh1cW/8w9p0ftk/wV5LAISM3lJP3SuIPkjds8E1XpB3jef7nS4CUqDfkGnN
3APVKVnbf0XeOL/SCTfgakzQvNUnWa5vqdNKMnBhMMIITzDvmNbo00tdMh8fjJCa
jNi74On6EDwVOCgwkkDWoYVowLjPwI3AJiZ5RN3SQ1FzBpzAMIp4QVoRRDPVL5+x
sIly6tFTI/pEOdNjiw0OvB6GMEFMIHdZTtdWTgYvHu0PDaIiq1Qbvy+UBMivTWy0
XEBbzR9O+uRHBd5q01SfbdaNDOuMY1tClm72spa4nEFIWJd3HgYSg1OSnMp5r4gH
wufuWsqtxX+hGtrGr/BLaGukvUz2lg3fwrs3dauqdlJW8Zpv+nNrhxNh0JS3URRk
0ozMOnlqwai7Qp7LiXU2MBx4lKaU4PYxy06GU8OksN4RGVbGmio4BzWk5XIYsFZq
He3iS3jBIUaGO8LOIfaUT9mN5SdaUrJPHwC6NzR7+BiMRYBQngqC/VsJShxBfs75
x5m6BeioDOgQPdIeBH9i7QSrFsX5K/JMQCAEEOgq6TvGXSTeqxAWoBzKzLCL+Un+
VLUUiBo1omMV3Ywv+EeMDLjd9t1v0JhmWQbXhZxOrPnz2gG6LJL5hFPuZP0QMiI6
GX4gTX+LLvy+JIKfDr3HAHbNBVvHjA0WZqHtBUAPg6q0LlygGxCoKErWbtEWCTgb
hWbMtt0jFTKlYLW1OWNlLoB0XK1vx4aVEswd7V2uCnCCqUY+3A6IYPoTuHgIHFCQ
o2XmmZ+wgEVYJfDJ2X7jIfYZh7ruoO4Tq6I4he1UF/AhnpWwoAXEBS9G7BpQKky7
a050RGaj86+AwDZKCa1BbIxwnYZUvCC72vw7eQn3+f4zQVgAgHg2Llwqt8H2XJyO
sX/H3nAP97b4b8RmUIySr5DLgTC3A0DARotGkGVjIFB65cjwYb5QBtdt5SETNDPb
OdQ8c1D1GuPdOQl6UDpvMwJ3r6tYv/02ZU2bUdXZpDrODCLiK5ZR9Zaz7Qq9LEdj
PpeZ1MEelmP06DQGdcyMO3uJu+XPLxyYE7i9RRJdljpie4Wo1QHvvRoSbGvQlqsC
kCVUi28hZQpGSgdqBCWzKZ6su9NTa9cEERkuYO4V0WpCAJ99SjgzyfHaG1k/lajD
H7i+M86ogMMw03oA7eWtHxm/vxJCsZs2y4GlP6Vd96KyOY6zcYFovZHnYf9q7v5n
rV1A+xIYSQP1WLTaP9BgLUOtX3SUrUKUR3sMu0UTfhSbXZkv8P8kd8KtxrTC/+Uq
Ln+C/sD14CTitrSXJkf0kOxY3qy5iaX6SNTOL8QWXbHdlorARq9Y1q0gAey6Kwyi
YGavsIJ0zwgqtFvb1nQqQBsdc18YOpOi3NM3KltQLC8YCSJF7hl00klX4ssu2rCE
POP8z//Cw7jfHa64KMpsgbQE7tejkLegG9hmf0AHp+R6QRqHUYKfYO+ai4lVhvHJ
LHeT0l11DhEebeXoHRymvs9SzE7zzk455Mu6hpMHZ9wZ19ZHjfbBq5s9Xug3BPXS
/Zl0SLgyoMt8n453OGXAJvNHFHd3QZ0GNWquVGu7lYciyi/mChQZDnVoziKMcJoW
0sEGqR+zmSORA8B5++dap4naRbjIC6AqLYKdtHh0H4nBC0xlF/tWonkczvcyqqVC
zlLJ4iwNUMCXGaX3Nq2FfKKIs8iG03aWiBh337XS5RdzQhaGCnIMnxYbP/tXEzO1
UgkIw0XILXEaCTjhl48uKuZXvx+AuhfqFsR45kEOGtoi0j/WmSe7UWeHtaGKdg+x
KYFWf4Fo9tJrCk65Q9LAF+BqRxHQ+DohOS+Qpz9SVU+EHda1OLirIfBbUe/fl3nx
VBPyNZe3F9uIfJVr3Hmy5OMeDBWeYDD9vITHlHdBETHsrv7e998sYYkuJM8/0J2a
wRbiV/1ZB9qbaYlZtspLQRjbR/V6VoAWpA0G7g8fs5tdz5EyboSu8G3n2jtMxjfG
NyWM3a19tJ1MovShgry3sUIxpqhsFRQJn53NsBkWehCWmy3kK/Huw7QI53+c9lKx
U8daHh7C/ykqEFL7zR62mOB5ueXX+tYKsvFq6fIS5AcgzIlkC4If8t++k/9dmPsn
B/7i1SGKzgTkH2qJXM4NvvNtaQuVbtOWnVsGFoHUyNy7Z2cg86kpr+XgG6WvqFtz
vKaPgeRBzjugPlap0+urgMxibpUcuOC2DRksE/Ly623M9wEabf/l3WK7AB8SXFkO
xgkDPUAVpBaN69DeL6ybMneh21H5zq4SwfYLFG/E3zh9aqE3P3ZN1TUaXyGK7+Os
fZMWDby5o+Jz//xcBnD5ds4kQsFYbhH5MVT31PAdlTqp/PeNlnqJnjNXjCSBr7/P
ownZui9kwLC20ck6prE6jtN0OuiVlXOwXr7Z9CpsDhySgYGjoyHtAaxlJlhoRDEY
mo24leenYkUiS3PRFLCjux3+n+7ZWXn6vDg1aXwq12rM2AVOxNXX616uKcP9+5kH
IzhJrQfajlg9vFAq8jWnWy3PfCuu0tN1EFF5zOjZZ6oag1m8XcPFRXOTS2dmj8/3
1eAecpvrJsmV1zjMP1+AntCbbG2AjIiMBq7MP4Y6/UYiF0SM5iWRtyq7fi4dPZ+e
lYikY52n3tIb2CwBcZGSLy99P1J1clqLlSJu98u3eCwbPSaUY5wh4RTfiLRunZGp
VsIm/PVVZXdnBGyqWqoRjo48H4aGz7iU264Bze26smqfw6mCaFKUSbaQloiCWu0l
IDLBFTmImP0i20+1tgapoHwyT0Qph4UqTNe5bv8Wc0ZCu6TF4AlfbbqYrNck+uYc
Nseu/7JY7oWapGdUNxEZgT+/ZLGPVF9606E8cf1+O6pFwz2qFlAWa4FglMoMmEVC
`pragma protect end_protected
