��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)����\VH7�d��:q��Z��
�'��Rl3(N�~`$�u�V����I��t���Y'��W"���<s ϓ�T�F?���-�ܚX==@c8�j	qPH�	��\�`���Y�ÿд�9a*�Z�Y+up��Nɕ�f�����4�e�͊Qm���A�|�v�H�v�Յ���J��P��M�븓Dp6���8Y��<�X�S��֬�9J+k�� )91���y$�3�ټ�#o�-+������s6!*�`������q�)�`��F�ldL~�j�xs�mI��c��I$�+uhv���~�6#�,�KXX�����0 &�'5����S���0���5)8礣6&#p>�Qu���� 	Τ����pe�Y����EG[_{��]�B�xU$PY�o�黟cy��Xۘ�3Y������p�UE��(F��K��h��P_�g�*�F�N=	�BR`}��cM��)���y@'�	q�A���!�/��k�.v�G����mڑ�Ȗ���R�3f�~]D�-��%��ϲ{�$.o�`T��q
-Z�rƤ� ��Q"������@L/u�$��TTj��s	����Zז�idR{�c����;�IS+�x�q��̳s��u蕝�N���7=>���L��Ʈ��E?���y��<=Q��8=)*�d-�I�����oEN>)N�R�k\��Ԁ��z��pY �t��G%�l�����K�}Y�m���#e����πaZP��=Q9c�S �d��{2Х��3+V���4�3��h��0��t,%I5�V�wf#��\4||O�|
9C����!!�4l�G?�q�_��7��gr}��Ѐ;(c ���.��h�.J�S��NU���Y�XO�Fc�1����Gk\�z��I�*";DH�ݥ��r&+H��EJ$=;��(D�Q���&�P�1�ѷ��tv*��� �L;P�0�7z3��qkz��,�^�����!
���b��r�j�M���n�b3�s�c}c��D���X����I��B�h�&E� ����R#�Y+�^�rw�����tRu�0�+O�AsvcS����Z��ǵQ��0_NDme)bxW'��]�Mh��>�	R��l�o��N����Y�ٱ
c<6�P�����~��O00�AI)��\d���B4���}>)W��B�h
�^;�3�<�=x����O��H�� 8���\��tEc��v;)���,�莥|B5�\wB6'�����.ȍWF>7:R�6�V���J3E��\��P�~�/��插3�<t�y�i�f����@��� c����WV����!%x�?ݮ���+�#6)�mP�]%������C���i�s�%���D�G�І��C����lMsw�cȼ�	Y��w>��h�S���OR�2J%�}�L��ff2x�Y u��� ��Ł�i���Up�(�;�ù/�}}��Π�[�c�# ̈́�}I_%�Ѳ����nA�G�eu�D���b57X}���{�W�ǯ���5�rDC���c�˞����r�O�+���crc�� ����D4�B��~��C7(��V��������!EAjŹ53s�#_�nE	��*V���D��Y��{�ޭ1�?�y"�XȽC�����F'����"��)'��w~>�)�e�'���Wr�X��v+b��h�����4z���e�܇p�]���%�9t*8��Հ�#=:��er�0�4T�3������O�[��LA��}�b[�Qk�~7�	�My�~?����Wm����}��C�.~���*ȴ��`H�݂�b��T�u�i�)������f��R3r^�3�4�ڊ�#�P�W}����teE#��Y���!�Kc��c�BpDN-	V�U�"�������/�ɷ8D���&W�KLD ��_0}6Nܷ����"�K=�nh;�tک�Ŕ�eFXA���Q(�.x�L)ȅ>ç%^����̈���P0a�S>6R�Ü�r�$f/�DFNd b�h~0������HE?G��w��v�@��lI0�u�+E����A��?�,B�>nK�~�l�q��i"�*�0Ę��ǈb[�|f�F�x�3�r��C'
�n���&��<���s��	Z���ٗ]W�z���y"�HU��z��3�R���Q�'^�s2'�j�D�����h=lD�&R�Gq��kV�����C l�$R���Z��V��4rV�u5=���������K1o��bR-ˠF�eKs���ؼ�8o�k�D�PFU�Rp�Y�H
�t�	�����U�)��ma��q{�B��"�
τ��Q���۸m�����@��F�8:��8�H�!9�N)�`�C�G:�@޹���r��x�����鎒9L�kh-:#��3��Af�e1(��R�|�I.Kq<��i��Et�)�:%#v�?���3��i��u��}+�x<ʪ`yT����f/[�T��F���׊gQ�汌:�X��6�R�c'�*��D���e^����[Y��T|��ѱ�S�Ɵ̙�T�89-�*̼�	}˒U�M��FY��m��3P��vթ6�Y�f��ھB=/���Pi���2rZ�+���-�x�"����Sg8|c���ih����bуj��ۯ�O@X`ZՏ6�4��8�;GAJtN�J�|Sq�
���n�O�E�����2&��.T�W�'�+�?�?Z��F�
,��Ҷ�{�5`�*���%�_��4��
�;-�"�Ԩ�t�z�?ѣ��J&P�R�O�E��H)�ݘ���0z{�R�n�������)�6e�_P�o�i�rxb�C�����Hb;.�1�ɢ\��(�F6D`�6#=��=;�:�(�g�)<;���Um�%g�{̱�xfJ��be!4nF~�.�i�r�#v�P�+L�(7)��3B��u�(��u�4,l:�\�rr�Y�:����8��9W���{��������Ь�����)Si���X�B�����Ͳ�;����΢|lm���š��땅O�k�d�7u��Z��2�4��;|�P5�Q�\����?��y ��v��7���Iz8�7.E��Z�Ut�Q�Ӵ��W���X�AN2c$4�"�b�����~|cޅ?&@��'�Y����������ys�wI�}�'"ך=�{��2ܟ/N?{0�����4ၔd|h��0�O �v�N~�s���Ni��ӓ�o�U��Wx@���#�=Q6%���$�ω��-L��M��9����L G���j�sx��-��+!�[��p��8Q˯�ct�������z�R �F��΋~P�:�*����?>�,��*�zʒ<���|��#]��Q��u_�EQ9��r���.�i��w��
Z���m�ih�w?7�k����<U�w]�jJ�7t�kFG���M�L�X'D�
t��Q C�ޣ]�٤��G����Cm)~A(4r�'D¸:=�m4w<+�Q@e8�ƶ
id3����N��M���J�ʯV���7j�)����Vnu�6)�@��֭�YkC\v�+ �@N8���M�C���&(�8��fp�ly{�P�7<�~�l����_��(l�s��Kt��U�ol�1I�-�m�����Jq��Jͷ�{�~u֨6�磯�4�V���a�Jڡ�-JV3ҙ��k�ru�3�C�#F�68
�����7'�ֆ����8���'/�	�Y�Ũ5��TJ6^����<�m��u�b���Qi5^`ӣӂ^�lcZ��<c(�V�~���g����l����=@����^z��y�m~��T2�2�ɭ?9Ɵ	G���i���Z�Ԟ���e{' ����D,��n��[���N�[4��@0�*~��^��ӵ�ę��ΤJl6����&>���5�q�Q���U�`��f����#I�(3Fm��ç�hK�%>�\�R
[�h��u���|�M���m���/�r�`)��/��2��VRF��	�	����\����j� ��;6��h9�q��s/�
R���/=����+�wVs9`���� 8��_~�����Z��݉F&3⁀�