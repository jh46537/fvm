��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���a�%�sK��h���/a�y���v��=��w�����:�y$f�*,�RA\��S����ћW;�U���T�Ǔ�q�0`�eѓ^����8YU?to�Pb�I�����9���������:����l	�~�Y���)���L8�|m[P��Z�ј�79Ӄ���e<���_�����^�2�����
v��;�{a�<Vx3�-�����ٍ��/�[�mg������o2����@�m�e�?ኂ��l:g(Ozl8S
�-�CW�gF�5�դ����>��'K�:���ϵA��8�l��X�0S����b&�7�%)����!�h/Sq�㾴.��"��w[�Xe2�.ƿm�?�g0ۉ.�*9D��>[ˬ�?]#��m�g+��;��Lb�W%��"�����n�F�`��VW��th��Y*�1 ��a�|�!D�+�iN��P���u'��?���ɍ���5��KQE��.υ���ݩr�#�x;��D)4�#j�������- � �\<T�㹓xHc�%c90_fR("��mysg�,cŮ�6��*�w;����sJ�I�Uak��,E��G4�ʦ}�KN�&�ۙ�h}��>�e,���&R��AW*�&]�*�q�d:���?���,����z<�oi�G� �>CҔby��yH���a���f�����*>�4Κ�[��S7���tML�W�z�G�3� 㺀[���݊��6�RP����y���%�V�16)PM�iX\\��.~�L��]�JL��"������6��t(OL�Œ����K{�J
�2.*zU����Or�CR�I�1 ����3t�C�UH6�y]���j�����n��{Vs�e�B��J̃�l�)XO����CŮN'Z7gc�'S76׮�����b˴f�8�ֻ����WN�Q:�V���� ���.R�;��Ym�&�}��p&7<�m�-��jsuR�sh�נ���)ZeZc��^�QK5�7h�4��0��^��W��[�[��5�rt=/����-�MQ��M��0���ڟ�s l�aMJ�(�_Y=lG�i�R^F�k�>��C_�`��m�#�0�e?5�l'|�4����N�t��r�x���&�'��K�v��|5a_�S���7�;T����}�j`���zsM0�6z��[��Ĵ������q/:�h4�j���s-2���߹����ylܿ�bu���ctX��6#˚�V! �W$��`A��K���9d�̕���7m�����s��>��'ix�Nt�����N���������g�Q���*$e<!�m�0���VY��n~�:��	�x�����'+�8�\�گ����q�6��v9�l~�|��aR���.;����rҎ�G�蟎�p�s^��U��JBx0�����=&�s-�i]�7oF	���9L�f( ��8�:x��5�kȡ�)�༿�Ǿ�<y�����ǱmQX` �J�x�U}`�&.�EPcJ�I%�T��R�p̝��;�[��ɔ�>zF<"��"��"R��/5�[%���p#�L�'n�Ϊ
$U���y�s@����<MQ����>o�jY?����7�{�� rt���+��`|Sc�A�p.�J��o��x4�v�Y�}�4�l?�͸�v��@��g"�
m>rY�Q�ұ���:��u�b�|*nخA���S5N��'����C6��h�*Kl��=��A"eSH8O��N�����V��w1x���k�R�}�C��y����^I�\�'�\�S������IÝ��i�g�K����~�6�|��65p�*���{t�P���ge�]A-[�2�Cۨ�"!Â+�$7f�Sf�).��Bd��[��w&$�Ƞ��bp0��M��/|޳6�Sȹ��J�e'�a
�*�A�":���1�F�y_�^�G
�V/��5\��^��(!���R<R��Ֆg]�X�cSz�+��}Ћ?q]��&{\����&.fMl5�Գ�oS���O�ڦ�g>%� �'�"�������G<$��@Iᡈ�#e��1��C�ڊ\�7>d4���h��4����i��=b~yO�B�dl��Ƃ��em��L��K���奊��>���a.��3_����}�]\�2��i�z��#䛭%���:�]��*nI`|�`Hy���=�ps}Z?���g)�B$*���u5M-�$��}&^�u�Ko��pH{�Q4��̳�l��$m���cE04�1{��.�������m�U�Y[��:^Kr����g_r!1<��׾Z5�~�ރ�b�:�YB*k%�lewN�}���n���~�U����L�K*``�����<M�y��y���[��Vf'R
j�� �b�������4��x��4��*9D�W�{H@��/�z�31ކ�F]�0�1�Ė�H�5�^~=�7�[���\��K���AJG������װ�sȣ����7@��{9D�c��L�=hw�J�y�)8Q�̓�Q��6���v��Ə��UK�P�F�q�as�O��q	n��e��"i	����z�K�\����7fg���!��8�Q%-�{(�iR�g�=^qTJ��!�9̗���S�������*w��c��>UCNRr�*�EA�H�t�~A��_T�_;�JN��tE��$+��;Qv�kU;j�% k-=�O�������_ TF�&����"!��a���fq���ؾF	X�؇2f�8*�0g���(<}��H,o,Ѵ[�SVT�`O�^�L ��.�d�۹���M���E�8I�V��H��y���$@E~�GK��4�>P,��SE"8[ެ�H��}QQBh3BP����j�T
�:0�?h�b��`=�:�g��R'�R��=[�[�����c�ú� ��*Sz�(�Lgx�w��#�h�����%s�(���]��se���F ��'�(�K�v�d����� mSt�M_k�(��a�
�v�ņb���Hn�G�Y��\xO�:���+T�_��S�$�5[��(b@�q�!��VVŬK,�U���q��bN��q�/N��H\��_�3R)�a"�O�z���S ��4���p����$��K�#,��1��U8y�[�H*ROP������ĺ� )�`M>|X�[TN&ړ
;V�Cxd�c��R��D={?`0��Ʒ���ax}Ƕ[�sC�j�oZ���^p��I�ְ�v���r�íi�z��_A����Ǥ,N� ��x�?�:�u����64�VO���0Dm�>D�u$�C@��'g��f�כ��YLϮ��b~.	��)n̚���"`�k�5a�h����M�P���6Y����}���B�]��Vz�D�yIH2����P!j��wd��-�<#��_� -J�� �
��{���$�#X�*R�qn�O�(U�`��>Ck��+�:k�r��"�hC��JZP̴�g���9�r���g�q=Ȧ��U����`.���I9_5��Thk}^rp:\Lr:g����z��7\eE��}YLN��	�=F
�p�JʹQγAǑ?m��42uɽwvF!d��Χ��*
j�Q-�ٛ}�����G�m �v�f�8�N�$�w�S@G�#�B�ߐ�%/�a�E-�b�^�#&��Q�5�@u�.cG���bʥ���t�%Խ=�3`��Q���N���l����'���h�dF���.��d�����3���	F�
jj��_�%`	y\u/�Pae�x(��z��p�c��h#�3�&��R�$I�X;�K�FE�]*IY�w^�����Fuv�;�Q�yb tIȉ\Eň@�V��B�67C �����`ܧ�+����!Vs�_mo�ĕ�w}�Ou���?τZ�k�3w�<����,����A�����aa��e�����[V��[/F��*7
.�Eq��'�a�簕�1��%�Jf8�c���n2kQ(k�Eս8ZX�w!�� -\w���K�H.)s2�
@9�d�+	#8�i� �yT�����_JU�ݸ�'|����I(K������?�����S����e�m��H���ԟ;�Hͦ��X��8I(f%7�:��x�/J����eO�iwx1w�-�h[=����ek��aWC^]�����6A<풳u�����|�3����`������
��_�I�iN���̀�:/@�;њ�Ϻڦo�L0�.�D�_�mc9+g���]]��K˘�
�g@���t�y�H��	�#/4����#<Tw���"�u�,	��R��-Z!��Ðgl	 �"U����~�;2ǁ��f�)K�[w��{0�٧�}��Ke�Ɂ���{���1V9�Gdi�b����B^~p�������b�������$P��������i0�a����adw��7Z���{$�!��\�Q˸��3�h�'�2����"��N��*m�����%>��[z�6�#$���Y��7�:�6�����N��[!�/$�����0A�����&p��)����~sV�B�`>#t,�����	6Toa����tqR"��X��~ǆZ��_*���"��m�7o\kx9,8� i�!��k�%@�t�V�����C��(DvG�4;PM��~�u%�y@�W5g9�n(mS�h0���Q#�l�G8����}W����vp�'�@��R��yh?2�`��8.�t#�Xyc���`j?��h[��b":�2�)L�E-����`�\?A�ܼ����(N��q���e�����sP�:���[�
�[˄Ff���-(���hiP|J2����	F�����9v!�h�q��@,n����'�!�ϕ~��I��=ņM�7����sd��-�� ?�\Xl�o;
�wE󎭏�L�3x���EFAT����sVb�b��Z��E˹�]L���S
¤��_��M>y�<66�,+�B�gQ�!0_�UF;c!Z;M���A�f��	/�%)UNQ��e�}������A��sV?�o�L�ܬ���H�ȍ��B�̈́fX��jc^�mO=�{y�ǵR�<��n�IlvB'w/�oD�-��M�0��"fd��G���5��,�Z�������:a�!p��i�s��jT(y�����S���Pݒ���5�ƍr��'�Z�\�oG�⤌l��Ȃ�j�f�U=�5��jv�m�qĢԱCr�s�����ed��۹Mw�kĘJ��[I3����xf�����(�@���]7�C�a��1�~���<�rU��>Z�z�@�k��2F<�9	^�{�f|b��y�L��u�>U2�F��l��q�E�A@�M%尵Ҵ�x�k
��
f �`�r�Z�=JUJD��!N+v��{=ɿ?L܇�w���F���DqU�n�/O㲈�iZJD�a.�p��w���$�s�~m禄:0�E�Z�ƾ3�C��q�bD���f����=vH 1�Ϟ ���CV�OC�MRj����
O�����OЖX�b_���4��6�E����	G�<���p��Wr#� ����ķ���F�׋���e���=K�їx3��uW����o�f�^Xm��Sk�%��I&ؖ�T���G>�\�Ň.�.<;�&qg�(�?��eD��)�Y	e~j���o����kEq��J����D*n�IV��s�U��5a�S��x�`sPb���3����V�V8�Y�/iF�� ���_�*�L��ء%�ԩC[��x�Py)H����e%�k)wxX[���R�x�qa!^BT܃%.�8��
��gQuw��5?�6vuL �*s^�E?��u����ϔ�{��SZG�}L��H���j�2)�����O����}L`�����=��f��g��@�sǠ=�N���w�dC����C�A|�I���c`��e�4�A�^������@�v���u�spG��`�p0���oy�<�Yܖ�I�����޵s�bh'H��#�Z�
�mrW	\����n���ˠP�����n��8�����<Ƙ�x��+\����z:���ǂ���8�"��hj�G��%b��*ŗ8�� !�y@]���
��B�s��r9?���d�<�G��jny�|`�R5p�"Uc�xβ����'x S�VWd3�{NZq6	Uo[��������E,���jem.�xk�Q�_�q�M��9���;�������y��1�ڄ��ǪX�#M+��_j]y|t��f�·74���<mI�����S�6��u/�),^�L��v*B�Ć�S�"������������T���j���i�u����JF����4τ�h����{�;в��8������z=D����u� 	+�5�V#��b�p �����a�J��g-���]�K��jhȔ�KKU��s:���n�|y\�v��������ۿ���b��z�>*����#p�,�i�N��=��&E�*I����hl�Ƒ��%B���5�Dh�������4�^�Px�����2�D5�W^8U�O��U��
�ό����r��2�j�LZ�S�;d����<C��f��D}0�D���M��B�M��� ���[2���W��h�[�W�;�y7�����4���_i�G��(�'�)`�Ь�>�g�o��0�X$N>�G������?�
=d��Ω�̾&���6T���/�[k���i��������<ǐ�ܯ2�q3�uu��6f�鵌�F�w�Nem�Nq0����8�q�ѩ�;|�����{�}Q���Ki|�Ę����N�J^3/^�@�T�Fό�����Ѡ¦(s��ᖺ�������ltqb�Ьӊ:v�K:���a� �<������mo�8���qd�w%���Gf����:i�W��S;!6���=�ٜ.�ݒxd��d�|TCo%���	�qŷ0N����Q�	��O�у�Z�U��6}��ςjތ�iе��og�c��9�EMW�����$��k�	� �O#������X� ���t�lN^� 1�p���y5{���Q�п��ϟguj!��/ �&f�Hz���5������P%��ko��۲�a�	o�Hv���=��FpQ�6��}O�#-u�n�9.��~��ҺJ��������v�Kc:�;��Z=�F<�!�p�FY#���z?R͆;��@�I#}��<���X����c���P\��m��աK��j!b?�Y
ы%c��u"\^��\0�}�JO.�z���+���&�Nخ�%��C	n&��L���j븆��Z�`�`�dJn��1�.�K���_�k,�����{����OT��c��ϱ�+ }��g,1d��Y�i9���X�e`�yO��5{� �J��B�Kk�%�3םJ�V*���T�E��v�(�6=B�~�gΦ:MG���G���F'O�e�(1�%.aHeE�k�O\�붚w�Ɩ�ٵ�	e�RإtX�IVW�9�Ʌ�2c����ūfĚ�<���` '(\�ug���Q�3i�3F*�'�;��5�8��� TuF�@��'����Μ^��؃�Bko�7�*����%I���ĺ>��n�cpWF+%�@���VhS��,5�4��()�:���MQ��c��W��T�xx2�\�3Q^���5b�#R�4��a�l�K��7��|)�-܁Ϥ5�G.k?2�Dv���=ﳟ�z}xn����l-�[�=8�ݿ�D���H@��;o�*��+��E5�h��Y�d��n� ���0q�eҚ�,�{AY�L�D�*�I�I��T�鹆	�<�;���ۄ��1�M55�A�C�������BT��&,�kR@S~�X��s���%��SĄ� �.Tȗñ�1����^�8F�D��q<L����Z������2a�9�ֻ[��v�4���1�c<FFw���%�o(�ؓT�uu628�P'Hޥ<���aE�˔�9�
��~d���[O$)31r�%噮�ᇮiƢ���1nao��c$x�	���v֘Z8S3�4�W&cdJ.��E_�X-�тe;a��6��6���|o������jǷ�/�����*��FRF@x�m�
B���s{�2�[�H�l��w�FS�P_��S�V!e�a�`��R ��a�`��Cũ��L��L��y�r�gm�6�uy'k��7lLOV��9= �l��<kއ���ȫ�{\[�k1-o�4��0��ammj��v�Tjjr4�W	��B�&;��V�7�4�h��F�AJ��]�Ej�Q�s� jI���[q�Aݳ�g[t��G����2>����ND�P=�4>B�u�����XpQ�o�|҉4��ӄ�ad�5�O��/em��d�!��w���Z0\C�v�Qw��m�eqo�ٍ��@zW�O�����O���l��~��a�oݩ��r�-&�l,C�$���B
c�'�g�8�QD�A)���#�~R1-�}�ڟ�>�Y�1�Q���#��9��ۇ ���xXq�kIx��8�9��'��wS�\s$��9U���1�okJĶ�8�ɲk���)�Im��VP���%w���]�~(�P�_����F���	�}��}�(��	���S�ѵ�D�z�����X˾n�p��S��N�������ZN,��jW�t��vx+�a������c.4��M�QGp��V�7.v��0G,US�����$c'2r~�U�ޯvԂ�4b7�ia�S��nM�
�-5�;�2=f���ku�6���'�b��1��4�����'{FEvfT�Y�?^˩ֈ�g0;��Nx7!���)�?݊��:�,�c��7��wbC+%%��E|N3����u {[r��ޥ��@(�,��lj�G[�ΐ#(CNVLs��D��.�����L�4C����\�{�"�C��,aK ����N��%M&t>lJ��-�~�F�r�WS]����H'�A�w��I�g�k�þ)��%?9�ŹՆ��e+9刖^M~���m����^?�Ka΃�	���t�j!a�<y�h4r��}�Bߒ=�c�;*����� "p`Ǚ�J��@��i��� OH1֞F��x�E1_���؃�LI����(��3����Xy��{��\E��rX4�>p�|~ӑ���çӜ�4��7ҿ�O%��Op����Cc���q'����Cb��E�&���8N6.���w�#GM��R&ص�<��b]�lSE�N ��7�^# �x�+���n���Or8`sO���*�����R$�9;�1TXΐ�G�[�C������>�C�֟E'U�DF6k�\�5\ӗ���t�8�{>G�Pg�I��иL��y Gt�K�[@��xQ	T`�CУe�f��)K#C�F{��	������.��]*��H���r/oM�by�J�DO��A}Y��~�w�{��/'k>e�;P��7l�g�E��2oj���X��b��oC�~�WO�����%����0�e� �c!7��y�sxX�GQ.#1�N�v��lw�1�D����h@3�Jӎ' c�\�������}Pt*q�X�h��yD�iV��UW�Gk�-�s���` �Q�E�l�7��vxE��gdB�VH&e������Y]_�j�f9AI�/��RI0�ȴ�l�+ϊB�I�3"��?/�:�-b~-��i�)g?`J����=�s�u �)TĴ*�e��LR%>Lm���E۬�H%<�&�TX��_�^�Q�S3�w fI��I&��a�aQ�/�+8�{�����L(�ə�K��dN�b�A�w�<8+u��d@<fOT�ē��z�@{��d�x	{lQʎ\M���o������X��f�q'�ÖA�2���]�6�$��O��Z]���[z��J�?���;�R�姶�J�䧳�[B�!�����X87OH��n�O)?u�]���z̛	o��0�m����<��Z���,���[�CO��K3��X�<��v � �M�����_zk����u(�oC�;~ǧv���so��, �O�Ī�&��V�N/�%f���J�j~�4Imΰ��>�'�Z���F���n�p�X0QM��o.g+��A��X�Y,}��RYٕ��8��p|1�$���<�!6���,cJ{�s*�E�g�՘a�Э{�6������h��;��H,��K鑖�]F��!Wny➧����펍�V�Y!P����{n�U�3V5�����c= �V�����w�GVl�$�[Ml�|A��w��8�1{�,�H�_Ϲ��z�h&bS�,�.Ԛ������ZnglC���g-������*P`�K��қ�]+4&d����x��_5����c�sx��v�Ru
b��W��Y���m�Vx�������S�!?�x�N�&��i}������/ʲc�;�}��<g��u�8
�~�7�Z���K���-��e�F\sK�M�v��^�l\���d�%��~�g��?���$*V���ƚ?���.VuR_�r�L�R�H�(�;9|(�F	��Ҏ���i�9N�wR���^um�&���J.S�!;P���Q�1ἝU�L6�,��ˈ�k�����P�Q����?�*���
 2kX��[��o
��ް\��>���#�0|P��bu���_{�L����Iz�z]��7�(^5� ā=%���5����O+쉁ON*/���uB��a+����ʳ��ӌ0q�N#�d��>KB-`�l)����w��yh[�BK���vo��3��U��4�����a	i��08�P^&M��ǖ�4��y��Jz�=�)Re��6����Dw��Ģ��S�}"0�H���Y���y"�,-'UlJg����/\t;���$k�R\#�T�*;=����9.�X\���6�9��asJ�v9�``am���{!��U�aYp�f[�B-ܳ>�AOx� �RԲ>5���K%;aફ�S\7<o�ޔ��w�BU%�0ŏ���-����=IG �<�e|���B~Z-.���(�83g�<i<	>M��%,�%�}K�*&5��g�d�����#�V��"QD�l�	-I��2iI��L�88�5X�A5��}�Ӈw�lb'�3��|,bL5������Uy1;U�;�Y�G
�э�jMv����M|�JR�.mڏ4+�Y�\�bsm�a�ܰ�ˑ��O���Q�"�`m�n}�@���)�0o�Y}^�jz�oC:8Ѕ*�o7�g�d-�����������������kKc���$@G�m8��=�.�uO�fc�-C�	���,����(����q��u�?�'����	]��7̖�IF���\�,,�a_�`ߟ���D����>�Ii!�M��:����Uɖ��h�Pz��G!�imXZc��!fLa!�����!Vƛ-��}��+��ym��t�rL�]V��6�G^��y��2�UƊ��NeI�M����h_�T��4ا.�9���ȼ'S\bO) ��;��&t,`�Y`{�=���󨴅��'�p���ޠP�G�j�J1'㍙ڑۗɧ�O5y�;�h�M,q��g��!1�?N�����%���J���S�!�	��k�5F��/�sB�~�w�z���O����$x4��x<�)sj�Ǉz/�tN����Z�_@4�	�o���n�9�R���'`/��F)h��5��*ˋ�c+�n��5�b`uTZ��'De�����8E���0��9.f>��x=�S�w'�ҫ��<)ҿ8��5��/���s�v���
��$�$�E�Oq맑�d�H�(d���/c��{����)����5�(�8�θM���!MC��S�j�����"w9�;0ǰd��C�d2W���<�ᴚ�������.b�顇?m�ͶO*�S�^��Y(8�?��Y9Sb ���%i�"���]�xѠq��D�|k��Y�7*76K��({���_4����:@u#�;�Z����rpqэx��1�PuFc?Jh��	%����H��Wf���
B���Z����B��Ǆ~fSc���rh��h��N%$f.v"H~8�����B���N;�����c��uX��d���7��h��!��]b�6i���e�͂�����3������a�Ot�P�s8��#z��6�8F��X�!�r���6�#ɨ���6P�M������X>�,�P�@��+C�ߧ:/O ���#dب��ԽfS�3k5%������]������v����87J�����QUR���{ ��� p1�޳��sz)*%q.�"����f�	����r����FH$9[;�-M�zc�y7�������b"ܧ:��*u+��G���sb���~R�������+(�o�sy���=4
�Z��k޽a��-U�֎w���dB�z�8 �9{�^5��EYx���'�@�@�}7 ��OU�n�b��ؘ�.�&��c��`���_=�ݻ3�a�!��-V�ϭ�z�Z��ُeCvG�����]�i5����MQ�E<�����RT�����$Q�N�D9S�S6J���������`p�ᡠJy��ai�|1ϳM����Ha�,����%��xZ��K�q������X�����P�겁y%�,�U����;�~�?ɇ~��U���)ӕ%�?����0�f���0�$��g�5�wKH�%�>"�z�4���^�Wێ�rY2���ؕHF%��&�իl9��+ᅉ[��c_�H��P��f���\^���Ⱥ� �g��9A�I����!�gf'+��t)�a�B��3��*]]i�
�čto�LvᱻG�\q拊�m2����M����C[kP�?Q�����
���G��2$tO���8p�c�[`��K;V���Цm3�,d��t�����u�8����&Zu�RTW��놶'}һ8��^�����f|z��"���������A�T�*P $9T��A��73k��Ldà&��!9�M���5���L�qE��E��o$Q�]2ښ�旣w�\|B�g�!��&
��c��]~3����s n�����=������9�b%O���N��������w#��o�*�p�C����X�i}�V�*����)gp�z%HJ'��΍��R�����:���7����C�Aʻ�Nׄ]:̵?�����~���l�����º��}ѽ���T�Ef��*~w1�(#��-ǐ�x�繗6!	I��'%����Z�!`��T�\���� �������);��ʮ`<�K���!�S,7'��:� �24�y�%ch�>��.�����TZ�,�3
�fpi~@Fc����2�6)�IG��#P���ńa�7�P�~0�f�Y"(����M��� ��[�Uڨ׃QE�E��U���
4�H�IP�c��2t�	�b�5���iJQ<��tRܺ
��¬��%
7Lhn�$%fPz����&}O�i�5��X�nr[T��jnoI�<�i���vO�!B��G���%������x���*E��v��F؟ }���kQ�щ;�ZV�i�����|���m��Ο~oI�򍘃�u��)�0�݉
�t�Sꕜ��HCb�J�!\��;�4��=y�G�j�%����̓Q���?�'�M\[H\�������P�K�s=�������]��a�*뇣M68�%9�y�L���<-g��,����6��'��pQ	F�M��'��j���ǹ֯,�ۡ��Q�/ͯX��=Ҁ�㇌�2���y�W�رu�y�1�^:0B�܄�iv���B��u�u�jc��K��}�d]�<��@oz|���KNB[�A�l���J�g�Ɩ�]]y�q��CP�]R�՚$��GV<��m���nY��2��%49�]�s�y�*� ܣ7e���z͠�n�.r&X+~���8Pw�֨���UaМe� ���j�����
��z�	n��=�N��x�)��$�h��)�q��ֻD/羐cɡa>s�5��mP��=oZ������s7��q�#o�}8��� *�����%qD!g����J����A�,PX&��>�����N?>k��ET覉��pG#OUd}"�u�ϲk1��s3!Sĭ+��i
 ���$�2[t.4+L;���V�S���p�h6!�l'\#�8���ox�`<p�m����mҴ$k�%���\D��e ;r�wn4+\s���u���Ş��G��������>����d���N~N�\��9�S}?�o��*�K�V�<�����OAI�0�S;&��&c{c�~��w�\�py穻�X�K�2����55.y�U�
�96<�ä�: �9c*l�Њޭ��t ���}�~1����hX�aO�?�\/���A�ߖ�L��o�{�Nt;�U�2L����7���28��ٍ1Ǟf.�NU�"��]kN�O�ӚG5�� ��(ZR9�q�L��_ɰ������r����;�����$�����r�X�r���6�'T�;�e�����p.*h�* W1du���%��h���Z14��/��� UY�J/�Bk0��~�Im����n��5 ��a���K�4�Sȑ��= M��#lz5�F)>�8*C�K�>��ܬ�����H���zj���L��Dc���6����6}�E�,)�C!p<���7��J2'ו{0�e,�V�|!�m��2D��{�����bN�zA�/��l�?:jCE-9�W%�
/?�0�I����y�ݪsM��vϷ�G��uxM���(�v��}ENާה��d�/�3�C�h⹼�%�{�=�>�Of��!2�-h"�46o�r��L=���#�����c*5[�h�������w�M&U�TN�&C��;�6x$�!Q!�3�2�\b��R�	�����Vk<��;�����A�nǧ��`[|�N|S@��G��B������uM����UFc
�m�v�cG�B@T����
(`	�z�CCq�s���Cs�*������ꥫ�d3c�)p=�T⒊�g;)~��n!&UB	��wK�xxQ5���i�!4���4���=E��c�fbdd�`�6%�2Ҝ
�(E"l&.m �=��b���kL���ҹI���@���ȽLM�_� ��������D�id�4�)�J�&g؜���?`a���;��΍_���U
e1��7��̨;��_cc�_�c8�.a�-VXj({��L�g��*��X�	.����V���c�$8R ��8�y�e�*�c�`S�QS����#!��k��k�l����r�-ќ�ɷ������f3�uvR
�~M�o���Q'�,��L��1g��E�zL���P�Q	F�iхɤ�C��-h�<��������U�E���|���`;<�~z����i�G���_	�s�>��}����9'N���c�hZ�,:x���ם� ��� ����>_�~���J�/ۇc��.6D��td���~�B��2d�ӱ�N�I���<]"ak�-���Q�c��U2�"�(NL���^�A�5���,v��8ʸ�^��#�ز��i��]�uؔ��G�\��mɆ��\�{�A,����6yx����d�3���m"*�$jD��X}f"�C��wiw���#���y�@�j@%���z^$�JU(
f:�,^�c4���#N1Ĕ�NejW���|i�W.�F'�v��r�P-ĝ���q�Ę)|<�b�%�qF�n���X��&GH�f�;Ӧ�?}�~`SY��AFA��5����Ju���>���sv���h��!lRs
Nx�8�Z�k�뫐��0��V���S:>,<!n��A	�ÈB|�B���ɳ�HxɅz�~�%Kbr��@��������K,�d��oL.�Ye����2��� �����3[�'5���I-�5���E(!	d���Բr7(���6[�e�&��", �=��/�2�(�N���&ln���.^^��I2=9.MU�$�Hq�]�p��v��ë���c7�k��^�et�㎄��p����8��pe�k{"��U)�S����gAxN��ʜd�Þ����	BC�����.�X�&)�Be�ZN�NQ)��AJG�_M�F��4ODW#,|��
���a��]��U�X���d��!n�az��`�ֵ+�qedY1D ���ۦ�#�y`�Qa0���,Ǎ���ԛ��ƫ��*��k�*ҕ��˪�9Ɍ@x��
C�������=t-�DV/�n55��}Ó�\D%�a��mת�����x����ᨊ�Nur�ibo�1yAe�R��k�jѡ��h,T���r��/�y�Mx��+��?�N ��sZXQ��;��SH[���}�,?`�RE�������_��[��Sj��ݔ�"����,���3��T~��Lѹ��p�����A��I@"�|�0S(sC4�P��ThZ�(��� �Lڰ���|�S��(lI� ��<@����-�T#�.t��u]*%�c��'�����Z~|Ðp����j'��{Q����݂��r�R���͌���>K��@��x�\�;Z�3F>DQ�W�
m^홯"��.��*��&�Dx3GE�z�/����ӿ4<�t�4�N���
Q��f%Z�c�/?_����݀�.{ɭ��GYҺ�3;?�v�I�G����,r�[R��y\[�?k ����H:��?gZC�����2IT"�	��ÄǨC7R�F��@[��0pNr�>B'�'�u�l�xH���SƚM&ي�g������,����H����3����=E��k�V������߻��~�W'new�T>�݋m)Gj�}�� ��P���ɉW�ˊn�f����䧲�8W��5�@���2�1�����t`Bx�.(�]i�|��YA�h���^��=[��I�V*�B�J�� ~�A��)�a��Q
��onZ�
߲��aV��!���X�;�-�g�w����~���s��̩�޾y���#�U������B���L�v[�����H=>�9m��(Q�����/58��kR�3�% t�?G�-.���M+3�]�|��Y�fFF��S;P��"%.1�<�k���H�t�S�ڻ�#цX3�?��ȯ(��� *�މz;�lT�jd>�>I�sy�oؗ��g�o̺��4 �z/oC�2��Y�	op4��]L�ω38˶�e7V�6����7�WT�0����-A��:�J��Ib�E���vwk����$7�����pQ��;L�� ��;A��T�o��yDB�`�`9�vz��*Q�J��U�36搕�b���G���n�6��M���2-Y�+rF����v߶rA<S��M�ir��C�p>��r��g��7&����L�G�3ΓO+� ���fT���vz^�)۞[L��L�*�.������KL��%RR�/�k��r�ŵ�yDQ�v�n:$`6ҳ���Hcտ�u��F滘:��.� '�Z 
F8�����)}��W�M����3x��dw�W�I�D�b���3le'=u��3���D?��Ug���,Vv/J���>����@[��,�T����_���´Lޥa_�B�׃U���	�e�D�v�
�T�v��.M4��~�B��b�lw��� Θ��V���"iF���]uh�H�!�zc5����G���/#!�#�]_@p�NS4(�\���¡��b�V��!�n�
��h�!4��p|�3E0D� ��˗4�?�^E�\��9�q�H\��`�{��N��u2HR�ʹ������>G��|���2ߪ���6���cȌ~y�ҙ+]� �#tޒm�Ùq�ف��P��1��z7���j��f4��&rd6�e3�4�v�f�G�Ь��д���[����1��%�:I�;���ү`|�۴H�!s�N23,�5������a���F��G=�S7�T5��X������?�9A�Fs�Zm� j�Kj�"J��E&!W��Dm�w�ځM�@}���27 |?�t��~�R����`����&7��$�+��R���pa�#�Մ�ఴ�"h-7�^�&!��[J�T���ci��Vb���Fͥ�J���/�2:���cul�$��rZ�`���M��" 2-J��w����u�a��ZP�F�v �Y��l�(x�H���-�L�(�E�JY�	��^�eXq�z�� C�a�Cˎ.bVJ���: }�MC��͈Y��PWA�v�FehHN���OI㵓�=�r�Fʣ.�S:�l)��:�����CT�;�_��@WL��ZS�T�NrvH���'5Ğ���-rZ��C+�;~F>������)βي�U�bK*�4ț*�wκgr��RfIdmb�++޵��ƓNi2��i�YAӼ|�KMdq�mBzdj�B�!���y�*��+8��?������B��>���\O�(B��2��̈�-S�/�z���������7����5���G�ʪ�����w0i�]d����C�R�J;ϟ��ϟ}Ȭ	��;��@��iKZ
�iT����ɘĜ�M�$��Ҷ�1.-�w� �����'������O�"��������w��t�{�6�;3�]��#&D�����O���$}&�2����g��x�C�&I�_"�����&���@-
��O�Q�+1�}ïJ�G��1]�8	F?"_6Z�w��%̌7�y�v�=��N%l}���+�r���ߖ��%�"�6����:�����Q?Dj���;��*8a@e�l�0�%zw��H�*4P�PyFCu�fV�̨��1�+G�V�,�s~z(?dm�*a������z򀟩�؞R�V(d2�F�_� �V��r�}mFl}��Ƚ63"����y�HKS��V��n1KV�"[o9Ot�]�	�i��5{?PrW#<�֒���� U�2|���Ht����u)�0"9�O��̑�&��n,Lݾ��~z����N;+E��&̔~�J&'�V
��ф[���6�3�t�e��0Q��l��Jw�=ۆl3|i,k,�N�ѲT`>>��j�G9k7�/"k����$�7���킠7�hֻ�B���S�#�(2����a��\����n�ћ���^�Ń(WN-:���xT�4���FH|�Vҥz�e��c}YO�z� ������
j=<l�v�^��p�j6I=j��3��+}�)T�
T�����S�0�pG�z$�wr�R/t�։M<�j?-�X�p�dߖ��3���m�f���{}��g�i�{����u�Sp�.7�?� z�ϔB���m�\~v�,��Єm�[�{�;}��5=��M�S��� d�����S�9|S��:,\ �	���.?CR��g|`����u��$ʺ�q%��0_BLX�.Fӄ�S����)���z�Y��I��1d,:���z*�|�^Е	MSc�8���:qk,a�2z�	����dj�7��,\bEq�T�h���~�e8&�{�{}1"����aR?dEC���� ��qDqX��_�� �&��C��z�n?_��,ʌm]�!	4��1�Tl�~!��ڷ�* ��a�(H�,�@��|wAO,mT�񴫚c�8�S���P�� ��N͐s�L���г��n��\����R]�ޯ�7vq�ߜ�B�OmyE�H��i�×e����	)���Hr�8^;x�`WƜ2Aߢ0Y#9s�'�������[(ǟ�����XY>D���,���#��k�e2��	c($�˶������{����Ȕ���M��ۦ�f�88��o�,����_ង�O���	|�p����~�~��ox\���7.�aBcuv�Nd�a�*�_���B2�y�Uz�������F���)��
n����
p�;����*J����&���g�7�I�tO���)@��<��tP4^�1�YN�d�:rS~���Q[���]�
���uF�F&O�'��-�<lg62��%;[hW� ��#�?nI��W�T~T���!��$xܚ�&2L�e���p�w�K�R{�(Qj;��G �{�G�㨕��M�.������YyT�Z�E[��+V����f�%OR���"��_[��ؐ�Z���<����j�Nj�d�����	��� ӏ��:1���&|_��э�BTo��s�5���TN'�k�gl?��(�^��'4a�wa�Y(��b1N��蛑jW���$�0+���	h�)�o�͍u�\7	r���h�G;�E��D,2V!��߭u�6�[�'E�b݃W�v�op�>G�Ot��A�xk~� ��o�q������N�f��W���+[2i ��q���=R�a�s#�M��Cy1v���r@�{�m6	�5f9����ꆯ�|�K1	Gj�R"=����r�Ǝ�P!�K���焠f0�^��h4�C��K��U���U�3>��xXG`��K���-W!��ڧ�ˬ����菲_��x���:ڏ}�R�(�q$�Y�4��(뼬��~IT�j�� �B�n,����+�c�q&><���L�l0���K���a�UB���3Go���B� �X���[�ƕc;��1�.�eZ�E��U��C�7X���P��L�O�Fݨ�Qe��Uf�0*��A�gت�Q.'/�wǁ� hPGc�yT� �}��V�]	� G�����  )�4c����Z�����i7<����f2d�qv�1c���Wml P����H��os�k�͎v<^��e&R�"��`,ޭ�Pb^�	vcn8g�~����$��Ԕ���R�5��h��x�vl�ݣ}Ŧ�?�rؔxb���	�|ty	c^(�N�^54�.�e���=�?[��]���/�/t�C���%�^���\�ѰV.�,�Q#s��pʋ<��3�!�Rg�/(�(Y�MU��^Em�,0
��)Y��7~5���c�S�{QjF�4du��P�sB�C���pع�N��^��������4A=6+qC�gS�}�\��64�X�� �,G���_4�R���e����"��������ꋦ}$>�M�=<����B;r��!6f%��5���A�G�����	C1T��f�D_lNX���[GM� �)�(1Fq��aFg��;ZZ�{��>B��o5���;ӳ��a�����#2^�ir�,J�BG��v�x(�aL���o)D������D�ozS�:��UU��0�L�Ҋ�?�I�MW��E�TǥlqO*���Bj K��P|LO���o�@��{�e�ؗ��Ob�/�*w���^�O��"WV�yZT���/W�f�{@> Gߘ9�����B�Ρ�p��0_��]�
���)F���j>�B���-�� �P'�d�`��>�[�Нdy��$'�[^��Z/ӹ�Bx?W<F�a(��o�~�d�H�>)���#o�7t�8�e�s��{:فb�~�c���D~]��L��P�.$J���+%P��*��~����HW��SNJ�ҡ��n!��3n��XJž1O�F٢$��.y��X>�;-���@@�C��*�1��{$��H�F�N���^�eL�YI���9₇f �+qsi� �L����b�wN
ϒ���?� ��c6~&1�՝����\M0�s@���Ԟ^�-���':�xk���?[k)���l�]���K� �.U��8�M���.7{Z]�7P����ى�%ǫ}�:Ly��	���h�/��*�8�3�e3���5�1`�������X`��%
�Uu�L'��"����%�ի���َn���	&	CB%x?�?��l]%ғ]uٵHy���X�]������e��n�ot��BC��sS`:P*���]' �ģŲ����a�(��lͻ�&w�N9���o��� {u�R�;hk��n(&�RG��#Ӌ�O��o0`��]|��]��%��u��[�n�Q�1��!3��i����>����5��f��N�{�EPH���'W��#��;�/2`,�7|PD��S����c��yd�:P����+ج�!=k�E��	��${ml���T��Z"�"ݳ\/a�[�l�4P�V4a�!�6��r�6�e
npy�I��R��a�U��Y�䏐���j����H��F������(Q�gt�"e̓1�Ӟkਕ}��9��1):��D��Y�Y����Cm% ��[#����Ć�A~�H1P�R3��O��X�=�4�����pjÐk7W��lX�i��V�z�g4}�Κ��7��.F����xy�#���w��4����.��X�n�*n=���hi8���L���x���qG;���.�R�: ^��,6�N��ȇo1���e�KBJ�7 �Y�o*�p���s�����O�p	Hݖ�Lt�Y"�\�����:j+��@�g���nY˒�%�ڴ@kk��Mi{:u7�)��͡c�%Q�m�"9d�=���
�1���?I��Ǩ�݌���
��22���&uF(rR�������q��-�}��-�e���[Oc�أ�;*;�!:�K�a��*��5
q�߯�7PI��] �̩�6A���]�q ���^ށpvr�&?��>�}!m7���QP��$����Z���x�2^�g�y����]<SH�	���&9�����e)��qk������[�Ç�$7t�D�:��Xia
p`�#��]s!x	'��c"v<jVq�`e�Hz��h��mf�O%�a1�(�Q��ÒW��d�7���1�����]��|�c#�w� �m�f��P� �f	k��/lgxO��Q�D`�eF9P�x��%J��@�uzanF0�5�S��Z��􏢝oW�|f"V�Ĉ1n�ib����V6�x	~FY��-X���s��S2�ę�9j)���=X���͌qL��" ��Ś��=�%��Z�3Ns�� N�g��r��,�w�w侊��mt�$Qc���� Wh
U�m����<��H�4�P�Ż�N�1�j /�|N�������ȿ�擢-Y������rh��,)��=K�|������
*pmĔ��z�m\�S^f	���2��y�q}��x�/�އ4�G.�_<>����Z���-4�>j��]�F���.?���qn����g��w<���ǶV��R��?.�Ƥ�����08,�����`���]��ݠ��F�Ո�������:ld?3c��9��{�>.���n�A���.�UĲ��G����B61y#ؔ�K���^�{���v u@"�,�ӥY����=��9�����}��v�BIF�R-��0�7u�^0&[�N��߃[un�df�lŸ爺$l�15��W!N���c3.�#5�3���$�ۧ;��4�K{Mn��2Y�0����,�'m��(����wm����K�b]i��Y?���`ܛ�ɹ� ~ܒZq�� �����h�g,μUn�Z��x*peS�H�'��V�d����α(�5�@�}M�_@��4Ž�$H���.ɱ������AJ.�.���g��_��1��$�D����#����yp��)��GU Y�Ca^�v<{���q�*���u*�Y0ydZ~g�>"QC�6�ׂv�i�_>|�i��8/����p!�w�`E��O�N�w�H�9�}wR��H*���\��U@�q�� �͎H䳘U�W&�
�+{Fw뭟���06��},�2�,���+���/���]���'=P}��ʆ7g_���P��{�P{���\�VG/��� ����I�
�?�Fi�c|��݊[V�\�S��.h�37�X7_5;�@�y��^�<����D�w�Vdz��X����;��Ə[�����B�ъ�g'��وNp7���d;V��ɰ�C��,]i�a��1������v&��A����ja��@���/F��.��XU<�&f~��EW����'hƁG��@�eg�\;�hy����N-��������9�k`�vvD�Y��B���䜠ƕnr@���;�܀2�$T,ġ
��~�l����~�z��)�<��O�	E���:����[�;�J�`���4���)���4k�E���R�|�z`ٯ2S�qp��Z\!ӑ�ɖ{P�uz��O��<`j��)B23~&�χ���L7(X�o�b��8sL�]1A���֛	6��k�?�������T��0�R/�]~�����tpk��������$d�\D�yB��b�d���/F?^�����B{���
gĿ
�oN�P��2��+	�H�۪�N�������e���$�RX/6�[������F�VG5�:/��m�M��@����zM�E�f��F�=�^`�'�� (�z�؀1��X��W�h7Ӂ��:���Ҍ<{:P����}����YG�5��_n�WC7�"��j�(����������XY.K�?3L�I�r�ZV$�����0�])CF������1��u8���Y�\2��e�!T��	�.z��!V�^���N����4�ȉpH�N���厱������F��jۧ�fu1f��F\^i����G�D��s���T�܁*V�
���,wz��S}���{�7�B���.`B�ʿ����b����[Ş�Y����L���RN�MwL^�2S������+r�"іZ?uH2��
�W�|��(�Ҷ�=)u=��ق�JN�=\Ђ��(�+�7�*��K�݌0�Bţ,ڢ�,G �������E��q~q�)LDU��}����/��*��r��~�_9���V
*"�s����tPf !��B�'
��O�rF�����x4�)T�N��9����J�'�����[vN1�)Ɲ���%�g⏙�� qm�Յ_ö:�_c���^��m��ވ:;�+ɻ1�V���l�`+̈Ͻ����3���e.42�!�a+�x�pt�-�[�-_��_s��cs� ��-�ÕN��<12��ڣ"i
���A�ӓ�E�f|b�,��)	]<��4�˂U9�סKL��nĢL���'D'��I�aa��6��AuQ�@{��!�]E�D�`FI�������K���N��16�h
�
u��F]Ǳ�>�����p�̾�ͣk���r	���L�A���k�Y�l8�\�9@$5�c��߀=w�F��g��4���F�w��G�T����0�N>���'t}s|X<�ɑ@�����Ї�]-���IyuW�|]��é��������]$��(b�+��G;/Y���/������a/u)I�Y`kO�VJ	�+�Ĺ�X��ʹ���ع �|*k�/���Z�ҹ9>t�#��
!}� �(!��f�m�f�5o��ߪܦ����[���`�^ĩo���|+�6�v/���#��*>St���W�Q�`X(�^��-B�;��-�G�V��>p��yyZE��~�T��4�%^���8�o��{w���8[y��J�O_��1s$�Q�������J�����`�v����L��݈�Ok��D����	����!��WFl�vy=r�2U1r:��� �iC	v�rG���t��o�@��8@��.����Q=m�f��b���=͔�oڜ��j�@�[�½p۱�)�0(�Q�YQqg��(!D:2�L$Ѐ�Gnc���b+�V�]K����ߒ�'S����-�x
�DsT�&ě�tf=��yy�v�� D	|�Q���f`��sz p+��AL{s�t��!��/�P��>���|q�H]A���>��W[Q�+1<9��k��h6������J�N�[��6r��g� �<�dY=����J�9�}��1���w�t��:r�� ��^ͣ7R�:��<huwZ|��R��f���Rf}��A�Mb��xc ���U�gA���T��+����b��1s��d�N�+����G�n��+�_�{m����/�����.�/z���IiH����ɐC6yB�7�;ՙq�m���ÞG�,���7��P	��2�5s|.X�7�j��n䫸����Q����2�M�D�+VKO.�T݃��>��ѐ�	<�٠�ߥ��Ό5=G�V�It3F]�uɏ���c�-`��x��W�t-�"d��F����[O��ڿv�"O1,V�)Pj�(7A����\Л�fA1_�8Z�	F'��#�x�V�ޮ�H��a���s^� ��9�z�g�M`0-�*��倽��K���i/F��V��L�D���)oa�Ud)z�fښ�{���2]l�������;�@=�a�}���t*y:2p�n��\�x�9�$�Z���e�~�[&�v����̓�A���)�=�r��%�Z�5�(3x5Ǩ�[6te���h1���y&?�y��!."#j��d�L˸6}��K���i�7e4 K\�(�A�a���7\�/ǘ�������HާVI/��!��l� ��v��H�
� �4���hNtTS�9+@k�Q�9��
��so='���pG�Uw�����t�ꔯ�V��uh�`��)EJ�Y�ZK���B=攡pXv-�X���2�s^����1w��ny�J�Ϫz���3��XR�m�R����Ȼ���v�sλrٴA[� V��q�rb�>'gG�Z�IU*P:�%]�8���oҵ��,���3Q������"�,�4auYl'
�����M"��Q��#��}*��6�O]���Y4NL�"5��g�*+�Ø^����^{z��c�����s}�X��D��_���iB�P��1�H55��*|1@�ū��R?�4̣|yg��!oJ�/��Y��5��lU�`��Z���3�(ʧ�b��OJ�ح����]�\�L�|��0m�Oեdp�ug�d����m�uS��Úz7ç��t->
x5�b��r�U�O1���j	��-jh'^8fY�M�Kl}r�D��بer��(��m��e��b>�#��`����ڞ�`�癄�K�"?/̫���G\����j�K��	 =K��Y���q%�Į�Q��Ǳ��Y����/{�?Pܦ#g����B�
��tE~����ˍ}���4�,x�	������g�8�H"�K�߳��?�F�f5d�k�&p�+Ŝ.��G��`���X$qX@_�l���8Z2p1@����KUpPo�5B��ݣj�'ߛ�4R[�E�S���8�_@���
b.JJ<���,/��.	AFty|ғ$y�*�y��h��#�M�'�u*��]��	�>�G쯑�0�6՜��Nl�/����KKE7� M��Sܒ�i���#�0h>MX^=�I��vL����)H��{��Ee|d=- �UϒIN͝��d�Z_޶̺�W�+;��c`Tz�/z�aa��k�n�#�����B�4(�C@j��!"yH[�d
�]���l�C�2��oz��	*�~XUL����G����8R3���Ϸ�c�a,�x eE��¹��?鏜����_�� ��_����x�=��r�,|��*�g��5�Ey�4r���m��ҕnOdJ�3b ��-$�´�vlp�T��f&�<�C�L��蟣��I�I��o	)N��Zo�Y+lOU��ur�{W�v<$��E��|3��{��)˚��'�i���d� �G4&Q��qGT����bS�2���An�ٷ��9�����D��B���6���;���f�ȟ+cF��XK�.��o �F��'zBn�JN�g(���,����1��Vȉ���Hq�q�&�o��D�z���l���~�QI�q�����w;�+�BW*,���ֱ�����#��6
B��A� 9�˪��[<0W7��./��fy,��h��G�����&e �����~��@�>{|
�e)ɂ�ʜ���Ԋ��p��;3��e�4�񷍳+�v��{AC[Iz��g�:�*�>"�(C�@�=�ϒAk�B�A`��01�%�i�<N?E�y�:g�92F@��)�5=O�M�Zk����ߪv��|�^˙<u�͈E\��x Ik<�S�j�P�u���,@�{Ô��X�k�S�2�/2�����q/�	rHN���j �r��'��ô�to�O��¸N�S9�G�aۛ3�խܯ�R�u8��3��݃�N��咬X��P6�o=k-���!Nz=�xLϱ�Ɵ"�,�$���į4��t!�p���>�ɽkNp|�L?���5�R~�:��	���M�|GC�SE��:��:���3!Ŗ��1��#z��p�Y��{ᴦ�zy����D'-�WŻ�ݧ���gc;��⣖�vT�z�*qY� ���Bu�/�I�k?S4���*��������I��Y�6!1�~zݖ>^� �x����;J�d$�)*֙�0�D��bvC���k�2'�n��q����<3����T�����P�6���Q��p���f K�bYqq��9*�ۇU.��z	��o߿�0����ۆ>�WM���E��QTb�[k�4�.�s�I������|U�i���:�p&�4��֒B��-��ꢙ�
ا�0OPj��A6i>���yz5-�Q��9z$��"�Ս�T�d�U��:�j֎���$�h�qhZ�����,�HA��u�(���֮��6�C�g^P|>oWhYS��/�P+�X��+���a�Ϋ&w�+�&�5�m9mUF
�R�6���E0�4�}Ud�[v|�'/�w�s��@�{�Ц�����?�2L�G���S�R���D|g�gڿ��,��ڻ�������g3x`�fRFM�@&H����Њ�f���[�0��%�3��w%uHn�c�Ӄh<E��u� �'�%|!���32�c��^�
*&�́ܘ �����|)����G�������ˍ�2�X(EObr�b�O'�zXd� /Q�El_T��vX��k��VRjDB��!��Qe��"��:y~ �����]�3�ڃ�������TW��99<��,A<�+��l�#�5������77�>$��
^0�#W��_0�qq/MJ� c˨���AA=��)�B�@���@�� ���J�\�|ϳ[�e4��(w���a��2��9�3���^�H�nJu��<'T�|���������Y-���J�>��Qѹ����

6��e$G�Ԫ&�PC��|���6�~`�J��S;x�Aޔw>����'�9�*]��JH�CU_�D]��
��z�5>]�NA�Mf��?Z@����kA"J�'V�%����+��B@���<�L7�b�Ő��<�R6�m˸D'���62龫En�:|�M(~q��u�y��Y0��a,�j�L�t����`�'r	'�$�����Rpp��3��]����V��0�ƽ�*N<�X�pƗ�c��95����h���4��/h#�@�;-GX3��wdM_N8~z٥�I�����(��^�k��Z�G:�d �����vf��~�]L���v@ ��C��uX�^�r�]���V1ⅱ���9���9��豽v��,?h�-j�b��X�yZ�<����[�Sw���BUJa�/�|�� ���,��K�$:�7�ٱT����m_t��\r�"����Nw���z�F;WQ��A�iV����\���)�z-:t������=zGN	���&�!Z��	��nͬ��:
[��P�d�p��Ԋ�u-��*0py�w �ʰz����e/I�[�Q@Z�5�r� �-��]���i�C���۬���e;_����t6�G��lԭaX�h/G��H�
Y����.�,��������u�Y�01��ue�)R�Y0�Ņ�߼��MlĦaݩۨ����R�@7��,S�_��z,y�G�y��v�L"{��c��r��`w�y��Z��n=O�]�R���K�.���h��G2�� O���4��sh۪Zd-pyZ���{US���gc�&���4������ޖ��D�4�;��UY<��ء ��0ٜ%�2j:�T�A��G��vʾ�^�p��Z߻�C	4T=���i S���i� ��e��^5��d�7瑴oTx*\����O�w��a���P]�-M�����b�Y�9���Y'��������/bEO^��?�=Q�/˷�e���^�j���%�GD�L�wq[.P
{xT>���_���2��^�Yr�%����ks.^0��2K>���$�+�Z�
t��b�6�7с@��jz����""/#4�j՚�ޞmg`�ai��HZ�Vb��{{!h�QF�^ԃg�@f�4�TD�2zB�C�(�4��ǟ���
� o�a/��K�u�����ȧ/ϱY�F���^��jeι~ΑvqNn�ߋ��5��w��jlw��bH����3e���N(=�V��ro��@�����8`�����m-��'�R%���
JM���>v�����E���U����!�a|
P/9/_jV3W�-r|� �� o���A��'	�B�x�<�=\әeF}�ҟ,�'�Ëڮ��:�8I06�1�At�!T��~�i$ riV�Sh���.����9���_I� >���L���S_� ��t\�
�m	�@�A�ZKbXz��'pS!Ic�	��ԂQ�OD�r��褼��/���%`b|Y��,�1�S�36CF8�U�@��6�~�ak�������j ��C��D���l�O��Id�����m��W��0�@��률Jj.+��sO�;�\KS�� UQ$/��B|��ג�F�ߥ�D�x#��9q��0!�p��(�K}��W���v�2�t��Uh�%�!����V%����t�ۼ�qœ���0�J+<s�����K�۶Q�ۘ����8=~�)st��K��;W=�m֋'�Ní6�۞�5�[