��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c$������;`�/ ��!�z�����͆�pRU�uz�j�g���;�bEh]\��L����Էek�?��&Up�2)P:�9�����W���\n�7߮�n%ziJZ�H�!�5hR��m���} }`	^��1�a2Z&�Q����?�&ǶdFN�����Ew�]��4=N=��o��i�Ժ����c��=׍2@�ϸ���)�œv鱨A��h�k�+<F���	Q6��:��/_"�D�EW|�݂\�7ڽ0��{�Ԑ��~�h���C�9���[\Uc�5����,�}���T<DDfL�7�T�V�{Q74&A�+i����l����tI;I-{%��﷡,�$ް�5�X�wŀ�+nc!�+��G�!�iZ�\CK��wKn
c���"C�uOן�z
�\1��"�s���s�v���O{3�|:�}LnF�9���jb\]Br^<k������>*�h��S��v�O�x����%�`��mH#�l�͍�Hh.�nb^�O'�5d)$����Q�����+�1����,�R����ү$l�g�O�<H�:�K=_C����[}����Ñ��4�dI�|h�f�-
K�b�i*$<�g��S�A��fl��^+`Ƅ��B�,n���}i�E;�:��Q���*�}�4�z��#�8O�zv�,�9��fd�0[#>��je��_Î�S��%�*b��6��e\p�ܒ��שʼ�� e^���m�M��O��La���&�5O���WM5���B��i
E
o_�}�BDD����*RS��� �w��6��}��0	2C�4H�oN��o�2�[����e�V�Lq�K*�;UZ���Z�Y�3��mQ�m�h���}��a�%���"�D��Kt�)�q/���MۥZ'⳹��OIp-�5��\.ܒ�y4,�1�%%hoN��d���s�����rK����|"���~���W���_	�I��"��P"�vcs�&@���k�����f��o��a��0��u�'	��x=�P��`h�0�V�	a �F�S&I�5�ej�H�(��'Yof�Ts��\�@
�N�#k�:�o詅E�vaBe_Q`�oesI���D@�u���'�g��d� X�WRT�������!���X�(8p��@t�J���ⰳ���n���B�����<2��x��ae�.t�������Q�� uVF T�e1C�B�G[Fq��sh��V�En�W� ��c0l��v���
1$��c��`H�K<|��+��\�]%���W�mH��>3�j�c݊����j������lj��O8A5�M\<Ml��qB#w�Vid4���,^�Ț����\�9ܗo5�(K�	�f�3Gg�gro�"z� 1�H����=���S����Ǫ` �(�K8sT�v�t,yʚ��Tb�F5�|�	��D�W��boB�wS�	�h���)�B�Ü����OybYEQ�R��:/�_��t*�[d=�M��G���S���q}5����.+Q���������
��@�� b�:�6������ҁ�K?v`�b���qhW���N�ʮ.�Õ�N�l�Ğ2b���X����aYV�^��Ch��Y�!���ue������|��1A?��ɚ%!�޸:) ��)��}�'���r��
�����k��2^K�5i�_F��f�y��xD�_Jl��Dq��aB(]��d�h�O�����r�$$�#��T���h��P�nw��s���۾#|���X^e�_I�r�0� ���؟�{��%�PdbkI8E�q� ��쪃Ϧ]�y�uW���Q�U,�~@s(��c�}ɍ�4�"�=nX��\��zn3m�1��>S��$�`�\�AŜG�E�E�7���;P�M��I�?���N�T�ĩ?<�ͺ�]�Ve4?qJ��cK����tD߭��2S�]5ZUP��{�/S�aum����0����,��P5����G��p2�k
1�� )+�z�ӿT<�ܯH��B��G�bry�F{����	��;-�L�o�h���6d�x��7�e�����`uY���ÿ9�h�7��o�U�}�0yL/�u�����b��(���
�'�����x�\M���"�]N,��Os`|�jNMg����J�&Y<��9�xJ#��6<�N܊;�[��BM����3������ujH���K*���~E��~��u����r��6Ͱԉ�0����&�[!�.��y��rME%��+6]�� ���~o�judW8�i�4�v�@z �q8F=��5�"�_�x�?�g��*龝2o������@����ƣ�Hܟ�����E��h�����B��Pn��#�K��p��|{�/�q�%���ٮ�����0����`<z�ݏ�$�]hl����&��L�0c#��?΢/���4,�<}k�ا�u`4��R=�,z���a+z������@��n���y%��V0����Jt�(�J�@� n�u8$ ����M*g�i�x�L8ګ&Ovp�>�ݒ�* �D�#܏,�S��Ƃ���uA6|��
Z.�QZ����,|�Jj���x?,I��:g���%k}�D�!r�ƛ����0e�k@ǚɜ��q:���{��M&�p�*n�T>�OI�����$P�gJR��a���������J���c�L�1-'�7Ĝ�
�oXE�J2��z�����C��T�!	��B�π\V�~%��7߃��
H��WT���A�xҀ�K�|��#
6i[�ї��r�v��}�A��u��?%Js�<
p��u
ɩ]ն��D�$��U	�č%�?
��1�wd.��q���2l�Y-˓��9u��`]�(g��q�G�G�9S�B�n"_���.{�,1��Ҙ�t�-���y�B�ы�xn
FV;f�s J�xw#hr���>ו@�(�y>B��?�t�U�o��i'eJL�U����DC�V�|�O_�4N�/k��N;��[��QE� 7֖)��ʄȅN�N��$IUWyWae�a�h�$+,��bK���%�2l��Y�v�G��'�Y�=�B�	��Z���M,ɑ��K2���|b8�dT[ig�n�݋ٜ/+L�d^��z�҆�jY�:ѵ� !�+`�H��
�D`�v��Lz��b$y�_�L~}�8��X�S=Ձ\)1@�S!��姣�&4Ԣ{��߹�E'+�����c����A��e��B!�k���#VbF{??��H4��q2�A9	B��l>����Xm���5�\�X��ߴ)wfT�q�����u���� ��*^��W?��qȿ�Ӝ=����:@���Z����gM(�s}:�+p��oÛ��7���j��d�'���s8r�;���0�!�:C��&SxΒ�#ڍ�Jȥ�	�~]7Y֡D��w����Ɉ�[:����G��D��uTc�jo�c���b���T eI�!�R��8V�=:@�1�"&�u�o��t.����z���9)���;���Ug� ���dh:u�δ8�m�W����G�Z1��>�ӑ��B9)��_��$�-�UoK�)3��3̸� �
0�q��S
$�-��	&�h�\h�P�ſD�����C�0�J72 G�p�Ȇf��
T6�q�8_�#�'P�2�_P�{&[W�����߁�W��o/����G/[��@����ϔ'v�lOmTI��R�pj
h=���wd�� �Aۜ�X%i]����%`��^f�\�C����p⛤�}g*Wfȩ�Nh<=G�"��K�rl�m�DT�=���|m��@(��d< &Uz� U�
�Bm!gT�7"�NeH�g-��I��~�k���d�ٰkM�X���JO娛����w�Ȱ���H��1�qI��v�_�F�:��]bIӘ¢���"B�as��9�qT37L����NɅq�;��b�# �3M,[�����-��9�4�a����b�\�"<S��Yp����	*�#	Q�Σ�n@���|`Ǣ���+ K��ڞ]�Ӧ���mS��<���$�	�G�c�6��ˆ�:Կ;�"�.cX��O���+,�ח�|��w$����ㄓ=�{זQHi1�e���	��q:����|���:K:�,bX���c4%�I&
1�El�]��j�.�u
ͩ�5�_�yV5�J1w+���]C6L'&{7
n�C���K#3����)�f ҢF1g|�]I����v+�*�T���	�S�`WM��AE�<�}R���I�-�	A���!�@��=K=j�x���!aU�D�<)#%�Л��֦Ơ����[�+; 9ֶ��2ah�(��`�b�F��i�U��D�XBZ�Rɘ�[8^�Gy�:6lV`��R�����AX���]u�L��-9�ݰ4�̐��(��o��":Y�6�݋T�}���.�*\���ݓ���i��U��&�� *�X���m���Ou[i���f���=��+��R%<��NNs�:&�n�e��]<�GZ��A�����A��A�0�N���dQf��=7CV�@9��ƾc�>��;j��O=�6μ��:�y��у,B�6�'ڂ^1�ˑS���b*3&�٭�����)dn7j���(ߐD&��#���(O"�={�8e�w�O�V�:V���3�@'ܜ�_8F��~ 8�{!�����$-���z�-:����3�ǘ�Y�^��O'GaP�K?.�������) �i|f�fi�!!�⟋��ڱ�Ŭ�"�
�f������3o-�}�"6�3+��7:����[j5P:�B���!D-�j�\*�
�f���9�&�36���X��xpwY��$���R��_#�,��Z��|o�b�-e�6G&"�_M�uXަ��hx��BE)8ɴ~�6���_AT:�xaU*�y��t�v��D��=^N�r,�R/�dϦ#�m ���
$T�d�B$}��CR���xc?��QؕC�kM~F~CE��r�ݎŢ"YX@���O����v��f��I?$��,Jݥ?�ȌB��j�-6f�*+@�,�h2�9Z�Y$��l��2	K�/�5}6-�[�-��QAKkV-˫��|i�Cy�U�3|��$��7z�\0]����b���AY�o�a8��
i���5?�Oݹ%�+���6.�紲�s�4�y