��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e�i�h�N>��v,�lhZ~��Rc�	�]^%����<��C�'�������M���,�HB
�?T1�7����qڪ��w�N�8��%?��h�џY� }`0|�3��4L�����֦�`a{'��D�{5P�W����#��S���.n�]���u���\$�Qk�F{�z	#K�%�gs�F���Y�Q�
OLƭ���ZӞn��y���&�V�D��t�H�ry*�VCaa�N���d(�DCG�Y}�����!�`-�f1�L.n�D�c:Z���x��hk@ȇ�q���&�/��B1:��������[�ԋ|�f
a�i���-#v1�/����Z ��.��O�k�C����2B�%����S�{�X�1�u$�q�"x���'���,~����u@�8E���vK�x�����U �+��x$�y�|8�B!�M�_�}+Ŧt�ʊ���R�����ݮ�G�|�=�����.p�~�:d6�k_�#�G;U�U����[6=FW�RY�cT����z�� �q��to1��b��(��6�s���;��	�۱�"6�@�>z�r]�v�f7��Mm��F
w���h2��pU��3a�+I�8c���D�[x�F]�]��ءP	�5*�A���dC�3ZF���$�Ғ�e�h�c��{H��(0z�����|���	��˜.J�>0�5>��K�u,�:Kews���:�G���ٱ�����Jv?^t*������O�1��+L�4iG��@>B��3N7`ǣ5|	���l�w�a��X,��VY>�<�6�I�7����Y�Eu��^����9��m�jb�
��D�؎&����n�����h�[�9��G�"�̀7-���J�sVN�