// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:45 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
X7IQIgotEsZ/hlWCjF2b9XdNNrlLtYWfgJZXY5jKXn7Yz8uJqZd8E/666h0Rltx0
CWVeaTYTizqpdZUTzlWh9j4dIBxbhqRzqPBrQy49cZ20pyzID9F1f+nyjWo6JYTY
rnTTREhikGLYzp8yaO7bXYR75p+BcBQyeHHZcp6Itt8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31792)
OWu4Ro6cRkJjoYYIj62pgs21CDJ2kLRcEJv6zQfb7YsJMzoypSuWZa91NiQPklBC
b06WRtxdr30Hb6pDk9zxdVq0NCLZdWOGrNKBn3xDFg1XIACIEeAm1vFZjRc+xMt6
cd02IdMOBsgq+GDXP3MCX+DcNaPfC6fr2XnxOymHWFZ2OHzTHW0TYlg6tCEHqCtd
+eU4U6LbU41tS9pi3YZ7gMDLlSYumqNxPP6zwjfZNWpgfIEDlOIisLZnXTv/CLY1
3fq7cLmxbYiPVQkZiHBVewZHc+dRaI49t8K0RvbnFtADecaC7CwaVBzkMLgi2vkN
LagJyF37NeAdcDpWlXXLE9DhgwaO1xAGtimX7bbFt5dAImKt6xKAc7hdlUt4lhq+
5s+Ndfo8jzWsClzPuIvL/hF9uhQJYTdua7pwLmu9DzxypiuiAWG5S/FWLH8CSYw9
c9R4AZs1oYERqmH4J4TpepxThAQBy5N5qCHqniJBaRNHnls7+zaym3RnDV+GSTX+
HQQpOg54QFrbpeJyE1CZbmsX6IDCLFTjLiCU3S6rl9IKwiImil+d6oWyjCOlxZG1
D4WnVkZ6laDGISreaqXHq1fymDhjT27Ux4jenuRP5o1TQWKo8eSjuzaG5rgr3+UZ
ykLVUb3ziCJPllZvbsUlrMC/ulryJChf2f7M9iQ9SYi555IfMwSYelu8/io90Afj
dpfUdAp5zIJoU+s9cur7inFN1uekutAqfjB/61zKXOttMg/K/NVCHtLOYQheqq/K
j835oSLRzBDjdTfgoL+UHX7Ql80FHAukmsXkXSRkacXAkqHKb/qvH9ENeajQ6wSr
BTcIsfN8wUUFSkbNP6sMndj9JDvtnInFyQLNA9qXID9WxWkKj2OvtXgPrBrS2N9j
MDDVSa6qzkqs8kfQBXIS5zKSsCwDcFDbKe1PTzkG96QW8Xv8GNXhOS+zzgdSuVH6
YlEw2LhEutPjW7qXNjVFkI/BCXU7xYUIHyZzzfqeVlg+DcoJdAP0TFUCV3ibIKvH
o96UPjBt8cPSAHL1bP6SdxJZqdfGxACIMxdgKtB4azQ29N8TH1srYU215xEHFDMr
sxidpkc7n/7w6dcExrujOdQhn39pULZGKk544O6QBzRI+xspnpnJ5Ne/p0NnJM7m
kwL3vIs8l5UDfdQhyHXGkX4/LqhkVdVixlxuf1QVd0Qfl99emP1lgtHwMqTo5Rm7
pEZFhlkGDL2qZg5p8I3phVtN/yBBg9NqhhFzJaQz8K2R/v8Z7x2RC7Owyib43jy1
VBGHEpqjxoIwMODa/mxQSDY6kE8+XZyfZE4tKMqdMR3ylmWl1CPOSvPjjjs5PiRL
enCKDe1/FUqLU8qIl4D1YFmGT/LXAM1reMGh0qCYc642Yn9NNWN0O8MgnQBIwq8y
Q6/ntj8/94Og0zcUXgG3VyD5eQ5uvgPoEcufMn9l7bXytD9VDOB8AKyjo5mq26AM
bold/RtSC/auEV59rkWyozR0QWS7yBCtam1nV+ZOD0nlRoQNYAt/4Hzke9DTMfbS
O2/0dt2WiyJrEKP3tJ21XiEfnM0X/ZiNKD12QM0JEyYDw4ZCpfFwyEsoCG2lvH0W
Em4gYxVNh8S0Uxt3wJBXdRNB0zi5+zDQJE3LmkG6pB7f2OC+bXCVRPdx9q0wz++4
oUSAcQxUfIkcqznnsJmHPW/obUZ8fMm0VG6h8g8Fy2+wa6oEy87weI3lRdAeIjJw
vLDUkIOboGXq+dyju3LfLNQCNu2DXdJ0uNkce6QPAV3Xq3VQ5acma57TFZ84699j
NCp1L5rOSeP2ztD/b7iBMysqdk4JHX+FPhvscpIGVg75AR8TjVaAdXLCHD9esHwK
lHw7PksLGbsrc1GrOK00zUfAla19lypTcpI+IZSbS0xZTDIKFabPxClzxKlLmjfq
raFP6Pz1iXuF7G+azSpaBQrIr5/f256VggzNSNGnhSeCUGRioNQJhz5yypjv5vpl
NhdctJBp064/ytssTAzZQoIWhdnS93pmn+qWbpuNOqYnQwkN/xUQSq67Cuvr2zcy
ZDDlFI+3D/gVZHLK6Xlmqtwo3jxc7rQnk5gLm7tKHcyqWGpbrAQqUO5Gr0J124yU
NLqbaE+IAGAuBTWIQXF/8ipz7wUoeRPpgFIkXxnWn7N4NlAcVFxhefe7ISqLa0zY
D0GPkqcn7nSZi3mIMvVDMJBraeuawnqr/tJVGKiV/wm3KJv75YtR9/llzfwXgzAl
EqXc0sbtKmOstVTXliP817t5xoCA2SVqFTmDTFNK7T+h2SN/rCwSVCMT/g1OVWhA
I/cnC9IIGbfWZSXMmRxaXQPm9AbkCCtdEpLpz4g/IVPSLXowUyblNsAIz0yNDvZJ
UYhKWI10RqwTfGEUVosLzoMBP4R+zWWyt77S8LBOi9L9OoSmK/lLxnmjbiLfJxHA
Gy+kYS89wtNpyn2xQzP3F8+mwg7pIJkTaZNyugzmW1J9GoDLPv7ZRpsTwZwDWdtX
3wyco23SNCo2j/ymenUWdp/lVTkU9W+xkYYS1bmO2EoHHTNoQPhtDXImau5OCODL
B/rVyKRGd9eC7TgZioaw5PjeXllzlcFhBnINSQ4KjZRtr9y21DyKTOWbYz+xa9LO
Q7Cabq97NxR4FxaLe8DHAvdDHtef5ItPkyk9lz4ftFqA2Y6l6iLBe6knEzHl6Q96
YUy9GwY8I/jHHtSJrXMDs8CS1koI6KUZU7W3aSsSO7YtOxfcjgyUkpgFO9HFvFVP
zLSC78t1TkdYyp5rp8Ht9cc0PJMO7H1FBM9lf7Mo4wN0is7dydqMaZLX9P/4exn4
MsnsnsPNI5ALx0wYNiBB3VF7QDj1cbC7rY92xL08r+/GI5E1nRDTcXjH4h+fGOYh
3Whyv/Cfcg1ZRd8XtCNbaTytVTV65I3t8ede5e/cBShLsfLFz0I3n7pBHPxIWqwt
N/rn1CigsGuL54Y4oDJHo1pCMDSg8cepT5j0a+3xt4+et3PCNSawn0ocFSfajjAP
Oqx3SxpdtWIgdewUsd8yissqlrwL9JxroIyPSrS1JaPKL9XkQqIaNDhGjIYlrjI9
GCE+28Smmcs9wgAh4vcCYeTQiDx7yFFMfEbBMab3dpbvik+RYHrgxdwzIVvyF20S
O6RJh9m8JQVPeCujw+kMPnMeEqr4DThgGgKcudWHSKPUhw4+sTzOR96prmnr/7Uy
d1qruXYP3BQBeO/MqE8rpVjlaEmJv3EtPz1hWQjPTZB+GQYXH+XYlrZ45V9sJsDd
z+9Dt6rcLgyklHd8BYR2FzIgFN5wYhAP5E/fgHt6tdIvNuZvwGKY7G2IKpDidATf
u7HxKzHAN0AFgP4NwhgiSAKXwruV6XAh+sXk4FxCgyN/s2uQUv6Bnd+WUkF5qQYc
MOqjaJXzQDFKmGSVOCGTemzvJQvjNv9Znva1taOkbs9ZDBqJ8XH+d4J0kSjpg7wQ
5ofGExAYIeT2dOwjw5tKePfgO0aFrzroTLTlu3YcLr/zI8/LvFDj65iXwcqWzpmL
i8KMbzB2K+/v2/imD1OEgw2Yp9vPaF74ZwUP9MJnDw2A4AIxe7n7IfJl8h9m9uRL
bRbZ5EVIOSW85+YUDBPotICSW8sDSSF4IkfBurcXNlbZpBB7ANhDfRA61RhhfpGm
NlFXeiEoUKKAgzQCs/cgRCyPkJEVXB2qgO9WWSMB3Kg/ECGKBO63OjjriR87vwvp
GIHL04yZT0KWiKhWoLqltAHq9n9kZ9YacPPvU4mVih/uk3nQhzz31tAhrigKjWTl
+xijEI7QfhdIbcTsXjj0+CIdUgy5Nb6wKVBs1oaTvfSzOWgETZGQDM/AWl4rj484
upeKBr0m88uTozjcXZpObDJLL4IXSbLJzRBl4S8lweriZ3Hh11Dp9mfs9pmA5MaU
2RM8n5RhWokpjqDRG1DdHIyd2y71qiZtIj0x3w6O6Kj1KirixZxN9Qb5+C9R4hWW
VQURRGuDGsQVMfeN4czzUvd45Yzj8PoeRrJ3YZ1bELLRhJYIo5oSJWdIMA4p5U3o
5iXoZi30bm5L303TbT97qZTNasW2BtTw/nto1H8qf9N8fOcVGJNjZBJEgr3cKazc
xbHIv8QgNIerFVHkFa+dt6M951V4BKvtDubtwviwcIteAiyo7FaDaaImoobkbzLJ
oZInULoFfbFcwdkOQBJhFJITR/AGorA0joW7rRZBg7721yzW4PwBjjnStbTDmsOZ
m0KRDqQrWU4/4g89wiJMhnN4r5eA6Rd4Vyr2UYLz0raAeTH9QJGX0ghxFuOOZtsv
jBYLWo+n34hcs87HuDzW3mJqdF4PZVYgTkEDRNYYcodH+94cU/gfcH4NdAymX1uI
5WwlFu4aXQgLxwo/iSxbZeR3eSsQvOOcnPV6nyLYliC6c4H3ItsbVXObMJPgvK6x
bdJAs/GyFOWMaq4fEimqWEj04dLKuXPJYvR0PweO46/bk5ElSUcx1cXTxum5zrO7
2+gOLz7orKkjhnx6W2IREEUK0FXDgzro9JB3g0fiPyNEAQ936ou8vR0o31TUoBuK
0/Iiidih0PIhBYEo7ZLE1/eCJdZvgc0h2Nv76bA4ierf4E2iOOSdsSXSbJZdgC50
7akRXW/Nr18DSCFgsxYORjWNQhx4i4RDWeJFyalKcDhK3DAzoLSIpd9UEBJzp5Yg
mMeDDDM0CMnn+bRdEGX/r0AuIXHjv51zlZKzjdNkhWDKhOeeg87B/jriw+MZo6LP
XvYYdBCs93GfqGw+kts+f7xYn+CWPBYx8f68LR3/DROT3zcZjM6HkAhp5kz7yvLi
JSdapFjhJ6Oi5erwsd2gNicco+/l78FuZ1lZxUJor6pGY5AyDdvLCsrtTzQwydvG
2vnmL2foJnCcx6eMbPW4FTYAasMNAzYMWsy8SYZYtSiGiEzpHiUYOmERQOlyObZl
LsPEM83VRNDQbJfQJGxwh1qYe9MrztBKjXuh/+nm8WjQBmCy0fCBU2vo2M5jJ8sB
TbdR2puwHAX6My9cBNrUJvvc8MAWiP/qIeNPTsljJDbsZNrWOzFvMke3ke1+rPPf
2PhE/Y2bdk74E2W2iDaOh7bHzs7M/+dOpOtZ2L9BghfXgr/ZEEReEmQ12XCOTQSE
0toYe/3L7HbvSdzUci6ItCJsk0VANKjQVH3XL0BcefyVPWNK+ePXM4rFhFUZjbVt
Gr5zsvEVhVdFF2UxzDH39uuuEUDY6PPIwQEDGAdOrhg+miTNOSzuBFgi/w+u7ebP
gC2Z8ZpCPE9IS6+dhxXQwXMUVgMcUs+Q0XEbZ/OkrOBv/VQiLIj6wUIUE7wWZqIf
7rZNtlOPRKPORJaiuvtJvyyjM+1SXxp9FbXCHD8+o/s3TB4HHdjBap1GMc1a/NsP
NJbLkyBEwodfOHrjmYclNXbIL1aZIOe/zKUtojxi5+9W7BxNFWcG/NM8JVEs2ch8
vTsHccDXu1jyOR6e4zGEwRizWt/PywqAochki+9sgSVYU+ObLb3zkKQe3V7IgXJR
8YienPVIaqYcsPQEKm+ksKpbmqp92E/yJ7fFdsQhx8qpLMAZIB4ihoVZ/njEypLW
hFD675ZGW3sXMu3ONgHcXCTDBnyiOeGrZhUADSk6cANGpaoSm+wYt9LqQFtu7W9S
vXUBArQx2quH3bvfGrq9NpcfUGTa6S1pB3sF+ksbOoeRNe9BYV/UnZh8UGwQXExg
ZOE9Hh88arAlCnPoT5kbczMc+5SnqaWOgnIkk4JAD4RpK8eq4Me6XbrUGqaidw+k
M+jOz/B/7q6ByTeb29feiKDRnu+CEitE1BzXmOWDPL9xwiANf92RqmLcpJ+EboMd
PpuVeSXTBZEaKDqtVe1Uox49BqUU4k6Wqgy0FmFRiEuqD4+9B8ZGSLQ/+hPzLos/
PvTsERpIHGfHjvTfBXo5/iAanlx+CJJZ3jBvy0SQ1bSub7/yJ71nUIEvWXqVr5fo
bazmJpFti9iFIDpoHUsXBlewQtPWln6gmGvV9NsJjSk6naenvmMHS34z+Aj+ZY/M
NuEaa7oqZjSjj7jvMuzpGSVrGRLnuHKQol6LB5S5aw8i0GasSCYwecl+Zjhai3I8
EV0I58YLsKxr30/W2O1btoAmRjIW8K3OmF//GgRsvajY7xAhDX6RMpo2GbHgfB2K
MjpbVb7wh4HiVJkKbUrKGubCy5CFbkJRxE4lTaaGzlBxFBTWdBaa5uGxJ7jaPAi0
Se8+AAjI105ebA0aVYpuBL+4HyxIady66a0vyVf6xXXa0cX+jldoBSAFdd3JZv4G
WeJwX8ucVcqhBRLfpTnh5mFK4x4h4WXDcpV+tqbzOcLLpex61WHGtTegz9LHhOri
t7Lsf4Ss4NpOUX73q+zmjLjbJSQiPSqqntYXRuyodtpswiGcLVSq9abBvmMg40wa
O7Hwm2WAdIDjZ5hATmPMxUCXaS8jEF4nZt4boM7hkjpWg2gcMhpBpSB3jKLMF2eZ
NkHl2weFx6bI9c5BknwaaOriGvLiP4T49pOb3JlIhj2LqeZ20K+8Nn+ErvIYNDMD
5dLaW3Er4efWifsgq7zLk8ROXIgHh1NbX0e+S1eI1TRc9zjsuUNzt6BPUsgT5uSe
O0DHYp8/LCXWFTMCRQLEb7ES0fYupencBFupqpXJMq+b00D7FRNZF3auybsRpBCW
KFUoSTOtPMkxXJ2Y6leg+rD2R+cmjFXFdnEADrdKqgPijedXSQJNKAbdNf6Lk36M
dV9oVAKyFD46Kw95Ep9mWuvcIc0xRPnBjg27j0IauzFnWVc4u1u6AO+yjVJAAZrs
SozZF95E7AGkD17oYHJ1PAMpger2jMGWI0iF84kRuHDilkDd8tmid3pYumohSnVO
uaAIjy8fsVX3hgorN5nJSNS2J4BnDpZ9Z4Sy5wZMi98FXrRqrycnt/C2IapqWSJX
JdQ9PxNkv8qYH3Ec3NeUj18Wr1u4xlv95kU9PHIbxOe+zYwBPkkzcmAUGtv8QUHv
RsyqQn/jsSLo+ch7+R9tHynF4FVARHyoT3jraFdMC/05+6xo59hyRF4KdkSJPubc
ZiA5OHtzaVKLCg2/fK3VCzLyQ0wsMbH3+i5IekLvtGKv6SY2lN/qNnZiMU7Uosj9
MroetZD4Sihmp8DEhUXWNk4CNojUTRRROSjmUM3SFXiwWFkG8xC2FdIXbpTNWN2B
/4oZYyIRhA4sSwBS9rnUe9nfEVB7WYJ+lKrVZ0Z8vSVoGnrydTvYX6OozAQ4dJxj
kIZEnJw7+/+Ws2eST5qpLLIwXUuhwyr4eVyYh3gXid7fjl6HqAzNdEu0Sg2aJuUE
pU8GzqQu2eGUW9ZPeZOncSVp579+hvszWwBD04tprGLsrR4KrabmcCi3elU3n3KC
d8dUgQMDSvnSn6achDip2EZW8XzTp7YHMN/3IUU4l+KFH40XbXYXshi8GWPBp0QB
4ARugfpv/odcFHIR76viKEJ/jP7kvTNHkB9ycRmgeZnZ6pZosE6//6mN7SZiuPlI
21VnmijRC3t5iKgDHqqCjuvW90+vQKtxtixrsMD8sZnOqtbf13JSO9Z6BKXRMJ48
EmUIBtPoPmShGRu1cRx8Q7eyR1nuWngVToUn1mY8zxgGRp5/ualoqSZLE2Zlcq2G
cuAHK4cjLVgPTLupuBjuSY+22cTz2WZqWLzyUYq5aDR44UvrPLvY44XJSe0ovhfu
E+JAfmOu1QjQI0Mj86GTfkxsqpi0bLQjt5BgaYuYGV6tguTtdKW5Kga6z2OlFqI+
SBxKs9j7WT/Ahu4CFlt8B8s1xeYDi2x1qBShwJQM0qNBj74aRpjPTT3BcK+b8KPN
LBkPl0O86BsP3OOwWDRjk1tI1wGNDj7ZPlnGSSsnhfbouk6LZhMj0KCTFHVNyo+H
okDz9qHD2PBLOJPzNvtA2SmoOX+xyEG3mfKdvTL4+3mrhtyrXjUcz7M3J8v8ES5f
iElyLLkip/0N33v5HDzDtoNQ4VFQFzazBe/Pp7NRsgugYBOhYIdKKLtxH7OQLALG
NgULQh4U+ZSqaczxAeJwqGagsaq9+tISo9NlM0SCylcWO6JF2nJP+2ygSnRTK4ke
gleK+xNgr3h6ZyLwibSSqvdrMIxioSyRE1KjIaDE+YRvQZrDQ+/gaGHh7VdnlFMj
AsjYuggAFasZIFcMqYq7rNOtA2/nKTvY46zU8pZi+nFu/YuRf1XnwBCsbL4kUcUP
399EXedJROMeZ0JIJPrTzrNFEEAi2sVrOWolTHjk7QYl5rcvSzkO6JruarV2F/xI
DH4cRfTV3AbrAfqY83CdvhLwWOYL/K8xzWPlrUB1LF0YySPwe2AU0NagNT3L3jj5
QXfOf5El3wuJC8TDQ+wBqbGAeltTLh8t3HrfLPkAWFlMj8mcDQ0qc4zQvwro2GUa
EJcxnJ+OFdMP7nIbFrYCpsjXLZNR+T7l5+2y5KEoIj6mI9Z1KqF4W8frbLFT/4Dp
kcrzP75Taj5lggS2jzZjLyzWfnwzGIBrqWqOevATxtMso4xxgVsY4LtXhopTEjpV
moAv4MAK63DJIfY9OykcL4JZroMEITRxvc+EN5vTK4MypFi+azHDE0rT+YTuiLP0
spk8qrwGA4BLevgCDw9pGcj7yBcW2vG70UzT8TWFgC27+yIX7r8TpuYcrWosxCoW
D5wHBDExWpc0txRdp4LKF9sCisiCl11vcl/jNGTk0v6qQH7B28OIHdBCKKoyx88D
q167srGbPqglibgV+SbI0PIxWmarpuRc2DZiikzfOmJUoYUQV2FblTkzO/KfLe2P
ofB0T9MVSYmTPcibuMkAqAOOl3Qi9S7k71RrF8SKwq0mnc8jfXpymbkpC0D08veq
uAiGfpNmgRznwjKMkE2jB7xvmekHA1BhL983eY65Lj2RlIUFgbdxyE7YiOEnIpVO
wpgrGDVHSrngaCz4eVBplbjbXKRdFhF5Ttz2RWth52KuMwQd0ea86Rgtw29K+UIF
EwsC9NB6Q7CsWI6KC6MaWSL7KpSA2U0y8JpdiHLfMlByfPJ/BxF4afheAIxVdzf0
ikaRpRF1fY4ezlKETi2PNHvc6kyuHDjRMvO6Y963T5TCPuEg+02EEnzuVTm8LvOZ
ANswGYRcBj3u+11knWV2TyEb5cnPt0d6bdfcLe3IJjuwcWOXKyDrydfgkL5P2cT6
G1sqYbYMXP6SOCjSJ8pRSbwCQQTE6JBCgCjsp6eSwFfrPRqX6vA3nQYdFBTSl64j
Q74yeEoEh2DDe658q2t6E0WmVF8b0bW8ge4Uvhj8L05yaxhBfAi7tun3VWo0UDJh
i8Vupn+T+Tt1L2vcO1KGyYzCtodGzU1YVOoNKuttKv0KwprqoC+5UBxdqYPzUfH8
PUmbqkj+NJSp9RFrRTp2HtOTb8nkzHpjb6ggoNT3DOP4iYR05G/johG3eipF2zEe
Q4xJq+znDiUUEbqfaHQibijYm+jBFXd8FBt1vuHBLto2kzbyxFRCiXw9UMNprRny
1L//A5dLWZuzftHOsuWM8Odb1qV5HG+jTFiGgCW+EB+ABESBttwXDJ7y5FqVQewk
7zitnETkOLTjII9jXzBSe38KdGN0k0Rn9X91Ss+jasZMXgyihK0XBdLlXOBTSpb5
dptcg1kVcTxqFHGxrjYa4NSV2o3kzvYKRCEJjJDUDUgdytfMp9Ocdt86qicJkNbr
aDsKw/+XaLdUbJ22xDBeOIDIvIi/eZSa4HSnU3d49q6m2n7uzP/8KswhTDw3lTB4
r+o4rOi3T2cCnLOVPwdF+APhRxCb5nFlJ/qhe1GnxDszQziIlTajs4QBq/mQxcJt
ONh24kLrOXkaCoC+farVBhYGfUrUsii8PI9ruVXXq8rRCj6UWq/o1/6kkDRxBa/C
xPJX0oGdoG+j79IUVA0nVkJCE+kWrKzUF9RSNcp2sdDO1YdnndJtcazJsIdppqyA
gjslP5Zh+UwHsVXP0uZHIQb9lppcucB/aRC/4P+dMIsDHyKfXQDO5LKo7WnP3D1c
hearAJSHAEopPkcutE5qJqVBLzwfM9PitrE9vikBKP1+KyxTiMtbI4tgVdmYGwzY
Y8VxnKJnKSFcb0iecSXz2nwwhBOlmPcrw1e57s986KCEpqK+hcS+zFQunODAilyz
NjV++qTPyglLC+w3pmSLDzEmG8tgrKeMMqFyzB0e6AnvT6dohM/fkjwdqI/d3vg5
+nWisQWpZNtOzlyaOoqpGSnP0Vvk5ItR2G9D1FvLi66KFgbPjo0ZZUi7RJpMSYJF
D/LgHyPRI36AvWw0cQC4iWc0pRejHm8FatUH5OwLTmExfS8dsj37B4SiW6tSkwVg
RTtcWOjoirM0hnA3qD0gyXDKytH7qhmsFwEISfJGmNUJtm/wQY82xcsa4HHw0ftD
kB5xplge/ArYuV9EdNWfLxZ/qot9ESNIT4geT4d8f8g0fjklP3Z0GVGW5k6n29ff
fBEiq/QVxGHzuQLtb93/Ec7WQ/giqDXdj9AvaSa3UnDSRzVvNTpb2hZ9blKvY1GN
4xSzB0xajg6FCHqhtNK15x+B1HeEjuAJ0L0ojCfG2kHkXeiQreRmuLh1jJOim0iz
99u3wSlf95Okxkr8sB8rgA0hAO/LE/WRTT2nMN/zO2APMlQB/gHb7wMsWK9AJUhp
luQeH7TNN0R7TAd9DLmzOYdkp9Xolus/qtBs+26boad4XQAl7MKHgpWIZTu+fJQz
9Mx4mEu+kYUHMAjEgludLDhN8Qykx7gbjvhAzoRo0q7KUoDUOGKYjVQxaoMnn97a
NQ2Coi5I1C/rgjL7UWOaB2IiM+d/d8h2zXyHaq/gb8wTLgh+bcnPlpueuSmQWs4e
Tse4SxiBJfHfNw0+jL2TShuHYBisGdNAUvIr9n8ErEwMhUvY1nNd09p6L8Wo60Bp
gUDO+gp4aYravb7j2YKLuehe1Ew3gOgrFhEXWbAoFt4FXMCgikjRcZpG1+jZV4e6
9Fofm5Fijz/eHjENuPuT56yBUp6rTN8YRL06UmozHarCgW+kW6xJbImhCFnXIozC
cqpCwNVLqyRQ+cUmDuzNFfYJkQYXSf4UtJBDp7YL+GEneerkrzkBmwTkDE8AbRv+
sdbk9eYskrO3XKKM6IAB071p24KBnGAF4Snol4gAKGYVW/l7P8gehkotyI7laq+E
/vkqQMZxG80HCR99pVLX0HVMZcXg9uphRz39H/4H8Bc6aq3bMwJBS/pBPK+C6lf0
wrVmNfa89P48NlGyw47SkSq5/y2PIRH+rrBbV+4cKrk2l7oyr/kGXCQkZQq2jWRG
dQQ02jc4twSKsqnpaCzXTfl5LQgpKZbzcyxUfNVjL3ZiBXQl31yHY85yg8mTaytC
FfjtQRbI7bbauTDUYc0TdXTjffX7G67tw8IAAEg9btUF/a4b7U3ywnf7couzM1lg
R1qcACqu81fY+t1EpD63f1WEN8b37FGsWRAuXdJQugEyEbSIaXu9GT1qcO3cAf9M
KWysl/0duYHMMFCnSCBSiPJrneRczDjZgPlLEjHzFuAlNfSwzeDJLh9m/KbRfso6
7F08arFSKaSzb+/5qpQM7drG6Hb1uOs5zJ2SsHjaUBWpN6dwc58S+XoegBCbcl4+
eGl3n2eKescTBvSrXJeoUku75sVFl/7WCm/rgkkkNtqw1lyzd/wU2dqXSzG1WIvy
uALZHQqOUJ0+3L/l1qoqo6hV2cM0hIPkdfW+3fdj3US2KNaG7K4apW2CV+UWdTI3
VGGimvunZsdSFhxwAiaz7jtq29rcr32P9Hl8sXj2CZo0u5c9Rn31fFCda2WE8Cvf
G9hud66H6Rsv+ZZF1dnikIs8eJVw/iMHxf+d66SSwdg883x/2zny4SVEGl62scN1
v0bFLdLjs1XE81ohkvWgqzFPTXRKvXo+1fu2LiaYxv4GDErZ2M7YOniAXEbngeDS
aculOnLC1SIK2qHKAsR25oDoXbw8pJIFvpu80TF3Fc6xTp2xbv6onO0OTPJtSBYy
9WlVzJVELBX2QPguQIHPbHDiBl/XX1fZcOQaHqovJIGcgZKB+X3/FffAmFLQGxYv
h0DzQUgnRBuRnOhk0ht0brvI+Jsn9NfC9wkPGhB/e9YocrvHsNc/yx7/mKLA3uZG
ox/VOjKLulGgiAU1WSbjOzBYJyCIDqOWoCAOPud1IrDXlaFoqH7Ryq1mHYppUEYg
gf6oQZsDDvV52pFAVES/puQ02vu4c58r7ixNT1QdiY3LnHQCy+5m3UUwBAVEzCZU
05skE0xhFUr0OA4nC9q3bHLH1CENCBEl1wJmcYyvdvwKMvxA62wD1OEN+8XwaO0B
jQrYnEi2HunhXjMmbo7tTtq8TfTYZGYmbC4NKrroXG4jlErJod9Y7Z3uLG+F0//r
tE6s3kihJBf5zjoExmGPqRb30ZWGIDYEnmZbZ6A7WypnFYkHSLWPSk7KvcY91jNZ
QDOWllZ5zHNXUB8cdFd+d1YqbVG0u92E+RICN4fVq9garMIW/52UA5X66HXu/6gx
ujWnTgN6pRtUoff4JMBRp53aJ6aCWfqizjOwSdDGpLWgTsXxmBuQekXhcIsk8+qk
4KwROVdkX/PsAN8b2pRgTpF6ygO/u4neOBsGfMRH5moG2iR+PIVPwkCTrbf+D3zb
CZPSCaBgRET911Jx/ues4rEiCkM0a41gozE3qhxxNQtV7cDR3lnQo0VunUU6DTx6
T2hzhefmNcWZimzpq0l+OmVnQjVGEp9L1u82UZVLHNxSyN8Pr6dN1jVfk1bTI2qa
0bVv9z18bKaQ8SaZixP97OkYUbk0QeSnHpSn2Hrh76e/WCxShJd1Uf5cLMa+sjUL
jquUUAMKg15SARLQ9AKTKOCXRPIoj0U0+QqABiQdGHV7YyyrlI1EE/n+yAB98IfC
re/IA2KbQRyb6aRqDwY8VIRI6EnLmUR2CmC+jMzxFWwxbbnbepige2UoFa0Uocq8
1qEdFTTGVJtPA/Lrf3JMxnP7e71HR0g1K7kbxCZ0mme5o9faOEuXeep1pRhdr4iM
NCozDY22KqxmRN+mWRz6HtTQTs2SN5JiLH9bNP+t4I6gUjAErKUTOmdf87dYVNbr
sToPZmlhoEqp8rNZH1wfNHvE3dd3G4xLpj67kpsCaIRAtBoZGUIUNSXCl8T8MP4r
MTw+mSQYSzzeJLp2qS9BvuHkSCcVbBdSsFxOdpUpRSaU03CEKCLAikdKX16yWuA2
sJd3LLmck3WbQhUKuBs6BFN4f3plLFGP9UrSg6ja+4q+XpFnX7IwudkGQlSNGDYx
MUQm8hPM6cfHHaaV4i1CAEjwXx63JpIuJqg3ctQD1YvsZ6P85e3hSIqfxP4M4Maj
EPPl9I72IIgV+D7v5sB21rm9GU6jqD9cg00kSRSwTT9xLbL22AZCny8+CLygBwf4
qdjaLRi+tcTNQENtNyLAtDfZtvn5l3/QOI9WtZGQTgJOvbsRP4FcxYGWMHY+HQcU
gybz2EyeDi4Ke0etjT33z0XOcEeP6vWCBjIRw5K5CbtHgQ3BE7n3lT6db2SwnUmY
FEA8PQMmjXm9M5vii64+eT5kh3TlG/kdO0pF+RjkQ/onQ3+M6jxbM4ngpU4Q/wDy
siZJ/fuydiqPKbPe8qdYehPFbOLBCRjd6fvsCzyuTprzqSMV5ACRyf1GwEqiBuF2
JwiWdeNQfqzGgCn7giG241hRoIv+8xUOAAwd05nPtrio/uj+8MGip7YMuf58g8/H
19PE2sgOHHC5tJcCxMJV02WzbCt5D7l3HigSfJzrMiaTT1rCtCCrS46wsXBUSJU+
tky1NqP9GF0hJF7YZCHW5is7/UFC9qGhkIOP4ruKtzyl812rgqHqyb+KK2Hu7rBx
ignvugNTyy3pvbFwl9rzRCPiN90+We/IyULVTbtWyxNSiPe1WzBG/+Qq/+NTStpW
4EK0Az8Ro36p62FkvOZRViFfRlBzbgKWA5/wA6SC9z0G1dlitD3XnaYbfsdha9go
neHnNHaGTkOLLdKfSVvzXYx7hO+DkKrSyJvCt5ALlvZoHblOx/2nkEtf18C3xd1p
ntc4va162VENthepUrD6vFibW2/LjU0vUu4UmTOSPXvsu4XEZmUiMwMmAJ2zEHbm
b2nixDvUai6X3/V893IxigbdHgoYGx9E3t19tPk0fUq67rNM/NsrxL5tiuagvIwa
Hm1MhdrpqF7kI7WRPktTqx1Ncmp4LZMCulzaY07gamzm5TjY3XpaP9eQeO4C32CT
CmRBuSb7ndJqaBBclTHbAWRBeTjEP7N3fa7aLyUlmXQuBjn7Uo2ahdXnQYd2iDyT
AklBNZyk2BvJZcEsNE6bJT7Jfon00eDUS26xxYrkcCR/58mdWFpeobdvfzDFBBv7
crGAH31TEG0+ouv7W8rR6kwUuYMxwx8WfdmXnq3/bcK/tlrAH2+W5hpNEpk1rE3X
Fk5uvg7flptgc3xmeM2/rNua6aEhZ8JCV3zsIcoA9HIDSAW0zOPhPCvJC02ISWmr
MTtnDb5mE8KzUVnYX03/USxaodmV4ysYCrNeCKFV0r62OxolW0TbZfKujUOeKkz7
QRQxn70kDWSy9HOyFVPDXKzHhJZfs7NjhhzMe1Tvqabymjfv3qdiuejCkJdnNbJS
qqVTrKk4glFOLpNlvDuZjzvxwAovpnESqaaoveCY49RL0h74Z7CWbBuz91kn4Y/W
GKodcfxS8UCwj/TO65HjkOvGjebHrGsGJbq4N0HjiccmHCj7MiNs/vYE+4znPwNs
hvLgRwIYp+xbw61MNsoz0yn2LuFYOBXDBywiO7vyeJ72u74c+b7r5PohcVc3TdLC
V6kcRzDPv/iXE5muaJal4P/EBj+XQOLzNc2ayE610AHzLUu/frpBo6CcuKJvCEqS
663FsZhfPZmn2oE2sc9q3QaaJuOjN+BrFFHIE/H4hCb7PnwKzhs1p/RJC6wKUWv8
scBmvHjkqAZeitE1Obo9D8PBjAZl5c9OXsxaFQBZ8AN5BOcoxng0kKO7OUKexEw/
yJaYcsiJK/rJIQFWwp/HM73WDXbKy+EnQDIqHJWMuE9ahHDg1JsVU+etIZQmQO3R
phn67bMTGg2AFtwwGoZWNj6J22qIGJNXvK60612d6Q/5abta+vZptD7xNflXKZkv
B9+5+ktugYDxcQR5oHMke7MQ+qhZ/Ss3/Ieoit//4I6YLR0ykVOK9YacoVc9ZGXc
aiprSvbe67Wo7l7CTX0Ewtel2yj0ELD8WsuiIlhu/erh07GMP7srtedQzqTuiuGS
LoDtehwhk6x8obSOd6tvj3hQOoeT0JfPIVaQiJbnCAwI9MuZNTMpJORlFRVxkD59
dmprL+G30uKSYGNBCu/yTp+94iZ2Bt0VcxfjRB/hTUERibZaT0O9eaBlkKUijS9Q
n1F4pUbJiysH9XBOSEI7vJXAi5l87oWUSpMFhYs42nyIcuN22epuXqK3LbAlYaNQ
Ra7TCi1KAZe/sQRWpZB1D0MZB1FYqPR5LV19SeNZNMZiw4hN5vIdSY1o5GEf75iz
ZlXKTBh8xTl8lGBqE4unT1be+vOTYeayiHkI7Ex3nEcpTOz3bB18ckHX6axdaGYn
jj9wKLfRaUOvQghEwBuEjE9MnLS2yOC14cgtuxry2TH6rOdRm1aE4CITc8EcbiY3
TI2tAoG//qcSA8Ag4k721sh7WH6188hNAtWmoiSFa38rUQxJcfYZZyLf2QhgCBs0
D4JKZCslZOtHtFZ+OVMYs8niReNI8zXP7EL5P7WLTm4E12+C2CYbS0gzEhT70LSd
RoL/oSwB6srb7YaAOMMy1CXN+Zmszb475m0oqz+O2jsbbCL4e014hg+ztt+224d+
AsuoaUqC98Gtf8SfqAZ8MwgIA8pS481yFFmgH+LnnsdujYBhdgPi5lJYOIS4ZkZm
Z9RolPCdJPfz7B/hzLSbNsJeiVQBpUVk9rkbqX40SfhSNt91kzq1+g+4xNqdi4em
BrKZ618lMSv1X/TZfkpFtYfXN6RyHR+cU/ZDimv+AcvKzSdUemZUvOnkSJLZ42TM
t65nxpPhpDz1dNY7UaJ1RXL9HCCE9fFrLJ6U1aTxuuafzFfLozXT6kM1xD2fEtJo
zgR/5E/arYJrDk2AmlloWLX2WmxIYZZEhWGq72prMKoUiGFHuiiGen+GwyJtMA5U
UEdFlhLr5/gHx4UBAu3UFIvay3bOtGLxWGF7uH8ffB+L0TsjH/h+LO0O0dW5F9HP
KA1UvM5VxnXVeyD19GhKwPIFNwksNKvDAYCpAp5+lXqz6AzOWwznaBgAbfbi0MUj
6SIjsUardCWSumXG0pu4deDpfNjlWO2kkmeKt95yAOZwRVfHhNCTvpK2ZIEg19k0
5WYIiC4lAHVM6tjDyhhTZXkG61ARIHU+U2qQmvbLeeAJfpb/CaNAvJr7BeeBl+31
f7QYC3aPOUGrgyRNYBhy999/YNDFcbRCXn7tdxIp17iPKb2IgQVSTP8AHxlBUVMH
9unZe74GpLCjUbOCNlHjmQ2YtCWUX8+Yct2vsTmB4yNKb7QC9TI+EPkgVD7iWT+f
AvICklmA2tcAKOswdanCkldPUiAq4B/wD5edCaKfNhRMDSfNZmf8RrVY1BMOi6xY
6IfG6EsXi94U7s/1vwiamclIgBef5xyRXOCqh/F3PxdWL0rYoeEle0rPJyLXvRu+
IV8bVL0qjm87/FqJGlnErjgEymavkx3YtHMe6flPrw847lV8Stxad1122PBnk+tq
/v7Mq/YHWnDaW4QAKdPsZrrI/fi8beWvjsHRoTipIWTZlIYf8jCHLWtwVFpg60ml
pKDnNhjkQgHvZcYm4WXlangEiERdhJO8wc27KMXfXGc9LBLjghndToAETM/lntI8
SfFPx6id+l3w4dSZ62tO4y3fFKVNILeXPqiqNnMYQ0ppRtytyynFUAvDJylDnnTd
0XEPBdm6z7xSmafqaw6c3r7qJ+KkvtM0smv0HDoOIatZII2duUJfx1zW0ph4wD5L
R4fom/N81pP4qJcmV3ckY4r+YI1JSBYgrV8Q/iAbshmS73vktPA3qqIFt8SZwIis
Hzk7+rvEXXcL8Oep1mr5gaccgJjmvGp3vPdozLm1m803BkSyFp/4kaKuydW+TdBV
rN7AErXqXVukK8Q62TGoJYCeEWNGAahgAfoCBDY2Egyn5DFzIbtEbwV7YsZFhRQE
hQIZRDUZApXK1audnP0nfVDkzwfs5nf+dfQ7+nNPupbM4NdOdDAFawLTn0AcaV6n
AbWtonde5pht+wc24A/lw2Zyb6fYow+/lLK7HCp6S7k2gVMXZjFabovtZcbDPWiq
rwJJEtlszd6pLae2iMGQ1SryWtuZEpv0+bIB//g2E4yUDqNhsuP8cW4edxUM86yC
GJpJFA6WwtX/sJrejcUShSEjGquHBZMO00OTggj+cngnYtIfYGcfMWCL0OsJJFaC
VKxmelHRjn/jpY+dahesSkFNEjbAxkuutFoohgL1GBr8GAGgykp2fOLer0YD/gOl
jx179hjdzTKyTL8a0vpYsowaAIsEDYjI4y1xrUIGAFXqXnHQR5tREkArA8Zqmyn3
+zJjKHCa8hbkOwbIk4YQBfGEAWoCzOqrhRoXEYoBQHRqrWszR68rdcGcB1Tyw2mT
6mynvFlzLc8fNu3M3WZfKKs3pnkkbQ6XpI7Kdd6ickG3cpsLDvSsOPfj7Guk5F4i
iNa7v/HKymnkH+vGs211LqzpXiwie8KCEWQdBm8ZysNTeQ/fxDZ/LWQ29kleaphp
6uihK5EDIzDwlHEk5vFwdSbR/1Q4x9Kkgm6wR6rb3pIcThHZ5s+v4TAk6VL5kjS5
/SCDH2+hY7+pPAoH1q7jNDCT2+ZFo653hiY+uF8p37Kx8myIk5KQjZ69Cs4xZmn/
eGay6fIGa9lgsJDjZu8q3NyC3fYaF4kWgUsACuVXgZhopTnDMz0aS7cZg8F+9Gue
TINfXQkJBr3mG9fkqqL2iWqb6T8BorGz+gKRKw5iqiVQRGTGCohQpwBkws845xP1
kDKHqKfCU3SLvLBrGY1yWXGU40SH3nbhXRuEMQz0w3J2ew5ttww5E+Q5b28ImOT/
HAs0icpBYs6hqBOETo/Bf43/A4M5Gh/EwWf5mJ7jCm2meP3SUxQqF8KFlvqY+tuv
/8FGf3T/owF6JZwksxrX8dq46WkePXloqPlQBFBWBD5iwBJ3Dr58vapnLM+KQanA
52xX6yR2JQVdAKNYyLN175tGBcuEiMVNDzz3TCuZxbRbB95EqRoV+LTucLHye+Tc
0SE1YDr5dATNrTn7+PJrQ3YBOdwTwgnAUT2qT/x4tqMhHX/g4AH+vG/BiIE51Nm2
jTmlc25Vjy/SI1F2GaMq/qcWGDYZWqkaYKKcbrIUbxJUJHMJucJihirCTIUM1p3x
BOgp3s/EOzPPRVF3XLwH9S0nm2d4rM6Mr1p2mbvXYlZzllCCO23lEpqUkZI8YfAg
uZ89EDK5C+DtioopB5G6VfEI+R9nTtL7LUiYLWeez2YFxVYJ/O+6trxOMo57+xWA
TsZvKyFzooI1hwTdbOyssZS0Y/j8NyX48pO2cBpDmLyqjwwaWpYbb9/znC2mUXqS
WwB0LtNpbokJ7S47Ca8bux3CRURxFxfM9frT11NsaZo30zvRUt/tYtZ/o5vV5rM5
on+3aQIaj+baCwlXqJT06eDBe0hyM5mv3sDsBwM0bukJPD48rEOZZtw554BPYnTS
P8SOBi991N1Y8/uDzcCMBHwjQRFXIH6Kmp52EK7F+qJDEk0Zu2HhZQ7SjycR8oqT
sL9h/Zq6DpvvMqS4Co5h/3DaKIkep0BpJ3KSI0FZZEr/A5AUiOthw99OZElGnE8E
ZB8m1wRDPus5rXUsaYXJZ/OFoKnV8loTC8WMBO8NNGdiFqyERocrYlXF6CDZW2tk
lKLkbmFra69uFLNa0+HifICeaI2nnvoNh46vCI/ZM4IXSdKqeyP3kKCBqodZVMrZ
943KKQzl4zna77aSfDdCwk59gecHa4G3shBQTvlB43xUl6ufGmiA431n8jGhIOtT
Be+GiK36MXXUIF1QiXAR0oI11btKVx9xJjKbMUL83zWz9E0TFLELV6TJHgfdafTU
P9pEC4TyfHKSKMWg5bBFm+D87XPyZeo050bJ/wpE20N/butKoLQvaA4E0m5czK66
o/kdPrwYtKAmvpGPgUWkZJ3uZ6gwu7hX3UeXj9eiLMUgo2DQ6/jawm/8tIBCkNj9
zLsMJiFPNHwwhIW0ROYW3t9LvRkkhFF3AugtoS6yxh0Gz2Xw+32LS5BZwp8DukYc
YvU3WoFPs5NDv4bKUuywznBdnwfHqt/Gt2Je6bEklGxTVIgOmpHLMst/21Ywxa4A
hnuvgdyjKQT1taifmdLtZG2rtjaF9yx/dqYOd3J2Ou7eLJoxCqX/sHt0eMQoXH0W
00iqTqDF9AEdb6cP5TzDDetTC0bjHtYD7+bQSonf7QXoiPfZI7/nOCv4eF5RAWak
n4L4q4OybzYy19aJkCJHcKxoD2lj8aoXrB2yQRS+GDk4lV9KqrVr0Jc3kjD1PxNu
c4zFOdCpIBXPUMe5efg8u9xzPCxwWKwuFjJX7bXwA+V3sdd+AAfYMK/mupr7Bwr2
NJkoRayRr86h8xsEJe1vtTUaaqdLf4CZVbbEK97yKpd9GO+u0BK7TrbsiSh4IRCR
aEKQ8c/zAobJJMTFAmw5UcfpuITjL7Bl8nL45tXi3tTWSS4oi8jPcbXHFXQUjLMU
9d6ngLwN08ZG/MsdCngBufLP2Bs/AL1LfPE2RyNS38vZc9E1ylaw/Mfu5Be0CNre
MgN4m7QhN2ux/sf/uIQedD+M4l41DnYFhFai0nLQ+63QFeRduYbW66pmwKGO5KXj
ygFf7zniUzCLY7WwdTGXTML9Vz1I3qgQnLMOuR68fgvmoBXJvyY1Z0uEMjdwdUAd
qsDtbRDzEItzDDol/4soXRLdq3T+6bikyW+QNwK97FFCuqChmx/QFmwJ9P4tqQFZ
n8X6dHtfkMvgZz49vdr2rsH2/OdbBAA4d7HBEstbbNVmv3RfhFDdUQWIya1W3ngq
Pw3Dz1y2szrn69DSX4uPDwX7IBryTzoqB3QkkPEGlB7gpZh+2tDqZO+Be1fbsygN
Peropy4Z01zT7TZADIl3s3a//uJEHzIWMzDXujkWqWyYjFOJqhJRrUKh4Ef/2f9d
TDUW6vyzUazdS4c3YpoHhHUTCXLnQ+fnlMeN7RRUOPzCAhMmlxBzVlkscEd7QtQP
bOdVpDzgVVAcBrg8QTIgLRDxX/rIWrsEHIHLdjvZaEIQR6SvlsEDGkcAUv1CArkl
Wp5H8B24T6WFZkWGrJ0j31xA5WOA2WNVH4URIIto7gAFY9QKx/ZNRpblhqtAl0lH
fdeapy14eIcJ775B9FuV6L67IUp0WTSVQP2Un0ADikgPLS/a/h7WynpD2qQKa+Cx
TdBQ+lAVb3olSHr1SYIiGJpoIimm1nwKdekNxAM5hRRVJSpk39yQfTB+/9l+YFP6
dwX8C9Xu+jvJOmBxw4iGs6uMnlsYbeQBkCZs4mc8EZhHk9a0PbTC+lGso5ZzrEae
72HMmzrEh9P/ADjZ2hpuwkClXN+9//B2MNBnr8DE0eXIQRLRIgJRgcXpVTPKqHzM
YghdyFE5AtfxUoe8msqpLR/3kLkSgi1AbuCtieb983FmPXLEB8Ulk0PSt0Rsk8tY
aervz4qgTMixyYsRYiver9vuVFIwrVnHAKKZNWNyDy+AAPs5/PamG9Gv0Q2+SlK4
VB3v4otpxX4VzGIztOJqTpr0ZEotoOaZa4tN7sR2OGWpRWoFWM8e82wYFrf/Edl3
Ow554FIUM3THU6uFNXaa5v2N3KZ14yV7HL/CAY4AHKGm6McjlIvceql8e/WxKqaC
DRB5utB9QxhyGCwEI8UpMzx5M4MHa2qQDEzyFfApACyB1O3PNSoxU+UnOPYyHvF9
y+CRk/ZZNmj3w5jgYjq4k0+zNgkvuEcOt15YGHnap4kJVKfbxa2qZ/uglBgJDNtH
XQZtBKOPLy8HqxLsp9hNAppTG9szBAyKYcdfVNNoyCtlsQrjOHTHTDSUp4/vQgSU
6/a3Yy6xAFurBWdTzueoFhAlmQQorV3mCPPGT6kmQ21zSIObvGYHRqWoiKxElNNx
WHrp5Un/vdszUv/tDgngGyYhOA2no15mtkq2JccFdHeYr4ius3aTohvaQ1/qyXCD
GuB7wnyrP47ZqJH1049jKi1tcRWFqnuovUvHs+K1mKYri66N4NKtmnYU2G3P8pCq
hfrbRJsbTJwZiyhpubdYeOpj0oIWHuOBPt3+GiKiZatW5pvuTgycc9IzISoSuTs1
jWRdHMOQsQyct8BU/01D7TQqPcqcm858FoQtO31YFLQRFvLSqE5ThzkC9vNc78My
NfJrJtLhAmQsMhzuXvR1qGW9bahNSK/hhJKozavWfYMDVze39J3BgBA/nE4CmQg2
T38vqNhbVU5aRJnPqNijM7Mj0kmG10HnBwksNoN1hK6be+2Fp/mm3UkKiWuOa0Bc
o2QUZK/ybhyi/n6ZJmBSX+swjBh7lqIujU1A07WpVtbcXLq1aY86NXp12wxH6bdU
zWVbMJsjSIrzrs9Rv2OVdVb3h80y4u3/uwYqdJzK5AkRlyeRutCD/WJi95LoRSUh
DRgSIIIoS81QcNKrb4sX7mYO8f+a7r0HF30DdodSBKHLrYEmW28vcF/EjWqPW871
J+62MqTmsBzoJiz3zVtzUn2Wfh42LEWqvyrCytyqrYs8tRhL2sHAEjQtW8FPUFPg
r+HwWFIX7c2lm+YMDpIMaZRA2kOO0P4WNfgm4Zkc8R1OfZjN+J2nPNofaEuINi/9
J7rz0Vm+4If9WCUCg86xncxdWP5D9bKZ2dxkStLYHVP3Y95x52lKsZU8EYOq33JB
zl2NbnRaZ7Ct/+PGKdPKaOyTq0YVCh3HyGbusSmoe8hSwLBr7bUdw+9RANKIb76o
xVNBRCnn4XlgWrnF2lbgnr4+7zBxAQsxrm/c583HpKkKOZDMiOdoAQgxF4JcqCpH
keh5jIKbuCa2tryhvohi3f9lLhRdAom/x2vE9fSgBaBDQ9No6chOZXDB0EtHOJTj
BTDlcf7b99ENIwkpj1XBsezzZ5+yiPXNDqmCKg2voDHJwZNC7lCpGfzFIrTUY4pn
O+7V6TDZgdW+MmMoqvv13x2ADK6FEM+pEjI6flGidDFYoyzFZEuHh29X5no/06kN
htFH05ndwaFB5yXGxxDgUdA/tDXBaroz4P/uZAfx+k9Y3p6xGbWHFMEPYoexZ3Hn
1j8tPHwV9YqNPgfcn46cby1+0BWgdb7dzrQonSEZQtcrIrZcROS161mw/Zpq7qss
Pf6IvXhHV4GdyYs1dcw1aHfmw9k48SV77qcfVIsCUE+W44Gm6SNpw35bpqfZ7Bnn
LQx1h407aOQqTzGqlwEAd+UIQ3OC0prgk0UE9Uwn7zlrM77eLnjN/RWO3T1cy7lv
5hoXBsx8XIcK3kvte1cDwanWSzWkzKiq+MzIbOUgdeHJ8BCch9C1s1rB2wzt7CWa
WETJ0Bik2ltYmVoRK1tvaUjgI/hc50ib90YpoTVfS6bGnES7v73C41f5Q7C+XcBC
QsOR7AkathM2bnj7rL3zfikk88fX8yloEBY5humxWarFbO/LYjDpTx47ToPAK2To
2FflRtr8L5xrsc9ddkkDzlw/OvlItCRZ5sbpxfUSxrQQDcA5763xCHZelsqlRr/6
yd/GiNBrQxcpO2feAZXh52p4V0lraBoGPcQEBHNFIgd3mJIPhzGtCqOTgWWkHnTx
rLzINVNiKL9O9PNI54YjRsZEG0Www+5u7T8V7v+jP2JpTfi7GavIOhuvfQDBh7Xb
rk1ugEtEUW3YwP3AUPhTCcqgbo6HTWQQSk68W45tfJaxiuzyi4aK18tzLuELXA4J
WYwTY6qlsxGzm5h4Q6bOgnH+aOBzZ7171FJNuvpn7XmeXZSobM9lnQxtfqdQsEEK
UjadFBWv0Vse61r4VIQ7+jPif5xr+qlu5yQmmXLuWTNaYJInud6v479PIXckU4Kp
JFvB02mi4ylwNCBTm/Oll+hOx0C6M5vRgRFdxi1eYNTeOSJ6YUVlTo+cPHUT3jI5
A8NiU6IipMwgy9KO/C4Lc5gEXD6aB3xOSXBZB10qZmeCFyp1I9BxIVbxdNaQdrTC
VnaNktKjcTRxSy1S2Zp23xmlSEXL4ZdaghYrHWK9trmMvETbCkP9GHXce2yewmGN
ZP6qfbbW+cC9dVYvFIOWaiDdZlNe9Sf5029zkVFrDDISA7Nh0jO85QKH7Bgy4kNe
RoU7AiulmwMo/VJ7v1tleGjyKf8ZijEr2wVz/kPxHnGcgU8HKndnI9chnCDAlryK
RUkeXBRTuKTqfjm0mQLR55yD6bQ/4j4sh2K3pKawutM+iV/x5xNVV5i7ytHOto9A
3oAEFVGk2cJq9a7NUEPPhZituGzAkAgDIA76anZxEFiysvJj2f9adc8MEgtw8hsR
HJPNRPlajuONyvZz86yOuuQLA86ymup1Z8i1hTVfW3QFWS1tnqXIJ77zIGzQ6vcD
Q6C4uLhvT8jhr0/o2Ixxml/2tvJ/beuT5xcNBC3vDbY/pTig5BGyqiieF85cmY9Y
p9A4xLlljr6vuqFLIW9RMhoPeR31DVgTG/OP4P/UoHU98byBr4YLLfV3guqE9Snp
4YpS8dnkp9WeXSA5Q09YZweHrG4ySjfnDpQ9WG8XtyX3o0Tu9VNQwXas/ZjlsVz4
+6OTl3nsj0yvihhNQheCN3VghMf5llEqSoJD9w6K7791MCFP7UPOgBY30LWhF6cA
57VWyvutTO/D9dU4Wi2qe1Mji3AtCSwBe9hMx3fNJz1W3nF+D4bPUCcJZ+nWIJxI
O9mMCaShABoY4kr2Ja1CPKQnwE1dizf02iiU1GTIAAkQYlTGaUNBj2rzm/2EqnoA
1PICiQpjtCeNlNxGJW6plZHMqa/2HSOrgeYVrFR4bsdVj1GJrBTLO5P2/giPjHIO
+ufXtfMvy+t3XEKJvz0RfkxOAUW4vdBUnBOOPsxUdjj05tEgsuJKX5nWy1kVX1qP
ustIrtjg5hLa7ckq/uc3RynoubKLG6fdj9Rj25q1iT0pPmb5VI1XlOt2HniYvS0r
Eueuk2m0uTYHrgSe3RmT6w8gWUE2XNoOVq6CcEmbdAwkHeRzsZ/t/sWE/mqGy+oP
xxfLFo0G7T75FC9HUztlovHtPIzhSU5hLna6n77cdKEEK4WWB1klzsPQTjcudU+d
pAYkW5Za7trgX4DCiP2jyqZfZzNB/LhzsjGhShkdYQ4TxoMiyvOE7cr2X6Xtu9bd
Onqp19Y0oXCJGbOehz5AJIFef7glNFftAXFPMTL+Kzex742ymswPISSTw996Ejgh
WAkhqMZ3QKfJre8yHhHv4M+D3ajZaZx0kINf0mI4/goIkMkC302lkQlFizdpUNId
R1MgSfqAZZgi1g47RMvoenFOJSiE+45LvhTAfHu2ffk1rjv5O6hU6sZ1a5xCzh8b
J2nxGE6X/yWtONetwdIybVq6cNArLoshNIud0Y0SqxFMGBNvp7CbjUxbfQkD43vg
0jXMVhInrPhdt2aGY26Li3OZ9FO99nJYtEVErJKUEOLhZZg8gBfnjTeBVCjFKx0+
00t34o7STii8R9W4UT7I2oXvZpT6ajnjMr4tSDQIX6phteZxz3h1VwGwxPrjjyCE
MfvsEhMPg5jGSgA7XkDi5TxF2HtRwHwfclvex6MPnPQs2QFvxlzM9eyHwbI9HqJH
uEHiqgLHLUZgBtYdnBmynaVIusC6s7MfeSro+uNWc0M0nCWJ8bREdnJPMbGmfwVX
1TXLkzavVb/QzoeEd8B+aA6qmD2ZZGatmAwI2rbQzSGR55xfpb9X7/hxRc1GJIzH
fF1aRTQQXAZLCBTrM3+ugBJM/Xo23d20UgW8EVX18nzY2LMdIdINiJn4LST2WyZR
44Korj5/2axCqCpPkNlxHhRu/wpyKg3Iuy2gqGx147E33b2bmV9KNoZMeQUDSvMj
Msyny2T3QBnokFyQRDJPB5D6MKB93GzT1JaqmbTuOJpOnKzZ2nHdbKelz3hCDBQn
KdzFlubXZcz8DrvFkUIQniG7u1dtaSAPadr2ZYMJ7fXZ60mx0RFE1xdKehIH5WWd
E4ZaE1TW/BFDgDswRbehrzgIRE8WwipTZrM9WkHH8nAYDvJ1shRxC42kYRcuitrE
vXy2rxLlupTh1ADI3r3srbPvdRYZcSHUTYLPzA0qv79CH5JFkd05ASNQSxGcH7tB
dGaCtsbSO/BW1vRNqK1Ih20fEjai9K43KZm9AqG1NV4IGRoBhV4Vex1neumMh5uL
9gZ8w9CQfdDGfwi9sUVfw9W4Eb5xu9PZsBumqmjentxrs+4ilwfN0cCKjxGJAJ2L
7LunTPLzT9VlisxWy3G7oKnRRePuERZyBtg9PIE+zThU4U0xp0jmzs4TdvVSuqGD
XKoqRWgrf6z0ESlbTQZ6IkSxY6rn6iW4BlWzsYl1JlEydKD76AvkhTdTpgOf1faS
1V4BAuylUfbkzATbvqMlwXLVhYU3XjmwnQ+qyzlaW01r9d6+djutcCze/neUMQzk
HRs4cRv5NOd3F2cVgqYi56DRYGy31s9If7q1HMYPUzqgBmvPHZUK228fAHbUhjDR
DjSI/nE5fZjx3epp1rLUGgQUwHL/KsrGRQy9/XOmcCMJSQ7rtz6+sIMjxZpvsIct
uXtRSF2sSnYSjlGGrZVq/OuS89ntv/p9ZZpoqLxwRJF85PP53GGgi85PdX0KTpDi
cZ7ZsJyAMdk7vrCgjOLpN92r0y/ozcCvy7KZvBbyGHHeJmuPLAaXJkKc75C80mTq
16nUZ1C7wRGUmMuawykCmiHGp6MuVv9Y8qipnhfSPmwRGYyKCMoMl7km2QK9W4m0
Dvz2MMWBqiF4NjadRBvZoov9cW2qns597dh30dDKdn5UQib3gCJjYR0HsSVa2ScC
1EzPVS6CzlImdaEknENqZ5MDfDg9q3h4s7FTcJiu8xrdN6BaeAyTZHLKLHCFEvEl
qOOmx4GaWrUtT61QtSha66cLD603v42I1NTJs17rSsrVP0CjbneF1Hl6rkIM712r
Z2pWfT6z4FY8BhMfYCjUQSh7MyJA9vfO9103rKd49RdPDovrFCTd1xmwMAc2M9iN
qLPpqKZrlDL3Kw0L15NTZi0dipUSdsS9dXQVgTJ5H7gcE7gvBkFZMK1dQ6SDAV+h
+L/6wXM/4rBpij2cSKAbP7YfrNHzn1vSDiYPBQemiJwbh9yXzIu/F22yFwkgGSYp
MrZd8Hz1PB1HSp/6yurTIcUlliwGSIM2aUEEUr4NX8wpOLHeUuQwzgTWxh2ftHAf
lnHys2asui1W2gTaOt2KGhqaChZSdvSuRIm1Zwa+XT3+S6zM6VTi1coDRNwBns/F
3+g/igx/2vwZ+kRyuUPGfsOE7KzApEYTHTFwfxHUqqE4qXL0opJmznFAJEUsO5qX
vFD2nbReFTmzZB6nKFst+fDW6Dubci3tYdU3F7ty6RSFrVKPGRRhp6ffg/YtJe4U
OezhNs5R39+OqaIX26h46CnDe+/vN+eEgDbFfEfBlP51QXf5mzI52a1KkWDVdc7t
j4dDF+qBhqUS4hSKq6ElDJh5xuDqRl9HEZURixO23Lsfw8GsNWO5FLEDN9zLL9Hk
w2CO2e24vCxmfCutwjS+1nYtKXlsdiFsoQq4AI5btUxLkRE4+ZccNrvLlX7G2Fht
TDCOCMx3zwiUk291CVNTu1eA0SDZf+PmyNqJ+NZw/lyehFKE9naP0ldBtE3aaHLE
XH+D3edGgicNbhQB+NJY6kTaP/+WTcpG3NxYg2BmNkyAlN59XXV2T2EMPHAo5NYI
BVNdOtsIogKn+zU84HGkz/M4oFbU+dShklArpLfDIFAxKTx6sBmrwm+Qsa4uYKuv
MAM31+It0w6+RzruAQztsYFMou4l4kp/waniOrzAVm3gdiNzms0QKNXxvEU9h3EC
VdufQ3Te8X5JuCP0W6cETNGLfOWc960UNmX7antZWHQo62t9XxsIV06q26xn49Qi
1SNTFEEyZ97aAEiZ8OSbxAncQQ9VeTL2Xhe0gMWS0YPY0Nk0QpbIIKPob1VfUAgG
Ctr68ZUX0XSXVgirprXJJhhK8dRD6uN0CORnZxmVdXsLEJmI7HdALnFe+KxS/hKH
FdFJT6PPcFLFz+k78ZHQOos8gWA76H7nAmaqOmPR2tw/UttIQRUeamalNlnLAK7G
UI/THNjVS1firE3qMIgD25xC041/i5lNb2B8NeXldLY0E7Dsvoz1YdEclxj2n/kK
4qn85nJp4hCL8UgQDMiArzUI8iRH2AXHAJZo4lZZl72hqiJYqIkvlvKrbbCeEhrS
v2lF7fE+k5eu/4mPsfoDpeTD6P+D+eVg8cwgDzSo7YwxWvi7HwSxfbixyTOQHMxo
LRkWFf9Bku/C7mrL7O4yv89fWbtosqsuDga6JoTXiYmx+FQwGpZaFLzQPg79qpFb
0VNZsR9BsIbrLuY6ZCcIYqZlVcikiqTdon+OS2zET1/urp+n1jKfrOG5XMQY+STp
JSMYq8l+w4ZWrGnV2Ifgn3C2xVGOFy3hWxHrFhlpInNiag2uDR3VJidxGuLxfq8R
SoGbQCOfg2xP0y7X3m3BN+6bFZdDGGXGtuqoO9A6lpMVktzZhBx7JvffkWsgEW3a
JRYkGDX6ynwmsgShhpbcIZ8ySAxqNKf5IneTGsMUnqTBOkYRZGhPxsjKh1WXx6TK
3UkkxdxaWX59LXHZ9UJ9GdNGQT5erxv6hoPdgmHtXXI6FbY8YAQtCITVCkqLuurZ
IVrS09MkYNlU03ak7H3kpFoVIY//wBU1XHUQQ1/Yl9jiSCnfRpWn/gyZpy2JPPWl
HSf7OMHvjxSDpqH0lyZMszxmGoT2060jBlDsrpNdKvMpq9SwKBc0YN3EMQg8FCOI
Zr4oxT0W486ShcQ05lkZFmtsr6EfsaVLT8t7V3WThGvpkAa5SHJBg755M96KgAGk
+Akn33olauVEvWB+FJ7aIUyscybz7cLaIzYHMpoxfgyArdakmiN0+vYrkAJ3nrX2
/Z/B+V7A2SSMFNOEyozstwAWmSaBkAzGBUShXLUUUptXCbHWRY/qqwgSPHgDd8wR
qa2YI5fEV/nrwelnH8cQnH+Iq+V1AR2K5fMVGi0hh8GFaJUedOhl/P/z4xqxyn+i
wZ5wTDVnWBRZpX4+/oLd9SHqdEU6QvFc4MC7dD3KGbihzAcv1K619l4BuaGnSru3
7Cy7E0BJRriETlcKTW+ADEGyKHoNcBP4dLqTpiN9G+f/7gWs6IeVD6CMw9o69WLr
LlAVE6D2wco9P5O2tjQP1MRk1fv4JtVUFbySUkpyPfKgmvg4RG9/nX5v3iD+cxpT
nPeyvQNMkGSKJ9FdSnQyR2xcDMX/J5pbr7wtYl++rE3Jet9cVpza3cordM0QTHqY
a/9hRO6S1H1DEIXrZ9gqSQG1f1zJIealiPVN7OJQf5rfqmFr+CAF2QIOZRtCyqum
JRNGk64whfJNf3VjToZGtujk+Ubir8p5PvbllNFRwUnAI86i+NBldgLHYeI2GlGC
O+QdxKni5yqQC62ksI4ujEpFcK5v7Ey1X6oDHO+mZu3VA6GZO+TTFo77thpOGHdH
frRyiMqrtrDJcb3TPNgrRIhZH2YFUOpRLK3K4FjwQSj7YlELv72Go40q9MlLrj3z
V9ZWMOsCip33EIeSm9UqzuDzvxnBwwr7FIjboRbUbo01az7w8I8V+HpwPh2I9dX+
8PzQjmonDnscd4Vey+IzNBYpm+DLBm8vjVLRSvaTcHi8kOvrSRg75+Sa3SKOqVtt
n/ZQTOxQwKXMUEk/c7EEJsA1PQGyso+Bj/yAnrk1fDKiJBZIoRPEKmBQrK0kuanW
POM1b3lhPiQhLO4K/a8zDJeO7aOClCXDawYF5qDIaC0vp5SEbZnfaHBMMirVpRGZ
xbcKvkjuy4jxiZWcpMUI5/rY9icjs4sK3rPct8wao4IMA/LutD1sqBzvrDHc9+Bq
NNIRvjGAkO2Y13fusw66gON9QoeqTRs09+XdMfwId46Bu0pPoncA5gTa1kD+t/lq
Z57W9owAfYvnwplXxhxPwc2VnJwHjeSyrwYD+ZRKPi6+LkOP1qUoncgOuwN4dznm
KAzRg+at/zyNauTqe+/0vLjDAmD7VV/lKfgqnPmoIACzfSQqwnsglpuX46JDBEYv
Si0e6tJWqohTAJc2YWPZ1FlbCSL5KBw0GbTq8estoxuE/TC9baCJrMT6S2bAQqSr
IE7NziyvVFyBFhHmEznFZE2lqzf8zGOfdhIGnHlRZcAUNDjV0sgp5R5FCRpns6dC
0jB2T+6M6EY4DpGHC4V/QU6keiAXDpJ8Pa742xpSeQhHCpiTjQlwRVs2J29oKa3x
ICOKLN2DbEvfySyvEgVurBZJWa1kTDYbOyo3g6oKOkJgMcve9qXEO4sr80cHYJwY
cBXDtx094BqFYZiQWkNyh9G5w0PWnES+nmwHK4NFdh/XGURCJ1rvVwUqFA7qQNF4
+VeQK8905oCeDGaE3KznFcwEEvNrJwWsF7aC5R4Ucu5CipqRSF7jESHn/Y4L0O8/
tqOEyMdBzmx4QnBH9vuX82pmaoasZQ409UmgJ9ibEzf3JKh45NdbN+gAZj4P2zin
3Sj6i0ViMoOkAvG5ILd0cmC50DX/jebMH/11AT6jtSdIGs/VTMF7eVLclCVxSeJx
XVzMfpjWIxBaTbYcucDTepBHNdtkicVjFEJA5UymxFvPtat08vhmKzwSKUQv9qql
JYFU//KlClWOLKlzB7ezHPet7iLuvQyEk1EyU+MwABWMNsqYNu4p+z2eBzHUrYdJ
ExiWDOBE6KvZUWGcb43siP1ekTXguWiPSBz2OpUfoeKUF23BQlIlt5WFfErZpKXe
yRk4dMGnkNWhFYQXV2UrmObCPbvEnAp05os/kSzQME1G//9p4aB9OKeeIIkpZ2g+
wzpyVGbW/giCp4NO69bHXY6C0YGObKrq9h9ckuRAV5Qy9+FsWE1Ydh97Fd3whesc
ZA0iAcqJ1NP7Rdkf/COeQwFBElclesvQfdTsZzu3zzJ7o0SWiSabwEdmGezD5oWR
BB/1p5pg2Xfb/j/ZJ+X9FlALOupWSE07Yi+3q2sFArH00bJXeBxtSYX+AHaY21eg
NBMkEx8MGn9qyXCD68NOvX2gsrLL64TgqKVMvN+4PeQMhANGPQA88lkjLcWz4Ok5
Evm8r6xt6e0VmKAcgLx4bZX3qIpRZ0+R5WVKDMwPlTgKudpk4nivdaev2W7oZfs2
PEio1b7PV6YN9iu5hewtgobi+qEt7HlTFbso09E7A3/m6PqSnMDFyMV2tXGdw6GC
Nti6pGUBJXLSWz+XzVaD8E6nDMH2uXnEH/YUzYiTyIxVqSAQeqsLB+sdnxDgmvIN
SV9uJo3VSkFekMckq/NW3AeM+mfT2Iv53eWhgXk7tVvU4eYfE57m7M9Grx3niMDm
kxYuby6GDmK+I9GSyoG8PkSty6XCts6nQSHlv409732kXz/kYG9l6nsmxM5U0/E2
gznqhLKbdRLOMJp+7LRkw2gKTWId/Llrvls9DUIPJa/Fwghx0RnJfVi395K/kEkc
QjWAs3c+j8498ZweZ/W27cIYYxEzBijHcxJA6rEtlIJzTNoprgRXd+VYOYBL5uWk
WQ8JuLbhBznVkT4dOh9RpjR6rF3lWZXYe0m3GDLkX6liEfB7bTXoTvSWsQc73xUI
BC7mfRlTwG8XI3IIyBZrt0RxtuXV0H0eG0AznVNScc4vTcVEpDGzbfMDDEM2dkYc
JihxO0Kg9OubRBML1tl+Dog0eINioV7M2yG7CztJd/wpjoFXEnwOfnNzCXX1v86I
aK3B2xjzcA9Ob8P8akEOzDTqQm1cx5jJ37eHkQwosbPdH2k2a4g11BiTFpJnf97N
0x9X+CGYOmFVQWvMOfjngZZ66kmuiGPG1gRy4TyM2SrHHvSRnJ7MKYhd0K+ZMfod
wKBoc7wfdSsyDs80LYVTSUaAybVsVfiQBb4e/w878YSoaEheAiI16X2mmBZfVSnE
SWMWjSYxQBFqiIeVszEOsjPe6s8GTO0LrCD4QdF8+0DXU1cB1d0IbhZGrZTYutP6
RmPjDWDaa9xMnphC/WSNQX7MiV5TG1Nqrkjgl6SBOIv1VatWbJaqHQd8LTo2Ta5n
BJMugyVfR7/mRDuTzhuN2oemzb7QMlA2y8cZjJvm6yL/bt6wyamPdXfEQHTzkkYP
bUk1KWxiiFLyRXdA6PrPxQrqjv4ixT+3Lr5v6lUfDIb6YvnAnS6TNArOp5z1rHm9
xyP56kWQNi5gRKp7gDCgDguHjy6bzO8pbcD/OEvmCgzaf4XWrR2R5kNuhCPRknkq
icp2+MJEbft9QoCmzTHcER33vQlnlADf8CQ07KxJXt9z19+uXA5gXixRPs+6Qn+O
G4XK1kcM6xZFUztTlXQLPcvQEIcgnXMdWQ1zCjK+vCDfIvwIzazFhwRiwj23T1zW
p1cK3zev0Fzj2dhr1JudxA7zPn+nVbzpU41ttROmoBspj2N0FewYhEkHOMAnDRAT
uUu4hr9fNCltpTz0oaKCaCXXS5Y2RDhF/qoofkbrQLjzB+s8LSkomxz0iB7fFPlY
K1r2+FHGhSPQaanZmJ4AIlcysoR4Ba0bbX5q0J8aeXqtQpN+mqDAsIg+2qJbqXkN
P53uNkeDNYOVQMbbslJ3gLsoV/6zhwKVN9v+A6jU9hzEb+JxPNTHti5tK5Zhn5CC
YjC7Maf+eua4xu6WrfA0dkhC2Qns1pZn53XwoAX6faShX1b7x+Iji8RpdH4Cs1Dp
iKW3dL/wVlEbsDHedWNmA7hFWL6XhQpg4R6fiQgeHkFuCesoUYr2O5GGIBG/ICbw
E+ndTA4DXLLDVwcSp+IBM2jOc/yGVt9sImS0IJM2FxZJnY+dN1/M7v2FyqInCDmg
0ArCJ4FxdcEzSpK5CpB+3K50bJd6HHxwOZIvYvSqA5sDdNTCq7dNIu/oA1npOSHM
8igJ8dbOjF6cKPRzEgAqTff6W6sV6qwgy/ij5thlN3Ht4gu5/W5AEbJPlPj8mRps
0oaABBscoDHzlwJ/cceeItuR+o/wxyMmxTEQAURWon/Jld9AMPW/fUEMCZ5u5+n5
QdqP4RqztCdrVanUCWcTCafUmpdolahYlN56CkBPfH1Wuop2qhFqTcAbUj06udCY
ixERf4K8vjUytbohG2avuzq1DNDmu1Yf7GdRXXr8a4ENWY1nS/So6lc4hXruUceF
zmNLqEWzxXNLEBshq49rsbn8RxSVRIuKKyUR4vRyIB4eTaGALUk3C78zTmvset4u
JHA/cXb7cfTxpmSr7aT8oySJwx60WVJW+oLvv2zM093kDyg81lMkCU5OTbHsV9xh
/QU5wmMEkQ5SLE7S8L3SetUEbfH4Ws2E9r1nGZEJan/W7FMc6vffO4dKpM6Jeqi2
kcA4UcFFskTnapMnPOVNCk5FAz+TNn1B3NrbH/8uJVXf7mgTu6HxdL17NqqwglxQ
zsc9eRhPBrmxszEtN4cHlxMx8N7ko9L2JW/RWPSLlM0pS/2fGC1ZkvG47n6onAEZ
Mu8KgY81X8CKt7LQP1ZmJAMj20aIFIkwh2+Z9OKgsn8/YiBz/B9GgWtL1Dl3AqvS
gaPv5SgCeo/N2v1rgkqe7RLwd0+KF0gV1FpWxOkRsuoXRZlY3R8j/nyUObP84sYu
MZRNhStSunkaj9fQjB1g4b37+yqfMviDQ8/P7qbUGg5l8y66nZ+on2wDbQ+BUX3g
5ggcPn0cfLgg+iIiJMfzb9dHxm+H6JYkkP59vV08z1cGlIzE71/ApIknFlP4SnlZ
/bh7N8k9auN2OnwMn3X+3s1U3VW6uHznW7BU5BrBq73c9fTPYzuHwc1tmFpz9XsI
QokEL7B4zPtMBHsWBcFux9Hhtloyi2C5rB+RTjX/qzJFf+cpoikibEG6su0IjhfR
y3EcI1N8jAfVQmX28Jra7AL+YREdTOoCTQEPC/rlQT0F41TeLd0dHGhomrcooIoi
Ci3dXWKyGfc3nW3iRYtj++Dg2NkQraDmaoi7HDaLUq+6ty3vOZIQCnuPBRpXJIxG
xe5fQw23TzKrrnWHoRIh7n3fb2q2AiF3DVg3TO+AHDGJnoFv0sl+8U4BkML2Kx+0
qtDurg+w3PQyn5uNKqiprCOX9nWxpKM7L/SzDJ91WSQAMgS0ZfGfvb3MnIX92WMk
YelaKSQ9wsrmYXtpSuXJg1X/e9S+Nc68mcbB7HG+haSn1EiXo5Tss8+N3To8FKt0
SX2MW7j4kdghKD/Sh4gBW6BUViFIH5dcQzShEdQvUtGG8W0vJTmhW3wMpS9NwHir
is1M8UJ0AuYPGM8G47Pq7NOkmxhtlCVCDt5ngk0BBYVNP5GGgMX3kt40cgoAEZCW
XVW8EJdylelJd4djzoylet4gYwBXRc6Qu3wT4/Up+dyp6Vj+QB+eVAEcrHZvDaap
qTE/7OVSAp8CXouVMZ3Dx2C9sHhnj/x0nWFsqcXoPanm704ljjUyZDFeJbOwC9ro
nSo7lpYv4Dm1Kvzm2g1qKkKPvjN4vCs50kOxwHCAjVbXlY9nCIe+OZ1Yc3ygyvc1
HPbwXH27aofMSsew5ZzBj4BOx7r6Ojh1c9hWngl9bj+HbyIt2aR5zHukh+8OPDEO
4gVCfUxBgVzjmuVwoaOxwx6ZURJBIRCyzSUSTK5hkLy4QBoM/PLjqPTzSEX/7lKc
O6g/Lggcz+pQt366Nen5jW0Gy6j9zz+4idkjn00qFEvBXf953nKBg3bCEbLD1M8q
F4Wnt4bQC7S5MO2CQg8/xMwrTdtRqUjGoshOisLiSAm7AHMUOOGDlVk//oXUT084
stWlADgbQ3HkGDWzYl69uXejFkQP1toNyUYpS2avzx9s/ob32OzTNziDloFoYmN1
Kjwvjc25HaQfLIr4rOPqfdZoQEZ9Y3Kz+HzeoOHHVb5myM0KOCBggU762lJkMyDI
rZilztWeK+wTq0/zmd3N5ImGb+QZJW5WQQcFsrBdeiJ5Lsat5XsIA0z5zFBT16zw
YGHo8l3lrXnbwkewrSvIF4dY0IED+MALzybJQc9eQXzE8tXpAZP+W9KtyPtbSwFO
4YmBpCKG9zRRuKipBfKXD2KCh5698ehKut3kLxRwhFItXDrmVdYg9rp0Zv4mJnl7
w/72JH1uL49LsiX4mTr+xmuPmsbNNR+hdTAK/tWgYXFRZaOAyczMhHd1L19COIYu
qjAopfcox7jyrnsNjkesZRZqV5h4t0UbWi9CbhgE3CF4hIGB0HBnnqnBkIxNtTmW
WitkaGTtcLZXH7chd5wMKe7NF4B+1A8qGVpju5r7r2kD3TiES16yBSOQtoRhSsQR
Zb9403XzasBfYYlAwLAPwBkfNkXDfv2cdjExL39AzBEToVeIVmYermkDAc++HW/S
6kjLgSTH5QG3YfGq3DsrJPFW7uLZU6khwlaipmMVL9exF0NALknNYyaDhr5Ny+LT
HkfkxrRiLbSTRLRrm93qlWN4Cr6Fd4p/sK1OEYIBl3yQV1S5rS1qarP7IyLB1bPZ
KP9GTDS9uEtAEiIfqAcmQsacOPd3M6Hlqz/iO8L4p4RN9QqRyAddWYVKm32Szphv
OSesW7GnobJ1pfzqQTSVj5O66bdksTVFxNSjNTFkhtDbrOjyndEQOYsGIoKWJXlK
wurVNeamKLxJCRyQp27nqvvwgQYF8dXIIBzNpCsj5aBRM8PrL2681EQt5XGfB5DR
c+DF4JeZxGr9Uq333gQSybHzXNMwFd8A4TYGcpy0NrNxLnJlBup+ooippTOA1YUP
M6k/V1z7/KJdHW5W8AeIrHQD2OAP3YA8Ig2fluTT9ZceuXZoljooyz5RcE+MGceB
wqMSppRLODZZvMptUtBR1LRRzzLgotTJenTbEOhNqxQWKdUP+8VOKA2HkvPG5iv5
GzHc1w08gRGRoV+4M3tI8CI1wMEOZYtChwpYJP9d/dG1A4Rb3dUsAtdFwGXWtHBQ
NOLLXL2eViTs4fGdzyEJaPXPTg1/VWoz0753W9otmQ4loDw1nfd9tIUQuJbRRQg7
MGQxruo4FhbfIjoi8jiQ9U+0CB4OvPNpxT/+xIrG2TGjLlpzXOXoayEsi8k8aC0R
znCNxxSiGYFEyF4iwCg3r+Vc8l8Nh85yBBbxQPfO7NmYrA/qcq1trHHbkI0SMk9S
hf6H6X0+D37VYQOR4RaOuyVVX6eBnSeJHPW3rryigEl1wNUNWBSGOqf4NkCbfYwI
gvcNM86CcigEdAtr1DtaKDh/qh8WJ/Cw1DRrk4jl2UT5fJyG7LIgZTVOjP+EtTUd
YTK1EVp/xJsCmAoiyhGQWAA2nM35eElhtr1/+4TQ6DXKfeyIE5b6xLP0Nlly03H0
1HmZjPjuntuecGFoUjztDAwwU2IY6jTnNYlRJYXD/ucBQO5HtjWGP/JFN+UKg5WK
eO8JcycIc2eh+z8dA8b61j4BfUNgcFFAW2r7AzCElaBh0dpQKuFmg2W9ziJ+5Tee
GIKXAoPIZ/mJn28BbgwsvrWeJHQo7Jjv6QbCYHHNHpOxoE84+M5GW0inHhlGPYcY
9wQYH+Bh5vtbHwMPoYghTc8h4kcGMdVVSdk4/Npd12ZF3sBITWw+ZKMzvnGKBjBL
ZxZfdlivQwWHBBKguhL1z2J/7JTpuDGx/Hub34Kp6DeKqzDouTGwU7WuiJp+U5kn
dsofPLsZEypXoBdRZoP/st0/DRryCcLHc7In6IeHDMjxdU0j0gzCvPMStlIBUXpn
d5ZUZk+DrepIEWqKWRjN/NNFTAcGQ545HoG+kvWL7Rkh0OPbMlZ7dCDuB6n6kNHm
+un5SN1g+suRo84NmATCqOWO1QgYedOZw0/FpjVqI1f0fl0os3FBlMOgPI8kNLLp
BZ34cI9fSY/JexXUCHI4c/xwK6iQw4+bq1+53duJmD1FdbX9FwR+vEXe+RNFdgil
lQw7EZ7dsgJvceavR2ApJAl6Dz2fHpFFnOvzCNJ0l3y96IyYzF4DhoRjZvS9KYyw
k8MnI4VWZ0TMien8Hn1dB2c2XZ43OQ1YEWD7q8TTJ9i6jUc1rSyZ7Rrtpi89P84E
dVXLeqhwPgDEMgPioGTvfEIwxpMxEzVe4WERK/BRCdobUml1gqxL/PKTjsLWK1tO
MwJApCjlkL4Ee2gjASQ2Hx8IZEEc+MtpIHKfIbWEok7YIFN6SFA9nLiYZFI1WMtZ
ojeeKVlgpgac50HCZyNF/YnlMAsi56QetSohnQbqBQk9A+jlSOEK06iML6tJBUjH
8gQ5yuE4UNIOuL2hQlFhwvoc8y20fNqMaRmdDdL/3xbd4VFkPC/+kUGsU55s7k24
8vk1+c93RZrHxs35FgzKkxTx2z0SpbgrLnF/BiVMipKysGX3amsPlxboC8+6Yl8M
hlwRA8QtdkxgL6lFnRuK5NXQN3g3ykookqCjxz1WlSEMNMjBL6SRU+8m+kVklFYD
1fuj+jCm7kNmXVU2MzT+WYU/1tk36Ffo5wrcqxjtIEE0faJ4kFJnWj5TCT8s1hbS
H4Eti0kJjUCPx1g15wsdoip9iMQ0ZWo2L6wkOaMz/rd9XfhBFatTBTnvPJOlMDI/
cKqsFSdoV2Yoo+MiD/IWpyAeDfTNWPc3sBWjUCQU3/C6SJiVRrknMf3BP/UdDu5D
V3CTUwTiv9e+gYR8h8mNYSBRFrN8FIklRdvWqNnQo8MKtC9AcHUHMFHd45McNj2r
X+4raeThuIHqhZrJ2hK/bN0AuQjd2NVqI4SDycjgCibLc+YqMm1jt7MYCnjHWvzW
8oeGeJZhXWVUd7/YxAM7JY393GhahSw3MesHj2g7hi4jnzEovsXjLb/pyOB9WhDM
gcLwWBEu+M+xTBlmpLX8J2Y5FhhbdVJdXVAkjNXBMgOik4fwYw9C9jd1wvYltu60
A1NdM6mcITAsnxQRMr7FCXd8+epYx1Ngkg/OUwBouv3b8YryqEPlqrtV1qwXxOTo
bZhh9qVwy0nUtGLETY24dvjT5FGuN6FT/jFLkVK/ZGAJGvwuaUIx4Xj0PqAOdnua
4vGev879vrWR/2zAeEATc28eTLwEVuenDZjbAG7hoBr0ltZ0A/fA3lblW8lm+KeY
vN0YU7aJvyTtSumywXvztF3ZLJJrJmsP6iXApCBO0GN/RqYbMZyEwA9rXs9QOQgR
FKmpy0z+GjezvwDSuL3LSS1lV1Sna0L0NB8/LZAV88PmJohMMmi4rjX05bJwrKCL
LBuBRRh+icZgDYHhuZ84G2ImlI3nX5GxZuSa5RnGs+TFGVf9rhNgIsbfVNQfoCRO
2du6s7Yglw7EMO59PPYVQQlwjXignAAUIBFQGRZelnHnSlTnw2MkogfZQ5UJHnLM
JAvF2KnrQuTNIppyYPdCQcGL1gpLkLKwSSNJXGci/uF4u4afO0kAoqzYlq0c2vzp
1XPjvgNMzax6jRNwyk/tHBRauGRGYaZXex4fZXbTaWeKGPIxLuCg4rx9uzF39tpR
oNmYDlL9WDA9bs3aZM5GXK3YNYDeeuvh8TBTkMGNUfuvBDfI9p6pDWetNEZ0NvHd
6x4ALWX5nlcswihyspHtRtDbwBfAE9pQQtzpUY6e2H97788PF3uwttUUFCyQYIei
NDEnE8uRzPAwB4IfIvMLrd7K4TKtkScdnx+gCw4zpm8UMYsnnzB9I8Jrgm0szlYP
ZsQOyT8lohzIcCBTfkEMEFigqEYuoRTFlwHoNWomOY+CwX8ZRN7BvUozmLyxEw1j
xrsOZ3VvNPBhH+KQ+xx7t9t4fC1xB/+K1qxkFizGX1Cne3CL+O59DbWjUf2f48yU
ICouo6qSbqoRyxOL2c4i8yyHpBfU0MlXyePF21ZreQp7PTemVQZatYEZE/X2pUJR
cgWAiZAzFasWg2cTEtbuANoMylYBdrajDyx6ADZrr99AOHBxSuEF6A4SlOMkt5ez
8Ibba9tC76YiM0O4F0QGMioNxoRlIQtN+aX7CuMjewOliO+jIHf2KUeZeL8oPgoO
i3eZ5ftaZFiKmVoAcDzNLOJaAY/KGTzn/h+mfUs2/yjmL6sNZ6LHli+dMu1T50B3
PiG/MStlh+25687zmmcoR6rfWHNz5skJmgB9AXj4YspjeySiGsZbRGYPez7JIMVi
dy5gb20NlrNgk8PjlZoCprMmyf/771vfjLYYvuNHOCUhhjxIKwq9vRvDV+fBHG1/
otQ8LtDBcMFRnN8tFz+U4qgbLl2mYNzq3is+RHgAypScbJ+z+VjEu6k6ltvT88MS
pGOXXk6bZPRpbFkfuiU5z79vcHrltKlgqSpdlfYOu+Me0MfWjbNjAar1Dnk5OJaD
6cWpp5Y8xBf356RKd3KJGNaw4tiGAmG4pbLEyBpdKoJQQ3dBaOt4mdOdpfBm5Gnb
GWuWLTzlDSUVIyuYXHvGnLOi/IhEWtE/zvgiFwFuwTXdogJ1o1fXOWgIa0w8+Hvw
hXm1KcTDDWs6OOUqmamHE8wWwXqUEDuNCwjm8xFu6uvSqp283nQDL7Ey+ZdKnLED
6qi1eSrQ1z+4SH2cLbxeQp8HBUwrtKL57ExFVtponMphsfdGSkA6zQ5vYMnvLY1b
VmWdH/Elc3zwWcghxn+W9Cev8sJXZYFetFGlBiPwJrejZw9h8IPeesu9UtUgI4V5
/7AgYfAEujUxgl+LwGyi7z3uM57FRQKKNHpR0YvMuAId52OySiBOCWr9zrsv32N0
jIwneMcxP0vpWbAV4vX0ROXTxbeT7B/2PxEPx4HNPhqxQI/KoXPMzqQX4/eFb+PS
I/IwVj+2kvlCQndvVxQhcuUEtvtBjHwBy/WJNuT7zm0y4oILv8Y52k3TfUokmi8F
6aoFNnjAUYoWx7g+d/mVjBJYtg3Hae4WKFFDZ/A5oB1nb+ixRWCUnrBxpTtufsuR
KZrnxKT3TtLXnifOoopx6PbsiY6mcwIqdZSFHhZfel0OekSJbmXR8okzpEsHkpQJ
Q+WKBJO+Dd80JJIsPMaUnhYzhcDTuaCjcSfIHi4kALbsYTFZ6nqisufrTVSfpEtC
9covpmpzNRSnbwrWVEX0mKRRCAaoPb9jux/iM9RB2AovzUd2aTCT2v912nhCt4N9
ukW4B8i35rI7eWqeN7p8DYve79LbBG3UyTz3dn/mnMhtuZ9vd560N3Z8Pj9RgVvO
00JH3//6Ymr1d9i7YQh8RG0kc0qnKiEf5IxoBk4VYZgd+UZzukD0nnPKodTyL3Uy
lOcRxERsXPBaI5Eky/zcLzDTxPg4U3hE7wSxYAhujJQkCdXnie5cpvTYCk5wVEMF
VVZIzCDmxpEJANHJi8k8p2dDkMgMbHVq2WYWzKUSKzhWkzaZRXwo2yRjF+SJcaDd
oC0+wQlmRD0d4nXG3t9zUBjghKWGH53XsrbMHIs5IQPRQLKtgRSbWnhw0KQfFW9N
RJ/EJFvhUIdWkzbQ8YJMrB3mwGIfBi4xoRCfxs+Qjnq0wjs6kjqo/dkRNNvXNFNm
bf0Ky0T+qz3fAUsZR+iaep9RAcGtpCYV7mdwmG2Pq2LthDYZlRP7paRkqDvSfLsE
YeWauE6Ve5t7xP0kj18DcsIRAAHot92RHgC3x0i4nfUAJl893ty1d9iNI0Z9gGvH
DPADvx05Xqw7nJmtxthdZIqwmqo7OVEYIF+77RlZZJRqRY2vy0Hg/VeWsyEW5BIs
r47G4O88b7rLNFjtvDpJiv8jxWP7fLubEtL5PPmPOztt2MBzmwenWAx5LzafQ0xT
6BgD0778i4NOxumLkbBs3y2vMTmHvmE3vQidyf1IUYIcPDdRJ9cl1sqbUkNfPJI1
aiIZFpj/dxOL4rGCB1jk7/2ZYQUnSXVy3Pt4iQN8ZLT/3CCmVx4ONcRvBzrOIRG8
iBhL0Yx4wIKxj/npAdMH+pbEKW1+5DuHbZhRJfzlvDblippKR1V9ncjrgatpmLx9
lxhQ3Sv/T7kX/WID0bXiCof3l6lNjdfhn5RubftHLfuriwr/vvKoFo+t2ha4BdZW
e9JCq12SPNQ0PmRPzaGhBmPVDmBrgU/c+HXknPgMQFsI3qJtm9LVu+qbaUCyIvKz
asZaz78u9l8A9KkF214KQL2xJ+SodMxSlIVNnDYpa2r4HNyRSi8SrdcSSCDN0drv
BdoL7+0jkv6vKWO9EGi8NNhXkirC5gq3oZpGxVrDrH4f5liUbs8MM46NtQesIPIO
1cRa3fk+P/whRJVLn4Jl1rC7PznFN6v5Am/uD+QqopMJlwMDDIe6No78CS2knB7V
n3Su8pW3SrBRjROslGe+8RMySbz0lmZdE2abXtRWvfrJxwRPQjqlmo/R/3WUdpJT
GicXrSzRksOKouaHK8UUgxGHp8TDxluVocGkQyx2U7rMkTLhKUL1A6leXBJunKvA
tKj3pg55UqJc0dDWpIPSyP+sfg8IjTzrlbqgz4tYRKk+DMc7vLr8ceaHN0ZUDfyb
IjJ4U5Xy9dMMaqsJvlQOjCZlMkKGJuH+c2zzORNrJRyJzTdG5LaSvV0fDxIP/ndV
mrxJ4cR8bkKtBTs7B8rNG5ySWu+Izzt1pWsRPV5AcQODmcM9KQJsoBo3YgDkd8ro
HVT0fnyJsZ4+wKaNX+MiP72o98Cd0ijQQZ95mtX8SAJTCw+/JVVEGSvRWEInE3+e
bzRYyFoHQuYxjjaE273uz7oeYxwQQjrfZSaEshbdIcP3K7Jtykh6bMtwE19tADJw
0WCFx2toMwUbsCjQtxgRcfjhsqrS4Qdq/GDsKAex44XXIVT5CV8mFy6gtQtp22RL
E9qwfp0uNZWeotyWiw/dFPUkcVrt+EH5IqH4ptP9EHTzQIPOL4O5sPfPQ9zUMhkI
vhrctgjhPUPEp8K1YQW6G09l4gNExx2cRqVNy/+UE4LqFh1x3femLSqtYyKwdOFU
D1nJaXDqo0tuS2+wPgu2wX9w0hrEmc5kFwMnRveyXI8NBs91E9GDDGOdIBwu3fhH
BF1y6Lsan2rluA/Pt7YKNOKUATppmDMF3LEeqEC0a1SQ3kRDoKOKwDPHl+Reo1cc
D3NsQNuyx0GGH3Nczzh2xaYNytBQsUl4Ohum+Of5YHBL9F+6bzRbB58RK5frficm
g/q9SXosodpkYjtNTtTmKCciJD9UuB7+M0Pw9BZJQcuHwqMueB0R3X8SD8S8we7I
nZBBF/F9s2pWNWydmwYka0J6+SY5uc/lgpak+vSQE4rn+h1GpD1e4+vbt+uMQnn5
SUZsz/4dsSJpSyGCiQ8stIQmIBS6/ukYSiZmGLE4Q6j39awdgWdbSBrAY0wRxDb5
MY8D8SU9aO4oEBTy1PbKdzj4uHDVQ717udmE5woQiczsbbVN9Fyd/9vg2gCKXyaX
PeNQAsiciOsRqjXLsdRQgt8Q4rD1OucEVjeq+aqDwQpwSnBrAIZ3tDbrKbXmqWrW
ckf6WXy+x+wwuzrfbrAjsF47PxaA7O8sqIniLCADJg/i6lhhqCQ4DOPkPOSvOtsp
B4kbKL/xe0604Cex8O4R4KpJAuB9aYBAywIQMugs8EdwVtMMaPZF5XeZM1KWShEv
102n6zPkMgRTtQQfEzPazpWsmiuWNN2pUvK/HjTgGsxY2GRrRO2WMGyQqLvHubH/
8Q+eJgm3nR5bEoC5CyOvkBphCazq0g7XnY5FKqtW+39MZnaNvCv7lhB0GaeW61s1
9EqmIc91ZMABGhHdyK3+utVBTAs3hAJROB+JZUi129vtjFTWqDhAoa7Mh4yD1EYg
Zb43t/qcWWrOvQQ+VfpnSF15Ll5Cj6SbNT5J/psjh3VmOfi6t+tLrbOs7rGxuJA2
U0FADg3q8lsd38cwrbGdoqZGXz7MK5tTvZdFVMmTjhHzmh0O/p9sQVXJSg2EnkFQ
bb0DVnBRvVQg2NqpFSVSKwKUS8S1sytfUxRei4RWMUean7VRAq43l5E+FTN0hQvW
lOwp1g7P/FLYoQZapxP+XxwtOJiB2kGjdeaM5QjsSkWZ0htXkyuEVnMRooMUuczD
JWi3ViXtFgbDZwtn2Cj19Mb9o7T274XuN3TIe1VvS404iEqL2KfnC/b3qqpV5yg5
zNCsKmv9NcQOPNFyc9hoI9OMeXrQ/3V9my18bHmtAxyoeKNRrLbx9Gcy5kLiL9Ky
ojnsTgA97VcECZkmC40pqCw31Ee42N1iU8BSdSVw/HaTJFJHZWMbOHPpmJ06N8tL
qPvz4JTkr/yU25gSyyjW7fwP7v+pQDi7DynzZVeXzs4nv1tqZ5QvyM6vwa/CGNLM
18c8OBHza/9sj7/dFPi0GkczEpvqw6+JjZBbTQHt0AjUyaqjgdYDxoQaHETSX9/5
S4v1B2NFXiNaLq1bAxBmjg==
`pragma protect end_protected
