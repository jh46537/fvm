��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�`��L�o.�/?�߈��Ubԃ/����N���?%�\*B�Y�p��nf5Q[����jh�M;>����]�UĆu��a��ה��¾�	��N�>����g3�E�蔒�r�c��[���������z��&RH�@r$W�:�]�u��&�`�.P������D�=�(iX׈��c�W14�Ґt%V��:g[��|����=,�u�3�p[�J���X�E�]�(��ˍ�.�L5iw�Q�Jj`=�4��}c���+05��S1��%�r:t�Q>#FX�>'�����=��q-}�
��ӂU��樛�O��8���in��%>N���,⭙�ƫ���R�#�"���q�H̲�¸����ٚ �'#1��@3�Y��`��Řw\2�v��Eh�5�7�%��˰q?H�rT��X�9���H�@� e���{J�.�Dc�*��4t�l��U)~�eT�Ӕ��m4�B��4�f����F|���Y� �ȏ-�A�hB�|��� ����h��3�&BG�慨�X(�\(�=��z$�J�O��]ͨ�tſ�&�<.Ϩ��d���ʀ�2��������maK}���7��L�21i�P_���,�)��?�m�Z��3��6o��p��ڇ8T�-���s�Oa�ܾ�Q�qt�< ff_��`���Yy(�i Z%�6'�0c�ڽW�ّ����L�ZeZ̵��AͯW]�u���_(s��l��pɗ��] ��0[���W|'5���\�H��Xn��4� ű��X�`	Ը�[k�����\�x*��j(��T�ǉ�d�R�M%Bs��D֎s&{c���8�Ďi���y+�H��6lxv<�z�y�B�*�_�O��zѝ�67�����i��r�%~�A_�;�w�B(����'י�=���Ӧt}��2*��R����,JpO�'�$J@jO�1�w��,��G�p��°
;|R�0�DtE��nq�բ�rO������3i[|��B�v��~9�4�{ug����ZMj��tx%
��So����yî�?�Oz�:��Br�䎘�]%/I����]K32�4��g�����ˊN�N�Y�h��0�[���+>��F�%ގG�/�i���w�AM,L2ֆ�<�ܐ:�jg�Մ��<���w9e/'�s~��i��0K���vPd*m����j�Rj�3�^�+���L)�4~
+Y̻!~�T�����P&x�8��wB��V�ԇjv�����&��vm�Ë}����j�"�6Qo_�C�!�}���/L�����06�&g
?�j�K��D��'�H��A��'�|K��.�^R��^Êy��.7 ٪|�[��V�-��Md������Ԭ^�.-+/u����/7��B>p��\�<̤�NQTS�Ly�f�E��K�%15� L���#�o��ZS��В�kR�%����.��v+UU	ja�w1x�@��< G	O��q���`��=�c�91&����^��}G���'}���!j�E��������9&��]>C�,��NuU Y�|���p���<�̩}�={��+���1�#Tݔ�RT��C �7��.U�0	И����� )cv}�>\)��xq�W�9��"l ��	$��B~��+;7CDם
�k�C��,�5�)�C��/��K�{ɕ !ֳb^&Y�(�L�Hܦ8te��`S�:)��Y�Y�+� ��'c�ۏ�����xc����TaBA%�I���4=� ��ď5��[zD�q�	eI�H���3��/FQIoa+�˲E�;�.�zv'�l(��R^���J�qpߤ�
~�����o�Z�+�]B���w��Xg�#�ĭ�E%#��,w��=W\ҺMi����S�^A��f���Zɻ����D��>�*�Q���"�}YI�й�{�
�[yÓ���e�{��f�G���`ߔ�7�T<pp�ϝ>�jφBwD�e,�J��%�_9�s8�La�\8�> ��-�S���$HJDs��<�q��3dL��E"F�xj#(w��XW�24�+&� �G� }|�>ɚDg�LS$wUO���ܻ�u��C}�4�O���:G*5�:c�1e}iD��c�����bxR� sZΐz��Ԝ����L���II����\XV/ӜD�/�(h�4I��҂��'��{�����/�WcxС�"y�2~�oà��*6��/5��Eر��M���ٳSg��҅ԏ�2g����ɶ�t}s�jf��8R�0�3"��� �w6p��xL\��#!�H\fWk�2f��w�P\ ����.�9����&Xȇ/9���VS����<��u���X��F����ȁqW��.�[��3�L�:���6���閛�5�9"���t$}��X��8�Q;�S��k|��.`�$���5�����b�) \�*8�P
cy'Լ��۩���_��,�#���l[̽|bo0�2�6�(���H@{~��a�]p̲L�ǚp�c���%�� ��p�}��Q��B�扂�	�'ɄDLџ��_��=m|hcjI�\�#�X�ő��/�񉽙�[)�/ɁxyK��*EJ�lqD3p�9�)���'�o'ElΣ�B��P�Y=�r��,���c��ҩ�诃��]��3T
�����px��u��)9M2����A�I���ه�<� �u)�;��*��������*�~jk����r��(z�r#ʫ.�=�\7�����/�Q۶*