��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7]�s��^T��N݃a�O�BL��@pj�\t�]@b��_9hÊM��w���.&鑄w��u��Ɛ>٩H:v�d���5�3�
T\F���H��+MG�b,��1���fI%fV�N;�x(�Eq$֝{|��
3o�^�܀�ƾuj{v�J�T�
���H��"��V-Z�r'�y5�����W�4��h�,���3�5�=�6�����}�T$��n�b������1�o��/��t�V���As�l��|�|�Ci.�FtXS;B�ȸ���C�t�u�*�IS�C�v>��޷�B�GK��Pd�����;��� �GK�W���)4
��=s�A���# �x�1�5!.q�z�e]ߛ���9ؑ���kQ|����;V8���j���5�Ւ(%W�ܠ���8�r+��Q�� ����{B*w��>���~k����4(�����*��u'�C��P�Z��f���.���$J�b�@_������ )�%L�`���$���Z8��n�{S�����Tt:�xQG��ڒ~ߥ��V/i�n�8�Ю�oA� ̝]@����t�NX�wT�9�	�	ୋ � D�Ǹ R`ϡ�Qo$=�6oL�������a�.:�C�|��)*ȗG'�tXQ=�)LG�~ك���kJ�\�_�jJā�ݼ�hK��H�������]C��1d'3ح�\xvL��]R/%��C�`7v����Ը����G��?R�����ԫBG.)�I�{ E1����*�n�ot��s�F��|��� }Ijɳe�^Ci���`
����p�+ia�����l��)����`"�%�%��!'��'v�1�QWEݨ>ڷ(g!�_R��*��c�2��&lQ��,�}\x��K��,�U�����t��8�O����?�E�e@a���3��<<�Ƈ�`��)� �E�PՎfo��--��߇�8k����2n�B,����V��L����ԑ)l�8}�M�!S-nݟ�\|یPy�fVF ��$��-D��1��"@��7&Ur^&�QPf��V��lh�R�:��}E�������Hb�SR���/]�P�5�܁�w+ƥ�p��i�ƥj	Y2�W�D}'�q�8s����8kV�E?��6�S���c��,���#,
�8E:ozF�n�B�Hv<���9g�ڼ��C�����8�7���W��;�>�	>L��+W�F�W�$ޢ|��c5bG������%(ymtF��2���5k-,|=��Yft�EX3�Ȅ����~���m�ou� ڽO=~��m��?~�%g0�ǌ��)�>�:��3TG�Ձ�A��"Bg�L��P���1š��y<�֠
$�ht�'c�:�Ґ*ܒ\���D�@Z^�(n�\�Y`�Xe
�ܷJO�!��	l dè�qXp�K�{Í�߉��^��smJ2c�ҋy�������ѩ���4ܾ:�����H�.��VoKe��z8Yu�)�J�� ��&t&#�����j}�5�0�hد:
�T�8��nUu�uN�ΐ�1*N����`u86�����ʯ�⢙�����Rد���[E�w�ԡӈ����� �Ņ��_����~T�r~P����(�z��Ã`/=��)�&�.I)}��r0kJ��|1#@��x�|bUƽc�9\��`H�f�'rLK��R$��k)��s?2H5(���ਡ��ѐР���K�w��(�k��q�u�C��'iM�e�Pf9�+ah��3(���F�j� ��i���@���'����
��â��᧸u�q&�Q�;l��|�#;�E/�k4�b�)zп%��@)�m�K��K�t�:j�߉�dЧ���:��Ά�����W<��
�?*L�~�s��+h�-�sZ4m���V�]������|:1����.���v�F�+^�����V���%'�^��hq�6�'G��L\4��ZL�
�߃L��ō��Vb��T>�Z�t{ɞc\WϴerM�e`b�]��w�;re���!F%}~S��>�al"IZ;ύ/��T�մJ�oz�XfQ��G�Di-���X��) ��G��3�|阳t?9�;��fo�]�E+�|�S
�PU��s�	�7^ٍAyty��O|o�Q�I�ON�>�v�mJTAۻan�<�p`��B/L2.��:zKCy!7c��e���*w4:�Dt5\���놑!�ß����:��y��"g#�h&E���|و� �>� A��v��h���/c���E3�r���Ȳ��K�d�ifgM$��T(�h���Vq����gR�dڂ�)�����s�bO	��[�
�z��	���>��%%@<_g�`��d�8�|��,��=s"��5#`	��ӌD�VQ/h<��_��=dM
Nlr9�`;�?Y����t��1R������sk��	10�������S����m9,����i�6�u�rY����	m}ks^c,�GJ�:~H���O��Ѭ���{�Ƽ0/5T�oN����{�`!^�+�C�~�Og��F�ޢ#�Bk���]X���^2M��;� `��\���0�~� >b��%Dwv�W�JP�1�\v�E�ƃN���Q#���U��֬�C��	٤:Pz�:���O|v��2o�j/=��,@�9m�����_窺�W��+��1�a�F-T��4���$H��ș����w�%�2�/�
�f�)q-Ñ�Ěl�لG�qInj�B���SwƏb����9���X��S"S5,	�i�<���k �,�&���MF���{��F�E%������2�/ ��*�U1��Y7p�ˠ�A5��b��N���Al-qm�r��Q�:��$�d&�dY���a@�z�-�l�.c�`mE"�a�1���]�? Q�|zy�Ꮪ�}�	������YvC���JXA�"PG���]��e	�^���x��M�h*"aj�m?|�����&��`���l�4:Gd��|�L�]�"�Ȏ�Rի9,#�!T\Q�љ�]fcE��[�U�i��f�4�=�C���?U�Dj��`B=
|��eE��5 R���Kв�i �B=5��U��za;1K�=�|�`�%��ظ�(�>>ˑ��##|���*�攭b��������R��g�$�ZH��ir����P�|�,���l��ޅފ��ϑd%�vd����Ⱦ"ζhp��6����E� t�Y�(��BQ��,BP;��2S�6��G��'�=��D2����V��w{ci���(4-{d��d���嚕w(�'Z��Ӑ��C�y��c�R&�6Ұ�:���l�+gsY��"��]&��I�o�Y ����c��N�I����9�z5�DA-3���!oG�#XSs.�K�z+�N�탦{��&b���lz��~��:Ƌ��2�f	�#ȊqQx(�b�V�P���t���Z�k=І?���&5�V��k���`��N
�ƪ�ޢ�����W'�L�UI�=&9�A�����mI���j��c �&8��;?󓍘S�v�ˢ��ͅ"bL�z� Uu�)@3@-Ã2m�l'�I7rL�(�_IA�,A�E%<~��⩴��U���_KxIY�/�J�f����:zTU�-u�f�#� _�QZ�:E��L�w�n!� �Jy��x,��rA9���&��XNnp'77:��U�ѹڌqddԧ�X������/p>6#�j�	'\�$���V4jNe1�s-1�N���Vʺ���T����iCX��_��`������j'q9��hG�X-yY��Ş��q�)Cyd{88%��&S��u��%	���Q
�b*v���83�`/P�ۺ,,�-[n����S\�l��՛>i��C[N~P���m�Ȓ;J�9��W��E�f:V�Ā*���8QqK�ohU�b�t��� Վ^�rL�c�ɎIx�Bb��
����'B-]�4��W�X�O�QH�^36n'�A�3�9
ۆD�� �>)�2�\a����o�Bt�$�6|��n�$�',)8�z� V|;v�۪2(�t������*j'�]"}�/Q�XYBA{��t�Y�<�,U�ǯ~�s�O���q7=��>u uX�r�1Z3Z$k>����1{0�ҕ�)���Y�#{����y�y���`�M]X�G'Oy��QOE�K'w�;��4A��Xk�����ds�&���R�K�����R6S����6�ösKn�~�tCK})?���A$�j�ho��#���o ��驧*�ik�����>Ak#7r�@Nqj�� ��%Cs��6vDG�K&V��?Sg�҉����_ ���5<�u�`�����?��~Q��T�>�h$�N�J�^�lw���`X(N��w#�F��M��@�	�̨��L�NƸ��YS��)2G
�b�'?�.����`��>覐�Y���>~t���F&]d:��,4���_x��6�����~���2�@b"�jyy�.7d��2U�Ӻx
eH��[ݒ)�Ĕ���O3ߌ�Q�)v�,��
7��qg���C5g�s���K�/���iܞ�>g�ϖ��/������T�2�(r��yz��k/.tԟ�#R*�"��
��Tֹ�y@�!��������{h� VO�C�&���`%�$rB�\�x��cru���/%�T�`~e1�C
d��K���
��1�zڿ~�C��9Ik�a����ե(�T�.�A���x�آ��m�O�M�&j��Fy��lLh%�?78$�B}[-ݹj�
���v�o��b&:Yg��E��6��Hs��Wl1�+�D�
��J�nË�m���Aڣ;?)���'X����A4�]^�3��;������5�6�}��#�L�'"2qR,B�5A�.�:���,��K)�7�݇Y��lz���ĳ�&w�����vwFr7��l=R	D��F��sxC0/~��e������:�9JM߬�;�]u��l;u��{�*��7��Q?�׭)�[kw�!�eV�n�Cn�|�:�*W��g�1��<9��ψl�l�^48�&�][�M����������-���	t4�(!A��L ���z�ˮ#lZdr�&M�ԯ=T�ճDA��Y�CO4K�|_I���~p�V��;7ͳ0|����1,�rN�H��i��i�{�.8Z5W�U�C�u�b�ňz�c��B�.� �����T|L���\��bt�t�('�a� I��Г�Q�C}��,)�
�V�I�I�y�G+��]3��­��_��(�t�����~�p���Q�r��0��t�[&T	��y�