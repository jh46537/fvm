��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw�a�[W;���(���=�+V0�[&R�$E�J�4d��4�6{96T�9b��]�ž�>s$Z2�������QK��9NW�=�xIW��Q��x�)���ϝ��b�4�ŋP&�C�-l?�LM��4c��\��]%<8�r�����J�ƺ��6t�ݏH�\�m7i��G��~�5˗����4P��op/r�������"u+4�_J��dw��Fh�)tJl+Dk�4ȷ=��6|�U=��5d�j5 �NLK�8�O'5����eu��3:��.!U>\reu$a���'���b>�feW�ju2�i�)kE#�:������!�s��ƞfd��j�0beHp�9�&�4��^x�U$Q�2�,Wϔ;�]��5��Ѝ<���w�&I�jxK]U����(�H|,����S[�10���}V��izcLg�x�2}*�r����3��?Zs] aXPT�į7UZfC8wq���e�db(��7}m��&,�k�T��>rĪ�, d(�6�l�o�rk�l���?�Ő�O�7*���Xv�;�㚫�E�+�z��,����=A���b�ܴZ�Ic�q���H�v!H)
�5���q�8ZO�&r��1��E\|�>,�]�n:�ݽ�cAn/Ű�����{l[0+��� �[�����Y�S�vW�3'��� ,�w�̆�!d��Q��
�J��M1#(��.��`�����Ыwdg_�I������%C܆I��4%��^"��`����ҫ
�5��[�"�$+RV�#�:#]�²�y� ��벉��jgpX[���@���r�}^q>����IRm��K����D�1�C��"o1����L����!�8m���%h�]�1��K�����5�i�芨��hkK�x��_�����VNaҭ��;���_d�G�.��0�Đ�H2ET���L�4�	Ye�_�����2���IwH��;��y��O.`�l��fD�V�u�T�U,J��K�w����Ⱥ��๨9C�렑ϳ؞!���M£) Q�D��v�I�����ks�p��gR�9~%D$����_qgI@���v��ۘ���'�3���!�Au�L��$��wDV^���� ���H3�a��:�V[c����@��Q��w��� ��5ڽ=��<A�i 4s��l%�l�n!{G�4��Y" �M��n�Lb"��; �)��A
�]ވ�8��IL�Ri}f9�;let`r;o�\K��@�~�w��m;=�C���R�,u=�k���6T:L����>L�7,4@�ض�!Xj,Z+�b��ю�?�R��͋xskȵÞ�oA׍%$m~��A����o�8��i]I�3l��B7=�ލq�?i�*1�xE+�9�e�������L����t<�$�(F�Ů.`R�Px`\8�Uy�͈_���6��Ĺ��>�t��!j�m�[�;k��荱�;d5C%e^�P�����04 V�I8�����rcy�װ���է�y �����gkWs�b�:���#�J���h�!�t�t��رY5.���5_H��j�3�Tc��
k��Ʃ2���b�
�$zߑ��d#�7Z��T���'�8�֤�K���e>���t�5�zʧ,O�9�R!_�`�wyZR��6�2b��F�è��JnR�N,�qY����d�1�{��-�Sm9���ַ˽�73�t�3,��d�����#��hV���o��jeV��^�ȹ0�L$�e%�J��*�3C^E�t��WQ�K����P�@"��>F��;#���i��?0�3�?�(p��Qg�%��iGw!r=��vì��(�~B��f�ݿn��2J�{e�U�[�9�g�!c�YV�s�rz��9�v'�i��P&�~�t�<�Q��nDU�7b�'VL�+�
Ӣ�c�Ĩ��x^�F:�D[�)���@�F 0�_ � �@ܑC��M���~�E�����ļ�����_Ee�U:����o1!��6����� �ۅ�U}��@ 8����HCC`�?��� �Yl�mF T!�vm��1Dh�o y<x�m���m�6O�}�U8�|C����xZ��2���RB-���+��h.��� �(K��3�\��%'���n�.�bd8�����w���_ʑ�W�k�b6�SS���6�O��؄��c��0k�b0( ���I(:�-���\�Rd����G���kW�����.���\$�k��	O��[7K��m�� h
��&�6l����n~_m�g�Ņ��N��(3�������CP	ֽ�����ܶ(��#��|ެv߭u�CⳎ[D���Y�X�Ia ?��,��Y�/�|H/!�]K�ӿ;!�%Su�,Tːv�
	�P�o-��n֘�����������?1�ը30��wG�%�J��K[�?�xi��z���,I�E�#�*�:���qn%����;��� ������>���U*\A=KT�`����)|��+m�:D��������'�u���2��=�R���>�v���S�9�P	�/OU�����4�{��������d^�N$�P���r����2�;ô��c'C���m?	 ~_�Ք T�e*7F�,=tl�r^^�K٬��y�� -mP�y����}�7>���u���"����U��d����V7���G�)	��
9[~��a�Mɴ�Rd�.�#��-p���J����^�6�?^��b��6U�� ��[ӟ���.c\�N��M�\̉>����Ǳ\p�]t�č�z���J���G�N��ܟ	6)묯��"�T0���5�b���dd�!����д W�׹l��R#���6�<�
r�C�Xw���AYx�m�^�m+�Wd �Ӏ��*�-�˼l}ǌdV�v4��1�	��~=T�~��'r�Z��^]	��`���Յ�I�s�׃/��I� O!>����~����G4�������61/g���58�X͘�V[�"L��ѿD�4:}�٪�����2t������ ���ǘO�c�������ю���ou6[p�*��[N�i�X�S�@���SƨV��	���]�Y�d��3�ZB%%��Ȓ�' a�7�ԡ�ɧ4[����`���n�
/�5���T�\���ǥR7�9�n��kY}����u�g����i��5%��0�'��Z���<4�0.�TA~U�>���az��&����y�"6~nf���:dCpF^�����BX\�I:�+7m-p�����l�����!��vҬ.��X�^�0����o��>@���P�r(��`��v*��qh��7��Y �=%�B��1֣��7���Z?�٤�xs��M�Y�I���a�Y�<�I���#��Xd���,f��R��'�)�ƻ�4n�%=7��.LI�kP���P��V�!�ݬv:��IO'��W	-�i�Vo3�t?U�C �;��|�c1�^1�>�����
m�M��[j�&E�'�NG����	:��I��S���DV{�6�q��!O��O�suD�:�Sk����_׭C�MO�S�N�� )��o=���&����2f������H���a�@�h���X���hhd�B*��3�`�� �R���������r(�">�Ͽ�߇7�ҷZ����i�h޻�^%oig�^��^�"[#H�M}�+D{i���E�q��<(p�A�8y7�
���J5�4fs�Ư��A�t�H>b����{-�Z�؛�[�U3"��6Ϥ8L" ��v�����W�˳%=��75����U������nF�fp�j>4��>
�o��I?����K���n���T���2��r�U�m�q�jL�7�;\� ��|퐾�]v�τm/\����9"I�5��,z�H	�gr4�)�-� 1
����3S�"�?��
�/~��FRHs፪�D�JL��T q���ō�k�#�O��q� k]����3����dL7[zE֯�S*�>nq��O,H�h��x�������s۷��CH��Y�%W[h$�Ӗ��8Q�h@yB��+~83?D�|k#�~댊�E��=?�t�wdD�[��0��(<����.Ă8;��@Vn:�B�7٢�8C��Z�qS���H���:3���M�U5&xr�`JwW���آ`Oţ8���v��%�E��<�,0�D�<G��0�Ap��<2�	Y��p����a����΁�s٪�MY{W��YĴ��/���YE�'����%p<��ϴ�Sٳ�,R�e��Q�<>U