��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""���᤬����[���%rҦ?��*3
�cӂJ3�l��k';pU8��+l�{�!#���Q���D�v��i�D��5���,zi��<H����uRBu zؼ��`�;.��16�W��\��ƚF�8o�~Q)��c�����`�s�А�����j��EXD޸�F�2.�#�,�P��f�߇~�1��.q+\HNF���t�χ����8�8����0MG��/���~M���5D�7bz5��LR7N	JcF�q�?q{�*�c�W臬������)��-�;�Kf�Z�������p��R/�5��C0�����lIXT}�\ޏ����!�dٹ}C48���6-�(7-ޱ1�_.55q��b+��6�V�x�?b�&�*^	 
�x��tk����bbOD,��G�
J}:➙�	�i`ֺ`����Xp��/������Ѡ �Ȃ��OlA7��ʐ�����Cr��� <4UŇ�!�z����|�mٷ��Ӣʆ�ՠ�Z�.HjFX4ړ�TesD<��ٔ��\�
	��6��q����e~��i����`�Js2�n������gd�4LW�g��9
2%�e�h��ܛ���B�Joh+Ḛ��ⰐMb�k_Ι:���%8$ۼ+3��q%��k�ʅ�����Z<"#��ϊ��|�I�ya<�Y�0s3��gr!\����):��o]���8H|�x�:k��F�W�>�~�2��ڤ]���& ����]B0��9G�|� 8�)�'D��_b�|	9R�ب����4|���Jua�8[W��,%���Ie@�#,N���{����-P+�?g��	b��P��#�(�,�_k{n�#Rw�ow�qׄZdH�K�s�"�~d�YG����-��k���=�Lg���.$a����괛��<#�p����GO�2$;
(��<�:gd��}z)S����B��󆮍��y6^T��9E`�)�,�<�jy�A�T$/�U��ɕFy<t*>g���jz*��6k�F�r�}4�`�tH��Evc��Le�[in�>��H�N~�w%0���I?�B��h��!��JZ��y]Ie�� ���f�L�+�XJ�i����Z�mf)�1\ ۑB��&+��`�=��g��>�wQp(�H����OUTT��1,�kS�=��S:����h�4��o���/vk̆p�x"�펬3b.(�̫��	��%_Bb��-��7�J��i"i����@Aq狍|4�oL��ǂ��S#�_=�}O����E��*�6��M�(�oA\9���:Э�e�sd�7���=�=.�`Vʪ�}մ]�"/ѣr��&+����1��i�n~���}���Ѻ������5�*���s��x���@It��ű��>ZTX�Q?�i���a�� ��M��Lp�VU2���7tt&�;�$��U��'�FV���T?{o���.'}P=e�����PC�:9�~�g��awn�k��Uf�	��7VS|>Dd�Mr�#��o�&�}��
;m���(���~c�(����t��v����A7m�>*^�|/���#=*��B֬���u��=��m�����4e��@��e��Y����b��ha�g���I��TW�5;b�^5e}�>��ġ1�H���ϰ��;�W�_��x��'��Tw��Wd� *5Vc��q�w/�>11!�4Ï��@�cn(n���:��^[z�ؖH	Y�P$GCWN���2�6@y|�D��ʚS�X'���0��ƾ���tK���� *e�a&^�<�QQ���cp�|U�KP
��v��Kp�g�j�7�����W���Pຕ�c� ��ӵ�#�~-�k�0��������|?���CVX �w[*�����u�jqe@�s%7�~��Нˤ��V]>�* ����SJ�ރ�t"	l�p��g�ډ�Ɂ��X���bC���J�x�[�D&{�"������JbYa��$Tp��@_�82�� iG��m4�lg�Y;�#;�������,��VQA� Ӽ�ɊD�1)�d��m�߅|4�4��s?��Ј0?������|7����;�O�m�	�I ��
IE74s�y����X"��Y����d��EMp�Km�5�ö���~ع�5q]O���>��!$�c���1���.�7��g2����g�Mq]T��R<�$�j���'�wDΑ��I��SC��e���w�[Zj������i�-�O�9 	$�r�dl��G�"Ѹ���)�0C�&"V�v���ʼQ܊����?�����[E	T�h��=p,	t�ˍe?�1����yP����,�jUm=`��:�1�T�+w�Ú	�H2���^��h����.s|���
�>Nm��������('�V�tD�Dn�5T��s�IR.F��-���7,��^�P� >&j>Lm�gY{'G����dͯN��^.M͡C����=��n~��ip���9k!��x>h���
E[B=��k�{�������s
z}�ލ��c���\�O���v��K0��C?%�����F7�}K��:N�����K��U4tJ���[����2Q#��{>~(+cչ�f���g��|O��cױ�]&�ZB��L�9���.~K����)��2cY��e�Q�c5�H���N���Q�"��+�!��3��_xg ��N!(��E5 ;)�iĴZ��D'���W�YTD�(�\�n��*W�>���%x+�U|Ac���V��b�ݯ������H�}K�,��2';��Z��~!����Df�"�K�LNy������+H���.�C,����]��l��H�ԕI��~j��L�@J���'��l�WA��0����@�c����`,2g����|��v�-�T}��Z�F�X+��r�o��U.=24�@��Hn�Y���T��|=�S!�]q�Dd>��s���m������r��5Ss����l _�Z�W��hr��3���ӱM{Uv�?��_	ܾ�D�J�8���Z�/4(�w�7�Ir���Y��o����q'A�"u�	=uodE��#:><,,6UlZ�d���������}íz����f�T��C�,�>*�
�S��<�J�o�q"P�{ ��-�j���3��)d�m��rl1�Eo��0չj�⇧��x�&Wj���>Y�)؇����+/�[G�h��n�
�����Lt1}��r�(�������}��L�I��B��"�M%2'�����$E�
��p��FřX���K'eh��.Ղ��C�֯޸�0pK��/4�Ĭ�Q�5b;4���}��2��J�o����<N�+�}%��rp�J���u>%�H~���lMVZѾa�(��T��r�/����xNV���E�<yj��JfW�$&��ZM	�/��h��>(ɄA%�@:V�V t���VG�w\&UP�P���@������w�P�la�;O[�Q{��ц}q�D<L�;�x�k�VM�{��ìeD��
����Deg?#~k���1c/p��6D���j��ܜx�,��I������q��A�h#�i' ;5��ն��c�M�`mj��F�3.���R���`D�)�P!Dۿ�Z5B6�c���r��^��Ș�����g==��Pg8x��SS	6���[ų����j7\��#PBz���c�D����E���o`[V��#���s�uT��`L�9�F!�.��`�ͪ+G��&���6^�Hk�J����n��l���3}Uv7�G�j�f]��g��� �qX��?O����ۂ����gx��O[T�_�p����ID��X�i?��
ǝ�b5�]�����*��F�i�U�J�	����
�~��D-��uX��(�$���r��u�q�FU��9W��N�0"�\���K������]��4��*$�1l��ZDJ�#�K6����sݒ0Zr��`�AVQ�4��@`n�rV�v�R(oj�܇��
0f�J+F�DJ�}�@
v�^k�Ӽ>�ĵ��9�n�]�<Q'�����e�Ԧ5��h*��"*��FYE���2d_��ҐcF�"X0��r�|�	;�'�W�~���UC��"��gb��W����� �v�!T������u��
tc�����A&xi0�����.��piqN��a�f]Ưi���i� �h3HH(� �Ȓp����ʒ F�cl�B��ٙ)<S�6CGԁ�c�M����9�F����i)� s�/�����nA�χ���e몆����r��$��1����F.Z1��;�Q��,)"�7yEg	P�Z�7�MuV�m?������=Ӳ�mU��(K�IdweO���b%Tr�H+�%2���@$&�(��1�f���A+���-�I6o�6VW	2���_�'�i��X�/�%,m�M����<@��<^c1U����p�I�&������9�o"2�����+w�E���-�ͱ��ڏ����}�K񑅊X�� ��ru��ga*5^�����t36&r�����Jlh��Q�e+�z�|���'����H|0� N#�̇��� �|���k�H��"�E�xҩ����N�B�HB0߭j����#v;�^��/&cO����Ĵ6�.(��CRۈ6�1�O����/�wyИq~�$8�
X��&a=�~���N�4y���'���h�{|��sZ����W�Q��\Q�x3�;A ���?	lP���-gZ�T���W0�[hjV��T��lDT˹�╊	��R��������)�n���N�[S+�~;�
L��Px����rq���A�Ԇ
w���}YK9���G#���0��9d�����f2�)��s�t/	R��kxFt%��0nr�8�EL��w�!@��\���&��vʺ��d|M��ZQA�I"+�����/�/kB��F�q�5��OJ�K����{�a�)M�f���1v�A3[;r�����&!ڰ���_�9[�zud�UFIg����\bd�I�^���LP�պ�F���J��Sឭ��)��Qy ��ڨT�d���E»���U��\��*h�P�i�yH�fs��N��w��b�n�h�����ib�kRٯ���o�{`��x�6o`=[x��OQr�^�C]Um�����Zc���!�8"k0b�LO��(��g����l�?�/݃���~Ro�m���j�S�b\�u��>�X�*�1�DV�E1<8c���EJi:r�U�~dlb�W4:u�����Pq�L��-����b��8�%v��>n25b�+�g=�u��l�~'���'<�^�v}c׬$�����5���k�ͧE�����b4��kP/�8�9�������=�N�NO^e�"����AaiW&�B�-�\�kY3����]�s����x*A�絔U�Б�f@��*�WZUR�ĉCh�TjH�}(��<��3$`1㯮����5a��(8$�#E��2�C�1���l�c5��%��G�4���3˸����|K�|
��EL= 
|���4��|��LnW�3�<}���L��} �#i,�z������{��6�B�:ɲ� ����#սw�rC�!�O�b�����6-5{�ǵ�!�g�Lp���Ȥ	�r���v.�3��YP~�3�/ﴝTJZ��X�/Wԑ_Xy�P�OKr�����L<�����%.v}pҭ�cƟ��(���/q�Vr����lI�kU�Q�1��/�X%��o⮴��yt��S�Gr���9��H�3C<6=n��頫�!��Ϛ���綾2A+�Yt�#��FA�Ir	B�xZe�7	z8�FcB�b���"D&K^���I!����O�A"Oy�>�]��j��۪�}�|�}��w�S7��<iC��}g�'e��,��!��6���qc�>�J"�8��3�Yw��ya��^���#R� �%����)Sk�bѮB<��1�����h���ɪD8��	�r_�BH�Z��O��Q�-4�"�]���^gMB1�f���at��)'k!�N^�K��,6G}�Ґ�K�N�F��ٴX�1�H�`�sT뵳�y"��Ȣ�: ����ö�RX�|�=j:(��Nq���J-�C˃�I��-���?���I��x5�U�1�"�$���B�lq�N,|�3c��M����ū- ���������hZ{1}��6��i��R�0��U+?'�VT���w
�e�� �T=����%�$�,�ϛ���Z��'[wZ(�6�M�/Ȉ� 2Ͼ�\R�����y� ������
*��������rr��4!��,����t�l�B�IgF���RؑqW�`��׽�u����g���������#����7��+n�ڒ�:2m���B��;gp���6��s��S��Q&MI3\Ǟ���b ]�����;�[��&@����눞��&C�:��#��J�׾���z�&?�$ׇc� /DT��a�>����x1,����L������vP��v������RR��t���F�� �_I�nݕS#���V�2.9��S�h������+ɲ�]}�W����3�d$���Pm�$��FK���yk������WPY��&�;�`����y%��}uɜ&)"4B� p�?��/��`���7��}_v�%Q��k���"��%z��������y�l�/��i;�6�R[�X^.��$ǾA�@Џ��)�nչNIFr"|�����_���5%kc�/�PD�þkL:��t�+��.��a6<\p�)�q؇�W��x�ޱSzu<��fR.V&����@�Z���c���R��ťA��>��Q�R6��0��n2 m��y� <q��gttr����W��~k�\�1)FSϥ3�|��䌕_gț�\��=K�����p�0�����F�\�.N��M�=��/���S׭���M�k�����t���^������c���� :7G=B�5d�����c��7� �[0�V
hO¼��a������bd���=!�H-'N�<�DfC.E�n5Q|�`������jkQ�]Ӳ��=��IU�(_7V�?]�A؁6��}N0?�����"ǟs+h7F����	n@���?b�
'_HO!��/o�ٺ�d(8�����g��u��?�5p�pu��zkא�g�T��K�afΙ��������ܤ���WY8"a��X}"�~ދ��-Vv��r1Z�+?� ����b^�-��x�7h~�#j�B�����N��pq�n��$�W������IbB��4%Î�����gp�	H�bC_i/]���I۝��-����y�L����Pc�e\J��FB�oq�����ŭ�/��4KU�@�orS%�b�m?�5j�R�3
fHq�2�nFV=������d^�BF9�Yg��~����w�(��z�;��m��Q�;�e#����*���յl�0��@�[��+��/�<W��×���� ��x~2�~�L�>�p��5�e����h�R����X��s���)x���s�Ay6`*\?��O��EK��g�@-&�Q�J=�����y�B���Վ�ߊ(�Nӂ�]R׭���kDN� #W��06�^�ֳ��Z͇�(����"R�g2�����d�C͐������R��{�'��hp�kH�����A5c\�qfی���8Q}�W���^� 2������@H|ގ���Z^���W_]�d�pnHݩ�[�a��.��}s��_S����R�h�X�_-��9�v�VN�3�<�d4dt�tgg���'T�؇I\n�%-H�T��E�u}��RvQ9G�M9�7���1,��hgv偉���օ��H�0x��_������^"��x���[s�Gx�H�9ؼ�Zu�T����q�������8,��SOLCp�g���N�͒��>�lN��a��~w9ΑE��X�-��e�u�]��0e��Pg�0����2���U�C���0�te��&ݺ�����Ԍ�;^�&�3y���+x���u��12Q�<�Y�1�H��S`�y��g�Ɲ�qiX���w���>d�}7���&���P���Ҭޫ���-��7L�e�+ܒ�,�1�" ,Ak����7�b�D-�\�,L%z���1Q�+���Ati?�RpK?d���6.�#<�cX��f���t)�d�:��~�+ a�7#[x%�l��jR61/ƌ� ��-H��yH�7�Ѱ�9-E�m@�EX; �Dt�l_#�`�w�����0�Ģm�\c&O�i����B"Zg���8V ج�u���VRR�5�'ѷ'����miO%�}�g$p��{��HRѴH���-��"MV��;�������[�`&S�m�?��vT��Sf�V�l6���k�p6s-�Ao*H\��������b�qx��;�?Mj�.�f�{�<�ve�O
@��j�����U�x+�?���\�6���KM�U6VX���y4%�=��Aok��2q�	W��?ǋ���JY�W7����$y�寗@�0~-� I�f��B).["{�.>w��|W��S����}иhCS�k���h�����@�A��Z�a��іӭ]��9d��뜹i���o1�o�/-�����?V����_1�\#���h�<q��R�$����=$x Mp��G��69���ѿ�~�U ��~��f�d�n>�W@�v^��_��ٝ��7,�w��Ŕ��??.�˽�Eq� �a��=}��� U3���C
�k[�7?ft�=1 &J�m�T�]����0�8G�A9�ũD |��4�Z"���O(\%wc�i�Ch�F�R`�	5��ài��uĄ���\�ֳ
��םJ��`�K���ʏ�߸�2s@F�@���G�"s�+�ǋC3yb�YZe[��et���W�H�y�
{�pb]�ö�I�n���z�f�g��@*�a����nbY�CqT8H5����nf�zqQ˨�FBl�,����wk)գ����?
 ®$9rҸ�����kB�b��aG��a��%
������q�ݤ*�B��Ĳ�[K�zI���ҳ	����B���3~X���nm-�\\�x�>�vt�d,"c��|nt�d�Q6�l��]\�"Aus������Swڥ.���ҁ��	��	r�d-Lxk>����_6P�&�ߴ��E�����CW&L���Y1N�nρ1	!V�0�\R���2!8� �A�����[�����Mig�m��ܒ���y
3ۘs���|܅��#)�YZڬ����Ԅ����n�u�Hf�|�:�L�[.̹8�C&�Z��.zA�	O��:��'��7U~-=G�=�g�K}������	6�P��_-��
t�j��a\��"L��k�Bʄ�9,U���+!�Z,���c5�m(�7q{�e��I��a)y��ylcؕ\יؽ�Ls�_�ȭ�E�#�Ϧ�݌C)��I ���o� c�~72!(mGN����!I=�Ö��Q<HaO��N�09-�L6p0(���bT�N��������C����3ʂ��|��6�X1�a|��6�m���3�V�[��}���
�x����y}v�].� ��T���<k�ܵ�E|�-�jǭ�
*+���6�-��j��'��g�;M:y�5z���Q�h��A�~v��͞g��l��gs�P�#ԅ�Ef����e��q��D�,�V��le���[��f]e�I�S�ztΘ�%�[�G���i�uز�@�����ﹼ��/�R����v�@i���S�!,<S2���?KNX�`vQ�����Nd=e���k�k�P��MN\:#w��U�G�e[��g��+��L�O#p��#�}����Z��8�w,I�Q��a��<�w|����,��USGρ��E��*�ײ�;����籶�u���e18�1�+>�
+�Y�z�xb�vE����IAhҷw2J�e~x �o\�� �豑���Q�qB�#�r�G�УƳ7����qv �T���M Lހ��E�d��(1ۯ�Y��ث�� �C��ie�Hy����D>\G���������d��*+���| �4���C��?�ņ�����*�_�_�#�>Љ��H�wv*Q2�pH^M��B���}
y�Z�w^�u�6�T���^�|�^�\������SMB��߁А(��4k��r��O-k{~�Z����)�|5��Eg{m�xھS���NΫN���v)�́��+���Cp���Q�c�m�7�ؐh�/O6X����_��M��x5�qͶIU�<|�1=�I��1�Q�JM�Ƅ��C�d�*͑��?6 ��+Č��KI)�a:RӀ�����"@�0m�
Bo��@`Ǵ��,6�W&O��@���6)��8|��S�ŘD�p�x�, ѿS��,��v*]`܌�������*I��*�5t�h���Y�՘�B~��bj �q��Yz�ЄݒKz��>Cp����6	�eL���,X����'*�;Kn\Df�~6����l�������Y?ÉniA;�祦	��X�%����|ݭ�W��v����=?' �s���b�fX1��DGu���->�q)��4����Z��V�}��V^.�̻U��>�/�o���&��MJF�C,IBf�j>��@>ۿ�W��#%}���;6�$B��N��j1�Q`�/^Ԯ~��>	���ԭ)��|�}n�Rۙ{�_$u8�g��q)�p�`�W^7�>�O����S"( ǔ[W�`<EM�����m��G�3OI)5���b���]�T���v� �]��g�����Y�l�B�-�겺1��`�k��ŪR1}�W��FiȲ\"�/�V�>�5� ��;z4=� ��ج�(��t�g?k��d�<�����C@Nb>�r�dU"�D�>� V�E�O��^��a�=�d/I�KÊ�LO�L�p[�7u�4��2P�:�2k�o��d��b1D0)�s��1���t�8���^nɁ<���x[�X����`�+,s��»�H�����imI�Ǽ��f�xR�tBs��*��L���z3�an2=�mSs��&U2�b��Fb'�_[s�E�g����w=P4��SQ�|�ˤ�|pSꊭ�爈��1iq�b_��㻬���L���*Y�����;P�i�����б��(��%[��:]�G�<様3������Ռ�H�V~�q �G;�qT�I�z�K��Mio��Z�XV�_��bߥ��H�R�B=ϖK,QA��ٕ2�2��}����b��,�K�(�A���f�=�ec��V�t��'=п1�N�>/]Q��:��C�{Mx�:?�Vk��	g|I'���x|@�(�z�/2��Lg<i���7���
�c�I�N���U��T�2� DZ(��mS�O�$=���E����a�6v���<?�����3a�h$�]-'���ǋ�)HV=�C��
�L�xYN�`�'Ԟm`��kpJ4@+԰
�j���E9ʢ �k��+�@��H�X�+Kf�ZgnO��	-���v�:=�3����:�:{��iZ�e�Q�hD��[Zf뱀q'li���"��nO���羊�̛���.�߶l&����@��}v������;��7|���V��_����|<��>�mŏ��v1������q�����sS�~�Vϟ�-�ۦc��\�7f��^�L8�{Q`F�I@�Z��E�18��Q�E	�-i7[���/m%_�}��^��qF�����</h�UN����N�g���X$c�i75�\c�gv@^p<�|Z��[q�����If�=Z.8�Yh��=�$W�^�:Ѿ�MP��橸�טv٩���?����0��L����?����Ԯ��jIu!��#)L��>��S���`[�E�X@fÙ�.ym3"��\o\���T�k���������3a�hf�&+��c�n����ͷ=��������.I(�f�t5�g�a���k�����eBC7�e���X@�t���`@�iDՈ�d6Ry=ٿ&Ꟊi�t�+�_��y����ȚB�@꿖%�?����P����;O��WM��ȍ�&N҆lb�*o������t��v�K���Y�iPGuĵ0�2)�u�w{�������c���
�5Ib��1�s��i�!��q��3}���S��B��tz_��w���d���"�n���8��
�zP۰�~�X�����І�����]���� u����]돷[|iJ3=\�#�g�,-�~d�&����8�(I��GN�_���*�����ɒZҧ���uo��X�ëtOo�*��M5�m��$�K�sY��� �RZ`fJ+�"�RAr�-�9�~��1~�z��!/h����u;'����^�ڨi#u3��ˆ���}}�D�;+��)�f�����9��1<U�$H-���M���f���E/��
>�x�E���oo!µ�UC��<ϟ�g|��|P��k*�d��	�+�F���G!�p�U V<F=�K��*?� ��-�c5K<��{跅"�9r�^ȸ�� ��� ���$&��`A۪l�Q��%��HI�n'
�yվ�\�n���p���B���(�7�J����Ɩ�N(����w��r�@7V푤�]��9I�
�Dn��7xGc�!<����F�s���X����C��
X��?w��W��AՑm`��K�O�f�1�Ü{p�Zܻ�k�/D�Wr�����n������u��rށ�F����(HIL����L�="�Fn����zm� O�;�R�O=�Z+�����\H�H��?���D 2��=�R{=��]�/Q��xL�"@�����k���yK��0