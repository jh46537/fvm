// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gsdoynqWzHpThcxPmJsg93ela2ByhzbJ1/d4/AY0k7qEHSZECaVNWzwJ1MGSul93
DPJmWFpsmTgjXCMmfnZH2sL1XfAmhvhgfCnpH21QBZIs0THIxKa3viovONVBEf23
j4s006LhI75z1fWDh2uEFKunr0PGkNOfoSLHxmLb++8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19808)
Y7yeUmSveH7/F69+OS6/Q+ZLLKd2UVcHcunUvAfW+bmf7ZpuD9lbaj15O+vOq8rH
hT4ZlyCSDF/bW2JCEnic1q7H1JUBjjj5CaswG8Ka+0FEj27xXfSd5jCIy3ur7G6s
rsjmZ6xR9ZNdDvDCnAB/EcbX/y5LQoxnzmjSGkI9Cegyr//V+VtylPV25CfjQlxP
oz1wGwNsjlYXooT10LcTQdjrbMQWYNjEdieYAa4FLRUX5cDhwf1BVVW+0X8fX9T7
UwTUDLLp0B8YEo7mI/ARxthewE5XVF/w8UPaFTkYbG/6gwcHJyQxFYfSM/Zz0Glj
mk1SI+lBHFv1JBoizDrk5/lgZBT6Uz08/Aa26ZMhmUMFJWqZAUL453QWzyefQFvB
o6bqzMhfmw+3XZghNUqz+o17i4erCf0SpyIEn9lo6hgOfHJ7IECJfAthp1k0KfUM
0xNZ9NqcRFMB85fMqKLIhIKNtz+YgHvCAKONy3z0/OLUpn114aFcMRltBTv+T6Rn
GASH5kvsQH1kZLRLWcpp0TMk7g2y+mPj/gGm+J058w3MH9Lnjj8JJHsmxp9EPiA3
cTglMLMzS0yU/505oCzTCKEb25VDjY3zLaBHFNiewyvjncVWy/UxQCs3MU7+JR5A
DipizlzmIB32Hm7u2XIuENwZwurgNV92RDz7vAEoEuCx9FKNit9wNouHDdUrEz9f
d/kVy1sAXf6lYAW2P4ZT/uZreZJ6BQWBvziOduomW2O9Dq9m0K6HgJOCQbvm0fZq
VXabsAcAJvS4GzxxM3NsJwnI2D3Khcj1Ya3C5bnIJTBBHYaBHdKrEo4OCrqwyQoF
xYjOWBQb4UdEiRPWCntg1dMieguRpLwOKIQBnQxW4tQ+ocWtFSDUKSAP6uPDYcnp
hLWfplQDxB7aH7XHWx57tCUXUVAonUCYwzRR9EwGn5JZaFotq8dhdcQp8ZDjMDC9
h509Pn1HxvzUZibQqgsTYQDhNe7v7ZSzUd8JPY3OveUxNG4J42CIaiosA7iMyWgQ
hD03k1wJCnQr/oTfaSLHTOB6ajWpD+pADzSVY4cg+i8gIHbnBTc2ziMB99FHITlH
Gzkr89umr7Oy7smjN/KgHb3GFXrKIrR3Nr8lHk6puQr07AEqOhY+hCmQFX++r+Wf
2J+tgYAHvPhykMsYQbxmMa/VBIMPNrfNQ8LjSOG2ggMhh+dkDsqqNVjVBKBLaxR6
/BnJtnd/E/Y16/NdAZkqrhax6xdif2OvO6DIS7qN6DVsh+TnGEEw/VX2eJ+nNFgx
AsWfpw2mDwTiNtW3sotsWKKjdqt1u0PY5OIogfOBOv7XLcg2y/1ffy9KPtKN2Fid
aotv6y9TW0Y/rzx36eWC3e2h2gGXa4lbGcmUJGcGYSWHUSi61FWf68yLxHOBD6l0
6nx70c4Xxl9/U5mWL0X7wiW6z0o+5PbcJaVlk0V61XbEzXD+zMPpP4A29DC8RLee
J3c0qkAlEgwJNYxjR73OiPBopSkb7nLOCXl4mbceX7LpNYeUODppjQLG1p9olnqt
+s27tZCJPOOLPS3oqBGbqZjtCRiW41gw1EvEaqahYI6xquCJwtneHvjUUiBVcAVg
qcQ2YdhlQzukOi4szTur8+5y+2yeHoox3ixSCulgspPKW56KgzKz2r0I9EvgbfHw
5SzTWDbE6UwSJYoFhThzXCk0z3ECpGclJc3NNaX79jwl5aIOeBrUriOHV4QVVzFu
hhGhXlyi+OFcXqYmNIO1LNeoZhFXWdWBDHKTBvtTyv3RNqHfW3LHYVGyJ6SmbyVW
F/RyhPt58n5Ep/TZj5HGlYCJkIDt5Vezc5vkVScmAY+jXcGphiCnhWLi1KW8iTjJ
hWuMz9m4y94S5gmgS0wYwh4Zj0Q4ZABd8Kejf9wh+kibSP9tQsKl5gAdEoTcEesI
q5/OblGbVvi230qYTvBrItG8RC57s+wT7fKfo/09pYbMZlOVqA0zCI9x4PAtO8Mk
IJKpkEImnGY3HW9Avl7Etmt61LzFimeG7q4HD9AUt/4iC1K4RmQW+UQs/2PPlCPu
t4waG6RKw+E8xw4yclxjLXKbN93iocjkodt94mEe3R4c1AE+YazV1AHfvcV/5E54
XBq3L3wAhBed8VfQibxT8f0mT7trmZgJCfl1cVtnt4axM3q0bkfbiAEHMffJdeWm
YX2bSJx0h4I0R9AFvttM2Hy1xNUVt84ed3CBGbogJE/+5d1DVmT8q3ey33cDqJT2
ouKHMBZnW7XRffn4/4Tl1QIFNjFSVfLmukTPPUaHMQ7Q2vw1sn5VAbN1GPMNQcgP
bqyIyU3if0Rdz/MjzwEjtS+Ac1UwKIyI0mZWITbthMHFjIC6Vg+ouo9NAS/WgxxD
aPHCcnuCzWKEebTAiYHwEoucnctDkCNQRdfbNbZfYj2egz0MaVJgsnxCdD1VPww9
95+511mXeX84b7HU34e4BMWMKz7hBlcDejbtQETuMDKOiASOaTQNJytulBUbYIwH
Bp/tfCngiqlaidCEX/NUGBe5wmGGdffmJqkJ8+eqzfFRi85H/c1v3tQOuIyhrMPE
ds2BZ45aPKcOgqgKgHgSTrIYL1yAFKp1gR3co5OIzQJCuMJO6s8jGBGPRK9F2H5q
SV+GQbxnVjXGpjKyLYNkvpIpCSYXZh2QEudeCjZL46iCAqTGgZq+bYYaTO52N/B4
okqnJ/SAcBGddqwRoieFDdwD3geWiWHJxyrduTZvOYuiKXx9Sqdwi0e/aEuqSaaE
kT33XS2dyvoHQxmy0Q/jtxCfQ6+1EXgs0GKnOXxndK8tENjV7LUojM2CJV/C/CxJ
ATtqDXz638nPE94iMG1bxxcvtbhCCQU3BYS0upfetQvqulvVMjDTAg7GeJVipbcs
31ciPNZiIJdglYIMDVb2x5W3XdcrQQNTOy2tm63w3caP4AHSBGt5ID0Ff5YBSnTn
vCtXX1Jb92yfqX9QjvOlSSx8/jUIo/xfLuNe1cVDGIffcV6NuilcrPCGKzupJMF5
gMxB+tezCtyUSrRvFQGrdbuTevwRKhgTy+ovqhZGprnbpwfhBEgXfA056u8p0pBv
eFP38nQ4J1ERecqRN51AaKvZXrSQ53oUZPqkoj+jyeqKhOc0PtBjb5nD2wdMqsqq
lQKH7YWJmruBDuWP2L0IyCySaHCvpmV6qMDObo8B/snT51MPufbLRxMEhginyCnM
+EcY+eEaBWcz9eSHwtz13Dvf8fWCybOU1vHWztR3D35N4YYbDVTZDH4xyVNJaWyd
GVoaGQ12SAumZHKvU0G/DNeHwadiuMt06vhuA6Q52jUNuSTOVI1EB2Ut+6gWDCGR
Go9ShSoO6p5ULQhcvqodoOD/wE2UI7Fn4Lxd20KNUBvV4sjb4Xp/+kFjFlBtwJ/Y
18o3dIdlzCmcJXri0ABZPlCvuoPTHBMbXA2DyM2GaxTta1XTOhL/nU7VIEuHwthM
YQvyDT1pE1dEbEsaNYSVwDksreT5EwpbLiVKt7wnUxkoFQ+xwxlXlN5cf073edYR
y3JgdhQWD97Rv/a9s8Y9iKjCgRl8yXk9M+VLE0rgFEZxr70XRdtL3nfK8dx8VSsN
ijQAzcTObcR5rS9ZjQ/QNznKXOs12IzbhCockwSjLAdF9aPuPJuVVfkQPA+wGQPs
8ihwwDHlgCW89wosMt7tKu1jihhDOm6B2iT/O6NeedxKQMbFOhro53ZQtyMNzQtp
7XP5q89w1PxpoA3t26ehKLmkRL0+vEdhFH6vM2LM6V16NqOgVMjOmZZOnwnCuokr
wryY7kd/F2S0oqfdpFdhFrwnOnp2ikxVCQ3qadrwOeCkMXQe1TRP/p+KMGY1z07V
Az2GamCejV2//xB47zgVanFCavtZCxEEKG5EJ1aFbuYp26P3Kw0+6aSil2BHhR3v
yZBu8RYr50J0qGtOlOLmuvhzh0z4+6PZZZJ7VpLsP2JbcdMcp5rfxUGJp+QGw0JQ
ay/eHTqRtzC8H9UMxFCdveS3ef2LqDKnVuM440bWXFuEfV5ivfMYSyObk3pzkZRM
8EKIG2dJZmWTKlAQokhOCDf79Uc/6HzgykvxSyRho5UgmQre+c40kEioveSvG89s
1Qht0T5AeDNtWnvd4Td6zaygL+cCIx2zW17Qp2VQWHkYq7XpUkYMjJbdmBI41JmM
nkNGD+GpLf0Sc42lQF63i2420VaQgJYfvUwk1c2Q1X9MS4Io78upIxYoXvuPxfF6
0GA1+7TCOtuZ3+RAlUV/cW4nEfJWcEvMdWJN7Ghv1s+98eCBcm8qKmoURuM9s24p
If/WLeKNBp0Bl81oEygJhnwtzQR9TYdmk/fXP3SqBZCtrqo+KRfVan8uhQ+y7E58
uouR6ICUGuomallJPNl3uyuMUJhwJwkbHMUc5nqVo8CF2vDL4SDZgvbna/n//Yu3
CHc7wDHtU882X7b7FglIJ9xRqLo95OFC05IyEt7TGtAoxMqXp1F7VI9jbt7XCKXR
RPoZ1Qa5WkWXRie8TiOv8afYN3ba5KpsVCp5v6g1npUTK96XC8FwpmO0U1gLbg8A
1TrPAiCQWVEefZuUHO0QQXsd/KBEcU6JHCCeV6hOY4hX7XFIxK933W+5tO5fs9JK
ytDPnkWaPcM6T84cz9CW891YYqywMa+4V9WW8gAT++B+5CSXuJScn7YhWp4V06mo
LYeq1dd0PprGHD67IuvfuIqdEV2G13g5qW5wYP39Py/kjjcGgE9EW7oc3ZQRihNT
ohI3GJ95TNEj2QVM2V/cm1WSX5xja6363Ik3DXALwA21GreyOI1pkwwIxR43KGj4
EYNT2HeWVLzwA7aGIQoU6VXiXkNBWuy1NX8AsON316A9NpEMgVT2VxbrkxC6W7fv
q0juxGYscqAyKn/KzB3BuYsnpS+1Unp3hABZTJ4GMkslYkhLrRErSjbCsflBPRQ8
3Z2FtaFnvohRLaF6ePljtfSYpAbzGFMBaMLup1K+MJsRzsSGBOT372AafnIiVb9T
PdpCaZI2RE5p8St0BgrQkwu7DigMnhhUD7AUzVLlbvoD4CEiERs486CKW0zBQrB1
5ywKFCnqwnvKnQ5Jtb4f/iUkTZ5xSx4PkL7s3N8aePSZbLUKEzzAm3YOlMo6NcdS
CMdNALUH/vXbR2+Eg1NMQB4aNaX4QLnNyV25P1d+b70sNucg4S6e/8XWV/UzsEzC
VKZyKg3FpGV6AB09ZjrvN+mMDv8PUu4cNJQLNeXjalk73lXCM7zaIZ30r8YgUv3P
Tmqi7I4ll7GztlwMri5JhKtwwtI2RGMEjjnfgXaUviY5YxpUmLczj7dzSS9gJW/G
9w6oJuyrMrN+Vpiw/Y46Z+Bwtm/06YXbkxC7z/158CUY6MKiurT89nJMLxukf/vE
tBcm/hgnKPsqmp1valilHQnRm32x8TK4gb9K7XLJ3FL9RpgjKVVTIXpF956bo7lj
P8Kd+auPC4laHXAk3aOCDetMz9S/V3Vj+ArchUKDgQMA5pYVvhWkqK+V0tU/I/Sb
YpeJtCbzsMW0vHx/LUH7koRLhzSo6k1V6i3HloXLmtp/5H5c2QOPxyG+TMWNV5N4
r9NI/uoULTFWll4DqVKDOiVMH6j76n2n//NBgKcJQo/ZQXZhmgKH51uxeeRCFkUa
kWazwDy5FuuhDt/c50cxZYDNhgkpGBeZSoPFIHRe70xldWzL8vQhPxoGD7ru2T/v
ViGtQoquQQK85u9qrHbnoubtyBX0dIucAyi4xAH4HRaslh1OPzwS5cpnYFy8tERe
OgUkwuYCwXNpVGxMH+zWiDDZl1fzbaFHv88CfacswfVKelfeD5xWka7LFxRjKW+k
+WB3E3VFcHQdK62H1vti/XY71J8Ewacy0+GD99+SccRSerOMd7F1/vZuR6m15NKO
XhHdxmxcB6vvDbMObLtJ9jsUcD4eqGI9HG46WVPpfJkM0AlYPDQ2OBrnSng4BHsh
yB80/uC68jXdLo0BLl32/CKI5kHzD4l/9WyZoFJbEnsvheEjC41PHt6dWsDR4sE8
qGjaMfbTLSyhG5fzjBinirkar44lCGl4KE0Q+jbcTjOQTJfFY+2/YNmV+9al+Rjs
ovzyctUJuY8NPXaXH8Sk14ccav3eXuEua0pjKqBEa6g0usLS6J4aaBs4vWt0v+wh
HariT2Dho2a2loLxH2HHwwl6qmORwG++QBMw+KHBQc8Pjm78x5yQQ7n5Ide5I4Ve
1V/BznGbUr8oHiGZl7Ats+/fYtUWLDUDmEj6QV52lFnIskT3FuVEDWfPoNFeGE3L
3NLy//06iGud/GpgxQDm7AIHM80Md8X3hZUn/GsPDv6KUXr0p6/jZyJjelv4tofU
gs29RNYpbw0Rb5jSlRlhT7ATCTrDrQ+duCOWz008Kq0kpM7EmBTavMHDJcJHuMz+
9fHq+sT6eyubFuD0N3wFDq9uoxDowXhc1xhP7sMnLpXdoVFFBb+hjuZI/6mP3NKk
tVmJQKpdTwHTEeFNexn/HgodVD4gP2tS611D6UXH4iwPJ+3mJz/3mKeA0Z373tUl
fMw6w2D/4bwAstCmbfvN807T1N+yqjct6fCd01tli5SnEL9/ZhCCADM0EVRq9LPb
CenqsQ8GnQqlAcbTnRuzjRik46plvIeHMwqR/INxp+MVDU9RUieyETj4VOKjsvLg
xEktw4vxOovk5XeBkL7fMY1rKM/ssOorDIpNmvm13ibUkx0HB6ie3K/PG3Rog3c4
LpYt5RUME1YVeG/V3vLB1m6DuwwKFNwa9qun/vyoxmEIFDjUx0dUwW+RP1Hpar2p
Jl7W1ZhsbeTV68IaIvlMucoAiJvoMiR0UdmFYlARjgAK+HgCffegyAuzhaiCJ5HL
1KkB2U1p9EG3nZhzyY1YHALpwNuQAEfJ39UIY/YHp4m+CvtdsezraxEp1rAHz5wH
mk3WnESriSJzmyrilmENgQ5NBNouCXAtTgHYol3abhk0yobfvt4smFiMx2H9KEK5
yxwj1+k0NdO3KIHKoe0Axv7FzGyp+Ml3LBbP8JvQUF91HpBVxE4jn33BvIzfh+ka
XpieQBCyy8fCiajaBd4ORD4yXh83gpgDldpx/n7WrWT99p/jmiVwO2/9RXkthEU0
SK1VePZ1wSZzeUyrq9ZDDRqnmbhMzO+FEqMdy1s3chr2os0VeIlS3fwLcDsfTYLS
S7SwXDMe7TojbBxuxJSf9PmIanrgkPkhN0vf/GiCXu6XtyZojaKHtE2ZpoOxkDm1
Ov0EoWLYp31DlQ76wdQDWEovudi2QhlriforJI/012WuKRu+9FShiRFWh0D1sfUs
YNNknuheT/9d5V8RtQrMvTLD/v/EgNPTv7MsZz5O0goaSeTvpmgmvDUxwq6N1ADF
Dww+tPsxjXYvCHEwJQqQsfesbAJ+fJjEmX+6z/Of62N6Oyavt7uELJej0GcJTDV0
ix7vLhECeMcIxCe1RCC5sPf0GSLWMxKDDXxWdsEU9zCW0JjJX7KQ3/GBSTV3xATn
/7+RP3iiziH3FBn6RZwUn6bBbpUA46mCKNk+m/dSYRYG5WZ0DT4Xk4q9DWfpDA0h
7KfwSr1dtXgD3wgpxEFZigXTkkibdzHAEUmMCM/4zL9VHeZGlD9UxSLS5ZiFjjao
dtfnMlxTGMkhV4+hsc9DeMXPbXRN/vHoZxLQS1pQf90gPOoGVQWkT7xdQzKZO69k
eZCRd4odbYNEZ1EDwJ0dVN2cRw+mJ5xHQatr78yzrintnIrkYG5HWp68ZylRDN0j
YSMmTlCWP7TqKymPD2narLSG8yN8YCFkHtn1Dij9IVJdqeVJr0TCAgQGzOSzSu4H
BfwunJDy7i1/SctE0VLfRl22CCOjcbNJEEn137eBbobvjdvDSHAK2SggbMKkYykA
fQqTC8o2tE9VswgMmGmLSWDCUmr+Mb9yecSH88XQhFC5hgxCbaVEVRcklkv7oieU
84yXt3+OnxNYnd4i3nQPT/5iqfvtULRi5AMWKDIfKKZoyrLvBoz3Pc6zxTsMGaL6
9olkZJ8J11L3kLD9FBm7Mt+Ubd6ExLG3HMEP//FjPnRS6xqxjh6YZYk7Oo/UwSVJ
SyUZV7KpXgTaxyHVXeoeJ0KgL2SnpGIblCajKaqspxgKM54HYqhPDJy3MQfYUraU
6rx5oFlPp4tB2jUi4cQFFZQYfxrHgozzuItsrRwx1YlD2+tFLz75If1tsqr4bVYH
7mnMgl8rdqBquPU7b/sR6ps/T2ULNPtpCQb89d2lBA/mxFuAXSOy/jEiu2NMyoj2
hI5wvtg74vCd/P5SOfIO258iZKt8Z0HiNxFQzRBeowtAmCuvHCmDpuY4uak49GBh
nTZuDtfczSX15a0vllAn0YBJmP1eSBdxJSXf2N3HXldpXLIKkE1XEOihqcInTQ+x
QMLdexbh55iIoQEaDHOO81IR9v8EJ9R56mMG3S3ROdDo0YbUMMHXAAUSoT16pOZu
3Q1BiWCX5hqMbTQ+nHfxmt8OcR9EFXCEYnaM4P0qG+U9rv4bt33mjNfqdcZt/nal
0nc6Xb6LKu8QjdEzad0mlppjuf9Na4toWy5GQbp2FPFTQYvBDQ+cJyiF4h5VnQp5
ly9bYhrPmAdMEI9FydMMQfcBdQHQ/eNCQv/2jX9HaXwV5uGqFQxNDQFgmjYu9mSz
/1n84myp6GuRoq9Fx+Rkc+0hPMbF9qfd2+LDLLD1WToATZAloXfKEGb/UiL56WEH
IxgArwhBjeoHYD2wHITvrgQQueZT1O7YmKqFYvESKdWoiuK4SmuGEHdzEpmKCdvD
Q6zVOcgzdvAaCSuk0kyJMS3mLIftE1MLSjL2FIh8OcGH/+JVrvWAqnGisdP8Zu4E
RPXTcsSsRBmnC7vZqKRSL3y7o1KjRUTrMY1TxY2abdntGW0E3UOzn1/WVPYKH5We
nLdwa6AL4rmVxiQvjWlawvkHJNxAGbdRHcKNB3izab5lQ488J7fOi5U5QRutCLKM
zQutKIcvxk5AadcFUELeYBGrbegDrrL6jSN9uJ7OH6jCubcKBqBpj+AjV7A5Br1f
nk0JQDQrPaqhAC+dXdOXXEwAnQ6/LMQTWhaGzspcUyQe2KP3MOoxkOvtF7mguqBE
ouLp6Y4rSVQli/jAWMLkl2jYNitIIfCXKv4Bl/aGt6ZCbCNedtm9Cw6B98rTA96l
MLb0fWnsLoLjNXotze8kzLAeywR/3ZgCtMYEQK8sZGn31XTB2FvatXLzWfV0aKfu
+Z1IJZODgKcyShFFjunhgyi4N3kmSzKVScNsXsQ2g62j7TuPgTTeIIL7hYgNdpgh
+cVdMadwwoB1vIO2aiJP3f7kmVcpD1g9IDjB4NHaVFQAW4wLlyR/IrPDI29czIsN
6DaVUD/+gnrNHIkK4ybSzCgb/jyllNRZRjmyvZhycEeGcmzWdVO6VNlmr3Eifokr
NrxrPYwdz1KBOGvLAIDaT45rZeHH+vNfxWPwHpiyzzIHbTfUHXl5s0qx+QSMPBlQ
gDSEO7X/HX9JnPpKz0hk347rjeEh/UnZTsKD6piOUV/ghDruypohEDayaTFFrfQp
9zpeCBmwc7JAi034irtCEVEgCdUwX2HfQltqPtFVTgrbCxPE7RaAdGro+X9eVDyc
UvP4+lG6h6yXMf6hJeIWECP5ubcdwaMqQbLXGtoTmQNdrhZUdLy6rcgdWysQRfUx
6RHtYyiX1v0C93C0P2JQDNI0/WTpi/BaNfMdigp0HoRwA++96l1KPT2S1clUxwf2
i65okICQF1iv1/DGtXRlYLgCDoZ+kuIGHs3pbH6otEyAdRK4d1GpgoQ78NN3doto
mO4AV4vSpA0hG/f2ID/nS3RwVX1A0ys7xy0SPLSYt9rlVLsaAVefG6aQA/7GFebx
ZWEr18IwmAUZkveVa3V6zed2SEO2uegScyfSE0zdI8KkGpaQa7IutKVcHldP25vS
EmlaTenBNm84SCWMDBvJ6H9uiXzqhprGwCYgDJ+l+a9fSQsOMM0IOMzQZVi9T8fl
o2R7oOn2568wUyLBT+UIN4fWcK7YkIMvYnJZy830I4v57yVXNMK+lBsfmcPV4HAf
beDD9auT+pORzTAtMLE2wvq/vk/qLYag8XbxT8KRb/d6EtduV7A5ATRMnAJwy65m
yKoSQZxawO9wPTKdec2kIIcGwvetOAuCioJA4J7nvMEKHXyLyQaC66oGfSY+LGpa
aecq9cJbddTUw4w39LqrK8IMkfo7sSWwTzHFzNcK/lgwbbsivl1CWO8WOcWxjRXU
1Q5Qw+msEPSI4T+yBzRk4aXfZZoA1RRYQPS6RhDZkdEko6ge2/b9Q9qGe+P5n3z7
L+Tn4IDxpb1q41NB0PbAPzUV33Xlif7ZG9xGmnX1vGTMmHD98/HIwbjL267x5ETI
UDP0B+i0kr7UDXIMI6FNASPpy8P9IGb2SdXLqhaWwMPmuxEg6BS/pXtXdeIkjqBZ
PayMYalR2cQnJaRfu1yQN03Xkp3k6A0oh4lXcHBpFqEsymulGugTwfj709TazSn1
ONeYMPdmYgAsMFeRg8gU/lPii5AKevYr+wuMmmNKGB68rhWx7dbGlSky5mg+V0ZN
NRLCqHulbmgA1BY1nha/Tcjl5RsYnV2AMIZ6h0ElC3oTS94fFbcKLXZfpjdXhbIR
PaEBUTG6IEkb8/8vv6cmVH1QIOHaaWq1hRYrITvnuTiRnilW1zV5+PU2KQFSfwtg
XQFRaC+nt1gtkfAT7olXiNyWBoepTEuBFA0/ruD/3uQtaMD0uU5DgrIgm9XfPg8k
Baow28/MRQi9jMNywlg13nrJK/pwtxk+6C4Sf+GeelFahpWVsN6u3Wre6MWwf+FZ
j3IYdpIWVhQfdySgr0sfnAkRW/Z8OeumH2hweLzVqtv0Sd1msCr7Y3CY5OcRUl6L
cpavbO/uddry+CBh5mv943N0SSorJNrjs/OyJPkpwN+yj72jSLEp3cZRgPQyA47S
DGaO7w7E6u4EMhvdcmZNOB51sZV8tHV1ngHAfSvrHn1NzIVcl4PdA+TKUV/ZPSBD
gFEn6ipPlL3UuQW7MruXXynzkrmHpE6qpusWH30qxS4qOHhe4QgwuZS5t3wxWtMf
ErQs0acXdGL3Ki0OPGeuR5qc1W9B5ilqIYhGadMsf/NnD/n0jxNgLUTsK/x13MaE
dHB7tDbU05Lf3fkGn21sHmThJNRZnoZucFp2965/lxd84j+dm8FwAi1uWKy9nyDh
x0+xWdAGOUxiBarnnr1N9Bdf7K7kEPTygqAb3YzMqkv4YM5UjM1SlLyJn/sw+mjp
AbjpPF9IQQXdTIatXWEyVTINYIhk71GG8/BOb4eQ+ZsvZ0lpc7/QldVKR8G12Kud
5tMeQAp0kaKBbS8C+77mx98u6HZHfSCUSYJsxyAjYeHbkHwtj+Px0Gwvk9vVj+Z8
iwcNUDjjZ929bO3OJE1MmVhLF/cvld4xmzTyt496sxNFKTITWEd8GpJ3YhzjteIV
kdfTbAdgrdB1Yt9iUOrZQaykeBEb5b3EAcWWatsZUiXsuzE+ryaEnwFxQaIY8bZQ
tqEu4rbXU1Iky9Vk2l6hajGJspGcgsrDVi5hR4NT3lBt4WHFJN3YQAbl0Vj6DKig
yqN2ZOPQBQY+0qIsjELhgJyApyFSonVvp0y/HvwjhTBFNnfKz+Z+LBJEI7y7Btur
t9iO7aq3Yulpki40FuWUU5cWdrQm4+XVXprjukwrFp4FwNSUxlKByeIvaAJVjlCo
0XSrovlxXVlfTW2ul3dZEByaIpycDtSu9+SMW//hX16gdXnf7wM+RVnxVrv/EmuK
aNqxW2ci1CshXLr7ulS11CPJkzHmhL8EED5cL22vzhhaNAzCAql5kbJyMWY9fwjf
YOzWlqzYSMjUxsq7U61k/iGOcEhNd1K/QhMhgZI7y0aVizRpMXiSNvfTOZFuYnb9
wEMJ6UzNbcLTSMpHcA185US1dE7kSaLVrtRR7mHG34S7awcvqeBqrowL3ecNAELE
UAxtmsO7Z0uEfyIUVVvfM6BptoQyC5KnmRQOejgX7xJ9dlSoCVjfQzSl8NyT93r/
ludJngG1zWNeZC1tNySq9FSNfmmEljuhYYpVX5qnqwi79Gn+CSM3dm+3fVwFeR0z
Z6/4DRCgpwVd/p0gHtgqDnFU6FCdUXX6YXvQOia6mNGqpQSSjAE0eEPpUo/J3pgi
C7U3Voe7xs54zvrsqHQTjL8Um44iVFTer/99Empas45SVMVWJAKhiNRC8WPYkT6H
O8o0DtyPxanKyw08QHkt7ue2Pr1clCvN7PknV95WHXhx5ML5UahqRoV4YBtEM9Xr
vIbl5DVD0inJNQJMr2eAD/yug49JPf2PuyPIJd5/NM4ogx9aZCYomLUMSJJPM5wY
xvXb5l4Z6dV5W62ip3cOVhvQy7MV0cUxcD25fcVX42ADZYzyRx+bzEGwqU8ZIzB9
9SFIhMaLevVWwgoKRXNN8+9et68bpa4nLybwVS/yS/YxQVoWl3kz+LAiMhpRFiah
tR4tg7uDfW4USFVb08A4SXCmqK/ZZRdnii5UHuS4ga7DpsniMwa6J6y7Z1H7dK0Y
VQKzUOi/cwRCZpc7oyEsLLno3NSaqFv9js6128FT+7vducXFXP6lvlL9xA+4p9YU
rwPbyqDD3KXWqYWLenocnIaJf9J1M4lBw0bY8GI9eR/PDv3vmB5u9rOx+pTKZhqm
lanH/iek09k08L7oAlzMlVaCWHIaeoAWkM75yrYqwoHB4sjEdEkHoteIZE3SCEOs
UFkQhOnBZ1Y6z8rABI1sTSCa1TTmCmCXqMGniZHSFzE8eA1Vz7gJF7ORFm4My9tD
CH3jcq0wphJ5ocvYj61tPbC4RVejPrAGM+O9Xk/2RxjcEDigVJAjbpT0WAY8+5H/
hDRasD/s1TXakTOMd2iax9L9oVPxAP0XMBEFe/u4rI6Z1w/Uw3dx3C6fp0h6BNI2
vi4J+URn7ff/vaJW99SeD5lFpcUkyF91Q4NkKtJLA2M0a5jGmZA8eP+Rvq7qR/EW
SMWOJowsivY+bUVx7MIG/aFvaj6210eOwi3YNRP6h1uIRTxsMI5BpT4LsjX6FtQe
VobDmU8H4FJk2H9nq8Ssc/KoV0B6kjJhoTsNOKaBW+8LBzByjQw60Oqk4NdEXPL/
ylkvzNqPN6Tyrbv7THJ+pod/3H0Oo+v4XaLw+nN+VPBg2E7b2bNRqRDDVuZNTV5z
67LmBSfrL4ZKMk6e45+7H/L2tupRPY4oeSLg4nBDRbWODN13Zwz1/Uf5JZ6vQicp
VgzlGdAv7EWAuw+YkEtcEbjNZFu1xxKjkINhd7RCLjE7RQbEDR+GKA6ss1O8friU
WkEIgmTwr8nmtfzrmhoMaFB6PPJ5SrezzX2MQ5RlUzKAP7OcDKYQ67paCXYN9X3r
DKrlgedvk9VfeqUT0CV5gIUvdzd7ih1mPXSd6boFcc+p54qPZi09t3rL8s8x0pu2
hhtZBx/mdiOmY2dvdZob/7GV53uPijlXLLtAmuGPfDP/BGcJfLbYqReRf9u5nVAc
49SvHSeIfOJbSYxPj0FOP6a9qfTaCp2tlOFPXNAfB0MZh/lky93QsB3Wsuu66YTv
fYqlLJ25EINyb9Kn69z/yHJOEVpDE09aQOj8fpNJYgrtQoWYEvm0PSFz5tmw/POB
yMN1ruBRMiNYSWEntdugdgp15MO1Z3GSc1RYTTDHpvrW7CSLZPZA8zwASiAXymd1
zHYEkV4w3ajb8lx0oTc8Yk16X8uCS6e0yF73VYZ6D9/9JpI1FExQzchSXmuqc25y
dZo9nvI5W/MBZD0ndd53S6TBxhJ6oVabuKPklEe/6DEDxgkSLtKMKX0TQZkK3amo
SgNnpKGsgB/tfzX/f4XUXRri6NU7C1RvHD3QFsrM/TfC3/Eu3oeSnKIPRlm/RRn2
61YM1gZB2a6x1kjnZGEaEtAJ8Hago+mDLX7NOuSQjJVffloO9bHcmpzgxhpOQeKn
cL/+uJAbTt2J7kKwnl7DruJBi/H3psiEvBY6yM2v3MFEsvxJ7nCwZLzCmm4FVm7X
ZwHtGcrYDvhsjJ2HmkkI0H6GsBA++P4RdjlE0tl5P1QOvP2ImRAm7f+2As7oCaFS
yGuk//ybRjH80rQGMnVJhhRrtnQZfrX3+PI92lLX6RitYkoup1pIny+jbePaGgT1
vlQws/Aa+JwCCQa9nQ/eDFpYfl+q2u+aSYPFC9OSGZXZm7o7E+QYxFhMZnd3HouL
ueGmFgebJTlF77PLfqpJZaFUQvCfCH1+nnCCeobG0dnlmhTCYD7jLhW+F+4jyr/N
RWPLgpbqnbP42VnMhBUM97LWAN8m5W/VW+tj+RFSeK7vAAyh5O8E90pM/1khN4gZ
HOL+oRcRA5uv8gBRJ5dfYU3I1tMSgO2b1Wn6agCVJ31Ac78rZ5vYUXGcsMRKiJzl
OsUw0gOTyUzKZ97JYM7X8Gg35ID1AptCCRhCpOAfZ8iTxddO59OgbvVlUTBXzmQs
ZPrVb/EGmus7BrDI1hu4uam1o5atAwLlZBGjE4m/PI3bduacYKrV0KgUYr4EcPIY
he1OB1WUixF+nntjndK/s2+/z7pC16kbKVYX76ULr8MYpdch7HrLWbV6F44JhYVq
JIpm5yEiiD4+brZY/jnwuPlEd7LdRr4EqX6aKasrtOfe5SKOln9wZvAAJVc+Rik2
055+MLmzv9jfZvG/618QCrDnH6RlHV+Y1KSwtOggazvnAjj23NcZctIrPSSr4V/A
NKIFjj31JMtAspzBoVFwl2il529ihXb677FXeQp46zY/R6lJOiq0rUZl1h9b6n2y
3aU64TfKZXrDwzgY0O0DoyxuTJGhXN2+s9OwmCewE9Kv5pdtVM/IBVxTBpEARilg
kjOvndDZLHrIWq9FFh+XY/JnOLHSPnKbdeCXap1ty34QGML+j5ODg9hXwdL59zPp
UN8e0XjV+V2wiPvR9+fAMcNLTg/gPQI2xC+8720PP1O+wW8v0+18jfjEJ/z41S4Q
dihE4WT5AxX6+fXIuY11XZyHy8JGvgmhi0yvT+eFq10fVD5jhRa2UtZ5jMR+i/RN
NxsEBdqVF5Np4iU+tOzFUUhjAb8oWBf6CTMs0JaDZN1pnMIIhvbakmNeiKE/gg5q
YbOopIRKliHjcSTzDudSdKZkBsPkiXCeOVJ6rRv4nnUnwAaU1gUgnAe4qRj/YoaZ
xk6GLf1OPE6dJ1zUzhLlVY1k91+NrbE5bBmsx/ZjR0WMYhnSCXtI9pkerMeWno4E
kFBETBr7zEeqLhvl2Ad+IBzlOQkC+HUQP4sB9AUm9BfYt/GC0yNczmH0Tx8/0+XI
EaxmzWRynRlGCSS45mMsMPd99VGT8LAtMfQkvoWM8R82+9noPh223C1PB2CF5XOA
7TuF8fA56KaFsn+raQB/hI4Y6fxXGpALovG516410qg4ZJOcxZz/jo1kzFUtmGcS
tWmu2myQ81Ruq4Vx2x/BRqoLO1gVAdjYb2peiixyMV/Y1l9QPxGstqmnA3oukzXX
PMV3GD137xjCGK7vnZ4o6m6ep8d2tbU0GnUdx8AiIDob907Uz8tTeY+pt9Ymlpz9
aBmS1PW5i3CehFHAF8xgIInMtf7dddWyoNO8tttrKS0OM/jTccLU3dnCsMPB9RJ/
JX/75A2GMbPl3PwaJgEQa3p3kiaZYYJr1IetDgXM9FtqNkKnUdDE3pjiqTpaBP4S
pbcBHI11CEmrBR+SdpU+mLP49+kXPgPxyedtowUtK4A8R8oSaoFhJypgavT05bPa
f150UH0LlqGg+v4UrfPAfGbw/OVgD6XV1DpcgixHw0HhSYgu+EbAT9YVjPZ1xXoJ
qyFwuYrIswfLaWIpvSwe89TtwGRw1+kbGIKzIREOxLWOZuxRtrxT7CoMIPv6SpDT
f8MbM+zjEefuPAPSeA2fjON/O9vtj/86Sl4q8BUazPbfd8xYEq50dxdI1wqau09U
ACaFoijYao4lyZ+GqwAgLLxhheTki+ijndjrMzGJrUhhssaqgw7GZPOYeWAF0qE3
RQW7lyjGZbgh70blpJ8uXy2q2HtCnwxvj+NRlrxRMIhvMiGHY6PKTnZFZd2Oepg0
kAj1uxkX488KxhTq2M5ZmjhZxlacYfXW49aI6Z7/9Qe2JmEDuH2CDcWRPSzil7Kz
1Go2PuDNMB1ssPCS9LSqm3dby1Mz3O+KUHWS2vknBmKAO3s9IXtWdx91DR5D5TUF
CEJfvRlb9+s61twl9IhX4S+lxtCeXD8EdNt5Ydxbva4U3Y3rh2xnxKVCI/5Y698i
j9GtCKJ2W+bP7KlHpKkNVGBzReeB/SzHFWjMPpPywxdRx6wkrfv1dtWunOE5oChV
+NIr+nPtDCfFXDMe3oO8SOneg+4ixBPkG6z4MdnI6Rfz3/4aSFcLyQ9ZMa6ZldzH
Z4ESZHq2yfuoa+w4PJxgpuEhfocVeMm4n9kpJOhKwlT6z0tV+kx04C2afbDB0Fx7
kiZoj+F3w8a9cvqvSfHmTfcnN5C7D7L6SWRZjOnkIx9hY1UiA0yTN+s3192UrQgD
0t6tMHGk3RemrcWuJRNGehBWFFIDPwhid3gZD1W0XDMCAJd4Y8irszYVw7Aw8l8t
3n/J4cOfvNHR+h/ZAHNv1YgjrbgLEEXIWg7KJK4UGyupO0zKKcM46HNDczVmSM/h
2ofwyXksnH4QwZUrpZZ4ll8i2p/R6sPvPDHNbmoijmULpdbrF2RStLSmC6hiqds8
eyap2mgQfEq1IfrF05P0GkVSp/mRKZWKF1xETTv296hRWdcDkfLwVWNa/4UvHd+h
sb65zf7Z0t0u561aq7cRubdcMeYrsoClzNex1Aq5OPMyiJeQUJTNmT4dks8O2Swh
wKWOP0hvUFPumIFupE6D0Rf6hEQwXdPeu0XMPjZ3d8LzK7BVI0l2qmJkcaVjqnII
BLnUlKONdKnu2ggx5w+Qu81KGfSxDH7JiCelI5WrBW+4gsdKxfDJ78gVlz01C0qM
067Su5qYE3ZbNpnQ4soTi/4JfiJ6yCcvGehkkiH6G62/Hr0B0jcFhuMaD/lNjEFi
Mby2emX9qM+5BrFAUQp9g7KKxnleb1CtpXw2nV8uub7HBeemFDp2V9VmVkyqbNYr
dREmL7kmG0lRNxz7o8l7xGjgAwuVtQiABvjmoE0oF+gnPO5WlsIMQw0LS+liPpLw
DAzMaZzqtfv29/UmC+NZ6cim6PfwRHh3ps6+RC13g7THbkYvBQB/41EW32A3PqvJ
BZ6b5fbAlIW30viaKMfRfwYBnJTcSsReKBAyZ0QJRq5kYQKqIsv1AoTfuhRkYAew
iSETRWNRu3dEvOUbDix0fKjbxl0ZSzLCacE4QbyBKV4d4flMLFjjGnmhTHx3vjVH
9uY3OxAmPH3mXTovWyqricvZcQKys9gbmmu5Gf+6Lxnbg2mRILGOV7rxkekUF9bg
HBwIRUt2BXBQadkDGRgaVHcMdhdg7tCSM+NqAGcLQWwmGhsE8hQoLOupAlr/gLho
dj/kQmcDB8Rc1eObPcP2xD1jRb1EgOaGcg7fc2/EKch0K+GIdwBFIuuxC6FiXFFr
51KkmVbTYUWNc8PsgU+aQc6cBiweLmkSCLySczTv4HF6F0+PJ10TJTVeER64d5+W
m9OQW4sMzEHo1+hfju4r/cTqE5zASfg94fH2B6Bu4s2Jf7z7lAbOWiMgthxCA//1
FqMjcwNvT4bMauZVtcrGPyq/XKUyPSaLSgSsosbIL/Gbmjt6FnJAaN25cH9rNf3W
Z0UDiCWJqjOJkoL8nzscsME4zOj7sQ6ZfOdJHTK4DS+DoXokG43e3iwdnWGbx24X
5pPfXQHypYl7JtRbmAxFZ+LxV/YbwhyaB24BKtRoOof9V0bO2fBZgbh/P71wkzpX
o3prSzYNILUg+RhMckdFjunxh6TOdghzhQpkHEpG6/5F2DjYKlvigMe/KJiBt2WC
LbNzMYBzhXwZiAT+c4ZEQ65BugbcjpJ8ECAcW0ssz2IA0POM5bNqXXWULiH5Gyso
R6wsCBKJ8nyQubGAyq71MrFAS22qqfVUPqSkjGbNAhh9T8t7dqE6/f8SJiTDBLXS
fIEsnjopKG7k9+7YPxEfSTs5cYOFW26s0uu6wlIFsadHsJHWTbzAirNo9R4+fr7k
PjoWH4MbDpRVMfQfuO4dkieWgeUw8Akl6NbfGgPik5y/iKklW6k9h9LO9gqBdNI2
Xibkk/tDzhZnq3mEVY3y6hxNFWAtIAFJ0PiFZEdpR1VFeKyQIEW8e7jEzN1ynnUM
0OCOamHbgm9VTGNL2ecROPpl3b1ZWJ3MBqvVDrjIILtSzkviFUl1LVNclmyDwoX6
muLZb5+JjDzqLo+1O7hWn1BFE0D1wvlkcpN6Vt+aMfEJPmw/cH+3e2PEMiWdtvgW
LyiLwUmh3xr21hbyWAKlN/J3MpCfhBZeCc3xS0+dIHQ172dkxs007uQ7V1Zp48qf
+IJLcssFT8+z/1+Jax7hm9L1qabn61hpxPASLT5MNBwgbaIkEotZWwfeXAFIVKPA
SMCOoUM99k2ailNL7O1rEoylDEee3ULQterQELH6Z8NqG2s0K/BF2tsRvVnDjbPP
x9XBvmJSb9qBBpYiZKoW5UDH8Irc/RuumW8STgNgseFPTots3wlKtpKL6TRRnrrf
k9ZHqPiX2d42vHvIsLjGqfQlURodUBiZeO8WqD53h8Vc5jM1B5TvNCFRkELbAvGP
vminyekgjCgF+G0fiGVJHHbCi1WTnsUpS1eOxZxmGhFrCRoQuOajq87VKQM0E3mn
JyY7UK2TwT5zvizAZ4TjKB9u0l5HMM+eahjQ/1AQfE0QnFS8NSYEQSG8POTlI6yC
sajjKSnGE40rPvl/8q5ky5dQapV0n4frUmF+7km3SeaMHQWSCDUvzyjD4gyH52bd
nTwl7Dh4Iw+kVW03JbVYx0zG5IHLPuy7L2TZTZ+0cIC4XL3W5PUxs2k8tBFUXwzi
PJz97tAkEUi79xl8lQB2sXwhj2Q8RD7JhUiWoNdjd5UwRKNP2V4K7R8wIdqI8IbE
RFFaSgmpVH/5uHkgThLueKFf5XJy9+SQ2udX8t798Ws5sKNVxHpRi4XA1xMZGrrg
5rBL9hH5cR0Uk6TTWsxnkjtkA9q5aFDtjF7Aa0k2lyEwaobDCpt9Z5I7y572DTEC
Ml5VNl3576FzG9KUSeF4pRN4g3Rm9Y18jpS201nTaN81cJzPe1JCTEFu+w96S2dg
U2UvXTJMSW/BAO7I8FGyTSjC9tHBed5wJE/PDdjNviwlyxu7e0xfizy0inaILKq2
x3q8bKxRxDA5+msBwwvcyTY2qxm3Mhg1YnNPbVZQW1jLHVEFEnKEKn4cJI0yALJ4
Er59BICgZ97BmHQD/j4ZRPsOH5Pl7VpumBOTkQcphCw2GcqRFNnyWNkluEL6zHd0
sno+9Y7v5ECRDbenocY/61w2oKvW+lg8G2wLagSXV/hl/D9dSaSnMJe9MZkd7qT4
Pn9Lr/nIxz97bvVAyxaItWYeF2MfjIbVX1WAXQibgzYWB1Ds4lB1lKVwvh6uqjZE
7v0gC1dgUyGYOZVcTiHfKLkybjtRrffOeGLld0hgpUFiWZrfAikibP99d5949+a9
sorlnEv9r1yPc3XtYZXEcdSTsdusiuMaMXTI9+6l7KYjnrCbRYboAWg2tndRyuV+
GpVtm59m76sFp8MH7XbdjY0cJIQB03oXKmCWZtR4iC6xKj/HgJJKQB0ApQ/LBdMI
HcR5JVxUAKU19UyEtPx+cI6DVmiHz16s7nMUflPKj/7O3IlQKa20KsJ3KN/j7b6h
YOhrKk3wiXI44if11dADh5iX8sozRrxrmVxGCllXjbxr7l0yE9UQ7/eKu4GllBrh
pUHTlwY5PINVIPF5KHy141tLCoiDUmrvTRtuKppOGCJgnnXqs2hvgU7Vw7HbFWuI
QNWKXB1XS8QsxFvitWTP8hnlA6d602DhRQE9knH65JfMc9X6HARt8TGbWXsUXYZI
xGNt5gw9xBBc6K3pk8bmXZfKtjFT9kZfu+Ra/qh0RvksK6D36b0IF/9zG1feefnR
g0HfKeEwB23q2RFOna2TVDgoeXfyb+9ouCE2YCGES9u5kF3D7fdtmo6Ra9kZtxFD
kCpqRC+cwJdOeUlwu1akNfS+n/KbX+3ojysbQRixzwAOSXKKgWcKTNYkWFcQqMKR
8387ABFJ0l7AV/6VFS+Oo97bkWFQQXgYgzl9UuiKMuk4Qf/C60fZ57IO1Zva4YqK
BFuSUzFefXS8Kp1MshQF27srKRvE8hOXIBaJTZDG551GHcVrg5PrxNByw7c4zVeH
5u6d0xo1ZyjFjYXaJsbAjM+v14dQKrr9y1FAM5fpcbF7tjImPvIjOpSykujYqzLH
uBZeHQjC8Bk1XRKxlLfwsPlhzD/BmMTydKziF5slmUquVmvSTCNEKBQnDoWBxdm5
IBC0OqdBuByzMf8WMu3NFr4vqzp4C4PmBcJWm7qvHNX2lWCB4z1SKTZxIHV3593e
l0EX7dfKrCYh+NCJR2WwrWHijOG+k7ma2reqWCtQCD2uHq4KnUJ2K25/ZkUNp35K
nTFilzw4asNls+HNaRFWM3oFG9GEtAupCod4hEDx2E9xqjB21gX0m2iF63370ff5
tg4gFWN3FL1pYDxNCC/fhjteg0Mmdb2E4K0o/rOWWlnl2t0CzFxAq+/rajxXnMtL
LWNbReqxFYXoytPiPjJc1cyiqzWcTH1jVELdwSCUZVpD7r6VlqhTNIUUZx8dGRUd
YT9UtHnxo5U5q4B6+ml8tqPa/lyhLOnZ4CxAqmmoRrEcMdLRtuCS/jQP9kB0i65S
l2/JmpTx5FU/avCKZ/klBWQ469zUk3X57Bm4RgJ/zl5NWcdiwREMrUOPsGdoh3w5
Jm44EUkf+z5RlfOU1FvDuRT+1iZSTkueTGaVYfz9PmHZV48Xt+rlEVcajHjJ+85m
p6nwVYH2WaxEXZNoub4OE72zlt1hrnmXqYAu5WCDAgKDQxFV+jHANd+4KIyDG1a+
51PqjG2HjiwY0HN0N2d5p+RaywWQ1r6xyAMY+gHyUNdYmuvqv+pRxjwf33bSdYKZ
ShkAkdZp/slbRjFJGUfrlRhzoqwut9nbXQHFRmD9OgJSBwPU8rztIAi5qQoSzax4
jLZQdqTyH/KFprj0bGAKHhX9hGw9JYC9bh98LWfq1xhg1ybdw9QNU0vmheVrBg1o
BvIJW9ynWWcp/yrUCEGbFGxyA9Fi5dVazefTYWp0UHIlIUJ6y635zjOGc1axna9a
6p1Am9D/BNF+UgUrXVX5zzwEy0bZF3St3Zt+o5KMW7GyRrSFD2z0I6cGGqB2iyc1
ZRj4/pOLsIBhwlxlcNQ4lS74W2gYeV62zrwIBqTEIoiViQLS2W1/CWqUscmO3hVs
5ZtAmwhS3Lx8i3bQ00ll9+mJD5kZBTzseHBMkwZQija1KPw80H0maow6867PJPqB
OZbEwNOBXJuZrtbmZIsmRuFZNIiFPE+NS+vEhc+I9fdQcFV3W3e91+95U0b4/06v
oCengdfgPfnm2SXD2CbXDhq0oBWt0xIuLxa8IUtabotmvBndo9IzrIxKkkI/KCXu
h+LxE6v2fJEgMjGGVn8BnzTEGw/j7e9Wwr3kRt06VgXXnDQkldpB7PJqrt+itnJM
h0lPxl07oLsXebmPVPKN3wX6ujHiRmkNz9lIVAftsuD1K18S7v8LPSg34iKKaWve
K+BP2XiU79J0QW9x9DgfYQVMYjfAgc/ahgt1Dtvb1wsmt4UMgYbZAqfOP/4relx3
MSlAwwYEWoLSsZtkyIH7TwoFL6nLCPx8NiE9k2gfraGvAx6qcpinCVVg7uq+p7l/
+X9/q8csU9Wd+kAtPIDQZ4qoynSRJbly6NFZHXrSwfDAJxdqQZ1h3YkJOPzGfo3j
eMZIzClmWzEIQX33/IML7+zAnM/c95Bw3IHIEmki5vN2GfifSZuVKM8+NQm2gVaX
+hpi0wJ5AKPXDyyji+guvFHcBqpRncXn6LpwipM0Yf1JFiGDBDtvlhlGSmjqDPOS
6tO/hpA/5SAXXBoVjkQ+BQBOtY+n+0M93MTJ73EtZJOve5mhI+TkCZe04MeD+Rnf
vi8KEL4UqEW0Mdb+BeuB+WXsahPSbF0EYSFps6TrRNBTi7SewNtrYRyFvqmhkDl2
5z9Bhqqqe2Ae/gRLbuE1WRVhZfVf3QjbtWFsJ75vbiaU9t9TsWcIGhI1EerqLfuG
I3enW3GhShohnNGhXdthJOfx4fCztTuOSxhbfuSFCdhx8N6AiMYpJW3cmWM0LyTA
b54iK5X+hTdBMvhuc1piAMHoDn7b5DAtrxIFTYokehvEG/FiFl41d2joNZNGMWxo
Svslu51Ntvsv4YDLLN0Ypd+V+io/kAt7stPc20LY4TghIWbm1hz+pZ50QEA2JVLK
YKnLYI78Bh5zfQEFVrIHGlt0aYTnlLkr1j9vjpnv1DJlnnTWdewdpG5LQhiqAPH+
eqR3Y4D1V2G1YsY4iGrVggzgairBGyZWhT0BCJtqoqM2JmqTy4hSgESQWQMkUlkz
bIZRMJCDnL+V1ukk2SlL2t7xnoCIglyf90YWo4o1eKTb0typTy5GNumPD0G60Lnm
5lFZKqyY/kmVCnPKBwe9ZaoQQkvzsTNvdzbIMRiKHqMf+fEvr89k+dXKsFzFj2/l
YFDFz+pgMFJLuZV83bQF2uSNp0PVoItEk6EE+VIwt4XjIKcGd1ySRRYlunbFYbG6
2CAWUPkKwkbWAnlKqAfc4HQrXCpT28bETudsyeSCyiHtlTUVTte8sM14ZKl4IavB
LscdAwbGjq92rpNh9FYIBMEZdk+VLYR3K+sQ0Z3xP3mTSXnvPDF3elZOt0T+Bjwp
uOMYZzWIi7xqT672rKm/oDZSj1WQ5cy+AtffYx4kEAcs8+Fta5c25LDpGDVYNui8
dTc6YeHfwP94/dbrUW2TRrnaA2TTgodQfJdx91Orohw3G9hAj5ru/Mo5MX9GlWzd
Bf7iYMKwBoRg3oO0ot23fZxhmmik9Y2EcEbqKgmLEQZjilb2omYL3zWeeQCmOGnO
tdmiw1npCosJa2/1rKic6HOy5MZZUwLmR56K6Kwz6YYZ50M6sBp89FYCFlvUdOQR
aGXDaF5Z6zSZFcjvJwYLFN/jXsJD3jlUQJ7G+LKONivk3rmF8FU6JoppKYW6C0kh
p0Tum9dMLugwDS82lMvPl6Zg28pdU5cCY9omodF6ZAfD8vgzDTI34e1GdzPATvLp
Y7uhclMG3IYe2DUrgcRBpncIgKoWSWCDeKYP7rnf2zkhDCAoXxmeIu9fzfiaUwAJ
olh69YxdfxkG/vIrjmg1LTz7x+gHQi6CK/+Rg0C1cXwCaSXWpuN9ED0Cfl88+/Re
TwnNe4epzU1qjXmIpamwJw847TIfqo9f14bCiNGHFJ8GnQyf7YcKPZuxvnfKgi2q
oTFsMRCBUswgN12H6XiB/4OsfdLZBrO8WXrjEH1DM7KvTumL3KFlE7rbcLE1RD/6
ZlIz6f2K8rynU/Gov/cFKA81PxBvSxnItePe/wCalqXQbTujbSVEicieUrpmu7uz
PvIizdhYf+PvisXInfPhCz4KA+5IQ85cRfOlz59zrzgsYADv3/LcRZPMhvVj94TK
I1y4Pukdry/w1fDZN3GlPVpqWLJB+bU08I+oAUjfISNt4JZCwg+SsygRNrqSBHOc
C6UGhvWYQT+qdbZPDDPTRoJkajAjyUsssScraaXaFuJpgooAdTIBPzW+TPD3T+Oq
Wl9ZzD1J+6XCJ7DIFZOKPg4eLn6BhvAtRIEf9nJFzqyMJXXZdG6ykgty0HhS6MKH
z6VrthNZJ3wKXy+IYKTwOPZH0hAsXDp+DtMnEIzoZLY6M0Qv4ujUGkjl/F6dGLAx
ydqc/srUCEP9LQTEb4UTEd5m5ewmNwPtXqYU+0IkI2VxWVRIO9ykiykYsVShSAgb
WML2F57t49Ri9SeXIVCe1pCOs3ElHpjIPJzmpo/RrPXFUMvT/XRyn1FVXCj5prcB
T6p/ZC1bORBdaTbQu9lFwckMXy5mL2vJAsb5r+AhyB2k9A+pt8/Jrf+OaP8PvFRb
Irj9dWZPIzF6CEbwjC9CSZnNv2EgbXSIgHPkoqTTaHkixsYMf4xT8VU7VvxyYkGL
2cHdYhMqfJ04TGff2nDtsmENafe4bfFMjdzWPVRTGQRQhivlB/yr3GCgoVGDh/In
VSQWJVoUMF4f6uTYH1oOJOsBuHPbWuZFj1mH46RCQrkc/xOtPt/weVUOReDplUug
61T5Cnx9soNogR/7bqyvAMG+/FFPx6p5G26yi2e+DzH5/PfpawIOmUV9iWIUQATb
ZgZhXrcLg6ZoqGjBx7gEatNTmlZMNqCFdwDzCERKGFKWAv6xYPMPd1pUT8MeBIzX
IcwIX+fEdavuAYurlMugds+nj75VeU2KCZdHzVRkyim4v4n3lm3+WU1CTpNcSc5s
65MwJMnq0XAupZp/bIawu8WcutooEC6+EkN3lIacR6F9SC3zleKH/3pfUON62FWu
QR11H3aidRPx6o4AaMWD2uDNmQmg3HTgxBSM+YZFPAi406pf8rXWy8W5HW6FfM3C
OOsH2SI/IJGuULNdXIYeEgJ+Nyo/3JWJ3zqAMNHGZiDPBB3UGU5IME7/QW2UB+co
tb9Fu6HFVAcEa7G89VDCOqHJs1hs+s34hVvUkXTUtH8MKLfTUxewYqwnuAI3lqQN
mCDG8YS9KWEvHO6sZC4AwL6t1UgWM9Oa2ckLwtRp1TislGmnyrhKcdqQwiDr4tk/
qGIa6xDIuXUjTJaC85Hy35fi1wASmfAjpqxNS/+cZj5egWp2jJq+oQ3h69XzkKuA
SObewunxT63QXcC3QjbP9dJOYGeVp2idmUYBqdq/S78++jYxjXPKu5kqzt5FF3To
AVYGE4zK0VZXTQXWDGkEZWvYTV3aOH2bst1bKyRHTt9FVKEP0hdkXmHkqT0PBZk3
a5hD1axHwl3DqbL6q7phGiktbDAIe5L9WB+c1GcaXQwfnGwQaLPoRkJCzFO1A1yH
RWn/cqdAhgzzhZRUXy/0L3N5QgUZ+QYRGlAa2Yoz4UmBQcx3PXmmba+RlNb7QLdh
idx65DFvjisMp5nQWAJu/JHDgNMonpl960vqnZVqH8OumgAY/6xO2bRfoCvsPDEv
U0sGDqIvZjA2a8rvMAHIHqvSx2GbY2qcI+MMT8Xqs4UOtoa/ZDimoKUf7OaYXJdp
3aDphXR3AxYWYVDPbmdtRcSTm90VNHrT+obyEa9Iu8g2cuS82zGOwNZkUBMJT6i8
8Emi1W6/2L8nVSjU1KatBkUetiA4L0O9a+ELASs7H3E3RJT4i1xM9rmyj73O4Fp3
I+tLL73rkJq7zXtVo0tVMqAReAo2T7EUhOXPeZexq0PrQ7FcWfa1Xxvi3pGqKWTp
DF/D9Kl8jB9xpSvzNa7Me6pMO3pFe/qn2Iuq/D9RDj/oPQGepKtSGCg920jj8/n6
HQdElZL0aBZyYkjDmuOYIP7CbDKgJnrANsqp/4sQ2szQi+u/d2I2l7/aauYNgqIl
7Pov2hhMEygsEZg1dsVwMkwmr1B/YUTNwdZTWNgNcOQlZ+NvtpMLUh0AMMKF+o9g
iw2nc7I2Ri0orynEDRvKXTGzp24IwfVlRvjr1+z2/xuL7HzFtFqh1436bOu7V5Tl
6nbkI2ZxRYDKKhpY5/vk7PtH1LkK3srOeffDYW/S4EdFr2UIXw5eVbk4k9mWGU6H
fcQvfgJ1WVywQEudIn2F9kmlJ19wNLWW562HEl7ogyyvW1bulWfJjFSuPnDah6UQ
XZcoAenvW6vy7v+r8dmkWs5hZ1DbMFfVFqE9wtwyGIP+2cpedzSWpjgIgNpSu7uS
MIydynjO+bXaCF7fTCGol7IW79GsZLtfV1a7bcA7kMM58ta8EAOqKD/W3t87G0cn
+Fa9JG7e5dYA1BM+m3f+4zd7joVwklXX939QOyKUisUzrkdjXM9dbEKU0dtaWVEw
Og69eY60zfrq0XcsoNVTeU8pXzjoxCsKkWc4ktv0ZxveT7U2UUSbul9+VKqr0jzJ
mv8Oe0uBJhhMLufC0QbtvFUI5lvyJhuJ4KY8QHBDXbO2FfmgxnJ69xXwx5cuX/Mg
yT+j10HcZ0ADOrgXqCUgvOb1pxogDhAsb1xVCqzFJACpwbw1cqsz355g0uNq5cBw
it66Po/oDA0uFDITEAijloRY1X9PTdV++3FAq8jM2/dOZvZUKNHfUW6cDWZRpa6R
mnyZ1RUyeqzBFwpBpN3nEcXd7bedCeKmwJaj7ds+Y+b6ZPlp0tyIYCtnLsky9YgL
66hwe/vIpK+lqJiUboF/MZrsbU+7aVggxVuKLuz8ieIESz2LfSefMG5ysCjWiioF
v5huYWuTiArdb3lAYcLnnuns1kfSDEr/4Tum5U3XAG4=
`pragma protect end_protected
