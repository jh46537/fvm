// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sBpTMd/mU7yDfxvzw23yDcR2+NDPpwzszDIDFmHWNjqtbJqExi9ijJM8Ko9zdT33
jqWCJXGXvuvB5GoD6aqk7RoIz0TXcRotCnyEZVnWhbdsJ7C3tpKhXUTLBkIOOmJL
ZElIhn4ZL53WeQyU43gfcZp1BuKk/0NjLng3KSSunkk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10752)
+puMEhtzyXDDlKucqU4fgsehSKRjZrzi7ruvJpZzvLGW6Ar8ZQWouMRKA1LNoQPM
ymo8seMxQ6bdk92LqCOX5Gs5IB2GOPkRRfrs+HaEx/2uSAq2rAVLKDnvPhPDqxFx
DhDugkG3VDR+tuG/AntAVdKEhzx0NimeKIcgYEa0ogL9wuTVpCqErWQGsD5e+qP1
WhaQ2TdN1J+XZbxJsCT6JsWV83pcz6DAwAGtuZYW5JygSFhFCN9r1osOOBzJbxNw
Vw3D9Vbel5oLtrPXzG+u/Nyo1VHCZG/Ig8f+qqG0kdoikB/+IUiNtKj3Z6ovJHeN
GUByeUJStGR225WeYegm7skm9xpGhho0YF6BAndSnlOewvlysRsjxwSbRbSGBdrZ
VPATA19Hr+CZVQqEwrLLtryvueVRih7rXl8oqO2QHWpKgAe1NYnWRydtVmS5QF+5
/dlgZKI9jE8/gA10nHuX5Thc9Cv/kcBBvhojtxmsX1XZiqQpbcmdHpjbQx6NHzRy
9FlRCZUsmpCmy8pDYJ7qeZ+QJjS6aeV/q7z7PEz/vq7qEqebIriYeuFtTeLgmWJV
1fu39LhOc2qCeCP1qjKHzpzT9ufqp/uyIayh139hvGUV9LRu2a6U9IuRIlLPVJmB
WJ9Wk/js9ICsqcRpVrZBVWnvu6lbL5wBkDobxgCsjmgMkgWOdOi8K+yf0biWwopM
9NB7EqxI7SZ4eg1NVpVO6qkd7RXSmc3QVSgjT+hIPkC7gxt6xSVMjU35zMOcdYH8
HIkqMfw+0wy5i3e3aiHal63dXFj1ETme3jZYc4YEgTnlm+3lwYb5EMtc8QRmgzkd
KEY+JARQSeYAAsmiDI/E4zzPUG3EN20xLFje711CsPzihZZkm/zVr4i4DiUnSb8p
R6AeRlHLI7o3chKqCxfBebXbCzkt/GKbr8psTUrZq6RdgEq3xfD3Z7RckBOQHZ4Z
AhtmMvn5isXTaZ5P1Mu87OoXwcNzMxwNvYdRhXOhicYx5A9W0V55dQjhwXWyF0KY
SilN728RWSPj4uS0c5T2777V9q5X7DxKmJQhsMEAQNcL0RvkbjK/iR4/HKAjlYIn
Hv64jY/PrdYikfuOeT2DfDMuUQGJ/i44HM0oP6xxjH89BJApyf51aiWhj3b23WVg
22gSoM12NjUJ7qqd06IflsDD2/NJ8iGg9wCuPzul64qgSo6gWnye/gly9KW9bH6f
BBGA8JD4+0r9U6snWLtYkCf4lUKhU9E6Yka5VuV/Xq/hMTfkMsowouNQR4V9eKY2
EikEgeEKYZDdPL+OIwJpcFXLACz7A4MQVfH5EOuaog6YlvYGJupkiX02n2BCBa5I
xcr0PCKw7czeF6diMF5H3PYnc6G7zhyonhE9zcxh6qU2+FyhVpr8z5VEGRY1sp/8
h9Uqb70le7r2FU2OXqgtEsl6FIyKUyWpOqQjP9ixK5uZ/8e1NGXcDRU5HxziTb+B
/VB1xoZCrofaM87cgXYKYEVt5xuZ03YsV3hYb7SeFexwEjU2bIpGsjx0DyvsyZG5
+3ikJu1DezqvyHBhMq8726n9wrsmKNjStpLxxTAuMBKADDJ6iuskxQV7UL/Gxady
T5pIgakzsaKNeStntZTdjSA6IG45/bSoqVcqZS/05fyELW0ydA0GsoRUbXj3rWdY
5ZZ+Lb+Gm0l7gsj4WqcIE28b/69kMupPkxiWCu71zJC2uJ9hIL40w/bDbCmzJhNE
udNI4bNFPYbD/Duf94GogNveb+qiXaJ9g0eVHfpxJJWRo/ImkAuARJtLU6A2xi3c
w5bXOuM/dKXSweYX45C+atUMX5UPJG6TuZ0KfCz0YqnLZvnN6hEWthGz6QqzG5Mb
m7QAD4RCtwbXDecFDPGdPzXX4gYtq2IgKHuyB4H8oKlr+rmeAdoDsCAsh39ifuj9
4NGUtiQoSZyPaiXh6HR8MlRWvtXldDxam6YLwA2qEU1sth2bAIlA0hEoM9kirW5F
EGaihFmyWfS8JTJdh9HQBjkXyFcPBYA9brzJadOdRwd6cYkhOPxRhylavsqyb/M5
PsVuFSPbrdBThbKXM5QzhZ4H+VEqYyK644wHQS7amxOZkCRoxeiyrdBbS4DHAqd+
eEmsogmm5QSa/Jt4ack5LPRJDucoBtUAdGA8P7TDD1W2W4FCeWTDJNfcvzpuzTCF
sGZIFfNJPNjgkn86DCXD2hYhrFx15y0iGnlU8WJZ1+ibOliZ5m1rpm4Dua4ffGq9
206SlRdxoHc82hMfiWjMP3fT3wkMoW/xDVdZ19Pge8t5WjgR+76+SFpbjAlNDSK3
4HKU+XwdeV1IfE67Vc8hyhsx5RtK+DB4m34Hs9RPMqy/MKMOuQWc1fKEP7YCfqMo
0UMmP3hNlc1zhpF3LvEoyhzKBXD4zY8e9xT2Yx3AprtN02ehVytsND4xgT6mzs5E
hTnwvyqIlSWnN6cd3u+WWw6nUoVl3hHOOhuRcKvbYhv++G7gKMGG3LlVBi2Sju/0
TQMWvLwd9go7fgkIKpvWID4vltN5x4c9ctE6Mg4TGWyIrI9DJn6RA6loLxrjFoqX
KG0mq/1vN4+FLwAw8n1GOvAOxf9smVnGvAFRsxbTYVGbboC6I0x38R8pA2iYHJTj
sJiVkh8RJ5KMIFZ9xO+7dcan8gQHp2XN4VHcpDm+2+ES+aN1lFwZUXL/4dUK6RyR
EGQkrMWeWfY7NQGNtiH/BR8JLBQx0GOcbtFZmWZl6OxsBV6ITZyPX8U4rZYa60O/
vfP+W/F1mGy3oacXbnIhMFRsrDHEWz/yZeSvUNIUavcC87lu1+fNChI1rfX0Klv9
vszi5xuxnCF8D3DrLwiyyhjJPvpo2CWXv84FSokAF+Q7XDpZ/z0xL/uKREp4VYeO
8lUhVnBjn/aBKNj3TMizsuChdhI7Iqj4IOZSnzhTCLqEUMP33apIFbAYuxqm1ncA
JuHT9+WwOLBFRidXF9Q2S3PsH0Qc3xJ/XQqWOMzLBc/U7ToaBOWKonnbbvTyCIEc
lYCUZe0cdflRup5L2TiSBacQmUxnh5QmM2EVFcFPz48E3Y/KkGaqymWjMmoGoDe4
A4ePCobEnAsjAUrlhuqVJ2cNBR5C9LD+IKMjLRjRuabVq+KVsn0tzroLrzrYyDT/
rZ5Pa6Nxi51u4EmKfLZ9i+/3JcU+MOis1OzE++gWy/B1jUt8zxgfxKnZb+64PlVm
iaStpDPdRYy8WjLJraDelcwk9o6kyLkKOB51RgbwLBqmz/WEDINspK5xf8i6cC20
ExBGS0IaiP58FFW9IaOSUV7NDwM55hZ9PrfCWix4wCBNMCYOr91g+38Hcl6S2fMy
wirS/5auuJPCdgMfxMS8tkaXDy7CF+Qf0EpCgStgaFHogwJ+4yuCfnM+AjGxe9Ui
7hWa8B+yIy5RwhgoKrFx/syFr0p0/i/EWW0flIclvyk7y8ToU/k5/JKwqJDYSPm0
GCDnN7VAQx5ssikMrviBK381vJ1uhIZdIVQf7asshR5gkwqLA9He3Jm8PHDAi3k2
Cq0IJ/kJPAxN/i58FUMKvWzxuj+FFGu9NFKCVkPmm687v7weStzafwU+dQh3xhsM
C1MFunQXJCkzqo3zUdLwRUz6dxY+xQQAT33AfeHz682Y4iGe1RJ5qaDYAlFnVUaL
tCsxuD0pd40B/EJ5VdicrxQnpl209dAlRLbamqLXGc4czpWVb2bGMqbHazjZAotH
3rfV9bEvpJg4NztfpzRXdyLKpvb7kuQUr1bx8OY52TuZcE/FxPWQlRvBR9CmqKlC
Bu87rZmpL6PiBrfPhl/7Z/frAun0ZS1FayQZtzbIj+XjuiyxLzOy2C44tPFjcOcE
0gk6DghhAzha5v9fnHJsIP1tdHzIbWXzBrtjKY4HXxFcjNEijlT7DfBOMdLGQXBv
yiEWTxYjQ09gSB9tDJExTN9SPqo4GfONpWKfL40BdX0WmlQJM42I1MaX+ri2suNS
69t2RevmENX3J+itT/oEfjwBz74fQHdin18RsFgGypdkTG9GSvkJpXcWwYBFTTNf
9VgiALeIsF6vvM47MmAG0jb58dTtMtXdiKDfkkhW4Z4co6KpXPj9hXvi+pyx/lFg
k/wWm2iGKp6iG9e/GX2STpM2axs9Ki9EnCb+36D2mZEELedD52Rud0Ws4RmJ4GqG
5eDlv0OnjVUOKjdHmq1dOzwQL6pUUoyfkFJJAABJ2rTaqbKL8vf1U3/lQRvLl/tC
s0rH78YB4ursUTKjSerH9GdkcVYM0Wgu9SQ5ytZzF0PWPLZMYg+H9bEN0IOnrXnn
0NyCD5e+OkVCsiqWhfyV6ouAmlWkwe2sN8S8SEY0bpg9cra11iqN5pgia9oaUjJ0
s2mWoWuyLIpkbk/kTKJAUdk6irfwkMEVTvstQq8kqIb6s8y+ImwyWtzmHLF9E0fu
8vMjnAHypC2C6R/ei8XjTxHuJP1jul1so2qZG9w5JtDLMcn+7L6za2FLdCiRw2qT
/5Nn0h2bRDTroF8ffnhJQgexT7CpSxYfp2K9qevneZG9XlP8PgjP2XW3UGXfDLYH
yoknnZKIvO/Bpy2+huGDflELJ2k2AAhNhcd3Ronq/G5Tg6jQsz6+fNNKmxo9eMIZ
HlbfIjOugXv4JkkEDrTIrPHMZEWntd4GPo2Nr18zQPjHLaYO8OXIQd5DuTr2xaQ1
i5th3pH+9XmePhSjk0qBKyNKFmKWEcBE3i1q38C27Xa1i2daRNLlwMrdawZU2B3U
WqL6Oxuu1loL0itSfrhmhxqSeqfmeblAyfJ3syhnD64S4pxnLz1D9ssgYGpKwJKM
bIKh31VP2pT0E0WJi5rJjQNE1SUDu/F/DNXKsuDAklZlZr3ncuWGgZe3n5PEDojg
8HGiNXaAxyACtziZXoFwHAfyTseRuL7iVN39lNrNVZWUKN9+xSbUY0Vq89T6rf8s
xR/9BuuD4o3fUzo1cloKd29ycYD+MqG8Ke9xC+Vc1a59kBbYfTX4rXmU/F2M1Sw4
Wpar2mqqigrtI6Fngydq1WOuTrdnd5FPljI8DoAovkorKfaP4FyPLtjg/JQU5faZ
+Zew7cr9I7um5RLseneCWt5Lh0u2O8Ri2Xxv8+AeGjWYPRgSTHsNWbnqNyCR8RqD
hJgClqZ5/Y1jm26zQguXWWVUOckFCI9uWUybICXkWDujNKhL2hJNvz8lp3aFUKSE
icpJ2EHFVuzYSwpV64v6Owaeft6UopYvSYBA7cswbuiaxMXlqST9ZUbZHCT8wNdo
ilLTeBuaKI7P91MUm+hHcUtJ5axjNTk+6NgjRj7w2Au/FbFXteRh5D2X/z42OMSd
nn3C6N06WVfYLH8l0/1f1Hitq8rOwnR9rdBjxWnZhQeaBUTdBbsN9hCHYTNig7la
B74kd4tPOBplLGJMjsfC6cmIBXJrv2rFDEaOCt1uj/BiCWdsn/BT9gpzk0EwUfn+
Iz2H6PglX3qmQ4wXZwi+bqEquPat4XefdHz2YtNCmMcBJRijV0jgeMpiGwqyW5nd
hMyWslRe5I/iXv1EnbfG+WYm6mT/W+gsp/aPxLdZ+Q3jBmeoXeG8Tg4uNeRel0hW
4Ile7uRf5UKzWiqNAIz63RyjhOvNcj9NDLB8agC6vJ+C1XERUhKmi1t360Flv7tC
o2TxcCafSddc0crQ+ISPbg+Sx/rXOa1GztlDEkBw5hqVrMGiSGTGkq4f08rulU2A
T1R+wTvLmPpQ1ZqOhf4pxJx1RhE2Mc4qm1aBIN4h4KxHphwF7lfxgDyrmQ6ISxEn
XHH42bjcu8XN9G2TPu67ftMbXdc0qNuQjRgdiYzCt/SIjXSPZvkSOn1cUw77ux18
f+5HIMPePI//b8YzePbuagZhTtkon5rw06W8fvDzQl+UqBuadqNAhGs5cLSTBtsi
3gleGYP0CKLbkxSZZKJUPgjvyp+RkHEU5puDJMN+bmpkT60flcGCD5DHuZNmsWj6
iilpoTENFzufrYrIfBGBTvQN/+UZVoI0B8afnDKQTk1A4okKt9/D9XrSZ8B29DCm
G3L/jnaeOAsxbmww6FsP/JMXWvwiQNgJKPNOn6J55it5LGY2cLjfaCeZo/x32U5Q
VjjT3aK7wc+BTYBckAnFFfvusKIop/eKCjgrG7s4oN0NC5Z7wkHjS50O6H9ySgFq
1fKEEEF8FqWnhZxtiNsR0lXDzczzTxa6gyzxLUI0c1CdwnJuW8B65BO8PxzTe0J+
N9l6RdC2I6vmk0pOdX+YgDjSMwCWvcvQHsNIpQ8Sh+/1nMArvAmdLQBbhZvtX2v7
+ZstUTcHo2dy4XcjdfBtbFEHl074B+rInhiy2RLOt1WUy8pCuVQo7vc/3F+FZEsD
0BrLV3bWYVjCu4X9aEI+CCGPCP/GO87GqOq7njY7KV+Hx4eoykbAqYrcIeZiLYIn
me7G+pCuWCwPc+MrnVHY62HtTjbQC1oLdYZcJ/VB3lzJzjeorMwaxj7/DT/By3Ly
Oevw++B/BIhQT7MhTTRaoAEv3suJS42eGRZLO12SpcYz7aB7A0wJ/qWRoazje9si
FocPfOqi3zwdnkIMVAsni54Dy4N0T0cZwVvNbhzbsg155MZp6IJ96Mtn2bVdX8gR
3T1YRnweR7v7rlyMdhf7aI5ueDvZ2tYS2AC6Z684b4X4j2tuN4vVE8ZdmiF8DUqo
m0YleA1ghd5Y2wz6XKa5QYm0puAe8za087CnfBrsr4VkZ3vTZsKRhB/hVa6yjwfC
jRa8MBMhw7nijiRaLfFsnjFwmxvGX9yH8BQesBua1vCq2FKqpHY1hKjYwUsle5cq
NcsfWv73xnGRwyOb26LvSPAZLOWkg0xMxTFmk2GWTXmWKsM6mqBwVlA3RxVWsDYy
BZhMoMN4roUMnvMCwOBq0eVKPL1jzb9xSTjTMaUYf+8Wd1h8dTuaFjQDGPZAPYZ4
ZBK1H7jwoBtWqjJdiDoQ6YBtir4aF18SwKHIvjQq6oWqyj9slwZEaCJjSMB4sWxK
JxAzq5pfsb88cWBdGl+HybOD05mEp0oqtv4v6fKZoBaWTtMxhOFbX2gs0X8un9JI
07lXZUmEc/rlRyWTd31ltDeWeYUZYos+sqkYaRvYxE0Lz33keCbMXQOmQSyrP/ub
/lQjnRwfywrpyfM2y4/YmHE0504MhvkTHaPSFyI4gviN4PHtUE00a3m2SnhF3xAl
KBZYGpOXP6MfBpYxq1bCNo/L85gB7VG9qwyLjKQ/3ySVoLU+bFnedASAh5bproLf
VZWAjIwZBAKs4qtTm8MG6j0EN+a1o4lERPCMN+uvSkWS0KiVjVxFnFVjfzyt1met
S3VkeVHMX9mgENoTDiV8yfXXGRTnmGc0/W3yipgYBd8ry5dNuudhH99c4VPR+Uvj
D4u74voHrJS4LgOnGSUSwL7A2rKRK4BAcvranHQIlgb45jHAJZBHGF3zzLhd6zWG
wKNDc6vvS5ZQbbz7W9R6X3z5lJm06hbRy3JT8ysuzhMKpbcGze5Hg89oXmZaxSno
n+aQTFW3WTjoXHP6dVQLVcFghzFPCc088Ml8/WORJmeKL2r6C3taXJt2Fy/mmH+R
O7dUvVpLCnaC2IB3QrwhRJzNd8U1zJ0tTEcDUa3KGh0tSJKwWaXSfZPCB0AW2nqm
1ZEszOTcme1KoNoeV3eB71/JHLJnRkN2Qvr+C4dL/fIcftDOqgo96K+sLp7lHVCR
/ZeStDQPuKujw0XtarnIJ9oHjawYwq5bLt41V3hJGMNIGyMuc6WSoqwEsl9gwnje
IVf5uXvVHAnCnwbgI0XzSsdzGN86UZGXv/vcipXad1GAsNlu2hYutCOKPozhhP1C
/QOYYEKhJ96IerQg/r/gugBlLWTtD5loc0nCfQZiVwN8NsyXBjMoELaCvaChAfsp
9wc6TxnIzswmxwDflpwmyKVjGG+TA9NOmx+lyN9EcGHHVT5by9pP7kVKOibqGbHe
MbBywKITXdQoEuaEcfeH6B/wGoJdmjiixMtjqeO1Z1qlU0ywYjIcFuMlRiYTocWm
ukbQLnXQrwPWHAD1NKdkKSSnNh75biENaKqhUlAQQ84Uhzp4GnXhmmJQc8U+y8bD
KIsRJ849wpKFnW1BQtj9pjbtJRyIf0Ra7TwJE7sAWCdtAw6efBc6ktbwhO4+Wq/O
plzp2gGQSou7GHJDcXY+y+fXgXFFiXrL2+YBsvdSqYYlRk/8oVU+QRZZXbM1Nk1i
/d2memtXVTYr0NXbDSh3HvcfIs/vn88pV6xBMN+P1UmD++RA9Om5TTq8yI6d6aXg
4DLuDL3ablWBYRnzKepT5AyhIsKWWdtCm4id7nRIunDRFjBGXV/7HzTqzMFO7FkB
ql/ooJuy7tBjTB5mJqnRjI1CUEPgj6J/H50R3IQA/GIwYfNiQPuWS8NFDO4AStWs
JBIPhfVl42gSufeMLmajB4dnzolyOFlM9Yi9qgFejSksIEYDngNTELMNkpVoXdoO
tdKodvdTac7ljo6N/N0CqHugV8CRn24jjL2ivRl0KAtetUZ71gCO8n7g12+GQDfC
mpzEHFcDEo77soNTdYjhj8qMcsH1YAXMIKKYhaHZ+KRZIYbJNrsxFMzJjAdyQr/j
uhg7K4U/zL7+XNW04/H8Tj4PqLlDTykFL9AxMs6PXP2phAmNrNrxP9tf4s5n9kdX
9XLEDrer+kEkFcKjC6JB8TQ7tfeEuRWwRUyQNXUFd5YfFSZIx17jsaqxPlRnQe7P
z5gI7IVgiU63mQTdfhvA4EdG5QXV/XqBJ1uNC7wHspmZmNBL8bLoEjfwz0hgXk2X
PcTNl87r7Ws3WFrveAylYVvhJjsiOjCOlyJyBAdZTYkYpNBkS27iALCSC3V3cSIK
dNSIy4bcmATZ/55pF6k4/E5+hfb5bgvMB36rt7fASORpRLIBpyK7/Vum/jDGsXAx
sQhj+RuX+KiFTmC28HKpqCEAWBKBdDB9iKxFgQTnd+zK/3SDasLs/Zq+qrgX+4yz
eBkQiBLu1TVEBLPK2K9hgj6dqc+rcsoXyK8RzH4M/uslGlKDPRBcyX6ZZySj7My4
SjhWEQr0WinrGCQEQPZzt+HQ0sSAbqNTA21NiLGiClfN0uoPA+exgTYdmeZTGh8p
EVMimug3be1YnXeVMVQ/+qGD+n8/ww0oW2kFeX7DEZTbRv6ONBS076/5VQM8v/ZZ
RdHgbjCuo2pfjtWe6Bxf6pooXYBSJoWkZmkXkw91AJHZHVWtPuMBcJ/uscuX6QJa
ZNVuDBAE8en6oCjZO1woj8D9h2pPNgtmucgOG0C8AbR2zSGPmrhnWj5hvP2/Ys1N
G/R/6UFKmOYsW9houZh+UpQKSpsqflknP567dvedttjRdpwnBGWyMCnSt/iMG+ia
uHEHvBfbxzBWrIMYBfQgv5FOYhH5r1+fc8scJa2wgsGcSl9tRFkrftgl6MgmFTcK
tFeCnxVAu0Ey6i5BpNdS5gVduz5KuIRHepSVbZtEfbCc9YTPp1o6/voUBqxNVNT0
u2OGD+lBsjcYnflW2l2XQDEv3lyO3N1jGxVJOue8dCIrBihC8Bph1hwNJD7gu2Wg
WGg1rwlfVnqA0kfQDtjpi1lW8HubGvyY8peNumcg146kAa+5oGZBm+yhd86dFZvW
at8WQx3U5EfAaulc5s+3lgNQ0/RKg0z+4yWtzsYZ1qkfBt5wWfGajiweQCnw7qGA
Lc/4eE+3V95VsJ8iBb+Rh/e7fX32xgz+xBoDy3Z5BICzx5zsaeofkvvv+8OfMODu
n0zC/TANnrzsNZI8vgCAu4ivOD/CZJRdXzXqzjp2O8M976u7sN5wdF6zYG3GeZJM
21Il3aGxxnUimQ6wEwoI+ux0gTY2cauIlAU3t/aQCJcEh4k9UmHw6rUREc0bnNBu
Gfx48rmS1XLb6cgLcXZCYDZDNsxVMLBrJdDrobNCN7Z5do8WVITK6ONRIJmaLZB0
4UhoWR8SHpjlE7F+Mxrb42OVs58qVhseaivZft6WwSQhDMgdJA+w7FWtaIef5/D8
5vHe6a7anpFOxN6T+6LUoW9sXBz0Nbld3yDWLqL4z5HOa/X3dySZzHePgqOSbY9h
b048N+ap3IjQVNexZH9kdk5DAIwHeZMCMcXGLimDNy2x3PvJ4BD3G8mgyFcOspl3
YWUYQLu2NHAkgiCooHkIp2gxSUVLW9CviDKj5GHFtwmm/AEiVhV/DHT3QUCmKzQv
2yXJ43wxwvklGP4K9rUeHu33ZolMxo3nLcaxwWcnaojRHJq0zgez2tBuCyTYMzSb
h7HpHb162sGSwa7OmPMbKqJDKfccZclagRe+1AQ0ZQWiPydnAdg/ROWbPcMMYlni
TS1qb5rJci4AdS9UItPQmjyAbHlk9kY2BA8YKOi9ZsGa3bY4BmtrZ4e9XHXyB875
yb4ogGJyaKwo4w8qkthYpWPMYFk8NkybEhO6dPDT5m/daCjZsltufQWfoyhidnp2
k76+UgCl3Tyjffu8nOkv/aRgweznaRk3lUUbE9W8l1aAFAYAEKmj3E5QdQwNocqq
juhYyvSO5mfe25hotp3o0SrMZslQVb5FRkh0Hj6PkCFfcEu2ht1ZTDmMaUZM304T
wvcScPUNn91dESm/3c7fxo2c7JYWi9SkKEjZBRgepMwB1kqPEuVljPnC0GLWfQns
wdlPJXY0XD6VzusD9meABcWHYcU/9WqAy8wb4sczUkyp/djxRzty9NVlAwkqshqL
eQvM/hBHj2zAXoBJIiAiR1Z3ejQxi2IO40TDfujdcDTBQjvMFalRwwMPXQ7f3fZG
GTYNYurrTzyPtNJVpoxED6kpDjw9+URuHJg4xJs9PAqBA+O2SQNIEkmddCdT6fbW
DyCJsOEiETjUxEymcOillmB54Nqvb++me/Ht7hfFTlYnz04q46Y+nmymvi1/aTo0
54rw0f6yUAQ89rsHuBjLItsN2uaZZr4WDArYNf+fkVv03LwDShPqRVMvLWIxGHSy
bNNnDrYhQLJ+xkhzzQQS2Nt4DgqebTJ7vGRTYXq7VPeJD/BrrjrVlut1/yIq9/31
OG2tDF/zVt6K2+H7poyHY+vHw0fwzWJMd/Z/9kmPdUBpWn1fyO1rQBytO8LdVroF
b+JRl5c3Wpxd2R5ONZBlBTs/EGBLKKRkpI/Jv8N/TGG10ZP3s42I9xjfSKivTfc6
tlWG/YoMG9+ie52gwJZ9SulsjrpkKKEM9gdGkaVwCvyoCwTQcyfZcV2StRhgpdOI
zKrQm3N6zgqIDiCGd8wIcg+Jfa95rjt8sTGbEs5R8Vj9fM+ptrx3/zPddz2IbW8P
4P60Aft8tLXfbfk5srF+bON/2hHEOQ2f7rwDojkuzfK8UnLIdeOrRSMbhrT3AVoc
68BGBmCUfDkV2n8LZzFG99BBW0QNowotXtJ8nvkfMLECJMuNUUmSKzPVXJmNoOCE
2qN54PJ0szw5E+CTsoeJ59mhINjdYTY/YqqzJCu4/0arvbKFQ6FSk64VfwFoLaFp
sFH1fGJBkb3AD6qGtxHn2b5BojJUbDhDxydHY8m3zDwHc/mdK6nfupZi/vq8u671
yfhc4ErMCgo0ZK/45FS/986yWZ2Lea+Z9Rlftx0h7TWAbbCoLWkNvn4ynr0OS3ox
sb/9aZ0wAniYve2HSMZ/Y8+Zc3og962QSoDMITg7SudIimXDnGjKkTss7CTu3MzA
48FP2ge04UHkwsqGELql7w4Mlol+g3CionrcG1mqf/dkUw7Kn9FFNp2sjamzlAyT
Z45b0RC710iDQz3gP0GS/330WA21GVghRwAGJwYUrGHDoZKr14FJIkKBTAyncD9n
7SEAFs04dIF2ZXmpyX7sLXpB6+UDxhkrW40SKYNJhUWGnUkemr9650rWml9xfGZ7
HUvj2pGlC7WXzez6UzCzAvnRNROFh01bggu4f3ZebGhQfAZ5bd/iRx+tf65xfnvD
Z6A1U2zvjtalvu/TsUVcRkwP26lNwYVsJyllVXuv7R0ccPArBOvgYdgNgpVLlWMX
p5OOgiLhVTRJlBQMnEs0IAi3cwWLeJ1stTvflea1uuD5Min6NpgnwXuM+9BULMU2
kJ3jxkv01yOtChy4rkd+U6cVPTE2qkRvF2TGTpC3Jfm8hTwytobsg3Oi+FN3/sza
l++KNtzLHHyembHgeVoTmACyMWImoiss1V38bff/t8obe98f6FqvMpvXaHnZObtd
LZYKfME1mK2VkJKbdyEa4QYVeVMXeUhWRAoGs5fj653BfOID4gDC4RKKeikO0S/x
DLsHPQFjcQxiEtyOZESvHpUxm5CYzife/JjEdAdQrlgi2EPBc3tcO67nYcPI2r9i
Wbn2OiRpsoH2WZcY9PXjVIg9PxMqOwiF5+EVAvRBgtINWTij7xJty1t/JKE3mvT+
c2eXMD1LRs1ddFIMNYhtyqTU4IpVALiM61fsIbgwnfT616TwONfGYNFBnxQCTiwR
cy/uDqdQH65RZ5DiQUhdA07TEFnUFe5PgfIZf+kvFjueFzIV/iUAXhpsIOdmWpeE
+Yj2asw3wjYWbwRnelZHpQU81xxajngkDGUv8VXY9ZBMHzsbOq1kLs6m5tnaZynH
4UbYMyjdaslKzf5DFwCnrd04EsukihkdECD8h7CHWP7VJOPYQg7Me9gkr64C2yyp
+YfzakQq5B16UniIMyy42OL5EeNpOUXPTvgqJnI4cUxLiW/I/tvLRXmaSIWOj/F/
fQxTRb4Hk9m4RUlBe3ATUG7n/RqjLaMExyD3nWmi2/faOmirt03RK8+4LdT8LKfp
RfUQRHDY0sgY0FCPlyxBC+nsfdv5bRWXtQ72wR9Yf5Ceag5NPCNQcwO7he08b93a
aFjhUX9TP2XBDxcnaVTtL9g9FvIewSKTN1F1/+5lBFYyhhCmCqXwhvohP3aKpzjc
10dNW8K7Kma5OYnJL68whmcq8c0oYZYAgH1LEjw9tJfXgSYgm0vfKmcsSuswkNAB
zYfQmPzrcgu9A6M8IdffkoCpR6uruggCAcUYChCnGnGdTtVyAgITINdjxWWGEC7t
7qjxlCJrJ1rjC08X91+ne0C+mIYx30fuYALF1FXheyWkw51+4IpFZlR4ZyYXbS2k
yDscKe3uo0yh1Sut/cwIJf8GeBdEjLi/8Tj8aNn+n/B/pIFurI/q7pcQ9TQOgpPR
DaIcdpd35EiwI28jxkbRr7TooWKHPNYDh2NuBon5Fqrginy4E4m73QQWqOOK0se2
gB/MnVc5a3YEMoyl3KkFkHyabNJsdznGYot8memF86RQHx8tjoLAR1yDL8la29Io
N9nk/qAknfBCQLrLoQbG/HpQsrWby2vgmAVqIV5k59JhYNsXlzf/OevwD7jXZJ0A
mNsC4tM6vpaTpu0YsWS7ejdf9I2W8zHHQtFNcj3W8fPTwUeZkbmEKFAXIDMrJQtx
dzNhJliVLX8LWSFfu4uWk2bSlypDUwCcSbSUUlDkcxGbkV94BD4CVkhEGdRKLz+F
dNvlM8UBdk42jqtFBRH19PVPi1GkhdvAExVs3uan+oL1yJWzv+ZyrR4oosXWPrvG
eYXTdrsynYzfhlZMqot9DiKAYAnavo80OJ0sRJt931Pjfce2eGBR+YimkyhQ6ekT
WOZp9oYkuDPREsO+32uOaihT/ykovrY3E1c9tr3NdDDdrGyQFJiA4alVuJhi6KxR
kptuZasOb8M13UmheNfaPAU2xNIB3nQ/fyvhxuyQCATB36Y1yKtMW/rT8C7M6BZT
x7P3D5DRjE4x/fDo+yjwUvQool2LwDIRPwXyqOd7AfL1b7kfQ7uj6BKQYsO6c2O8
wLfFUNtKeNTSVj+568ROzjnCqpy1yA50Vw3xq/41c/gS+sg6OCVR2LJDZKHhBirA
Hw1hwe+L/Ae+mwLzLufCZGR9eNH396t1lfhMzzf701dI9h7r6iYKAGgYlGwJYB/A
wHm+/g8T2lu+pFdRekt8QGe0pK0V8zvGyRgvBPpD0cS/T4H3iXJPO1NsMYBqaA5+
8BZ/SThvi14jI0QSfOp8hYJMGr8ENmR/NcTyvAUnmapTl2Q8cAH5e28vxwnra8Ci
WWKo1kZ58+Ek/Jtk96D9RfEIlp4Nmer6/8CGLCpG4lISK33JyQaV4V3u9a+K8UJ/
6m6ZR0m2tIqgiVj4+HVBDkinn900ydvk8rJvS79rqvfWQTFmLFpqSKmqQdrtOMSP
laboaDGT/V/r6iui4o9mdkOl6wKhaZL4VKvrIV3eSnoPDH7j60EkGH5tz+SthkKh
tvZP1DGr4GH+cvxWo+c4rguB45NGB7u6qys0pBYBP6Jr3XoW6srBKp50vbz/jDhv
3dgur//Ov4NYNXuYZQJs5iyXvaCDGDeYiVyiq6AhBdDUwkdS0d/HHGHsMCyB/gWq
`pragma protect end_protected
