��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��S,7*��a�.�_/I2/��m6 ^g�ԝ�Zr73:6�I�e�B�#P�L�a�!e	�v�z<�,��$R��%#����� L��(��6q�[���Q�%}i�W\V�(ª�S�	���>�(HM-�4�Q�K�o�dm�������OhؾN�G����tآ<:��d�e0�*f��W#�n��ty&�-H.�?F������0��Ei��f
9�D���������TWU�{u��J������1�[,\ 0b2�:����~頨2X���Fn} I��'a�)���TG9P
;�F/UVnZ�߫>�ls����降�ܓ0�Pk��Q��%���j�0%�̕�-f��H_�ۣ�:��ֹ�5��}�{��]�P�DlP�.��?q]�_���)Ȅ���i�u�-zvN}5(���"��â*@���cGD�4�Ե��e������t�c��/��˾|�Ph
;��LK���xR����.Df{}��N�6�)�q�Reo��#���D��}�Yx�4��sZP{���V����G:�&L�q�$+uJ$_�T$&6��=��}+�Ҥ�-?U�U��c�����f��ڎ�!!��N:;���Ĺ��`ݷe����ׇh��4�E������������
�)�}̆Q�����2����ARQԁ����u���ӯ��p�5��Cz��(%���]���7�����<��	��K�mTmD>`/.��I���c�tp�� �='���~40�D�I��Yn~g���A��CM�upש�[�n�"l���WΣHSV�Q��A��~άmڼ����|�Q-P�.�q@��8��_b�+�ejo��o��!Z-�к�pi(~���KK�4�t醦\�Iǌ���0�)?*+\�z��]�K��z�׉����j��r*j�V{6Ƚ{:�A�G��&�sL�`���fV�T筒���|�^S`|��ҿI������YCt|�5S7�@�*I�[��t���(�ݹ� �K���G�[�l�6	�h@�#_"Zb�������ɶ�����o�1P<�r'Iګ]Tc�f
I4�~xس�{�f�i�,���]Ƒ[��E��E�B�L8mP�
8���(	*�Y�t�:��!>CМ��� �|��c�[Zk1���=��*i�ML�$��=ԭ�A�l��X)�*����Qe�x�	YdE���7=c�Yh�!��q�%`;9�4��AQ�]MM��i�����]���{�໕����6^�_y���,g�γY�Ml�\�����S�%��Ц�}����=�;c�2RY��iy$*�cŬjt��"_�_����iԌo	ë�_������
L�O��>���JwK14��?�-O��}�7ٍI��f@M4�ΛJ�V�[z��1�u����X�}ҏi�p��sU��;@�7�O�I,M��[t��3�n�@� ��Ir�2c2�HF	�0�[�͋�MzQ��I�_{f��t�q�a7S��#����������r��Fe�)��ͬ�1�`:A{���yߒ�~�����Vi��Sҧ!����3�˫n��x������A[�����c���"��D�]j���ٿ��f���`k3�ި���5��	����*��������Y��Fj z��	p��DИ=��mO$�MQ 4٭%���v;~��2�6pRD'&�Q�C��?-1�3*��0�̋�C�2kI�f���%�5�k���ҟ��:/�S��q����dG�P�"��Я:�2�ƄMuT�R��c~�֯K*��Q5�����T"�"��H8�������K�����Z��v�*�0ӺI�W��\hJ��	sH�&��6E~�?�x�����C�&ر��8Ҋ�yđ���l�	�r=-���?� l�����.8{Ip�ёO�=u�Pq;)g�n'�zW�zٮ������GJ����Z �R�3�n������Pu�>�'\��9�<���Gl.��89]_1�S�O-�Rk��N+!z��q�75=��l�UW�����rjK�U�Nr�*#�}���ەg�;���$�r�|z�"��39_'|�p ��<씦�j6B�wm�`�O��EEz�O���,���1NyD̶�H������B~�Kxԕ�~���<������}(��Skn�XB�������U�.&Ɨ�z�̃Y�Z'��i\_��9��V��\7��3x9 OF�C�'���
�� r+FY�%y�RD`P�ǐ�X�J�Nf���Y���khʁ�9@|�"C��?�)H�V�2�����D�����?�/� ����$u��:V��P��G�1�¤�����t��}��;��R���G]r��[�Pغ��D�6L�ܻ�����;73-°#�A�~��րF��5l��z���j����u|΄��"uU���\5߄��X��ۍfڨ~{#��&����`������'Jh�$�0[�	���DG% �f|��u�ڑ/e���D(�V27��ٔT,-�>V���l�T�N�fX�B)��&ϙ��hf�cDưv���R)�7v��϶
���[_E*���D�<2>fڕ�����$��F��i����+�;��e�]��;J\w�_Ao��G��!sMmМ�Qaì^�W�h����xbfԀ_�q��`{��B<��3�����:s�J�I�A�=Ǹ>?yK�"���g��w_l0�,����0�c�t$wP�C`�g��,&ތht���y:��#�w41�$��m���$x��KbR.��e�+�a��n�L��v��@���"�^ZI�J�>K|e�	LF"��d��ɏ�r�jBj�D��(@���I�Am¯ס�P��h�D�`-|i��~�]L�,��aϞ0�Մ*����D���$)sI������_���<�\ ������!�ʜ���57� ����O�ˆ3� [���&X�?����5��X%�O	��"wT7Iv�P	Z'z���7��9!i��;�K�����x�r�B���6&�0����{����,a��M�#��I�NO	K��%�ݤ:`3R�+�� ��]6?�As�ϸ��p\�cl��fl��L%a���	;�E[���Ԇ��W�WpX����ͮ�YW�gX��܌���C�Y[��L-P�䭄4�>�����9 �%f]�Ru��2��pz]���dJ�WC����Q �~���#M��3Cmq��3,T���;�0� ��ι�M���;*@��dʡ�&��H�a��[�ņ�*�����e�%ǿ�4ʁ���l��K|����|@v܅��,x��S�ߦ��,j��JNi8̏|U-4�6x�Q�D^��#��������m��F�����T�� �;�UJe�P�_%�T�����IrL��>�y:zl*H�T�����#��)w����߆�y̙o#a��>��[�w����_u`�Þ���M�G�v	������=�y�}:C�uf�'�z�2�I:�< F�Mtj�|A{�Z�(+|��q)�um��B����_�F��o}:�Ú	Y!S��H
jݖ�)�.��2��W��``8��H�2�!Lapsz酬�(�},ߞ�|'@B��O�Ի&��O�:�L�b�z*B[<�uQn��B+O�b��y�(�,H�T��>�D�X��P��	S$��*P+QȝBY���(�&���*E��5�q�,����բV�H�Y�.�Z�<:�7T<��N©��Q�"�BJk��g;@4�I4C-�EPa�2����5?;�H��>/Α���}�}�|�| <ɭ�x����A�ٙ�aM\�ܲ��ё:Q�Z��d��Ѫg� 'k��L"�t���z�G+�SYNw�o�F�w���y����MŊ+z��EkĜ:ml�".D��i��W	�����.��.�4�x��.z����)j2�D=�U�t�Tρ�9�aX�7�\,����D��� ��
���Ӈ��*�]��l5a�Y/\@�4��ԠQ�fˍ)�K�=+̌|�i!@ؽ�ryy�I�4���T��~u�sԳ?�z{e�A���̧�z*z;�⬏-D�ﶞ&�gʬr_wo���v�z� ZI�4��G�	k�Y�!�W(�D�O>��F��b�4���weƾd���(:��b'4���F��<�8R����/��o=�:1�.��;~	�Q}B����̛�E�������_���Mքw!^T�K`jvi����ym�b�-
V	m3�j8�q;E7m �
^�J�%�.��4J���w�o�:~�k��`�A$�$��;���7ʏ�%
#�Pl�[��p� $l�E��P���̾�1P@���B6��~+����U��c��"'D��'S�d&rt��= 3!�)GΚ�b%�����&Eg�i��8��]]��װ4���Ul�\�j���m�pV�nCk���w�g�Lt���3 #{l'���g��b�Y�
R�ߟ��L��i����Bjc0u~(ɹ�>d�2t�^q^�;�ʣhS�%�^=���gn(�Q��%5�xTɑ2�.ƄY��%��׬�Wl�.Ohy޽�[={��Ε�o�$�i�dB��*��w���O��MD��T���=U5¯�2�W�gQ��{p`�(�H����d,G�MI��Cc��;,vq�O:��v��+C޾��|f��g{o���Y�j�9X� H�_qp#$��J|8ͮ���
)�Q�/�/�P�hE�v��2�䍄��T��Up5�xؘ�e�~!j�9���������M�c��G
��#sQjv�i��Ϛ�5�ܠTCX�5�;$5���>�Ve��@��}�2�v��U'ā�*ʾ�}�C�Q�����b���v=�q���J�p.˧P��"�,BȠ븷����q5��U�[6��M�X��>rD8x��!�	A�L��bzU���y�\��6�G��� �1�b7؄���CE�Rޔc�k��=F���}���y�s©�o@�Tj��!Y��K���)o��ab�m52چ���ďP�lIJ��H�*uR!c=Й����VO��� C� �Îǁ裯w�*�5��-�L���}�'΍�6,��4���T{�To3����H(�۠*F��7�8V��#���9�l�[�7
0DكX;��i9�F��xX)��@h�ȹ�rN�b��(?�3ev@K�xTp
��
�I �9j�\7:ŏ����i�����X9O` щnêw��l�!}����J��N�t�����(��q��zt��{������v�����c��Њ�1o�/�\U��W۔�,Tu�V|5�tS���� ���n���mI���_i�Ť�g%�����o�tAk��5,G���	}�}(�h���*Y)������C���Ö�&�lGߍ^���nATG�1ҥ��9�6b?s�A����v��o�ޞf_Ĵ��Ʈ�KH��ᝯ,{#��oӜ؜:�����e1�6��GZ��^pˋ���<�iq���}~F}��a��:iʙ��ȯK89��eQ��Nj ���F-:������e�+�ȉ�Dt��W��뿧Ko��\]���q���*M�p��v�M@� o�jx�����ފJ#~��
�xw�|�M˳�OS��
up�bu��U!�v!��o�Ԫ`��d��{�A9�p�f��Ą�P�kL.
�D���-*���L'iK��z�CA�;���/R�Ϧ�_���F&8����Qr���"M!�;�ay�i�`�f���W��� �j�
=����o�,*@�|6ʃ�XBo�I��\cS��Z 1Y���t�I%,�e`����zTl�ȃ�l��
�z��8�+���; rv�8��"ޭHNG�O�彍, 1M�e+JO#^�>�
�T5v,>��%g��ϫ��=c0��<t�	Yz���|	�J$�/��~���Z�~��Ԥȇcrr��b ��dɳC1���Rz���NEl[_��l���}V��3[>���wm)K|�6��rS�����_l<���;�d)�����#�vl�=�+F`��Md��߀L�-�˪p��:��N���AOR�n?)n�y<�8.�L����k�r%����(1���̓(��Bm���)Q$��
�ل5ϰwԆ1���K�Q�O��.μ.��/l���t?�jzCɯ�S$� �=9!'�N�j��F�dj_e3��b,~��/3�eTܭgI��JZ_X��8I��+���s7C��w���M���_#�?��#2�;�㍖��oh��!�,s����
�dX�Hz�s%i�61����5�������I�
C�l���}nnh�]��B��tٝ�#�aSc���4�S��*x��@�/;���8���-��(�ua�nIߙ���g��:���;$�lǇ�/Ak�j��<�z�8��R���߅�s���/]��J����x��@���_���e	5�)�b� ��Q���t6A����4��Tf�ɰ���-�������'���S�28�zn��o
�A�"~���51�u�4]��3J�<�r���V��;} N�l���+�1�L��~��^	�@��� 2����wԕm�~�I�,1/-ʆ��M��IBU��08!�ÝNK�cyP�f�ߣ>*Ի{Q�MjS�a�l��p����4�b���&S��.�����~�i
����K'ڒ�ä���I�n�]/I��.6�si��1A�Q�u֎y�ÿ3��*-�Sn��-���dP[KG֠��b (D�a��1�e��j]�:L��cw�W»O�N���N�א�٨���[��0Ӭ�����6<$��pG��WBɁ�A�����!"l�g �%@��,\�f 4�4�<l��!��9�f�O�
�U�SD��0�� ��2�t_5 �B��YB"vM%��$l~k������Z��~p44)󽺁�|��(Sh�E���@�v	'��q��n� ��=��xx�C4�>҉>�|M�j��0L'��{y۾��>S��"��r��z������W��M.ɞ�,Ѿ���O�?��ߍ�+�]�E)� �͟�z�����v��W��kPm�T�F7���R|6�v{h��F4��#�-���lI�̘��d"F.��:���&N%�'��ݥ�}���Z���f�$Bl�=�M�Q�Lh��I])l���"�|�ȸ#�9����F���o{Zp)��	j�'���E�{��T����֑� �0S����_ ��⑅X���	��10�E�;�H�A��x�.]��J2[�6�Z��e�����=���q�� � i�ͯW�e�ʭ��\<~%��y��t�]�چ��� �h�N���D��`�V�|�0Ɖ�,B�/���|5�g~T��� F��@}Le��G��pb���'��������|�}_���`�1|�{`G�z�>N�|�M��'҃�@��yv���桶`ٞɒ�����iyQ�B��H�����[O.�0���|��d%8.k� ENo;�sQ'�i�;�>Q�� �>�D���=%~p�R�#>U���XS'	*q>M#{��CBN��0�r�R��+Me7����?���k�}�u�ydX:���_g�h��w�9X	Vx����f�� X���l�wng�磄���P5?�p�['T��f�#�<�8�Y�wfIz7���1W�!_�J���s�����-wY������F0�.��*5-{��z�!�\���t5}�����^]����.8��FhI ųyj�L=#b>���ٻe�d���P(�2_��4�qL>��#�����"�"(��Ωp3f)c�P{�?����d.�J���j�����n��ƒDJ4�D	������f-��;���YD�a�%��Ǩ��k�#�͗%9I��Ć9l�%�;Qh�^������=���Ù�9쩛���^�?.�6�}M틽�r=���^��Ъ�$��!�	I�j����&�	OGI��e�K�$���L��qL>twb���5T���O�Ԓ=�-}�� �A0sF�F��E��X����#'�p:*?n[��u���|ҿgҠ"��6.�B�_�6�ߣ"8I�F�lr~t[�L���vgi��i�9<(0v�O�Lx�l�0��D���%���I��v�J���h����1`Z�>�B)�0|Ad��QʁBx:x����	����-��bK�� g�C���|WDٚ�<&k?:�?�dP),�韨��Aq��t���[TL|��R5�茺(�$9,�3�FM�j�nO��IH��>�c����4�j �堋Dg�̒����j�l���Q��c\ۮ�
�y�Pֵ���p�4����A&��މk������>�+^���3��UG�G�XZ:U1	'����|���݁�g���.K�����;��$=�̾1�����h⼉
�E���?g6���i-fK�=�[r��98�5�v��X������Ge���@+䍝�E�)v�l��4�!~�@=�~�M��i;���F!Bvă{���e�B���&&t�T��ťs�.�_~-숛4�Jg1Z<.����Ca��"}����jƘ�k]AW��=�dCp� 4H��	�!Ī��v/u��6����zr{db��e\֣�KS+��Ӕ�;Г�8��O��ʄ�J���l�Lz���I��5��Su����U��_u'o��)h�ݝ�o�Zٹ*�7|�%��$ܘQĒA�d��v ecB�g��
�q[��8ʁ*�S���'-K �<NPl���(�tN����◎}�� �J���d���v���2>��O�"����?j�h���(벨8K)�Z@S�L��0�݇
��-�Je�Z�i%}^3yS#YIMx�޶�U�`�(��f��%�K���^��FG�ŵ�F��c4t��0���ly�:z1��q���5�h��H��,M�pJO�a�46@'L�cW��p�{���Ȕ��y0���v��&dI�O�u�o�ɯ�L�Fʓ^�8� �8�3R���x���e�xl&�ctu�#�f�`�ҋ�M��A�gƼ��̸�>�+l��I���`IS��}�,m��I<�{�˒��؝=��P�>���jB����v�7�o��"��/�lm3���<��m��C�5�Գ�Vգ��2An|�r���j�#@��WF�2~���@fq��wW]�E3�4I)��e�ɩ�耺����!rTτ��9�?�>����n��^0}?��|�ģ�"��O�""
���P������w}�g�4ց�f�N=43���ےZV��Ӯ�sey����%`�`�U����=��v#�~������9i�3g_�0�}Mx	^e_���J��\��em_*IEZQ����GK�=�eM}�Dg�����(|�Zj ����u�2�L�I��-ڈ��G�����gb�"���MS�l���� ��Y��{�
�|:��]�g�fN�"��$-�=����� ��s��&\�4�c��G��������=�РR˲�*����&�Ű�dKa���j�.Mc���s���k"jUC�&�~������?�k���Vy�%W�:�ͮ�T��)�\�gpý?��H����[&�E�v��EC��̞��Q�D��A�� ��&lFQ��I�`�tlE��bOI��[���a�9�j]���%�	��F)u���62Wk�2]X�aD�P��}n,\^� ����W]G)7�	^���~�Dx#���٧�m��!u8����\���H���ܩwC��F{枸[Ϣ��:��@�뫶�C��(��:��<u�-D�߲X�8�]��J���K�܈
�Ϛ�p��W�>b(Q܊�u���Rr�tw�D�,u�C�@��?'�?� �ɑy=���T��`�`i�K�9����$j�(Q�N+���r:�Ɣ��7Tz��6BT_zE� C"s2Ygf=�/�ީ>��1��7��W)0#�H�rj%���ގ�8�l�4A�(���ǄH���TV ~� ��|~��N�
`3����"@�UK�f���Z���nHz���
�\}<5�� LX�!�To���F�>ı�5?�}7u��J|E8ь�B�j�ei��>���O���so���y^HQv���^�;FԽX�Z�~k��Af�d�:8�[��»4RI"��p%����*�y�p�9wCES	���s��F��5��}Y��ޒ/�b7���'��+on�����U>�bC�_ԉ������1��� ��yɢ՗GmʑN��T�#�����x)j�}�DQ��ѭl�Γ�-�1��)p��^_���lj�ۆ�^��.X�$��g��B�\9
�%-ԥ��9����>\����i<�@8���2�#��=BoٔW��沲���D-�bn��K!���+����M��$�����ҫ�b��їUWh����,t4p岹�G崓��ۧ%��!�m�x���r���]�y�o]�
�<����K���	
x��Z�F�p~i�� k�M�����������Wo߄h�Th������ޡlKj�?`�Y}�(ϳ^�PRe��/{pT��*���҈��¨*���o����DN"rй,y�n�p�}�#�=�n&�'SF62���:�κ��eL�ޖg	A�k[�そ�3Y}�om�tTX�#��76�* ��b\�\Q�ӛ�?|�O|)ʰRB?0H/"}���ԡ�����\�2+9�E:�I\}���i�)�#֧��1�����DdeE��z�ƮdaV:�mg�o}���~r�畹�_�&n@Wi{t�3Y�� �	��.�v�WЯ�M� �²�O�A�A���]��	��x�lv�@9z���:�p��m�e�5�$���1���:�Rd�kjg����Ϻ�	UOw�Pâ���D�:G�QF��ӛM�Ei����wڵ��mˆm"3���K4�/$��yM\!/�*������}�fɳ[t�F�!�reC�5��r�#��+�
kp,w���j1��2�6˾«�� ǆ�%��NMI�K���{��B?Z�a�_�Ƨ���FX�u�X�}s���܊�١OWZ�;���cjpp p���� ����M���[��C/�r�(w9"�a$���%d��c.�}m	?0�X��S�,c�w���0�|���������3g��т7%P���7�,�j]��2 7јPL�O���tvv���/�����#�n�Q歉�$V<e�|�)/ټ��l:�+�O�펆E�Y��jgC�?0��u�B�Ǜ� ��X�7�ϓ4�!{��BnfΩ|�믜�R�4t�_n�B�멷��|o;�,�G!���U������<����DD�E����B�4���'���6(�V>���G&�M��c�-m�^}-�%p�tl�/0���A3�Rj��q�HQ��㸋�M��P�Sx@�ݿ�r�X*�F�Wi���½�X�Bkz�����7h�`0̜�r�V��?܆!�E�~��Q3���l������������4|6�]�4ҕ����-��U{���Fh9��R�qa�� �}��a��a�{L~;�Z��5έ���Sֈ��(�Qd5k0�#�W���hU�[$-�?�S�c�T;ѐ��\�<EU�Z�5`�{�w��K���5�F���a�T� 
�'��7h�4�&�z��ڋS�H>|U����rB��[�K=�Ļ�� -k�ab�G�[��Uγ�A_�܇�� ��VrU_�5a���4�z����u�%��ö��]3�WuYy��4R}�c �Dq�7���!`�̥�ی�����3o^s���;��*��ݜ����@�dP��"��a�K C4���k.���n�;��6�ŝX�"��������ט�&��U��%�()���i9r���c&���(@�����+A&�ڬYt�,�f^"x^���Mɟ��gy,�g�s��)�a\���$�!���Ԝsy_�0[����
��n ��l�3M��g
^�BF�1����g����2x):&��U���+�(��g���g���M����*!z���j��! /P.������&'�|�4*�j��݄S���e��.��R�T���H={�=&)�C���lYaU���d�?\�z8���DG�9c��kyM��w��V��}�Kp�=��9���>gl5�����fEj���d���jJ���3��~`ď�Xv�Tm{�Cs��smF��R@��D"�����M7�����!�T��wL����v��Z���8�5~@�	L����g=�!��0�%��P.��Y� o���^�����<ʪ�A����gd���)��S:`��$��k!˚ӈ���l���a�I��3EЫψ��p��C��?��}Y���@��.?bN���۶|̟��Lԫ��1����dL 	X=3I]\�9OưR�=AL�"��U%����a?e��dN�V�y8�p� @o-&Y�Ҙb���ծ@h4�u�.�T�ف��J`���o���۠E������P�����\&�u�2,��\�^��b�a��;,����	iK!���e��A	V��V��aP����¸�`���P?�o�;�SQ�.��s4ؕm��B�'3�o�L�ޚY�ٌ�����!�%!�x�|���e�s�*W*d�+��'����*@�S;�2�G?ő濣�Pt��È��v���n�<j�u%sv�g���TK�w4I���o9�r+=Wb^�ӻU��y۔܎7��o�;����:{�|\kh�B���l'd�i���?C��H���Cle�囑Z{%�:H�ў��d5MP�FuũPd`P{Ѣ���(+Oz�Tf�	|����C�����gOb�9��Nr�'���X����vEFr�{9�'h��� ���ЕHQ��;vIo����Gu#R�"���qyN9���=e��wY�馊���Z��)�������crqM��P��fV�K�{34i̦�� ջ����C�3:�>��f��`����1�����Z:Ωr��O.�g�~v+�Y?Y����R�:��`	��u��-r���8͂�m@��6�w�]5$��;F�����u�lCmAC� �f��^4��_�#��%c��M���e2
^����f.f9�gh�S)����P�Y+�=�����ك�	1���Qj$'���8{�F"Ąd>#��IP��Qw)�J�
��w j� �(�@�3UPK����V�� ׽re�蚤Һ��`�>bS��r�I��i��<P�(�w�&k��x*��
�p�e�k_����G�2d渰`?��Fu��egMw����X�������R�D���e
���
���R��g���d���qU��ʪS�} T��A	f�U4؎!�6�Jp!��/Qdx#Ҟ�p��T��r`�6[�d�R�:�����(F���̗�,��|�z+�b����Z��i�h�t�|Ɵ{c�T�F���Q����׸ȩ�"̫��ס��hpa��}r�C��T��hp�,P;M�FɶY��C���G5�C����p���Z �5ķ�����%�0�q����u�FI� ^!ݡ%8��;�L���Lg�ٿv�Gq �����ub�%>7�j��������H�0��}�~VNO��V�'�{Fʕ%o�o�f��&� H�|�\Iq������S�(�7���(�LLa�-����U��|l�LӃ������6�«��΅��Z�2����+�h�)�K��hy�2{2�Gk��<z�o�lf-��]�40Ү��)~�7��+���c�ǳ��m
�@�L�y�������(<��Te��+�8OP�,����P������	B2KY5b+<���{" ��.8��)��ڔuu�MdZW���d ���b��i������
���v�6a^@�4��u��uE�YwoC�)�b��u��O�@y��Ku��:7�!W	��Dά�|� 9>E���K�Bz0T:��!�Vk¸WGn�UP�y8�`3� ���]����+r���V��-����x��:��JAd�"�}Tc��F��DNz�YZN��g�����+9Udy��
�_�:��ƏQ���r��� ���y��5�㠑��v�r^I`.s�2ܱ;����	e%f�Y��8PI,�y�~+5�#�O�4��W�ǰ�1�}�d]�a3�;�b�n���w�黣+��[	*��m<��l�BG��nvq�>c�桺yx�'�fkl^	���g'���zrd��$�f�Ԉ<�e��D�֑�R`��Z`o�K�����q���p�L��H�	�@���@a�G�����s ���%H|�}NX�sz��]�#�֞��RI��O�%���Դ�x�����u#����<�F����x�I/d�z{�L�$�P'L����9�bt7	L��;I(���օ9k���r�cp�Oih��}^:	6�ߠN;�V�_���x�r�­s���qgY�&nZ�;u����HN�ޤUeȆ�P�ў��g�����y�?���rkG�Ն�;��mv��*�uw�ͷd���L���#��(o����_B+���$i�We��8G�hl�|C�,�tW5%��4W�Q1z�K)%h��;��&.U��'Г�Ɯ�(*�߉X,v��_ P'�sө�}�Ɓ��s�͇I{ڹ����,���LY�^��y���N-v��%���+�[���O1?��'�T^���
0P�ӗΫFl�7��<�xR�E��K\?u[垆0�yO������䧒3���亸4��˵a��pH���蒶BOqo�i�΍y&*�� \Hʖ�m^���9�B�6�eI��R����Ij�[��������v�\M����GAR�h��w<�t.6�%rYL�D��U�zUFy8���# �Ԅ`�L������D�jWc{�V�����쬝��1�yt���P@^L(����8���NyQ�Yr�t�<��z�#��k���uE�]�5��W\F��8<��Ŕ[��^JH�]8Tt7�Л^���!�μB}��w�.��許D��`	E*!��#���� Gy��k�5��ҋ"+ t�߬�)�\���~��Y�4N������ ���~V����)�u��|ml�-�ݿb�2� ���*��?��iL�L �{�o���_��bC�1���ҍ�8*+ }z�L,�*Y�*�R�~�L��v���wG����/9z.7�mjGr��u��(6��
~	�`L�|$�;� �����u`(0L�L.�M9�[K��C5��9��y�E��ض?0#k�{~\t����;Ģ��0��1h�ی�d���'fl���E"{`,���2d/q%��WO��[��q��̎p �j6_c|�pg���B�Y#<X��k3�b�/��*���!��'�*�"��_�,���h��l|~Ȁ��21m����~~�J�.m{D��$8������h���7�h
�����ޡ�m��]|�O�S�m�#��b�rJ[2�O�OٕO�oԮ��4�	4=Q畮�����Iê,L�
6����)m�g�I�u)���W�k����T�A�jy"�'n[\�l���o^9)��AmT���T/R3��t�~���\?��AJ�6�p�:�rg��7?��,�zV�=��$��˺Q:<�+�F���d�������y�H��Hq^Д���Ȍ�F1�� ���P��a%�,�2�AЀ��.K�O6A]��4Cs�+^?���
����
ތa�X�w� v)Fm=T�#�JV�����-F�o5X�P�`��]��
M���w�~�>��(P B �Qrí�TT��\p9�*3�ë�j����O���X녈�+6��l@e��%ȷ�<�N|2Vy͉��TӚ'zҚ4��3��C�>-z�k��3/�:���x ���`κ�Cl7��3���+j�c6�(Sa l�EJ/�อL���<�0��`�Ma�♖�S�N�����Y*�Q�v����<k�xƮt�#nx���M�A�����~]���a������֣=���T?��\e$Ԅ���p�{'�,B�u~>'�ީQ@�����Sye��ܨ輨�܏\�d�% �����v�K�UhƏ���?kc�X�^����u�'|�����A ��p���y��͞u�.N}c� �$Fr��@��<v<��3���l]��ؾO�鼸W���T�	_�ܝ�8V��a���ap��]��~Y�"4�k�����W��&U�k��ʵbw���d�/R��r̤i�[�3%��� -~e���o6��f�3�`��[�0��I$U�zm���ᡊC�7�Q�_��T�梅ڣ��(f �Q�H��bzT���j���]�L��0�?%,lCNi�*M�o�K3A<�W�\�MR�����X�/�Ϩz�ă�P T�n�vipI&�����䝱쵎�c�=�c��^ Q8',dv�������ֵ�{*k�g B�I����_��WR��ߖs�6[�z1� p�͸>��."L�Ou6�k���Y�dG�<ȋ�xi!B�n�����GB�k�{��4������P���1�ܼ��Z;=n=�5z	����d]^��ql0W3DV���D���Hg�6���2s�����ϑA�.��fY�~]�����h;�Y�b�h�R�L��+x�#x�b|� q/'^.�F�!�ڼ��X<�d/�FP�wx����֧C�;�:t\�&���H�#��.��YJu[��ҕ�����%�vy}�}���ΔJ�FZ���-y�Ièv #�'���c��Q�0�v���p_7nTm�S7t �h�"��k���q��_� �Q���f�
a�~!��ĩ�o8^��(N!�L(B$0cƍs`Ϛ$��F�����&�l�d#�1c�kց���>&�SQjO�B^�A�%������3[��&J���4v��3���:5�=�=d��� ��N=�v��'�yY	�y�v��K��SK9
\^�Õ�����}=��eE��i�5:�a��"�����_���B���C�e#-���<U�.?]�e�caN��]�H�I��`0Em?m�����������?�q��Tvf(�'h��rCajщ9D2����R���5�[�����I���T�7�V<<�*�Z<	�VT)w�(�81w<\1S�V,����iL�AL��z���c�!������ֱ��հސ���������[��Z�ǃ�FY�,��Pu�,݅<`A�<��"(ι�;L�\c��p�1�"�3� e:���H����2�xţ������!����� ��rt��M0����(�}���?�״��ݠ1�>`��W�C����X�2��<2:���2�-*��f6�T*5K�1bQ����t^}��������+-Ľ7O�L5����eaɩ�g�ImZ�~v�^~�g�4Z-I-"m��+f�V�B��A���1�>�r(׍n�ɱ ���5��*2@pe�ȼ?�%�C��$�A%&K�;M�7��`��A���ߦRJ��>���h7!���Az�a�i�ގ�Pvx�M��9�YaAG~����.� Yu}�ZP9������i�X���bU�Yճk �(%��˥|�9U��J����ZvI�%I�YL�[��O�슼c�)!��*��N9%6לB߲�Or�+�4��L�N��?�E��lӶd��˛�6�Q_p�efq�N��^�¢@P�9�ޟ��AhyDŨ�Y5�-�=.�'v9�ʨ�?�F����:9����S�4�"�.��:e������o�,������m�\�G��u�HD�	��7�y7�@�3.���Ihʯ��x�00��N�=S�Z���ߵ+��]4�O�:
k�Rr�Q���E��~����xp���=Z9 'և�}�ƕ�I�K��R���I�47H}SaS��Π��.��o�x�ݏa~�
����Y�c1f��e�����Pf��]�%(�J��b-�4�}k���{�����?���c�9�,L)��	Pي�2��uO1��u��ƶ.3Yt��Ԕ4�N��Ԫ�yȴLsjx��(�P��Ĵ �_�ܹ�=$,Zl!:��$y�����)7��(��z����t��A�ʫ_.%ݎC�e<!a�Pj�����L?��_]��{K��$�|��9�s��D���5�ye�$��۬�x( ��5�D��!�$B �ѢTo[�s=���9q�*߃kBU�	�N$k?�M�)#�`%UsO󌷰%{6 ���`����&o0�W��Mg�hiG�늪l�\���Y�)(�S�SRc����Ԗ����va�0�P����SF��!m>�U�M\�K�u������.��e욥��M�EL�б���HE�C�*����q�qGm����
R�_��{� �2i5/F�|��h�|#f �;/�Q�^4�}�{w��9v��5P���:
�+n�'��ӷ��BP�����^�Jv��$g����������M�����Uӆ+��]&CI����Fa��.RVTq�	�H`@�W0s���[B�@?��6kX���=��8�Jl ���\o%�p��TF��e����*.8��A�pG��¡./��B��>����ڧ�����U����@]��Rs�$�J'k���z�i�y Xl������T��E�A�C���0uP��j"�X�(қu\���_�MA�VH�L�0q�dh�l����������擲�)���7�әu%ā���zB��9��[�f���XZ����H?�����l�ko:��&��t�ޒ\��!�N�}2�6{r����h�J-F��#�H�p(n^��Z�
]�e</����Û�!/Q���4۔�$�*�z�%�����t�:A���Hr)�������>+�;F��D���;cb�*� ������ :��$�\���r�iy'K����o��\� rQS��d�ZF?7o2V�jHA2�VAADyϾ���\	^X�N��5ԋ[颋Rs����ѯbnr�Y�YQ=V��RY��[iϨ,	O��=���]�a`��F��]��[��b��қkT�{C*�1�z�� ��"	���� ޯܯ���%a��95��M6�m��y�a�KXdk{� ��`P��l1Z�&��'�v�|P]/�Z�����D�ʥ�Twp���q F���c�8Ҏ�;�@�5�����-'ݛ=��/�|fЕIh%�֢�o�w�J�X�tF�#�u<�dp�ev	��4��ڷ���'¾��
]�w�U�����\�/Ż��v �,���������L���2nu�JwxΣ#�j*����m�W�4.�<��`�K�R��[���l�L;da��I�|��^�D��������Ho��n/�϶|��������2���*����M���BXBS�%��l���-�Ϋ#��{����v���9�IBU�|�!�������߮���~�F�
`@3������D����"\��?����[�����v���`i��K����4o�Z"D���4����I�vQ���&�o5q4�������?T`z�8#����G5�ɧ��9 �9�U��!�m�KM'6z�����J�i�@O�)a�����;3��Iork�L
8���ܶ�ƶ@��ݫ���`��
�s,�&Ȝ�,Y����ױ4pWM���Y�,ʕ|���C�{�/O~>ǵ��|V��K�I�ϡQƢ M-F���dD+���H�.?�q����m��ޖب]'�R�d�;0�ۺ��2 ���/�����+��9�o�n,��W�G����ٓ1?N��O�_k�Ӻ#�qJ��Uӵ�����P��-,N��+��y�?ΰ$$�e���NT[���Tޱ:�k�3/�(�)��~�hֱ�}��l�F��ئ8?h�[5ʸ]��7������O��H?�iu	��|� ��'�U���E�H��0m����k]�=3�������\l����������P6�|�H��}��I�4!mW,¨@��ހǡ���|�H��	;�wS)�F�&�F��`�a�&�`t�	�ei�@��	�W�~b>��D&��5Opq����a\��E��	�@c�^�f|�@P����>
�L�K%)é�s5'Zl�ک˴��ö�L&�H�`B�Y.���$�a�|�k�FU6�Q�V�ک�����I���і������R<Nf/~�	Mt��G
��.D\Ϟ�| ���� Q{�y����?�{�>B����Z[��v��~y�l?�E�I��F��>�1ř!EZ�GMƫ_04u���3�/P���2幻�j�
o�+}�[� �p�Z%˩h��ǺA_X�1�3���Ҹ�{9�qثZt�����w��$(G��(P���#Q�rE��Y�8I����0�B �#qS��i��~�b��zJY���x������~؛��i�$��S�ӭf�Y&>02��Fnl��(v�n%8Z-�z^�3m�3���̛X����:Z\��i�4�p�%9�Mw �s�QS��KV.��/����p�֬�C.�N=�E�(��r)tF�h��\�; �w��c���cuQ8�	��׺�%iKSD���e%���pȁ`�����.�O�ߋ���!)�����IGվ����U#/p�>�-�.��y��{gw}9&��M�r6W�ni\��E~)
Ǐ�b3}�]ks{���7'l+»���w;u��bi�����{�h����͔�a@j�w���O���g���[����܉�/����"<\���~�\iu�T���f+��������폞]��L˸���G�O@��:c8<zg�Z�az
V;�HcY���\:�)h�y�M�<����ON�p���P��ު�p VB��Q�"��s2<�w&?��P�W����R����F\nb��w��u�b(}���O$F�b�c��Lz�m�"����'��jIn����Q�-�B'/.ϕ-}9�2OWP�ΜV���Æ�����;dꧫ�� jC��P���hNy�
Ϙ^�>��N�(��H�u���3��C�W��&O��D�Zm7�>��b%����D���s�^���A�����|0>/��b�r��)���Q
=ɻ�#��� a}՗7������i�\~K�>��a� �U�\v�$�X>���Mݥﲇ����j��O�d��.i��A'
*I��������Ř}t^S�W��Zn��h��6q�Y���+˺ �����"�j�ô�����'�����uo5��ϒt�D4���Z��r>��4mW���S��|-���@ {L�g�g��U߶�	鉨��R5�X��Q�Q�a�j�����r0�/
S+4oA���}� S_�����[��������:{��2r\O�F��Ke�r���>�C�H���λ�s��N0��9d��Gބ�.��ip#����_�����8���(a��M��iC�s�lU�� ��C�pBM`�߯^�s�y6j<��AU�͐�%��k����>�� C6��GlT�zٔ�|㺔�!�ׄ�� ��&z}m��V��N���i`�Jq��l�Q���$��ĳ(w������H���pԟ����sa,S���2~�q���� 9N�|��\��}����l�D�nl<�o}ڴ�Bg�a\c�j���93</�3������P���7�8�64lXj���ܐ6Q�k�F-Ha*%#�2�$�����=y���|>�;1lVgfDb`K�9!F{
M���)�����㥁���d$���{Ys��1�P���]^�-rK5�	J����Ra��t ��$SH��^��5��9�T�IZ"滋�����ՓM��f�F}՟M��'����B� Z�{C(�	؂#Hⲏ^���5��w���Y�@ZQ;���T�# D�v����r�䍑$�e�əeHXYA#�9�!�צ� o��Cʴr��J��s�g���.�Ā��=V{�Y 
��|�-*����u�u�q=G�M�5����D<'G��F���z���,�a�mW��r6z �ٌ�_�~�,�Yj�al�Ɛ�.l�����Z����=渃ȣL����q~��|,�p�������8�C§w0H'ƽ��� �E���מ��h'��EJ��Z��X��r�_j��֚�iFf�$vq��[`���n�\�Z��L�
Z�/�3�N��yԶ�Zt�
����	�1�-l
E��z\��;�`����1��b��&�ҕWɞ���O�� ��K�P�����[x���+ԋ�[1��k�1�t:�a;b3:Y�j��z���<����r�d�#�lPtTB.�Xvb	>j�ue�9�`�i,#�{�{��N�5�����}C~}Sx���P�B���av\��VP�a���0E�����u�h`�&L����M?'��ex��ӹ�NkI�#����$�p7w��Y���?�O���3L�+fl�`��g-j���h-��*��D�1u�Ѓ�O��_�����P�ه�e$�L�����+�=W�g���ܱ���da>� F�`��`��6�zXY?\�S�|H�V�-$_˫J��+�^W�p��#� ̴h��Z�g���Ƒ_Ϭ�!C�r)�@��Ø��*�:2�fI?��I��޸�av�d]�H���l����T*-F��D�L�/D�����n��3m�֤Mw��g	S9Z_T0���d��>YJFǨR�,�O�q�->��q@v��
-���8����fzC�Oa.B�UP��ڧ��"�H	��3��(T��!�+T���&�ke:�Q�>�S�/O�'�Y��!9�o?���lT�B��8-`#yB�\H�H��2�̰i�� �����teQ�x�����ϐ �0}��%���� Q�@P��W�c�BR�Ƽ��� �Inzl��@6��,-�?���ll<wo~ϝy/z³��.�����s�'�!���:Ճ�3�`�{�5�ş~O�>��p����H��Ys��9 ����Vqe5��x�\,OG��|}v��M�h$�M�,�3��U�+�aw�c�	Zo��+�����B�������7:@�8�krHg{�#x���K�fc�gyscI#G�F��fU���fxU7��J��	Q��U-"cu�s����vS�Rs���x	��O���3G>�ԗ������
ͅ�#o"j��`� 9$�����P�!�j��dhi��oru]�q7П�.U�%����W��E?{�f)s���\�=������H~�Zb�*'ן2g�\�{x?�HH-#9'���~�Ģ��J,\[%�$ �nb���]!4|�Zm�d� �?��Pe��I~zl�yd����"�J�W	ɂni��6�\1��TX�=��F��'��-�V����q�syS�a�Q��t=�s+o�b([�=��h���c'��U�=���%���D ��2��؃Đ��5ɒ$�p.%Kc@5�idF���$�:��+uHҖ�{N��Z�Wbߎ@+�Z�S�E�P�-W���c�y5��]t������t����U%��0s�+�����d �����4ڶiο �Y|��fB)!�����x$+@��(҈�a3q�r��� /���f�$|�eV0/&$%ld��'�� ���:�T8%�z6j��3�n���Mb]kvw�H�8����T�:�{�XG6����!�:���k�n�s�څ	�'�0��;��˩���NDL�ѫ��+'����5-�����W�i[>�Z��_}���G�Lv+�-��A��3�p�yD��?z�8u�B�3S���� �����B�P�yo�C���	|Ь�Q�yU�$�X��}�NbAһ��w�S�<�`�+T}���w9�g�vd��\	��y���ow��� ks%)����D�yT�,29x�d$�1�S�}l����r�����D(��k��笉0��8����h��.j�B��~K���kfK$�ٖ@Pӡ�j'��3�u������@(��k� �*⸒�#�e��Ƴ[e�
�<���8o3-��G�eN:��� �E���Om�.1fl��2�	�+�Bm�xBA�8��2�d��,�3+��d::`Y|��p���
�T��	7�C�,�E|�0���X��@,�^�GrG�XPSU�=���\�{L0e�FY,���u��K�m��^X�T��ݏ>u�ol���M�a发�Du²Y��?k�<Y����}�.��uQ�E�� ������e���q���I�ẉ��<����x�zd-��:0�"��S�1�!E��� ����\����p�/M�����^w��\'-f�i[�F^5�Q�-��W9�"���u|^�:`E'��@b���"`Y�֨�=����څ:l��H��6�3t0Aks>�`�P��Nj��~�h>mx��VSL̨,�`�x"u���iވ�Pt��w�S��Lt;�ĝ�r��ϩL�Q_�Ke�]���>lg�	f�5A��L�޷�@ޣ�%^��$�{$[�l����Ɛ{�TZ�w��zS_��0��1sc`ť�F�1A���G/C�OK��<��+l��w����+��6�x��M �Fe@��p��n�/��͢���*�>������t��4 Jc�Mm�s>r�`@�G~x����9�)l��	y����g�8��`�O�^
}3�y�x[S�H���I��9CӘ�2�23ӊ��ŒU�:d;���|Cm�Ȉw�*��3��Pe~6[I��D3L�Q R �c<
f�������7��$�*��'zREb�����_�Ĭ
XW����Y4%���PO�0��%���x�$�;�r��X�y�.YB�;k���s� ��Ey�(LT��tP�G�P��	
;��llrq!�$Qi8�:5ߍd� %�nI�@ԫ�������v�f��&�>&1����MFU�UQ�3�5%��.|Mh��s�zo��f�h���.�*�`RP|�>t��WJ9��;�n?��� �p�x6eo�1 �����jU��������WdS�� �_��>�U��ɾ	K#'����Q���'�"�çu0R;zq>��X�KȰ����d䞐�.���Mb�r��1�n����Xm�8A����\l�W�=����>�!�n �tJ�A����_��
5�N�|Hd3�R��U-���W����lm%�ub��O��B�lO��'�3v+ʕ�����?�݅y���-��D]?��"՟R���|���7���hS�8)2�,.���.j��!�1w-Y�
������Qo<ߒ�*��jr|������*�����=�?����(:�4��9Y�B�����Q��>������Y�ۛ�u��Ǹ�Ӕ�(���:xh���tX6�����SW>��06s�Z��y5�u�k8aXK���F�	\5B,!{u8�G8�����gJ�6@����9�DMUW���5)���3�%S��_p��p&��J��y|��1�m��������ʋ�|�ӫ�ՂH���$�:���>����*Z���%c��)]��83�a���q���ˇ�nxR!�®��
B�0��E9�,��#Y^�"�J�޸f��:�����p,�R��<���5a����{�^p��[R,�������n!ݏ�^��:H�?ްM�,p[%h�ˤ^$⫪����3���x*�pJ�@y�[rnD564a���fn�A���GL5#��g٠���B/��w�ӣ�%D�ۮj��T�J�Y%���~�$^���5�я|����޿=�3��O2UR�rx�Zұ匔����p�o�  w�b�o7y��!�U�ZN��?�٨9C�gw�٥�Ro�?�}��m1�F8����/�Y��BЪ��+e��0p�o���
S��ʯ�MӺ!;� v��W��5{_�,�R�.x+ $^�9�3@�Լ}z'lp�֒�� C�2�m�#�f��UϏ�����}9�c�S��$�teM\�����������C�e��� 7N&`����b��s܏���j�����8��N�ʐ���"e��%5��Z?8��W��Q^a�Nr���w�
Q�F'���D��K���&C�9��kE����L�?�W��1�N"/�.��S)�U}��A���C8�X.Pǃ�,/FVUssD+�V5@re�5�Q%֕�P`y
��0����Z<�>�aۭ��p�^�_0�q�v��!�+�s�g.j�h������lyG�k�PI~��R�I���rƻ�f8$��|��@(4��sS�R
�e�K�J_kSڝ���>����D`�g0c�ȸ�d�Yf��ݹ�vj�Z�{E�#�ݍ��-�B�v�%�"3�f=�(D�"u�M~0��WRdw%2]�eQ����5��q��&{da�{�"Y���}������c}k%��N>�D@(h`� .�L�"tC�vmV��ߣ�2�8)W��D����9G����g��ʘ����g��Bc�.U[J�RG~D�����������I�4�0X�3���uN���Tv,g�8�a@�n������_�r��5�X�	����������W�ɠ��/�\�^�E���*3_������\�!ߥ>�E70�I�h�_G�]v��`�;[�z.3��]_��?�t�os	��+7�h?�>������
����2,�UH�4%���\�-q�n�HI�� ����G�c���`B�_�(9jW�s�*c��'-��##;��:��'v7��m%�k�����k���U�;2�Ł�-�wۅ�@�"��V���x�ӂ�YO���p�o�d����$ �u�2�J�*'	r��n-�俑惍�1E�TXY����[t���HU8r����;O "Rc(���~ඍ�(�Ԛ#�=�B�Ah���b�pP���s�% ��`�&�Y+��ѩ�_���8@���%�X����[�!=6��z��K�S
�h�ɖ�ŝ-�{n�}Q�W�p�uf N}.&�Jx���`#i,?���7���b+{�ͲR�B5�W���{E���\sl��4��2t-̰�Q�A�H��zHUr���yʃ:
?0Lp��+K�}P�,�-��[�#��+�~�T���!�N�ŋd�[�����nibU�OϏ/�y@'���b�i�p)*�{; @�Pr>6_��R�������i��ߊ/e��+v�H)�mR-ԃWzP��A9gzOU��I�Z&e��Kd�yC�ϣm�B#�p,
��i�X���f8�:=���\�'ᨶ�Ĺ³S����Ķ��մA��,jTCQ�E:�P��[�����o]	469�ʾ�u��4�ڜ��Y[���\�V�W2d`��R�vΓ�����M��Q
��i�����MF!�kGq�#��Kt�t�+{��"�cy���}c���޴�w 0�.B�:�JKX�����:��=P$>�����vr<5O�����on�}�ed�:g��(�6��X��Zc#D}�遶�y}e�^���	�\���XnV��1����%��H.����ŧbZ�]q�&�c?ԂQϯf����n@k�.�v)��N�3�)'ғ�P�[6��G�	��U�pnS��]�C�u�eZ���F]�tl,.kc{�P�]RU�+��mc�zHב��Ӈ�w�θֆ��m��ɫ��8�9,�_��[��s�PZ���*��3\�9&U�J�0xaBy�ʆ��W)]^�1�P�n�Ӿ��uᓻ��.Oz��;���;-�"fO�aW�O��d�[��"�����h���iyJ�;p�R�`�I}vļt@|�8t�7�J;�s���I����q=��h�e��9&���`l
�_�>*:t�ӒCJRC���U<����|��h��;�L��@��Gi�yKռf~3�&�'(�P|�����>Y,��t<�Ą3��d�G��8ps��.��n�>��tz���P0C�iи�mnXjO�b�� KE����.��]ѫ���0g�;)��*z��z̖���!D�����?���2��-�#CH�n�s�H~<�������|���8�W�~/=�\�L���DVŠmc-3�ns��L�Zց0� ���*�/��n��:�W�{�6�~yBm�0B���>O��fY��<!(7r\��0M{C}0��+��sg��f�iX�[���QY��*�ӆ ��T�D�ϳ�J��g4S(��qEp[��>�N�ِ�U����/�ʐ�8׭���D�5M���b�+sYS�쌛�ο���yk������1�.<	���Ki��B�#�D�=��r?V��������d�\ V�*�G�fg�H*�XO�/͸��D��.�����p����$�
�x��gX��(�����1
�W��y�Ю�S�}�'> Y4�s�Px�\���f̷õJs:Tͧ��/���.H� ���i37"o��~H�g�R����_C�`}e����%��� �)��Sd��,�^�_6F�9�nǦ�_�Y}}��1_ۍ&�9�8��%VUR���d���*�P�$��_�t�]+͓�0����j5,�����0y��C�Kd�� >�>�=��2Q�g�to��cl�V�u-5�c����0�@0�`��k�L&$��'�T�K�*r;$;��9�4cM������L�zzѲ��T�e�'M�]+6� �	7D�ؒ��9]"���/I��#���9�Ų�'�����������Xq��0��^��-/w�Y�/����B�z�AʂQ[{�)�'P�%E!t�� a���+��w��Í�h�e��|,�:�{��ާO�;zDJ�`Ӎزpd$n�?~ �I�5t�$=��A=��.&�f~�#� �K2�]~�'��e^��M��͝���r� рC�����s.L��_;R���#���i(���1*���B��~h<N�ΉS��ɤ�_����y��aOx��'�Dn�+�tnem��L�xL��:)�H?��&��rn�~�.�L$�x��̒w���%�O��z7���A�w�l<�\ʌ���;;�3^�̗Qܫl��\�����0ʭ�h��Ti��VbǀpX���J������&9Qj�D˴����[�C*��'8����y)fL���b�Tj�̃J�o��f.i��(�
�uW���]}�$1�(�m��+1��qN���z���wF�m$��%{��3!��v��:�Uڬ���%1lX��D� ����!��^�oy!Y�0�f��4`;뤎�,������jjIo<������x�p�)�P��=���ʹ�Ï!֜�삣"|��\e{�[U�y��ٹfX/�cHv�@�����s8+3��ɜ�#��an���w%��A��R��w��{�|I�Sg8����ͪ4'���(����&��g��1�L 竊�����
��-6f������K��U{�Y��֘a}|fW�)�8 ����gwk�6�ϊi�sk[����8��`����q������;X�����"4`�����#��T��ܡ��D�ͳ�~�wХ?��!���l��p͊D�E-������\�=�O��R�ڮ��>�n�c�iŁ��A� 8A������v�#M������g�Y�-���r�/���'K1�w��pmy/}7�Ȼ\] 0��0�ߧ����Vr���6ٞ��D����5�dw��s�[A�u�u�����C���4�2���l�t�h��你A�/w+y��ljW����7�;+�{�2�!��u;-Q�zUM�?%]S��b����)��Pֻ
H��@mOD�04$J�dГ�v�T�v��p.�\@)n���R��Z�@��=p���!,�o��3pq�Z�� ��3����Z��
I�C6ց��������&ޏ�Ҙ��%r6s�ߙȳ�3��V~�ו8����̕�+Ѹg��v��&�/����7<p�=��5�{�,����&Q�7����"��Psͮ9 >�i��}E?�������<��؆���.;�o#�I�~�-f%����|�x�$����T�"� A��U�h.�ґ�[<��0�vX��oP�F;�*T��hM)�pƐ�Y� �vИE/�6�a��G�C���`}���I�����a�mp�Tx�ꈨ{�&�d�h�ȱT	#����.���i����Cg��ǁ���&�������Dxi��_1�.�����B"X�Ct��bO"o�6��YFEP��*XYnJh(��\�o��	����H.!��2�6R�p+��Ppj���Npp�Ǭ��4��5�ފ��!dS�I����CS߹F�+l6̧YݏV(���T*o�PQ��d!8�.V��wt	�H�9�>��(��
��@�f�~Ω>�ӉԑuIA(V��i��\���!��C�H}��x���2�1�} g}��v%�z�ʅg�o�6��aty��"�GM��z�t�k���F,%\��?�o����0��Nܙ�H���X���đ��Y�e7��)Om��vlLi��=put� ��i)�)�8X��p�]r�H2Q$��$�S�a$ ���a�^�	a!�	�r��G[��/�5Rp/%�]3�z ;�=%UNWF��J�����Y�ct���Q��:U�@�|R������9�S��^�������~��޻ޙ�Rh������.pE^���p�X2��x�l�`9�.Xbf1��2��X<JGN#�	��4\���(�K��[�Cea~�#}${˵�"��*��z���WP��3�͜u�Nrw�����*Ӄ��E>E�?x��HZ]K�&yE�6c��lI��d�#�+D�-���q�[:����<ĝ��s��<ʖ��+ }S�8�>P�,�fL.�|�Z��ӽ"x��@h�>�:��#'�����n���Y4����/���k����9�m�y0�YPM�"�_(�18�"a��_4���ß�������IxSh���Ã��/ߚn.�(�� [u�)k!��zr�L��p�_����Z^R��p���jj&HY�������'n�uuN�A�M�P�ϖ�tx��,�k�f�����1Q�(X�X�Q s�x�%��4���q��%O���"߾�a��K�!@�ƥcq";4^G��Ch��w�
C�a��y�����3��
ez<kd��zv@R/ȮP �U�~�����83��!���@����~{��*_��g��[u]����c��X���2G�C�;�qM��c��ٹ V���{=�Ie�q�&'� ������Ò%K�D���<�k3�r/mL��zΎ�s�!��D�rg���g�$�f�m������*`��0�U�#�K���S8����C5Iot��\y_Z���u��Oqw{ϐ���ݏ��ɤd]���w�!X�u����f�,���֙&DC�8�:��� n)R|���1٭�Q�9���a��ï�:�)���T��P�W�د��7���M��vn�?�R�� �"?����!7 �1ڜK�[F�dK�4:j �ͮ�SHn��e�Zݪ鲪f�2Pmj�����Y����[�`_�ǅc��2O�����Ep0�Ifh���ϓv+8�^�xjzL����<�b+��bԀzّ�a�';���_�u37N~I�^�:��� \3�fu�NFB<F�C�9��!��Jz0 �G�H���+�ߤ�
:��|�o��fA:N�\���:���]�$QC�tbtk��Hd"Q����'�.x�^�fV�Xv��Ht�<A ���z��1C�lN���q&�@�7�n�&�_]�1���0�'�|�<�4�a��t�`�}�S�����Z�5�]��t+��=�t�l�di�M0�����e���j�����V�D�@$(�s�ʶG(_ƅYV����%01|�v7Aoe8_�ۭ��"�
��3�в��dM��M/�`B��c-\`�
��e<˩���oWA6�v�l r�v���rZ4τ����(���*YB?K��UDe�@8�y��pUS�o�/"��&jG�����	6��]�uQ�Y��߉�c�Ή�is�@�r�jqR{`��@/$�v�5=@�]������i�r��j%[z�%}pȫN%UI �$���c'��,<L=�2!X&j�3ו�X¼I�lW)� &B�_��k���wH���Ϥ�����M�P�x����K�o*2��%��a��?��Sd�\` :�L�z���1d�&!V��VA+����6:�[Y9��}O/�3�J����: �:o�l�{Q�L���$�i�[�1!)G5,�s�P`�6ʃ<����&�C��X"N�h��73���>�o��r�w�L3���;"4��f���R�t��]����n������{<��0�Quf�%�-*�Pi|ݔpg�}VR��pe����%%��y䉳���8BI�!�fU6���-�X�����:��<�w���uzy|�(Ĩ�]������aP���O�Pb��O!Wge�ْ��zQ� ���o���3�Db��7�Ax������Mm�4�`m�橜?�6��c[Bٛ��h�"�!EI�=d �7��ߦ0ՀP%m4�u<X�?'#;	�@�=��t��tN���Xs�dE�U�hn2t�j,ǡb�.������]��bkZ*�����V�\7"�F���\���ͪ�	۝#	ㄆ��h��S-�	Y��)U��2�Y�U\��G�+6=��q)! �	��j�D��I�ǿ�ǨDf�WEЩ�a��͑;2}�)��������N�v��1X���`���w��O�!Q���>+j �D�E�1��x^�*	��^����/�.n��ۼ�^_H�1�;mx���G�(��'g֍�6��^�ʧ�&�f�g�b�|>ϻؓ��ze�Q�QG�N���M�\�g;��I}&:�i�^?�,k.������τ�|[��4�R��� .�d�jwڶT�ZW�>�٫�ݺ�Ⱥ�*Ml�'���l��+�ށ{��[2��UH��D+��bV�{Q޼�����`�W�t@��\ +<fm�?ev��"�
��[|��A�`Αo~,�Ew���M������t�p�Yp�j��Q��t��3��;���l�nZ<)�ͼ�}p�����"Rؐj��<��s�P��;���'�^-h���u���S�e(�2cK �r1��;܃�ld���P�(�+y��*���eE�#��`D���M�Ɲ� ����n�g9��?�\�k�ia1Z���Y�be�V(UR�#�z��֤��! <�'��j���Kp�0�y�|����H��͓dzS���l���d�U��c?���*On�DW������T��ڣf�����%� f�Ң�˷l���ݿ��'O���ռb.Q��Q�Y�D�K"�
#�4���;I������6���ײ��n�2�p]p�#��x�Ml5�V��c1*�.��ke:�km��Z`��w9�
꼿��&G_�e%����:P�Z6݊�ŁMp��$FCo�d="�nl}�������j�l?����;[��(����H��!�N�vm{��g�Fy�υ��aq�:m
�t���5N�9��^D���k^LG�$�?F&�hV���Q���,?�.�����VE	�K/��p����
KVQ��sg��ug�u��E*"y�������2׎*��3Mסw@(�1JN��)�jgtq��#11��A�����ÓбQ</:�57ڞ�(X���K�4��v�_�2��mU?��DfM/�ɦ��3P�褐u �L�VOŬd��r��:��qĚ�]��l�LseM]�|����]i�/80����4�l���o��8n���)%��UE/�yο�}Y'�6�N����D�����G�q�i�˘^X����5����)�M�&)���껦o�ݷ�xl��)�$�L�h\��4��(YR.<�r@��*�=*�(Qr�b�;��_I7i��T�C�Lx�F�g��[��eOr��@��S+ ��8q��Ά�J!y?&�h@��ygcT-+|0��*�6ƻ����5��a��U�p	��%�6<�����v�'Q�h�9Zw��Hb�gj'�&e���U{��+�g�W.����q�%�$�G���,+��K|ޑ�hu�b���ϲ�����?����T��{��q}~�e6zϽ���r�p��B6ܒ�9#ٸ��r����!�o%�H3��6�D\�\X3ūqA��oF2�bR:�ܕB7|�#w�Q�kky�Z����jL���_?��~n�G_ q
��萹N�R���X <+���8p{�x{�&���{���T�S���͈�cL�q��.������>�QdN��Y�R�bA�k'�j�KӅ���z��);�Q��l�V+�{�u������ᰬKa�N71�,�H�SL�� -�vQ5�r_:t�@��.�©�I��|O�FX�Y2/����PZ�+R�+��`N�CF)-��3enu��X��B�督�+ڗ-L�ˢ샇�*�c�36����|��ϏLa��@��#e��7�B���v5j��V��W��;L��	��k_G�����=	$�I����<El��̰���|�'D��ꅣ�Z%!�a�s��x!�d���ҧ�|�/ � |�I�:#_P֞��C.��̩��<��l��mF8�\�0XQ��+|�'��(��s�gx������&��c�EJ ���}��8�ٮ���� ly�f+�(|6lI�¬ڳ�y R�r[*ˡח
rz�q�yh��1�Ϻ+F�w[��C�T���21��������
1%��{���b�5u
Bԇ#|7T�<G�"�!�n� ��������UF������z��M�3�w�xm쌡���+9h#�蝫��d�_�������Z����GT2����ߔ͹D�+V�p�wE��u8���|�Cg��ϭf�F�&g��U�Μ����n3��{��Ǭӳ�@Y�&���r�"���1�~if)
Э{�$�� lXD�V���E�'RA�5l��ܼ{�u��W�����"%~�ݒ�%�y��(�R��ˀ�w�\q�M�q�|E�#2�s����v˘�D�_G�yf4�-]�k�V{Ȳt����q{A䞄���W	�!R�7�l\����Q���u��`Zj4 QV�K4�������y���`L�=�Z���М�O@��QnR�
#ݭԒA�I��� ��cC2ס�J�R�?O��sI���R�Z���M���*s�m�i��±��|��e���w��#p��s<�[����
�C�Q5�6f�4�/����X��|���@\�����,-�]�]�]�V)-�c�}����{p��n�e�6]&ś5�>"L�����5cE�v��n+�;-�]ǈ
����)�1�w�R����T�~���j"��r7Ң1��_���$�"�g�*+�eU7CH�t��E:Y��U��M��R�em�z]�K�R�}J36�����*�N�����g{_���J�:'J�ÊQ5f�k�AU�l9�bCD_�CS�{��bxav����Lڪ���� U2������n��\��q1�5�9���j��R��<B>�x��Ҝm�@\-i�ݜp[˲�]�,�*��%Uk`(�t�!�OUxs���9l��5�&�yҭ�+�GY �?@�oFJ�!7�o�8�*��'{U�Ds�҆WK����]���F���ܜ���"��AѷlC�iiA��oLiԳ��|y�5l�����NJ�=�Z���R����f	/��2uf�_��/�)�'e�����F_�`J��t/6�þ�oy4M���ק�>ݶ�[����Mpc�".��rmλ+��!��R�B7
�m'�U.�g��2��K���e�P�]��J�	'�e�冾���*�rZ�f�5�F����{�y�2P�����F��O�d�aoˏB?�A"�߄��%��sDp���V�u2�,�Q�Q��&%6�:u�r�U1Y���o#c'���)?O]ūѾW4�\ZA;ء��d�Tg<�}�;�?f�ġ���5�t�Q����[a0d��%̽y�͘�լ�r���_�(D39A�wRK���`��: ]�ן�1����^u�
)��tEz�A��K���P9���<H�ϓu`���.�:�����(�(oJ��\�ʄ�N�.2W��O�������՝D8e���e��pz�Jy����\	��:�ʻNm�m;GP�]�f�zB� �-�$k>�L�{�c�@H�P^h;*�8oG�3xw�
�X>������D�c���2�EHs$���7�(�ex��AR%<&Ow���G����=V��3݂�D|��@�l{����$�Y�6�/T޲r��E޺���Qm�,�a�A�u3�p��~����?؞(Н��%UJ8���DH_�K��PS��ie�#�"p͓�F���v�x�\�qA���F7��J�v��hUK��oQ+0�5]�1�ܼP��1�,
���p�NL�شsd
��J/TeWxtx��ˮE�8�w�2=��c6��� Pny�v*����#1�b]?f!�������	�7KP5A������P|�^@Tc��Q>W�������ȎzG\�e�=ATu�-|��xެ��F�*�	��+tYZ񺪒Go�����9�Q����x�� 26�j{��;�����eƎ��%�Қ����c�Z@��lIj	�y��g��kQ6�-�N\�1_
C	%�M4%�q�K(�L�i<Kj�g)�a��m(�`JU�?<�h�ߒ�N�{�[�G\w��a]2��V�I�����Q��^���]
� *TR&��#Y&#���bD;� sQ̑y����݆;��E(�1 ezO��ObYa�� ��i���O�1
���'x[N��Оܛ��<����ߋ�#��;5���q�g5
�dg`O�p��q��G����+���3�t�]9��_Xb�w�wn�D�1z�Yw�q;��\�ٰ�F���� �� D��{�r��z�q�Hl�E�{/l�:�/IY�ؗ*�@�$�}3(a,5�����X�2&4�¥�@A�2�ψ��^u��0|V<9����.T���	�����~`(&�a!��O�j}���T9�j-wnR����S�ϖ�ˬT���~&o�Eb
6���j4g\��T�`&����K�(���	���+�3��`G���Pj���OBG�%��5��Ek{�����+UVE��Y	۩5��)`���F�i�y����B�q�<�ZR`W劋k��@e�:lltl�2����FO�X%we;�;e�͛�{��Tcu��Ta澌�$ 1��W�c�! F���2@ԧ"cFxj�/����[�a��Q0q3��Ya)�-Ͻ��3�d�>##�lb���/=:*e���gP��)��h	8�h"��^P�͢����|3yj:�o���ܦ���S����אH
�me��Ő�M���i�Iӎ���/xz�Rj\�&�Mi��[�>�6�%�\@�lKl,p�{=�hβQ��"�� �&sTN�^�V�P~���P�`�8�������YV�o�����0|z�-�<��0��l=V) �>O�7C%h>�4@�k�X�BgQ�����Ю)�[/ũhV0��Z� +�(��3>s��]KB7%�u�6�(������nL"������C��GK��sz��t�T��[)����\��g�rtR���\��vwGa5eF:%Q���w]Ơ��4��I��Lµ�U2�c{"g����*���W���$K��ǌ��O��Z&R�3)>�C�x��r����~�'-u�:U�5r����\e�vV $���9�H�L�&�p@����_"��~����_"� �?^�W�Y����D�R��$�Gٲ�%/��Zn�B�}]�Ks�s00�]`|-*�f4S^s��#����d�̈ s�&?N�	�v���"���_��v��h:WA��z����]�iy=�e#���E���	?�eә��+t��}G�Q8J]N��ݘ���Ђ�&�Oc���W�!
�.g�+>�w�#74ɑpR{[�
��:�Kfcg��a!	ɘ\��XWv0����w���"�7_���u��⻫_��>	��{oJ~/��)N&��%����V��������_�o���|lũ�:��%��>�KZn�7=,f[d-2�`�����"�����C��c|3���i�����n�Y"U�����pY)��piz�/�{�k���(�S� ����NL6���q8YX�_�ƒF�<z5E�us}r����A��
C뤁b	 �k���I����5׽��Z �~r{pvxdT�p��H�wb5���o(�Í�49�+L�E���g��E�:G�F���C/hx֖z��/�F'�в�]��G`bBj��L[���..`����rk�����	"�ޖ������	��`�x\
���Γ�g0��L�;�z ��\]�.��@4T&?�@nQ�c#;����c{J�+�+n��0�-ŋ��`udK|��;8C~ƣL���)Eꡟ���|/�A����؟�Z����&�׫F��V�D�L���6/B��4u����� �F���:@�ရ�.��jM`���"��E�o�*R�^<X2j�9c�3X���}-`
6;T�9o��v��[�B�-�p������!��0-�1���e$���囗��;D��(�~�҅rC.�צ?<�(���o��1S6�3v� Ln�D��֏�=.�a]E�`�
��g+{\�q�N��_��a�	�Θ=�UW�����}�h���"��p%�ΈO��@���Y�]~A�Nw^IZk�>�ޓ6\Rei�]2�`�.��!KY�#��L����䯄6����h����y����Kbq�E�m��
CDI�V�J�	*��*��"v�	ئ7a�%'�l)��y<�6@AX��a��2΄�!s�(F`!i%���շ`47i��Q�d^-�Ͼ
曘�V�ً^��o{t�Х�	�^�>.6࿨8ߧ����=��=��X���8�Vx_����@�8��H�������+v
�=ʅک���'��xsW^\�{�:��im� �ԅg��-��-�
���]�?��I=l������N����]�\�����"Ox�Τ�"����*׊��� ��C	+�!��F�
�Z�P�g�������ԕ�(�����~��3U�DREn5���7��ϱp��h;��l���Ko�'�&�?b�[�8{��-/���ɈΏ�J�0C�ؕc�--\0�j2޽Ï'������%�ږ��[ k��n懥��]l�P3�v�ng�Щk�N� �"���"�*�;"��xk<��<K�fñV�l����U)p��d>�tTN��2����v-]b��>�?��G~���)�!�x�hsa3�5��s�[n��0�A2*[�!$*��:� ��,�qI���TC��f���M��w�=-|�Ͻ.X�7�d��W�ī��.ÊC�=�HW�|4zY4����(�󸫛�cb����/��9�gͧ�XU��9j�u�[˚=�QY��&���&v<�{GT���9Uۊ02oPn�[�Uxq�M �D�T��˶�������i<O�y�'�$2���U�/�h˥/$��J�BFζF��;n�yr���eoN�^�F��Е�1!1e��?�]f��>��<<��1]B�k�
�͡�1�ߚ�&�t�X�Ee��/���$+��!ϡ��ݓ
�㘽c��p6��`�YU�� ����S�5��Uz(�G+V��ro������x�2�:~K8��<dR��PҮ��n7d�N�z� ��nSV����`�5���t�2v��{�ؐf�&���'m(b쥝M���TO�<��'�,	Lz�m.��B��� h��[�JE��5׹����C�zҩr��s횢c���) F;1=����ֵ��
[���(F�oGYZ<��|�^�^�jD��X:uZ 铫V�tv&س�~���[J�	�"��4V`���y�o����J�l��q��|�OM-�7ȡVf�:���D#�Q�ĉ^_�Y�r�a���^χ���SR1�)$R=��)�ve<��������M�U��CCV�(o>�V�Sc}�O�}�_9Q*�c��!��_��+oRm�����W�x+v8#J�iJ�T샏�I�{��Ō�=f���S��+*q�cU���m�!�O���˛"�  ppg\#O=�m5z���rh�*Eec�&I�}f��J��pL8����k�-&l+=� .���+$(�D�uM���jD4�"��w�M&	�vw�.~'mM��_s��˫��4`W���
|�4[�Hn��Pa�M0��V����(�9��,�0����4��Jz��Cs6d�Y��iR��H����]q�/AqG������1����&1�0�F0����Li�� ���f�v/���λ�l���8s�ճ%9���%N2-U�}��ubw-?^|s����ts0�=��=�K�<�E[̾����M%�`�d�I�Y�VNC},��\3�oq�0���~���#��J��������*�K��"m'a�-�$����mBt«pۯ�J�Y�NE�; ���_��-� Dn�1�hb�4^��A-�a}���ɥ��ݡ���1�$d�j��_�\�n���Q�U��	����9XIcKy�|���%s(0)aM��#��;��в�G�"J4�r}E��n�*����q-���r~
�PEC�0s�c�{8���7a@�2;�JbI3���o��g��g�{�xsE~���v�q?�`�R��JzZ��&���"a�,Qz�K��y�rL�˸�;�L���4�ق�i��F#o��k KV�[�~*\�A�E��2�B=��I��������*�8_0�e.ߢ��^]bEnfWK�����R�zN� �>��y�0��܂�}����`dƣ��W�/I�ʇn�6�\�=O���7�X�KB��-_L M�_�*�Gۦ(3�,����D�'~��#���G|Օ@�
[����~�i¶N��p�a�;�b�[2�o����1ɏ!����_��>d������|?�'���{{�''Hi&9� �_�TZp�C��;V�O�]��/��Q�Ͻ�muV�l�%�m&S��X3|!q)��C9�l=�=)8NB�-0��I �����M�:8����$��`h�7�֓�u+���{$u>�+������m��� ��G���r������G_�-4��q���^*UkV0��|oD%���)#�pF"�N�)8�E  ���Cɯ̧�v��T�"��n#?֐�$F�԰�������ګ�@��6�4I幡Gq:���M2�6~#��q�R�NW� hr���7z^���/���(���?Up]�=�j�� l�n�1!��E;��6�.�%��2cUl|�'|ܐ������㽁�H��'��Xq���������,�B��ϨK�b而$A�פ�G%���P�3�����|�	�L��@a��[u[���U�XI\к��¹s:�ru���k�8�~����^ϗ�VY4T~��*�(�+�w��reH E�y�ӆ��*�������,�Զh�FYjR9�Zҥ1�r��M6�El�/@5�q��
Z\W�yM�`��p!(���{BM�F��|��} �޽�qW��ĥ6N�i;���Ս
��EX�6���1��7�v`�#>����1F�ɦEJ�](0N����:f�G�X�@���t+D ��������@��C�i�r!�I!`0\��S�1>"M�`ߡ���T6P�]!էh4��&�p�Z���%Id��*޸��3&դP�q�7�Y� ���%��,�|Jz��y�4_��nH���[�lW�>��<��C�`�p"�c�
���1&�pq�q��f��BJ��c����C��E��9|N4�05o��y+@R!��Z:P�'8qlyV����M{M ��n�+x�V՞� �����R�O+�7EO���s}/�P�H@Cł��yc3�&{���xC���'D�/YQ��P�|�����5�H�NR"���ND �$���,���뵋�fbT+��X�$�2t]5����Sw�x�Bu�p�c^�%֣���͏ȷ(�'r�rр�Gn�a�<j@J��!l����<�}�~Ku&O�������`�jM�`��V���+���:Q�qR_P����'�������I��Y�1�(Q�rfy�q�����y�ej|F��5�]�~��PQ;C�������YK	$�Y�q�����@�Q2��H��$Qet�{i:�ص����/H��Ec�*�l�Sz�
�Ņ�)�<w���s�������j�&�Ɉ�4��m���
��m�Zyr��`ekk�(����J5m|�:��0�K��-�Q�����O�1�$��ꨀ�H2�\����r�����GɎ��d�0���=��fj��-D�f\�Z��Jd� �Bғl<
���]�i �Ը�P�[s��*E���<VĘ��-'u���q2�W��Q�$�%�٨�����JnW>u��|�Ԛ!�̉]N
���fJ�E�<�f]�fM�!��vO2����0�@��w�����c�����ZQ  ~������d����3��Lp�տ��*��_;[i���S���^��*�/������껛GD	��2`-�w�2��G��J��v��'s��[	Ł5�f�MU�p=�/�-XY��7� #Ԝ��oBO����~�=ٟ�- U4�i�l��!�yE�G�cW��g�D�xQh������~�h��S?���X2e������t5�Aĳ�������Z�����rSyw`��ѧV<9'6&���8����22|��p�~�]ʥ��X�7a|��8��<{O�����U0&,����/���ً	�,��|���}������g���k{�2q���N(Ϗ���{�X��h�c+���^i��RH"�c;�������NA�[�:(�C,��hB2�`B%�jn�{_H"t,�l��a%8&���Ť�`��~B�MBiR��}*>� ^er��J\6���ꓺ�z����L�e�:��6�6��4�"2#˹U4��Q�;춟��)�Q���~/3�ɍU,�n%�F��I�<��2`���?N;���Z���fz��u�:�]����e�+姕�w����jz*���>>h�a�������Ɋ�
�	�s���o���
h&�x.����m2���Wb%.�fS��n�$��5�h)Ƿ@ � Y.���Y�L��-[��g�+>��i��;�^#�9B�fp�p>I}@��1n ���5T\ӴF���WYИ^#W�`�@}�iw�:��u��[PX�EJ��y��o�\Yy}?y' Ҵ���6M�U���}a~F8�ɤ�Z�S'+O�U�oKK[oj�y��@��ڎɹ�)��ܥƍ����e��d^�rĚ�)v��C�B=�i�7`�@��@I�(�z���K#Wp�y�{{Qd8(�_�����Sp�7�F���Q�5璒�L��*���	�H>��������9��Elqς���^��He���0��Ha�c�!�	:�E�����Py�s�pA��n�dez�[ܼq����!��0j�m� �V}\�@]Û<�i��'�s�'%�`�9���_��l\�S�Wp��e�ϥY����O&
s�f(�$����k���]����.b�m��.B�=�����b�R�8n���ʹ����k�y0��)b5t{1'�N���[�؂�=S�⦂�^��i]̹�:�wt�Q�n1��s_�׸
��\T�����=�'YT�v�`q���m�RF�% �H��3�x��	��o�SN549��n%����@8�lK5�EmU�v_�/�`���<]����!$G��ُZ��S�u�᫿	h-�<���JHF����]Y'F�~�
�K!���'��0��o���p)��~eܷ���غ��nc�<},�N���V�XOiſaWX�^���6�u��kB*#��(�wП��	�?�7���>�F�6�����^Bb��6L��d��|��Δ-|�fә�v�Xw���.��ߔ��?�I=v�ܡ@�s�Op��O#�q�Jx���_���O�����L��&�Ԕ�>s���r�}w%,��+[�S�L�GAM��+�7mʅ���P� �rjU� p��{���bw�`2�+	"
p����-Aq���b2<�ʝ%��Z��$=7�����/B�oy�;d�%N����"5���f���V�.���
?-�V��=7^6���JTCI0Wٰ��/k�r�h�<�}��~�:V{�c�Jl_2L]m��;|OH+�����&2��&|8�s8{�g	q�����<��������T.btl�hߔmt>}Vٸ��R}�޻.�{^5�:���O<i aU�l�"��u���0.����)�	��V�^c�A���{Mk��J�˲��f��âtz0{)_���/���mׂƿ���MT� �Xy$�8qZV��NE�������CY\PXY�kǢf�f���l}�f͠o�1�L�tu〲,��eR�9����'r���DTwy�/�㔘���ƾ��8�ʁ��ǣ��*x�(�*�������.-N!i�K��� �@���D�l��p�����!g�=����.�I�?�+��^و8�E���s#�T6�=>�����i� �(�m���⹉��NN�ON�2%8��`������@D�O��+��"�&��!fZl�U�9�N�^]$v y	���ߒ��n��@/JCI�7����܈R���Z��Ƞ��� ש�W����*�	#���'���˯�W���a��UG�q��+����i�_Ɂ�%
��PB�Unl04�C&)�EȠ���3�w �ʂPM!U�f*'F�Z�G�4���R�"��܉�Kӑ5�RV�ތ{�h���f�$�F��^�K]������)��rr=.l���z��k��S��3}�m�ш5ܙ��s�Ob�r#��&�P	�iZZ`5���7Q�)�Sٝ�����;���D�a:�f.��h�t�c\с�������Ym�X�b�3�'3c�%��R�'�����CA�S[�>^��*q�&jf��XFｌ��u-�t�� �N��k�G&�6P�m駣�O��;�P	�
(&~�Q���:��Aq�E��g��^���o���eT��YD�x%�wۻ f���4|�F�|A1"G������:��Y�T��1ln����:|K2x�:�ׂy�@.��k��A$$���Cl؉|^�/��w	��rk�t�9p���R�GK7Gx��a��:��Yv�v)�_�ۤ�����y�ˀ�8BO�j�zeU�l����>Y��CJ�?���̼h�n�_D�Y��C��4��������=�لaپ9jU��`��N�(�	&g�9����*�4�7���|�N�Mk�~9g����H�8���1*�y��P�� M_�%&�0:H��P�<��K��3� ͸P6�E�������I��uzA��˄L�iZt�z��{�2m��3z�԰~�j���a���ǜ�"�At �>f�n����.��@���(;�����QP�o�1��ol��3:��%FY���=1�1���L��bԀP�2t�e'�J�b��pdI��N#���� ����!Y�f_�g�?{�O��3�J�yE�n�� Ά�s��koħF"�۠��_���c���I@���~�Fy
-�ɾ�J�o�����W��O\b�Sv�`(LC`�$߯�7C2�<kߒ��͒�ќ�!!ƴ�>��
˭��Q�F��y��������*6�늂�>�R�`�)k2�.�ۇ�i�7>��j7*��<�B���Q#�䛆)ϣ(x ����9UBAZ����]��+6{�����W�{WR���Pۨ�d�2I��0;��K��Y�L�5KB�|�������L"�;���&���,vQ'�%�l�L���S-zkQ�F����[��o���E�0�0�(M��<��_Օ�faih�S����r�ĉt�o�}^��h��32��"�2[T����.m^#2�"<U2�h=����34.?�9Ct��]��'zs3͉W?�vോ�I�u���E��e�=�VS��W�M�P�Z^��~�/����^k'a��@�ym^ϚG�|���y�0_�}3��Чqݾ@������P�Ji���纔�,�f� �g6^/��?��t�%%s*F��=��ξV#e�k��Nx�<�1n���E��C�)�P���j%|f:��7���5� }������J��tl�C����m5���<��W��oC&*��b�u�K���Yц�IT�6�1������̝�`dW]�xsM��SPqjf6��<CG�]AfS�@���۔�1����.ఝ ��M{��|��*����z��@c�GJ�㌗3���\�z,Z�[�R[����"d#?�r���§��&i�'�����G��ic�����x�TzL��iI���«[8"�Hm��J�L$�ʉ��H>�e"��ߐZ{\R���h�?�ʩ�{mE5���P��!��43�u*Y���F�%P��8�������'��p����H>1Z% � �R\|g#�������|���h�Ϸ7���qR�,ԡ�k��Ϧ7�=���w���XcI��1�]��u�dǛ�ykZ��;�j��EEY_Y���5ft�p�����U�x��mD����>V�9�Y�S�Vܐ��JȋJ�:ϾCZ�?M�A��-�=�T�|�6Q����[�M)jeC5��ˏv[��!�D9jk�Y�~��ެ�,4�`
cҎt�.�� �f��]��.4p�)V���tO{��A0���_@Y亷oKg�mW�p�5�*�ʄ�jM�sv�V�F]{fR#;�,!yᇾ[�$9��S���s��\���QiYc�8tY�*�M-��-)�O���#.�+4?���)������I���ǻ��6�AD�R~/!ᖊ��Z2�PK�ԫ��K�0?�,c��k�EvUʰԏ�4ѽC��e������d��$B��7"�U`�Ǜ�j�����Hf��G���dx��r��߰�H^��Z�1���)�����:������M�s�]�C;L�\ܜ;4b�������%�V�e+��|S6��f!W��_o
AݠKcd���#��\(��2�@���������h���Iq85{AJ��Msۇ�6@�O��^x�O$B���f�MIe�7}�{~	�%����}
T�$��7�Ph���q�gf����>��8';��) H\ʆ�����o�Ě28�t��V��B&��*���%y���)�<8���|�->�}�#��|o��4���!�ˎ�8�p.��l^%.��_Y�V^����%�J�#�!��ҹ��x1���Jnu�!�a(2p���~�uz�{g���mp�j���)�4�̩"#K�A�T9��c&�u@�N��
��ƓU���9̏?��po���>㋋��J����"9s=_9��KŬ\�R׹9�X�Ս���u ��?>鬁߉{�U�`�s��&z>e�1� �������E�_���j8I�pj8Q���� �P���!ׯ\�՝&؜m~��s�e��h��%Ir�ޱ���4"E��dT4���:�$G�J�3��~Q�r*���?'��ղ���걃�퀜��N��7�҃U¸>�ZH�a��@*ק��둣0��䷝?��)�P_��k*��;+1�{�)`-V^2bFU���*e�F��q:��J��9�K�3(y �_�h��8�!Y}���������6-rO�q*�D��;
q�^��PϟJٿ��7�V*#�q6��g,R�������r��yϫn�3�vkD�`Z:��;��� wGT�#���_q�i���y`���d�Rw��cl7��=2�F��4n?J�.��L�om�?D�o��>�|�<���jE�Ŵ��q�Gh�k�z����:;ACm랣��5?�r��x��5�qT�d��F�ŭ�N흈O�~P%k���W�T�)�f�st>�sA�����B��y}��LUl��!օI�%���w`�#��~)$��K��5ߵu�8����'ϟ���Mi�����w����OM�֊:I����w|�ҋ������<S¥6����1�����YA!7��D��T�(��h�)�V|Ђni3}��S�i�������]nIA�C6wf�>����
�q�d���6���8���]�p�����=�o�ƋQ F�Iؘ�*�}�@>��:����E�]�V��'$��L6��K�}!9���"�ڦ֋���$i�G ��N#��Dn'K{륾����`�NQ�
��-��-�}��$Ti�dҐnȔ.�bz~�����z��C�P�`m+�y¦I��&g��(w��!� �&~�#3.ښR�d��=�����+gY�-)}%��{)��sa6���WU
,U�.]Z-�7^-��r���/��Rf Պ_5%P��:h��e�>#PA�}t
�.n�s9�[�E�^#��li�T���`1�G*B� 1^���r�U�Kj;�H&�>�� Bb�����>��e��CIC2��x�(�������B�<��VI"d��<P�V᪵�$��"���â�׬�S��mb�`w�K�N ��D5Ng龉 �oT�gJ>u;���8���/�ݰ˛M�]���OJU��օ�'�<�V��n���Y]��H�M�G�-�~}J����U
ǍԐQh
���4Z���7����5���Vb�m�%�fb�����ʣF��% �=�e� 
��"e�JD�w�!�h/aCP�!�ӑ�T"�GW�կn^�S��4�N�;vd����sR�����=�_>�K~I����L�'sM6N�|(�I	q0�|�iY�����tBF_�7sV=Β���|���62��⚚a�G�̴~O�҃��h=�6��.�RI(�lD�%���`��.�>�w�3�1χ�e;Á�R�r�QčhA�/��w�8��l&ib���8�9�AB�4ȟ7sEӊ��m1���`�z�u�����~�`+�ۨ�{0�F�P��91х] z]��ro��d���3�;���u����x��.���p���'V�s&�0D������=����(l�t�/R��97�Z��΀���u�^�Nu}�x�.X�^�z��ɸ�u� �XV���ށ�}�qɏ���ӿ�LO��ڌ"�w���Jb$~���H7l�b�)�*����|e���;$ӂ�X���\�e��!0��&ye3�;@0G����=]��^��y�}��T�b�OHv��n�j�!#|ߌ=�ۆr�V�U C�5t�� �OA�eix �3�v_U��#%V�����(�q��rO��W���}�u�@�tJ������euL�mQ���9��O�E�z5wiWzp�/�Wg���%�Ӯ��o���}����[}��(���W��Vej�����sKq�,\��0��n�VZ�}^�ޑWJ�m��@�J\�T@,���u|���B�Mל�7~|�6�F����O�X�ȟ��VT(qkN
Z���''�!`=��3��ɡ�~��1�Hg�c��j�0G'���|&
�nAw;�-��#"2OU�O{~���yN�=Wt�"�lp��C���0�Q}�����(9\C�� Y���J ���l6љۮ�����9O*g�M�4w	]��'���/[v6+n����T ����ݷ��EfϜ��*=ǁ ������R���'ɐ�,2�p=YTN\���5�X�w���+���r��x��zk�^E��J"�q���� �#����=�E �h2�ˉ*
�6���� ?�}����O�#UC���זؙ
��X�Վ����X<�$1W�Q�?g4������L�)���o��Azq�S ҋJy��2O\�uXYӾ�qi��apa�3@ՋD��N��(8:��'N�O�MA$�XP��5ߓF�X����I!��C��Q�D����'˶Eܙ �ϯ�I��by]A����O���ΧnG&�^qw�D�25�ю�q^���M�4�k�շFTF�a�]�[O9\*���
�?%Ȍ�'�
�^h	_�ژ0�B�:L� :e�X��F�[ݭ�ق1̈́6��U�S�Ӿ��+U�a�>��v��n+`g�ԉjvBتJ�P 琷��%eh���>��^#*P�Yg54��X�I�/D��+�@ ��Y�gld��!�X�S:&H���6XN�3U{�����2C`h��9�B�����/-r��W>>��H�o��WP��I���� (��m~�'j,���&T�3D�eJ�U{Y�|�iS�����w�V?�7������4�Ѻ�����wH|�b�Q��@�C������T��,�6o�K��Fhw���5;��!^�v4����U=%A�}��\�gx��W]$ �h�E��=`w�n�'�B�]�z(ޑ
Z߰��� �`Afj,�m^UA��'��-P	y}p��4�����J�:#3�{�
�Z֫KV ҄?�K�rt��o���Z�hF�Is����I೶!:E-:� ?�����E�����,�b̥��-�:q� ��mE
	O"\��JR?'vt߈��:2-L�3a�xi��9~Z>ʏ��AKb*n���Q�a��nħ�O���Њ��P���=��1yhVh������8�)�<B4�6���ΤV<�Z�����cݲ��B�np���֔��Z�MJ�a }���%$�������'�/��&�>���0_�W�ƱE�������Xjt�\Ӊu�@�2)i�뉓�d�ë�N
�Y�q�3Ym|_\tÁ��,{	^姯�E�����L��|��h�Yr�%f��9�gf): ^���d�y/0���u�^��,����s�@N��dD�%΅�����I����̌~.h	U��"���������'[�c�/]�>��Gt��F�D��1ӗ
�$�b�a��gE/I��E-�
5mtN@f}����9�t� �ߓ5s1�<�rCI���o�z����`��o$����=�39�7���ح0��Fs-�ۑ��3ӽ�fMj���#���B �hD�EP �|^�/il���mqE����#Z��z��a��#��8��ݢ:\�=S�n�-�.�ыBn[v��VRDCׁxV)Ju��ؚ��ؙbnEK)5������+��yH�7���?u�[�ɳqt	'ߴaC뚘��T�<�'��JЃ��`�4S�A�D�G��>p�PF��@�о�� ����/d���]7��zt�y�׼�Z�s�`����V�<mgO� V���h_v��,�#���r�0q IG��vj��e�V��@v3���N��!m����l�_Ϙ���_?�l;����V�ѦA}�,}���Eky��#�o���.�m��V/��R+��/^�0ɹ'��f�#c����T{z��WZ͐�F�hY�xkQOA��$�Y��'e�dF���Z:9ĹY���[~IN�@k,z��5�j��C��r�<�5�{� �
�86H�5qX�TMƉa���q���0�1�iYw�O�u����ךہ�������s;|�;���;��;=,Jb�lvt���IiR ���ik��<yiZ�#��X�F�)���2'w�Ti~���1*��w��r)��T�7VpF��r;X��YR3��;L�R]ڧ��m��Z�>\׷�&���i��J�<��\�^s!�Q�L}��6�n5m��)7�$-�Pi6L1R��-��t�F��h	%3��.��`�������j;_��c'�-��$�(_�2=�}�U�l�q͌�IaI�o����d2 ���I�Л
�)��-���V��	ė�z�Bu��ED2� �]�A�=b�N�I ��?�׽��R�PT���Op�9�e��^�&�8���<�an'+�dI�u��J̚H�qO���>�-2��DvT+��t�����kھ_�a�`�T��g�|~�@��w�At���������u�~������pǉ�Z׏/����H��Y�֛)��U��W��Ͱ����V���I�mYJ--N�м��v-d���4}�;�n��yk��;t�$:ǳɯ����68t_	�z*e:=�˫���4��.�M�ծ���ug��}�i<�o7(��;��!��f�h�*T���0�o��L-H9H�����<�B���~�h�L��o����(W]5��� !�҈)�R�3f|l͵[Z~3>�P�iD٢T��I��Z_��) ~�=�����Y�tHg[h(������0���
��T�w���=!{�y��t�߃�1&bR)t!�U���`l��2�ubP�YSڻQ^b�7#���as��8����5E�}1FLC��ᑴAX�//��P\3$�Ш�D��z!�m�?a:h�o�p�k�"ll�j5xzƨ� bR>��W��ߢ ��x����5rB� ��Qp�L���\���x,�D&�m$��[�SmR����"�w[q]C��QM�D2��xϪ�19rB�g�A3�/LM�x�Y��߳32��i隙��ÏS�� ���ӧ%�I�'�H2{�Ի�R��[�,A��KԼ�{���n� ���C���l<����xڄ�&)o�U䠷.	�G���ɳ ��s��MC�`V%�w�e\��q��ċ��[�:K��R��[0nH���_�+�m\����P���'��� :h��9c��J�LZ��p��h=�x�X]�ʵR�L�{d�	��l���xb�uC��u��i#2������/����e�r����p����t�F}�� �W&��V?�`�@2�$Z�Z3��dْ��I�cy^�������f@�ɬ��ȩ"�ADb��hQo?<�f�w��<�0(�ϸq�B4#b�H%r�՚��L�5�G�`f&��t�Z;���p��xQ���Π��.���hz��2{Ft�HlTYWd�&V��L�r�;U��.k�j���\!�0q*n��;�K���� �^ V��B�{=���p�M l�Q�2IY�Sh4� �֬c��3yoс�(:����4q�s�g���	6�(~����a!�*�>�6�qQ�ܶ�
���I���}v�A"Bv ���T�ail?	;G�����Q�$Mi~T�6f���8��w��[�)����zD��sN�郹�;D�a����P�~t$�+.����P:OAX�,	Sp�"�;�E�j�<Z�<����> =E��E�~
�Cƀ֗��S�"��DN��긳졕c�&�
�W����C�5�����
'$�aw��ɺ����È��/���c_O��n�������Sٖ�p���e4���c%w�=�;j�} ڷn�e�|�]�����g{��H�T/?=�$��y z����Ś��}0��%��uz��G��塸���
����,aQ��ݞΡ��H�!UR)��)����ɜ��z�Ƿ��J�8�{��_��b}�&���O����@@�¤����ty�Kc�R����߸ �/]��D��9�n��l|N�O��_H݃�۟[Ts�H���_�0�	���������G���J#���y&O�����g�s��ArS�ke��Z-h!��&����|W��i��\^w�&GNmՄ�Ԝ����$5�(�4 T����7�c���C����?7���
��f��*�C �pf>*;4lT\Ʃ�a�YL���i<�QM5Y� �tzouJW�.�K��,����^&��[�2���I�)���y��5����?��H�R}w�J��;$��)YeL��s�y�I۠�'�D*f<���=7[�G%�dð�0�+Zio�����"t�����w������JV��:�aR��?�nU���l�S]��K���oa&.��gF���d:5�p[{#���a��9�N�*����l7̧C���X�� �K9FxV��`k���p��m�[���4�8�̭�URذ$DU�02יD��o�P�����u��K��Slۆ�`Ct\AD~���%̒R>���5�6hc���ؖ+�Rt�g[FI�dJc�j�1�/��	����MYz�]���| du�f`�����yG?e[��p��Ej}U�D)�:����A�6sg)a�I��� �r<��m2^���}�-�����8wlmj��z�,+a<]u/)n�
xߠ7�22q�A�u'���˖�HE5�-�f(�1��)�x�xל��c�>n4�����y�9��	�,a�}
�rrS�q�;���r!� ���͕>�����}��l2ϭ�&�0��Sk�|���7���
^w=����Wq��4�jm�z`�fH������pG�?iY����l+���.V��"�hi{���s�ܕ�~�:Y����;��F�VDC[���A�=�K��_��mӡ�հ>
��>H�ƺ*�Gg�U��j7)5��"��3M����S���,*}&);����Bw\��
	�4��dt�X��k@����p�6��`_�OLĸ�/�Ĵ�<��ˑ��!� �/|��˅�O؏���*��a����*�(�ܗ\�r���_ U	��ǲ�D��8b�vnLBfeH�Vx��8�굻�Ѧ���/n7�j���^�~a #�h@�DO�,U^aV)�EY�e�y��Q�n1�4�2u(�f;J	NӰ��#��8��b�Hv��E;�xqA�C��d/S��^ˬќ���|?���م�D2���R,�)$��p�����Қ+"]#��>4[L�䀖f/��g
>�3�KJb$d��k9��R|%!6y�+�g�o�5�֘d[�]�\M#�c�?��`��.�+`#�u�xՖ(X?��hnWZ�u�!j���V�����Ԇ
���T�O��Wv��+U�:0�w���5�-J5�}"��O��;;]�e�}	�y���'���%m[�4�7�"��}@��:�.��X� *�sjh����]�n���6C�]��X��:>?����^����aV���KX�:xU���s	�vE�ӧAk��Ri�ͺ@�Y�h @���L�n�jn=2kJ��L��E���@.U�}�M��B[�I�ꍷ���
�g(�w�7� 0�e�j򐅻�m�^����!(�댏�w��f��(�D�_7�7N��Q�I1Q��$&�5���I}l���D9�o㣺yY%w���?���K[�g�9��=�H�}�鬅E0,`S�� �̘-?]Q��H��v�8��p,J��S�(���5�k����ƞD�a��E�~�j��}F�6�🎶L���ꁽ��͍��\=x�&�	e;PJ��F���`����w�%]�A���b&p3v%Ƥ�).b�kE2�^48���A��2Zvd�ڻ����χ�"�<W\ɜ"ϝ�{�w�,�bBk��i��b�����6i	f���w5���!ɬ����3��ˉ�`������6 �sO��t���U�W��FP"G2Q��TZ���}%�e>��5���=�r��~Eu��p���8���\�<�.��C+I��~ot_ȺP���,g�Lg��02hީ�s��z/H�L<J�xOidۭ����xd�N�T���K���;����T��'��T.*�\���?!�0�}�粴�=C%����mM�����^ib'
Jq��o5�xg/_��L/J���N���9�J��lA�5K ��(��{b�61�[@��ؔ�Xv^�uޞ�� ���o�=u2�Vŭ%D�Kk㓦����*���l������m�,\�c׋9� [��$)e֚,�5m�� )n>q�*G`���}�"h�?<l����_�����7�i�p��
���J�8]��^�~c�4��O^	)l.R���f�OƘ�@�-��~*�c8��_��N��� ������@�z���m4�mYd�J��e\�2요�n��͸F۴�������9x@��e
ԫ"�Ǿ12��!����N?�����<�k����l�wJ�M�P"�W20�:�#�
��} �=n=d$b�;t��Rf@!9���"�:ˀ�[r`N?��/\��D��󬧉qȺ�E���S� �F�-��S
P�Ġt��Ӌ<��\����qN����5mRq_7��?���s=��P�U�2��vPƗ\�'����5<0a�X�4�T`;\�j�9'��l���jҵ%���G_͂���0E$ј��jӫ����$�)�x�����#l�������14y{��R�1-ii���u���a=j����x�kCN֠7|�7��yl�5t}�I��Y�h^1)�1��)_,�Vrd�D@YY��ܦ�A�0�>+&�����_2�����ͭ:s���[�ɵp��NeX���A/_�o��W�i�d�2zt)��!ɑ<�{�G� mB��mV��\ƹ�`!���h�`���5�-�YK�2�M�=l�:�:�Z7j[�j_�p(��;��1���R8*��.r]���^al�aEKwl�Uy=]H6,���J��,�Vɐ~�*���{�SUk��y�\!�6�^�C�*�ڍ��i9���0hG��A�[J�ܼ�$�����L�vC��4s;���|C+���Y��'�!�\��)R��<������Frur���mٯ6�>�<��]�xmSˀ��s�ұ:- [E�0�1�V㖽��\T�m�7,v��8��Q���)�#�g�R��-��R�&[[ˣ�W�-��>@���C=��T��u�����1�Qdt/��T&
!M�':N߆�6鬸���4:R��L ��hY��qaKo��Ppjޓ7��@6�|�Qd���[�X=
�7�ǝ�f���Zz|Z�}��+!�����H�P�.;fWG�lM��)fi�W��Ԁ?o�+�����U��2��:A��%�#��ߤn�c�BbX���;��n\oł7�%�آ����z��DV@�)7S�1�'���~�~T���s�1��ܐ������.I�w�W�� ;
۟��m�#S��LIfN�@}'6�5e��sws-ڛ��!�n�$�����/c���	l,$�޹V���*�x Aiݠ��V�E��✭A��ͮ��t~?ZT[9�j�ď��o�m�%ǹK��1+{	qN9�ߘ���3�af~L��fG#�Z�㯕�&���[K�?b�5:�CE�a���$7a�v������dQ| �z�	�ӾN�E �c��g�.T�X��S(��I�̾7�ޮ�z��T�J\��y.l�a���W��Y���Eⰲ�ek��}�x�=�0��(,t�w��-�zGwAB�°�N�Ye�+���-
���E�+��!��̋��$sc�	rB�������g�v��s���b�#��J�������G�
O�w�1�2<xJCRV��-��K�LsGK+�4-M�}�Z��o��Lk6���6������9�Òo���	K��>3������C���Da.0c��b���P���4.���2��95���Q�'�� s:h'���#_%���ᢦ��BI�v;k�������՞�je<�ؓ�v�f¶��f*avZ�x|o�?y��&�9�e���&,�b$��:H�]��t h�ME'��:V�)��u����Ҩ?��+PX�,u��1�)�4�k�)���>ؖT�] �����#��W�������@c��3�F�}�j���n�j�X+��:䒪��)\����ٙ\C�x��{��nfJ��}�Md�b�)r��ܗ��]�A�6m����yO��pv����
��WC��5��B\N��\�r��O�	�qD��,���*5��o��*JkPY���B����Td��Ҷ�;s�󓋆��&�w�O����΢"�l���%��(pxr_�gy�?V����F\4��I��B���x�md�jP3�{y��S}1%p(^�v��P7&U7B�%�-�]�b��b����/����&k��<P欖�H4]�8����NW���7yz�����܈���.з�;2%��NU�L��²�`R���s�w0>���j*m��6�԰pY|�),�ئʰ���!@�h �!�ikW�8����QN�=�;�q�d/�|��S�t������E/���g�{g3!��T�ܶh����������I0 ���&���u��:m���2��ߣ�a���vd+oζ�z�nqn���b����G-*�$��3)@ ��o�;�^9Ҥ&��`��W�lϗ�Y����e��>��o�
%�������\jI��<.���3G���p��!08p/c�R��;��V1>Hɠ
�[r��;z�UFf#`��QՁHV��s��u��B��rV%���J�C�J�P&0��Im�|�ڃ�y��,�I�����A0xq+�px�@*�Z�!͗��_o	�	k'|�����Km=���;��ف�凞��4j��q��@b���?u�ݯ7z<Ɵd�z�.p���b�Ot�ͺ��N��b7�ށ� �Y��J�wpQ�R6S�����1I1�}�� *-����#h�5���Y��ו��c�����$�dAY��X����=���V�Л�D��j;ِ�>ޗ�8�.i�z�{���A�U�k�=B�n5�y�Ns���@-�L�Z�+n�64�1H�ʃ)��%c��rVkH𱸓s��c����h0���)���6w��d�]�����:�:�arW�����:��6�H�����_��(ƙ�ĳ��$�k�Bi�Ĝ$_�O.V9�	f�}E�Ki���x��!ל�Q �������qi
���wc�UU��*n!� 1(ZZ��K{���W��;԰)5֗n��q{G��V��;(��i1k�v��!%��.���h2�Xmȕ�ɏA^��vb��kG܌���l�	e9=�Zk'�8�=Ɖ��%ا��%���y%���������p����d���=�Gfg�p�b0Ė���E�4Hc~RY﵎�xX+d�L�$�$V��P��h�,���+~yDRt��4�,�Af���8�q��<��5#1�s)��r�t��j���i���F�ݢ z�]0��|��g��ge��9��+�:^�s]�϶ն���x�*!?�-��g0P�]s��`�s�o�r�M{t��:��Js��ǜt_��\M�p/��G�sP��50�E㜀n��M�e��t�0M���e��/��ߌ�l���m���U��"��h�6�~jR�vHT�E��~o�Z�~;�&vt|�K���h����e�nY��J��僭��ӡ9�'Q��b,���
��-����g̉苶�e&%�&@����c��%��&�H!�=�p��:7��g�����[�pQ���֪՛c��5p����Ů�6gH���S̑`F��5��/�1'BZ��75+�3GN�������f��K�L!�� ��3]r��s�l�kWA�q'�k�3v���z�9��~�k��Ǥ.�(i���\f�D��?!o~��P'��Z�n�B¼�����R��3bЏ~�r�$AZ���RD�{̼p���l#7��P�
ԥ��i�hO���q�u��FTh;`
���i�p�m�o�g�Z�><�2k-�iU��,����S$Nn��8nU⇌����p(�0��@���uh,*�c���˺�s�}����I.\)�H�^�,ύx�I�S�� =��W�p��1I]o��:��c���;'t�q#�,���i*nAH����wV���C��)� ┊o�c�}�o*�9� ��8����>�����E��L�%��{���}Af�x�V8�q)��	���]���ʙ����..�����2|PvV����^摚���~gs=��o�}&8=4�4�M+\N1��q���G�X�Z�x��@� ;0Mz���#� ���\�T�;�+��L_�y�x����塅�3�8mA�.�w�h忹�]��|ʫ���8�{�qN�K$���d���r�qD��p	���+V�ҝh8�3C����Vv[UwGZ�xU��\�9(�M�vo��������tK��dL��{2���Jǚ�������j����?t���Ъ�mUL�!-�t��s�o)S�4O�H��bҖ}�Nѷ���݊k"��z�(ò4��=�y�������]����O���*|��3��vڇ��X�%AL�V��f>��a���վ��/��(���ZC���d�d�J�u��[A��{�ua�����E��M�����wQ)�;3lZ��u�:�@����'1�e����BE������d��Õ�X4haɗo��4� ��,����������q���)'���p�O��q=DU��ױ�0��i�#�������M��}�K�i���V�I8OP<P���dU*�� d��zeI��@��(_��w��\���r�J5 q'���� 6�óY�fE0 �lw%ԏh~ �Z��j �@�B͐�y.����w��2y�c3�i�KBQ��ֵ���v��m��z��6�=RV��;'��E����'��A��s��բ��@���>��%�����W:���Oi��L1N�F�p0CB�+���9k���G� ������I�-�p�Y�Z����J�V�����;t��s��a �O��lj�����A/����%�M���N���Q�����������9
�5A;�"Z���,�v
;���q/��㖑���G���������e�i�zѸ����a�1J����bn�^�Z&*���AP:54�e�ѯY*�=�́;���S�QfoUPhΛ��C?1:vp������3�.[�P���󅒋rd�#ag��#I}}Fx9_�/������:�ɯ��-�W���)˧f�=�ٗ�$�ڮ�u����P.��Ί�&.�"�g�\Je{`�S��Uz�K:B@�بm�R�Zr��N䯱��c����}t�}�e�s��8���N��S"x0��X�Ɲ<]
t�X��E��j�w����jS���	ڍ_(m<'N�ZpC�p���,N������J��G�o�W{k��X���5ܷ�����a���*��50Q�? A0��r���wV`榮�뮒 �kV���a$�kŞֿ���KU�,�=�����[��a����U��Z���7�Sy������o7��E;�"4WG5���$�;v��Et�P\~?��u*�:?���d"y�!���i�hr����y�����}��b����7��(&�0��4����=�gy�*G�T5��WE�f[��g�n�ߑ����Xt�ò�*�ɯ�y�8=�� jN��g8���!��H
De������|��� ��{��
��0��U�+���Q�^9�~E߸�]��0^DD�����ˢ��,����1�D{������XꓔdDxL�A29&+�QH[�P���Da��hy����z�-�;+��V�� !,xÒ���M�{�S�Պ�S�e��)ƏǇ�<�m�*[m�8�X�B�n����7�B��_�٦2���G�����_�c�*����,W�pTo:��}��h�	1��E;��B�Y��0�p0k]���Z�w���oݾ�:o�9N��@���f�h���ޤ��S�¾�B���M��&�^0W����Dj�en�h5�*1B��"<I ,
p"Q�{p-���h�["�� ��<�q�^�e�g����	[���O=A	�'��? a��&��瓊s��1��|��<F���>ŏ�!vuN�� ŏ�˒����`pē�^�[w�5q�4$uU~.�/C�C�y:�-1-��ż���*��zg���TS�O@�4},7d�	I��(�����"��̷t'K����a��S.��	�ɱ.7ӧb�rl��9k�D4{l���q�����Q���IB4��ef�`A�o��a�V�J��5��?�.�{Mp,~QX���!̵�x/raܝ�t�k�rٮ+���<5^�����1�WD�¿�yQ~�)?���3����<��Zx�:�q�\B}�����A�]��{uqd�=�c������p8������sjל@��"S9��������Q�2��h�Kߋj�98��G\�U��Hr�Ok3$�*�p\��_D (ӹ�[G�V/ݜ��'���N�2U i��To�k��R���W�u�V�(��8�^�P,���=��g�5�Y�>���_K�����ӛ#A�YUXSs��BQ�gnv��5�`^�I��ڧ�/�:����gHJ��̼P�2�6�s�J9�"���sЧQ_f�j��Y���������s�o�>�j�4�]k��m0Z�w�e�wP�#��皜eU���L��zL=�+ѳ�����Lz��kjd+u�ޤ̫�#/�QE���O�R��'�q�,j���x;�܉�~�c�Ӹ���EXPR�A�ź�rYH�\�� ���;�9���1���{g�v�bY`T����*T��H=��%`@#����6�	Y #g
G�A��u\�¸���g��-0��q�9M���Vja!T��d�?�=,��Q���]/)���+-�������n//���E�!�l�=�TB�YᑒJ����n��&�0}��*��\��聧s�l�{H0K�f`�O�������:}q�%�,d�yu���A�Vk����*C�Ƶ}+9|q �gZGO�#�Ol;�8X��CAK��*D|�a`�ZQ���������%78`}.�*U�|/f���i��A�$�תY�|n�zq���7N��B_���@~�2P���q�W�>!�����1��Iv������<\�"��&I7!]ڄ��S�nK��g�L.�&�\I��4��nd�������k��c���O�x�O��S�10j�Ş��V�!X�<������5/��L�@$m�CPDn ����!��ͷJm8X�Q��Ud�T]�@ͦD޵D�'��GU��f3t�mِ#
�{pr/tXP� w�6�,�]����-ȷ�E�p
��z��>9K��5)�Z��zdA	Èo Q~��YK+k��6(l��i	��3	�����CT�A�W��W�2�i3�E}ل�7�j����l�/d�%�{�5�dQ�j��"&�p�q�ւL\0H���z�E� �� ��Fv6�M�t<�e���K���?�~v4���e��rV�����fYg�!�ɞx̽������$_�>㗑nf!ܺ����Z=����g�Ac���۱��NX���>I�f�������5���s�	�H�Z��yN��q��9-�V���$`�ɣ�˽S1r�(���eHtaվ���������޳e�w���^�d�9cr%���+J��56�v���,��?�`zj�;�Rp�'��P<��ʉ�3�ę|W��P�G���ݍ�ڀfO2jEd."x�83v�����_�*3O��x�|�Y�i,5�e�,mc2���I�oU�|�zVԚ�g�������}��U���:��SZnΛ$�������+�����~�������{�0�����
�u9J�2��#9���v�z�(\�3�P�>�s֞��0������'Y+~TkNM���Ud�	I��+ &�W��U��#~ E�i%�@XӉ�=�m���%|/KՄ�RR��.řh2�.<�����x{t �����[�;�KYT�z��O7p��á��$�H@�&��[�Z�R`��>*Yݽ�?*�^�/xB� r3V�s��͡ļb�P��F:Ul��*Hm�3=��Ё��'#�I7U�Q)�0b�J8��bpg\uY�Ư-��$9
�>���;��N�8a|{wC���5 �d����t&�	�3L���]2{�j��JO~��U\�Jr��U>;���	c��L�gu(��-��A���>�`�����P���.^�<´�hK��?4�dU �O���޴���\�Z�*�P��u����X�_��IL�-01�@�%h[Y�dz�g��/73n�[�h��4^чx����'�9�>:�ɄF+=P˿L�Kӆ���ǶUR�m1����?��T�x�,#�]�5]�G��4 U�Ae��薆Q7�ȻvD0�W&|G����u;�9���C�@���rn�����ޟ�+f��Fl3�)��|е����嚷�h˸�۞�ۅ¡�.d���;S��>;&Z�Xj 
b%�ū� o�m�&+B�C��Pr�:��Bҧ��K���ޕ�z|i!i���[G[� �z��o�ie�����ҽ+p�SW�,&4tL]9	]�$S6$�Q�K	_<�&�]ZO(>Z��Q�+���B��:w�q�K�vF�BĠ/�0�����C�](|yu�O�=�4�."K��TFy�=@�e튎�G��+__���ı>U1��g{�u�@ݱ3�O���L��op+Ć
��M��F���E���Ю�DN�P�\X�,���Wya�B�G��[����3�j�L� _��҇T@���>� Np�M��|���ALz��e\mKcZn�JQ]!�U
N�����/s/�n���S ��?׻,�\��K�4J'&�+��e��(Z�e�uHj���|I�4[���W�A��#��Uxs� ]]�q֨z��l�L3#W�XB���zB�ĺI$:I*<F�@bD�?O�?O�^Mj)BM��f	���G��54K:<�'��n����\�~�p�8��7�^p��׷�d�s�,7�#�{#��RI!���S\Kf4�Ĕo���%�c;'���֘���ĵT�
��ILެ�F���lS`؈j&�
���H�R���?H��]qh4ץOJM���L_9^��&��b������Cm�T��Բ?>@�}��N+$׌ͻ�Q4kަk�Cr ���-�#��#�)�Fgw�a���,��|d����& ej�0��ǜ�$�P�<�mٰ��C^?	���"�8)��E��m�{pYv���Q�"�wL��
4
0�@���W��O�M��!�J������u��-z$��)�w�v>���v�6���b�i��c��,��6�韙ۉ�.U@��+$�6�R��jRN���Sӝ�`�VpA�����N��S8��ޚB�����ۻ��-d/ᬉ x�,�j�s�LEF�P�cJ<!B�*��DHF���}����n��y^�� c�[�z�ʗs*�����K�c��0s��H-Ku��1�閩����8r+�碾���om^o�d�(�]�D��Bӿ�Y���m�+���Z�����R�o;A"m$��!A(�z�N�z~�hV�Q�m��ˣ���+ZSn)���V���:�V62Z�)�����-R����
"��@�h��b.��5����Y�~ܺ�P�ya<pa��k1�9�Ɉ�e�Jg7F�*���	+��`J��?0�2V��` ����W�y�Y�P�ŷ���Ѝ�6��P���Ȁ??_��f�CB�=��9�(e�5V�x6����d�9&�S)�%�w�mX�7j�S )�n�f��6�"�P�� �����(}�'��SK����0݃/pJ�é�;��U�`�+Gi�:x���ڋ��/R�� z���_�~8 ��.��o+���JY�}T"�BMU;��?72v|u0��ˮ�4q�<�-��,Š~�~nb=`^�!]g�l"�`�S��ŭ�Ex�&k��!��F�<,EYY�U~^H+LH���injy5�����*��{##<k��{�&2
�]���O��(�$R�rݎ�b���S.�+ݔ�,���?���I�B�K;N?��XN��B��O�L��=��t��?���S*�g��{3U�mi��Sa=x�&\��HChz�8�!I"��=e��&�@����Ǫ7,�[���?��VC��$��2M�`����X�L\Q��a�D��ųFAW���c�V��վ�bEv�KZ�oc )	�g���|�P듺O��{]�M��8�u�CV�Ox�1{Dmh�]�-?�w~'|jd��*?��5��9
y�� 	�n���B8VZ�`�� 挫�ch5����;:��џ�1��x�/~\� jM�]�,}�j��,�w����ywg��188��Ki�"�ɬn�(/�xFz�K<4�Kg;Y�=f�)�L�S\Ҳҁ�O(��ܒ���{��;dh��hyɦ8� T�W+ђ�@��=:��&h'�Y\շư��,h�oevm���pauE)3/)V�84ލ@�����C:���
Z���`AP�j7���xʪꖴ���G�8(I�24����S��#Q���m���-�K!� �.��i���u��0���2��=-O�=Ε 2!FÁb,w-r��))%Jo�����0�w����-P�4(�6̡g������l���|�O�IV����Q�⚂�P�,�z�j����t����S棄����)'�A�v�᭘�7��\?��5��C8 �ծ�z�3��q���+�J�9�5���l�]}��&`l-e����2����0���+ж�FX�$��8�i@�E����O}�}��������G�9�=����HW�T��� ���7m�N_��L�����w7�ל0�)�=N>�����>�ik��7�I�Ui(1ksb����(Z"=�pz�@i��5s��ph�">��b>]b��f1���z�P�.:U�_~�2Vأ䓨B%�G9��0��K �M�wvNL�EyE���R�Ք�ߦk �L*d���k�~qi�+��"�!VZ��1�w$����~�s�d�̫��[��������HIŞ���ރ��G��!�։��;����]]\�C[j�d���i��O�;(c߹!}�Pu�de~��k�L�d߽s��!��p�i��g�V�zS'��?��ae�l�W�r�	A�t�N�G�3�9��`<�[,*�u��� ���PJ-ҋ�?�Í*U$
-��ӳ4�]��פ|�	d0tBy��S�?GN*�aһ��Dk�W�[�-�^!����SR@5˴�������r����-�S\m�\ڧh���k�7S��$r�`5=w�E�^C5�� �Iv5���&�O�ա<���#�|߲0�t�E5�C��5�uT�d3��q��ᒠ6f���ϟ��r���p.m�x����:�=B���k�����{�z���-,<�Y�@a3Z��
(�U�usp��T�=��J4�uÒS���e*X�T�=�i\Ώ��u�148�T�e�Zij���&�Am��w�E��%�E���Vc��ћ�6��rp+�V���e��D@'�*(�S�*t�AL�e���/F�w�r��(�;�=���Ђ���|H�
P��NN�n	s�@:}-[��δ+��(���Z:p̼���=��o��B�����*�]w%��	�qߒ����9_/�!��j�-�?K�A��E�6�����!�6��]�GSv�7�Qi@^n�"�%8/U������ɳ��*��m�������3wP��is����3$��P��$\y����O�0����#�tN�������!0j�ie�Z�:�U�ȟm}9�i����^=>�ِ���.?H76�l�[�߼
G�%X�Y(tD��f�GHf�/��T�]�//��Q8��x�nV.f�&$I?M��O�*S��h��w�߿��D��	��?M��<ٌ����r�&晒�ızb��)��(��3��Z��y�����w��He,�.�#,��u�7*�i����*>��o��v���b�9�KD"�6��Q����]��#r����bew$��	o�2����,F@n�5�=�p��$H��F�0kƨ��?�
�X��h���_�4Gs���]ghPGi�~6�j:�r84juGu ���猿ແ6e/��M���ۙ�
�"P�+h�%�qF��H�*�ES߁�3�۲�˛�1[���E/�x/��xZS$a�oU�
�Q� T�<Mzk�i��DV�e�P%:��0>���"#�mn�U(/]D�pS�Xxae۸&7���N�����yh����<��Y���;n�ݷY�{[M��A�ᜈf��Ѐ�u!��%k�?�c2�w�L���g�W-%�p)�K�Y܌(���j�Mso�&TM
&��$�6��s� v��Pqoꓔ�GF�[[�Z�5����S�3>}ӕ�;N�>�ƓF��'1@P��k�Vޜ�h�HTGS�u���Yss����@y/j �v̶o9�UP�SH\�G�����@�"�0L��	�J�FtWJa}:\F~T鍏�c�	����.�Ls}�OQ]vl�G�D�J%�qL%�̈��>c�2C� ���[^[��U����o<�/ɞ[�jAY�ΚC���9w��U�2�"�\�e��q�B�t���H�u��F[�+%+^6?����o{N]����f�X��_�/��	<���h!�s�ߍh[3�
ᾠ��O�9�>� �tc'�z.|F�?\Ѫ%���x�����Gۦ�`���d"b��D΅��m����Ҁ5A�!������s�|6�QiN/�<m��`��=�S�.��H�\C��o�0+ۺ�lcM.����Kll��ټ�"��=@%���Ͳt�˵2��Xn�˰t3v�2[��3�H=��#�G�A	���E�Ya�gS4ES�\��Z��Y`AH�~�+��ZQ1T�e�m\�S0�����������ݐ�� �fz��3O��]v�*>@'���Jȡ�J��+���J��]��#��#�,4z�y/�F�['���B��y$8J)S~F~t����{����������l����"@��gP�)�/�r ��܊W.6�5D�-���lY7a��i�h�<�nnEs�#Ւs����)�SUg���K��5��i��^���wu����e�Js{K��A[�4-~����̘*�y�^ދ��T4T�v#`{�* �1H�z�/���ڂ�_ԅ�WW~���oBZ|i�z�(k0	�f��a["{m�((k�K29�:�dM���]��02���+Dj�Ŝ��>K^�D�2�yCQ�8���>�pS��ѭ��X�f6[ ]Jӟ�&M'7����JHt蔺?Ԫ5kC�M�Vg��o_H�Pդ�<��U��(	����ΌδܐW�g���-�/p@�4�(je�U�08�D@)�deN�7b|�����-��IwD���	�߁潔Ta��qo����;�B#8)rV��&l��y����P1� �SC� 
��S?}�%���Da�LQ��A�-�NC- �t��#~�蹍�W�$7��G��n���aE�����c��݋�q �﷩��@F7p�H�FP8ӵ��.��/31E��D�������l����#2�l[ѷ���U��X@��s��ف��4K��<���� ����|ۆo�_m�|y��~0Yu$pK�I��w�m���=��!���xO���{��j��XGЌ�?�d8��%"��A&��&s�O��[,�C$�Gp���13���/�G4�/@v ����옻� ;��O����CE����C
F\)[[Ze��K2-2xXh��d�E�WW�2��q���Z���K��2]���<�^�ӂ>}o�n��3�J{��A��*U��&PȎ<v�9�o]S���w`�ȸ��/�40��"�< ��g�&Z�����M�:�
����+[������c�Y�U`0�\|�[-��|I�������о��t%)��.At�� �����W[1������3e�C�E0 �H1 ^�VWҲ�wxt�H��Y^�6�39����O������7���c��\�ߧ��e�/t�����K�`��3��Aċ�L)��'��S.S3,���=Z
����'�qی�@9�d��P�g�,���Z�B-XX������������y��(Ȗ��r(���Ef��/ڋ=70V��R��H�ğE��6���aV@�U��Y�ʤ/�6���k��o�d��F�r��7y~��n�fp����,Q(�#�,i��e!��b�	ge)��578�j1�A�L]$�ȃ{C���NWw�/&� ��%΂�I����oӛ��x� 1,*���/äMͯ$ډ-h����a�^�'F�&,��h�	����?�v�;�'j��l%��[�*�Йr_�B�Ւ.q
����Ck�m��wR Ӽ:Nq��(I�xz��U*���Ͳ��A��2�]v۫��� ɩ&(g5��r���$���1}H�4U
YW0I��lf
�[�=-�7B�,�߯ۜ���9c�i�w�㜩�"��~�4D�� ���g�����y��=X1��V?l��,�Z6�ƙA�EU�Wv�G�)���t�]D,g�����D=p���+Uչ�kE�@�W>m�s����-�T[7�|��b���F�Vȿ������u�w�}���&��mي�0?�2O!�CI���>"��e�c�-��-�1�1��?�&�Y���ٷ Ȑ2�	
Q��gW�/.|�lk�^U�J�T5�?\{�hz�-c(ٌo�rX��&zZo�v�BT -��Y�h�AVfYu����b��U�ø�L1V��J��ch���2�!9��78F ����A����8��o���hˇ0r̜��i^Xp�?d��4%ȑ~Ë5*������:�yk'�hS��F�C��'F���3���	{ ��[^��K�Q����#
o����r����ǯt!3�ߓS��y�_}.����y¡�QןI�1^g��
���ۯ�����.*�+��	㲐ļr�1
����;�r�Pa�p�����*>#c�V�"�_������OQ*�����wC��tiN&�;X�؞�x�(�x�q�2�7���	k��`rM}���(2A�lK���:�9���%z���،]>A�u
�4��E(S��;f�S@D��4�K���Τ@A��8�b�X�(���*��|�cq8�{9�B���
my����a�%p�����Oo��i���D6:a::5�Ezc^b@^�3�1ց�i����~�A�I�,��{�*���m�@�$tU���4�nccm�r�X#0���Pl�ڠ�F�����e?RD1��/j0��=|LTrL�������lsF��`������J� �_����C��_�����g"��	�4�5�C���.���򘟉��#~	�aA>:0׶��j�hp�~+��1����ݯ�_�L��7ڛ�h��[�(wڽ&�,F��2��+�Y"��`�ǲkd�j�ء����ƝwP�+�X��$mqoc~jq����')Y�䔮���)<<�b��A�gk��ӯ��'Wʶ�Z�
 �S��:zRO�:TJ�����*���N��ڥ���!7K4�� �=��g���XZ�ek�o�-��@�o��������S��}3#�L��{�=���5��=g�N��A�9�f�bRض0Z�&C��"���B�}�7;�������"�����Ҽ�� ,�H]�N஝�&�_����M��\�	Rs�;4;����*F��%�$F0��_�FjԲrn�9��E_��pXN�`~S
K�Ú:�i���(hQ���$���"Mw��2w�Ac�{F�:A��2��X[�k	h��#G�*^� �Ԓ5y�@M(���b��J�Ȋ�״'be&����$~����y�?�a�B����'%٦��~tS~����>%9&�������C�W�QP�_ח�n���_@KS �I���&6)#�[`�z�sD̩�������G�[��a� D�[PΚ�J%.����o|Ü<�k��s-�`:�t�2�WK�Q5����RV]�?��AG����.P����Ȟ��=+8`�
g	�_�[;���W�޶It+j����ʀ��Z6MeK�� 1W"9����-�U�9E-1��zo.P]��1���q��)�E��A��R��hC}��b�>?fC ���z!Tǹ��c�0d<
�͛Ei�}�N0n�h�͓��Pܫ��LJ# �ϒ�ܪ�g�̫�Z�7���ˈ�(fPNW��̱�����=U�?4�m��IT��R���J�=��]b3���^����O��[���/�"��%��$*�
��Q����īi*q5��~�����ᚄj���2fJ�%�#K��2
��8vdaZ�SԳ��.��~W�K~朇�ל�x�N��yc�i�uf�������-:�yh	YO������)��@�m���}}�{�x��'U�5��g��:p�ׂz�V�a*#l5�&�f�4���f�Ή��?�����ђ�^���ZPZh�\�����0�8�>s\���x�A�v����>�YM� ���1ֿ6B����@S��d����8�ӆ��~g<�~�N�4� �)��iē�IN;S�D%��to�Z����0�{�9L�i��~�/�u�T�R�?r>���"���#�l��K��y��O���tV����V�����͸�����2ɑ��2L^������ȗ�%;��b	��7�[��r��9���:R�	���+J��b��a�Mo*P�i.e�����f�j�aM�>��k�*���o'r��0ΐ�ԫ�U�+��Q�v�;��+���P��� �aK#��>q죋�3M���R�ʟ����q[u;Ⱥ�6�Q#�_Q�*�D��ژD>P)K#G����rzh�:	́*���m�nκ=������C���q�mW/s~5�a��<����ˆe�wC�=ț��=��tx����r��+u��E��~�ѯZ3G�FQ����I`3�*�ƣ]���8�,�#����I�l��*Ki��핟��Y����� ��2U�������B�9��u�`��!N�"��k�,\/��:��M!�])��S+�\�F��6��<�Y��
/�w�;����ҵov��-�EJG��DpS��
4�[n��(�6�{�npм��y$���~��െk^�u�/�[_A>��8R0I0��H%�B��3�\6��q{g1ý�q�wf�l�P��>l�<�-A��	Ӊ��_��0��~9�/�:�>p�Z��Ti`�vy�����v��=�5�MG-��ӡq�0v�͆~������h�\��U_U��`�Y�\7-m'?�?G��	V�Y+e2��-ODe7s���Km �򝹓���yp[e�/s������%�����M��ftS����%�[�#Q��uR���[YBk�2�8���d���ґqec�l�����&G�$�Z��=�F6��-v�oñ��${�����5�PGd�������#����2�:��;�;��m�͟V�%wK|�p��-vL(ă6����7��lP����w$���7����Ɇ��-t�v�w@A����P-1���"�������1�.
��zCi��ӱh�S�,���(��'�/�:����S�� �X���eW�DY��dX��HKy8����E��Kp���7���~J�}�*�V���>�8��@����RU�1�b�PT�μHL��h����K,�O�b|���<M������9oL�.��6�y`:ZϚr�6/���D$YYm熧ǖ�3H<��XĜ��f�g�{b'?o�A���Ȟ��DK�
zM�L��=S�"xr~,���`���R�Y�J�aq����zSr����ъ{��Ou���3N�n���ۡ���</3�yT�x��G@����p�:]�����Ԫ�'�G�x�S��n�G�<s���JM�͑��Cq�EK����6��t��oV�ǎ��b�����R������;2WK���� �����>x9�=��{ҸąN���OA��>�P�
*���~t�$�?=1��$P�9k��$'��-���0��N��F[�.��ͨ��6t�Q �
�:[�*�!!��Oib�ꔞ��v��>Z]���%�E[s��[�rBaiU�i���XĦb:}�������nt�TA����L�B7�H��{�.���� *�d��_!�8�	�:e��V��s�v�~A�D1�cu6�z'�C�������x*{����|�]�(8܍Z��"�x\�������aTBE	��B��[�\oV{�Ǩכ�Eu��|7�l�hr�.��!@���E��~7�N��|9�`6��"���"�T8AJ��X��%B��pV��"��2!
r�w'Q�7;W��i��O��0\�!�sC(�p�{]m�W�on����榚���Cx�yZD�bv���eNB�|��*	H�a���Iu���|�U6�=p���wh�)�WC^B;5���e�XqQ&'�h"�H�W(�J�B�[�S�mDŵ�FA�&����}D�f�e0�:}�����G�N�媶�b�����K�)I���v�U�]6�q�����L���DK�����&O�<��\ݪ�U(�< �y��߈�0}�o�'*f����큝�|�jz*@�s`&8��PD��o��Ҿ&�@!���,�� ��yO
�|.V����2��z��*�fO
$Ջ����S��S��n����MG<�]��'��t�'������wN;�����~�J�7|?�}��#Q�I��rL}ϯ�_�ٶZB7��/��i\*HA�1�JIp��#�p[�gŲ�A���޴n�k����K�Ճ���L\uX"&d����	�,\P_,���h�6�MC6��:7JL^�;Jԇ+p>�:�־)mA�$�q��b%}��\��W_t��/��'�C8D�x�m�)f�����OSj]p�<��U�OG�-S�ϟ���K��:�49�C�7T���#�Qar幚Ϊr\ʻG'�B.��T�el��yH2�shJ�F'���3l�Vd�Ή���K�?5e��S�ї}�Op��"
���$*�\,��f�E!4J���e9��p�ٵ<ޞ�0y^G�Y�`H�H�f�oS��Lv�{�X�b��-"槵^��QZ�S=~T�rE���f!8��I��� ���$ ��ϥu���*�O���b��	��&�o�,�g�a�2��ٮ��H�A煌~#eO�������
����R`&O83���r1�S>���7Fi:���G���?-���� d�K[�KM��e� Aw?+��������5*f�*�
��O�U�C�D]�`9������B��>V��29��ՎP��U��8�}�ѭ��o�@.�X�-v&�{�Y��\�����+Tŀ���
��J���|b�uL�h�*�
n�X��v�ث �>'To���d���۳�_.����Շܖ�w� &�]u���V�{d����`Ϛ�4�G���3P*�Ҫ���-�u06թ 8�_�g���2|��}�����*NLf;/�t���*fPh1g#?�4�I�����'�*�?ܶ������c������y���$*�B���m,m��[&Q-�g���2����Z5�nGM�2�J��$���ʈ�]_Ylƪ|:+������\�[Y��o�!g@��7^��e˕�2^�}������;п�!k��7C������p�`��IP�v�fi�6x�ҟ$Ԟ8�j�	���_���wp_��G�L���-�Ƀih�X��н��.$�ۛ��MP�U�̩�_�}d)���`�on��lP�킑��J��W�w����[-�2�mؖ�I�ԍܹ���
ML)���*fvO��gQ%.����x
��6��  ���J.����uj�ns�H1���9�zK1�OhЧ{-������qRq�]��D��r.�?Q�Ϥ�O9V���,�u+hX&r�8�~���7p�s�G+����Y��x�(�,F��J/E.K����B��yw�|�0����Ī����="�@an`H�%�E����O@(��":rX�ӳ� �IbĬ�w���p�Z�����VpR��3ے�&�wO3d]?Q���"?�0�p�6��R�v�v������Z����Ƃ]��Os�-hY��=�_$1�}Q����nhI����nR����)K�+4�4���5c�bQoG��l���DBW}n�@��4�M'8��[z)����#8��M��U��Ȓ]Ǣ�� N~�e��&=/D�9�lG�������� �����8Jw����1���bj��o���BN�4UL� �#)�O�����/�����r�bʍ�a]��Z�f�����	��PI�3�<5݄܎1�߃�y�\����ݣ�|.�զS��pD?|�U|A��h��~�a\r]�>���F�ż��yw��eݸ�zb<2C\��������If �귻I�N�_�!��^Ri��Ҽn�P���1��'�	�a� bݡˬ�8��&�D��kuT|�zx��K'�B�N}]>09܆=�eL��b��7댰%�b�Lox���UK�-��D]���n]�������}-���c�C_a	-nJag�3`��F/�N�n���d�f:D1r� �(g�yP�e0u�D<��O�O�m�G�峃5���$BZ����x��g��[M˥��o�
mv��� ��~>°��&�"���Y�}��XQt��K኱����d���~5#.&�U�.\��(�)��d0Y��r�PLR�`l��KZ�*r�x�HPP~���cZ��G������(�?Y(E���ZٵE��5W�1���4���փm�\����~s�!{������2#�B�5$�k�#�7(?��� 8�����JXVx'��wis�L<'�a�4�}�6灮H�՜@��̈�$��������Y$�[GŇb�2�ro�����d��Y��=�8�sA���&�~���-|��'��]�V^,�jI@Utd���҃o��!E�)x?�`h�y˿��<1kS�������7Wh��6�%���P4��f�W��h����7�N'E^Z�1T?�����2�n�����l�W;�w%A�"� ����#s٥Fk|Ǣ�����9^���25�ܢr���g|�ˌ9%z��ܖ�F��aᖒ���e�����9PBہsI�����ڹ����V��$��3�O�Jq���펚��/�բ,C��q�s&�T.�o^hE��é�4�3R�	�)��
Q�~#z������R�9j���ђZI<��e����cQ`��?��(bU�'?.ڔF��|��1�)P/��J���v;QC��Q��!)��5��I���~	���3GT�w���»�K���l�������/]9&:f.'�}D�൉��6�Û�[q�٥�}����Sш�v�g5���%ͦ����y�*/�m$��xA�d�Lc��� �K���T`s���T�tp��K�vҗ_1�x�ͪwڂ��+&������@��M8�ݨV��;'��X��4��c�5���������r�;��x�{y��ЋA�`;Y���"Q�����9I{L^ש�зBy��b����ܣ�.7F@}?"[�ٕ=й�"�����`�rֳ���㥡��;���嚀�l�%WC�[�!��D1P�b�z������	�;6��u��	�f��A���Stl����5<��L,��ʳ���)�话'5�y�:M��K�"p:��r�$U"�ҙ��Zٸ;\xK�P`[��0�աy�������	��G$�b_���%���0{%�} �ht�[�t��@{���68�����c��s���O l�8d݋�a&��Vi�e���g�І�\oc�gk��DC�2�0J�"��E��4{��×�j�9B�}ڶHZ������Q3?E�+7��d:�y/
�sٷʟ���w�u�7�KF�
� �qPگ�ԗ�ke��D-&BP_���n�Cvzy��h�y{)�&v������,@���iЂ�Ow�<�M�v��Rk��z��Xf�e��g_|ں����yՁ�>�y>+]n���0���(��ܔG���\!�n}����F���⨛�Tfٱ���שzwI�;qm-zW[�%��S6��Y����\�i��`�"��9X�r��i�̏��^���)7#Y����{�#�J΁��Ss�R�4�VJ�.3�"%]Y�j��s�wH˺ͭ �.6߭�T��V�3[oB� ��,�i'Xn\nP�:���P|�nF�H�㼑u�(u�iwΦ�_��:q,^D\p���0���I�^��*�=:O$!kTZ�8m6"���7�N2�fT��T9��n�{�l��Ez�����9��>?���{�A����i�g����Q�����Ǘ]�I:��eO������ -t/��:&z���^�5.�|���1eK=����Ǆ��8�Ԏn�_��P���#�GQ��d^Y�)Q�:a�#ār�~u,���cl�;q*R������n{;<ΙE�P�X�#��ե�M���2{�Ogȁ�QZY>�;'I[�d��g<=�̠�i��o��~��(#��ǒu�)M�r^	�.���Gߔf���1U
8Nh̞�yĒ���e��p�E�y���ף���
<mf�o�5I���p��MKɉm' ��<��O#in��4ϖ�����i� �T\��C�W���������';C���@��:d�����u��n�@'o�.C�ws?mڊ�a����c��E�D��c]I�G�<H�>��C�w�z�9.�s�Q�):�}��!ÝW����a���1�p%O�|7�o�.2FPOi��޷��+g��Ξ࣏(�>^����n�#ɫtfW1��/����̗x	I��Ʉ!f,��؍��E���R���5�1H~cբ����s��tG�b���z�y�r45�b�|���䕿�@���*��6y	$:ޠη{O5��W6�Aq�Ϳ"QOy�*�㣢��_M|ğ�4Q���x�����5:i�#o,E�1˟��ѺhH���$�H�ו׹���7<�\�YpV96̖(��hG����*���G��P�)Pc���gDߐHt7]��6��N���)�H��}�����/���u<8������H��}���Ў���Z6�N�{�:q���T�s�J �,>�3]��Z��(����� �z]L�����_����"Y��R�.��C�Z�$V*���<��b/�r�@&�)I]U��sЌ�/���$��DQ���T_l�0�@.�U������S���䎡�� ��,SJ���f*?F�����Wm��Ś)]���Hh��:����|e#�J�$6����{��dx9�Lj;��ai�[������ر��Q)s�3�o��J9d��.�l�)�cY{¿:���z\�z6���/x|��s"�MoDzX�agH�~����5���U�u��qS�\�B򊐝��S����N\\q�������s��Â�戇_Cб�G+;�z�'r�|����C�M%�o�Ȇ����0X�)�̕Y��g��4M�=~�#=��1�M�e~�u�2ǝg5���b����jp�)�1qo�D�.{�4�o�*�X��%�N�T6��]?:�T���yw�YR�LN�Q��s��W��F"������o�A��[�s�̌ �+����
�5���h�{�2��=,fesw�4�:Ƥo�P2Fm`]0az�=?�3�d9]o���%�(��+�_�H���e�vi���v.���U��OB��$����<�5�:��8n�v���Ⱦ�J2bX��,�9�)�5=��4-��oo7;+�*&������y���ÿ���J�d$7,��Q]s�!��"{߈��q$,�Y$V�M����H�n�d���|.���������gȽV���	����Le}�Gh� �[Ď2�[�U�}=�qdr����j 	i�A�6^宲d�る�(�\D)8$�
U�'��P�`��?Ø��0z[p����PF�܌���L�N�=z��roтm������OVw���ӗ2 �2��w�+���w��s�ܧ\�<7�Y5D/g_6շi�5��_s����heh��>fVh;b�':R�C�`��&0w>SR]Y�}PU��U1�K�T��$1��i�]0�#:��-��]UuQ�Ks}s��p��b�����]��L�yhl�ēB$Z����7"���ȭ����20�}��xZ[�*\8������'O�R�����@L`z�&<JW�� n�[��Y6sN�=��N��jO��|A�N��>!s����/���ޔ�됪��6�:��+tp�Y�m���d�f�m�TD$]e���K1�݁8�K'^<�Ȫ#[��!��W�<p��f@���CN�%���`a4��Yd}����r>+0�.���Vh�4DW�W<�2���-�hs���N%�Zx���)P�l(�`�P5&��D��L�Oҵ��o���հ���6�|���+�H��=��<�{"/:��q�L���X͸MJu��C��m7���9�^gvk��9�8G����^;F����h�:�X%/ �=P:�����7wmvm]��8[q!�����Y_��0�i�o�:żA^�Ś݆T���A���J�F�G���&�jtUv7�������4��ڣ�yQi~Ͷ
�[X��|Ѷr�6ky�K���_HM��g��� ��0�I�/�?ԁ���^�!(�'kW��d,�L!~�Y�m�g��������SP�����sj�:L��5o�S�.�#�S��5l���I���.��@_I* 8)�K���V�8g,����lk���%8#u�0�Px�@@3p��ׯf���\&�]��Pu���`Va��<-��QR��%�p���J�?�Dv����1��f�5�~��0Z�6��]V�4[dY^��Z�n{?���zUB-���Mbިb#I�jO&iv�(�8Վ�����4%��&����%��J�g��w3]��!z�=է3w�t�X~����V�A�� $��2��q�쓜��w��$2�bN���s��[��H�P�� �$>^S�t��݀��!�������=7�}��}b�j�A��9��F h'�z�u���,!Z�R���tz��:RV��������fȨ]%2�����=M��@!��+�a�������MA�����6�@���O'�
�N�Ѧ�V�waj���Λ�Y���>Z�g=85�>.3���&sn�S����k D�I.���ʹ߬����2Uj�4�%��86��p��U���q������L��A*���N�ԡ�!Ls�9�m�QoU�!ʦ���lh�O��A,���Zt���<�'Mq�$�녒`��o[���R�]���`&�Gsx� I0[5p�d��خ�i���E���� ������ر���W�-��}��@f[-n��w��o�	��Ɖ�(u��^�M'�p'x�W��?���Ot��:g�|t��d+?�U�)�_/�\w��c��'�uy�"�dq/�T���(��I��5�5/ƣ�N�!�X�)�Yd�T�bu�/��q񼜖�&�bP�J���6dp���t��;�(�� FI�1<��������������X��@��y3�~���CsO�?����lts_'?O���3��"�_d��b�8e
�Ж@~7�n�����_lN}VKPL��Xr^� �����$��u����1mP��tK�����͟_�7�`&!���.�/Bٙ=)Rg�%B�u��p.�[>�ݵ{�|���V��@���W�<[a�P���:�����4���B�~�C'.u��
0D�qq+ĉ_ʢ�/	{���ya�m��:�_�?$HsMؕvPӋ�z���x_��A4)lK9R9�eqH-��p��k	�����Xr?�u����/o<�����\��$1�>+�Ey-�g��~[ձ��&���q�`_�$}�Hb�ۀ[�(�N������ӕ���oM�����,'n��V��x�u��hT����t)seې�B
ķI�b�%��(�>y���a��r;	�^K��~���I�h= ݀�;���]_
�KQ��H��ݶ�=g�@;{N�*��Q��g�˷�Q�ƞ�M��dS�is��w��y����'�4�V�~���97=�Z��ӥ��8����G�ӶjnJJ�9�5f���|�&��I���RAw�N�Ϝ�ʛ�)ȒGW{*����R=�_��>Ͻ�r��vp#ҽfs�:֪�'����4V��\��ƞW�	��~t���tH3�}��G$_���"��mW���!ƀ��7%����DG��&T�,���ӽf@��>��JB �������_�c8���<�T0L]�ꇧ�����^�Xҙ~�a��cY�N{�,�6��|w=����+	$�AJ/�V�|فK,,�w��9^��6��Ü��o�=��hnW�"�ꦍU���0mG��
����܎B	����W�|V^󗑿2��$N�E��0i���2j��oS��9�E��g,�n��V\�@���-OT��Hr�o�����_&@{Oє�7�����P�l�N�r' ����jf��,�t��ЬY*N�(|�,�A_
�[U�R���a�f/C�g�v_~�Gq�����,U�p�����0Q=)�2��M[��_�ܩ�N&�����3�^��<�᜛&��H�T�&��@������a����u��)��,��/����4Chi��(r�Pr8}y}9�՚��?+o�d��n��hJ�qpg��1�0�]ƹ���»�<���xGS	\���R2]'�3��.pٱ�9�Lc��|���A^�0��6�S���m
�^��&,["3vT�dAwV�ۙ|!�e��c3�9��U��#S�\x�-lM�
����X)�M��	E�qH �o�=p8�Zuc�#�v!�qJ�F�־���	�K�h*&�!h�r(�.�ϪLAl����Ay>"�ۮ�\��<��0�fGd�J���%͒
(��)�H�Q�:�c��z:�.�@H��ap��IF2vf]&C�=K���	F�f���P ��GYW謌����XY�|������vR�}��ޢd���*Oi�$?{s�������	C
�&���s��X-��J���@$�p���#¡����� �Y� �D{��j=��\�'����2vG���\Rn���������~-��D>�s�M���s�m�:�>Ȫ��Dw�VAq�$��[�}nP����j������`�ٍ�'�V7c��=^����`�b5��E,f�M���`��I��9-��k�{��Xz�"�"����������q�8���
������RK���3�5���+V[q�t��,3g��(��7�{��-�2��>����ra���X?��h;���Tu`�ł��i�u��5�e��!��;V\&�x��dQi������Q��x$�Q,Ο�4�h�� �|�J�Z �}~lR�� ��0�+�� uW,�ɳ���ި�~]�������3+����$��2!5�-a������b��d�jՕ~��F�mi�T����7 �D$c��x���{l^&2���� Q�j@��)�nj�����9�RfRy� ����vsՏ ��$���ʥ|�A�h�����
#2a��C��]/���nF���V�DU��t}