��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���q����f'����U�S-Կ���Q@	�Z��*���������=�0 ��w�t��n�^�g������w����3����{p���I��'�/�qޙ����6c�r!��
;QN�A��,�sP;N��@���m�����eg��,��gm�-�ߞ;�"���%M����SP�y��,Z�}X���w��mBS�K�8Te��5#��
��mj�:T1,���1�����d_8���Gbu�h�$�_H/�Q�)��G��v��_3��z]�L��p�IB�4ݯ�z	
�{�r�H  l�8��p5�#�8��E8��A!(o�R���.����?���CY���
�F��f�9�+���q.6�i}�c\X�p�F�]
�u��z��m"�E�W��\�D��J_��C����ǧ�(C:�yFnP>�ù�ĥ���<4���V!/-e����`]&�A�5F�d�br��*�a��������U"#��ܘkYh7�����v1.���������[�`��[�x��n{��j�����jipj��U�A�|��q�a�t�IU�Gx���/��Q���u �`ڙQsp�#C!T�X�<�/���1Y�=1�"��5i�f[�7�t�;�߶� n
����Cą��W.�(b��k'�5oˎه�W��44��������Ιiɢո�ڲ���D��"H8u�Si[S��a�4����Jv^9�o�w��n"}N,��B���>lۥ���oVy*��_%���NkŊ5��80�TN��w���g�>."�$��?�Ñy�+�{��d�c��ʹ���������9�d_���k�IG�40�=_��g�T[�K.`�&�؈�A����h�o�}��.3Y��s}}�Z
�{�%f��-�Hͦ$y�a�/�1��܂��(7#�pĶ��m��u�xaYa�U*�����&!�g6gN���o��I�Ž�J8�*�ؤCxghl�x����Uv'�0T
�
I��,Ԉ	2��ᗃ�i 3�@(׸�\�|*B>p�ja(�?k�{^�z��鬳6j��XA��Y��DPۺ���ə�&��χz�NuQ����T�wf�v�t˔�l&L.�E�H����5T�%��*�g+k�Aω�U ](~G�O�־<g���)�CA�'���%�s��f�S«e#� ���t�G����q��k��z��[ā�m��]���F�:�0��\�W�i��6��O[�8Gz_���Y����D�L��������2\4~IJT�4X���U�ъP}�ɮ�z�n�U��X�}���W�o=!�¿k���_	Q�
-��I����������	W��W��f;?s}��(�e^80Y�"�{�����i{E-G��ǫˤ3|�'�U��`�N￥tγ�{�Z+������(@�� �^��f��v��J�����@| �&���A`�Ӄa����$�=Yއ��'y<�'^9��~�fƭ�m��ص�H��t���R��S��5K:c&X �`T���C����_���ʶ�Q�a�+4�g�<��7*`�?VV��?��s�Qs�{�'<�|b��0|�M�ҜJN��ͻWb�6�1Q��c_��?��#�kH=���8����X��I�6H�=����iM��M���] �}>;�4F7N�?�����r�Ie���w�� �l���D��8������Q�]���*��
e&����"�7w'��U��o)�p�QG�	�'-�ݗl��Z���_���PF���O˗�9����W��bI������)
Ѷ��"F�V��R���[�'�-��I�@�b�KB�y�c�p�s���#f]�<ؚi�GPx�iMT3�RҚO���jl1��	�u��z��-�G���!��+�J^��}�ٯ�}�0jk0�ZT*��ϻ��9��"�0-F��P�f7=��ԖL5��p��~ �؝c�g獿���Q`8ȬB��w�\�?�h�^�ϔ�E��O�M�"�Ț�)2̈"���"c+�c�S�o��-�ɡ��*K�%0ns�*p�)@|�7$_���VSgf$�%�Q���pPU ��
��5�D27p�iN+4ҽҁ��0J��:�b��MC�
�.'�zǛ;�t4�H�@#Z
���%�0�q��y5�A���O4ST������u2��q\�&�-�d�X���p��d����P����8�kܸ1Mz�U� 6ʽ������ϗ�(4{Q���[���:�������d���+.�S��K�K��ӡ�a��dx�!w!�dp���F���J��9����$����s�j1P�8C=�S�sE��}����4��#���;�*��ĩ����zs��*�-K�#R"�(&ЛW�%���)��Ͳ�}�)�+�C�aɐ�n�b�f-�xw��H�������J�š��}$���Lv���ۭ[��ОjZ)G��S&��w�v��l�F�E���-�)������ڀ��S���Q|`�"���QL�C2V��uh��G�Ր�4s���(d&��ZW;S<������������s��h��nQ�����[�� �[�X�)u������o'�;3>d_ȁ,F��xh�P3f�H���z:���2�"�5v_�����Ѿ�s�0����;��*� ����ГR��r�'�S]1݃pk����e�ޜ�&p�0J5�_��~<���q������z�}Y