��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,����۝�gW�Z7��?-�h�wC�|0����Y�C�PbX �HN!Z8���9C��>C\c֗�C�e�[QD"4驑Gu#t�K�]���hJ2%�9�=�xJ���1F�̢�;�#��anf�-[�K�:k�%~�K�r�,.�h�����S�0hZ�8��s�E�h��}[:E~��k0�tbK�+ޭ�j)��,�cL���SN0��tm�� ��z���DP܃���g ���9q��Q5�Dp�%���[�����i`6��i�Wꗟ�ToH��ű#��!�$�G��t3m����C�Ǡ$W$��6�ě�\�����:>8��<\��D�z�y/�%z��xN{� ��bśp�)�O���q� �<U�7��EOYk+^1Y�m��g�z ߶"|O��Ӛs��lkU�u��_�\�V+& T`��*K��86�oh�Ȼ4�B[ʞ//�w;�Rfՙ�����ӢWPa����}w�iw)�����I���?oAl�7�[v�騏ٙ��z��=0!ɻ�������ț��?e�����*m�MN�ш��b5��E%�ž�ҕ���g���^Q���X��N�(�䅩�>'���ܥ=8u�F�z��D�{Ͽj�){yܢ��o'�,d�RCf�j��bځt�{lJ�;�Y�\w�D�lFxv.͖*���ʷ���v��6�C�k`��H�l��#"kT��2��zd2S�N�8-�'/�CJ��U��;=rĶ�f�����0�+��X�U���!W�Ŝ->)`L�'���r<�Ô�ƋΌ^<f�Of9q�o�Z"��R��T����Nի{�_1�yC�@�$@�\���y�@�2�(#��`���k�if��is�F��ۮ�؂#�a�_���o�:�e��}�:������E�Y���5���S/&Ñ�N1@!�SXp��s��xg���wKC�>�$s$�?t"I؄�A��_�P���[u�>�$�(w������	x��ۿ�j���J���� �Jx�t�nj��/�G��p�a�L���c�V��k�9��:{¿�q�<\��1�v��*�N�͂���f�m�����5ӈFlU8�7�}�V��D�V�g���T�߬m�jp׷��Qc����8� 2����t�u�{��4{eYp�[T�@�j`V �}Q2'���U��H�.V���Sg[A��q����i8.5u�<�H����P�*�.�	CV|�W��dz�OMa]e+��t�{dP<�>� �Wv�����w�E���fDN�����~w<��#����7%a���,��o�e7w�1���{�]׬RbK��k4�H�97��Δ��y`�� ����	~��E��!p��<�/�AT�Ҵ�5 X:H�W�5�w3�����Kp/՗H�L�6�H�h����MO8,}�"�1?�����.yR�V>_P�5�?����4q��*�hc�ǌH��J,1�1���޴�1WLZ��Qw���A	DaG5���8�����-sm O,�e���5�Է�k� 5�!��2�U��ykΗ�V�Ҫ)�DLFZD8��i  \no:_�������h>e�/]j�'N|ݝ]HdiJ�吟qR�	�!��a�Ib��)ш5.�߀�ؽ�,��fwOsg '���/��C����?��̿�cW��h��7g	eP�l k�㕸|�hƚ,�3Iq��� �����|�����hƂX����,'=D�D���kC�3x�h�q!]��J��|��.�u�	��6rоO�:���g2��S�/{��Un\��G�zG�PͰ����D�Qq*g�8���,���Γû�,#}ZVT�]�ջ0��G�7�ps p}ƌ����҃F:���!���H�8�,�*֧��Ih��;�lCJ	�O����r�_G�m�u(�����׶�z[�(�kn�\=BD�7�;䮘� 6&�jɬ���'Sc����hH1z�|�s_����c���q�$ 9�/1#؄���>��n�ѫ��!�(	��ʙ���o��$����e�{���^�x'o-8=��Nr���x�-l��R�Z�W�'l*�iF�>����ߚq��?��w������x)f��t��V�kQ�gc�Ŷ 3���Ę�Ef�x t�Q��8�Kl�~?�2w�6{���8���(���
<���`<lg��`5�\%O�����	�k�O���}�Y��y�1�I��}�:��2|�)\�V1)�~���y�#�����Js����uhטR�e[��e�?��o:��w��C*���|��iUf*�L���B���h��8��v��Jȑ���w,�(*��uC~�Z���|��Q����0����N���R������/��.9��_��
�+���sڢ ]l�p��L?P�����%D*��a�n�@��X��)������Mv��6(���z��э� GaP�,�/ׅ�y�뷆'{�#7 -���>G�}Ȣ�i��ggO@_�����x}�@���M�җNC�ۮp�β��#�,��ھ��6R(g$5��X CzH�C�3y���M��ׇ��g�f�99h¹�X���0S��'w��\��o�+6{Kq�Aq�T�6Y�i�]�������E�B�����Hms�0��L��C�X�����6�}:gD$��Y���V�Ԏݧn��N�2�VV�,�׷]nA�eE~kr�I�2�q,���Ō�[JMKS������pFxR;,�X�ה6^uq�/�&���aON ;_j��?�/�꾪|(|�"Pl����U�.�Fn��;�1ZH1v�����MC�����݋�X�I����K�������F��@̀Ӯ;��aKzz��hHUʃռ�M�nލ]lL|\��xd��t��v���|
�������Ƌ��%;�k�bpߞ1+��p�[� �<�v��2P[��h���D˝�],ɼ���r���U�lRM��~9څ6s���L"�=�2ې۲�F�;-a+�d��i�����@�CJ��!�Z4X����T�dѿ��5�����x��\���֧�ܻ,�6�g�5OR�"Β�K�!���AuM;� ��"�:n%ܪ^�wB����F:�e����%�(l��Ϣ�3oV6ʒەsԬiry����+�z��D*�R�L��R�'����&<���S��U={�^�ؔmxʂ�>&�.���ˁb��
܁^��V��.<��:�\�m�9���(�<E�E������%�Q/,Sꌝ$!�����bM)����I��᭳|��"�=�	�A^��뷇�5�˝:��Y������%CQ����we�}
��u>��0kD