// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:40 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QWKMiUb12cx34b5SUHZ/btqL0n04b/GlLpV1f4g8ghoS2BffPGKMYRXkC7M07Gb/
6x8NJGCwNZlF3256kkRFJvi96bM8RGpzFAhmTlljZp5ukhRiYG61Lq7/PYeobibq
lB2JrZl20ijryafSlfV0yhXga9hj934e6vPkcPVx71U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17120)
2iEvR7PUzgr+4Q3ViuSen/SvleCOAiAbpOWm3JbHs0mbxpDwy3P/V3OGXlSCb6mi
lbNtBGP8FTz86cU3CoEeZndhPwgU3aXmFz13CiYM6h2rbV0fuE+WCLgPYMOYSP+a
ZViA12XeLh3mioSCpE6uk/AHpbzhGPgBBDVHla55GBtiDcdmLRcBkFnSc8pS4P4w
PUVd0Da68OrF0ZeW0QfcIvUS7aUTAILs4CWgiHamC+feZy6g2pBqiDvCtDO8TtI6
otgrnH9xIzt4iRq5ln3okDSAcfzFVtupFtlO8Pk0q9aJQEsjjP5dcu7sHajlQUce
d4tqTuRVMFmA4BEKH1cJNyfkAbpCCp8e3t2jIWsrgDKXpV2gLxDSPF3TP7f52PcY
zaRMOihlro3N9VtYNacanYA0wySWtd0EzjhV9NyHTBNwvXYR45vrpyUZjz1LslaP
Hddl5J6b2FqqJQLvVFuAMlIfFh+iDXqVGgf6GMOQGPJImtRMvDo/3pZMEQS5Ucm8
oFl26z26liILjalWZlHQjZDWOHeedJJGnKLlNR3qX2wPhWJUO0vkvzPuBTwn5wzr
AcMZSQDUIol46tDOHlmN7WU6V3zjw7P7DcnjqPUCsp2lvTiCni1hND9pMrvHwtoC
ihW0d9lr8xFfatw7ffRXT3FQebtJsAKRyb+j9FMW4MyPtdT5Ey/nsNJD7WODOtaT
a1idlHfZO5uBjcBvfv3+uf621Vyc4Swh6fPdg0TE8mrQ+3mHk/DgkHlrvHy2xSW0
8TVc+sKJZLvFpLm1u1lFs8Ix7m9pvhqgTes5Jc9BhCfIVnWW5/WZHzBg0d+6etX1
262i/Iytjp2pbaqU1/L9vc8f6JiMy/3qhe5tGRSrDKcm++EZkSs3lEUJgIIdc7+Q
oyy8dUk9Pj3BkS5xLnRybK/oq8rVG+yYngtwGg4NqsZ0WB782+gOIiS8U/1R29SB
SMdlux9u9PfGAS8+e2y25W/XFBEuCt9QuBKDRkd2KB+7V8PPxyFjJzP4Uo1Cp0zJ
MKE0ZTOfA5HJuKd69J3OsOhKCciXfMQgFiOO6JQnz/VMcqDLp1Hir/M0TOHVEg9A
nED4UnNxpZ9LQeEdXgswaApJGXninRcUDseUXt7vLHzuxmhMYIeP8T0ptBQlffyZ
aLpgsnyPgdRplD2pjSJ79JcFtzQcLPJLxC2NQbF7PPMzmZd9LFTKuAfIAXugoIAN
g7UgoMqhBTu0n9h9g8IrQ8QSx9t6o9Fu75WeSj3JKTDZtexSvay1ZfluW9eKFbRF
DTnw6N6I/14kIe9LBnDygeo2DjsOxBQa03JtQVm3HUa7nIZjyc+mjrOuV5ZZ6Pni
/NJb5nsUvmziVyUg+OGEUy59NB2IkeUXPXYXpIuw0pIFlKn64S7w/XJ+oo7Z3dvV
Vf3o4keET1QaRz/itj4EwbyG3vxPad1WCLmiBD7uKggong4BJiGKYwlLYPUK/TNp
os2l9mFxVMe6pa9FMxquIuojJ2Urw/PxkECj06h6ZqEWLtAyPgCHGPPXyf45yvbl
+oKewq5HrLrlhzxgi37ZaIKBwrW//jkBaGzmW9bJGREE0JdDX7U+ammFLQvidBm0
NlNZTXGaXHpVtBPaZ3fbaMCqir99uK5gro1kr8yNY1wN7NYbE2vkWiWexIMbw9zc
fD/IhbMdWXR1Mxk/FOZ8kzdNMPSe5ABlQPIws9XHjUQ1zCrTrvuwdLYlQeAUStUL
gAdE07ERRASRD93N4SYUKkdyAemCW2wYaU+yIxlkLCnDApaMt6KnCD3ZUAQrERWr
CTINLHP1e5tzmAdLv9lUe7oMUD6c4oNM+3GFsgfdEulzxGlfxww6eefnNuMIJuZP
gNog98uJ1E5/ylze1H3Cxt312UByvnF5DRTgUXFAkNbjiFh6ZbtDxD+P1MxjlR6J
rjAkCNM9/COqr4CgEjhFbAHKlLEYX6tu7wI7fCFImDW5Efa3X9BWf2Os60+RF27Y
Goum7lv8IKe44JDzKJFYHflZbHQt2n/zot5muub0gFGDprJEGTCQl8TM+n1bJMMj
mNyuJWJTUS3hWL9L3P+CFIyfKDadmgdu5z1AYbQDjDnQNrmAGL75hLsnDdNPG6Un
tBO3z73omATpX2C9LOUS3gWltFWDy4oJzejzJE6k0m169cFgvZQOLvE7jKnfcz8H
eHMtvAqgXRtM+SZ6rrOGEBScBKofZjLfy2VXveyYTGk2HUmOwq3rgwcs6LvdtrQU
SdN87yX5mtzryGJYzwfCXHL1+yulK+GJ2Dnx0VgoWA+KTLJ3Kuxe4+9BusVu5yM4
12QF/PtYdYccHj4+sc7Veb7KwS3s/kJELLJiMH8209I4bwvK0RFbFIf3ZHTaNm5n
OoHdUbXT9d8hUbAvpz+yuIofw3y7hUOTOH/xVOO/5/qMMtT4F30A5U9wYx2LjBka
03FovtTzx4cn604kKR0ARDw1VZHadWTBL60mHXFjh14Jo8AkuRnllVY6imHCHtOF
he/Zc2wfkTAFPoV91wNZL/Zev6ys7osEk/hLDRp9sCtPNVl6H/RjD3EUn1y8hukw
52aW4xGoUFyuBdx1Wtf1rzqKGAWVMcY0ZMuiyX1kKE5Ej43Uj0uFbKR9B4/TrDb4
iUWQzWCI8SoDop5Z/6QGbvR2HsnSd3pP/0neqN+4V2FBjahJ/D7HlEnwlAxMb/hM
WmSVDqYnwnyImZ9YySuYG3esfvuRB20q3XnwfoUNGBtQJsfBJR0dqvvVPi8WP2Sk
mejskaaXM4U0m+cG1oVkPD7O19GeoGkBwdRCe3vOkXlZFFwe+QrCz20L7LBDjHLZ
DvmUVMJeUNq6TxcYqsx05OqNQyYEv+wj4cThFsl4OJGy1udLNYU+91dmbksyaZVv
imrX5cs2gD6RYjiEM8e4gkmTwgRCSzIowtQGe3DcXmV5yJhm7tC5KVeS2nowh7Nt
8V5oiui3iWzfvfNoRpelxVUjTLXeNGGu5hMtF8Hm27lrv0t2RtXpeBi/T78gkMjx
LjKRupMeFlih0kHMxOXy1zru040tvv1qfItJhm82vart9cni/N2JsZHMNtno9i0W
ieo0/kY18RnGNlZoGuoD5/M9hNj2jPriJy4xs3tHSLSbjIlzk42xOObE7W85VyF7
rCj0cgj8mPzgEaY5biGQMjzTvDUAmRUpI8CBlvUBBfLjq/hhTEQIm/oYPuqEUWw/
0NvHKgOWfwW2DTpkfI7ZZkRrGlc9QIZPZF+Gl6xEdgmyx0oV5HWA30uWN7WyzQrD
X8SSgAMgj2joBGOFc4beyjF3IBqeBauMBlLATx8BvedDPdzzse5Ix9HRmhzMDN7b
oLVvYHAfu0OOke6+aFEfNCtXaRMvuIytH/kUK0dnHr4CN8+t2Mm/L9Qko7jvMELL
aPset7YxO/p3E4z2z3cIAdH6TfLjsaQWqCi8fJgRwNATK7tbyrMuIH3X3jXFJJ1k
RrShDfDhJIuisaMEeB+YacmrfIdezMLrM3tZCGpO+EjXUOx6/rTzEV7/AG8cDLcg
w2/qvkKYAASTLLPvSfZJkHb6wiwdD8wEfTjq7kDbUSSJyklhXzC1KTYku49H6M2U
vSkfAPHtXyLHTYh7L8cz8SgzdYoo9tyYjMx7m7xSw3FlLbi3gUj7o0G6z05/IxZe
poQzN0tHAoZs8/0CJ5hUGknISN7YkGSjAYGaQkOokilzXn4bLgcaOI+72Of3H0KZ
nALw42/9OEtYyJMOUQAHPxnqhkJSu/PAz+46+qlZyfg8uzYYwTiRvmrq7zUwH2sD
QxUBRlKU6bTPwb0NvZG4XpWoc3ajsVR8yQqvNIP5KHUoKIpRHhUkO7ywr0oOiAU9
YAU7yfk3REwA6Zi/oXZ3qOjKXXKM0aRT3My5EeUOD2lkD0YzAEIf6LnmlMMrLWwH
W7d+4vGk/XOkn+YiVUWD4Vki3RubuDa7N3jyJ0QvoelVagyBsWrb8orNAOJvDeR6
J0IT0lBr48ktIclHtzgLj7HMNSbnxdwGmWclu1wMk45JafaICAVfy0V6HjNb8uau
TVdp+PZxTUElX4Sd/QiEJ5/3/5COOA7h5vo+EnFP+pEXL0d6j80PBSRgNG60V5Jb
bOFF/JVurtd1EnuxsykyRjb8tL3x7rPDBKE5czWW/Dx2/hriwlHQpF+mvWZZccLS
YaH6WqJ/UZnnYGN9Xus7/aa4yadchZuaKiHHKCigX/tCmAS2YA6jXJjDIN4xI1W4
T9BFTOJ//zRtXJq1qDjLKM6rW2dwGn8jk6EzXT1JxatVmnoMlxkA1cPpJc8nbM72
kOO6Lox+hHcVlEuYmIAdJEwodGWNMucgGO+uwPzFxS23Ei5UXfksPIftAJGHQXZ1
xYUGd9KEnWA32/DDSZimxqoIbsffapnw8f5YjVvwtNug84gS6tcvjwPHss0/sp2j
G3Pdds+YlSYpmyt7gMv1uA9YnVyoFfiafewP0EW8kGJqriA2cTZM7KWWDI+lZwMw
gQOR+b7SLjLbLHPD21Y4osk6r7zptQEYzCVj4Le/ui3hjnvfdMsHs4K1Y3CbQVrw
HssTQG6SkErWL1sG3eKjZ9WBRmjsDE5UnlDIQSwD1hvqnJdQUENwJNE9ZbWNaKQp
4jA+ktBO9tuY6ERM39oYWHNEurUa2kJBqAkc2ubOZhjfq1Xfef5X0A5Rlv4u/AfB
fu1LHJdEHdR5vbxD+0SLQ6H/jnZIOiPMt2vIN1qUS3V2UZvlLtsqfrvKOKhP4pSR
KZN1Nanaos4feVbctreKNakMxPO1hlcuCMKj4ijTEBJBKr0Xnto2Yj1kFH4YXIsq
sl0Och9KIysyMuR/hGYdT21bT4gPXMEt4zZE1HiZdMczKG7S5v7z/cNmmeLHMVE3
ZqC5Pivm/jDPMR7qez0hAag/BnjcQ807X1s00ushnLhyqomrAYL9DWpo4dvJwnAr
Byh7AoyGoq72tQVnj675EmJuWqL7JFd/FgPlAcRP6Yf3sOHRXJ5C1+om//gPQUGx
PWCnqrnnTEv2dcCXe3K3sjwJKGDO3/2WBwmfA0b/IxfnR69JHpSlbzYuna7a2aCU
Dxm8CwOrIosCAexYs5ZhXs81B6kEMgJmUbI1XnJKSEUUzRUqRSgTqRZ7B6N9c2CI
UanAWbqCVV3hBzESjgsgtdb6kzrcyJTunttAhmxJbtoFah7gmb+E9dQmj5S58nTj
RIvG/HITFX+qZOyIU7E/OGyAjZyVBlgkk2qyBT2DgNT72SDBDDpDH7OG0MfhDJ3j
fe+PaibFJcnZMLgnDPSj4jbpWDTKuwQC+OfHVIY7sL9Uqaeo8gWtuduLjkVXV7GR
gtqq6bSqmIgeaNL2NwHZfLlIoCettV2gTDY+sFCI8OPaoTTsXuidITShnFsz+KL1
e+5gBC5TSPOwof+3BMTXqnIhfZJ2K2wiaUhwHNWXZ9ev1+pxW+zoA5c2F51IJY2H
lXr8jlnIkh68wRLar4r66MxoWSpIbF6Tcd0/48xEIWxyQ/5IUpd1/Uu8QhltpoSf
0cNFlctpNO0hdQgP+/SgsaxKq6ikci6FD2+bMLGHhwKG6okxP3ckgAC5n3RmlXXO
FWxsFXKlxIhmncNZGPjxzLxGF8+SxNNrOniU8HVIaxPm+ouGP5CknXXVjlUNPmVi
2K11d1bfD1PF9Fr1MpwnfJ0Hr/n5AB4IyDXaG2cW3ZL5bpv4hIWnzXV43MfZBZ1q
CjvO4m9S+l3pLrA0uNxKh86CG3/z/fZk7GuLL1TD4XJGp0H2UQuLycY5LIAz4dFu
oSFBChbS5IicSGewuVosPfHHUNzYH3Y7zqpky1ADM8tFDDKRqKP1PqqZmV8ZB/Lj
doq5v5GKKjSxVKimy9KcP8aJjjJagh7nbCcme2xU6RX/E5+BjWUltX43SS0TCyuX
VYbChedEK8wkbLeYEDHnAYW9fjtwZJBSthSXis6mlx9OgwKEdi6iEwaLtuU5XCQC
esIzUR8LCvmGCcv307wPAaqgmo3Pp7vBaCbK/gv2uvpg4LWXZpZHo7eOhnrNO/vI
k3Fzo4+Coho2OC3FwhJJwLelRo8BF6p2STAYDsRpOTcDBgHVkz/Bu0xhEMzsSFoO
AlBXRMcPq64mUteDfPFlJ95UncmDuyP15Rr+KBCvt4RIees/vIfGZh+5m5FUgd/t
7oa7HgEckDSdweIwGdeSRZGf8HNZ1yZy+kevin2LS2M4P8bwAJBluTxjql5jestU
pvkmf01ee88e0i+M8M61vn2qsMvAHzW7Jag9OOxoCnoceT9c8kiQs9NvS1K3uJ4p
pnVfrogIVa9ZsQpP0/RcWqsMpzuuYkPqDhHpvmrKUY3x1FxEXA2tSpM+uDPEny2m
nk41kZWMYiJdswC0Ir+WEkSZKahRokQQnaQMnPQg5hjLAoOwdywaNNnh27klOkLL
mZghahQhNOqzLe1q4AIc7vqO16arwNQ+J7iZiQTL12Hw4tWVlHYNjNzFYOYjt4Dv
0qNbn6Oorg7s/FNFMDZvOZta2czHibrpMSPx4UmPRTw8yQkN8JWjJtjdiG/yseKL
x8EZfm7NKVMY1+uiF+5Mc3JFbU6vS0KkKuWa1rvPfrMaOT4yta/mxPY84Gb/AwdN
0S7nRdRUz7ps2H20W2gMUN6NXXvmpZHv2EFOiapEmgNc8yxYflYwMAsSedny/1Rh
iR7jEUI2gLRsoyf3UJnD9rge7+dFH6MOJVpfdr4yxCFQ2wepayn9pOnGv1aoZMxX
4h5iF8J71ezKAe7hCEZ0+x4rLC8bNswsOoBulsA1MdlUYKKPbAoUb1KXH238p5rb
suCgcXx+gzX0Rrwz0fGFlRKFMwgxnMuzbel+aDo0rPaVzcG/4eTpgJ166fYfdN3f
1FRDRVV1bEKvIxwaHeyH1e6x3eCDyuDNYl9XfQCuOx5WTBapRB7DE7dYUnh+LnDO
8v2Lps52MzNBhTybMFjI0RMVEaWOyMRSCnvkn7QXx7qQ8vKXVPnkXq6gOWLfy0We
1zlCg5TwQb+9usehHPRcfb05OqnyAJIbEY0nv4Y6viq1Nz1dhZqqX+LJCsqiXvIp
nwb10Jcw5/dZ6rPivD0H9TWdXp28cCp2/xWHzUfgY64eoss9S9i2GAoHcMkmeVOq
Yg3yd+pKNDnDEeA1OM2fpDkHC6wWtEXdeVp4rJR4006orC/Us6mXeXnZCCuVTHxe
Pg9NoRnb5IRvG0WUB4cs5ONC6BttU73yfNgx+M4ePgYi3TgNCuSwK7x0CKe7RIwF
tqYiSVvvSR9P1oXQEG53mI+rQBzWHZT224FPBgulrp161gw7mx0gVuqNiXcxH8Ov
NrTf0WWVUruOKm/N1FbZ4z25Xwid0AhnBjTSFLiIqV/LhbxUoFnL3OE7SrLlVyAs
C4hltj9jr9NxlHR85QEiJg7wJLeXUjqq7cxtn71zFRO1vxjRIj8GE9JdgicxyfD6
WGdmyPD45p34O0EN65FWcxzuNG449o3X4JBtz2eRe1/DOrIciUt/dCVSsDlRM0O/
ANZfkc7fPsUj4cIFIKKTXm2PAEArUWaiQLu9qpSBGow/0bB9R6CUJakKGWzwxWxW
ebllBUIE0EhafaSfedRBNUcqNgjkTXoaL5LUIO0sWqPfYvq2Hnw4rHjINE0//F0G
nqD4YM0BjL7z2S9dqaYdLcoQEow1HLOXmEcPLlt482VkG3d4BEp0B2LOUMBEi6Ab
5fsxtdxH0NXwew5TIjoYxOflpKWX0v8U+lGpYJq4cjy3K+6ws6jl+dXyn9GeogZl
YBxR33lxOI3pMCJUXWo9bmSXkqEsrQJ2LUHoe2ZVcOkVSWeFimImKAq7zVCZiPzb
rDSj+HkWoJxPJOsfmUsyGc+WjCZzmc1D2+Nwb6OdE8C9wOu7irSYDw5dP7AFqKBB
7YSf6WeooNd4rEGrTZgj+i7F7cyQ/ovwGQiQWFUFYXIuR3AFM3uvRF42JC70LBN5
85mm9amLujKRThBubICkKjPLIf+eKGwQ4PJkbRXN3NqQ6KTmlmv5OJw6401gDekh
e86WKogw5o1HJ5hugtNYTOJb33CWVOI5lJLiPU206SJKptR7zFPCyk6h60ANuVYZ
9aDZXg5iy0jGgsPFsc8PkTQmMykRrNjkairhd7eRxrk809ca/i1jeQX5Vlvgz0Sf
47t8y2Zwl/kfiAb7+Tme7D64g0X/RTIQjEP6/4kGEnEJXm7IdUjJFBoNkuwZFwCi
4caCXDySZ+DmWnl/uYPTnX5NmQsh8JyxOR2uMxYI0691TWVD5ca+JLjLV1JMQFB7
91pIu7mpG2t1mzF6D3HCNQpeWJP7Fazf0V+GNlaJOEY+BCZ1cs//P/ZAme1ty3vE
bCFZ1BAMv1wOxLJjQIBDW2ThEeNlirOxnuKNbzgkdIffTU5dfzj2Urb+kN9Q4bMK
GwfYSsUyKTY4NtWPTSbLDfZuRufXOXRkAGemCkH9zDiQICbEYBzXq1HF3gWq1vAx
bzjvQuzH2FWOT9osw3Q6vnHUrEabXB8l6dgnupyj3+1p7K4e9Xoa5G2pbTb1+AX1
pL88kR7UXgDuFddVrRyLdEn3ULMy32rSAiMeRkN6kpgz51kpgrWzX0AVRqv5p8aj
zO0yIbA9Bnz6eQGJ36w4ecMl4vgTE6hvUDbejSgQMg4W4kp7lPMH7Cf80ppHb0mn
K5yxJzSZFlg+7+aSUPEZk7KVUVJGJoxuTlcX46kCLNDPnwiPNtXTv7bdniz3mC+k
V16PWwQyJBRRCoGGYwSWM8/boRDrlFp3bUy09GeO3dOeMo1Cy5GIwW5a+hEwFkIw
pVVIuI+LbS+HjwmUcQ/T9a41IUmvXFVoAbAd13UkB9G3hPfOhfooI2my7Nn/yxT6
YYKlzb9etNt/NNeWBBSZ8nz5YbN9LZxzo5VwfXxUhI7BD5bro31wlyoluTkmtYky
a5SqRlTr5a5HC2Gp09klWzGA7RBVlI5/5bIS6wu7HS3Wz/MAp4UHWGyvf6a2XuWd
ZqeosvERXXiIveh0lu7N72MmfJg3i4FcuO3JEdPWCkidLe/AJIj0FEu9GS3ECSD/
FcRlf1yELG4jjBFnrRdQFIewXV4Hx7fBZGSGgHrkm9LPkpQqGQpEFU2nrAgwXd8y
hnXlKs4+v5zQLx14G3pxHLNHDwADFHUlVuzrhb5Vv4Bo9w3KYsnDFnILsRSge3sX
0jOZ3rtl+YJ7tLr3ohCUAhzxPd89Hm2sD4HRopWq+XuarHl3leHABetCJNd/fR9L
GRx/cF+wrIhljbdtrUs7tUSe5flZ2EZg9WglPHDn8d3fHq4Xe+h7mOFLWglypg8G
8FxL9TCTDEfsQq9fPgxm3RwffcDHQfMWUsuAWhET6fHxHOF1VfXKwTgPdA8gAOyk
oimBqQaYIea/f/LThpfXRJT/d0U3spnx9RBndcyDhLT3VKdqvwozFTY8YRDawj12
Zj8A/DQHZe6PaNM/ofTm9ra14SuPnC1CCDEn1UTT5Lw/wod7gQJq6ZHpHRTXH5v9
KULvmTlJaXm9iSy61dqNGnthAmLPStyNLO6emPIpuDa3Ctn/p7khcVdCMLSCa/8t
4QCm4a/XVe4k19pUG4DllelG/OFZzbSYB5WdOEbI3xrbF1cxRTbpnDhBXjJuEzCa
c1Sxdu0V+Fm3G4/Wew7esYFTO6aotsc+/RVUjHuO9Kd1EV/dipT7jJdmgaXmWRxM
he/PjR4qoSaVWrmxQfKTPdgdSblYRGTY1HgfQMGHb3jUrf67pw1F9G8+U2DHjj7d
+BFzast9tv4a0PDH/OAXT9BYgWmYBw5wNyTwRJcr7UadeWin86gHGDyrgtYcDLd8
HCB4+faY5SE6sxHSDyT11LPxuUji+PoOXkNloJwPLCpooLIkx1z0y5xSUAe2LiXs
ltR3ndNfFhTVRSLzjK5QIJBUYyNQX0MuNEm/shG+1xOYmE2kugeVZD2S6zCiiDDB
Mw+K6KWK+rXEbcg+QVAd2lLO9PpF7Q6DpUtgX1p04AsB1KEWYulQ3SYOgYg2vEY2
Z6HvQsYs7AwGtN8SCfdDcVzo4TZ6Z8HWBVVmBWUx3glgCymEb74SoBchi+xxPqjz
PM4tHpWfRzQ6ebfOHh57vnee79BXeg2/wwDYcbYWHzM7j0VjqgWm0el+2MYodQFY
X6K5YbAtk5REwhVhEh8187HWm2xGCODm0djrNcRY1sUqmYSf6iqBv4VDR2HQ4LHJ
GOVDLCG3cj+TSW6O3dsrMaX8DXh1Y42UMWSlZYoBLldJlZCsrxp+jGd1kacP1pMZ
E5XaTPFPEP2O3tjRU5ehEJxQcONNA4i0aEnAJhcHIjm3I08yAXLkOBHlbidPbBSU
icow7IX8TloDJ4VrVApcPyj0op3+zyylHuk4iPgWEGpLDoWnvs2HBrVlSIksSfgP
gMj/ozIDq+JqbY8okcrWh9P2YJyLmF392jkS2Xf6ZUpHjbWrhL3rnRESv+hVgHET
BISd9yo4tIqwLUUX6BO4NmBzciYugOfF91AzbZrZKJXTnsy/mToopQI8F682Pv5n
avFGzN9PPZbKfdZ7eT2dDKGizlD72lqTZh+1qGnUCzNV/xGMot8UIxWd7DSer0Dz
Cov8wtvrfX8Muz1N7JSd27QmuCzeJ9jTa65x/aOzZRhbmhLN/0oayPH7hWG+0hWe
fs5Z5o944fp1AGtvulbHbsIKDax6F9+Wohtw7dVOrStnGlIJJpLFNBahfNJQaE7H
vGmiPuLr9pcwp7pHbNVMNcGaUMLTPamQYE6uyzkBMYzRmDvLqSs6yBQJNHfsZeAj
djroCBy9LZTMPC8xVRsLT8gt3xjXaJsOG84slDyJZs7aq7ucZlLtdzAxuV+YLGu8
5njUM+yKLO9UkSTjq8wi5Xxfv1FC5cGjEOgKkTewruHvitscYK8N1tPGtRb9FpgX
yK3u/a+x2SUJ1gNzyYrp4OVSWouXldSPXzk9nRlhHq7Kh3PIIMbYQjYbiKuOHv1d
Zq29QrTbwOHwLyxkbCZILiMffORmKaFKN9wxHsbflJJDWMHkdx+snqdeozFKpGat
pcRWkYugjjgD62u/o9nRiIibyRS6reSRPKqxojv3chux04ZWUuS8B+dQMnEiKd5Y
dLgtrtXA3GR/Jwlt6hq4HbXhyJ24Ab3lAPVnS34ZY+H2549HNrQaVh+pIn+1icc+
db1Qf+8oxZBAjhy02ZEqwegMA/mxySGDhFPqCmeUAocerA+lmdoidhqaedKokmgu
HxUH1wkvWwgclpJDNPPRrHvQyYmobVK/NA7gWTyCsySdnXgWWBurqKw5tKsA77MQ
RXSVtz7zCkXk0W9SxM412vzzNUOlLU/01xu0tCNZSI9foM3Lfx40fFYjCBVi/qoz
6wGcIN2oavSnmEeRSCjNgmhO6bUNfkZ8PRQ2kyIWLmVt+FHycxG0fvTxtZhwVMMK
Hsy8fpOIITWbv8XJBe06lIUCTh8oNtPOs2EmGFiYRo4ymtPWUC9SAsf6w8F+mzLw
3D7kR+Z/IujH6p+RFpzvZ/Mogp+UD8nVc00TXs1k3DQZyB5xHfdiVqmtqFq/vxbj
H91TwjVua4UHCnBaGZVdQ6b2XnRXaZVYEb2/v1H6lNfiaQ9WmmLwMsTi5/aPJpj4
+fpW7/xJ1M+BqFpZVurd0fXkF92ljWuBIvUWhUwrY7l+vTadu1ng/i12/hcqbPsg
qj6SxtYo5Ekeg4cRNKMQ7T17gmpFKznrcXLov7g2EyHbTibK1ijzRMm+zPFVqfn4
OzZNEtdGz7wtdaMbY5Xm41cQEdudMyTRWHGntjzTQiF1IAJD4r8MlH97rYtE/y3O
1hIHXxrzLf8lN0GdjYaQ4+IFNG7krp/BclcN88RlBhd6KOUQsKKTW2OBnmh0BiJ7
Zd/BdZZ8P+Hjp29okQ0jAY6AeAScrQSqpeaNOn8SB+VIxaG/ap+ho+dSZYnJiDN8
0y6SmH79fsb1Kh0xgfi7RO5yqy/j07I97tr2Ip8R5/TRqn2RFct83Trd2Rw8H5ju
o73gXbj4jXcinlaOd9bD+Z2+YeVTEHBHFnfWmrB8yXPHiVHiVB/Ai67gjl1vs2BC
m8zGjM2iv74+S7pwdooutbRMqvA1FVQfE/DR3uBNFSY5/Hrta8NUFVfCSLIwBK7/
LHPpMkz+GBVbyRwF/h4YMIK3Q16mIo7lLnDXigLsos33HYyXvKmpt/aMEEmWDTUJ
ctSWTXJ0LGQCWmWo3wg6Wu1Pv7/hEJt+qMQaE5yqlUajHPVaQawaTfH7FUBqpHoT
+P4KnI+Nu1rFa/CrbezwZz34M4dGKut+Dei9D19CToONT/AI0X2eVQe/9iB6WY4K
LI1fsJfI9HhaX95jqROqh/rTe8h31FwrnayO03x9P65pzvzfomJvy2ScTXFdVH41
faTmxHKlCKPuxO9w7iR6r9ZTc5ynWIsD8SSzXkhwqisb7+XH7g+C8tJfJryu2UAA
EhsskKRIb/vCm66pLI64xgMc8qwtqDk3YxSBv82hQ7P4dyztFc7KulZmQTi0HmSy
drVZhu+A5o8VhZ3AFYD8p6kgn/hI7PqBRzkUDEQJ6uCkBIvtYpnsMQo/SxBCokHU
X8vj8UJxLkVLCuCGMKEo6woyZ6m6oOjbWu2nkDx8RJhZR0RjCHRtiPe/akYQs6WU
y54bAsSDoEUZVV6ZmqOgiCYgZPpFMZFTqNfhKYKL5PYEFbIET6V5OcKMh3Sw0FWs
ai7OntfR2HbTP+nmAnHhmdiXZX1Ska29wpM/pSbV43aQA6+m3jvcn2btVVn6sJzM
nDjI2FNONgNNagge/DninK1nleJ5qoFp5a2qsRNRLqYlBajrAfP5ZQHmEt2NHhzc
uRPaPVXdFwKtbOH5ZAKSqLZxyujJI8ogDV5dfuMp+96DGVGlBwAjNor91q3/hRvZ
LnPAUM9Yicjb0T7AKbKPbMBVyibwOAay3ghundomt9d1AsyDtHWXWU3gmyTfrtHL
X57Xb6IFr/8FBJOcOHRp7a4MukM50bHPGB2lFvlIwr3jaiq1eZ16oD6BH/k7ZwSN
30Tq51W+c31oz0kqkDxH4QwcXqyHwZw0E5gik3uiWfiuTNmyt0LwoGwz2aAEPTSc
JL0G50nbGESMV3H/J+hVGjXnf66rGr9TjKJJtIJMIR87QDMgRAywmKJC8LH5uOzP
8l37UzaASTvfH6nIPOVOUZoikvbny6wEwDVpwSuUx2F1bFO7qxFfMsPQcQh/0VyQ
J8JDd+orwnC+3LVG55faii3VDbaM8ElhaQ68t810vUhr2oCfQFo1/zEmBNlrUon2
iPL9IvRa/tFdsQQsFkc/5EJN4vLQ7752U+NYf06zE+ad242XAmBw7HvDIl4zNsSX
0FYkEOABmB3FEh+u3sv1AC7WLuWADCq9e2j/GvuERazzYts7tTsatWT3nTKZxnza
qX61ZHS0R7OXoPtifun8GKEMJ0IsJTlNSnGYPac9K/aiu9R+twElPf1Sg4qu+KLr
kjWh2phyT5wsiASmK85OQuDcKWuLgXdF1B34lfrzi8UgUFuzxlEdV357Kpq2jlnK
zXTtXQk+TL01VjpnhRpRLQl/QHuWO8F2voCRLOpz/hgJm8pH73URgbq3cNSTMi1U
RdghRF3XLISIRSJLeCw8dInnfDU4d2tGcWAeIwjnNRGReZTRYnXifBavDZvferae
ehVbNhfXI0902qpjtfyR1pQV9pZA5b/zTlw3BpMgnn8/K+d1gY6i0YztB2D0KIp0
2EsYQ/f947oQleK9kebwtvunqxgJP/rZVsrH97FtPCCA07K9dLMEoGgJlQjg2HkU
0cMsNUGH1W8R6VBxwX0yZdE90Fg4KIDqsU/bxwfXFSEN61eXq1GEGvkMQcvTsDmc
c6zRFMWz61CMPlSyvTII3GbqQjuJiELTCi+tp1YWvIA3M7MZQqr9BhE+GwIgosnH
rxOtJ7OK3aB742P1rtYjASadq9p6bzvzf0KZQhDQf1l4PraOaZ3Cu1dgDVai5wJj
B4Wl12Ny0OBEmBPiivhIWwjDip+mxNpYnDyIqwHIvuLPWbFKngBz4j0MHKOEDRE+
y/g2+S9hbNenbia6IF3GBH2Ev0Yp12EaxNiL+2bP+BHe/p68g1SeV1YLoMWCZajk
f6K7I7RFtb+24ysIr8wLgZPEpEKpW9qPacwqc3VAkqKiJrmYfqMPdqScDJCE/SBJ
rW/15MbmPEXCB+3xdCIY5T+bsIgYTW7kCdRpoHGRTrKUWfMTjDVFGP/3UfwusdFu
PHVs2Msjfst2ZH9jDL4pWdSABOYjw/u+U13Iwjiol9xFZmKW1XEaa60R+lpW1GcN
P1hJPNVXm3oBIQqr6zcERKyNc2esFQhfkVPYL6+YgZFykNVNolgeppoF6EBduFm+
RqQVeGhejKTbj11LBsTQq+961mJGayfYbeHqr/QMX5XRmHwoSLPHu5gz0P/FcZiQ
1AuV/qXGCMsGfBnScmoKBsR8NEt97BJ0+vJs5+hfQj6SHTaPoUmo0eX6CF9ijuxB
KKt9MOiPhv6Z3sTSrvbUCh6EwhZf/Ol9fwl/mJ86zJCZKjyjpSwNYin5Xv/rUTtz
SnUWaVu+bivnio5DKNH5QtkMy28At4QyAhQ18oQgYiyguT1KrWDI23Zdley/FkzQ
G9OxjgatYchLdJap0k70PQnUvB5BV2SEFUv9hlz1uWef7y4JiP8jG691kmXmTAu5
O4zcrzrRQjeMDUbwKWZ0tvk4LJH8cQJMe3C7WxXDmPGLP5OAFltWPmx78lXgzZs6
ips/y4hLVq1lfScL4Rhxbnbg3Xo6I6r6LKF9jSjsO5f6X4UTKgjHW/BK2ZkZllYy
5RJjE/WdkJyyuHFnllF7A/UqzUCBG2BcWyRzXCUls+r6z2O83ieV6zeiRP37nyKx
g1fe+hP1yUSW8RMFXU9w0WhphvSMxhFKRGLwgXM2ky56CcA+fYZcxeKWNhI+K/BF
/R/kJ8l+Zl0svtteHmkCNFnt8FrhojOKuhaR0U7/0ak1wtlo8iyAuV3XYi/bgPrO
kkYng/2qnZprq3lmBJnAjpm5ZB9MMVtLYmg6GNqeXiHGg8bngwXmKxIE2LHx+mz7
inp7DAitnuTVIpnhlYZmYAWuyYgIK+6eWqtFvU9hMyvOACOFmawTBmPwJcC6mHZq
OVWjRB2Xe91LsHeEQIj2L+ZTUiSOpa2fsLGR7lKwufQYtUNy3/KG+HzbP2+wSljX
9aZsLTb8ABP0H7uGWaEKE5WWNxSFs1a5BUfxkuxnC+M52YAJp6hpsxawvZY7Kg5E
vKoORUmTZMMkndJaeVZqp/EC/V4s3bk7fzoixhP+hQ5vPh4bMf6T3uMOtQ7Dmsr+
IVawIq9+DH2OGFR/GnfTTCz/YwetOqG9mSYx19ZaThWqnRRevHb6tnHoaoqFq9XC
yzNcU+HJGV8vsX/w6hQnIqTcnMLFV0RYqdmITrmWak7GP3Mf2lxJevL2hZM3qaja
x4BFNMYJ+oqk+Xlx68jwqG06nxbTYqQiACW2CwsKsiAu1xDgqOht3UqJ4n6Icmc5
Kdy25+7YqI02XjSsVWjBUN4H8MN8p5LNzNq6YKw8gwmv3rurOv6w9kd60T73weqt
RmsoyZGzbq3ecs9ATLgeTuCArj3DMVqaOUt8UYI7y2jIajM6IOpAF7iKuUYUnXsj
Mspq6vJB3/WzqXNeSpkyBTSR0BTA0pBZjPnW1T13aRTxTih5BXLb7E68TybAzsTl
ZkvKuLBFpNaiagyh367U0tdanpgqVmLSzz0wfvczBy6q0Fj1Dbk3Iamfztj4eGL+
IXBjAOIi3YPI+wn9StWor28FJEofXqOEL5W27AxA0fQko0Hl5COxWp90B2lxXLhp
9r/5EOCfuMnQzyWMVfcySMjcy1ICObNJB9+3g9XsrkswRxH6n6WxPOjlou1QLaOX
7RuwLPn7C2DByudHAaHjkW7eqGruCMUMQ4XPGktLt9H8iDIss6j0nclT+2vWfBjS
+AhQUdgmsmts8SCM0UVgvLT4sN1M0r/Jr/DkDDVS2BAq37B6thC2I2AoZjf3cjmG
zBZ1Yr8WT5RejYSl8M+fgqxgc6Z4wneuZhjbSOq44yIPUP+LvpRRc7HsGO3KdCED
mbszSiTT83MP/OsDAnALCpoHh4gYDOw443KkCPjqIoCG78Y5DtAY6pWg90f8nC/Y
TlPUu97Acaw07TvN8YIQlRmPxHObSmRkNjEuz9ZVUqz/alHYGjH5uRzSOKzLi04O
rn+Jl7ATLtcRIkrPje9JoqAlQ4Wo3D6yOH+xH2TEy7rb6Np3jjX0FZECR/DJpdYP
kfVPVq+7Ozxq4wL966ur6eWlMMZoiQIwdiuQ2bIzRcCEFOvOk7vySWv1Gko///eX
tVR4lDRkJ3zFM6JRcSQeikiYRZzmL0y34+Me1hRKg988s47VhyqxEffK/jwMr0Dh
yt9RSHPRgY5wq2O6d8sCFP75dlKx4+0pwqlYILNz8fghOFxiIlAvx/tbIFHJSU48
xVV4+zyAy1YUaZKM8bm+fsmDu4KvUZmMnKPhH6zkEV1teCkeiSvrXaDhQvDJK/2M
S0baaU1YY+fsqC+ydtgFKzD43Geg6zV8/3iomiUQry0WTE+C2VQ6xkc0XXd6PY7w
tRxFMe1j+srO2zX63JnYJV91kwQyJRWt8e2bR73DAmWVUoRzdRVPWTBlDviZnBZN
7EDDSu4hMCp6NcssmpD3j4TgSOtkuGugHnSGijCQNtmGN0pp9ws7QfJgRFAnG0gc
lvqFhh+znxJNs1MmiVsde8MtsjUK5zETgBexeVd/+a1QmlagQM6ZqYwwLCKkGi7Y
NnEnEkd4Rq2xb+921FWGvElfqntQjLFK/yoWf1OlQSXJVwEJGh9EP6gB8nOkTA7r
ugxNiiACQXkIG2YJY+14BEjCGIDShdcm6DIASqMnOkMX16V6QceuOWneC4PHc914
nA41616cEpeQKRcnVeU/g2ZopS6BrtmDRc0jZm0HktaNprMOSohrCp5elzBYYazz
lUJwAZ0iHwnjjz46wzVRlKliNgyLWjCP+jzUQG8+hpojqb0fwMzuCPCgdExl0B15
JlvrhfSe6GO/A296tthYfnFYI8YX8oMopKzeKmEh2Brg5oLxWFKBQ/cJomr5MIdh
4lMRxvol2PLEDopTnCcgAzPE0FicH/LcECxdIsKGIDY701nBwfTLO8XYdCXEJdqN
oBsGRd7ni3zRNQB4fBo1jIZf5HtAaDZV0MvAA2GTDiBEVQvUPDC1dUp3mdPQelM1
ob1mEC2B7mNoSQEWd/1i2ESwrXVW8wjPjVtlCc3s+DYwbDeF5FRVSOWC1nTo9yP6
QmanrCg8zJImJpdl7AJs/n4LOZqoiOZ4HEmDME9kSLDyj8PIKss/VSeee9jXVBjP
KpK/GWAG4nqsDgf8+5ARmKY7TvsAIMuU+X+Z9D5d+TV2zqd5HrlwZ8w8UbV4YYjb
x4XNtmTab66uDxO9nJvoktcBjDvJP1Orbkc5x18vj3A0lmebPMRLWc4i+mT5w4vg
8/FuydZFhQujQU8iJPImo1Vr2kc/TqTNNAalHyOCKkVOSBw4854poGbrHj36FFNA
0nPtKmWJplB0D5Oqc6LNubkmdAq1eTAgQLiVJiL6DizlFaZUFDXd0/oTLUjsanQw
yUkycWlZ80gyFsvkBqAyi9VJSor4vjVlnzlkLnYx3ZkDQbq9Ju9TVD/8CYFVu4VN
SkL+tHP4YXZVz5KwyC4pRjN/hprUN+qYs+/+UPOBXPmuSmmWtX6yMbOzFBQF5xvM
hcaz7hUIHwsyri51N7MlGUDcz+9FqDjJxzgoHnSlcSyJj4ROygugltc7dBdVL/qs
EQ972iEWNWYDlpKlRNWjDaLcJj6WTf2wx5YZPsASQq0M/Gr8syz2KaZRVK2p5Ykx
TWjV15eiS2hSaZbQA9GSfpePVhefnqGAm0xrNJ/1pVSlQ18ADj+UGt2Mxw44zxy8
odbFcjGe512yIvrxLa2GjVgq661vvo3Xq2xsfwlVsAmnHn77Flp/Aa6FXRzJOMbc
8lzUh5oownz5Hd6P9u0PUz7Y7d3btqRMxGTiVK/H/BWtMganC/ETWxbvc4l9p8RL
MDwYYNil+oVKrV2RA6hLMuEyItNsUkon5QV+axs4BBXhPFvgdzjH7sdDyaHrOA3C
5wr9/W4Esq/g5Ww/9il9xIXTv2Irx3+uOjYY8JfY2XEfpE8awfp7uDDO8UtSfPs3
7hHpCcvcjpBrd8ZnOx0+5lWQkzxgL0x7B4sIo7yy0ipCFKhSKRX9/6YwiDRswItd
fOCreh37wM5r16hZvoBTOPZMLON1Z4VK5NxlHNV8SJXumiBkJSlKk7Yup+a8V7va
kpOCRcuylr1rgwQuu2y06O1wCKAY1LkhNOqmHZt8e6+7sD8uvB8YJgUSV5CwteFK
ATMDPNxpHVCQ5eshWjGsrWLXXEFP8koyitdm1zc7Nx/l9ZQ9vz2Ey65TQOTEvg9K
7FV3rt2c4E9vBk9pCV7cJWFezBNLz5j2LhioPfAt6ZrDaQ8uz///HZBPdvO9IX6S
ZUxNvNVOCmlg+qe3wvhhykr+eii+IyYkIJ6GPHFUng3zSP8wMTSfut48eJTYxU7r
B25Q9CfLfIdr+yNwROgfp7/m/qv/5EVPFIM4OIU88ByahppBoFRWslRGnn5ze3x6
oO2jrcm6T3ITiM6YBW8G+W/43lWAJckgqkFOsn/PHk8kZyxG4W77wfbDzav4CPSQ
a7X57r5dtHQ0r4vcAlI6nM7OFEOmdOKZ10+8/FFKzVC2i6ywIAltkowsjtmwVz2L
omE6zZOoGtYPNZgQvOy5/CVqoCWJzI+Jk8IU/NRU1sxidPhTJw8M7T/VqjTsWbOO
PcLjX1kF7pyNZALT5/Y0kTwAZE1jvwn/83Mm3tGVSy1za4N865CGVhcuPvFWK6hf
PNvocIhV78WGd3dYnIqaYJiyHqEIa5DwTJhVomXKHBL1sE8bycn6cFY3j4uqBzXD
KaSlpv6DGCYhukKgJWskPe1UNx4GKDo8Ie+jfTXOSS83D5m6l6Xuh283eazvWxEU
O7hrbkupAGbPu5a5EhUxnK+XkvwD89v0+ahC/Oc3hslyvaKmrhEb8YQLtcEeSURo
l8b6R1PD++3X2/p07VerQhJWRJJuNiz6GDymvCqC327lHO3bn7OCL5mAHvLDJdV7
uNpZwYTXv0hwN5wIZW3uEVvhYfle1VZbvicsNAJgyMbWO2Lh66xiyoHdKbRmBBh8
1LaQW2qlejYZNw74hlM75hWagiAv8+PA5VCnkJlY6TSY3k83jxLXeh3akTJfSifq
/p3ticainTXyhWWWU25vTw8TFI2b+/5kABl4cPmDiPavXmnwMqFA5wnVpX0yjEu7
G6wMYtS9LGYX1a0SUwVL3zafEixGJ3eoJ4tUkNp3di23RlevrtDNHeGC3sNa8RIp
rLmh6TnXziTEBZcOuStt9lzKqhVcyZHePQ/+hdAYilkBhXxz80uDoXVOYS2g829l
Z4hFwRExv/inXiiSZC4swAwJHVEoa5q8843y9R1rF0+PRV1VzKNCfNGJtANatu/d
54++rtAzumaB6ytgI86OnTldu6hhvW3ocvgM5ySGjlzQCtjO1+0jNwu39ddCI8rC
4Y8C5zUQ13i7G5WkBOHeiixEvMd2B49fpFgFlTW9QZgO2BaU4pyAE/QSSoDrPWvp
jgWg31N7vP2C0uLoYKoCXevZILak36uizYhlN2AFZZ1CDOw6QCMmXsZXAgdAvMMA
EnjDACBYDYgr9R94K5+kdMmTOHIB6zMoCMS0SYz9huFrpD/2d0XIvsHm19egf3SL
DBDcYwtdP9JQNELv+5t1PvNnasPs6UnBHLHBkUnnwCp9xQqqRwyHYlFtOYkW+1e6
iBlAm71hIO4UXAdIx5Lhja7iUSVOgoVG7wLWndrR0L8NnpXYKv6meKsk4wXdjqA3
n8TRmPrJvtniaD68kbV5rSWLi5RI5llDPU9Qhxi2WplKetsI5e7I8ew1lNqtrhH6
h18XQNui5DInAzErv/60LSnwg/hVXxfeu7Lb6rw5fhVP5kLvRk13cXNsoqdsmbeh
Yk59JrG8hadgQYNxq6YFmQBadh2cYj2xkSCoRZYb/OOnXtS5l/+pKXZG+ntrG9qj
NDNJ2aB74dT/K9cyy+MfIf5pkFaBsDulRohEffkNAwqwXFXJI005BMcDmm8ByfTE
zQvnZH6TdaC2rI5PrnqhucE1bvJDkgpLTDEJce1WQr2UdFsqCDC40DPMEb2ZFDOR
PvANCVgdRZPfqLFaKe/pxofo/8gh6D1HIaIx8CueVvF19ULUe2O/vslDmIlgib9b
u3Z7JP8/5yRvmRgahlGWrpi6GnuBamD6o+8x7e5xOIyXEAWE6se7aXxruys92FQP
tr7j1DAMO0YAax4PFsOsWOB3+UGxnCS0inT8SRHoYrjKG5OW0Gfuh7Ck9t2WiZbU
HLRZQSDJesqS+2poonEQtTMiO5QW6Fq5+di9aqqG2ZklSoZCUmABTdrNKOMIZA4e
mEU1fsTuJwcdGJIDVgXgMy3Veso2fZ1wuXPnoHy87C7SF48NXuMTOZaXJtOGzCZG
JyqPuMINsiX53bu1Ftsbcj8+9OsTUNIE4ahrQ1xw4SCeVITO4b0v3Q8SKwTqGBJ3
/WAdyMUUOWxv/3n+KGWFAgAqiiQzDAqqqZIkdKbd3/rW8TLgSweMbS5RCvZa1YX1
Og+0bLGj0shIANiMKIPcAi2hMGOeSHiNbdWiIBlIilUBmMyfVWnFia/agQfvrWLM
aT0D/wTB3ETFpkyxaKUnMBb3KcaeVK0sQ/cP92/bFC4qWcFk+OwChJ1LKMbRyl+q
+jXQ7Kz6Fd/5y+r4+SznWGAs74b6WdRkKkBl+0zHbDLKm7kbyvmqAos55R7EW6ck
XTXNlKNjS0fxyaJ6rSAmSYPYtMZaV8YwZ8C0IuctlEL9Mcx/6bmGVQZ947IhE8ts
vUVpJY2PPLfQjH/vkL6rRiEsl8a8AOKq8ADBxBNIW7xIzijK9ZmaCpWcWXdJcz52
DjfweRRuSyMtxWOaYJ75LYR+HuqimcPAOhtLHTyT/LHeiD0Ltdt7D0aWEHkQyufs
R9GhCU81dgtLe9MIbXIlz5VnXb3whniru+zPCGsMwdqvaz+w4XAy+/mDDjXACpDF
G6zmU802StwEy9Wek0XSTDEQWu8IT10bS1ijJ82Ky5w5G1hJHBaXEXaUqKdwD6kz
UTW4Re1+IbcwXx3/obfUNqlQ0fso8pKLds3hJa3vOpguriOBbiklO2mZwwGQc/7q
dcOWar2KGPA9zOSyNv7feodYAphJG4dMYuT5ptHBjpe2zPDHn80nFCIZDRqjALgg
cb7BGtx9Qs+WoJcYXv+BBv44rzLwazUllo7F21mZb8sSfF2ao0tu1Fd7Tu6GuIux
gIEusVZWcoFTpvYYgrQ3iXr926HMC4uzkT96LjbhE0G+a8IN2HXTAV6T7sMXaLdU
qsMe+a+lvPWovaxUNubQDfgEU5DA6G7451IkPrwcYeBvmDqKX1F04cegVNQaOrlI
px2RYZMM13k7an6o+BtDDF0ccwOsfNMnWkmdpbsyf2W9nNsqi72V9Gkd2fUlXowp
Z6Tp4/IdSI8kRfi+xhFUOFyyyJfDqbxhfIx6jZXqkoUDakdVmRwP6ISRKBK7HJaD
1yP/udSklLdRipl8AhDOigKtnVAZQNnghT6rbuwY6QEByfKWIoGo5Z24IA0n49za
pew2in1LN2PuMHV0qPktiZ64xESAtTgOnho/VCIhO4TIbvPoE21ZlG6i2np/Krv8
OcjFF9NyWN3XwcOekYKCQULu3xULF+o061obNrE4CfT7Ci02vvkKZB2MGhOaQa+L
V99yHV6i2spF1Em6a7idyUHcYRM5y1sQNa8S+dMwTZg6asdNYOGmubzStStG56HL
z2lQiNN1YM6BK36g1WyBaTw/3lu4OYY63NYPPEpsidrgUYI/fSWzDeOaz5VkL0f0
vZTWz5TEryIVR6Z3dyQwmi7vcPIk3HTwh35y9VTbYVVBHZCqyNM6r4zLsswvUz02
wRTDf7D8XhAqCOhfCDNH+joBa03uQy/FWlBK9VIHI0KpW5MMKD3g80xH4hA+HNQ/
ff8zNetFTkLjCwHqdb7u4L1BvOiv/RirNXR5nG10IPkJ1h+kZAPuYvLvWAH1TVRH
gWl7vyIX9ES9tmRioSiwYfMm53LXHjYA6mAij3nFS/zMjjpNOg8nSY26yUtVeGzb
WQtQL1Z7+KWhAx3lnRWBDfJ3vWW9jc38f4Pa97uNNx6tcZ6eelqsi79Kv+Gru6ed
fqUj54+mVnajqk4zEh4lPLS1akeY3w5yuvFbn38g5BupRR5T592VYgTnGAoRj4cz
KTKJTU1d2grpohD7ThZN/kAty65nFl7fmG+dGWbRaeVxcIZzYK7KwSwlYEAi5BKM
97dFxYYtoFAnGiALJMOW8mi9m2bET6c8Hf2wjug9n+AXTtIp6yvMEDfUE7JrXzSX
lDXs12fmskzhOWVlDnsVq1Vyn78Cdle/A8OjP+ncCI1KkWROoTnq1Jp0HSjM3Pey
+3f3RxjQMzm2455dsfKiuskvonoEEZT8M6xE0gLfkUhKiPiGeBu+dJVNqQlTz3Or
6iln1k/o8/DbFq24q5EVZz080XCMIEsx9tf7D0DVYQI9n7852yZJcmgI48w/dA4n
jBRj5N6C//IUuoHWg72H8+85LHwuGzMmiMQwnSZ4mJZNRixd225pxYrhD3F4nm0L
tkH7F3o53KDgr1zHhSJtKge1+jIFiCt6edhjuxEenhoGomWA4Dnw4uKjE++/cNTT
DKf2WP9fth13u7cNMgyuTQ4ghsdm2i04RxMpz1m5QFw=
`pragma protect end_protected
