��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���Ⓞ,B�$t�{����c�,�-��� k�4�	��[%��B�?���4��\�@e-��� ���u����'᣸߬Hӣmy� q�`L�S�L��-|�,���Ξ�<j�����̨O��f��U�,ﭵ�h���voҭOu���[�)n�g*k�<l��p�l�O
��䂍F3v�N�X4�p�j�7���6�x�$$9�s�=����8I���;Oz�^	.�r"�ɮ��;о8G��Cu��ǑN��������灟48�fڭj���B��n��g]�U��lr�R�d|6a݌o�J-�;JWˢ�5a��Y�M<�.H���Ͱ���z��i���dRI~��PZ���Y���RS9�z�Bx��c���C�N��&=�4�^�f�aaY^�!=���}6b�&�q���{g������ {������b��Ӑп%k�@e�&�;�OMZե&�u؛[۞�R<�#��Z2e�]!Y��A~UX���F�������r�0�Jl�
���n(��$���/�Q�+{3
*O�����8�(�[��wk��v�����a�G��_� �x ���'Ty��T��D�3~�7Ӓh�ݻq�~ʍ��-�Ozb]g�~��i={�`�=����?���W�~�jH�l���&�ƶ��z�*=�v�������24fejn�NŜ�5r��-/���m�
D��v�Eǉ2ĭ�.�܀�Z��,���"����į�>��E��f�ڹ�M4��*雓�<����A{�v ��V��~ggyOER5G-�B���.��83�&K��X8��uC��L&��3{r�d#-֨��a&s��B"��O1���}B�f��
�q�w3�=��~&a�S�F��=�U�������Ř�̘���Q |oэh�9��D `��P��n��̦>��~E)��h.q���̚A��ex��Qθ0r��J�B8e	�#ݷ��������)9Z�$ϴ��M���3y�1��������CF�_Kg�&��z<���1�3�H�/���R��S��ڡ�e�:vz���B�S��-"�KM����ͦ�o2b�����	�f�	�p��*/�<��og=Zs��*�T���$�U���+��@�[Qg�$'����Ą�j�-�y9st�j�R\�L��e߅7睅��Ԩ�Z��{��4��_��"8���*o�ذ���/�a��}p ����慪��y�	:�E2N.����n��մ�{����;��9���}M6x��]&8����<��\&PCyի ��Q�2�S⧘_��P�T�9t\Ȓ[��e��i
���Q��!a�Y�iSm	���?��*x�m7��뭷B�D��튮J��ճQ�uT��������֟���o���+��Xs�A��K�V�kS��)#l�vф�1�Z�J�E��������_E8����e���ɂ�
�w�|��I����^P�2�����} �����:���h1�k�.�$�P����~��\mgٷ&FM�}�J������{)[y��`�,F(8T3|��c�43U+�3�� h��i�$�T #���)�^.a��ن�J�-Z�2
2i�{��ZHAc���_{k '0nj��u��R~��8�˥iTA�ɇC����6�+��o��5@~�=�A�i���[c(�֕�3�I�b���
r����� HE�H���j��Ĉw�hg��^���K�0��|��r��%���1ח�Լ������@��Co��,��_��}{������37}�f���w�e>�y�'�S�}�;���K�[d�9��9T�����a.�dL_O�'���)hh8I��ah�YR�{�;�j&%!���rs��C�uä��ĆXk�ꃦ�G��e�,1��"��d�n�,J��o�Y��,�2���?�t'�f�-|�7��i1
Ol2a�E�'q�eMΏ�N_�>\�ݧ%.������S��=�G�x�����
yTKR�K10���o#�!�w=��0�p����H����Yҙ��߂����-�P�!L�1�O'�J�#��:��Kɫ�o΍�?��u��Uہ�9��
��Sij����� ��d��z�X-���I��AV�lh�(=��Z�Na�U�����
w��p?n t��˧#�,A?²=Kgí�sbc����j�A+�5����N�6�w��G7�#Cx�*C�1�F�՜J�לH��Ɲ���/�_!ڮ�i���נ�'��Þ긎�q�$���̌fQ>�~ԟ~IU�e�Y��/ M�x����4���7��+@B��ߚ"���P��Q��(��=�q��'��[� �����y��|���8.&�(_���Q�bi�F����$&(|�h��"��rQ���t�0��,Ic����U!����*Ju[�w�H*�ڧW�o��n���i�W��(��i�3Q蝠f-ᵹ�x���9h2��T���p���X�2���A�����4zآ��[MO/��i]5�i�Z��c�ٔN�۬�	�#��t��c\�/i����#�!&��fa�֞Ų�o�j��'0� \����?�F��\�����z�5�4S����_����q)�{#V��0.��*�J�*�9s���L9IA<�;�}__,��)��3�4�=
�q�M85�o��h���bf�5G4'�����xZ�S��P\(2�pR>hGO��P�[���ho��ݧ?����y��N��П~�9m%çJQĆ�0��[eӁ���m��,
��+q)��qdEw@���C�����+!"5
	+-���p�$ N�t�<H<�n֗�mX�O˶���*���`���D�*BA�w�)x@�r.�ƑC\�d��1��ѐ��0�3�J�̆�*㽓7��E��kTnlށĜ���c	�E��]p���b�������Y����$����.h,M�T���=BJ�<���z��1�|�o??�C��l~���>������mX��H�Z���\٘����A���8$x�w=�z֘��lR�/K�+h�FeAW���� ��02�u]��>g���RXt��ݨ�S��e7�[���h؀��2ZJ��l,P��9�<ӫ&s�l<��|��D�J��l�QmMb�|���~:��w�,/b&��vAn7P�����F��qi5+5�L?G�/D�
:V)�DD��%�E��5�Wǘ�H�|� �����J3
�� `{9/��EZ�,�U�|AS�U	Bk���2��RY;ւJ��n���p���Y��]�L�GVz{"��P���t*s��N]�R�"X��,�����̋�*Ь��b�cE8�f�B��n-M��3В��x�;ww԰�Z�T�����F9�Hl�� �������HH- _�Ԇ�/�ˠ��ux� qˌ��,�e����]�<��l��e�~AR$�pN� U�b�p,x��5C-R���u�����tsqR��&��u[�s�w�tRP�X��:�L���N���ݳ�ϐޕd>��Q���&�v�S�d��}�*���Gp�C��6�U��h�dI{ȻC��q��[�Ǚ��ǡ	�_�:L��bN+�c�UP�S����M'�,�^ߖ��\�u��ᙙ�\w���lZ ���~]�~��`�HD��k8��.�O<r�5�����w'����'�.�	�&��~����:w+��#{��J# �\�p1Do\�7��;/�Z��\��L�o+I�]~�K��rh�u�N�p�s#!v�R*ȱ�`�\y�J��|�"�r�މ��S���A��;��O�oN{�U'�����'�fG|�����°Ύc��&���&�p�`���׮�8��;K�;'�6Z4�:�P ᦑ.PZ@�Gd����Ϩ6��gƟ0�y�*����+35�XyV�gcU�>��廤EY���:�^^��S�4鋥d��� (� :����� ��v{Fp	�Mnr36�ǅ�C*�����^�.\#&	��/ ��A�JT��GQ敏��ա��&'��d�D	'�}��^dypRC�a-̼9w���@-�H{*r��Q�3��y�R�J>��ť�{��]ͨ)�Q�8p�N
�_�{@q��Ɠw&��fl�\3�o�-�X��
�wz�%e2ɟ��%@arm�Zbl���R�H$���[0
���RR���b�%4	AH�f~���@o��o�˫aKJAvKs�4f�I�?��>�"�,y�`���O��eəB/�o�J�p�f�Qx�bVH�'�R%=G�c6�?����s5a?��~R�d>m�0N-5���XC	�X/�E�?{-=���.$bD�kr��szէ���g�1��#��b�����"}�Mh�Noz����=cĆ(6��Yi�)�����~0�]�>1�f�F�%�eJ�f��4;>ټv� �_���y�g�7�`��QЇ�VK��>s}Q J��p��wJ(^����هR-L��:˔� n��?�� "4������qJj��'t���&��@�ŋ��4a�Y̺V&zvFZ��-��E�.�Ą��bk���L�!=Um��S9��Z߆��j��~p��+9����AkWl!�����w�5�$�9ݱ�.4y���+<\�A�"�An��N��Qj�Q���,���=#���@�~Wc��Γ�h�Ɂ�mH8����Ԡ���M�eH�c���޽s�PVN�Q�ٶ�F5T݉������_�Aam��wv����)徵� g�m���d+�+m�6-C�񙉌h�W������h�
�r�v�8��K�=n��]n�w2s��C�OR��bH��n�f6F45���D�,�ReU�DL�ۇG�xXI�U�e*�&��A ?c�U�ZԸt����:�$	}��Q�NMM�;��NR�w��t-zk��2��4�VNр<��#�#�T���y[�m��@�³�s%e�Y���gVDFXr�a�qs�C�Za������-�L�ܥ�+�e��W��W����Fe\=�����\�t��"�0�Kcy�2�4߹x�(��~"��X[w����ݛ�Dtn�<NG������TN�V2o�j	vۃ��B�ea`�본�=$���`�%���� �5�-��7������^5$s�V���Yg����s+�S+?NA11_U�B����T��-���e�<Zx�N�Hgh�D. '�K���gA1a�u+��H�#��ߺ�j��?M2|N�j׎;n���z�pO%�M�d���S�?�����]��s�=�+���fQ�NQh�U*p�Gl}n	��o3�y��uclR "���8w�?ho��b}4���f�(L��)3��EU
kzc>x���ӎ��|��a{��E(�I䃔���Q��jTa2���x�H� �@/���t��4Uv-�Ƨr�ߘ�	�G�h�tk����oK��} b�_O�KQ�z��l���P��ߧ��J����3^�1W��!�~J�,��9��ڶ2D�����3�&��MxU����ϙ�h0��c��!��â��@��Ԍ�;^�� N��ȳ�쥲���?�:��4�;����T
훪�����˶M�*<:N\�&ͨ�x��������$+�D~�P��0b ���뙉��#�� ��Ê�tf���_����p�^Ww���� �zD�DbT�1��#� �ce���ʵ8���d:7�R�ï�ר2�Yp�N
�P� 9D�OlV�4����QDBwr]Xo[|i���I^��iW�@���	Ý��'~`�*�ݣו{�~�X�ꨬ������CCGj��E��)|�'e.��&����0J-ԝ����?���$��%C�*)i� P������C�:��T�.oZG>O��ځ8��S8��7����O�_�l��i�Xg}u<�b9�1*L�L���)~�=4��[���,���i�t+0�Y��u��=���\|�
+Jr�"؟�k�D�2EF��I��������7j��r�Cl���� CX)�>��_p,���*���/�#��q�>kz��p�8U��y��2�E����͟�W`�(Фj�\���8)�
�>��I�l����Z<z֩;@Rʚ�@mJU��*��ha�2R(1��6ֽj��]ŇPj���(��	b����=Z�*�z��#����ST��1���z��~�=����=������o�Q���?HC�hu$I�ω���M[�lr8{V#	~AME�fQ��E
��A�R4��.��7J����
�$�*O|�����p_@��(Ӗ�*g�N�P�DVy���vvӄ(��gq��r�B���
CY׃�wp�؝�8I��d9P�ߙk���>L�A�d&*X�����Qx�����_W�aW�p���U��yn��0Ճ���q�P} gb�tX�Ƥ��=[��~��c%���m�)�~.k,끢��7�5�hnD�$'�8��6'�T��9���W���(�ס��5��Jw�x+�<d[�G�����RV��ދ���"�'�$�xEu��^��T�����:�1����;rH֡I!�f�e�AΎ�������{�q_��&��\�z{����#L���"��G�)M4��{�d?�� k|���<���švN
ѵ���&/�a�N4�T���Tw�y�� ք���܊@ڕ��n_���p��^W��O���i�J��q[|PU��!1�o�Vx%�IJ�۟#c�D����"X�xNШ1��c�EĮ��._�T��U�b7�o�K��}p��愰N�N�Y��JN./1����'m�ӷ��x��^k�q"��e�_h���CQ���n�Fri�sn���Nj����,I,� 1X4ľ˟��b�b�D~q#HJ�,���?9�ݐB,<�K�{B�%���j�5��"޻%�W�/� cMN� v%�
y�-�7���#��ƍ��d����4���[&?l��̉�.�UKp����aR�Y�@��p�܉�9s�ޜ:%��!��K��=���#�&�d\�\��^���ǀL"1N|>W�זf�w���N(L��{��j��������9�CB�,E�FwO�I��uҸ|at[R��1c�!�h��fe&���%���Y��y-��״-$�	#tþ�����YPp�b��8 2d�5�ԓ ��-��A���jX�11�|D�5�_~���e���v�o����|\*���0��Y<3� �ۿ����\�e3UȒ�Z'z���Lg�,��N5�g��8�U4��R�֗0���.
�=�5"��:-�s�Ɓ&�����0�<b��fY���kÞL;�1t�y��|r��*��#�[+'l[Oo�w1����#��\��ȨY�~@B��Q�X�)�^�,��8n)��q�L43�I e (/6�\�H~�����Z\��Ӆ�p�?`�`�0皛�Thl�.ڍ�IF�,V~��;��F}�*�L���~�>2q�A�7�����7���[��I�.�a�a��{W�����P�6#M*��̞%8��!�k�H�nR��-*:D	(��\\��2G���T���Q�2�b'��qkp1e�R��ó��s�	r�j�^�Mb�&]���;S����r���E"��j>q��FV�]:?��[C L-�ݲ�^	<O>����6����L��^`V���_��'��j�[�Vg�?�ɩ���TKᧈ��tK��#͸��</��W��`��}9��`��&�u��k#�-*��YE�u���No7��i��㕒I��:W��!Dk��]��m=��ߛ-Z&$��N>m5����N���y�|O8l9�'�z�D���n���;��
��o��'z�:��Zku�/N{���	td�j�ç��V�*���1�9��iR�D�?��NL6�v-?�Sc�������ໍ���p��@F�KvT�-�\�,�ѷ�ZZ���-��!����g�(�=3=��g���/��:umˉ^��,�{��{�ʹI7�-�og�:/��� ��J�qm}mt�IZ;�r�ꪸo�Ḏ��=l��I<5[�,��*p�԰�I<���&]3��$`SY�}��X�*��v�)��ػ�'�d��ڨ���+w��kM1��O$�M�0P���Bu��V� c	�i�?Hg�_Y�w��L^B�U��� �E�U��"���Kfdx�gRy$�t��A��ޯ�u�녊��eCT�@��FN���	�a�3�)�/ڣ�}��ly�XH@�x�Y�r}�hxҝ�n`�s�ʍ��!�o{�k��BD�ɂ���h>k��� ^� ������6l��ᅺ۲���F��i6f���A?�Z+!��}� �4a��m_�(�$�g�ƭ2���4�==�e�^蘽[�T{�t���j���PL|: � �� �,��G�"(1��&*�a����iG���Id	.�9s�s4)��z6��z��Ag����{�����v�"����K|����DW��40��Ӯl� p�h數��q7�v����x�O��ߤl�۽U{�t_�𕏶AH�[^�Q���"��bEҔ�jPK�8N�6O�8<Mt�B4�q�0d"�w�-Uiu�䦚����Ҋ��;�ru{�}2��,�.�T�&��^CYY�V�g5ޟ#"]��ό{��A6����n�q�DT��2ʤy"ʓ;8ۨ�'� ��*բd�5Iq��Ԭ]�$�N���u|�i����~���V�Ħ*���Y���I$�F�E���vH_��L誛>�cx�,�@�,�.�U�^�;?F�J:ڻ���]�x7K�\*�;Uᄁ���Ơ\H�'����)4���4(�.�l���_�a'���Qhq��@-.��ԧBni�q&b�oP���V��r�
v��h�Ic����R\�%�W���ym�, ���ߴJ�ƀ��pǽ�h�r� ��q}��;�cs����׏7�Y�Q��5bb����&B$X�)1��.�!XL�s.��)�״£��fr-eǐ!8�o�\C%�#v�G�}��WI8�����s�����`<؋�r��d�A�Qk�^��JzE	��#c� a�M���p��E����%,����h �K\=+$�Z���8� g*��l��w��Fe X��f���\�����9��w;�|��k���1mv9���K�}U�����p۾[<u|�x�rk�~Py�����42_6819.�U��̾�j�~=��HuwcO�GH>*%#��	����/�̹���\�mB��E9w1���1Vs�DT��h��v���ׂp_��*f���8��q!C����O��Ư��lb�f3-���Ux�{�u�-�� ��>�-9��e(��/�Q����/_E�)(i�un��d��'��[n�v�Z�I!��M�`L},��u{i���i~�N_Jg�H���v��W�Hs�馨�E�i�H_ƾ�[a-`](�$*��k�3},�fY)��ޞ�H�uKq��Y���N�N�
z��҅�F�c1ئ�bh-H�|pd�5��/�R����'c���d]�l��B�7~MR��cP�b�:�m|�1'��G�+t�H���暪_�h{D��^�����z�c|+��aݳ�>+��oF�(7Kʉ<.x��s�^�{U���ߺ� �F~L.���x#�̓Q�����5�E�9~<-6;����r�z2T�ϰ�
���}}}QRV�j[���A�:�8Fn���!dE�E�`�=��A� <�Q{�A� ���=4:A���y�� ��*նf���A��j�MA��}7T���(�2]���?8:py�S)�1��0�葡gq�R�G�b��ۦ2��z1��T��:��������}@�u�=�=�����h^U���;̔O����n0k)�%x$�s�E�rf�� 8zɫ#�o|�����Syl��Xb�S�Aj"!����/�����R�q�>$�FҲGC�=�:z�@�XՁ:��"W��G��ˢ�i����2~�	��|��n��	k��n�`P o!�+�#��$�ƈ?�n��smQ�@�i˘�����`�W��.'{�j)��=7����a�)PUIe^�P3l�/D+���0��)yN��o�R҉ ���K�Ғ��*�
����(Z"'2}ʉL������2(X���E{ݾ�����*t/k�H<|�.�F�Gd�9��s��[���]�NW�Qb�b�����|Ô&f1�,���>V�aG�W�ζ�b����GX���zb<I!j��#�Lsu����z�z�5���΀@��Sy�
a\���WTn����ݪ�>��ِ��li5,�h����'d�;'H>5������U\1ۑ08�ȝ�!\�ɖ�x�����; f���L��x���Z�Q,Y b�k���
E �(��Nɐ���$�U�
�����T�F�V+�����Q%���tN�k\m���8v��6=+O���Z|�	�g�GMޏ�����ZP��)�{@��� ~�����5�u�����f�֬�M�8]F���p�$ʤ������@T[�j��}o��B��z��zcJ R������S��c{7�>�.Y~i*X̘�i��O"?h�%����� ����}�'>��bƨ;��kC1ݿX�T��#��p��`��i$����c�a�F*��\0�m l�o��^_g����u)��2w��(նZ��q�u=UZ���z�N����V�_����}<�>0�����_5�p���K�8���c1�=�Ě��iw�.@�To�G?�	鬌��6M��N޾o��^��w�+�~��]��V��x<O��L%��P�sj�e_w&ę'x��c�k�P�
�Q��s�Ջ�E����gh^y��������͆�g��rL#*�k��V&��3�©?`�Bk�`f�]$\�Y/���Ʀ�Q%/&�>���WSY�	fg|o�����|KmAߌN-�س^,�C�ҝF���5����l��馔������13�H%�	��v��S��V4������2O�LydH?h��ߐKs�8����,i�m�e�m�$t��*l�h(��s�c��h�N!�*�j�!d�F�b|+J����G�ַ��kZH!5X:Co�"Ĵ+�4�o���p���� 6�����矐TEV�-�:��4"�'1�L25�LkH�_�Q��p�=�q��/#w�׀!�D]2s��Ǧ$�鐀K���(uۮ�zy;��� ��h�-��x	��!���0��(a�BOI@�����F�2^�:�uW�-YB�h�)���[i�e4�K�F�(M�������=��&+:6#=���ú�q� ]�t�K�=U$�_�h�v�Nn�_���F����Q߃`ݛ�Ng@�ͫ�H�K�jQ�i*!�F÷ZۯX0$�<9D�*m�c3|�}T�l��O��@8�J1Z�3�q"�cN��)�%gሹ �����|��9�r�]�~8JR���&��!��G�5i�B�.�<�vY;�[o��
�����z\�F�>�6�"�xr�<���5`���u��Q=X���@�TzDt3����O���"T�z.Ҧ�p�,O2�CU�;٠��L�k��m��2fm���^"���&�"�N8�->��C�*�h�ׂ�Ǵ��zƴj�������R��S��1.�>ٟQ��TXQ)u�a,uB����z�����%�5��s�(T;�һ�5���UY�o�B��	½���[��C��ƅ�c��8�J�>��6�7�T_5�=w�K-\�q�Z�� ����7~��77�f9}w���iωw�M����U��"Y�޸BP��2ɶ�ٸמZu���U�L�\��U{ʆ�Hږ�>�n6L�(�rK��$��H+�%�{L��L}��֐4�ai ֖�iO4�#:����5�\
�3*�~��Fq���w�X����JC�e}�c��ymM�4V-`� ��QR�/)x� �W�s_\RŖS�f&���^]�ac�zm�\��;FE�%�:ҨYϙ��,��K�d����½����:������{�F��p"ª���Y:��f>W���c\�����J����SE��o8	4��4]�Q��F_�>��B�4ΤB��R}g�d4G%�?2!�+��L)��G$��<4�.�WE�%BO۳����Yf�n��,�ǡh��&b�*�RBc�Q>��l�%[^�����|p+��B��� �D�p�Nu�>e�|���G�;|��WNa�HN�g����w�>+��.$��.m�I`��� ����)��)^?E�p7_�o(������
5gюl�X<��"��`RD���0�u�Y�s���\×+�Z����c�lNU��c��"�>����5ZM��Y�4�Ԙ�����D���'y�5�_nn$ʮ��:#�������,��b�`��0��V��o��j�`���(�@��� |�N~@��	�)o��0����}�_iT�����*L(�M{�*o��=ԛ��!��	:1�͢��,�}��v�­E�U�|���ՠk��ca&�wV]�Y��%�Ƕ����`��:�}լ�WY�\M)�rMi��Y��K��R~y��s��*!�K�M����M��>�b�����Fß���BY|a�];�=���,��yq98��DC�>4��pn�1���IR2���E�,�]E�2M@2}�Eְ���|�0�,p�3� ��D<L3�;��b����?^�XOp�mǼ�V�z��4�x�����|Eˎ���"a�]z�HR���7a�>אV�8��ŘŔ��2�����Ԯ+E%E�άν�w!�d@��»�la
��"�?��Zњ4γ[[ aH�ӿ�F����n���G?q���ѱD�I�=�g���h����_���<;��k��s�5»2�
����#t$���U=|h�\՞�>_�3k�����d_�z
0�����q�g�VI�ĭڑ}��F��ae]�nH~��t��e)����'o�(�8��0��ݩ4���/z��Z�X�3Aa�I�J
%�]�^�P�}�eh�F0 )+�1h�7s+�� YG3�� %�`Z�e�i��sp}�Jχ�����1��#HW7-I�C���7�φ��qc�*����o
���ZPw���Q��`H�{J[N]/�L&���E�i�.� ��x���r`�ڞV���Q��D�r� CI]ߝ�s���U�&MS}0 wJ.N������\�`���H��)���&z��_}I�&��0�p�F���A>�]���ͫ�]O=	�"� ���z��&�U�z�����d���9Z��"��啊_��n��k���ה.M�҄�=�c14�7�^,�d5��F��=d���!CG�\~d䑧9n�^�承u�lB8X��Pf�Z���;��5j�������U���!�t]�S�q��> j,�P�g-l���1WB���qM$$�q9�u.���j�An�V5h��s�3��^I�[��o��:���yOMV�g���I���i6~=�6�!��-15MJ��b���W�`�~E}��#i��NKl�J��!.��F:1�y{-�"��R:w��8W�92l�i&6�@x^���ڻ脙�3F�S|ݾ�w-t%�z@,2G��]����D&������b����@ ȕ����Ͽ���B�7Y�m-�K�b~�~��aG�QH}zGw�y�����3���Y��y����F̘NWv^�-4��3�ƅO�:i.MC#Q������k��GHn8���\>`��$�ǹt��}}�<��TW۱z��N7oiۖ]�)u����l��5��hҀR	�Y�&�S��M����{��J���h����z�]UJ2E���I4�,�L�����+�L3�P��ſ��z����?@^�oy��h�o��L���d�5�؉���s���2��r��9mܡ6�{A��?@u{8P�Y#Ϲ�E�"'y-���Z���W��,>�_υ��0/��a̬�*�G�%��������tͿ�ڹ*�9u�v)�nY?]�H�	���c�P���ź�׮�PJ0wu;�nn�����`�k���ބcp��kw=ݡ�FegM�K/�X�v��%�v���jR�;m�Sg��?��-�9Y�V���AaR
7no->���� �igs��d���)- �}�5�m�b��!�w�����[\����Y���	���׀Pb$���]6(�k2X���4"����,�.FV9�`g�C����H���V�r�Z�:��U�w�u+�+M_rP"�2�އ���&�w-SF��N8�����o��`�����J@����6Ͷ��Lc��0h�Ўn�,�j;&�)s$zp|t��;w*:P����
�t�w��u�].��� ���˦N���uj7v��8 ��\kf�"J�m�U���)ȭ�z+B�p�;&��;�K�9��a��I����~D~i���)��"�VYy��f�1�EXFd-�5�.����䪰o�͎-�h;�i��nLh�YQT���i��-Af|�3A�,�Y3o"�XHD�ه�K	${�O9������$m�JU3���A�y���!{C��z���܃���n@g�Fp��}g���=L�D�x�WB�����QAl�-Q���.�o��Sw�x��F����ܫ�i>^��/_|o�P�*9lPBU��"�*��}��"R]��.���5��mh��8C���g���:DMrm^G��AuԷ5�i��&A:�B�ɜ�q�dnN%&?�0�oigǫ��Y"��d|bv��b{��ө-�W~��������V���6���\եS�}����%�O�N�<Ӫ6��1�0��z�r����p5�@Q�K�r�L5��(�HS(kkOu5	j~Ԓ�dm�oPx&�{^�l��̜���"��2b ���?", o*0���:�[H�(������3%Rz+�FEF��Vf��,S:<;K:�j���V%1�ѩ�q��U�6�q����X��6 _
�sp�y����+-���oO �/�b	�зe�m�C-{��Zϐ��w�<Q��@Ȩ~��K�}���a��C �ɟ�1ճ.�+~��4���TX�& NL`
]MųB`d����D�C��IR��CaЮ E��|TKPr Mª7͉�����I�u_R�y���{L޾%�Ca5p|��\xOpC�|��
��m�A�?+�';��HJ���//�U[��2�mG.F�dG�<9n����tbΫO�C�2^M�
Es|�z#��XY���ߕ<?��"�jX��x��E�""���W��rP� ox���;�'�;\��c� ��	Q�T�7�\��[/~�(��]�T-6�`>�j�'ahW��ixr�����dH���Bף4�E����6��?�5��V,��8�Dc�����o�c�ӎM����6�G_�h�{h�������~CZ��9\s@P�L�r�}�g�,	���7�7�h�9�@T�2�$T���.�����BPl�l���l7��0.3�2S�����e%f��a�1k��S�2���%{�� �M҉���3��љ�]���Y��\�yү_���yz�vݖ'ӵ�)r��:�tךv<�����A�)]cZy�������Oj���I����7��\��tI�I�*8��努C�U�j�t�(�ж�L�EY�9�Ǟ[���4n�96�Y���N�t+�JYCR|$s���ț�6�6�@�ࢃ�{&Q\�8+��I׊Ƃ)uGH(cBR?�K��15��+�>~?Ƥ��h�I8��0��\�%���2	��τ7g��v\ծ����=cXoP�[`�>
���xk�s�*�8��>4��9�O[(����0�2�z%Ѝ������0gщR�Yb�����������W��w˸������̃�N�� �ʿ�P�L��� ��y�E����~Z���_[+�����i��
m�f�54cg�V��4�]�K'�Lj�tP]�V�t��]��kދ�[�麏Q�;](J�����QIh ���f��;�nf�<.:_z�?�Mu;�\/�h��B�)�)띹݃�i'A@�����ɰa����L��e��#$6Λ:6�Dy�����������a�h&��,!/�L�8DN�/q��(�-�nJi]*���'d�4w�Q��[�Y��Z>;�<����Mg E�2������n��ߠS���>~�3
��1�9�;L5y�:Y"Z�b��h�����`�2i��̋d���eV���`QR�N�)(��8 ���V��_��౯u�r�~#�-O"f6&���ߕ1��qbnc��uk�qt�N�������qֺ[U���k��!}�3�v�xQ��~3{��څ����*PY{YZ�w˸�����z��V�3"��YAگ W�C�۞MjO�llr��=璵�|��*p���*�q�S<���C�4��'�1(�b�{]�J����x,I2�V��M�*K�������O�a�Z~����cp�.�4<ϻ��/N�E�v��qI��B�?�-��G��m��Z �o�� Qi���#&��"�ܴ�&74\�h��W�"3�|a�V�� w!\�0��&�ܕQB:g��64$��ܔ+
�/��4��OP2a\��E�ܧ�����4D��h6�F{s��2j3�/���z�&L�'5YN�a����b���Z!�q���C�q�p�5��G�y%GUc���`W��I�iN��2x�rO�Bb8ǔ�sMo���[>3�%�����fH>�EW�"`#�N���L4�`�5|d
��̬ۯ9U�H4(\
��
m�*hjd8�&{��7��Ux��Ғf��d�O�@y�y�����%_�J�r\y�%��� yY�s�G�:��_c�͟tdR�p*9��e��L��J��-R�ԫV%�o�Rvr�>9�M߻� ^ %L��$F��!����.�����s�~-��]/��:�J���c�(��?����f�����e���RE*��иoT#������\ۥ�ܬ�nl���Ed��K��/�58n&ud8�aE`��me�Z`��<���|R�ͬ��}���pN<4��xϧm�@�?n�K����f�w&�����R}�L��̌˯�ܾ����T9)#���at���R$w�
A(=��T�C_�d[��r��|	1�����(��xoO�Y��Vu�Q�4�d�:dl���SB���0��5rzҌ}ѣ�/L>	,�)�T����R��`M!�J�WAg��w�`tS�9V�?�ڮ�0g�V�Sa"�/�zl�;�=>gƝ�b�L���g�W�Ki҅��m��]{o�A�K,�E@��&Xջ��|~ޫ"���70����)��כy�`�e�,��Τ�{Vn����-�ӕ����ۣs>���!u����p�a�!��(MM\<��µ��?s�8ԣW����_�ż��~R~3Ѻ�I����D(��7�د����<,��.��~����>:��Ū)E�������S�sy���ocx�|u�����Mv�i���?���d�";=i�Rc�Q".�#<{C�z)��
R�jP�����n�U�����x��)�e�簋Sg�2��Ƥ����Ɲ�����d��|wھ�*��-z�@f�"�vl}>��k��!p����g8^��L�x*��ǽ7�X|�bk�_�!
��O[�S��ǯ����,�m\O����<L]� ��v��� ߈��s���z@l��G�����N�}
E����)�`�N�hg\?�hT���$s5<Τ�X���{.�`�m���T�ź v����qU�gr
�?ɸ���)qAסʹV�3����*��s���XI��㨋k��8Gx�_�;��s���z�uUܯ\u+P��_zr_S�����3l<.מL4���.�x�i맹������㾹Ma;�k�~���4=�Ԋ�C�,5�.ִ��-'�f�BӉ������
+���2��:����`v&B���CT�[7g8�9:�$��;�D٬���0��CF��������b����a�t�A�f*M��֍�{E��8T�T��A�����A�ʻ�06�,��i��[��F`b���~^�ް���}A�t�Bm��	ԚH�}l񘅬��/~V�nD���߆��t�T+��p}�#����շ�lUn����R�7�S��q_{1�7|��,{VER	�ԁ���f@�
�1U�*4a���%�mr���5>��,>Ҡ woJ�a��Pn������J��^@z.�t�؉1�p���B&8T��NbD/wA��D�h�>*3��1=	�@D����%���m6� FM/?��u|���!ֿ�B�'Q�;�u1I�'�l"2\	=��c��g<�m��K,��A~�;L���m��p��w�?w7 �`U�r$�7����]��:�d��3�Sl��C<5u��O��r�~�`H��� :b�5�����̙c��-MzZRG�������Fj�n��4�g���cЂ5Y�Ck�#ڭYWp�Zbx/���*w5��q�	I1��K0�X���!����|����5�[���VF���G�n�N�d�z.1��q#�웦�ڷ8V(e��ck� Tt�.kYO��3�b��|�{�1��2 3]ȹ�N4V���*�%�~Q"ڮ�=�\�1�� �h�"�+h��h�S}�=�������協7�Ӝ@��0��G�/e�0��%h��kČpYՃ��a��/6]��e�r����I�C�<`�7�ۏ6�`��՛=�^6�aO:ʭ��W7L��%��D�&�5i�o[!��M����W�U�a2��'�u��2���
����N�f��x0Y�g�(�G
H��F.�Ɲ�)��[���f�X(8%2Dל�~KE2ݫ�rk	�vB�e��2���	�l[�m^ 