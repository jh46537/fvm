��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7]�s��^TC#�yM�g,�%kڅHе6��&E��1gm����J�)d=(����3#���H��Ɉ.tc���ҧuq&&���:�
#wH�t���+�b�;�$�O	g'��E�6�Ҹ��h^"�KA�:������a�Y���2� �I֕'�>��%#M���yB�D21�~�	Ez���ĥ@���6��[(Y�+�X}��-�)�$�����5{��f�|1��	Ɨu61�i�9���u��{�7�_��ol}�C��k�Mi� /����r�U��L��o�8u�#��!ɤ��G2��U�,������#�� �g$Б��W�h��z��IF����&���o(?�i��C�S?�LY�Au/�`̙p�*�M)��h���o����;��B0��s,����d���?!��^�'Voײ�8X.v��k�GsQ�rY�K��.]�j#�yT?�v O����@
֐���t�cR��Ħ�HOIIV�����t<c�����<��8I��ջ;��8��~{�ˢ��=ѵc��� V%��䤞�V�A������S���)�����j����S `�nkC�x��<�"$�k��_s��7~4�pu!�VO�����Kz@U�Uy>�>ɧ��<mJ����u?z���B�W(��=&�/MjgڗS'A𞟒��:+Ĺ���c2CU�������q�~��5�b�������+��䠏�p��;�	�gzӟcO�&xs��"��q����F=�Z�O�o,��,��I��e��i�,b.J��_rY���P]��{�T|(�<�5_"g{���j@L�AqShi����y-�+C<��/ )G�m��z����'�r@�u/�l��c�T���s�h.|Pz3:�N/aux��A�6�O�IM{y B���%�+Ou�P4Д\D鵲]^&��W�r��Jē��4�<�?(��2�7����E��AJ�qMQ4ي�Ӊ��_Ԧ]ܶDNx#!IP������Y����\Myn�[��K��rjvp��gBXw�._�U��	'"v`�L��0�ȗQ�nF Z��^���)A���G�q�NS[Nm�~��
���GT��]l9�M��d��MYjgZ��:��������x �s?���o)Z���Σ���T����1^,W6a���N�)Ԍ�,yS�����9~���V�S�Y���;s��0�����'l]�5d\"�P�m�d����'@��B&��&'��r��Q��T[�0c�i�;��#^��,*OerI߭��E��h�}u��Rg��2{��l�du�G�:P��z4h�5
B��l6
�1��M��Wb��n��+��rp�6�|���7\��&��ƭ���}�N��j�������YXQ��_���i�
���iz;��z��S7�7N� a��y��/��h��UΡ�g��ҿ�]Z�V�'S[V�,]��=Ddg|��U��>��s%���_+�[֟���撹�'�#$���@Y��S�Y_� L��iV��fV��#�����v�}�o!H�,�Jm�DHr�A�ɰބ�K�Z��#�3+����f�e�BW�|�j��U�Ļ���)���ѷT#Ǧ-�DZ��P\�<��!�3���ޓzruD,��WQ��B���i�*�<�K��?Q�Ŀ�V>0���yI�@�7^nڼ�6�����|3�&�c���b�.�q��}����3�q�/E��+~�N�7vTb7���	��Em �*K]V��:$ܐ�ۯ��U�X)�������YA&�Z�o����+�L,epU� �-�(*Ox.�|����vٿ�n�Ȓ5�XJ�F(7)�f�����Y�H�Uk�
�\�2����TP&�F�E��c�����Q�_�Y���ʤ�I�_y�V鏊qذ�]���^`._Ґ�P�!�	�o5���M��m@��Ȫ�A�[6����;QSI|GD���-�&�[^��j�ưK���c����UtH�C��pC���h�0I��"��̱q����"Ú��������;~a�=��zQɃ�YTQ�KV�g�HNM@�/�[���cs��p7�����8uVl��}�X�tg��]�_d7X>���Jp���s��>O�_A!���'-�*���J��}*�s�{/E�x��;G���
|��� �8[T1fgj������g�����XO�{�	C�ڳy�|�ĝ&aK��[�B%�Y�<�+�9�9��46%���2A�;���T%�ȁx`�E�'����J��s��; �H�!c��S�����\�K��U(y�o�hC��;jΕO�~��k19`�*�E6c,��INOt���R0ͮd	�MM�S��Ã�Mq�ZK�f�K@�Є	�겇�[�"']�L���z���%���TJaj�k\Xɇ��9��<�!�@��������b�'-����2��o��0M,�H������*�t�%���L_f<~M�,���Qo�v��)+7�$�F�O�0��M���ⴏZ'�v`��Nѯn�!�-���U1���9�����rtj�#�Q�V�1�~e�[�E��'b��pذlr)��y�m��Q�R�wY���P�]<��Qqo�%��KA[N�7�J�1����NpC����ꂔB$�/K��=�M��'?��DͰ�$��O�w,`�A`���l;
!$3�HA^�n���o���ss1��`��2s�0z%I7SKe��}��#y�e��YҦ��:���`��]G �@�6$���~o�O�?�gWdz�6��6z���J+�Q��qh��i���.#�dw@о>+���m̯���ˌe�a�HT���`��;j� I�����c�f���G2�<�'�BJ*�^Ccsy}6�$ḉ���Z�7iy�y��4��`���s��i�t��Z* ?�U
��� 03#+�������䠂yj�wЄ&�(r��ķ������T�U���T��/�`f��uѪ�ӻ�=e���vW2�� ^�9�I8��|z��Hn8@d{J����8#����Ӈ���c��L�&���p���ѷ�f�qS/�a��e����ș�7qn����̏�Cw����}��G��N�cs� T�jK�VPh�ݽ�]'���x��>:�$�S?>(%7�+DJ�׀�zm�dЕJw�ˣ���f���ag�HT:s�ѽ��Ո������'о�7��c��\hf�ˉ��%߻M8�vj�%Z ��4�TZj�zoԙ<���4hޅ���*��[O��;��u����8OZj��>;�ÇS��t?XZv���=���k�@��(��i@1[��x� Y�7�i�>.���2�1���C��;SlPZ����?�>�
��D����T�|��d<�z/mh��D5��Lɣ-	j����mTgD�4vF��G��	h�H����9�Ms�4�������c��u��rVv��,PT�@n��oLks:���w#���H�tO�@�@b��g+�?pDV���쌧^L;�p	�w��Dx�P�$bE��b�F�iA{y�K�3��i�p,��cǇ��mX������?��T�x���ʫ�t�>sJ�z�Rq�n.��:R
+��F�b�O���ÚIV|V��%������,<#�!�տ���&����OCF'u�3:��~��$j}T��~9��J$t��|�u4����Y����B�c�؅�J����9{��\�������"�e�8�0~��'5:�T��sOG�J��aaǳ� ���GA �Bѭ��<$m[@�A�.h�kb��xнt9���-���I J�8�}�}��L��ݱ�{��F��/�)���R�������+:==Z%�Ҵ	��14�k��D*�X��z�r��:?��!
,�,�ѭ~�^]ʯ�5#�zP�������F�ճ�W�%�23��ŌO:%���WۆGH�@��+S<+��Sr`�>41-R�	\��щ�3�󊤚D�j��F]�[O1)ˆ�ˆt�y�S��w��4�����5�v�JU�g�~�[wGh���Ea�C�����>'Z+����
F��&�pE�*�؛��v}$�p�ЫZŭV����.��$�7�sn���\ߊƀ,��ݘ�U5����Qܱ��<��m�~e0��1"������H�@7d\�� �]g�-b�3ȵ����,ؙ��:S܍{�|E�`oe1}e�觵,Q�(�����(i�.�<�k`��=+k�rk 7w�>����2,h
���N�;蜵��q[\V �k�l�U�9z�
�3���䜧P�zbC ��v0�[1�x	�rJK��q�ƅ��X��A�{������t��!1l�E�N&q�t  �����C&�~W���%' W�.�b&!�YE.��7=�ǵ�+�!�]ì��k�k/��������?������u7R���	N����R�D�{� u�ѡ{�5���x�c�<P����g����yIx�:��1F [���G󼿣|����Q��J�aN�e%��n��%U]}H�Z��������
޺TK�8�+�`�h�r�2N$�\��x���Zό!K\�Ajp����B�V�0�E:��u7T�W/��cHQ�;L�fw0}��x��M�	�d5���*(�� 6'�����b@׻�'�������u��g2/#���6^6��M����7�36}m��rqB�Q�ʤ+%;��h��h������ZXMe��� �@�뜵!2)cԇw�G^d?�s���'|M�t{$�V�{g��XŞ�a{@���>����䦹��6�t�<��+'�ҜW���_4VJXA]�C�~��O�{5���G}!�V��I���t���@� _���W�xdt�C�q�w����u3X&m�5����|�ʁ��?��Q�i'�'YΑ:)��Xj��\�ϱ	�_9��dB�r	R���fRa�,>�e�{5��e/��25�GoZH�B��(	�QKK�#}rH���`3
�Д�-}J3>f��wY�`���<N���	�H����e]��`ша�r�B]�'t�*խ���>�� T��︐u��R��ij�핤�W
�V"�2��VrIZD�̪O��ʍ��:�M��Il��NIX5N@&���d{WV��5Z���7O;^�Z|n�4����Yu��GfqA,�b԰�G�5��I��H�������6 �zCU��d�R2T)[@�0����8)>�#�M3�pɔ�:�j�i�XXl�;�qf����T`זdT��D��W���i4��e,CQ�|[d}3��4��fϴ~sջ���MJ��/[���+r-
�~�e]�a��)�$�tF�����CR��yA��v,�
��v)ir��ses��p�=L���$۔q�s�x^�"fc0���=i�~��7$́�V��ai�l�����~*(V�cl$E�&�C{�hE��q {��t�����9n[��lez}�I���IM�8��B� 8��g�We�l�{����48���/��MCí���)yN�T����(6
B�R��r$5����|��Eߍ����R���3'�V�"��?Ӿ�ld���xN| %@_w��@��Fe���Pf����X��<�g���Y���y�T,�V=�u]�M����7�P�@���#������0\�1IyDr����Z������Vf���gב��<\}��KbR�����%�m������J���4��A<�>�/��@���p� y�H KB�ղ6� ��Ot�zQ"���\�Y������w