��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�k��&��Bvx�s�!2����-	�C�o$���%��e]YC����td���bQTTn5��r���]��ו������`��r	��ڈ^�5Ng$�]��� ��ڷ$@��VEbs,��v��a1����UiYAY�֮�}"�ɛAJ����Լ�N�$��Q�Z�����I����\�9Z
zd7���<$�
4;���/xLUd���\�נ����{��?ҿ����8Iј8^�6Z�,z�7]��Uj|dӣ�����vE�����{�M>	�V���_~v���ܡYQ|{s�a(�lK����,�>T��3\���,e�US���c`b�()��+!�H�q�]����CV���F��^�~F1� ��+F�H7�IT�!�S�K�-��cW����=��8!EM;�X�ß�Z5���71��a:�CȻe�(�;N1;�Bi��[)�{��c���	/�^��;����N�Q�e`С�5�E�+�:��~��"�?D��H]μ6� �SgY��!.:���:���y�u������r�J�
K��{԰ֱ��.�W{=�u������蹖3"�J�'U�a���Z.���-{$Gɤ�rg)�!5i��杕؄` Nн*�hu7X��\�t��Yf��GE���of��sqR�3QX�Ѝ�����Ӑ��셎�m�4�I7��[�6ܙ��?�صw����;���8�wO���$)9q�_�{.���<�j&X�Sjˈ���|�y"ܕ*���o�{��5Va�,�=$�	γP(�]�9��P�f���a#rɦ����PzNTZ(ZC���jk$0/�M������l(Ҥె=�|믗�S��� �Soj:�3/3�0������Ng7��C똸���q'ۈ;�yŜ�oi��c���t�>��3���P;#uRH�aE���T�.�{���Z�RA��L�+|�.��I=��X�t��|[s���X���@n�0?GA�l6���i�>jC�X<�K����4�m�A,X{Y��?{���R��g|��D�E�9��s}53�m�V�'Bgŗ�z�r*�RG�ۧ\#Xk};hP�hΎu.�ܩ���<}�@�gA��҈�v>����/]�:?�ȑ8�����)��ZO@>��1��}�m,���	i1��zG����^K�!3��x�����3J{r���2��v"��×���#� ~O�Z�k����N�F�e[йH��ѱ�O9/��B'?��z:��`[��Ԅ-sK67���40��`c�X%i�W��yɋ�E-X�y�X��0m> ��s�A�i� }�S�Piӫ9�,>�L�ɣ�Bb4}l�0�~Af�D��,��fy�����&���t EH^Z��
N�3�T�e��ԥ�Ѿ%�X�*�.X�4�.��]�;�8�5Ҙ���������C��Xi�Il́ɊaZ�Bl!=��&�s ���͒NT�K�_���8H`[2фyo*n`'j6T~W����r\�6��a��)`��E�ɗ8'����Q�����a3�/�c������à�^!�;1���/r��1�wR!�	,����_����0?�Px9������ٔ�SJ��9�X�B)v��d^G�Q?2&������x�"y��L�.Z"�+Qфٍ�J����n_�?V��(6X_Cm�;@�,��Xf��~���,��%�ŒHz�o�n0���v�N�qǗ�#�X�Ҹ�g����	lvO�!NpI--v�ݎ�l����q<�4	�w�wQyB�l�o ��-�=S�ϑ7؊���^H*�tp�v��uW�׾(E�x�)���g$%_J�ߪ*s>^�w�s�X�/?3	h��U�&�sKm?��uE�$�f�����(���y�(.Yq3��A��!A&�'�1P��A�꩖ �V���.��@9��b)✰X�])r��s�@CS��>�:��d�2�q;kHN"�Aز��q���w�EI<��rOi��?W&�!.S���%�25MԾ�h��ax��¶`}O�{�J�B~A���V�r^gN�b��ۚ-3`��k�H����*s����S⬉L�u��$�*Q��80���#QV���y�b���K�@��mg2P@��YaCK ����60����.�ؾ&��z$5���)G��.��������ۭc���(�X���z,Z��b�����`�����i*J,~�#Uk�6K�9_1 ��h�z�&`������Q���3�ءX�7�xc�%�j��b��m�>T'Y��wT�� lB1���%J���+p���C��Dh��1`�?ו�a�!)�m�]���G~�����I�{�g��Aݨ��ŧL@�}~�*[�#����R��y孤$��H�V\Z����:��h�����z;+w�v���<	����<ެ%���F�����@�lع`�LNc�$���j[����Ho�>�N�29��<��D���dY	șu�/ݡ�|I~an�4c�d:��vY�2+�o����֏
�9 �����l�� ��n��#��C�gwNYc�%��#�iW�,��r֍ğ�l�|�`܏�'���&Zʹ<�LG^%�w���fȩ�9p�>s�,��J�v�WH�0K��b��$�$������B�oLR"���xM�c�Tky@*/�GQ�'��ڌ7E��
=��H&7��({��}K	����&�Si���㖵�|����A[�ʜ��d�s�S�5���U5�n��'��:h4�nR�S� rU��<������`���.J���Q*��S�5�>�,Fh��}D�;�*,+T��wterkn�;�Xθ���Q���!Wb� .�0��˒�I5~Ĭh�6��NfM5�%)�\�������и��@îߩ#��5�F��hm�RJ˵�*d	��9�����j`�+���xʢ�Q�6�dylc��ZA�������h\��T���w��G�H��LE�1�?��6�uX��e0�t2�y��@��s� ��Pk�04�sU�`HO�B�_��,���pQ������g�[����t(w���G��Ge���b,K�иxsˍ��pW��h���49������d�)I����8�kA���D��ʵ>��!�Dҫh
\oZ�}�M<f�+��Q	����z?��Ab�[)����PL�6��,����>.����Zx�OEW�e�:��0�Y<-b)Ћ�ئ��@�_/�98��Z�f==q<zJ2�=�=�v����z�%j	��i��6��IY��lY��S�( �|�j4�A�Yk�''i9����͏�D$<���ī�J��A��L��j�2S��i�'tx��6�U7����`��p���DMY�0a�_{��!�nQ/i��n�Я��p ;�r�xx'�iȹ'��P`�υ�R�`���u'n��iX��s*�	�~���Ȱ%��Ze�D�5�D��8�bدjAv��Yv��8[�8e5������x|�-��*){����[�jo6�����gL@���W����YY]��*�$�$���I���3�2�6'�6ք�f�&���\[-WJ�k�<��^<o5P?�|���e��:J�Q�8˅�pS�v\%�o8r ���;f�g���w�p�`�a���P�*������ �?'N�/5Wݲp��姧�<u�P�
>0" �u���gE��w���Q*��`q��{��%�Ǝ˱S`,un�M��P׵�{�gr͗1U�(oÛs7n��1l�-��kn�r�%����{�yD�V��<��H$��b�kJ��$2-H���Y��W���!����ԫ�� �z\ػ��5����;��Ǥ����ėm#���A��G�}s�u��=2�*M]ԃ�Z�:[���N�ͼXܞ�O7�_�]��{U��A���_�|ϣ.�j_ ��������o�XӨAH��_L��)���� dLF#����b������/�O�5���(}��K'�fl"f&_d��7�]8�:��<u�zj�V�����H4�mob�X;y3;�w@�\=-G�`ػ�X��­�u��r�ǰ�&�n��%y<����u�?��y��V�4w���g'��5ƕtN�D������Zɨ�w����;��S�U~����r7wz���<c��7`J�v��B �u�a��x���H�ƾ;P�͝�[rw���v���4��x�i/���=AI�*~Ӷ��,D���La� 6XP��EB�7�Ah��؋�t΋TvK�֠<ln�C�=�,�%xOR��u��Tzd6r&Э�[��y"I;TE�R^�9�+��͑�gX��-Pɼ"�'*�;�3�5��.�/�0��m��f�c��봓�6��݋;F��zݓd��=����zr~�<�R�fD,u�KԊߕ*����꿚Wg��~�!�?Zn��ǵ��IO&��繙� ����*��9+g��2ua��" ��A�K�4��	uO�T0}�>{f�ܢ� ̀�A^��o[��e�6J�b�yJ��9�aߓ����BN�S����WgO�Y������U�V�`�j���.���k��	CX���(L�6���/��Y�~X��D�����r>Π���~�!��(��K;Aں*��ЌC��]�[���v���F:Y�\V���H���$�0��#��[�v���fO�8���!.s:
2����;My
V,p�gL���(��f��E�$���2�V�G�8�Z��孵a�Vܞ�"7�Ͷ���u�ڜ�����A�Z�5�*�R �k}U��f��4�͈G�Y=������S��%��2H��1�э��uW�MY[[�w� ������^
�Ij5 ��Y��ִ��v��p��5�e�70���\��F䣪�~����rME�����b�my!��{L���y7��.  �9����O�<�4��*�dg���{�=�;�?-<���r>��>�7Q�k��f3�k ���$w�R����};���՚޴�&zy�:}�V,���,*���R������ˤ~�Lf�����ì�Q�&,�>X�+K�W�*�qє2�D��0 �=_��m��>���OJw��y���wL��"&3��K��䒯���Ύ���^&*�9�y;�2LJϹ?K�q$(\Z/%v^OR,:��P,j���f���[��+ʅ�����F�t���f*�78��t(e�i	�w���4���V��"�������Pu�cn+��U$#lr�T�ζF�rt!�?J�I�%��fj�2��Wʑ���3��%����BV��|Q��,}�f�ͮ�c9p
�P����ߎ\0���ɭ�^�s�Py�=� ��2�ʱ�����=c���@���4S��=���؟*N�w�3]
��#�tH.�\�$�ʢ�N����?�%:��c���L/�^Rs�^�2����&r͇�"G�k�/�4񉍏��I��}�Ht�ƕ+U�<����dw�����ռٹ��y�E�i>_����L"'Z�L��ȁ����1Q���P:T4���)�ײ'I�:n��kx�Ŀʧ�u��ZfjF��H��A{��QJ/�&�X���6���V����~��NIQ�^t���x�U�YV�o�)N|{+F�q��u5���S��%-�Zc���\bE��iiU2�A�_������
H$^�t��ݹ��U�.O~M(���y���X<��,���
"�%>si0��K腐� (&�ٙO��ox)V��[�2S^���_zP駲�������]�
'�"�7Y���".����Uۥz��(Z>��QԵu	 X��G^!�RI^��G�Y9Zs��tT�0M��������{����&��l����6�>��ho���Ю�/%�l�ɘ��b�D(�gI��FD4���@&$��P��0�Li˙�&&�0�2�Ft7���<�z$�h�p��^�>��7$�n�8�BE����֎-Y:Ba'u�����pq�= ���	���s`Ѷ��u��������ts~H��4�`:��T'��fiիs��X�*��'�����i�d�ĳ\E��DTǅ�ʱ)�vT�^G����T_hϾ���J�\���!n7�Ɍ��﹠s7D�:��ii��zLo�U������]N�c.�BZ���Lx��Xwj�)*��
��,ȏCmLJ
 ��K}K2�z�) ��6���!5g�̥O[Ҍ]�:�/�"�
Y�o	��D�W�_��ZV���`�Kοo�ǥxx�Lb҄"�%4��b���(�Op}�N��v�&������h7�;@�=��6���b���ƅ�)�L�`զZ�L=l�����6n��TmJ�M"� �!正)��݋��΁�a���:���
0���<�9�� ښ+���wY�f_�M��\��ڤ�L�����y�w�(���&��r�Z���ߜ��H����AsO�:D{�����������\��[��c�A��ɺ?����l���&_H��%�����p�|5{P�!F��j&A�rqc����;n���18^�U��J�`��*{ы�2~rn
��덻�zܫ�]z��m�f���� �ݞ|���]gA�	+�d���:���[O���z�	��g�<�֣���e/�o�UH��P7����ɽ�g����@�l��A+.J�~r��6��،��c�;K}�Z7siюDj�ʗ�u�2���