��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c����}�����°ȣVZ>@�#�����QW�|�i����#JM[fsW�Cu�6�9��U�?��#�+�r4�B}�a�+�M MF�"Ҳ��"txOX���q�I22J�{�|㹨�3�x�w?�Pbx��Ԋ�;NK�	��[�\��H�@�.��y�GPS���A��,�V�l��O��8bz����>�@�-��7������M)���yg?$g,��R�wΕ���z�`�O��ogW���~�j[L@�ɗ�/W�qp�����8)f��x+Q��_���ޜ���q��&�v�89c������>��QN[��p�-���睌OЈ��>k�+�ף*�U�M+��Z�wS�<n��6�J�ݢ0Ɗcl{ ?�H�����_��I�^�V����>.�pt�ʚ5�Sr�K;�g�\��}B�T. R4���j��}5*�F��(U�)M�-�
ah��*'���r���?@�F��*��?�;Z�� �ܫ��I⳻�4����Ӑ�k�������;��f/3:�Lgx���ZQy= ���$�y�_�he�t�&�a��I�K��V�XQ}}� ��,��wYݮ�i��x�t)�����(ū@5�Sa+
ަi��t��A!�:�k�u\'L߾��:�?�"e�m1��,�����E"���v7�T����1W��q#6K.�[2����'�%����@2Z5���2"(�ب�;fY���M�를z ���{��T#����àA-È�E�N7���lZ�f#�U0��ÊF:��
�H�5,��)�ʦ���A���rT��X7�bEw[�Ů}���������_�:�4�t�CC������?_��kj�b"֔<����p�i���œ���+�Ǳ�V�cT?1ߔ.�#����Mf;cޏ?%��Mr/���w$1�H`��_��l�E��0F����g�;�tOH`%���! ��g��8TT #�ڶ�����Y�\���P���/G��ק��Z� �97���T∙f�!όK�D��l��iŪw,|"�]�DwVi��u��I��F���T����Ќ��A�p>�?��.I��>:�y����[�z��Z_P�4� 9�ؕ��A�x�i�� ��|>;V��ɕu9�|2@8=�뾇p45¿���m L:)c:n�W=��rP�6��a+~[)w�P�:� ����B��2,m����nw�=��%NB���G#w��v� ����n��AwG/Z�dm#�O�̗�.�L�w�Iy2�k��Z�'!ʳ��g'�{�D�D��?����+WS�3gl(�a=���M>lW�	�"Rp�.�>!lm焮����l�{գ-G�I���%��57H�0)~�XS��0��vv� L=�֜�B�t[�%���������?u��(-D�eqn���d�4�c���z32��Pe� ��b�bi��8���K-��'�y�u&5Qh�RH(�h�z�s�K�d�J���t���/��>C��S"U��c�x�E��r-f�
cO�
�j�*�?�y�o݆Y`PVGD�[<7����8IS�����Y�*o��;�����6��|��UuSݧ�o�
�{���YW�;F��]A�ZY����<��iG�(	����
&����Υ���S�ׂ�	&�z�~3�U<�M��4�ƣ�a!W�>��������� o�[WhףiՆ����F;�?��QEg�/rB(a�,ؘ"`��KġR@��3S�d���y�>���mPOL�0�1� �6�/���!J�JV:�IP����J�������aG�"�;��fq�0N�Q��ja2������K���<W��S�c~TU�K�~1(G�w�J$����g���0&G��J��/���#��K���e��1��h��FuY�>_�ڱC۱��i_q(W%�۾����1�h�rHYp�a��W_�(w]�Y>�Ǣ��I+[����3�Z��e[� ��� ���ݘ(oyQ��Q����M��i_�c�N��\r[���ie��K�#;a��X	�}���ḻwh��9�Ӆc���5�CPI{p�]�F�Yf�n���6����{Dr�Lp���͉�^?��/��L��O:qhf�V�w��rO����6�X���u�Z�kQw.����gYS5*Z���OVlMďY9Lk� h"�~?�kwD��P��ŉ.T�������P��MBP϶���F��D�Ί���-�r��������	�݇��-���Ւ--��k����t~��̕�+M�^&��y�U���i[���"�09����_�s�?�w��A����{0W��/�j%��'�W�G��il�������&XH	9_[�:w�~�!�k�ȯ�0�c�jZ1n�!���O��������[6ܳ=u2Ρ��Y��l�_Y�[�s�0�+��(p���p�\��SĚ$���D#��H�&A�*Js��ՂM�Q�܅E��d�+�u��:�����"Y���u��l0Hf����z�o{%~��}�DC�c3[�������l��H��DQH����wK���V4��Ėh72^o�h������I������Qu�p�p�-��ʚS/P���l��*,$M�n"�2����}D�I�C��}bv,�к�GL_��Wjjƛ�M�u�І����e����[�?�$/ U9�G�Z"_�g�`}�:�C"��V$&Xi�=¬���=�׺u�`�~�X|�T�Gq�^�����^�L�@0e>���m�U��Xk
����E(���ԉR����K���� ���Ӎ�X��݄��q/nYf�K��e��S�S^�Lأ���emyp	�!��<�K�y��ۚ��D��]�~Μ�i���?r�2��nt�ט�� �"f����ԁ.P�YRL�@�$�������#q���'o�HS2�!�;3o�$�Q��';	����Ŧ�#fU�7;�'������3�О��������q<{�*���� ����~c��H��	��WNT�ntM+��A+1x�0���&���U�v�|h=���4��������Y��3�rg�AwI�jd��)ߕ6yc�1�I�9���KӃ����i���B���^=ϊΛ>�(\�� ;I��o�x���3�W�@�{�$�sۮ��S��[o���֧�%�k�؄��љ:�>؂���d�M����&ë8>�1'2� ԝ cEܠ��&���[�qu��� ����'�K����H2Tp�߂]��p�'��B]�@Z�}�S���JoN,�y���t�ώ�2өq�$�. ��Q �4T8۔�aX���d��$A�t�%o�#�`��?>e�8���"��oI��K'�����l�)U�bX(�ȗU������!f�a������Ț�E��WعɆ=�i/�`�P��qV� 4��e����>���r� ������M��u�|ar�N����7,m��|���cy�|4ɫ4K9��SE�?1��k�u���W�9�Q�=�g`�צ+$kۓ�-P=�}��d�r�Ma+q	#R�|8�7SCi~�}�\#1[a�F�_� �s�,D]:1Ы���m��47�g��)B����«,Dq�-�5�(�\6\[̷�c�E�Z��`�2 �b�7�AK�� am��V�9�\�	�|x��E�13�d�����^vEJj��U��aC�p�,�ֵ��`�����=ڔ;�b,�@K���bt�qK�oEG$�:��	K�CQ�'bv�ëL�f�9P�ќj]3R���f�E ��
)�C�!�쾒x�7jE4��cI�!t͒aO�(�1r\ظPg`�GS� nD5�!�[���.h�=�η�d�1gy�N\D�վbT
�hq�ȡ�wb�V���y$�����	pF�d�b�?zP����gL qe|���Տ��T۞)���S�:�E(���Ґ6/�'�����㘬e�'�1�����k�R�.-J�jY���Z�	B�P���.'@�64h��\��U�u���r����=��2��b_m�f�"H�ަ;t6>�N�ެRW���=h�j��kՒ�C~��}n�p���NC��m./"VT8 OŖْ9-�[��x��@���]EM����� -�t%��Tg��	�u���?�lRɂ���3^{T�%_�s*����hQ
W�$��҅�.;Hz��<+p��Q�x:���TF��n�=��W�HV��š�g�=*�LeY[���*�MUr���դ�7�D����1�J���"f�E=�����z�0lN��q7�w�Rz�Q6(m"��&g�[u��2�c�?�5��,� �[5s:6Ps "��V����R��ն����f�?C��d�d����C�	�@�l�5b�#)E=��^ Ku�����*�r�ɠM�~mq0�黨��7�h	 ���%Ub�HA��[c6�TYO�r�TZ�/]MtH@�p���g2��FA]�=/t�'3����/�q|���?�@�|�/F)m��V69��"Za{d��K2�|�s�Z4$"|+VO,[�'1qn����~+'��"x�.Pcs�EB�}�p���mOE��'[���:J�afz�����!\���?�ګ]�J��r�ߍ" =�0���Gr�����Ҕ�d7[#ڲ�]I�d�y�k��ՙ��R������I1"p~�p�T�>LM�>;��OB�e�s����'6�\H�{0G+��͇!{Jȱ`OֽI�9R�����Θ�@o�VVɆ5�]�Ay��`�
T�E��^��� �>�`zr�`˟),ɋ\��~�Qw$�b�h��VG̭���ᵣ����j�
V#�C3�tC�m�>i�J��T§}�5#Ê�"�i�2��+�b�V-e��wN�N!�R�Z��ί�Ϭi�Mc��-���|V�1걊4�zSJGKTM*R�Ws%e.�����BC!EBZF����UEY����ݼ�����XM���:zXJ�w �oǠ�b��7�=���Bh
f� �#%��`&#�"S�4I
b�|�_��2�n�*�˽n�A�L�9F�@����h���eM֤*)�^��ʚ�O���ݔ䬏�8�l��:T�@3d�$�*�6Qdw �i��g�߻��1#�5*NJ�5Fhu��ck��ˊ�$ɨ��G���,`p$�>g6TR���Ov-Pgs�Z��$썳��HQ4�Oէ������f�����K�w w���J;�@�q))�ؔZ@����' ��xOo���xC��T/Aێ]���P{3�5�+Bh��Q�`��`�����$�����Z�e�(���I����TS�t׾�1ҿ?M���R��(�e]�����mn��^C%`%��,8��ߎ_�?Mɉ��]N�)�;t^$��	0�:g��,��(���dg$F�5kw��%�P]�(t�-n�R�s�2� �}��#�QHF�X�,{O��Š�|�'R�I����iR0�z4Ѭ����\���D�f�y��B������'@����wE����/��E����4mIP(*Xw.���%{��lė��;��v�����;K����X��f��%�K.�����*�O
0��;K��ԑ|瓬k���+�@�yh�����ϴ��a���1<.�'�_�
?�l�
��?�c�7|,�ɥ Ø�w ���=�s^G�Ca&���BX����(q�;_z[� �%��I�F%#jYw�M<��gz�y1��<B���Ţg�����b��2�v��@�p\��-Y/y4Mec���ix�޾�K�l��+�wu2^���2��H����Mcgм�'�U�)-)��u��IL��tE�wV�j]�FU$�^� U5ǄG��l�݌���p��R����A��F}�ځ���FP$����r���X�뗴���P�{n+{O�c��j����P)kb���pO߿��CP�<c�dq��`\����0�s�]�]8�%���x�u�l�v�P�l|�uJ�a(��%��|���b�j��]��n��tI�.J�!�K`j�%�S	}V���l��FL���y��IPi`��M���w�3P�E̉@�)Gy���������'%��3�VP.ޞ��J�GV>n�.m�wVa��!� L�a���,��T�#IP���o8���;:�K~���+RH����Ժ����{�����W:�H���{�zR�q`���
�ų��U'@&W2�n��ܰ|���~ny.'���?4��3���CF�$V�
c�pe�Ğ�T�� ��.3A��:ԯ�-��э%��_��H�uZ��ǆ(GA#�"FA���
�F�<��I B��k[c�N���n���p��3��Z"��kV��V�1�S(b!�蚑��F�1����#N8��J�D�����}1h8�Q��	n6�ͮ/͇�=���uU%����8��	Y��@΁