��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�%>��1(-fR�6��Oؽȏ�)���V��L����W�H靠	��*�0N#�"�z��|kVL�$�lLp�_��5	��'���%�Ƶ�"Z��ݸ�3W'r7A�Z��`�]99�����::�1vTo��/��a�#`����%J�\�=YM���42�Ο�}Ǫ�cT�c���~~_.ӎ�n��#y��	q��̾��4�d���l���}����E����֞*���
o�8�?��M��0	(pv,���y�ۉo���M� ��e�P���{+S�
��2 �&����J�� �\�HU(��JAX�@1R�P #�����0��B]��)A�7+n��r*^�92₂�N	>��x�W������-�{�/��_�X!�X�@�=b�:�0?ɒ��0w�Sc�>C����@?��,�Q�"�dX� ��+�i� Q�Jp��fp��Ͷչ̳d�`Oyy���a�$S@㤒R���UJ嚪!����G�"��6��~�d�|�AQB��u�&>ƒ*������ILn�Xp��F]&g�^q_N�B�cz�n��Ҍ)�X[���3�r��`�xΜ�:E |��wҔ4\`a�L~�k��v�#����W(�&�*j�,����N�GWi���<5�1�Z�M�"!(WNk_��T�2׺�/l����=f�"�`	[+���a�U��^��?���,bIv���n��%s����mF�n'S����{���
3��o/rI9n���SP>�R�]b���5=fv�Āc_�v(�Gs��BSMD$~�����l�(�*�~�6�3P����M+%�������Y�Z�d��\8`pfƻuk���s��1�&�S��/��\$�:}��(��[��M���M�IH};�$ع�~��]�/�OT�R�}*�<g�/�T-���|�5S:İ�tMe�(r{l�����/r㓶OEMމ�νz>.�s�s I�1�����L��1xў�/(x�%�U�3��݌Q����N{���?%ݨ'%�	���cTy�i;���o��n�7=�\*��  �.��1�5�0��Z�J0��N���4߱3�W���+W��e�@�U��9x�)�8z7�p=�wy�o��N�_j7�yqs;e�TR Eܷ��������L���u�|��%Y�mSX]���p��M�!��,�7���E-��[��bBZY=�ri������F7@��e�9�{[fVf� Q���{��-�a%ђ>����r��jN�S���s��������6G��p����/��F�Zc��"۱lg�!���%�tA0 [�l���{�� ��V�p��ns%��_�n*�`}��y�ۄ����O��Fa-��|MQ㓹C���G�Vٰ�����l*zj_��r�!�io��Bi�iv�<�x�>$�.6�2/��f���vB�l.f�����L�����h��6CcY��&�tP�E+��f5�D��fh��a�WQ�p
�_��Dw�"��3��U������S�mN
:䖠��L�y���]��T�o��
�u��C7�(@�pw)�&���'�s����ҚD�R��;2��(��Tq?>*�l���z���C���=ϻ�`Au<�G��1?������.�g���-	c��nn�?98M5zcEOޗ���t��+���D�?�y��Y�,L�҆���~�o�GԪ;�o��8I~�"��r%ǣ�փ�.�lP"_���R��������G��D�,<ɐ�V��o�=�n1����&����[�!F�Έ@�� ��2�qs��m��C(L�qZ��F�!��_*�'�<ǵ3��\�2�`�;�K��YG�����-X�7[����)m7��/a��Ǻ�%��O56~5O+��S5@
�����z���!�ΗR��?�?ZZ�͕ZG�<��yJ��g����v ��˽=y�e�*��&��G#s���\�AK� l�B;Fo9��>��c�a�t� O�,�w�=I<�"L���h#�=)T�<t��C�F�c��!���g��1}{xaN�J����k�7(G�Gw4�����?nH�}͟�.��0}����A)P�	@5�0\�UUF0w�vV����x�x"�߮2`�e�: �
+�M2%Mt.m�}b�L�q.�:��幔N}S����*"'�f��:�4��.�7�xdз��ⴉ]�0`�"PwaK�I�˛���0�0麖ao������W:�+-�6����)�53����(�,�I5���z��+ޭ�/�ع�����h([Z�/�ˋk�d~��V��V��5�Rت��c
4UL*<��>@8�^l�{p%*����M[՛�,�t��
E�6ųa8<MN�[�~F�/�aL��0�G���!�NM$����8�3��D���O �bq���^�`Y�8��"V���G�321MO�a-/P��p��?�D���i-wtlEx����<P��Rl�� ��-�8�9Y�JO�>�
���vh`��H;��K?���饱}fh�Z"k�nu�킹�h	jd��`��	+�B�Ґ=�Tӿ�j�3w�يd?h�)���+�!������	�,��/�c������#����GCTɡ�I���1��52e���uf��a$�_}�Ղ ����F�Q z��Ջ��|���B�V��������a�l�go�
;�@����_����]�QF?[��{m��}�|D�.��;�����W������la����ND���*k�E����}�k�@�^����2:��D��̳e��8�V�<���Ɲ �XC���m$>ke��-{7ԛ_e���C��j6�֌tG3%�O'�h���qTRz��6�^���4��-���k�oG3
�bT�2Z�Q��=;��S�ʍ�/f�a�"Y��������6������f�`E7U�?��tU�G���^8����{����2�&!��M]\uӰ���@15�_��胞���1�'��d�V���)K�`$�L�sf�p,B�	�{����&o.��2[�E�mB5VhU�2�Z�/�W�g��#C�|��M��?��('��H@hJX�c���>���J�G/��Zq>�7��N�L��g�˲��!�����^[��Ŭ"� Mnci�%cߍ�-%�$�ۉ��jV�R.���%0�(T݅�n�G��*,��ۊ<R��Ge5e=V��cT���K2�V����8��4��U9��bu��S:����M&��'����DX[��_FR����A����b��XF���7Z��g�Ţ���E���^�p��Wc7󂊓�A��}����q���n�b��o�R|��.�0f���7����}��t�N��tu�$������<8������Y���ȏ�$��PC���xW��_R����mh�n��q����6r�'�jf�������i��d{5C��!�K-�RVP��&��x�
:�ܬ	TZ�Xg��P�S]���	n���Ѽ�6���t��6_`	6J��y�]�P�:\�5��6(h9H��&n��	`@U+�������r�'!��C����N8�ۈl=fHL2=� ��5����	Ql��\}4P���KF=;ϯA5/n+�@�+��g'�
��%뜹��(>����y�"R���_�HQ��@���-��[Z��LSlH���w�k{�g9���F��)�Ă��������@�RS���4f~<��d`=���m*@��+ذ�� �(&3�I��$�N�6#����bqWp)��~肯���xF���p/e�&	��g<�����]�r��y����~��'!t)>��o��;ߗ��eM� �z����$�����#�����lH���[u��69ֿ�����#-z2:���GR�1�\d��΢���E���/��`Gh�3'KXM�6I�C�5�4�a,N�7�7VWr涵~�I�;9@�}1-��o-�'�c"H-�82�v�8gh/�͜�?�������F��E�,�c�0�t��}eɥ�1��LN���b���-Q���~L�w=�^�7���/��2�Ѧۄ^1�����<o�s�nS��4�����C����p�\�W�$9Ԫ[����Xe���[B�ܵ�t�+"�͢QE^��c�ZR����gZ=W��ͨ��?]��(��]��#�.8�&[��1$�}Zpr\��c	���)C��Αj{r����3�9��Uca�^M��Ã��i�utxp�i��?������yo:��=>SH4����І�Lm=�ڙ5�}�� �I�U䣀�v�w��4*�ÆA첀���k���<x�'#N	�4/��{�񪕶��?�r��%1�ף��1e��'��dC�l���+�#x�ȡ<�fKb�S�1�:ξ�/���������k� ��Nz���D \mb�=Y�i$�.�as�2"�����z":�P���	!m`x蠡���1���L���a��Ϙ��eQ�is��/�E�ό��(�m]�)"��+�s����q��{��{nտ��ea��ÈlER��޾N\�n>�Cpj��|����0��2�op�����q��.����`���ͨ���	׶��7˅�t��-H/b�8+mE.�4kLH�K��[����,?��єy�ٔ�����F6(+�_�����㬢���5El�f�Nz�l�����Y�q;]?E�?�:qA!�R�HV���#3��X�	���[��S���V�+���%.ZF�^��P�4؅`�t��J���/��$_I��y9������ȑ����޴6�Yeu���� ����Jd��+��� �b���֮����vmp��s'���T���\&p�#������~��'g��6��h-�9�Su�k�o�Xؿ!ǵ}����S�R��TP���+�����!P=E\�.(*�:�-�.�/@�8
T��xw����k��Ϩ�]��]=d��Qӱ�A2󍧀�.�A�ɕ������&[+�3Y�ά	�Y!/�fe�yn��p��k�E�(�׮]b�4͒��%/�a3����yJ���&e�dF٭=v�����:��/��7[��0E(�c6;�[�c�hP�4K�`^r��d��$20�M�M��������6ɥ/s"�� �����{�Xj��ؤx�����k�H ���㭳���ϴ@�p��?ֿ����3�錈Q�3�) J��1cur	=����`�?!fK����3��8�	�h�2e���k��ul�z��Q_�)�V/R�q)i��RM�[{ͣt4�����OZ�a�	�
�З���)�+�-��H��*y-B�����J��M�⅂5��"]T���E��B�r[P}ӷp�*�HRL����Դ�$����1ݣ��&����F]3��N��c$˻��	Zq�=�b�F�<��KI���t%dG��:/5��R�RX������WFLk~~�dآ[��I���ϙ
��)�%����٤-��=?�IkN�mA^&�M;���Feڏ����A���(B�g
':k��X��fOw�-�w:i�q��ը���g�y6ug/���͑g6�ҢjRL��.vl-j���~6�/�ڐ]&�3"N9���ƖJ���euF����Z��� 