��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<�؝����ɂ<������!R���kc��azZ�DQ
O"��� ��Y�u�-T9tg�"�l���|�8���n���7��3&�����9"�v��tk?�u�{��U�4��\�,�F3�	��0]%�}wz�k�0�IBv�DyA������=�Ӊ�Jrm��}^TcR$9�B�6�5��ѹ��w���W�8t��3/u�L�vpP7Ͼ�\o�j:j�/��1�J�$�! �G�v��mm%g�ū��$�W�-�S:wXZ�57m��d
T�[��,3�K#g�,zf1N<b���_��
�������V��x�{3�qȡ��&��|� 1(���跪a�U�Ma��U�s��_�i��B{�l�$���(ݢ]�]�42�?�t�Ie=%Ԙ�Wj�=�����zx#�e�
F��>*��J	^.cY�����VW0b�-��Gː~��:&��B�W?#J�ki6���wL�%�}��;��"�5��*�3JA���W?K�9q���]������}�
���M�n��C팉������T#��π���=r�}rL�����>��pr������o�E}P[='�V|L�&FR'%i��]:�wȖ�y�؂�k�}i�՚<�ʏ����g�լ>D�yA�� B�bi�^&��$�D�cx���]���)�e_\e����G�|������?�Iu=��R43>��J}�s�~�P���	�0��,?U��յ|vy�`.��q�q�d�0L��U�q��^Vvh�0p�l�;2Q�1`�e|���_ܛ�����t���.+�x6�LiI�>��5�*d��[|��O�5�%re���H꿇�B7
������kO�K-Ld�{>�Rl5��ð.���H��˦L�~���RF��z�^`�su��љ��'�1������}��|��5�.%і� �X����x��TdKSXP�̩����|Sjy�~�~<�w�?��ى(���i8�Yt^-Ï&PP����-����d��P�8f{T����TI�(m��LA�7�Ȃ�[������D�SI�fQ�ą1g%47��7��Tl��@�� J���ý�^������r糵�[�$U��}n�-�S��b4��&�����ZX�?|�v�1A�%i?O���&'~*�R���ÄmM���N�xy1w�;Q:A=�P����qumV�8A�c�+@�EI��y� ��qy�#k��c�!잆Bu-�T�����yA��OZ�G�� �o\G�W[�G�M�Բ���Z�A��"i��O�	�)��ZPL��D$R�������#��F��V�J��ڝ�j�m��3pm5�v����U]f�3�w�.z��X�!6o��Y�`�����1����o��"m�ffJ�w�� �_?���8�>Z蕎�,����	D�<[g��#�c�:�h�g�h��}�����(Mf� �~� ������~��Ox���2Fė#��d5���2F�|X���*P}9���
�OEx7��h��]v���Vgǚ��=o\#�xżH�Q�+/R���`Wz���0ƻHst��Y�$�)̯�iN���"sY��v�ǥ{�o���������J��Q����>պp�aG�"c4���wh�m�)9�8�൵x��\FL�j#�c�M�X����ٟ�]���9�q���&��?��ya�����X%ר��A���4�� �������Y)4h���k	�p�~JE4ۜд@�A�#$7Hl���X��g�H��u��S�vxfb�D�L��Ɂ�j�����Ȳ���I�[.�R�w8�r�'n0�O�M}AF�������i��Ϥx'�DΠ�Z;��
��G�Oa��F���-7�Hkb:MX·#�f$�Y�P0�v�{I���e���γZ��9�_�tQ {���@� �T��s���لA,M f� ���+g=�ˤ��m(Clwm0�.����4,���k��b���_M���7�����i`���)�"�ߟP��Q24Jl�(��?w�;f(�k��
��(��[lI��ir;HD�:r��׸'O� ��N�,���5i
�t�ujf�s7�Yv&���g����_����֣��)�_�gd��m�6�P]��o}�.(��Ֆ�,)�ƀ
�Hj=�T���(����wu�^_���q��ēnҥ+���[�4zQJ[��f�h��y��;��>�����Â���ζ��6�F�qu��y�C���x��M:BRR�G;?� kP���{XJS���Rҋv�d�n�����n
�Һٺw~F�`"nU����� � Tj��+tbA���R���7nB�b�ð]=�te�Z���/#P]���t5{������g#C�/	p&���h�_ ����N�.J���J�@�W�Q�VD��m�VH���Џ�4�hoc�c7����$����ۚ_'�_��&���n�S 2����\4�lH�q
�C]]�p���y�y�_W�u�1��60�%.O��Z�8q�PS^]دN���x���֮:��W�������X��h�l6e��3\�,��Ω�e&�	yr�T��u=�Ã�J�ř���Oҡ� �.ȡ��p����F-$�/ %��K �c��0U�Kn��gY���8���������󡸠u��:N��0���X�@��u�e�.���=���f�x|_B������KJ�J��'=���&�Z����NYp�+���#�]�jLx��k!����9`��Qi�^�;Rs>���Ub��*?�������z&�M��v�#�Ñ6�c�!�ر��T�}g5Ole�,L��D�~�͙�sy��,�H�y�h݁��f�5D:��WS(��J�@l���U@\,���&�i��Ҳn��Yu�[;��NiA7fti��KN�=��Tx�	��K��`J�x����!��R�Y�+��k|�kT��}�O�w�Bs��U�)�ΧI�^�]�'9�JɊ�0����Mf�:�k�Tk\���e5�w�ۍh�(��Hˤx��&���آ㠍�1]��8̱�9N����V�8@Tlk��ķ���xӃ ����y#b@����&�}���E�%Zr���2
Q����q�wE�J�c��"P����|���o���%7А����@�.ܴ���&X{�N�xau�̷��j�ϡ��pe*_ZL�[C(��N���;�v^�c0d�Ñ�zg)cdzH�7=�3O�J��e�M�;#�a@�ٍC@���Q����A��h^9F��VYu�V(�DVUv�.6Oj�f]�FcA!��ŨwXg^�4V)c�1P �L���U�u��Ia懿o�Dta;W$��ղ�����/���psت��!�I�+_��_Aב��"���H�p�LU�W��,8�	$�N�(�vT�@FZň}�Z�
S�o�Ȗ9]�C��2�Jv\���@����"�Ն�w���Ȯ}!J�4�4�$�wļ'Pu�]=\�|C�gc�|�NW�I�a@d�1d� Ba}8�.�d�~�vB����BF�d��n��`���ܠ�x2�2?Vm@�ӽ���U��ޭ{�a���>��Lfm���\��5fT�,+�ei�X]����h����p���w�r�Z�q��������2s�UѾ&#�R�Fr�K\QkH$�䙌/�nP�3=�e��J~�?NM�_B� y]m����c�`񴇂�"����"�aP{ӓ�����Տо�SVj�o^/=�����W�~a'�Ǝ�26����-*0�~�V�|�>ש8,���*���/��n3ԖCQ</��@L���}����ه^N%�&-V/o��Y��3x>��s�<c�T
�-V�ݳU���5 �PP�?�N.�����B��q3�ш;a�*@ݿ���Wѫ׎o�k{�j�����R[��g�VF�1&|���>2J�O�gY�Ƕ���7�<?��+�fn0ɂ�]-��y�-�*-���lՙG��T9��ln��|EL��8)wY_
|Ue^�g�)]܊�ﶶDs����@m'pu_�eWy����:�y��2�œ��ʬ��
��!���^�������UO][�&�;?-|z!�h{G�؏L����ƍ<��Y��B��eF)��=@P#�cP(~kg��<T��kn���TS���V�W�]�p�0���-Q'� ���_��Բ� �j���^�s�C(&�&���B�-Sd{C���|!�o����=0s�jkŅ�yk�(I�:u��P{J�``)�c��)HE)�����vER~i��sNf�p�6�h5�o��'J;��8�P4-[f����z�����PmIa�/����!\4��H\���q�k~'��j�`��> G�8��ز^[�F�͌�V��I����[v��ȡkKP@"k�� �V��'n��L��On�Zȑ�N�ڷ�ɚ�8ں��sRJ#�VF�}��&�1S3�֗�q��aVk�:φQ��p�a_�+����#<�sꠀ�^��c����ڶ�b���H�n��kZI;�+�/�zrr��J��@��ȷ�vd.����"�*�諾OuS,-�g���X(0��-dNbL��ޫ�]���P��:��L��ߒ�vG��f^�8�ϻ2��j��q��S�	e.ږg�Z�t��oS����a	��.j�:ɹq��,���@�n�Y��,/���
O_%�1��ȣ�z�dY
+6�� ���}w\t���,[�Q�5j!�<}\0��p��8�g
&ߌN��yzA�s�Z�Jbaۂ1_7��W�7�5;�T��=��q?��Q��<�K�4�o0=jT��UbZ-ZH	�I��vD��BN�&�눴�-����
���=�����	�.X�^��O��,N���Y�nI�
��RU!��y���$o�_��4Jw�h�;%GK�q��0�fpE���\MR�%��.� 0�r�1��g�u Pd/߼ɩT��"7	��$��(��\���6:��%��qv&DiL�Q�w�Eځl`jd��I�����޹#C�))3��@��;]EG>�

X�9�4��2���T�kb&�cS-����� �ݸ3��_�q��/3ܛMb���?��5'c*��xvG��I+��oYcN;�{�,�L�}5)�HB�~����x:r�BX��~��Γ�L��0������nMK�}����{%Y��#s��O�,q�T��D~w���b�"�����J`�0�Zx�r�0�n�L�����:W�GPg[$M�V.�KĄ��~�|� ��E��-֤Vi����Q�M5;ɱ�u��ȈSgnq>Ń'�*�Mvv�H|]�����@(�Cԅ�� x�gkWkc�����lۡb�s>�6B�'��Ai:���:��rSӰ�7�D��X�ʦ�C�a��vtX�H#���<��V�����Ѥ"@�D�֝�� ̗)��Q$���XR�D�h��!��Pu<QӲ���sB�A5�)ž~`:��y���$4��z���R��[]��]((�pK蚒� ��޾� @$G��ޖk&_f��q�h=���y8_�;�,�J}m6R
�!�Ŋ@�^�I"�#Sٗ�/#�+	ވ���e�8-�����$z�!sDd[y�ʓ�j���D��
~�9�tP}��}��-x��ѽp�
�����N��m$ӱ{;��[����9�f��n������`D�]ߋXa��̰sDb`�A2���&�:�o��w�H<4�,��r��
N�a��@Қ�T�Y&��+��`�w��a����'�-s`����:�iTz�j�SbgJ�җ��rxIF�eT���-�s���{90e�$�P8.�"�}y��+�o�i &���f�u���ܽ �,��CUܔJ�8q�L��v�����9T�|��l�k��o��k�]$�_G��c5Bzg�en����7�y�V�=�&�ul*a�&�w��۽ ��&�E;��W� ��C��δ!]��!2V�-�F5�:}Tļ`����+o�wXM��[��n���?�1���XoJ��h}#Q%&��9�� �l���8�+5ű�O#�l�}f��^N@5��GM����~�b/ӻ����$ӨVvR7'�gɷR��p\���>�/�㘓�{Q��XA^��BtK|N,����kDK0CV|�I��p�����*b<�K��-�iCpɞ�=�$����I	A�HNRP��n���`5T렺adR�y2���%i���Y7�A]=�{�đ2��a�� , �H{�n,	S�K�Sȗ����󶓸l5���	�5F���|�Γ�&1��h>��3Iτ⑸�+��.�a�P>�J9�Z�ci�c��n"�e���j��6��i������P#�b�����Q���]B�*�o]P�2�q���V\��/^հ�>�?
�@œ:�/[҂��/���f>V��g6BA*/�4V���l�a�/���Q��Q�8jݩ�y�s5���MdC�"�P���Q<�Q!���V#�βD��%Y,����|�)�S�V$���v86X�1�J^�{�?6�F� ��E7����a+`�L����ӐN�vU��5?j��	/�Y�Z�D�{g�U������
B$\�L�$�}���&Nι��7��قS�h��Q_�m�ǩ�Ļ�xǞ�9m6�ΰ{?����[��t��'o(!+S%����� �"���I�%�X��ܛt��<�c���i�ޙ�Q�.�.'ʂ!~]������#�$��}}Սe�j��5 /�O� �&�֋i5�U��Z��q�A�ǒE�Z)�g��F�y-�LJ͠��^�s�}2+�L���Ŗ.���<v[��a��;�r8 /h����=l� ;�T��R#�nd䕯��������B1߿s����u�,L�V{	K	�,<Pah���/,˘%�A'(r2�1,~�����~{YM\��DĀ��i���]�1�{J�w������ӎǳ6�d��h�)�b훿{�V�	N8��?ɀ>�	�\�7�)Qg�Tv��⏗�k �?D�`ܡ���{���/*�@�\�חm�EG��2�H,%4�t�I>���g�	w���l����=��{�>����78��#2cg��d֭��6�6&��we�.�t����7C3r�W�E<��w��kŇ�mS��:�y��k���vna�D2m�98�x��)c��pV#~.WX×��ȑ@�úx�-�����`��7������	�O@��c y|>\;B�T����%~2_� ǎm�K�����_㜰�l�(��0�8ڥ>�V>�f@m��>K<ޘ㭹��
���<v�2.�sf�E��#��������V@���������X�TQSؽ��IaqD��,�i*�����i@$8(W��48[� ���l���^���(_��Tl-�aI^ ���L���3
��l��$�aH�x�"6�D>!j��I�]�]��-��o�C~�(�~��Am#�ٗ�"��n���T��b�dF"�t98Z���d�4ٶhF%�Fӳ��L���j��ӊ�[��D�N����j��Ǎ�z���y���yӅ^���B��bЬ��*�a�T���{�5@��½ß�`���aEum,f�[�>�������Dw�TZB��)��j��P���Isl 0?H-���,Xhp��^�ω���J-��U�����d��Uu�jks�v�h<ּ�h4����G�U�3[��?�&�tJX���)]��!X���{J�����.EU9����~<x-��"�Rt�����G�`�ɟ�k����'	�H}[{�[���"��p�FF-�I���&߁�r!c��ur��i����!��L��R6���c� �U� \	y�B!�S���Ĵ��A_���q��5�*�2ݲp��d��Z�Q�a��݀�L���8s�@�&W��9y��W�z��ߊ�02]�Yy^�0����Ԅ+E��?&l�	��[�.Q���?����18�I=���.�~���v�����F}-�t{����Z�X���5�<[�sOk���L���0��#�3��)�A�O���?�n�O�~�üio���>��Z�jK%;�e;��^��h�ە��tBH^Ǔ7� ��w�r�߯|�ʕ ���i���F>d���yA�}�%d�Njr���{�U��4��#�*� A�i������u��[��"O��oc�1���l���%8��G<�S@�攄t�'o�ߣ���ZE�ڷ�6u�c�����������]`�&�DH��Ä�p )����z`V���޴VawE-���4'&�#����tE(b8��S5N%'p&*2rU�se�D���чk�|V�Gni���y�3B@4�~V��gNB�,����W�����7�7Ӎ���7<t�����l����Ea��wSW7�`i7��;>
�B3�����&%����O"���e�OI!�f@���#��Y������'�=�~Ͼ
i\͝���I��t#�æ�R�?���VfAUP�!l?a��0Vb?y\l�:�mr�`�� ���T0��,L�� 𜊠g?�@�s=� �lnў����Z��/;9
�`sC�@:X���';��83u�ܜh/���[��с�q�z*�C	"�Ⱥ��:U�GӘզJϝf��$�!~�_�츣,Y�M��T���J/�E�x�eBfo���=������!�OgBb��mc�ܺ#�O����l4I�B~�x��[4���v̻��ull:�w�-�4�Q�*88�R�Gev5������2X.��IM�%k/�-r�O�g��g�q�L1�'
]��>!}�N	��V�`&͡���Ũ�^'���$�b:A�vA���Ԉ��j�7�w�%������U�+H܂�<b�۩��n�@�=q�5�в�L�F6���/�6��p	�"�N��������ٺ�T}�E��t�Bg�QdI����f.�P��ⰖBd���q_��3f�$��"y�̡�Ʃ��D_7��"k�;Y$��e�a-�U�������{��L�lR^�����IJ���s�t��ؙ���)��D�q�n���~��{ge�P�bx�u�l9z�d�J,�뷐��|�I�o�Ne��hm\�`�J�ô�AT�!�0�D��֭!�[�p' )H&�R!2�rUh��Cv��LƩ3ܳy�~�p���F<����X49�LW(˅�oeᏮ�9 ���� 6ޢs�Tjda��7��	�Y��<� "�R�?�	���$q�~��F:����<o�Nډ��p:��R���~~��.U��o��т��G��MҬb�tjgY��jя�pMk+c��hI�)���%����%K����t�R���Q����
����Gw�4i�v�a+ҾA
\��E��n��~>1
�=�����	��I�e�D�^�s�4d*qzy=	u���P��ˈO��w�D8N�(��VPɵ��UN�F>�a���B��Z���`���EUm1���]f�`�۟l��)����̔�ض|I���f�3��:�R	�2���w�n�?���'����o�����rЗ����.�#Rg6���)Z�Z�:S�7��*Q�r���l�����:$F��Y>�+��v��̻�u̓JGK�|h����;�S����#�V��mD���Ю�5�̩4vi�5pl���	�Ou��@�f�0ӓkt2�̚�Q4U��_ǯ�E�����:(��&��.��_S��^LڡJ*�*{��g��W�k
5���Ov��3���d��Q\EU��e��[�^O�cBq����
e�m�)R����9Y'G}j��@ �̺�e��/֤ġ��&��~��d���8eҁE��2���\NY���FEl��_���w��6	������4����o��.�l�a�E� �|�C�Z�IM��WdO�K����){���.h�ހ���}| $p�Rg ��_
�j��Z���ZRYp.���6����0�xV������ki�J�L�dÁ���#J����٥��A]� :v޸���JQF]j,���,C�K�'q;ٝ%�dZ� /��
̏���9�C�>l�S�����.�;|8�6ZP�J�u�ZK3�R�WΨ!D՘�=�k��f�:1�(���[����sX��%Š13s��`���h����&�����2�5@�!1���+��Iͅ\��]aG�*g�P&���r��;6��Kȉ!>�9�L���-�?�u�}9�ZjƗc�g�A����B�[f��H���[e���3$�T�蚏�h4aq`����߃T��L��Jy�nwQ�MQ�6�������>��`H���O@7y���d�C{7�T ������fDy�1��D鲺Nr�K1K)��d�Z�:ބ��q=X�K���Wu��R�%�ހ�m��IȬ3�G�0�CVȧ�M��P��+`�{XE��Fl~mkQSDR1R/=MP0M??2�{]V��ý{���'���o�)� ��e}!4_�]�� ��G���x�����C��7r��������bAy�0x{����A���lmXj��SQ���k׼�R
��}<~cKG8�,���t����M�,�cM���l����aJ�:]�����)#���9o-?��n8�҃϶IH�
����Ft[(�(?<3�ͺ[v�f��ONR�5�]�#pf�R��]��3 V؛�'�V�̉M���UhL�C�:��0 ڲ���D7��e���q��P3����U���
7P-}�C.n���ʕ+y`���+�����q��d��Q�^�����-م���IPq�@mq��?�[l��a�����1��q]�����M)���b������6��7���K	5�0ET0����>R4��Y�6؀����6��*�+/��	����:�=ہ����B�ɫ �����sQ_f�<D��x��.w�Ba�"�1M˙�&��&o\�ee7ClD��Ս�@�7��]�q�,kE��������7擊I��0zYf���9� jץ���v�J�bC��~@|��D�����"������w�HP)(a���.ﳎV��F�Q��^Ub����K�5sЂ���o{-�p�/�Pcq��P,�������yRi���RI87WV�Q��$�e��CQ���gW1�N�(	-T�$�
:^<�sa̄�3O��ďWQ��!�� �%&�L�]�f�-m}�賾��l��ٮQ�n[�+qy)�!��B���I���nm����=�5�`y��O.-��*Y|?�����F�%o��Bk�F}��Lf��+�dUl�����+���-�|�faͲ׭cc�C�٫_̇��|!�V�M�{^������ t�P�%�2�!�8z��ʱ�*�e3��7M�imh�ޘ�rOvpv�b�e��94�J�JRBw�L.!<��j���Il胀��]y{{Z�rջ��cP_nWI��Z|��<~�*�zI*7R��Z��	G�a�4(z�PG9�2.��WP��+�k�ڳU��E��vGI��o��k�f�'��d@-\tpq2����G-�R�͵�.<v�d�a�0V���dr�P��AX4��ڮ$��� ��c�F���@����_06��~�Zܳ���8�NQ�iK6#E�M]��O��4�S}2_��3/��8f/���nϾOg��<՟�����X�;I?aa�2O���v�z�P�q`��5U��˯����t����n�y�I�d��0&�ՋI6O�h��uHB�OA �v6��G�KR&=j�h')��
��������V
�������~ S�C��<�r_�6l܌ǻTX���}�BB��x�M9��v�.A��Z�����Dc�u��rz��*G�x\�}G��I�A��[�o�yezX�����oDd�aa7.P2pLy��� �K��n
f���вU�)�����h�m|�m�36K֘d����96����^��.ն~g��P,�u�8�-���PK.��w��&���淯a�r�[���W���h�s�=�!��	��q L�X�e4�yǾVq�9uW�z������C�iC���,Bo>T[��5�=sm���[}ffA��� ��Ub��`��(h���������7�1�L14��X�ٕO�dy��L4.���<��ʮ6�Ht	��1	yo��%i3��>G��W��~^��85�c�Qߐ�~�׏�Mw��F�9�z�X��{*�m`/�3فȴ�����	��3�vڿ�#xpO�W~�p�����&�\���!�"#dy���fS.AHBM�*����������W��尚��?�K�y>_�AmRW���i��b�5�kC�`'QL���Ǭ̧D��Ҭo h��A��b��	d%���O�0A+U�8"�f����е$�N�-�{p�X�=��Y(@0�7{�'�E%l�[�@����ꎹ�T�*C��H�d��~;lf� �z6<��L=��Ʉ�y�+����G����N�����g�;c��H���"���OF#�-�f�P͐H��{&?V6�:}��_����~��w���ݖi?�G���!��uڜ*�3�y1}��~se}��#�Ƚ�4c
f�[��V����<\�������d�n�F��2�r{'��u��)>�dk�K[��o�,|)b�VR��Qy���Ώ�7V�5��6�W� �L��lO����S�l&�ܸC�O]��5f�z���w�.GӁJZ���	^����t�[j|8PRb!�m�0R ���M��p����AS{&R����'\	�4�\���@��H��m�����i�a�/�h��	'�c`o]� jL��Wk�N7&��v�Y[m�����"\�}@��!���Y�h<�N#�fi��d3��գן���t��"ܢ�ݨL����U�\V=��q&ʣ�F`ZJ�L�2�fB�����\=3�	���A�e�:��S�*w�]Ҝ�S>ؤU�˟L�ߗJ.X5���$O����+O�֍���7��w������i;�`Mǘ��}�h,e�uj*7CvR��vt������y�����$ñFL�p<��1�I�4Rf&�^���B��N���E�,���yI^,���I� ����MZą��gP��6��F*���cS�A)A��\v�x�;ߜ�!�hٺ³�8���g E\V[ʥ�J��炮I4mG�5��	��uS��n2ъV�Q���B��0�F��.zV�2Q�� m��@�;�¼����6���v�k��5��#F"�[#0��������9EJ���G;Øu�~�3%���JFѳ".(�ǹ�7�!�9�a�TF]\�f�w#��\8'X �r����
�&ۀ�h��
�U��.�o�f�]k�Ǝ
/�E㱑)�� Ib�=i8��S��e	I�5YX�:f�I�hc���C���g�.�ao_���)����:$nh��[W���&�~���(hD(���@�m�'��9 �eζz��Q��
t56wZ�$�k�v0��A�Z'P���M&�2�ޞ}�}~����3��g#E���>2*	�sWh���M#3!,�P��-QUo�N3��tB�_E%򝈁�(:;�r�4��/$y|��9{4���%J����"Z��Z R���:OṚ��ћ/)��J۶�8�\.	���[i�}��87*&�S��4.yW����03�_c�u�T[S�P�Q|o���c銸�9p�1��,W��q��@��D�� ȫsA*V?��x����R�|��dG_)�r��+b�r�疐�*Z��X8�T���:�g*��?� �F�5�/UmUS��J}���xӿT8��X�!��
=;��4V�c�B����,�[m�}F퐺7� �s!o��;�D����pI���o��bZ]�e>��H���J���������G�+s_ܔu�����r��cvwɧ���x1'G7�	��\3ٵ֥���qip�ꝙ���,�Y�qmf�*٦�n�F�����q�L�w��I?�oDp&��c�鞀���
|+���|z#�0�aSm�4���2�%X�xm� ��t�RA������燱��T�o�����^%6��I�]�'�)�a4���F{�U2E�Mв�J�.x�j�,�,D��b�í3�y������\���rj��7�2���ȅ�����n$i�$(xX��=���VD��a3�:N����@��e�Os��>�����/�0l��f So���m������!�<��x��J>F1�M��Q��Ҁ�?ձ�n��a�%�}�^�����! KAwSz	n�䚾S�8���x�j L�`a�ԭȄ΄�����fx UK9�#B�Z ���M0�6-~c֛d��S1��K�_4���R����z�K��(�-/����/^c� �ǡ���t���c�iT���g65���ڛ����)ޝ��@�P���me����<���TNy�.`��l�r\�cw��*��C_�Y%�1�a���242��Q�S�=�^�AE��|K�z��؀�j�$`D��x�*�&�n�W�0O_ӥo��<�����Z�g�hߥNN��n;�ʂU�ʁ=����[�aQ�U�BM�E.qt���m�8x���翄&�����w@X6�����C�5��
]y��Yd��;A����{��\��d��QCi�/B��7�8"�2�����ק�Q�z� $J��	T�_t	qO(*h�MF�(S�䭰�����y�MD�n��Q�bM�y; )���}��` ��+�yV�9�3�S �z%�R0��Fe�!,�kuPJ���֠�"���ɾg��t�dEVA6u.'�G�����S��K]�x��z���Z��Pǀcƽ(`���E�i�E��i��^�6�	�2<�б�Β	�r��i�bt��I���ҁ��uV�� ��(r�� �O�9�r1���od�T�9����Bk@a8��-�S&Z�L�C�� �rIJ�P��4�xD@h�=Oᜉ	�.�k8��^ˢ�xD_�1��#�KJ�o�����H�6�ˉq\���3p�ϑ�$�׌�SB\X̸��]HRC;���Y�����@#,�:�d/L}|�+��m}��ZS�\�f��p� �Z�q���$�9X�N�L���HZ��(�� ���V��U���G��h�8E�����l��d�
Dd�,��yC�⬰�ͳ�1*���A����O9yp����S�f���rɵ�ޛ�����5�p�C�,�f��e�^A�{=�}�D�vʩ����(�=��?��bq�
��ab�x���e�h����<��놬�����-���_���y&t��	�Thf��ɘ6?�h�3	�8�e����/�qd]�is�*��
�ᦘV!����_�z}M�!x�=�����`@���5:͂K�9��&��nC�s+�L0����mi��ـ���щ������q{��1/.�ڿT�۸�؛]:T�u���g&'�����>�,tyi��/�գ�n_�~���T�z�wL�Y��g����$l������ `��M��"Zq��z�;��������Z!s�PD