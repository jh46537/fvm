��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{�8����dOɁG=槆d��;U�4X*)=��9��� �>�J��e'�G�׭X�1���u�x ��L�HH�un��D��(���_���?�j @���2=����7ԉ�R��i�Bx��;�~9�xP�+�ٶ�3�<��Yh�t4s�$�'X�St1�B��u�uwG@5\�.B��w,ɧO��E(��uȶ��*ZP�8@�rͲۣz�t�Vz��oIS����@+��_$�U��m�`��I'M��������%bR?������B�u!0�	9��(��S�ph��<<t�G-����g�?%��'o_B�0,mF���Z�WB��x��h��&�Wtn���$>�r�H޿;H���,��$�ʫ�]\R��7�Ep,�rp�a��U�ڝ=����6��������cZ���ck��j�RMpH���yp��C�ח��S��k��hl��@�W���W«z`�@Đ/G7�S�J=����!0%�i��!�W���S�5��¶�fu���H����,]�N{���]�(�v�ѩ�	���cA�+b�x������ f-��Ϻ�8)�"z����B�CXN�B	��p3�_C?F����f�TG�>�c���R�Љk�
���%�7�Ao��$neM!��@/ajb�=N�|.��c+Y;�c�7`�%�v>��������WK�y��������g{aak4麴Q��렎ƻx�I����F���s;rVzt�|�k)�������w�|A�*���r/M���"A�8�Gš@�2ؕ��u�+$\�)mx;	G�_@�&�«0e���J0>ݒ����:V�%�~�H=ң��������N���N>�pխ�����-v���1�v�b�]�Ӭ���$ѷH3���J��<�y��ȼ���]����c�(�[!�X�8( G=�"A��ed��lz��V�H�^���r�Dc�u_�9)i�J��%e�z�a��UX���K�����+���3WT�j�sl�����k��!jJx��o��ۂ����JB_<���S�O��@�=r�x�QmJ**)嵭{赭���8N=3[�2����Q2�E�8�����������*%"2��9�~q���FZ*�^�Q�C�ư�߰v����Jɻ�ǫ�L���y���~ �(���D%�k�|)�\�z�#���V�4p�aH�ʇ�<����Q��'�L(��̃��a܅�r����C L`�U�5+����A��	��UqE�1��֧�B���D%H��E�/������8¥��'���a�2�:'�j�9�*��ٰ�<T�g}E�Id��˕?)w�mb���;sUmC�]�S�^V��:���/e��G�NNp"��J"� G`3>�6��'~�\*��=2.MQ�����ZV�: �
*��qH��)Hd�-��r�p��8��)ƃ�[�7�g+ ��w�tx�{Q��[SW�����ʪs����R��A�8�3���ҹ��t<"���x/4�|\��;`�lɑ���:�ڎb��V�'3E;F}������L9���(s�<��L�n��p�.�<Ƃ[�����ۻ�,�,�Ȯ�Ϧ3�F5qM�BE�K��d���+oD��GU��P��2�Q�"�{E�h�@n�����O
��Y��Њ�c/�ئ�z�--�$�-9��񭚙�s+��A�s�'��QV��/��sraa�9>��H�b$1��pF\��~�R�4N�ց�&o���K�� T��K���4�2)�%z`����x�Vo����_���t2��1��H��L��u�1p���Ȓ|�+�s6�F�l�l}�4�A��ǜ ^I-н�\��E;��7�������G�`�B�?�T���x@I��l�:֖�\����� hh�};���<��7�@O"߿�OV��}�L-wqtu臭������0i��z��b�x@Α��K;		��﫾��q �oْtgp��{F)������S�R��n��b���%�~rtMw-��G�CIy=U�dNw��W��J�����	Lܻ�Z�~R�<�Wڭ��I/~��w�����_)�'�m�f0�!e>��@,�IY"��-��2� G��]F�[B���Nb���鱙��Ǵre�\#C�Ք�"ڛ��MF��#Z
����l�H�y�*��e�o)�pE�͡>���F���BQ��ȼ-���<�{4ʘ�X��>e�UB�6dtߒ��(|W!�iG��I� -ѽR����*\���\���8Б3�R|�|<9��b�n�|޽�S&c����g����(7Vn&��N�v4a �6��B.�Ҡ�U]�:Yb1���R��C�G
Æ<�&��O�Z�����l�B����J`@�p�d��f[ǝ,D{I��g'�t�C�Y%�l�=��1jI�y'7ѥ���@1���B1��og(�Vme�u��hނ�S+]��v]�j�_2��ʔ�����b�8��8F?D�/�a_?"�a'N�*� AOC��4|6 �Z�~��(��/�ŏ&�ȰzN,�5�@{��# �$��-緕.�����[�����5��!�U��}����/��'�|�ۈ�@e�æ�t#-j����Z�����B���N��n��b�,�<�?�J6��vx6�m���� 
���m1��>3"S}ۅ_�M����d���-C,M�nQnmIe��#s�Y�9C�w���4�Y(v����3n��@R[��L��G�AD���?�DR?
��W�GFy�宿��=0/l��nS����'��$V����.�Xt1�Q�?Xp~t�����1Lbj4�}{n�JV��z�Bir|��&IO�?�pD��.ۚ;�Z�t�|�F�N�����U:D+�Ǜ4�('<���]�u�p"�Ό��2�Ͷ��.�P_��v��vG�XP�NB�G��/U��羽�Bml����tx9�y�F�S�Y62�#�����(No�4%��{�Nީ�����a�`�&��@�ݟp5ZЈ�3�!��Ŭv�C�F����>/�����cK��򤕽oPj:��
�^	'sn֫�H���TV4�O
ej:����E��?e&���Q�Ѓ�I�Ф��~�&��T,�R��3γ<�ki�`_Y����2���m;�,�׷a*o��?���|�cE�K�����'��_�/xC���@���hS5s����4�Fܤ{��pzh����^q���{q�	D��W�=�������mJeTL֔6���"�"몑�T���.`���6��ˆ��Z{��{Y����	E�S����p,��M�+�8����g�bJ�w!/�~$[q��m^Ӿ�)�t�۪�9[��PY������tjl��>������ؒ���`oe��v"����!���Oڈ΢y%K�4DL�?+��poɊ������t��H-�mxp	+2i�_��:J��q?3��cG ��j�CK�� �85���\94^3��B�<�~�Lo��g�4��Zi��?��kt�K�x�{��"���p����ht��=LJa�g5_>�i]w��޺��#����(r��[�7ͬ����� e'��yA.��l�����O�=�`h8����+�R���1-�|Le�1Hުy�o]g.��?��o��#�)!S-~;���.��j��p���ѣ���z����w@�[�����Ζ���8?'-}�{�[ ^��6�x�,��PnN̳ý9i�&�X��gc�/�ΑnC"!��۴գ8C���;jV>�/�,����w�W9����R���L�yWl���.s�����5h#E=��I��"�p�<��p	�%`֬��tm�(/�t�0���G	�|�@�u�|V<̯#D5RAV�2���t�/y�'�"yP�����-���OX�L���N��C듖�o�L�6����%�aL��%n�qML��p�x�	an晉�i��OM�!�դg��$Œ_~����/h����"�1�d�Y�*��u%�%/X�ւDlI����O&��]#� �>]D���GRkm4ۺo���e ?3Fz��w��V�Y�7I3�N���^��3�P���s��SD����s�˙�!s�x���|�'$�g��!��c��+�tR�d]~���F�y˄(Jx����6�ci}�p������'Dϴ��	 B$��Qի�h�^��,+���9��٤��d_�%@)�Ž�ðV��[A��y�Ô����:1?!F>#)�����\���ʤ��
�ֺHW�BJ�*���K���q�%?A5YI�e,>h��n�"��GXs���0��Q��t6�/q ��l��rek�'�XfԹ�[�K4l&�tXA�)�}b:w/�1x�U��/�<���1Z�l�#�BR�����F�:��}3�J�z��l2��'���ל��F�aZ^�*�Yw�#ߊ��e)�2��=�gB�ɇ
�$�p�`�0�����>	�Æ�@=�k�����Qvj��)y.@�bG�(�kc)^�[^���a����!F�J��m��N��#0�,=��WI��r<����ީĩ]��_��0!�B� �j�bO�j玈\�	��A窑���$9F΄N�HF�5��&jPP�w�PO�U�Ϸ�ԃ3�P�ߘ���Y�'۽^'�ż��#p��s�z���Zm(ז�
I>��߱z��/.R�^�~�VA�0�`�xo�<��+�݀W�k�J��E�� ��FD��8������ˈx�
,�"�wz�F����,��B.�Zw�Hg���a����i�*+�~=ͱ�J
a��x�qG���0 ɥ�^���O��ZZ�`��z/���Q�an$e8�kf�����z���4��Z�㺴n�r)�����Y Aȕ�V9���<�|;��Y�.i��P�5Q��Ԓ�"�({`[�4�)	�lm����v�d&������0J���~aW ����j.���ۖ�E����\�v��X�$�����sW�'a�|�c�m�_��\��1��b���P뀗�*N-5�,t vQ'�$�Ey^/_���|�ZT��^ϔ{�
���Z�R5Jsq���b�*��U�ǖ��!�"m"F�v���b��%Q����?q\Z�:��
����0�93�`q�<�w��EN7N
��)��Y9W��[����2�W�y�W��K�����#}9��BQcP�_S0�`[�h�bٙ����_���Wn@1Ŧ[B���P�ŝ믓/��۶�A	z/���j���o��6��xŐZ����ӫq��H�d��" �g�C�X��r?uk\!1��TE9�)�����#�y��ZgB'O��}���9�v�
��H3C�q�0������d�ΐ�hzg�#s��s��n>�a)���aU�_^5v��u�[�3R�����">J����❔�W0�`��H7���O������*t�s�Y0���?��g[Ъ8G[�LoJ�!Vi�^�o厬�T��/�eD�[֎�o�j��'�+��q�.<73��)gˈ
�[��+�Dl��x�<ܵS$�R�j�1N�2�!�5�e��:H������8{+��o�3fU���|��0#��p]��e���q4tB�)�v�����`�1�I���]&�0�7Yh�3#~��Q��I/h75X�
�f��#/1���,䈼�%�}��$�?7�����d��Z(���l�s�Z�b�}�'����@K�$aE����u��� �{8\�W����NJ����%�1mm>=CW����2Y!py��1��%�
�1r/���+����t|�	`�P��nS���$�	�f^�?��'MS��J��?!Xу٢�6Q�n��֬{�7��ȍM��h�-1���Rur�� �wv؛}�?B�P��ǟ�	')u죲��X -� #�L@��Ii��3�X�9��/Ԥ�:�vY��2��@��08r�V1d{tDv�ԻA���1!&�yo���;�����s"�9D�C�����_=�3� �f�%*�}C@���s�y����h`�ł;C�Z��腚@Q�̕������	m���\���]5���;�Rn�E�-�zm��v����ZWI���ޭ�,�Rp�3�l�h�˺��k���N�I����Yݞ��$ �1����1��d&�b`v��,"L�e9��	�� ��`��-�kW�TM����wT��ɏG�j�튜;�G s5�UI�/\��DT�;�
��9��&uV�;@r�+�䧠��x��^�H�6�\�}�y�LN*�(�r^�m)�W�_"T
G�%{7�� {ũe{�(��q=�>�Q`	�AT�ٞQ,w9�FɊw� B���/L�. ������T��o�2
��]����Vh4��e]FR2�_(�^w#����	9�95.c�'d[��w�[�\)p�5���bz������n��ښ��qG���"{#{�هF��wjN���m��v]�I�c�����s�����F�H�����Ԕ��������b;����f}���Gcٸ'�q�޷�7,fG�D�Hfa|;�LV�cR��fj$��f����86ޕ�Y׍��쵓��W0�b��3�v"���!K�r5��]/�p��T��bwz�R�� ���e��/�|z��HJ<��z/�<].��LF�z�vimQwy?�xJ2rSpȬ4�tg���8�)�e�$q��ET�)�ܗ2g萓2�j'W�?.��MF6��z5���+ւvV���O�۴�i"����w�VTW���=
�
�ω���i���+rN���v��Q��6��^�!zTή��6*HO�nI��j�-]_�H�T�B�[�'���πg>�fݶe�=���C�x%��hv�����$Q��'�G��k�j�8u$�pq�˸s�j�s����H9}	��ݓ�&��7�=�?Z��?������B�&ncڻ���H+X�A�B:T	��Jb����R$C�C��w���F� �8]P����da�:��L�1��*��pI���:�#^�x<�M�����4�l�[k�G�
f�-�j�o�� ��R����>�ҧ������O8���/s��oZ����������)�cZ�G@W<��bO�7�����a?lC@�6��xVEt���jܒ�|CF�8iZ9݅Pl�? �q�R �}ǩ�����@���%����#�Ȩ��D�~T���zgOε�N�?��R34����=��:��b.gM}=���Ô�����S���?��8�b��St-���9��yqfM����48�R>Ţ��Fn���]0L�m��{�[s^��T�t�ȼMO���	Km�3\��2Y��ֿ�vMq���t��}��B�-�Ϧ[s�V4�E;Z`n$E�/&��2��ϫ��Rkm}3IC�o�2+g��E#i~��d�I��SW��s���.��M�N�`��N�k�)�.�vHr�^�c��I`��VZ��W��Z�p�s1'�J��ّ������>d�\��y��>�[ѦO, �X�E�Y;	Sv+��j�B1��w�8���w9����j�D�����D�����۽`q;��%;��m]� �{�r&����������<���ӄ���`������t\����p��ڐ�5p��i�)@�\�2-�$�\��rG�E4,��=�u[W�b�f�Wrј�B���^O�Z$k���*³���Y"��S)�Бg�%I��vg��N����]�6t���[br�����S���ΩŴ�iSF�f���Cpn�2?��Vr�RCu@P���w��K0�5��ʷ^��;}��V�5~w?m�w1����x���D�{ɰ/�r<��s�3}0�γ�'��_-=����qX����'�i_b�?�AC&`���{�5x��By���{/v�#��������h��A�Ƚ�͚$�u	��d�g���ط�_�&�)�a�ppOq@N�p�]�Y)ݏRIޝ����3>Ѻ˖/�𸪅b��훈A#�!�~ �'ƀ��\=��S|���(2t/#jӑ s��Ul���y�Q+��k�[����9�!�6�B��omz±NDH��y���f��؟�㛙=��CЍ�rZ�C�8�:]c�TL��+�R��72U�7U}i����[�Y+�$�.⢤��mP��i��_��t��D#�xc��>}���5��[��tD�.���>���X��$�9;��G��&��X�o�PC���]c�NBk����~��./�7bѴ��il�D'�Z�80(�Y�ڬ��z4Vn�V-D�)Q�]�x���降
O��/��O�L2��l�~�(b(�����1P�O��n-h�D|����$t�ơ��&1����9:��{;H5�'j�W����]z�"{N��F������!g��@5�#B�ለ�/���_3�a* �Pz�'�Dm���[��A�e�7,^���6�1��V��n��0H�F��oc)��T�)�8j�LBZ#��D�lV~��U"Qh����!�(:���_Q�b�%�k���s�jٱ�N��x$�;�RKy��pM*Jϵ[{K{��_�,,��ݧ�h'�������@X�O�Ma�蛱+����viBh0U[�{��s�� ���=b�[��������,)3�3!�����h_�w����T�l�?�H���[�7�V���k��6�.�mۭ�q��5�+��08׻���5�b�̐�g���Ozu�S��/���oP�{JF��`����v�\*,yZ����e������X���