��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&���ˆ:�����ˏdE�;N�bh7���1��&��-��+�q@{ߜNŵ���nש٭G�4Eɛ&���މj:�/��h�e�3�{�b 9�৆H+����K�mgYSZK���e"���!nAp]�c�� I��$�mdD�Q魰d�P��S�@����j�UV�&^;�	) ���]��E�/�7%ma�ٟ��Y7ﰅ �nxn��x3y�!m�]{�R��+յQ���W�!(v�$P���b��!���aO5 �R!W�?���[���c�/��Ƃ�ҩ��cb���;����k�H8R���t�X�t����o(�Pc��
�JH��Z�^N���g~:0)�ͼ��χ0�H/�a�Cۘ�ش'�����fc׏�mE|���oLi=�����	y�>*|)�ay�u�z�dz�c.�a3j�ts*N�.�T}�A���ĥNǐ�j�I�f����`?'�4�@���!hw���p��Ϲ$���C�x5vӡ��Vs�R�Z�t ����%�j�����y!a���?�H�G�g�k���s�(�w���zwy��̶A�(�v���c>��,L��b������ %�0�<��5R-���W�[���C&�6�0�����޺�C��]F����]�_���@u#�Ke�|�f���=_����3b�郈��(�S¹�įBO���\Fŝ`ݞqN��7�N/#^�/ʳƹ�Xv擧dd/MM|����d��� k��}�s-�cn��4鰕[��^#�c�A�	�]�y�w��3[�ghnW�w���Q�[%��V���޸�'l��g�M�s��t�Vf0a�j�u5bt�c�Z*��A�5�(&8�y�z޾Յ��A�/��h���O�%V�5��?~A�A���a�%uT��r���!z9տ�F��_3D1��ѻu7�A��Sk��N�?^�Q�S���~s��a�Q!�',�'J'H�s��0R�H��4�[��l����Q�S�������bmz�y���Q�0�mP�����6�7+�fd�5�L�M9x�<ϛS%�͓�P�'y��"��R����=�Z\1�,M����V���L�@p�g��?���d8M���U�a.��gj��7��0BԾd!��{���x�uQSUM��Xl�ج�2�1=� �������K�v��� ���������_���!����4�:6mQi� ��+�E�b^�����d�s��e�jrC����C��X+�uXJ2naqs��u��bѺ�R�7s^����mmK��h�Ҩg&1+0;�f{���"Cc4�Ԫ��d�s1��X�l����IaЋ���3��Vd�����摭[^*Ȝ�<t�
��q�F`�������C�oq^Q����V2{�ͤ��|z�yᥒ�7�\�/���)t�R8���B�g����Kme��>��E�6�	��̼y�l�E�JjB����4�i�(�
�'j�q���d:�	��N�m�����]-K+��^�<�� ���fʩ�I���,���v���;�nZ���=�}�<3��m�?�R<Q`F��#G�~���[;ڤRg}��ZMIk�;����3ss�,Ѧ���>)���U��cA�(4u�d���-T�	�f�/C#S9˼��?������b�� -(�:���C��П���癆Ot��Qe��0I潆�nNl�$�m�M� ��-�O+��nv��~B�I���s~&�k����X������*\���tx;S1�5����G^�&�qDf+|�4��ӽ;�N:w�� �j�*5���~�m�g�T2��i�N��zb"��F�d1�W����=F�S���x�>���u�`[2��c�9��MC���>	M�W�f�F��e�ȯ_6@zd��T�}� ��Vǉ2>���Fk�&w�L���o �$	�t$�2Ln!�r?�e$2�; �/(_a/%���n}Hq�}�����b��Ň��?��x�e "��==>*�������*���y3��D���Z�����M��@���Oq�V�5��!�����	]s�9�o㰿��s�B�?L7�Ѐ��:��gF6���R{2A�VX��?O3��o�C����*��·.����-I1e���1�Cf�v*��`(�r{�d�� b�)�^�)1���=��$5 1�1 _��2���~�][��t�3�Z�M _��7E�Nh��z�LP�<
5ib�r��/�L���s&d�dp�>��^O�'7�!� <F�NM�F�)�[ߍ��Oi7����&�?5�����J��=�5"���?b��?�d�r�����*�l�$�A2��.}H�O�Y�ᥣ�����%1$�XF}�Ϥ9�3�9��+�W��.�o&A��G@���3��]۽3,�l���F��മ��=����Mh�C�Έ�t�u~��"t^��8=".�L%��U�����>���j>	�w-���sG3Wa�/�0`�[W
l|��5���iW���4{1�mz� l�4��W���̿���$w|��`?7v�s)�4�ס]�>cn�rK؃&4W�a��\}#��J�c��u�յ�?��R����j_q��b�"a���Gs�D��	Ͳ磈�&*3�pj�k�B�V�O�ݯ��GJ7����<���vB$ ���_��8������	~���teg��mPURͿ[��͇v����ˈ���G����i�El���:�'�<�Q:�BUlb�R��|cܚ1#�b�ks���aPLL@#k����X�.�7�n:�3�BDSi6��5��;�֥wUf�y�^�?���.[CA�n�w���,d� ~ +첽|,)�6N�}JC��J̯̄>�
F�9��p����ɲ��&#4H����4�����Mq,��8@��L
��p�@�L/���"����X��^:�l�B0�%���x�.
�����B7�d�h��Vq�h�<�0L��hrx�T��.X31�D;�����nS�]��6�f:�6����q�������\�~m�����i�}��wq��-�Dk���Ώ��L��D�{���r�Iu"�f�'<�LfU�UI���d�a<wc �ov%F�X�d�#�\��^�]M�h�.�@�=^?-e��1�	�G�_�(�P*�_����v�0�$�h#p_�;���J֐��kn6o+���e�4��yԡ��*�ܙ���Ja#���b	4�2�gZ^613OC@-��;.�oI�}(@S�æ��p0ꛕl2Ŋ��������3bI�Ǟ]��W��W��^YF;������ xR-3+���u;��"}�����_��j}U1�ɀ�m�ZlF�	YMŲ]��ٶ�R��囋X��@��v���~Qtcͺ������~6=I���e׳
;�M��j���4���L�-�M3J�XK#]Os��;@�u�����~wG�i�a㮿>�/��HC��WJ7qQ�.�W9Q1E̤(�Ke� �#�R�|�Q���?��+�rcM��5g޿bh$��I�;�2��nB�9+���:���RxK�M_��O'���:	?���ܣa*'�@�ݯ��3�V��.Ԥ[J�DaD0T���46�Qj�]&<fNSB�$OG���xQ��C> Y�L�x'�43pܦw��@�(N:�4��2C����$�vw�b/DwOB~����.�������kkK��O,I�]b ��>|�u18���D�*(hQ�������-���h
{/�i�S�>��g��ObɃ�y��0���Aa�ajT�8c���;߳��8F �w&U�y߿��� �g����b3�ɭ��n�`T�UҲMdtd�`���?0�+c���kfC�����M� �}���3��J�,���&Ɯf��7N�����@3�n�w�[����ڈ�u��+�P\S��k�Xl�����A�s��ud�V���!Z{�����J,5��\��]@��)�Lخ���#}���9��� �Թ+ӳ<�X1i�5�3S����R�u��v
V`����?����Τr>n���s�Q��+�\瘉&�ί�'=+������>��>\ˠ��
9���׎�Ȕ�]�G�_w��!�@��߈,E�����KU�ע����ȳ-�K���a=��%E�ۥf��ᙼ���C�V�Qf���x���i,=v$��?@���%�2a��$�>4P�a�_�k�j@�b.�}OT���bbT�9/�L�[f�a���Q��֛����&a!I/�!$�2TnYA�]u/Lu��ru�:�X
�Tx�����¨�Ϟ�#�Y��C�͢S߱r5.�k�vI);�[&�Ѥq�#�1����<u�=��p]�	�`&��RЗ�(P��կ&��^ZY������\�&�n�M�Y4v��Z�i/��E��Ʈ����-��">�I-��J%�����uGZ��uO�]%��:��R�N����8�8Nc*�\����s� �^�(���<{����
-��Յn�e�ZD����lDp�9��h�_9��(��s��JL��$�Oק	5z�K�^KYp���bgt�ޡ��y�I��م�Ҕ��G_A�ٚ�=`
d��+o�+�[�1؂�yH������C���ű�?V�P�?�^�1�طÈUq�X�b�2��ر`�fd\ҟ>�(��qP�f��c���f��	���o Bpg�M:��%�n��]���O�#�W�D{��t\�fǺK�y�� ��%b�w�:?&�\�9܇��[�3���w�	|�n�'=)�L�?j��e�D,>��)T]
����svE�x2��Ì�=��&H����ݩݎF����Z�e^�n�Ͻ؝+�}흲y��h�[�������"E� 6aPղΤ�Aէ�Lщ�;4X�m�\a<��2#�;�T���,�\��?�p���`��Q��V��M�>���;ޜ]7"H쇵���a� ��f�5F,��A9��k;���[��J����|�rq�����ϐ�=_+�� �&�C2a�����c�	��BnI(�FG��#w,�g��?�YN4�\&~O�҈˝Q��ϓ�����;�ۊB~үT��*ܺd�QlL���x��DDd8����;C�����fY�z���+�0������4��F���A��vo�IVc��ߣVj�_߭R־W�uG�㣦7>h�'/ѹh$���ƭ��}Pg(F!���_@�.E��X}�d1!3҉)���?A�BPu�K0�4�M�A�1��+J�T^��:5
ٜ��um�G�^�|kl���؂�����N_���2U�BG�[��m'��(
&���v�KEv�y�������	���遚�u�u� D�߱#OW@�;5 �w�*~�0�[��$�������q�M����"�#��G��E�R�36T�^&�[�k�vo�=7���"����B*��c�	B,�\�����g�&Z�طR��V��@����,����sv��r�Ecc�p̐�*WOk�ڭaĀ����/��9�#�N9�;J��<����4x���[�ƌ�|���f[,X,�7
�*��y���,�KD��9�Э�h
����>\��%���+tͅA�l��ii�m ��!c���n�9Ǫ�P>5�W� ^��>9'#�rғ�����\ne��_2�:�ѷ)P���m��B7y�r7'Y��O���B�;&�އ5-BV����r�e�sWb�O�S��%������I%�ZM1w�v�qd�ZJ�0�Ԙ������w�P5v_;��1�7��M���/y��$�_�����0L������ΜvF�Q���d}���sj���J��T�a�|�ޭ��� ?���K��SC���FJc*�����u����F�[���գN-��@�q7%���SU9p��yd��r��޷ýY�X�p�5�fw��n�<�Nf�<�w����*�H�z4zo+1[����HE.L��po�'y��K�K�MK?<��Y����9{�:��tlYx@<�DO�+�c���!��%:�c���8L��{qTԅn�7#{�aK�Z�ѕ4*�zb�7u2�܈B��Z�1k��W�z��J�f���b�#��L�E�P�/�zp	ٿ{ \y<�:����-?�;t��v8�-7Nӈg�L�m�s`2=<N7G'C�l�WϏ=�(�5��R��~������x:�a��Qt��z�JGjr)���?��|�� �~�d,|�Ol�m_�Qt����������������Y�\d��zcnb����i�/K(R(��'�<ʀf�o(��·�o �˗�	7�G���mʚ$������k�p�t7��>DM]�(\~5���Q�v�w��SK���xe�3B�O(|D�㝉����P�hD�����{���*vJ��5�CՀ�`�Z�	r=|[?=��9��'�
���=Sd֍O|���7'<&$YXx���n��<�B?x�eĂ�ϛ���a����@d���0xq��_�k �Ϭ�1�"��Zĺ�wI��8w�.�� @���,���U֏��M<�&J�PE�"p�u҂Ӧ/�����Ӈ\ ���p�{���?�+?�^ul�DC��7�I*Id"��+�" �ᆪ��t:�H�
�I�ز)��M���S�j�W����2�0�?����?���4ۓ}���T�W,�T�,�Pf)([�����dm_e8��J�W�,�纳�q�x��(շV��YO�z�eZ����-q��^��Y� On�j�7Ь��ٮ��=yP+?}E=�$��?>�F}G��V��{Y�{ŞI�x`�p!��F3��ێ����4���/�XOS�j�H�Di��1 ��Ѿ'k�����ns,�Z��ݸs��@.���j˗	�'�7J�Pr�Y�}��̇����C[>��
��Oq�2It�����A䌛�s�K�S'>aiѮ���(3jl����f��V�҇p�0E���'o
Ts�/�u�����¹�l�����܃��~�A��_:a�V)���L�=8��7NG��`J��� �Q�x�͑ŉzO���􋸑����)��4�=@����e8��9��$*�o�l	v�'��K{��|~ɇm��
�x�#B\`���ii��	���ʀ�$�]�6�_�|K��(��k(���'��,²����kl��m^��f�*˽�T#����/����Z��	-�j���P:�mw@C�<�!qR�k+˒�>�s�|3�F2N #P���_���_�;�����E#�$�y����>v��&���{��!�J���c�Y�!�O	�Qa�D��Z��6
��E��3HU\U��5�ȸ��p��iB�Z9��R������D}��n��_���P-�tlE����T]ȅ՚tʒ�H�C\�������`�R��ݳ7G�\�_��	�H��F�}�u�g���;�}��9�x9�Q���e�IM8#�e�$��,���Gԛ�d��izp�y��{��.����P!�Ir[˷+JV��(�9j�y�%C]C#��($@|��]$�Y�?�#͸)`=��z�eѫ'*K4a; _c{�8ԓr����q��{�/<��T��%r:��{�e���A��;�CD/�gpo��_m�'�<��Pt���Mc4!y*�'�s������n�k�m{-a�3M@~�O��
?�|�50<���[�J�b���l#��u~+��(�jLxS e�?�婑N��m���������u�"~��ji��}�|i���?ysĹ�p��<��nԒH���y	9�N�������u^ю�y 7�K����㱱pu��,b5]I�_"Ҭ�����x�By�d)��6J��1���ع� �-�p�\`�ۥ�nw�����C�n�xF�����c����=�@Q��
TE�V�Ɏ$t�� ����v��VnHn~c(��s�6��u��sT����6�Y���H�56#�,�|�|��y�o�@�`P�G�.���KD���bi*�%�(�f��PP�fBX�!An����+����ZxI�Yg��< jtx$Z�t�X�Bt��~��b����W�"���z��V�浫���&�)0�_n2~��"c�yo_�J�c����W�vDc�EJA��4��!A� �rv�n�p�c岗f�n�p�P7n�$B��ͩ��b�WjD�x��`yC�q�a��,�X# �?着��.��=�'��r�~+���G�w�1m��B/�Jy�x��i_�U�H%BB���b)��Id�������s°츰�*t|
 �u��YC�yL��%�v�*�{��8}�LX���9g�]� u0,�/F|'���e�U�N�y�L[��?�E�[�0(!~1�9ޤL��l��7<�w����[n�h�Trb<����5��N*V~�V�@2���y�̒t��M l!���y� ���H�2����
��Y�a�h�
���[�l�w���~�_�Q?��K�)7�U���M|�K�����x� ���!u&5v�[*�{�����O�fCgc��S��Z��Q�F�,�O�7߀�4��DF�o]�,��w�
:���˼6\�3�
M'""3�Y�DG���}�M�N!��td��Kj���:��f�j,hT�Glo+����� �����\��������);�)�@3p�2#AlH
f=Tw=}��h �1[_�ྒ���yod��)h�'
�û�4��է-���T�Y Epߦ�����`������P��m��k�ήM�W�_��͘�0jBZ��c,f�]��b�hr?boN�X@���=mXE��Z=M���� �����K�V$:�����{d�ɒ����ORT��P%�Ǒr�iۭ&����B����=A�S�}gh������v�C�3Po�
Y����P�*���.N��ȬJ_a�c�Ƽ��) ռK������`
������\W4�N�6����+�����)~`t\�U��0�vd�I
Ύ���huY��,�w��y���[P�@t͊ò�/"\Y ���U->����]�� ʛ��������0���蟉�)8�?� .s�8�X}�;4y`'6ѓh�S6uែ)����������W��F
�w�[����-��[�茂�/VĕΤ�QÎ4�-JȬ0����7�M�%�����n�p�O�/aJ�NIu���v�c���J0��}�$�

U���4���7"<�(KGz��&1��$�L�I�C���6�E��OE2<7v29���p$��[�d�������W��{׍ism��w<���\���a�Gy�q�
��zۨA�I6E&o�9����ȹX�uv�1673h��s��sc��&pp�d�U�K!�'�I�9+�7P��lP~Ň��`z��e�*-mx�"Aőʰo�
9����S��J��p��ni[y4��7����S~���mJw�-B�h,}�l�4A�ε3�=���ޚ���vi�R7����b�C������m��Tc�F-�k���s潐��a0�A&��YD ��x<5:K�s�C�Q�|k[ϺJY}q�s!
g�C���u�9�JHK!k�Q(�tV��ڪ�o�l(�F�X]�/� Clĭ�O0�N�+�%	��@�Q�@�o"�x����K����ЊL��k;�������T