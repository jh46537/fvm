// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:32:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BxdLPEWEPzl/ahZhxZ6Gw4x8xHHKSqmoMgsUNT/KInBMknf6Bhq2qK6xKbm1NVJv
NXFNmkZpECry7KQWZQn26MFMYwcEaCxMETCU0tLK5WR9s7vpuMSHuj0s6+8iHdH8
x3QS/qB85tRZHOOmVIgwopMQQl18PzRIM94sy3s6amQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18944)
XjJnLmdTc1cLqJ+WDKMJPpv616OHI5cUazFTDV+30q0M1w5DSf1VsBLqraFXjRXu
22gL6qukTWk39QgV8dM0kc6c/rOip9or0bNdDD8PdJx0PCEo0TimLmbu0Incfg+9
1jUTC+kLUI287Trje9nZmbL15qLaNBBpMp/hmX+RO5rCrQIZLzIFRu7c/UfOAkIg
UeJGxkJkG6TjhPPrhnbGryvtfjF6aZ3N/apbymkx+bH0sDTBDF3CN01yjhHOjvWt
Ykq2hGiwgslsd1u+YcZLHe3NcAIgDy2GWaVOUfro89eHvdD0o+pwtBVV9Thkest/
MDL3rzla3+dxMq7eK7G5S89k8wBUoiuSorS8EHnvISGCd/+XiUwO9a0ZWZBxP/PK
m+if3b9/zgKELbeFZd5MfSBAE7DX3L5r77hHo4wz3X+cZoVpqzzySHENCEGyISN6
YSNBAHuWeyzve4GIB7inOBCjMBmmkdVTIiDUd8f+boOsSGJluhk7vDHpzPosKUZi
TD44i0BOKYIbW7ufNfJCSBjYdRpV8pvu77+dCFgAHFSesL1KLwlDtdVf6cPSHGYa
wpp3PLUU5h5hEorTijvnhOI8Osp6AKPMnd4gzUTr9PTS2zes0KHLcYtbDhbtVSJn
xtHRdg9mI7bnektDsZQz967r67wWwBGxw6uq8ILeZiWskG4ZlEpnPZGkO+h1or9L
zzKL1yETuOPT1QVvveiME/q2X0VAHVpvlZPRniV1+SSRI4rbrLR7PkvMFAF6bak6
pJGeil6L8Wr/+ZkjR/8tJHEDq2DkUplsIyxKBz48nuWrb8AVQXRwGuIk2fFu4amc
ifhPGifp8pvBYczfXGI96rX0oQQdOJgo+jItHfWLcXQ9tGn/wn+nbtRxMB/I4KPO
hVE/Aith8OySqbtWKepP/6oJxul6pAgBEcaDffTDRJr2Hip8qiKumV6tVVqtlASo
AQQ+bHpC0DVtHRotTZV2ii8l4fxpfcxRBhD1N/wrzA8yMd1tPU3pNoD4Lm1lk+sY
aV+U2yjxxaaqywGgrp3XaTLdxzg8Yhcyfw0by/K7QuXv5XPNIw7uYMQiiAXDJjvM
3ZRG4zNlOK8IeRog6aFwYShaj6E7xKnEfVJ518iVtXYNxcfL0PZd9Fz7QDOKISrt
2zfcrFNUEi7ekzAIFs2kiIsJhfywAlXSTpXyOptvPo0C3Dc/KpgCLJU1b5KWYgt5
N7upR6lNufymNJdFVmBw25COXTDwCEjoxg0SOYzJ3AZUql2/1Q/2uWZSKlP8I6v6
h2EPRGHPHUlvP1KSKEfMOE3hAFz/SxWSrWrWtrsVgrPaCiq21Yskg0hASBKLg9XH
2XgSe+mywKyIS3nqNoufAzzojFlfsNgQSjgcevz0El4ji/W3Ibgv9Lf71zW5FlCl
4nDSJ4xm0al+vmseeyqG2uqq88NLj10my+v5q8s6Rvq8Q/kNz5LIRT63gcrs2d/7
ojJ8CctKgR/ibwQ+m1ZLFdFR5iozxC/wKhMORwGp7IT2jzeipWPu2ptXZLpQ3Eya
REHRVsa7YuQD8hz+UH9gFYNN81V3Z9MV+3mecCkzWZvfU5whJEayDJeoQZYOxzsF
3W6wzE+E8lRgNwThXozEw7dy6fkS7MqnRCxCCoZ7wXzmC47zrbfgEryoLFG1dK+l
DR3yxKZrPzpAEgNKHTGBx5xFun3ODCHGDq3UVbvMjkUP6lHUCLuBfI6ny875xD3j
Eprq5e6Wp2O0pdGLhqKtWOmAUeme+1dQO8+vh/+HliWo+OtU4+Yvj/LFK9mUY58R
rmzRSsbBlXBJ5KROeRDeAT0qWR9FGkAYBlWNhjkOSRx7I5oa8GXaAKxcsfec88W7
Tbvsb2clK6xorxCrEnqEho2UjY0hUAR0YmEg+EhpMElNpHSaZERBSvR9YRmmwXeX
veBbvT1hYrHEJr46A3GNb0XqHQXCPaD0H2GtochhUmQvyaiBIGnT3MI7b+jBBgL0
yV1MGTLRgiSkJLj48dqyHffjRm5l6CQVRAa7eL0S3BdxzzWv7RAs/OiHWQGSVpOp
wH2b13gSdKEH4g7q7C49TO7ORvkfYpT31aEOAu3hgPtUnmatM81HB5/5y4xC2spd
3sSIYQmj65dYawIwO+zRDUdSEH9bk0MV/Ukt2gMYkt9F68efQzRWl9it6XUgyQdJ
7HXmlxQT+cyLHYElSEQIDRg8Cj1sB9uRy2kx1js/rfJoQyp/Q4mjOzTx2yMLwrj+
NsKuE2/sUZA0TNoTRjLMuy5vTZnl300R0QN0cdyGOFVIsx+0pjodvcr6mxJqSXhW
BrEl2+Yjjgbx8jZuegyWoD6/35H9cwis+pXZYZklXeDxP+F8ose6vmrdDgUU+7MX
YPy+xr0vgZ7pXdeyx//f4El1y33WL8zwcjx1UBFVqqqOPWYGmwvuBzCTGbVwfA/N
DY8IfYsqtR9Jj5HsgP1Sz+mFftBW2FZyh16jCS3+WDLoicGvaXJj+XN7HY2aF/lq
Z6sPZXn8vRTAWV5IQ1nprY3+d7ww+/GWdUrP52zwlfZma/Hq5oDh/XbaA/C51PIY
a224DaPor9AIbRQcndr4vyafP8aDQsN5c28yP2CDJsRLcdPuBuHQXyzw9T7tZ0d2
RjPcPkgT6q2anx3zYlveNuGhfSdrudNqJ18c3OGlA47oBEBBFmuL58aMnIcwm9dz
gNQXyHt6JFvRn8cCLLc/T30ItJT8Ui3GoT06n0XkswB81WZ7ic+8bFlwTROM97bS
45WoUq6oEo6Eme+mL67xPiDY+yQBh2aq3kmAFAIppo9VVEmGdwZqQU+iKQmIf7EO
WwqUVlG3qzhxWibKMTTUL65nhjnCM3CKNpYxxJhealEQa3h3JZeKboRaoCP7D/rp
zuhpH/lh3GEkXQadsweqiOvV6uH/qetpBSFmehBRKYuyXYqYyHyZbXNjTaqeXuN8
WbQ2PutfKdSc58ATTBVNvDDe/crZ35GpUfLsMin2tyfb3rXo4GcLxkVGAiPT2t+1
mduRvuMQHER6Dsh7NxMVpdJm3kjmtlgtt/tfal67B2zEj+B/o9bxGghLQ25YkGVt
MbSN5Byjjy0yrKYuKQfZRX0ftnuGebTSt7ng5VHhobfeyjxV2cwL9gY20su0TZ/7
XZSdLQHAyGsgtvrQE11z0SEFu2QIRTQ3sNrPc/yHNBg9qbDgspaLCrAJMgC2/qwB
063oisCcpY/UPhwB3845O/8yFeDRmNcgSqEk227hucNPKqNGsrbUcTIwBPZ5d/KL
Tye7ccYopvqIsPKieKhMfD21WNImhvcdEEA2wrPhTxXPtlYhu/exLK+VrrMsaGXJ
r24m4Ku66TRfa8J5f2pgGhbpEzMsyD3wrvisqNPM70EOcVz8d7qulQOpodxosImd
PCfwWj2vUc1xhgln5M3DRiuFYpXCZ32GjWrggUNhwU3++yGl+S0SBA38LKmyNP0c
iHtkEu9vNeHnTRpUb1JKZSc/XgNVMRi8hVMi4DGcEmxgRqgNwBY3IjAupHxApaCP
yinwM4j+Fxwg89LeAJmIOkJ91sFcA+x3xVIsEp65ssnwJVJRRddYD893c4JYxzwG
CK5oREUMHLhMsJyW7qyrB8TVs9iCoTe8qCIMkiEOv4ZPbdhtmlVo7cXEY4NWgPLQ
kF3wuIdHS2xLpmfs/87HL/1NHa2+rlrLKPBkWqVpxnkobrUWwkxGOeot8ZaP9T0d
KQlkED7Y8dMP0NftH0XGcbCg2mnqpXQXs0boZjZ0pJVmfWsfSNfQxHkNw66Bv5in
6Hx7H1qVHdY+GiylUeE9vd8P4Y64F4DMwwIKVQktd1Ks4ODGNcVMEzLkeQZdResl
m5j5RJBZ1nCu7/PS5OLWrcdGGY/kRiUcaTKTwrXE7Jr8vblqWYZ9X7eQZqjZGBZ+
jauf4bpb6dOPYRytcxs0fxollrbcx5HdPcNyviABjHQ191P2GzA8dV6rchmSV6Tq
sxWdgzLGZWVbKJaecYd36q4a9cpv7P4+U4FHLonlzg8o4/sZuHgORS119bwBj9Zf
0a6hbPu/3csEMxJRZWPkRCIg0TOKSIHwmri3uYugkV+OVEqIZdny/jUweQO04HPa
8hFgUkOQ8QMAMd3cHws4gwX4meHReZMpOjor0GnhSuZmWguLTxVA1rnEOItwWowe
bpRn+w/1DsbQ2jPBq+nzBceLp4CZpTgk8xD3aHDD489r2s4M7NMRbFHMuwA+uAqT
US8yYtu3ZTalxa4g50R01jNf6z+uwrE09ivOLFRDROg7JDecDD3kw6osPlhnKCV6
LKxIAY5dmJLgwqbqoprk1Yfj4tNhbLtNPs86B46lbCyHTwGsV9qXFMnUS0HgpDHK
exV/rXwlWW2bYaKegRMtBTlIHUc91tGvfRKHubf+k/7QbYoQSM0NHCz5mTa942hl
GCH3Sb6TqnX7YZ97AwNAsXt0nSGueLSdFpBHVDchQfo54yKRTWCfqDCd06Czx+JV
3sOgSZKmqGT4HAf8GyBRykQsZHcVhfOKM/JgGxXNup3XXEVrWOASTWkPJAxoRcM/
KHvcTl10T8oaoEMsO9OWfTbGw96OYwHxmxXnFtyJHAlfhU2P2aqdcYpLkacmrRmu
vThelbt7RFJYyEdmyytLgoOJ9U/Vb9+moDFC2uAntUtT9xfQd1xDtvLhnCxWDJ9x
64KkUgIzFaN67bMSSBy/8YghafTIl9Rkg4Ey4KCfIcUmawhmLFEYlQVlJV4XgRpb
I+RHPkGCOfw1R4FvyZo59mSyrbRNPQ3R+Y+ebb/a8hJsAAgTFvMV/WEafgHRoVCx
5aG4DaFW5Pewn3wwLd8Q4ufSfPiZTvBGpRwiqedz7DBFHXb9iPlwta4eGiczWGmD
nktcJKUwCv6Pu7tVKPRa1r2JQq8sYJwAJEBTH5JmO3bkJ94olvhMaATgNiv17xhe
tC0QPyk+v+3QTMuBNPKdQE18SlKlxtrZT56VK+B2yobDaHuijile2oCRbLSqQ0Ox
gPqiw3rTX35NjTjmJrNTXoaYtAhR7vbEM0YMkYzejlMrAr4pSPeRwel2SQopL4CP
rXBg2ETqr8kYxTzrTsoFVvqFqEVhcY0979kI0ggyBTKynoD9nPT8YAJ8FYYJcdc6
dLW+Vm9dOIK1AZmftkeVpNROWJx62deYdpD+/lKxkEFZFOlHh8xcF8wB83wcdXti
7XLFQ0dixZRn9JSKIbmIT21WjG6dwfQKjMmeeKa+Emlh+r7+7JkHBGxCxSRQYiuV
UMnEhoNRujQT8gb9YU76IETnIXgH9Ee3XV6EtzWmmRYtZzFKxezGq8aTQeHtblG2
g7f+VS9ceNXKelWPGpv8LzLG4Qw5rQwjO+FnVrQgY4Mn6rDCHOIKQzmZ/2aPpOYJ
/cYPUYnpJlK0ZIS8DFFafx4a5HdBOR2CJPYltqAzGcvcC6NmRZL8xzoDzTP+5bpm
jst8OccLxzr+KVYERDy2kWC19rcvVhe8EeDr6QA+5u9jdjJC2wlx6IiB/O/FkVNH
9QGBdVJZhL7BaH1tc/U9klbOyUsuwbHwgSM5LZ61rbHa8+DmwwSQeEXuVCnb/dDV
/TSjyl+8Pr+aS6ilADnPLiuL0Z+GOjHXc7I/Oun1CjuK8dOUjmd0F2KsnPVHTnth
p5LyLBHXFO9d2cKhCkMu0N2Fh56Hg9OXtRowDqm1YVXMz92X03NKaonnnlRfruQu
h0JfrTOWJJ1WBO8T8+PgHLEWJF5ljsxHMkPXnHgIL75XgCs0sGH8OFHVdLCPUjY2
AaH2UnKATenrfvDNSXOrp6kHR9fB+VAbPyOGw//5Yb7+6OaIMLau7OxwZ20Rocwj
U2SNiuE8la8Fi7jvghlNRlwmobWzIyUBeoIsT0Epqmq2Dc60D2DmY/8+VVJmAL5A
ok1hjr0Qyx+9Kgv4Eug5kttmIpIwQMCue8end8FAY480HBXpRZjEGYtiA0t7N4lY
EjfJSpckXIVOUHrl2G1B6t0wpVvA4E7O+xUGVlylvEkIEAerLG3m9eBe85E7eC8Q
SkJoHbiuY6iksDGUENMhBXBtaNDg24PX3QTthaFNFgy/NCa8Elx25EA/DdRC3xqK
xPfUz4eY9xYOCQcKBmgIovK7Ad2z8SePoNlybWzz/6zBBk+OupPorILujdrFDX1n
Bc+Opv+F0qdZy7amXA4P97Q8ZH1Wq2GIXQbHlwx7emzMqJ7IEk+hlMsiadyi5R+e
+nFSQcaNJQJix8jf11kEK1H/nnGLh31pA8/kkSX9wFKpaP+lpkooCs/1v1zAcD3w
Nmp457PhbmbVOZ8j4XWnbd7A3TTiJ0HuOc7Tb2rjxGFH5Dv3WEP9mofH5IjzLfiP
5p6qrE80zQD2W27ycHvXvcCV2knAP6ikVX19nJcpgmLmKnLpV2A/o3l6cOI+WElA
NrkXjshYcD6RTd4DDn4QTUeIlbHKepME5/s5a8rcx7O44zM+RSX5PCrU04iM3imW
wq/Rhg7lKz/knfwOIHWev9kINSkdX14vv47XyZR9ZPvtU7n/C/8xwZSTvxkgGdL+
6eX+s/v57cYS/PVs1YlKtzbXPOeZjdLZKgX8SMwoiTz4Jw7wxHdFdVJTWaoTmZ9w
7vcVGR2Uv/1U9KXdgc/hhmmiOYJe6PdEB3Hs95HEE+aMfoOrAbiuY7sVYt9MiB3g
Y4In4XJgtMI2ix2O0DZxLQCUHgK4/pURNcoAt0ChbdD81+T853c0JdNJgNYp7Mg3
M56LoeM0Z+GLoGA2xWsTTDQ69bjYz3v/0fJQkas0wZPFmH4Yczf+9sVF9JiN4j/O
cyUfnh0790wxQzMy2YKk0TXm4gfxCuk1oJ4rR8sdPqvc5RvZT7YKhG4KbXs0hkzB
a/FAbh3HW3KUmX2CvgIWBM3h10dylrlJDiS7+G+nYFlCgYpeS4juSn5Tq0VW43vC
ksIo2dSliO4bUc0+SnFZnWyo9dTGZ3l3X6u3klhho5YLgDJCfRbBzzuYLojC5CzK
0q8VfdJ1/bierATvhjlZsf2lio87v3vqC7dc0SnHJDh85Y/t7YxrHvD940vt9sSB
TxB48nWTV/A1gn090SjaTzbF1U3XAlgDkAideCt+YD2VKCGt7rOfHRKMrnj5VlhH
u98wycfiVo6Jf22hBuka3/vBG+nObPmAFUHblmdvenozpzAaZIqUa9Vz3t2qfd+q
nIIqqRtB3qaise2HjqMwM0S4MR1aVacS8iKpOyDiDMVret+fYKYt1vy0MzTmVaC7
0lXkXl2SMP3YREoIMGD8qzYZ2Gm5UsoHC4MXaop/gowpN7tNHE8/Sj+Iu1ktoNoG
O1MHPIwn+Pf7cRoKJ49n50U/ZXQSAxOEj6x0WZoSrz2xYDDH6suLGRncIExYP8W1
tmB2ync9h8ngPYyb4aPlDatAvWXT6fkVKC9ymhtLw6zHo7DAJGelhhEqJErOkdCN
2ZP2P69cejcyGizlzWfFAVuge6Pzcy95G0Ypl/wvjjPhX+NqOwc1sIK0SSQB6PSB
tqWsZkVnngh0uAVoodT23CafqoJDGJLuKjwGb/+kAcBywQcSgcUcnWTultO1NP4Y
Wh30bOSaf5XRaMTFA47GmFNswWGJ/dImqsD9IubNZtAL6nCTW/BM/GbKyeLrqXJT
2xHeKTrW1pKQko/5OIS2j1zFxxB6GtL7A5LK9cTBKRxReCzo7A3Lun5YcR9sr6Wy
z/U4prK3T0NmuvACvXraut+LYyHqVz2ankIexFr1kqbd1zHS8dhGiMCMCipP8AvR
5XFugpypjcb/beUlFO7D0O1FDcOB5tVEbVE8sFW2NSEhk/eee6FVoibYOz7XOJt8
aHRrWdzq3QURPvwSyTde6SeyJwz+lEIQwzNllF985dr2eKRnXCp0mo8qjfqkoLjm
KIWKfk2Js4UiIHYXq8WRXGsb44f5eWaSoxCcZ1EiiX85u8jNzWDJ5ybzvpYBp9hk
CgOb0sbvIIg3oy+jR4dAYKw4H9HXoSnn9ysuqMAnx8AYtP+RSkfyzrsxojov+yDh
80tIYZDzw6qPWYiJcvB3DXqKUkoNkqjvEojyDI3gaxCbV892b0sPPhr9JdvsK7XI
ADZkuE0snJpc8+/EV7+VfoIu35ia7qLd/TCjxv0JEQn+c1CYNHZiUUGeXb5SGoBk
2F1UVHcn4JnPr4fSIbU6PA0Mpp3c8/WS/G8vhQMEkWaHnQNF+/30HsyuybSau+qK
3I0Q98pWjr+J6LStmWQvuVc2vxyLsuk1nqnZxj49EYwqG5K63L8aD2wl6ZFKsRyU
PzQ6hTzk2YJMgvwU+ncy0pxc9LWjc3Dp5NyQjhVag9ejui9ZfVuOYsQITzDx4hZA
K5E1xVIoI4T7AQrwDcRhMWoLHUb125k9wFl96WVBtu08hjetBTqL19lJLvLO5MC3
mf/fmPl9mBtCg2P3ulZ8fa/8PuvL6iE7hCXuhPrli/gk/ByYQsH9zzMBDacsgpcO
9j0OHCDFndo64WWNR8WcAbzeroZ3dcQ+MnNe0mV6gbDUbhkoj6KlmSEUqtNJBi+T
w1j99/PeOb823KDGlHUz3CQTi7sxg21hH+SnkZoEPVPZ/IAHmI+5QpBIJ8rs+smn
RP8AqnKiISMeM39smoQj62FcxjY1V+CoMRjbl015bNmL6dQcOrAZKSD1g6bi24K9
zwf7ADfC0hdXRjIGgHb+QTkNqku7Fa0Q1tZjp/GfNw1LBiSvZVuyqV5GN8znOTkK
ZjK1rN+ZAYGG5DLxBpu6tpwjnVqkBxjW3IRn0/DLm3rC7N2geVHvkKyLQi1etXoz
KahvsjCSfONQqqvyB0QtCSZWNyfwbMxpDrXhcG21c376K+KN9LvPB2msL/VnZ62Q
M5KIF6phzEYtoCmYJgEPKxQDSb0IgTpfN4AwBB6D6VUtNEWaVhgkebgWeqtIXrQQ
qsTDpp1G4e0HLQMxOuQLZP3UUcRL4z7S8ZCw75EDkbbKMy7YYqjfZw2teo3mfr81
G/q42UeATWJbsrCYmMFlnPrhZS6d8XkVDvRMpDmS+So5G35wEb18onmrQlGxJAnJ
omi5PCC/ue02kMJutHcu8z2uRNTAfnHfzadEwM1YAJFqLmPwLNCcNCuxuns9l6gW
lC08hnOworg6bJE9VPOQzhMelA8Y2JMxsl818ZWq1RW9Su7ngGoIVfJoyvTTTjKg
1k/MFsWL2U/3/ViS/vQ2rL9pQQg99FTSuX/z7U3Ls4uuFvr6x/Q4zyFOZ1etDKOO
YKVOtKWeGqtACEYPydtecn+f2ba3Z5FTI9syjjsWWhihlfkalQ0bPKJyOvG91Nci
cq/AiVZDojHocZrp9v3p4BN2q+TQU/0fUcw2nWG/NxQ6EC+wRndt6NbNFnDXcAZo
+3bUeWmJPuIivhev8UETUDgUkhtQiq2aBeVX0mIvlDizmOtuBSq3X+2gY64j104R
bCJJeaEz0bBuuSB58sRCmdjkK/0vf6k2Lhqb7kgRrW8FUH0fmh9SP8jm/HHp2uoH
6O2p+nVa58q+JUFfxsBfzRXVvx8yg530EmKHlutawpUazCa85FQrwrsRMvlx23Wz
otoMtKYmpAGdfegir8GukRnSTeeu4Gk2gREjhkWzbcMw1VcdKGbLbJwjdjuzKrmh
53oWq5BlNcokUKFkpky0Hd5vWxOoLvxWv/aQEPMEiTCnjOuRpD6IqEvNo239xPmR
c7oj/+dzhbZE8iPgLsx+0u+Dm61KVt3DLabtJfYHcfwHxEr3eq+rbylXRA6SvfI8
oqhyOL5ynoDH+ButNNbZYJL5VJMOCH1KpqWYqHfv9P/vB3haSLiRq/Ds78YXKkEB
BAXZMpVeb32aK41wNuRbRXREPhMyAfeYzohGP2Z9BtRMdoi7fXrDB3fx49XOLmdX
0f4BsLjpf9haswOcaYn3yJkFxzrR4zdyho2CDjkimTQYtUfEteJyn+XUS2bKK5Ta
AvMZutg7urkVFIZEIyNUbBO7V0w0Nv6hyg5Sd05cagapQUtVRs+/bxchVCQgAnWV
RhkrxPUYBi+SKmzxTvfOsltl3zKFdW59jbxU/WtpvPpa1aLGyv66UA51mtP+75PO
D3ttGEz7Pn3+pYEeSIT3y4RNIu9vvfrBVrDfq2OK3KbjvEPJFfPIzgJTXUkzyK0p
KFkMNqQMWLqS7gBwpGDs+QFNpMM5m7chKc06AeUpzto5MtWY6yPvQZGTqlempSLy
qEjU5yxeGNODh12caPtDjYly8rNPE4wVqBo6/9EPqS2KoraNcDIcdHjPEBkEn3va
gLcWCCUMZT3DhYoBF+pXUB8sD3mhrZfeLnPReiV9J1fn/T0LMS/lORucj0fYqfzN
nszf6qmyiFstT3H4FHtG5xZ9FKNcgKL4cDs3Fseo07bSQeaTj8Koa4+dvqKtUbmO
jAkC43c+Gj0i7SqTGOe0IcwCRThX7M/5424i10J9RZvyD0T6b//DuQo8O9BzTN+A
Mavo7KHrCCec3rSIUjmKM1jTSPEbBb35aaLK7bk8imkNhRRotpe3bsxgo6Vfbz+S
gDpUwjrJ1rFMOTABE4d2GDrVQSynCBnFo/OC6XzXLk2XBb8Ah9/sAY/N5mP8V+BB
Z5iXb8bIhiNB2RikhSZOvlxxULt+YeeUlILf31Wt5RqYxjiwkReqOwly3FLlGZ8N
XexjAVLCAlrbu4Z9HqpR2q/RxwbDCruHR4VHGgRIQLTOaPgi1UkQJ2Bi/r1peFah
j/5eqkt5lpRqtCtMONw/kfjQcLnknWweUQog/XpCgtLZBwzef7iFTcIp/4s5I9ih
XysVJbC0xu3djAIylgjzODq7r+fMvtAc38Usf/6y2nzJ+UM1KD+6ShpgGH9EoPns
MehXiwpKz2w/GQ0E8LxdRn/A2MyK9zesp/Q79eJocFj3K9RYLsKsGygj7DGuQCB2
wFRw9zaP0SJIQ2PLEK6sWO1O0uj2H+SWLzmLl4tmp2xI+DM/185MEng3OmozlHP6
mNdMA/EAiYvMU6Y7Lz3FyVWE6n2MvN6k63tQF7oCueF5v2RRNsMlrmVCeo810Q4/
NPV9zC2uYrnxHh0Mawg1FETuUlSA/xTk0U19I9zpSGwoZ8KsIGnfp9AOacf7kdWs
2TB4HpebuGGIFfsivIlhRXIYhO4zjNAcV5Uh/FKf77/a7PyHcOaR4ZAZ24ppvgHR
4dcnryQ8x3zg2QQeaqBD+PHMLCLldC+GFRB/FUqSb7gSPeGQHc3HaQ26hnv4erB5
SlnhA02p7KZSGfFxBh9h+QHBir58PKbIbZL5TdfMHZuZz2eSO9QkBb5ebJBmJ+6S
8phKBS+Tlz2dk0q2YpRNwLhEVAwZn+aO4OILyUm1XGW+IQy20bY1FYF8XEgq2P63
sTasuKTib3OGMKQWR6SWxdzfeUDFOXKqGT1cT2+thmHjmmABpueedUBHkYP/ZLEU
HAxX5oD6r9THMFuRss3kROe4/rR5552xp67+tsuwkRkcM4SfMtm8tF6XUiPxsHEu
WsWMYgaG162rHEvOYgJrUfRDq5WSq4dKB8Poj5XEUDbuG0SDanCvBOvrkjICZyI4
zybgY2+eZCQzCQYDkyfwouZL59pMViAcWOin3j5WgSuSVsSCZ9toE0zC8Aj0qog/
/FwLcj0ewG7zat/l3XE91h6oo2Ic+WMeMHzbk1vCshszn/qYHQ8L2dFJ/QuIQVmt
bwJNYjp9r8qI2gwVoM+9lWwoodvaLFKELkpOKDcVVsaqefAnMmWLcjrUVRk3TwCv
hXVkHYtVzW7J0cH/usAFuDcQpKevG1fBxZgDGYYAnKAYSJ9c17q0BOlBL2V0OnY1
tHaZ4Uc1/xmAm1cmFLvAahPhKxItEDUb39lMuetJLEmWTZJK9MKNXmWYMwYO6e9J
Ktf+NJe1cr+nt9bBsX57rmgxNtWQxFlNCmvo8CnViYlwAaOUwifJYetezCFvJilA
13eAqB2eucWCwMh5LQqTpe/Ei3JSe2SS7Zyc8RdSXV5h/BRLM3vJHHFre7JjFo+F
Ha4cXpzxQe0K/9iNmXcgdnxOlkIzgpYTnQQVwWEPHmhOHQmwGUBQDLNd2eiNzZ3v
byyXxpFBjYqGa3XwM2Dxkx+rfQOa6eWFy93WCN6LKKUW9omRoUTu79MwFsVV1/Hg
jiHDhFJ7w7/mtnsXmDg1WNglXCu3YxcDVPTqxB3WYgGZhquQMF6SZpEYjuy0gr9Y
h1W2vGp9oAVHE773U2DNUZWu2GSHZqwfQx9KMyLZURy12vjX3fBcerHUre95ow1P
OU+rOUz04wgI3KbwSgibYc3+f00a4eVoHBIIHexn7dEyBs5cRegQdqbYTcAFIgGY
VoU8FTsYWb8QWTkBpLtUt3FEzPv2sr2TuYDy2QtKLif0JsUvFTdfmN1pB3LgJ6kX
xps5Kft+m1u7Edqm9rLKiFP4Wq/hxxLSyIBSvs1OPOaKsJi1p7p2zLHzpakmBfEz
hHtlZEXp+Cu2FGMAEx9BHwCzzULrZB/tMNcnX2V0Lw1loIVXm/TgDm87Ku2GynR0
ZqRuvZRr7fNfS56TBuBEUATPydoeETMMST3BPcVWriUhz3vXR9GCEYT7+Ksa9B/f
BuXXVbBJvyjMFXnxdSzh494SUeOX9pYnL7GoXGbAk9RNSrA8+uqxT1oSLJuiaGBg
2hNdIWXNmrMxcpFI9egaS15iU+BV0mu5MoeJIXz1isiEd1cKpKGqbEom5LyNMgJF
Ac08f+QJ3y5xn0KufOzer1iTD72lUdRZfZ7LWtYemY0P4BvsUd9TbOwj/ddI+y7n
g3i7mDhH2HgRZjh2sd4wjyMcuwgQ1Hg2nK3rPGcU30lD1rTENR6ZmGidQYr1SJQW
r6MpzAriohZVIhJYvLW3AMliu9gcrZs5zSVoHNJ3IMXj6YZmI/FLyvmhBcUH4FNF
SNydudWLeyKWtb8HBRQL8nT3cYt+DLcRqoo0zPQDyeyHuAsGOPAkWvhRfjxEYdll
iBTg7RKjpX6QMdxM3Rw/Ww/SYNVac15zC0959yX72HD6DcAbwUyXyZ2RFhtVolOk
/ZD0a0axxwAXXsNm+C7OoMR4FgZ8PwDYRMRY8tziCbFIqRlL6fDsvHKNkS4BbA79
qOo+Wcu6mpWtsIsOgzqDo7K8H9W1AhLuS/EIa/aWTP8ZT9I5er3ia5wjYg9U5Jpa
OO3ybXIHDdKW+AfoAQqNuwS3KOK03v3MVbwwIKS7aRQNVVN+Wnu1oKYia3Ia0igM
8KZScJ9URg9Th4mcKuYeLhsWQO/d3XV7yQzLJl+xEeoVqktibz2R0IoT6mD0qr3p
Jmf7yDJanZzApbkrA+fqE3wHOJ809OssXNYS8215W4EQTUoe87ZQx4DCdXeYYvL9
3BISi6FfCrRQ3pdMh8MCY31zrQLbws0FQ5GWwWi2xAT+CECgpD+S4PaBxAjMH8ua
8V7ToHpAv0j0OKV1h8nE6NXdz3rnD6TkEX+RH2xYNGbKw5uPcRg4OUosoZXF1Vkq
GJ/Ix2WefFkrA3nrAENUYOinn9crL61SeHPZW/K2LPeSYCZKwiwd5pwFiCZiRso+
Z//6dVePzluiaw7vmZL53JwAk8D7vTi+4LT2CIEEivgdXbezkA5rY3ImerL2hERp
YemzRKtLairlbmhFhjTfopHnuDZz/3KToWzmSouYGNXtP3mp64ynUC7meTsnZ+cj
zzY1ANFJXEkEkecvF/o4+1dyEwEJq1DdEoN+8SiQEvWKjNSglxSJzwOsPJQVhq/D
y7+kDXhYga2Iik49kTcGURmGa3iTvIvh3cIAWve/YBHnrhteik4Loari/kdkcGJn
JOCMfMhjaJAkYxlDgY3alnQf/swVzOL9ceJsKTUovuJpjQCuysdkEoBCgZAngzPt
dGc6fDfvoSuNbhloOmdlM3QeN3b6wUOIUp44NcLEwedOLWG5AEPyqT3EL8vCIckw
VZgbb0QLa5KYyxrKAEC6wFIeTXKmUypg1RVRWHM6FFvjJrUB9Du6WZDCloHXBZwz
+c2u60wz+2mW+KDIy8VAp8mEZBasMw1SEtn0t52q3GlzUoCGXxb3IPK+566Dm6gc
+he2kTna4qmwNf7ONU9H2z7gh7eswTCOd8lOsPK9M4XN3yF4TRIsgAhXdQm+xAcL
KPAF3T9qQ1fFGZZOgCssYFQR/GWUnaZk+Ny0EHqK56IiUk9MTD7UnlJ9KQ4uas3t
TVW8VkGVEIP1gA1espDhrB0dfXJMQfShiIvNtEeReTzI9HQcRylt1Kl0lLuNs5Kj
Al28nt2cb0ak2mQUaY8PvZBa0HsgplrqdmS2bgPaxqUpZfbBVJr4+dHkosD9tBNr
3MW2eLIvncUBk7FURqwC6Jm3DF9SjQSom2zsmj33BRCd9ftGYzLT9BEOkDsn/bb6
Di8JCygwdjmD9g1U4l3WxISoS7k8arMIJQgmZufarKX2eK9Nc6fnIIUb2wj4FAiR
oXYFJYNQnBt8vYqqtR9SWQBDgBiajiSHlrrNe4c/9VxHO3aBXkY/syrKiIfd3RYB
iDjy/2KnrpLX5cNppsi4kOI8KfYU34AdUZJDjrPOQ0HWK9j85sl4GvjLDI/rw0hp
gSq2kHABd12D21S60FfAs617PXRtgKcFS+g5slu7ESsFYZrxnOLV4hS9ed0SE6aA
fbCh5R78yu1Sb7tycLq1c9nAT0RIsq/eisttxyeS/cCRVBM/6Wy/VBVyOvsDRiaT
HNzBFq5tQl4owJSDrSKFxf8ON9YyScXrsmvpeGKeQkHqEKiv79qfB2CDaEhQ8kKV
sNYqbprtJVr/XZQubAkDbkFlarVLxsBJs40Vpa3GDupYI8azDSbllrSVQwecf9rR
Nq1Xc0rdPUkt+yE5ugtm5/KTnuG+YVHX/pNILBhXYv2ipxiwg4NjxfBRo6Hy7RQS
kWrvybkk7zqx0IMbWw4bt4gkPgcThmHMOnGuiGcTEqs00iwH190cnKUIRSW9SUUx
JJYwu68hqhntH6eX+NJTiF3mKMIzGLiELDMzt2XaCDYp5ioYSJX8GT4VwWnnBPVw
z2Fy3rpWiw70zw+d3YbXmnLD4C0UBefAYn0JynFb8ejFEEvnzfp5kA5Xnr3oLwpz
bMxQYmQ1HZCvtz9Ojh+ykZrpruul5HDDqVRvlyOvYUV9X7joQYhU8LOoM2OFTaHX
gLr0cbHl1rtSDdQfOYY+VinsdgxbpD0wwKOL731OLHoToLNnAU+9c60RlARFqQLh
sJKer/of/Oi3p5SknsF83//RIHP95EZbwrShn2GQ/ZzLtp4lrsRRjKqWw7k8sSeM
3hKO7Ib5plWu0Zm0b7TJhC+7wP7W2L6M5McHOPJzSV9jJEvt1Z09SgEpVB8Nx0D+
rK8tx1NfbJcoB9cEVOMjPZa9qa1jhsSdDc5g3pg/wRFB/9oO0SiZSJbTtmRGVHzv
sLPG6EwJN96HMWd+vCkStRjsJzH79zddPrA9Usu4sGYUvln4zJTpSa1Ez6Di8Rjf
yWR6THyHIppw1vDafeGiCsz5UXLkrdnH37lLfwWxss8H1jCmRL0Qmg5XpAyJG/SK
Myn61cWGuueUf+gbyeySKe9H+ab8QUZakVBg3E4WABYxKgRr3mRX/0CC3lc4Y6IJ
nGlAldlOC98YvtvbYDq+mNs9+FYuyfFikqtOnAB081ikcgcDVdUYkUNORDxMn47J
boZnSDYTFJQPh4B/BG0Ql/dfXmn6lenceeDNpzOy51deKueYJ8qO/Z8dZR2xK0v0
aQ2ngnrEhXjcIlm8eoRHsxSq9JGTFrrHgxyZYQDnYMb+76ueDfyfBAFkyo2/taDl
9S/5uBXtAUnC7ym81y2ghbibwHTXzSG7msO0t5SZPiccu23g34A6oJMRs8rCx4Hk
5q87Rx37TNXtFlilOSt3WwFxcJT0O61KDZl9X5uIPRrGtWVBJ1YV6eU+Vu7Mll0i
KzsH63/1LZLymbao1U5cwq6svYl3+Y7ua1oDRAX4apsnRjRrtb/8b8v7BiJANYLA
DRNiIBXlQ1zq6LtlM5r0G3ZGd8E7htlWGFPLSxReQLys+VgWFJV+a5EB38PiGhHB
5NgH3M+HExev+vBOGgWVQclac8HcNEbW+ILDonV++IF0oxzDWch11QUIJzQM0Uvk
13IRfAp++l+ArBkbbR2LJIFkYmpZWzd5GJMgLQhfJdxVmFb0dHFlCSzNAd5JV+lf
RwhL/7TflJtUGuXVbszpyYOEspf670D9hmvR388BVTFMvmSuFq1P4wJ6FzoTlAwQ
GCET/6/iGvvyH0o0tp36LI6i18ZR2QASKapxE8oiB3ZyjDMI5jqj4gJ+30FGSQo2
lzWCVfXunbfYe8oHjobGI3BW2AqmDRpmdXBOzNy95NTGqbhrkhIvzf2Wi72Fpc6l
fmI+K16PSHiW8+nEGcNmpqUHfLcqa9Vb8w1UROLfFlBHBu++lJKjJi5zsV38qsq5
cHvPJLrhcg32+Qo2L2MNdK1iflDNvRiJVEaQjMBXcHstYFaTkI1vNI4JFguqjHZn
pIDJuORSieJ5wXWPvqzkxajgGQj0wdEo485N0A1p5QOgPDEOo3W8qTPDu1N2atJU
gvOFNDpMCgWFw0Wf+hk8OU/+TB+3b2/ov2d7zjb6TZv3OYaaf4/VF3sYXoz317QC
f+t1icVNviHjR0C6Uw5X6BbOB12etsk0Af/o9xWMEIuQ4sWdxEohyfcG3x7QXNwp
CPrp4HGVtp43beYWs91DWv0Jy6Ge0GB0Scb5Fj3ffYjaobJCbxqhalDZdve/i0l+
4U38vTIWUxz8trG84nRCjsXZhko/a+2S3srdMvPxn+fTLp2z1vvIUFvnpEM/9fpG
dQ4OKZOpIVof8QybhhMiKyRw6QW3C+fZ7mhv0TFG5Ij5l6vxpqkTcTqyJSuu4zkv
g092HrfvaXKl8STx8zUWyb2ePnoUahJzkkqXy09GetDPAoqVTG5fTpDXrbhxiKgp
txX24mW3u+G4EQx3GsH90NY2PfZuDrJRJYQ4uPVI5zVA+ZnIx6uqFRMg6VmIeK89
AUIq71ZY/NZGXupkbkltEpLLdZMPwQwhZVatnAuTjeDXc5NfoOeDR8aOnHB4n0Aa
7/T87WBgjDwH+wiGqJB9uPUskHnt0K+m9T5n32bNVuCxhF5ttGiZN1uIYj4wPDZE
3qsz/FMND+ZwUk/kfrGco1rnA9IiAlM2uXIlHTyXqpk+Fwk4KP2DirkZ2fs6OQsV
2ZqUAxrJ6DGiASDaD1hcH1/PRW5T3IjIl9k4CTj4dcLvTFc1X8SMMczAjRgNutCb
55VAJI2GUgaN92Gn1B989tK58a/WfGFZXyYZldhpJRlxSmUpnUow27efKsEvZhSD
cqOfwXPcNSOMRN8KKbnQaoCT+GLjgyNByCUz1urdfgCSkVkkHWurPzVET3cmhB9l
ksd98N0KgFPvlJ7p+AssLofzX3FrUjFLTL4D1dQTgW7anqyfHwzG49Ke2+nZmx17
IhRou8fkHbtTJWsmZLbQg+DNYFTBfy4P2JyOTpdQEXDAmXPhsmmm/Bp5rDw1xTCB
V/BdHHU0eYi3qUBByhZ6kfURfk9pH49EpjMsCRYkf0EGG3o12fX/mJRw5mExAxyM
N3Z7w+xYMG44qXIkqEQn36c6ADFXKtDUThoUI42TkrTsiXhK2PZfFbUxayjaHAWB
ZNeAZQYfFpcVeGxMk+cYsLor/rHQlO/1epZXVKg6kJFihh9xb4kallSq3bK/pkAI
kyKe6wjEepxNs7uUlO1+c/gRUHl/VT0iJxEBQFNBaF7S97XXBimmcCH4uy+z9jTP
Jyay5ylxYTP1wl6vEggD7UsrV3UbOEAEOhIVouf8I2VE4ae9PUYghx+dvuDEcCZx
ysHZeYN4VdmAgHTYfGumHE4mpizKOjjfm8RYtSCRqlTmK0lrQ/LYFaD5eE/MCL82
f7DwaPJh+dutdXO5V18eOh6dKKHpzBNBoMg/5ZSYVE7VOeXE4Fos3jzncMUI36iZ
Xb0KX+bkozqqHZ9Rfvj+8MnZXPIFt3prlPiwb7HJ+VcPtT9bVQHC0cvfIlKb/3NH
cTT+5pvPTjSI3QyiAkR/AAqdh7I89C/Vvg5GRCsd/YUIrK1aExOMLuVVr+U50D15
MW4+boXuTQBse8g4p6HmIhKIC/H4KdibUM4QG78KWnCgnHXfyHIgHYt+yM3zGeef
G8JTtNHTtXVtjPNAugtlQy2VN1jm76j7GBziYTExQIe0GvnSwM6gYlmIrMd9RMN/
RfD9EptwzSezWnmKoTi/82ZaPjbStyJrKIS+kIIcD7AHD/LSCH/+U7wEqmyCQUCC
YYePs3w1SiZmQYqsveukBjHchQsS/jcr4mmQRGTKMcLeA9u4IcBJXNbYlIDpPLOi
B4Sz0zODz8gQkF6VAGWit7KaGIFqVzW3VYYVqRTgt9uQaGwCAfRfRwwIVtG1jOkO
wvug4QU0/NOpBamwCPWaX+4sehVYbjcvP09VYYUHXBHY4G4RsNxNQgQVd4xFm8Y5
cXjpX7JzlbizRUtSObzsaqc1SCDnjZGNQpZuahE5XLxqZXa04MopcFtPMsf/MS16
cKtV78iRBs9nXnnoBrU+IgYiOmf2KK00tcPs3xctz95aSL9ztDjredvsjpbQMtfg
xuXxxaUq6fG4MkemAsp1YGOpXWTqqijck8mv2uxzkNMfMPwH1PvFjAlrAe7xwGyc
JE9ioMeHFkj6yRzddQjT+mBAQcoZ/WkumRRj7S9uooG25rva4F67s3mZCvdVBN01
sbRZ7osQKwR3gE3I2IYKtWGW592BYTUIEo88L8QZoV3iimITetV/ZvbLB/Yg+Ryy
4nAZl4SRRwXGbsOuQuTcpOsIJydOm6DX9Yw+vn98feH0RrN1UoNJn8CVyFnxi2jN
KzshJ7G2oxRxBemPZ4FqtN3O66qtzWloTAafLtnIW5V5wHtSwjO23ZuwJkMHifK3
v7MYSKBnyjFadh7+sYQ2vTgyx245sh6V+eMHh5YAaTdKBMnxuPocLJViE+HhFHG3
fj3vlIPntdtWEgkDGnOXtk/rDaNCvcTnnXTmt4ssvA86lXXfuv24RdpJ0u714h/a
UWYf7G1+nDoKo24N9mD0rdCos772bgxEW0jnD30mrtD+QPARhSdQaiYU7s6vRAsV
hkMn3yM/V8j21W7dNJrn8DqXGTuXUHTDXhO5b+qxUtcb1NSKK7x84Ty52BoaBync
xeQO03YzdUGJT61n2EyQoBPd+u0kJvM5PE1sPSrYZQtFtkyhJngRCad3jSp8igsF
1Hq52ZtCc2scDL/UW/EkjD5ll7C6dT8h0Ww9hoP6OQMKx7xdBJVStI+xSZbgitZ/
ymj7jnr13lk3jCrtUIkYnUrK01LFoTThPps/JmCZ4+YdO57ppXFIhell9E3zFc9w
N5IlTG6cN9K2tLwJGesIO4ctQZGMxxm7P9YW82ElW2JNeuCr5Ol5mxTLJWMZsuRG
tgVkNDdnIGiPUpCPtAv2l8kIr1e8UaFUAcuQVnZO0/mydTCs1NPH6xw8+nzpdVbP
gmmhy7s5khsMFQLaLv1Wvmae4SrpL9lj00+AC4hVjEeJUBZ3lbE0ZtgfQdGWTOjn
T4pOg8S1dO9oOnjjlXxJEDFAp7YEKxxNz1RLPF7/lUp96DthrLSpbmSzoUs2yS3R
Ug1JtbrDfG0Ws35vtDFeKO3oaxpMMSRXxYfarFHQroLwxvvbyT+CZjsXcbnIpPPW
aGny8N3u6OKdY4icm9oAwyN1H1ghHBNo23u3UH4GY1T4cjflOzEUD3B1wuwrs22w
aLTO9Swt9dZvZqU7tXFoba0KbG4H5HwGo7o1etLQ43c9VW3nuOtsMi+Vwfuirflx
1EoWkahoJO16F7hvDcJDR+0L85VHWqKA+AikjQVs6prErGqZFxQb3mmpG7sLcp5m
VcESTZUmvLKX0J54t7Air5BbFJ24B8nE4yqYZHKrJpi3f9thfwGCDtw1iZ/b8H5R
KmvYr9bidl25Mwl/+qEctHaNtgT15f9AcFxH9lHrybKEeyawFjZajlQJkwBCWOpE
wI/Ab/KGo8KVfy8O4BZxcE+xatf0Atfo1Tx+KxJTtxqL8w0lT2CaSt6CgXXU2VIx
e4aDciDLMXSr0+7ZVu5L9k00RxvEzA9uDNaezzGv4o4KdyvtjgBKrJ2hcHUNlaSh
k3skIiMOxwcLsHC/FfT64p8xadRrPwHoSyRU3lXtpgvWbdl2r/NKqfhIHbvWQy+M
NBwXllI11tlIX850vkd9nFbXmHzH0vavwI/L/Egi7svWunoACgjkeKbSOXs4kW58
s2pOHCBSktIKPmpDCd8/1Tfdf4Qtt7c2350ArUSOXE4MIFtJubs/kBTQIrPkZGpM
mujNa1rdg7ar7L/D7Hrt/7BztAL0dAiHJhJYspEdTajEF51a0eWrEb+932/5MTI9
K4tfogYOpiikV5k1ZR+JSkOKsfIOflKy6VDpZhqjWYZNuNgL1OjjB2mxH405qbA1
gn0z24Zuh8retrJM6ZKsJrGH7VbE6vQ1g/npo16xNrbyLUiOSDgs23z9MD94Cg69
gluGmiwZx+w1Xd7KHQu/OaWQMgHx7DIQo2oEiY82xOmXv5Cs4MJP2WbH91gZxV3F
g4p1B/RAk0Qg/i5r+cxwZBIiLwBTkEUrXDG1Xb9axUV0I/5tV2tHsCS5V3DG3iiO
HYw5MrdM/twvFJcclVDpMPToGbbASfFvTvRpuJeGEINdIJVqkNwkeHXPbiOQKhyH
G5dq56nq/Vtw267iws1MKiKC2S/sJKPYTEM2qPUW9rw7hFHEjNaSBMYEn9rHrVHW
o6lrDihujWG7mYF/4glsMZibSAUDvZ0rLtGoxv3g2w6dhAyZ/wornrswl9oZtdGQ
aE6fgL42eV85fMbRTvCNB0ekn2iZoqy9ABeEg+H5rTn1gnPN4yRS8Gb8dFcnBXaB
pRAF6eQGoQZTLH99xK6sxwq1GPH4+hotu4CAllLK+le/tvkwSRCrwgMpcf9mK9hX
St3BcgBuCh3RqDgnDxuP95Ar9PkGMEpUoPmZxGB01sAiEfZWco3xwR9eHJqAQYPf
eM9CG/mTUjL6+EniJ0VtjzqADi5gSsWf/S5BLncEbZIjX9opGHadK1PEHCK8jUxH
vO4h3WJLUJc8KZsaOCkHtYq6tjmvaAW0lBAFmKTmrIqllrV0mel3gbjuzu9qWGtF
rOep6Mt5MEvwwBviAf5jev2vpWkdsMH0UwpfVbaT+4awrKnjMIW7YhlIbRSj7Cbk
1mmCQ9r3Yv65aTrwWoTvniC7+6+SLZk4R9PfSIC3I2MWKOu7t+fqSeDWFhzAus7h
cMEF43OfjMJAf2hkm6Vow/8U28NNEAZFl+TrfKM722tQiaBr9y1LeXT9FpQy2AKT
auqp3Mb4uuBgeKTlqUmtxrJb0zk7Vn28+hfPBh5m6ZJZp6l2L2TrsLXVp3N0Fy1z
Vjvhj2gJ2TGnOBS4BsSs37cMO8TuKaGdqCjR23uDG5YJSTtrL8XP9JY3r0uvigMh
wAa7ZWZChr55cjos953bZz5fKGHQ3shkGfIzz9Yxd0pnpOsPOQfLHgyV5b8JA/Ej
VnNk5vUSNFfaNNmoLSCMX9/Aqs8zbJ0t08gliDFzGZRymZP21/InckVsRl4nWOOL
0o1Yif3a3OqAzQ/Ewv8ZtzCKxnopVE5WWrrZpBDuN7ivhxXPWfQQUEbV30Q093VT
rTK6g3vmba0biUrpyfa5j7MG1HucDuxydcqMdo8Dfgc6k5ihYk8BCkxwxvu+/rLS
4U29m9iE6hxTAyQWr8LaR+lUKEULM6kmjiW9VWtYh+kGtR7cXfQUHuVu1pknNfAq
t3VBvPpctvuxtEcG/IvJKBdz0gfoxySXwsuB5XI0Iug/WfVbEAUjn6efDIsQrOBw
MtZayYtEIJ5sWOzFd31cxUvK0PVek9GL1/vqp3QRaoRhK2cdlPxyunz1vBTFtQW6
CxrIhbsFcMx2ibNK9ToCa0j4R714SkQA3UmYzEe2/Ahz7e2O67njyi111zE1bAOU
EIY3hW8FBzy3n4Rntxgmf0Z0gr8fYGLCXjnW0M1JMX8BaO4kBU1+sO+OzA7r1KpG
+wV2CQnmXmA5hMy0WhhcyaEvDIqX02zmjdVnDfr1TiKVRwHxx7b8ehQRir46u65D
UJvDuZYiMJpyOnEZqvGlguCi8l/8mhxCBKFE/c9J6uxf/7Er0oQTRK1EW907aI2c
TOrk0/foTeEGaE2TE/TG7OVgo+V13Qf7JH8nMX56JlopHHiiaDgf66oJhvqqG6HJ
4wcm0tUsR5yuzA4M94JoXRkqf35Y84xgDqsy2He8tLo9h4mK2pYtOZi/g6kOPjO0
l/8YDCAOTUpUqwq0deGer2a52QwnJ4cCntTX/QkRhK67qfiVmnd9QKLujvWXN3oJ
syQeY95+YY5KzagFk5Uy1mDd6PdrrDcZcV2fYwt+NP9eeckfqnAUhFhwzNCUp0aM
gTF+16fSN2Msfpf0I4hhbyYatpJnJwr0c2IRmqmBhalyQIQKoU3wyeW8kL4Ro7vs
tN7gh/UEpr3//39Ue3wpyrvb+1suOXYOqOCriuGBcJRoeZfOp2aDeyqVKhPq0KV5
d5NF+Z+99FRiQhDbu4x6VLe2J/3duXoViysVZG/phieALVwmNb2Kj32NzpeQ4ASu
Leg5b9D97hmxAiEvEauN2YDhbASoPQHxnfTrboU4YEoZRFU5N0bXwH/KPox32qOP
nQqEUFc28e3N+L8UWKAgCFvsI5QT8x4d2ooaBXjCnAyOFFE/0kUfkuKr0TiGAECn
f3hQCxDaJ+9BVAwlDsYyXpgiHtbviBkyR1uUy6GCNh+HfN4jlXCgT0CHeK4KSuS9
Pt/N4KZ3ENOTQBcMA3tZ814rv604kwP5Ku7bI+TgNyhvXDtbjWP3cglVfrKADD5B
+VgBdcSs69MEDLM/yZ3aPSHzyF4rf+GVudABdVfAq/hVGRiMWq6hUnybKfB5y74x
BNh09JAdes/vXnt2teVk5UgXmIgvv09jHQ00KBdnDJ6PKiflsmvrITpA/4PnC9zd
RmrjvuBKlRcQMfQkBv6JjYPULDd+CuJp0tc3CLQZdpfxffwdFVq1pUY5DUnwK7+Q
my7OibgqaajE9Vk/nclaC68J6jDMj+nU1/m6apiiDQP+XKtBKQudpR+lcZoKcR+D
VvbjBo/aOtT7ufdObPgXUKXSq0RD0DGiSXPu5xF2FexLZhzAtP1u+HeiwcuTRnln
KRVwWzRfHZg+fOln/04Ny9LaH9f0RiNEp74tUuK1PfdcZdteuhgkrZGci6Ij8q0a
x02VYk5qsL5zpZDGLDNz4Shy7KiJOz6teZgtnhkM+xh4/nD7OSbAFGiv9aumjgRM
davZ7vWKnVXBxDs5pD4a+LctR4lDuHYPFNuBfo3t63qoaLBGw/NlAgdAJpl/yOwg
2OH+qR1FtdkfTbLcQWrJvJMauHmPr9dxNSIiUaJZphFo3hAECy1uWBdoe34qIpLh
sldp6KJtm/6xp1Qayc76gCrggL/z1FmK8Sra3oK2HVfmw1Uz0aineF0D4F/cIUlh
81/B8yRX2iX+mfAUgTKQgPcwGueSUZDqFTMpYUAcbDrjnVPFF2ewH5CwA/bnVs12
+wWL0TYB4yLW2LiLUm9MaLbFHLka/n9dnnEenJ7P8C+7XKg/z8eDjnj4xst54Szy
nsYlGYGIAXjEb8SKMomdg719IchUFr77qjquy1uo25UA9z6ajwJjl5wi6PlJwS+c
p00B9CfKPHZmlMaQYR6xBMh4wV8SVQScnBJIf0uIgtnt2mKRhtK3uggfbLxDtlB4
hdLDGK6+5n7K8Ue0aJiwQdUyUpQNJt6uQsDrlf8ljTFWYTGlILhzhQlmYRKZs+23
E6kGhqnylZTuMoDbA8/MfT3vlD7iXrJSyFNpyZjD1YUo99ldXfdGFsJOkPqZ+EdE
cficctzdEIiDal6GzBh9ETofb9+KdVcngM3c+G0dBW51f3GKV2k32rVZjD+mObtf
d3BjLockAHXY2hZjFPoED2m5V+RoZ4Ut3yrPzk6yuwcNxeX6U2weuiHMkm+s1XlC
FNDyW6M5nvtrPrswvZYV3N85FVoSzrLYGUzLwzuqhYE/Q7MPzr/sihq9aY7Sk9bX
TdNmxt0NRjwhOj0RulsY2WryExaFhnh9FmFTJ7J3vdS37NKqBvKnTYJtG1ttbI5C
S80+fHTu9kvbB8P9aLdfoiiorDdkW5QS1KVP57lJJq38kM9bpn7GhhwqHHvrVJ9S
+7O/JZ15DPeDg4ditVW+JU26iEvV9XckaOK+OOUvlsmAwbuogrX+UpmINCsY8v6A
FTcZH+x0aNMDYmIxZpY0CEAH64X0ckWCn+HCgq5WanArwsBwYZt3Z2yi4d6ie75o
1ztELUFxVc/3Vcz+M63QZ6YxzGDvpGpvWCeOYaS28zUIVJZqer1w1//cOF/cpcbY
pgEIAJOqXkzBGHC7jd5QQge+UNEAmbumExlIq+Fqrfuy7aw+S8Kid/OEmm4zUog3
AiG/d1NFA6lFcTJ7ThHq4qKBkRhFoKnHcXX6SXcXMMZtPz4c7QzxzKZW/qLS7eMR
pswVEa50VBk33dJkkk4AFzvarYW2d84LVQVgn12Lf4BA+W55VisRTZP7jRHClodn
Fha9q6kbV6Tl0YPV5ty3Y9XrQZ43aCsNAcexanhPZ5Nic7U04UWwMQmc0P2sRbvT
5uSotIkDbLqoWcZWS/QOFjWA2knUVq3xREeKCBK2Xn/6HFl0h4pXZPOPES4NnNCW
hBOABwr7A0yMeg4wYT7Nx67xS7nltZ58BbGwjGQoiYTeEz82UqYAAjBTAtq/cTBf
6wJ0JkL6ApJsE0oxjuHeivIERcIgrWcp8x+gKmsvAWUMoQTrOo09WPuCDd4ajAAW
QpxQOFkJiseUOlbGZZF4cE6j7CKAMXV/2num40HWYNK5WCe5SqzWovG1o4Pj5hBQ
JwFtUTOlLRU+ZSqBhfTDRCL/9QgLgmIRwFryi0WmIZVrHDPEbpAMXS6jOz00aEwn
mA/pWZuNE8OAdfs0fIHdgPewDr46X8Cb7LmJKA574xW1KZzK6EPaEPr5Nk/OCxW6
0j0LQSZwHBwNx2hi9Wlz4rrQ5/SOfPH2XdcRhjE6uSqkeJpC9Kbi5FK9gLqNR6m4
2QRd21iOwefrW2mJPo+lUkQZ0oA3F9dirVCLaRwc3mvWlnzHBurDc18EM+16VYmB
ak+opUwi4Tr3Da7jchf2W9X/TQO1dWddpLZAieDojo+0u0qUd5/zGnL8OBU/B1NK
egbbLQsNILVdaDtxm7GRSA+o54CCdWICl/Gi35fhUvU=
`pragma protect end_protected
