��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb��N�9��8�
`J�t�+K}=Y��-��.�1bSA/�\�1��Qr5>ڇ�֑����#J)�^���l�p�(�XiP�q��m*����,\�j�DYk��f�%oxy�ɘӈ/	���4`m�$��7���Ȍ�����2��$��:�>&J�����q�j��I��S�� s9c����֓�&u�iI�N8�E�;{��Z��Ԍ��l��F�#���V��od�yCW��I��F���9�HN[r �vE$
<���������z�B0*��p+��އ�li��0*6 j�9-kw��4�1Qr>�3}��sگ��>k˰(���w��w��/JeL�N�vNr4�΁4���ge��SX85u���z��rm�����Ӷ-BC�aF��E�uT��N�Ă��z�~�6L �1��;~c�{(���3��p���}r���ޠ@��&$�b��-\� s��Mi)a�_HO�y�(���i�Xy|Q�e�Z��� ɚ������JP�7�I�����F�����H����[8�;e��-�@,YVY��~�)uN�G9R�3�1,
���M�V��8��-��]�U��޲��٧;���Y!Žc�jd�.sQ�y���Gh�1T*���\�{��V� �\�&~��ߨ�c(���1�t?X���F~�ԃ��ܒMk4d�:�ϕS�k
V� ր���u�B%L@"{$#dH�Gz1�^��<���V�A��u-��:ѵ�C�
���A��p�J�ǝ`�-�^��������*���&�nB���� �Hj�sw1Ħm�1*�}���8�q� ?-�PMf_���f���f�<��(c���`�,�&=0
��T7�}Uӈџؙg�ȱUM7ԷW�P��u;�����h��@~5�Z�V�+�~�C��H�*��[��#,2qU�� "��|���5�։�|8_q^ߐ������k��	��2���UP9̶_Eƺ���%�pjyh[�}d&Y��և|�{�.d#	B��h��_kpd�Gb!vf{<���\��������H4ڔ�/tX@��<�ܓ�Me�!���z��qX����m�
�/��7rd��z�Џ��^>�cZ�n�b��CN��e���\�[��NBҽH#�gJ��߾u�"����`&?�g�K���)SN:��2��pyN��ܕo�s�t����@2���z�����3���λ����
�ZA�6�T5x�:\�z�b�lq�Y�KY�IP ����#�7�A�8��qC��O� <�  �OR��aR.Hط@5�{���e�G�E�{̞�/�Z�b�.~�W�$��oN��Ɖ]k�&��&-�o���o�b��{��A�%��N��Y���i<r_��Gq��#TmD�Ϙ�Fr�tʾ4�עYt5����(���	7p��������ynõ��=�Z�=�֣0��w
���WU*��s􃔙0rI{f|+��V����G�+3ηۼ
D3W�&��6V"�!yo�?���p_�]#}؊u-8Q��j�'�oJ@�|06#Y�Xm��7���ϚU)��@$#�B��Yp�5�dkKl!$1����S����tB�,<��K9�e�y V��ȧ+��_��a��0>1��A(ᯅx]�����4�'�sE=(�[֘c�D��r�����7j�	J�G0̫�;�,B�J�&���Gy��/��˻���Ki��p���Q��PP��֡%'	�4^#+;���O�J�����:f�]+PJ��o�6�'6����v�`LLj%W �����$���Pi�]MRCR������`e��s�h:b�]
*�!8J�,�	�B���7?����{^0�f��U]�(�^��3�Og��)ثJ?��,��i��U+��o��6��tg��\h�!���1����H�/a���"�Wx,��,d�ޯ��qF�ݪ��E����!M�%�wR\�a_
���:�:��[_3#�V���#X�)�G<
�
�}�f:�D��7e�����X��Nwn��a��i-������%����Z�8M��h�E�jv��8��pJc0��u:����R_Cv�X�����!�2����'�g�:oi6�lz��B�V����y���-�zq4p��0.����tN�1Z> E*L:��4j������hD�Cq%�u�I8�"IL�Կ������ùq�����^T��W�^��h,�%�����e���b�7+�q��q��΋�����*q� �����Q9 ����񒋉n�d���G&x{6X��i#�haѓ<��+3C�=��z�ib���QHՂm:8�i���CIШ:F(���y��k���v{��#���2v,��P?�+�Ꮉ3�T<v�ї�n�tE�GD0��#|Ol\�����on-�ѭWՀ?��k��;�D���~�h�K����/A�@l<�]fWr�BD#}�Òu��Fm�&��i��޵��s!�ʃ�˚=+F��ǵ&� �x��HR�����) C�"��%!r}�j&�)i�;�~3j7u�i��&�1����4>�~�����Î�b l=�&�\bpm��8eE��'[�=25�y�7��M��L��2UO�ټ�Y$�����m����I2X:v9�-y��Z�9O���J�a/z�>F�dZp<�y{�"�ͭO:�s���݃�ZM	k�v�&�:/��	J:��$����Ƞv���6�|����?����Wx%y3�R������RS��5�&�n��2�_�SՅ*S�����|W�u�_R�pmX��y/������C�"M%ʿ����XRf��(���x���9X�a������'�e�F�k��ݘ��
��Y�Ʒ�c����%�7�X��zk��^�\�;E�p��|�	��/���kcy$(�j���b�n<<�������*Q���#|�{��	1(:�q�}�Z4m�bNԂ�i�g����y��8����Y�@�VZWQ8pr�
]̓�Q(H�g��ҴA��KXx���+pU��UZ
QY���(>	���|&(�mA�֫@����s� Bu��8���Bf����{��3A�k$Q�t��������^�w��d��ԟ���^�1B)���z��֘ k��}C:���_���z�0U�vН|mW�-Ӕ&�]cE���6��a,u�r�:\��v�'1j�+.�AN)���<��A�-���`:C�ZKw X�M}���?�Αu	F����\#6�M�D�� �0%��-�-o{ǁj�g*�̫;.+:�i�"�����	�A����5ۤʽ���SH����OHz��I��
��_فIʧB"�c(ȭ|�/Z8y��v �j��%{Sr���?�
��G8���$��hS�Z	RF���U�a���8��<�A��$��F_Rs�Y�_��V�w��\���-�.y�=U�̡y��T���`��ߎD��P����iO�ﾺ��v���lGq�]B��%=���a��d:]�z��p�oP�۩z9���.��k�b,�%�245.-��qqR����O��- qW��(uH�WG��a?h7l��l�����G��� � �3����򉯹u�\J:l#�t=Epu�g�뺛0��
��X��S��Є�R���M n�r�:@Gj�A�g�?@�A��jE̿���.n:�󿜹�����ؿ�mP�d��D�����֙�t��8�߽�K���;�	I.Ө�]��E�|��Q��<�DTk��:����z�/'�qxK����h���%��u�\ ���?�E����Dd[��1��
��F��ʹ��Eym���L.�#*�*���YH�X=�K:~�����S�-?fl�����9sU3�hR�b��r�B!�;mq�kC`��8�&�/j��ѐ#\u�W�ĭ�W�ק����m�Dig��Da�l���[0��M�=��C9�W��n;����kQq끇\x��e2ｩ��;�_ץ��)%[��*��Y>�G���Α�4�'��N5��;z;���d�Z^<�A����gUD�%��J'e
�f�Z@�⢢��պ�������4|#م�tZV���!?�Õ�l����R�����l���():��_b�ȨW��r1~"Ե
gD������=��z��Q{�@w��4,�]h=l���c�;�7�@y����Nk{�~eE4�t���,Iۻ��e����m��H'T7�>�g�5��)����;/���v�=�ɸ]Z�0����"�X.3�eȪb������fs���X���ٟ���J|x�nܑ�� �|�'��&!-a��O���ŧ(��8�gγ���Jb�E����&�FL;5s-����d�n{��1>H����]���\}Lu`L?(ZU�ڜ֛]�MJZ>��`&52������0���ɳB]5\�~ҌnZ�'�^�n]�B/����T����0��뛚�V��h�g��b;�WL!�A�vbjaf�s�ss�jB���᪄4���ܥ0�ʖA���b�I9#�f�X9:���b?@��-)z����?ǃo�����Q���[߲��"��g/Om ��G2�}lٻ��+W�p��=��)��|G2B��Ơry�_�N����u�!�G��_ P~P�pWl&�go��͋�rͦh�gҲM��6t��8�Ϝ�c�T�V��[M�:3X�s�z	lťr�oB��b�^���{�\�P`�p��cD�w��25����Y[�V�a���� )��<�'���7���|o�lx�jc;�E��Tc͓W���#�$��E��Ul6�q��0�C�K�JH AO��~�Ʒ��Qѷ�'j{�r��i���Ɇd���>��0g^�icLYAr�ϟ]��9���p�we�F@O�xdSk��'���!>%S�Q�+wWc�A���!���SD�]#F�:�a�|n*-����.��=b+�Ia�In��� �T�[ TJ��_�������ӭ~����YU�F7�����S8a�G�(�������ӧ]b{�!be�"�6)O��g==T\��t�"��5��.�E���o�q�����d� �ĥY	1�;c�����~)��4к1!|��H�ѷ1	����	�%I�]@|f��gc��D�'Dʙ��a�='�̨5°����L�Ӧ��إ>xiz	Z@h܎���RxB�Kr�Ur6�F��Or�)�vE�Q��$$D�z��8��i��o%[�.��D���Lg�(�8�T�f�/�Y�*w7fB:/Ŀ����哊D>IM�����|�}���dܷ;X�%���E^��H?@y̤?J��� t7ARu��qiC�A�Q�߳V���+FBO/؂r��0�	[㶋ϑ����|	)�`b��/�|������z��B_�(��	�c�lL��2�BP�"[��C�?�l*
]I�>�о�b�`Ac������;�מ��p(�՗¸h��������fe�Bw ��;��?������)e�MS+��?�d#;�-���.޿���)��:��� ��
����p�'o��0t}��jȖ���w�so����:~�ڹ)[ɕ�V7���~d�5��E�\T?)SQ�a��w;�}�h����T�,큵���9��`��nZ佨�1KQ�	q��9{V$��j��9�Ѹ���UQs�i���UA��5^���kY!����?8�Ξ�;GMI��3�W�DԴ���ǎCAPn�Qd�	�_�]�o:�#�_a��@�S]�Q^�[t��g��6���h��?Tq�1�k7*�.�R����s��]�
��u�H��"h��B�}��r���@�a�
V� ûL��.!�;0A���#���vR{9�a1�����`�f�6��2��8I�S������*G�2��:�-��� �h/� N2F+�f�^f���j~��R�ۦ�^��G,�&T�qJ��k!�n>��?�cn��/������3��Y�a���f>�p���1ģ�tB��L6�'��ظ�1#��d쟓�.�%S�)m�^�� m�����Ї-H���W:&�b����,�S_��-y�����9(psd�Z�"n~0D�R���T	#(~^�SI�Kc���I�"��u�Ev����+F��J�O1�!!?>��y�t�sc��>EE	�6
X�%]f1f�@�2�CFVN�`j"�D��įfK={�!�)��ߣ$��;+�`4v���iވF������b���i��4�5�p<Lu*C��ya{���P����í_ی�b
3�[17)iy��i;���Y׍��'⟶�u_�*���}u��.�o?óZ |)�`O �����R��D���E�.�/����Zsˆ)�S��Q'�q�p~�7���u��x��{>�P׋1��AZk�5��b@��o��$���1�%��)I"'i���_d���VJ�m��)�p����+$H���zyBnD����+��
Edك��)	���}���;�z77I��*)�W��}#1(�ݔ��ұ�V�gM}��E�K(q��1}����v����O�}�c#�됋���+��r� �wnN+�����W����8����ݪO��?��ՠtg|�X,]��%��/�"V��	7S d�]�-�/��)��a9�+�gI�M]+�m�
;e��2�9��fƺǧ��Z��I�Ñ�ܔ����0�D�P"*�5A��#�ŐPc����1T[��tq�4V����ڙ5\6ю��d��>f���0+Zj�L�ìKp�#|�q� |��[�Q�6�c���&[裹L��IbGf����L�n����j��$�*�]���hx���,|�R$6��S<�g?Fe7d�s}�0��ֈ� [������Ⱦ�82��!��4�U �ʽ�@1�i�Dw!C3����f�ͱ��s�{�F%j��gmq~�cB0��%�R�\^C�MR��H��B�X��8~\J\��DZ�$�������=1��l�ЌU/Hڛ��4��j�PY��4!�E��Σ�rS���#e��Zrc����/*�Qa�U^cr/�6)u5���x�m���IĞo���Z��-���C����I�H���#6�]�'z�]ٝ}j>	 Zy�:���6;}��F�_i�Ǡ+Y���!��e�ԆKP���`�,�y����#��w���ۻ��L����3�Q&{M�����1_R����+��-6}u�>��+��I�%"P�S�)�5j�R�Y�nA9��'x�'zm�9{���^W��E}0�������ӎ��^AP;ز	D�U�=��غ�+~�9��-PgT�GQV>lNr���/jm_� 6����NBWm�����Y}-k3rrƇ�A96����h��Z)��ַ�����^�@d�i�rrC�N�|:�2�o;���σ���F�c7Y�l�5ܘK"Y�ڍ���\Fs'e׶��aTv)�A�y��\�o�$AL9g�ׯzճy����3&�oa�~ҡ����3U���[h��)����[
�|s�mE�kB�
`�c�����L♠��C��YV�i�g�����(�.�e�ӣ�e����\5ha��=���j4+��>Y�����;����yc_��V���M�D1��QT�I�5%5���{�%5�����f�n <v!��@mX�?\2�?;���y*b�:��p"����ʧ����i~B���Z���4+f�.q3��[�o�P<��X���t�s�(�¯53�X֓���� �٣�Y���X���=�&Dem�$U�B�,6E��?����3v�)tz��/���N�ތV�7�Tu�偈����k4��NV;&:)��(��B�g��gb��Ե��s��<@'�z�I�F�ɳnsv��<r���h�oXX�C�Z��(�Nn�?�T���-����y�C���^6���x�xSf.��q�YAV Tn�ow�q�C�g���^�p،PΈ��_��\��2��h̉\�]~{�i떏�U:�����>f�@u)�,h���٢W�$��6�0����� !ɝ���Lhe$�)F���� �jN6���<��s,���l��"Z㣂��3r�
�}OU�����Q|���TWD5�*`��O��禮���,\��Z����hp��8k� m6�I��3�+d��.���kb^u�9Ts3�4�o���D���gN����{�|���+���B$<�ޗ,9\��"LD|Z�Q���ߛ��߅�O�^T73z�ԅ�7��%��3���l��#C�࿞7�/4���6������f�xmN��%u1���9��%)D���ԦӠ5z��1�A��"i�ܪ�9g�>!0_o�{��R����l��Cz�-X��7�O2_���α�M�X/U�(n��$"�f�J�:x���R
���c��0fK�ǈLϵ���z�f�8Ʀ'�w� ��W�A����A��4�U�Q�/$�3�UXR��`\�Z̈́O��[��P%��'A�_1 q#|�XI�8�bft��S���}'�o��2��w%	`����2mc4s�F�q� �!$<�}���acvms�Zt�Nu���2��"�cem%���Z�񮴙s6$)�s�AƩ0��ͦ���&��Ea���/�(@���`���wB�\Y���S�y{��Lf
F��~ ��WQ�2*����h��u�1����ˣ/��g�M1#�+t��(��r�^��!̵34+H�@�}�LR��2���$�G$��o�0�+ojӱ�&*��b.�L���9Q"'��N�u���(��2b��ɨ��O��/�bN��Ax�YG:p.�g���)Z��.��6}�CHjv	 *��T﬘D������k��c!.d�G�W��Jm�Tau�	}�����0z����_Q�#~�V(KA-�x��|� �v�Y/�`ȅ��Q�k	�����à����P�}�#�#9=�?��Ѫ���|T�y��&�ט��K�W���U��&j��v���_�N��u�u�M�򮒂ˬ����g�T$en�4���:5q6bR˛�x[4���q��1ҿ�j\'`ѐ�n`��A����L̈�7�6p��Im&QBی�u�A�@�WY1�a��]=�o0�������$�@�B�+�[,��O$g^X"w��e?r�"˧�W 2�$�S],))E�<:��������k�&1Q�{�b�ӧ�?[�ߔ��V5`^�_?N[�4�`�Ka�6T�7��BS������l�"��Mb/�����8�,:��+,��W�ޮe�LE�B"v`��G��b���#�#��h=�_�@��S�s�y�Bй�~]![�ȱ�O�"{�1��q �P����O(��ϒ�S��֓�7����y�)�0����q�I���|��<�w��,2����2�AW�1��H�7����ǘ�!Z�۲����XOr�(�{�e���U�X4Ԕ�O|�@v�{A(?�K�xH���did>� pT�yu:�P��&qH
��Ғ
����8V�/�I�XY�9}��������qx���,~xL���}תW�KN��d-�(��[���r�z1�1R(�V�ɬP�`?�d�!���j��s
�z�I==�8�����p=�T��#{bZ %`A�z7Z�t'�� ��\���ZNM�nZ�(B�n�.�Q,'�v+�Θ���${q�&�Y��
��`r����]��T�n$�@��m�FB	���c@�� Ls}�ԸAV�Ӆ,�!����.����C��,������ �����s��r�����V+��,]���f"$*�jΌކ���Ҝ�z����DD�$��EЦ�k��+�e��v�ԓ����4	ߪL��$�I���
��q��(r8�==�U��o3Q3Uf���VgD�'�@�{j[B�|�_����2�fZ��ʷ�rX��p5�86�#�����+�m4#D}��|ڨ�B٬K��l}(HPύ�L>�1&�d
�os�;��F0���CئjV�ɊOql�hhc!���PNxu)�8[s�m{3��n@���s�,����,�b��3�c>=S�1$;<�"�BL� ǅ�0֥�D�吏,ɒ����|%[sh�A"6�����k�0~�VT�Z������6> R�֮'!��[sl�w�'��k�_Ʉլ�N�0r��O*��vm��S�"spCU�3����Іg���V,�������,�6a���]:#*��7ߋd�6�d��� fl)#��+� M}C�q��[�@Gz���i%[IJčs{N�5�i��o{c��X���>��;ЩD�ɉT��n�����|S�'S����&�**!W����5󬮾�r��j�f"��R��\��#�tQ�cN����u5��P���d�sC���ƭ#_����(&�� ���?��.�����㸇iP��	h�|8au��C�n7��P�q��i���܅�*������M�I��Gۚ���ɍ*���;L��BrM���DgQ9\�d�B/�R�o1��$��[ϗ�p�.�R̎�� 3϶A�(ӷ6�y6���q9��g���.eY�0�$l#�{Ic%����G�Wr�h:��c�������cS�u^�ש�l�-�U����+�B[~<�N��	}b�p*�~��Y�2��V���S��_�T'I�
���N���F�/����CA��"�.Z�pm� >��j������`�`3�Pmn06���ظ�D��֦�*.S����/%:jG0Gj�v�A�_f��ìK���)�&=�����Ĥ���D�_�h8���!ÉZs�u~��5Ŵ����.��h�a�I�P�0!��X��iNւ_��`��}>��ӬC"����}�I�&�V����o��'nZ�u�P�D��wħ#!`ga7��]p�+�	3E4�+;g�C&���&B�N�Z�����'�$μ�^@�"/�P�rx`����� �-��f4����"K��G�����M�����&A��)=�Џ^�~�FH*���4C.Ź/���S��J����~�1M���в�Z m��`a�hMG}a:$H�%��~�o8� �춁	��'=��Y��jM�s�s�A7jŎ���&?����P�c�����!�?�������\]���F�7�m#�p!����½�I��tF|�ZTL٠Q�YRV?őy��fZQ\��~�V�1Yf)w���?h��5�P�T�ɻب⮺�d�$tSYk+R�v���F!��Ӷ��'uv󱚌��1�e%�Ϭ���A�z6�R�ǣ�&���H!������f���b�
WFw5���IBɬ�WS���)cRZG�ֽ5�T+F�Z  �����iȔy砐�A	�c=b�@V�����i��iv����\C3~ߞA����'8��(�-�!��C���A�ы��3:w|,K�^4Wd��dڷ�bI�5�e�������G�G����Q���mr��A����Έ����y��6S��ĥ�a:`����Ky`���k�i�|��oN畼[]i��v�����"��;�~5��v��i2�t%8�h��I号��-�#�5=	F\�/�=߄��Ed������fy�$T�����2+���@��gEȘ���bm\
���8�����)\�[Ԟ��zr�qY�Z�H�������q������:poC����x nsϏ�yYte֓N���H�u����z������3b]�d8�V�;Ԩ��P�l���X�R�W�L��3�	PtY��$�E
,�8�*ȇ�4&�#�ٟ1Wf1}�-7�e	�l�m,����bouV.8������@��!, �nZ�C�����s�v��Ac�����5Ax�H��Ť���\i��.w�w��q���e+q����o���F+n��gH>3���r�NY�?����1��ɓ�����;N��&ڕbc�M3@��$҄�!ؘ�T{u�Z�oR��q���5%7D�O ���l��E2�شىYy�����0o��uG���[��5�&�7;���Epb�d�C�C� �X������g�潂*�]�z�7�Mb:.�w�3�w�ʲ#����?�n�tX!ۿ���wA�`�
�/-���KF�ٜ��(�}/ T1ip�\�����1�Eu�g��ڷZ�2���;���ЦZ�S�L�0�W\د�B����4٦��*���;L>{l����������.?z�UWw��'�Ogn�KHw����4H�ԼY-3 7�"�-mt� +��g��Q��(iV'���:���/:�����>����O%Qa#�_��'A�+�Ul��=�fR�z�*�S��$6�JNn�\y4����$�3:�ʓmE��	j�[ �w��9xQJ;��n���%	�2p�|U)�n�GD��'Ͷ(�c���IV,D�S�1v��\��W5��.^*�	,]�:�Y2<n�}N���2��i����dܝ�+��د��ФI��\���8BB"���䩩����ێ�	1Eܬeg+i�K)~4z<|L-
WOY�����
�Me�p��3L�C權�;��@�L��C�t�z�x^{�)�|���l��q��]��o�Z��H��Y���o���87-d�D�"���u�jY	i���r��,�$�Kg�<*o�suL�S%Ҏ$Zy�����Ր%�ԝ�$ve~{��f�h�S��z����8/�բr~��ѐ=��_.��( A���6T��S��1p#�/�䷕r4P�+�>�<~� .��tǠ/�3�S\%;R��a�V�H)��Rأ�0���L+��jZ����q3�kes��O=n�k+���pv";����H[b�Wy,n����<݌p��cW�
�Gy+c%l��WV����r�����Ct*���-��=
(�B�5UU��D��ct�6٢�0?����-���ͦb�6����e����/�0pr�a�z":ڻ�04�3���^a&
�]���7To�~,'|Dt�oޢT�ʓ�����]2��tx��ۮ�n!�t��Q[��f�v�/k	[���s��e>��c�����f2�Ib{�^'��e6�s�fXT��yY�:]�|Z<�K��Ft'��RF�-�3��O>�����QM:ܺ� p�v8{uT��<�'��nm��?KC���sH������00o�S�"L�cM�i�w�������$\�����s38�%��(o����9����P��;���5�����##�(b���'��W K����F�JЉ�� �� en2D%�:���Ǖ̸m���+i���*�P�?��8�x�P_�_�`*쀫a�Ҋ�1HW���%b�d��:^�������7��j��C�=
Bb�:�bky�l�7�%��c9�DЖ�r�$�k���D6�pC��_~G�5چ����R1��`T�	B�U��/j˿Z,;tTd���=�|��o�GA�5�xO���F^����.(8��
K�}�7�T����F��)�]C���[5*���`� xY�8��i�8S�ۯ5.�s�"D�gQ ; �U�7��FK����\�Ѱv���uܽb��i.ʳ��󨾻x�e���M���Q2�%0�oJ��eɱ���"XӒ���2�E(���Fd���1	4�A����d��m�`��h&��j5��M������
��R>"5��f���QL�!�Ǔ����;
"������}��U�'s2����/a��'y�t�h�m��*!F���m!)o�{#��o��a֐ E�u ��)�Y�]�qv�J����J�ӳ8������;�0�)������Zs��6�!�*������7�6ɫ�:@3��||���h��~�_�~�[�0`�2E��eHom8��	l.}\6���y�&ul T*����NTN���>h�[g[�T��Dq��\/���<L������x2y�T��H֓��[K�?���J�29�F���C���8tG<�����ڂ�r
�-^��U䬰.���!� 
��|�I�8J���u?�^�Z!�_��.=�.��S�b�o[.����_@�'�T��W'�Rd���n�"ϸGZZP��S�}T����.t������O��_D�)4w���l�AGk�4h���"`�:m�	*�>r�����N{��E�v󦢂���s��� ��3��׳؀{��εRj����(��+��BI�H�Gt�;�JK�ت��%tb{�=��8����e�j^߸O_1��k�&�Jzܧ�v1���J��:d���Q����UFMt@�q毣%Xgu�s9����T�ݺ�#�m�C�
�Kv�ɶ��W ��bʡF��kl�e]˸�ց��/��s%�F��׬��h9q�L?	���n1j��֙�Lf��#<;��;���U�(�"`��T�Ң���G�Þ�&��襔���_�]�kz~�q�L�[�ġ��ˇɕ�L���?S�e�l�?�kq����Ē���z���
�Y����s
+��w�h�0� ��^w�n|�����A�}O�����X�z�+�͏��w,��Ϝ��T���.�lP_�F�K��/Z��R,��>��B*����l�8� �G�F�3(ݐ�!�2=��݋��Yt��K��q�(F�P��Yt�Lig$�V����/��Ҕ��a�\�k5��EA�]�v��A۞!W����� �)����s@�Q_��+/��9�,�<�J�!;�8�����;�����M��U��.B�㟬������)C�8��6���bC�ã�2r'�-3ɂ��(����V-������
�y�y�d�G��&3�>r�(��O����R��Ʋ�j�eAUL
����`1Jw��ׄ�59�N��@��J#�� l�ֹ�OL
���ocֿ�p	b]�J��2���@�_�s<�0J֕� �kyN�}���#�狎\����+E���8��)�T�_�8� R����ȇ	�#!�E�Ï�I���aWN��&��7�5*�J�
<�k�A�������!{��$ ��}wUEx���RعzE��-�x3����ǵ�����Qv�{����Y��@���D��KQ�m0�w����DV����/+�'�Qr`�ZZ��hx8B#x�xSHl��;[瀡י�=�4ب�IEE�͐��4�9�
}N�%��A�:70�]r��P�1YP�4��s�'��B��
�>)� � =K�x$6��@��Imp� !|	�@���{���C[%LP�k��������x:x��q�dnr�n�2kr׫ؓȅ����|g�p�22����V��9$s2L�B+��X?$l;��ߩ�S���	Q��ܫ�3�f��IF���gO�T��Z�[��".�A\��V��T��C�@�eh,>;�	����F��ys��t��*|�!@.�ˣ�/��dfsS����T&sF�'��K�5���xk� j�nIa��(�ݽ�:�P�s���&�9'�t7��
j&�s�9�N�W¹;3��]�f���LL@R�K6ڪ��S��SZ��M�A���ʅi��w�2stK��[���x�n�<q���$ցZ�,
]�u�;��F
is�M�����:�'LF�K��3f��0�i�����ڪ���Ц�,��;�#K�Fb]E��_�(�>/Ia�!mz�+�Q�M�}y:�
���3�IN]�`fP�0�+�%3��N���^l�	S��u�U�M�%U&�D�%�{?�e]|��7c0 ?��v���f�ya���1�ǳ�O��m���w��K�Zd�S�d827;Z����"�/i(MQ�ԟ����͞ �SeWuo%+�0�sh��J 2��|<�Q��ueo�r���I����`J��Ԥ��2O���M�a?^�E&�=}�B���>�+\k܆��p��1;��6.�����(�}R�ď+k
��0�S����p�}�Vq�������
=�(��)b���*Hb��g��ZtI~GJ���e 2mV�8 �[W(�qp�[��u�g�����K]����	XF8�Ŕ�����~�֫�4�=JSᯉ��p�{I#Hև��H;��ʤ���#�Ht$�9Y����X����m߿�����8�M�#]��՟���݄o�I�g�D���b��>�8P}�)���;	����2����bD��7�CVh�v�0�(�_�k��_4����s�R��Z<2A����ŉ ��y�KDߢ7p����v(Pp� ��`4�����Z^�
���.L��~/=����_�AS�*.�����!-���0��^�<Iƥ�p���U�hc�z��x�ij�l��_f����C��Qy�-��\I.��t��U1�c9������ f�ii= �'I�� ��`w�J�G1�Y�~�s�xP��d'���a������DA�1�1L� ٥-Xy�|Z�h���WP�"{����"v����KO@�oR��K��/m4��L�{���g|��*�$K�h�_��m��f���GK:�ۭ\�gWti5�i�ˈ.I�UGF�S����%C���9�#4�I�5�0�������t_΍��بgDL=J�"$}L�q����'����݃$n����FP������"Zd��C�^�&H&V C-)GW�۽�Z���2��b4�8q�~����}�]�_�"E�'VW��14��BT!e�W�=/���uB��8
�\���3P�K� .�O�>)U#c���y�i�"/u��]��u���xW9����t}�����m-4(���\1#��:�D�����C>���Y�`^�;���N׶QJ?�������3��f�?�[��� �Am�vѝ�Z9�t������xG[�)=ƿ�+�p��=��+m��N�1<R�B2��I���E�~�┾K�îU� ͕5ث��V�
+���+�޿x�X�<�LQ@}����M���<Ƹ�E���F��o��hǻr��o| `�\���"=�����J��H)^�3:�Ǆ�<�H�o�Z��WԜ��o��Q�Q7�oe�tb
�x��� (V����)70�ܟ#Z��aM�"�v�55}��f"?�vh�$�K@�4�Z�e��4�K�N�x�(�rH�UF=&���
H���d= ���P�����?��K:_s�X�I�:�����Ja3���KF����9����@���a�>��0n�x�w�rc���O����C�pe#��@y��ls�\~�h@ +B���-������P�˶��z=(L,�v��.� k"���PC�B_>ނr/��[��Wp���zx��$P��
��Q7ռy���kp��� ����Z�����J0p��aJ��Wz��0gk~�!�ӊFRi��?'���#Y)�uA�H��ȫ�Xu���1����m~��zQK[�1wKZQ�?�x �TzZ��s�J���M�<�V8����ZK�3N���uН`��,:Ħ�3
�2��� �0�s8���_�;����R��Pҋ"K�̇9�m��zBHAE�h�٭��+�޺�O���Rj�J�n���۸����ъ�9U����&����n6��������T�3�a�m��D ���0���&a��Â�	Q����#P��2���޸60w(���e��b��_B�<9�(���je���,��DՄ�o������.��a��q�7�_����&�Ȏ���
h'��9�p9s��+/��*��d�J����9����������6M�I��r�7ʺ���
ꂲ#�O,�S��ʦ��Q1� �f�ں�k/տc`
���//7�I�-�0 �֪�-���m�����+�M<�'�]����BLĪeY�:c��xy���haK�8�[�eR��j47Q#�:���+�ʂ�]���ks���홓m����@3��>8S=T��0_ ��Ai@�VZ�O��x󤗮g������\�B���tۧ	�������Ϻ����\T=�kw�3��cP�E�E�(rS&wx���SB�Cj�G7[�fۡ�Ɏ&�5�&[���a���v��3�VH|�+�!�����n ��D��F� �=��dR��NW Eԗ�m�H�]3#�Sx�T�g�K��D�gZ���~�����A�����O�4�T��i����1���d�!��ֹj��^`v?y�j�P7�>ޑ��B��֊�t���_�Iow�h1C��t�����D��ߪ*�5�B[�|�e���� C�5�e����a�)KUc���7�hۂ�0`8�/XLhUY�+S�3�tL!����X.� ���s�E��E
�/��.���i�p[�[R��9�>��+e>�e��ih����U*Q�ylS+
:���~[���C;��� �цx�~�M�ۥ?p�-�6w�2%���	�i�Q��2�r�}q�{Ws�+j1�����'�?g��'��k�:�C�l�+q����g�_��m�����FP� )���:�P�/��Lެ*�Do-���V���fz�	
�W<�>V�-Ջ�Z���$!�)!��Ă��c.�hͧk ���Q��S}7��B��y��N����KS�[h�� ���|Z�PW5oi�lr��d����e�U;z �hex1�I�t͠&MI���NkR;HYˈ�nN0���<P�5�[��������gvhFT�����H�%�m�Zq2�xѥ�\��X��>+�ۻ��i	�W{�&V*U�gAy�{]G�Kӗ�i�W��Ba]/Z,g�#NL��Yj!F����Y]}�ݼR�

��j�
��	ROIP��1H�M���s���(��c���6vo4NN���u���!��_%��@����C\��d�x��1I���&�3�� �]=�����(5�G�����	�c�V�㿃�$`='(0(��	��H"�M�^�kH�H��C���د��R���ei��K�ȎC���b���?�������[T��_|�W�����-�����mn�PG��	f��DmS8���UE�F�	�>X	b#�z*��v4��Iugo�~�zmKW�-�7���Q[;D��%�8�³���a{jeZ̞�� �,5+'��ڹӂ�����<Q��a�$��@��L��E�:oǹH��-n��
ᱜju���^{��ۈ@��}��1ԁ�9����R��Ps���yV�o���~�F�5�Y瘏��|��ײ# �����O���Ae0P�V�?ّ�e^R"��?�2&��tyg��R1<��)<n0I�$�oz��I=����Yܓ�#:�d;���	�]t!�8yp�Uƣۭ�~ �IELO�#�9I�vL�8��ŋ-m�xd� �ZZBn�K4�;#)ڶA��8X|��ƶ����)?����G�9}�W�����'��}��
�-S�c�<|%��4v�AXu�RJ�X,Uc��D�O�UN����=@��1����,#��9��fsq����-]D��������=f)1G.���BTs��W1����j]|���,���@�#j�Af����������/��r�h��b4R�\���������.��X�'Qb��?P��^�n���qY�Sq^6e$�L���ǣ]^�Q:m��w"5EѸ�h��+g��7f�&�n�k���2��U{d�>���1�x��>��F�M�SC�&��� j0LZ�����R�P���������a�!<ϐ?��'�������T��+�;��`������Lf?B�t�N��j�������n�R>'u�f5�y��ֈk%bR���,.�Ό��������Xް�x$�5YY�:��!�gr;��[�C�����y��:��疜=����I�<�K�<��_���l)�EJ���i�c_{,�|��ՏXN7;�t��jѸFιhP�o�G�˩�҅/bxm0�	��@&��wٵj%�{���su.��븠��S����|!�I���۶{N�fxSF�h���&d��4,�P75�����蝥���������=X�	kҐP
rq�z�u��a-�յ���--�/���)&��;��uZI�3��_�.Q��ӟ�4��r/mP�g�r�֏�����PԈJ���<W����V���Z�)�[c\��H$Ő����6�D3ݮ���F9 �Xg�`���w�ɡ��cڨ��^�� ���mxGmw�܄YI��=�P���і��3e�W��@�(�|�M���<F��m�x�%e���u��sr܅�@6�¤0��GT���� ��t� ��v�GVb��J�W���֏ޖYJ�����u����ٻ5��ι��1y������ɸ_�y��T��'��fp�΄z9ںݵ0�֯��OX�$�h�Z�s6�́�%]��������`L1	M����C�V���3���*��x4���º\P� ��t���RU�B.rr:��=�o�L�.�y�܎er����M��;�(�_[�*2��-�٩�C/�����P[�)l�RV;˟]r7��2�e	}�S�$i�v�?�:�s!F�y����^)U5_�:уk��	N��,�qtW�K2�Dw��e/�,m�ZV1�-n�F.򌘥/���1p0���Ð4��n�P������w��z��9Y&b AF����V����1.�b�(\)lxPAg+�mՏf��FdM�^��Yp,�W��q/���"�x�+Q�����mfP�D;'VA�~TlHqBh2d%k����"_���D��`/�S�Ҫ��������#e�m�X����ؗ��oҚ~��j0ؙ�=��L[WpUf�/�8����"�a�ut�����b�����1�?u�g�<oh֕���A_�H��3���P�8�ԲL�­H~68ڦ�ɕ��K��m��}�?�Fװ��꽘���@�4��[������B!�%���0����Z�~�����8����F�m�Ox�C��Yg@���+�aj�酺 �[yR���2���	�T��ټ�j�`/�e"�LC{���*��ԋ��0�l�Ԣ��������(1�xC1 
��hW�����d�S�4��2Hu�)����ά��J�2P$ђ�+����
'�(qK��28r;�����"-:{mf~�M�$8�����Зj
⭬�L[����q��կe�����m�<�,�H�Uu�	)2@�{�T��z��O	�E�VH��%S�W�Ct���=�ڣ	����]i� t���	=�F@A��[���U�P�D��� ���g��~G`��2���hH��0>�"}�Z��e(a$ɜ!i���y�nF�޳*�Jt������'�8!�g��5�[&Z_��lI}_��m�2�t�uv
/�������T�[$�H
 �VG�~h\ú���b=u�tZ�e���,]K���z�B��í�ڇ��Ys8�X�W���%��ќ3�N(35���O{�	�'�R,��Ӧ@1��yp��&�=9��bf�� �,d{��Yo�(�u�KY�p@Ļ��1�)��>pp���R+]%��KD�V����q陋%�ðw�F�,o�1Y4�TH5.e%�����Qʘ(q[}zQ^������{�b�<X�JB����t�琫�!�f=���j%:{e���'W\A����r��EI��xF��}��[����QD�9�W�!��	sA�ƽ���.���uc��͖R��4�6�����-�2%��\1��ۖE���)��� 8mJ�
V�/[&6�8��1^�gh3�ʴ�v���������,7!ق\l��1�Oޑ�j�����^�
L���I�ߦ�%MC��y��-�?��޹�QP��H)0-�f�K��r��1��e�&�;ޯ=W4�����ɩK8��W������qW�*�}������R�H��y��<�-�P��+3�-E���}m}GF.S�kY�d����o�hts��jI^�)��[�/����})�|:da��=*C�=��|�{5f��FD���l�[i�^�8���ha�7�D/M�Nt6�D�O0 F=t���͠�w����?#G�2�
�?��@��B�]qw9/<UZͧ���Ij)�0$m���=�Ed
>��%W2Ɛ����}�is�
YQ}4�11ՑNԞ$D�aL���q�f�ٺ�n�'�_��|��\�MT�)h���qiU;�؃��Ҫ[|�Qdڄ(�lj����i�x
^��9�H��:����2�^��k��$�� �HZI��=
=��������~�:�wz]��A{�/b� �8�~.����|S:�WDDn?nG�?��(g��b6�e�Vy	�*�Ƽxe0�hE�~����9��jt��L����>���	�	� U�\n� 5@L�U���Ë����8l�����1eTO��J�=V�`��?DO�<5$��\Z�N%d�>�]�⢓|4��g���eکXu/*�63b�3T��5�#���Z�8 3�t�'ĒA������~#�d~�2(k|�`+�A"�*���c�ѧ(a��(K`�]�DeEx�ݽֵg�:����m��~�����e��1F#$��< d_�d�|�-.E<���Q=���+�ZbSZ��{�Hx�UԉǏ�9��&phv�а<[6%~;Ԩ�4����!p�|X��_�9��E� ܔ��r/�=j��.U���\ɕ��dC�ѧ�+o�9T�a�]�m�̔r0*�n��[�w�wo�i���{�	{ŴI��+��;�K�#B٠PI��k����&4��?�7Z�ٳh1��oP���Vj�s�� �-�p*��,�U[H��cy��.����_�+0���n���)��;�W��ϯl�A&(�-��N�۠}"e����N�b��eI��6ň*�׮�|��hNՌ�[�GӬ%����	e�]��e���.��+
|G�0c��L� $�*P�.[+��6`L�m~v<��M�J ŏJ	*���b$�.0�6&i�;���"�����@���5ճ#��~JO�v�#�����:�u!��VF���#����'��o�-<2Oh�2:�Λ ���������M���(��II{��au�`��>)�����&��z�B�"zit��1��D65�v鼐�+�#*�����Vn/'�k�6�#D_.<���Zz�����9]Ik�����jv��_8�g!�2����#�TWz��4o(tN�t9��$Vͻ�����|r�xÙ��5�jC߆d�<�����^N,&J	m줖�2��k|�I�DcyE	3Vϼg(k���������t��O���Ey��'Av~b<D�9;��Z��ڇ��|{�pK�9�px��Q��B_Y��.˄���WQ��I��h�z���: i����\�X �lwq���Z
B ��{+S���*
/*�?��b����M��yWߍ��:O�HuI�K-X�з�M�ݐ� B%�LS����*��:�x��y�����I�V1ߓ��+�yήB�U��>x��r���T�8R���j��"&�#"`H�U�8��I
H�j�zΫ}r�\�-I��b�ҋ�,��<k���߇q��Y��N���K�	/J��5>��ER�N�洜{j�l�Ez+B�ॺ�����q�&�(vu�~�|��M,���m#��$n�M�� R���oj8�K�4ڷC"�y&>��F�ef.�d�����W)�����e�"t�n��OQ����8��Iǌ�:�$u�Xr�QN%�5wJ��ga�'�gL����kf k�%;�nR���rI���O˓6y}�Bo<�ߌ���={��}M��.����,6W�վv��O�hC\��O�ֻ󐂷dwT�C��։H����Fc��4�s�𔓸@�յv��ͷYvۧؑ��d�����"U���W���D�#;L������z����<���<�_x�~&r�����sd�F�.�dx;����lZ>!7}#~�pK���$]F���$����F���~!OF D�[ 4��`�^}5����@(YuϿ�>)��)v�?{7ߢ��i��ܲ=f�S���{���&�c�'p�����n��(�$��M�5�%(խ���@My�X���ä��@	>�p�t�����A�%;��O����qݗ���� ��@has�a^���9���#)�ݐn��:I(��H�=R	��5}��P�gT��Uxv@QV�.�`����)>�Gt�ĸ:��t����kV�/�nӂ��o�w� ������N�F�t�[nѾ��[B�d�K���i3<)2�x�]��5����9�x�k6�7�9�ē��cf|���U�ά�$��ng�=s��Z������<��%؋�j֬ԍ<��ڐ`8Wݘ�tw���E:A�p�����)E(+��^�G"3Um�\�v�"CYʷ�o|�x	�ꈡqc(�+s,i��<b���"&�WF�4�5@C>��Ґ��N�=��8内9��-!��o}/��w��Y�M[�w���pN���Hό �G:��� ���{�< \�#0M�ۻ;�Ӿ|h�@P���� ۊ��~��zsx�v��ӱ�p�?Ex�) �-���������K=fRN�6~1�ic+&�����G�I�-)�c�7�6P���?���|T�
�lJX��A:=P��+4̀��_)ӊ�i�
�W0����:.f�fɔqKR'tkV&�*�*:�JL�_�}И���ଖ�vZ�� k����Ҷb(�^�\$A뒢�ߘ}{d���	�:�v6���O��UϞ���JT�h�Y9XфQo��hAsq�3��|t�%E��7�?��#V~����Vؑ"E뾜������w�i?Q��3J{D=!@��c M�o�9��b����B��}�4N!�56��P����ef�����.q*{z�<t�)�^\=��������ƒ����G%����h�M�X�:]�Sz&��o�P���L./G��#�<�Bp�@n����"?��-�ħZ�	�Z����A�9qXdP�O��v�B
3" u�j�����r��9ɣRI���p>q7#Z���=��n��I�z�Z��p83��l�0�B{)�ů���P���W���6O�j��l��<�tej\b�g��J]f�!�YQ�;3F41_����J[p��a�D��y#�����������ޙI�|nv(j�}�O�G{dv��AJ�}y@��ۡT��%��6N�̮�_J�h%��-��9��{��Q���
�+Fӈ��a��0dK��ȍi*}J� ��K�V��h�x]�K��Q�����;�:����ss�+%��*�X,g�Z+[��J(�mN���>�P�<u]�_?�Zb�{����߽�}Kk��]�1��w߶>�<�;�\-se��@<�)�;�(���Y�oyQ�𼰕���D�Ǿ⯆C�>�2XOk=`h�ݛr�ai���uj��>~Z��¤��	ލ�"���oП�W��ë���=]�yY�852�k����{2|���urZ&�� ń9XY�x�4x��ps[�6������⥵8��ےh��Uh�4IJ߫>��Zl$f���pP�V��&�+ 'l̉�k0�EɆ�\=R�eCvy�F�}�����Uc�Ƽs�Q��f������dJ b�\ٚ�?�^!ʗD�)%�������)+���[��r'@�S���%���zb��K�|��'�ۙ����pU_��B������f�=�eN�Py��+5�ͭ�o�o��p!���2RfDL �fP!�o�n磷���Ƃ�I-�;51S�')�}���0{|�s��|?���5#�*�~W�A���LӌV �
NI}=��lEb=E
�KP|�,���ѩ�<��E;zޣi��>9^"�_��gd$��ُ~�>'��ڥWRU�b��U[���Xg�'��!�E����p>[��	/	�N�yӪY֬ \iP�?���^8�bE0�r�	oS�RX`���R�4��y����cS7���5��lc~w����W^�	~�j��i�<0&C
>��fMK���eĚ�l�_"���p'�4zV!�!-�Qۋ�/�~��+��Ax��	b�q�8ᮬ�G��#�%�{��3?_������k�����IM�s��@�& ��H D��S,r� 5��v�����F�"�*WkM����vbՓ�e�^U�`��g+kchP0jSZ�;��a��A-���|�$�|c$�̵�e'1<���$&	�nOu��=��}���S��U�+瀛�V)�1,{���a�/�[��Q���́o���A�op�*1�������W����R���ha|��5y��D
#`�,E?1a 0K����Ԩ���]��k4Y�lİ�IG��q�|���jw��([�2���<4{���\h�٥c�~ϗ�*�g�����$�	�r�yus3Vg�Ю�����a�'�/j�)��vH�y�k$"�)F���[�dҴ����և�|��������<M!M�F�)��ّ�r̦Z,��8�@PK�T'Lwi���s:M�N2�=:�=/|
E�~��Ǣ��B�%-��N�%��;Ý����=:sB��h�n�rM��,�Д����IH�>�MХ��<�P�eA���\q���Fee"�8�Ya�Ά4�ˣ�ap���IP�]��r��绡*z�S���W�+d��RP!_ iH墩���c{@�}�#����O�u4�t���Y�W�Z�)��� +��l�������}R`IB�37�������]�s��p����a��Ī����qO,XK[8����=q��y3�p�_�6-���%9���-V�X���>�$5��R.�E���l2!����O����S�8iy��D����Q��J>axE�#�`=���V���i;����b�K#�,�tMb��PiE�2?�3U��������Uk����'�%4Vc6frq�;�P<��>f<>��F-)��N�$�$�L[ Šk�ܦPj\�RV?��AHG����Xw؀&�s�s�Ew*kZ=;�4$�G�ʍ	����[�Q��� ��d��m�q|��=F���ǫ�m�3f�[�^W9w��"�>Â!t�u��x���N�H�R!G���,YQ�48�modV���$a���-�E��Q�(�p��쳟����F{�e��g�IR@�9O�j��.j ��m�E��l@���t����3��+���ę��C/"P�p����}O�<e��-錓(P� ���-"=�6�l=�L���R����H���q�Qh=����f�n����>��w���LI�|�M�%u��M�6��J{�g��E�	/�譩Z����9�"ױ��dH2���ġ�3ݨY���cYg�?�d}�|��a����3+���<���*�.,� (�A��O�\j��I{~4�,�p���-��-W�kKZ�_�a�������r?�1�n��D@��4�$�luL��Ys��A��W�fr��A�X������J�zp���a/^zQ�)F�v*�c¡Ȟ��2c�]5	?�ҵty�%	��$���^a�E�//:��]��"� RP}P��[�F�*�㷫��\���JQ�BF�@���x�_��ě���KK�W��Z���+D%��]u|r�E�T�N�Y�ZLmg�����e#]
���Z1�
N��2��a�-뉘�Nw�j��;@Ph}_W��*��F��8����>ş~k�ê�o|�g��9�w������� 6��y��N������?X'�9�gxΒ1 w���-�0b����?LpB�n��P�����rZ\�4��U��'$>�h_<En�`�� ���_����u��A�$��4��	�?x�4�qvv>T�ȢQ��V)����zoe�u�ş��w��67�x�]��>�x��B��)Y��A+/:���֢ ��ܟS�b{��K���gπK6�����foN�	{�8�O�x�[�SIg��3q���UiTF&<|}Y�bx�b�X�8����j%����)M�+�S��K ���N�ֹ"JM�(=�[��q]�cψ%��C��RLA�
xNP�|%&��%����,���?Zn���@��b�G*+�ưp�R���P��������S첞~����Qr�p�6�\�+lD�VIǜ_	b-�ڭF�\+�N�2��W���`O�)!V�T+�!����
��� G���.n�	�b��+bwZ-��뱱�
=o=�z�/��s��,��^~W��Z�bkG���	�[���8P�y�ʯ8�@�O���A<�bz�D"�n�P�L�I�5#+�<�3w���<�/�dl�b�pj�&pKl=�ڰN/,��yC(�Xr�~�̉�VK���0� ZJ�(��=�qjG(�W �ݞ
ܒ��4>�����!��~x=�洆ƺ�%V��^�:��4q �tZ�GtWU�ǻ��>X�����2WD�҈s�w9�
��V/X�|޶$�TTUNZk����7`x��%Ȏ_��3�HP������� �|�l�tQ�
=�� �{H<�UӨ���,r�C�+Ŗ�{̤���У���Zr�{��<*�Hk�C�w���|���nGrtn�:�&�dTF��Co��Ǩr���c|��ݟ_{\�������*"T�}�7�M��@j�e��M�,3��8�vl���M���i�ݾ�-�i6񼕊�{��?��d|�3u�������������Ѡ�?��z�l��3m�@X3]Ԛ2nį��hCT&���UJ]:/iQ���̓
�,���f��� �������c�BI�y��0	:�AՕ"L���V�ψ�q���_���z���Q ��BʥE�?w?+�M�%��c�"������`n�O�Op9��H�b�Z9OUd�e�TV؅���L[�mH�")�&T��`g-$�u���@�M�2�xm��r���z����خ����.�3p��h悃$��A\L`��d�-�U��9�Ze�\�!�=�ʓ����l�K�v�������3�-N�Ar&4KZ�D�Cҩ�
 �V��/�.��v�%prfZ�:l��R]�JP떥�_�JT�3)���d�'�l��v,X,�L|� 2J�E��j�ݸ ���zf����-��&SU��X�X3Iüp��şx�!Hw���g0Q2չ����x��=�a�-)�q�U0�֘B=os�1:����	sc�y�|�%�^Y�X,!r�wG���7�>���B)��o�.�y�6��<5��w�
v��X ���T�d*t�+7�bA��oy��Z�B,pF�m����z�[vt�(}��I�R.�y0�h�13̐i�E5ODń���5��#*����WI��c=�v;�u�we�&�Î
3���F�pl����%R�J�IC����Q�"�\Z��iB�(r�÷�f q�=��+�����:)� ��ԆV:��j1�sEsY�	�Ґ0�(+[�^��ac�i�ѻb`U$��Ό M+�	>�A��_6I��@�1sb�E��Td�� ���ﺠ�u�s�8_��m��ZtxN�cď]n��Sz�O������n`���O�h*KH���W��Wq0�o!(wO{��w� ��m�k�J� ��"���3q�v�cQ߶��B��BE��!n�5�CH$�'�w��F�a>�/_fSn������%f��Z�T�A�p������:0�dQ���6��s�*�z�5�;���5��W&��U��/�JH�7����ͻz{���~�$W�7��g��DO�� � 5�# �n9�0#y*��%G��,���=!�ǿ�d�T��t�"FEu��7߶lP��`�?Jp.�=��`�I�T_�Q*.�	E�.�����>p�z��(�Q-���
�xf��+��J�ys_��������`��B_���;�H��z"AeFH����p3�ͨۚ9��6!c2��d\�ݎ=��\���ծ��<�8ɡ$���:t��x�R�>�7.{�0�b��a5�5��H�}+1��lۀ��FC� N�	z3�J[����Z@��'	������A(״�S���OD!��{�0���n�yJh��\"_��S�����Z^�l��B*3�<������[K�r��?��U�1�@] ѻ�5���O�ᕞbx�ȮXv]Yl�#�h��t=��z�ݎ:%��$suF$饱�
m!A�{#(�ˣ�]�=��;��+�H�2R 1��3�n?�8�`H߿�x=5�D$�8�ո�����o��d ��d�?��R<�I>3������q�����"P����.J&��)*)�m̏��f#D�2k"@���S=��C���[Eb1��6l$a��l����]qf��9�i�`UK�؍y2u�٦��q��F��+�{G:��)?��yŉN�帠��l�J��i��\|�;9J᪕n��"�Z��Z;���桂�,���b9��$��SS�a�h`����Ä��Pls� Ô�D掭�R��4�b���/YѼh�+�v���� �oV<�50d`��j2��$H'Z!HX�#�`HH44&%6�A-��@=����#��;nM����rm'$��]�7�Y���8���h�Z�w���eᐎ�º�+j�W���0~�,�)Q��R�A����=E(��m��Ã�g��A�	˰��������y:�6�@�;5��>Wւ�Q%������A����X]T����p��]��L�W�ܱŵ�o߳��EG��$\�g�d~Ǫ�*����[�1�:�¹��6/���
Y�����8�����k�:��s~Xo��9��8�e�������f�I.L�z��"��C�Y���x��g��z:f�`yAF��2}w;�ҜJ�?��T�=�?'1��C��nZ��2Bb���e�j�34��Am�	�/:xf�ׇ����!1�ACa��E�C�k�`�������meQ��=�85r��V�q���{4	����s�.����H
G���#���؁���urE���g�.g
O����1��}j㳫kNtv���vW��֕,��Q�G#�.^x�|��+��� �uh)]�#K�?��&�'� ��M]w�3��z�{*��_�;N:"Nqa�`-����x��c�pm��l.�mK��)���N�*�d{"�+�.�x/4]��pǩm^�'���=�IEɔ�D�kz��^<�6�@3�(4M�W������X]��8��N(�V"��y8�e�� KT�.����lh�p����KJ7�?`F�ƨN�"Ю%9u�ᮡ�� ϛ��P`��]H�mCmuFt=�
�C��#����[�hp��϶�]o�zA�G/WG�Q�{I�p�YO�˺Z �P���F����@�D*9([0��M��I,��f�t�=H���w��φ�T�����!0a3 �킀�p���[��C4�4M�0��C/k�g�Q�A��9��wy=��s�11}~��K3/������.CL{�')9
�̬�PHv���PxJJ�:LG����{)1j�G�����Cj׾;k�1�E-���"�2@��:қ�9<	k�Z���ם�?a	Z�ٍ��e:�9�
^߽����k���� �{��C��v 	
�rA�F��_�_�8�ͩ&��hST���:�h�i���_�Atc�T��e/*�[J��0��ic����cvu�(!}K(����#�#k�����b�L�Z�hV��t�R/Ƚ����~���9�j>���U1��D#����Ӝ�"���D{�j1*�rs4{cǙL�n�m�G��И.l��P5��T��7��ש���W+Jԇ�8B����,�VL6�|-,E�7�Û״�.?��j�z>tT����_�� ��dme��p�wRw9�l�:��1��K�����W���	H��nN���D��|:��S�/�7��C�V{ge��!wfi�oW�+���t��
U���^y�@ F�l�F��ö�l�����(b�'�#�U�w5\R�����>�P��y�4,��4��"��������>#�������P�;Vo���2P�&���|%N�V��>�8��<\g7���'�[�m�l�A).�[3qU�Z����ی��u���Җf����%1�����9�O�<�,e�%(I�w��Jo�:�{��jbC�%?"ژS��:B��V	���zZ�m/���U�rQg@��ө���awn�y�x�Dׅp��鯓r�wF��nh�~>�|)�3�K����hq�= R.����1�A���R�~S��c�G���K��k�X�fts�)xϹ݈Bac��ךV�u��ЃB;�X���������_M8��O9��/�!3��������u�1?F���`l�����>B(�Dˆ�V���I>�y��X�I�j���=����!����D��p��\��T&|b
���!'�.G��1&l�&����{�/����t�`I��������b�ѐVb���IQ�NO�чL���sa���Hp�_.��Ԃ9o��d������3G�����r	[��"U���*]q7��$��}]��o
!`g�B�+�]V߫c;(&$�/�v|?������D0!nە��;��l	���������-�6�$�Dg��tJ�BU�S��px�a�K�$=x��0&����O� CÎ�b���<X[��~GĀZ`�E���=ǿE�hfu��������tQ,�mT���{�⁣$�C�}���lܡ������rRe�N��;�+.��O�*�)�{q�U��g�-�؎FQ`YA]h����6�M��>�7IB���&�v7���pȏ_*;�2i����5�Ҋ�NX?�Z��5�N�%c�_�<�ǣP�r��!q�ˉg��h�[z��wݹ�d��\MQ|���B��MN��K+�^$�>�7�����?����u�`�b�����,�Jc��Ȳɹ7/�`�SF�j�o��Ic�ƪ�^.n*���TڳY����G��	,�?�����Ju؇T�DV�����X���z�b#D��8c��U&��z�5�O$a6�d�QMp�$�ɽ0�z���VY']w@��"[B��ڽ�34��{F�"�_�EZܞ�M���!���q����!)4ӛ(if�õ��s�ܞ ��R^��]v֎��Ze)�"�@l��컖��6k/���h
E��CF��lzD�*������Ql�X+RAe�47�����U�X֑�Cy���K:�sR�uU=���HUB��w��e�]���_��k��S&�
\�<I�{�
�k�IٶY����?r�瀎�ۑ�e�Y΂~�U��X9�gq<x2!�u��T'M{�؍���_Q�d��#_q���"{i�7����8{�r7��;l��<�:cPCgg_�/tK.�d�-'*�N�=!r
��G[��]/R�*_�
}�!3}��8��$~��s#U���c���~a�������*f�r�x��q���1�bP�Ax�#08�1],�(��c ��,��D&���j��"��R��~���*��o��P��I��1�v��)b1��c&�rA��F۷�PN�>̀5�J�Rۈ�:�%d�3��=���[5���I���׽m�{�S�������"S�V"��lc��N��kL��]�(�d�J8������]#k.5��e��b���(�c0�`�O&��J�sy�{a�vSq�����8�X,�/q���{T|�?3�Fh�� �F��'g<D`1M����|$o ��1u�1Cxp%UL��T���4G!��u���	�|gk���/�B�kET��db�c:*XE���/��7�o�=�o��l���E\R00�>���QK�yNGA����t�]�Ph.�~N����q.��}�ݨ�Ra{|#������%o�v*o�g\b�Қ�����[c�f{B��}�k@C\Y��)A�y�֓j�н~�@��d��7]��JS3­|bf_tQ����voj�벐a�Y����Qz���� 4��G"mt���V���ЋƳ~�~f�2�����+?�1|}q�R0��>)~�YD�;kEӫK���]���Jŕ�e�>~b��^��6�@��bL��5?�Y��]C��C۰�>�t�Ag�y��8N�n]*���}s>�[v8�G��3C�s�쐨^�?�	�)�W}?t6@-��2�P��k�Q�Θ&-�Bw��hGԄ:�Ű���b�%�U�y�ga���ɶB�3�:XE*�)Hn�I_JU�Mh�����#<�EƢRO����̟�Ϝ�n�*��ӌC�d��;5:$�)���0ͭb�v��|��K���wk�6J�3�,jYup��q�=��ɛ+�:�E�o;H�<�G;�!'���j�3�xKu=��	e_�)E��3PK�է���*�2����,K"
��%4[�r�>kERo</%c_�{�5)�8��i�Ɠ��˰*B�c
�!9�&}�Z�x���o6^���9�OP����=������h��{	��F�n4��2@��[mYw�2P���R������	נ�����=n�I�%�l�lU�u*:=y���w�+�� &3�����hǖ�ɶ�c�	a�i�۟���0�uŵ|K��GK�ѿ�6TH9� .�d>�K'4j�GY�a��ħs���	��q�P~˺	~�����b�YZ�M�ݢ/8V�V,��R�x�����恮-����
�%���d�BRe�� !�	v5�·nB���G�/佢)�X�tRi?���C_`0�U��JY�Vb�c�+E��V%�rF� 7˿SǦ���9;�)�9�'E�^-/���z�҂"���A�9־/�h(��tlQ�h]�6��m�g�Z�F�o�^ђԶq�١��A�� ��i�BN�S|.�}e���*����sXќ�Scn�-��!i��`ɨo��EG��w�� 9���V�̀�����[�FF�!>Yl��}��a���׼�09�������6jU=JO;���%�ƨ͆U ��	�q�>z[y���v?}�`��a}�dIj-	��)�D���C�b�H�ӗ��^��&�S����Ym���E�*��)�Lec& jn����Ԧ1i\��6�3�+�+	Q1�������U��$5�{c�\�[4�H_�Z�i҇�E�(�ey�{Ӳ�0MnW��i�[�)����{:���z2����:BV��\�����BΕ,#[@RaL�}�zދҺ����a��il;P����oN�7��a@EEqX����~�����7b�Sر2S�bl���ȅq��;G�'�#�fJ�7%a���O͘9�D��%���C��H;���<T�� ��&�����i ��������-ӜwT�V;����~���dy��X1�z��wv����� ��D��o�>``�s���q�nBJ�B�T5Ie�\#v�K�P��z��w�O�H4�D�:D�T�;�JJ��J< X�T:��u��d�(`�z�J�o�X�4>j��D57$P<��'�>�@�>��@�CZ�/D�KV
db����dA"C,���Ld_n�G�Rb]�z8�9��kX)�v�`�Uv�\%�Ɨ���V�yų�����-�J�AoIpX�3Ƀ�/[i�">�(�>�[=yک��S������G�އ����;�_�p�.ۂMJ;���
������;3e������'���A��:���(CW�ox͕�\��I�v����z�u�/���#�]��s���Q���6��U�v)��%��'g�d��th�V����g%����'��'��5�[�Ĥ Re�2�Q�q+"��Æ|���	?�R.��������v��`B�����������4W�7��g�� ��Gf��{��M� ֣�b�S
f7���!�i��Y�����0���3*'>�F���8���&��1by�ր8�>K�ن,�e��#�ap���L6F�
�
�>�iB���M���,��gD<
ewOU� (OQ�-�e�J�F���e���S>�A�b"���"������S%_�6J;���'����Ez�?��kέ<�����;��i��3�J}?%�"N�L���]��.*�>����U����w&�b��H���&���,�J��|z���-y?�������l~��#F�SRCI/� ��mpEd���þ��⩿��C��8��Zf�`� ���k�,�>��;!A�`v<�W�����R3�iaL�0�MS<��_4S�Zby��6���>�S�	e�]v��DR�w�=�y[�:P~���N�����dBzT(�;�[%����7X��3���a������6�Wj@Z�U�S",%�Ǽ
��~W`e��T���P-� ���NҋC؁�o��ʒvW^jU��t����4K^�wZ}�Uj��?����nρ�|Ͼ�i�z�4_QP�>���E�X�y� L��,J�y�j4J���� �U�Q�3�G�
�D*z)���_��������3d�5��֫���4�`���Zl�.,U	)�v2
��݁�nj��Ȋc}Υ����S&����^�v-�|c�1	X�����ahh����VZ��
.Q�ډS3"G�Q��>���
I��=`\�������_� �%�>����
������j| �з�Z�4!O(8*qt=�s�H*�?�g/�K�V{��k�� ��y<e�� _L�,��U�f�V-�O�P(���IQ�AY��&��w�Q������o�F��g'���a�q��mʹ�B-IQt�7���u"��4�wu�!����P�K?��0��-�7*�C!x;*�vI���({����+��gC�\��h�g_�%l�����{�����o���9��Mo�'н��8���*{Z�_�4����:&��I9&��Z[&$�k��ޤ
4���O�t�~%ZmNF��OQ/�X؞F����n�^�e���u��Yv��Jy�1b�7��!NX�~)�� U)w"�
@F=@�7�mL��瀭�{"��qdgx!�M�SP�Rm�Fy!������vZ��b�A��1��#�xxu�+t��bv��;��0-��kQ>~��w��`4_��.�e�8l/��χ���X�<S�p0��c+�Y�r$��f
V��0llA����.�%"�?�
T3��bpG��N��F-�y��b}o,ˇ�0E\�+��o�޵,�v�(_=�1%
7K�E�)İ#L���=Yl��MqʅX�@��>[f�ΊD������C${�w������stǡ�/�G6���_tU�5��PQ�A;}�$	�m��	��n*�!FђPG��G�Nu|8��M�T�^\�wo����Ą�ig��Q�ڹ�	g�#����>)Q�h4R���oQa�nD�V�^�� ,xj��.Ƶ�� ���3^�^B���9}a:p�+N:q�����B^����%�Ļ����g���W�O[��?x�oN���OF���Q0i,�?��{��ug��4��Դ���>�^���Ќ���-ce�ĺo�L���HN�����㗪��}�M���{[IX�T^�[xf(�
%5:c��eC��0=��DVۘ��:'�Q_M����|�|,Vd�_�Jc뚢���ѹ�����>�'"g�&�j���}W��[|�v[�r�2B�`m$�_�6�/�r3�ʗ��l�'�ޱۯ�s���B���:�(�#X�L�ۖ]e���o��]����z�V'������vLЍݞ��?�q���D���y�Ը���`b�9z�= �����_�Vs�V�ѽ�8+c���_Q�$�����^e���Qΰ�J~�D~w9�|�(��)�o>r,�L(dq��Ԁp])!�:��K��F�(}A��:7��G�vt�fܕ��B��P��l�\!��^���kPILC�!�:�-��Ȁ�e�q!�2�� �j���($}��7��K�}�S�:��ɗɵ}�<j.#']���pxt��(��X�}�6$[Iޙ�h-o7kkԂ��p� 9����/[�Z��%�$bA�괩�]�t�s*���-��E7�,	�k�Ƕ1�]y�;F1�o���F��Iޙ�ܺ����{�B�X�R��^�������y������ ��7��?�
�N�a�W�muv4��-�zH]tm��!۴7����a������7��^"���ANŊ���X4ܓ��W��!�X�$������r=���U4���8�m�:dQa�ZI�=�,��^A�G����y��e��|��n/�h 8>.�I�\{�׌y{Y��^��n������0��'�:�e���J���Sb�����C:�r���/iۃ�TI~��V\\�kq7�h�����y��1��8�VK�O�		4�P��[�D��Y�N��\�J�/��Y��@��2�֩q�6����}5GШp?��Q�Zji1�ʚ�w6��9��_��oPB�r�F�A@��2�U�ػ��!T�!�v�ǭtZ�ҧ�Lc��.Bh#6�B�l�$=y7�z�d4t%j[�R��+��(F�8fݱ�FK��"��s��d h�9r��R*PQ��:E%�?Q�yJ�e�A�'��Լ�GS��(rOs�]~�m-ȢRh�����)���||�z��SL���D�ק�fx6�~@tѹ���'����v�-)�:j���t_طWd˚��JY�VaI�6��4 �X��6vK���� S����>�8�!� %�T� 7�?��2?�uer�\����(��tF���C� �)r�t��
��e�銎��QP��D[֌��� �d2��l���)J�pˌq��:���W!IS���!H ]��˼��o�lF���Ƒ;9�
�o����ڠI��*)��"T�eV�]�&v�^ؤ��K�:A  �9��Ǭ�^�A�1C�9��֌S%�$��{AP�|�0"I��� t4�_AKU����ʀ��:���9�F"G6�LE����hߠ����
��ai{>�(��Qz.΃5����F�Ᵹ<>~�qYHi������|��fӡpz��^y�#�@]�#�v_�}K`��E��ݢ�s'���JһVS �(: ���)R��
�Y>�f�{���'�a�/N����ժ�Gnd^Y*�9���}
8"�k��DY���H���a�ʞ�m���m4�:i�(�,M�R%�`��O��RT�AG,J_�r'�D����Gb7Э��V����/�!k����ߓ/6�|�Tkج��Q���C��dXs���s��҂�����lH����c	�?�Lv�&h�G�#(�3q9�~g�`���yv���B�6����gFVG���\+���ܮ��!�|����x,�0�x�=v����A]e,��y/��#����]<��1���aX'�B���vG��,2�:L�K�����2�܎|�Cj�`�B�i�xR;8���w����$X#�6slϽ�${8�&Z�S!������yg9F�6Q�e_ ����H	�W�� �}�F�5h�y_^�z�
�Ū"!���(�R��qj����P�9���Ft0�(2��di�����{������)b�35S!�2���qa�� ���s�r�������!lLߏ<�=\�{VJ`��f�'�ʤ�$M��L2�R	 ����-m��Yu7�B�y\�S����Y�J=r����g��̏�n�F�,u�'G��s����������Y�KoP�`U��*�6�de���f�����	(��/��pkVj.�?���I_�P��f���e��cv������Ob?�'ޥP~yN���-T3T�ګT;�͢.��΀�W�o�Kk��ޠѯ-7�w�l�e<�=>����/DU^�%�%}�R��v�뗃H3�C�毌\��/r\���_�"s��*�3��n؝��[E��!��9b��v6j0�����)E�����XThce"yWǀ�,��<c������|�B�4�kQ�f7��	M�tWpf�-!#�	x-52��9̹��S:�X��M��䕗���T+m�VG�lǹO�]������&o�bE�n���]%n������"_���7IR|�
�e�E�>V>��b�ަ�ӟ0[H���[g}]�H�7��"	��Y\��ʟ�Zc��-�~@V��	�@�4o��!(_-<�����e��f-���i�x;~9�6\6�4��Ӆ;����6��΅#���l�H8	�*m;���@�'݋�\G7���竫���ot����o�\�(D7���b�!�WK!���E��ax~�29Ou��T���1��f�+�f�F�X�퉛MG+���O�go ��r�ճ3��	w석����:�F�k?��9x5�N\�9��~w�]�#c魸�����v��-'e�?��[��� �d��@�I�+F�L�,?ă�0n��G�Z�
��M)���V�ů8���f���b01^��0D��}�{���U)iY�6�c&������
\�f�p�N)X���@��8@{WlSJ�<�Ï�e�:�h*($�����o)����f�0)��#h	���������s*2C�DyR)�g{S5��[^���2��0����	`a�p?��}p7��8K�ۦ�>Ht,�=�UxKw�Wz2�y�w��f[��$��	l�j�e����k��Ew�
�? �:����Ы�˙0����-��=q���hU���eJ��m��i)G�Z]<?u�cS��t�*T�mq�E�w��p}���Ԯ��;iީ>m(k�t���OO�_�v�.W].�AD0���g�G�[�^i!.9jS#F��Dl���k=�z�n�}9��S7ͽ����KG����h�2G�i����?2�уV��Z�
�^�xI��21��K�D���Z2��~؆ �gֻ�&���Gq�9s ��W@~݀��s�l:;�`���"��{��H�GѮe|O�v[��4����8�^�Y�������( p��4�����_��jy��* �～�N��Bp��C}�k�N�s�Yv���7%t�R��}�6=�Q�� �p�f�ȻX�	j91˼-Vb�^��ڢ��\�l`��J-���
REi^H�C7�[6�v�Oj�Z�?S��aM�����WWL�`��C����"w;��[����4O%'~����?��� Y�oY��Z�-D��{�=���o�.��� 9���Z���66�����!�抉�q�sK}�t���N��qZ�ÏC��eb�e��ESdo7�8-�
Ə� �5o�`��Ez��#20?�+���<���r>�l�w�%CX_���8Y�~
�UfC{o���;W�	i
3V�Yt�ZA�r������1�Q[�zC�������wx@�b�����L�A"��gԄ]�kj�������c�>�`N���4R�C�@�DGӒ8k5��03�/�H�36������P(�_�=`}��[v�s"SP�^�+�aO����?��p�2YX��,8�(Fa�V�X�!�=��q�F ��A�h��S~��h�t�1�y�W��e��LQx�D��v+�}��T��g�33%iT1����5x XL��2���¿5?����`����L,?NH��R�i1��i��C�z]{��t���Z:���� �*X�A?�ja	I��0�/��!�*ߌ~�yi.��'`E�̈�v��{�w��QEzg�O0���c/���wM��N��Ya,P�g��P�>�k�,y� v���ڹ�'�(Ts�fV�N��]y�}G�P���/�j77�dA�W��"��p"_h��S"F��3�8�Ǥ�8��-_&%Ԯ짆k�T*TmaB��%}IuŤ U���c���:�By:r�<�����T(f3���2ķ��2w�'���js�0@�8.�x(K�g+j��A��rV�e�۔�<ZvK�`?�U[@�8Ggх9,��N��{��X����O���V �+���+��/��d��D�Q����1���]�UZf�=����& �]fjڽ�i��c�����x��l��^p��$
��ѩ��r����B��rx�J�k�-XB5�c����Z�\�1������D[�����K��I�����f*�����lPN1��w�9�簲6/�#��t;( ����W�l?�o.(Y'��ڏ��ς���j:l|�Fs�Q͌&�W��)�9�3���d�-K�
[y�9� ��1,~��!�~�m,.Y���N�n>0�(���jb���t�9D˖�]T��3��Q-�@B����L��+�\H�O��2�i�`�0�V,�NI�D�����8ɯ�^�̸De��m jޅ��~���t<���w�"��v���;���d��K=Q�I�
ubAd�"�^�F�TY�e�{������<(�ٰ��2�z�&w$�!�3$fvԨ�^��$(,��v\�p7ϼ����]��L�NFJI�1B�3Gk���׆">��&_��SrY� �I�d�)��S�h��K�n]7���_�&ElI	��N��WV݅'�f���i$��
���NJ�P������?��`}�s�j��0���f�3V��JJ��f�U��5-�a��������)���m"4������6��7�&7��0�h`����G�~eAn��Z.�~z��θ['
o6�k��"o&b����Q>1���\腦L�G�ʺ#��6�`fY�U��:����؏�dl8e�SryA r�y�`����~��M��D��M<�G�=�Y�~�1�����g>������oy�x�'���%ekvI8��]���$����a�*�ɠ�O�.ڿ��5�w�Lq>�>�7�c�����t	�T��Z��X�g�.j�S:vb��X�26� ��-����]��m�Vz5�
cת�:��#S�6���}b�c׽&�]�w��$?�d+U��z>��^h�J�wI�I҂&��}��<*&Ӡ��M/7{*}������-�ڔ;X�m�[�߉�:Cp~�מ�n��Z)�ľ��OE��}v�P�F���L�E��6�=�A��W� ��P�زĖ���)�)��ඟ�3��XP\��^�]�;A�+i��]=9�&��#��N�X�0~�į�O
��v$��lyko�z�U~�o��D����ڐ%�S�[�-i�	Ƿ'?QS�p<�A�;#)��yԍ{F��i���z}l��u���<��_�����J���+�S�M33��x��s��J���z�i�8s��:�]�m�<;ڡ�#-���\��Kn:����XC3[vF9�\�����)�=�*�����_�[|�`I�K�k[,���j�L���$��1�Mb�!�=�}6u�Q�yx3c���$,�#ң�b0Jn('�T�w�� EJl��9�i �Z���ser��R�Yhf�E�3���4����5�iz_oz]�8�L��[�ۻ���2,�o��`��