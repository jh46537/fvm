��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&:l�x3�[e�,.Ϛ���;v.�S��-P��P5��3���G�ℋ<�Ք�Ia5̲F��{F���'($���gG�>�����{D���0��v0qU�8!]^�3e�)��#ih�CP�5m_��{gm>���H�/�E<�"�s�IzD���T���Y�+e�a���C�gv�/��Ψe8	]e�i\��LRՅ�x��?���8���:K��;=
A�S_p]SI�xq�|Q���N_D!�oG�{
�2��·�a/ȿ�����X���UhE��fq~t��-�n�fMIW58�l�h�tȲ�+L�ݰ�id%D�W(v�a��X�N9�����.?�q��I����B�{���=T&[���2����c��9�C���͜�$��z7��m)���Z�g^PvJ�G�e+˥I[Z߆[ji�äa��,z3� ��7y�(&�W�!;�N��/Vػ����������*��8����^�j��A#f-�	W��G:�gmu/',K��=�q��&�2��Rb#���5i�F�vn+���O(�\����M�p�<�^�j5��n�#Nin�X4�x�|��> E�qtC/�(!��.�P��׶Ϛ2��v|$85_�ʗ�R[Z����PX�2�l?��P5��Ӥ�o܍gYyn��h��K#��B� �Xk5��ųt(��W�����*��Е-�Ѧi��e���5�F����a�q9��rN����������ĩ_6u3���v�7�S�rr&�o�1��)s�ɾGz4��F{��G1��F�����-�/i���9�q�����W���ȅ�9:l��Iz�u�����a
rD�O���B��9�!���%g&a����rWA����F��SH��+��X����5DNy��S�ࣾE �"F��^\���KF�(��M��~3i���:F*���.���%?�q��0�Յ���^ģ걒o�6kY:�	�tO����Ǎj ���D-�w�zߞ���Iiٙ�ȐZUk��Lf�녋����X¹��_���q�����(�_�r�|�����:
i�Jvк9g��l�~��H�v��&}�U� �F\�2��2�6������i-��ʭ�-��Jd��� >[��/fL  ��T��	vR�����+�=D��lE�7%��3M�
*d����V)��"�e�k;_;�(0�X'9�"���'��|�eۣ%��Y>��*w����C"hs�SOeX-������>�P_��`kt�0�T�0vv��c0���$6 !��r�j$Y��u� �
%>�{&��}j�Wd��<��SL���@��r��H�?��X*��w-b~�5u�ٛ�ƃ��^@�Sx+m�g�ٵ�*h��#TG��)�58a+��o77��F���H�����P�,���k���xo���L�a�O�Ġ��UPP$#�?'�����Kަ{8��e7u��j
����z�/MT���?����,�u�3�
:JK-$P3Y��~_���n��q�}���m�BEhy���I#����yv��3�|c�mR&O&�K��#�w��g�%7.���x�����=g�Н���T���W�:����b��������5�) ��&���=����p�8����G��$� ?<ry'�@@� ������U��l���!���%��y�;ϳՀ��#%��Y:���-G���]�
CplZ K=����TnH+Z�ڤ���DMU��4�$g�`�ٮl`�)�����@��(0�X&�Y��N �b�m&Vj�!��c�ۋ
i_�/qN�G�Z }^��[��7_4l/=u��$f��5����E�hk1W$���%�~�i�v��U�v6�{�n����sL��w��3���rc�]�����)��s(&D���YDC�l� Z�"�!�|����
~��JV�3��+�N��F$�$��Zni>���r}h(�E�����GDpƁ2���T!�%y��L����Κ�֓�Tӽ���-/�/7�ԇ�G�n�LY��޸�UD�`�xVq�]T�ʆs�1��#�<�������[�:��rOf^6�<K9�*JM�'�\��������0��m�.�ֻ����_U��?.5+�Ml$�i`� t!�N���� �Ҕ1�C�$��u�h%�ĖZ7 ��۽�Q���O�\��㌚}��+��۲��|(��d�c��-���4�`a� ��:��@lv�E$��~?�B��W�`&T���庯���� �hyOc�{E��t��O��a��Ƞ�iH�.e�b�{o�S���ϕѝ֢N_T;L:���Vݿ��:�3fWs�+E�ܞN!����
���!�����+E��)����)�Vw���x.d
�2�!R���頩R$��{�c�H#�x�� �o:�_pAZ�=t	��:����mX 1z/���#(0�{ȱ��פ$��@e�&����#�0�
�x/����
���_��X��"	�9�	��I��O��VB)�B2;$JF�6�g�gW���9�9o�������2�@$�Xcr(�,2�8%��V�r�)o
�3�k/K�'`�%�'�AǠ^��Lgϲ*=p�]QL����k����j�
yh�%�%��o�-�2�k�G�P�C��&���i��(���*������p��}95�	z���z��2��Z�;�x�Q蓟��w��S�4>#�A�'�_L�k�8e�q�~$[zk�$�Y������a�$����k) W��g�tX#W�o+z-��ƀ"*5g?.G�����Y�|p���O����7����n�������vy�?p�豧��G�n\u� g�LS@x?D=���v����>d#�sx�_i��ʄ�4����Vi^���J�we�:���M>⯜:�?��ܩ�K}�#�bź��o����{�9��Í*��|a���,[b)k[�&,�uQ�-��*��+ �
�m63��6J/�� �-~��8*�"T�kl��2 ���#���`c�z���\:Y�R#S�`D���sr�e�7����^�Ǔg (�.�C���薄�-��:`�ި��%C(u©�^۪�x�r�6�Ye���n��K������x��{���$��L���]WA/�'sx#��ᬅ�^�������T���$�|6߬�h(ƁKs1�����cˑ�"Kτ�=ڣw�y���9'���J��
cl��\3:®��w�H�Ԕ�u�*n��[��v�˴��:kZk�e�:�</��Z��kz�Le
�����!�5�z�^���π��L�R�<������4X�~rFثTK R`������D�`(PlCXҺ�[{*���,K[`�u�+iso��	�6-��_�ޙ�-˥��6eI��CImu��Vq��s�d���{�]��v�|d���y��Xx�In<�"�Ek��{C�y�3.9���7kz;V�;R�N\�ʀH�mZB��=����1�9�R-wP_����S�x�?����B!��Z���նI6V˹�p���]��V�!S1nj�x=f<W)/�%S-A��p�?���d��3����m���5�z��c� �[}����d��������l�T�$Ηc�ӞnewD9���
��O����t�y���])�@�D�&̻��􅰻�_�Rd��^d��f�o9�Z]'�I9�,LC���@�A	_�%	�cO<�?	�7S:��;�C."�#	_�%N��t�(ϸ�i
$%�mAc���K)p��M������D5ϕ��HqKLo��y����Rt���)�H~d<l@w>�B
35=�n���V*��T�}�WY,�/�d���i�e"��C�)�w�(��R������q�c�'����IR��릑}����w�B*�Id��7z����l/�U��5�p_AV�W��Jy(�%���U�P���b�l��}G^I�H
o�{��_E�����	B%M	}.��V~�e@�"� ��(Ȏ}
���1��Fw��۷��/�cܨ�눁'��Pй��#!�6����z��mM�~��+ܳQp��Z��Sm�&��,_�s�\��O`�k�l>ڷ�#������r1~�����_��w���ė�A��	4S</BfV��0�a��g�OrT�z�'��{��r;����w�)���X���F0n}�"�˭afyz�רOnנ�z]F�;=�,_O�=����-�02s ����U���r���Nr�h�R� 7�TS	C���Jn�j��)ML,gv�\��lW���v����$�3����tr���p��y���m��57|�<"�eυH��{��м�q�hY�Hp}�/�?�l�q��j�[x�����cc����:�uJnf���c����.o5�iO��&���AZ{/�$�	���I����c�\�{�x�
���ֹ9�{�Zޛ���Sh�������t�t�#�/�P{+�
CCՋ��Qf���Dr�`��A���sX0P@ה��`&%R./�6HZ�]�I��u��s;)�;I�y�,�>K&v���o�o�c�i�����4Ľ����E������Y��I,psazW|�\������ub��Hs����)���v�h�����=�!����Fέ�M}Q�BY@7((6���&����mQ�.>�_,N�)��D���Az��(��s�M1be��Wo	|�������u�twqp��<Yn%�4Aa�q���fD�%�=�f���aY�Z��|���wh׮�Hr���	��W;���8�cw�V��U�4�F_��#1�Ÿ�,��u�wS�e'�Ӂ}��N4r*�H�z 	mr����p��v��oԕ*�i�8�~��ϥ�B��/v���������[��9���*Z�Z����ո�ٸwt[xJ�a.�z�Y`��z���#�N�Z:�U{���Q��A��Q;SV٫#yz�%>֞��;���ud��V��.i�Z2��v+-�뙀K�Γ�2n�$� .��a�~kc���Ũ�,�P�:�}x[V�I!k*���(9-��*��~-����-=���<�d��z(&���;��᜹a���4��'v��1`'���YXl5M �v&�����mq,2�vR+L3}a+:��-r��E����\7tRh�S��J��Fó��Q��HC�'��㋼�xa;?��<d��:0�jbr���n�o���z|��%ɥ���Ey�

�%�N|�ϫ�z�%�Rm�c�oU8d����f�SN{�^�ި�::W��C�x�`Z���`�l���Q����2pC�W�k�����{�=�-�ڋ�i ��"vm�h>��@5E<�09�/� ~��u��v�(rL�@6���}"!9̍c�d�i��8f.��V&R!�Վ�T�n����Qm"��7��� OF�aL�q5!�H���oѯ��0�jh׸����e�mەL�<d�'�(�VT��0���a �j��@^q�u�2�צ}E��@��ܙ�#g���{�����U��s�U��|���Д 8��syg�_n�`n�\��r|�
Wsó*�t��䖹�+��:�)c}���`�P��&�5xo����D9����#m#���"�[i�B���.�Nι����i6�19�& �3V������`IP/l���א�w!#�g�3P�p�����&��/��0�V<-��P0G�d�ar�˖��X���	��/�!��e;RUb��R�N�쬟|& ��Z�# ��;�R���a[Y�l�ky���%A��5�W���*���sٹ��]��Fn,���]��C$V��o~��B����͊�yj@�0	㒬	<S�[�]v���.]Y�țxz�Jj^1:�|�b�uf�*�����5�Y�Q7�h��D�����$��@w��-K�U|U>;d1'&�SH�2�����Z(FXQ7����'8�L�l�+��FL
j���=���B�a�Z5����$1�������4.������.R�q@�q?��I�3s�~���#�|�����p