��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)�����z�-��8��;j�7�c��r�����^�cs��1m�)��9��`� ⛠��$�!�Ψ~��,�Cq�QΪ��0}��4��������,��hEi�����I
�&�'_�KBo�o'ť�
�������rn繵�K�\���W¶ო�i����ps�p+�sjD���R�H�W&v1&��s�FT������=|qYe΀�m�AՕm�I�aq�¶�՟u�ZT��q���ԧդ�W���.l2ñ��o����)���<���U@3ƻp��&P��14�$6VF������

T��;���y��O�خ�`]_̷�%���[�r�� ���};4�~�ѵX�M5� F}j���
��GJ�v�6�\��W}���q��#��q��V�N����P�G ~3-�wJ�!;r:hi[C�o7�\�d4P����+O����W�+�K>�׬H��>�%� kW��<���ۂ��?��MY��=��������ӟ�WT�}�䒸�VRQ��#�^�V�t��?����*����֟B��R�>���h[a�si�>�4V܌��LĚ�\�l�)��TvA�0� �se����$��'�\��g3q<��<�`9�B5R����^=�?~�������:8%um=��%����%d����0!tI�]*�&���v�eeWQi/�Ϩf{�-� [sNx����6U#$O$�;�[��O�_s% ���{K+v�ݞ���4�_����>n��6�$�4:UD�|�
����2K4��@\K��.�P{�#N ��hս�sN���YkZ]����{U�6=�UX+Na�@0�����1R�z����X�M��En�%C3�6K#N��!�Iy�A���D)���3�F�,7�v�V�*m*������
�rMK6VT/�d�N�جwm�u��7��M1���;U�9���{�������6�(
�*����}�[�وJs�S�`�/�U#�>���V�a[݋��^ܙKPRFpǢc��m�'+�. 7gt)חA�.k�g�ȡS��N�M݋�%�����u_�Q:$���U��(3ғ-�z|cI,��mO��z��j��r@��c�ϕ�lh��5�� ��d��������H~x��o��ބD"��Ǡ���P-��!�]�F�
�P�͕�I��~m3�=U6��� @�/��&p1��`qF�����i��V�lN�JP� �����d�$�a�f�l����:����
#���7�{���HV�QM����`�O]��xS��Wh�5�(��krKW���TK�@6HQeEz�OJ�طZQ:Y��~�(��vH��x�z��e:��7�뗾Y\Y����>'#ݪ��+��^}`MG̹�^�r5��������\��R<�H�Ca� l
w�i��`ao���,�_�\z��!���h���80;����W��[�x���r,��L^O4\ނO���Ј�k��Y���I�ETP���Z@��� �n9�������􈱯�8&prw�o�j���s�b��$��4��<�*
�b{Bn��\^��a���4��Z'�/��W��e��v�t�r�T�VEÇ�\�閍�J���i�p�������dK��+��&�b����������F�4ю�u��ꍉyp�?C�"��>�޻�D4S�R�L��4�{@K>�&��6�Uד؀�/��G�("p/ �����d��s1e��݊]b��qYX8{�-�fHH�,j#\p=����G!����%�^��u�Ч(����" 97��ЬM�p���K?f�m�&M�����ρ�Y�.�<�`LA[�2U�VT΢�j����#l�B�<�E��Nə���ޅs��h[��w'd��Xr�*X�9�����f� �8��:>J&���W�.]�vPNP��i ݨF�n����j��yq�[��L� 2{~:͎܁w���*ܙ	߈�!��!*VIY���_o�F֟����7�^����4ˎ]/_��E��=���ƫ����B�����;�� 3l]��'�T�o��S�i+�� ���hJ�E��	;R�a�����K�jԝ�����:�j�C��Iv05�����_F�5��#���`I{2����ׁ%��=ϖG�	�7s����5�
/Vs�N;�50P��o��xAnAWc� '��s�۾vVpu>x�)v'���U�5��)�H`ذ�[e��{��+��OǤ@�����������a:T�
ͱ۾E!�p�k�hv�,��n����~��0jߌ(����˙���?ˢ@oԑ�x�c̓ޡڱ*U�v4Ven�����WF�=fOc�7�}�7�	P)�P0׹Wc�;����P���q<��0S�Е�gUT�1;xydb6���=Wq��Ұ_�\+�d�C妕�)��M�i��ZM����`Bg����9���t���Z�m��K
ֺ�gc{
T,�C��a��Z��a�8��c4G��0cõA�D�/���f~;~_'P���RA��6��R�� �ڎ������#���>����T�5a�Q����,���1a�A��7QD��Ǎ��q��c�+�y��0�� .�}��y�@I�@öo,��s��P��(O�tw���X6��\��NMU�7TU��z�gbZ����%>�C��d�
���^A���{��b/˿�1��Ҩ�.옻/��X�$�^���������J�fH<��A� �3�2���w������w��,�s��,�u�Vi�����K��@��a����I^|����hZ#�1!?GCw�˿�YZWێ|F��_|-]�|7t.ʜWq�L�`e!yj,��P�t�>������sx:�'p�f�8x0a����uޯ������!B��m�N�0H��1�om����G�sh�<ZfH��Pp�BoH�. �-zYH���+�D�q��M
pݾ�x��yOy�>�<�Ӭ�T������xg���eE"j&�T�?5����1�}�p9�P,���P�`3Ym=,Z�j��B�
 �>am�B�([B�	Z����Wo9����;��%駊�N�HM��k��2&���)���'�j��4�����6��~�9P ���X�4���!�� ��bw�o�H>b�M�?#^�2H�z��]�%�� k.(����'l~��ε�7��&�0W-aB|�`X�.\5���
��܇�&+�������>���6�D����'h��28Z��Ѣ������W���(~�Y4źg�b�N�¦l�p܄�~T[�D��p��eopB���.*���Й5ݟ ���r/��l�2�+��'D�JZ�j
k�i�7ǵ��^7������HSle'�ʊE����:���HD��h� L�~���×�>��D=��wi�9�h3���~y�KQ�<ŝ#1�o�!8�2nE�_l������>��p��v2�qv��/�H�s�[�η��[���{R"6�su7��) ��9^ܐH^�Zs/���c�:|�ڲg9~��EDckj~����n0������IϥU�i��~�ןf���z"�����BV*d�\N��{�F��&8���nXР�\����"����"�0��A>������S�=�����H\��"߄��-�^f�l�m5L�5�o����eQ4�\ə�ڔ�݌��W�/��Xn�z�=�,^6�ȗ�= �u�9�N�?Ck
�̴��@��aqt?Gk�J�F>��0��}���Hq�՜�\��L��BE�%`�f���)+9�������"��N�������WR̎K�������5�:��������~��%�<��e�?�P΃����(KO���'X�Qp>�p&��9�����C��jq"kP�(^hQƽFn���B�p ��Y# L�W����w�Ŋr @m��y����.UZuI�
n�r0�~ߊa��"f��3gO$��$���:���>sNyv+�:���'V���d&�Xȴw�4(˪��:��TG}��+�7�8l�e3>�,.�`ZD�X�����vkr¤�mcz��Qv-e9X��%8�sX�|��$�o�(�FJ�������1���}�z��0������5F�l!`�?��p$���$��q+k��,=��[�qJx�3);�I���7$���T�~yei�mIi[ʇ'�*�Fi�A����C�j5MLqa8z�V�����{���I?���ƣH�7x�A≵2V�\���W�з����ǘ�c�����v����H0P	vE�+� �0����Ш�AK�w:<��T��{)�Bpi���5��]����q�Bfk��05�)��wP<�ފ��"�n/�i���<��� ���)mee7�4J�D8N�a|�ө�W>���ێE��6}p����x������u���&4�� ���	�P��Hct�Du �'Ce�?d�}A�W���6�)æf�:h萟<�G�viZ�Ξ׺2��������u9�RwR����Rq�V�_@���
�Z���QX�<ǲWK2��xҊ�6��vfQ�ƭ�-�s=�/A�$���?zn�m�Y*x@��A�����RA�wQ~��t�}Ih��O�j��^�u��"��F��I$%�����m5��Q��Y���)M���8��v'��S�o�a���́��=���F�~u"G���ٌ���1N��/���оA�.�(\��"�x�P�m�5F�d�m/� a郆�r��7K�%�D��eɣZxl�QK��K��˦2pe���q�o�Bp1�A*tl����a���0������m�gF(�!�%h���j�@˒��k�����M�Z���ſ8����m�"|�z�g�-�����J�P�"��/�|��mk�b�n��i9uqC_�E:�]�~�-s�p�`^_F��B�1����P5�v6z���&;ï�����	L)aw꼐�I%J�t����K H~�U�g $=�
NS�A����'�ak ���5P
��OZR@�T��:�m`D�BT��y�B^Y-����w�ij֌���};9̧N��$׬�X�ƒ�8_��Y����sVE^��8���;�����-uԁ&^�V���e4�F�3-����Ѕd�6�0��"��-�kt���=��V�����������d�I�:[4���-�t�b�{[4��;�_ji�zS1z<���]�
��XX=������@3}��ĻP���y��%Vو��{B��������o��(; ��ն�<������,�"ŷ�7����1FQ�L��{�	Y�` վ�є��LJgM�<��$���Ӵ#�!ɡ�N�|,�'��l�	9�w��De��i���D�3[��]���֣���X����(�݈I�B�����.��EVQtW�,檷������ m��1y���v�苝7H��=�~.O�y�vh�����,�'�V���lu�j1ی��}i�hP�g�9��o5]�\]9���s�������)W���7��ԗ�*�;�Z��'M=��8��j�fV��*P������b�@F[�A�&7L����A	�#O?+� M�[UK����i��F\�\U��w^�
�� �d��#(R����iչ�B�<T��[3��著vF}g��g�U1���V)����<9v�I�-i�����a=�W�
а����!�"���#ZN�aُ�#��Đ�1n�9\���G�_2 ��o�Fǹ�])P�e>�������T��m$  ��E�g�3�K�Bϐ��7v�5�v�1��r��R����Jү�a`�Z���Ā(&)<j�x����KU伎S@HoO���ק�(ܒ9�G�~�Մr�I�SJ���}R4&�à���
�:�pЍ�Y��/ԕh����d���v)V��Y�+�d�^��?��������2��Ls^�����pz#��p��.i�=�sQL��u�_�Y"~��S��
k	T��|q,�K����n#�smV���X��v������8W7$�9�#x;�+���r�ǀ$�=r�b	��=���H��:d1��y����߱�l���d�h�_��N&]d�\]�#����w��q��K��E�3��y@��H�ǔ��5����.k�a��"ʃ��ڪ�3�0V��iљUsF���Y!M���D�2��K��2��(�T�S��_�Qe��X�Qo�����dm���j(���2��d�g}���L6B%=A/�>�����X~�1ڼya@���^��J��O��-g5ɦ�dy�p&�ja��h+��OvW9!f:
EB�ׄ�X���M�O�E+6�$}�޷*�O ������|<A(������uC�q�RL�G}���$F�� w���@�zӚVGQ�Q鋹�K��,�b �@jЭ2n�A�oSh#�K��Z��Կ���n�^a��^V�65Fg)�9�8A�;�����uIC2s�3ש��s{����U�������^1d�s]�)��׹�C���ߞ�R�U�|���:���֕F�`"����9��Ø�ۇ�D�}�M�����]?��	�2B�^�N�n!羥Bo�	[	,�j�]��������X��^J�ɳ�LT��d�KH���V2�����5N��A;����tZ%�R^,��%X���C^��g���@�M�*o@�����hH����"����o�X@���x�Nx��2��ɽ����>�A�����,��*��f��D?��[,�	J��?h#��cT����ř*3�9[e[�:��/��
�RH\HVt�Ŏ���Yތ�p���i�}�A�
7��}#��GE'b��Z �4���$c�ߨ����>8t�l���-趝�lVJ?�fw�"�F��lH8� i�>&(�u��p���F�x��h8�ϼTQuۻ�Q��*ޖ\�%������'�X�)��b�2��x�l=�H ���Zf}����Pih���O���5���r�v6S�5E�T��'׬��<��׍�5O�o@��̟
���x4Wp���{P�Rj�lQ��A��Q�v��BAߦ`sgx�Y�)��zR�J�,=�����%J�%��p�d�Y�FdA$����`�P��;�c�
X8�=ɻ��0~$k�����T2/���W&�| �{3U g�t��ɉ�J��fj�
"��%��8
ԬQ�]��d���c��?>��PH8�(�̓K��_�(�E�"ռ8�<�0�.��7��X�]5��1ƾ�˔[��h��3J����L~�tz��໐SHL8ò8PO_�6'�fIj���s��q)�-��u�+P�b�O��G`9:d1A
@�cK�)�����s<n�a+͑�C��� U��Y�C{��`{��*f�v�gE(���3��s��R���3eY/�%N�����)�%���i�f!��q� h,:A�I�w��M(�;����^�ٴ\�$�ۀT�4?PA�
I富-��& ����&ʳ� XU�$���d��w�A
���zϚ�[��õ����_����DX(��d��ݱ��2�Hܢ�S��mH-)��?v��H؅��5�=��"MG�&u�����O��l�t&f�2З ���"Ne��弸[<k��{�=�!q��'΄�g�@~K��J[��n�F����?Ѫ8�'���������0A�9/a])�:�ӯ$Z��M���ߵj?��V投7��7����n�VB'�n��˟"��˙�=�P���E8�HH�N��E]���k�=�莬G'�OĐ=g��yT}M�H�`��pyӤ�m�A:�P�͓">I�?��0[�]ɜr�}�{L�®��V�h�?#Jx�%>� #D���}Y��e7�L��.&l�J�7�㪼����!r�{ۈߛ��7�ӠT���eG�1a������6��)��G
&�c�Z�Kޅ�8�|�	ҙ�?��H)��8��c�`4����Ɋ5������iF���+<}A�]�}���1ln�ye)���������O�
X�f1v�k[�㙈*���N���.��-^��lӣ�{�T@�1��b���MӉܤ��:"�`�G�Mh��	�d=�'��˺h U��	>�K�P�M����7T\&$�����P��f��)=|���掬���1s����bU �||C�y�`@����.�{z$�vl�_1��@K̴�ʞ�^�X�
�q�������D�=���٤j�9D����lH'���G�����z��lPV����j]�����"�N��l�i>��lA90�����w|�ܨ�k�7ĬB\q�ӭ߈���(�V��r���$d��lt�G�pVI�~OC��[�i9E��q��a�Q�A�1�Kq���:��GԦOBZ��'e�.P�a<�G[GWP�D����N���݁���n�IA¼��R8�vڇBG{njj����>[�O�zu�xVDL8�g�"�Qo�A��Ƥ�����xm��ȅM��Ϩ��{ry9A�b3�!��8�2�Y�5�">,�4�4%]�?Y�s����x+?��IIVs���2� ���x���be�Q2�rr�wwa�	�i�o˸_SX�3 �\Gh����U�u��X��w�ŕ�L��nFG�<��6�|�6�1�
����n2��� ${��3���씹�aZ���2�+߼��	��8��"�\-<J��#?5Z}���v�x�����0Zb�3��������}� =mY�9R��*T#���]4��8g��O�
}����|S����Z+��؄��C��a��w���v�G�/`In^7�Axi��T����4o/$Vf��������d>(|�������$x�������cx���Y��:�'����-&�fUyC��ЬM`��ƅ�㭟WD�����?�Aa��l�}���B��~����B8��bF�ڍX���^jb�\,!��OX�2�\�H�^X����$�Yĩb���t��'���ї֔\�~�v��2�8]n��pe���֞��'e��`�0�a~3��{�Q���Zy�rו����C�U��[�*�w<��T>��{�)�o�Ya���3���;��f�Z�~�1̧�})��<���-�1��$�!�s1_�ONff�J1���3Y�QNzeP���鞕�z�3�E���r��1�~U�����%2j�R��G��
��譊ϩ\�֏K��=��+^xN1N��S={1Y<i�6�<JD7\H,x�v	��ne��К�ds�/Y"�s�p�(�����,�Q�����$t���F2l|FU7M��%&+��ob�~k��b���\"Oj�A�;��v��n�~p=V�2X&C���At<95�UV�3ʏ^tS�/
Q����{�iN��GUEZF2�5����(J�O��������}&�*eǽT�Ggu�V��Q��K����/6KǍ��Jw9y���7�f��s�<$�Ј/���HL&}��/αZ��_ �r�w`Q�j��d�=�t�i�u1��P �v�:�%�n�U���j9U��Q����,:�Y(� ��2.cO�-�ј�bU�+���@�ۋ�ş�����ǒJ<��L�Ȗ�:XU��.��Kw�� }8�ь=����-������L���V���U�':i��xI����!�+B�������&�qi3��x��*@�5����6�k�`RF��r���L������Ģ�����a�<'�M���ݢ��.�ϓW�R�0�\�2�^4-2C��F52�[>��fdM�\�>K.���7��"(�ڐC��o-X1���.;�"�U�������8T�D�e����w�Y8��7zk���=�g5r3� ,�lt@:��v�����F�SL�)t=�.uDBn-�Vb9I�:{b�=MHý����q9�o���n��Q��I�e�H;,�6o�;���	y��m�k<�������!�f�8ѓ�����M�~�)B�AĞ�ae� �,���s�4Z:>�(}�K��m��=Gp���D�p�w�]��0h�(��6����)�j��ͦT�.3B��n���jĆ_N�V���ʫ����a�N��?枋@H�'������T�?�tZ; ����팞���)�ji/�gcR׬J�[R��S��|&w�����b���u�h���3D�,0-#�z��+~хh��K��46���ϝچ�̆��&ZN��M���#��V@}:"�]}��z�4�_��8�����%�R%>��l�/O���p%�(!<3_���v�D����k�h'/���Vن��_��㔾.��PA��E+�;�p.���v���0�Jj��ק�Ȭ.FT�]Xٲj����'q�-@!��m�����[`-g\���4�H����r���gc��τ�6y�x�x7Uа����Fx9�+�����W[gR�Œ�����{,ر�;3h:���JAP��O�-
i�]q�M��/3���(ש��<�e�����i�����avB�9�!�8%.��O���]+�"܆���d��53�I��� )oUf�g%��G����ā@�=Z:$��J���tB��']��J��/�3�Y|�f$�9o[��v��y�>9�G�셿+�Vۏ���3�MIv�n�X�f��@����!$F�_�Tx�5+]э[u�ם_uc�>�r��%!�3�,�7X�N4���ڤ
��������n��ٴX�׏�wu�CO�ꝡ��L�KI�,�a��U���Z��5������<�d�������w����T��p�	��}�#�(g��	��~+�� ���g���&�	n��"�%s�Ů�a�N-(�u5�do�����1�r<�5�g��[_��@�t���$�a�������V|�¹�?�E���}\C����</�V�C8����0����+X�����cq$���� F�&�3��4��w�خ����v�[i�8�e�Xq"��O��j9BDPo��DoV-,�|��P������)��n�Mj���^m��Os��yYl\]�B�k�%�����.Eh�,C�4�W��[����)J{�:RiR��V�Ai/�;�A6�$4�=�޵�WIl��0N�x�	�6Ԝ�DE��^wc�|�v)����㲋����]��t@�^�a�^[::6<ji<I�z�]t�� y�O���!@�\����%�ahrH��)����'�w�,��?>B��/<ɸpiTۄa1�Pؚ���d�[���Q�Z�]m���r'6�jy�G�f=���iW��#���k��fn6ˆ&Im]�ov���</�n�O�%��Uu�#`���w!�Aު6��u���|{�uh��M�1��㠇J�� ��2K�\���	�d7(��7���s�/�Ofv���������e�-�p�ZL+l�����=�nzγxć�,�=�`���x��f�W���'$5Z����C��
Y��@6S5�A�I*-����L+:��F!���:���=�?I��J�n�	��u�	�eJ��a��Z*f�������E�H;�.&�ѣ! �1�pkm	:�82��Q�p�}�A�&Bb3}!�38��pI�3 ?�m	)U���]�����/+�j�{��j��� !��=tB�E�!���m��+5zeG �HM6����9� Z�+#A��Wv�I�9�}�hR^4�+��3�i%��)	������#����Oo�uT�4lF�l�_+*djI@� �m~�PD<�S�����8����;pB\�TKn`oe�&!gv��� kx���bS���6���� ȍ��5=�W����Щ{����ܕ������޶Ư�+L8��@���TZ��N�%���(�ɩiI~j�ܳ҇�|ᛞ��c��ʠ�V!�?����?�ӯ>Xz8<�A��^���$VT�,���y`��7ݗRb���0S���yG.�EH��J�؍W��o�"��MޔGoJ��$����hQH�j*Ǡ��ɰo��?�h*���C�?g���w�'�O,3�5��b<�/����"���+ A�i7��
"�/`%�߾��i}��Z7 0|��1'��j�,G�R��2X!dc��~*Z3��ժQ�6�ņ;֫%��V��ϳ*���!��u�|n� �r	�=��
��X�#���v5Du"I�;��)A.�_��Tۖ��jA�a���͂�j;�֙�o���Lʔ�Hg�fU9���D�b���4EB���G&����~*/$�S���B�1��YsA���[M#7�&B����>��; Ԟ���k��3�Wэ��W�8����M�C��`���n�d%u����+�ȫ1'��-@�CJ�~�8�l]�F}"�{4W�G�!��<�$lxZ�0�'4�>�a:;��H�5��L	��}U��Z��T�x_��qv_������}��� �4�t�/#����i���0^�/ddtR��u����=��%'�r'�"�>	����9�w8n�h��!�(d6��;o�o�àµy�A:��:V�?$��ߤRs:�� �ӪA�R��T͸��/��
h�r�� '[s~���Y��\���94��R�gŬ$�B����_LCp��F����>b�،�6��߿���I*J;|����<��n�|"w��8k�����T9%5Ph,P�g�o�OvQ�)�3��af�K��9���[��.Z��Ɔ���*�d'�m���G8NRU?�Z�m	�����Ϋ�
F�F��@D���ށy�J��t�(-/�Z!O��)��&
�JW���uS
�S�*?ڍ�;Ӓwa��G�Jሎq��-�W�=����`m��������kU���PѮ���� ��q��юܹ���Ƹl-�֙�<��!=d�.���F��'n�<ḯ��{H�*�����8����L�19|�Fs��[�+�I�Y��� ���o1�j��/
��ʴd����p����x$���ڐ�0y�|	<��H������b�Z$��±4����Pg�y 2'���1!��e8k-H�3Gn�}��L�FzR��`�W�? ����0|)��9n���pY���C�P[���È�@k9�{x��2
�=��C�̃xUȗ7��v�f�?���ש�l��}ͅ�*���B|K+g�m*�nM����C��l�&������i&�ju���
Rz�8H�J�8����|� 9��yuǗ�@V�bPuR(�	-z���y3D}���j�&Q�"/-Pa�a��8�bp�gwW�H�a��i*rr|���B����J���΃z����s�%���.w����u�y\�q��.�!xz�HΞ��/ŕt��u�k��l�Gə��*�1ݷ�bZ6܏�@Ņ[>�I��Oާy�d��$Ҋ�zY��i����G�
�rz���B�N�_l��3da�|�?8�ĳ1Ѐ�i����P�U��/<�ʣM =�[���W*�,��PN��΂��ڠ�(s7a����[i�����3�V�n3m�Ah�,��
GK�~7�u���Ѕ�e?pVu g�Ba��,q��A�L�b��u��q��С,e.�� ����n�=��O#k]����������ـ\�r���"1�i��a�OY�%W�*c�-��z �!�b�����\C]5�nTb�Kj�)��<�DAG9lB�c�0�>.��ͤT'[z�0a� 5*U~Kx�W5%�'(�"��VAȏB�x�F��=p1�p�uv�`B�.����������@��˅��'�P͝�m����g^�*�ؼ-D�l�E��RT�A�F`�i�rvY.��Zv��,�A�]wq��+4��㞬�� ���|���¦�����0O�������Zq�R�a�|� u�3�N�yK�VS��u��Yy�`��F�}!m	}FaK��j�G��Ƥ����q'R��0,2@2���x��v:|�cKa�`L�5�Ol�T{�ᢧe���#I�=O��{1ҷ�I�[9�[��
i	�?k�u�0�s�8��"��z�8ۼwg}x�،|2���Ff����^��w����~P�І�6t&��K	ʷq|��N=��0e|�Q�
�������:a��ĠZ��6��Gh(�|?X��1�|b�f^����p��7�V� �M(�Wo��<��������B����i���
Ie�k��!������ך��n�8�ݼ|�P�6�td?[j����"�\���.P�|��(�kK�Za������(�,�@��Ҏ�5a�H�K������@�Â��7����{�w�t�͸,܍�S�&I�	A�6t0�]���C��z�Cp���oR���9#8���i���05j�-�"��L�����#+��)�!4��O}��/l�L�^s�G?L-|e>	�y��Z�]48���pa�#�t�P�1�T��'���Zf����H��n�c6��Ж���,�+�Ԫ鑰;:f��7}��<�-�����3m��07��W�ɬ�����@��������A�^,G�a.���	�?�\�=b�,aI�h�s�ɯ"�|=.������|���0h���I�(�ڄ5���?���J�a��b~h���z^���D�&���̦��G>] � KՇ��nǀ�fc����dC;ot�)ꈚ��#7���Sf���qD�Ö�}�}�(#�U3�S�d�v�;F�|�4>����;=ǿ��>a-�j)2n`���ȔS�9���
�_> l� j tc��[$� �V~���'��`z�)G^�:ه�Iʷ��9�<�Z�u��E��M��T��e	�|<g��*�I��g� � ��o����x��h��fH��-0[a�'�K	�g��N&j�Ѩ�Ӱ�GP��<�����+��X��>��SR��.G���k�]�{P��B�!h57�wq�ˤr0x�	�%���}*���>�Ӝ�j�^�O߈��$��;|��|�X�Br��<�ǀ��	����	�ڊгN-���p�6���x;��3��Գ�4���:T=0�I�=`�#�
�7N���#�n� ���A��"I#S!��͵��^�0 �"?��em���E�Q�{:�y�j��(.@u�Z����v�k���靊�q���p�u��(������ū�tr'��Ju�b��[��}�_�ܼ�Cgx_U��4H��vo���}�J&��χ~5f�	+�;YӍ>|����?f	�T?�Ӿ��#��n��o���,0T*�!��h�E�S�$jBg�V��WIs�{8
aj��r�����Qk�����e��_�=j��b��,:Pd;c;ͫ]Z�����fA^��-���n%�A�H��J5/�or^Ea��=��ӥX�jrm��Uk�IQ�"�X��nFe�L]����2,�n�Cv��^�#x�}���/U ���˂�4?���o���|��h+zX{�QA�#W���к�ѝ��L!�������f�����H}j�a���x��}P���=p�~-�3����7�>GP��݀s�E.�Y������6,9<SOř� ���ZO��z�0�un#�+�$����ck���Hf':u춛��>,x:�-��V��>����C�����F\k5� ~�����RM������8�6���@�	h��>��+2�����s���E�4�}Z���7��}I���|r�}����޲ĕ��ƀm!�D�5��(q���>B��:�ȱ�}�H��e���P���dgU�rq]�����A�{�.T���}?�^��O�/r�r�stƉ�"�i\|_�}�W<�;��XC%��M�+
Q����oD��t��}����H5Pǘ�U��9[���z[�"���.pJ�`�p����45�w���DEw~�������k�UZ��NlG��   �.���u��ߝ��__צN��fz�@��)�2y�0�Cy��^�Y�f�1_�H�UU�:=��(=R�kP��슏��?�8o�?�e���v�ЁK
�jJ���q^�(<�u^�3@����]l�$����<�@�������,_sS�YX��!W}2?��r^��/�z�e�J��k9a�[�z������z��y:�VG�I6�-񩇁Ü��������S��g�y��`�У���m~e������1�E����yp2�w������'�cԽ�3����oi-}��P�.x���B~����_N������6�ȕ�Kv����q�r��h�;롁�V��X��IxS�����oZP��Q�t�-�!IW�1����w��;��~ T�����#�l3�Cx��RU�kɭ�
z ���o��I������H-��K�q��u\���<�o�J �ھ���	m9�?L���)Ћ@p/�d�xݨ�����Ӆ�6���{/�D��Y��c��ԍVr�c�r���(= ��F�4z�e`A�ɹ�H������Hj��y��xX,�}+6�7��W���G�/4��b�r�?ܹ�{L/�qHC��"���|��+��?N)�R_� �qf����R�Jed琜�h�?i���lԎ֊���#�m�-��]����;�S��F��M��]~5�M�1c*��0�6��\[ n �BB�3���/Ӵ�Lw�j{1��uF��X���cr��ʖ�߇	k���	_)1���֣��[���rE��<��/�d�0{π�q�X��">�����E�7V
�ʒ�WtT:E��6;Y0B�Y������͛M��~���8$^ϒv�.�bFB��nS%p�9M�D�����wg��a�%z��Q1"x�Jd��NeId�k���2;C�/g��]��IzS�;H��w�C;���~��d�tݛL� Y�옠 
��*՚��>IM(�xV��.��i6��*=P���IF3��i��l.���j��Y|��PSh{��;��G����U^Ь�K��쎕���f��?�'�z&��L6�2o�[�0�	3I=Ґe�n~�א����٤+�r�"]��..$�!����j�1�Gt��%�MH9��/	��X��,��+#��7_�*A��$�U��u1�|>i�kRw�$A�oҪ4�5������L�+�r�BJ�+� W�H�ׅ���$Y�����C3�� T ��q��-�k�E��4���*4�]��?w��雦6��ǝ�/���uu���G�Zg��J�D4}����B�����N��*l�q����pBA��UH�1�� gfL����5[c���4�^#vo7�����l�qЫ������aF���M�ƺYD�0Qݲ�J6��@,���*��FR[oth�ȗFa������8|҆DC1��|��}�$�ՠs:����*����'���p�Tx�G��"�4p�T����8�Y�r�_q[L�.y�i�PH�&�&i�����Ϋ}�Z�����Ɉ~�$'�uf��v�k��Âл��>ƿ� T�M#�RT��S�ClK�Δ�a�	��N�m7��@�{�.�H`a����[�<��)y�]Z��9��dҡ�����('2:,)E�9GQ���ɾ����U�$dN�=������Bb0�0���kw�Nt��~J��y	B��2��gw�Ąԯ�5��3g�%k��W��/�~�S[�������#�ò��^�_`]��$�!��Q+���#�<����`qD�/����9��b��%O�J��i(��!�(��D�'��'�%aW�̲
�Uh.�f�*�摖=At���<����^�Au���9��a]wG%ׯ��;�nR��9�.�2F[�yC�׮K�h��6bs��U/����\�(��jHR>	�t���4Ե��3�2�)�>�"�t}����\kb��]' Z>s�@��A����}���as�K	Eg2�7��b<���|^_n�Oy�nj�0�e���P�5J	SO�f�������/	4�go^
GB�(
�?CN��X8���XKC�KX��oU��^��5���Ɩ�8�{��oِIBoj��s;Y�2>ɑ��rDLC,tzE��g'WO����]؎�}+���yLb<����/�=��m�@r.�M�����aNuG��p�i�4Ui�^FW�4��%՟��aL!��#�}$J��>��ʶu:�+��tumtQ�A�y�t��]�'j�0�il=����7��sH���y�V�
�LS�P�i\p�����^�k���!��Z'O$�����pz���GSScnW[�}�x�o�*���jf���.�~��s����{�� x�Q��A/�i{w3<I�"am��D���y� ]�2�KU0TE[�j�����!N�e%d��D<���ᐥ��N��s͔�3Ҳ�L�4"?6.l*<��)��x���D��f�
.���"%�k�
sp�� y�ꦆ���X% ��n�������+�q9�)��f�����,�
�� �A�^\I�aގ���]��wu,IN��m]�=q?��-/�&U���/��61��M��icz�O�7��RΝ�5'Q7,Z�Y���'�h�;�$e{w�M�ҹK
e����T����P��O�Ua�V1hq�����n<���\E}2�Ͽ7'����O^� �S�&�%����Jgi���&��_1�3=�$]+
�O�?���ſCw�rV2�ߗ�{�1	����dOi� �.�"3�LU��tM�����X4t��t��z�5�����^�;)U�o>d��B�B��C���Z|�
fT���~��^�
���GD�u�~�ӑ^֛̊�@��i��Ts;�e��{>�~t��F����ȯ_��Qߥ�&Cݣ[�2��Z��X�0�!�:J��J�
>0 �/�a�Ϫ�j�f���ѣP��b*K9x�����K��>5�_K��P�ێ�&8��?�d�}?�X�/�.�PuR��4@����M�2K\��8�A
���X1v��D.�
�㋰�M��9��*�(#誵9�ɯ��Bέ�����"R���#������<�J�����"�	�M,�-�cj(��4����rT�^@%�:�����+C�|!L|W�$�����%yơ�`Đ9f>G�"�Kj&y`az�E��{ ��ַ��?����#�E�6����ç�g(��S�	��L���3��G�A���\~���[�6����*1Le�z�sGD)����͘�܊`pM$����JcD�L��v#���m�r|�}���!�2���å&���7���?65[h�'kP������c/|��le��C?���C��jwU��t����`�X#>�S1�-���l+F��
�~+ tHu��d�W^è���׌��&`C�����Ax�B����[%X���*3���u��Mz�Ġ´
J��%�c�o �.��]?w*;�yJT)w� �X/7�"lfHL�=��vȔ}E�h�G�uܫX�<�gPG[7K�����ŨCԠe$�\�_� xCrRt���u\��g���� �;J��k�p�+g�|�>Ǹ@
|!�g���ڤ��jX���al2K��l��g�5l/��d���d�#R��̗~�/RE��;��x��wo&}*���,�D�R;i�GI5�e�v��
���Q�����"�`��1�@�9U/I�U��1sߘƱx1���Q�t���@�nG�9 o]"duq G�N22�p/�.�4��;W�?�����J%y�̃O�Z��ṛ�K�M�B���V���8@��ʬ��]�>^~�-b�:�J�g��H�P���U��<�����E�0�0z�԰�6��+$���^^}�?b�:Q�8Be?�O0j)*W;;�!�la�о�D֧�'y]�6�a�ߖ8��xRA&�dq�[e;	���-�?�Nm,=���IP&,*6(!tG�a-��q׈�D�Yӯ8��"gQe�9j�»i/{�ǘy��,��;��F5��|":��$�;�������4Yg��������V�,= Q�m�w���!3�j5#�Q�%(�M�<�0�]�6<��,����W¸�|��9S�O��>���l�!Fj��jI�܀�o����!$���u#{�S[0A�TJ|N�;1��N��|]�1�����u��%�.���A�uƔu�s�]�ߥ/�"�s������2��|����xq6���n���ab2��=�
�ݽ�Ez%���H.�ҢA��bϝN�岵��>*N�B>�5{��CiF��!�P�yR��Ȁ
���E�\53��u
����F@�	YH)������q�c=?��i�cOV�H�go�<����MgJ;pR{�j_�e�����@l��'��j%U���>m�f��峖1,*:GT���wN6`!ޞc�T$�����yڅ��G`E�&�UsЦ��M��ͣ"��e�ĸUxi�%A��}?��9�lPe;ف�ǳ��4��y���fń������X�ܟK�5A��d/�.����a7��myb=�t%�"u�ai���Nx]��`�o�ٷ~�כϥIn��7�1e|�N�KE��gKDg�|��rY��@��c���
pzx�ú����S�6������񨒺��y�������j��*�wٳ�@�	��U3s:�6�ȪN�'Q�L�-JeF�����`���:��]q�uז?3���s�}//Rݚ�)]������(]�e��m��
��(�y�r^���]��ؗ�ծf�1C5���cr�4�BwX ��ARM�\�:�{��b�L�'�m�@��5��Ѯ/�;��us�z�ݔ�d�'�`�䷲��3��}��ֻ:Ir#e�,�o��6����\��d,]���3d\��A&��� 3U�būe��^:��ا���]B�0���î�IF����x�0n��Gڼ��bC9E,XO�����y�M{{��7��m������m�%:������O~p߰�ש�uKR~.E�\[�J;� ���Jy�5aE0��9�
�:�j.������r4�cP.��O�w�x%X�c�0�ԝ�(���o�
�T:D�˩&�~8������g�[L�a�vO�U��MQ�AaBi)�s<��|�F�OK�sR|�F��s�ގ�Ҏ�-NYjά˚�gP����O�nM]r��gi�>s�Ɍ��q]�EvO25.L0����&.�}��~g�����lt�ѹ��0�c�?Їy� c���ӆ��a��T_NxX ��*K3vF���5TG<:obl����~�*��p����(Y#�va�+1�pW���L���
���qD��d�!�r�Wüv>�L�.c���8�0s�7S�y"�Lm��fr1l2|�p�����-:��576n�.�v��� �T@`�W�Np�i)��4�nC0<R��y�������O���ł~djyq���+��[�i��^9�չ�坣��S�@J,ꟓ���yNy�M_�`ܸDJ����м�������4��Ք��9�����%7Z?����}���1y�Asٺ��Wh��q�1i4 S��]�8C�Y�NZ�-MGƛD��Aj�27[���
C�I��P>�{�ۣv�q
�߃HIdH�H�ujO։��s�Y3�bU�S����{B��M�h=�'�`���B0"��k�(zx ��������b�Vֶ4U�9ܟ��M���'�SmǪ|���y�6�a7�gK�_Gc����p6'4��F��#��u���Ti�6����j��75���@�Э����_�T:R�_8+G@�R4W�g��m�"�V	Nz������w����"�դ\dK�P8�|e )�Z���hD�,���Q��&�a��C����_<�dq���cCi�>\MOւC/�<�<�TW���P{tEѿ�н"9p��w�ߗ*��U� n�Ki���1�RV��r�V��檧����_3��z���=�g�J��iX���s�~/�l/�T?�NN���&W�%^�Z���X�}˵����uo;-�m�׫}����(D�҉����РB�
׮��G3�Z,f�km�dv�)�-���kR����K[R�<�@v���.c�m%��J�ҕ�6�7�r6-��F�^�0���ӷB��q-s+�i�s���>�#�,q��N{W�d/�c/��V$��Z�L_#�M]�����w�
��P�:��d����Y��#6R��_���M�'�:���5D!a3�^�q�{��p.=P��ū3Z�&�޷��)#cȋ�>� �׫�<<�:�7;z%Mc�zLF�H�R
_�)�Ҏ����f�;���x��ӄ�9�Kw��#7�-�V�����y}r��	}����r��%o�
c�O����,méFD�
F}���F���X$�3�s�\fnz$^�W���2)j㖒��\|���e����Bh��B0�Nؠ^�}�Y�����I��P_K~Pd���IfM `��~.�2?�5cYQe�Ol���T�f�QG� 2�)~S�Ј�����f�gjҾ�#爅y�O
ѧA��1�0ȫ;L|�T�Y>��⋮[�����T�3�*O��/Ba/��wS����H����?��(A�w7����>ӡ���|�p7^N� ��Kl}�l��jl�\fҊY���T�[��G"��1u��e�����z�����mI�����0�%}��  �ER�Ȗ4�E,W2u����&{c�m��ADa��Gh:�u҃�n����u� 0J��)���sv��욕�����Ĵ^��,��$k��#�[�v=��n+�\��,�e�R���yt0*M��dե�E�׉nug��
��P����L�,L��W��9c�1K$Ƹ��@PIn�R�4���=!�4��*@�1�r��)h@ˬR��	9����N�Y+�xJ���O�DJ��B�|v3Bv�6#b�����%�S�+j�]6��ټK�$���;�_�|Gè3��+:�q���a��-e�qPz��ѐ��Le�$V�<�V�qt��T$�Y����OS?E�%�#N�.��e�t�h뻒�N��P!���(�V�c� YXd�V��e�@����:HY�a�����H������������pV�H���� ��Z�Κm��h5[�/�P���G����P{��3-/b;;k�VE�p���C��H ��S���pr�:z�z�|�S���$���ذ3��D�'	��ԩl~�s\2��#;%����3u�	�������;���U@��[�ǯs��n�\�sM@C��/�3U�72xwsI�'�Qԉ�⣂Kd��vhuޜ^6y���ܰ�bl�qf�2Emݘu�[�z�z�+FK$�͹�u>�QdZa��(L������w���]���������rҍ��O�|#�cE �3�t���ͭ6a�7L����ջ��$P�)@`�5	*��bN�I�(�N%�s��rVm���&�E1��D�����9�b���['J�5)*>�%P�Z�?�a���ǭ���O�t���W�6d] cP\��NJ�T�
MK��iz�:s3T�4Ȅ�/����6�����ұRc��~=��*|��Nҭ���_�uBT��k�:t?�ifgYp��<��=<\�L��?<���e܆u+��S���>�������a���"��Hv�\R���!�[�-#��`���
��U��s R�R
���S1����T�(�]>��H����̲���{g�3��ڴB �Y)�h�{���� ij�*�y�<�6�P�B� ʺ8�˄Pϟ��]�H����8
�Ȣ�����v_UJ�3F��\�i�xy���B'��}.�3�"��b���"�7𵿎�v�MTi��P��	��-щ�ZL|E�/َQP�~�$!�=R7T�>�8�[;�[��<���A�j9ş�	FeG�	�yDO�S�$�bY�M�O!���GF �(��O!6F���o��z�g��?v�XH�ž��[���F8�M��o�rU�dQ�����
��z�y�~88PR��ʶ
k\�&</�ΰO݊�@���KY��J|<4#�{�m���j��O)��5�˦~x��L�ҁ�����A7,��+��Sy�=����9�g��z����b�l�:hs��F)B�B���u�٭w��~����0�P#"h.�