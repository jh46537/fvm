��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�I�X��a22}L����*����
�	#�A�<�^�Z-�gB�(q@k����>���g��Z�ݖ�Zy����r�4AU>$�N	��-�u�u�'N��
c����(ቻ)O��9Dk����K�9$s*{����o��������2ؾ�E�c�r�Wd#E�K�#R�۪��h�?Ľ1h� �wy�9��A�^w�(X-�h~kj� �^T~.mj��%	�
H?�qh-[`_� ���L��e��!�������ڱ�����3{��:�<���2�6�_ 
MfA�70/;�p�P��RT�[�@K�a����T��Ҟ�<�<����Sb����$7�B���i�颼��XQHɯ���T���h�b
#d0Hb���쾖���(���"C���w��W���L11���� �:dY��O���޴z�Jc;�D��r	��4�����4{���I�����fk�T�0j�G��	��g�zW��e��9���$У�)�Hg�n��$wG� ��6���>�`;������28��i����|�U�D���͏A|��8���#F�6�� ���oHz�����w���0�40o�S[��xȠ�ZKʍ��@����,�Y5B�̄����:��Eg���[�$s�����1U;�X�On�Yk��#,�`OW��O�ܹq]��Ax�':����fu����&���Ǥ�c��+z	A\��u�����R7c*��B	�<V�S ޱ������f�2o��]���^>.!��$Ul-�`Vq�Y�jE�u�ĩꤓX�}S㤋\��R� ��l�?!�^������M�ۨ6ʊhN�bg��큮D�j��he�½�5(^�������w_�֫���\w��N��U��n�Q�T�2>��+9��oH�fJo%���3��L��e��j5:�[e*����0ϗ�pMo���&*ݯ�J[���N���̏�U�� ���+��֋a(����� ��m��l��K�}�^u?T�-ڷ5�"F�f���i\�8#���;_"$�1jJq�t��阦pİ���ŮHmM5���q�ѱ��`"X���M��&&Cs������Ѩxe\xW�Y�+�e@�N�2���r�:,�,�{���g��/��?Ҋ�lO��?�hԃ-b�w0r��>��~sԭ�1��~�dU:����J��'=�sy�)�Z��l_}��9��㾪e�tZ��6���&>ͤe�E䠱/�'�����6�&�|�Yd@pk��7����>Fl��#�b��O`���.�%�8�N�m�t��
�.�)��J=���y�?k1�^����)�q �(���݅�2��x�EV/������u� zVEy	�����r�c6_W7y���.zWrs�B�����,x���A�<�3���LH��Gzae4���y�H요�Q����U�$=���8�K�Hz��vPБy������R�T數#z�ч��$�k+�r�`O��\�86]�fy���g{>x_O�Or�C�Aǘ��Г�3�.ԟ��J5����&���CQ;��'�i���,�n7��Fx�P+⑏7k��Ġ(\=mdu�	��cx�ʠ���ǎ�/K�c$��C�KW���Y?��<Y-���p�~� :�X����K>?� �p; ��[��O⯀�nz�j�Y�� ��$��?�o�t_��L����:it�iUd+Bm%�"|��>��h�-<i#�Alv�3����u�В��5tr�y��[���ȍ��E�������6��L���u�l5��L��|���1F�n  b�a�4`�����k��-�����q �2�<� ��G�`H��+�S���ؘ�Q*��*�S�䅄l�����r�T��ysW�>�^K��~��N��9<�u��<S�B�
���h�f���6�a6�L����+�Mw��!_'i���~�������h�׉�3�����<}���H�z��9�Bb �<�8�����I?�4͛����SQ���T9�Y�K���e��XW�Tq��M��XR���	f�A��ķ�wG�<OXx���.���������*wsy�1~!�:����"�5�UɩD�{���~Z:�! GB9��1�5�A�w��)�{���mt��Z(�[�V�9:�˴��y1�;3:���ǥ�4���"�Bj=N����M��o˸�U;�v��4����k�׏��"&h��At޺\�L��Zw["n�4(���S"��a'�l�ӌ��ݧY��G�����<�3}n�d�|�����J�����:ƅDB�=o�;����\%�C����:�lk�,P�������ƦP"hl;^/�b�eҷNU���>�M�K6Áo�QGH.#�ш>tZ�:�4i�"?,��Mn�0�Pz$��wP2x' ��pn�ZpU��E:��m��}2�\U�d�<g�K;�=\��ׂy��g٨V�/�~D(���[I���G����ʚyax*���%��*2��_S=.B�:�Ȋ@)rv��u���0p�0����æ���M�]�ܓ�#����"��51��#x3{�_ l��Y�W���^�9�!g���%W��bZ�V��k; ����C�,?B�8д�&�K�k�����~����`ku�^�u��!�B��S�m��k�D�D#i,�p���3F�-�vU�Q^���2 -> J�T�@2@���f�p� ��6cU���[��������ʦ~�yɊ�i�T�?	��/*�fD���n|�*N29���;����8�/�:�ⲇ�����v?8�4��ш'�d���5�'�](���D���~�A<xD����.�ip>�O7����=63�\*.�d�^-�hL�(�ɫ���d(�b	�:jtʼX����j��9Լ���_l�De���p9�TI�@�ه� ��lu'<���t�����TP&m٣�2i�:t��p{aAz�i�og��tږ�&^zՓpMҶ|L�/Z�u�}�3�Y�ᝪ���z��.{3�T��[N���'x�g�h�o��ҩ��ВPm�i�jDj�ϬD��-1�ry��U�-�t��ǚ0/��3u(m$�It?��,>/�ʏǄc�t���KSX{�H���'V�Φ�l��n5*і��*@�HGpi�ϐٞC���!�1W�"����>�-W���ˉ�9�-�J%�F��M[:1�~��h�c�z<p4��r�*s����0w��n9<18��_R����X%��eɂ��~�f���Ml�"�Qx����*K�<�Z<_����G3�7|��D����"3��n�؞f�M�9�3�XOq*�x�Jo=�oo)f[g^	�0܋c�TB4�1�^�u�����)�Щ>�f�~��Lw�k(�|�i��\���\ʌ�������
܅���6�B���ii�����X�+p����z�~�v�ǖP���e�&�-��ۺ%�x�Պd�ѿ�Y�<�7c4M�fZ���S�Z����d8J�"s?1��	u�l�xB�����&����_���Ǉ�C�Ac��Y��[��q�qS���C"ʳ�j�+W����۪�+$� x�ɩ�#���S>b���A�l��L�t]�G��`@�^A"����Ѝ�b��RŰ�����[��j���E
!�y����Ҹ(U���Ȱm���}'���<y���0֫�VvD9Nos�'���ןB�A� o�������B� )3��$�Iep[ped�Ώ�d�ߕ��?L��Alʹ�
�f�����Ҭ�j]��yϱ�e�{�����i�����'Xsj�)�&0�ڿ��0KЧ��;9=?7�i���i���a7Nf�SߥA*t��� �ㇵ�e:�E�AJ�M�H�p���+�w�v>�����G����=�(�R�T4�?o�xQ��P���h��Ƨ��g��Q��&�w�R���������X�y��6G��V�S�_�=; 0�o�ǌy;M���Z	A,d�����C7�lf]d�K�p98A
��֠�����qgبbhZ;��k�)�M�3��w8���Har������"�J���W���W=�X]����"c/���CѧW�$(�ՠ��Yo4f��.?���;�m<�Y$�0�>uĲ����4۝�{�h���8�(���'54������O��prfZf��+��eӔ�k������`�y�5�-�i]k��,����drD{�9:�3)�@��E�W�v���E� ��)�*�VN�Yޥd����kS��SF@Y��|�%��}��_������z>����o`��m�Az�z��;2�I~��d��T�ӡ'�(�)���q�j�Z`����që�/�'�}?��Cm\�����x�����V66���4|i��N,��V�V���vT�h�������/LB�>_���5ڌ��גH���pM��!�\�P��]�����v�}S0�$K���7@>m��:I�E8D�#l���E���D�wd٢hp����i��7c񣻭vsP��+XR��=n:��L�z�Y0su���b�U���D���,fn�aZ;�I��)Dgo�,��e��C����͈*L�����>~��0�{�T��D���t��)G�i;c~�F��Y�Tnb�1��춛^��Lw��F��M4}e�tbd�} �5���yG��
���LS�m�Vv��� �Vd.����!�͵ �9X�AN%v9�&��Xl��-v��b�P_ã�·��R���>�t��ޡ�x��� ̧����II�̇� �3��A4Bn��\Z��|��JԲR��˛�����yb �\���F�d��}�*��;�X���)�|$����W�ݞst|���B���Y�r쟂
�~�2>I�@���8�m���m��D�2^���1��_kGd�ppʘ$��(�6��a[����[��֍y0W�+º��׻6+Ϝ��.���g�!%�µ�7�ٲ�?���mm�K
�z}�H�o?�C�߀W�h�0ER��ni�S��(��j���n0�;�~��
o�K� ?�