��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���q��՛������@�oa�R��Iz1A�#`�ԀP��Iqh�3��F�`�ҥ����c�
K4#����ge��T5��G�z�4��R��\3jU�;Ѫ.Xq��d���D��nmac��V�ܕ�;�)=�(?0�י+�k�襮=�%�YO������鏷w��>�s]��6�t�u�;]��4���!����q��
1�xF!b������.����\�2�X���`���~���4�k2Y�a�w�7=�E�u��#��_f�g�:�S|.�� �֞/^���J���,\*��p�#�0k�|
]c(��7��ȩ�'�Q�	�kR-`~���Zk8�$'��x��A1����Ko�� _'-l_���\��
+*�q�k�����V�LZ\?rŮ5�xwpP�V�22m��w�j�{!��;�Fs����]U�ӂt0���ο[4�\tg�[Bcas��r�����2�RJW��Z�E�CEi�(l�9�bQ�r�
��1j��+�'!P5��ʮX/Ƞ���o��ns���Bi��5�k��>���5 )ڎ-l��HWz-Հ�x�N�������4�qzl��q��ȆG@�m�Ww~Jgv �D��=@�����	��ꪢ���3c�~�@3�[ �zu�.�z��5�7!x¼(��ɞ��9:=�f�� $�To��ͱvA&30l;�ӆ{������uj����	��A@��[�?�-~Ũ)w��8�XR{7�����_i�3(��S�_���"R���;dB��.9P~i���e>��kޣ�m�2�̳��Ay�Y��HDIjiN������n3�-LV��^ٌw�>����e�G������]��L�*�8�h�H�Z佊����,p麵�H�^�?M� >'Se�u�~��xKs�Yg���!ek`�a��SS-��)�*��e4ά�ޜ�L�^8�61���3&P��U��3�~�$�1�2{,m�!�Ix�O���A�H��AҜN3��\�7��yO�s(9%�vP� -�G��}�4��6�%��n�}�#7$��Q��jZ��@�
�����&#��fG���,��L������9:�z�ˠ�_��R��CT�'�K�l���6��&�F�N�_U�p�m-	��n	�JT�aw��Lo6*��k�6@6�0-HC��o�i_#v~�K��q "@���8W"R�J+�:�<��T/ɲ8I^'ېxa��(pԴ�hu#��ڢ��p~Y�JgMBZ� G�N�)�sK��5~� Ine�O�bk�oʈh.��G-�����+��9l?}�=�tK,�4��r����;+�:���fW�P��2ɶ]����/r�Vo�yw�M�^�]CA`�D 2����o��,�Q8���`�6ЏN@2�vek�����|��.� �a�{��C�N�d��yC,���L��S�ة�������O^�v�A9�ba�28�;dV�RwGZN��"��)��ݸ�f��چB{9~0��8:����C�����r!/Ę �E�ӅNc�i�GF��&�(�%���z�JpR���tN�6j�D�e���0u���J��43!O#�:�����묤��΃;��ی�L����ĬY���{�����b�>�y��c�����(�W��obWv�-��(33	���>0d,��)��%6Th�4���)�~��:�`��$p�`�оê=�Y�0���W_)���<����R´��|�R
��F��Qǆ������qbo�M���B�*������a�+�y�o���N�.�t��=��gb<O�t��{S�Q��E�4q0d�A���ݦ���!�X)�G��+`4+{�{�K1��c`֢�]��~�����3ਗa@?��p8��`��ʣY����P����U��k_.����v=���(�9d�i����@#�ԝ5x�r �0�J��Vm-E@݁z�M�eѦS}��N]Bb�Qޣl��!���QX���V��?&���_;e�����*��,���I4Hܬ���4��l���ø,͆z������Wt~,m�aK�8}�ʇ��z�e����r�-�3P�#D_j�O�Xv6e��L�S��ד`LИ-±\k1�T�e�ch(�#��K��3Ug�W��yH��5Q���)��Ĝꥢ���O@�u�L�A2?��Ea	���`X0��Z�(ć�̢����i<����O���g�ɘr)^&
 �+2��W� ��0Kי�`��I���˼=���2S�0��O'T"�b����Y	�_���W?/���
W+;32;:�����D�U{�5m5l�ƐG�6��iXj˻�;�b���+�t�a'�I"��!��-(�
��"�U�i��n��e0ht:�ڀ�HW�Ƚ"Z�U��o�Bl!�S���N�[c���(�?�`�{�,I��j�`#au�$]"�a��ט�p�v�/�����	g����1��c���hi��7{��"�D�B2wt�5˨��q�C zJa�i^Sw��3ğ���P����Kg��8����4�?$��[��7�[�d��Ϟ�,(Vx�\��/���3�rv���k8�m����j>�IN&eK�KQ7nE�����~�aS�����6v)\۠�ˌ�{�E�I���__˜�LR�������� h
 �m���T�g�������l�ߟ��������0^7�������&vlyϟ��Y��:"��n�b��A����K����,�:� ~�H x�ÂD��e������ғr�Y��*bh�/�R��8�_����ۏ/�M&$�':z�y�S�>���9�1��x�c]�3���"��zg�1�'��AQ� /���5�2�`O��0�Ӗ9�贔�����P�ĥ�풩�L�����$hu��Z� ��.AD��c� �y �m{㧐��0l�d�� 6�Ǉ���Ѿ��;�|l/��eh��m��CA����9(%[P7s�z��L�.6d��?x�x�i2����M��0!іci0�M�B�p�b�a�k����#�R	x�~��̟Ѿ_�NFJ̊E���?��z�������Y&�(g|��5|)����-�l���
����@�-n�g���=�u٠l�^�����1Xy���U�-T���j/L�7����z�!] �R��([a[s�Fu��K�m�g�Q��8O��������ʋFc��<B��p����������k،�w��-��_{ej�� �!>ւpL�kiAR���}l6�4��4�ϯ_�>�"�h
i0&�}�i�1S��)4�YcB���B*�)���D���'�:�"Y�Jy>���nMY7����{���� C�8�#uxIi�Y�x��ͽ�
��r�<�kh^ZO0��A��V3�9��D�W�3��Y��o�B���P�m:�|K���u�l|�ˁ19B������m���5���H�������z�3����-%��|n5���e�Lq� �y����+��ʲ�rq/�Q#Wz��?p��s�����'�
h�:��9C�6��o�Ka�r�ya�D����v��U�Fg}���hl�r��z���N���mB���B�S�82�*��<��6Q�����0����-28�ɲ��ԏ�h��[���4��J��P�)�\S@A���������5�^�d�Mg_
IMƒ�ֽ�x��8��'�"9�8d�*`$�ձ.z$�d?&+�Ab7�	��]&i�,��� t���{>��B�V��T��r���)"toZ��n�A����/�=��G�@�t�uZ�JgB�'�D��2���bpu��R K�ذ��!���T,>@9��)׀Y�aݼ����:�����O �h�~q`Á�GXH'z��5,6��hSFR���MuW#èaT|1��/&��7�",��6�E�L�в�N�kH��C�q�ݙ��)�1O�������a;:��B�7Ǹ��[�m�e!S,k�ш�#eF�#Q�(�A$E�9�'��Ö�z59��w��z�_�c�s��H`��8����o��NZL
7 c���
D�-��p��t�����)~�g�V���?�Ǝ#��� $�{`�[�>�iopj����.�FI����sT�����+�Yw�f*�`CP�����%U�����O���05�P*�uM�́����<;�|x��Fk��Hv�5х�}9ʾ{W�Q�"��� '9�J��QiH�8�f����G(4��^��),��b�)�$��_N(�B�Nz��6�@�rNvG�9d�.��HҢ�'{1|kM�`_p���؎���6���,1�E�����N�����S�������:��5��QǏs��;Կ�>u�.��}�5L�f���8��  ���:���y 4��^@R��إ����0X@�	�ɵ�����E��O��f�x�����O���f��E�)�8[��p���!��C��Yv���ކe
��¸0�W���i�&e��sul��B�2��Z��iDdP8�de0P�jT]�4���x_��a�8� !l�wG��4��s��s��m���⬅vkWE�o�5��;<���ؖ�þ�Bx��0�)(o�⢒�fMa�dk�Ȱd���ɥ�+�Xڬ+{�a'Z�b�_��\QV�����?�9%�f�	k�l��㼨��ZJot������f�*|�7yۺX�(�F�C�H�/��'�_�+hv(J?6�4�?�i\�B6�o�})��D3l�����9m� �߼�	|��.f��yN2�sGDn9,x��{�g՚H,���g�V��V҄��Y���%$�L�m�C���wm�.�6t�*Vm�%�wT��?$�y�
����cK��ݮ�H��J�v��F�C�,5G����JM4�B5����}6-¨��EͥH?�U�)Ei�6�+D67���9�h����M�rlHL����62�h�����o�w��_$ �`X�8wN[>{|�a.إD������|6e���7ޞdׄ?��J�Lj��\o�����_�����ϖ��C�
��X�2ɐ�˼�ڜ�fJU4O�� [*�.?����p��~__sK�D�r�S
�� ��(��y����A5��V�8ڼ��z�:eQ��]yee9p��~�������2�/�uU�Y�,mj����ɾ���a!2����#�b̒�M8�4"SWB��͖᮷�I[�{"����^��إ��	+Î� �2�ɨ�d��!�b�Ö����X�'�D�k0��蜂N�Ӣ��@�5Pg
A�9vb�Mh�k/`-ce�5b�Q�8kOj�k28�RXȊ�bU�)p1������r�y�9�sC�=�&|+����Z��6NM�<+��a?	B�=��B�r�}O[yML5X��TFP񶡜��WЀ~�9��@i�:���z&��jzrw$<\���	�^=k�M���0�S�~D+�6U�$�U�a_���!&���3���DmYn��Ķ}i\ė��sE������nk2g��������؆��О��k��v�)���u�?��1�P��Ѽ�@�c
�$z�zm5�|���%��P��.Z��xR2�#Of!�GYj��;��/�aV%�}���>��&G6}z���H����e�����-�bт���x�Aj�w=���v4x�(�rI��b��tk����zrJQ=n�5�P���wχ��d�.0M+�^v�?S�
�=TGR�����g���^;���B&+�ҞH��gV�3�d
�՜`��VǓ�� �E�Μ�c/e����ue[���FBO�Zs�ͬ�����"R��G�Ƶi	O_�LC_N�������e`�ځut�x�Gѷ�-k�y�@Md�:p��Z8F%P����tu�f�5\��ۓ_��'�������ym��w���!�'�CT�b������v����u���&B�!(��y`��`I���Si�JF��P/�N-�z��ޛ"��j93�Iz��D�e��Ti(�Ǣ�.�,ܧ��V���^-޻7�@A9����uo�]q�o�(�I*G��fQ����јJ~��Q��P(0Ƈ.�\�48�Yx��D���sE,\?�[Ji(WvV���ydL��N ��B��_����H�E��YX浓D=����2�U=j�S�	��Tr��]W�ͬr8w�ai��Ĺ!��ͭ��X�ꥴk����~=_��L#+�#5��v����&��x�����9	C�����D62�`��o�̍���
�HX,�m3P�K����?Lݥ�ir>�#�&�%�R���*T,^���C9���C*�l���NU-���A�{h��ƻ�p��4�ʹ�JB��`�^�85 �?E�?�ꊲzX���:;5�����*�����S�(��*F랁��1A��Q|b�#��lB]a%UQ\#{�%��B�r�Nr��N>��Z���K��d��l!M��O�K���(p���mANuL�-�ZĒ k.�W$�kf��잵��cC��H�y�����H�4t+~`��@y�yNL
!�wL/�����f�'���CjL�Irp������_^��j���F�?/� ��B�t��ѤqwR��[��l��OY�!X}���|[4д��7�Yrsc��)�.�μy	���N�-�"z�9
\�n4��*��B@�)ZLd"@[�9�l��� h^P"#�����J�.iߗ�Ҿ��"�O�2Q�)筨J8�z�}d��W��tn�g�~�=�n��1�R���3D
���ۊ�Ӹ��2�M�I�!s�i����Z��+#�*��{'FW#���B$g���ix�[��I��.9u���� >w��j��s�n��{Ѫ�FBs��6��;}x�;{]�ΕuJ��4��/�H��r��O<��B�����`մ\:)+������݁����Ps����Ae�i��4��]E�t���v(��݀�}��1������뺭cW��܆�ٖ�� �|@��p��R���Cx�ޘ�e�Þ��U���@(��G�Ƹy���k��sm���}68��y���3��}ۋ���.8����ӈ�Z6"�r�*�8(�G:��ֻ�,�ȶ���-��4��j�R�*@����{�'��!�=)XKDt���~��L����.9�����M�SS�����24�/���d�Ly03�[�Mf�/4T5�%�� \|�1grx�[N?��2��0�fm%���&�Vb�J�;��*]]
�@a��&	�(=,k�5�I�r���C��eer�5�a?�5��Q�NC�X�xG�eG�j���Ѳ4�(�E{ �`��u�Z!r����8܆Q��ZUa5Z#��Kd�x�`�.����VA��9�����'�e���/�|�u(L��E���k	l��M���#%���6E���)��r��Ŷ��:��*R�fۀ+�]�a�H�ɩ��ȐX��9�V���Se���N�]i��H�F��q'J�a�$�j��[N��
K�W�u�@S͟�>e�#�JE���3KUM)CxH�9�z���B;��b��b-#.f5%�O��M �Z7�����p" 3(+=��&+��#4I�um�_@��Wo�`�L�5HT��*��V<H�s�� Y����y�J{N�����ksX �zA�t/��\{����lQ��@$�C���?�����0c��t<`��{�<
�<�CrJ�5z!/Ai�&ӌ�j�7��5*뉋4����$��C����&����$��#=O"�j��z����
:��g�k	�<|hs�]A�m���99���ޮ�TTC%�8��9��ʎ�b[J�vl��c�=Y��c�7��xi~#L]=fz��c�A� ?��Τ����BX^�R��Aq�.�;�B�.�{=/:�[���S!R	�k��7�S��{9�#�-q�v��v�bJ�'� U��6W��&�DP)�Y�E׹,[&zr��K�=�"�њо!X���Ҽ�Y݁�n�3R�bN��O�
����x�E7�Ď�k,j@KQK ڹd�����E�e?�]	D��ʈ򍖀@��K���X)9��^ LF���C�@��:Q�#z�3�w���Uv��A��+��}PK*�K��3t�#P�Ԫ8���M����%lS�U��m0�G.Mc)V�%������}{�ZZ	~����S�������^�y��UrQ`���T�9�/�q���Ң�%��5�vz>�:��$���`��N|�#��3�/���ڌ�"�3�am�����s�Q�-"vQ��،������Bt��yB�Ƙo��&Jg�"�N��u�?��bn����Tp0��2��x��|��w+����l�řx�;t�	Ϻ�;u����^��Q4RQ`o��;�l�f)R��1��R}�/�uh`�h�~;��w.]�0�7bq����3�$�f��N-��?���xK�Z6'��)�z�j�7#W7��cW�:}Us4MǦ�+�� cAɄW��d9�3\Z�-i_�]�<nT��*�F+f�~�jG�ɨ<�  B�Ɵ�-��Bh2�z���v[A��VS���B-��'����[��{����Υ����SY]S�?2D��+���#����p���.7ӣ��ب�X�v��t\"҇�رѐu'�K 3�QaE^e�P?��6��y�,��!d�2��}�82)И صW�>׻q�O7?�����s�M(�a<o�L�m�GF�n�YG�`ï*���_yg��AJ�E���
{�X��I�R�� �U�oa>c�c{�s����f������`��׾P� �剐x|5�]K��*�.�߆��>čڹ����J��3E���$��Y�P�A	%�8*Gd!��wy��)��%E9'OYG��Ǌυ;�P7A���I�J�t�U���h�19B���To�Z���T�T�p��0�����VP��x[|I�Ζs�H�Q���o�e���Ӆ��NզC@��=�Nw�*�tN���m���p� ݁²�5"29���^2¹sIj���9��<��͆��j��QR��
�R���t����Geۻ�|��2%1l�ھ�+�q�k��L0����(�!��<j�����r�%�J^��D?�[;�B�Ր���/�}Ru�T��ӂ�����h������s��Q��D�d��N���w��̌7�}a���0u<��E���G)�[aV��"����sl��L�n��R���ΘM+tir�Xc�MϹ��?d4�V�D6�WGc[��t���6$G5���c0f=�������:-�D�"}��~5ك^�C_�Xĵ�k�?h��*��̓ �I�C�h����zu��Z�%x ��W���*�3ĜXCĴ4ỳ����y �"���#�y�҈��A��_~n���t�VvK�5���Z
rҿ�>f{�'lK��2�r��xG(_����8��:���]����Wxdj,��״��5' .�n�5��䱑T�}k�+U �yA�.Q����i�>G�V)F�NJɛ����3Ceݿw�E���7�ū�u{�S'U�X+��ŋHUeq��O��n+��Z��ѣ=5C�K�31�HV�1`X�'��mtݯ�^Ƨ*Ѳ���n]/-��<�욼ot;G����R��~*^+~�K�N�\�so�t���'��'o==&��A�����uik����g�y���v)�;j׻�T�9�8��]�u8�O�؂���y�G��j~n���2ᠨ�Dڪ��|#��o�t%%�X��H��lV��M_��g��;4xMd?P>#��(�/6�{�R�\���A�?�cR���^����ml�#��z�kնb��W��7�+Ÿ���˕]����-��7x��qE\Yk���H�
{��Z�RN�[,p����7J¦$�B�MJ,�G�������.vI�SdA�J�
�� �O\��G>�����p�SS{v5f�i�����l�?�&���r�x}�;��6�؏&�yNa�~\�7��`����X6%_Et�?S�y�����w�̎��@9K<�5��I������_���"Q'~�4n��Tdn�((��#?Y6C�֡ ��gݠ�c8By���?xw.�p���C�sF���x����t3܃�Q#�ȡ_�'R(s�*?�keA8]RAEN:*�O���|߱e�4�-�S���������
)=��.?�6kz�m4"8W��8�M��4��*'�(j\�݄g���z�X���F�p�^fO�L�<�|��2�/�\�j0�����"�۬}�|��E�35p�.Ē�'H ep��Z4�lW�B�����ٟ�QPc7-\�
�t�K:܋H�M�����l.B�y���4Z�D����q��D��Q��2E�@���l4LO�V�W}���q�6l�"��f�0<e&9�$��#���qp�L��������u�TnK{�),�C8/ŭ[��s�X�GfL̨���{mU-̬��F h7'�~�>�;���