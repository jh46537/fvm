��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z������{4��� ȽR{����_b�Ǜ7���`Ĳ�v3�ޚx����8�C^J[*��A�8�d��O��ìiM��䠒s��zTn�^�+�^ u�?�JUTQw� �C�˔��g{���{����/�R�dASxY��1t���5i?[�4�RQ����,����g�V$�r�-����9;`	hA��g��O�as��G�	��}��Gt�y��� {&�ȵ(�����OgO3����Q���~m�
�5쁄�e������ѐ�s��{܎���94���b�����ÃZ���2z�Ƀ��2��W����>� yҷ�lҗv "����W� a?_q�u�0��ȷw�~A�`����3�܌�����*C����t�S��A%�ܤ���"�d�c�KrF8`�����&����Pmvg6T�~g���p�<	�̅]UÙVngT��׷��р�/��fW�T�h{�����KW�R9i�Y��퍐f<0���w���z	귬�������a.j�P�g�%�`*-j4K���b�x��]&6�y3GOZ�Q Q�
pWvw�FR/�v�-�j�c|Pa�P���d��a�C��/z��EQ�C|p�K�
���1#�4C�q2��F+��Q����3�vy����1N+:��z������9'#���5�s�f�w֙�����Eur�?0+�kW�)C��dV���.��_�Y�ܛ݅�#_��kKF�4�U�D�$q�e�y�UyڣL�dMسXwR#6���c��_�g����?l3���tȷTeY����2��GI�yE��9�5@?ǆ2=iѬ��Yl�C�?_�kIe	����i�Hϴ5$���y����Lk����h�|V���L�&�EP��g��,Լ2���]3>ɜ�>���t��r�d�d�qf`g��^M�e��RG�|���	�л�F��_3�n��u�-K�s��#p)P�������Ԣ�>u��@���L@��=�Z;�'�S*�'�}G� �ƮF{B[�,2x���;��5 Bȝ�d�"B�ͺ!w��Q���d���uC�,�(�(�pv�	��2��A��\]��'	!��4�l��sm�F��*�!���n��'���qz�>�`�O|���èr��M(x�e��(_�����h�4�#Cu�.��q�@����?������m3Dr肜nF5-^��0-jE�uYJ�wб;��M�f�1��^�'���\����T�,��f�}�3��(F�Ď*��J�nT�NU�s]�AA��~�h�/n,��7w�o?fu�E}�k��1D9�S_�C����{�d�����ۭP�H@e�e~,e��#��Q���~>���a�{�ƅ=�X�]�����瀍��bҳ]XH�/�J!k��Б<�fƗ�LS�icmV��Ah_�Y�����2�o 	���h����M��)	�<y�7T8my�������_�7���2�U@
FriШ�B�]�՞�y^ܸJ�p)Ґ���G/�p3g��v,�5(��E�_g���*@i߲�>��k��oB(LN7��4���@S�Xy��%Bhgl\`�1����>������IF�W�"><�K�"�?�5�"Sp��u/ݥu�S�e�u�������r>4hC8%\'�X784���)�u�r ��F�;IWd[yH{o��.pNJw @�+\�d����z�VÌf����sv���	�����.M��g�����g�T���i�ø�p��VNA~*�<[d�/�,8p�ݳ۵�!΅9�DXu��R>�FK�5��6�8e���B�{�&��/=J�~���Iz�p�ь#�Eڲ�p��d�ؓl��WSj9m����Y��ٶ8��0��/�L�`<ɞ���4���U���8�ٿ��֒��A.q�5]ɟ[�23TgҨ��nP�F3FF��@�c��<��_������N\�S(f�
���[�v��ܸǏ-�m�P�1�)�U�r����A�C�?����4t^�<~)]=	ߡ�����/q��l�X��|b <���֥�˲g�FRWbE����t9���6������ʁ�d\��?U%���<-�?� �`@ϯ�%�z������FY��fY%]%�ԇ�� z�?�1ƚ>��$
�k�ON�, >p��8bA2#� �l��b��xq���Ҧ�ʯ.� �_�ni����[�R��?��Г�c�1TǴ$��\U^�g�8]�z��on���`���&R/�a�֛­��
T��6iz��F'=�tO�W،��p?У후N�Α��(p�BߜA�$^��Y�P����C �H�Ӈ�+.ua{Kc�Δi����/�+��G�E��Td�yP`�7�)O�V[���F�2l�v����Ԫ��\�=$���<����3}�ܳ�r>*��q���nQ+�S�ܓ#��	�(\�0�$��
����������y�[)�W�/:�Ycx��W��b�!�"ib_Fn�3����}��H8�v��=T�͟�k��"��%?�IB*���?�Ϣ�
	Ǘ_�O�@�/���������.��fU��g}@�h>��[��/J�:l�Ȁ]/x�;p�TM�ڳ30�p�R���	4�̖^)<�6Ѱ�~�e�F�x�Z&���s�� z�0����������3��K�|]jo���z����!X����xy�H[�T�O��$�Q��#��rss9�xO��^�ԫ6,���Z�.a��8�Z{,պ����:�C���,�Նd�� �Σt9��x�PrM�CJ(��T��º�t���Fç�����S!�moB��dġ����C�h�U{y$��oF&��R=�v��X���Y����đ��G�.u�c:����5.�G!��FZ�����|�vw��sJ��am�1w+M{D���Kh)�t����Y؎�pR�u(��]Q�~��BسSb)8Y�>ʱ�g*~�-�6�{���Z�����8��H	��[=���Kn����.������zhu\�[)�xU:�7�v��䇯Y�OH�+ʫw	p�����G0�3�MWrVa<�I�!\`���*��,�J1����W�~���źwF���"C�=�m3ŗ�]�*2�"kb����vP�y!��-���$
Aׄ�����w�w5���@rn�)�.���P�ęw)�#f����Gy�H*��pY�$7C�w?�'`:*nF�����1�L&ᐯ&���WyKtJ�|�Jo!�f?AI� ��-�%a�� βOE��ᩪh���5�g���A�a���^���A�������P�H���1��ޅ�1���}��z��\��V	��؛䗚Kj�җF���H7�Μ���p�Ǡ�~�θr���o��A�g����K�e��Gs�?lxM����l�4G��P�M������/4&Ξ��Ź�g��'�2yOe�c����a�8ā����;�+Q���{,~��Y�~�A�2,\�=OR����iOzѯXM�Ѐ��qk84���i�<�u��mB� ��R�{�� �Q�]R��$ߦ�d�k9��cәϘx��R��+B�S9���B�������)$�V�4��Ѧ�K���XRʐ� K�)��Y��T9��e�O����a�F��/As�U@PԚ�R�h��3ʪ�|U�#M�&�Z�8y�mu;�%�rHm����w+��*�����i�����f�d'����)uVp���{2S�U��@�������#X⍷� �񭡁��@�Q���Y�D��k4/�(�5�!(�k���~r�y���"S�-���4äW�@TƓľ�1%E��٭�����Ԧ�lۋ��L^#�T�T�k$����N�/�N��|]��TZs�4L c%�s�Oήz�>����xG�XE��И�p!�B%�od����`�8�4%[���*rw6� �ѐB�Nlc�����xKT$�U�#��؁�8�{�8��lqc�b��_�l�>�b�:�"�	�#u4���V@4heἉh�~9�P�H�������]9S�-. l >�`øj

.�^�=ř��ƕ�����օ�>SO�[���sB���H�ϢDLyh�L�̄�+�b�m������ƌ׹�=(�}�.�Ov';n~<�n\�^[�@�]A*Y\ �m�_Hz~�q�\���i�\�0�p�#���7ԱۡC_ʄ�H���V�U�7�w�%��&(�^�Y�3��|)�9��Gpx��]�K��ZVkz'�&����2�)+N[_O��r���F�!sߒ�2��$���V?S��@��Z)�{M�\��Ԇ$=�	�y���A��ۍ����܇n����'��Px�v	~��r�&m]�Y)h�!TZFb��[��yd�Yh�hJNrq����Q67*'6���4�$�V��f�4֘���;՘K��j�D.�7�Jpȃ>���-*�bI��|�hj\�.%Cq���gR{�C��?C��B�v#B&�l��m� ��$�X���:{��c�@~q��k$,+b���p�a�`<-�n�{���"]�	Æ(xEZ���]0H�@a-���CR�w���w�jq�v;�u-��P�����U�r�͚x��3�h���J�7}��h}m�X_���Պtlw
��aWw��AC�irEmL(M ?ƻa�\6�Q`�3K��C������[��?x+J�ǻ\�����K��$����43�O��#�(���9[�e�Qi$)�5$�IS��gX{R	dɀ�r"W	�#��A���]�8N}O�7��u���f�J�k��>�/���$�0t����y���UE�bB�J�N�j�d�_��0f���sK�E���]?1Up}��v��ч�� �ɸrq�R}����+�"ʪ��{�IΛ@�o�q::Y��tS��?���-u]��LZ�	h��xwd{5NG�~C�~9?��	h�T�^.�Ft<�:�u+��m*���Զ2��q��z*t5M�'��<{c*���'��'G��������.J_�=aeG2JB�"u%Ƣ��AF[1Q9��9���5�n���)�_�@�֒ݧDfuV�I�]̆��`�j��0F�0(�U]yv+��}�l��p#30� ������
:�/�P*?<_[�_XL�Ϩa���HsY��z|w�a۶Jlf�R� 5�rV�(���ESªЬ3��0���=8���2Ȕ����r2b���#�+L�7�B�j���Q��'/���3�
��AD��������;>.ׁx+%�Y+:�t�\S�BK���!#yd�!*	����>]�Β�d�9>ADE7\H|�}��w�kc_���������6E��7�
H�EG�EVM狜RCY��~x՜�c [V��pz���U�ȼtX1���3������Ļ�N����y������x�:ڇ� ���w�0lq�R���(�1����G3_s���P��%|�1O$m��+*�O����/�ri��Sb48��t �
�5��t�*��.�����xW�jj������8ZW��YC�6�V����t�8�C��`!�C?K�?���5���C��-�3���{q��5=5������Bn�`��%&ð���Q��WB�D,,�k�?����胾|�	9m��Hu���^����G���R넷��8R2��MjpP�'K����,U�H
FS>ߜ��l��,Z ���͝���
<\~��X�e��5ɴ?-Е�&��}Q���~�U�\P*��u�U�m ��t6.Bj�Gs#��u��
��4dZ�=n�������ϫ�u��[dm� �?��䳤�M ����	���\�nc���PWoI$M뽂�M}���-���wP��O�t�+F�b$�;�ʆ��<���Ok�ڂJ"VbfJ>0���a�����ޚ�6u��57����?֣g��m�\�U�qW��6��;�f	4�%&2	�ddzq{ ��H	�Ɵ�����]!�~T�a�ꪋSU��7��	A{��!.b �.@-�d����j��`�g�S}�SFE����h��F�K8R�´�j��O��񤼝}D@�����ז��Wc�Pϔ�2u�!>�w�CCRW^�x�~�֛-�y��r�л�̯g�%QCaĦ�h��������>R�R�\�Ǆ�������o@?�a�'�M��L6b�0�o<�����4�_aH0m��*v�a�I��8e�©/�+߼-�.���^眥���I�we�}�O�����9�`Y*5+/P�ݖ>�R~N� ����;���nE��SB�itCk�9	 �:�Y3��F�
�ZU���($�E�^e޷�~���n�/Nz���O9��d��v��U6��N�)q*�H2�`hZ"_絆��L�c�ɟ��Vg���g���}hG�����-"P�i���W�=�^���"�9
��^�\膝h�y��
��`���'�H��w]Yn�`�����	h�ֆ���;=n��T�xQr�3�
]� 	�&K���>[��^�L��$��^�[��X�^��`jZv�iܐ�#�o����뼒Zj�PGG���������1�0���֬&���W���ͪr���]�a�`������M����V�84ֶ�KC�&IkM�ĠDÛvk`,M�_��li��N�`�߼�\�!z��UO��^�~�P4H���v(�X��"�@W��5�:�T�/Yn�*5�1�+=ƫ�v�C8���'A��� X�0����<g6�~ꙃ�Q�Aک�'Kz�i�g[�K|�lX�~�&õ�<����~��>�eD:;����F|�_�pԯ.����-���%�∧��u�;vMt;�%��u���l��ݚ_�O_4�Ç��~Q9E�mhV������a���(H����FK"�Q�4hT��oa�����d\��B���ϟ��M��X��9B��p�\���dQ{��� x�}9�~x h��=����,o��ȓ˾ΏP�{u��A�!3�v�.~�0|��o���y'��@�DZ�� b=�=��_��SR�C�0�KY�>A�9�tnF4mHU����C,���i�#�P�u4��N�)�Zn�HP�4�Z��"� j���{�5;�����Ϛ���1k%��ڱ�Y���)�a��F�R&4g,�����؍ ����Ta˙�{�=��}�K�H(�,�#����w�����e,��|�p��@ǚ��:z=��9����w�4P���	%E7f#K��)%�W�[1N!�7�N���<��C�#%sZ�-��@��͸�/v���K�%�����OAf�a~N69F@�!2�ku0���Z˩�83t^�. xr��g/�9zV#�:ϼVC'�i��=d,9
���䘱���qT��fg,+g���`���
c '�q�m�) ��1��|�jB�*R��MU�+e�_U$m�r�*V���#%'_	���-���|p�?Y��R�Hz��Y��-�@	P�
�_7򼏣n�m���Ԣo�I��|L~qϕņ�������X@7���"Qk�jϕ3�x��aX�n`6gE���g	0�w��O�[����J1��x@�Wc�B/�0(/���C�N�8\O�51N�����}AR�Ы�5���;zi6��Օ/��'tpeWj8A�z���nN�#4D��gx5���y�h��[S���E�9��R����n��ddVbLo�rc"N3��Mn�ߛ�Gfa�u��x�H����D0HA�P�fDQ�),�Hh�+е�7u�یvF����{&�r-}+.�=��j��6Z�#"U�����q��^��J^����AM�Fn<ۖ�W� �-� R�
N�a"�ю(� ��z���}2dO���]��e�tcr�0�lL�/�ꙬeU{+�N�����??�.O=��������g��0 ��7�	�/�f�R�B� �j�Ⴎ�1������䛄��B\R���z4���d u���0�Cp����n�cJ�qԦ-Z_>&��
��zw�6I[=Ӄ��Ivu� r�Bs+�XASBL���ᗫ�B��+���Wk��/�����"��k5B�X���呮v�E��At����y�p�x����k.�<2��L��z�w}�O�846�Q��B9�Px�4��R�s�� �9L\U$��GM6����C��U��|A��n2	�q��;�[�=�R�&��"A���L�ܭ���ɔ�'����4����q�����&w�
�Ǔ�/+8py�/�b�SW�7����C���&�~���Z��]���_@0�V����Z�B_�W��I��:�WP�r���{ӫ ��=�R�Ny@L��A|��Q��B�X���O!��F�YL��3Z�7���س���^�Q�����Z��+r���!��0�Ao�����L�d�_�<'�L�g���=���G��F�oAr�C?�1�b�5�}}+и���N�ԇn��}�!`ſm�b�'��'��kz{�x;k&JT����<����MD�&L�6/¡�!�P@�@\��I��~\�t���1���������$��Ay�MH�f��Mg�����B� ��j1;P-f�-������N�+I\�{�C��H��.�*�i��V0}R���J#�
��C�'�a��jP�%���$����^���S�ᘞ���x��ve��r�:|<��<;��HG)R+E�U���*:!�C���b`S�Ρ�.��T|�7ji$��R�^p;�u��%�L!��V�����o7Q���-��+��C���� ��<��&�]���������/)�`TA���x}���A��A���:6:�K�'c���mOu�򘅽��.cn��L�AސSE|/ZQ�!g?��a�Eb~<QI��H�Jږ��\��LX�LY��r�ʅ�ń�E�q�W��8�W��`�Mz�}�p�n���iO��{c����O��q����U���Ҥ�I9o5��6:o� :e��ǭm�peD�h��K��X��y]�oI�v�C���#�}8��~���oTR9���v��U��^=σ��o�8G��y��&�~;��ÇG7��3w��:���x�
>pC6�&�s%��fF2���4||9P7ܠ��-��7�����+��FB���8�d�Xr;��)�~L���ߜYAsWV@����`)�ǘ�{�����E�����!�}��+����w�涴)��XK�f��~G@�s�O��'�����ׯAxx;ޱ(�,V�//Hy�w��{����=��xp�2)��n.�%z�+���OM��Ç&@�6�J�I�p2}qPR�F��r��M��`!�.�V�1L���'L���v��
�)𳏨-���	��yh�#�r�T~��O��G.� �w	kS�{�ߜ���FH�rs}XV�5��Iz�֕�;�*=�%��Y۲qO���o}؉�Ѓ��4�,Q٦��#�w5��g���A��^Njs�&Y�$Б&�KR��Gt5i"�r�~1n`,���[y�#-�bX:�Gw<�<2����{#,*%�9���Lg����xU	2�$���f�~�3���DS�0О��쏢z��R�eb ������ z!�w�_\���O}�'�{/�k��IN�b8%/���c�5��r.��a� u��ȟ�pI(�QRόq!T�<y����W^G�{~ȴs���*��U�V�!;D�9�m���MjY��������?��I��u+s��=��w�@{� ��d�p;V|x����.M�94�O�+y�Q�U���#��Kwaq�W�I�����[/�u�ws��Q?v]h��^�bZo.�������t���c��d�~��or�_�f��R�Y�*_E���D��J�_���Ioݶ:U��-��:�G�#Q(8��܌�?&�� �W�R~�]$#,���e=����г	QE��_�"�j\�̅] �O0��e�m��f1 �v:�o�R��Q��c��r'wr9=�r���bv9�v��r:���Qzsӧ�I-A�9��'P	�H���\u��uWf�K棑ʅ]�`�}uP���f��q����f4��9�{�(F>��G�MF��Sɝ*z�l\AĽ�4ԏ�Ԉ��t�t�8�4=M���t��� ƨ�}������:D�Q�$X�xv`_��0�I�!��e���z��
xz)���v��N	���>���`r�1QFEH�[��q�8���vXt��c�0o�Jެ���Pn}��&�D�g�������j��#c����b�<$':��K�B*&j�<��g�E�Rjn�:�;�y?�'���-�q@k^6U��� ɉR�@]y/FB`��|V�1��<���Y�B(��bw�E�����g<����fe.�mX)�����/��]���溠��і�nR%_���x�^|�N��0ۯ���	�y�+���a�D��o�7W�^��ˊH|Az�I�~���E3,����R$=B�׌���h�t�f-��k$� X�������Yg�
ų��I<��j������y�����ʼyH�|ƾ������;�M&z)��qF�.��x���x��
1�a���-��
���۹|z���n�#���h5�K��@��A�����/���]A�xo�J���Il[mW/� �k�E�?����za�����Jvs��T��N�"���K�FIk�O'g a���ϨM�1��P�(�ϒc4�ފ�B���m��6<U�29�h� du�\��H�)�e�I�9�f��z(3���ɵ������%��8�m�n�F`D΄�W���kֻZ�4U����Z���C˙0�Z�C�O��\��f�QܴൃS�ۈ�
���R38�Ͼ@���)~��[�,��i����P��t��\a�(Ce�-)��Tf�TƼti�r�N7�@."�<�_6�����<I-Ͽpq늩uMo>yd�i����`����g�[��G*|��]�����(>��̀��[����D�7�H��߉�C ���F�kvΞ��h�Tbf�� ����:9*i�	����F-��k�(����P*,��d�Կ��#\w�b0�����6����p��0X�-�;j�uV|)�]&�tv=����w�(ࠄ|)��.J�2?��"��=�X3�b�
�y|>�ٝ�6J�je�a�h<�mC[8f�����)Yޣ��=2�?0ld��#"1*\G�k�N'��"x�|d�\l��	� ={:���k��L5����-L�R>W��i��0��^���}G~@��L��֙#2�K�bg17���~ �󪲿&# ������7�	��3��+�2>R����%�9@��E�8���I���PO�z��iW���a��CT�Oc�!g��~��4�7�|Ii������`V�]�U}F�5v2��5> !�r@[�r#�5��
_Q��}t1���P�S$O�{��]CR���P:0i�6�BQ@10��Fz>�\��+v�����m98R���3��Ti��/V�e �PV���i����&��;]�\L���Bb���P�Z3�I�X��9Dv�J��On�K*kj�ɮ���""�wD��-�E/<�f@M��s���>yA7�Q���E%	pb�7���<%�X���ˮ"�i����5;C�e��P�d�a�%w�!�O�;*�d����=���E��?�.r�*�!��{�d�O�L#��~��.u�s e���f0r�#1Ξ:)l������(4(]݈MKr{�b��x�/�2���|�1?�~7N�ХYc���f�0ؗÑE`�n�:O����p��Q��<�8��G�HK�H/���}@7�����']���_�)�U�QQN2���{�z���ٖ������{��DK��?d!lި�36j`�-
\���Z�$�85���#/���[�ה�"X���͑ׂ�J~ɐ�%k-a|Af%"8I�coh��] ��v�q'��d�}2"���pq��w�ݒ5~��j�P �Po��"ff�O�dEmuC���qg�W5��w�J�ʻ�Ό��iؘ��~D%;��zT��F�C�n~���'�+����%�-Xw�\��B)^m�~D$ڒ�~�"���kSkLþ�B�A^&e�ި��ǚeB1�W���w����<������|�rU���V�w^?*��h��m|�5;�]���2cQ���-�(���/kz�an�i���iZ?UY�0i���7��s:w�.+����T8�~�+�v=�	�>U2⇶#
�bΥfis���mG�zv����F��_�~'��9<�H��q��$�5S�6�`44�OȝЯ�|��\R*�6�&����u�(`�L�-ZĽ=0��q|�{0����VQ �q{ņ��ؕ�]�����JU�}h,�'ҼUo�?-8E�Ҵ�4�F�����)e�>ŔH��4O�ZE����'(EUs��9R��e4}�/�E�ɖ��n�c�L�hP�b]/^�ti�fd��yV�u$]��FU/ݼ�;�!�b%Mh.B�\����L_}a�$�Ih^�*\�N�8�Gݣ�~/Q�Z [��B��E�[�|^��*3La�1	���f^B���^YW�k,sT�=���.�sw&'.�ˬS�R�Ƽ��ZT$�|С�t�>}
XÜx�	�f���673ZؚE�A���U��� ���?�0HQ�
�"W,~&�;M�
����ː:1֕��䥭䄜�9��hǥ��.�&A3|���>��M7��GK��N�Ӑ@����d�oŋ����ɣUe������*���s���gԖӈ�dX{J�t���k��F2A7G��U�W�N�7��_������]�����QoQ�ܪҬ�7�VH%���*�fW�~���~ꁬ��*���V� c�҅Te��ə�v�������"��uϵr�@�.Ī^�5TlQ<��٨a��e#�KQ/�E�㋞�s�q�Z�G������
V啦���WH'�s�wi�D3D���Y�p��/Z�I�DM�LE���
@lHE��g���g�.��pO�U�C�7[.̘�}ﺵ��O��Q��A�}�I�M�J� ��{��=�+J��-Y;��S`��6rE�7���[ő1R|2�����V�\�����M���ǚ��&���!�iҢS�X&c��X���3�u^d�� ۑW�ܯ-������KƠ�/viu����Y0�����D�����P&���p]�z�2��
v�7GGH�.��Ӌ=!n�9�v` ��ܝ��h�^���*�<iz �}Al3;��?r�{S�D�%����y9.#W��^BIxq`�Tͦ1ԏ���Q �	�OK�H/�2Y�)2������y]:?��0K�V]=�X7�]ԝ�_/��>�zO��p)�*[���E3�sЈo��v�^�����iX�xGr��Ҝ�u��o�{�ׂ>Frm�)��=����X�Ӽ���ya�J-�����熹	W�iTIc,��`�=<<'�'���;S{�����dqGz�h-��l3'L�vUo~�}O��&M�2u�d4�^�v�=�`�ӳ)[gq�]�tZ@:��E��K8�y�Jf�~�&���Z���}^�����R�Q���������E���{6p�sj��gϛ���Ou�87�v�UD�T�t�"?���\�F;��{\�v7b�A���߂�4U��X��0Ca����g~�P��/�ZF�������I����T	:��8WY@-Wa����:�z�i�='=�7�.�A���s���_�f>�:ٶǝ�Tߦ7y����n5�)��G�?�]�dצ��΀���ƴ�Q���/�*��C/yUΏai��{�kt�"�[���`�(�|�	�Ua�R��W���#B��e�-���k��,O!�*��wzl�Ѡ��Ht_��B�J+q߄��:���GQ����)Wh'��o�d4�'�L�',��4|8W��yX憙E�P������߅R� �ߜs�d�J��6��%�����P�o�U���B��?�C�I�$��M������yN��k���aZ�I~c�Uk��::��=)�E���sKL�t�Rm��
�Ͳ���x�m?����jJ3+����>�ej�������*�V��zr�{��
e�O���X�q;},C��(,�"���i`��A}���bx;�a��dC�83ن�d"u
��q�tz�D�k����$j�2���k}�K�~O�M��$D$s	�W��6ԝ3&jUā��4=�����-��S���^I�ۙ�W����qO�@09����Q�a&��4�H�+
��G�y?�	[f�Xm>��U�C�#�
Al��!����*�Q�W��wND(=�̮���7�P35u*���'V�5��+�Y�;]���-�+�W��_��J䶎n��G����28���S,b@�>���ry+���f��9b���5��^���3(骙$~4���~�T�Ŝ���@���=�	��zȭ.B���.��h�>>�6��K�*s��%y?�o��6��S��q���A��{B1阞̓��6;�%|3Vl�D�����*�>kn��Q�/�8��b�$�707���I{X�'D9���|���ۄ�[ �������I�����6��^��C�=��=���oa�U�eH0�&;_&��Ȉ�U���۾m��ئq�������XGD�?e�%�J�ۣ�2q��G2���Hf���~���#����/;��S�>P���ٕio���R�޲=s����Ťu��(�-	�a�_~���
&�r~�~l�f��ɥ\Sv�C!6�Q	�G�~�����Q
���9�"#a�x엿�Nץ�gi��3��c��h:�ms��cxJ�[k�r@�Q�]�Y���9.�0T�� *��8����"�1��,J�d
�9���M0��Mҝ�0�ӈ9P�I
�g\�>k���͒u��x3ҥ��ϩ�)y9��>,��Hq=�:�����t�BA yp'V�=+�9���$��_� ?i-.��@<g��x�0e���F����tI�7ߺ����-X��,�"��_X�L+�Q�	E������ˉ�8������;!���k�iA�Q=�u�Y?5XVy���J�r:j&�7��l@�#o�G���»G��ĭ�/�u�������l�2�v�7�)��/!}A6���J55�n��xJk�HS�����U9��[c^B!4�������#�Lz��f|Z��$rV	>��J�6�s𪃉�E�%9*��H�V�Ī熖ˌ�F_��s���i��8�����~i#*+��&���Ģ��pT�
H��3K%G:�/�p�M���z$)����xa�M�H!��9�^J��*B��K��\�v �G|���l������>��~�JAu	`��n��8s!�C �:�vϚnN��4�0� �F!mlRc"�s���U�:�H!/��LO��!p�$�%�OYk�����,5���B�/9�v��}l_��7���X��~�e=/o��^BI�G�Q���R	Y,�=b�U_G�
I�Zh�ex���O�����طa�����|����6��BU�m��(ˢ��Fع�[>��,���ԥl�8B���(æ�,�;�"]��XkT�BI�ɩ��;��[�L����w�wة^�F���KI�m���w�}������{�@�:"��\� ��p��"�J'lۻ�Ņ���^��'2��Q�a�l�ؙ�>�4�y (q��v�Bz�S`n�Y,^d������[�ȷ����Yp��T`צ�"ά2��Gp����t�Y�}gv$�h��Zag��$������h��� 3@�s���������Ա���D�\�\��X�*Pn��!kjfm�<U�r5��"Sv�i�؉�!u���=��q�?����Љ1y�Ъ�#������lE�1(�����;I��j���b��d���� Dj�w .د;-�L�O�`-ǟd՛�%4l��)I��V��%j����-�{�����%�S����u��R�����l�ѵ
��5V �+�0�Z
7��'���j�-N�7fcL���1P��K����J�$����$�It���N����6�m[�x�J�l�OY{�ak�)�s���d�;r�t�V�T��˝��?�On	`c5����ҏzH�I}��?��d�=a]�om��9���,p��(�`1�(bY��f<�S�BĀI����T�{w�7�FZ��<Qӎ� D,��%n��N���y�X�֖o 6�>A�zľ��A|"t����DF�S�|���_�������Hss�;?�Z�_��ge8�Vߗ��Q��+1� ܫUϫ�3���H0N|�G�j�Ni���������(��Zz���Bl&P7-�4���I�|)�1q��d�?k�~mPŦ��¡�������]�����i�RS!�XA?]q\>b������]2�X�f� R8|)G�A����] �N����:6���Ʀ�
6F�y�?�K��^�b��7�䂼�\�.���	�.Ep������[��&�#�_��{��x���~R�s�N3�/ w�ݟ�rpuJ��Y,&��Yv$�]��Bh��4��A9E�Lv\���k[�³T�|�X��^>�����'5�������n�W*�%!L
�!p�X�闟���L	��Z�B��N����nYE~��{G\�A?nȷ������)Kg~s��؛��	� ���TQ� ��dx&u�?T�v��{v�(<&>�	�.Wp=�O^n<ae-�p�9>n��j�N����1�Jsr�\v�����W��Ӌ���'����P�I��d����SM(�'.��fcB�����M����I��|�xǎŠ�Y��3W��E\W�H2*(���
�1h�l=�T�o
�����z�k��|Z6h��j� Aj�%��w-�<���h��ɖ��q=��؆�r��_��"�K�a0 =Ѣg�
�N��U���4�2N��m*/YO�G.��G��e��kn&Ì���SJA�pi֝�}42�M��7�7��)V�'hҢ�b�޾ݎ@��� ��3����������[N`��K&l��oϘD��2n�!h9����͋�{°�9�\�����I?ߡ�/I<�?�@�#
���$L�P��y���m�y{Ti4��%�{g����\(^��6y�E-q�d-�P�I�=������]lN��m�*W�H�55�.a�R}KL��q�˓m�ϐ��!�2��`JL,�sG�^C�er>A$�!,A�9�Y������ڣϓXS��j��)ubc\��G�^�߄\���� �Ou�c;���J?�|H�ɇa��E���I"�x��b{h�t0G�Z�.��2Y�*MD6�;�����eeτ�)�%)���G���77�	��MR�~B�V�Ӳ�a�]M�&@�y�9�х�7M'8��,z>]�&+FZ���U��~̋k!��O��j�C$���m��;g<����Vz�O�oyW�U�Mm�O��f������J�a9��/���jUQ��(ϋ{�>0R��SZ�ۏ8~q��K�m�c��.sI�iM%}��~b�.Mzc�Iql�!ܲ/Ra�2�bU���͑"[O�O�i}�D�Y"&��C�S;�d��4�M�{C�bh����i���l�-B���bߴ��`�ѓ���65=_�a_��o���-+�QS�����H�Ҵ�*XҌ$Z�����m���~�g�(q��.bsVc�L�;%+\�_kK���}A�Mm 5�,̃�ѻ��nQ����|H�2h -U�(U��t7�>�r�S�4W|� E����N���AJ�bn4�`w��I	�7�R?Y��xHD��x�3-4ĉ�������J�s�<<f�Aj?��s-�K�`API�h��ӝ[��M�%%�%�!�Ij��=�7܅�&������q�"���kާ�1������>����1Ю�cu��_`�-�����Rc�<4�m��#��:wPN���1#����	��+U�q��w �h	g�J;�b��;Z��|��I��W�X7���`�I��
A�t;!�M��֤��ALH8��:L����ӕ7^��J}\s#HyE����x�IB;W3�,Wb��ʞ�{r�D6���W~�E� �Ȍ�0
q��!(OI�p1
���v���F��W]OyWD5Xہg������3�ȴ!Ԍpi��U$֔�`$A��WT#�aۡ��͢����D�Iv��`cb�e�zThg`XV�V��^��i^[۞�����,.����şK���ӥ0���à����H%����U�k�,��LV(?xJ=}��A��J�&�t���>"�׬�J������	�$?|�0|�
��T���u�a^�c����(��H�Q*Z�Q�/	���Ë�[��*�(s�+��6)��B��r�_ TX�o����.�Z B�0��u��N��[�갮䪘�����H��o6P�Z>w���p'[�����gw���-�q9&�CJٕ����R��x~RɓR0E�����S�L�(9v�vkh��ʆ)8�u�7y��QE�'�\����a#Q�F�T��/�5fncZ�%�S]	ÐmJ��y·�p���>��'"<];f�VP���,�uM!e�z	��=�����`ZpA�]Wh��6nr�x���|��s������&�0#^qʍ�K@*�t)B������9M�2���vփ�n|�8<������8|��J�� ʲ��:gj�ҧi}"��B��-��F��n�k'F!+�-��vI����^Q�l*rWF,�o�;�G���2�T�����̣^'��D��1��ݲ����!g��Z�8eV�M�>i{���9�h yN�tc֨{A>�������M��g�Hѻ��9��o��~<�v�A�ߘ¯��l>�'p�?u��GTٮ_/a_�z����X�B���G�?+!>a��A��8X��`H�{Q���[���޷�]��w��C�(F��$��h�S�6^.��2�z�ˮU�ə�u���|1����\*�Y��I�`N�at�J��4b�#ӄnh�s�n�ۓ3B�̴s�|lg�y?u(|�Q_}��e�`�5���W�zC������Q�
�!�Q˃���>�yߣ{a���"-��.0o�#����T�ΏK��V�i����h��\�5�:'.�I3��J.r>f!�5�'��&�Pشȿ���I�ǖ�8��lz�s#g�¼@)���h�U��sb�V�4���2㩼�K:[�KX��ۄ��p��r��0I���
L�N���ː0�0g�Ck�ɒ�,*��	��Ly�b��,:�K�R�@����Z�>�0E����2/�j��:nI�G����%=r=<�����>��j_�패�����k�Ӓ����BG&UT��+ؒ >>zږ�/�h`�ݱ�ö�&b���35ܮ�OU�^ǀԨ���{&���,��^2lD��T����7Aj������ڲV�M�PS)���Pl,a�*�Q�Gt�9[�����a��ؽ�.'l�_h��5'����PY�-a��(0�PY}�`v ,Rk,���1	�{wG�4�n�mͫ<*�S��"�@�<�?Y<E���ӫ�bP-sU�����.�`Y�%��{f�GEH���/�U�~ ���o�u'(I|fv�PMd� ��w���8�M�D"t��J���EhR$:!7ΧG����[�a�4*�g��|go�,���ݮJQ�\�dɴ?��_���i������"����bD�]�m 1�*��;� !�l�#�,�~Zy��z�<W�~r����h�(b����bv������3��Ҟ`<�7�.�Zw
�K/l�Tb���[��an2�uq
4揘�˔�4i�P�	V�S9���L匄R�J�/�`]h��"qPێ�w�sk@��IF��ckpv�tی�ݚr�r���a��FO�$��?b��I5E���S���d{���	��Ae�V�����}w���Z��\�JD?�Z��- ذ%��H�It�iY}��`^d���rb���\�:ؓw5�O[CL���T��6��\h�)YM�ŉk���C}0<�硣x�<jv����)�����P��Լ�Ǉ�h'K,�/q$����G�\��q�-$�;+�ᎬN�CT[a<#xZ�ENc�{�	�dl*�[��]@��
�L]�='ݗ��A�C� 0�tZ-�Ȥ�����K�`%D�ueBR���/� oZ�0 ��D<���|bS+ ���(=�T�ׄo�GC�v�=��ee��h	B���m�yDV���Ȧ���<�y�n2�=��F�;O�m����m�qI>�m���R��5n�`ӄ�O�1Ȕ�Ҝ���R�O*6��1��sfs�����1��+!I�$P#LK0[*�3��7�������v%������ .Y9P
�L��@P;m� b�/�ĭ���	����Kz"33b���?BWy�C�~�PY�2�c��?���ۗɂS&	9$�S��m}�����t�`s�L���°
�:���b,��,������J�F	��Q��v��XwO��."zlO�>��'2`�[1���<��X��ĥ�pY1	���'�̂���6ƶX�(L��0n�^�ߋ�h`������T��[����t3�g���m�錻W��
k�g�i)@��ynr��"H*�o��؏���SN�|�G��yko�i�����[��Y:��s�d�A���n܉�դ7:��'}oGS Ҥ���L��7֎�q��=�Hxm2d{�����U�T��^ձ���hjs��ÿ���_���O���NbRm�!X6WH^������s��l��楑ƵВ=�Ӥ�X�w���,�8����� D��Na
�I�f�����,��f� 4���6���,��UM���M�;�]�������&[���)�~��cM��;.$�Qć�h��J<���Xv�����_����6#$g�Ɔ�O�=s5�qC��9�����jQ���f�(�.r�c\v) :�d���v�\;�.*�1�+��"��u�ܒ#�c��ڸ�kJDc����F㴾jS�>�mvĭ���̀����U).SG�mE}-��:��"��G�M(�eWp��+c0lp�ި5[����������?�z�s�O��y���k�;��ކ�)SC��\c���[(*���Z����$��8~|7�*`�
fq_�'b͢��&�����)`�D� a����RM�<^w10d�N�L.��;5<:�"M���I->������2 MB��:��Х��@V��Nm�����y���u�|h������#,�=bs��+�g���8�&�YF�q��e�^)�f�9�kl�v�m�&�y��xC���>��r���r�C��of�����0;�O�N�G �P�o�������O���t���!�3 �}��|�2���=6{$Y*4��V�"�N�����@2}����nP'���=�����g1ˡ3�ӯ��?I�,nj�9&G�N����6��z6:�����c�vhk���+�����14���x#�+��;s'�ؿ2ŽB�0bb�*e(� �ú�ojDt�z �c(��
+��1b���|���\��	N��L~K��ո���_b�����0�N�o �tz!YU�I+�T�k�[59Ln�l_��S*��\����s�4������`N�D���ͻ֓Z(�|��vSA$��/i�z*��``,��9W8^}H�����_g�I��j��^��_�t�HK��:���ʺ4�$�ve���XS����y�O����V�ѩ�\�xf��T� �N�j<�������wwF�R��q�֯�f�.H�c�¯T�T��2�����1	�|~7L��JP�a�:��oҲ&y9l�,�cQc��!������C�����M������	fk:В_��؜�,��� MB[(��bѽE�1^�|xP�FK�q.5����"T)t��"�x�z���Dgf�J����M2ϵ�3�i\]g�����Cx�C���J�m0x4� ֈ\ P𶔦D^����������r��3�� (y�W�HUN���G���{#�v�>�2�*����F�
SjE=���������(o,���|<k�	��T��i���FV=w�v����	Ce�^P�\� ���5
��!�U}��u_�k�A�� P9���`�5p7n��Y�?	 S:��\e�a������ǈ.bO�P�+6��NVV�"�k="k�x���T�y*SSg��~�"�AU�V�}�<tQ0���)�5��\1�֋	�ÿL�q[�b�
�H@ӓ��h�|M��SU�GJ�����UA�!��B���ܧ A��'���MhԽj ��|��G�z�㭽�(lIQio�4a��`�*@�_����-�k������d��FŬ5ή1zK�w��~.���wI�߾]��a4���p)�����jӚ�\%+�}�S �ݰ�a�E�q�U3�����JO�����p�(MB�=�݊��A�c�F�ׁ4F6��ؔ�
6K`A`@i�>\N��u$�&d���ߧջHNY֞�H\_K=��8&�%&�����p*�y�n�\�XQ7�<���G���Bw���=q�e7޽���{Q���f\D�78m��X�!#ο�=+I��@���$de#�)�`Xw�ڻ�����KE�a�>�'T�H��d�tx������ǁHZS��Z�C� 5L����˲��VY��P^m��x2��A�?$��B�k��֩f����������a�L�?�����CM�
������\�` ��䫺�ͻ8�y�B�9���m���1�(���m���Olq=���UD��V�P�;^�� <&}i��ad$*FÙb��i�����Ή��@|�c>�_�i���&�
t�4�hY�Kb�_���k R_)Ď�	��L��ނ���Rۜ���M��'A�ex�!�}u�N�y(B-��6*�i��w+��Cm|�];�M��4Y���I�.q�s���2����-�^����B?�ؒ>^��
~Ek��k�o��P|�h�y�"&D��%vh|Xy���5�)�zl�4�`����N����̲2��h3\=J|�(��P���c�u	��ۼyؐ��X����r�H��E�STyY��X��#��W�[Ym �����"8���J���c(ϐW��CU��B�V�ʗTw��x����Ow�2h���D����S�T$z��Y��Eq;�Ek,д��jd��?�e�;Si��7���  �x��ٿ_"e-W�6k�r	~�Xd�|�|�TR�.�`j1�z�w����-��;�����_�����fz�U|�S���=�9���k�J$5s�Z�тu�%�h��D�Nkܔs��]Ps���x���.��
��mkb���ۑ�oQ�O��� u��io܊��v�X����H��}�Td��PwRk����-�V[�������h�:�.�}#X�������/��y�k
s^����d}���ރ��%��8�����-	�򜟞�%J"$��w�Rm��-�7�]���0C�fL�w��p
V�'�`�r�1���u}��z)��M '�g��3�5Tg�l�4���s[�i�����x��X*�2<B9���]Ė�	�����r�m�;gH��uO�N�WJ�8<���Dv��	����UO�2L�R����V�� ����q��*^%��`�te�*��Qn44� �h�q���_��T�����b�j��:��\���T��^�@J�C/{�"����B�
���>@<U"ъO��f�Y�Z�b<�b�z�J�5
�"������g �B�2o<����y���E�y����1,p1Q�\DԶ��P6���P�}a[����l2�[��~�z�,h)E՟��p;�cn�&g�P�;��4;g� W�?�0��n���7m63�"R!ʀez̄�
��;�^92�xR���`qgϩ-t��W�պ&l�gt*�
��疶=5Og�HG���a;��@7�棬�d��������^�O���K� ��KA�����7���)��	B���?��:klj[�T8�R��[��+o���t�[73e�`����,<��' �:q%�-<o�E�5]���p�e�kS]���2���u����� �����̶��魀������\�,}0��	�;�gԼ�3���	!q��R&��v��)�=g`�5��z���@FW6���YUѹ�.������-MlZk�KS����GW	�6�3��Z`�L���(��/����4Y��4�p���L�=�QA������ �U�Q�^�-�'���:�7�|���h���@��]`�e��K�vl�~Kq+#^��*qgg���\��E�|UKa ��fhgP��8�m���S�S-�\W���ld�~�V8��X��S�D+��^l�๒j���K�Ax%kd�}o"%Ar�����P�[d-Ƙ�+�ym��m:O��>����������h�p��g�,�ˌ�NT��*�_���#I�9��B����% n
ﷵ�6izeyȈ�Uo
�b6Ԟ+�B���>n�Q;�1kxU0����Ė�*S��u�V������o�w� Kƽ�(�Ӗ�S�B��x����7�K�?!C'4����j4w6�ѫ<I�
Ǝe����Gz%lS���
�"��a�y��&�H�ڪB���!�ho�p0a+�a�2����>�6�Æ�2t�G�@�#�I�q���������f��݃Ԟ�ow(�Mk^}9���%�"JޣݢEJ���Q`/Ъ$�����p@��ʺ/,Ү��8@�Ť�I\+>�Ǳ\$._�U��vN5�߲��xZeM���!�e�:�����6�5�	NoHEǊRs_�d�J�H<_ƺU��hLXԌ�OY>�r8�p<�]�FR�^���oN��Ԝndm�쟇ySo}�K�V��dy�ÐH��;�&�T�5��O���Ld{���/�Y0=�D�↌�Wa�r?��6~/K}��F�ur�z��_J^�?2%>l[rƊE6�+ºI��oN����)!��9�ʏ��DY��[:�ܽ�����%�ڼbP��(v�5C라sޡ��h��ru>"�� �ӏ��9�ĈC�^c	��1> ]iz�6���h��^a�����9ޑ�<�D�fKXY�a�� ��Ն05�5h�8p���>��}��Wi�B0�+�WNR4O� �$��9l<d��|�eR'�so#c���$�6��W�Uw�A��
к�Ul*k|�8��!�G��<��ݴ�mZ��x��;贌%p0�xjq�O�^��?�Z�n���;Օ�<}��_����}c�,R�PҘ�0�x������v��K~�Y���W0���LVS�/p�: 7��I���� �^�}2Q+X�7h3�L�L���,�Ȏr�>x�z�ŉ�0m7	`���7�c��nA��T��k1��9D,��7�M4�b �i����SWS�d@Lp%��_�h�]���DdJR6TU�}[8������|f�p1�0@~��"_���Yi�Q'SuL(�=�>��RI1ke���m�����+�>�^1�Pꢜ\���J����� 5�g�߫�"����zY�K*	"�t�`ɱԥ����A�ޜ2s��V0�.>�,-a
p˶ צ��":��pX�F����/�
|v 	F>x{O�01�]��>`2�S��y���<LzNQZs�l-BA�>��G;���+��|����W4�i���GRv���۩�q.��J���V�:����K�	4��������K�J�D� G����(Ȭt�ӏ�5�_ի� O$,��d�N�XH�ș	+�,� ��S0t�b�+x�ߛT:�ë}N{bhW��i7��f�v�嗢M��!�!71��s���3P��*V��`���E�R1��"�.ٲ"˙�N�i�	2���cɻ�U�~W$j�uT���;*ӎ�F���kN�]��4��l��,
��%5ɬq����x$�ǟ������v��kh_���+��y
�V�
�����8�_�s���Յ�1W	�`�WXl*.AM3kDH#������k����Lgno�LD��y�{BK�}�?+�����H��&�!��S�T��A<�ٰ}�"[��2�$�@l�j�M(��������a�wg~��x~EY�u`���������)xdc�@�><����O��\���;b#���� � ���ʏ��K�3c '�~�U�\�h,$��=����3����N�6_~"�1Ʒ7���6�g��bV%>�'?t��d��&�S@�Z�Z���=Lx-u�/|^�x8�=KZ�3�P���Q�������ˡ4^�Ԓ s���#��/�KY?�ބ�h��B�~Q	�v��6q���!Y�Q�i����~¬��-��+5I=�˧��>��Z�V��k�2 �@�-��{����Q�ݢ��k�P$f&���TR����^��l���#Nbf�N�~	�KC��7ϓ�![�I%x;����C�aO��%�����3a��(-��>��nᔺ9x���=XMGI�� rC�$w�M����7�ـ>ya!����.���m��a��bv8)\���	GRy�W�x����=�,�v+Jy�U̶�\�T�<������p��M�2����;N�Uqh�L�� ߔ�I�N"�J�8��**
�?��>�w�o�c��7R�����)Mܔd�
?:���P�3ݐ����0�M�pf��Z�����J��˛�]��2�*	��l���Ga#��*Lg8l���fF����&��;X�J&M�A$��\.T(^>��C�i��ދ�Ǖ��u Ϧ�w3���,����}����O )F&�������בU��X;kN"��
!�p��*�;��H�6�	{e&MX, �"�}Q�il�~���	Ȼ��4���ߔrj{?.L�xE�KQ3��q�(\� ��о��`,��̈́���^�6+~k�Ϫ�ѿ<՝�ƃ���bނȲ>-MU~t����Á{��[��[�!�y��֕�i���(�;B�|%^sr8�s$���՟��Y؁feN��a�<�Zi=�h�dUl�5����~�迠|��N�:�BE|ԁw��[B�6�KR@�H��O_#�~��w;D�;	���Μn��n�i|��$�Z�p�d_\h��~H�w�ˉGi���~(3��'6`^�	s&�ͼ٦[	.%]������?��~A%xwX�!��K_7�]�4I�<�j��ЊR�+w+��E����0�z�?Q2Ա����D���|v�.�h��F��{��K̪��AY��?$@=�����q�A!���<�c�
�U�U|���^��<��1jB$�S���*�̆�ٯ��J�JEy[h���n�7�&0�m�K��)y=Z��t�a��uŁ�脻���Je^�zzɀmU�"���������
��4Q��!v�~���Ù�Kzʛ�Г�t������U��'���t��4�R�]r�wT�U�?��(=� �V��Wk���.�^� �:kk����"��Po�:SC�?�����/��3��-���������'�ֺ�?���0L��ͅ�$uꚜ-g�Uh��g?V!� ��h[YP�G슌�|3z4u���D�=o����_�X*͔�xg�) �e؈��cI�J�U~�Q��k�S�[�i²��c'��LtC׆H6��r%S"�Y�f�s��n�Ử�c�,��{H�iz}{IhUZ���v:3�TzY[vwI���� c�i
'\c��~ZTt��=�4�sc&�(����sX�c;�e1������N�}�J%�7!p< o�s�D�:�ʈ><�3�֓��u,�6ܝtoq�o�Ө<�_D�J�-�!�^Ȋ�q�d�r>�V̨��?����]�w��g��04"��(e8Q���L��j��F�?����2��'K�jnCL��wD�	���z�W4(qH��";
w6��dʼ��~�)-4ZX�'y�v;㵼c:@��
^Y�|z$�*ό(�����H�F���OT �V��G*�u˯*
�(t �=&������\*��������I/Z���\9��mh�:um]_��	���)��r�N��$\\(i{�c�!D��
`H �-!C�}���vݟ]�.4`!�^���w�g����1��0v�����f��Ƚ�e@>vZ�/��i�b�ar�|�'�c��Vg�H�-�f�RH��܋-����U�y�HͅY�\|�����q=�~u{Fb���D��U��=�EV�>{�P p;s"�Jr�C?�m���&R�M%_c���F�y�GYyOUG�J�ku�f4l/t=i���:Hސ���<�l�T1��Q�\BW��gp�ʘ+��X/��	�h2��f��B}0%c�t|p�7G���v�'�i��E�"u�[vI��WCE�֟��{运e�MxG��,��i;p�)|�«��x��d�|��:�{�"gsx��/����oWZk�(K���^uW/�W�YĿ2���C*>t=�iƭ �$x��	���l��i_�y�JSb�{��"���5y]I޴�F��c�_�qQ/t��!��z!�F��X�D�)
-BR�eHY$-򑎱9�in��Y�Y�~rf׌@��q\��4��_�S��#���,���܄�)֡Y�g��B�;��R�_�F���TF�|���FvEeD��c~65!��4N%o�.�y"�w�N��δ@�V�Q��Ĩ���n;#�?��:�KX��
��v�\�4:���� �*exa,@�Ůa��4H#�"���-�iľ�������-Z�YpA2�)�>b�S���q�Q��~����e]M��Ns�I������&����=Q���sg6���ax>&��L�7�R��;~�^�qj�mF����]+X����t�$�8v~��o������F)7+Oݴ��g�]4����цՁymi�g���-fa�����c��+ Vl��M8�JW��)�O}#䤳�����U������4f��!<��Q�撿��PG��F��$q|��P���uJ=����	m���^��`S<�����g��=��ѡ��/�b�X����xe��'��n6��.��Y�a$�������JR+(�u��es��Okx,_�@+�tt� X~F���h�,Zh���w-F�e(;	�B �_�[F��9#RpW�9��fH���d3� o�OHё>���	�c��Ӊ	O���lOJ��59�oU�{8�_������ɠ���j�1�>>�-R߹���8�M�����Q��޺�o=sf��AxF�qB�$�a�-�w�A��I�Dt�����2�����d&4_��S��s��ôY�/�5������u��, �U��� o�?i������yh�X��eO�[���¬\3N*<���� �x��Zg�^�G�b����Y��-���+-��Б���i���(/���kT���C\T�3za99��c�,�����;�QU>�j�!d���bKW�Ri�8n��kahih~���*��̺
�*������Ig�V�M9�z�Y�Wכ�!";Ky��s�֌E�l��Zg��;�@8H�^U?����j�uM�^8<'1S�ͭ)@�9`�@L#C���Fn��eP�LZ�j�v2�Hk�N
�-�A��9��C֭�{���j#$z.홰���ctk����t�^SG�ŵb��,�e�+	A:m���F�ċ�_��S�S�F���M'Ys��Z��T��]��8ɒ;�D�x�/��xI����:i�o���n?Ц�&�I:t����	�F[vY�̟.J?���=���\th���9�o��,Ғ��?�Ο&5G��XMtft�O;7�u�Yx�� eP}/-�X���v��w��ؗN:V
gj��*y%[i���7�{�&ɘ��qC�s�aO	N�\�(��/�j��a���%�=�!�QU��t)v��J��}�ouq��E �2�|���*��Q2S��:i~��T�~Z�}����hw����'ܛ�5UҊՑ�˘H~Õ�WL&���ݏ�ST�o��^;�A1��7E��w��"�����E��s_~_;1$�\��� 7�Ex�q��S4`�F-6UP�l����2�%���в�����p��{�@c� �?=E��JՍ���q���\�U�L_}�B������aL��E Y~S�( }�3>�����z`��?VL������&�\dV�C"v�*6�g@XZD��6)v+d
��+�����,0���)� NSG2��3z�c�ip�����Z:mZ � z���D~,�)��Ph�C"�
@ia�e&j�tg�_��&��\o��D��K#�f� �?�{]�2�krE�`fDg*�E�m_���7`2�"e��3oH�w��p��HH�L\;웞D<X��&}�ܹf�ף<� ����of�c+L�j�R����S![c����J���5�fHw�����������gԨ��!�� �3���C��2��Ox�]8�01>��`���c����_({��XBĢӋ'�wPʊ�7��~Ww��_|~ ʆs�v@6��T�]�?��4��M0�_�9����G�(����*�T���b�c?�K�<�K���	��r�j�D�W�'\�<����Y�� ���NC�ݣ���L�t������Lt`�q��	��ͳǸ�k'$k�8G�hTȤ�^��R*Au�u�1��Y�`��佲�)w�6�k�X��ϩ�'���G @B��:�C���\A�+�)7��l�NF&��z�q/Y��P5dn��g'(X7K�uV Y����7wE���uA�[}c/��MT�h+�Y��l�=x��Ӫy����9(G͕���/?�Xf��f/F��c�ޑ
�4Y��,7�t��:;N�Ж~j���K�����[g�b����y'��KN�Y�Vfi����^����Ée���%�E��8|.�&���ʞ|(��E*��(�S��`Q�jp�w��x�	ܘ��I�����Ŗu8�s��UU�s�$�[��B��jr�l:��gL�G��,Ov��*G/[���_�#e�F����f�Q����!������ak����$����TuU��7�M��2�a 8>�F���~�nG���a>�ȧM�0�o[�e.5rＫx˘�,f%?,U'���ҷ�`��Xx�NM-�g�t+�d3{	M��u`WT,��n���Ix��A'�9���=s4���՚7��4K�Ff��g���؞�X�{����XPk-BZ���������R�9&�����r�9�f������1b�Q����q]u(�h7�(��T�,��u[�8���&�	�G[Uɏ�����"����r��Ɔ!����Db��]�Y+�������Ɩ�B�#5�nE� ��\-�C��W�^��j�8��I��o�%�1q��lѫB�U-�7$ȁLB��/E��gn6\Wˏ�����K��o�4�<�M^��~"T�t��g����s �Gnˀq��Qμ�����^v�&������M�7'L�%�1��:���@n�`�ŝ�+�Ұ�ڙ7c����7��]`ҮN����9���҈�m��g��GnR�y���H�Ѧ��w�4�_����=��`����c$(Qy�d���D�5<pGF�&'��Ʃ���!� =�V��o6+�}��艤�\֕Ҫl/�)���<B$.�G���k�/��zu�'��f]J�H�p�,��1�-�1�.��<yrws��,(�",2�+阬쥙�a.P���=�t����X)�����g�ݾ�ꧦ 4�	!��{l7�0����REZ�)��bAI4>����Slrsu�J�M�_�%J�t��w�a:J��,��w�ey�FU�����?��i� �S�4�������b�V��x(�Y^�։�\h��t	����.@���\�pFn�^���1�\�b��#���%2{=�5�Oၦ��.M��F�����rЭ�G{�K5��-�z�fE��=4�>��<� 3�_{N�(6;%�'6ݟ:�ɣ��<7�r��(�PJF�CG5Z+�JD���E�~�jW�w@�a&�K�����z��2���������]� F++�jw��Z`��}	��Cqd[w��lM�r���^��Âk�&n ���`z���F'f������Q�YO�P�HO�$��Uxst�7��[ek�K�p���C(j��'_,V�%����2����+�9�@!7x�lz�X4� N�챌�Jzj��`(@�p�-����:#N[e/�IG�W�^�2�=�{W ��!ĚLj�1uTqi;>a~��Y�؋�8�g~�\\�\F�q� N)���V�v ��n�=h�����t��d���tr:��AP����@�t|��{O�x~H�3�Νɿ��f희ĳ���<�H^Ope��:��L�8>q\#���8*���eST�I��N3�Q�\	��L�@�L�� =Z oo�ή�A��a1�2�	|�J�������G�-� �]	4*`i1�T��K����Qj�ݣI�~������c���]�6T>1x*�ʚ���c�F&���}8�w��K��.?��P'� ��-qs�x�R՝�ޥZi�M[r��npL%�F�hGM��.����z���W͵*��h1��	[���_d7s`����"�V��"�Geo{6ޚ����r��9"���U/!�Ǵ�L�qu�5��|�<K򴬣��05V��Du�bNKJ�5襹��M/�J7���{�����v�ȥ�qYxؚ�f"#��V�4���L2����1s���"do�o	{J�OT&�^3�ʔ�\�V$�W�<�l �E��h�N��1�\��l`�F���Xr��x���&s%��K+�s�ԣ�|C��d����]?e��Q{���Y4����s"��odg��Cmt���͓X�l[F%b[rx�@���A��V�@'�(Z���~����EA�G`+��j�P�bLl6�-�ʦ�n	�;�;'$��Gp"��/s�� ��5�V-�z��3J��<�jM��8��w�����q���jNz"���/4���S��/i3���Qs|�,	4��	��}�I �36��O_������o� ��Mt)��.Dn4��G'�|��I�ڜF��eߕ���_�g��H���"����f5P5�7I
�s@ڊ��ۑ�J��Ɖqkh�]pUG����Bb�$/�<����:�,�vg�n�c�S�LX��?���я&]��K��ߌ6�X�j��w}��mvίV/�j�ʾ��[u�h��f���ς��X�9'�-���F�dw��q!p��MO���\�j���
�lZ�c���]�5��_|����=[�����>�gh�0���*�~KP�ߦ����S�cHjg� �I�ue�(]F�ni�P�n/>4��z��&�����>�3Q���ؾ3B�����)G�+d7�d��8aFy
�+$�vcE�x@�7��Vg���]yq(�wb�����&���s��on���}�!K#xh�G��F7���r�~��Ԉ�� %���dw.*�JຫA�ߏ�ͽ\�u�h�5��5чV�F�R�L���S̑Ak����o�� ��M�O�mV��2k?d���Cr�Od_w"����]�:±�$�k<i
	f4�簾V�b'q8F"܄���ꋿ�����Ne4�N�G�(��ˎQ�X&'G�q��m�4~K����9�+	�2�x�%���ThK�kB���p�1w(hV�e��f;���eX$�s�Vu����z8��hC��fЦ�A��L	�?s�벰�ܽt��B�v���1�fS�U<u�P�q �fR���\�=
*��Cs��P�����=�>�b�����C����{����Нi[�Y& Ԅ�cQ���L������R%�R���Lͺm&�l\x�Mg�J�$ޅ��НB�W+/h=@)�>X�W^��}��9��@K��T�f��ӫ�'���l��%g����@�����j��m�0ò���WÛ����"�tZR
yz1��}��5�y�\t�I��m(rť<�i�RO��aP��:#�ǎ-4�����{���;`,5���ι�v�1�Ӵo�<r؇ M�<WT�O��z������)	H�">�F�4��
��iq��D4��0q<��<��AtQ�s����<K��l��m@��rl�`D�u��x�{������y�^z&�uQ�#74�&DVɩ*\�	O����ae]�5��,Ή��O�x�C\����9+g��,��O�e���xh�;���'�E��ʬ�@��/�bD�-�%\N'��?�n����0|x��������0�Mϔ LcU �Ŀ|.RLC
j��u�B]������=r���.8D����ӞM�g+�E�j_�[	 �[�X�n����Y��0��V>�P���,��@/2k�f�#	�8���ts��^����O�zɻ�~�gLI�Fl(�o�U�A`�z��GGK�.Z�=��e��w�@��I�6�p��Oz��:dE����������G�qs'�_8o��(9���,?�m��PQ<�}c�ӷ�{!,�h��)b����F0����%��N�b2Y���.�UHZޣ���H~�i9�lA���4���G��y�6f�C�7�M��d���2'�c��Kuϔ�mW��#�ԙg㴭�K��vҧ��^"�p����Nt��c��o��n��F}/o�� e�U���Zl��82+�#:�����]<���O������XêkFZD щw�>g�c�������q+� ��>����8�*��jI��el��g��l,yW��\��k��s�䄖ǔ�"H^r鿓&X���S8�{�w�o)�A���힭:7�}����l^Ym�uY*3��*��L���9�<�a���b���7��b�6X�W��[ȧ�T]�q���F�<�d�B
pS�z=gT��Bwc�H�?	H��&�H+���fp����A+pQ'w۶�p���I�ׅbEE��C"����2�sv���rɲ�}��F�S�.W�~�ҳ���r.Ѝ�R�|�󖳲��дO���}�Y��B��������:���p�b�b�&Ku֭U@U�t>�ʞT)��C6/��k��T�����:VrW.�J��f��ݕn#����Ii��T����I��'��U��۰�g����?4�;�}��I�Ac������~����O��@�/�'+ez"�"B
�QpU�"Ч&��?�@懢��CO�Hr$��V��vj��g���1U�w�cC|UtÅ���ω�;�
���d�X����E����G��8L,�̹��<~Q�A�/���+R�8�B�#m���7���ZxC��D��O���a���S����GR�0P�`��&�s5��t�t䏺�$kr�	sK�@|�=���@��Q+���oq���'�@�C����a���c1κ�P��,��W��M���ٻ�!�8��F�	����[=]#=>�V��4����f��-j�A�mR���i�n��xܯ�$p�����d�Ky�����?��@�5]�1`�����+���b&��Ed��/�>$��Q�Lv������Sއ02��2*�2�5�8��n��} �2)�O-pG�_��AH�H7�W�[�\`v����ű���8�@g�v�YҰ�`�"��`�e�앁c���b�����j|t��&���s}�������'��y�a��ZwO���C�tx��3*!J�M=��A"�D�P2+_��pf;X�c
�Ŋ���o�'�ychoZ�	ȗ�=z�ӕ�Н~�@�_�do�+Bkm4�|�>��sN�����+
>K�&��u��@���Τ�İ�Z�;D��
���	�;cJ�{m��tP�}	���#\��W���(��*Z�K(H��~^������L�4:h�x�k�<jpVA�0���c��>ݘ��"��d����'#��$�]}'����O?��i&�~@l�������D�Ɣ	E7nη\������m�G�O��ݫ�ZNC���z"���1��=��kU�5�N��	2��tua��K#s�&R�R�e;KI��%�M���ߣ��Y��~�{���z�#֠2�k�;�}���!w��[KH���b�Kf�U}?�V=��G��ƌ�I��B�"]mE�p��<C~~�3m�!��o^�7GM�%��^�Btm���.�+߷�٩%�(��z�F��`�{��k4����q��	�ݎ��n��o��[.X
�)���9ҋ��Ԡ��Y�8�u�<a�;�!��C8�(����D.�XU5��BD�p?�f�2��?k��*�3d?b)J��r�d릝Հ��70��c[�P�LQK��E��p4ec	T��V�P0��3b��r	l~���G	C��𥯮b�>��DSFH�����U�o>��6�o#�UT��e�"3��i3�0P�j�Hc@1��X�9̀���
�+�3� ��?�`����i����!A��Xay}ׅ�Lʿc�w�/�a�|Cѧgv9:�٭��C
�Y��T�$h�gAtk$k��c���Ŗ#���o�����|^���P���D@��aN���s�~@|�d2��s���憵��������"�6�Tx���"��2Ch�q�8��$��OQuO(�^��8�K�ښy&G� y�v0%�ElW՟�����6�M�
��^�ܭ-S� �r��N�G��K��L.���Q���I�)��?S�I���/_<�bj���-��4� ���K�Oua��R����{M���0C��W�⚬{u=ݶ�}�u�)�@&�`)��]�4j�$�HF�(AxȔ;oQQp'�Q/j��O���;`�+#j�I�fpAy���%���4B*��؟���h�������f3�b66�;y\�'�V��;(�B�-Fq��xI3r;��P��ɏ`��� p��ƈ�\�AO���)p��m[��������N�ؕ� ���,S�T����=������lv_�|�;�2_�{Ȁ��`^���e
Bo��~>�o����)�-ʋ�����agt��7�Z"� �L����Y[ �UB ������Ts��=����'�ُ�<�m,�E\5u����G�[��]Q��`���M ny�������N�)0����	��Yh�
�E��3"���
���=�j��ˀ��`�"�����ZB��j���T��;.'�'�D˖��Q�v���[\�s��;5זȿ�(A�e����w>�^�rP��47I���'))��[��!R&��@�G�2]�"��gW�eŋ���f� 5?$�u�� �y��T�=T`_ѿ��z��`��1��1�q	�
�>��x(��ö���pвqm%mKc�W�_��#^v����,����d.2��W���U�,<
��
��>��\�:�7������'��&��Q�RN���o��$�x����C�3���+�"U��xgR*����0�� K��Ās�;sUm�.R��b́#s^����d���m���ςĬ&��W(�Ę�/1x�jz��,&���_���~J�'r~;6��%�A�[�<��Y��ë�b���	�"���A�3��%�☽x�qӥ���Z�~O*�v�fz�ywY]��S�����%C4Jk�d��� ���%ޱsğ����!����@¨�|y(m�M�?@ִ���	���d��w�J�W��EN�R��fڅ+l�|L��d	�d1B6�L��=`]Ll���3<��ar�j|x�$�mq���CYO�޴'� ��rF�.J�뚧�qMp'u�=`���A0,�T���j���L��0.�E����9���gM^��[c)S�������|8���fDjKcF�P	��E�E��,�W]��L�
/ѵ�п� ,�7p�+i��w�v�E/�P��m���v�ź���ŋ���OБt$~o��]���y�<O��8B,Zx
�=cP�t��3�J�v�P�`x�G�X�xr�7[��t���=4���r.A�Gvh�Bkŷ�B���e�[|�yp�R����ѵ�S�=�'<65��/AV �,2H���AS�y<Ï��1Y��i$�}�F���Z���"����fο��R�y�F�(a�G�ުbHu�����F6�Z��&�5�����$�����Kv2��4����w���lK[r-H�o�T#�$T��B]�\A�?+Q�4�&GF����v8s�3'�ޣ>b�ǉ2z��xq�����h3hK�@�STG[�5xIe�
�m�@LV��B�EU$R_����ߤ�N�*�X��F�m�'����/+?q5bjϢ:�O�x��V���6��m%\�Z��wGǝ�3%NL�x���ަvE ��A6��=+2t��6�ز-2-V4���L)����#n�aVsn׫���T�L����L��&��2;:[��
��vD.�Q���`�낰c'�Y��>M/��N����
��-J�"J�.m��r؇ �R�8m_����	���_C[(3u�,�c6�6���RA͝����ż�f5���)��e[ �TW� �Ҏ��|D<\n�!nI��Emg0�F�щ+K]��_%V,�h?+�'���Q�
�mV��&˷�'�xiE�=��n��6�n��I!�UUK��A�$��dX���-���_�l�g�3(M
�����;sx�
��M>�~O�Ү��߻�]hs"պ=�L��C	&��-��E�����cp�v�p_>:R����ɴTl�<��'fv���Gi���fN1Q!�^�!E����q3X�v��*�K����&iS�<�	��m���8qn��[ȚΣ?��<JĞ�T�tH��.�ل(@>>̃r8��K
"��"�hq=����v�����P��v�V��#0M0�*�C�.r��H��q�jyV�.� 8u)ZX������u(�]�Jl���uz�C1CntC@�vnJ*�Jgt�]��x���Ҹ&�HvG��)��~k�XFH����'��V^H���۝�eA�e�CY���]��ܛa����R���$g�fwo�w�s
��n���W�G��%,�O�������~n<�k���	�r���������l	��y�o�g~4�8���U���t��Y��n�L�᐀���]�a��^H"}}V�Gay�Q��$�i�w~�զ����U-?�k��j�׌vN�9 FX?j�|t�0������uC?�cSٵ�
e��U�h�j�R`�x]��Y���,@����;
m(D'����\Eq��=$tO
xS�0[�:�SU��b^��=��k�S�!�D�MR��4� 0Ur��VTTX��{g;�@QeG2������@=�4�]^�z��?�"���]P�i���9#�2]�hW_��3��;`����=���j�A[���Zt�~���F-0�2�[�A�C��7�D�Y�n��^��e��J1_q�솸0	�I�_�]����U[J���ߦ!���샇*[/%���O�x���W���g�8�^7�� '|q����F��e���<�e��s�����')��Ȝ,�T��rޣ�z�E���_XbE�6tP>�+��R�p����Y�%�������r�F��F&�k����1B�����X����A����1L&�������1�Rp����׼W[Ƌ+1cs��PV`�4�����բD:���)q��PYg��/�俗�De�ד|��z53]N�ĭ,`jQ��A��H�{�W0��T����l\�Q��*�x;Aͩ�m*ZPHCF��t�4�Ë噮��Y����d.��j�'j�I��]
wC���aڪ:|c�y��`y(/@H'ڹ�Q��6K��0���	���'���9��~��4��i�����U�����~����koϋ�X��d
.R��^���j��$�X�kx�zTh$��W��j��&_L�x6�
M��RB95@Qpv�y�]��?_�F�S9t�<�w�����5���iu�R��UxE�[0�-��P�A���3��dn4�a��1��Y]���1���x��`z�LF���'0���Z��3�2K������ �G����˴L�f��v=��X�J�Nnƫ�ަ|ڏ�(e��L�as <x�T%��彼ߤ6���j�0��,����B�-�C��Ԟ��u�$��ʒ>�ܵYU�֗�\��`Ȋ8��Kڷ��q|U_!�P�N�nO��*0\Y��I�Jt';�@��+�4ݡ�N:6��݈GW�į��ģ�����&��k?�
�]���W�`���(iY���,���z�)]B;�"o��g���(L�Q���a���y�01KV�e�[�C����A�3o9�!OE�����)<ur�,!DUa$��	E�m�kQ'�L�Ň�n�o(����b�E��B���&��D���܌�h|�uE{�V@�0ǻ�/|�=&��R��ƝA��o*W<g��< ��QOZ��M��i\�t�sQx�P�J�р����egpl��KHj���=_�xg!��-�^�~��I�6�9�K���$��m�H�,�/'l�lۺSj,��'��ݐe�D�6 �'|.���0��׉ᦠ�̀��.Ks.Ώ��.=��N��ȉ�-�$-��BKꍌn��:\�d�+��{��*��Ou���Q%�����iv�U�ĺi��$��Dt�*�*�l��h#ː���|�!�h��:����M����؁���h�V^�g��v�&Y����[���M�������k�Ms8L7v~�p��xC�!�ާ�\�c�p��vK#C�s' �O: "s����7ߌ9��2�Ӛ� x�p��B&�d���kD�aQ��v�8$";�Čsg+���.m�|��
i�5<�Z�*@�O���DY���֛+a���1���8���vnA(�_:��ԯT,��7��j���%E�߽�
aǾZ2�=W7fO�`$���KP���������K���wj�b��tgC?\1N�(B��}��B2ig��6�;Ri(Y=(�ԍ�N|<��������V�J�,�	���Z�����*�?ߥ�*�?w���K��D)����}	�Z��鍿�c���b��G \��^~×��k��0D��2�|h�r#Űz䙜�O���E�Z�����5� m\��&b���MY��}�Ɏ�i�x*���]/�׸��S�w����{o�ƨ��ؐ�M#�ͷ�*Y�v�雖�����8��{3��}����Pg�w��u�ֆ[�k�h�cPw�ă��PyqD\��$C��3�S}��=�Q|ʗI4Ks.i�\֡�I��e�-��t�����W��5N.�`!W���q2��.�Rip�^�v��m(�F"�|�V�	:��W��傻qn��V����e��?�7����y]c���O���[�#�Gm��Gp�֠NEk����{���촯�ȟz6F�j\��AoX��i�T(n+�״��l\��.@x�T�Q�I�-���x��%��{U��[����kv|dZ2e6HC	�m$�@A^S^��@����+�^B	�Qhi����z���=zq����=x�o�����K��'aM��`��tW���-�/J���
�w��R��A�r�Cކ\�9�TX�����`�}�X���_G�H'R��Vr��
�Pa��`!�ex*�;�I���9�5���QM���p^��$M]��@**]��U�>+X7�����F�>���&/k�+���tл��n�����\���t4q�kQۯ�����-��e�&���h��D{���d�j��L�H�+g�Ѹ���ѻ ڱ'��`���G�%(��O�?�a���Q�k��w�dUj^Nr��NVܖ6��)�|+k�-�#�w�e2��VB'����If�����5q���-	�P��P<�&"�0�r����<�� %�Lӓ�.��(��L��N#U��A�E6����e]X�AP���O����K.i��)^��h<� %L[*���miz�Q��r؀@�L�pcz���t���G�0Z�����`���dI���Bu�����eth���%�1������6N��I&?)��\�xӪZ�������P+�I�F4D��i���e�<Gc��e�(�_�S=�U y�@d����a�x�W[uUY�[%��so��� o�+�Tk�)L>4oId_ǵC��5036���u�I/����=��OČ<�f�lwpVQ3�̂Uki�k�`a� ��}4��z�CX��ؖ�� |���5\�����@yIX��IT����WRֹ������;u����6֠�z\��"2��}�{��<�I��R�?1ue���,��:��9��@s�[a����S�:�u�=�I&_tF��]&
Y-�s�8��L�\�Wmt�V�3�&>�����xS\I��r$�8�#E�7�K��V	Ɯ앳ʎm���"7�ҬL!*M`� �Lcd|;ĭ��<+�!�G���.$0��4���I�X��{G��8��ar��"a0�$(���<K�h�ֹ���:]j���I�n	��LKt;*�Ħ�Y��c���[�"zNc�;ˈi�|�R%&�{f}�15Ժ�Qm5F;�h?�uS�Wk�j�^�1r�&%��R[YE���t�@�^�o�Q9�@�g�`"��gS�C'�7����QrS���{��.����xc��Ci�������S
���t�-�2(E]	{�j����r�-��&m-�@u��XptB��>)U/��Zr�L5+{��M$��9������f�����\��imr��q�Y{aQ��J��32;�~�`���w��u��w4���M�g���5݀S��sO��3�n��Ѣ��>y�߼!T����W6�h��Ik�>�!��[�k�L-����!x�XNn?ÌZY~̖����9eb��Y6lj%GO��!&�et�Q�����c?AW`!@�	�	�h���*�o���W>gnʻ(�V&C�;)��w�~��%zμJmy�1��j���w��F�f��e��	c*��;�=��Fհ��%.���Tn����ģ��/�GA���\�{�SN1���d4a'��L�����i�x�o*���t�BC��Xa�������:+(p���e�o9��Ť�R��]ig*ȸ9��i'�`l�G[�%~[-��L�$g��. S������`d����{�����F���i�S̺d0��K0�u��~	�R6���n$p��3R�����t��GE���\7{���5����XK�0������6�'�@Xԅҝ Xa�(	�P��N�]_�� و�󥱣Y�x��f-�Ժ�_��(]���~4�vUV��d���� ��iA7�s��ɮ����^Y�#��`�I7Fu;�.r8�9y��ތ%���M������ ���P��^���S0��"t���1�k��(���v�kU�EG���(]�ZV�@g�W�֒�!wm��/#�a�G�R��&�`]m�)ˬ�`²x3��_�2o���*��- ;j+�Y�C����/��W�#�*����W��QA3P"z�(���-��po�>�T���N���g<�l�������ƺ&¬�=S����T���ؿ��[U
Bk+c������T��R�޴T-a=��������_��;�	�O��	�;h���7��Mn��8�3!kԳ�� @�V�=�񁰋Ra�9�o�+&��1�jw��vP�ds�2�u�Eh�
јsq�۫ܶ�vY����%��{�C���y�#y�\�E��ʕk&��ʿ	m�*�fZVٵi��c3ww/P˭|�|�|Q���ο�p�����{�����i�Դ�j��i��&��P�͛�m��Ѽ�����Q:~�U��y�~-���:��J���Ös]8{�W*�?~�%���B/�C��/_D�����p��|�F�=��[Ó�����D� _��ji�a0ģ:��9���N����æ��7�n/��	�4 ��85�A2T!z��]ލƘ|]��3�p�����cK���6�]��)��F@�,������jc1�D �,v��+�=AL��
~�I�I�6{�@��w�<F6%�g+C�$zɏ�w�`�'���?h��G����*�7�R%���$�
>�_28�*Fj�ݶ����R㺼3��H�գ�?�B�BxC��� �>_��h�ߝ������T����o~�k6�W�u�ÕQ����8�?�K�����|n�#Y�W�hs�	`�3���J�
8�{�w&�Ƣ��_�P���k�/�OJi���w�[YN���d_�.��>���P������qE�LLy���p�x�H*dy�9 ���dq�L%ui�hCWc���X�@��0��*3N�bP�~�� ��tc�dOZ�<P����XXMӶ��Mޗ7�8��D�a_�8�`�v��RE��{�&�\�Nz�Sc��V�޽ʮ6��`���ؿ0�Ul=���b륍���;X����A�X7�D�Z�NGɔ����Q�i��B���a� �\��*d7�n��!��D?"E5;���E�#[9�2eq�Z��^�	`���VF�S)�4�M�[�\��&pW�N��dT�H�5Y/^���g�4s�Tqs&# �Y�s�5O&�쳾�p C���Xa�6�ʞ	vRF��4P�Xl*�O5b���y-2�JRs/�����~}
̜��R�����#�6q�s���S�wxxO�`d��UҀ�<�~�����L�.�G���za��1p�����\<3Y���ů��vd�Ѣ쾤��Azs���x������O��;E������>��X�%�� �&yA5i�p}[�vQJEr{�|xp�V��3�B �r+)xI=4`�%Ȗ�Z�&u�*�ǣ2䈈�|J��5}>�>��e`->��$kŚ���"�Ap��?_��X�����z�dM�g���;9�h"�v��6�,��ҿ}Jq-7Wݸ;��tx��s��28�C�:�g�RtL���2@(Q���ְ6��.��:'��=t�o�k*oh��������t�m˧&�ݚW�G$#�0U���Gl���V����Hwӌ�C�����uʭ���3�9�lr��R WA1����U��r�Щ?�qg�H�T3+YI�<=�?�ǭ��l}H���i<�����{�O��q��2 8�C�g}ԑ|��HÉWB|����C��D�ʘ	��V-8p��(AeT(��u�)F�A��؟{y�R������)����Χ7P�΁U&MBW��<���'{u1w��x��
;z�8�y�XYe�*�C��2@׭�p'�~��%���|�J8�eS{|�6��fR��87�*٠���oW�
�A��P[ǤG������i��4S�'��e�8��B�$�}ڒH�$mI?(��̑����
��{k�ь�21A���&H��N�6=4?���>��L]8�����j0"[��:�� ���Ԥ\s�G{�D{M�:XV�$\�Mn�����J>s��m�0�:�flN���1~���-���Aq��k�^`�)AW����o��oÉ����ɓ��t�~;�/|��aTec���ٻ΢̴a��j,�M��l� �`Хb���ZV���O�i�/kЕ�)���+3�J�ȷ�p'�6Au�3ѥ�I�?���]�������<�_@�<]��y����j/��:�R�z��3a�);t�{���ohE��
ꂈ >��H.��Yh%#��6�!�q�%�V�������Hx�:Pm{iP�oC�`���n#D�%ݚ��?A�;"�g���=���aHh��Xn�h3��V�j��g|�����r'߱������}
'苗p%,TtH�x���#���p.·�8M
�ʃ����q���YҲ�Ӓ�\�ua�c9<Z�_r��qƻ���G�Pk����y6����U���h���MV$З�Z1��⁷�����@��J|�zSu8h5ELYb4�ȸā�1�� �����D9�H;q��	�zOs!��eHK⋠٘h,��Q���S�2�s?i�o�L�<^o��� 6f����t�>@����M�\�jZ<ʙ�k�6��
%gb����lNҐ�O�b�*�U93E�w���g����:���|�׷�mE��u�m`bb�;op?�F���7�野�Ġ��.�׫{Յ���&Q�0�|��� n����AP�w�ʅ�#އN%�@����o�4n|��9���xsw1�7v�p��W��: _i�A���| UY� Ԟ�x�D�Զ�E��:bˮ]��5���4׊��]�CN�M>��$����pg�I����f4$��u�^	?R�/�����1q��gw�G;�/�����X�`�.��7�&Ǣѭ�}�7��#q�9hubP�}/��=?0΄#����|�H���{���u�mQ}$Z;���=�`J��՛1���w��j�ap�Ko�19t��.(]�W�s���3���-�jx��������Ϙ����� s&�����&�ɇQԤ�>Ox�������O��d��h^�l������(�����SkLu��"��r�D�-zr�º�k"�� ��g�=�z~�8.@%[��e#A��a��7�;�-)����9	�X^v�NA��Y���������E;�����!�;�5��H�1����v��z0��%��S���ߦmv��le��M�ww���W�d'�<h�x��!�H�����xf�|HK����n*���$��m�J��n�:ĳ��S`�[s�B��*lz�=k��\��xq�#�IG��V?�ˤo,& p�d�3M������������׫~K�j ������Z̹���%P��`N%��dۗ��c�O{����uGe�]M�.�}/+�:�F�Q�'s_d\ChzN�״�$֒�8�'���b.���J��E��8;9ڿ���!1�M�=��P�'��D�>Flzl/�|% �/V��oz.Eԏ��K��������߆���3�w�]nwi�������:间9������˴p����w����"��34T���;:�^��$����B�����DFxr�~��

�L�E��G�����^�/'<�!Y'_щ�F��_MK3��p�l&�Z)�yG�x���n*K8�ͻ��3� G<��Wkw,ʛ��w�ŧ��6 R�4�/=�%��b���/K:sCC�)p��ܲw��opN���k�#t T>���GLo��~RY�;8�?8���2�i֟�[��(xf^#�bMA�4�Q�dH���k�ئ�Vj
�h����fN�|XHB�n�_O{�����ߡC�5z'bg �٧½��U��c��p)j,o��CJ��[]��vyROG�A���(��jR�N��ݞ��P��!�JW�f��G�z� �չ/Ra<1 Iǫՙ���ʰ� V�	�k+��Rr!ݵ�V*�NN��{O&v��n�p���G����� �Y5�˨D�U�YA�b�=�kT����.X�+%��p����0�����m�1x�K�� �Ҵ����o���)�,B�K*@<r�$�l>f��q`5��D5A>��S�\jiY�"�@}�����]��R�VѤ�� ��v	��Tj��1:�% �QE(�r��h�VuGǰy��R�,&\EZJ=� 2\�0'ZJPp)7%9Sѧd*'�3X S*�{כ� =EEq,h$�*��9 �TL�ʭd��'�@:���Tr�I_�c�s�p�ېV�6�ISx0A���B}'%P���f�gm�Z��^1T�^y��tB��Y��BA�����ņ����a��K-�O���|��3`�d��P�H��_���+e���J2�&c؃s�C�&�m�|��׽�yXCQzs��?5����G�a��f(�߈c�Ϡ�oې�k#�X��ˀ@����n�y�`^���6ـ��p�\a�1�j��e����r�OBͶ��m�[��f�gA�i<�:]N�h̅��-gD�0BTj/[}�V�#&F�+��~�����V� �g��zH�ń�K���!������C���2�u�s�%�ѽ���%�~}�����U�8���GUU�1ձ�%_H c��F}���k�ʴ4����-a�$�y�p��1���80�8'��'�T���1P�����L���`q����$���?�^L�ճ��:��s����.Q��� ��֘��'�;��1�G�$��{p���_��	�<�X����d�	�*į���mM�z���'�R�u&�(��o�e2����t%,�̜[,���Q	����y��N ;?�q�e�TiQ���NHK��-��ZW 5&�d��ôKƛ�,O)�31��ƅ�~V`����X�]%�}�׽"�5����b�o�r�4S�c4�D2�WU�yͧ�X�ëv=:�:2Uȓ��fnW�c���k;a���%�f�82<�� D����G3!N�${+r�9�#�ؕ�Y9Jq.�Mʬ/�^�s*(_�n�m�M�~g�(G?��z�]�z�ƀUxY��&.kOop���ζư#>�.Ȥ�Y�}��v�-���v���\��,������	L�L%h?��򩀸s��]�G�Nx4TC'�h�us�_�Jl�B�ʠ���H[=TO�&��}��hb�*��U.����PGGw�5^��5HE�M��dR�],Kl�;T�c�X�,Z����$�m����]���U�S.�l��e��G�~q"_��t�k�ay��[��J���f�0b<H/�s����t~��0Pԁ����qƹ�hi����\E����]�;b��Qߞ��uV� )��)_j��.�L��j(�b��#����,!�ZW���̮8�gQ�;+�c>Ih�Ct/F�ϋⲄm�/�M֋�ҋ)Is=3gUř�^ǚ%Н��zlR���& !h�Y\�#���Ǚ��	�Tb�T�$G3@��1�����EWW�#)��p֓��H�C����O�u�@��:�`��w+ߗ�(P��$�'u~�ۈ��!��M�&6/�9�:q��O����[w�����$�zQ�%�)�s $;�o�V�����&�g����Q�(�e���*��㇎0�f#�<S� ΈC +��i�������A�ց��5ƚ���ELK�9��"R�7�H�N��q��p�f�>��)>!��~��UP:�	]9¨�e}�&����S�L�MEB�����L5�ǁ��ɮ��D�^u#�������5� ��h/(?�hv�0����`���Y�ں.���Q����.}v9�:��]x���=W���D}��CT��ώH�2q�1���G橐��a�ZJk�C�?���:��%�]L�OC²I%�TN2@���h[������͒�Bǈ�1����i<z^7a[>|����;��2m���K�V���]\��P����Kt�a��/S�)Ԩ���A���I���Vw��o)Q���� �ԕ��	+W��O��;K|KU4��a��9�3`Q�l�ANR섈��h��	��>���4��n���x�5h�>�<w?`H|E�k�^C�)J��U;'�輴:eR�=�����wt@\�D�	�u7Ğ�j�2�gz�XbFW����`~Hs�r��7�i��՝�n�S��V�%�&�Rg
�F�{���D�W�߼^c��48��
,[W���_�e��W���1tD���<N��}b2*��v]��r2*? �S�I��ʺ��k1Z1��f����N�Y'|����N��T�pF'끔�q�l���5�O�$��R���Kh��ηe^��(����JC��l���WnKiީJh�����Q%lsls��զH�ʌ���g�-��@I�j~ĳ�A-.x l>���G��Âf�8oq8c��ק��J�2�F��ս�5V��vFM��[斶E��F��n-�z��Ʈ����*EY�)1^J��+� n�#��t%�8�Nv:����	�tÀb�!������W��l9�C�9P$�N�������{!J��PO�z<@r���{�v��'m}�a�3K�rM_������I��$Ű`yTE���N<����Aw��7"�'NjV����Qf�WL~(�n����2�u�r,C������eR��s/;X3@��e�5X��n�%��-V��y�@၎d�K5�Ǆ.,�Ln�WJ�� /��y�V���Va�5���~� 4�.������� ����\�kO'�F��)���!���
�A�������Pp�
�t<��x�{���߷�����_;q�阾FK���{9}�������Q�N|%q׾�ʌo��·��E���Ǟ��c�Z�Zëp3u� w���0%9��R���%�0���������i�����ޭ��x��Po�������M�<w��ٍў`X9 �_O��-������DB���V��b=Т��JݩA��������ƒU��RJ1=�����]D\ej�#�T&�ǳ��S�:"=@��ku-P�IR��)�E�$?�S��6�E�@������蹘�7��븤�H�<p<e�غϸh��v_��S�5�{S`�N��_Τ�
��f&���Ʃ�=�����(�xTSA�����))z]һi�~�@n��,��l�c��lO}�$F�?�p#��Jc<?���=��f���mn4Xeޞ�VͿ�6h����u'��]z`n�@�̾S1F�2��Q��yh!�Jsx��lͩ�O�ǘ�勊f=h������LX{���؞�G�� @�S|�TN���n!��S��ݮ�U����R,�½����,��ض��:]���H�Xj��5�9LTQFt%��k�B�|j���.e@l�|su<���D?��0';G������%ɂ�lYvn�V�{����#@�=� �.�����%�S�#k'ˇ)M�3d�{u8U����NC�����m<���q�E���R���0�
�77�[AͶ=v��/7����v�&�%b���_���YI�E���D�Xd�B�}�g>��k1��@!vj�h�*X�:�c�?JO��d�Ř3�2��2%^� YvS����⇏��3�&��L)�m����6þ�ґ�@��Jw�7}ꌯ�\N�b| ��Tg��fz��k�
#�-�<� Q�2aK]o3vu*s��Ot~�#���/��Pcf��P&� �v�lŹ.d��b���̓L���Ĕ>32TP]BW��mw�Q>O��I�~��B@��1��T�"^A؁s��^p!'E��|쒗׏~|��ݎ���@�8�ڌ�>~�"�$Jv�L#��>�j������w�#,/M�u����M���e��k_��������S!��4 -�a7������C�tl� ��_�ta���n�+5�ĉ�SU���/��	њ7L��2���k��3w��C�Z��G�h�Y�h4�-��F�c������i/,���p�ڥ���#�г$�ܜ�hL\������[8N1�z�$�g%����}��)6�пq&�-���Vg��d+�LzCd]�Fw�:��0C�.�(�M�h�U���aZa櫉��
j��c;� �Ȥ@�Rh:�pB�&i���3���+$mT���sT*+ڧQ���Ѡ�i��qO~MO�bN�fфU<����7��M�Z�iU�zse��̓/_�[�AYc�p���(a֓��{�ԙS�+�.��� �h���&��gk=c�R+'_�a�.}��f���e�tL�Ϳ��d�W��ی����;i8��~@R?�ǐ�<��3D`#�
��?�2��2��-��G��w����*Ntz>��1�5�P������e��R=VJ0�#K�}�g��c�[ݸX!��:q����me��w���P������:k.�������@���Ղ���Z�)K�kʕ���<5u4>���� �zA_y�[[1�N��u2!Ec�&lh�*�xIF��2��27�݄�:/�9�t�K�'͏�gf�N��Ru-E�9�u�
F�!�����	�Y���c��|?}����H��0&����)a*���ݓ���dt�
�=��ѝ��C������/�5^2���(s�8��)R0rp �פ�|�jf�Xfn��</��ێ���wzy����2�~�J�o����L��3r[H�����w��mu}]ݦ��$:L.�7ak�z��$GD �z�r!Ѹ]��:�0q��ݙ׾3��U}�Z
�Wu1d��3M���8����'�9\�<���*M��ݫ��2�5��H=e�w�)�(8��5�nu��SU90^�$'yMp�T���+��~cw��Qo�P+�pP�t�6����;^Y
ۗ�s��#Q��<�����uD'f:iz���M��5]NRm?��v����UwU���Q��z���T�>='fGh��5y��ӛ�~U��F<��g_"������v}JA�iF�v�g��M4�������f��y�M���c�q3=�xc�,N6|�u>�Cю�4��h��h��I?Zz������;/�g��%�n�˽�ZÐ��w�)."��mݠz�v�?6N�E�ic�P��L�?윅�2i�D�2�>�w�Jْ@ʱ+>Q�B�t�Dliu��E�TE\�r՝��<c�ϒ`�:U��¹yx�FPs��l�N�����6���]�Ns�u� �?"K�����w�$���a��;��I��?��h52H/KrAz��W����o�4\ ���=���{���C�\^ګU�e�e��o�5�Y?���{\���>0�D<�o��<�� �yTvK�}��x�e�6�?9escE���f��s���ӌ�2��0�����j2�CO�t����^������Mh�ǪeXv���u`�	���>+ݕ��ۑ5v�0s�;zes���� ���P11|�Z����wr�/�扆!��P�*�/�'{�=���^B�/'����&]�uv�<����G��J��2��:��ެ��}%��I���ݘ
�M>֧�l����Y�/G�c���Jo����������G�@�\"�׊���ߍ��P(-�+Y�`v��*[:�A�wt�Q�ݜ�+��~���q��`l�N|5�D h> �Z
�j�UB��%�o��2j�f F��e5ܢy�%·8Fg�)/���MG]<g?�hg�w�z�-�n9����Q�,���Z��P~[;`���;���O�#Ȟ5��E{�2���OXpͦN�-5�I��o�?jc;����%kĪ��t{�8B��kfT��E���Y�������?.<s�*���+z(�_�,\�һ�1S"K$�e�rB`�]�f��83��`=L:ǝb�5q4�A2{�a0�I�Z��@��wV���s� RF8m������4�6/��{OAB��G��E�]�8����%�d�1X/���X-��bǭ�z������Ub�+N�8�g�8�}�����I�����.7�O�I����t"R�x��5�ݠ��Zfr�<�L)^�����������vT#�B�vk����O��^�}��y'd�۱��}_ZW����+Z `b^B,
ʴ�3��N�܁�V�X/C��fӌk|B.^|&wJ�ŗ��4L�O��~¦��&}lċ����Os�4ɧ���� ��n�%�Rc߃{_�/#7=��p��b�V�RoU�<�66𦖣!�G�Ht*�sã��G˝ȏ����y��11�ۀTc#dd�&���i�vZC�!���&q�8��4�չ�W�>O�IA$�������a��!>U�$!cGu���@�H�9�� �,�4R�6C&�M2K_�RiQu�9��!�� ���^�!V�j�����F6�F|�Į:/�g}�k9/g��(Z�.�fߕG��jp�'	ˠ'�n�(a=�m�)���୏8I<��S��Vw�����Qa#逸Ϧ�p��0R,���w_P����5�@�,.MG3Q���F���>�z�m�8G%v�)+H^pr�g��cIt�~Q&A|Zp,d�&����Q����S=�t0�	���V ���g���~W�5	px[�,
��F�^�ϙ+�K��k3����r�Q�;y,����Cf�'�A=�[�&)�3�X��j^=J�!A��_%��-8AanpS=��6�6�)x��,�&"�V��}�J)H�P�&B��� ��c�֋�0j�����G��;$Vc5e,�
�:k��ɝo�1�G܄}&#���ry��~�g3�8�ʢ��JP����~t"uu�xB��a
Z$�.���k��;TkzԺPUi�Q�3����r\_g#!�f�;W��6er�;�@������	џ��|\�;��q	Q�Bj���/ �6<�v���9m�7qإL.b>��`������� J�e�u�P6�5�]^��a!�M,�[�&Cd���C�Du�
r�S!�/�A�`I�DB���%-Y�r��'��g;�Zt(�c����J��p�J��yoiB���ז]rS�2�F-h��:T�n�����"/d�6|�<q�ٸ��>�j3�&�ܛ�E�r�8o��1/4gl���+]�f_"��BLp΄�|ݾ����ƤC� �gq2;D�2,��T� �f���!rd���ʬ�@Y����t
�`s�")ZUi��XmQD02+1M��� �a;����Ģ1=������ӿC�SШ@�@����3���\%�;ĭ'�@�t�2�['�'�	yyg;��r%�p=L��e8N��s��#q���b��&GzX9�������m:���G}�"����:�|���v���Gg`t"k{�W;>�� +�%"��Ƙ�uSO�_/�d�q~L����a���;������sH	��}�f(üA|82����%/�����5~'��������O�k2��b��bL  ��� 7��W�ԥ]9@�޺�g��C�����ϥ͈�yNk��p�s�9�9q]����׵3C���;�s�����)K���%�������|_�jR"�T��
7��AD�ő���\^��&���%�,�ʛ�x�co+��P��:k�mH<m�j�8������zw$c\B,�34}�q�V���I�}�&��G��b�6Y9x��o�]a`�;<K�Τx-5��y�Q=����������x�(u�ۘ9fi�'�Ҽ�Gm���9m�R[���/��8�?/a����p�D*�G��B��OV��]c��XWܦ	���7w���q* �A�=w���7z���w�`vMA��8�����D
Q��)2;ܖ��<�� �<����GJ% ��w��m�à'D����K��DX�ًts�ІΆ��.�so�RZ�+�g���A�ՔjTڂъ�|�p:�s�����B@��(�u��Z+H��dwX�ru�DUr�����{!s�k[��sy� ��j��?��>t��h����v��*�@M�Y8�A��N�#�H+���+�+���!��J�~5N��|���K����r�
����+�����Rk���nG��0�e5�|F�wg���2�Mf�F���>��##4�?��{�i]������=�p�/���J��_��M0J��G�g^g�|�zQ�e�D�{� �~l�xC�v�h ~�d�2Ϟr��3�"v��\����}�ɋ�&�0��5���?6l�x�:;�W�� ���w=xM�p@����c�����6���[�2x�v=�/3��}O��B� �-�7 �>#�B�X�|t���o��;Gu�[�+���T��O����s����j듨0y���[*�'��~��$j&�.�и��5�Z���X�]gR���o�|�$F3�`�u��s%�=!�qj�M\�M������?z�r�JzP��cE��@��}�ģ���ם�����+1Z�j5�ٚzE��Ӵx�@e�K��~n�\W���i�MZ���o�mo��n_�q��o�J��3F�r�*W��Z�����L�l�*d4<1�0��~:���{�^��.>=t:�&��tX	6:�~N�9T����Ȭ���'c@��/5��a���S��_)�uM����U�$�`o�kXf��x�)��n��M[�=rP3#�4�&?�B��ǟ��6�^B�?w�%�j�����B�!)H���7L"I����l��hvO�*�^Fl�����l$ʂR�t��ǽ��Ψ1]�Z�������-��bY{����i�T��jG,�U��BϘ�C����Ӌ0S��ԡHY�C�%�����V<��)%�ZZ�Y�4�ꘀmqg+.�-8�^OZ2AK�c
# *<��`�ks�Lԥ���qY����<�eh<�F��yOg��i!���S�����jC���g��b�2�u�|-t�&�m�.�Z����:r@ܶ܅T����󹰩�1
�b�t����nܰ�4��П�9v�]vɁ��}�{^|�w�!K^n_�ɱ�_�Ul�]����� �W�u�j�]��u8o�c�p���8!�HZ�3��ԏ����D�*�P-�ӈ|�On�B���-���v+2l��]��;��~Ʉ�|��J٬�Aˤ+���j�,���A	7�y&�ݳ-Ym[�9�f��4
����׉!�7�}w�e��ל�]�
�d�i8����3�)<��w�#Q��܍t|'Ҵu ��hJBW��}�����7a�'sPhwQ�`��<�LL���L��Upg�m��L���u�Qx	��݆�3����̓E�0��9�#>koz��$o�%W��9��bz��4�!�m�����Ӥe���*��-ڷ������EN5>��n�����,y] Z�F�g�8�#��^Ş۞d�7��]׸f�)1��;Q��o6��BE��|)E� 7R6"Y�d�0����a�O��h���=���7����ޗ�?YN:�8�v���r+C\qTa�����%-R����H1�LЍ��%4D��Mg �����i 
��sPԣ�C�J�V���txV���$`#�H����l�O� *�X����c�<|n�+z)ډY��6[Y��i0z�S�WR��ln����	�h�<�4?����'��AE P�hd�j1��e�8�f�T�F�����\���\�Kֺ��pt'D0|PT,ZxYP0���k���FaV/�|ZB�Um�x2����!�'-��j��,�ЩӒ�^}_V��*��VyS��sϬ0:qF3���t�g���i�Z�B�Y~6f�Z6�OLƓݝ�+dg�����܀e����XH�e�ʨ/�+{��p�;�E�Rv}��x�U��8��)5���7����3g����=�v��vJ���BG����KW們� �����oW̡�r�j�SO_����6r��l�w����pQ�*�	ؖ!6�~��j�{��F��	� 4�D0�
N�gTkhȇMX%/[4d:{��^�x�A?�fUlh����xi�_�|ZT�hC��aZ�8��j�+J�h�+��3��d�֠���
�$D2�g �XQ�A���7V�Vʱ0 �}�-U�?#ʯJ�
A�o0$7��M|2�Q��핧�lG�>����|ȑ�8�O�\3����u��Q�][X�\H�u��3j��a ���,�}@�<~��b�]�yz�X������P�&����L���>գ�]���i2�ܷ����F��'dL����x����@Gg�R`�ST�(N�,d��yC(��F��'&8�����?��E]O���N�J	�&�G//8 �Z�DK��xKD�m�cu�f�R*�i�5�(��W��*tqI�A��4�(�:��"��<�vm|���[����Z� #f"쉷�g(��o�s~6STF^��V�q�����s�D��L�AD���l\�Q_��<_D����(��?V
!(g��<*`;fa39âO$�74~���/�ew�t��Q���4h�:�b�yU��Ze3��L~�B����Ӌϡ���&�a�y�����u� J�!�n�gG��������,0"}p>�@���=�r�Wϒ/�ߍ՘�3L����1LK�,BE��ҧ|X�)�0���� 'SĎ���;{^u�I�yU��"�]��w�T�W|��>��B��iߥV���&��5 jۿ�N	]�Q� 5#��O�G����T�M�Gp)�#/>�������G��ꘗ��~����OU�U�uWd��=�?���F޺��_�v!3����^�&�I�V�9�*r|KM���7���F.��a�$� ��Me���3�ι�S{��9i���+�14�M(�0���:��;��Ϻ�:�rԺ�9�E�Ka�����m!�ˌ��̦GiN�����e�5�+vk�0�<�(�F*�@X�W�yzϝ�}&���J�P�]��w�~9����kZ;N��~:����*���,�Ų�{M��j�o2�6�ٔ���
�J�z��K+5�ѽ@3gWot~��~��C���A��oF��)�F�0:&������ҎzG4j�v<9B>%��ks��y��.	 A�뇇b�K�&��6ʅ�S�_xrK�c����iф������Qlʱ�*P��>��Z�ٰ��^��Ӆ��b^��gn�/����D�*��8E^J��C-��w�Tޭ%j���m�9̚܈M�T��Tn��e����b,uŇ���� ���,i�^�,�}�"��0��@o�M�2�L-xG���\nr1�8D�����F3j������,ݘ�	*�pD���_�{�-�����_�ze��oY�.�C@dJr�X^�GZ=�IVi^,@��qѤ�F]O���<<�rKYr�+�ǪN!*W��P�"C�h�8��H����QLێ�8/{{�)Wm�8G��T�h��r�����vx-�L݈K� #&�E˫<$,�3̡$��8�i������&�"�R�u��˹�ŬGp�{-��z�=.�J|�3Pf֬��	q]�Q<��[�wp2F�m�όS-M��$K���iN"Z]�ZQ��j�
m�[�FI�h���\.Ⱥ� x+��"���RJ�=a[�oV'�2k��w;�Q�(`=�����^Q��i�7!���KU�&0�P��m���BLL����ԁ�����
?X�\��>��L ��#����5�~�`,���sS��y�h���i~a�e0Цh{��ɂ�ysn�U�܃�Ʉ�d�`h�����DGz ��^�"����~�\���B(V+�=��Rȹ�.dغt��1ƣ��7͝>ZW�� �� ��'���L7y�OC+�I����Bs.5�ڜ��>xX���M_D0Iʎ� �]j��[�kkV5Ь�i쒳���%�2;,|S��HG2�	){±be���x�]m� �&z��+S�OH�Ɔ�BF4�+�C�t�;�8*VNb�ceoǃ]���P�Sk�b�?=Z'1&՘Y7���%& �)x={��	 ?v�dji%a��Ǥn¡�	ȫ��˸w7����EM8Au� Lb�#�K����؆jҴ�vh�#�n�o���0��m���>VzI�`���`�U�+pC���Cw��sщ����^]����P�31ŕ��6���~�F��5����6\��ڽJ�z����+��J������3��`h)��W��Y��(H�	N��}�/�J�
�2�|/��DQ)���u�Ӗ����rpAH�sӌo�rd��J@��2Kا��=[6 &A13a�D�%�C�����C>��r�t0�[2�V}����Qf�z�"C�8�����gs���R�Q�I%�B�a8 ~�8E�	`�,1�2,��7�0���u���mL:�;��u>�?�1��O����.��9^$|��L".�y<� ����݊�jߋ����@���jn�7�I��nm6Ze��ڸ"���vvy�L��3.le������W���5Y}�dO�k��6����=y@ �Mhysu����a�O�U�(�КW_��J�ˁFh 1(�C�@�n�<;�z��&�f����ll|>����XFf�fGJ�.�>hG���'��G�4Ń�F�M�81��J'�#
�c���LQ7;�"��о(���N�;=8p���^0����j�F����^�Pu�..���#��E���@��4 *m�:Y�[U$�����^�d���,����1�8�8�p>�����&�������{�${���(&f��6�C�ӊx�i��S( �hQ�6�1��i�N�xm�a3Dl35˺���cPq!^LuC]����T{-Ϋ($��	^�N
B(ݎ�
*��9Y�;D%/I��nж=��Vă1y��e t�j/"\Z����Su��
s�N�{����G�&�{���P��K�c�7�G5���JӝL=��7��P, �ǛJ�֙{B�WG1���:�f���z��l#u�6�Rŵ��������a��k�x�A�!����$H��N�w�򴵉'�#0�����c�� �?���ڦV�7Pu�=���h���t�!:�}�X��>+�a�Ya䡏�1����Uc�Ȳ�B�����KZ��`�'v�������ȿ~"����S:����G�	
v�/3��(-��joN���@I�M®��Z�&,�y٨%��W����M6&(��܇��C�'��繃Z����:��@c8��ﭓ�0�I�u��qꃻxdT
Rh˩����r_� 駠R�+�˛g  ��EO���F���"��5�p�5�A���t�m`ϯ5V�˼��h!K�U��V�R)�[>X���/�^�5�I�'K��^c�n���C���A+�K��5'�4zY�z />.޸�Q��%��f�ܰdh�,�ڂz�A'�PZ��G}��	���9}0�C���w��[����������e?���l�G��~9v�n|1���V�@� 6�:T���������emv>���X��)؅A�	���K��eG�+��]Y���Ď�m�<�M,����Qj��SD��8��	���1�&4Oa���$�zٵ�3��?�	�X@��>+-�٨Aq+��Q��C/u��h܋��b0�'!��p����+<[��x [���4%�'Y�0����>��9��ޑ���I(��͏v\��6�ڊ�h�f��=��#z5P=�Z��bKx�Tf�,����9#G�R����`�$��w�2QP���3r y�=�;�7��Gk��gB���s��0}ϳ�CIz�=r�ZI�*b��a���,��&�]���Y<�[sz_л$�oM�t��q�*�V+hg���|~覭f�c��d�O4d"!���5��ڒEU�o�z�uf�y� �����!�ӷj]�nn=������?�r;�)�O&�_B?��e�\÷�g��r2#*�4�ԫf<�K��/JWWz.�m�:����v'��^�Y�q�ʻ�(�v@�DK���7�&ڤ�?s>{$�wtF&��gſ:����GBba�$$!�5S��	#�Е�_���j�J��Qd�
U��?���6����ra��t���^����N���L��h#����5hf'nl+	�]�v�ш�F&^�p��:W-���`m���4�S���#��s�:�6�خ�b�vl�BD�tX�'��rpߑ��r)]�֝}ϵ�Z����X=|��/KB*|�VR�M�U�e�%8ө�t�t6�U�Bg��V�xP9e�F��+����X}v��WC?��H�"Z�6�{��NF�{��F������\����j���ۏ�>f��'�9��$�=��*�g���|+���SI�Ӫ��݁�s��ʺ����ѻ��vՐ&��NM���Z�9U���;�����z�S&��=K���L�Hс�J�Q=��*z_`��tm�򀀠wkE|���88��6̘����4&Q.���>w�TߌtO�ZvB5C��9�gP(��)��7i�Ȉ���	� ��YG�Z�p���Hm4��A��n�)x��|\�U�ꌃa*%[�shX��;�T�b���1/FZU+�������^1jIG(&�;�$��fk�b�ZG��m�V!��ػl7:��¹>��7�g�0i�_V�:��;�����,��f�%�v�%$��q6��>�GZ_��1�}b����\0�_�MY/�*����n���78� ,��{,e�X��ѯG���,-n�/�8��p�'(��db�i����[��PT������Gr`R�s�ٍ�d��̗;�,�1�;4L�i~�f_�eT�U6�z��,~D|Q����\k��z��T@�^�����F"�̋q�;-���Rt�T���8|b��(-˞��cvM�2� ~_�����р!Î1:]9l@�G�+��Pi��(͜о�9Ҡ�4M�^S�Z&Ё�[���գc���;l������~u�1y]�����\�?aF!<�#8���4^ �|b�
&DF͆*���i�;����.�����A���{�&'��t����7ci�˝�nK��W�Tɻ�z�#t��� 񡚿���ȇ�$)Er����.���F�	᣺覇	:�܄�A�E�B���Y�����][B����� �b�imǧmcd쓖)�)�4d*T���F��ӯ\��ₑ�4z&5�d^�QI'���M�^**z��?moHB4�T�ZxH�w6I�,Qg�����+|�b�V
H�t�4�wLg��
��H!{�X�[ž7�|��feQ�.ˎ�^w���b�xw�`�C@[r����=9Έ��$%Ƃ���*ݰ]	��U>�Z�Mg���n~��=6�c��^�7*�����nw��_������\�����0�@j��6���8{�������5D��Q����A.�iN��Oy�KS�QV��l���u�?^ʷ ����M���2��a�G�p�Ǥ��"h�0����A6o�C���Qz�`��?�HRpԌ�B�AE��h^�Fp�����~ݦH6�`���8� �q�S�~�,fVF�޻��B,�
y�C�Ll��&�%$��L���;L�wh��2�w�5g��2T���>�T�䟭�T�P��i�����F�?b�/�)�e"���[t�d:���<d����U�HaF�}m�0��㽕�b��
�e^�%��4��[9d�ڇϏ��l��!6������]AR���	�	v�CO�v�/��N�ڌ��o�<�8ʪ�4�h욬�}T�v��q� �"�h��:y��qT����Q����l��m���B]5����|��$�bdFO�m��h-���Tl�[O(�y���Q[#N�]-�v�)c:��]�6�3�r�^ �],oKT�˗ ��h�����x������v!�^%�J[�V��ֆ6^;a)nOx��Ѳ86�ݮg�_��ezX]Q_��hk����J����^�d�/��N}��%�w{�&D!0���W4DPX1��
�֜��b���(���n{�{�o�����a�\��z�y ���'�т���$Q����_j){L]��wu���"f����[2����E�`�q^Q.ф<;�B�� ��}u����m�zI��J�NP$]e����r��^|�g��p!%��o�*�Hr�͢� ZP�9W�5�k�50��\�y.�%4EH���	A�,t/�	k�����	�O񈕚Z����cCE|첨ͣV�ȔZ�6D�d�k�g+O��2<w��㘅hd\	�Y.q6�'jN�i@K���(�08H|�ѧ_�%��Щ������4d'ĖQ�������>*�6u�\�;�"Vc�b�hp���\ZG�g��p_�m�m���.���g�;�V����;�'С�p�b2�1N7���p��&����L(�Q����c�v�!�^�������j�m�XG�����������<���$e���}��ĳ��_���e���z\�*;��n�,��c�� tǧ+���<l���<C#~m�\�n�,d�B�A�w)Mm�_�,�K����i�����߱-@P�Ei:�͙D�'*��y�˽���^ZW[[�D!vO��;�m�
�1���a��@]�YU����+�Fݱm��m4�ל|����u�~��;����^������o��7�0�g�\�7̦*�T6K5B�}w�=��l>���)�|����d�B�-a��&��×|��R�M�����s���u~�fi#
��w���="�@���d�>ꇩȅ�'+�ee�5M��H�h�B�?*�-aB]�)��M���;�D�����h��w��H���V�
�\��M�@�$I�HB�?w��|٘��������EЇB��R/7eWS�ׄ��¹���I�~d� �I�늗ؓ�t +��|�����h����w�R�+t�j���9���G#e���g�%d�g=Oɼ��M�(0�e���O�!KB��
|���NZ�{�-�\t��D�5����*�1==}�ƫ]�(�0޼E�h��G5�K7��_�� � �>a��,Q�]/�w����6;0c4Ld��2��I��*1�])��[��K2�ʝRB6��>�U��[Uxz�{#.��ً��PˬGh�]�YU>&���pvx�tH��.?��L튕VGU `��)�,9������!���D��rႫ'�X/}��=��?L�BR�pP��ɮ���*��i�i|j�x�p;�KFgZ��J�Q�וB��hIZ����0�N��������"f�O�ڍ�ؐ
���y���G������nS����W�3�+pR�y�xM�=`n&���ݐGРR�ͲM�w��>fX"t�ц��Y�����w�I�����^*Jz޸�f����: S�Fv�m`!�w�+�R�1�&9�<<�#goz�=��Plx�������}e���U�9*�k�j���Uv���L!D=R?��mP�T�RI�5s�]��Qmnu�t���c�B!�ʈ�<�W��K*`�W��1�p�S���m������*����,�
P�6�PZ�>q��yx�9��b��wB��u�P����zgX	������;�QȊ`ml�w]� �b�f��(6fF�����0��ַ���gC9��?pllP$�x�^$�ؑ֝�ݹm�pM2y���ߨ˺�\ˀqaG]hN�g�.���r�?�6U7XSo����)BW(X� �݈�y(|��0�A�v;_c�¿����b�J4e���˛ɫ	�$z	���C�ĒcČr䨣�������>'}{Ύ�_���^_۔c9Dr���T�h�����N�U� P�ǖl���Cg�0t��,I��ݔ}TZn�g%!lP��r��e"��H��Z�S��4f�v^lb���p$+>�nxZ+Aa�z�=s�8��7uR�|ɃX�Q?J:�}��
�	�Mpo�U���^8��
blB�m_��Xx�f�� ]ԕ#B��>��I"#�O�G��~��s��?�^`ز���LG�A�fOތ;>mO	�ŏQ퍗$�CK�14�\#�;�E޻C������;(C�9i3@���أ/fYRY�0I��W��j}�f`��L|�)6��e��v�'
;D��Rp����{��6#��.#��Rb����ReوS�Q^=��j�='Na��I��A���#���I�����s��\�Q8^��z�>�tb�s�M��A[�l B�����?dB���Kߢ6����
� �񰧹�?Gf�>�f�9���GA��eB��Ȼeڋ�ғ���a����Ay)���e�_�b�!�r-X��� ;&X�#䀐�~�
P�>V�ue�#�4��r����57R��	�yׁ����i/XD\�_�dS�.�r9�q̝�UMv��J/����>dW0���J$���]" �Y�����h����/R5DJ�r�e�t�3�]'ܟ�w�	=T�B�d&��Q�J|�r�@ F�RHZ�(8͒�L�9�e{�^(^�_��(���~�f��O�mPp�����j��`k��J=kǝ��m�+���������is���{�(f�+;�I�T��x�p�Oӌ��Ǡ8Y���<I�(泈�؞^<2~���t�쟲����!,��Ra���-
�Kl��^�j ��-��ׯs<�rAr����D��J��}̬�i;P�/�������D���}���lкx�B�Y���U;x���Fskj�����L�k���}S������-�й�g�&86L�tJ�x�mؓxMi}��)�q��CrC�B����.����/��Hg�y�҅�j3
u�%��l�.�6���5%�]��S��nk��ѩ����⩼4p��_�/�>��1P�{���?���_�h���h�4��-�Ў	ب�TӬ��އ F�N�|���`�9��;MB��a�v���"0c��9ay5	�����f<�l_�ջ��KT�I	�X�.[[�@����}9�M�H	W_�8��_�!~n�e�j�z�:4�բ��|YhE����k�zޣ�e��760+1	<�oߥJ���j�|1�I��/�|��hJ�8\L���#�g�ށ�qߊ�[���g9��,_fYQ�_E��I�R��.:�Yl-��	�����L���B�f�b�_�@�)�pvs�KZc$bF	T���5�jA��$��|$v	Lں���KoMZ�IC38.Ҏ"3�����а×.u�5ۋ��Ϸ��za�g�)����}��6�̙d��B2�bP�+	˱��g\�Ȩ0��6x9�B�專������j�W��򴧼�r�-X���k���/%J_�!ʘ��2��L��'�T�>�tStM�@L��f5x=�܋*o����3��*%2�U=h�p>ϙg��(Fܦ��uj���o��x�\ݝ�j�-��{)�8.u.����%	���~бz*�WWz��P_�������A��<�'^t�A}��ϓ�Zň0�/�] .�v�y�2�/DǪI��{�36�r���@���#�~�;Qw|�ȳ>�^�g>9P���]�����;�a�-�ʵX�I�$G���ڄ���:̳� ��
������Dև���Z��Ňb}�1=�!�
�U��
�[#���_�Q��}��˺�P�x6H���6�]�8mS��
+�Cy�-⠢�,��d�b��s)�$Xc2T$˳��D�(섾e�	��}�=Ɔ��p���uaSa�؋ͬ�:��w�
��r��!H>$:�n���U4""ƛR�Ol*5���B�8�]cv�A�,�8b�!��3ϋ� K��"U$���L���߀�GcƜ�h#N���5}�gE�ͯX2�>2���?x�&��RI53��҇b�]'�o���6n-,�S�9��6�}by>X�;U����z6���D�\�K��6��`ت�38Q�n�
}ys.#AO]�z�Z�ѥ��1����Y��S��I0e���fSm�;�{�R��� S�-u}���@���{�>w�\d)���[K��8r��j7�1�{7P��E���!s�f�}z��&�Z���nAa��d�-frO�
�P K�kſ"[�b��J_��<;	l��ٳ��i�[F�03��{�s#�>��n}C����;�3�.�wq�}Ą�7��*c�xh�t�&؂�3V}��->��\��˚+{�%K?���8�;f��\Xi.k^yQ<e ���Ϛn�C�p��&����ˁ���no$�=�h�
ٚ�K	Jb�y�:��8c:�=t޴�ݶ�ӂ�
��NM�\�1�}&�K"�Ғ�����7����@e<�NT�%pBkgͤ0 3���L?&J��:.����} Q!�H%}���7B/�ܴN���^�Hv&��$R�:x���r��9V�a.�~�J�+��NjH���@%��Wrܲ�ͧn�Z@���s�����O?�����f?0��ŵg� �կV�7ܣ|RQ��H�h�D�����f������z�	:T=B?�!��!  ��}������l-��y���wc��N��9E�Y��zʉ����������dτ(��?��
\^��]m��t�i�b,l�l����A*�~�.-ڹ�`l�wt7��^P�2g29n�!�2��ˠ�H�B���k��8߆�|��Tm|�1�z�&<un�g��a��X �.pW{�Ѹ�f�����+ �G�5�I�Z�����jpi�wN�&N��mh�1L��f�$�ۭ����vjا�'�(�60����YfSX;�U��Y�ܧ�$U`/�[�����u�L!�l���&$U�a4����@l��vf�%�������7:�C�_3߷EwwȾ]�K�!��IH�Ĺµin��eZ����G�r�*�/.`a2��֐�˅��
Y�s�ہY��B�����z�1=�E6R��-��~{�o���H��؁w�Ȃpf�S�Ǝ�����n�f����7nv#�Ȳ�>p��ڄ�.y #E�R��1�iȹ'»�y�4��c%m9��-w�7�M�3����.j*�1��j�i�����B�LB�&�.���
�_L&�U#'D�M�PF���M���y~�>�z�j���r�N�����eM��<��0�%�`�LU�~��b5��w�W��|Fu�h�VV��{�p����`O��׌�3�y>sAq�M	�����4Z����2Þ��.�Ϧ����Y{����e5�̴"�����XHb�2�S�=�]b���lЈ�*Tz������X�;�d�+���/��U�rˑ�5��%GU��⾁"zA�*��/@��^��z�l�i|�u���9a�?�w�Y�
A�e�'�L�����DO���rkO"���0��e
�s�@щ��?(���e;.
Ǣz��s	�K���JL�n�2�e�6ӣ\ڭN�t���1:��Ӯ�9�e!�\Μ�5A��(��d5MHbɣ��a�ǣ�~���f���v�^' 3 N/OW�Yc9^ �3}%���7��p"�T�]rv8��/���ܿ*β�F��GEz�Yx]�[}�;&S��;� ���J]�F���Pwۀ-�VN��}ŧ�������L �D�k��.(3�&�?:Z���!������$mg�r�.ͯ�&���G�r�R]k�� ��\�"�P;����F7J���q��F(-�P��-������j����_"5�^Yz�],�-lv6^h�$O�lktި0��Pq�l�����%�)X��*^k�:v����А�|���4&iG�K������E	jܨu����q����~�D�
�xm<�e��L�D8��$j�K}Տ^��?r<��Iǀ �^�*U��`$v��K��]��BZ�Ua�@>G�"�c��cf9�p?����JG��R����u��fɛ���߽瘯�8�Y�NK��	�s��|�Ȭ�<�2"�S�~i�ӆ�r�2sT+�����	:3zmJ�a�#܅ �74|��-�;�߂J���y�<�Up��;)�A@)=�@#%� =dۤ��9h?Ƅ<��5k:�6@�i����w�N��@� �L��,I��dQąۤ�e��?�F�J#��W�Cj�iށQ�l}|G��췣@	��i*vۑ3H91��1�~]��v0�@��(�u�i	R�`}t7��͸gvG���m�vIY�-�T���$]5�˨ŷ�'!o=�dNɿ�bR0�$�-�$s�8~i5��+��n��|&�Y�{��#���I9�{G�KݻT���$Iiy� ��q��uo�xP0W�Wa���;��ï��'2���6��_D��p/R�
*��Q}���� }�|S��ȳ#��O�V��3M.N���*��	
�$��?�tLx��ֶ1%G�C��qA�F�7���t5��:�*�&��+�.�Z�� n)��G,�L���]ET�:$5��x����d�{���큚}>�Ic�p�����L��[��3�#���x�'2x����iB����g򫶤j�~F�Dt��u��}�(�:kF?��A�<�M�M���ph~k�95`�F��G��Z�yp���ږ$��� �N�XJ�vY�Kt��qjG�BGsP)�[`�VS�XŊ�b+�����2�p.��.��MJ;� ���II�#ߡ��2b�J�ߥ�g,d�E[N_	ڌ#(��Vґc
��"���LDK}�\uw ې��n Ur��������'�JCЉVjx��9%ǌh6�콙���j�`��6�(�)����85q��3�����Ϸ=?��@��M���Mu�MkW�:��z�%�����D�����jn�>��!x�Q���*��0zڡ�d���5K���%D��K9䑔�43$���%�@[v��mxxֲ�>X0NN�܇����p�U\x^!���2��W�����K��o�����Gն�l�mh����6��r�u՘[։�����g�[w���Me(1&�#��p��W�F�e��|�2<d��Īl��YMy��Ъ!�0�a��_���
7��T���.]�!�$�r�C������"3�0��U��,A��n�z�,���U����)G�Č�p��N
����O>�L֚��Q��#�$�l+O+��g�1��qΟž�l�~A��ʋU>��^�,�����=�L��晑���T����o�Y;�~�id�h�9� �^��RL�F�@	��Ap>`(�p�Ȼ���%oi�U/u2�
N>F�D���5�&	=��Xپ�i�����i�S�{��ՠ�[�qhn���Y�`��%�[��G9�m�oN����1@������+<�̿ �I�cX&�7������Tq��j`FF	��y��8����t����7$K�6~�&��`}��֊�>F2����K�8��V�1�P�G�f�ٰ����I�����a��l�M����z��uj�A���&"�;J�=�����VQ�b0W.��T�GN꭭#
��C�Ĉ����WޓVY�B�ELLVBɀ=��F�_iV?�pA���ܲ�-t�T�b�0�T�VN�N� N�bd�>#E�N�]x��mJS�������P�<��p���>��?���c�ܠ��?rWƵe�F%��P5>�g�LJ'���cJ���Aˤ�]�Ǘd�������h3c��,�q�A9��2l�������i#g7�e��m��)��Um�UB
�ҝ��G�ϫ����յ��&� �YV\h=��WYO�Ỷ�@��g��O��;	F��4���������A���}#���D)w��sgJd:�2E��f�Kc�=&�l��a����ո�*�R����_��Ix��j|�&б]�pC�Ƿ��,��U��4��X5H��|# C��xc�pQ.leT44������*��x[�K�5�<���wq�k
Q�	�j�����GN�u*�'Cr�7�ć�+�_�
���1���I�o"9/�;R�^����Р�i�Z�
�f,Af��^p^�"^c�LE�<��<4G� �қ0�?�ד�`Ɠ>#f^��t��}��⏊sTg�v�7�}�Ey���x��@o�����(�c�l�)IWel�J��l%����q�^�tZN�Ys����|o]�}�Qbj�-�'{�d
V��NQ��a=Ǯ��iĒ�3qX*�y8k�Ov�ex�2�>,Lٹ�AH�=նʃM,9+B>���co��_��Q:#��˫���>�TQG�ݿ�dڹ#�嬺-A��u������q��ov8�%u^b��RyF)�j���� �aہ`���.#�6���K=�i��lL4�p��ڱr��WS���>b�->�\]�������Cy�0���]\L�:��k�o,�ܡ��shך�z"�N�E6:�8q!5Z�"U
F��	K�Z�	]�Q����_f�avCQ�4�%*[M��H���S?xX��\��K���@�3-O����c�E9�fR$�ѸIf�V<�ɣ�t�v�U���\
/�D(eҾ�YMM<|0)9�V��{G�d�M���+G��ݙ(Qn�#�b� p�n�Qq��]�t�Z#�!h��b�G��d*  �yf;��c��]lX��W�p��9
��e�,�M ����,gM�1����	x���Ϥ:�z��֗ҡaT��#��k}��bi��[t؋�v\Jt��`�����	�_|���I�۩�*�de[¶��5\��SI�MR?�>��?~��e��*L�����R��p��"C!_��68M�J֣#�ӦV�i!*G*��fSF��VG���_N��*�KꟵ`�%;:�vn[��Q���J��9v�������k�-.�yN66ϴ�`/�[uPK���Q�l$�?�ߦb���G.�IV��e��@�������}(����WS3[l�eFZ��!�Z�$�+1��h��z��L#���;�6��yE]�Q�'� ��~�
eq����m���U�>g����7WD	��}O$=��V�֪A$v03��$���D��v43����Ӫ5�V�ً��{+f]�8V� C:%���1#��;�(��άm�[f�����\��{��-�����"��<	�v��ԏK�-���Λ� �yq��'���XHc��hL�%ι���Ӊ��X����'19]�����8� ����G�1�0�i�?���ly;9Cˬ�>� ��$zW@�Ŵk�T��	ͅѼL�����p)��=�T$q��Q�Ʌ}=�Sɼ4OP���{Rڗ^f� E���E`���\ZI�@fa"�Q�.�g��Rm�Kʩ){����<�	q��� �B���pc�(
�����p�-����:i�-�m�Cx�U�R����K?�?�I��sk�Q�QOU��K�ٯC�Qa��AtJưO4јW: nֽl���t?T��V�����op+�l�����H�Atƕ^�	i�zYPq�>��i@˸v���r>	ˀf�:��=|ό�����jg�>zA���Ќ�kh.�<N@����|��%��j�O�	=������YL�P�ĳ���#�R�Y��Ys���B�-2ag�nm�(��B0՚�5<{���FB1-����>���|�B{��������i5dN�{V�Scq�qH��R�}����<�)��y�W�]}B�PJm�F�����>�
�|�i�=���9C'0���I�ӳ�<f$�F4k�(�phxe��"��Z$����z:8E����
;ƣGu�y�'R.�ʖ O|���q�)a��ǢUٹ�*�)t��C�(C�,�S��'�� �Ћ1Db�#���Vm��${�-c�E�L�z풁�nQ]��I�MU�r
�u�F�w�h��o���,3ʚ��3
�?����T9�(S���$dcW��U1���4��;���H�í��3��oy�D\jr�tY5������M(�z�մ��IX#Z~ޖ|�iSr���;�U��	�Z�PA��8P=0�6�q�O/�`��~��t�DA��x���K;Fq((U�%�]�=酪��vzq��&6�"a����W���]���D��>��	Wn4�L���}�KX�S�(��M�\��~�VF9�p�GD��#b)砜��}:���ΐ�<-]Ψ��lD�|1�DL�$�[�p6r��Ր�� a�����t���h����V�q�Z��_��轍�_c�~	��@�7_�-�5eu��zϖ�앫���8��<�#	<!$1�:���X�N��Us̗�1l�D:' b��2l�Z���;�s�m{	����I����h���=f43���_�)x�ŉC(���<���sV�\�kg�fxӝռJ�Z`�_y
��ř8E*Sp�m}_��j��;��(r@�3�%��G���`U�0������XV�P��1��~����$�Aͣ\��
`�����!�(�?�P?�Pn]+\�l�p ªcXm��`ȩ�L�t[�;]R�3��i�p��A.�&�q<���jD oOc��0�D8����T'�W�J����^��] ���Kk�m�����-SbI߀C{��]P���b�ԑ�6��̌�G:��59vE�>k}��H��pr{�z�uY��Z���,H����y��t��ϡ���Ҙ"�sɠ�P�	��rM���(qv�����9��ةѣ(CE��"Rb��yw��N	8����p��u���I�r�E?bi�O9BP�����}H�^��s�2��N��Ӳ�lS��F���Ψqo���vO�)^V�aP��l���[ܸO�A�F*^{]���r�T6m�m��Y��ʤ�<r7I�����[�]����W"~n��j�>B�p���6��n��|����}Q�7�%d�]��Ţ��'����#T}��֋&�A��@3�$�g�l�bO�m �5�0IFthjL2N�IV�"Z5X^Q��#�~9&`/dю�b�vay�3:�z�GY�Dl�mŔf�|�@���5�h�ñ�m�6�X�@�٢�l,���22�2���i��v=�1�˛���yP�䛲*,ÁV��i�Ŗy�W�ۮ�\J<����uڌ��mu�\iKʪ�A�R�,5f+�@m=�s�YL��B|#�u��V��N��:��ӌ�^dN��'Ek���GM�� m��P��NБ$VU�bޱ>���f�d���	0�,�a\-��C�L�6�Xy �������t.���2����b�,���#��2z2Q�w�{�-����(����S
d��������X;�Yvm"ߟ�$�g�m�	����N�>�3Z��5D��4eCg��;�]Z�=����)���N늞̌!"Q�4����9��n��k���<v}CA��@�����7!IN��I����#�	Bɪ->�3��U7�a_���,Yy�����Lgw������'�&+ի���r�Q���z:ؒ�C'���U�%쾉���O�� 嗗��E�?'��0�5)�Vjd/��p��7���LȭLCM��u�|�B{�~'a�$##�Z���@��8�(r,p���t�I0�M�g�<-Ǳ6�o{Ik���}8�,�"tZ�s(>OTB��=z� {b�������'.�3��GPa�A��������# ([��)�ߦѳ'�K1�:�g��S�9�S�[�u
۴hv }��SR�V��ߞz�Ryt��By�A�$��g�f�����)��5�W���!擟�r�rT��N��)\i�F�p�h� �1���?y�
 H1@��ȳ�$M�(���bgF�ޖ,,�bFb�Oa�{�λ=������hC�0���X���Ŏ[��<�}Z@�XA��V~�a؍�Lb�~ZQ�A�e�7����]�y�+NZ$v�z�������KYR��,	�jO�̇s0��UaK٥��?�����ț��F��؁�����A����˗O�L+V������N�1{ZD8��0N9Co��8��7�2'�>:�稯�������a��M��X\�n�o4���	�~����'Ƽ�r
�/~mB�v�Q.Ok"Vѽ����D�7_DK��Z��zV�LV��jX�����ߩ]sx43�eY�R��+�������$�h��g<e%�z��n���@��J$����e���a 9U>���`�P·o�Ac&�l���ǃ���<�{�p�@�f��A�M\���|[Z�m���B��F��~wX+[����r@����PE���VE5��O)m�g�@��Y�h���+X�6�'�eѐA �׫�ș:�	�NS0Do����xs�×�"1�:J{S�ۑ1�Z%�)�I���<ꩡ�9��t��	XD��װO�S��{1�5ĉ��0L�_Y��*C��R�q�L���6A�}��m�8(2�С��k���¡`�s��z�|g�Rc8���o�^�CG���#<�h�ܬ���y��W5�r���e{�@�-�v���'�uwu��GP���S�-!WW �c�o�ԭ.Y*ϽF�\)��sn��&�$�F�MSs��8?W���8�8ğ2�	� #���� Yd��m���>�`�9P&kͬŦ7Գ�yEX+	S���E�Ci�ỽ���Ou7L(�utA����}�&{���o�:��A�ze��<�	����U�U�puԍ�T,��i���'uO�`\�1�ñ���sꇟ�G�YZ�5�?g�򢶛�n6��Fg�v�u-o .����1ռ���n�M^wZ�}fҾ	(U�ͫ�G��7�� ��t]�����7?� ?�G�&��6�*��v�}�a,�~�k�j/{���QA
��4��נ���+��C,�|�٥�������!%��r?K@F���r|��������hZ&o~4I��S~Rf� w���~c���d��?U��!��)�2!�,�
{O��㕕�b� ��K�n�$s�l��h�e}�!����s�F�Z�䃟)vMeD\��a�f>w���A5|pdJ���L����qa����z����?mK��<�F���yY�ZeE���
�/��~"0��+�OYR㜷)�b��g���,̥�`����U�𥽁%�-T�-�:D�WU��Uwd}t�!O��}�����G3>�U�4�wJ]�Z�ޤ�Üc��H�4�� )�V�+��<��q�g,�c��@��P�VS�jL�z7�cӧ�w����)=}:�G~�=yh�X��X5b��:�)}�P�����i&x��Pd�i>��Y�Dsq�v]�y"������L��������7V�{�m2{� �N��C�,�
��L�I2�.*�j�3���09����@�bd呦U���6R��'��hm�TZ}�$��1�>�5�����{����`�$���F4�ٗ��R��b�yS�Lh/���(f�f�C���Q�dz��KT�~]阹t�qƄ��0͐L��2 ��xG�E�ݴ~$X�fD��[�g���]��!�:_�_7�<�)%�\cT�$N�F���;)e
~��إ�#xLΜ^uV���㰮v§r��{9�h(6�*o�B�ҋ�E���6f�L��Ǻ~.a�IhA�i��~�xRK�����;\�%"�����n�*"���FT�=�b�oS!��b��n��k()�],|]OVIS�V�Qݑ�dH-4�FU"$A� 
�IFM~��x�QO�{D�a��:�lj�v�CBC1Qzh)>������eI�zӄ�8}�U�ͺu&���۞�ļ���f���W�4��y����<���'��W�s|��ؔA�����Qd��,�P=]b�X�F��|�6���S���93'����!�.<7;�&n2*�l8��#�*�XQbLBH(���j;TՇCn���x�;�8�|g��O���X�iM0J���5�N+������Q�B�S&�r}:�m�?��Q����q��A=�����YWߕ���QBX�~+�ݲN�IS����6��X�EO��u����)��e��{�Gr�֢{}���8D\�sbO��m�D�.D~��o��m��>V��tT�X ߛ�OtfqS�M�G�1ʱ�99T����}g,*�Q��.D[�`�R\���4C%��H�|�g��V���j���m�8�ȋP��{�uq�ݪ��c~7S����*����G�J���{�V�E&��x�uWr0_P�b�8VJ������_�bgd��':��Ď��a�>G^h ��m\�:��-[E�c<B��%m�vB|>5��� ���S�T�#�U
�X�zz��kc-З  ɬ�X��lʞ��2� ��*��pxs�W�蛝��p�a�H�������E��O����$)�!'ɦk%��<���ρ�	�`���>\2vK
��_%O��;��O`����b"W"�[Ci�������ϑ���#jL�$�8�ð���F���E� o�j"a����7�7N1�*��AMn�Y����6^z
�0�y�	�~�/Ns���l�ИC�)����:쏁��o���н�����^���z�Lr�T�?s_��&�*��� ���[��=VΗ$"��Ԇ.π\��G�����}!x����zNs���8�ވ�s��<Zf�ny���q9?�ު�g�C]���D��1��Ы��6�T�����d[[2[����$H���z�5+�t�c��Ozǁ���Eu�^�-���S��U�d-xiMSPiz9��>K��s��3�>F�*�߭��lҏ�x�q���	�#=����p(�dϖI�!�`>ae��b�n����MTUٌ8x4�/0y�6*r�]Uc�}�}����|��^��M^o"�ߢf�4u����a �[�,Y���87rm��O�!�U8b2%ε��eM���1|�Z� j�vy7�>pY�b)p�W��O�Xhζ��h;oՎ7���%	q�t8K�-�)/��߻V�#�
x��fC�/�Lض��M��r��*�p����S��
!��-�T9I�]ފ�3Ʀ�⊞$Í=qD)����Is��S7������P��!�;�SI�����1�O��|z�9,M�f��c`��ᩋ��ܪ����X_������T�`�?��9'�Z�6�"ՃV��x�Kߦ�8�ٱ?*.b�w��渒��h��j�h��|���h�N.f�6�O��u�~������G�c�Vm-d�6)x��F]��N���F�E�7��j^md�5�(��r�"̤9�~�1��
�L ��5�R��$:%��$��&�X�L�G��9Ad[@8R�Z�}@�e�X���K,�+��5��d��	 ���T�f|>R�\.?\ʑ��0c�e�=
����|F���K����9}~c�7~�' ���F�hgȣ6�o��ǅ�~5�����x�-H#�}k��Ɠ왥���6����qX������`
��59�'i�N��ȏ~�(���e2��r�N����or���D�2M��'cE<9��
c���V��s�MΖ������l]��@�3[
��,C~���d�˒i��$�#=���_�&A��}�,�Zq��s=8w/)}e\ gh,�UīW6�\�N>�"8�U+U蔠��U����6�$�o_9��(��1l
��l����m�x�F��j�i?�Q�XS`B��37]�&�j���+��=t��Ǖ儰<
�q�*�~�1�3@?��ߪ�S�V}�P]�7���/��O��)3�>"���!M衤���Lǵ�" |o]J�	E>�`�l�ʹ�{���A�s9R�f	4L�ϏjA��������t#9?��>���%ONdVfӞ�<*�ܻa��8�oM�����и����6G# �7�B����W�[m�\�q_�y��%�T�`>�g�ټN�p��ոJ��ڧƜ(X��w��^�;-+}���>��$ł�ʺ�My��j&�B�p?n�e���2�����O��H��נou��3��`�g�vS��
�;����ԣ�p'�ꑾS�Cۘ��C����B>}����;R޵<I_@jGwܓ$�'�d6�����xv@�s������Х��-Zj�ޚvŪ&j�v��1s ��cx��v���{B�)݁G.��Y ��gQ���a��;?ݾ�-|Q��=�5��U��}D��?Pb�D�q��u���3��!�V��,���G :�ú��!q��Ҙ	�dB�3��]�+����hN �hDd\m��y�C�D�ɹ�m3�Ƕl~q����_��⬓�(���S�}{�P�g{S�-w�u#w�*���]�[�$���N"��߁�N��)��@"�~)�jO@�Hw��æ����m��7[ABM�'��l�l���;�o|�7ar�gƱ�B�[SrP8�)t>��&숼�;![�7�*�G����C��|=�M��?�}|�h�Ƭ��@7�_������zE�ws|��D��9��m�r����~�#_7_� ���*nቷ��zI	��>_�H�!��<�ޏ��pveM �xS˪���H����폿�����o����Hٶk�c?6:���Rn�낞�Eŝv��KX�@�5�tA6+�'DD��$��~�����L>��<���9�\��9z˖�Эw[���d�{�c/�H�tu�� #Nn?�c�F6K��f���r��.�D�����"PZ��i�X^i����3B���0���_vc�0�}�+99R8��'�A]����Dn頑?��C�T�E%��*]��4��	�A������iH�!q"��o���x�;�V��=ր�9!�y^Z+��D̺}�X �g��R��vJ`O���j�"{���''�?����ʯDo�ZaGf1��s̓#������|5\�ldc�ɗ>�/������WV���Nb�_IR�h�Hӭ<���(�Y��Lt>;ȭ69B����t����wFX,n�<9���>W�ڹ�pq�.��4�腶��¸��gN�j|q�+ ��@n;pn���vff�<��z�Pi�b��=��J!���|�*q��ۊ�ݫޮĴ� [7Q��_�5����M[Y��F�~3 [  k�|&	��Kq&�+%�?�RF�#��HA	@��gk.՜U:��j�W%�9�K�k�P7-p_Ό0��>�S~��8�Ĵ���P�=��}D������k5'�S��0Uqw�����"���B�0��r�f�a�Xv����:���T�ad3j����D,�Y�Z]�q�O���b��
�y(:}��u�Fw��\ (�������j�6�+(8�@ؒ�i�q���͓V|���:t�fi�;vG{��� �d�&�X2��m>ug_%�"+K"�mZ��.� XOe��\Q����~�vCp��C�ľN��f̋A��Hlf��<	 Z;+��yl�>M�_H�k�������ţIݼB̢?q�vq�s�am�v6������X�{�	Ҋ()@ӌPh�=U�s��|�r���S�2��I>a�0�]^�t�z�L5 _IFE�8 ꡁ�DK�ӳ'ۑ{�Z��^좝?�T�b��4l�G�~|S͹YށL���s?��H����gD
�_�WSE�2���{�`q ��g�4i�����f�v�����y��-�>��N]o�m��*Ԑcҡ�`8��;�ۣ�;����2�QJo���gR��{�{ӵǱjL|.E�E[oi�Vc�N�����r�Ĥ�Iby��mт��m�I�_�c����{��a?s�����8�A���T�o�z�9�[jo���C��3�٤^��Y���ή5|�5 �V�uE�#8�-ȫJ� ��R˓[<��PNy-�)B�P�3L�LF2t3���_�Ԛ�suU�<�����m�-ѷ��Սɰ����B����U����g�|������0���v*22����i�̷h���C��� ��jzp��$q�ͭ�=��ސ��0������AU�"�%'Ţ~}������r�Q��b� އZ��#զ@�؛�$㥙S���k�m.3�erp��X��HO�}Q&�C!}[r\��Lߙ��NqB?�=�uB������	�Jo�J~B�Jښ�x�Fq���̄^F~�n�!LL���Ehc8q���%}J���D�j�A'�	��5�m��|�Fdŏ��.]a ,$���M�,2�vʕǾ�y`���#��qnĊ�n�ɜ�{˖��}^�T�� J�߹��4���@;T��q�/��|D�;�t�'q�nܸQ�����f
�+<�P�nj5IA]�!��#�=yo�MQ�m)e�N 襡������Lv�Q��+e�࿛p9�� K5����>_�VA���e��l��1K���Np�=�@Lo����v=��R��4Z����S���ù#��K����w����H�j��
��Z+d�_R���j	�Xy���p�5���r<V<��T��G������a�٭�C`����P4�t7���]>Һ�'_C�Zm�]��)����GJ�矤M,o��)�M�_�,�kAo�<F�]I!��M3v�B����ovm�h�I2�#M�G�ITH���֔���F�ph���<{�����BR��!���������R9�q#��;��	�|���6�n���f��6S&2S����ޒ��H#�0]��g]��zPuD�>G0cTq�DG�;I����Cy�؂�����JT����A�?�*v�!�oQ�N�:3��Cn(B�*KY?P<���"���%]8ue�_Hn�&Ը�$��ʤM�Ȣi��$cP�~�koHo�l�D(�@Y�$i�S(���W�/�<(

�b��_@`jL�<#��2�
��/�)7�����Jg��CT��Уׇ����䂬g��U�^c�n�����&�4��g��2Fp�S��=�}�5��.P�dG/�����oW�(�<��,l��*H�&+���D�~jA����M���u�Y�k����Q��Vˁ����m�j�U�ض�w�]�~�掉h�o�/B�̉;;��m��Ե�%�s&dZ^B�ӝjIj �5��a� ��<�`5oq�����̩���=y����vc�,[`j���
{�@Q��-��@KLE`,�x�צa���^r��;���?x��Y
x��4�,��fU���k$c-�;1�ׯf6���?���%��Be��G�*����T�m۵���&w���!��H������.}�-��� 4�����UV����R W��`�s~B=@!�
r)Xs��k]�a��7��T&FB����'����	��\[4BjO��@`N�d�S!̹0C]�\R�����nc#/SP��/���,W�+�5J+��PK�~
�@��������h���߰�/?�C�c�����غ��}�ވ���:[4w(wU�	�km*�b��i��㆚���S��kœ���A3Y
�.Д�t��f=���;)���ҍ=��n��}�T����r]���lK�:���b���׍�p�?������O�N�mWv<�F	�V�]P$�;2Y��`u��H���ft�ә�侗� %�<h����ibC�FW-�
������c�²�y�vP���p�[��o�%:�S?�Q�MLK�MM>���g~�v�^��h�:m�O�Uͮf[&�i׺�����K8U*@�7���A����4U2��k�5-W���'�=|ِ�[`yAڛ����mE~�Ω��H��t�ޤi5�T���f��Q)�`X&x9
�S����4�i�," ҡmͱ�(Mk��5u���=����h���cQ�`�_�4���{���T\)G'`� 6��:mxc����~u�nk�r�ዢ
 Y����	���Y�6��gه��#�w2v�At����>�������tں�XU�J-��6�F	��p<��
�BNa�O�c���w��C����)�E�[{�%0=�B��VC�ofF�e���0IEĹ�r�>D��;aLi:u���K<�-��Ю��I�=��n�_;`��V��x���M�`f�E��[�01 ��$�~D�r�Y���N3�4GZ&��~�\)&�-S3TX^�Р��t�Z�~Hvm��z�)��P��W5����v(!�)����H�>�u[1-]��r�g^�A�۠)%��]
��ҏwr��5E�2IXB��Q(�&��?���Y��6���y��K!�U�}#O�ɓ�Z9�^d����߰��*����_!ɗ0�A$ڽ�y���Ύ��7�vD��z��L��5F�~���X����z哬1�aN��!��K�à��Km�kv[�{�&me$	�օ:�����p/'���"d)�tf�T8�/��`ێ�	Ҥ�g����&0ic�o�*|�2���а���j����N�Z�N"ӻ�77�ˀ͚%� �����cS��3UJz����5�
w�!P�9���Sʇub2:�
�����-�&�����zU0c�'K�D?���0.T!���GB5ш}��@[�S�X����(Q��K��(�[;l+�5[��j|����T�%z�M峕P�a8�:�{(Ҹ��B(���Q��m7�%�Π'�N?��հE��X�G��c`��׹ٝ�ؕ�v����,�jr��Qm��+r�ˁ���jc$q��P�R���a��ߒ�eyZ�Z�%�w2��D5x���?*,��f+�ܴ�ئEp�B�N�����o��=Q��G9��w��A�H��	�\W&Y�~y��'a�u�#�Wޗ�WW�e�FsI!rl �TG��� C��z4j�Z���c/��[R��0 Qi�V��{$fU�:1iWψ]mjY�d�0y���Z�1�C0y\	�p^���+(�����H�?5� �8����\�Ր��/~�Q}��J�[eG5��%�><Y�a뾞��[K����s���O5�E��8����XZ,*2t�Ҏr���$<N:�����~��"����������2�V0��tI!Ѹo9 <Z2^G����_%�R�.{g�cڎ+Ie�`_�~ "�[Zpyb�Xܩ��}�*�	�&�1oub��ܹ}���t�K�h�?�ˑA!��¹�|RL*���ض�!��ҕ�z|���m����
��J{�	�%�W��T��̐��^^
�9 �W��Qpƨy@�#,�8�:�:M��w$��~�B0� I��t�������m��H�&LF�`��#�ږu�l�-K��WՎFqt����s��`j�>3 �ͧvuO����G�t�p��KꄝD~�"X���D�b�|oz�H��(4�ݪ
��(I!Ne���\�����R���B/0:??Tɞ���k̗LW�^�%a%F��2��ۓ��\ʝb�Y�"���{ጼo!C���UD6'��{�w c��Io�*N�9VN`�hSu��՜��; �1�*��v);�0��@���o=�=껳u��� {̵d�;��M蛱��<�ﯜ����Oj��b�آl���O���c��6�e�R�,��W2�ST��%�a0}�8KV��V��'ȉ^����g# U�Yqش�.۟I�
��+�i�H��� {#�	�%�;'dPK�/���J#Q�u�"�,�E�\A6��oQ��-��7��"Hنn�XGq��2�/��cz��I����G�9��-���HL�v����F4�/�a�/��,����ᇅ���
����� pS����U�V��O�ͯp<�F���Y�a=�ׂ93q�]ܳ��,,Ӕ���	ɗ���]!{K���r����w����0`<����<�@ �c���x����fu�;�x+�c�ᐄ6s����-O�\k窻� ���5��-\W����ƨp/��Z���)��f7�rS�����]���ɗ�v�xV�j@謅�D���7�FK%;Qe�e+�M�b^i9gн赗����֋��q�
ġ�i��w����Ak�6� q��h�{�m�_��hb������K��(����q���Ӭ���z��B��~�Xu��z����+so:ĕ^�v��<�rn���"��¥ɺ������Ld�I9�=��^����KLU������94K��Z:�^>�N�|[خ�g
����+@��1c���rnEa�m�@�����TSnu
��M��N�^BRɒ��|��m ����@i����|��Cк�91߯7��V_���i��� ���z�c'�G�-`�S�������\�~¸Qyο�G��n����cq�R������?H�}S�����a[Z3�/��6���,T!,�g0_�&&�:Y��)�,�}�/4ϖ�T���n��Q����v���L�%u�C��mc tgP�	��f�� ���-vx���2��_��h>�s�"ņ����R��"�@"��j#a1�@I�GQ匨)V����"���\-�D��/X%Sԏ8��~�!���^CM���TJ��O/���ɓS&����q��Le5��^©��3�M,�j�-��	��<��6��m�����~��!Do�aY��R���tW%�b��:���V�>A�[�mUr}=��R$��X�
��-����.������D����Zmw�p�B����|;l��3m�x���!�y�}EK	qcW���M&Aэ������H�h�J��8����jD�9T��^)���p�6���s�u���gj|K�M��Ss����юm�N��1U���+���CD�l )��w:�;��N�Y���\�Б�=(���1Y��i�.��������g<��;�hI�R4�v��E�Xx�g�&'��0�ժ�K1����9�56�*&Pă�6��b:�b$gx4�-+����}��ǟ�64������":q/H�p&��A_�ԡ�PE@�u�jKWYGs������<���`/s�sϬ#�6�0&�I:˓��& y��A�Y�����g��n��A�n
���.���L��;�G�8 �7�ڮ��F�,�I�~�{����=��T� ��>���To 0���n�Y�;'�á(�1���u������*�wP#.)<����$����C4���Yee�<|ߞ�p�ja{�om�Ҁ_�Mi?�a�O�sI��4�M�(\j�l�]W;Ɩ��"��ȁ|C����/

���ӫ��c7�ю��.����{RxP��\����Lߣ�]'�,8]���+e�ϸ�.WG�B��5�a�^��w�5:P��l3���.6#�ہ�2"�c��f��28�Rx��>��F���6g+�jj� �)�{�NS>�{w��v����'�<;@wَF��3��v����Џ3��I������L�Et^��X`��F����u�#���5t�f��#.���V퐏Xi���.��"�fzB�X\�*537fq͋t a�Љ��( #I�l��k�<������s�އ�/��u��Q���A�x�_4��F�0���[�'���z:x �&��za�����-�C_�GX��0�~�mqe}���C��;���.�6R���N��9э�������d��׷�8�g�밅2��W_�FCZ�0Hb���4bH"\<��> iu0��2�H�.���.!�ހg0��f�N���ѥ�r���5� T��+���/A��-����wr�T�����T��H7RR�?W��'gV3@V4��x�����D�A]Q� ��Xw���B,]�u/��i8�硉�C� ;�XBw\����S�9��-������+�"lS4-�~2�t �e�3��h�B(}�D~X�4G��|&��_,����CT�Hʶ��ő���~׳"�xL�} ����r�+�`��L�ݫ�>Z��)`�Y#�;�d <���Dkv
��Ƈ~��0Y��C������.v�m�y��Z��y�v�=�Z��������(5My,�b|� �#ҠV�?w����$}ŧr�*Z ͠��wnx�x�><��c����(YG��\T��R_�C�$�@9��?����#yg{�ɠ���RJ��u6�j�)gU!���d;�������"ƽ��)�e_a��~ڍ��|b��l,�vja/���\�=Ljڠ ������'-ZZj�b��������Q9dՐ��s��6^��*d�7���Ō)Q���W6�􇴈n(�:{p�J�nZ�Hx����]y*oE5��'S�B��y���m\'6} �� 5��W����Y�@;�UL%��oV���a�٪3�s.O�]{�Crg5-1v��z��C@t��r����K�KY��	�y�$�ݫ#=o�k!ˤ���W㷩�6"���BF?C��̝���h�9�xt�l��<%7A�RH��ۢL(�O�Ƭ�x�שh$����X���Ő�U�<uV^������7Z�`G����8yw�P�Ғܡ5�"U�����?���ڴ>擎�US{$V�i���r35���ЬR?e1�^̣�[�+E4���Rs?����Bj-�+e��#\j�7�MWr�}����~�-���P�\+����UN*r��g�&���B7�.!����<�y��ن=�0VOi{k�+�����GD�W	�-;�i �z�X�Р���x_(�m��=����&uN�kGc�����jj�E�G|�&H�bKy���1�k�`1�J��A�&���|M��n/qV>aF�,f(��1ԿӐ�+C���I>�����Ǧ9igL�T�_����t�1y(�,�5a�=.��`�s���V�z���+�a��hJ�!�c6
����<%����=(�7���v����{����*�Y̑��}1#�`m?�plj�#��0�"ҶYw�\F�o=��W�hϑ,Nc���f�\tPz~�+�S�X���%�,�������ԔQ�t�~��7���uU�y�S�֬��N��7{N p��l�P?��`DMh����<�U�Z��
��]=>x�̅	���v��R6 Ne;<�����ʓ�%̻���y���0�_M��c�F8r��Ż�|�Υ[����c����E����݉�jHtk���G���}֌������� �D�a�r!^Y�Ѣ��]��L�SA���}M>�y����x:����-9NYD�C'Hp��]����s��P�V���>D�=�.��Qa���`Co*��B�y�����>�m����_��C��q���J*d'��P�x6��b�
�ڄ�zl�<�B�����R �R.����&*e,Yf��3#�
��`q��ڴ+�e���W�?L#���w���Fn7�
T߆�%	�á����Sr��yM��O8Z>�<��Q�(+��(>�7X@K�6I�ΤfE� G��x5��-��R��n�Q�|�,aJ?����Ir�6A�AxSz^R=�U*\����V�_j'�D?X���Dj����ax�w�3���<̘�$��7��)J�U�=,l���'��{�F�<�o��oܳ@�2��࿇_���@��Q�\E�ٗU6��LO��n8[Pd����̧�%X����MFDl~l"��Uǚ�^��C�,�Q��=$�2�w�s���O��.sԉ�<��;x��c1��[�R��V���_���k���5�3ZǉӤ۲��"�{�!�.��,%�C��~W���GC%�X	�8N�@����){�/��k �K�s˾��{4�kIu�ea���~�n��nC��S)#s!y-)}��d����J��b�+�
C[#Jcw]
��u�:�{�z��-�����O}Ll�ExP7uR��	1b�9��X(�����:�_�i�r�L�������s�la�B�
���U��A��]*_�Y�Τ��~�:��6,�k�4�Y��{��9P���t�-�v^a��<�W|�fӹ�"߬U� DŨM��W@���H���(�e=�w�k1R�}*�����ƿV!Y�z�wGsb�=�w��7�$�."�;XE0Kg#1R�P!���)
э*B	��>�e���[T	"�k���m	�I��%'P�s�-�\[���ȕ�{�*Ʌ)�!8�49��9^�� ���Ops���y4���8˝�OJ�$sy7�b�΄\���Á^�G"����wA}�AA�I-�>^�tjTR,��M�i�(��X���g�(%�Pzo�
[��K\D}]*�� V���$c�BT4P��&����BS�m����&0�<b����妧F��^1�9�w��u�����Y���5�¢�j9��Ta��������p� vlr4�'PO��������[2ե'�~�Ԃj�H�˦.Q;2�����ƫh=�QywX�}$eqK��I<B؞�G�O�ʉR
��8}�E^��ZC�Zc+�ӯ����{")ҭI���z��BK��/�Xm�z�O���Cqa�*��0���p��#����Ǉ�B<)��YM��RYeS�C$��4�sy����	;T�"���;aX�WgK}�w�����O�˖�bsʉ���W#�{R����թN+�����jt[B����;��T�NT�KM4��9��)�ď���.:���Tk%��g��h|����Ҵ�G�����e��[�x���i~  �DQ�1nG7z)~��_�x�F�������U/��I���z�� t�~�׾먓|��0�i��� u6�6�z���Ey�r.�uMF��#c�U����tZȎ�Ni���"r��S2��W�/[\�n(�Õ�B8��+�S�g��y$�p�GF@��K�΍d���KA��J�����|��yy��/�P�	��H���!U��c�0]�3E���f�0�M���E�P��,I�>�#6eRql<)&-�q�i "��l6Ŧp�(z~O#e�MC��vd4yˏ9	Xh�{�FШ4W)>�B����5�~�6���V�DX���D�'跟U��V�#x��,�&�󀿻U���Y�h鉾U�ʧ�v�=����{���D�)ق N��U�R�"���%v���㯀]S?�wA��t�AFi�h����J�cj�(�B_^j��k��y���Z�t4,h:��e� &��KY&xS.�We�,����,��M\����tV��j-�k7�Jy�`������Y�#ǧ�h�N������W����tC�b�F��e������Y6_�?��(|�W��vn11��, (fhe�!'20`3k�9�M�7D7�1̏�(5P\��
q�er�(+�(f��u˶�7�.�P�p"�q����8��a&���D<��Y�j_T\��i�����WZ�dF���w9�.�\�<�����T��������D��C�k<9ᶯ��3�%�?b�j\�i4�\7��v!���ھ�&�Pl۟E.|��Z	��ۓ��0�0Q,Z	����.�dg��s�Td+���?�;�T���`����'d����H���S�X��c��b�ޣ�V[obR3IM�R�:���l�4<wάy[�6a�ʩ㎐�`�:�y_]��V��K�҂O�>�K�Ϛe��s.s�,�,l��u��������|�mhr���Dz��Xх�g�D�ϴ�Kg�Ǟ^�7�4ј����T��μ�9�F��'r�`�e�o���-j�$ʑ��V��B�5?�v���כL���}丏����F5_�����	�x�����	ޙ$�`V�?�ڱTP�|���&T��+�������Y�������o�v)�[��tb~�X�����U����	�	o��ke$$�"0mnM�7ڜ����+z�K�+_N-�w��-¿�;j����&b����n\qfCS��� k���w��R%��]��	7z�|���"P��W����~�7[���D7U��8F����T�N���\)ò�g��a{�]7w�L�����Ն����1x����%�= L������붞�iƋ���.0J�m�o��uW��S��&�Mn�/K2��x�sW�#�)u�Gh���[X�Ǆ��8���j-���@/��e�k�,��Z�v��8~\S�h�-
TS��5R�%��z�B_��x�H�rߨ^瀁����W�3�ҖX8��$9�:�� 	��haӟ�#�.��knsK��Ꙕ��ڥ���	m����������'�qg�����z�	)N�UP�yH���'�#x��1�� �ņ	���@lI�ZΈ�>��a#N��1!5N���I7�/5���%(^~�u�5VqL^j� *�"�>!򙃶ސ�Ƕ�<d��et��2�k�R�� >�-������$�|��1%��^#魔U����m��¯��&���=VI��<5�*.5ݨ��T���56�>����_rq}c��E�T.��@+$%�1��3r�KP���אL�+�	SI,�*>�EͶr�ك.3ZozPH��q�\!��OKN��j�&heŔ�Ȑ$�U�Ӯ�s��[����T��ckqڱ�JհF�2|�l|��q���cm�r��TcwuF�[1��aƄn*�/�<�9i��t�0ג�/^�H�����D��L��1&��S'��*�-�`rĢ��낭��y�)�ٚ�Ѱ�~T���E�:f���D-ށh4/�g�� C�h!������f%S֙8�a�Ta�%���ԾP)�0�a�[i���+�A����?��kb,5^��,ҫ���Z(�Yf��{5��R��U�U��4_d�O�RtK��7$�Q�a8����(����i�?�&�����(��a��T�������d��,o��0$��㶟��ư�,O����z%����g��ęC09�Hi���Lߑ�	y�ɜSD���O t��vgw��L�[�늑4�4��N�j�5ۃW�aW�W� �#!M��x�ȠnZ]..�͢�?�C쥱P���ʌᖎ�4�ȥ8E���p���[�wdB�P�<���E�q�j���_��Q��F�I�mB�V�>�2���8�˱�@]�K��o���n����H�:�ZX��+4x��]E���Fie�x��ᴎ�X� $o�Ā�N'JC�C�@�cQ���4w	�.�d jV�X ��s�^G����=UM��ݽf�&�;]F�}�_��և�p݅$9��&V��x����#OS�'��"i )�K'�)�T�A��F��ӍfZ�B���I�1܀a&-0�����?i�{d�LDt���F}(�S]�r�9Q
��5d�0�-������6�����[t�5��<��eۭAK}Kɘ�'#	�]�������.=痕���!�_��^�p��]n��<5�j�i�a�����ʬH�`O��Z��T�U��5�Q�@�%!*��OVSR���G�++>a�1{?@U��3�T0�8MT��K��y�#&9"O=WW-�*���zb��A8������3�Ctm�%:"�!��x�O��:���t� `�7t���j֙�zVO�&��+M��<H�]0E�wR���LHf򘂤�����I��^l*i���]ou�6�[�)���tV��1�U�v6��d�ʨ��R��_a����PN��d�fG{B�j���{�(¢z��$Q�V|r������[đ�d"A%;������WV^�S��xc.�=����#Y,����p�p^���q�c�N$�m9ɦ�rD�� z�	�1o�������Ҡ������m��?>p�Wdp��Ah��Ԧ\BPl!�)[Hy�~Bњ{��Ʀ��5q��/Y�U������7nni��cwPIN��e��F�\���־�f��g���x���K���&8���ᢞ��_l}����3��>�Q��t4�ɯ��@W���oN#�ǲm�͛��!l������mi 8]u{>آ1����l��X!d�m��!�d�@'>q1\�x�6d��I�hMm��՘^�Mk�j/���̮e��g�e]���ڭ`�|;�0>����WJ�����*���n�S�#U|�^����%\�C�� �X�e� ��N�Y�,rͰ��'��AlWN�"S9�j������8���/��CM{vN&��xg/7ô�ϹVP����GǛ�
�9&�0���J1����kq����Kܬ%�ئ�g����m��Vj�D��Q�E�%�G�Ћx����� q��a�~t(֒`j�V�}�Ł؜���s����h��9�ɚ-�4��0����&o�,���-���ֱWP{q|}ȏO�prB2�� ��k.bx(���ꮖ/Q���5��9��zz�@��|:ڥ�s��cߩ�K�议����;+u٩J{���
g9�J%��Hk�A�.�
iӜ�ql�{!(_T����愠�����Jl0:+�x:G��T~T�����K���E1�<�l�o����FQ�<܈�8*q3�{Q��G��+o�H�Ϥ����,#	��(�4�*��U����"��'�^@Ǜ_��2�#�}&�8)!+��~��'ʐKҵ�[���U��#;}�|�̆6��Z��xףk���H�^����oGp��ӫ�&Y ��&�=�oq��E�h��87- ����W	PC0����Y�����B�db�aO�uI�6A.(�}�Xt
w��?"1�	�GW\B}��W�nM��^��8�U#���c��1�N�Rh��W q�u��)�������[4�Nc�y�������X���N�ӥ�VI4Ҳ|L�`h/ ]�@u�B�"b���zǀ񼣡����"$�/�7'�24Rj0��%苊����g�\��}�D$�a��Ss�q��kg"U���D�<2(*����7�9o׎�gn�cӗf��)D\���������pv>�L~�9����qo$��co�i�Àu{{��٫�E��:�a�_����_u��I�H|-$Q D������Φ������]9��6N�%b�`�Jl�ŵ��fRU�Mg}s�N�Vh�$�欱Lt�c@k����U�p=!ĸW�2��q`n����z���Xh� 2#g|�7uƖ�3�b��!)ut��l~Hnr�h���ah��C�W*���c]F��G,?~���k�o����w1wHbVlt����.�x̣�����i��N
t�!�oyvPu�7�:��6(����k/�>n�pA+_�rjB6�(tܱ7�O��לV�2A�F,�9*"HvB�z��n�{Hb���,��w���K���ʇ���W��'~��̌�>h�U�w�C��
��]~�$��}��D�3�j�=���d��x�,�i�����,��ng��J[O1�ȰvG`�}�G��%���sU,47Nj��	�v�x�v�P[<�Nأ�.D�1k�M�*FBkAZ2߲��6�/�_�k����/
�	�s��h?F��7�e�mJ���-�1`���=��3 �}Ĭ��M<� %���JRƋ���nS1�L^�x�浛�]ܧ�%0N|m�?�yNu�4�@I!�Q��j5Y~�&.�����]���/��O}�#���?�G'�Z^V�8y�f��.39����:n��$ETT��7iJ�dT���3�0]<���;0f��M�3��|���##�Ph$�mTC�ݴ�9?#��}$������.rhlt5��q��9u����*2.F/�����H6)��9���%��c��A��h��Q<G7��SO�~�A��gr)��xGl���;b�Fi�H�q�FN�~}�1��z�ɀ�w��EYK�ȋ�NZ���E?��Z�\+m���R��̂M#����`�ՒU��-�n��,˯��+����+ ��2�Ep,�wt={m3ـ�$��G���΁���_E_.�o�>��v�*"���rm��������!nx-�ɇ�&Ht\��ÙTg��g�U��E:�fz��!G�a���Ͽ"AA�����ė���4�_P��ݭ�9�G	\P���/z�5�hes���%tߴv�½��=�,r�ɳ�.���'h,E�1w3��Pק,��V��/{�?���E�p�}ՅJ���1��G�ʫ$�~JR�E0?�\&j�`ZТ��3j�%��x�����g5ȕFB��f��,�#�0�J�+����.S\��s~Z�>W"i��/��Yӧ��1mi��<�Ϋ���!`�z�CϬ��3�� x1�В�����c�}�����S��zskoV�����L�s�e���c}t^/��czm_�#r������.ԝ콵�O��1��Jf�J�E`vݠ��/�T˩V�E����*g��bʮ03d���`���_���;�"�1���z{�U��4k|8Hw�'t����DҶ�Fᥢ��E�H�EA�����z���l��zT�N��}C�{�^�d���7Sř9�7΁J�,��8��l�qy� ��E�!��Q��/�@\0�~�)*�'�����GV$6^��BQ�,Xk���S#2���ϧ�ڽ;4���3����k����K��=�
����	�fe�P��1��N��9��G�4\���BWP��*��ԉ����6�����`��dǄ��ipj��X� 0���c�>0y<ja	*�r�?;�>Y$7N�움Z���P�k��k)r��a�o��-7�ob)�C� ��>���um�����X8��}�ڏ&��Pf<�$ϟ�PE>ʡF�jN�c�A��a��ػS�O� }���W�r�`� .Z��<���Ć�z�Ē�Rc�ڗh4%���G�ٞ�h[�;�M�4���������	��n�?SMR�`�gh�l��?`-��ewGp�5�O���0�vP+[nH3l�kyh"�׸��G��WF���~R�^�s �(�$���^y��&����O��G���h��Q�os=[Q�����U��:{�K�wY��p�R1��ZJ���̶U ��=����bs_��uk�E�Mc�
�(���nr�옆S�qaέ��ڮ�*
橏"p��5��n`�2�Z�J�Z��R�a'�E);b�V��DP��.%�\�'k l����pc����ZT~c����4Uj����'k�2w&���ܗg�_�·�yơ˘C�G���u����	uH�spg��p�x��s<���9gW�_`�$�dpۛ[�J�����ׯ)�䀺�i�|�d'�j�,��������Q�j�i�C�S�ļ��M�%ڻ:jZc�jW5`|�.��|�d$����gy~�%�U�<��(W����!]�`����%�۹��	�b�c�y�V)�@_j��!W��ٵѣ���$s�{�(�� * ��������Y�!�x��;�3���U+��R��hk��>���n�W�3�"��ѹx�� (��ۘ$6A�L+�
]5�R��A`|<��uz�t���kYMb��
�;��4R���y�ȟ`H��XNK��]�F`��i��Q*S�tJv0rx�z퇋Ӳ�j�j�a�tzYKHYW�vj㙬��,E�N����.�Y�n���V����V�3�ؗ2���ĥj��2����%�p���Z���⽲�~1:��ɺ�P?�����qAJ�7�]͊m����/��M����=�O��͌���nl�ͩ&�[����p춏@h��n�#h�:=+F�o�k��c��L����+�Eq�N�2`U������~�VϿ!v�S�)�FZ��E��H���s<y��(�(&|��X~"��l�-�)iTt�첁r��)���m_/J|��
�o:�E��]|��ii|E��N�,d�X�_MJ��X����t� {=��1s�8���I!�%"o�.��jhl�5�����|*J�d�Q�>�6�،��ϵ�s��t?Eݣ�Cv�Somm:=9��g��T��7�CT����#ɡ>�#S�0r<�m�OK��-�	��µ��$g���P����RE��ڀ	h��Y֘�>9��w�ea��4�X��re���헌��J������yh?�K�=Z��Μ��c[����*�"'�k��uK�Xr"WC�Z �ZO�R)1L(Eb �^E�=�)}�}�UGc}|�]�-��BW�?�b��zLb�ZK�U���P\PHw#�=�5���ǎ����8�%��I5r	���h���z&��3��R�[ �<ƇH.�J�C���1�w1)��';����
v���jĨ�O�J�g������y[XO���������/}���ō��l�0=�۔��� �rI��0���b���[�m����6��s���F�Z�1�SF0N�S���v��]�)���х\u�8 Glo��R��H|��%Mܧ������
�2��T=Qt�v�?G�J��p��-By8�����c�p���ђ��z��(Գu�����-[��~ ��֕(u�*��_b�k(�'5�x�n ��~�m��L�>lI=?�㏫�*��ٲ��c���:��\"�e@�K�
�v�t��lQC�ۯ^J�tʦ�0U�+����-ݭ��B��"ڞ��)?̘�q[kN�X�����Bϐ���(,�6(���|�}�Vޞ���O%õu���:|�C+. ���ncJ���ƿև����s{���SM�����D/�XҒ	f9��p�c���\5��2'���� >�nYUz>�'��F�Ɠd���Zn�2��s_Eh %*��`S�H]��N!�Ǥv�;uw<�?+A>h�]F2�a��{��ܴ�|-?U��Ћ�&�'���oR�&[)�/��
	��K����Ț����4�� 2t��\���^���6�����I��o���o��;�A2�^���o��bh��?,MI`|]o�%i��͔[���L~ˣ4Pm���A,�8O|JE��u
�o,��[�Q�-O��r��@g���W�����?��v�U��-z&�&F��j������>o��	uQg�f`��qӰg�3N���P$��_��=F�O�l:�寕����v�$b�����~�Q��d���/ļM萹g~�|h��m�zd��w�l���v,x>����?�[xae;���֚�V��8�hGā��h�c�����.�S*G�h��������w&�|
?y*^����"�. g�W4
a���p�0������ޠ�0�A&5p  ��;���~��g�6�֖�Ay�x9K�`��_5��� 9=�(yU�5����mj1���<���-�[|CZ�Yw�4N\--���+�:`&����z���)�x�$F�V��������{'����@(�����9-g1��b�c��u�@�"���b!o��\�%;B}����qɠi�B+!+W#�-�% s�JY�:2�y!��Z�d�˄��)����,��M��v� W��\�}{Bǯ��`�\�y_����Z�8K�_>�c�� �~��~��JQ�}�S͂K�r���/�ZDQ�{�s��,��f�Q0Aftb>�hr
Js�`��MlWHo���,�nMOZ�X���#Z�H˗̂u?��ZT8��c8�[Q){�mO�P�F�"m�w�U�����Zq��Ȁ G����l�V߾2	�M@�LP��us��X���G�n/h`�/aU
}(/.�~����Jr~�YW\~D���5ߵi������h͈��D�#c��*%',	Tr9g~	v�Ꞇ�2���D_dHa����>� 9Ϸ�N6$�8��4(���1���^��`E�w38$���DE'+b%^}������t�&�$�W�?+��<(i1Y�\ˋ�T�2�p���ʂE*�rX�L> �y%q�Q�rx��a�Mb:��۷�2��u����IS��s�� �^�a�	 Ft�ظ?���ھJ���T�?��鴵��\5I%1��Kv�i�\������970RAم/Z>J=�Mc=�D�&ٓ}�
t�Mr2���p���1=E�Fl�@���t�J�<��GP������������o�>nK�,�d����T��A�3��!.%��8!8h�{N	VM�H�/rd@���P'0M	��T���\�II_Ĳhnf���e(.{��1��� C7P�+��I�d��5((�5�)٨�[���i�5&��5�%�e6hV9��L�HL��s�4� S�5�Hw5,ܧ#o�F�"��ҿ6\+������>8+8�%��WL�Μ�shgP
'��@�ڭo*a�7=�"^i��p��T�57��S��M��8!+�Ӄ�a�|�EVz&P��HT����gŠ����K�����g]�t@��P������!��&X�ط�㬒4�;/�$�;��C���|WD"��L�:�
�׮�J"t��� �E>�j˄���͠��o!cY��� <��rM\i�̰r0�JE"��~�~��Q�5&�$K~�~+�	8���'n�픗PKC�ɜ��w9�ϯ7�F=ܢ��䩁��V3�2���ZGG���X}u�.��VD`��Ki��xz��2p/t "��a2FT�M�\��#&
����,,_�=3+	Q˜J���h+!�9|�x�VQ��"�q�<�r(�A�9׮n#@�D�^6\E�LpXG�,X�:��@<�<�[��^�28��X�0�}�|�S�$	/�K!�M�љV5��Z|�q��>N��<`7.��o���b@��ߏ��^ ��q��.&6��55�͙�Ԡ�|Nifj�]��?僗d9�¹�unc�b�$2�a����1�Gw`�Gc6z�kT��@�dW���^oM�tWk��$�iY�r�'nZ�x~���'�Z��b��=��P�d9>{�[9�Jx���$��C�I��E|zK��Y}��z;mMk�����_rtR����q�,2�;��HN���{Af4�-���Y퇈�ښLB@j:�v;�S�/�7���k����7�{��/��&����=5��O���i-\�(Ǔ�`����>7��H\�'���σ�mR�)��l]�{����C��J���������ox+������o�yf�S;�^$�>n�Jm�q`^\%;c�< ������ck�W����!$~0�~�?��vvΘ��K:U%�
�
M�����>�)�V���v/�����"��Y/o�������6i�����_Ώ���Qϳ�W�Ӂk������V�ROcNY2��VM�~��u��^?t�}�������x��L�X-)y~{q�T���#E��Hubq�z�Xf��.�ͳ?�J�'Nl5��,�e���`��s�Q���{����h=	�mѿn-�X�V�6{<Q����)����N�g�l$q'�Ķl~��M��v� G
��A.���'���G ��F�I�Q�W���ކND@�3x�ccy`�0�Ky���xU�Pb�|��i�/%�]8��m?ĜZ�G=�A������&�\c��!�&g�G=떋���jLU�_�W�6VND�W	��]�,�� ��W�)/���
H��7Im����*x穚�{X���!`�"�g��3�,��Ig�\�^�g�[��!%b����m,J�V�a}�w��b<�,�]�@>8���`��p�,�ߎ;	';��j�;:��f��V��1A7)jDl�k����L뻶�
9�]�K5N�����T/创���G�QeRu4i�!Z���wu��Xb���:�F�A9&��u��5a���%lY��}�i)�o�^
�R��/fvGG�O�`pK.�=�-B�%�<2Ió��	�lH>��5�@֧I��e���)F+y��w��á�f8�3�TWICWNmW2Q|����4t���?�$��s�տQ�c�<��#����;K����%$�H����x����s0l�3�Zp����������¹[=�I݃��҃�pڠ��U��ޖ)�q�{��v�eύ�3�@أ�">w�jgb�7�-��ʰ�jg��_-���?�0=K�y8$���֕Y?�{��q"��k�W��8r����7��gdOI�� �����#W�=[�����drn"�$��#Օmvt�P��}���:q�)ł뎌��2j��Z��"M�Ay���	���k�E�g0T�7��B�&��p�^�����2��F��n=bآ���m���:�Y���9���9�׶(�4���9.{_qǈ3 7�$ &����}�gXoUHuw�+�T���0�E���Ǣ�d���Nx��m�){X�Ĺb��\l'��m���`}1����XY�W�������Ȥ?�6V��C���7ؕZ	v�[)�]A�5T&�uu�DI&qx���v��5�+?	��q����?�u�X�5K#�K�+->�z� �AF��N����nEXx���2�ӡ�ǡ��Y,�J��K��a�v/��DN�Pw�#�ǝ2�݅�Z�UF��Q�����]��d[G���5�{�u�C�y�V��V��U�ƽ"s�糎�X<�~�V8"����?3���e�[|��'L�q!�=��Cb�Z�)u:���WA��3^��	g�եl>c��hl#y&���,7:6]�G���ԏ͡�4H�y��ͩ���4�ɛ��Ȥ�Ȳ���հ��a�N������۱�]Т6'��U�����qU��1�������?�'M�v�Q�8u	��zN=�%�"Pm��U/7L,�c�?��Ls�ϳ�����z´����S�/?��"����k/զgoh&4;X/�;�w���քgN���Úd�V	g<�M�-��ǵl�c�j�\���Z<���6V�D�yJ ��1�6>��݀��e�7c^���׻idm"O����7K[��!|��V1K��c�z@�8�~	���L��`Ţ�X�ը]��x�NH,�ٗ�1�j/sRX��Bhd��/}��s	�3����b���JT0&c�?����p�į�3�X��h�q�X|�l���ݮ�jIr �]��M��&��Dֽ�o�(�KO��s��4���G�iϊ�q�ar��������A�jѐ���Zq���Z �m%q���]M$���Gu�IPǉ+�i�փ9Vp�>S�Km~I�y�h�(lD\,�Re�8F���m����Hhh��;��]�yq'�'֭�Sh�B�JZ|{�H�����fQu ��6�I ~���ӑ�饺t��y<f7f�YS� �C|��(��ȉ�h�ɮl����]bC�����ӘHM�LX���v�Wvvw��⒐oݶ+1G�ïTF���jlYiKYa�6<N���3�K��5$�I�O�V)������F��tZ�݌͎�2�)w��=������(ZԐCG����b�X��	�w��+��+��._4)�躏�i�.�jV�[�P��oE�t��3�;?�5VQ6	�� ���c�7����j�	3",�����pRʵI��1a$R�{|�nԒr���ݰ�J���?6�/=�0��z��	�L]@���V3S��2)��V�B�����}� �~��A�Yw�Έo��.dy�s�gJH�}��iy��N�g���c��׻�+�@��g�)6������`p�-Z;Ϸ뛫q�4�!��[y�'a]�t��O���~�J����58�l���44L��̔��ht|~+R`y���d�f��{��CI*����|�N���H[�Z��E�L�VO��җ�u����ϙ�P�������P����5��EN�Z(!���2�2J��̷�`�a�C����4�>��)�AwsW,��m��	����(^sJw��}4�c�,���W�V����l�	��]Z�������G(�_�|#�n�U�B�S�oNC�%3�ă�Ϳ�`�ބ�R!<iރ&�xAՇ��s*m�r�d��v(�EJrd%�����ag|y�'eQI��ڐ�i*`س���Q��Lq^E��� ��w���T��]��#;`91������M�l�E�8�|��h8U���o�ָ0!W��A$�z;Z���^��%�Lל�Gg�4�Z�!��9��'�t�sʗ��'>�<�C3��np�Uf M�M�y�U)pvM��X�#��jP�o���W ��5?�m��p��s�c���al�5T�{���� ��A�mu��K�0���
���wroܶ�2���m����A>[�݈ym��O"�T�]f�<5��n�U�դ����r���˙��H?����5o��N�'��i��V?��IB�ڤ-��|ْ���z��k�Ǵ�M��t��1G$	�a!�u7�;�k�l$-�y2S��`�:�*�D���(%�W�p�v}O�,��#��s�H	~A�-���>y�/=TV��$	�4�I6\|_@y�[`���`J�1H�����k�������xse���D,=<�Q4��=/PgK(&���HP�>�<�Z�ᝉ���u~�~	�~���o8!י g�T��ė}��x7��x�h^��n�����=���-�>���"ϛ���q��������yNN�0�J�Ri���BCzA��Cv��1�������������^��|�^�y����t<�kԙ�I���4GF��d^�mfᶇ������O��0mw����-�`�����(<\�����ryrn&�=�kf��TSc���Y|�"	v�g��MZ�Pa������R�vY���ǈG�i�����Ǟ�hR��|S^,m�+� *�!ʂеX�g���E�W�x��y�Ӱ�)Y]���J�@Y�B� ZE����Iz���5uˬ�0!;Qf>�������\&�\����fT�:���.a�kBp(k�oz����yr�Mf]Z��ب/�B����AY�Fd�*P���'>��>d���֨A�v��(SXQ
��l���ֲ��X�R��f��iT���^՞EZɈ�H�^:_�kWlm� 3[���Չ�)P�xV�������L��1S*��L�vr'o\��k&�^z¡��r�m�i�K�qY3�jW�IaG�{���"q�2^�.Br��z�٧N<��衰8�;�sNkYH��CZ�q�;&�]���F@�� ̹����b6WQ��"��P!�2QGf];�;ao�&o��j�ab����Y���
BU���O�Iz�D�k� �x9~��tpUT�K���/%|�y��eQ����cJ+Yf�������[Z�/����l:m{&,@`!�_J%�SR*�ɖM��/���hŤ5O����x���U����-I���]�.��z#ō�[��N�D�1c����A[o��Q��-.P��07�f����ƪ`-�[��glB��e �iy��1�T-\X�.������*tB�.f���ɋZ���j�s%Z��g{�함U��Ц=�:Rq䔠�|���nmf(:>�b� %;���	/J��wPJ���D��ob�	�J�T��?�u�uں��t;6�AB�hV���mmC������y���N.��_��O��æ�ܶ&~�NGvU�Γ��9j��·��tt���3�;s���i>�eN���ܠ�f`����t",�$Eq���{�M�
'mR]8��Q���[��{R��k� �rxܣ�)�\[����Й���X�A0��B,������ܝ�����(D���9`�7���3�k�����A�_J-���S�*�<
R,@�Gb��9����XT>�R��I�O�E='k&m(i���Lad��R��w���KI��@E�/����k̸F��ة��옔���x�MCh8!���7u��㟛] �����T|��b�U�4�&b��(���~��	/��Fm6�����P;N�/�c�EkMa,|k�L)��1�=�辚pJ�+Ǭ���$�ʺ`�	�|���a�,����ꐰC��9����ld�h[������O�4ب�� �ƍ���ӦqKG��ݠwЕВ�-������P��i���6��T�ij�r��مx ��]��lb�r=��$��@��?',M:�)��V1�p���0{5?�6i�f`�מ�1Eæy\L7&��z�O�Rd8"���)^�nWM��܉w_8 �;����#`Ln�NT�Y����l7�������.��[wau!�\�^�9�J�,��2�z8L�!���|�J(��c�I-Ne!@(���N�_��۵��mm]/�;�8��б�O("u�~p�/�Y�_�����s��$sR�ƻt�o;J��۽@�iq�U��>�)� �}$'8�	� �5�me���	�=�vg3��z���\A�� _<�����i-}�|
7/�y��eBQ@x�0���N5�E*�Pc�i?T����*����؍�z2E�KdY�pwH��6��DJ�p��:cO�{�5�����Ʉ5����F(kޠ���*��
�l�6�Y�V{��8
:a˔<�V���������U*�<�8��#+ߟUOW�d�з]?N�Wb�!N������t�V+&kzn^k�|���BU�y��̳�(�zOk�t�`0�R��G�S=���qK��h	��F\*�Q2Ы�V��'�Vk�y"�C�\1��!�GTMd{�������N[�?8�l�D3O`�-��_ՙ� �w֯�)ھyhǚ����Kӓ��/�<���ܝ�N�J�<��;�u�����`b�FWj�p_Ƀ��\��qAL�X����[��6a����*Lg{�� <ल�'�]��g�S���M��>�JCQh勞��[V���J��*u`��1���� ���I��@W����[��ܴ��L�I8�����N����i�_�zp�ɴ�\����l:�G�s��^!�oH��:�S��Ŷ~+�:�Z�P�ؑ�x
�R�|��F�_rU��B�Ag���M+|���.�y��\3�o]�u+�yh�;Uot�'1�x�:_S^�42��� r͙�]�4`��6L1Z�;۩�W�*�qu�������X�_�^ǖ��F�d���9�pYh�*z}�����1�O>{b#ai?�j�զEd=
�	�����R���H�c����t�[�3DWJ�Y�b6��]=U��K"t{H��^^�Ӝ2���'� _u~#�7�_(z񍫝�̟�_�o��dz���~Qn�wCh{���x�u��DP�W�Օ�CM��($G��KZ�yZМa?D L����C�&l�6��r^#�&�.���ď�6��KUMo�x�!���,�0���_p4G<�0�����gv�����F�U�0�xaK���D|Z��sPT�{�9����hG�:/R�E!�-F��Ej��t��Ydm�����/�χ�Y��]+�9� �1_��G{6�B����l��B���)Ǘ������P��;y����,�i�79B�%���{#`L�����r�蚵QM&ؾ���E� �V��;�����'�lQ�/��V
NTd�t�0o�H�ս�q*����A�������{�2�u24ěiPBlXՎ�5�ǐ�Ff�y�1�Jyȡ6dbl�$�ɥ|ׂ��ꟊ��C��ao (�eC��H5Ɵ�Qb�f��#<ι���B?���A,~n���Ň�9��<Z�dұX�	Se�$#���ohy����:�i�2+D�m���f�E������$d�U
�_�0�V�F�Oө�O��1�Uo� U�'V�ria�����#���vaҟ�Ι�o@��{���&wC����� ؤ���)?XF}�����n�4�Z�7���'R�5�R�M�~0��bI�*���P=�h����#�X�<��� 1���ҤY^a2�nx#�Y��b'�*� E�V���ʡ�(�A�5�<һ�!��bA��d3zx��}����r%��`W�=��*^^rs�x�h=s\�k:m����P�B�\�쏃3DAJ���|J���;Z�r�/<[ .IL�E1�XG[:��|�O�_������`��l24/��fͳ}U�U�Mz<!B�Q0ͱ|!E�A	����6r��M�Fgt;-f🗇��Z�M�+��_P���{8�D�SˀLL7E�/XNU��h���:�������_AA�>�aN-0��E~�y��b�O3����H8���4�v�橷@L��!�^���Q@ Ȅ��(�� Y�y}8�}�Wx�C-��,���3��2�Fn��l�/֔�E��IiI5�1���eg���](����}= VD �a�z���$�x�P~�����|w�< 1��[�g�:6�)�O�����EnH�K �N�)��5uPan�p�LI�nZ>X�$Cb���H��jC�s�$���S�((˖7��=#���K�>&�9A����0��:�~�l'�aB��:w����X3,�Bx9���h�zn݇�N/�|Ej�B�A;��|�g(WjX뎨��@�ԡ r�V�)R�hN�=|���!59!S��lP�|�.��v�t��8f'�D�?�糚	��"�}d&vA�����5 ��ͨwN�L6�r��ZbH=�0��3�^;?�����hlcBl���n��M�K��Ω>���i�ԸWpG�}�#�P{��A��H��(,>�\xf� *� ����r�,�-��مÙ�΍��v{S��Y{Ϟ��Y's�ܗ�4�A M"�Ł��H��Lڻa����|�P�5��q����V��sUܯ�<O!�{���X3[��PA�`�)���ߪ#o��֞��h�:�p��h��������u�*�'"
����OuT���,@eTB%��2����,���n��?��;�Mw��y�W���ju^B�#ߟU�۰���ر0�[��0�9CYAN�wqǼ�/����mL�[��;��"�R��c<�&g�O�/����\�����*\0�Oxt�z�s>��OS2f]&b��JX!��$:��],�Ht,��w�sJʓh�.a ļΈ���w�0k5�6އ�P"hqu7>�Qje�c�ft�=�Q�f�:��{�~]J���&�4.i�'�����B�H���=��wLT#�5RW�����'�md�W����ļ��"RAͯ��ÅyS�	�}0��P����s�+;g�~���ٵ%h�8i��8��3�i;�H�}`Q&���'��B/�5�Gy^F����
��4��X��C�
�N�68s�aӂ�X6�{W���*�#y���ԥ��@��ZDS�P~8��A	� l�J�]�2�a��]�ܼ,���Ex	��P����͐��8�h�N+����{�P=��rCO6���4l	(��x��;�B��`�6_�Zw��s���#�M7R{����K��Bð�k~���a%���Z�FՉO�ݾ:��R���?tEI��Oĸ�[���𞭺r'xʇ���3�g���K���8O�Ά�)�'���
��Is��͕5�Ud
z��M���P�1NV^��D�v����?B� ��v�������3�lB�����r�w0�`�F�����tD��Oj�C'��	!v�s�����f���2�,����9��A�Z\�s��1�.X�����};�7�_^�z�]���x�A�P���TZLW��&�ؗ�$ߜ��b��!i�5(\>��MͮgC|�0�T!�v3]�F-D�L���C2ɻ������r��<\����l�i#�Y4+7'����vކ	��r����'��Q�B���A����mZ'
4#�L��u�c@�ƉE֒�y�JY2�X�^�r���J��h��M��ڻ�tɏr/�W�x��wU�$�Ao�ό��*(x��uߋ��p����� U��I}��f�O��bl#�߄�/
��D$=�e�s3*���W�_LsU)�O:d��]�9��h��L'�a�"Qni�g7�p�G��\�lpr~y�=�Di8�����b	�l*d���,:v��8	�8~��M�E�z���ij;J����߸-H�U�)���&�Q4߶)9����i�>���o��C@ܫ�RLDZ�Qp���O���Yk�`��9n�`֖z*,����m���A��:�*՜oOD㽖V^S/�JrB�!���~� �)�1���EQ�oqDm��w5���
S�XË� �u�Ysz���P,��![�gW�F��j1F����F�ǆ�z}�B�'|��Rm��E��7��\���W��쵌`߾3��)�k�������&��q,�j����-a��}q�t跶o��}nm�ڱ��{�r����]�X6��ۮ�H3��D�wa(����
p(��%�&�N�?5d��IZB������ݖƯ���"����9Be2�.!�Nf�TE�����4.X�8ܘ���rJA���b�7.R�\���N:b�|ЦP�#�VY�#o��$�K�V�j�ܯ�ZS������y�������`R��jNu��a�@;w�^I=�pW׽�n�Bo�3MF��L����Rܜ��e�*.�,&Ip�lr8J2���䓁·,�NH8�iP%!K���s�6�^Z��d����躖��h�l�J�^��W���O�8�Ne1B���Gu4�T6+�4ݥZ�Gxw��Xd�0���Gu����l�pR�GjO��DZZ~,|yG�� p��bW��匡
N!�Cb�� 4Ӈ͟�LZW��h��2{���yO�r�(�D�$�id$W�X=�2���|��H�$g!���� \���%,E�8rO��-ԚVk��Z�O6fT��n�2�Դ��g �.qm�k9<t�	u���e�9}$�X�68�����!S,�4�H��'���(�����VY���Z2��w'�[ҋp��pC+���Ŧ�t��(,�N�	�_>�+�����i�e�>��c��ѯ�-o[�׉=���Ũ���b�4�����'a�U[���UYU���^�}n��FIL�e�~TӀ��7����v�/!��СxgCa���2�;�rr�<}5��Ӹ����rY�j���p��V�o�1<b&����Z��%]}cI��x��P�)_���۳z�����9�������;�7ʘ���]_`�E�z(K!8w\����N����W��G$ͻ�z֚��	U�j5��Qnِ��R��n֘&�Ph8���Pd�B<�y(��4=�<s�f�R�8�p^��^WS��AK�ٗ@�	QXF0�/��pl����.[3�y��f-�X]ؙǌ�l]�������*�>�uRZXVjF��1�lM}�^�d����]c!J7i�Fg�Qz�w�g�eq�wwT�?�l�Y@G_o|�<-�Y��@��s��=͸�aSv�O�\��;�4=����k:m<�jt�!l` |���K}dYaӲ�q�1��W���-H�ڠ2$3O���t�s �ٿ�b�����/����������� В&Y�Q�N{9?_fu֫ EH_��0Hg����(�����<�G���Y��w��]@�_�J��7�q?2^�Z�<m?���!�J�k0�S���pc�X��Ia�%����zbƴ����Ҁ&����7]<`�����R�����I��ց�y�k!�F��5�譢^�[����� :buQ�2�pl����t��~͍��+�q��=/�@B�q��k������S>�(�HTc�l8N���t,b���L�r�YE�o^��|�J!��3�b���-E��J���<�s���P����F�O���ioa^�������g��{��炼��>!�j��c�#��s�R�u���H����q�t�=����n$=��}C��G��^�c�<{�O�<�a>�q�:�hw;mU�RG�R�KǬ5b5��e��eg����H`a�v��}�]��1x&F�53���x��="�h���������i���uU�ܕ�6��E7��S5�,���������-�G������EV���/�H��U#�z������$��w�:VO��,xZ���.܆��g'p@8Ni8�؁/��L��N���N%�*2MR��x®��P�?-)�()�cΗ$�Ý�R�G1��[ʠbę>�%1Kʢ�Gq�^РC,��u)�S�6�^��Bhiq���&R��\��W����u�A����"�1�:`�oR��yp��Ӿ`�O.V+un8X٭o8��Z��+����Y�Uw�&ug'������5�k ���-����X�%j^I��s���s�<Z)�~3_#<qk�T�x��ɉhs�Ğ�=ܞ\�}YF��Sv�n� Ի�maX��W j�'aˠ��`� r�_��l�ѧ8Q�"�$�g�V3���ɇ�a@��?퓽�>�;Œ0�p	��j���cM,���.�
RJ�RJ)N�>x�`���7,@]���{Z4���Pʅ7��n�|�#/�G��z{��M��>ȱ@>��}��7�쾊�i$�}�SB�p����7�T:�F�s����$�fĄy��JH-y#4�N)�Z��'	פ�6����dO�1�6]�/y�l%�6"0�����1���Zy�)f��
�b-!�g�9��lDʼq�.���ʕ��;��<��.ٯ}�?_�@����"��z�?�hX�ob�k�Hlz�p3q�%\єqg�
|Df	��	Y�j�&�D�m�4l{����@�$9���<��b %y�x����TgEɫC����"�R�����F��Çn������q����0�'}�a�����n��G��;#M�co�+��׶+�S�B&��2��gn����N~\r�[��HS���a�-��0,�ȉ��4�;��q�g��	�N־���$D�����b�Fa8 3�I���	�����? �9~���}V��4T����V@�\`�9�]�/&�� ����|��YU0{�)���/��!ZM�-܂ӳ$x��Ò,����7��+�u8�B���sI��>�i�1:�����[
MJx\�����P?��k<.{;j��V���S��}X�0XJ�$�N���V�R?&����ܶF�&bɐ�^�U�a����	����|�J�=��p&w�R�/��������f�0����v?�gOi�6�1|��뛫KT5��g,���odJ�:�Ԅ�&��~Cˠfӡ��TW+0h�9���w�؏�D�o7~/�V��}]��_�Nv�͡G��VP�����q���s, �!���b!�k����ĥn]����r�"���B'�2��z^��;Xmc�1�=�����=�j?� ^�0���\���?传Ѭ:�/���v���D+��'G�H�,%�;�;���xE�����%
����J�p�d%��Z�ø�yv\IH��r#��1���]�%@M��Qs���sRȥ�|I[��F����*��:&%驩م�r��6� �oHb�7q�Y=�K��9sWx�4P�"Ҧ��r|]KV���(6����ms��{uÌ۲��ހH�e�?K��&�j����"�u�d+�<c�>g@�S���h����B?��A_�0��g��aؠ�t��8�m����?�QT�\;�/5��s�}>���my�0�A����s�_��^�NƦ6eP�>�v�߂J��]�*]���PT�����=�K�ᬒ���IG��l5�f)ؑ���|�$�E�c��#�և4�mO�_�$�:
�d'a�+�B Eo"��+�����I�$)��n�i�c����?��=�"��]�������b�c��H�RVsRC��<m�O�= ��B��j:�<E�6�9:�A-�
����Kw����JM�a/��C����I�	(�-0�DBB�H@���!�XbS�Qț����ӝ����7t�ē���*G/��%QUr_��)��N�j���Vn}#����$'������R���	��Ƈ��u	H��z�DhYd;�ΓnFjݲ����q����~��{�Z	�up�*��dI�����ok��L~��â���h�������K��ɧMz]�.9��ȋl����?3�/En�E��t�:J�����Ϯ-��ΰ�`���,.gj�T�ڐ�S����'{W��vA�b�.�{9����W���=�2"�?SZ�A�OJ��:��J�/,	}}�X��i�s���4\,8����p�Qg�k�U�qS,�#}-N-l�`�.�1��\Ӗ��;GF7���U�U����Y�rY&<	e�H�8�F���D	@u��lq�&�2�*�F�Ě��Kt%�^���F�GP[nƕ�H#q�GZ�Z���-�,��K`%������N�3�Nj]��7�3��I�8D& -�����^��o���Xk� 5�e��y�wԈ(ɹ�\�]���
��I��c(
��<S��<7w���%�n�>P�p&@�����=;�G������gԀ�F��U�F���W���4���Oؕ�\��|�ͥ(H*B��m�M��|�(�|,�9�v�dɁ���!������e��=���0�P��z�4��t�섈�l��"��~�Ͼ۫���5^��T��ٮZ�.I���':�-�R��BC)��4��8�v�A�������ϰJȠq1M�u����#9�&�؋8.��4�^������`5�ޒ�sO�>c����J*X�$��]?��N7e�O��VR��9r �̶��W2 śC����+N����ߵ�?yfX� Q���oAn=|
J7M��B����5n�2c����;���6 gc�3)Em�]"V��^l��L�:�=��drנ0p���i���6�:�ä�V1IE�e=z���&}�>�~��xw�>B _X-���>��xK�jp�2�RG8J�Ā�
Na<�}� D����EU���Č�? �A�ywv�K����D���T��yk^OC�]�>I�����]�l�^��� �;�()��9���Ƨ,��|�>�-hf����M���,|
47[�e���.r.1�Z��d�֖*���u^6���}��a��o�%
��X�s1U���}K>��J����AJ02_h�~�膝ip�\֩�U��4���/Ѝ�>n�CyM�<��i3;�K�'� �����5��Qn�̴�E����@�I��Y�/��,!��2�f�LBr5
�(�F_���S�z�T;x�3��U; M�|��9���C�ws��LpD�Rv���ϣj��ɖ`i�eŗ���[mo��^��'|�͂9�^��'��^�9b�4�?�W�%0�^/m�P��2�a(��gs &c�)�)=�ܙ+>gF�ʬ3��FEcI�4\45��9�jUZd�ǥ���}��}�!#��_�W���T+tLQ�b�,���O�����.��e�~]��&6�����x&�w>_���;\&�=�����B9��I
�06��� T������8�j��c����CH��y.��`P�i��E��1J����2$�F� ��T#ǟv6�'���ˀP=��oOe�E%�Y�PkY�nR-�E��K���k/�I�Ԃ�"��n�xVDpT��������ˆ���R�G|�P�6o��ɣ�xc��Q�3��+��_�AVr� �5������T��6����Kp&�b(6D�8C.�}+����X2⮅�îE���x��Ls�n!���up�t��i�@'�;�a�?fј�����u�Tas����#��!�x�������� ���uԙi���/i$V�V߰S���-�1w�����h�^b��$�pv�V���o��<��a�)b-�ˤ��ޜU��߂�f�z;�?���6�+�mی�ԇ�ap�Ko��#w�S��|��߇���`��\q ؂=ײ2q����x`�>
(�)��.z��_r𕿓��A�-&� �R.� ����l�~"�V�OoH�K���GY�8)��?��/�壓�|`ֺ�(�j��\/>[K�o��"�sz_U1�-�PӘ:���w$EB��a1f@*�'���S�����w��ȸn�?�,���WbQ|����r�y?��	>���K��� �r�v��$2�����`���
4����:1��*x.�D%0�j���јŋ�J����cI��pHYw���7����}G;�p�����|��Z+X������;��?�)
`ZT���!�I5D5��g�ҽ9�-]:E<���R��R��Ρ+����h�.ː������d��޽`v�(����3J
�����'G�>]!�����ζcN��㪒Z���<��j��NYo�iC����AB�4�h\��}sqp�g��
� ~��6�dX"���"D�
�h�L�/Zs{��y�^t·���6�d,q�낸����p6�E�P��07�z�,�R.r���(\h�ݎ���nN|�����z�2��;��:m��z$�5-)��F;�X&�$��Cw=�9.'ch�x/�ו��T�\�%t7}��*>ɳ���w,�p -!H,����Z:���i�?��G�X�M� ñ��p�R��tu茣��W&�of�ge�B&�d������
�f8��U&I4kyx#{*���Q������m\C1�V(U��<�\��n+��������oف�Y�u��2�7�u�d��v��e��3��h��b�����>.���I}��MP}4Vw7����<%��YJ�ph�t *
M�s xpF���c'_���e�e�N)���.,�.�`�MpF��hwE�����|o���`*�!Ȳe4$�ޚY�7�onxk1h ����-3��':�u~�욹�V�eJ���G宼�N\yA�nD�剐����/Ufʴlu	��5�~�'p�����}�l�����k�	�8��Un <a�т�720jJ�p��}�^���|�D���-w$T$��$��T�9���W!��s@�B�KW�S�E��J�n�F�mA��k��
�	\9�\���0�c+�'Qx�WV��-z2�����z�˭y��ڛH�,��٘��z�0)���L�[ 
�(�҆b���u��9�(5�	�RvE^���� 1���by���_�-pH������n��r1��*��a^�km#�u��j��E�Ӑ�%�^c}k�mKb$�����:��k�N:_ma\��%$8.N0H�>��!���p�iH�l�vi�`��,�ò���u����A����~���?�y5�YՌi~��q�I�"<i(գ�L3�cv!�~�2|]��U�kْA$���Q���UM`GC��j�Q8�EKz��܃���K��YrG���Q��|YF}�����̭C2ԑIѸ�F���$y^��f�����P��H/X\մ��O�:�Q�Vg��c'��2oW�-:��~{Z�QhLh��H??�KP>s�h��U۵9C"�X�u���[;(���4+���漶mI�;�0��@/��?����-sx�� >B��C��<�}uh&M㹻h.݂������U�5_�����c�!��5=�,�V���A3��,m�{!�[j�����	|-�ُ@���jkǻ��^������OK!Ezc�&�Hlæ��d徺���7�P�{�h��|��a�V�̡BN�'O�r��K�?��fmI�^��oA�]��{6���-��y Z��E��{SU'�D� ]����l�bb�m ����<���nw�)�'Ş��}���NmO�a�ɀO��!�h5K��شC��XXNX\6�{e���mW���q��f��7�'kN>A���[٥��t�j(~�[���r���o�$���mU�T�e�01�<������3��e��8�y[fArk]^�N�F�}�;ϩ����ڄD%��ȑ _���I�T�i�E�^~���?c.�s������P+n`ϫ{����kF�O��pf���a2Ẕ����B]*|f:l����a���`��e5�_�Ni��l���݂CVA>S iԄ��n��EJZ	=��t��ߚ4�pR]۽�v�^q8���#�w0W��t���;:�{�o���7�E&6g���Q҈�����[;��.Y�ej}�a�%1-���F�t�Ԛ��.�zўZv0pC�ݳ'��FԤ���4�m�b�c8e��S@��W_�{���Ю�}N��9B⦥xu�$ؤC�*eD:�Z�ӝi�2Tq/h�݁��r�wn�%zw���x��38u���֨�V��k�^	B~��^%mI��7*>���<ӰF0/e�ݾ�f��=	]P/ ��q0���a��Pq-_Oj�I�d�Ϡ�k��I�G�a�l�N�;��HǕ�GiwL��i�D���D1l�u_���O���i(
m����G��n~�\�FZ8X�qAU��۲�*U�6��b4I��Q�o��/�ùZ#�Q�ʰ ���YW�7�Ј�;8mL1���?��z(̀������[&AMjĢh��<G���iy,�Rg��<�����v���\B��z'A�.�|�,�!T�^��'��o�w�Û�4��ѓ7�3��Pl�N�Gtw�I���~�^TP�Iz�ee�1��_�L�����]���Z� �!���K�S}_�pv����{�Dҝff���~����,�#�t���Ν���G��NC-
��	9�:�>7Ӛ���B[�P�_��I��_�	�&QU��k��m��t��5(� �8K
$V���N��G� ��`�h#"�5Qg;	�!�V<�J
s!�TPi��G��^���Б׸���? �J���B�!wQ�w�a~:#�ٙJ�Qg��۳BVW���Gz9.k& ��{p gE:�����$�e<M�5���8i��S1��pՌT�d�T��m���������Un<�%�u'�3�	��`���0��}#��{gY�o���^�Vz��Rh)^�k�A�K�ĳ ��|9��2�������)� �p,�^�'���� w*&eg~�p��Ȣ#3t=P��T!��vs����c��cz��"Ӗ�U�\1�R-b�|�EQ<%G�s�:�N/4�-,�:u�o�\_���j�>Ź���מ0���\̀y�;�ζ����u@Q�2�2&:]�-��&��n;ZR~��>� ���Oе<:C��'f|w�f��2�*���0��?RmI�=�л��/�@�sO�?����r�58W����Q�;h��&�t��"��}�+��*c%�\��l��8n�Չl>t��I͐�}�o��tZ�qi�����p�$O6�~k1���q���g�.�X�
�W�1�G|��B���nO�W0��|<��L�����0f� �ص�b(0	���[3�Qn����ȟ��7�����>o^N�+��2�-�5K`���̦��@�[�A�6���]�9�I��
�H]4Sf���{�_G�s��?��8ݸT!XDA)��}��hP��n�;���y���I/�e��t��*���Vi7���H�����G�f0�S�#�7W�5O�C�:�1��o/�����鋊�@�uT�����H��S�L�S_u9Z��I�86v��*�����d�ٓĎ�`�RV47���Y��Fv���kLܧe����wS�G��6��-@���L�����21ili�����b��.]�ܳF���("̏���;\B�-`ܻ��Z1`�q�:���{p�9`��F��~	@��c��j���n%����z�E�䞏�r����ѧ�X�N��lk����b��_�e�����+�@ګy^~�
�\r(��D��G�mש���peO�໑���v��`���� ���Z�*q�f^���]��J_�9$������H6�8��=ɧ�z�~mmx�B�0̚�&)<
O�k��c[�V24l1'�69?��m��� �$9k](�	"K�ߌ8���o��5zbΘu�|�c�C��ł0���n�
��̵���İŻ#Y���#iu��o8!#:	?.����²�Y�y~k�*&0��sύG��A�@�'�+d��QUb4GT����ft p��e�E�� �1D�޼�Y��<z� ��0e���j^���W��t�8�]Aw�x/X�WnH���DG�ȹ�G�"�>G�`6�4zV`��jiٸT-�$�[i����\����;�bDU�'���)�ys�e�ڵ�*���L$����b��C#��~�ݒK�5����3jV�T$T�Ge���Y��F��3�7�b'�o��Ϋ|GtY��,�b�fL#���H�bn�X�r��-_�������o�?�NI5�31��l쌠���}�f.�����,[O<"�*�miB�S�ً_�^�; �f2��p��:p�j2�3�>�Bm����ͅnb"�{F�a��dp��h���񸗺���9Ec*���5����q���������RL��U���M����@5փ�q���L���)�{p���]��Ë<�AK�B�'��nQ킭+a�Ccu>�F�*��'�H�(��x5�&\���G�~�߷��s�Wyg;��Dy/��*

�l��<��Җ�fR�Oq�X-��v�{�`��8G�F�xlM����M����G���g�c���)4��{�ۂt���rʳ�ˎ����[P�1�%�Z������4��c)2:��b։��r�e*f�o��Y���� ���7#C
??���Wl	*�EA�=}O��CS3�hW�W����;������Xq��Iz�.���;728D6�d'��N{�s:��Ŕ�U6d� �6G�<$�{����R�}����0��~|������"�B�8�ާ��,�� a��UH�!�abK!O!&�zl�-�It�G5��0k:�6	u���a�sG��v�!
�����-��	�Ek��!��,�̘�H|�m�薷��%M�D�3 ������S�.ӓ���1�LS`�D�PY�F�/dF��;����x�Ջ�5qa��8ͮ�F�� ���$h�>Mt�Т�"�8��_����������� �2�)v���:,%�}�p 
ql�>-p�{�=���Ⱦv?�b��9D8
F-1[8�\U�U�]b�J:���):uI|QB����$����I!Y"��<��9���)17A�j��0���[ܗc�[/,GP��w%�����,��/��"�O�`� ��غ"GJ����6��W�ӕ��\���a�v�L��7vO���#���%�Ɂ�v�Ns���A5�gU��j!�cr�?�dl�W���p�������yw�w�m���L�~�mB�؅�.�5���`�_�*��$�]m�T�^}��������~^^�G
.�=}���L͡��s�;;a���9F�e-�N�o+�ff�݃�I��J�Ќ�IF�'�X��J	uyR�$.���^��Rc��2t6o��ۥ+��}M�\M���5��v��Mu�+�[ec0�-Ɨ�<�ShY�����W���(B���^��6s�N��l�Q'9ɪ��Iۺ	-�N��&r
ߑm�sz�Kk���+g���opT/4������X�yn�צIէ����h���Pڥ	�V��6�4s��8�������"^{� �
�S2knP�T�_�I�&��1��%cs�����wmM�Ɲ��V�g�^�QD�s�����)�X�euq���ms�s��f�G���U�<w�	��l[�Ä��RuuΫk�پ�8U�J'��dAJ���h��2?!�"���,���JN��qQ�p��Ţ�>1'�iEp�cZ;���j	E�
Z.�rA��F����[�����?�\��k�y��u#l#��	��p���`���
�h�ZY�4Y!��~�\w�]�S[L���vC��B�i]<F��m�@y��F=���״*���PcN[�������I��><'?�5�6j��{�r<b�g������`�g����ᘣj�u`��`����o-�"N��e0���5g���@�U�(ƅ�j�:	��iwVE�C����m�{k�῕��~�Ku�׽H���GH0G>���89De�� �'vv U��V�qXɯ����A��$B��0�]Ay۱  k]!�ZM�XҲ6�����m�X9t[� ����r�����&�zm�rt���ɯ��R7�X:��B����Q���R��\����n����x�'�������T���}��ѕ���Ǟp8���}���\��ͼdA{v/I���`�ȏ�}+Ƭ�o=_9C+8�BV>�g~@绀W����z����4rb�Ut���~$^���a1:<��$X^¬I܋3y��J�:�B��Q%W�b��`��kη�-����![�&�PU.�����*�[�ʒ�������F�uF�����7�L��g�L�f�x�^~2:f9j�+Έ�Ŷ�?�QO�֒�j��Z����s)������j��uI&֎��	�9��T;T�g�@��j�Ю��<�c����f�
���^R>���=��d��?����T�l��`�c}xdYB�q(�O3C��!�m?���<�c$�{�.�>^oVj�k�hJF}��(�Ͽ�1��~ܺ.6�L��^G=*�F����v�g:t>�I�m���N�߸V�ђ��S,'�߳���u�f�C)�;��'[��i��W��� ��A� J�-�>&��=mY��扨�^j�V��6a��6��7>w��l~@L[{�c�9QO�	���A3��0j��]�K�i�O�"7����Ǻ�'�m*u��|�kЊ��O�F[��uy���`S_����8P]���WQ0N*�
�BkW��h<��p����_����1؉����,�1k�Eg�zج���������R�2jq�F��4p��tb�4�����o0I%p���*kH~�����Bush����O0S��G�dف#V��p��A�y[�A���WQ���@�6@�ѫ\���%�pqK��P��Pr����c)�2�჻[�����t5қ��î�א=�X�_�Q��#�����	U��o-���-!��v[�KK9g�wju�$���,�Y�K�^���S�Ĥ�Za�M���^�� ���Ӧ�h$g����ޓ���>k2�;���c;Ӭ��㯒�@(�Hɭ����MG��.�vERTR0�tm���2��O���K����`���`3��j���e�s��� ��걕跽͜fe�t�(�V7���+�"h�X<&n�if[�MuJ���E�l�"�:�r���@�ެ�1� �Ά:�[����ZE/jeHai^pºE�[�F�P�L6�䚑�9L���6?�ַ¾��L��siTx���Ã�=����߂z�6Ί�?_�RB)������������jey0,�4��4�0N��b$�.[@HõJmv$oO���Q�6������{tH��b^ �aG���G.�ՀHa�=����j��Yd�\�IG����S£֥Ձ���}�Mh(tP&�������9^�4��Հ2w�����0̄��3�aR.�m�
ħ0O��@`���u�y�5&� uk����1�OX�a��zFd�M�P׸��I��2'�08!��'����'&x���m�='��'�*� ]:C�":eVk�^߶R�r7=�6�R[�r�a�� $l bi1&r�����8L�����(�|#��5`���
�0�I���*�dKq��{3��r�ߢ!x硅Ҧp�fV�o���y8��航`p���a�PF�$�M���c����<#��./J�Z�Af��JZ��^df�_��%��\��AD�Y��sGiTKl<�������6���s�w�m����:������˞;���=]�ʎ&{M�;�]�Pr]��.��iF5.�!c���De�@f���y?�ݳc�q]�����C�y)��/}EE3���r��E�B�м�t�}�w��;_Qkx���c������L��R� �E����SCK~0/q2�]��T�b��(����
[�\��pny��\'��wV�X�	�$�	��m6�df��B/(���}�u^ B.������ZLv b�<j�#ۯn8�i�j6��5F��S�n't�{�W�6\m��(�G�d��wz���@FmrSǗ;���\t߰�˚%w�et>}S �!��q�>?!�÷}Nk%J1�_�m��nxՃ�:�Kd� _u�7�1.� �C��gxM�*@�3�#-��K�G��0c:���r��z2�c��V{���P,6�W9�"�)��8��jˠ{�z�2%�<�XU4y�?n�sxBÄ�11}��sU�.��8�Ū�1���}�Ah��x�DՌ{5��W��6z�J����|�e�*��cB��u7VK[>���ڏ>�<Ģ�J�B���G�	�)�0L�l���:�������;;W���Cp!��%���-���/�y���j(b}b�_l�D@�z?8�؄'�|����v�ɍ�ZVC�d!q/��kE*ľ�	ː2$�M��)���q��_����S5䊐T�Uv-����M�GtSy���W�*�
 `̆K��`�d}`���/Ȩ�:�"�d^Ч�|���]$�$�H3�\#Ő���<���K:����j�_N�/=���tS#_)f�P5Cj�v�P��cm���m��^�n����:�3>��(��ѵC&|C��~e�N찴s�*bC�婯�9$Vٝ߱Ã��\��˛��=���~)B��v��[���[!�;F%NT� 1"�����E�h���Ld����6�G#�*I'9s�y�G��9�c㜗$�:<�����=�f��ߨ�Y��\���E/q���l�j���L�����w�7�O���O���s���)��x�[�XI��&�Y�<�wE���­V��Vk��,.jB6`�v)��?vL+�B������aE�]�{�vv�},o�茞�'d���-��8e���%�5^?�� 
�x���C��w�BleW&sւcMp�"f%���v[����B��zg�����kI\PE+i�B+U�k�}�\����t��ޕ�i���uiyz�Q�1%e7���B)�+���{���O`���?�I��q��`B��#��B��@��Ņ^��YzH�7���^���x��
!M�`R�8�um�.Ty��q�п��G��*l�&�m+�� 5��y�-ʯ=$-roSW|���� fBt_+2!��Y��M�����׵�]�W|������g��'.�-d�zS��χ�6��7Ԩ���r\��	����j���<]qq��~�E��0��R}� �) QЃ^��bV���ߌ͵��5�R0�$��)����r�'�zYC�Ϟ���<!I�/H.�~���v����~�sX&��%�_lNDØ��.���騥�V���se���rޙ8�=�SJ~#��t��0���Щ\����vf|{��.�%�)�p\D�a���X~L�2�j��Db�~z�P,��_+"�2���i�������)�3vD=cV7��US>>�[�؇~?Ԁ���e�|��-,�昡?�l��$a�Y��,ϟ�-�9�D�c�>��w4z��&���r��T�r5���,��w�5 �\Z�Y}dI�զN�����o'�v�r���/ڣ^��]��F8��a���03�UTogh�-z@�b�PnB,X���d�|���2� �ʍ�-]=����ޜ۱�cMJ���J	�Rp�l�����ɢ�f��B�VU�7�
�'�.��1��U�m�%?�2��5CA��ѧ�,������[�)} ���7����,
�����{u[�I�sW5M�̛��j�NB��-6�V�ay�E�u�YPa� ¤�
�G+W�7���1���
�l��"{�qf���i�U5�$y5n7��!�q�G��	O9�tH�^�f�b^u�G�XR�j��~��'�,u�|U�˓�0�$��ܰ|c(�_c`i%�ZB/�b��/���Rm��*�c��*��@����WgE�'f��v�.\p42��%�I^-H=� Z��"����ї��!�05ͦ����Ohx���H,-�|=��&sU�[z�r̴F�ڛ��?X&��7���=��g�/iɴ��"i5>h����R~q��XZ��B��d���"��A��%�$sm���Г������7�$C�{l�9n>��v�w�hމ�փxG�H�@�ZMmp���9e�M>l͝k�t`��L9X����R�/BU]s������d�,a� �� ��W:E�k��xөu۪Hk�9�[*H��9�.qXE�K����"���цo��-ɛ_l�:"W��o��W�bdt-���F�c��r;�*�����ѵc
���ڌf��#�@�=�W@�$A����{�A����A(�;�c s�X�]H�s�G��
&8�����ϸv}��b&zv���Ų��O���|�l�%����P[y���;���MN-m#�a(�%���cC� � e58��ɣ Fm*���A *�<\�Z�ٰ&�jEJx�b6+�p���+��F�6��J�LL�z��&J��	����23�H���[��}9J�2#���N$^/��p��OXV�G�jTx`��D�_�� �g�%�\n�Vw�]����[ �c�	�T�q��`�&��\��U�4Wh�Ϟ*�t�����������r��A���!9D�7���k��i�]�|�*G-ˑa4�k�~�1K��Z��̤�����2�հinQV�o�|(�$e>M�u�7�h�bۼ[v�/7���i��`�ޝ�H�P)^*���A!g�o��f�SQ���f�b�ڨ♶�Z��Ӆ��1U��x���vw�$��۳��}���T�[��F�.ػ1�**iZc�,@����օ^��l�C�C	�ĢVC���l�,/�����M|m����j�2:����|Pܾj�?'Bq�l��X����/{�1%�$��u�#^~���?~'|Y�Q���{��w�?D
�%s����9MR`&H�ռ} ��TԔ�n�IQ���n��a���
���Q�]���	z��
��R�ض_q����5�};Wl?�Nn���	��0��*kEU.2#nS�MTO�pź����3#Ag�y(9���NS�s��CoEAN���AoM��H�����jr2�JB
<,s��aUw���w_�n+���PaV����)_���(7ª���6�o@d��tk(�\���	�2�P�	���<�t�oo���DjUd��Q�wܱ��l��đ�Ն̈́y�q�� �zi
^��f��?��l����L 	M��� Sy�5#�Ed�T�;��:.`^p�t[���FW�m��|c3��(Ty
Z>"?i83�=�Z��{���{Y�vQd���䑻���&�`dpZ>�1��^|����aDNl�.��hep�?m♋����o�(Q�u�,���]z�?���f��H\爣�>	Jȁ��2��2��=J�:=oԮdb�L��R��W�NIy�E�B����0�����39����L����H9B7{���7AI��W�x>���_����G�'����l����G�ս�_; :!W4gm��N7t{ ı���%���`�8�Wh'�x�#��d{�ƭ�(�5n�f,>��gt�2�AVW���<g���m�+��� �Q-+yGaE���S+��}�Bf}Zj� ���>���d*)�� ᧃ*�8A��
�>b��*�q�� ���|�H��Y,�7a�ۘ�z蟷�ÔO�rsӠq�T.@M�L�P���b��ꡃҲAB��+�ҝ+�.��%�֦^�Fd�]�7y��
砸FKI/�~�C*Fuܫ]�b̹�-��n�9�PB�,�����������e�m�3ͽi!0Y�*`���(m����`,ћR�2K��q���ļ
�	{����/��1�S�6�!"}(�F,�shK���Q�Hӭ�l5��7�}d��_�M���Hqկ�������)*�����&|.�#����C?�~^�q�ˌ�Ε~�sWr�P��ƇߠΨ�wI�������]���'�/����]��6^>��L���!e���?�w�L�<A��2��2��3��x�r���P�S�'�!r� 
�ᑭ�k�Шa��� ��ε3������z���J�y0鬍���қZ���^q(`d�w��9�c��6�9KZS'��:�ч�.}�'�^% >��x޼�X˲�,5"���Ă���AO�}P�Rd���4i�~/fu_2�S�O����{��m<6 �^ps� 8އ�W�rUc	
~:����{Ɣ�í��H�5EA���/6r�+�qaoid���%���*;����-�����?���B�y�4mZ��m�g�6i�#+����	�O#ĢC���>�35��j��S!��iW������Q3X��L��{�@ٹgIX��p�G��@v�!�z)���i�ő���_+��v�g�؂�Ͱc������A?�h���x'T)-�ZmZL�C�iG��w{�Y2��ږ�=����������It�@J���U�R���om�b�����"rH��;(��& �C��'Z \�p���ORha���"T���L��۰�~���H��A/a6% �����Y$�+K�	  �כ,�6X�V�`�x���w�sC`������*}��|(��H>dғe��2^Eh��g����Rk��0�	��pi!A&Ωw�(^�*�~��k�/ �u�i���J�d/�=�*�������g��Q .,��#�!�$�*:F��hN��=�ۜ���3���LM+�|�7ᱢ��:EZb�pNѱBhG�šN)�Nи�Q����[�U4|GK�fco://-����E�Wf������_y��w���;�w��
��t$b�x�NG��9̈́m�����j��F^W���#���~�v�f8�P?� ����	�����NG��� �����.�H+��������MH�%�+omށ�h�G�\�.M�)�s��u�b�0I�6O���׺ͽs�kU݁EHkYG7���7�5���=���14�ڢ?�Q����|-����z2�9�@�n�_
��O������%\�N�'�G��Zֱ������t�ރ7*a����G���fK>Yy
Tt]4�zu����t�Ȧg��ɳ�w~��R��w�+逕{0��y���)x�����G�t;Y ^D�QUA���1�s�Nw�q��E�4�F���'��vb=���	��m�mU��5�}��F�Q1,�	8��!,����M�mf����
�w���@hX_^�%��
F��G��<l'TY�[j(ƀ�u�/�2���U#�0LeŐj+�&�>1)jOs@/u��-I�}���Q)��w��[�MM�����靛�@5�>H
R�2��G�W��5N0m�M-se��r÷�e\͢QJ@ ����6���$���+��߀L�_���}��I�����(�%o)4%ʺ�������x�������:2r�P�xU@�����𘹾-�˼�(��>>%��d�>�Wm���ym����-h�������	e3k	)3ϯ ��9����R�;�RHL擇�.�n<W��|�|���Y��\ء��?`�d�[�.΋�N�c�8Q���g�@8Hw�1���(� �-�_47�IĻ�N�7d"r�@��w }/�sE�����vzeӎx���Ҷ������RBx���']��8�A�Chbr��,��oK�������G��r?�[�N��X�X�c�ʩ�K����.Q6�p�����XoM5m0��ak�֔��3b�������C�Q�3�v����|���M;�/|Y,mu:7��e���Խ�R4W�-Y�����q�[E'~����7�'o�����C� Ԏ��M���\c�!n�V\f�"���pR�i�֌��b�sWa_ޠ��c#[>Z�PK�!}H�ymP�'��☺�x�k�`ۛ{_sw��R,�|��0�ka8�8❒�˹�s��I!k�|�z�3�y�FS��Zr3!����v����3W�L���`>�_�٪d��<��^��[s"F���R��i��:�B��@x?4U})T%BxwռJJ�a:�8�
�at>�D�~�0���;��6��#��SOEى������@�њ�9����:��4�"�M��Y�k��j�tۂ�v��-�F���g=��[���}s7Z����m�6��	�N��O�����1k}��ܵ��7΍�}24�h����T����I�FZ_�f���L�:��6d�g�$�HZ'^�ѳ�z����/?�yǦ{b��2��pv c��XU�ā�e�N��u�2��y���5��µ�T�	16r�(* حU�.��$���߼�-�X�"({??�1j׶a�w]�t��)��j��1X��T�y�ǣ�m��\�Z>K���O�� U�;�u��D9<;����{Bu�EV-�\5A�v�@�s�-�������d`l,����̤��Gy�}��)��Q��T�*�EEh�0�yq�s��M�'�˦L�4��=ڲ[kQ.�RayEo+6��2���S�7���1hj�K�'�"���q�`>�_/�d+�ϻC@H�)`�,*�v�����4�
x�R��HO�S�h�kV�ؐ��(��m��֭PGyݤy$�؎fbAb;�Wl���Y(jSp_�O4M��z@�$��ߙ�0}�(�:x���i����T{���`/�#�(�&pUi���Z�͙�@2�	*�8%�m�#r��_	�^U��S�mz(��tF����`�J��'SY�-�]5R�V^	V�"�>� �b����R���w.�CvD��ť,�b��������]�^�m���X�}S��̗�/C���(�� � �������ӱ���@�9�j@)�:�}��:��)�BV(���n�si
�}��ۑ����T���T��4��5RG��	��b6�a���e�������![�XYN�Y�y�2 @$d�'�C�@��.['�R���~��"c�u#U������3EBm!�����os�v��.0�{���]�5�O/m���3l��г"")I��^��q��ۉ$7����v3�HS���Ȧ6
����D�]�JTP`�]FCB�瑍�������f5b��������Ud�/z�'Z9����x_3k`P~��P�/VE���0��A5�b���M9�����ź���M�K��KP{y�-����8�?���Y��	��|��2pp�I����#2�b����h��ù����Ѿ�֋�RЍ{��44zP:��G�֙e�ޛ�H/xv��P����z>�0U}��xz�ρ�^#\�ᨆ�a���w�O��l��K%(%�Y_Oϼ�R�����I��'q�i$��g,�? j��fl�'C��i�$�Fg�h�O��Ƀ3�K�˪g�;tP�Q�@#��|�h�<��aA(�#j��}��wNrN�+�
�#��ԾA�Je���'M=�&k�>~�Z��4�+��L�&g��)�捱c���=L��������,��"Ch�o/�6�M} �/Ϙ���{�	7ɠ�HPt�">�����b�����J	2��ri�p�560.��5�SY6�^W͑YWU�TQ#��M��Ĳ��qW� �r�Q���O���HPL��%�X��;�#�o$�Q֔������r����'�OYq��Y~����?9Y��	+�]�2U�M�x8bB4w'1������'��oD@C}����=&Ʊ�L[	�(D؀�>��`X����zgB�o�EX6h q4�6���yw;�K��6�94��< �M���C�%�"l�8��C���+��w	��V|�����t!�Fg	&�G��r4 ]�Бْ��<t5���X�a��5�zk�?'�Q�	���]��E�m���joc�$��K����[\��E$��:0����N=��
�f�fC�
2��v\�s�>�a��bk���m�-�a����� ��B�:RO �6�o�m謐�^���F.����S|�ȳ��Ce��wӶY���z"��}m'�X-��+�Nk�w���|�_���[B&\C�o�b=���Ou�z>km5c���kzDVo_U&O��K�@>E�$���['��սj��(^�
���&j�^��x���)	��� C���[��a�C_١�ff��q�w�I�5l
�KԘ�Td.�;����P(h��<	�v���u��7�H8�m���E�%S2�tE�A@G���S��?��պ��ZU�WhQ\��H���C��x��=n��r��x�#D y_��:%t���q���j��=���f矴m�<�C���|>�.�*u�[���������zq�.r1/�[{���L'0z��߭���ޖB��d�L$P��NB<���z2?.�n7�Z��#:C���1��ceԉ_��ZG5�����kC	�A���?	+Kr��.�Ĳ6����g囉�ށ��������CC�'��}�z`��yDN*����U�R�d���QV�F�,�)�Yp�mT��n���o��X��W�j��Y���v�)Q��j_,н�Pj|TΔ�5���j�{.�8��ҮEb�{��r�Gk�x���]G��H��JJ������d�I�D(;�����wh�J0p$�Ӭ�	[���b�1�c%'��^�3YcWXuzE�wB��.�Q@E��ξh+�1���V#tK���Ǫ:�ʍT�^-P����\ǍK^<�Ꙩ$-V2q�m�RV�2�к������b���T�Z]R�3,&	 [��ᇯ�>���V#(%�b�4�ܼwE�,!yɅn�I)[J�i�GB>�&��
i.3rA��L�:��\�_��~_���֙��"���=_�~	�-�~���P�q5]4���H� �y.ѥ��z��� !$j.�l^ʐ���쉩e��E��&k���R?Y�Hj��%V�{2$.6B���L� ��� +���N
}M�{�}��:�gmniys|)�Jt�T�*�<_����vH{S�Bl}]6ی��1!���^B�:�4�c/��v��2Q��G9�"�#!����}l)�Y�ʿ���d�|��#qaf0Y�{��vV0�]Yڰ�Ib�.���)�p�	��2
��Dݐ}��5��'i��0&L:8����%���
Y�ؐ�\G�BBݿQ�lE�Bj�ب۰��ĥ�JrbX��5����(ڇ�b��[f uG�,�'o��FA�*svw���-g!Z(����M[�6�Tx���������p�u��(K����^�N˳�o�b*�U"�T�cԨ7?s� "�af���+s1���U��%���Ԋ|G�.��P4kƂ�(��p2��_]ͱ�`|��7���|/i9���Q1ܲzq���ۿ���U����C?�t�<�{���'?�Q^�W$=���?Y�' i>"3+�S	u��%(R��V,z��XB7�}�kzQ����X,b�~�*�ՑB9/8���T'��� �}/��%����P�{n@BC�
����Q�y<�˿NR�z沋�鎧�@���{���m���r��S��5E:<	k�FQ&,B˧0���'��н K�j�؀&�.�8y��9��ƫ��E��݊�d϶!��[G� <%��J(���y�4[�"\�HZ���c�b6Ⱦd�k�Z�*�'�\�B5[�Dft�����䦬��
G@IYTT8%=YL��*ZG��6�B��Tp�(P��0��0離��ϊ�d]�$�����L��dѡ}�I=C½=��-,��y"�N~C��f��M����zs,``�5#'d��yPJZ��>�4�иی�o�߾H宄R��D�����s;'!AY@�=��-*\����m.����s�u�f�N}��!��B����w�v㺪��@�Z�~�Է�_��=���MXUa�����c��9��{=pq�ٕ�i�t��	��V�!� 9;lL�B�UwY�f��${�*���-�f�B�T&�5Wdx����� $��:燶�W8�xE��5�>��*nut&κ��)c�+����zH�7�'h~~N�zM��Tk@�p35<*y�T8-LFaW\��/�>͂��~[s���,��!\ rԵ�[=�X �rK�~�w���h^�r���i)"Zl�s���=r�"���V�L�� �MU�&�W���&�T^�ʇƮ.��Ă�s%�:ʻ�~FA��Uzփ9�ڻ2B�3�]�P�l�����F�#A "nׄ��������RGʼ_
���j�YG��MN�?0��QKK�����)��<v�Ș����p��I�t�m67�|Tz�߸�P}�|D�>8z}�����1��:�0�H�W��������}�g��
�{�o���ׇ$R5�`:�iHI���w/�>O+��[��.��뺒�"��&Pj;؂@�� ��u�;1��V#<�rT'̮�b��w?P���u�M=�@�X�2EK��Կ}7�B��3�g�̯i�]�[��%���^���5"���w��B�%���.��dU5]��Ŕ}� $�F�"�p� ���K>0����j5:�T�&:2��QC�ֽ��	U�꣧�,\�K��a��i���#�
H����u�[�Z�G1Q�5pP0�U��E�fi���
L����ޢtW�2�E����/�HRאh�}��ƭ���qq1�eÿB�0l��;(�|h�FĜ�v�L���y�Y;z<g�f�_����r�.�ޑG4��ߥ�i�r������To������3��z��'۲�r*�<w�����s��>DM�"�@3�'=��uGu8iuR�+w�Yq�$~}ë�l�D�P}����eV��3��?��*G@3pE�}Pcg�bz�}���%[`0�E�/
�j��ɫ�XwXL��r��H�e�K�za-��d�/�[���N�A����!b�ƃ%-���C����E@��������o}QX/�Z�D��\d>��)ZK]��+3�&��q��x���zi��y�I�ͮd#�Z��/�	[�)�7�(�˙�.���݇WG|���:9��1�2��8��}���� i�H�
�U��*�_r�>���ξ|�oy��Ġ�9l�P0�,h�G����HqF8!m�K,����'"�u�h���S/@5f|V˘Qx,.bљ�a*��˴�`�%�/SY�/�
�
Ad;/����ᐚ�@+kI�bQ�2���GD��� @���a��<`�i^ݔ�$���Z�ڔry /��s<P�Y��|Ρ����v�X�D,�Xm�s�����)�/x��� ^K�e��}&'0��0&���Q�� J �0��eC��L��+�o��3�6zlX���e�n�1�1�F
�*��O��+�ߓ�rAΖ�;�Z��(��,�L����,Sݭ7�<��"��h��qdc�#zDvҠ��*�����>^�U�қ�#��
m{��(/�w�`��3�Q���hҀ����%��&��Yn�(�UK�魍R�ˡroZ�������;?�V#���P�c��|�{?�n,��rށ�,#	UP;E	�&40���2�<�������&�U���Ȓj�!&� ��H���� �m�`�*���"_>���c0���玢A��p���1����s��H���%s�P4e)��$�\/ ��
�+_���.��W=F$�H�Gt����X���rwf	��IAa���`��ζ{��]n�n����
s�	%�!R��B���#%m����|�Z���"��5��D���v��f�E�l�G������7-�s�lJ�]��T�m�ˣx�1���y��X7�鍔�-eAo{��%ǔ�0�z<�fZ�%R�5�LD.��4��>����H�upG�>`�V2��G���u����嬰P]��i���Z�-����Ƈ���
d�����uV{*R.c����1Gx
��s�;?L���繞ي�'e	�+fN�Y�;M�FAx�.�Q�ݾ�����f�Pۺ4��W	�����+�4cP��I�%���>��h��+r�F��C�� 0�ى�:C�54����������� ��Q*�%��v�OR�-LĻ�5�������c�o��YYc�.Ѳj%S��s|*���0�Z�6Uꩍ!�f��e�vE"���T?"�M��n�CLI=��g�h�{�JC��=����,�"U�J�!��s�P�R�R@�U�1|�Rq�@���8�.�|�Ӥ����$YkK��ijD�p/-�Q�x$CW3�}Du�z�#M�țр�!T��(���:y��� ��T��50O��3�dV(�eu�7̎z�ǠO���U�@N.t�s8m�a�5%$̊Z�����n�ٿN7`��Mܒa�W�����3f��������({��u���.���BA;���wؒ���S��H3�[� meD�i*���AQ�_:4�u��o�i@RhfZM�s	q���V�1�R˶�c��oje�p�(����T�"q�E�x�l����1�2(沖x+}�3�(�i8ߺJ���ҰS#n�x P.z���J��AZ�/(C��
 a��l���A.�/��	~ѢT�ΠI'�
��rH	��W�Cm����W��1�k�{�F���"5U�bE5ց �x�z�sW2���h�
�}t���5>ߓ�E���s��X
24�+P �hTH�VR��U�����	{�����:�UH�Y�z�}�V�A�t+��������.G<ߝ�a�9���`ң���va!���j�����YB3.� [�@�&�m,�+{��.ZV@���M8G�f���SEշ2���u֭�Y�z	`>r�INOg����)_�
��~��τ����DU8ҏ	֘Ƙ�a��n�AN1k�I�a��|R�������2�XM��2����ŋ�T��*�Ij$��-L��uwL��5�vm5Ϭ#���Q B��)JE��Zו4V{=��s���z�*�t�=u��C� 4lgų�L��Z�s�һ%��M�Fc��O��]�J���ȳG��L5ށ������(�Z\.
m�	,v]s�:���Q�n��	��!#��7����m�6�oJw�I��v]�}�"Ƶ�ӃX�@�HLr�!��a;�N;!_�,�\�����R�~�����>��_>K�o���;��U,U뺬_�U�z�	:� Ȕ�4�ܿ=�	b����cB��7����������,�s�`٣��a*8o	*�è����B�pydjw��[�O��܄�y���{�V)Q����������n�x�S��l�x��J�	f*Ȁ�S
���;��l�އ�� \6R�p��gaU��z=GgGN9��]��!3PG��(��;KU>��r(QU�6��Ug/�2� j��Lsb��5k'�����R@,� ��l8���'B���T��|X��6�p<aP��:��pg�>�8o�,+X��6�&.K8�D�)

P�{��4�<�]�X���3����35"��`�4���W���
��a�_����\�6*¢�]I��%tPҰ�2�X�:OOQr�kZ�1�h��%۱���0V�Hny�ag�n������"W���r��s�0��dr���Eh9������ V!�`7=�&��؅|�Q~B�pXrEq���/�gA�9�/�[\�:{��2��Γ�$��?2��!��G�%�[������]�W���R�L.����ᏸ����>��q*�ȩ��&�=�ӑ�m�+�7w�SyhTB�ֿ�s��SaRʦ#cϺ#K���Lf90�m�~��i�zZ�x|�p\
x�	k�u��=��C������Dz���?S a6��!�Ƨ�eF���ɹ�ʝe8l��"S�T�T�,�.���8�<�=_D� ۙ�q��fB�������Rn���;�M�v-"kw��*m��]�ug]w����&��.v;�I�����>�7wcn*�+�P�ċ,�};Tmp]>��� 	'�D��%�,i���'�޾$lQ��T��G4��J����_Q��m��随_z��m�pY������;��������m�f 4gF��^�WU.�d$�����;(�p �<�v�J��Wǎ˃GU2�a�4Az�99��K7�%�݃�c����j��a]����.�KM���X��I}'���
��j�"� V���n $&���	:���p֊��`;���?5++�'V6h�Ϭ'v��8�
J�%��7Z�c9BY��
xy�8�98��
��-'��0��;����E�=�ȋ9�x�dsՁ,��k�EH�qnw\�BٲQ���N���w%�iN�`U��@���DH1��n��@3�����'Ě)FOy�;_@#�����x�Ӏ��*ė���Ɉl�-����N:v���d�ք������R��Y���좨�5�y�$b�2{�q�=���W�j�˃!��t���:�qpX�T�G����t\^v�+���V��A�[��v@��j+�� ���Џ��q-|^P��Tn'w9���uu�z�t#3IZ�I� �g���ҚD��k�R�?�\����'p�[����^嵮�n'3~Ub5k���������|?d��':�c��	�U[�ƫ��r)�� �����d��?qQ��]��m�ty�G�@s���۷iZ�7��4&��A���~FF���%-d�����r�I����jM�QitKʸ�olQ�u�D=�jR�s2��$z<^A���>NV˻���	d�{kӅr�YDVI^�?jq�1�z���Nߑ��t���"�{.�le�]�@�!=+q�@ھ)�$2�e�s�[R�qb�vb �O~̒+���C9&�Z��+�[��*�Xi)�y�����%�~1k�MƉE폑1�b���r7��\{st~���Ef�oO��y��~�<dG������1r:q�3G�Ȫ`��3z�Ǐq\V3��yк*%y�g�n\:xLP2w�\�J�XHo�
d�F>����9;���$A[K�:��j��U��WiǄB��Q[S\Q����t�Z=�؈������ ��=C�q���l�ף*�Y�+�65-`[��A3ʃ5Q�-���!S����sU`�<���Q�V��>��������J;k����0�S�kr�A�
�>J�q��1;)B7�(�X�h��a��r�;aR������u���W!���<��z�2���G^����=��Y|W4�aJ$��-ф0�m���i���f�E��0��:�cF�ܪ�]_�E�#"�G���Η/^_x��:W��ȳ�U��&��;����R�-�X�ÃD%���q?���d�cfId|�ׇX��m��F^��Z4�+	�AE�  ���mnA.V���zu�~�4�Ow�����3"��u=�S��]| O����p� �����m��4�Q|It|��̺��jfou_T%GܤJɑdύ��m��.͢�K�sm�z���[�xg����	�/�!z�6�A����k��[º֩��4��|�"�̼�LӢl�I���/���[cso6/J�˭"1�ozPo�K�/�[x��M.ߟ�@3Y��}��έ�l�n[O����T9n=C&��Cx�$�0�uF^V^�֎1R�i�����2��\��kT���Q����W��l�\aTX�6*
������^���%��<&g�cIl�s�U*_�t���3�M{�.��d ��)�-�?���_�5E�i�sO]��㫎bI'*J+�qs��o�b��X[��k}��ut�P�P�*��^E�'U�k���E:��v� �x���A7��쟀�~� ǀ@3��{���)(.�E�`h��m�=�u��˝�?P�'�pA���I�L��IL�Lj���G]��\bhu��"�%FF�5v���୺�.�w�B��D{��;i4sYF����)�v���+�#\���0��%q9>9\Qa� [�}��� ���]M�uy	m�Ւ'��IF�h{��?���BdP�9D��AT�y�tL��N����"?ǣ�_.� �K�!b�����Zv�Q@kzv[��������V�D�mQ�`�q/ܷ�)�Ҧ9�?�o�T�������^|#���Z���7�I�|�a��|�J,IyBg�h�3�y����bH`��`��G�6t�c��恦p��U�|	����<�d��Aiq�:�e;�-fC�4�W/}U�� ��'���d��@d�	��<�T�l�`>��y�o�"��2���k�X���C�����ʨO/��@c5gƕ�%z���]�@7�+��&�\�O�?y��[v(x�r����A벥������Uau�%��/�rK��ܯq<��F����Q��|�0�m�iȡ�@kLɹ0/<4x�i����'2)�%07���c[�خr"MD���g�me�B�e>,<EGE��C[�dg��=��B@Ô��x�'�M[�pd�_Źv�s�N���(��͛���"hs����LxyNt��	-������.V�=e:!|�D�w���u�����Wr?��wVx�����"����3iN�~�ܺ_��9��+�J7Ab��a����%xt����=�M��00�5>����9�]1D:wZ��=ϑ��u	&oR*o�/��a�������E-O�ǽ�{	��P�r	�O��]�<;1c8��}L�/h��-R�����K���/2�+���?4+Iɇ<h�E���r���k�����㽮�|��/�=��r���nI�Z��z��7��fpw�1����1�)AIuX6 M2�r��{��
)�F���K~�x��@�i,/^���tz��P� 3�Z�
.�Um^���O$ tO��3Z+��0�?G����	z/$�4B�U�ʈ�ԝ9hiNZJ��|�#���>��1Ѩ*�B�"Oy:̂s�t�0A}�e[FȒn���8�/�琖hn��1��r�R�2:Z���{��F���\ub�,��">�<οr����
�j�]�����lbU�nKV��,���:4z|AK�f�P�y<����<��
څ�ABZ�8�(aw�@^qJ'�o���q��ܐ0`%G��(͹��~&�����ۙ����B�`��7h�:?������Y��w������x�n���bOm��j���"b��U]��ϋ�����!XM ��M����x4�����K<*u��wlU�c�U8~����f`Ƞ��j��~?C�NZ��%v� ^��cI��+�=~]!��b�9��\(�ΣJ rw��}���#[�)����3oF�m͞���,X}��{���"����]�s��L���b�ԇ9���`�����F`���з�����{���ч��K���|5�!�����y�WF����D8e��U�e�e�4�E�&g�>��`78�L�J�ӝ�q�SH��-���s[�Ų��w��uֵ:��]���p���k�X������0���e��2bc��Z:�L%��)q6�o**�.椇q�@���)��qDʑ?���}��1���Ux턮��)��\qxW���/F1k%N�eͪ�u1�W� F���n�L��Ɯv4�3C��Ik@�9�]PƦ :��{���^E��1�t�­��%ܵ�`:&�J�l��;�>�*�#CY�g�*V�'��F.�����og�O���Yq�_f2.�5�[hX9�tt�?��e����ʾ����e_�r��荐��m�\	�[�4pX�m*�h��ӓ=��vjش�1-#��f��u~Z�s5����s?���xWǡ�lUS��S_-�������>��g�"H�5� �A�!��w���>@no4�<g'x0mǷ��<�s��СC�E �����=����,��:o�2��I�&Q���r�*k�׀8��2��8�+_Dd�ҳo�R_��LY�H��:F���\K��&�������^ �a�u���j��Z�z<f���s�]PiQ�!���07�dUJ��E"W�}���3e��G̽�fbX���3�Ǚ�����j��vc�8{�a�E/&{\"�����ߟ+,���O�~���5����Q5�=~&�5�Ḱ����z@��C�A����[Q���QKa6ddD���^z����o��>Ԏ�٪�k���R�s�M'EP�0��@I��x=*:�v�}M+��SVG
���w��圄���'U�
[��|a*z��o�|� ���t�1��t���7����H� �#+���iiG �-tQ����7�ɷ9�{L{�2�,v�v#�Ĺ(�̱��M@��N��4����� ���ĤuiYZРUf�k�hN��_ϭ+q�$VO(�Q3O+�`5�5V-�`�*�Jr����,%4���l��q���1U��C@TU��&Y������������|��v��C�v�
u�,#�Ía�Hr��
��si�0+���	V��ѾJ3Fk�E7i;��`]h��G��o�W���npY��Li�����'�?��2&Hw���լ��<Ρ�:�>Jf�):d�S�]�L��x����h�/uh��v��6tz����%��U_:>d��q�@<�a#٨��Ɇ�c�)�A(0 %j�c-��Y2Wc��s:<������0�``Z#�\�3*�d8�|�f"�Ŧ��@�a��w�$��*3ThC���;����g@��\�V0>�
���0dU�I:UOo��� X�J���L��F�vo��Y�� �'�o[�|*�,��rB��t90�P�A����k���(x����*�~��W��W���+�e�c���w�������uD��?�8��n�'dZ"bg]�ǧ�*�Z�|�+�������B�#2�t�8XEr������ħ� �����d��G
��Pf��㙫E�g�	.�~\Q�<�o5���RV�$����zq-K�~\.�:S7�a��0��� �[�_L�/�?��5$0�h�i�jv�i%�R��vG(=s�u�PPf}�~u�ب^�c�]���5��ʓf�:�?��`6|(��?�c*��V>�X/y=H�w��\�w=F�+k�!T�n��*VK���̨~�:,��w�pSn@��U8��v7AϽ�%e�B}�;A*�V:�D��PG[��"ZT{'G�deth��%P���a����*��]����_(�&c�����k�3(���i2�껟�Q���1�V,+}\R�8g|&Y�����2���P���I��ʦ/���	���B�U�/����;��F�k���@a,�=�l���
ʿ2��7����>>~M�M*c0�4!?ḛo	^�Pe%J�
DDX��@�B�g�tq�s�w:�u����֣�J����J6�x�'�L��U��γ-��J�@Z��̃F�7Pr�V����G=|'Oհ;�PqcҔ ��<S�����8��ل����EY˂���+Ud���ҝ�w4Wr2\~~&�~�+�h�Z�Vn v�z���3N�W�%]��6�5�lھ#x�0�$3�2*�+���K��Ƽ��
x�Xh�e�^��,�a�Xx�]dx	�|�/�'l��)�g���}*���_z�v4��&m ��4//�:�^�_:~�6�cn�u�Źj^@Y0��D"�5���Z�j�7�ϧ(��VU���� e��_���Pyo���>���#b�?)3¤��¤�c�z�:��2�s�g���:S<F�D�x�^0}�*���$B���yI�P��$��f�7��CBY33�(51F��<m�!�H>?t���G�h+sC�J�E�7��������Ó�j�OY��C)�Q�����	|��C&��'���4�FM�}+�� &wes�D��˽9�_G�"���u��[�{ >��c�t���LX� ��Y{����b@)夶J3�t�'dP�im=<�M��+�4���G�\^.ޟs����Ĩ�B��j��X��� _*�Օ�p������#�^$7vܳW`ܝ�+(0pXah��*��vH���6�A�9#ø�
��*lȼC��i)4�l��.Hg雪�ud��j�ز5�f4_�%����F�p��fA��e��S�q]I�o�R�2�"65(\��=�-vZ-S���$�̗S׾��(4o �����#vy��<�r��Sx�|»���e�B� ��j�<�����m���G��ؠ��&�Oz�@�o��f.��Ϋ�?n����q(��.����m���r�,��*J�֐1����?k���*5�?��Ww_��g4oʕ	{�ǇF�D�x�XivӼ�&GUl����Or�P*xM�F��'_D�����&_S\o��d�Lւ5�����J%������:�ОͿ���3���i�7���@�Q��~7k?�
����k����u0��+���O�_�aK���#�W�M
����d�s�ּ��4�������1K��'���=� �33�ݍ��r�E�(-�JwC��r�
���^}�r�ŃS�	u
���n41�Ѡ2Ҁ�Y��I�	6��G^��c���{��H���L����.��Av.���	y���%�F9�*��B��k'�1��+k|��z&B>�$���y;���~����&�
�۝J�Ao�kt�G�c`B����`i� ���	ٞ9~@O�/h�M���>�-�����\p֟��D�Vv��X���FW�8�vd�͞B_�H���^9�;#��<�j�]����z˴fP�F���u���Jt�g١!��k����<��Ag���07��.CN�` 7�w���G��3ٰ�r�A�5����2B|�b���U�W��N�
b��}]��"0�:<g��nV�4���t�:���<���[��w�j�?x����WF*Hr���?|�����1PPHV�.��9*
Κ��K��0�yad�X�) �`���x�0?IS�li�|'4A�g�_���#<��gȃ��c�Ú]�r/k��˵&� �苽c3� "ٹ�V����q�k`�u^��79u���ԓ7;�B��g]��̘ۣ��E?�8I�Ϙ����3Q�hߍݧ蒁=KO�5g�oԧ��h�`%�L���S �A.֨L�|��ݴ�g^ĜV�"�A��q�����N޾�i�*؈=��k4��+!�Σ#��y��bQ���fr�+�i��2��"-��a�]�H6�ҎL�����;���_
X�~z%��2��m���lڌJ��YK��@��IR_�V�0ն�a�?��
�]~�q�j2����b���s}W��}A���Ԑ�:���*i�M�D%̜m�g��Z�R�;�H�f��Y�ց;�a�Epʹ o�F��b��\#L06�Mڔ,� ��O�_f�*fIPZ���l+���`��'	�?[�\�)�
��k\�#�k�Ɋ.�ZJXs���os³Pt0PB8	q�{oa���?8y�@����=9eV�=�H<��>đ�l�V�V:]���/�|s*DB-zh1�1i�s�\�Pva||��n�W���S�_Ku����q�=`(�]���	�-N�� N��Y�*���� 2�_������<����oT��;^LK9(ď5�=����m���bcꂈ��c�EZ�[e�ó�9#?����ַ�r�d�*]��emO���T��qR,�a)�P�4}�h�ٗ��\����q��fп1/!�ΗV�u\o���G�jk���d:p�,-⾩[}#�-�A�a�=�nAH�h����iz��"�q4&B��'��Z�sV�I�1����V��9���;����Q�0=��DC���{������(���>Q[������a�0[d
G��R�:�ي�d�/ �
�.
ݐ�m�s��пoa씑��sd����Yኆ?q�WG g��VS;k�(9o���=���G�f?������n7����x�� cI�;N扜�?
;^�ϡ�=��8N)^�mu���(H�b;X= {��}3z-T�u�%�O���N�]�A2� s�p�X�Qg��ֱ1qM�@��9�7M�j)c#Iq�ߦ'�N�ū�� �ܴJ�9h�'a�;�m��aI!Ok��]K��6�P��� 5YH}G|����?j/b�n�k/B�x�g��r��X��by:f�Ҙ��x��zY�ê�BW���㣵�,���7	vF�.�f�>�Z��.�H�'՗��O�;��P\fsܿ/W��4�׿�D�x��+��G���qgEH����A߽���C�E� y������p� )a���	�҅YK�`�z�WJ��n0\�G�Ll&r�K�8��͵Z�tb��L�P�g"*��ƌ�˖P�-sceD"Qun����\�A��V���^�?���U��-����H�X;ϔ��B��zO��d!0"��T����B�?B�3(�������eܸ��8oypx!GM�L	.B�q����҃�5��ѫ��me�����%��O-��&���
�ӝ�0��x�;G�����ǓL�^Q�t�U�D2�fK)�y���6"�fk+��A��Ĉ��.xQ�E��[�y�U�'-ΉWV�:���O5���jp@M��cG�T�@p��Ym���\�8��ń��+��QMvw:����nv�����3�����"�t�+�ݩ��hD� iZ��Yp��ʱ���m�f
��]>�G�/w��6�0pL�;�H�(���"�ћ@��������z�h��Ц���<���Q�璣��������Ж��+(�-W�X���*����uӘ�\j������ֹ�e�,o%�C��d���N������8�T.���*Vj��g���������xL�9r�^jmvh#��c0�w섐c��H�LC�!�e�F�l��r���ʉ+#{�XNZ� �1d=�m;��3���1�YR��Y��?��Җg^�QX|�73M�a������*+�4zMus�={t~�gb�T�ae���.�.w��=pi苶'�^F�l�]Q�c9�֥>X��G�웃i��	
/%״ȍ���Z
�Di4Gٝ_�ƙ�=�:i�`�?�XȖ ���Qg�Ln_"�I.�B ���zʄ�a�e��H��w����E�u��V@�ґ:5����,��0?���N`,�
H��.�}�A2{FA�,	� ��D<�P���ߢv�k�n��I��4�V|%����6v��d�H2����1�_,j?�Rc��ȟTD�cI���"�*��MCR߶�o�n���������Έ�h�*g�!�)]+Z	���cͅ����B��"���-��j�r�� �ъ��eՈ�	BlUl�w���)����	��H>�+�w�S�)�ES�80��M9�eH�['��GK�T�W�S3�g]������G��PYz�.��7�����.�ы�pS�����	i����}(8l�+VV�<�*`���O������wzȏO:�4����e��&;%q�U�R�!���I2M,�6)d����#��7B��\卨��y����K��z-�h �����Yz�u�]�)sd�こX����@��ɢ2%O����BTuA��P�V;��l��	'T��=嶘V@�Y���4�J�^6:ǉ����9<��By>T@KQ0���'-�nʖF�~Y�v��S)L��j���0~|ADn���h��wҏ����G|����;�	P�0\Z��-9�@�w&8��$
V��HWV�N�I����sUd�q�\�|W���;�7�xa[n#	���C�m؊�'�]A��]7{×mxN��I�Ix�u�H&,�"p)��#��������zOY����k7���,����џ(҇ηMc���wD����,���LF�_:hA�Ҭ�tSYy��D�e�dA�g�6������䃖*��[|*��E9s�Z�}��H�k$����"�}P�Z�HEG�ȧ���a" 8�jJ����_hl�q֤�v�8v��Qܖd� ��	����L*���ᵴ��>B�a���i��9��1V��.`��g9y�����y*TW�K���ckM�w��Xn©�[��Z6�?%��Dshި<%	���涚�.�ܔE�|W��ӿ�jYo�d��҉�$F���!�7�D��)m��l��/�繰J�+ ^e����+ݧU�ׄ�\����abF>�����[3V�;4B�@�G0��UD��D�#t�>�����f���>~ޥ�R�]�Ļ����X���D�����L��_�AԲetA�����1vJV��<�֋�Z�ʏ��=�|�[�{�4�XI/`X�΋���杌$����s��T�:���I����(�"��|k����g�����sf�����	F6�js߂}���$io��3��V��\���b��.܉$�W��^��ч�;]���{��T�, ��:��m�n��RP:$�������s��R�����0�f;�#u��t��%oH��/���o���l���8�y���`b3	�}�v�����t�qW�vN������XR�_cV��D������K�[]�wK�{���Ҋ�X��^��0!6�1UM�՝�N%�[�}є�z#&&)×3ud�/w���p���a�U>%!�����'��2�{a�r��t�1&��Y�31�6!�Yg^�˹)O�@���"_��ќ�C0��ճ_���Ə������5��{�AƨW�v�D��@�,.�׶����� ��T;�4�rU��f�Nx6/(�!�@��R'���F�e�]�~�உ���F(���U��i�GV�d����O/%G�!iT{�\�r.�%c�0����-O^ҥh��9�#zht�'�nQl��	���w ƽrQU����
�]NKc ���o,�@3B'=��f�ܛ�d��Y�"ޅH��ר׀�0!�a�0n��;�pj7�כ����V��|ѧ��+y��������)M�^�Մ��g�5��;�JM���^pY�����~���l��w�0$
`���|�"T��%E��`��u�	Z)��g�RH���Z���`�N×�R���%�9�� ܋��66z/����[�X�>>�� k��͵��fQ�u�N����_Yr�9�K���`����_aܣS�vt���L�ђ��?�iA٥K)و/
{�P�%�j��+:����͔�hh�Wm�Lf|�6�T4�d�aY|(�<������0I����
#1N��׌���ᵲv@��r���y�J�N�r��\7f��2G���%PV�Uf򹋳�.ՠ����νvZ���κ0�M��48\��3':�kZI�)�)�|����Cmp~�DuQ8���hjI���~���D��Y�L۠��W�&+ۻ=ݍ���92ۖ�q�2[��� �HgV��� :��b[�l��� 3�}�%��%X`L��s	���85��,���ǇR[zm�D:\}���{�fJ%�lQ�E�cp�q��i`���X��y���_�׻�v`�,���o|��Ƨ��8�e|�Pj\B 04�.a��[��n�A��%ӕ��ѵ���EX|;�ޥo�X%J�&J���e��Y/��Eد�O+r,�� ���e���}�I��5߾%_<����m ��}$Q���0e��]N�.��S.�!Cp
'���T�$�	d�h�$Є��"�������ii���[�M���-bd o�ح�DKcV��ަ�C,�<��ifk�Ŋ2��G���`j�Y�Bs���O{«B�	�R�����������0��ʩ|质Oz�3�X�T���IQ�)����)��@��f��ĕh��Db�
�!|&5M~��rd����v��-`�1�OwBCp�0!���7� MM�L���Y�W�z>qRR� B�Ӝ[���F:>�\�E��zDF�B����r�pY��H�OU��[ߋ���C�M��"zىm_�ye 6� ��uk�)��)��F�g2�͸4��6��| R��g;p�xO�٠zC�hS-��Lߗ]��\�^�T |'�k��\r��>��:{�u�ێ��r��%�#s\,��-z(��-��3�UA�p)�����3r2&�j�H,���&�d@$J�o������jop$ñ��f���Gq�3o��"@�����|���Q�{Y��Z��=s�A q�a���Ny���a�����Rs�t��� ���8������X�;NԬ?�a5��b*��^�����.�7���Baީ��SϪ�3���7���0�?��d����V��MJ�Ou���� r��T�>��V��['�)A�q`м����1�5�t�6��̼�.	:�F"f�(Q��:k2_B�5�]���/�s���b��������G4;9�F�X|��O'�PUf�fd��/�и�0������%یGvp���P[J-�{z��V�c�l��v��E���O(��z�v��Ӣ��f:�Y��7�P�8fm�DK�LT�դ:j(�bP%K���S�âǢ:�ܸ�U�ڞJ��8�ɐW~	��aQ�%/w�*rq���Y�t���@к}����F�@��u�#e�jz{�aQ���[TU���X����8�����!@�Yb�/+[Q��N�I�\��dG�!�
����Տ>U����<��Q��%&˼�/p���(^��-?�o�v_�k�q�����4~�&m3�"���7h��٥?��\�6l�[���<��P�;�G�����>����EH̰����a��~sP|�l�ֳ���k~��n��kA�,����0�J��cLB�#U|� �� ����`,1v*K�@B,�[��:ך
s��*B�]�i@�~N
X�sõ~Ur'y��T��L���7��rʿ�@~��V�F��7����ģ��x	�2����p�I����'y`Pz�F�/_�ۘ>�H;$��Z�	Ǳ���P��w�FSظ�>���d�#��Z%�ª��EiO>��&nE��,q~�^sQ��-V��+��
9
���p�&�V������o��P�!C2/ܙq֧���&�����Φ�v��Wй�ݰp�Ӛ���C-���!ҳ���H���j�`^#K�ltB�:7����%:�X��)�o��Wt1�ha�����϶�(�mB��6��yw�����պݫL&���Q�P�ÞU$P-7�C�R'��Ѫ��d����.?�?��y�|ik�zG����'Jr��h�}&}�?+�K ����l��җ�1[� k��lآi��]9�� ;�g�Ɵ����Ӿ��o��b-ã��*8d�v��i�|O ���'��$+oՠX�M�>\�Bn�oP�s�_�D��գ�+ݧH�5���i5�$V�����F�d������$�r �WK��&��~4
�yg�?oF�1�h_q��0P�W��Ez�:�M�
��*�}dʫ��$�?�/�����?]�U@:
~"�
����|h-�֫���X%�e�,�A�ܐ��/i/'�1�jݑtfX1���$��0$߆X��Rd3�'X�51�a��M�7ր3�������6���RT�81��9������\z��"��l���\��h9k@�h׻�X�Ci f���1����
���Sy�g<x��0yH�T��m!�c%`�֕��(fJm�}��X:���+��"J��Q]��Me+l��H���͓��_�1���}7fȼqo%���<;��jR���bB}�>����|G�3�D{��\&Fh��>�d�,�;?�����B)*l6~����#w�N����Zr� cE��NQ|�_+��ةG3D�0PB ��YK�{,y��
����i���Ҟ���5A+E�8�\|��׮�D�Ť��/���	�������'@��ݘ5S�t�v]�)aMy�i7�c��k�uV/\s+D�C{�'���Ֆ�6�!�#��+�7'�y�K��袆Ѹ���Pb���.!b�J��� =bբ9��By:B�:���గ~-��(!�@	��K�P��kVtAL;KQ
ìh޴��C�m��:&O625�B��<���u���u�sآW�?Yr�ͯ�����:(����]���<<v�M��U���Ci�a���X�K�'��cl���i�'K�y���k�"y��R�8a�<�L�Vk��	e�ɗ��T$����ܸj%\�dH��G�PWĖ�ý$�R�o�{���=�B%�$��ר�`��_��s֯��1\T��}�8J�X�>�G�3�&��Z봄����I�|k�v�i�@��ޯZNȴ�����y�yy����g���e椭�W�B��eD��*�;�u����H�/?�r0ޒ�}h=h�@����-��/\���R��2�:��9������HB�^�7��m�j��K/�_������Y�w���b"��V�3�h�:I��
&H�Dn��4�k��c�m�()���$��HIk���M�H-����g��U��,��c��9ߑ�Q�d�P_$�uc�t�<{_������&�Re�W9��n��hv�L��C=����)8�,#����k�ׅ�]JP�MW��c�03+�%����*�ڭ���R)���.�.@�em��������1B������v�Y�����-(�op�{��`Wt�]�C��Y��&ω���hk$,��w�8f⟇J�q$�w*���^j�]%O�:�!ꁠמT��¸��8���b�`��jmiwS��y�E�£��^{�'�t)z�=�}]�ø�1ϕ�P�	�){�{NkI��$�ۡF<�x�F��)q������� ��Q�n�'.œ���0ͶA��f	.Q�-P��e����Vp��I�s0�q�Y�2�r���\��z_$�ܓ��dzn�� v׾�]®�����o���I�9gj\+UE��߄my��4��ŽdÖ؍}*9�}�����|�����R���-V�MG���1��G�X<�-�nh�\w�+
/��L��|��\p�}I��O��5�e�XhH�>����-�d��_l�h�uuC�>>TD:�'��:�%�&i;�y����:ʜL�t�WL�����"��e������-��P\�ë��6��qOɎ���Jy-4�])��%Č�<7�|�s?lHcw��(`�x?��K"�<xz�N�u������&P�ЂO��/?�	�iA�rV�g��w47��VUનu������YE:�����t�p��܇e`���G��A�
~��Ŧxblk���^\U}��߅���G�0�l]�6>ޞ�~ 5�X�� �]_�PԘq�dP� ���v��:�����&R��Q<�_%��kmj�(r��*m-%���n�{^t��&U�tD����3�d�k��ɋ&�Ϩ��� >ZH� 
?6Ы�R�#6k�'�M��� ��e�����= �#DE�ħ���h�Wa\�:��pAT�O � ��h�)� d�9ى���E�YN���=9d������.3pȷ%��)���?_-J�Ht�lm�Eg)��Eo�(���=rO�?9G����@VSi���-#�J�O�
n%UGM�X�WƧ��>�x���:�v�=0 �5���)�$�}3~�c=N=���o�@�4�h<P���@��(ę��	l$�4��5w`�S�͐����vu{�Rr5�\�}�w�O
��6�U�������]�̳����@a<��7,�Y�����2�mj?D?M��]���C�.ܶ{]�b�6>Ǌ�'�ݼ����vd �,r�����S��T`t��v��}�Y��Dp]~UA|�-��`C����ޖp���Ql�~������>�!Rh�T�|E
���'+a���b�H��O0JL#����L�QW$��-f��n��y�<�_��Aq�|�K���� ���dg���K�ߕ��_/k�\
1�� cC�$z�cTN�@�����ű��l5՛>42��Kj��ze�H��B�`�`yN�����Lv+��%�0�+q|�d����׋�ZM�ݛ�����sc&���w�u����]����cnC{��
.��3�L�p�|د���H툨HK�}�p��]L�jd|����~�����Ε7��IM�%��X�M�#�����*��^��f��!6L��P]U��p�Ŧ��CF��/���c�$ԚݞQ鉳gL��j,�r�!��,D��AN�W+!,��tۮ���c���G������z�q�i#�8K���?���x�K[uyhU#�C�Exz>΁'r7Hc�C�QS�����Ζr������J��6A�
2����띛��=�y$��_<� �f��c6]-œ�^����ҡ꼲�ы]���ъKhH롌1h��,��xs
5ǘv�S]� ����xg���-͐������j"�p�c����	�CP6d���B�%�f���LV��d�,u����
B\�OfUE�y}�27û�>M�un��8ҋ�f���;u���8�C�-��Y�l��U2z�u�Ĉ���|����]5c�[-��j���&��a�f��#���o"&=��r	��[���XJ�hUԅ�`�<e�V4�B����U�k�:���y\�/Vv@H�nEr��h��KOm�>CChq���� �Ȼ�<Um����c��!M���D]��`��u^!�� ƺ\��H�]"����+�m[���`Q�ϓ7aT�ao�PO��'�e����)�$y��?㒕�=,����G�g����¤��(d��SA�X�����*��29 -��U�
.�Xl!�+���&,�JW��M�)x�n!�缲bL5�UZ���
��P�;��N� B�Ehڻ�o��"�!��.��n�|�.����Ň�jN?'���٪ه��C�P֞椶�8W���p����,��5fW}O3a�����6*��S��4�b5�Kjߧ�"�D3��ʹD��`��d��͵���۪_LQ$Y���*��N:]e�"NgyU#L	�ˌ�����0����8,n � 2ɯm�v�\p��6�Ԉ"�2��E�c<pu�/���k"�dFds�%[oR�q�������\�W���8]c�Vy6�1y(�{�M&{�u���
̙���]�j�S2��������$v��!~I^�n5Az>U��uqs��;��� ����v�UT�-�F�ض�><�����!���;RK��2y��(�uԣL�l��9��H����{�R��d�۽�rI��0��~��h����������79.�t��ϧXܟ���WxހOW���`���*�����
�,����h��(X�=z��G��u�# .����j>"���AMk�C�\����w6-z	�ąbirem$؍��O�!�V���b�x��-������zrת��s0��齵�y�)j��P���k��IdUu�N�p����7K�l#�Lo33�В����#�.:��'��l/�N�hsG82�ӱ`ͤ�(7u*Z^����a�9��z,�6w^��֔�E-^K�q��K�l���1��ATn+�����0*�nI����;�� R���O��y�Q=-��z�F�R�p'�0��-j ���c�%��gy����tTjv^W��)�^-tG/�iCi	d`��n�c��'��ꖍ����YFG�[~]�i�($�@-����" �J���(����u%|u���X|� B�,I��W��?���B9 ˘���,�$�a�0F� Q�>��`4���F��V�T�-`���Qs���d[�Xdzȵ6�`��I�{V:��*�(a�z��3����:d�4�'��<6����c���9[�nn7KbN�˚��>����}��[�~�n?�;Q�u���b3O�o�*t���@{�'6)�B���Z&e��#Ζ�hj?	)ԃ'�tŻ�B�v�C�Q�� �{����l�0���#�Ik�_�q��-Y�"�VƚDC@���5<�|��T����S�z$��3�}��|$���򳨞�߯ I�W��b�x�:=��(�Bޛ�j49!x�P<)쒔��r��r�
�O@>x�E��0v����I��}�>�Ì�u1�Yz(,Tth���b�&�v�$��G��f\����V;�p<��Yn��I���^=��羲�f�����<ik����W�ϟ����ř��F�hg�0�,�$BO_<+<4a�5�������2��'�~~ �㋶�y�8C�%��m�ע�3����a�8��� j���i�HՅ/�K�f��Y пr����,&��!皡�I�U��ǟ���Y�	E��gPeM�Z�σ E)����kb`�|e6il�i?�f����� G�8X���'�CWK�%?�����j�t0�q�ֱO3������w�Ծ����0��{E
S_��H;�z��+R�]:�xZ�0�hQД����5*0
�����&;�loGDn�ھe-/-?<��d�*5�Q�\D���Yc�80� �K3e��TW�Ϝ�9��TJOg��:H�>eRS�G���s�j����
��	�Va�z���l�4l2Y�J�,SJ�FPy���L����z\���|�R��!G��s���ɚ�}�	^���a5���)�K$��Ge" �6�s̑�;,\	*مЎ,��Dh�=�/�N�{�,;N Uz��R'���퍟2IZ{�.I�ep� 5��Sui�3��{���t�g�n��q��
�Ie��I��؍g��:�5���7�I/�*�[����U3����*�	���dYN8K���-^\ �O�����7�	��1"F�%���K��3�*v���R9�~z���ε3캸T��rB���K�*��[􍶠}T����#u�g�>�s����5�`���x6Ή_|/�!=����P2���BNt�_̝peV�`�U�_����6@�����S8Ű������r�:Q���i�l�`�Ȱ@�罴��E��'�%iy,~�_w;�	8��"����d�J.�㐀`�Y/{��$��#^u���8Q���� �8G'M�4�,ɱ��R��L�Ŭ�e��	c6�c���b�r&��؎��6�Ѝ!S'-.>�W) [8ZGԡ�(�{
gY����2G]~��UH�p���X�����}kfDt����'vY���%��4�yc�P��2�}�I�Y��ZlN�/�I	fI�k�~ ��KH���v� =�����Ni"n�q��Z����z��T��y�*���c�j	a�fQ[}z~���G�c�r8��P>��c�8���H��q�ꦘ:�M��R�6��E�°cbAG8y(�)�x_��ELEٰ���8��*�9���ʩ�3⌀Y �ؑ��	b� �}��*M��8���5�"�����������3��.�d��I��V��0�r5}�[g1;���C@D�\�H��[WhI�aB@�lSNM��z��4>��l�+��1*-5S����v9���\���<����B�{؜i��������z3��g��4�����Ԁ��oR`�T�����z�dh,K�Ǥ�<���5�]WA���	�J��Μ��ܕ=(��.5>_��K�p���wi2O"�d%�8Z�ve_��&W���R������j^[fXD������j��TnU9u{�P���U����+gx�lDz-"1M���������vi�|�5 �-	�s�gq���Ct�	dE�9�"h�˖�$Nc�C��Nm��{�(}��A��s��~�������#b��er�	_>ߐ4�0V{�#~~�_��ۊ5��ٯ���"x�|�)��]g��I��Tj1S���:�VF��o�	�%`[M[�k��(=k����U��R�$��7tM�s���Y���G��0t:c�Y�"$���� N0���]���]����̡��L���
o�Z�J+���uh���/�B����?j�~u	�����51�Z��u��B	�m�2N���ߎ���ʋ��s������1�r!`vV&����'	��E������y@�7�C&5�c��wt8�rn��1Ѻ����v�~j�{z���K(�7 �C o��f��(CLE" ����(jP���/KE�1�ˑ����ޚ�+����}�\��(&�,�~��DF�2��W4�H�b��F�˞q���BE	����@��M���Y�p��0ǀS#4R�*�3+Xa�%��#�M�w)���s���üSs&zrg�=��]xk;ҙ��F��,'�PC@OnK�E�H�R���a������q�7Qz��ɑס����c��T����V�:��!�k���`2�3[�8xi�-@�B��]_v7���1���3�&�Z��O� h��!��SIw� ��_'��2�pQ��ţ�O�\%�ך�.�CC�<����s�Zo[u��{~s�e�.�����ME�T���� /XF~H�dm�I%h�ҡfa�\¯h�v82WT�t�GQ;�#_P\�0���P��ɟ��BB���LY��0�z��sGG0��.t�r��Q��I3%yE?t���Q$�s�B�
�Z��xn���Sr<!�A�d^>��
�p���ޔ�tP@��tƭ�T?]ڙP�T�Ց�����*�w9��������6O����恠��GcD���>�,CA%� Z����E��;��x6�>ĝ0F"Ǽ��c]]��ǒD_�MO; r���F�u�Մ��N���?���3���s	�%�G`n��τ�,lO=̼bF2	���eP��'F��m���H�U���S�� a�x��.j�v�;G��(�h����KoM�1I�ơ�
�|��QV��Dc�/���_��w�&��2�ԗZ�1g��<�7�Af*P��������Nw�"�6Y��P`'��s�{�����P�P��jL������	A#�@��Y��M�&��?�`Z/���j�)?��参���0f���zep� �钕� &�50�W�ˠ�~�m2��oŘc)�˥��HQۨ2Jxt�a�^�)�l׌ ��J��)�*{��rӶ�2QUq�#5@m�$�3�NQ�q��O�b�Ί8?��nC��]�Ewu�����.z�F�����{(@n��nn�D��@�H!�>�}f�E
�3ː�b(C�KwP;��U��c��
b��W̚�XW_�O�k�i`�$������_�g)d ܙ�c�z�,��x!���=[.�$5�+G^4@�7�aܥ���S� _�h�=%t5��Ǚy뤢~��X�J�p��ڈ�m�r`�Є���T���谽kt��h{0	��s�/����Ku��d���о��i L��d5[�����Ȗd�k�(��N���~��-�k��1������=[��?'�!3[��v��Ɛ �9�-�O\F�9���uRG0�3�wO��xj5syk�/��$4�7j���y�,m�8,I�Dj<�[�~{���J��=�`&��ee��'/(:&M�0�+h�i�t:=��˅�Ъ��n� ����_^RM������aCu�������'��f�?�"� ����;oH��Iy��vjjF`8�+F��C2#z<�� ��'.h�Ԯ
�W6@x`�����p	�̅"s��'�X�0
1���?5�K��Y��PSԫV�杫z=�S�û-
�8�݁t:w�K
3J8۠�������~8@�$��&`y{tVh�H+�S#���V���� ����f��á���d*�8X6�
��422���p�r��L�)�mauzBKh����v�>e��;*l�F:�`�,��0B�i6�9�Z�!�}�9=����e޽�u���.��m��F�|���Z��N5�gHV>����~�%�o8�T�B���r��vӖ[��>���95�\g�Nv�H��X�����AYi؟;�:�.��XF���(��M�m�\̜�2��گ�Գ>l���gN�3�v=�Fy�� 1eN5��6!��>|.�":����x�%�L�P��;_cr;�K��V���=��.ܞ��"���E�Ԁ�tGH�Z������iU�81���dQ�J����2��4�{e�\�� +��۴/��	+w�xNz�l��:0[ePJC�i�KA��6��ϼ�k�坯���sNrC_t�ǯE���D7t�F�h��֖`��(=�\�_�L���� -#nWf$:J-�7 m�2΢P��ͱ~��U�G3)�F&�[�4<��t��Z�u-��MT~��ê����GQGK��w�`Չ�h𯜨�v��r��1?��Gt'x����ǫ�e����:5��S%J���t@�ō��¾P(�%��8]���Vџ$_o2?�蒻�Rݰe��^H���6�w��缣f{�W���/�L)�'�+����+���� <t��s��>pd�p_�b���"��)��D'�W(֫np��Ҩ��)���VjAY����tߥPvx�
Tu���������4\�"$j"�v��5E�������D���̨;�U�t�.y~��EUv/���	\ʽ%���^Ʃ�$CD"�WWk�	s  �/;�6��^Cǘ>x�fݺ��_���O�۱���:`��)��~��?Cy	��~��|o�S�M)��R���ωb�Ϣ�қ�_?
r���� �"]���s����#����Ǧ)D��r�M�I��]��klBga�^%�y�R��B�Ot�1����'tx+L��a��8�'�9��������v��P»���g�h��U�@̖�u�r���a7�8�IM�h����iX۱Fz�����DY��h9��T2k	��n��>��|W/>'e�"L 'q3�u�ꌦ��3,�w`��S�����4�%����O �4-�a�Z���<�t�-�&C˃��$�|u]��4��8�fr��h�^\�N�/QY�US�?n
�EU�6�XSzr�#��m9�=��E��Ҵ��'כ��M�+�A�ha�n���*^Xfn�{�+6�d���=&Iq���ӈm�����$�>�K�z�;`� Kt�c.�n:�Ί]{@�`]iZ��m6�c G�nI�u煔�������a���~o�߼�ZsP�V=P@��������S��zGq�,f=_�p�	��O���-+�{����v
�K����u9�T������T*��11fxQ��PP��T�F���?���W.ڟ|�XY����eYò�@�N�i���~p�lGSd3�w�-;�JR�ïy�I�O���,���P��zoϭ���3ޮ>��Z%o�!Հ�����-�=�k��y�NtH����Y�	/hk$�mV�䳉M�mi�\�+z��q�⬻4Џ���u�큏w�Flb	�z��ic��Ji��kMJ.���/$3&�8;�rJ�0V|��[�j����W�֯i��UE\O���fO���)Xhʷz>}��q�TQ�Ѽ�Mg없t'- Wߙ����e�G;#=�����C�N�S�p|�֚B\b|l�rMD��+��-	,����f$�r�M=oi�E;�d鋕�]م����WU�n[�S��8TZ�����X9�8��ul�}e�a �B��KT�b!��h��E�1�iJq�o�.����v�^��Q�����k�y4`��J�  8$�Do�� <�Q(�q"�zC.�Z���f5��3�K�1�vl5D��������!)���X�kt��i���$A�n���[YB��$���8��O$�xio+HBcg=ڧ���;J�\ �)�Q��l�����y��Hl*j#�~8��oih��bP}�h�1�@Dsi�Ɔ�׆��-i�f3LEQu��YjAHt4��Lws����N�����y�u�>������Ψ>����cOb��a"ː�D4�8�c M�,�e@�RSA����s5��!<*�U�.r�V�:�~�s��B�D?`m���@A:o�O5J�W7W��v23����sҔ��� ��AD���X�<-?����fW�~�9@;�WF[�����*�i�6��s nw�~�������z@�k���9<'h�wG��ن�:L��̔3�2P��p���C�i`�W��~�dO�-��D���>�a2`ޫ�y&�[��l��uAn��w������h@G	�f��p1�4��O�����[;ZP���?E�*��q} ��@��B;�\L�a��<���j�k���f�����])����gj�y�I�Ԛ��0j���'擙�j��У徿v�ό������i
DM�_c�y��V�1c�ڭH<,�s�ퟚ�L��Wҍ�;���&P@m +'C�"J��$	ӻ�=+�N�\�Qm���F��w+��R�j��?�d�Pu����� FVw���ؾ��� 
�3_Q��]p�-RKB3���T\S�l��v���Yԁ���J�?>��S� ���:g�P�~"�*ۺ�ԡ�������0�Z"�jB�C�qP@��.0�$�Jw��J��V}�����lVK�v�Mk�����5�Q:���E�.�4�u�!T��(X^��~@Ev���p2�S�	A{r4��&����p�%]Z�\��B�9�/�'d���A~��>�-�̯[�#�I�D�������Ӱ!�
��z#��&�WD�'�wZվ��������u�$~"AP���amHC ��R��v��x*V��>θ��8,x��b�h_h�|�����{#)�l@1��q$+��I;n�_�_s�>(O�i�`�ȶU�_�oxL���T��R����8.�M���_;tr�x��{t��ß�/m4�����lUgɲyh[�aO)%|�qI)2:~���}�L��dp���NBJ��|�2��*PfE�g��<�~S�J�ۨ=�"�[H�8��N����wP�tQ����	�h�8G�TI��Eq&�ê�*-�qs��]�e� LZ�i�n�Gx�"�^�8�����y��x��t�*�ݠ�ݯf�I�)+,���jg�Q�,t��K��d�
���?�o������%��,�s~0�>M�� �<;�������|>?_N�c���K�oŪ�jXK�yrqꘊ��lYz�{@�u�v�)�!��n����>��+�1���Dz="���p�^���	
�bIYQҸ�& �ZZ�\���(�\̩2�9�Ǜ�v����wi5"pH�����,4~_��.P	T���^�_�|h�[�s�I�x���R4�ZEO@X��fF�Md8+(�3��ŧS�9Pb~�y��U�C�lR>O*���f�b<(S�����8��c���Q�{0��_?,�T���8O�e��+��.�J���z�q��²�y�Ĝ�I <��Ph���[V�Y��X��nR��)�$���С��&`��%�j��/97�8���B0��3<�?�΂�M���� (��R1�j��:ͷ/�߬[���c�iWM=4�	���ivؗ��]bZY�����.[��PM͸���Fݙ�?Ӯ�-&81=!���$b�����.��)�͠%�8 o(��,�{8���}�3�ϝM���1w�K�t����-��0���<������a���}�/�-�,&���#L!K7�����csly��_l2�¡�����2~2r��Ȭ5�-R.��i������86��]yCO�4OZ�x�sU!�9�Q�kP�̷�"ɖ�D�����` ���g]>�U��]��qX�>,�:��8��U�8��"-�Za,K�-�>�-�Qm0K�V�W���TOW�56�Bx2��Ktj����V�C�zS��K��.�Q��B�O�>�%6���9wa=����p*�&h]�xC)������l���sw^䃓(Oӊg2�o�-lX!���{N?2d��%���$P�8���(�צH�v�/2�i�%�F��q����KL0/Me~�\T)uY�bZ�_
ZWMxr6�2�k�����AtG�̂��׼x��H%���hgJ�>H����;w�2n�bꬺOWW����(\%��ݩ�J��(���Q9�ޚ��5�L\��'��m_I_�sI[�����S���Sg#_�>2�v����c���8�z'����
����Q��7����e��u�9���]Qc��0&`ȶ��Ŗ�G�����N89^[ș)�͡	��F�7�_���O�fym.<��("�
p�D��-� ������.�a(��p��^6�,��M��U�	�!b�2ӏ������5��y���"4��c� `����w�L��k�Y)2��P��˧�r
���%pQ,S�@��M��|��C�^�Q����bv�\�COŠ�lA~U�!�A�l�~;j��/n��1�}-r�����uQ��U�	�� O}Q1����*��G�
[�)m.�׬
ń�j�����k̉�UX⣬�IO1Q���H�,xBɄ� �b!�fw��h���ja���լ��Eb�H��aMF/��Ƅ62d=�?:+C� ��r�|Z0�g�� 4_Q���G�;��\��ڼ[�DF��	�.�횔*����$���y���,��/���Mm,|�<5�g(/A�L��y��/������p_)�{�hHq�$�R���4�3o�Y�n584i�	LS�ͫ�K�ZJC�bW��m;��L����W�F�ظ���0�L3��c��\��VUo��ʄB���tjB�[�{M@��DL��|����i�φ���[/n�w�'�y9��ɒN[G��ޏ�;1j�DV��=�����XU"�v���J�u`�$��Pp�y��%�	미f�-�X}��΃C�����L����K���/_8HD�dgh�����%�!5�phgx��R��<�Ռ�����&
8y�3�W�(�v�T��MЫ=8¢�
9�i��lK�Mջ��2F<�P�ЭZ(@�>���=Y�L('l
�yRm�!��<�I������O_�����,Sg��wv�o�=##�!�P[��j�5I6q@n�	"��g���]�8��k��(�Y��*��s�=�Y��'
c�r��h.���C��Ov�nƏo4/[ђ�5II��Ė�O�bΧl �l�2�\cP��t6��j\�I��/�����\=���%�*�'�_(US��ꖩZU�/�!%��h��W�)�_	�&��3j!�zW}�AR���mK��Wؤ.�)��?�?�<%�ϊ���)*@)�⨗Y3��Ս%��,������ 0�Z*.�i�BA��d`��C����oI���Z ~^n(�Q��մ��Fsv��z�K�罁<>K\���soz&K)=��	�xdj}%Ȏ���G��Bki�.$�d�u�J��޺�1��oq��`l��.Zԡ��T(�v��L%�:%Fmp/_C�yxШ��辞���κ� �@8j����=>R��\.�M�F��������/��a��-L�M��X�P��'}����Nl��0k*�V�X��7iF�9r�U���>3�:�����mMԮ(��͘�����b��<.�կ,���ښaoe���5t��Ap��(�g��[EkTn����Ԃ��m]
�Z���u��'��`#�0�� �����?��k֣�m������g �e�y�A��ʀ���N�1�~�Q� ���h�6��v p�X��i�(�Չ�����4�O��m��ajdY^:�O�&��X�K�!mć)�:h!F��Ox�
�!!1hR�C���{��P|�t��ZB^S?��),�odJ#ˮ�lc� �9��������I�C����H��7|�&���{���k�ia%��_�!�D���c���D�D�Cq� �
�"t���cp9��yK�� pS"��MXFd�[{��G|���)�GB�)�ԫ؇)�H�(���ӓH�򅔹�K�3h|��~�b�ҭ�/ݲC/l�#��N�BV��|�Z8������s��:�O�*����,�zNni���ي��F�G^�#�?"��,wHА[*��8K�+?�f�T�-�խʜ������@�*���!��O�{��L�VyR��h��i�$J)�:��u��k�D�GZ�D�JpF�� �li��D�T��;lc38u�Q;È��Y~���+�n��<n=��	d1�M�I���3ѝ��{}�ŉ؋m������q��pq�_�f�!�?���
!~RU��@�Xݘ�R��Z����>�S�H�(v�sG0��M;=�àW���a�/}K��^���Ch���:_Bo"�����ל�4u���O��x�&��:�w�<��VP)�VPAP�?A����b/;1ȁX��ם���� J+�yxK�C���uB�D2;�.qPJ��Rg By&��<��w�&�]E������F����+����N���d�(�G��3SCA�?a��}���WsZW�g�>y4�D�NYtG��t�1�s$rf��F�C�:�*�ʐ���9ֱ�dt�6Qҩjr����[U({&���!�*Y�k�=��B���C�I� �Ό�����:�o�q1+aH�r>�W�}��B�~�]H���i��iu)�7�ŦeH ��yb [����$�����Y�`b����"Sj�v��@�<�*�܆���*d�.>VvU��t|A�S��ejd�`#v�4	-��
j� �+jb�y�S�_��F{�6�1uS�2���q��wAc0ɕ�8�m��˂%��M7�LΑ�htn0h#��3@�)��=�Y�v�v[�����gf�g�����}y�8��vͭ��;ã�(s�lkX�	�A�T�t��>�%~b�
���4@⻐���n�l���7��N�.�$of#��wf�e��5��n.C��X^��ۚ���^{?̑��k���0K[�w$p�8)5�BM�q+�<��M��*C� �+�}E�5g��|�ɈC���/�C��%��(Z���� i ��`<����&z��c���D���e�$�X���>��s.�/L-)M^��w�y�j��z�Mp�q�f�d�㹄�MJ�JUh�v�f_��~�|HY�So��KM�^BF��w���Ug��4��s'�G;W'���,G�R�
5��MlkZ��"���kQw[�����e��oJ�-�]��ti�%D��mlN���6�J�ػR2t˨*ʩp����<ޤ�Q�v�r���6�0�V����������+�/��ɐ�
�U����0�|J�7��F�wh܋�K�u�Ʈ�����pg�q�gS�>;}y܅�ƺ��������Gwt�S~��<HM�<�Б���3t?���G6X���V�����,��(/u^{��^>�_T��Y��v;�(p5�w���6���o��g�TxA]����6P�C^%5��c���pZ,�N�s�twۈ��S�wթ^��7+��TKAR�f�]󧚸��jƔ�'9`��<g�B6K���N�����#�߮�']1_�:!��ͼ|�ߞ�%�Pת'W!ﶘ�x�qv���L��G��r�����p~�OJ��xb��u�x���.sO���7bB��G�0/���@A��|g��taxİ�]�nN'��S�{7�D6^�����J_�&{ �m� �@>��?��8'�	�pYL~K�y�(�?&��R:�\Mw?q�s��7x�����W�8���e$݇/�`v�x}��qd�A��ͭM����;��Q��ME��-�w��N��Ӕ��т�)�����*��������Ǵ��1!��`:�������|�M�:گ+L�������u�v.�8�1�֩$Jo(ω��Mc�,�L����cxb�[�� �(9��")찔�|�b��5��N=�F(jC�K�\u��,I�W�0'8�/h'�v�oR�+N�t4�P7���z��}��."��*&�&�r�����s�I��29rڻ���Ɖ���}n�F���ڰШ�A��0�P+��T����6,��Q�g���ɤ�P8:ĆG�r�@�!�����9�O�x�|����ط�<��[�O�g�?�uP2��pNH͜���gUe�]J����<sC�%+���~o���M��R?�16M�U��"u��k	����쾻�M��fs؟��������\��:����l?-�?�[@c��KRb��dH��Њ��Y�T�̗1�-��A��"��$������t�b�S�S�>�� h�H�$f��bs48���U'��NT]�Һ��oQ9���=�D_��$��)��ʗ�Q�7kD�Cr����CЧ�0���i���O��z� `jD���W?6�����E�	��a���~�����������;���;��h�L>5`= �������v%�	������-�I DyD�]���#� �Im��#Rq°{���$V��6�JNH���� �媘�/&���vp�:$iJoG��X�+�j��-a~��0���	uɄ�+����-��BQ�2�Zl�./�_֊rDC�<���((m���F9���i����r�^�!)Pq��q�m�:��͡dN2(-��zR�|�fj�����ad
	�o��O�Z�F�{)�Y��2���y��]�6#r���e�f�h�S�MH T�@awD��s.�:�x��D8"���$�g�Ul���NnC3\\rt؞p -��9}�j5BƞV��+� ���p�y�X�Ji�&f7N��a$�c߽��r�I���'a\p�䩰;�J�Hm�L I|{�����&��W�c�0-�P� k�k�&�xLs\К!|�T��d\c�3�׼A��E�(�%,,M���5����d*l�r���n.����S��~dRq�Np��	�r#ĥ-ui�m�2���2u_��ѳ7����1O�"�V�|Aʾ|Rm�x��/�;�;�� �h��.Ɇj�������/X���?�<�10�4���2�5`%s@I�/���6f/��J����"�|+L����w^������7� @�"�S"yN�hA.��l�M=t���Hj+'?��y�	�0Ti1]��]���k�攱��8J��X ZKBC�!�{u�LH�@�#�'�Y�h;���WW>��Ud�|A��)G�	��|��e��J^&\~�q�/CE�q4�?�$A�p�c&���Ś��EZ;�e�m�TU6�_A�J�tj��F�^6#����5Q�6;6��jf/���F�y<,M�Bi&��vb�0b�CU�~愶��^������UN�I�#w�2�91�نnn÷�c�m�,��9+�#�7n�!z�k~�C=�3Y��_��I�YͲi��R��z}���9P>�
�2��]ٺ�*U^D�oW�����U���<:���z\{�3�/��П��-0T�/!���Tp��t���L�&�T��z�L��m�������Hه#��c<��	����$[����ݝ���_������5�^�(JPy�l�������@0A	�X�)�s�A�e8⨙*��G��9�)� ���!��/�8	:VbD~frز�͡!�����o׾Mq�]��"4��o
+Q���l$�s��\��5rWu+�k3;�y#,���ח�ʐ����b9ۨ�z�l/����5ύ�+|/S�n�jé�<.,�^�w.|�gѱk�X`}tM�Kx�0<=憳n*|�j�)��]��9l��+��;&3*��j��FB�S��.�����Y7þ_�}<(sr�םl'}���f3a��ъ��C���ur@tC���p��))� ؁'�h��n
TZ��CƢ=Q�.�A�1�d���${�'��V��\�CM��O����y
./��'^XD8��5&��� ѓ2t{��z1��k�l}_��_|[�f�wo�&�pYͩA�9*���)$P�Lwu�m�RȓS(2Dn]������CE� �j�4������l�/{}h��3n�S֣��c�eQ���]��O��-kJx�=u�穉Z�-JG���\,bT<_^�q� '"�W4��N�ΟE_�:ʱ�ΌSm,�����3��l�tϞ��-H�pH�P�}�x�iqᤗw'���?��V_���#oe��� �K���-�'^L�HQ/E��X��tu���F�|U�D5zE��=�NA'7�+~���^*�t�����'��cy��#Ү1��xS��6f���ξ}!h'�<[!�+/�ag5�H0qW��ٟ�2����o�^L�3J,
f��ԂX�AI�X�!�4��~�z�Y"��b鹲���s�n?W�!�Um�C�����s"�r�Z��i͝��K��Uv@�T�BNۋXF4%�;A�^V,wOB���j�l�|���v;��%��jR�����A���h�<9�-���\�5t|����X��0x�j�S	��!���� �$��@'B\�KY�"(�YC�;�*~l���+�?禍G6���Q�q��䄾���5K��X�v�_��_�#���d�}ߙ�h��i�z�K��hu>��0T�O���ń�_�����+p��X�A�SL��>kk����.&
�'��j�������E����'*�l�Z~a� ��D b��(	Ӵ�Փ���ʡo$ݙ(���n/J���	���#��gy%��F�;��(�1��N�����ᵜi�W�Z��W13�	gI� � ���ݎ�̶����ui�]��O=���c��x�ʳ�T�(}�.7:�qC��r���.�<U@�p�oʟI:R6�c���7u�?��q>S|>S�+�H�G�Ѐp�c��٘>�����2�5#�/����s�-��he�"��$�'�Ro���L��KY���f%�������: ^�0C��ro����km6`�K� ��~u�M�>���l����T�lS����и6�cY	��־lL)��)JY��E,>�^rT�k����׍�??sK\M��t{�_܄Lu�I�L��<�S�G�sԋ�v_Q`��ǲ���y���;t��g�Z�k%���!ElIk�8� �C|W{�
�%L/�0���FO�.�u�qp�+H���B�Jڭ��!�e��(�I�����ӻ�p�@=���7��Y�S�%��B�/AF:���	X�p��P�I�0,�K�\]���J�-��s�B�� /�@T��j�~smyR�m31�Z����C�*��ʧ!����ؼ"�`���Fm2���%��|%�P�ɝcB��ʺFU���(�- �|�3�&��(q�m137s���~h�����+�ٜ�������"A��/����$�U��-K�]���M]l�b�i�1m<��������r�I<n�˳��V� �$���f}��M����0�����b4���������v�S�0)�g0��7񺝣�\*��)y��d*<�}f#M�fS8�nh?�ޮ�"�ui��az�?`S�����q��h��|�����הX���f�k5��X"����.��ڙlW�g�d�c�m9�3g�:I*>�4���ُ��VD��ź2�n��߈��g&\��ե  �N`^�G��l���s��{q'0��O2��KB۳���!i)�c����
X��]U�^F��R\K[n�-�)��'�W� ̻0���d��!E�H�^�yaSU��7��R/[y{�r�K���[�>�M������%퇇�de��	#�0���0���<b�����#�	Ǐ��\�lt��b􈸹�]޳��hr�W��{ zo�/eB�pŁ׼�d����$o�O�͓�Xƺ��Q���S!HC����S/#M���������������Og�UU�Rtf?r��z�jtt|�[�o���C1��	Z�D�k��q3
;�v�
A(��T�C�i�F��=�Ƚ+��g�v����L�.�8P�l����l�@�Ȝ1�Hֶ�!r�V���t차,w���������9103+,�W�q���8]�C���,]\`��	�%~1w5c��lYf�&�Ň4����ĸ�ruΗ1��j0��od@���U���w�B]�E�)tM�Z��M��K?���UU�r�������2H�Q�����`�t:�N�������6��b鶣z�&���=�(���`O���h�.3���ڂ,k��w�?X��U���)��?b�,�;��`��|�g��߼߿:,��AoDa1ǃgr�p{Zu��r�|���Q�AD��"tw=�Q{���ͽ����PK{־��6�����#ۍQ�!�2!�omB�+)t�5I8�m��$<�Ħ����.�_5�p��bP�8A�����~ y����a���
�%���׮4_���1(NAk���gC�o�!��M�z��#���X�Lխb���,�������D�����E�<E�lZ��'E��xX.�/%�^E����#h�[	88vR�!�]`\��F��HP�A��Bj�e|#���2��͕'�h��Ņ�rp���&IB�i�r���x1�t10ߞs3���#�����O�.���_1��{�ྲ?�o �eά�_eb�A�,v���"b�w�����iB]�I�ؓSz�v�r!�tO�G�����7&|�>4|�P��V���^�O6d���iZ���>�=��o����yL��.s\(ZO
h
�g	��.o��(J��
X� ؾ7P(��"�:���-L<w�\PCu�S�ؕBH.��z9����KFi�im{"_M����T���j+�B��x��K�n�\vqne�?��K*����$_�^M��0����Zp^}��pi��� -�"=��wa����U6��179$�zӂ]	��w\�H3 uzS�s�:r�酚}A]�bR.��g���C>@��,$[�����Z��ETޖ�GyA��&f�Xv�������>�N����*3�K-,�
b'?����>A|�=�}#��IcЯnl����h����~�e�x=��}5�@��2|5�Vt����D��D�&y�2 �K/�����w��9,t�,�iH�&N�{X��S^��Pd��AqՄE��ng��O\�J���%�|q���c��P]y�x��o)�@Y-�+�w�\�w�ŭ8Ú�\/�^��}{F��J��P8���}��v�7��������Hʙc`d]�6jt��|�+��F�����M�t�U����� t�p��� ��D��U�Nj[��[�0
C
1T����niG���ҁ�6P�ٻL,>�i40o:b������d��~%��pʈ_�\�<4W{�tu�?�U�����oҍ=���'yo&?k����T��3���ψ��j�e\W
�3bM�FQ��Ci!�lj�������oj�Ċ$��D��MS�|l�V͓(� ��y"4�v�����]Zb���c�Uc'�}(E����1��Dg���i��%#�"7v��n�	[s�8�(!�mQVҮ�.��W3�NW����Pu�ݷ
���[��2̎���LW4�g!:I�+ig���W)�3�؁%�1^�
ʽK�裗kN���B�� �����M���Х_�����a�9B���t\VLX�~��5�1�����NV#Z#/̥+��@(�c���,�vb�Tj�O�W�M�_xrcv��xu$�v�9�a�aߏO�S?��I?�*��lV_��@�9���%�}��>�9`*��8D�Lɫ=="a7����ՙ?;����X�I����A��_�7��#�p+��+����N4���R�M�_>$���$=�w?|�C��wS�Έ����-��6,�D����륥�:�KN��p�1�(�ۘ��c$qѪ�T���wh!F�3��*�#Z_�x��#߿):[�[	��$��^zT�J}��0�A���轿ge�}�r
�*��e�X����0υ��p�/c�@�%l|Uo���a�P,}�I���gKd�3�U0��ܡ��<�<K��렄j�_LB�'�[�p9�6
�|��j>#�!�ת I���m
t��J�T3�͈3rG��__b����8�c��Ύ�	�%���\��f!�&Ǡ;�_�T4q�2_^*�0�#�M��;N���gz�~�zЊ� �Ѝ��ZjAnE��՟x���X��;�)$f��~�\p��߆��s�V�QxK	���y^ԖX|!g<@5�j㙽�SѺ��=a:��q�@Zya��K-p�OPl���~L�^IL�3���;=�W�h�ăj�ټ�J�8Z�V2�/)�:�����a��������D�:p��#��
���W�A�E.�C$�N �q�И�9���oy'n��QR��D�'��or3����\�>F�i�c���)�b|��h-�������J��c^uT^�[�pɗ�)��AZ_̴��!�`ƹU��R1�?&	�^=K��Hǣ�6��k�p��b����G�z?�r�}q� #@V5�;L	��ɤ/Ձw��"6wk2�>��ig��8���
}&�>J�y����n@�a�4���Q)�*
ѯ��0���N%T�W�@iYR��=RW�tz�E(�²Z<v�ҭ��z!α%j9��μ�p�@�#�I�NIg��+p����"��?4�f��~e��K�h2��4,������(����J��$��V�H7�IzD
�vu,B��Ї����: ʙ-��R/ �6t��ٓ�<� �)6�(�v��X#HD��2.��s��8��7�ʆ�N�L�Z�\��4_IH��:Udpې���%���W��"~|���Ԩ�ppfڹ�hJ%�4�Y�1��j��B���#�B'�$X!pi�T5O���U��$
bE�X-�u���(��J/�]�:���=S�)�� �����ul��tL�:XX����w����׿<�_KV>*�� �Ϡ0��q�M��lb����h~ʇ����1�X֏9�VΧ,O�Z���'g��?�17q��ݷ���%8`�+?��gڣ2����;�s��#���K֯A�჌^����BkN���I���1�p�P�eE�O�����Cq�*�g!p���Z髞�w2�cPWyB)n�/ܡ�:�ۼeȝ��
�E��Zy�5�p�x,M�����ᰆ�㏄KX*�,�����F$�\�6ߊ ��k�v�x��/����6o{�OtaÊލӻ��W�Ɂ��ˢ�>>��b ��s�Ď�^v��$ͨb�h��J%�ډ�\o�H.i8�!+�p��ƣ{����$Xy�es�~���ާp� W��#^�Ԭ�]E�ظE�H��4�uϏ���Fsb��j���R8��p��N���0h*��Y���xA��e��M�pT�I�u��.kQ�y��E]Xǃ5z"�h��9|ת=U�~I665lk�>�&��d�7������ͮS��m hG��q]ɏҘ	�t���l�8�����>��O��J�셗��r��j3Ca5W��]�{�ti�G��Vp\���PwO�v�ӱb:�4�n`I���A
M���S���\�-`�3�1���MtC͎�0(������
���v�X'��:�Bg��Z̕�� =���̈	Zp�_�9=/�L���Qj��u�%˷��Ҳ���uc��Pa	�HD1��bE)i`����\ռ� r���l�������q��:���5A43J���<M6�L�)���ĮP�~�N�z}t�M|;|7
��m�׊Q��>�����v�B֢%;o	l�Iwr�^�|�����gd���e?�v�/2��^1� W��K4��ata"�&����:\1����:_ɾ$��_Ou�������9Kv�Xu�jV�	���Zp{T*L{C>��n7�k�ܻ}�X����-�+�� TED��]@Y�K�v5z���4 "N'xy^=s�������B�=���{��E%��7����ݿjv�