��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�]d�L=3	w5��?�N��A-�5�P����B�[���훋�^b�sG(�dt�.KR��:z��X�X�8,E��c��DA��G���\�9��=�����*z?��'�]?�VUv�.���Ԩ0���L�sB�Ξ�U;�[�B����gM�1�·܅�̵�$����Q��^����W�M5�}�<`}�]مڦx�|KW��(`G=2[�'J��m����5�E�0�d�ܩT�I�f�[9���wt��f>�eo��k��F�����Z�jz1���(�+־876�����O��|"��Y݄v ��#�<�;�dWZ3wP��3�Λ�v����6ě�M6Ш]� �ಳ \��+��1��U������
����$8b� 0h�H%˂��>�cxf�T=qE�Dʱy�B���	��cS��4���f#�7�i4�(�t�l5��,�/k7↢dK_�$x+�}�Z���]vr������'���ٲT;e2-E�Xi4c'TŬ}�<��o���<��&�<*Ȓ%�w�|I� ���b���	P�W�HM��Npsl#E��Ÿ}���D����|LXr��E,&��F��t����+=�,�Rtj�,�:m.)�+x^G͕n�;^�3 �&�R8��כW,r5��r���#�i�T�|�{`� ��lF�/�&nZ&�d�+�)��o&�п��TEWrꖄ�w!��bh�����$ˑ�b��*Z�!�lȽ���,��D�['�v������SC�y�V���Jm�	�}�᪗�I�G�K�-� $�(;���L�D;'�;�JcF���Aש��yzRܴ�)@N���rH-�d�=?��g!�]��b����TI������2Tk�`w�e���Z�ƚ��]#�2��&0s���(��b��4��yT�W��Ρ$CX�ER���x/a�A��$�x)�`���+�kтNr�/}��x?���1mL��/�j�A��Bq�}!/$���ϒ���� �``�{(�)�Ծȥ�9�<c�ND���B�Z�>����:����=�6���e)��]���n����w�2`�E��j��U�a�g��\9�^��hڢ-��V���8Cp0-��,:��=m��O����yr�w�Jx���\Lv�<�ɶMH���:O��S�tîU�!<�f���M�Y���n��%9?�z���Q#�5��x��)��O��v2�zW��r�d��)@���"���B�S3+��3��>�&�̭(!��!H�����aM�!=c����<�n���vc:��W4�l�#W�� �w;��z0��(��_���ͳ�=�[l>vf����9Q-�e��U��}4&�
-B���ц�~,�#���3>}��	� �ij<�h����E���AMV�CT�����9C���w���^@0�cNLt毉|�2d�@�\����΃�V+�C^�ՆȘ��^0��Mjy�>�[/�*8cz6i�����n�h�91��)��TߙU=Qc9��9���A>X����G����D��}X���Ir��N�?#�8M�v�v��Lh�?�cd욹I"�dD�#�6�:�%a�|���xamQ���B0�h��$w���k��^�$��٨�Tw�o���m�Uj$�y�m�s�i<�d�в�?�1z�8��S��s�0��~��� +Q���;Jl����;�I�?�[��lJ;�J��')��K�WW��l	��9��=q(i����z^� ���ieL�ɋ>�2�+�"-����@d�C�܆l��v�䙥��+:��\�8Q�]&��0�NfY��EvR��Db^f�h^�f��>����Cp�z��Rw�1ظe	�Y��`?�&Le|:��s����kQ8D�ף�{鋜����+��X���Ky�=��J�&tޱ��Z�����L\��f-t��F���O�&�#i�	 �Ӧ5�f��@�8�OYi.�Vpp6��t����>�e�+��<�ֺJ!�3&e�f��U�߭NpF�Ng����tv��m�������e-\�x1�c|�t8�@�X��)��fC�_����U�&��y�0������_i�[L$����/�RYNഔ�)����P����O��*/�؝�pA�m�+��k%��P��ܠ��ߚ ����� �9��g#��f��нt\e���%k��Z�@󤄃���2&1{�9�z�G+�a^M���G/H{@FH\p-X�����e$��kc[�pMFI�=	�#�+��oc�u� ��k�&��zB`�<�4�#f�
��4J�� ��^g�(C�0��T��?�ɽva`����l��6� f���6��A�=K�����6���_����̣j������^;2��V3G&x�^�Ʊca���:,�b�������bdT�h�H#�S�Y�lp{���p��=(�*��b��&.�D�&P x8��ğ��YH����;�.�֯\�b�V����_�q9"�Wd$�/[���>���"O�LV����K}TH�L�0�����*\�I,�B�
%�9�|�N�Z�(g��N�xݿs����&j)/�m�L�	`����x7�z,��iJ�ʧǰ�E!�����J�Y��I��a>�!��ʤ��>�*�/d���;4���ߜ�S��x�1����ST�E#�ڗSx�r��V�=�I	 �OU�����
y� ��swȁ�Z�erqM��GT�<v��>�ߔ\oAnx�2]�%)�^ykTE���9f�����ѥ����'������}����Z��ln���rw�d�e���Q`o倦�?�؝⧻ڨ~����`��,�8���2Em���ʃ���~O{�M�+�S��~�|y��
�\qr�fg�:y^�:�r�-�S���`�|�4����o��V��N��d�_���\h;q�Nq\�Tp\� ��Sc?�"��l����s=|M��㌻i?�=�,�����`y�<����Z��]�����Sgj;�絋�*�c}�y�����3^�5I��)��R)��@&����m������U��LpK�$h���0]�NI$kMIŠ2�N�}S0qfr#�D(0��8��3��<x��8��A6W���`?gJE,HA�����{����	��~��J`�9#T
@��c��qZ����$9)	~���W���6$�T],�1��	ӵ	"�:�ÿ�71?P'0�yZ_Y�"��<+���Oo�~�6�,&_�\B�h.�kJY����$�:gsKL7`�N#�v�)�[�5�bmES�����5f�	I�zύF�c4^��'aB�8$6lϚ+gt4��Uf��<Ӻ��+"���J�>Nr�X�Rt�@�{�������+1�g�{4B	}Cv���
���i�����;
����p����'�Ԃ�,�B'YiX�eAy��^Jɹ�[f1I]���Z~ZS�*Ʋ�BYW�;����?A�At�=�b� m�3�lΞ���C��'�4H�aA+�#
��txN<V��1Ȏl�:=����}:���l��܈��S!��Kx��c�^���{=n����s�(�SY<D�hz��=���5�3!6�-rn��,Y�}՜m!5�J�[Υ
��1@���
�4��c�Pׯ"��m��wh[�/�:f`��s���ٵ�`Rn�"!��,]���P%���h���] ��G���{��>*Wj�#]�l��q/s�A1�;d�b���[%˺���h��{��!U�1���D��A�V{���JQc�k�B�xNRhM�5jɡ�b�je��?�~�_!�'ࡇ@[	'�t�U	;�xF�]{�UKJ��qF���@����.���W��l<K|&Ku��3�F�2�fS�fiU�ͭϰ��h	��r�^�{GWcIa�������הR�������u��
.�ߒ��#4���6oF��y��ԋ��S���o������$8��c�� �T��6/��ѽ��8���8��"�5!����LgU��C|�٧dzz�̰���D���'����S��S�g��IO����6�/-?)-���X}O���� <i)	��~�ı����nI�ueܤ�n�!�����,S�������9�q�?���`)��6�rЀ'=��@�H�H��\�Pɧ'���%b��ڙ鲔��?7H�&L�W�%}�M�;�a����h$c��ad�^фX��Q����s�.	~���t�LYF"�(�[�D�����@A�rjiX<�A���5��-�~��,��1q�{�n�����{Y1�AKs��g��X%��'#x<�8]��E,�����bX�Xh&���O�6�!��ܮ{[W��:��X��	�G���%x
�-�	v�B��/��q��tB��j�ۀ��~�l�FB��y0� �ϖ�1�Ĭ�K���c��wD�����O��ݎ�+R'Y�cƆ咝�Qc0��P=�)�&!"��ސŔ{zd j0�� ��Z��"��b�_��
L������
������7��W@zZ�0�#�MN��R`�̭��h���˜�S��3`yp�qe�ڒ�����.�\�%R�ԞS]��o�I��V2�I��SX����w�MM_�f�E��T�Ƥn[]��h�A��O����tC8z�7�N��;�<	/�17T(z�*"W�����욧׀�oy|�yڎ�� A���\Q�G-|l{s���և�����)��9��4���u��j�`Wҷ2Y�moT�L����ڹ+���k~���8�Sit��e`gQ[{�a�Q�r��c�9!�mmh@��í$p6fB�t�KTj����-�^��O�(�$�˗��ay,
�]���N$ 7�?��ɺP���\���#1����^���F`v�Ԑ��K��˲�� M�4�l���&M<tȜ�������!�::��;c����i���;=��:i�Gܸ,���k�2�T�x۪��v�	8��*��:���\O��:���Ӽ5���E�}a���_i-�ɜ���gA�x�2̊14�9"�d���#��Y�\���e��R⸵(^2��o^/��V�B��3Z�$����#z�^1)��$�ŉѬ�Je#�r�)q�v��Zr�S��C
�R#4"[^��҇�ꮎ�G��g�b�&ϊ���>1J�����r���m�}D����B�Q"� NZ�E2�cklW�?�/w�U�;�٨"1غ-;�`F�m��x���#%K�[j*;����s
�;_V��>���t����
�)MX����vθj�'&�\���^(#kb��N�)��2*�4�=��Q�Y X�\ܐ	��M���*��l�6�ȣ_F �q�q��{�"��6����`����T@�!�M�&C�������p�B�?��&#��%���~4��7]�,}t�Ad���~E�o�~;��� z�Y^1m*�T�Y���BP�*��-�Y��y��^|�E�7{�k�W/1?������O诱)�6�l#�f��J���r�!����2.���c����������t�r�iio�X7�'�-?B��LrDm�����(���R��[����4j>�ž�E=~R[�FӦ��y
���*��3�s�0
��Ȑ�E��EV��pU�hC�)��=�;�����h�,�R$�䇶u�~�����V�7�GH��n9�Z���kk���ߧ9�>޿Rێ���Jh{��Y@a����6�Yɤ�@�j�m=|�l�Y��ܼ%��O�R�a���38H6C"Ih&	v�����nҌ��ӏ�58�͵�G&�"��8��������=�(��Qs'�[���G�����_F�^�-���Z����<2� 23���>l�0����+�[����W�{�3"r�������Hڧ���fcy �*G�����+��)��j}٧Od{��GR7��>�����{��j4�QX4�Y���:H��AGh�|P@x���_,��r�יF6�>}��K��Q�n�b�|�X'
a���̣ZM��}ÂP�"si�!��Y�?u��q� ����H��D�(:/�Ye�]�&e�7�lYW<��:?D�}�]dUA�G�p����@�D#��T|~B�X1MAU��ȫ?�I$26:�o���F&���N��Cܒ0���r�U��5G��6�ب^�G|���FzV�=�j�R�ʺOV�gr(��!���9b|syv�c�g%�S��V��}��L!����Ǿv�/̧�y�Eϫ��#��Td��=-ӝ�y�b���UG�#��%'f���J칻C��/�G���������|�V���~XF�!���.��䊗��mx)��8�7�p-�n� �l9Kl���I�Qu�밉ʈ	�q��;���}��j.��N�����]��ƨ�e@)G���d�h�Ϯ~��)��b7�#d҆��7f�^1�3Q�v՘��
o!;� �>��iyP�"ߖ定��Lh�2�Ksc�ϧ��u`=N+h�(M#(m��6��N��ӓ����@�x��./�����dZ���dB�L� �&�Ņ��6�qh����S��:D�w�_�r����_�v��Q�2�j�D�����=�r����9|�$�W� V[��FqT�d1��̬���<P-���;x��Q%jr�ʅA�E���؛R#w� O<��o���ّ��\'�^�a�=��ZnV��Td�Cz^�R)��,�{��p��W$6�)��X�U"im�~�9�s=�%4xV�)�X�L(nj��c���E�*��LӘ�iZ�s,�6/��p0�iZt�١U�$0%�l��3���A��</���AoU�szj͎~6�J(�rB�{w��T�O����<�@��Z��	�O���l\�2@�1�v����LbbF�wC`�8͜����*T��@���DUo������T��	�ʹ9���ZU+a_4�߈��7�G
_�у�HDG`핷a+��w����
�������=+�;���b�f
�#	6��j�1I��_+Y�R�kf~2�fK�q8�ƕڨ�g��ȝ�&�����7�-�COO�r/�0���2�%C�
��I�܏҂�����!b���<�BK�����e+<�di�&���En9�Sb�)_@[A��|��2��R���PD�F��ǌP8�M]���|�o~K����,I�ĥNT�C�K��o`���ڦ{G�w=�����=Y:c�F�J:�s/T�!<�Y��<3�A�MYdK6-`��լ�ߙ�8��{|9K�z�R����$��D��|Ly˳�����Q�qS��"�*ԡH�����a ��'@��²9O}��0���i"3]�MJ<"Z�2���s�g�б�p����f9�\5�R�iY|��%�G]%Q�t���53ϡ�l�+��vH�x\c�(8�	Z���?U{���;�p/(P�;S
��!h�� �ғ�t[��lj���{
�'>�%9rE1W%�3h�Bד
�d� C0�i��۰O⼦���)��DV�+A�E��LY���N�l%t~;�2n�E���(�V@B��ѹ��Of����X?ո�%��r���l�˭#M꧌���<��]�9�@X���\R��u�]�� >���`�^goٗ��!�׳\Eјw������V�6��\5�v~ �Քy.��+�mf#���n1�6�ѦQ����m_o�4��N��9�u��4$�NIO�oc����NTl8��h�1g�4�t�4��ȓGx�����u"g;�
����;i�Z��}W�Cyݑ���C�x�n���G.m������)	TQA!�)
�B�`����#a�A��v7ß*�7��V�Id1����R�\8G�w���t�r���#mo�K.�_�a��#�[��jCv��~���vn���+�T���{��t���z��/�3��|��i�G�\h2FCuHg�fY��!_��a�0���"������uaH�;O�� ��ػ��F� B
���]u٥:�|A>��I�i.��m
��`��"����;�~Ӹ���.����&�ú�k��bM�j���N����/&TQ��`�}:�E8aw�v��ڱ*ss����4r^S�Z�=�Ŗ$1�G�,q-�g z�����e�������(���H�W��ō��c�R�`=�� 'U���>���Xw.�C�i�f�a2)Ͽ �)����/�T+�M�l>��~�&r��[�Ykar��T�
:����9Ȓ"cO�,�C2��O�^�����
)�/5It�Qy@��nrG�W���Ã�z3�r'���g|����7�Xy�#�I�f$�2t}	@�xlԬ��~ˀp<�c.��$�%��Eb�T �J���Qn$����bǑ�mc���d��~AA���Jf�q�,lDm򺰼ipL+�f�9�= dt��j�]N�:��(�3֚��F��,���'kX�#��>Md�$��;�w���H�Va)R�%W �@�������j	Ypg������Q� <��T�<Ǽ��|^2��Y�u�ǩ���L� ezw4�4���G����O�ܻ�X
-*է�(��%��`��y�`w2�m�3�ie��O^�'�h,uE�.:/�����s�:���z�x������~�Gp)��l/��G����"�q�w�?(DT�J�0S97%��2|�E����\�Myx����%�q>��4c�Ky�z
����cz�}�2J�X��I�W�Z�QU�Y�R��,�4�N���2P���U�?Jq�"t�E`�i��_�E@���
��v^�?M�6���[g�'>'�z`�������LB�9���_1�h�k���M��?�&�.#�de��*o�����A�2�{�n>؇&AC�^+����rPz�H�|�v�a���_Ҝo�3�BQe��L�\�m6��c�H�䙣��L�T��oŭo�
iLe�ޅ@�z�/0�/n_Ff�s�[��ơ�qB��ԬM���h`���Tٷ��]/�ܩ�)5��G/쎁A:���}�5K�?45K�Ӣ��!�r�|*�S�0���+9~#u��7N�<�Q�G_e4��(+����P�����4�F	)$���$��7��_���Ϗ�(gbD�p���͛^��n�?ׅJO<�pˉ�q��sl��j.$Z^.+�c�(� '>���Dv'gW�@A�Os((��s�gᙀ>}���P��vY�q]�`Eh��P�q�j�tG�.� ����glѱ3��4�򩁵%+"�2�q�D,Є�LU����0#���#,2�#�6��U}����"�\������irk��Jm���Tr=̑��$2���Z�����em[ߟ>ǆL�G�0]��������3�@�f o+�h|����yƯ@[!U:��D�B?����b
g�DE���'�@�'$�@|F ��ª��F��뾝|ͨۢ��,<Pp��FdN��x1Cm0`�<zF�Kyh#���9x��G�lo��E�"Ǝ'�����C� :����y���Z%�=����w0��aZ���#)T�z[g��^nEf�r= �Ofq�9�Wc���Oyht3k��"R��/  ��u�NsM�W�*���~H\�;KY�y��l�����>'�`�AW/"m`�!����[��I4�Ri�bI
�������Xs�-Lk9Ԓ�x �C[ � [*��hӠ�}v�(������9F#�Xe��I���m%>L�9���=>���'q�����-Ϭ�y�0_3p�y�X�
f�dv���Up�_V���]�\<�he�e�78����.)����Ua��`�n���������X�m��Mfc�E�AJ�"x�լ�qN����/�b�j��W�Z��xFB7
.\��#��(�R�VE�!��ċ�����9����IY-�+���k|4	ro �.(��Z+:��}��tR&�^W1�԰��6�]	��������[���:�ƴ�Q��x����)Uʌ�.�e��J��f�Z���Y��_�R���d���?|��9��Lm������4ž�����IGۯr�m�F�����,	�bw��p��˧O{l�5KE��m�wNS:�{N�P�O�f7t%P�9g�ӫ�$�OIL�a lv�	i�vI���2p�K��~�¤#(��[֙��e�4��>~�=��M2o� D���גU�D"_ܹ�h�na;����l��M&����K���P���,Jt�G�jr��綺�;$G X$'tX�L�U-��1��r)�Kĩ��]@f���s}�p@�Gw*�钣 =��X��BI���/�'9�kN��e|Ϩ����Yq�ˊb�Af�32Nu�Ǫ�*�H�eIL��)���f(b���,��r�~㚭�	e����9Bÿ��1�%�}�Rd��6a�hݶ\�>��G��l]{?Ϻ{$V[&��oXOV��v,�o檈(���4㔵T���l܍
:�0�?�[�^E���"j����4B���;j�kO?ܗ~�
�<8(��8]��Fϩ�yJaJ�q^	p���Q����Ɏư
@��j@�S�e��K��hSO2{=�))�tA(݅&<x�7Po���٭�A`R�@���X��VÅՒ����e�{	�۽��ߊQ
��r�� �?^�HFz �Mp�z�����, �3p*��Ax��U06�tpG>�p�եhv��O���ٮ 2p�
�׎j��_�0՝�"}��h�xU���v�z^�K�Vu@w9�ޱ^�U��Ҙ�E�7�$_�._���Ҭ!/����-����#� ��������X�\X쯽C��쾅��2�˸��jEm�'��⊬����y���OP2O	���Xʉ�����|�fC
��i��ǌ_LfW���Y�u�dt�b����)��C���0P���(��F�H����u���
ӵ��Y7�\��JK:$�w�^����,�n��G�ao�&�
��dT�E��p����$�(Ο$�<Q1����g!��ŧ@���#�sw�~�ʗ�%� �7D�f��A-�k���`�@����F�ZhKs�v͏"z`p���fq��-*'�an{�*g�R��WÒsذ� ��&�Gz��G-!��$���ʣ�
�ڪ�&���<G�CK�P7ж�@��b]6���&)S&G��t�=�Ƽ�mZ^Cb����~�V3���KWn�cI���[jBgT=ާ���_eQ��9�oQ��Xߛ�C�΁�q3��T�v�#�1�,%�ݚg~��+I�?�ǐPqigm���lf�6�ӦN�#KL��:�70�ֹ���U���҉󾷰��)�z�HQlv5΄<qN�-yjWCr	��܀��jgų�l�\���')��Tp�h���zT��� �t��/1���&a�3�4mK��uQ�,���艙ܟ�Qf�i�W�C_�%n�id.����Ak V�}�
����و�)$������	�^�~�B70��>OX�F*&�Y�r�s��4LU`��z�n��F��	��V�*~C�$��C��l���HcW-d|���n`xLm�gr �݅�`���+��:�gE�H(�M�v$���� u�\P�%�q~^�&$�T�X!	:���� ��݀�������(����(>�,�'��ĲD���/'���l�H���ǅ37�~d}���38䴸��E����;��n���K'�\G��w�:��mm̪�l�Ӗa-'Z5p��~LOI#���1��\ D��"�L(����m��k��Q���8J{��i�\P�&zA�L�q&��؛����8�љ-�mE6�!泵Ϳ���3�C<Šf�nq��f$+18;�E�ȡoq̣ˑP�����G_^�5¢��u5Bx�W\G7c��34�BZ��H
)(��P-z����,�"�!��
�K`�O	�\.�UHԓ���t���uM��1˚����(�ӄ+����ىw�1�~fE�??�43T�z��u���O��G�n��}�e}4x+��������|����ւ�c�z��H��s���A��h}������Y�m7��n��  F��8{�kFP�8$Ŵ�1�� ����z��g�}h�*��j��NVP��~����z2?[�C�AiO�����J��z7QÅ�KB	��z���:�Zo5mm^x�X�xڋ%�� X{�����
34R�� j
����}]i'綰��*��xF�A}��2�N'Q
Y�(��[Jp8U���uOo�{!�������1�A�gA?�s�3D���}� <��e�ef�/��Ґu7�c�+E|�q����z����I|ϫ�T�:c�(�);SC��-����U�m�y�	S��A�@[���$k�M�3DAVY��ɶ��L�]�v�1�	�� ��3W�o�=�^zjo�K������$��ֹ*(g�E�*���* ʸ89@�Z�z*�/�'�Q�:Ѫ#��vW�����0Ѡ��Y�2�>�K}�z�6����#Wk�o[�U��w�P���	R�g��o"�3��[��E�fy{�5�[z����4�Ȃz��e�yiB��@	�bCg�Ko��<=�q����NQ�0� _i��>Y�Hଡ଼fg�PҘ�t�M��V�E���� �_�r�l���͵�9��I�}���������Y=3��q"ס�k�^�f���֍��җ��/��yi=`����L5�+e6��R�IJ����5h�߬�T��Sql�t����c�k��#*�V�p��JE갪vU4�8I꾂kw��BL%s�&@�y�d�Z͎ ��>�F�g��n&���8�>�����Wmʺ�Yf;S\��1�*�*G7�5�Y��O��w9Ñ�Z�u�A ��c��&I˱b�hOΎ����e������XA���I��3'+�QI̵z�FoT�s�V������|�]{�� ���~H��u���ϊ���02a�K���,q[aIX�ԯ)���W���$h��q�}�d��r�b�L��Vq��G�%IN&���n�t��/U�o26��$��{���m��0��4ys�坾�-G��$����B?n�'m�^`곯��݌�+�N��x�J�"u�"X�j_�fqt�+]Qc��YɊ�[Z�_��s�)P�R>�MMMx�"�2��s`Pn��j����"J�TaQ������c\�h�͇�}a.�iO��{[��IrQ�p�hbIk��ٴ斗��ѵ`�4��G���[.��n��������U��J��'T8��� �����Z��	����H���A>GQ8nZ+'�����:J�nXג8JMZfTl�_eVO93w�K[�8/aÙ&ߖ��f����D�Y}�	���WL�yM�p����� �C���?�������W��r�����g>�-�4�㖩*��t��7�|��kH�=�_��p��WX�zn�@i"/�|�U~��@�����M�2ǆ^�\���V��ݟ�ң�
��D-!�I"T0W��CWw�D�!(��>4��an�q�Ƥ g� �a��Nն��x��{Lbd����^��ui�q��%�ѝ�&HDhD��~b!6ʥO�Y�0鋢s��Xa���&>iL�B3DZn6�����)`�$?Zx�v@���l�ے'��,��;��SW���:}���,w ���4ؼl��;�9[��0~j��9:g���l@0	3f��1�����u��}�wW���{`�U?��qo@����ɉ�"����NSm�u_9p˼����q����D��E�ҚB��ڌ��oJS��[,��
��{����t�r��s���}��}N���y�������"q$��B���	���-	{�.�{���ʧjr��)ޓ�:T»p�5�-�F�w��=���ʉÎ���5�ϧ�2��B_��D������5>��Hl�]e�Z�ʫ��O�-uo�6�ZP%�Ë�0B�7�Kԑ䆀��0�}|������{A �ejR�=o��6�7�Fڢ�R|��_tmW�j��DP�e��F���r�3
X���z>�48���������`�����{G��z�<���^��p��Z� ��=Dóq��մ!/}��T��%Ͱl��~�0σ@���3��s;u��Ѱ5=X�:���A~)��-S\�sKM�z=�,�=+� f�y�.2�{�	���t�:����;�$,��uU�1�x�:vM��nt��+^��8>ˎz���yc��<�۽�]�q�
?z�������>j��i��-�����u�����8ܑ�}��q�e���/�	���S����^鋰3�U��y�d�0v;t6.50?Tɸ_��U�W� �Q>�I�!!w����)
�?[Z-���:���0
�F)(�L/��hpTYPv���c̾�=�]��r���K�%�04|�$���!1b3���,���Q+�H���:dR�I�َl8�$�s��N^z��9��M�+]�\���w���p�MPB.�`��uoa�!@��Y�0�R ��!Z��)Y7�t%Y�?M��a�ً6��&_xS�2��kn����l�GF����BR��M,�J?�-�D�E��[Ǧb���|�������A����l��d��m�{f��ͭE�fH��%�ټ����)vJ��2���˅wR��_���*=��/�xJ&��UO;.��a8wp9cj�Hܭn�>I���uFJ6m�f��s�	:���p�����#_�4�����`S��T���x`9�����#����z�#���=�ߘ��������1��Q�O�h?�|jr����4�~(n��G�Kq�$ǃ������
�j��h��WzB�iG�?��Ăte�3މ���|�Q�X�1\��~U�/�PD���+9��Ů�Ie
<�Eeo7vڞ�@O��G/U}G�d���F�C2��I���x�C�%�����&�IIJ����m �	���������]������o�ڼ�X�yI֕�ǜQ�Er��������esܼ�ɧĠ)���
]}�Na�I����+ug0h��D�R��fӌ~]m^�^l�'߻8ͺCD�>]��ahP����ϊ����Vl�7�������hFq״����n��"�K����kc�F��z(� �r��t;�9�I�$�;[>��4Z]6g��+��A�������=K]�}����&0/^ZZcQ I'/�ٙ����o�CU�C��w]n䏙��Z@\bї�����>!q����ؐ$������I`.�b�d�X'A�����d�;#��Kax�bg�(e`,�x��s*5(���}V{۝ԙZ �A"q��>��j����:v�d�$�kLU��н����ˤh��!� O|P��#�� ��o��Z�I���2�	ըc�b.ND�)5�a��Dꟸ/}����������W�lvaZr�M�fӝ�[ik�_���"2D��!�Y�{�W���6�&o,0�ׄ���1:r�<����.��ni�ӻ3$~ ��r���D[+8� ��jU���廿�+7R����s-5��ܫ��gF��3Q:�
3��
i<�%O�Ģ��wwOa�}��v����g�a���<�Ŵ>���8�O�{�t^T�G�(	�;�m�1��0P�9::��=�k���.�?,w?W��a�n��Շ�RH�S�9Z���6z���5�[747��t�Pvvǉ���CF� J)Ѓ�Z�Њ@8FA�e��4�z$�&���_��F�H�h��#5s�#�ؼ���@�WYw�&�դ_T 2�5?ԍΗ:S�;}�y�5-��+l*73�e�e�b���������i>)_�",�|��ua��L4n���FU4��&x;�Qt`T�^3�k�|��6:�qE���D���W�Z2�b���d��]B�H8��?�+`�9�_y}R�?	fNΩ�0U����ÿ� �V��Z�	�ٛ{�A1'�8N�&�����7��NH�)��o��ǁh�_�?����-�O�C��d	������&�Y����I�#��h� ���̩'��h(�.�MR����WQ�t�/��M|J�/��~-%�K�b$	ԯ!��'}Y
`�~��m(���-[�H�a�
�"�x�<�& $�\Q���DD�S�*zn��Wܭ�`|�橦*ȲB�C��O������~/۶ՙ���d�Ó�q�P!��Vg1*�����t	 �L^���=��Z��<9��+}�A/H�.WG�K<[U!����B��iTvۙ�|J6tj�ņ�$ŏĐp��	�b�H�1�T>�q��k�h�����D m'\��v�����G0PC�4f��ڂ�{�n-����?H���)�R+�|�?�GT��u�υ�e`<��sicJ�$b��z��|t$�[���M���i=�\�j\1MM?���OإGױK�w�9�H��j\pÎڪ�Q����؉��]vŉ��mVf���Z���^oq�f���o�:�q���Ee���ʵ� J�f`��l�^�b��T�*!�#��H�=VZ�8�D�.�nu��"_�308�^��"�@���jЎ{�t�H����i�(��H�;�he�W��l	��ɰ�K��R{��d�
Q��X[�Y-2z��z�eӡzt�e�i�.�i�(��$Hctw+!r���Pqz3�`�s'���]��`x��`�6����b��O�y#�;�Xתؗ��%�"�fj��^��t�e���Ҙ�ُV�1K��O�F�^msS��	X��!����K1B� PuS���A���3S���1a��0D!i���v�����F_w���(� ΰK��k2,��� 1� ����=����a(��P���$��~U���9n��I��0�"#��6�Vqdk��|���%���A��(����/���C3|����v�+�e�}�I� ,eɒ�|]=օ��B�� �MO%�R��(8����z��a���[�o�����
�g�54�Xcu�xת� �T�[	<W�<˷��.D���w���R�E�WI�ǂ�n�0�w�����f��������<\�lv�z��E��Y�^��Ĉ�cW/���u��x�r�W��bK�j}� �]��>�6��6~t�ؤT�5�:�~R�!���Μ~m��m->��M�Kh�� �"�ή/!쥶��i�sf>�ϒ��H�k��ע���zI��{�$r�&�L��WE0A,>�U�o���G ��A�����p�^|�ANi��>(�r^�x~�u`��sؾC��nIĀ���P�+�������oJ�.���7כG�f��@Z��T��o�/c�E��D� �I�D�4Pr|u�(*M���*��c+~.�A��u�ݎ���b�'��_%�Ľ���qWE�ԩjjhN6��,��!u#�Fz����0M�Cg��\�ԽH8���}u�tt˷A!x��-7	Ђ�S&G�L:�����{P@<m����qg=3�e�]��Ϋ��=Pkㄇz�<F�O$ q瓨zFBr�������K
Hށ*h1��vW�MlR�ʓ���_z�p�	57���e�O?96��ԓ�He�R��"�uL1
�m���R�ӑ�\�[��*b�A ��S��7�g�<�_:X���B����-�����-+J}=
5Ԡ4/�~t����LO?W=�Ϧ:��K���*��t�Z�YIsLZ��o�"�� �[�@ح� a:��m�ҿ5Ō�1E�����<�;�L�	X��[�KDR?vwFܹG!
I�p1g��3}���x_y��:�H�T`:�;�4����!��͵F�'�0�'(�"�$�8�DhX~ݻ��Z&ᘲ�9���@W"&�v��p�Wz2{%��
��5�,zsd]+���9�S��.Q/���TxqdE�B.�=��v8�����PI�_5�*m��A�	)�v ;a%���5[.�t�-H%g��Ǜ4"�a��Ao�<�L�>��٤���<�S�����[���я�T�^����u��Q3�� �+�D��f��� S��M,�������ZM�n��F��˗�FcU��N�s�����\����'O���������R:%� �1�Ks����q^�&�3R����c�q(�p � y,(�E֏�QUaE� ��ް-����,�l�,��P$(��Iۏ~}]#7�~��u�RuD��`��u�����PI�w[r4�[%,� hk�a)�J�\��t�o��$]N�zU��2�Ya鄞.3Ut`���1^�l( s��h�s�(Z:���l�x�D_��K�Ƒ`8����+ק[+{A�gd#��-~��`��L	e�q�\d��fP�J~��~�"1tVN����d�[���̋�v�N�9Ϭs�4JC>���1��h��S;�:�'�����l���8����H�_�tf�3o���q6��k,˙~���W�x2S�G�t�va]��~��7�= B~ĜN�udv1��ܮ�n�O��8��	m�	��">����N{�$^|xT ]倎������@�u�FU�~���|�9r���u�d�9� x��V~H��n���%����6���M�1�&J�_�#�S��4�e��;c�5k�,��96��Ғ��a�׽��w�Y
yv�HGK�n}�|�a�/;L�q��?��(<��ً�pq�S���7�lU����W,K�Crq�>��{���#Z��=�
]Ψ�yX�M��D�D\�1�#z��H �&�u���=	��j!ם#���]��%F���sC�(R�(%P?/����ޤk�"]H��s�T���R��ϥ9M[�g�\��u9x�ʄ~??��@�I"��nN��7{d�i��:+ݚa�v6�!Xc߲9���Gj��K��)�#Qx�iL��rk��)�ۊ�)�"/��W��C�eV :B�vD���F�_<���(�Վ�9�+���6��=�F�y���ϋ"/���n@$%y���F�N��1k@~v��u�@F��o���r˖�jt��Ul3�剜��{M�m�w�,�o��[4T��'Y��O��l/��{��Aƛ@����U
��w�RC^�Ĕ��`TǏY���}��5͂�ݨgMH�n$,OE�����f���V��r�G�G&�ɇV�qx]�%��$Y�0?�ԄO�J>q\aӓ�K�-�h��Wz�Zi���rV����g�3�p��l37��^�k_ș��o��>�M�I�m^�K��TfT�����P�E�$�ҵTTr�׍k���ѧ�#l�͡��m�©�9��A�V�kE�����۔���\I�g�FT]�Mq�還t�M��������됎�]�~j�Xt+U�ՠ��a/�&H���ΧV�\@�ȷ�E&UsJ�-g�|��Ey��a��Y�� RbDV�+&���(�����(;P�ڶ"z=M<�?� ��lt^�GW��uJ�k�:<��r��;G0V���d���v�pn�!ǠV�Ƙ�+@��|X�q�VZ����6�����>���^��ה7��@9������1�Uv���یr%{|F~��܂"���1���*Ό䵠�L>�E%;e�}�@)�Wd����Q�!Jkv y� ˼qӽ^i
IC��A�$R?�����J?�af��Js!e�rA�j�����	?v��zz�dS��1�*�m��9�k�j:i�<4��q5G����2�.�0Y�F���x|��N�p�C��n����|��q\J��\m̔��a��@��GD����������N��{�&�:=����6�u����cм��,?B�R���Xy�B���JKŌ-��%̽��j"ʤ���t)��׆���iJ��u09������7�����l��zY�=1Ƣ �3<��=��b�mg���$��K��%y�ʨ�]���*��|�Z���j�u��eoΦ��O��3AE�����8��G�1�:5s���;��@N����I��ӫ;���ь�X�q�+ ���6�5U���T�Z�1�X��Y��Pq#~nsOpۢv�봏h��I�5	L��o6{�k�
4���(� J
�x�؀G����҂r%��p��3n���;���ظh��}�Or�А�D�7�֧�7J�����Ll:Ԟ�dF��"��B�Ʃ�����(8C�W\c�6��ꭴ�K�v��U1����8�樨m��I������β\���6'���&�+�/�2a�z�㉿��rdm�
�[W��HP���@w��o����&��5^p�R a�7jF��T[kg���3o�"���^o�ѷ��k�/�|�[:+�1�Wc�޼OJ�*�ՔH�(�2�gu�g�UP0q87���Fd����
�X{���+���So�	�8\��.�_���Y�ҦX���]B�ntQ�jd���h��ۀGɋ+�<2�Ox�,==V��f?�x��
D�c|���(��w-���UKL��^_2;':q�d/q�BΊD�j�
��8s1���67���_�D����|H�6�
�	��zP���g��y=���4���)��_^C��|��w��g��Edܴ�L��E���_�}n���%��N�/S�����71�N}�O����!3�KP�fr%$�%zi�s����\�┬�J$T$��'�"�?�{O�!J��h�.T���	jc�}�}�O�L[�,�~�A�����j�M��(G,vxfU�����`��\f�yC$*Ra�K�Y�]��h7�v��~�;w��\�t2k�z�X�-����=��e�Y����0�k������|i]�B"��J����]B1�	���Z�D��VSc+�{fC�]E�C=c;G-�_�b�:�dD��I��W���,:_X?R�ZN��2ʐ�./z�P�,zc���T-���1��k�f�Y9#��G�(��롉�±SԶ#oB<�Gr�qxi��JI���Y���U��:q���>�5#7�b$�\1�VyBu�K��ڜ��R��`u< �z�*\D', ��3��k>	���Ӥ��
)��2�1��Ͱ���7&Q�H��9�B_`�Hm�ފ��A��*$��Z�b�2��ȓ���
�(����8�a@�8ZK^�8�����큎�*ﻡ�C��(ݯó��]�Y��"`���4�p��J;X 6�����=
���M��9�d��o'm	!	�(h ����֔
��?A��џ��E���S�h[x�:�M��9� =��t���n�G�O.IS&��^��U�i�[)��]�c̞���S�z���N$��Ō�+LU��\�]Ò���DP�gH-=&p�!�	�B���x��@���������AI�0���mo����2�bְ��m����a6��s�u�� �Z��X�)b�>�@�p��Y̳d������c�M�T�(�jo%0���i:
�0��p{.o;nd4�����Ɣ(LP�E;�ߏ���Q�����pfG��S�,�h��V�!�gsG9�
�E�*��2
W�����C�������)����f��~3f�8��/��-S��،c�U�IEe�q�<�Kvh��N>Qx���.i�a����2
�!n���^=����!��#�,
0��>� �����5��t~����~�ӷL�f@����+��6��.ӵ�������{������׼�l�s7B�'aM�5�%K��I%�}�����K��O93�>q����آ��`ϯP�l�,�16a���t�hU���6_��!�:{�gX��G�"���<���u�Ku1��y\�	l�� ԑS��f����"�8!�O�iZ)0�;o��侻�O�Lsl��M��J6�xS/LX8^1�d�w�U���D,��+�d}�c1Z����+r���pg��B*��$>Z�q��ON�m}��x���4�{�_�]�&�frgM������3��7O���x��TCx���$�X�P��^/��nD+��"�el�*R�؝#�����r0��Hd��c������8,(ɇ�������R�����>r��8�\�}Ҟ�y�1H�"�yn3_!7�-��\����jM���|�H�,��c.�)kSK:���(%e*��`w9�7�3|�w�}������XQ����No4�XpAr�^h�0�N����.F��TO�~߯~���y���֖�:�k �q1Z(:vG�b��=��2HC�"�H�������W�dlu�y�Оt�!*�������8t�
�|��v���3�-���i��f�D��Aw�̙��۳|�o��$*�>���E��4ݏ��_
��=�tXrF�A IF	��p(m�/o��_8��RR����Ҕ�-�*��+F_�axHN9{�X?�xf&~�E�	#��J�'U���	޴i����a���u�K��b$'ދ��ȩw��>HQs14K.�I0��{#N��>�ޤ�*��ÖI8!m�������w�#j��QB@!��N.Ө p�_vat�R6���|k��*Ƿ�܀p�����J��u�gi'�$��f����9�Ѕ�#8�����J�����r�)F�v�y��$hڛH��"�X뢎�5\SY4	X�����&���?ݞ{�p}�<qM*��A(��4�	�x!�����0���PӉ��Zb��]K��a$������jHuk��1���N>2k`��~Vԗ�� �]���8*��mu#{2S�h^g�/���� �ǡ)�L��2������w���W��ɉ^�O���L|å�gz��gںژ�h������)���%��C��A�~��$K�U���`�>������_�H�8ƍ�{p�5� �)�M)i�
��Q}�����\R]?�g�%q>oWm�Q��6���L<ۗ���yI�C�$G8jiY�O���l�W�3H>�|��g��W�oC�B1I��%C"hOy�����~m׾��iyD�X���:+�}9ѧ�������I��x<�
/x-�R��$;	W����
�?[���5�:����jO��g)��R.����R�����.�,]%
�1�>��/���{�.���F����v�o��N�|4M�	����:���?S�_�Pw�B��S�e�&�����6Ńɦ��6�m?��o�\�����E���r�dx=J��`T(>���i��ֆ�\q)ӿxp���b�T�I�ez���h름���D�1��H`�����:v�,ڼAh\Ō��F��\
Ww3~�i^�o�v��ٯ_�a�iU��������*�n�B��f��ڽ&#�H�T�����G$)?z�`2ċ�[X?]Wj��g7��/��7)x��G��
������T��&g��ga�����ﭭ��	g��?�+�<�f��r+C� �����[���ȫ` gdݍ�]&�+ᝰ��D����A��1��=l��m��%�L��[zv��dJ�C��9�)���H�\{��ۼ|�.a��t)�Jض ę|�|�9���6�ɣ+ᥜ�5���ס�7�1���]��w*&Z��3�3;}��1G��8��o��ʾ+��S�?K����1��iKbaʕW�R G��m#����2����A�;�Dr{� Ƀ�l[�9�Pp����mx����]X_(<�y� ��%�ӄ�C[k��z�R����C�ހ�p	�1kVp�k������ʔv��ED�~���Q�J,�M;�Cz[�ֹ
fh�&���#��I? �c����ݵ¹��R�4�Q?St{~ج�Krh�3KRF�� YH��	i;�.�pеM+x'��z�N� ����δ�٨F��d���d�ZI�=�e���oq׍Z�E��s/�6Ĥ5:Mk�&-R1� y ޿^g��BJf�Q���5�r溸	��Ag)T$�;��Yt<���4�"Ēx�i������I���H�j��Y�:D�Kv���u����;tT>��c����+َ���)���vn7�Ʊ�6%�����{v��DU�$�/j
�w�Gq���+�|��6��'b�o52�ǹcg���u@Qy�)t�!v3��uKL2� ��?v%�	�Nō:�Hg�ؐ��i���j]1��t*;)��LK4z�\�؋v��A>�P�)�q��J]B�P��w�4� Z8Q�rZiD������� ��P�Z���LXV��ZEeL��n�p���$sW=�dXb�:�-
"~��Ga��f$���c5�K},��#�-:���nt�S���r���~!���k��Jo��uI4���?O�����z|1��<WQ�f�o�ҁ7�Q�ۦq�
�,������]�66&A��<'/��`�a���C8>f�4[	�`�41�xԃ)3��4Ş:�;$��b7�˻��:��bh���]*&]��m���ު
$�-��<��l<>�b�V���p���J �w6'�؄�ߐ��r��]Qƅ�s�yM����\��j��J������"iV�G��5x:����=����Yz����"1�)�t��pr��e��E�UL�[J�`	t������ڵw`3�"�*�x^�G]\�r!�2z}�C�y��k3��[E���XlifǓP�	#9@�^�+
:���Q~D�c;�;m֘���X�ȸ��*�������~���6��������p[�8k��X��{B�H��ԃ���$냞k�e��x�W��$���y��<~J�Ct�H&������_�*���N9(YB������X�:�a).9�!?ExJ�,�dj����h������O�(�Ìw	���t)tg�Ż�C憭�s�U���tX����,c�Ƣq�2<���g�n�i�6m�"2���!`y�#ЀtT#+�T�zk�z����tH��Tɦ��[��k�^G�@��bD��P\FFN���|!<�z��������Mc�|D���9<x�
��+7��7���Uc�z(�H��6�I,�Hf�)�5��M����nk�4����s�s�i_ewm/r�C��*#�!�0z�năڒ�`|A8.���~���*[>�d�kiW�_ȶ��AK{�iѠ�<)�>�{���BF�1��I��6��~�0@��9����w�ˏ�$=�*
\yh���l0�V�	If���0W��]���ӳR�����±�Z
��� ��ؗ��p��]�=����O)?���+�%4TZJ����$�#!��{�`���g���0�}ɩ�z'H�`����E�[/�o��C�s1�R|���t�+��iBr妊�*ն�����sG<ڎ
}���ml���2���D����﹐�AŅ4
�iX��^ȐY�a6�����}?�ko�M�� �Z��㏩S�x2Rԋ�l2�����d�Ӣՠ���z�Қ�����Q?����>S�\fY��+:^M0���$�þ�}��[so��[��3�~~�t���\S��j��h7��\����Tc�� `�Z��5Gƻ�j1���^~E��{��к�$q����[�X4h�-�P~��	;�^��]jfl��C�/5�n�tA>�e7��X��U
�+��#��u��Xѓי����L��?�X�/��NH�[9�CK�ВZ�a��a��!�kYJ-+y��rg�06��2���7.�IWd�x�&:�f粰�N�VF8�FM�	w��W���p*�Z��&ӕr�U�L6��am��8�,���W��L%D��g�ӹ�w�����Y�9�z�X>pCX�j����{��>g�]���ӗ[	�@�����kϬI�S��=��l�[����[�G����'Ԭ���#���
_n����I���A�F����oZvu����q��:�,���ξ�dB�%�H��1�FC����[��r�?3$��[���?����c��(��q�<����Z�����N��F�>ƪ�Z@�p��)d��q�"q;j �s!-n}AƢt��^��`�u��®k��m�����p���H����,����;K��E�~w��K���|�����:���[�����b���s����H熏-T`w[�_t�:B%�ł�s/��-�M�����W&��3#3�˩ohWp׀U��d��Mx��m^������`^_��G$�{٪�����4���4/����|���lN�U6�9~K�މ�q�>�x��3��@���$�&���/��7�'�0�P�xˎcfI�ʾ��g�_��#�0)Q�4C,[3�uδ��;"0�L$C��U�Ҫ�>E��mh��_�!�ʹ\t\In�t:�?����s�;�e2]�=y���$݉��7R��G�{���8"�}����_��2�0�g`�0X��v��󘱲�?\�8=������w�ț��a�ܤi&[���G�Cx�T넎c��̵P=���Z�b�-�S��5�lI����r ����x0r��a��O����P�?�����5�u��ʹ�Z26�ڧ����nF��%����g?L������Љ�`!��]m�@����iS�~����<�� �����u mLЦ�!�����f����e[�Z��R�=tGo����gY��H��iC���'n��֖�o[�7��ü�,F����=�Ճw����|�ٱ�N?�Js�.r��9	��_V�(�*��&���"��)/k�����p���aƧ'l3�n3j�x�]c`'�?:A^]���At�2E�E�K�T|�a�?����!ݑZkpYEQ�������>p���[��_�.st�L��4?fY�����ݺ�fS������b��.�)�X"�<�|����C�֍��A<s��Tr,��H9&?^�y�Jz��$�	���X��Xm�n%ǈ��V%�Y�^�'[C(�g��6����ǐڅ	 ��1�������;q�2�Њu�6�B��쬰 B˂�(�7�t�f,����'Vm�0��tG8���k[�1��БԨ5}�����T{�()�W���1�X��G����o�ZLvh��$�%ߢ�.�a+H ���½c��m٠wZY�3!1�@��M�R��(0g*Pz7��(�Z�.�����뭗�rU/����)�ī�0�C��^D����b��P���`B�I�������f2������I���@{�tNe����z�i�������ۙ������U�3��rj�ɥ��e���׌DZ����Sf��n**��BN����SV`>���_c/���7N���Ɨ�+Ӥ�0� ���N8����0DT��.�����.$�zl��]�O�`Uwr(1{2O͚̺
7 =��h�ۧS�?:(7��	�l�XE�s�ʜ��狠
���б�Z_���Xn��n��nM�x
;W�V����"��+M�Z�J�/M�ӹ3��>
��u�`�p�,;P�\�k8��g���&�ԠI��No�&d|�$F �yk?x���fɌ̅ΩQ�Ʀb �``2��Dss�!��3&��$�P�c	nJ4:(^gܴd�,]f�	�%oJ�e?��[w 47M|����D@�)��C
Ց{m�!\����m���sNQ�L�S����j�rW҅.	(&i�2{#v1uh2���.䷰�gXa3=���r��K�]Ga��V�ݷ|̧
��r)]�E2��O峐��d
��M6�����ߋ�o6ƅ*��v�}K���-��eR-[������8��[�R8�"H�g�c�I�,�H����P�S��~�E~���H��&����@xs�ө��w�В+A��C�tc��]`t��������`b��	�R��d���!� ��P��M�����xQ>�=U���Uo�S5;>]��BD䅛�k`n�N֪�)//�<�����+w��r������|���rR�G�=��v���4(.z,����蕵�	��:��T�Uxi����T��-.� ���ȃ�aV�p:<w}�"4�|Xl��\/�g$�j���l���3��+�8�|�{���J�{ 8�!��}��s��yq������g^iɽ�~�c��XX���k���(MN�=��,/��)���ύ���L�;��q1 I����[[�i"�<�܁Kq��c�`�^�;4 F����Ճe��Jkur`坆�RvWP���
8�Gp?'�N�X���@����:����I�$Y1�D�^+
Ø[�T�I��}K�|��-P����:�
�ʏ97��N���8���V��
`���~L6�l��W��r��!�0.��88Bi���:Ԉ�)�
��b��˙Q��.�Db��r	hh��ak�ZՍ7W�n��ѝ�/��/�����f��s�݃*ùZ�񁓸L�RrHj�]ߝY�"����Jji���j=�U.�yjK?<�h6�z��A��y���3j
t=]#ԡ��>��-�:�AJ�v��%hcך 4 '��ZX�y��T���ݍR��Q�Y�S�,=����yP`�z:C��3�x�������ן�����~x�6@^�j�C3-��R��ֺ����ߌ"K��ͦ�S���}�F����2_�=p��y�}a��a�w� 7�8�q�W��Ң��1��c�X�_�0�j�����A̔��e�­ŤQ�ͩ��To����6��sP����v�xL�wړ����"Jf�:P��L�?��A�3W#쒌Q����*	V�U��~����[����xiQ.>Q��@�� YH���U�]��5����g������v i�y�EiR�C�m2��vp]��~���HE�a���d�x��`�|
�,B`6e���2�/?S���=Tk0�,Aw�ݟiD�}
�l�m�3ND	F�x2�n|?fj�e����t�'r�֎�V�B�6�D|�8��"ޥ�t�+;1O���9t�yD�#��1�98�1�KVn�`��.&��n��� A�h؈㘘���]_֓Y����s�n��in@���Z�Gd���T���w �����L]i!�v�#;K�tmn��dG����F�Hp=2$���!�Q�^p�����Y�$钍)l�}o��k��Z���C~��`� �Nӧ5��m�_W��O1���7�*ǆ�K6y ���9���.�����@X�Ls��Kv"�7�rvD�!p�LԨ�����ό1�V��F�a�u���c���M±�4 c�]�
k��-{n>�+Ogk2�跊M���#Q��t0�G���@��{T�lU;Ƃ	ii��Y���*;������Sq]�f2����S���Q�b}1%��D�A�yH@�齨�Xٙy����nSn�U���^F�+�����F*���&ɜ�	[4ܖ�=j���k�ݷ) K>�ȗK?�z-!C_U�H,L�u���q�Ms�HZ��9�6X�4H�2O��"&?)9��o�-��ѻ���ޖv���ƅ�nqMq_�+1eY�WY?�
68o�D���,o�m������KP��"L�9(�%��eT�s���BSn�$�I�G��֩S�˄�1v^���uN���)F�{G\��D�Y^T�K1���gQے���[?���t�P�=�{�jm,����ʊ�5R&`��K�l'��j=[��ݯA&0��(�QK;�j):&������pY�0[&��99��"۞#���u�bt{���@o��t�p�)+z�˓�P��¼�>����A'!/8�~�D�,�ܟ�	[>p��.B��x�w�v����Q��P�z����<��hq�껗�3X4��G���؂�� bxy�ԩu�f�n��ak�P�?s���u��]�
p�	dO�C�L�4��C�QOB׵��;��l!�Y�P%熨o��JS%~2ʎ�:B�O1�z��^��s �*���knS�+�/�^Xy�h����Upʘ���)��*|���Fעϯu�]����j/�/�5w������1݆�H�oE�L$ە>���6��t�FZ�>�`&�\�G@v��5�n�"��QMy;��
t������&�M�����l��{ǫim�����%_���E�ƣ�3�1P���d@�2��$Q�1"sGibwv���V.�@���K��1�*Xb���! -�5�U���ϫ���V��n��;�P�uk�П�]U��/����p,H[߳�}�c}Hȍ�3�����U0�Q.4y��t������KU���Q�zBa���X-hPY I�N�U만t~�@Ȉ�����QHe���(5�{--�DO��M͏w9]Y5͠��0<�Vhy���j�/­���P��&�F�2_�Izr�V�q�~N�F5'���.ڐ���_]�����n�pM�6�~�G��
�9~�)XK����}, �N`6IC��&#�r��[:��G�#�*��&h�w�j�ʭ�ez6���9�;Z�ݏ����2����"���(t���C��)��D/�-f��9�R�
`���b�x�>x+��*��$pϧc��<@����2�4��(Ϻǔ�pE�%�Pؘ#��>�$>h�@��ej݈����t��7s�ot��*͘���m�R�P��Jԑ�T˯�����UC��w�"�P�n�b�n�E�W����3@��p���錨�(g�ۗYi�a-H	�wO�P[g�R������.�b5����҃����@p��"ڗ+��yPT���������?!��6w�.���@X��^Ӣ����{��ǙA�A��m)Q��t���Hf�V�[�S�I8�7g1�g�O���}O5����bE1��P�.���!2g֯T��d1zx�<��;�P�Jf���d�T�[y1�¾��N�=;�Z2yk���Ւ��sJc@v!�F�)_-๡��NN�W9����$j�����,���b$i�&��@� ��{	��O�ܔ���,���{�ZJ�F�sb!�bHv1�
�����UONtf=a=I�3�z􄁿K�i}��FlH�W �u߹��u�
UΚ78��C��f�Ӕ��.2�+��U��	� i�A+�JiC�9C}��:���!�I@	h� �cg�uC�;�bstd�z;���R�p������Q[d��1ze@S�6g��ة�ZN=g�NT�%������CN��È�S.���g�����»Z�1�3����UD	�7^�֕*s�{��  �Ձ#�����K�	k�U.g�:̍�=�
�X0����:�I>��w��, ����G�:f:I����[r ��ǵ�u�z�T*�J�װU���Y��Vo'�k<�=��˲JJ�Y�Jj��c�8h犚<�r�/��
��LXU^�,����_{ư%߂�#\!�LG�ld��eB��+,�S��&V�4�k��;������~�˗�r*��40�f:h��u���T`�Ϸ��]a�+6-��6��%o8Q����-I������p=���]��a� ��\�~�^{�[,Ga��6���1�A(�����@�R���V�!�ܔ���D��E�V��9�n�3=C7-���K2�w_8�ȋ^.b����%g����:�w��m~1j����S0q����Y�^�s��A�{���w�c���-�S#%@	�9n�D�y`,�=�	L+�>��d}�#Lx��u�~3'2MB���EE, �x5c���6D���)8ىh���F_�?�QH�d!ݛ7���K�1�����W�',8� {�Z�I�&R^��n(��˷Iqj�`?�[��SD��1�Y���<x��z�ޅ[���	wv�:���~���㆜�e2k�^�+��Ӽ}r�cD�����[b�D���?���n��?6`O�k;�M¥�,F���7��oUx�O_9'{��݉\�b|͖l��{B��8��I�5)���/]V�^��;�n� t<���XR� 4��J�,zcJt�U��w�n�9@�
eg�qD�NSi�9���bc1x�a�!��?���-��u"aZ���K��Ts�Y���9�����;!�fs�<�I@Ge��۠̋	t8�1�^����(S�DG��w:�N��Go���I��3���!��ĳ��֢��� ��� k�>�-�^��Dc?�L�sj��v-/�y�#����!]_}a}>���D����e�:����o�k�RU��'�oV�����(Y6I��&�Ϻ<�##��8�O7G�R�E�u?��TPl{S,E���F�'� =,�T�&a@ ����,���tmOM�}���4l���q��T���:"�r�V�P���8��x^��ԋQ�#�2�s �y����R�������S�9���ƞ�y`�4�Q����:���:S���VW,j�6B��;�S��>`�f����E�˿�e�#/�0�;���Hw��)1�,�]@6�mq7K�Oag�%�Jטg�[l+�\�[I�.�M���R�U��n8#mM_���iR�%�Ck�!�\�L�a��2��X��$�ehq4	j&�w�i�)��%��^��������}�^Sgˏ/x3�/|��9pm�s�Mp�r��Rܣ\��8r�ϟf<n�*!��K�o�*��B�W����`��4�1>ҫ  ^2V�f�Tks{�l%	R����*�rTGv����	���r�{z����%�ϓ����
!O
�a� ���cu��:��Z��"��_���0iЀ����;JZ�]�	�+M�
;'#�bz�K�N�.W���V��z*�m\�Z����ԟ�^�ZkU� ��f�ѾD�������Ǆ�|S|Ay����CET�o�+��� !�G�u} R�o�h|p�Y]�ӌ�}Ws2������)��?��,4c��sw�����ȍ�_({z��͒���@�Y� $�ak�cn&�zPN.J���E D��-LW��`���淦��l�=��2L'�g	̳����ᔭ.xEՆ
�_�����로Ԕ	~L?�O�'k�H��xn��3�rX�N:�����x���-�I9F����Q���HD��j���K��;����"��2��3�#��g���}�O�"<�x�ӿR饢�>�L�(�4�v���1���f �7l<�>�CsY��a�+�z�����ey��y�o�Ml�&�?Z	P�K�v�dg����J��iؤ.s���5�̴]�+��S�e��f4 �\������׌[��)��fڜ�G23p��
���1��`)���-q���]�ַ*�`tЫ�����b)�06�"T�chm�cr�j�MV(���TJ����}�*Cp���9�JL��>d���Iǝ� �K��9YlIb���W��͎��+G�Cs&��Gn�����M@��j�>f�n{����m�_Q���t�`n��)ao�����NBYt<`I�?k�S��Q��#w�[0i�Ttf/�^�5PPu룖Z�kj�4� PK�1_��K��I����x�a*Li6�ȪZ���J����캜�Q8f[Wbʺ�2�}��).E�o��,�}�����t�R��5�{s��[&db��>.��%$G(s0� 0���&�s��?Fr�@���8�܂<Єd8��W�K(�q��|1��`��g�^]���Rv��!�0x�2dS2���������d�f+�Dǘ�:t_�03n[D	�ϾBv�#;�)\� ��v�����x"�w��謑�i�%� �;�R��m�����)JJ*+�Og{$Tg :�d`.�Z�k�¾ʊ���/?��E��VD7�|��VX�����`Q����Ďk(��+��}�,v/�~���Q���Q��NP4Z��O�) �����z�6bb�(S|q�.�&AA�s}�S���ϩ�En�h*ƧӉe"=8��"��{��7�2{�#��5Q�=��\9�F�^� M�61��`�n�j%wUYS�t�!�I�&�$я�V����a�-/�T���
�[kgf(]�a���k�e���ڀ	�ZΆ�� ��*� fN3�Y�ڋ*���\y�o�+R"O!)�ײg��j�OGc0h=<e��������n�Q����A5��o�f�CF��J��`�n �#��8;>b�b[d�aO��t�EnU��wQ{Ȃ����"$�
��) ~�M(���<���6	�$�Wge�Y͓���al�z8�S�0�҇ً��w�_��+<���T$"j ��!��mwDĮ*81�ɽ$�O�at�r���_6��d@ ����R��h�K����u���U�חO��8������s�#���S�7*8��_�N��&��2��N0��6�_,%��1Pe�ϝr�|��A�w�k"^���AL@c;ưs��Gɓ7A�y�H��l4��O�W&(�5P��ORٹ��ݗ�C��h���Ď�Dkkx{�E��Q�X�R�pVLz=�C]�L���Z.��g�|�u��OYm�y*RZ��jd�Q@��$K�}��0�yl��Z[Y��/PH�������т	�6|�~ο=�U�����{�3���6n�	-�ձ���V�!�,��r�޶Ȁ��y����w��_�
0��
{��9b��h���Tg��f�3U�N������N��}�z�{����,@�=�o��U�p?��N+U^��+cH+�p���Ҙ�b��>C3���m���AQb��b3[������h3X�N��[s,�__�W]ԝ�=
�!�h��̧
��K-x]]Z_+zk�q{{��gD��bQf(���P�8^T�;g�EY����.�U��)��tJ����e��?��P4�������iX��s�v����s��S�8���j�1Ώ���LŰC��3��ѝȒ�� �
It0,��'�E3��Pܙ���5�`mI�ֳd`ܟ�{�(c���)~ؿ�My���j�X�e*i��O��x�,W�b���j��@��t����\_	P��P O��J=�M �����@�Yl�U�C	D+��Mݸ������7�%���O��P���:��%�������{s>�
�㴳�[��۳�P/�.R����̆��ꈉ�r��Լ)��P�p�[|�~OD���;�O��is��l07i��BΞQ�d�x�ᵪ��,Ɠ��!
@����-ܮF�t���i�l������VR����v�א'�2ZxL���;s
|F o���ׯ�}�6ɺ0�=I��w�������K����~��|�.m�l�%�i�L��`�H� }�Ц�`˅��������4�:{#����Ꜹ�5Wb��%�����_�5T�	��`h[�υ|����a�t�71��tS�|j`�G���b��*��FjML��g�?�L��^�%�sS���;1���_y���Ih>��P0z�F�������B�J�_d�V�S�a�G�=��I�nI�-1�ػj_����ak��ڢ������a��ǲ�ϒ�%f��h��fi|�����xG�0���e3���ZS*�9Zh+0��|�+�V���6>X!5\T��M�b���n!el�%=�g�`�-�GZ�i�n{{��bC��C�N��O�y�Q@.{���e�Y���ԘUF�g��b�N7�c��C���'o��-�P6�#׬��[��[*�9*/����6����e�"��=F1�