��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQl�E��*����XR���J̕����u�0�t���P#�_�Va�^��(�u{މ)KY˞�m����a��a~����p�I�l�����q� ����SA���ɒd� ��U=ϝ�g|m��g��ͯ�\E�昢�*�_�5͔J=���R1GΈd\+G��K3�Rnq�?����7b�X-����w5�LPihot�t���<�&�Y�C�O�&�+z��H(��akx�N`�bX���V9Ƴˎ������Ւ�̌�1X�������g�Qm+E3ohЩD�=�?�
�<�&��&����Ґ�Ħ�@9Swm��#�Y�f
���;�L/�Wl�|���
�N&�ץD�upo���s_ɶә��ɫΥ�%��-���K���n�K�J�"��d�h��O���,��վov�Լ�dii��p��)���e͔��u
ؒ�����R�z{�8�U�u]^��L��ɝ��oJ˄c�{�����u��&��2�2�V�/@o�8��N!�ã��/ܡ��;5
�oR���R��P4ep<2���3�u웮��{�eh�<��_��]�����y�4�\�1��{��$Q�ALT{�
eKf�HCM������9A�[�iT���b�7�
[=sS&�R���T���r�H���T@e�wY�L�,����S�!��o�:�s��ւIc�n匱9�i8 x�$:�VF����}V|"���҆<w
l��Q?J�'-u�5m߬j[�=6�h��Bx7��������I�<���l���KT��$<]�^@77��N#Z\p�Xj�S.�չ)2q��xY
�����&b���4"!K���?H,ĥ)�&a��{��*DC0��_�.�`���,d�K5���:��_��?���b���Д�*�f����s���tD}|w���.��#�	Ox��fNw��-M�d�MXM
x�>��s	;�[�T��tI��>����&��*����'�o�b|�X��`�:���Kp4�u�j�����w�"�C ��S" �k�~��l�>��aɏ/����h7�p����`X�|r+t¬�DTk��J�%Nj%dޕ+|�k���@!E�VRʍ�mL�~�������
��ߓoU5�d�i�	NVc����h*q���7�Q|������Iw�M���Y�^��*��B�"�Q~�֚��<�b.�s���v~�@:�ANYgv���H�>U��wj���[S`�Xe�3"���A� T�f$Zܰ\��G���,�z,����V�C�ŝ��̧����Bd�?�p'D�Qt�UF�v�+�c �z�\k���8Y�����d�!���C���.����z����������c�n��ޗ�n�bh�C-�|�V%4���8�@�Q�hF�1��}�1��!}�����,�5͂X�{Ir��h������1����v�R��^#)����ZM�9(���E����������v]��"�9M5�.%��PX�&Mh.D��3��VI]gH���v��V+������GV-��+�]��"�g;y�P���ϖ5��<���-�u>k6���I2�˩$��c�1%Ԏf���}��R�����ч�z�$�[љ���&ʴ�NX�CL�jk�L����m#��2�`W��<*�� �Q�<��B KNC�ع�vU�Y����1�t�~!1T�dmM��A�ġ�^�h7�:[���eD�o%p���he��оj,�>��_Z�N>�̦!vk�	{6J,�uweIm��,��%Fh)k֤�脾WM����	`HH?[����:#Wԛ˚����矟W�XgQۦ��	��̓P���r^T�Ԁ��C���%�(��f��kȕ�	0@��'���3�j�2[� �\�_��pޚ]�kD�R��:܅gS&.�@�t	Ib��Y���O����Y(��n�[\8�9T�K��i���J�4�������C���ɧu�iLE���~r)̈́ϱa^���ʫ.r4�\��n�4��&���A�<-u��J�	l�����PXHj����N�A ]��㯂�L��O�0��C�~���}�9YČ��7������p/q 4�_�K����b?��k���'��5.p%_��S�P ͜��I:���L���G��/q�y({t���#F����,T���@�U�� �ǶOt���>K5Y��N��՛~������� 	#�����ž`��U<���z�-	;�P\@��*E��KI�`�3E��jKa�(�B������t���9׋��-�X|}E(�9��V�������L!�6��f��R���ǟ�Y����OU�Y|]8�5�ZRN����|.BO�c=A2�x#�,�F�kt)j0��0���q��$K��6Li��Y�'��_�'G��T�n�	�/ߧ��'��If����R>Ű���<�*Y֕�1O��J�֕nw�ML>��r�u��B�_�✪���Kxg��.���sy��m.3-6Ȯb��<Xyj��j]��#��?7ܩ�����{����[(I�d�&rD�)�;͓�3�]?g�J��5!���r�A���<Q1�'1�ݣ~F�
ŉ�k9��tc�"���[�̈]��×)]~;M��Θ���1�&��e �[o@�ЭQ""���JEB���@����Wj[�T��4�E�"&��=QYy�m�Pt�a>Aw���ij�1��ozP��j���F��5�+�S�Wb��! A\�S�b(j�����s�����{Z��?��k���^&���)�R8���&���]���`��=*A
�b�t�U��ZV FR�ł�E�:�!U,�H�%�xr�A��T"���|P!v���cN[�r�^���׏s��6������kNusM��E��D�[v�]�K@TU�2�,ʡrI?K�iT�5�ݜMӔ�׳��������Q@	ώ�ɧ���(��X�7�Qt���/��U��z��O"��ď(۶��H�ׁ|�����Nˀ ���6H�<�����#W-Фn�]����&���g�j'��x{��)�ʈ.�����ދ�އ����']�|�3\DNÅT�=f�ז�O�s�!�;d��;�b��2�-��<��ϝK�ɢo���)<b���)��$�u�8�~k��)�a��q��X���?�o<9��įV�A�_���r�?k��,N����.�{.v~�ㄬ�4q?��bø� �	t����u��(M՜���݆�(�]>����\���O������(�GF���x�LW��jpr
�CZC�Fs�����Z����pNλpu�S��=J��%c'��{[�?ELG�Є��/a�~�*w�������{����#���P�;�3T��v�їR�쒠9���?-��4*D;�9W/�񶣿M�� �5��O"%��<�}�-t�*��ZR�.��H���p$��"ݖ�e��Q+��_�^�+L��b�Ll��5���մS�j��t�n���Ɉ��J4-�!����'�h�B���&����4P�6B��+���xih�yu���:�{�>Ѱ��i��0V��D���K90�1�Hh3�?Y%�ۃ?JR80!=�!�t��m-��U~����p�9�!�Q�����S������vH��0�@>�3?Ic�H�D�$�ѢlS�,�DeD���{�#UO�J�1���w(��u �����|Y�"�zw�b��(��mGf�.3��'NڼnfAX���1Wv2���?�a��قWR5/��ыM�2�w��.�]]��Zv�@�cI`��b�z�s�B��A�ʘ���u�Y��yQ�"���5���(i���*T�� ɮ�J�����O�'�+%���4�l|.[o/�˨"/�>��'I�H���Y��.��(� ��CJ(�S�F��S5].�9��2ҬAO�ɛZ"��h{xD�\�v�H:4�ݵf&�U2�PM���I�$�#����O�d�L�@�\jX�`������8����C�� �n�ٹ���`V�6�/�s����X"�����4h�f�
g�Y[�(�co0p5�T�A���(I��{��m�����剼�~�,�-|��?�*�}������c����ǎ��>W�t��?R��M��@*\0Ha�U��˹�6�	���h;BΔ.kZr��$H ���0x�al���C��b�8	�Łf�t��)��~I�"h	����]������)Gb_���e^1+�X3K�j�d��U/.���BNE����fߴ��V��أ�W�nn{R~��j]C�����L����$�E�0K��a[�G�ݧ!���z&�Qɯ�F�kH����B%l�4��׭��\��K��ƬƖ$i�z�y�k���\��k���[;�c�p���~�i���A˙���hJ.�Bz��]������3Ȑϰ��o�����E���ʨPC�6�g��\n`�@l���
k��������e�4��6m�n�uV�V�'�Vϒ�b�~�X:$?_�K<&6:�(yIt3��0p'�F*O��M� ��Qi�5b!	o��X�c �/��Ȝ�5�K"���^@���k��dt�E�o�S��Ǚ�!�Yv�#.4��=���$�ki\H����s��q�I��?��߂$�\�8���L��0>TM�͵�ͱ����ca�p\]���<��8?ؾ��4���_�k����7��`�9�`�vgg����i|9��Q����J̀�e`4Xs!$�H�b}�ƥkw�m?"F�o���E+��K��Xg	Q ����y�b�omC�W9����t�.�{&Zb���TJ�s�3m�b�M���� Z�NHm�o�Q����W�[O�2��=%`�u�_��L�Tpݺ=�l��� H\� ���㸺�![*�~�'�J�{���GN��#�E�'c��o�6���i�2��'y�|�UN���Ӥ&k���a+e�M���I�ʈ�`3І�7PBHy��*6f]��-|&��l)BJKN��a�\�$EC���~��.|�.�&����KgVx��xEd�߉7F�<C�4��xmr��*'A{�1�1��XU�k&�'��ReX�Ih��c�^ġ�S�Yʤ
)}��o9*��-j�