��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0�����
����'a���en�,�=y��~{��i�#�sS�Z�àx�WW�Bg������𓇴r�b�ex�Wv�c���V[�4+9o]��\�S�������_���]U��J��]2c���L��<e�@�&���jX�3r|~�SrOa�{NR^����y�R�ΏD�|����m�'�m@�q��S��Ƣ,(�jݎ�4��>X���w�j2�)M��&�wU�=�a�;�k����K���b���ʎ�\������E�\��,D�`�������A\]��J�o�A�����^�.�c�mC5�h�9����N�
�.�C�!�V ˘�٬.#�]�	ޔ.�⏩� j4pTMt��U�uW#�����3��ɐAw����/5���C�اDt�����e���#�h�e�W��QyG	��,ct��{6k-���w�Y&=pK]kS�g7�̝WJ� �
�Y�X�K���L �n��ӡoQU�Iy���r���o2k�aYDx���v~WX������+��xe|F\u�R��0?ked�1G���U��'i��Q8{���=X��c�H����Մ�t>�
ޑ����肤%�n�ˎ�;��|�бb3@�yh��CD͢`�Pj|8�&�lD��Bd�Gv�\����J���S(�J�{ɺX�n��S=��/XE�|��ڊ�]4D�P�����m�D=1�	I� B���~p� +���j�-��2��X��o���Y��z�ʀ�	������>��@⡢ęKM1�:u�X��b���xl�ܖ�2�J;�x��M���� j���i�u+jnH+n�[Y3����y�~�{�6nk�ʔ�$O��7�vڧ��������c��43�V!��B�ܝF+���� �_fZ���z�n�5&���� ?ڧ{�:��k&bv0ݘ\�4��s���e\R�ł�Q�yN����/��]-�ѡV�^/��bJA$]3'UW��v������Ft���>d�X�aPp�jj�^w�ih��PӴ�ɵ��zr�!@���F�ڭ�D,���:r5���}�K	�޶�ΰ���֌˥�p�[~
�j�i��_m�Z7Ø�n���.YT*&,�8�� E�m�N-���h���{z�T�:Or�^�3��*ј�Ǎ+��l1L%���ɼ�q`*���ҋ==������%cZB����j�0׹�R�ZPIg#�-�����*o+�ꝢlV�t^r*R%�d��߯>���H��Q��9�Tl�,�����F���B�Ty��Ou�h~�F��J?��m��)�wEsu$bRF�9���s��ơ�C#择l3�^��f��]�	|ߵ����H�ШH@
qU��\"K��=*
��A��9�f�8"���쭫@0������B^��f*���)Œ�>X{�=��]�wh1�j	b�Ig[so6.�ip+D�d'��c��,`{�ir��
˭i���͇����cm=\E������
����Hس{r�呵��滜�M��b�j���nE��2k֡���^� ��$���U@pqb��M%���/��e�pQ���F�Z��]��~��.����72��!�fT�nS�P2�D�z�eТR�5	pn�҈H���M�5���e�D�$�i@�[�w�K�#-ɻ��������� Ej^��!�(ˬI�c���}���y�,����m	1�Q��mU�Þ�`,� �T�8����Z�gߐ���G����dQ�(ޙ+���!��m Hh$
_���=�d��kݐ&��Ų���Ý;%���	��Y����,�+ҡE'k���Z\�}�%|�k� PYp_pۑ	�#`F�� ,�tr�Gśx�����z�K�e��uQM�j�Z�Р4��U0��<I�>|��s�#�W��?Q��!��;�͛w�|wC�p���������6i��,��Q�w��7瑼vW�c�6�_)w=)���G��"l��F|"�"W�zͭ0O�M�DB!0��Q�-䫤%����������P2��(3���#���R���!�"A̽�!>�#[8a~2O�c�pD~��Cp,/�C&�[n��bj��*O� G,·�ԁ~>���!L:?��:�Y�+5�6i�,@p�(?x���@���c&j����g��$�̈́.=T����M�/öY���B�<�!J�4���7?�\�Zfj"�T	*jnW��Q�qƍ���"t7s��������
�t�c�:�u��{����?��T>���Jz@�M����@��0_SD<�U��!�k�7����-j"~>u�7~_	�n]k�.����i	󼦥�0Iб_���d��4h��uT�J�,�B��M2iM�%{{�6^�2�@3y�S `�5�G}Y �:@���2��w�ߤ�O�'���� ��X���D螉�-�&�s��Ӈ��1�֙���˶tv0�v�t�j��r���ҭ�����\�?���R�4{�:>���i���ԛ��j�T1}���q����=�H;��1]2��I��R������C��a� q	�T��t��!����Z٩���I��Y���=n��'��4p�hYi�	9q�g���~U:����t��,o��Ĩ��_uJƻìޙ%��P2eo��d=���B����cW�����4 �
��g���c'�g��!7� ͞i=3G��G2�4	l��.꟨��}�~���qm�κ�I�\; \ ��6��å�5p��o��q��ii�W��D�)T�����b
���¼�w@���y��8el�kA2mt�]�����~H�<�ݭ\(���aw�F�3nDc�]�i�Ү����^��w�Vzl��u�_|~�H�f�J�ȚF9tu�o�=o�)r�oڶC�5tH<��7i�Y\:)�\aU�A����2�۠�f�MI:b����a���Z�R�j�芨�fӄ�.T`���B�G�(�K��R��m!�ie냒8ۤ��� \�=���0v�-0��YC)[P�~�:[��y�3�;�7�i�4�&���1�/��qfe*�qp���F �y^�z��|�`��ľ��)����?��sn�h�BV�F$��6����)͹�j��F/�?�f�$�t�T�o~j�C�\��������J��P��\��8�5��DuYo�g>��u�%�$hGX>�*%���P%�`~Ѹ�eVM(_3~�8Q�9#k��H���!��wr2I�Fl/�ppzI��q
���[�2@֠�i
�u����UE6�W-g9#3,+c=��~��-��MY�o�2�6�����Ƃi��ݴj@�1B�o�0���l��z΃�
�������K��Hq`���k�5z�(4��ŝ~Q�Ib���(�������(�W�����`�L���cb�F�;��Ts�Op+<o�G�������;��a�T�Y���ס�#�=/��s�?:�Ή>z����i(H���¾�O:Y��f"g�)AF��C�� 0O@�j���o���7��5YkM�{�0��`�̪�������0�S�aBJ�[�BI�X�W�Cl���B;����c��[>�w��{��6bX�Ef:��,-kW��eNK;&�f5����%�&����n� �x�a�_����ɩ��dsZ? 㗧[q!S1M����������`㨳�eJ�'��	Fw�)�zoC;O_���{�Q��qr~����_�VI}B �c�(o���"0�����'ɉ"�u�	/|'�`��,ū^<���Pk��`�5��Y�tWW�Ϯ�QH�l��-ǽvu�pc8�scY�PN���'���i�e�2�8�7��ehX��n������r�[Z �7> ��h�u�tsY�����K�Ϸ�,\�2����8��]�d,��.OOS����W�M*p��Z�G+�t�G�?�f�u�MM/4p�χ���a	��%_^��*���]���q��TT(�R|�[�&_Iad�Ń�xÚ������5�י�8�<��ju�	�ǵN7�q��7��#ѝ0�pd�>?�L���jt#�^���ӂ��������j���O?�����=HP�9!e�hF�������l�#�J����r�R���BAe?�x䜡:������%�e�b#�s<vK��Ϗý3%��O�ඣ"��F�R�3��E�*��ԫ��E_5�5RS��^�2���=��g=,栺m��4+��'��r
�T�f���<`Z�C8o��dFB��͇�8�@�G�7���&��k���4�sƜ��?2%�+�HR(��7-GMrrM���Z��}RQgT��5�X�_�g��x5�e�y�5�%���V�*+� Jn��{	�^�����i��H��J���v����J����0