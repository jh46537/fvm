��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���a�%�sK��h���/a�y���v��=��w�����:�y$f�*,�RA\��S����ћW;�U���T�Ǔ�q�0`�eѓ^����8YU?to�Pb�I�����9���������:����l	�~�Y���)���L8�|m[P��Z�ј�79Ӄ���e<���_�����^�2�����
v��;�{a�<Vx3�-�����ٍ��/�[�mg������o2����@�m�e�?ኂ��l:g(Ozl8S
�-�CW�gF�5�դ����>��'K�:���ϵA��8�l��X�0S����b&�7�%)����!�h/Sq�㾴.��"��w[�Xe2�.ƿm�?�g0ۉ.�*9D��>[ˬ�?]#��m�g+��;��Lb�W%��"�����n�F�`��VW��th��Y*�1 ��a�|�!D�+�iN�=b|�A2A����x���DŶXW��{p1��Ƌ��f��QBw��G�t/AG�<ki����ο�%#���G-nih(��Z����=td3���XSGr�� \�p�n;�&u��@���.����$����P��x��p��ˆ��o�5Eheup\���|��o�z,�T���%�+�5^���D����f�����HY��
����	d��$)q��#�W=���n9��))P��e7I�j+��#��_~���Sx�y�&PS+���gΝ��n��9�;��-�vI��4��WZ�uGٿ��`!�2��p�D�LJ=�E��{�2����������p����'��]f�Kh?�x� �_��ú?`y��9Es_�����嶡KFF%��菚0ٰa����w�Eű?���WM�ے���ˈhǎ}�P�ߛ���T�$N�W0.nEY�I�R�
^6wse ���$w�=���PBM\� ��k/d�h��<�u�
�]��~�K�;�`�DE�_7A�����(�X�be��l9<wR�F��,�������w�ǅQ ���̱c����!*C�k��7�
���*i�|��deDҶ���%�ŧM��+�I�F���b,�Z
7M���y:9����in5]}q�}x/�̩bf�;�ך���h��+��a@u��'��/�/�4���t��T6 ec�Й�J���>�ȫ���ӌC�s��\y����M��_��4��un����8��J�%I��_�s�P�7��R�B��I#���	�E��<��C�R!�"��踙��}j.>�RBT��غ_w��.�:e%0�D�~ڲQ�g����*|�T];U��:!���`5�S4dU��mEd�}��c�~%�\��]��8vt�$(Ic}��wA9�] g7��6%���Rw�x�������KgOʣL��H���c�(�6�[j�8�[��8L�*���[��'�Ʒ0�>˩W��:EP4tm&"�>���Q\�A���&!X�{G�	ߧS�}Vs����I��Ļ�:��A1�6����2��2�,`y��Y ��⎫
S]w���V�c\4�=+�aE����z��m{��7QƂ���z U��1��|�M�[Ƈ�z�M"?�]�xe�⪑� �~�t �wPb8а>�g�ҡ9��"�r���a)�h].zٜ�#��E~�
z���<܇��E�����1�2�23'DE��_�g�8��"h��.�՜���J�F0��̯y�CJ��P8 �H�21����w������ǀ��������autp�_g)`δd�wc���h9�ݔye��]��ܽ�%%�����W%������MǴ	T��� ���TV]���iXG�>�4a��(:(����.� X��gk��f�K���Mې���I���ϊ��K�X���[�L�ğ�h̗j�>��d@�D��E��ꗏ��Yc⚘P��Og C�HO���be��o>t�,?5<*���3�"h��éO��MD���c>̵����5W	B8�֙��6�����M5�n\-��\.{���&�}�%�����}J�6�q9Ύ���=,�	��]1S���*��4�i�Es0����E'����}��� e^������i&	���d�죴@�����7&���c��e�\�O(ıdO��Z*�M��I��!WVҸ�(^	�Ǯk7c<����{�Wɱ�гmH��fЩ����F�+{MǕ ��G�䷃Ə��2�J
;�>:�̯"��rM*l�`p�OIh���=Z�X"�2d��(�~Eʑ|6V6���h�8���-�hDv��0ed|S�<�E6��H�� �z�[<-@��#l?)]j
!��)|l�`��|!M�AC	��R����"F�����a{����U��Dʅ|�bq�g��I(7��Y<<��ʅ}W����JKU�L,қ����?��Q�Ԭ�:",Q����s�P��Aќ�+��iڳV�$Ѥ��]���
�. �nO3����y�3���R�r�%T�(20�&&��Į\�������+�k��kT���o�r��I~��o���\u돽z`��������4g������M^��]ןiqܑ��e�����@�{��X��Ff�@)��A�  �<��� �3[��=τ�B��+���
[Ճ�@�L���/[��c���!QՒv@;�d�����R�='��m�r����WS\OB���f��	 ��`8��F�t~��1N�z��ݽ` "5�KCAsG���N�{6/!�
�r�'���w�!Cj��J`��D�p�y�$f/��I'^&�SY���߸u�A�>'��������R-o���Z�U�+Q=��pL���\�ʂA\������o��'��� �Ku��l�c�.�� �֬i7�NG1��B�(d(���]Z�V���`lpt�=�$NSR�[x������S�nW��֌ �ַ�f�T�N����P�R�(*n��	)/�Tz(h+����G�N��ȏe�}��i�P�ӞE����������.���l��K�������!�-��Phw�"�ug�Դ6�f��.5iY+d�eo,=����e�~�L��^߮r��ڍFՕU�C����d{�ۃj���uJ-�aB�iJf0�H�ȁ����c�I�I/%**d,E�eoD�SX��ſ:�k �����������KxPi�:p"S9���?%�Eht"��e_�����F�먞̢�xO��u��LYl�+���V��K�B�Ü�*'�v���{G!�=r���uN6�Y�s�F5O�$'��X'-�e����T�N�x.���9�MߧXY�v� _j�"�)@ �Pr	�{\�о�4���M�/S����C��a��yDv��99�o1L~��<�<�@� ��(�����W�f��۱�e�/���n�k_6��4��L��ا�;����5!�Ae�/�!8N�J\��h�l^�tB?pb#����v���9�������Q��r�����W2f�z��:\�aS�P�՚�N����Z����0���)^&
�*q��R�DfOA�L���[g��ŏ"�P�z��ݧ��ijo�w�;�%9ˁ~ K�� H�V���d��֋�J�����v��D���2^ƽ�ӌFC���~4Vlx:�#GɁ�� �
���r&��p3���K(Zy��~ɸ= ��8W�{����$��k�!�������d#%I�j:�l��}�����X��ui�l �̒�YXsV,�4"���Dk��j��/w/��͹�ft�}�]8=���S����s�LPr�P��qU�����Ƃ�&'�QuM|�OfD!�+���M�#�s|�o������@����Ooci�n���-������T��ٰ U+��:�f�����@m�Z �0j��툁<Э��h�'O�F���,٢�3Zo��/U�4r�NE�� �&��R
��g�]�z��	�Hĸe�Sn�Ccdڴ 5��S�d��J��T�^�t����Ϸ�&��〣��-�y�w1��X��uާ��p�q���`&���@�ˌ�>�vm�Ϡ	�{劖W��h���V����������X�a/�u�D��S-z2j8�t~>���9n��`�d�o�<Y�����$��o>���a �E����j��$���}E"��'��ቕ�>ټ�aM���Լ�xSn]�L��ڬ��őw
�P[W�x[W���14�6��j3x[�դ2�T�z���%�"{��W�u�ⷤ�EHLzɿ6�nz
o��t��F�ˣW���2�� ��J/GE6EV��79�6x�P}u�t��q����w�f�7�-K�����RA�wJ� �.ѫc���u\Qj��V����]�/Tp?}
;�������f�ٚ(t�]��������#��啕ߑ�z5 ��ǜ��v�"����(̡�B͜~ɻ�c��vNʳ�8�WQ����²��s��ʘ|.#��yr3��W�`��OIX���5RR�-g�	�����Z`c��b+qy��������^�ǧm�h9$0��z�\���&� p�K٪u�I։�������Q *���?|�� �¡�
D����{,ĭ�pv��3|̼˶X�u6��d� �V�q����߻F���a��$[�]��lo������ɿ*ò���xOa)��e?qI��M<�M��TA@C����!������X]	�naȄ����VҘO<}��Yn�)����Ɋc��u �j|��L��nS��/%����2�p��՝�[mÎ���iU=�������3��e�K�dG�]�Ȉ��-)�x)�B��?`B�X!�����8�f�%[�'(L�r�����L���6��;�؈��C�����&]�n�����&�`%��M�O�f�?�����P1��!�U��hg�3���Hb��ix}�&rWC�p}
M� 3������nN`�=��I�k~���xtX��1����JU�^�o�:J��N��8�g+��)7�K��It��c��/�%=;�P�ţ2_�,R�	�IX²�>7U7\�M#/����A��o�CF��(�hcN9D�9øb���G����9���܃خ�\U��˳���8U�P�uo��5�o��A���j=�LØ�8��y����5����c*U5�;�)� x�̢��2�m��8�.J&���g�����½9�m.�7QMe��$� $!�����`@N�cK�� ���I0s�5�z�;�v�1�4o�Xĵ
&��Y���8�~��׾�I�T�F�~���K��a `>�*�L��Ҳ+����ι%��i{ƥ����ꡕ�a�o��1."�?�w���&�>�y<����*Ҿ��/Wu��M�.�J�����N#�H�(�{��Vv�%����b+N�($1�5e |���'Y{h�N!�,���ȱ ���3�72��Lh�cH�IgH�?���W6wh��J�h���<����ͺ��G'Z:6���?������vnx�qrB�LN��tV���
 �����;�A<&d��<@�@_X��eY��M��S9�5��}9k��R"3�5�3B���X��ӎG7U����`��$)�h
���V�=��QjI��m`h.D~H����]\à0��-05f;7'�C����xk�E���>Jv�5�R[��T^'㪾��K�a�ߨ���gr$3�
��m*]}g2�7�>mU�%�y��#�]�PXĒ|.{z��]y< ������o��C���-]���B��k��µ��ᚌ��nߌ��`�9��?��T���*��d�7��/M����zy��K�<�l����
�P�!��*�`s�nq�H��*�ء:��]���@r#9 V�D�Y�G�hI
îˑ��-��%g��菡�1ŵz{-��n�� �A��ܾ��X�y��B�;�ĲP76� ſڪ�r��Єf[���d��lη��EO��i�ym���0�~�Դ!�-�P�WZ3�Y�L
j�;�
r�`x|M��]�pA,�4~�@�^B��!���:T��[��	C-rMDS	�X�b���r��>�5�@GԂ�s;@?��j}�ԑ��-~�x��������L���+<1��z��-���7���)�*� ߠpVI��C<�o	�I�ED���8�kDM�+,dէ2�bg��i�Vk�)�V#�^4S��:��$��Jֲ���Y��8���}6$/�?����( ���"*��H��X�ڑ�����G�q�U�7�6�vk�a9T��C��Q�DSiPD6���^{��#���O�)W
�X��a�M�?���1r����aބf ]�f��h� i��-��i�$nWZ�}8N��ӛ��5�h�ħ�xk���R� �2i�O����T���ۙ��Tw�oi�DO���^{�!��L��,��Ɇ��� �AG�«Vo{����7r�{���G|�ࡠς��T�>AIݣoV���P8w����_K��5c��o�dt��ܜ��B�h�M�zn}_>�'��jz�޿	�Q�v�@~N��zkl����D��&�U�a�?� M��������w����s�EJd�dD�����zCy�t�=��|����6kn"��T�r� �,D�|_+FԲ}ce�<���(O6�[�j�'�P��X:v�4G܌4o�}�o߁>0�f�QƧ�WZ�d��P��s�ۍ�J�#�Nbe:H�CP�̵{TE-]���C�T��$s���gҢAATD�fl��g�"�����ik"e��'��iJfڽ�zأ�N�Y4u��r���F��
|��tko��e�Q��O?�m�bT�=�K�v:�+u��F��̏�\�����7����M�p+@��X���8(��mVW#֐j0���*P��⣫�=� cr'0��jȦ�����'rmi
v��q���hu� l�%����Ê��|i�r�]���5p���J|����[���E]�W,x;03J����V�ݯY.ۅ(�x�C	<>�F����������}V_��5�hA��C4�\�q�����_=Y �}W��Qd����~�>z��Υ��:�������!�M4g�Ў$� ���^�S,����νG���e��A~I�`h(:��S�Ǥ��߷S4�|�z��D�i�r%
��K�J��}ى.����_\�o��'�ƅy?	f��:�2�<$�1C���9��@rX���f�G��q���	��uβ:K��qeݷ�\Hr+e���%X͡��nU��:V=��rUw������U&�୿+a�T@�C�.x2f;X��B�G���N��&���\Hb��D��cx�y(�UX����E�պ;����f�����L��FT��T� �R�ю\\9
��/�=����=��}�¥W~	�b�y�l�D(ca���z�^4���>���n>�9��{僾i���ɿ����U��,�;Eg���7E�Z��;Ry��W5��ڞ�[GcP�"TyW�#F��z?��^�g-%�cw��E�o�7�,�]Γ'l:�,SSg�#;2!?6�s1l^��p�~�fb=g��t�[S��\U
�2>�;y"'�;C�BA��^չ-���Św�|J�K�ӹ7��~r:��А��w�a��f��\���Ǖڋ�g�3P.]0��C,�����e�G��Lo]^���Z�@2�X�Ȼ4tl�V�GP��/�A����}�S��`�E��6`�y���`���)�S�c\��~qz1Yk��Z���*q*��Q8X�P��#v+	1&?ߛO�yŲ�:�+�M�9"a��Dg�wC�穬GQ<\�`��h��3c��~�p���Ay��{�ۻ
���c�솇�iꃩQgW߶��:�Fꩅn�����;���Z��g�dI+�gM~ߎw��{}���ɪ�hPj����n��} ���(uo��,�q�lH� q�X�i�N���8�:wsK�#�% �~B⸦�ɬ'ת��.���N�+^�d��j�����j�g��9X� :jsy#�Ř2!5�ӯ�Y����},��$3C^�Z���X'b��r�c���6�*�({@��ͽ+�c �;S�t٦����P�NP�N�\vO���?+䗣�^�`�a�|J2c��lʔ�k1�E�w�6�P�_�������X�Y�z�I��Z�����Q�L�����Єq����?;%*�_hQ�I������h���u��y�(����;:����lg��o�$����D��BS�m�
�sgn��=s��<I
SL��+�|�}��6��������!Y���s��'[Ȧ>Fd.���P�U��?�+�x��w�î)�C��[nB�MAύ����mMj��x�p�H	���"~׉��C	���c�/k�����֞���H+"5Q5�`f�+�WM�ܬh��6��Lϭ~����3�:����v���>J��l��.�y;�����p5Gm��g?�K�)ںM��ʂ���1y��^lRh�0�s^�DiBuAϨ�s��+��z�Ʀ(�o�!�v׃KF�D��&�Y����j�:��(b"fT����RA�"�^�o8*�I���v-�|�̗��'? �R?�B�Xbm��PE�v��Q/���T�l��M���!��Jf7�%�ѫ>���������OS����R�^�s��t	��N����bR]�}���႗e٨�J(R6�1�����4�)�m �I6�7��;��G��R�� ��&m�����PVP�Q�0u����*?a���Pc���<7~�m/���k�SQ�H;a����U'��G>�J�zP�~���7��}<�Eh��8,Z�vj��VT%�8e���u�)X(Ī�(��|jZ�A�Z�u怕;W������Z��˒�	9rȘO�-{�1\|�5�E���.u�Myx�0�b�T���91���KW���s/}�[3Y�qK�~ӗ�\�>�C�������[V� ��(�\Ć.��Vj 4�rZ�	蔋M_�o�Ұ�t#��W�Q,��|�0��~~�շ({[R�-
��*�'��nE�q�W���Y͘`�x�h<���g�
����yqkH����R�f2��Z`�@�ْ{l��Q޾��M�����O�M�0�T.�'/��ݖwv�{��e�A�f�f��0s���s@Cd���W(`�,e���2!r�z���m�i�TJ4c"SF�W�aB;G�;��U�����+�Ւf:|���q	�����|�f���Dg�^픱��Ef�:Ƨ�;v��-��0}Z���s~5�������K.�`=S
����q��fP8WiV{�����*��*��9|�~��qlwȖV�������&�i٫m�rêwي-���%��ߛ��Y�Qrx(�Ls<k/RZإ!l�VED�Ϛߩ�2цjj�%�C��
ڇ[;߭.�Fy+���5���IM�_��U�vÃ[ޖ<Q�$���붝J�����ȐB��dt����Cd�]�����m���Ax�����t.d-��U�R�Ie�-���\���;¾�.��1��y�tQ�Ut�����
42b�Gmm�B��V�\S\�k�z�XOk%��ANl�B*;��F3T��nb�H��w�["�6{��GVl�"�l`�G"~@���=û\ɮlL�)R���Vq�Ü�KƸ}(a��J�݉�eG���]4���ɒ��~�k�9�ؘ���g���9�{&��69njz$�m��Y�zu.�A����l����җ���������	Y�֠&%��gy9����Z�p�ex������+9�z�X����2^�	d^�ʡX��41=ݵ�������O�#�@I���ńk)t���jk�#IռT�$��)ɴ��(,-��}�1_b����(-JzA���7��(Z�h�p��8(���tJV�3���MF�8�۔sk$�u�4ב2V+�H7�Ç%tA�Z;�ٕ���k����ň�u.IM�q�g(���~�LT�,{���~���?hw<h��L<wc��gY�m��Oخ
�`X�!������)����'�oO�2�B\ ��øaw��L�$�N��#5J+n�R���	b�鋱C��u�{�zk�L3���x�FK����ֹ�]�0�`�,��9hB��y4�9Hk�jzB�G�����y�,9{1̣퍸v�^�u���;�F����&:��jV�В K�(���8�a\�W�W����ΟtS֩�2����.Zsѻ�S9T�� 2��W�=��Yc|��dM>�~��uu,W{���h��hm3��X����o�H7�ᶓ���=&��Y�ټ���c>����0 d�o���|ȦQ�HK'qܭ;��nR��f�Eg*�!e�	���2��b_�]ڕ�_����I)K��H�&�x��u����g���%����h�:29j�k�k=��uLns͏/��>�������Xte�{��r�+�U1P%��+����"��o� s+����Ͽ&AN�'��n�%g�ӆ��f6�?��%�G�-I�*�ȃ(,�Z�6MO4���-�:�
��B�PҐt�8dDКhe�Ո̼�5ؼ�L˼�t�1[��h�.8�ז%�,L�a��W��(V�w�(�
d�	e/�nhT����^�6�L�-�0-��
t�N��g0X�nj�E�8�Cqw�RP^#�t��4=d\�jCA�>��}!�~K�m�ebs��@��5�fy�ҠF�GR���+nR�L�}�!����$�D�i�y�;������v*k(y�����O����;�h��� ����dm���Z�bi(d�
B�i����xW��F�[͋4�l�a�J	��g}B�T�C�o3*�{���ŴÖ��j�X��z��VQ�-����2��#B�#w]�2�GH_�>�k]��j�0�I���gM|�mYe�'d���������丄�*�Scs%9l���E,^��w��� �lX��\�r�tL"��N1�oX8�p؊V����~���Ì]��2�9�ޭ���˵�ͩ�Z|�:�O�d��Bc	���r��K�#K¨�L�{>�����-T�e��7o:�^� �q�ˁ�MR	/s4��Җ�:���z��6�K|����Չ\I V���%~*�;r�[�?#���T����f-;��Y�0��R��8��K����0��ּ٘u�*a>����@[4Zl���w���Q�˹�g�6�0��ɹ�U��c�==y�xlM��z���CW�Ӱ�5��-?Wc�[U'^"��}^��Zn��6��d�롛��C_��Ф�E�]ש����v*6�jİj+v�<���[n�"�C�QLX�L��۹��wxDM)7�S4L��S�y�3��(o�uoP�C��� 4��. ���^��ĭ��lw/��|����ct*�c�@.���{( 3�f�&L�ӪO��ߩ\m!�ߚtn̎[��f�4���i���pk�R[B0��t ی�v6[I+�+�!��9�}H �e�yb�İ�eB<��tD�IŠ�@���m�Gɏ�섯_nC�U�g�?vi�1�_��z��|%��>Y'�b���� ϯ�ԡ3�ss^�E^� @�v^���aldj�ը?@��`O��y���xs	���-��dW��v���S��fh9�Pl�df�*�"��Lț����gG���^|��<f�]���$R�����ݾF�������My
�b8��pPM��$���O����0�R�Tn�y�Ӻ>��>����AA��N�&p3G�o��-}�<��(�|~��a�=}(~U��n5��9����˖����o�� �=T�V�Mz�n���u�:�`{�̬��� �t��t��N�:�4\{�(Z��s�'�xqk��Ƃ�G��sV��3X�x��$ZP�_��7lGa�7���Y��h+���#�g��x�嵋�#�B�ƺ���h�1;�au����i��Cf'�´�0���b��4�o~XN�pPo�c��mo�����o�� ;3���T��w�O^3܍˛p�L]�*��Xg}S����; ��q����������A�����sS4�`�Es;�j�by������z���=�iOSƽ�ءF�DS�����{�� +��l4�P���z��@���IU��2�"����C˚��S�/FR�T`����J�E��Rm��� q^�9�0CF*�X��H��tI����&%���7r�$7DэJ���Y��%�O��"D�3��Nl���b�D�:�aE��^����}�w��v��k�E�Lo!�N� �҃�	�/)1��nI�_��K�/WQ�$M�%K�����¢�;�B����1��fg L�^F���g~��XpV�����cBP�Ւ������o;��z���(�)/�W���H��O2U��\���$p^�O���X�b,�;1u!���Y�z^(�$\���X�"�L��T>��D߅�L%bH����S"2�3F`���n��������c�Xll�X��6��+�n0�di����tEW�.	\�~���D&��(����J���b!�G��A����2�~pq�'2�q�p�����%ˑ,�Ƣ�K�zg��Pg���r��}���4ۈ{��ȃ��en-#8e�I���H�"���'$k^�Ɍר�M�Y�&y�v�ͳ�"WS�A�^:�SM�'�)�Lo�&;M�E�ܬϝf�)��c�v��Τ%�hb��
�2P��|�7M���U;٦���1}��L���	<O0:0C��A��@q#�"��ڕ������f�]���Qa�T�|�z.�G��,y��|�{v-a����|?Lg���4�O� Pbsw̃��On*>�_���W������Gsb@�_3�9񁃂��R�0r +� �Vͧ2�Q�I���3��Mn��	�^�]���c8"��<|�W��{��c�ҋ����Cp�WB(�V̂յM*��&�]_E >(]8۠oJ?P9��?[��l�Le-d)!Z��݇�,r���I���.�<�k�2	���������{F�nbaO���UR���<Bs����:+���bi��]�pu�g�d`�#�&�Ԭĩl��p�GYE�Ŗ�-�����y8�,�����yh�G^R�1\�.�C���ф [��fG����R1D&N0��"@�y�ŇK�s���
�n���|B��\m���6eX�>����${�ν�:|�_CVp�X��m�d�'�ȊM��e�O�D�2 �&��9��~^$�?:I��W"�&���9C�X\p6�������GƑ��(3н4{#�D[)5"�R��2�����Fe��e����(���A��i˾.'�ԑ�j��ؐ]��Z3@��k�w�Ӱ*����[���!�I��셓o{�l\��.L� �n�2=~������l��77E��H�l���3�ż
"�ؠP��Ñe�����f���X�L� 3�֮b��Q����CL�#!3N(~�soIGi9x��+/��8�B\�N��s2B�+
���P�`wa�i(q�ˇI^�L7%Ljn[ȸ�.�g6��)j�E_b�Ag?�5^�<��Lᵥ��&�̐��Bh(5UB�ѯp��\->���[rrJN0[K�g��pn!O%.�_X�.H�@/u��m�6�����L+W���G�k�OY�Żz^&�e���?g�D��VlNa������	�&�=2v���$l�������w��«��l��tY���*��|���2�|؈�s��L۾��d�c�N��|e4����夐#ӟaVI�殖
���\��e�ׇ�Jqf+g8�!��"�%H��1����Z�nm(��CG�|�S8;@�'�.|~g���&��3���v�_�&��9-��b�HiI�t��OyZɶ��Qgv��u��A=i�Q����j@𥡒/��L!@{$0
�W�ܫ�	�z��|8ωJ�[��<���9bK>�GA-���p�6�<�xi��n����H#��Ø�u%-�Mhv#O11�KhD>���\Z4T�I��.��ΩU�?�Ƀ�\�=	��]��sq���\���nO㙤��kO��L'"�Ǌ�4O?r���zT�Q�g��
]���'���".�e�,nR�`�je{-J��=�kj��?�`>1
XOX9*�� *M���o{_K���N���;^g,��iZGy�DC�0/���vf����ú����W���e���ޥ�쩱JKDK�����ӛj��h�������G�f?��
�nw�n�����|z��b,.G���ۦ�I\]�h]��PM�`�D+ᅁ�)|oG�R	Y5x^��h��b��^s��O��,�Lwù	���7���R�k�3�=mL'׾�!E�#�y���(C�'��`��|yfc��0�,���Ml!�f.��*K���ﶱ���7��[ �h���E|�����P)o��Υ�]�ȁW�����<��1�"��$1Ɛ��9*�j{���C���ɗ���)�k�<#�@�M�H�۝���̓Eg9��9��+�m=�a�	�	C�ߟ�sq��A
̀#�z%��=�_��EK�R��}�G� ���牜V7�j�J،@I,����4J�z��� ���HlBz��P؞�V��: K���߳�����똋M����u�QC-fY�3�FY�fe�o^΋���'C��(����&��'�HWr���ީ�hձop_�W~S턽rE�P7�V������XH�`�G��_���������3y� 0l�*��
,U`��W7.�re���{�%�h_k�o��!L��%�ۼ=�s�LH��4�u��¢��3��6�VoKS�Q� ��l^�Fz�%�ߋB�!5�VFPp�c�t�<����mA&�/�G�¾��6He�ch����^�d�Ty�5��k�)e��� 8`�T�i�ڷT������U<����iGU2�D�N��0� �@3��aUj��}�t�w�3��f5C=5��홻�8@�~ "Y��	U���O�i:V�Wc=���iPi���+y|��lą���f���D��o#��c�X.5 ���شͻþ���Zy�ꐷ`3��='�
��L����nD�3�b?Ĩ릸�y܏��Iy�W��C����V��\�J�s�o�8��tj�N�����͈_�\S#O�q�S�Q����9e��8F��2D�-�����@�?�D��=*p~)�"ӵV,����S����Q��J��~�jJᙞ����}x������Zw�M�#�O�Rw=�@H�Bk�v���J���e�u�(DԎp�z��q�o�	�4c���U����o�q���c�$pF�^Qd��9�VJ�S� -^�TD_@P.3׀V�&�-9ĞL�`?��I!"3ٌ��~No��g�b��U�-Q�D�U��a\�Մ�=�N����M�0��s�t����9L5��?κ~�S�.��� ��]��,�)e0RI�A��p�{Vy��rg��� ��><����=��1���g%���빹w}@�b�	�
�Ua9�����  v�^s�Iͭl|����N�[[�ɵ�.Nـ\�'�,�I�Q����'��g���wZ����I.R0d��K�~2��xߑ"�s��5K�G��F�a8Ԅ��·6��_���Οvc�n��N�����-�ڮ��(�n���V+gd�Rj�s��̬L��l��-ٖ�# w-���F�ͧꡌ��a 'G[�ITG�$U����0�5��������*]O���&�BΊE8O�A�a��22��i�T����SOm�Ϧ�3�mz%�}i	�t�5�R�E/R�bȹ#��]r�
e����pW�0��&4&�n˰)�xA���7������CY�:�1m���C��(��m/���ID��n�Tt�7���v�ۼ�\:'5ѣw,̲��������&g��]�A!�n~��ha�Of0�gi9C
 m�����U�*&�ˁ���sn-�]vN���s�����|��