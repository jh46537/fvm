��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��ߨ�=�]	7�N�)3�M�Ρ� ��B
�i�k<֐�1(�/h�"�+r��ҏ�X�fИ`��6.[���L����Sg�$|����x���
����v�95|b�fUw��e#���`r�|�QZ3E�*��e$㩥�֢H.���a9��[��}h��P����{7DI�y*��f`�K�>BW�{�����z��<�	&u2��<��q-F�zB��0�t�c\��L��U�Z���T�u�o|^��G�)�=�d�so,�yr���o�L1/�%�o ��)X�A��f�H9=<~�/�f�ԑb��ޝ��X����3�5�_�O��AX��ˡr*`�}�1	��83pPR]�B~ƫ�ug�D����2�9� �����/E=4�pzD�<QCY^��}h[
KV �����{��g$_�_@�6��F��7c��m^�<E��"��G���e�j0O�;X��q����ۄ��ˍ�Zo�@�J�?�,٭�'�P�� �e�������X���ԁמ��TӱVl#��E�1at�Z�����'���H>�=�탛�^�\�l���F���博Go-�*TI�-\(�:�����:d#o�Ű�mtmK�rc��?��a�:Íf�gR&����č�Y��:v;��2ϵ;	� Jq3z�m�x���S|ۍ��[O�:���~ŷ˛#GZ�/���o��<��|Cl�ȹ�U�� l@�c� ;(C)ЮS�܆Y#�@���H�shn��Ȏ�bЮ�bu�.�y�)nC��ypv���s��x-�u]�����])��C��͏��*�V�Sx.���3�e:���ҿ�,���� ��B�S[����� ���7�XmE7����Is��O��*>��RJ�!�b���䙸��j�ۑ�q��F��de�-��(��~[)6�ϳ��FXK�߇cnN�Ƒ)�G?!�jz�`s��^C��&�\��� q^R�y��C{O� w�_���N(,��!0z,+������ ��A��G+���f�G����$�A���K����$nMy�˓K�x_��Bq����%,�n;諆Rk�TW�J%����6��9�ma��kl�h�&eU�R.m�%RPRWΩA���"�Q��~ r���:x!�݋��^G#��:]��M�����a�q�5	Ő1���͊*��@�0Y�`P�ݪ1�1S9��&,Y���f"�wb=L���J�R[��B��N�=���fAʝT�
��LN��xm�7�}��"�]�wJ_w�+i�~+�Bu!�*��@��bB� ���œ�{��W��ß�5��1�9/*�%�!�5g��__�?��KH���r3�-f�.	Sw`��VS��֢k�/��6�y����p��T�U�	�o�Vh�%���{*\z.5^�K� _��2!�������*���R�V�PUF.�p�7M�D�C�1���q~��kod�K:�&X�	��+�ؐ��i3�ܔ7S���mSu�P7�,�yz�#xw�&p�Y�V��d��J<ަ��fׯ6���昒��k��C 6�]�#z�8����7��O���o��ɬݬ�N2�d)K���D���if��U���QR�o�4��Y�5��P%��蕱�Z� >Ȃ]]1�RT�ĔҨ��77*�<}'&�$=W���pn�)��9�h@����W?�w��%@�!��q�����N[=gm^$#����W<�k4ff���$(�������W=�Q���A���*�N�^睂׃-�S�VW;��/kɨ' �&˲�="x3�Pݱ�p8�+wv�����(�mr�q��ҹ&��J�7:�P��򕞞:�R��qN�ib����
��T��knWk�ON��X�+�v���n)�UOH~����6�a��Gc]��7O�dT-�Fϗ ]�V=;=��$3k��#��ZȬ�j:��H��}��0������~�q�$P��N��z��p~�ކ�l�a1�@�
{�E��A�}�)e_8�{��4J�41�e@Е���C�Z�],��a��x$@-���5��� )`N�WSfV��!�t6���T5�i;��ѱ���l��B�ƫʼ�g�{�mrMv��g�~+�S\��$B�A+��3CttH��P%���ݣDq���띀�P%���
�(���
`KAG����ôHQ��ȓ�<��aͼ ��vס�(RӘ&��N@������c[�V���86�	�0��s�Uv�Z�2��S��=�Ɯ30������P��uL��U܏���,�aN�X0?^�.ʅcC�B�v&~��\A����g���*��3^7%LRQv�@��3�c�+�=�R}/�5��q��"�T��U�� �3�E�Y��O�����6�8ڻ�ȰěKL�R\`���K,[�H�L��?24�9�5S��P����~�nO���z��ɍQq8�'Η�W>�mW΀&;���ǣ��e����~,$��8< }÷�^&Rˡϥ���ty���6��"t7z@ס\5GK	��AWnӜ֊�mz�Fҥ�0���C4��&�c�>�ܣ��]��~^L����^�����wH�D�M�[��t=�����v��č	\��a���}���9��>���i�����U�����I?{����l1zS��к�Jq����M�D_�!�f��V
|�&}���@�#���ygQ_nq���y���v����e��]n"\$��{���	*����EݪژI�C��C{�L����*.��Bc�ƣ ���"/�I�$.[��'�}��3t�׬�Y��KY��)���Fq������NU���HYgX��A�"dSwC��o��^L���-������9���t��-���P�4�Y��o	��AS�P�&��:���~L��Ԝ�G�ؚ�b~���bI��.�z��k6�u~-cE��ʪ|��3_����x�;���]�jAf�(|�'�8]��i�^�_Z����6�xUs |FM�Bc��	���sk��c���r��vʅ�DX#� ��?�1l�v�4�z�f*����=�b�#��U��@�L��	���?��W@�̅թ���<
���-9�N���3ԇ udp��FmŽ�J��F�8=��|qd���gj�@������e~�vyc"���p���]x��ˊ�D����粎���[�+U=����X+1��M1�.�@dd��^�J�w�gO�+Xo��Ě_��Y$���{%���J������#-�&^��z�zPF,���C����[Xq6����1�C���s?�� f�u��q�
p5�s6��ԯ�zsv�>JW��m�}a��ȧ^�G��A
e�o�^�^Ѥ��/o��b\PȲ�`�aUPSH�$N�e�6.HD��%'c-J"F^*��o����'���*�a�:;��U�u���ێ�I�q�fv���VX���~�m�g-�쇇в\g_�y����aܿ��)F�V�``wxZ+xML�J��������?�Q�g/���̑�P~��e^-��x$����w�������B��Fٕ�~�>s>}�'+�@��b�0����b�}
vr�ĳV���"dʹ��v��2���+�;lqV���g&������x5��\Q��ɋ��ꩠ
�"�^�{Y�u��߉S���\����-��ݏ�>��L�i��"�=��� �?����o�k�0����k�����[�D���&�L���/��	�*�{M/.I)^rN�pW��|�ã%���4�	���q⢛Y��õ#����2���j��X��^ǩq��N�=�ھQ�W��RA��dK���Cs#U��`&�ED*�~"�ʆy��|ܴy|�TbL
����F�t7A�}�I@<����g䆐w�<PN�`�HwJ�t���(��A���?~�������f.(�Pٵ��6r�r]�;�gq�6ʠ_zd��٨�����W��h��3��}@��Fs�9d���]V��^#U�^2t6q ?���?��CT`�c�H�+/�XI��b9~[i�aN�l=΋%������ת)����߯sͷ���BC��Wn�-4z��u���VL��Ġt�Y$4ɍ	x;L�}�ky��뭆��QY����;���1\`7�m_a����� ٪�?)���QJ��b�:�!JdbSE��:G��;|R/6y�o"��n%��#*� ����٭y�f��H���p*Y��~����{E�i��rJ7�v��3�{�D�� uy�3�YW���$�,�����yY�z�VJ����,�x���z��������= a(>̡ȸ��؇�W�V�m�=Ϗ[|��+�M$s�>��!X3�(�r��!�r������'l��k����4��&��}
���>�����j$��d��a~kWR����e��ǚ}]�B-����0���~c}x�|
�%��X[7*2��b�Kp'���#�Gx���}`e�"M�糝ٰ8�2�KMaf�V�n�R��KN޼/����.�*\H@*͆z~��v�1G��}_=�^�H<��ERV��[������k���:�2@H�����?��-�,���<�'u� ��a!A�
$גT�q�>[jA��Q���Yn�7'225��ĥ���.��^�
��ǁR)NT�R�g��;�� �%��k2�������#��8U4��!�)K��U��.��F���� ��ycE��rW�n���
oc��VyUrP���\�Ḟ�e�p���8�!ڵm�k��5V �u�h�Qxk�X��w�P������ȥ??��O�
�3�>Lr�n�2x9�Jۀ�M��J�&>#
�s?����*�>�i�B���:EnP����H��r��W��W2���6��9�n��*�"#p����A ^!�͓����zt��`T�|�yP���]N���.��8�N�iĥ�2:�}�	-`D�ؔ�ЮO=o�g��QH!Rw1Ϭ8��2�9k�n�����uP���f�#ߑ�v� }��V��c�;��S/��3�'��p���G�f#�b�޸1�r�w!P�jW����e�ㄟC'Ur,�T����&���B�<xl����zY
Ӻ��g�E�BfJ�39zJ5�*/35����o���\Rtf)���4V�d^�(��4��A`S��o#���#Cv�yzI��H6�������e��)�x�Of��!�ma��@�<��嬯ㅭ��T�H���X�/LL﹔"|J� +l�+@И�0;�����G�Z�i�6#".�;A�B�܍�߬'r��4�"x�yV��r�����v~�z��)_��c��l�N ��lT<���P�b��X69��%۪�Jd�AS�a�����5�L�@�	������܈1��p'���\x�Xop��'�����--�$�*�\��q����y��O��E��Pi�)
tzڻ���̆���T*Cl�gs�WŇ�_��Dc�%i�:�&�K���lP��rT�����"S�,���3\^�&
��&�~�\ M��#t�B�,�i͌rzߑ�g3vF$�LnK0��d�EttQ���͏i(�^�h�Z(��x��!����-ĸ��*2����-�q��V?��C�oC��^ d�����Y�+���$*��<E��ut�/���r�y,2+����z��$q����z�:�tc�%����x��\X->'�0��Np����m_��Zk`t;6�I.�^���I��z�c�F�:�]vQr|��0�w ϕ������ͫ���.��|�j&`YȪW.���R܁�t��vq��O�I���[�c��� ���j±� .B=�8!�(`x� ˇ.�v	�[zsC=�$�<�2���J#�2ȾEH :��A[� �3�x�١��������5T�2@W�%����HG���A��l�&ҷh�#�\Ը������N8�g�����e����^�4�e	��z����5��Ɓ�!ѥ������Ho#!꿁v�訮�W~W�z	�-��L������=������<;��[g�??/�10�9^^�`l�+�����O�8d�
��[�Q ��1fjϷ�(�~�(`P��U��0A��m�n('?� �L� q-u�ަ��~b��.l�<�G���E
��<&�]�|G�in]�Q����gצ�M[�vuv����x�E%�iK �6��73��c�\��5�� f�V�,I�\g|�3>��J�<i�IbȄ�������yK2Zz���������p���"���ڊ���| �N]^�&�����F �ט>	�9�XM4n�N���fe����'��#�ss/@���J�62jД5����Nݲ��^�=�8���eo��aBfk�?տ|��T;R�t�����?GU�����i:P�E�ޒ��cY�s聪+��Mt�Q����+O5>4�B�udS���"�.��ɐC�­���Hۓ=�G��
c��+����I�.>ȯ�2�&�m>ow�i�}��,Ws�ј��>a>J���(�}���.��s�Y��J��%A1.)�"~X�q�(q�0�����e�LĈM�Ӭ�n��皤�V���)�~�G�P���[毢�Q$l��������E�k� 1��y2�qMj���c�-`j'�)�4��(�����C��Uϊ�!���U"ӡ�O�+���(9�%��s�26+~2{�ۣ�?'���#|e؅W'����}ZS�K�S���v3՘��ʟ�RAUw�_�����V8�|�rdUr�Hp�
����Ka�:RB0�������i ;����)�~��v
J�ڧbD�u�� t� ��I���e��p���s���ﰌTM�[�dN�[f
�[�;�5SL�J�9?7�=��t�1��_�������92�,�[%�4>1�B������CBk%�"03H�q� (�C�j��m�� ��Nt�N�j����U)����m�ҥ���]�����M�"������ˉi<C�>�dw�0pE N�Æ�gP������bͲ�����
 WYB��u>��bR�dU�kc��$6G���aE�j8���S��o��0����ںnH�p����wc�#g���~)ͲH��x�=��5Y��k(S7%
�p�;���gf�����5�+��13nn��fo����r�@�6�D�C�$��n�B@�%��c�<�:Y�Dw���{�y�������U���w����t`,ٟ�o���)��p�$�hԈ�5�-y�dې��wX�籜-T��NLfn"�͝ oW�K�>C
ѼY��[��?�Fȕ)*���|-*���R}��7b��m>���0�`��7�B翙�O}Kg��2��������:�Ǹs���,��dQ�*�/(ᜥ-�ک7��{t'}lF�4�G��in쾊���p;����&%����,
5�
��>���&%����տ��L#�A�Y�]��'��"(�5Q^�$�o���~{�g˧P�C���,�+�H�u
��h ��L����h(!���&��Iދܨy�땫n��T�lp.��+�ʦ�nhj��z:�@l.T7$3�h6�6m���4Cq��r��PYܦ��S���#�d�[@��K
�@��*��.k� H�	�K �Ć_ꘉ����)��֠��25v�Ѿu���?��t�[*��틼�Dp(�D���0�v�HF7_Lw/�\t9z���27������)��	�A�
)x��\Lu��R����t�L���,_� .���Bƙ�&yL0�j������rr1 aADd�V:�}~^���u��S54F4���k�'��0
Ż��^5�x򇈱�c��sw#0���ڌS�U{�}zcL�
� q��*�i�%�z��.u��q�]Q����t���u�b5��zF���K��DU�!.ng�~�na0@Jt��<<>fhy��uԼ������%��Fk,�O�˽�eÿ�J=����$�%��v��Y[��t�k��Q��������~p��[���wi���q��9��/jj��N���`����0��8F��(ٶ�}X��˘2v��1��t�s�F���h����_G����k��uN]/%��=��*����������QsChD+��e1����q��FrS?iǞ�,ÜD�	�m�(uS�t07�fM\�����f������Tx� 7���gh'00�\�Sf�@�#W{lI�y�)pD�8K��m�"|����B*��aa�r���B�x�����	���$�myr![]�n�ZW�^�Fe/��9�Jf�/�&�1Sz}�K����K.ѝ��ox%0~/إtZ�,�s1ϗK�\����W�9���	i,ʾ|ef�3h�v蛌&^��S8$����aVϥo%*��<(�s��a�(�6�U,X'N3�7�nqLX�5����]j=�љ�؊�ļﵗfb�H�����Q�z��/��J���A��,d��C�^����u�PCŏ��X�`��g,kvp�KWC���o���O�1��v����U�+Zh��zh�x%��?W��CSK͸)����X��4�p�$֙3���������Ϗ�$��/ a�#粪j����N_�T�K�.�|�P�c������g�m�$�р�PmK��+fLpIj�	ph4Ƴ�^$�g
5߬�ǉ��֌؟��r��TѲ$�j�(�֮��"�Ƙ4ge(!���)}8cRh���;����-����4�R���ʬy����u�Z�����������Z�t�{�&|Kʉ(g�z�Y�����]�g�K��~
�I��U[�q����\;��R�v��:��h�w�ukd�]_�EQ��������-M��J񕫬ZDКtj�Q±�'y�4��2�}�%�	��LP��#���@U̮ص��c��i#��8��{Vza�P�vԄ���ק�-�FU�EӇ&�.����'x��� �L]o��x����|��R�
;1��������zDg����˛�2H8��j�*Ŕ��ě�<oQ�IN�d�J���(�E 9v^{_L�\"ts��fqY7�F���<W	�y�E%>����o��a}�3H�;yz�m�uHSN%N�3�Ps[j��Am~v�7$�I},�{a]=6�.䎶�v�ۊ���-��~�Z>9��1���r�{Էhlv�er0�ͳdT�;]t��*Kv���A�/�.PE�㽹5$r�嗽���΀��E�9Y^Y+��J.%�(��B����p�GS��ױ��z���iJf,vҼ��W�:����ͪ|2āY?�o!�`��[?�q��a�I���}�8Z<�� �}��6'W�F�ڼ��Z�`���F9��f��<3�h�7�w"�M �FAkU��n$�%�Z�RRt�Ipbv�k�b�&����&�	{|�7�c*J��h�gM �d[A�����(X%�:��vڦ�E�g:���3��$�;Q�}J[]e����.]��9`�ީ���m���7:!A|��m떎����D�&�c���g+�{��H�[a<��?��jN�ЙW|��R�)��$0�7�ua�6/BW���g�T�d��%d-|�f��99�iW�#�րc�L��A^�a!'�D�Z�I�E�� ��|��^�������U�O��K�!��h^+L�I���?�"�
u�`$�9 z��u����'���Xy���J�ތ�Kpk��(��2��9�*�Ը�^9�Ǔ�0S:����~9[���i�8G
%�Ff�9�$�.Q��QR�L���g(�zB`��5`G �n)�n�tIi�.�N�~�0��<�/�/�e��\`�6�
�k�e�eP���ت�q�,t=���F���1{aE>�S����&x�VC�=,5��B0�dn�r�8b1
�P3�+��%��qa��r-�lU��ڎ<v�ݙ����=Al�Xvݿ��|R�k�o��Pս�����iw$f�r,E��� ��6C/�l"�u,<<ށ�Ǥ$*'�-g"H˦�9ܞP1q0����)�֧G�������PAF~⟈�;��C5��#�{��`Q0C���Pn��*LÅ)��{彊��2`���������l���3BnX)����T�$��<��7>q�n�E=�k�d���l�{\,iq���:��m��qB�5.�Ĕ].EF�kUhK�vH�	�s�7�*c*<��K��UUhG�:�Θv�2�4F�H�w&	���՜Fʹ �S��U�ٟ�X���R�T|Uk��ïq9��#�{&�����o�ҦCJ������+SH$����q����;{Ną���3_��&(�G�j�5�YZ�12�8�r_^��>��%O�d�ЯJ��{�#Tͩ�J
4_֪��b�&�	��b�]�� �*U���_p��To�u�V:���QSOş�p2eDe_'e��ӍlQ�t�g��y��M�b5�n$��X����#��-���= �ٰ��s
�Ո�}7�b�ckbR�0qZ��Q xRTE�Ʊ��P���ֲG��0*ڗ��:j��9�E������S4���z�/O��D�p�������X�꧒^���/�Fb���x��S]B�9�x�=c-=����X�!TWR���{�b�}S'�O����u��N�Cb�1ȿC)k�d����£�����P�%O'"ы�����W���93���g�cz�&r�=_��D�K��\X[b��?�e�KZE����0����,D�Z
UW�'��-]�<�,�VIf��$�V�^3<\~�E֧,=#�s�@hbn�b�i>ȯL%�.+�A����>��hI�顙Y(�4��\���ʜ3�MGT`"�괢_�z>�T�*��S�u7
c2�ݕ��T��{���F��p2����]	K��(����I�.L��Af������c>(��-��5�c�@g�X;��k����E7��O1�t��~LC�x��E�@b�^T-A\ЂWd��3��n�_���d;��t����:�[µ�u-�}��{
(&k�����E3+[3��a����4��ž�@2�p�e\��	rA���� @�TN'�qBVD�6���j�]�&@�����l�H��,��[�"߂��ٵ�{�FE��ʷ���Z��U��TV�4J�7s	BS�)��r���¹aͺG�1W��l<��(٘m�LU��a����Wd٬��M����W_|�:؄�Թ~��^�ʖ��9�� �y҅���ʔ"U#�0ln	����L�̏��)���� �C��B+�9P@�L:o�UR��ruj�uQ�3�+Y�t���C�+���?�@lu�
zz��o�
�Xʮ���B��-w����V ����{��GO��b����c�if56�m�wI�B@n�P{M�]���b꩟�_���wG6�o�`F�͘w�W�[�^�7�=��r�C�2)��_ڡ�k����T���v)��o�*L���z4�G�/�j�ζq�Jw�P`���(ǹj��Zg-��UX��������q�v��bun�X�������ء^��mT�N�GEpa�7�O�I��1�ޜY�u/�/���@:"��l��6sv_�ǂU���-�U���t�x�q�p��fE����q
��n�y\�+%1�B��tݐDђ�<!�E.���eG7ϕ*�,�d쯱g�%9c.ux��S?2c����X�x���s�!��e�����R�9r;#|��T�~������6rc�0�A�|[�M	S:Um�]�9uJ\u�U%�Ϸ�E�K�����z�@�S����HYd�t��u<ʠ0�1�ɷu�s��w�)��֋�TCnn�&4��f�%�9L�\2�-ʬT<2S��!�H <�P�����r��)ڃ�?���SI�f���nꈅ��D�;�� ��-�|��yJ��b�bG������J�<��h<���Id��W/��(��¾�tZo��|�o̓m�ڸ�v��T�ce�Ϻ�"p�3�8�o����PRFF���ڂ�bF=����	����4A-Z�uɯ2�.c��t X��1
�jKf� ��k%��myv���:�Q���(��}�r���C��C�]��;�w���ge�܊2N���f�Y;�:)��!�:� ��5����|	e�>����Ga~M�
@�p7�O�m��_��D��H[�Hг�4�F��3��Մ�a�#~���7�6&ZA�{1�R�͛h�dS-�IKe=���m("�T`���@=�V�%����|a���7�2b����5��J
��(����T��-�V�gi��V�W��JPW�Fk�sk�8����&��E�m��jm��`u)�9z3�2ON�)�w�ï[�����d��	���l�������+M&M�oyQ
t��k'q��鋺_���GHr�X��ᥴ�z�A��.��� �!:��V��t�2�Лhx��&z/�t��$A��\,�D��W�|)��
2��3��~)H9D�ծ��(*�I^��ŷ��T���^�e���!�_�>���$��Wͦ��]Ife�J��>��\�Q�$�a�h���	rٞ�5'dun�`P�~Jb�����˻ )�� ��ig��2N���'����� E�9�l��#�<�N�>�M�N|�}&F*��ů'!^G0e�����JI��.����3*�+��8{�N�z��V���6"�y�J�K�*��h|z[&�a�h��x�݋�Wj�N�����w�C��=��A�ȫ�h�qx�P�u���/�N�6|`����J���G�G��y
�M���Iq=R3��rf��aD���0�9�F֊����-�>R<KLx���NL�AL�:�:?�����0�H��g�x�����
u;���>�F31qK�A�UpY�J���1{�����nY�p���oq ��i�C��lX_��^3��'尥�ح����#�q��uc�^!7�����[hCY�K����4��]�U�3�\�k���@�qQ���?�c�{7 *����ϰ�`;��;�W�;L��b�
Qޑ�nN�r������aU�o*@H]�U���+��#0X�O�% L��� {�{8m��^��������Kw�TV�pm�)�c�b$xmD��m�訄Nȥ��@`��3(��H�xD��A�����P�N�J���~A�����_�B�R�%��;��I��43�#���յ`�΅N�Pጹ\��ltH�`ҡ�
<��L���.7�kH��V`f0�1�ʂ�X4��	 ���r�2AW��Y��K�W��t�!�?߼^}-�\��A���:�8��ڙTS/'��J|��v���5���&+u�"��!L"Ggm�O��R��xu�<�`bą�se'W��W����"X'���ψ��8мϋ�Nv���nؚ�
{3�!{,��O�1%)�;lF�����˟�;t��L縈&�G"@0�9����oJ
��QS�a&/��Q�H��A�c�d�0�ʎh1p��X�����p�M��Љô9Փw����1r:_&�|�;BB3�s1��I4Ie)yM��r�@@��RiT��r��6��-������±5�2�����}����p}ʿ�$]ZɄ�ʢ�6����	Z#�-�MH�{��f�ɥ��g���C�L1ór5E~�� ����'?}A�8_b��!.��O%�Jt�V�h�dZ9Q�o��'�p���G��//�Ho�ur���A�!���@l��f=8Z�mũ�s����묳�h ���k��!�X޲�]�5��f�G3����y����,��1�=jN���^�����W1��O`��5�ޖ9S������:�4���(	ٯnp��7+�Cl���`��x����?g�aỷ�;bm�2d����Ѭ����%˝���
�0���;�I����6�!gXe!�������v�|{w�D_D����ٺ�H��2�n��w�U؟����v}�a{\���u5�N�'5���;��)�����,Bb�t����KpR,�m���w;�Լ=ȃ	�F�Tzl8*�EB�>��ı��/�[��:�a�<�(���iF�k���d�@H�	b�+ ���o�������I6@,���yE������'�3�-8㹫r4��.�'�eΪ������2q��l�D�J�6���<c0.6��b�c��Z��+���N{愸�.���U��^�Ț7 4]�I	���oGU�\����b*������+����n�Lp�%����/LM":���5
Bi�;���!�ۺ��V;��%4� KJ�y����ō�&1"��d��a�ɁF��x�<h�F�yN9�X��}NKG�P���Y��i��Uِ����DE78/+��;6 ��U>��m�|��ٍ>L4$߄�;���1r^ �(����y+a���%"[�R�x]�sj3k�:�ؖ�]�j;s!�����J���K^�����y�4Yh��O���]{;�צ��po�km�ou��Ya�����!�����i�A����l�s]����߇뛖�h�q% ��Ȏ9����.~�dͱ��?l����-�'�n5��}�u['�ޗ��������9��p�pͥ��56�%�c�i2

Ӳ���v- �T�:!uU;�U|0'�oؙVr=�j�PF��UO0yOL�=AK.�G��3�}ϣX%
G�G��S�vw$�v����BX2�/�R ���%K�p�����d���.}\5��'K!����9E��*\�d(��r���������I�Wwz?ɰ9�j3��W�j����T��r��U�ǩ�u��Z۾��ڑ�Q�0�����wFv|:�vJ���O��͠����� ���4�ΉN�Ϧ����̊	K�D�,�˶�]�/��cH�nʔ�z��jvy �{n�E)���e<j�kܣ%JƯ�^�v~%Җ����x���T��nM�f9�8����
��P��l^�{d��:_5��������g�V�(+���~�g�M^x�r��<UOf�"Mo3D.UF����C�&�"X�z�U0(؁ov�:9�fJ��n�-$��0��.ǒ�%t˪�%�j�5f(�ċ�>o����uVF�D_\V̫?�r%� �<ㅐ'� ��$Z�1s/&�2wǥ]�*��Y�g��p�.՟��6F@(��aH0uߝ��g�:���0����,G�=�9p;�:*0��]Ӌ2���/�yD��TWr���KI֬2�)�{6?Zlj�����Dc��s��}���E�b���(_&�Qy��"�b��X@�a�%g��`�����ݱaP�!u˱���@�^��,tyU�c7��h~+^3�zS��jA�j6Zd}��E�f�����2�n�ռ��s�P�9$���%u� ء��w�x)L���9|���/��Mi�k8���a���
����"5%V��v^���5�Vd�Q4�ֵ �f3���fWY���W�ӷ-0��-�_��yp|"TPU�%>�dB�ށ�%�[j4�hG�m�hqIع?V���/bU��4�f���U ����O���7�[�ɭ������!ͭm'^���*��<�d�S�[U��H��"���2�42�ߒ�
J䟰�8B�ԳޗRHGW0D|����7��i��zh�@����Ht���l�lm�l��9y���T�jF۴�q�i)���١��;��^�@������Z0���am��~`�,�H�)�k�\��ۚ�'�ta�+o���u��#Y3�T]2�D6#���uYH�U���:D֎bfz'����3a ���?�+ݤf�0�9X2E��פ���#+�6�!�Kyѽ�A�ĦT���,�����`�jJ��4t�����(��E^Æ�Υ�F3z3�5ڼ�gO�ķZ���E4��54q��IjO���r�ey��=���#;���$ypZ��;{_8���7�?����f]l �\Sgh ����/�^^o\�Lc�4�ޔ+*6���G �M����)�k.q��m�$��'��U�Z������Gs�|Y�'�S��M;:"u�~y�P8�N둶ڒ�D�2�Gg%s�,ߝ����j�t��P�J^z��Z����גN�|'�J�m��p_�~����4o\̌��M�/R�|X�믖jV�7�t�ɚQOH��WU��Y��T���VI��c��S���?�O� ��8#3ر�6x`��
��{u��n�0.�j��F�@WX ��2�y���D$����-%����F��,�~�%8��T�
�s82�ْ�,Io}��M�(<�f���V���?}C��ʐ<�b�Jʙ�aI6���Xz�X�J��� ����BE���c�y�I�,M�Z #x9�5HĝJj��<����{�u�W�{�#g�_'�!�47���( )!ɛI���\���Z]C\G#׫q�USϳQE��D��;����21c�B�o���8�@2����sqB4+��%YE?���E���	�������`�AKB��
$��>��X0P�s���d�*5Ma��A�P ���e��3�J������p�M�����l`�$�J�=�Qܟ��W��s�y��^����=/G��4�?��	��(�6�������!V�Z6�����b~�ޫIIM�<��x}���S�k�q5�nl����"�!�T�w�*��?�A�������a��+��U[��^�Y����]��o'$��d�duQ�4���.ԥ��nE&�v�*=�xV�^�|տA����P+�����X3�Kݒ;�Ȳ��	��Ut��Ί4E��}uW,@�}���bɮ��9RΏ�bH2,KLwN���lC"62����\>��n���4�!���v��GV�r�R#�WCn�q,(��n�OXO]�5�`jd���QN��A�O˖
��h�@�E��i�+��t�����}�v��6,���i���ps����㯦	�eaL���X{�8O`�d�1QT��fޢ��mhĬ��p��釥�R5���B%�e4	�s&�o�w�5�c��P7xM�c �	"L"ՙ�&���0�y �[�Hd
�$����g ��7xZ�[�t�z[��*g�̨�����T��ԛ`Ao��R�q�EW���e���������`�^x=����`����]�Z'����f���v m� {S�;�qO.p=�N�þ@��v�((��$�v�ф�c��$�T�X���Pe�k�C �R$��D�QUu�d D=��om�e�>ͦ>�qx��<�+i�~�^Tl.��EԦf�'2q(�r�`έ�Ƣ(}c҇�*��� �}�u-.�nR0�]:�c�gk����n�o���jǍ>��6��
�ʆ��?�-{*{($}ei\���s�a�+GJ1����Sޔ��q-6�5_�Aw�Ķ��HK�ɢ-��rh�O���nѢV���(!x�r�}�*@(R"s����q�[D�@`1�P������,T���'Q.7S�����C.���S��D��d\���0�ն���N���Y�R����O�$qq��0���\�d��'�Hz�9#���F����n"��p��N,2 6����U>g������a6���#��N[(�6�Wq�G��M/��7x���#E�0)AM���\o(v��|sx`G����ю�Oi��F�>�uSO�~�2�Pn1��ۮ�ķ���S�����S҅v7)��A4:����sW; 1�����{�PvjO�?��D��Ignu�71�Ix{��8�������\���t�Du�%=�.hyn4m�rCT@��0��2�9�=���,FfK.��G�mЈ�w!�ӻP�E�gj�r(���d�Z�0-2V�=���@�]�ϰ���5�/:� �Fw�S�VG?AK#���Cc�^vL�
Iêb:+�M�7kt��+&մmAq�����/�{���)�Q�Gk�tv��\t���u�.��v4"VV��$����:�����t���8z�mB�0jA���3	��DA�H���8;�����L
���:b������6�3�L{�U�b]��Z��	@"㯵2��$ ��躈ha�sؕ�+Q���Fi �2�Ć:�v��|S�6,P�]-я7ĉ� ,�锘Zo��T\�:q�t�� �׵ N\Җ�����{�_��=���������]"�7�K���dL_z�8��V�>�`��Sb*Q����M1���&6��l��8w �\���2���eR�c՗�)��P#��U;zg(_�{�آ˩S���Lb��ɿ�}��(-YW}	0ص�%�f,�����vO$*