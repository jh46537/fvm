��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{Ns�ȭ��+{do�;��F�0�S'X=�2�gП�5~�T�/�y�ZzVQ��a��ФI��y���x�wl� -7���G��A+@�׬M�����rK.�|�[�\^���I���!�-5� �����ƒ3���=JM3�=�(���q�$$��e�4��~8?����
n8�,����t/_���ڈ�s!DZ}U�N�H�a{?3|p���'or�;B!mI�7]$��J��(n����i?�,�h%��_����ӱ[�q0��72����"]`{7%�\��? ط.�wq�Cվ��P�BapJ�.k\������}3L9	?,�SR�n��O�?2�>�`�7h�.�����m2R�4n~Ah��r�?���Yݳ��$�O� �a/}??ǒs~��8���f `|��a40y�	޶C�&h,�7
 �{v�����)�q�ߋR��(�FF`���2ߨ��R#�~_��mj�Q�EU��0��D���4��;��
��Exx����+�}��K��'�R����{U�V��$�`�VRA�?�B�>���D
g���8$~��af_E�Ю��%��GY%¢2��A:�����ȫ��R���gt�n���W�pw���r̃U�iJ�,�l���h��)4�՚�=h�Q����ȈE`"��^�T�:��J�C�<�X�u��.[E�'��E|6�grbx�õj��%����R3\�[Y9�i�|��e����yA��7�itfBO�#Jr޿�@Mu��5[y�9��f�,嬫��"�������.(�Bh��c�e�T�z�������|v�M�g����4�Bߓ�t����CZ1l�B&b)���B����&O7{y�!�\�W��[�~����D�=wd��%^��Wm��I�zlh�qu:R#�7iE�!E�kSzO�^&+��0��wa�[%��ٙuǾ��[1��
$����׌kʩ���f�O���,\������<�֙�xME����32��i��j���GAM X��ƒ#�18J\?���a�Js�^��k�a�2��?��S[������[@w'�l�TX$<�8ic}���3�~�(b�l�!�o�
Jp�x��yt��n�>���\i(���� �h���C��(a������!m�U��_�%�x�Ĉ(`b��w���1���������~�y�b�lԸ�~�9�g��u�2���}��p��k��u��]WI�"A��_���)W����:R���4��K"��Y���y��"��ǳ�"�;�:1mN���D� 7�9a�E��&����,�V�G���a�Wx��(���K 5f���+7�&q.�~�0LC��A�:� �F�XQ�|�Sd�O�$�p#%ڦ���/J]{�:I�m7����ᕩ��3��+m���?�~��-k�? �4a�1�����<͐8O�6�oR�N�0�I�lC|RH4��V$l ?"���<�`z�4'e#oB��ͯ����eZ�c����n{O��n(-K��]:�!2RD$�(8����&�F��"�Pv�6p�Jf�:���h��fэ�
��Fi'�f���������� 'l;�`��\)U��yTh���������A�dXkJ�1L?r<ً�����v=6��C�+�>������eѸ�\7S�c5
/W'�fӅu�qo55�'�*�AڅK�z,�����_3fNI.g.��Y$���Iy���-Q6���<ұ��\X�����vҝ��z�5B��R��]����ߦzA�������$j@kG*Qw�;�,�ݨ�j�k�+�7!q/�dM�k��&1��.�{MVg��hV��h�>���[��R$fI�8���x#���P��L����7�ǈ�a�*z�A�mo� ^�����"b�5b�TwU�Wk%���5be���������R+U�?�8���X$���(5I���p`Hx��Q�<M��n�T��)ZఇZ�;���U#��H�Q���;��/��l~��c���F%��Јc@��l�aW��:��m�z8�E)�:㢤�^�4ڢcmR�x��fN���'`����k�O��I��cM��&��ޝ��zf�ea��6�G5��e�p����в?�)V�d�$Ű�?mB�.�i��q�;�1��O�sË'��~��ENeƯ D���)^ D)ظl���)��V��A����ל3��h���q�!d��Na����e���W*ˬ�tu�j:4b�9&��|S��a���s��GO :�z��J5�7�T��,����C�)����,O��p�?��,����#���ݏr�\-�'�8��)��B.%�m�#�1YC��_k����UCb��qQ���ܱ)6���3�B�(������YԳ
�7v���)Ħg��nZA���v�{��"l5�?��\�C`�d,-6&��|�+ f�5kc��������^{rdjv	w�F�ӡ���d��-]f��|��[����3v*\� ���&��KFG�O�s��56ۦ-ݙ�.砺YcY�ϣ�Ї!d��Y�dv�փ����9��tp' �k(G*�HuU>ǾS:W��A��g���:a�d���yXkϫ՜�Q�XcQ�4A=�>Wk,�&wʮ��_�m���w�|#�!Ȍ��{L�&�%4���E^a�bD�s�	N��;�ʢ�r����K4��.iVu��eK�kl���q�U��F�Ȕwʋdo�v)%�˯q�o�C�l�?�S��[�q؄�g[ֲ(vS)���O TJЂ�8}:��O�?��]����(?ī��AR[ޏՎ