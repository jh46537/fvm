��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8��A��t��
�]W˱�ӆo �I{�C3槏��ff7 8��6���7�Y)`6�-�7,!�=�f�&Q��"�qiK���ﳑ�ɃnT:��J����""ӜJT��Ʌj����uo��]B1��IJ�P+p���Ү�r���~$̬�͇��!��||�XG�@,U���56=�t�we[�Ax��mԧ3C�d�u!�R�9У�X�c�m<>$y��l]�
�tf�?�� ^��fdT<�n���r��s�?��Z*�����)��Y����:�v���c��0�`X���}m�z0\)	�/O��Q�J�rV�SK���&�v�!n!	�!��z|�M�%.�.�\��R���Y�q��CN�`"$�T���9�w{��˙�������m�![�Xxug�i/�~����ʠ���t�s<<��3�54s<���\0ΗT����a��	�ֿp'����su��p+��hN�#l'�I/O��fiUJ��,�����m��l�0�=A��ݐ3���25>pE��S��������nDa�"9	~4���h�K�aS��'�B:\�`���ӝ���C��a8a�,���*��;�26t[ۼOCT�PX"��%{�k۴7*��Mrb����:ghl��Aғ;'�;�"�^$��z;ާ�,OU�bK�H,�߉2.a�N�cls�	y��`�t�g�N]	�� K��Eo���%w#�A�w9�0 �';V��:�[]�ׇ�G*�/�3�~��&_�m��>����
h�Ώ}BDa���x���/㪷\B\ 쨚.�U9����"��mn�Ĥ�������8'���Jm�j�l� ܏�f7*�gH5/�	S��4�b�/��g8���������LG#iq
d>��V�o����}�#�X7�`BE��̝8��j�T�r�қcA�\5	�JG������G��;��ym�1=�P�������GO�0����fs5 �3Λ�~�N�K���`�Y�g����Ć�/��`nH�2/�U����I�Q�pC4?��Wu>��26�ps�+ŭ�P�P�js`����y�����ߊ6-����iL_뎤0V}	Ѻdy���j��7�y�]*��A�ǒB��V�d�5�ݟur�:�!/h.��M:���oK:��E�P-z��BD"�Ϣ���_��ȣ�p���BȾb`c��j� ������o�M��ʰ,�y��}t���M�a�������I�2p�s�4��+5��2+�+���I��k7��������@�^j��/��D���kqdߧ5a��8��T>�Uf*�TR!�������Ǚ�����a\�|��N�U|������g���Xa��8f,X#q{�W)]ݩ���P�ax��֩���.�X8�B�|�Kͩ�t������X��Et��H�!��t���������r�0'�<-%?�̞���5����(RK�!ڿ��U�7��4.�I]��;�u����ed�0Ԕ|b����9m�59{��%�:	�rp+}�4㖦|lc4�k@.<OW�8!K\Ƣ����Bß-{D��釘EM��M������T:��M#Z�j��:��^�	�2�4��k�R &�	��-�瑤�TN��p_t�����L�wP�BP��3�S��!� �*�9�&W_�[��b~kڒ�g[���`��SWZ��$���<
R��u\����-�%b� x�Qt��uZ�f����t�*�սI�������C{�� N~H�d���֫\�a�w��U���4���`5f5$�J����fES�Q�����[	���1����%CZ�`�ѩ��Rc�>o��W��]��ħ�D�-J��>�=��(=�q�|ۙ+�A�F����T����{�~1���0���ӨO������Ș�T�#�f�l�:��V�n͆[eyӸd*�hT��Z;��$$.�
���a�$�#�P%��e{$�u�#�y��>�r~"pXi)ffJ�{Ʉ�3���+��I��W�/H{;%V�����
F�l4�������H}Sϙ,�$�	Ѷ��<~hs�J��X�*�*�X����F�������FLSZ�(��ݚ����۱f׻���6��������q.�q�HK	+���~R�7��t8��`�֘�vv�ʋ:�WY�9�)�!+'m#�9����3�?�R�����N�z톘ꆻ��� ��D4���:�A&O�:�,���ȸ�|r� A^�[����ZV�Ұ�GC��=BXF�j�-F���4V)��C;��7��pA-�|��7ュȌ���R5,�5�Sq�Zؼ�B��	\����z#U�'W,r55j�-4���(���|��-K���[�0O��Cϫl��/����5Yӵ/�l�p�A<�g���\6 ��檥�-�x#�?����#{ytPk�V�h���4�QN�	�d��)���mTmG,���xonmQ|������ީD���R�����w{�7���%������0�)M⚤y�͈��!��"&l���i�匊@6�QV���^ȯ�ӎ]�2�Ջ�Z��0�K)ta9��+�����m08#�fTX��������;^iܩw�˧RO�zCGU�[J���OLp�m�5���y�s0k�IZb"-T�>�I�J}�+������遖a��]�*-�/qySp���ؚ�.�Um�ZR�_<���tl)h;��-n���p�#�)͈�@dPM��q��Ʋl�-�gӌ5�{�@K�-�\�cT�|�����o���h-�k���Tt�T�H�rZ�>�wBe������ː��y��*sBHY{���ZyM �W>;�3Y�m1M���Cy%WzF�����dy3�n�^�$(
'��z�X�6H��D2�U��x�yd��d���ڔ���z�������&�[ |pXi�������M�C�r��K���f�w8��О$�b���μ����Q���I����e#<qA����n�(a��`9g�$Bi���N��,����AuL��v�49�
[��~�����aC6�u��������YԨ�z���"'l����Ʈ�0;��ʧ��Uc0Ϗ�O���Wk��Y�4�)�X�hX��1�H!�|��d�1���C�-�~6?A�[���b�>�� �;|�v3?�r��l������-Q��E_�ȕ���k�Q;��j��O��,w�����^��RA�Z�=�І���Ӽ�H/?��z(#����n���(1�۾�;$bP�4�RQ/�t�����#&�jl�ɫ�Bvܐ͑�L���Ef@���bO��w!C�
c2��ܻFo�=�V<Z���#��mGK��$�;��:y�{p�>����`x�j�� �d��E;.?<g�R��N��X#�X5Wq�:o`#6(�3 뙥=�{|��^ M��� �2(ħ��è�	G�8���4��*i��ɬ�'� K����<��Y���伴�L$%֕v�#�l�Ev�r�^N�Q�i@���x���h&)f���P�	�ɒٙ�ߖ�YMko^:L8]C��	�Q�E>=�>ez����ͻЃ��H+f�~�kլnM]p���������ݛ��[R���b�·A�S��<�������~�Bc��xxgX�Z��v2�)�fے�L���!�5g�1W�����V���h)�r�^q��_ ���͔5���ai̆u��v~`N� ���L�b�3�\x�u7���ӷyD����Ǘ��>h{�@g,M��9��rOGR6R�5����0��M>�d�D�X�[��~��y7�Mim�@z��7U��yBs����N��+�5l)�(��E0����]�%ȫE@&I���<x����QX���C��/��%��f4�����V�i�+�&��c2��-��W�l�I�����a��I2}�>� =�:GbU9/ϙ=)�"�3�b+6tſӁ�ٹ�:��W~�U`�Չ46���-�;���yK�2��N=k�&4��j���?	2W��f.�=�-��d���%�;���� �4�'X�gOy�Ŀ_eA���R|Ģ�������1jS�G�e�V�!!��grz��J��;IQ�+���t�������{%T����0��pŇ<V^6�����ֹ��d'����8�}g�-B\�����z_sqdRu��Tn��d�g�*���=c*���P��H��@W/�' �f��9�o��{��+�����ާ�G�&��0��2\1W�^�z���o^�,�]�s'���0��gq�����P 6Lt���oa~Mp_qn<�`�I�X���
���%��d�5�g��i��=��xj!D�
��J����9�y1�2�8
����$������Hc�4���,��'Cap��n��(��0bS
�7�}R&jh�IB�UO�(A4��G�v¿<9���!�GP�#��l-��,��[>�~KQB��>��z����{T��k� Y"!���5�\AxrY?2=ݏ��/��^�C؂�}:���2H�\��|���i6@���!vKSPf1B�'s���@�_ĵ7,xklf¦��༚*0J&�hUE��Ec�����r/<��S�idUr��-_���45��e�p=����v�^G\���d�XtpЩ���� (8UK�����⻉��G��P��w��Y�2���1��֟"�z�V�9_ף�$^/�����ZЊ��#�($�m�.�\�D1%�;s�A�:mZ�����ȭv�B�_zLP?��$'ޕF��O�`��4�����C��+� ) �rn��v��m�]8NZ���KL`#�B�4'h����;�!�u�D�=�"����G	�덯辂��^��P�C�;�^fE9��Ջ���Ƙ� �y�"��8�E����}�9�#W�ͥ�b�-�SSN�h�W-�w`q��YN�뢜�'�{R��L��>�X�ֺ���h�/��/�%��D�8|����M �Tb�)T����a�SL�l���{���K��˛ш��y~pJ�t��K��d�����;/҇�8g�oZ��)���6	oo�ӐH p���F���A�+���˿	�!C�?�<N��þ�y��D["
a�DXͲWCXV���3�B�>Ҡ�-���Ǔ}��(F$�|�ȐK	yEIǷQnr�ף��j���X�M�K7���O����'��䙛�P`���L���,��]z�A�/cD�Sn�E�>�3��Xs_~��p5��� c����s߹���T�5u̢TEz����,����Få|�䉥'=�+���u�0W^�F��*����P��:�=u6�C�{`<������e�n��������y;O�E;>�׹C�D�oRƇ�ɌU-�����
�m	SC!�zE(B���W5�MŢ�����k��~s�S&� �t�1Ěhܐ��Z�WG��Pb!����w]�G���h�Tb��F��EYi,�F��k�u�d��B�[}��[�u�p�^��V�a�,M�u�M7��%~y.�'�����%D7K7m���!Y�n�<�0)tgG�&.��=��sWv<��P(f���J�),�<\҂�?n0�$�s?j.��mv��~�?m��pʊ�7�y.��|�X�
Q�YX��T����_���x�r��3��]�t��oP���k:\	��Ov�|6~�=ʹ�\�YUȷ��TV>\�Vp�P�_�^�1Z�\c�?�p�DSA*�$O�+��xrz���o��~N��	�s���mfp��S����꬇u1#��SӴ����}"��4ܢ�*�0M� �=Q8�ڗZI�b�@W����E��.�>¾T=U���D+�}�N8����"�W֊�����u�a��AR���t��T9F|��󋾇�MW|�d��l�1�D��"��* ���:ոO�z��>q����{�0�P:J�e(�ة�)_����'��gc���bK��O���ndnZ��I�\ӹD,��a�����ƥ�ZNt��O#���2)?�08	?z���,7*tq���E��p���媁�Oc�B!#x4���́
誉1�	|�s��o��1&,�Ɯĝ��&�41t=(<�a�0����Hګ�?������8&��"? ��|+t9�g*�����)��'��#��a�:C$�ω���#]��V���k�8��M�*j�7�bX6˒~��j��㿤��	XgY�{.G.�9$9�d��V�sv�;�Y5��<�aR�0�Xs��}ͣ��<�$�C+��jʫ�1��4�Cj�[��s�b&ϔj�ӉY�E���yPJ�^����!�$�E�l|b�,�]�Pݸ�vH.�b��2�	"`|��#DNt������ފ	��g^��;�ފ�@���|��|�73�w�f{�&�/7�*���X����r丌����������x[.�O�6��VC��S���+<��wN� �}��#H��p<
�z��85�����T��d/���P������@����q�U��6��FK6�\=@'{���	]�SM�>t��.�o����;E�����},��H�w�X�y{��e
���k֨�`'�|��ҳaY��23r��Hb��t1��a"�~���6c)׻GPL��C?���I*؟_Ӫ�A����j.�#�]�\�e�N�*���HS��Б��IaI�v��9?a`=i$y��o��&�b����n�53w�0���k�M���+�J��c�WOG~ե�ߠPnl%�l?����D�3�>v}��	:���'!WҦ�r����
ҏ�_g��L�Zς;Jį%P#$�t�,��%ɓ]��s�\G�a$�B�E�4����͡��+W�"<}�b����!������~Upc�F�~���[6���dn0��rw��n�'`�T�G��Rh@�|�( ��-����e�>E��Z;+`����п[܇?�T܌�t���dfi�3*�)�-�/Y<�v �(���X���^HBe�K|�dB ۮ��p����f�}}k�m��i�R[Ի�Yg�@uF?x.>�h(nC\�*Ɉ7�k]��`!�B��͗�큨�|}��"sf�4s7��=��f;�����/{yٲ�BRkp>ѹ�1ٽ�hEv����r�`�'����h�qYW�w�ށÅoZKCꯪ/��YP�Ï�K: �u,��n.�=%UI��N�sO�響�Tg͌�P��P�B�����Զ�"�807���ȆW�zg5�z�=hf_n9 �[G�0����7��a�T�S�<:ʼ����q��e�8���4@�Oڤب��O�f?g�q.}�#�)���}�TL����,�*pq���_�ݧ1N�v�Q춷���6&��|�i��F�J2H�ɴ�T�cҠ�~5���V#ѹ��(���h��h:���jw�6�H^1���1�-��/t_�<5�5��˺XTiKJ�ζlg0�+���O,K�f��y�^]��P3A[��+
~��>S7e�ն������W�ܥa����Zw*e��?�dCFI�!����p;0r��G�$��JIw���~��˼'��V^�i,R�kD	T�ѬjL�*r��S�"qM/V�n�@/_��#�tC�#��0�28�ǟ��X�٬cRs��mJi�{�;PW��*���w7��%잗���R�t�,��[����V����B���V�Rp�~G&؟{h�eN�l��b���j'��d"P	���f��b�e�6�O�����#t��F��7A����w8��S_j���o9�L�2��������$t�R��y��c�'��9�,��lW� �a3gX�*bvm8yT�ŦO�K�t����xbBQ�~�����?ʩ��Y�a�y�	Q$g��0����N�~Rz4������豵�	�	E�_�
"��6%�]<��z�&E9��B����Co���e�
���w�^'S�C.AF��D��s�r�Mü%9�`���a�Y�íwQ�-9Z8h���:�Y�r�B�]v9�0�k���8U^C�I!o�f�ME�������Dh7��Oe�T]٪r�I=J�9�fOs�.I��ikL�U�7Y؝�㈌�t�ݰW�5�s���{4�@�U��]�H���N��;��	B� ����%G�EG�@�rTP�YaA���9ԁ~�n����ڭ��IYƫ�gvf�N*RTD]��ڙ6��?S!�?0�><����Gaݸ�ێ<x�-�AZO�v�v��\�!�M�p���X@/Z閷� �����	&J������8���NZμ��E$ ���Jj�r�����v�({�I�Le�h�>�5�L�M�������x^�h�+�Ab�QAhL���^A�GՂ���2�\b-��s���N֑���2���+��l���5�Z)�x;�X[����)�9Ō�w� �4�W	A�JM�WB/HJ�F�����\�b3�M6���/�L� j��⶜�6�����X�z��
\cZXZ�.y*	��=g"�@)ҵ���>�5=��:�R�TC_�7��K���OF���<��/템u���'
!�S�En��/L*
̈́��P��|�6׈��L�"�]��YF����Ró����p,�����lX�w8�[��'3���2W�?&$����-�ϝ]�O�l�4BI��u�NeDIcc�&�<��?�`�R+`b �"M�On�AMA:��#-sX�o�oJ�]��S�2I`|���]]�T�vMK�g\^�_z��W��}ez�Y��<150���e~��1�a'��l�;|A�����B� n$_Æ��Cؒ��Y��"rD�S����2: ����=Z@��-�89[q�$����n�߫>㱫B/~՜�eM#�A�@I0�NGgl���>�����%1Ȃy�w���rԣ.�h���	s(�`��������!����P5��3�W�*c��,�MĽ�Τ�� .U�c�<�����i_� �<{�8���� �QJ�����ʀj��C\i�(���;�&kh�C[:�2�#���b�����/��Y��.�	�s:�(�Hg-��D��J������V�i+�eC,�33L|��Q��|�]�)W��k_ڟC*�ކ󺜴OC ���Y������ֹ����� �:�j��M�2�!e�L!^%�����Ǆ�V3�a��̍�#��qD�"��[>��{���xL,���`1قw��;8O�k<����}O��F�hE�'�S�����:��8'YR'��XH��>��3�����?��QL�4?�2�.iX����;����6���#X�������4��S|���ܛ��ۀ�I��kI�*Cn�Y�]���C�i;	�\�*$�HA��f)�41M�=��D�R�7��1���s�[U,Z�{�QŚ�w)̍���J���|Iv�8���8!��v�6�xQ�@&ȭS�0e����ʵH�Q�-gk+��dl����h�B=8��G�rm9�p�gM�?��r�l���s^/"V��Q=�����A��n>�$Xi�� �	���V[z4v�@�g���Q��ߌJ��>��+H`��	�9\"�O��܊��CW7]�����B`��Wq���!5��I]�ݦ�� ��ʅչ�N�����B+ضl�k���Qr��n��h�S���t�(`#=�j�V�D�M�p�Z{��L�����b�(U��CM�I�n���n�ղ��l��y���̝Ҵ���%���n�`�ӽA��z[N{C%ɱ��4�Q�|˘����h�aN�mo��%]i�S��j1ʏ��I*�*�tcӽ�Y~�ت�v�_�:�`������jf���E���h|����قm\���k�,��;l�T�����ʖ��g�ɜU%j
������J3�2�s��6U�-�tS谖�,Vb��<�Gc{
���ы}�]�=�iR�i�{����7�tѝ��%�iryk�.+Ѝ�'�u-Q��:�I�4��"�FN�5��C���.{�e���/͞�` _���;I��!�/�`A�)]�Z6��%�۸��Y]��'���������-8�׊��u�u��|�[�p�GW�8��%Ώ�i�Kz��#��AAB<�mfCo��.RH͐'1|�Z�p���L%����
?�6�NQl��j�EI���z��<�۫� ktȔ�I�r����4�ê�ʣ	�͡td(�udQS�,�)r�91�;�ti��O���<-��x{k_2 f�9�	P	{3�G濤�(�= 7�c[;C��k��N��5��|U�U�������=�� �h.0��R������lqk5����ܨ��~��u�qv�cɪ�B^ �9I1:���j��M3qlu� ������X�&�[9$��%�f㔩��s}R��;��chy�mp[�|��:a�&�r����y}|;�`�����@�1�?�t�����U`p�WW�޿#�}<q�$&@7]?��^0g?�����w`��!^|�M��7Oc�oΘ���uk����(�6��a&�+|ߑl�EKj�UBU��{t�<����)��ah��2�.ۣ
@$	 �g�p�F۷!��Ka*���js��0*[],�4��:��\�~�X�Q�5.�R���eE<�(���� F4B�q��*P�-�t;�v���\q�m@�G�~[ !�Q�z���n������:�N�{!
�4��M�6���	�z�,I;��]�AR0Ĕ�s��[���t���ИE����cѝ���.�/~���z�h�=���Bz󄃃�w]]�}���]Tr����q�jD?��S1]^fy՚��sݤ�b$X���kM�Rec�������B3_�E��,���1���:���=b3�"�ْ�~KM僘Y�,��f>#5����6�-�=�X��C���<)GE��CU[o�܈Ί��]���9*�Uݱ�S��&�#B�d��.>)�:����&��7�Z�e��2˴���M�x�~e��y��'���E~1���<^�$p����mLϬ�,�~�x��R�����OŐ����3]q�c�
�m��}t(�Y�3L�x<���[�~3o6 ��c3�
kכ`Bq���Z��������e�j��!d_��*���Y,�<���T_��6�/x��tݴ�%[��@n��.��>��MR��R�U�C�V��n��;2D�AO����o��kq
����Z�VDt�����Z^a�� �]:�p?p�Rp�L���"�<=O�C^�!yf���E�|�f��U�0R+;��+�-�a���h�8��nO�'G9�%��1�[�樭�x�D�P�K��Ah�\��G�|�x,��Ą����1�	���u
������b	8|T�mc,��Pk�m}G�b7�9���T�D�����R�����\�.��ǣ�$.O?���;8���D���\�b��zg9�g6���:�rO��� ښ��ߝ����k��'&�z!���4<Q_mE,뗠;���������E�jϒ�B�CУ�"�户ZTS	�����ʼ�i�VQ�G_��y,�"�4+���k�!�%����\n���s�أc"�^�K�i�rr�A�(YV�è�»H��ǣ^ݕ�G�J
���u�eF��>έ�O��������ǖa��%�^��o��B���f�
RO�~1���!>#�����'��-~�Ɓ�L�� �J���0P�DR]��h������Fȹ�~�#6w�KZ���#äu�>&�c+�~S+�m-Z�P�O����eh�i�`���������z��i��X9�z�%�a�]���\֦���荸9��;'7�z����$8�4�^r��Z��q��_�A�\��m��kq�0ۊ��qA�:�&CG)��u�z'}�`�gvэs�
��B<�M����
,�9<����Mz^�I$�~$k�9��E��S�9�`f��
h�bs����"��rŻ3qio����x����Y�HnN,��<c���[L_C�[9�Z��{NR�V:���}
�-~�XB�n�&㭄s�[}$��*v��^پ:�]�c�����#+p7�+�u��zb3
L�0����:R���������&�pg�C���o��������r�P�r�����#z�Dq>�3�f74�\�|���f)D~��>���A���	�w[��I��H2)
2��.�x3��fc��+� s5ҬHJ� �$�v��P����0��0"	�_k�B��� ��T����T_����9�c�f�shC�����6H����kNÊ�j�m>5����pu��� ��M�J_o(JW���v|D;_����J�� #@��������iLyf�����P�{H[�$�q��a��+(g��KȱO�
�M��=qT��D��-��T������!{�5��`�Ԕ�F��|�'��rhKf���ojz3eA����
�}`5�|�/WJٵO�>W��Q����7C޽u�M9�Q�uaJ�T\�p�x���L4�{��S���Ռ�p�ST;?%�{���W��s@�5��4ȀGt��*���x����|�"�6�ݨ5O���	׾ ���a�v���|E���8N���(����
��C	��G�kb�ݟ��Ngs�N����&���>���ff������٧��T-4˨�;ٳ�0�jǨPzd�>,;b����|�b����!���Kg�''�O�OsߒB�£��B�O���z5w��G5gfڤ�B��,F�&���	�8٢�hƫ��u�t�٧�٦7��}$=�9�"�'c��k?�(����s�`�}��μ6�9�^G���Fr�Uӱ�;��1!K_�X#�+)C?�-��+?Y/��J�P*0�bp��M�C�;�^(׀,��ث#��ʪ��PaZ|�m�X:�����cr�ަ��M�3��f����1���Y���`c�[J�A�Z��X8	HjnW�"���Gn�(������_r�b����
{~[hyοnV�Y]�*��WS��xE��V˶Bb8�Y�!�5ǲgs�����1y5�^�?�{Շo���X�J|.ک]�%�Qr�|��:�e.�&mL=}%G�v_h�*Y���.��$�\l2���i�g�(	���JU�t-�O�E�,n-y�b !���x�^�,�3��O����z�i�A33�*��i��Jf�(����-v�#����^h`M"���\���{W�� M��ҍK�{2��cCd�a�L j��4��ذ ��*�(�y����g�h5"سZ�(fUJ�r.>i<:E��_�mA��/b.��,̐?'��潝%G�l����2,���-��ö)�N��UU�Ýe���)��Ü"[�7����o��Ɍ2����U�d���
*B��6b(U2?غ8�\GL���g_|f����n��ã�9��&t�e_d����������FA`/J
q~޸n�#��C/�-h�P件��Kj�<^�/3��+PW� u�#5����@y'W�d�]8u��?��n>p�� ���H���+#X�kA C"�m�%�D$zw�y�
��,�I��oml2'Ϧ��}&�g������:���g�QF�r��|N�^���t�97:�sS��K��FhS嬧6+���*��*	,D1��q�E��z0|i�S�W���vZ�&��E��;('�:��ٷ�4ڿ`!�%��w{�әDY0(�*�u�s��Q9TY��W�h���S@H�.h}!*�:��]A���M����,���Nc�<��	���!��@Ӷ�) ��yՊ���}�b��y�p����Nk�h�.w�@�Y�0D|Έr"�{~�r�x���1�fޏ-�0[J�<m�=.;T�@��Qǹp,*��M�O�`@YH���v�b$I�~I,~��f���0Za'�@	7A����~*���T#L�BB�`@؆uC�go�TʀG
�L#�Y� w��J?�j."�zޑ{�QE�p�qm%���_���cJ%~�if
��+S�]�,�t
�X,g'�:Wf���e���m�r�
�A�y*�[庽K`}��V�83��_{��2T�����d* �צ�4)�U��9U�˵D�i���2<_" ��A���T_�_#,U�Ң� ��]�>o�ܓ	�w@�a�_��F^g�N����z^�ZGsrg���� �+R���s�r��'�gG�y^r�m %��b6B7�x�%��9ϾF�h��ag8h�l^��IM�(z�l���r���l�U��{�|����T�e��7����ݤ���N�սN�ݳ��[0�G���NN_m�N_|�����}z��F{Cӕ<�F�8��Y�gO`���,�yw!�Co����WU�K�\V��x