��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��)Y� �1�c�{�C�9	��܈Y!����lJF/C$d,�V�<�.
Ւ�-!S�h��n����X��ѢS�R#`�ǗG�ݠE^�^HQ�JDbs��:��y��I����@�1��'�1�Б�4۔�K�s�~�Y.3�L���G��6���<\�.�
�m�܇��Q�o�j�>�o���L0��8_����M5ZN阮(貹��.+z�9�Y�]}"t�(&{?���s3�!�ii�ߎ�u�+��S�,�mI�=G�/I� -�Ez���xp�󴽏�i7s�[��9���?�i���m:eT�!��W�T�Ì%P�Y�M7?(�V��ē7�=�@	��$����ֽD�(S٤�����|>
LmC�r}��?]c���r%����D=�����h֎�	)C��k���ˑ�;�,E8��5�'��竣sC������O�X�Ur���s�ە|mÜ1i�>�;W��I�%tő�� 4�YdhV)R�,Xq{g���x��_q��ť�K�D<���U�dMxƯu�&8�C���ʬZ���S>I���F���e�B�8!��C���P
��Ȏ |���W�����g�������h���n�*1���~s�+㈙��Q&:t�$|a�>�%��X��J���p���_��`2j��](�S(t$�(k�����Сt�v�-�}�$���0=a@�ʎQU]3&$z�^�m!]�l	���Hg�JΨ�W�[$��ά� �уg�������_6�L��>��z��
Z�/��E�7W*[N�� \��z9�H�-�k�j�/�O�3l`~�ج���J}�V�s%�"��vέ�Ut`Q@�h�^�sX/wN�)��8{K���US��~D��D߉�����\�c�Bɶ���K�F�Qȩ�=���7ΰ�aI?�|l��1����h�&���kx�@ꌏ�=��S<��xY*�?O�����5���X��}���g}�O��3K��X�0�`2Ae���L�^��y�`>�o��GrZB���X���ɂz5�T�no��Fiʂ�Ĭ�n���H�8��+�6�q�[o�B����Sۇ#��������)8g�0�[J��>�W�Y�	=[�:[$��Q�{ڱ���PA�(�{�[���i
E`�ߞ���k���a�X�z�I�*Yoְ�����]�=��0������'�:�Lu����&�AlfC��V�'0�ꒈ�����]$�G
b�����>�*�-q�P���5���k��[�\��c�7L�vl)=T�-��G�qe@[��*%&+���39���s��L�Х�Kc=��V���7��}�%���������z���W.
�ș��T�8�D����{��6�e��b�?MC�/����u2c�u���-޷����	����A�DqGXr�Q�����G׵L��=ѫ���t���O��e�~ES�~��-���f��1�X�v(�)�p[N#��C�
�N�5�T�q��������GqPu�@�(�R=��e/���d$�bs�)�+&��D]�q}�B���wYe����{j�_�?@�;�uJ��>a)�߯�FcD�M*ya���	S�;�®��w
��O�rs��'6�6�pK�)�N��)��7

���9c��.?��;�t��~э2M'Ա�J?z�ʓ{�l@�Ε�?^��je�ʖ���W��/�&D������q;z�����Pӷ���F�%�����;	�TMD��k�f����$�O�ò{��:��o�Mx��U�����p�q7�2А�I#�#��H}C��_ �⡘|�F{�pFODjP�-[��$l�"tS�տ)���y^~H5��Ή
\Pd���V�J�Lhk �6��b낫���&wZn�|�H[M�҄,���h.-�0g�;*����S�1��jC�#������� �N)f�=���Z�$*(E.�G�����(r���=��@Ō��7sV��w��(��p�CqY#���\�iI7$-��n�f*q�5g"ū>Т��<�P-���yj{�������M�Q��R*ֺ�#�|=	���[�N74���x�d��� HqjpE���<Ob~&�3 7P�G�΍������̞�k�+'o��\�YS��d�g������d`��|�k�f��w��Q����'��(��/xוl�x'\�;�_q����bz��M�'��'�k����2��g�&�ៜckZ�A_1	�f�BH���A+2m�أN����O��i��܏}�kx����M�T�u�[Fq��/���`����R����a`{��`JKipƅ�(�O����F~�׫L��$cQK�~�q�/��RA���9-��̎:H����HG6������@D=�&X�U['�X�Q�L�R����[n�9c�b9��@���C�/�#��a�e�=��%�������1_$ꅹ�N�c��,T��!M��>�B���_��+�T��s�֘��plt�ѭ�+.1�s<j5J|�H��	�P���Hw�6{�y}���o�����6)�Z�¥��E|�-�R�\l��ڡCM���CL��:F�`xxƌ����Bpo��<b4��U����sp�%��E�զ*^���!�)�h��ʱ��ܠɎ{����/�?�sˉө�U��mr�(I-�^
�����4E���L�ňD;B~؜�I�uB`�t5ݠ�T����a@�
;G�q�E����x���1��ű�k��ر�+��E���5�.4���	N��S��b,wk���������҈k1wi��#Ct1�F��ho����ׄ�5�.��0����_֣�Yd���O?�ϋT���E���$.��ᄼ���.��5�Snr��ZY�3��ST=ZT7�h�o����5Ǉ�VkؖR%��	�'< ɫѱLl���`Me��N�]=i��j+��c�X�����L����p.���G����%F[�!��z�:�(����>���؋6 �n�_O�(�������2�_@B��ltȊ��Ȉ����ev��W;񮾌��Bx6q��_2���Ϋl2#��!�5���x!\bA�)O%8Pqm�`�0Qk�=ѢPRo
4e'!��)��F��p�Q�V�Nu�VCdop�y�9��)� M6f�_d]/����+8��F�l#o�=S#��KIiڦ�_�4��a���*nD������B����V��l�`N<��o����c�ҽJ΅�R�]���C\1�ÊI�H��o�Ǚ{�1����YoG��bS��J�կ�~�d�L���g���o<��*g	��.<�^f��8}��=KĒ�����/���+��?&,�C���
{�Iu����W��Qo��\(+2V���y��b����n�~���߬PHסc��@���ʌg�ҵ����,^��s�� -ё��Q0�4 }˅�5Q�(/JǍ������W㇠�k�ÏWs��ӝ��r��H�����G$\D?' 9K9�(�[H���zz�?���7���A�@�|2�J<-Ϡ�&vi�?9.S�w����6�������*�����`�\�Ѽ��_qR���.�T�gH��p�f�A)��X��B�����|-��Wٜcu�(l��:r]5m�gҠ+L�V@�E�>�V�/n	����z���.%$������$��*��n$��9����z�~%e�0�p*���/������x81eM0z���ϳυ�	ʶ�]��<_��Ejo�v�N ���}�9�?/r�F�9V=���9��>:�H���-��7��9�#�z���m�%�1Ά�'`�*fV��R��yI]b���y�Gw>G�)�wQps��,�OG�G-
8�
]CH�'�.g�� ^��iI�Ǒ� :i(�N�:���qt����-?Ό����	�H[�G���m� ��b�R��,U.sʰ@�&^BR�u�[�*�c93�vZx�̊V,�;�@�t�
� ���yF�H ��V�p�����6Zk����IW�����0���ǳT2Kh��.,l�7���IZ��U�o�2a�\1x��S;Sl����e!�דy*6��#��4�Χc��i��c<�Bn<Oh	�-ƿ� 걀-�.6��_�u��>�i���q�|���\�yKSuqiՙϸv�����``����T6�1]������}���]�����<�0��hx�GGct�>��Ç?��*]uO�Ԑ��H� ��0��=H/*���l(���-�c��U�&������@��1��Tò���^�#��-�!��[�<B#LXZv�8e�=�D�'+���7B|�	Gނ&0X�J��~<`sHT^$�hw�AE#��>�O/�Y�A�'��Q�\��`���a�Qc������U�`F�DT(՝Y7�l��l�A]%$R�0����zR�d���6.���}:�Ӟ��Rn��-����fr_�T�H��vG��X'�ߣxab�-���kL��b|L4��^l~��!���,U-��4�7.~�1�P���7�g�Z�|v������j�o��XZ�`/�4�����J���p;���{#S��p�S{0ά�Wc�33&M���4_����4�K�P�^N�(�h=���|dn�� �,h~�E��=��9����B����C����/�h�:ֱ	��4ocg��r�yG}��R;>�Y-4����~�O�t�u�V�GH��3r�}(<��N��C(�H�y�^'�C�z�/�~:?d,�S�B��jvQm���`���dy\1�B��G�����F~E���{���Y,j�w�h��l����- �7>�97�ʛ�;
K�ĵ$�s��ƃ���9iԇ�]B��3���A�u���)oN��L �����	t ,]���,���D@:�{�sѯL�8|}��	M��	c���&-��
��O/��}�,|���_]A=ګ�A!ח�Ʃx� ��~�&���4+�����ϲJ3	�]��r���e%�
�f��n�ل���R�	w��R�� ��{�Y7�c�MѥW0��=G� �L;�s��V��c�	1˖�l�����5[�M�tF�4&_�n�0��*��`4�(r]����g4�8��?���|�b�|RJ~��&ru0iJ`J�P��|�!*ӌ�w���b��m��/�@S���)��
�KR���HGg�ન��9K�2 ��z��u+ظ���,�>�3e�'�Ay)9�f�����+:d㇗�!-��f�.\�J:��̦�� B�gbк9;.XK3-"���W��=:Y���sz�t3�C�3,�]���9��W�{Cu���ze�Uwȡ�L�g�[ a���b��5��V��,�����_�|D}�t⳻k�� �m>�L.`!�#;h?�5̈́u��:�ˊ�R\iz=y�?�X�F+I>�b���m�fr��:oy�^Ո} �?�9c��1�{q�Q=�:��6 �{i���J>?�%F�u0����bu����܎���|[r���6.M�䭮��
����ЬϘ5V����1{#��l���y��u w�Ы����z�o�_}��������	e)�/���Щ����'<�Wռ���npB�ݍ��$A�����S"=���-���P�����j��/z�H��I>���;ݪXCL��M+�-�5�٪&���|�w.��N
�4��]�=X�-(�>
�Q��*;)��n���R�w�C��j ��_�����c��}�qG9jE�����5��{����K^Q���c$�)i��Ƙ�:ɇJF�N��ͧOtgr8�)]!�8Io�~HG���j�m�ػ}�={�U
��i�Sap�N�Y��H
?Ar�����M����*B��:as:�V8?�����-(�03#c�~�oA�*+z��O|mcm��p'D�g�o�	�>�=�aۨ��G�8!�ȳBŋc�6���WY��ue��OyyN5�7.pZE1D�����3�L\ǜ
�	;���g.�������>����S����l��e�y(|}`mH^�c���Ck�ws�	M�|Њrd���J�����k�_�JNd7D�j����]=��4�Ӽz*K��mצA����A�O+v�{��h�A!a�6
/���{-{̺ޗ���,rl:��e�^�)�5�H�B��(t	9��JX���Q�J!�;@����P�7ؑ���NR9�)E��o	��y<�lUd���dsY��ݶ/	��q!	'����S��e�?���/���Ds71���۝\u5���0��[��YDQ`��o:�Te����Z��a��R�q�Gf� ��NVr���1࠷yUj
],,�u{B�RقE�Bʹ�ɩbG|�J5Ƿ/ڵcb�j��]�J�Hֱ��k����nie�ͦ�{�n��G� ���9s��KM�m�e[n�ln�kc�&e!N5�j� '}�oQp�3ċ��6�_��1+Å��������gK,�n`�	��c��(���N��d�k�x���%����Ĥ��&ꨰ<��6�I�?��U���xe���M��O��B�Y�9j�@�-Z�uC��u��l�$�r��/Xҏ�F}���9@��
>���4s��7�+P�C�K3�C�M���u��+��DSF�<��$a�2�T��¹u�J�\ϒ�C˝� �:Jg�c�Yو��|���e%8�
mڟ���ϵ�>1��#ב���5{F��k�U:&ٿV�۪��
��#s~Az�m�X1ݏẟ�>x�]��o���=���X�r���.�#b�bU8��ƪ���)z�ԓ�C�Kyr��Z��?vQtV���-CJ����G��g�
����g�'�jH�g1ꮅ�5zњ`�b��zD|:6y/aս���5K��Wt28u��[�I�_���´�aha�r/��}Ͱ�(�I���I�x(ѝt�7��/u�����7�ʼ-Ȟc9e��>5�e=���ȣ�@�1�����Uj���ے��7��3����7������i�_ċy:(*@f{:�{�d-J�')}�N���{
� ��Nͦ�k٣����zw�䒩�6u��8�5X���2F�X��M׏� ��[�#����'L2�y�����>tFs[�N�g��[�h	��~ʱ	�z�A�%�� \��?��ޗ1��:3��U�IJh��:���da��R�����u	�=W�w�yvz�uֽ�s	~���){)\�/=q�Jf�;UD�v�lT��\][[z�T˖1���v�=��ߪ�7���+���g�������.t�w��z�����B3-P=%�~ڌ���)w?o�\�U7�2ۖ��M�[ =ڌՋ)����=�"���׬��l���]�*�7�`a6뤚�TҺ�dQ������-��[*�V6����s�xV+(1����~OX��N8
[�;5��R L�\b�9sWX���6M�7��,A����z��B@���!�8ny�~�C��Jw-�Z���.4B�Q�����wa�[�l`��L�c�#j؁�t3 �%���-�Z��01�T>��P'д���mP� �͚P�c)�ږ�0k�.=~�_H`e7�P�U5@���Zb�8��P6�5���;�F�$��;l�)��؞k=e����\�2��$lF���E�d��V�k���:)��@Ё���c����zK�pM� 2�
����+�>Ǣt�χ2��F�kL���}�xı
����� E�I��6K���#��W7�>앵Pv�ʗ���?��v`l�\AIakIO_����l "�61�;�ǎ$[�/�Uj�L_�>�X���*�s�3��}�%��'^�=e�:����Q~�p���K�A�s�Y.�"{�֨�q�{D$p4�~�Ц𣮯��.�D.@�s��':��<��r��ܾHUC�nh����X)۱�@@_ݻ�-����8�_B+u,������5�Vh��!�*�z���fW�kC�'���x=�*�eqK�Vۥ���9W���<hzR�/�	�M�����b,joS�6G�VPV���!�> I���\?��e�<��{�h��o�\���<j�^Dz/6���v��U��e�j.@t�+���V�.M��S�#�#���f�'��ۺK٬\[�Q��S1��>��f�uh��B�����K)X��6$��4bL ʬ+����7�y$N��xD���̄N���5��+�t��r�9U��Z�u*�����d��Е��C�?Z��.4�HQ�:O9j�p��R��uФ-��&WQz����9�I=��MBD^��:=p�T�QT9%�����6�OD���l1o�),�훑2Ez�ⴈ�=�g�75��F7c���U8�_	�l��fO�p����^��I�R�lQ��:�;���z�Hh]��cz�Y9�At:wN�B�����Ʃ�ջ^��tp�^�J`�x����ƾd=�d��� #.����U8}L7��[R�<_B�L�Y�[�GH��r�F&ԋ�!~8�ŋ�Ǜ@��S�KfB���P�U��D��K�_P���dmO���c6�\U�-r��7֘��//�W�a��x\F����̮�#,(�D�cD��I�f�d|x��x]�l�G�F�Fz���)E4*���>�m+C�Y���sp���t��*/*O����1[���i�*K�����7����;�n��u�A=yI{~X��(/ݳ\(��u�F����l�Vx�/S��P�ﶘR^��h�{KO���P}{t�����je?H���pV�7��C������c*�d��U��N���F�Z���R%ag�:���퐣��|
	�t5�ώEW������r�Q� �2a5�e��z]R(N�D��s:����쬴��¦s��%�Z���5`�G�1�w�P�𪻰R�Թ��O��QKy�;���1g�������y��j��O�*,��+]σN���Cr��#︞f��K�*.'���<f$U��T��Ҽ�(M���=�\���Q��@�u>�I�����R��`\;DI�5�TS��?�0^�1w?��H��c�����R�%��{B���Uv	�Z��Vp�z��m�$��������/E���͘�=y	.��i�1���߄���fC1J�Q�N�.`��M�Nf�M?Qkm�(2h}>`\��J6_Z�X@��:e��ǁ1n������~c�>�f$��ו�%~�[V�W�_<;�l�/a2��=��K��"AG[A���܍,?"������!��,�6p�V\n���b�o��{�^�E��r���ݒ�ǎ�fW6v)LuJ�L�g����|n�Lf�W�xc,mTs[�������y���Hc���c�!��؇
�������(�\��Jn0��O!ʉRD���@cX
� �7��E�����s6��}������C���h�$A�&l��\�.po�Ŏj�hm�$K���E˃�?AE���W����%�A"��;����ҭ"���uw���F�fS��RYWH�A[�eO{����7��*���beܡfR�[��m�X"��3�`�WAw�-���M��1�H�u�#�z�	�ҌA8Sؕ�[���*�F~j��վ�Eܠ�a.��2><W��a���i�)W�R*�u�R�kf��Ʊ�B#����F��T�4�&ԏ��xѻ)�$e�L�1^�b�$�ЅKf"�G��P�nRV-���Z v/4Z�҅#��V�x��2 �I��yg��fP���\Qq(1�
1*姉/z������e%�s���([���Fs��>e����+�b5�DbyewV��cC��V�'b� ��$?-�F	wI����9C����c��.�Ѱ�9h���<*
�uA�N��S@��7�\�01HY��^0�������T��G��%�.l��/���*�ER23`ت���A�vN�JśC �������U��[�	D��1�\������'��e��1�u����<��+��?��������z �wg�H��bL
e%%�M
t���jm�JK/׼7�d�RXV����Jd��,[ ��� ��6rR��r�}Y��3���M*��  �T}����v�����*�Az��5����+R�S=���8�b%�C����ԏ��% �l�E�}����cu_)��K��Τ�o;+}cc�9��"|��v�%FC���~�`c�Ɋ3��Հ��B�|&�HЪ�K�6�~�5���	���k�gwi����ǓbY�9l^^��3K�j~�i*��pFֽ��h�%F�8GO�>�y��<�Qku�h�:SoIĈ��$k�w�2.;�T~'-�����u��.o�l�X�� 
�?�-Iw�^�/2�2<����u�͒����Z���y
�!�زh�:J�q�j�nc�M�Y�m> *�����|,�,��h��?*#����|��T���V���]�/����f���+�_u@���
�U���Y�y�nD����2-[j������n}g�t7�00z*�0H^{Y;/�w��h���2ȅ�j�A��j��vDN95-xY[+�T1�����!���3�����yH?�,9���J��d��<��8*nL�̌�ޚ���;	S�i��Quhh&�$wb��;�<n-q�h���ՠXZ�h���1�'5�tl�N��vN1�������C]lo��ަυ�!���DR�؏t�����*��s�� �.��͚T�i?�K�f���\Y����ˑ�y������f@����1@7��\x�z{C��P�ƽ�N2��Dn|�HK����Y��<1<"��" RSKN����q�GȮ�����"Eo@Ѕ�_���x@�������CS�T^�X�4l�"!��H���>㹐�{KnBL}aq|�Q�9�d@����=���)&��5���<ly�7�5���!�"=�T<A,��8
h�~�dL �� dWZ&�6�����
Q��SƺL��3(?�)%��2p�{n �z���j=t��c�yqr��&�]م��a�i�)v�ڰ�w$�@�D�p�csy],R�\2���򘯁�z���hT��['�A��G��AP���z��Įj��y�E��.f�J��=�}��ƀ	�ݸ�.8)6�h�������[�L������={������*T��#��2�"-��Z�}�J$W%֋l����[�:ȅ6.гYΆ���x
�=��<>v���L��S!`H��(�~�*�˚
<�J�g��_�3�(V�J��ή�n�0�\��&��t�аS���Pw�6 *z8В.�I�f� A_#ԢU��(�VL�5/7�zzdq��{�7�#�Jw�.�5�>�h��7Eڰ�pAG^�G]�u��?��ܠ���۹�^�l��M��k?jQ̒�I��ٔ�4|C�T,���;)Y��\n�����-�Mс�֝��	Wj���<ZF3Ľ�1Y�$\,�+^>_.����/ȕ�x�[���-��F|��
��\X�����,���!>��v`S�ԡ�2���K��<^��)zP=.k��G*G:�E���c��*c��#����b�Od�x*aG���1'�*%�n�~}p�� �ֺ�̍��J����B6	��O���
H~!�����eX�Cp�C&�74zH#�R��?��6ldBBٙl�<��z���e P�L�P�:*�ڒQ^���M���ӊ�Wk&[Fy�9&'Pt�	4�-���8�A1J�Oy"q�d���s��(���}x��H_u��F�i��zr����٥]w�fʶ{�>����
���#Q����-�ͦR���8��";�h'�ڄD����gV��}�үb�j�y6�~]%r���z�5�V�Xg!��^�o�t�n-�6<8���@w+;�&�b5����@��ݭT��s�kĞ���SrO�"�j��Vp D�ر��!��8�Йc�f8�(��k��$�{��g=�OX}$;1U��趤��4F^��>g���~�����u��B�p�O�/��r�k�#�c������Z���$M�̀(��N9�aEJ�BS6�}?�ɡ��6���S�+h/\t��W$[��<�k����;[UH,�O�����ݯ ̺8��T��p�t<�3n��� �� �LC�ZVU�FBV�,{��j����ӰcWM�Ӽ�ݥ�VJ���G��G���b+��U[vӈ�$�_��ڳV.p��xw��{�|��3�a��r����M�����!wT����UIr�֓���+��lT�z��$�O���?������(f1'�s�qEͪ����a�oy�Y�
�Xb7
s����!6��a�.z�F֍����4�m��OQȹ����EM�c���5�.�$���O�f$DG�.2�đj,���(�hn��Q6�9����r3�������!u8�'i2��~�nƉ����z�����x���o����Y3���=�!*���a$Ŋ,��vT��t�@)�4���P��/خ�)k��}^-�za}��v
���IDaI�F�/��P'�&_ ���6Y���ڋ�粚G�<q�9�E7�����"x+N\���x�^��Ѓ-Ċ!$���|�`���.A0�r��w�_�1�6���CyC�[*�n>�ԕ`Kl5�S��wt�'�fc���I�*3l��.�H��X�J�l���e#M��y d$��.�y�jD�L��o��G$ӹ6�����~3�Z�&�
4� 'A\dOW��c	x������e�RVA�Ĭ���o�j���3�e���ܐesN&2OS��)wK�����|��.������nYYK<�m�d�;+f�ܵ�s�L���s��hǵ��#@�H�zI������BS�>����除PWO
��*�lJ�uoN��2�o���C��#x{@���3�D��`�W�%�O}�<pad���^	.������0f���B.Y�̯���$�)��}��������(��j�5Qx�B)�:��tTi�yQ���C?~s���w���[p�6��e�8��v�q��p�R(f� ���d 
s�O-�H���p��b�4�U����.d�ֵ��x��l��C�/2��}�SN�i�K����[�˾��
����}q	O9�{Õ�N�z�F��_|���-T�V:MH)�Rs�:,����5�6������I\�,�)x|�ٶ�D*�0\rĞz�C���FB<;쇌��OC)��+��	�۰�$����f�N@�w�����մ�wӎ7BC93�cX!O���I�E"�Ư�&S�u9<m��9�m�W���x°��\k
�)����Ji=+�|���-�;6�Ђb���jeQZt!G�3�ߵ�<p����N�-�bf����	����'���2�^.L�c�2���g��9j&���L�9AϪ�KQN_��-za�.�_Onx�ݟ. ����i� �\�=>Ki���d#���&���P�\��7�y9k2Pp�y�.R�X�\����yJ-l���\&A��de\��/9�kͳ��Nng>�{�����P�8���}՝�4B"�"�X-�O���H]ʨ�q�oI��<��^�_�B�{�]H���T��5�W(Ix�BS�#$?��z=*��_���%�vc������ED������|A�����Y5�q*�@2p�^2a[���2��ݢ�"���g4l�~)�c�|qX��Ō(h ܑy-�B�����-/��dyT��X8) m���3����I�suvr��ۮ���QbchU�rߜ�v5�����H9����6��G�3�V���mZp}0�>���6��'�:�
@��ɑM��?Q�V�S�S�CY������59��S;-�ag	Hx�o�~��rl�i��]r�5��_��z����%��Jrk�圾La�&V��ߵ.��1���ga��.6m��_j{p�-ֵ\VG#n[�￮>�G��Hד���ۋ�*x^�4͘,=B����ɲA#�1�7^AI8���13�B�U�3��H���A� ��@:���S�E��*�vh����yx�n�E�]�(
cT7��n���i���D[4}G�#%����{���,��s�aN7z �uǗ6��7B/X+�٫I��Be�s3�4QX2�Qq�{X�k�K�7
<L�@�ѓ<d-�o+h��G��Z�%5� �Qx����L>���ŭd����'������c2:�_�x؃���8�[��(ӓ�M�es���*p��oE����:��,l]�x�����ʏpmh��C��P��0 2ӷ��ҙ�i�K�g5���Bߒ�n��ٜ!8���������l�.�Y`��<�댭Z1�w�c�HPB��
`R�ϑ��/��ʔ~�"��T>�*f���r#�d�`�E,Vɴ����p�,ڴ6�
J�Id��{��Ӳn�O;2E�黭(�|β1�U9T<��@�x�/J����}b�/X�3f
����sm޻�v?_�ע�$�g�m�:Cv���R���s�9�� A�xptƵo+T]W�(!-y�kq�ڑ��`3�q�x`�����,P�����Q����--������C�0Xup�K�t%���/�}�j}��r�������	�HN�a�9*��!e1��U�7ڤݳ+�i���e]���z7�Rf؄Ż�.�&��)T'��%S�2��ϊ[q�#�X<Ο�
�<4p	���'|
C �9�Ք���k���k�7N�c���j�Ǡ��{i��<��<��~`�=�+�R�JOj�c�����5H`��R���O]��Q4l�D������N78���-�Ӻ��sUB;�����y��7����1���м{�o�cю�5���(ȸ �̐&�'f�tof�, y��aR}X��piԄq\���ڤJL7����TL2�0,r�W��F�%^Gm��Eom+��}'H���!���:l��#!�_�j����"+o��7qWK`prݰ�zD��92�M��N�)#	�J�_�����>3@hVy�5�)�X��R�\Σ`f~�=ue�b�r4o���?F���U� <�We��"�&�c!X���ek�;U�a��\	��$�- ]G�Z��-$U����su���z�Jw.���d�	H_;	��D�'g���$�d%!�@
Ab�>�r��@(Nݗ�/<����+�]�/�r�" -&�L��s�[�S
��x�k���i�\��V[M�{�҉|�S��vi춾	�׊���g�+gs�(�U~�#`��<U�!F��.��`W�����EY�c�6��A4�D,�P�q��@&$�Cw��ήC��:^������]�n��w��(D[[�������6!����v������k)w��{���4��u�D��*��~�!؃X�7��/�r��.��;�I��8*�:�X5�3yZ�����%냀RQ�]YӤ��L��O1�t�%�ė���ڠ�}~J'�6Dk\\�a����=Q*��Ec���\$G�!�N���'1�c�
���cV�a��&m�� eaW�$vQ9��~�S�˞�c�KA�EH)}�r_�b�'�T}t05����=K���4��d�+��S�A��&���ݲ_R��n�����+.���Z,�%%变����я�f�������]��װ���j%�z�#n�]pI�`*�����i>-px�w�d>�OP�� z���$x��Hd}qP҇,� �%R,�E�VWS��{S%Od�!W���٫P)�C��C�F��V4��f��]��C/��o�|�.I�n��9�`��1�aY`��Ů/�F�ػzg�(��\�n�E$
F���'�^i��/��������EN���r䴓D*�o�E��O= �� �����X�Rl[���y�>[����XXZktj�{�Ӡ��
�k��ZD��MJR�{��]H�Z�lg�=��z�o{'/'�^݄ˌxJ<"�xyQh���e����;�ݶ����5F���YdB�3��m-C���:=����׹�_0��g�טx�K�9�rS=ǅ[�]���J񿈡/��s���܊Ǚ�F���t��aS \~�~L�/�皜c���%!%+gK/�oF� �3LtVU��6yFNT�x� ��A/�� n�˦��G�A|�!W}�EuP�.H��Z$3(���Ox���JSYc������ A7 oT1�&�A������R4"A`S��3�R��)~�1R5�xiC�x����'���o�Z��K����ud �K �W��K��D������b�kvNI�������[�;T���]���v�ȵ�.����>�n#0�̾x��|Yj��|�H9�l)Ի��H�� &�ަ0��IB�ŹA�#�����+�����|*�4��*i�.1����1��b�~ZLM��g8&V5NG`|ن�6A�iL<�_�(/;]����G�񝼯�Qt�If������2@	�������+���$�{�l���窔�4x|�>/�ë���;�n_�7�j����+1�fڵB{p�0Ś�<��Q�C<=��U�����-�<S��Ü��	�胏ʫ>���J��B9* <j�Ԭ��^ι��r|9�buvX�(f�=N�꥔=#�ݠ�����b�d9�Pߒ1s�S����B:
,�[9tԝ�ͥ���� �G?��?AA��e���nN���gژrZ;E�������A<�쪉d��Ds�6�o��VV4��*.������':>�8z@����F�(L�dB7��u�rg�KIݽ }*	��w�L��UD�U6�ڄ���R�� �0��t�y$:�`�Kv��ut�u�<+"�S�:e��c�JjwM����O�Oz���@�3&Wq����y4S^FK�陏qDz%��Qюm�3�N0_ù/�v��-X]	�5kiߐ �@S:��|���V@A�[ܶ�`����Z���4���
�E�v�#���p�����S�h�l�=Cl4Nfs5Fl��?l�t+"A���tK����)v
l��9r3f,O�JXmjU6_AU�Ƣ��*��W����^�X��)����4<��"�ɓ��˾�Q�x�^�l*ņȋ�71�?b���>���2��R?"�Af�b�����܄R�/i/;�z��������
��1�!8��M�њ1J�Hq_�ޕ��`,��Ѳ"��OV}�aZKb�������Ƴ��@C
��I�����x�8stQ�@Ә���_D����}���ͨ���`�dD�Ĺ;��F������{�f�����CBL����?Wٌ&��8d	W�6���j�^ jɶ[&EwMs�YxQ�~q�?��d�!��l�Q8�Ω>����,�2��+�<ř"a���Y�T�Mh�:�8Yw`D"�?K�1��]�TÔ���o�h��qr����u5�	�S�?üK����PO��{�k�#T��p�
b%QX�	���ʌ *C�$O?������ܜ6��\?��hb��内DEV������j�2
-��<½�Bv�,�
F�ɒ��w�x��K���K�ѽ�h�"<& m{Ȃm��Pm��AIKT'JXσx������X�%X�{T�]\����#ܩw����Z� /iF����^޺�z�.-E{y:)��	�j	g�p�<czm�� ���ŮM���Իo��1\_-�cOf��u���p�`����D�a������S��j��n<q�H]]�����+��C�^����c����o�29F�̃�G��Tdص-x�G�ۣ�}�ݻݜSS��-�&^SC=�[���M����gL�Hf5s���sT��S��<T����J)p
�E�X��h����'/��9D�7t�W��$�wa��^��-�
�
8����-]��ʶ�e�����	Qn�a~ݕ�X�^K4TG�ǹ��z�#�(��������޼��D�D��C֯��#j��va�o���ףO�&�-�'>��I1j�k���O4�c�_oRىn����'���o��y��F6w *	UX$\F��a��wV�o���%=t3�k#�}���y\k@��c(����ڀ�:G��gt�����Ӑc�T��Q\|�z����]ʜ�/� `�l����~|>R��\�@wV�X�[���+��a�.���x�t�j�p,�v~�]+Vt�����FzU�?�c��a\�5�A9\�_ޢ��,ɜ/��h��R���E��}\Ru�(�7v�*�H#��p�[S�f�ld�M�3_ ��DqƲ4���<�4����ð����,��5o�\�h� ��-x2�L�&��k�����n��"A��}Vɹ._�s���AZ��^��Be�V5�T@���F�rc����4;F��/�};��O�)˃��}��*D揩���*L�{�0U�촟�։2lӱ��ź����髽_���,���my�1W�ٳ���hP{*���ǧ]�M�0�P���Dc]�p��7��s���O�B�zs���&f)�;��k��vN�e�o�&����}�*��f��*l,d�O��#�0�=P~�yH껾T����[}�ґ���V-!F�`�hɬ�����K9��2Q�~�iYx����=r �m�@�7�}E Y�Q�(�m�ؾ"]6I��.��Z����2i�*?�b�4R��[�TL�� ��p�A�)%P���F'7 W#��|DS�+v>ռX����S����̚�ʀ�p7��E��E�-�W�e���k�^�	��g��1�Z��p74�����⭮q;��Q�t�ƌ�*MVh�ꗓ� !]6�e���ڂ�!{jq�z�z61�6��҆?6~��kD���gꜺX��HWu��"�. k�=�d �q�nqE���=Z2s���U�"ပ�!�@�B�-���:]�`g�4�L� K�k�6P�[_>������Ԕ.M�QoM�VA6�W��gJϼ�+Ąĝ�]1.�0��!_m��)h��E�>��x���V�`;N�{��X^�X���%I@`�C��C[�O����):�KA~G����'[^Qo��v7�@�EAY(�Z OwUvlu�;"٦�a��0�4s����<�������F)�Z�:�ds�3��h>vBG��� &v��eg""��y25�����=�q�C&B���h��8f�, ^��I���k��a%:�_o���f��)�s�E�ʉ@L��S��=�b�%$�����n��ei T�[�nOq�O\����<F����]Z*Ƒ�=��"`�sO�� &T'����1 �7�X�}/���?�NbA���Xj�A8c*T�_��k���Mژ��l�|��:���I��߼p4�-%/��)��)P�=�
�F�^>(�G*����'�/n�\�#��5_���9T�d�&�p�]���C�^���F~��;�!�j⎊�8�8���5�Ͼ�=4Ģ9/0�w!�K�^��Qg���:�C�C���괍������э	d���e8���'w
&7�A+̱v�`����w/0E��?�<ȅ�wpm�N�3a�	so�H��"�	�Rp�����j��Vr1�l2�'(v�Î�چ	�Z�ȉ9D;h��H�����O.�8�}핏PyJ��p�+a���ξy�C&�ÿU>>U�3�U
z2��e�9:VՅ(1�sl�"��|�� �F�(e�i;Y%��76s��H��g� 	M��Oc.tߕ|!���"l���D�6��K�/*w^��ߍXy�n|�x��ߗ<W�vq|��2}�5A�Q�Qx�����q����4=����͒�ؗ�Q�.y�9q��I&�[�j0 � =��������C$z9=D��r��m%���u��v��Ͻ�4���qPv�~����k��1#��b򫼱J��� �*�k;*uRv�es:<ŌPS��q��?����83�o�TEa���=!_k`���q7Ʋ��c���1gxã��#%V�����}J"�/�R��S۹m�^���b���Lĩ�}_��Bv��+̉���V�	!O��ӹz�ɗ6��E�7[X�D�����$'JbB>�}���n�h�O�Oo�����f�jѴ��g �(��*�x5N3��70',��K��	��.��C�2ZR�@�0��~�I4d\0�oà_A׏XP2�1�ZROJ�U����F�TC�ZB8�K��}z�2-H�Yv�f�YBw8���K����H��z�ş���3�ؾ��.W��pڮ�`�r��T8V���fW.�ze�f�6:T[���dV�~���yx�=�JT���en�'q���*"�0��
"rwyW.��O�@�^R������ڶ�>�;�1�2���O�*������,�Pr �Si�T�Ů��f3
����$R=��o�\�Z�'Q�WS~�h��H&\e�/����d#/�B��G�4q{ۑa����3R� �(�ĲF7����p� ���]���H�v��+�p)�	z �.�������T/-ױ�n�AR�I��h�ږ�l.qLz��<s�g��p��צ����g���c��\L�L��G9/�iZ/G��J�07Ɂ��e �!5�j-'��~�wGiW��(W�|����m�"
i	��^!<��mwR�rN��]�/����h�����!�f�Bx#A���ʰR�ep�L��>��X{�k�P��'�ؼ���=�fD��k���GvAC'����9V�Ɛ��z#�Yjg��0�,0�5~�S�	�54)g�����V�r��X�t|@��|��J�<���Y���w���9{��� J2q ��C�,�
�1gC�j�/��)���7O��Fb����m�]m��$�O���YX���9�r��(�67e�Xkxiг+���h��oA�����i�&v=�
@���Z�@��mW�m��1�xA����*d��
�2��J0��"�Aw�|9V��B�zn��^ep��¢�0��+��	~��ge��H��%�z
���vr��~�������T8Q���^֊��Dң� ���i[��LU?�h>�5�Ϫ�bk�Yne膊X]�	�"[�U�F�+	A�4�;vB� 5/���^�^���a�@�I%B�=��O��YCԟ�g����P%3�W�����_%�+�� �d�X.�$�k�����qڏ��sBK :�!T�<sR����$K�0���ye�e���^~;踮����� �&pW)��/)�����'/�
6���g���y{�@y<�V��~���=�4�����\�b S��Is���te���8�j͹�1�����/��z��S��sX��E�֬���[����3ER7n<m��Nb��P=�I�ق��yЗ��πnv����va��}��$y5�V�忞:$�B�hI�WX��1-q�z��� .L0Ӆ��0���Ɛ�ކ1�%.f�{`��d):��<�CY(t�[mXXT«�)��8 ]����؍	��>�9%�=Ʈ6X�T��� �>��H�8~�Ơ?O�M�4Vv�х�K��if&ӹ"�"������;���c�k��>����(xk�����@���%�+5��C�J�ڂ�m�-�^ސ:\�����>�k�2�EO8A�bΟ]��`�;X��<5U+�g�A��-�yd*>v��(ݾ{��>.��Ǘv�x,�Yi�v�,���o�;��RZh��I�kW�6p(�``dʒ��4S����r�#U�f�Dज��<�ޟ,��&�QH�_4(�0�D��(~7���O6�_I�ݎ(���7�j]$�Nf�r'��D�0�JZv��4D%�#�׮�*�����6��{��k/I�(Ү3o�Ӻ..�(������7�"��� ��j�2��T:Ր}l
w��3�>JY�'G�YLb����y�Qk5_������h��`�˙�@�����i�0WK.&1ԇ��,]B�B�QH2
�<b��[�N&_e 4�ӥÃ!| Q�H�~�3�ڹy�l�!����`�a�|��Ì�Zp�o��,},>��o��������8�9�����V�ʝݹst�o��x��h�b����A�p��^����vX�z�g�-��%7�G�*�z���d	|߮C�$���K�ID���K!7�FA&�t�r�bF���ok�\��|��r�nJ��8�=�r�u#`�(�)����+n�K� �nYCR�vw�U����8+�);�&�\�.f�1J�<�# ��m� ��@c�Mߧ|�Ӆ����u�h�e!Ōs'�"be��jK��SLt6�#�TO�},K����C�@�g[ekS���|�hG�\��؆��\=��ܹD @�X}�E�;-�\G���J@h��5�K�/u�y�����{�f^�g���y�᪐�J�!�cY�A8A��+�g��n��Ŀ��5��h��c^(�7C{ 2��n;9,�=�5x�vkU_]�N�D�cX��f���MR9�m�&
V�
�f�;8nJ���z�)�ڛ�Vi���<lz�ȫ߆PJx��j8�1Sxb��F���y#�<����$��!����Q�(w��1o��A ��LX�Rmi���R������E N���@,�|$�}b-uC'P�)�٬��čԋ��+��t@�F���p�3�����+��?��}�BWT"�mX�H(W'n,J��,�u
��N��d�J��׺�t��fOre��/�O(�"�i|�3k�%���z�/e�s؅��j|�Z���,̟O���c:�ʖr F�����c�K�9ۧ�ԕZe�n5���"�s��֑�&ucm]u�&=I �V�����I-c!����e� �q�YY���h�US�[�^�§�$��]M_���br�v:Lw7.����5o�&�m����*Kǿ�C�
w��x�g%#��7�A�e����iԆGy֡f�U�0�W���H5�e�
}���g+U+~��^�k�>w�H�>��0=w3�FjE�Uo�oA6�|��2�M�$H��VsA�F��ڐ�z¬�����ƌ��X��jT_X�;�w;�����w�����@�޽�P���ag"T�	�υ�HFD�I.���י��TW�L&���	]�b�b��Z���7�4�)�(&����ʳ&;T����dm|ſ� ���)��&}n�M&��%Sv�)�%�ݐF>>�ڳa��Y�9�V?@03fC���`*������� $�r2y}4cV����̲��Yp5&�x
����ך#4
~����������+�r��m��C*
{�T���d�#����`;��$p��$�6��$0���-,��V��j-S�oK
Ց�!�Ϭ�D.�7A �m	֩'Ի�%�|\}����c˷r���M�}KKu�\��kd��~o��i�j�����,Qc�L6�-D�t+���gw%o ��S#��샄,X0�x ��r �5@������=���?|?�~��_sj����y�r����G�t"b���Q�����a ������˳q�R\�.L(��%�q^��lV7m�k��顣�}���G��Z�N����v�7��C
\�<,�!r�/��f�8�ȥj�>�l�3l̺#�_�Q��޸��K�1}�-�����{���K��X8Ӿp�C�D�a�5ߵ)�R)o�w˝.*'�P�㠣���8�U�a���֠�b��/Y�|���¼�K���{n��	
D{�z�ilp���<�-yf�����x��Y���:D���;8�W�Glf��1��=U�z�+|��b��&�g�m��C\ ��'xP��c�NE�T6�\W�F�2Ԓ|PW�\�?qg���Ov��/�d8��d�" +N>���H<>��[����	���������f�Rz^�3I����,-�B�0ʂX���V�6���p;ݱ�Ok<,\�"uT8s+ 왹��d=��
���w��9��v�ݮW��U�\�_-h�6���wFM]��o��0��p���w�h�DF�������S�;��b�^gh�z�U�����_�R\6~��]��o����CO�����\h>�7
`������ݙV�����	��VAhR�-3>]�&��L�${�K>(8��U�s�Jl&��>a��n�X�����k>��?C)��IGEk1�i�����x$�R!�A���|[=�������$!���Rf�]����bƈ�|X�l+,/ڋ�H�w�����0���| �O�=��L�o/H�u
��ԟxT�� ���������M1�I�>����4�1�Ճ���n	?f�?̩���#S�n'?3��I��V��W�"*�=��Y:�) +�{��\^pe��ެYR;��Z�ڪxM�*"bS-l���X�rԇ�����&�D2u�H�I%<�Dk��k
�f<���l��g�rn!]�e} L�b�b6�\���-^@�+�u{���lA[���M}���Y�i�@oi��-����]�1Y�M�"rm��wc�}�^�v? ;t�Y7m���頦>j���;���x�9v]�Ҡ1�aW���И�*���-L��IVy���3�2���㘽��_���I���T��8��o� �2y)�-�����M�b��H�O�B�\�V��p���=���ձ���"��I	�?���r8m>�� �`2v��&�1�����M�5e-8@o@�>X�7��h�D�!i�`r#/q�&�)4��p� ��*���FL��W�a�������3�%Aa�0}�PQn�s�<���$r$�����kw���!�UHI3���T��m�S1���Z����#J�BO�*�wF^C��ڼR#N���<}��ȐNI���D�Do e�v(��*Q,�4�H���1�D��f�髻���EI��!(�Fh2��R�����h����T;�j����K�F��f5�1{zz�9��l�\cؙ��y���g��؍ ��bQ��A���>Z;)�� ���{�#�?0�9��oJ{Lָ��!��EBU�x'�/���tf�#f�M8D]lW���DE��҄L�����ۼ�������G�rT_z����i_^j%�R-�"a���^ƶ0R�?�)Y�~>��cufDR�I1%�5���t��������3��'�ʚ�b`y�W��r�~
h���2�c�-K��m��'�b��	�Z��ۈe�i5� ��H����h�tF���[	�^�T��j���k0���±D mI��ǜ6�Q�	6��f�[�U�HC�:�.��"6䱀���(�W
�qP�Y�C�\C��{����KHsH%��=F7�Xv�g��p;֕��pŧ}^��& j
���SSeUD��y�}�����6}7��-�N~U$�5Α�e-�Wh7�����/���a�3)�y����=��D��4�rp(�����O����&,�%�~4��o�w3���8�>��z�t�*���ں����@l�O�!K�1�Y����A��]u�������~���WM�-'��E!�R�$���B�⬦���A����E>�Q����;��m�/|���a�A�%���V^���]M>B��}!�S��Z�5���u�d�^�%,�g�-�d&��#W��Ê�GO0i�qb]�h4��1�+G�/�U�>�9�QV!M���!�f���@n�l�`�^�F�&r��w�<�ABi'��$;P(��}���,U;�A��lr:m+�H�-��vT>0�z�c�^u�Q��}#:)�PU:T�����8��E�)��	EA��+�u��)�����u+n���/��&���#%���A��Q�,�f��$�g�z����#�RH3$1�{a�6�"��壈�̋�d�[6:z�i}����S@�`Y�q�]}�W2׫;�Ŕ䘁�>zxe������u�0�˘bo�H>�紑�
F��ҝaYN'>��\���z�k��2}G�@�O<Շ?;۷���T��ǈk1��;a�-7*�ɀ�U�7Ck7��G�]�c(*t� M�#W���D�}��+���G��Zh	k�P��C��z̴�f��%�4��ۚ�X|�T���Y�#�bC4��*�%ve�~k�DQ�́����o4P��]a�X�< <&�kt�R��]����vpS��?a��8�"	�'2+��֟yf� ��Ԩ���H@y�H5�"�K<��C��ZW�nB����K����_8?�r�%��
�3����ɘ�Q��)cg�:��ңE�M����J�}�P�O�MK�Wc�������UB��gnޔs��W��f�16H �,��`h�E-�.�̌'(���V�#i���K5�s(��р ��B���e�N�MW���Ntu������Kq]	6����iͿ�#N��'+��R������B��O�<�m��b�59[�M���+��j��b��w!�4�i,v�a>f��tS)���07bj�A�Z�T�j3U�_&�ѷW0�~������4,�\0U��4e$���,��m�
�!+�
��9l�240q]I'1�oZW�%�s!�=�pZ���b��U��ʸ(��8�� �s�P[4t��`K��m�ˇ(��!rW$Z�ma��j@X��'��8���[�ù�����"�{,��%0��.����z�ݎ֌S�!��6�_�!&�w���}B�����=�$��d�JWȭ���A�f:�ǮŸl*��[���L}Gr���o!��i#H�<i���9so�}���n5�^������L1�IU�T^��|��6��ˇun|�����Z�΅N��V3���U$��zº�{�| �M �(�S��A0/��_�s����2@��w��m]�� ��8�
�����y��J۠"����+IZ����]�p1N=veِ�׾|��.�e?@,��&_���WmX�Sp��i(DL��?�p��o�F�l��|�Lx��+t���8\�Uژ-�5�G&����+�Q�墹@� ڶ�.7a�ؙe3�Gk,���{{�Q,���jAeH��G�����e�C�吙�@I��y�i����P���{Q]�$���!]���i�a=ኈqSYGъq6�zU�����w�95��k��vf�����d"/�^���9���.��r�
�i�c|�\�eݯK��E쮫���=�FǺ�+r����ɔ��8�ߦ�v�#���P�7=�P��CV$tӅ�/k����E��v���W��N��1b��V��+�/kM��B/8%'�t�c<ds������j�A�JI-B�o:�e�����cb;��:����+8m�5HX"0�ai0A!��\9/�ko�z��P�F��仾g5��������N>���xy�޹���~j|���k���A��BJӉ�csc 6����t�8���ņP�}��)��	��+e���J����K"&"-� �Q�S�`<��Q��xS3i����8��_��Dz��?�������$Z� �ާ���`O*�?�)zW �#q�w�EXq@��o��m6xx��ҙ%��T�ҿ�4)�������$0\9����L��|����-n��b���z��;�Kߖ��:::7�z7���`������k$�!��?"_:L,���#yD�}��|C�*�Q�z��1F"����G٩� ��+�Q�8�a�!ֿ�ު�1g4���Ӊپ��#��f��� ��A�Ja� ��M����rxI��t�
L)��t�"?���Ui�eΠ��!>F�!�~^�)�h�R��B�; T�1��0�Ր�J�3:��#���2B��]���
�.�i���4?�u�%�^m�~�egl���F�?\V+���q���U�M^ZCݹٜ~��k��9N�n����ѣ��^_��9J���c��������7��c��t��𿧲~�鷼�ꒁ���2��,g�����͡ǪgC~"R��ٟ9��H����M_�H�7�@�b�o��Aa,
���v|�gB�] �l�@��螨*9d�*����ڔ��gsF��ݓ^���&�$6�_~e�|"�<�{�!nEɺ��G��~XP����&�����U�jOȾԥ��X��= IX0}u�j��
�38���PK���[��ɬ�1��u샋�)�y/8�G�G1X�d��fX3�@�P��Pi��a�ā��(��K�/ �^�t�&w #����#���i���lʕ�:woz�����b�N��յM�ۂ��@��b���)�b]ګ{r-=&���GfS�A�O�駶OL���i���N�[N�j�����v�$�T*bR�8���\�I�_����O�&�S��G�_�M��y��l\�{d4�&"pX	U�_�.2#��u~y��o������ -��+7���trP�����VK?�x�s�������lء�����eCǂ��&?ŗ�O�ٍ����|���Q��j�����6#��ُm�8�H0B�vE�`K@������G2�Me!�u���=�GU�7��p�=�p�����U�r��yr���U�)���Y��>6���Z\��)\b]�;��+$������{�͞g�����|�(%���E��@R/��jY?�Rk�� DoY}�G2Yp���Zp''[\���Fa�/*4�.� ]�C��� I�an�� �j��Qnܜ"�#?\=�i§}{�R��g�Mf����O1xy����@4���������,��w��>����5��a#�-W�#�o�B>o���IՃ����#3r�|Q�t0�� &~eL��1,�y}(.���ߒ�Ŕ�V��J�r� �9q0;�6`N#ð���67ዓ9��ۺy<��{:r��Fju�8�A�F �M �Ǥ��]E��˅TR^�-y���ದi�Au�rӪe�0MW�� ��a�U�Sn��z�s�]�I�3V�#�yb>ۚ��d�{g�ҷ�B:�B[����L��o5�T��1ޥ�\�B�)���]%|^a����_�"�W�b���P��~;b%I������8�{0���C�Sa�3�U���M&	\kK(�C���FP#�f������W�U���Ұ�:pgb<�A�����i?��qF3)�T�<�y�8A���_�!�pJ�nǻ�[�:9!D&r�l��Pa1tZB��c��3PlI���bx�FIn���`�_���n��xWHu��mw��#�gp16�.(�w���#��0W�I*#
����~m</�,@����y�J�U�T0Aw��Z #]���Vac��aM��!�NU��a���{0[����zs��Z�6��D�W��
A�>z����i�qb��\[e�F1�m7���1�V���̊^�xqq�p���#;ڞRM	��[д���M��]�d��%*�C���R�}aT�Vٍ5k�a�����R02��`Z�А�Ef{_w����L
����_��Ƕ�:V;���W���R��8��i�=^��`"�8�NND1�56V�Y�+U�B`���?G�	�o9�пЂϽ��(c���ʓ�Į�Gx�0ӥ���QԼ�$��!,�z�ɯ�U��Pv<���9�suPe�����/a� %sXRb`�=��\oyfڄ�Q����~�YVn������?�F���6 !}�{i��,{�	w��R�<mw�v��^��
�X=�%�hp|]���@U��T����Df�Z#^>��sF�I�\�=!���j�z���PaY�~�^�P�jؚ�cO_��c�O]M�<1h(�����I�f����2 �R��,�$Ǥ�O\Cd�,�6��׳�WD'9�;�����K<q1�vD!�(DN��p��s!������z��]�QV���c��B	�)+'�֢�D�{p#!�xK�_�`����0�����'x�@����>Ww�hǎ4d�����irX
o/���@�� �_|�Fh�qY����p��r��C|2�Dݧ	3~�����zX ľ��\�sN�~JG�~���mR����}*�C���۾���B�.����㄃s���ґc�IO���9��aP�ƙdH�X�B�3Y��Z�Hr�ޚJ�K�*�D�g�S��"WK���}�s�0��Ֆ���'ά�F��r�����B[�Z�K�>$��Y�U��3�p�ݾ޻��p��z����^&;Z���j~n�X���0S�2��� 9Pp�x:�T�\���/�5�>��Ӭ���V��^m��;�ԛb��-ID�����,M;�=�I�Aa+�J��j�a�j�5Ŏ�[�D�}���:�߻a�C�݈J������kQ��j��d8�.K&\uT��h���u����Qw'�̸�6�t�Rͻ�P�
%ݿ:;G�]-���+�����H���ϛH�� �֍����Ĉ�她���A��kÈ2�v届y�y����>ʫ��?	M�I�g���Y��$s��~�@*[V���iv��պN�a
v��CjB��!�@TI��u	��]�G��= �Tl���p���/魯x��	�B�ɗ�I��l��E����-KU#b�"(^ 6�J0Pn��^pS~��A��LZ�g�1=R��9�����9>�c�� ��7�G�-Օ����u��?�AIM��F�3��Kf��Z-I3�s>�9}%Ǝ�����m�؍1�ۛ�61S=�?�C�����N<�8pF����W#���9q�d&�·"���1Bd�x*��^��q囬�6�T�\FQ�Y��h*3nC� '
P��R�o�r,s�m�����C�ɲ#�� � �קdWm?�v����ӏ�dq[���j/�of�sг��r�!�?)��vF��kH�\}N��ļH�:��y;AҐ8���I>�|էC�5��I�a�В�h�3�	�;�k2��*��c\|���F�H<�)�R/JAB ���� '�"R˪���,��1&��"L4�l���Q�3�زW�'��f��#T��	y�+M����Ylaҿt+�8P�G0��B^�8��<ŰM�{+�VK
�Mq:zb��h:�'-d��`��8�?J'���(�#�o9#��
?	��V}bW�|�JD���8�0։m:����8~ ^xiP��]�;�3o�q�M��@ْ�p��O'tP�z�i�r4���o1px,_]4Z oÓ����^�K�f�r��K@�.���m��<g:K�nDv� �L��
>�����Χ�����E�(^9=�?>uܙ��%7�Y�Z���쟼5���،Z?��܌/�<F%QL�K�.��J���xތ+p�y<Q��ja���B�=��>�tl��F��Z��'[eޘ�tL��$�����C�����bêP���z̜U�~��p%��T9h���z����X�����ddl�%*��E�Q.�	�q1���ʬg%�Lu�����i_j���^�t&0�\�k�U>Ւ�S� �U�l������b���[lϤ�/ܪ'>Z�	��HS(W pcʙ|j�]Ŀ�$޷����\vfB���<u<��ŔJb��Ax,PX�鐧Ů䤇���A�sm��&��G6�M��J�E-ʕ�Y4�*�}6���Sm#֯i6"l������R~^�V�s�m)=��g��Mx�m���nA�n�)׃�1k���3 ����^@��w��`~w<��ٱ�$aj�ѧU$H0��X�T*W�lЬ���.�}�u���:�G3����p��-NvCJ!��E�vz�s­��XO�w��ʚ�HV��Y�w�o� �����բ+�E�8�Ԉ��0I��9(RX$��*c�����m�Ziƥ�&��.~�Ը�?R[-dlF7bK�RȐ�N���������B����yct#��l��7��V%��K��R�H��v���F�j��?��R���ģ��BA+N�S�r��������0�>��x�}�!4Ø�7�=��,�\$����jA#9�4�@��MD�8q4��^�@���F���<[�sɆ#>PX#�w7Y��}��-�����|D�oaTF�vV���� ��i���bg c|����yU�ˎ0�}s�6���e�����L��>�%P��_ٓ��ǩ�6���DWx�6����N!H.�މ��	
�U◱B-�yn���{�B��j>L0��ؒZW����2�vo�:[��F�c�S��~�0x��о�E�&����ϡ0�C��頃{�K�S�/-�ɋ<���FWJ�d0�yO">^���Pߗ�)P�ԧ�b�?��n������v�o���.Eܪ��4�R4��r�=�7!������f�E�Uf:F��,v6 ���Bj�|�WH����Q҃���'�"
#�g.��.�.�3�����H�n�0e���P�|@8c�/��p��x�r�:ɭ��Pf��9YK��BR�~�s�Xa��#��m�=�HN��+���$h"߿�ܝ�R�5�Z���"iAɤ���D3�nUsVY��F��Ŷ~�kZ�df��VhQ��;{���Py�pd������Y2�v^�I*2ĖO�f�"w���JD��J��H�����S�t�ʃ`��N�X����m����݉6�]��t��*8����6�n�`(�Į�'� ���<���/�D�&�cȻ T���G��6�۫����M����p<%������.�A�W����׾��>�m3K�}�a1�KȭW�Ş|�پ�FR&�&S����!�]���5�R�t� [����/)�j����ǹ�M��(���5h~ӂlD�����+�����J1T�2:�>� ��
�;�{����3�u�7�#vo|���ġâSW�CWmF>q�Ƴǜ���^Kk7�����?�=2�@>R	�"�x�U��s3���Q��Sض��/+1@6x��1���$	�e(��ѱyߐ�M�Z�Sh�E�W����Ő}z�럳5�è�$���gI�6Pݞ���>�u��̑+u�r7Oc�f�Ýs]ϰs���`Ů#䍕�L�;�>�^aE��� �iI>��@�މ�R�����3
�s�e q����j�{��W?�fod�jO���c%����j�L�?_���m	�)ؤK��_��<E�U��pyӜN*is�x&���Q��H�%2xrQsSc#Ei��~E���0TY�D0V����	B2�}��$F\�E��
��Z����H���p���vf�ۢ�����X�"��r�0�V�����B+B#�O"-�����lC�͑�}j�[	~�D��Fk�"�s��׬���-`ӫ�%����/mP������P�gX@�v�'��`t�We���]�٢�F)A?+씏d,)щ�8� -�F��4���U��:�|5WxH+��L�#Ɗ�zMCT����\�/���btտ�6�6|��T/dH�m����5]1�;��lҀԀһ�v�.3amq���������������,����` ���E�|O*=��"^�.x��4�7{������i�h��6�~?�Hj�q���[\���6���}p����kz%¡
������%4��\�ŀqk�`���bG��"�Tr_�r? ߙL^�Dƈh����'h�?`��A�U�tK�[e�� ]��H���Q`��%�������z�������'����f҅g���|�i��n�b�D$��GQN�o��qo}��1�*]2aZ�qD�@���X�˱�)��De��|oZ��\��L*--D��O�����M�
_��p��0��\�~��k���1�7S�/���[EA�̋�y3(�~��4�#�L��o�m��N 1�tIÎ`Ū�r�� ���@t_i���rҥ���z��:���S�]�00��sz��=��W+I���]6kw���"�e営GVƊ�>�e�y2��U)����R���Bc�b�$,-1 ��0mǵ+�)�IK�O�!��;��H�ЁXX����w�p���:��l2��~�Fl6�P̡���ƙZ��B8˾�ER�=��{s������:�������Y=�����Db˟��V�=^rA?>�Ŗ��Ö��+�uRPoK߼5hR(
ſ�LV��B_�}��(�1��>�w�D�k�@�,�dU���Y~ga�㙟���a:D�r#�yOU���㱠��S0�`����T����KBۡ
5X�s�m4<�=7�����@�dʷ����9zYmoȡ��jf���4wm�������'��#7���P��X�
q?��}˪LBc=�<���N�:�$��G�f����޵ N>�`���'��j qX���ԏ�%�Y��0
�ΏX[�0���D�"#)����M�������R8��[�܇���2S�b�5|���5VR��kr��x��^_�[]z%'Zpb?U��Yj��>�X�,�8���(�UR��2�0�>!s�d8:l���������t>."A4�=�d�Ŕ&�\���&dS�bCegh�g�۹j�M��sm͔\<)��EE�D�;T�9;��#����鵞��2h �����X����{�����ԋt�Q4�j��N��.�0����:�4!��*�9ȠF3v���W�υ\`�o�礞������TW�޼b �lœ%?ؔ��3�ޟS���&�C�/C���$��ĨjцP��a���G�$�r��Jn�˜0Az�5���f�n�J��}���j�K;o5'0�k�@$P=�6
��+�q������N##��.���� H~�Ǻ;
�ѭ/�����yK"��j���X�r�}>=��)h!�m{#!N��u��G��KQ��»	ezk�[	x,V���u�C�9k��:>�D3��3�ŗ�:��>j�V���,�X>�7V�֢
ʖ�8�[��h5�[�����,���;�0(|��^�`MT��%lxiF{2�y�|a7�KH$��n��*������`$����orY��˲��`M�.��}���~j�H��j���!�$u���2:i��'%_�	O"��V�B��w����} l�q4«Uӛ��	�4���o *8�~�7���Gf�ؗv<;2�n���3\SQ�E=0���W�D��>d���Z�$��m���=��C)�D���v����`����Xi8�P��g#,r���������o�C�CR!���4�(��:�Z��A[7N&�{��=r���wY���U.~c$�k`h {:��jB�X;Z\���{6�7W�/c~vmX���2���m���'����Nn4OH-�  ~��W{����E�g�D?���Z�ׇ�5�Y�v�y����[5�n/"7z��U���
����F�w*�}K�zc�*���%�M���?d� ��b�@�r&��Ӕ�W׹v|�VF�D�-v0�@�N�4�Ή�ob���U����]�4գ�&hn�!�A[l¡������F�k�����r{TGJ�#u�Ba9fP�6!�˰1k��9H���`��Y�P�sKS�쾦��Bl�]>�WK�f%��A��0�������^m�$uCQrJ��[��b�!Jb�s<ͅ���H�>�8����˟����"{(,{=}�' ��>�ؚTN��m/�&��qhX���:�%*}���������Ղ�7���3�%Ew��_�#0],�~��[H��7]X�INA�$a':�OI�Y�?J��"
Ph%3���c!��g�
=Ȗ����K�/�a��R��6�"�ߴ�@I|���!�gNz;����q�5��Aڐ$�aX�O`QJ��9#���$,�2���D#���]�S��a�n�)`A�G���{q��PΞW����%��t�uא��-����⬻
�j���hj��)���]��6[�$2�Vh��ʄ�����t������%:�B���o1t�=�J�� 7g��g�^��}s�>O��F�܉���q:#Qږ%Z?�V�� =*�۞a�s�@��T��i�>�`�B.�s��aLoV��DbwR��'__><�ǜ�Al>5�
�+G}a����[Y�e)_R I�]d��8��$�X6i�"Ϡ�w\�0F�u��H$����Y��0��V; �s�0�����Z�\�XoÎɾ�Cυb�P��Z�A��1��Y�#Pl]��[�1��}E��%Β��ê)D�������:1��7϶��2vɗ��u��V��N*�4�?}@��$))���]��pTV���'����!F�����=V��r����!y j�hp�b�Ajma��Q��,�z&�݅z{N�Y
���	з��B�^Z��/��#kJ-lh��v>����䝠L u�Y��AV�1p�Ǚ�S��*F�6d
[����B}����I��<]16���	�ecZ�س!
}U��w��&F7B)���"1;�RG;5�Q��R���fX��=�,�d�#���e���\�y2_�K��R�����#��̠��*��W41�����D��ҵo0O�AZ����$T��+r���i��V�{J<U��5M�e���3���b�4C?�2��F�b[A����>�(g1�F����s��j�P_%�B�1�9"^+��u$r�Hz]��oG.R0a���tJ5�������tY�V�&��Fxi��/�E�d7�.�:�#��w|$���g�!Ő"��x��uez�t���4�(�)Q�eK�&��G������Iʓ�{R���V��8�tYn@��
���b�d�vh�j��1�\��M-!	D�A-I?��c�X�9�%��v�L ��B4 )�+Ⅹ#���f�6��O �]��#=l�c)y�Ԑ�x�'�\�UZ�5밪���'�Ea��Dy긟Tܥx���]n�Ԝ�~������F��;l�IE�@�:�8	
��`o)���Cs�f2{By�v7�@/���_�<m5��CB���8���_ɜϮ�ɋ2��"�w�'�ӕ���lxғ��?A�����0I7��$O�dS����]v��l��E買���MU�ۡgv(�P�6h�՜�Z��G����>�p
b
*����m��]QoVY?����qkc�.�3ʗ.n8t�"v����ul&����z�FY����*d����� �j��lb��e}{JT�&/(��lV�#~;l���յu���D_��;��]�iV�qPp>EQ��p�X��X��a�Q�vr�f��.i���J_�ϲ��d�LI�U�Q�t.FrH�ցU�c�ނϡʠ�����Rq��g�'���֞з���&��P�ّ�N��*�^�>C����sb�j�)��'Z�Zٗޡ���Rnc��9 f8�˽�
�sP�~��`dZh����/Gîɞ����d�ǭ�G�<}8����R� hv�N*)���C΁��)�F-�0.��o���Q]��Z�4*���H�D�e�#����؃r�&J`=ns킥�~�t�w*me���p�hJ#����jv
���C�L�>2�+x�K�$v�s�1��ڿ�𢾎KR��fol#���lj�.HܼF|�����T�KI U�Z�v[u�)���a�s�޶�7VKS������΄�N�gG�a��;�q����<X�Q�N46��ЇA��D��'��0�/%�Ƃ�5m�j�py,�l) i��g��YX/w�r�=���?I:�J�td]֜y[r�֣�beV���{�Ƨ�pZ��3( R���,8.���It����Q�؁�'A��g���t��\�<�Y-ԏ��~�*����8A��\�\bG�P��,%,��s��Ϭ��K-�^���!�5nç��NN�}���9}�L<�3�3K�����@��T*��us�IG&�:�0�Uo,+`[�n>K�=n,��W7[-���m��ìDs���q1|n�;����7�xa�5E]�	��ț�v��95�9{$��W�&4���AYH�"o*�}�r�M~����y�S�����1����Rg/�
r1Xنp�zӚ l�;�"���듪��kh���v8A�[�ޞ�>X��H'�:�c��rp�5�bDL��p����[�p� J�$�ϙ�e�Dh�͸T�'n$��N�rJeG1E��ߤO������Pɶ��.�^�.	q��h	d�mn~tw�����=��(IV����(�����]�@�o��8B�Ya��$�^Ǳ��b"���f;tY��̈ğ=0
����!$f3#�'�ɣ��H�g]�ܳ�`��,HK�i�J��/�Vώ=�tZ�:<�����]�s�z}���e��%r����Աva�.>�NR�<ɪ+��K�c}��g�X��kq'����j_M�̌�A-�Y8�N4e���-�a�i�=��&w�Ε��&�7aN)��L�.U�?3>�^��|�6G��eZ�Gę���Y`lJ����Ԍ�B���^�6�����`ᅰ��Y������y�]�K~M�M{U�7͊�0`Gz�q���nL'n���W��܀�s����kʮ���1au����f�BnN\�A\ĉ5q��r/ԿL�.��.оB����{�1(��>�?*\��3:4+�γ+O-��'���s��aB��}�+4�֛�ʱ4��؁�T;j�A�g�㠎=�cm��V�q���5pu�u0���;���4���i/�8r���6@tr�0��#�Cmꘋѩ�I�+���>�3M/n�+K.��@^|�ty;�$Ϣ�\�9�e�wq/�E��{���osSP!WB��.�7�̒# ��LT^񺅚K��݆� ��l�78����s{�,XFtu�I����l�h���u��7=g�/iL��{g�]>.��������&g��'8��#���U_�w��T�9/tbVf�(P���$��~soa��Ni��l�}j�
���!���v��ͣΊ���8�����#���;�Ɏ��j��쳉b���3�ӕ��Bd�q��ԈRϼe�����Ȫ��_ִ��|��m��&�_���@�DGw����
�!��)c���= ���o]b�o!�z�&