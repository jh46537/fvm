// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:43:30 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MYc2ajmQidRdklzEP6tkKA7YG0H6rhv8GlVwRS7B0BETQTCjoaGiH6ZsbREzPP1/
b4j1GjOYZZ3xutQ1ocYskGSqBm5JBwy3fr6IlaQ9rBHuksxVQ+PgMgR+KmkFI+ky
uT9+p2414dsIqjzn5EFLyidKP7y3qxb7cXcirH30xzo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3056)
RLNLs+dTToZGwmqWfX+eaQRFFvPqYqUV+yi9K1X+iWnkRjUA/EyG/+mY69gXYHlN
BiSlvTWS+sCNlg/eoq7T4PAOXK9B/VZH8qkHx8ACjydxJK2lC08vn1tWonr5XtFb
ZVRyihpjs/3plR2xkGHZudYYNpomsxEIZQhhsHMvsZGOufX9U5D1LqpeTOBhXajq
JfRXLVYk8t1u7Ygvn2dk3lAQfslPo0teHqwtOGsIM57Vw1iEawlj+eAB5/1Sm5lE
AHgHegvhKdBOzjQ4b6pBpojbAh1dKljf0aJNMApPzQZLmRrKBCEN4E/rm82ghgGZ
p8jfgO4Y6LHxFz+BIkxEbxc2Ay9JB9V7GU0L21Ff9dLmQtETbgCkAdvR+1TeKbGQ
PFSeVvVNn3D4a1RSDZHpUspcqSZ37asLtYlplhtbZ/4d2+7LIVt3dudurJLM3acp
E18f089cMqrKfpBJCl3TpZT61T81rN/by2KBAEqqDVK0TOQrn8uNxv4pnTCaWYow
2AuduqHCNmx09KV1N9w1Mwn3sISvWYjyuE7AxgCxp0qtHkGFbYKtZbr7pAW+XMmQ
/pYH8fqsILJXmhO7P9r2Em8msQGM/rmKtDh3auNviOMiRdriJG4DGY0rwzYwUXPd
ylUQFKaXtm/fwJThB+kKkTfe3iExG8MTmRplK+g1ScoZV4SZ1wpeonNulyf6MA6j
1f6ViDmlv5OF0uotD3WrFi7WAOJeQM+D7xiFQrcX8Mdwn5M8LxRA3CsNCu8H6t0I
zM+NrT0Tb/8guTC+6CSIKQGhse/NZl33K25uUGP1r1Q/Ffrgdel8J96xTc+Sw8PH
HwrMHBkELdpIlGjcsN1R0otUXi87DkmoAaMd0VshEXO3jpgG8OgY+jADeFM9juAr
Vb9m6wHVLmncjkpDkCt4ihWIHHz+4+8YME+lyWAdp/u+LMQyrAScG8WonaZ9Qu3U
7JZ8aVzoIplNWZHq7F+/ibaJARpi2S1qs2HKLuctgOnVnSs5v+kDnGMEzDGnidCz
4iqYjSDbhUFei5cfSE9PXcqgSu2bpQNZ7bjljw75/nDaujUHbopQTavYV2dBvGdI
hUK2twGBV1gIR7iM17qVpK2nVIzBGJ02Jg0M005qUTtGDRTjyQwWcg4+LC+dYacj
kw6YzZfsyWJ/wtQo04MsU46+TCQV2JkFCHIwnzQCCnsnu6x71RwAHvwUTo1ieiq3
x+P80l4im/2r7VSjLJL4r48CH9nP5CnC16cHhzl2Dv1KnmR5h9iR6s5KYdVH10zD
ozkx15Gn5fKPiV4UaEWAgfWFFhEoZ+shy059v02H3MQ91Q6ORAXfvtWmKLY7tt50
ESvWeB237ENugvfeHSOG46e5dTQbG2CCcblv8GDWyhlleCWOZVx6qRP8GmGrTG6u
t5RjrRdou6Vf8n9kVsy5fih0p+fVgKCVn6agm+0RtY6or66P3iql9M3xV6hVEVcP
lYaQxP9Igcb3aBeVxk7GXtHu9uYxefgCbhkIAL2fgoWNbEPOVBMmX+BXH/6qvZYN
zPyNVRB9chbpsLrR+zmQfRyaiZF/AACX+MHqcmEWh+AWl7cqAhNBz4TUsCS7GANt
t/IcTk7xj7DieU1yN2D2El7orDYJ9KBzlgvFuFRzOLHHxwlm/ppQcDTbnSmptvuS
X1Xam6eWosbXYViWHaSLtSE1VoTCrIt6r7VNTGbCdzf24EEZCVNwxrQmUCVC83sQ
AcLwFeT8T8Rv+V7xWI7CBF8WtypDXCWZctNMK0cqLousRLk/OCO2NPe4Dddrz5vV
jcnUAri353pjKQko/fYnkkL1bPjHYkd34EmzXJEePm4Hn8uiTiVjqUbTkPeYHGTv
+ySxAFrq0A92PFEdjiC+3yZ1rRyOCbz9iutz4UhrnXlnBf0Rg7Wy7GBWcG2uiPnt
A4hj+l4qZGsNJTMP/MPstwaVgEyb013joU/C+KkPXqzzy6M+8O/VvlNHiXwHkAui
QJNqBnRS59huqC9jw1eoUsUeKhSdcdx3tKvns5+bckxHpwqwEzQyXvrI8iLhEcq4
6t8XW/dafLggBkMA1UhFzQQsE7J5qv89Y4dBJ2Mvvv5kJONedVWWM84/eSRZ2cni
2AVfR3LIz/XVFs3seYnqfx3dnas9jgcFsBlLa+H+O15YaPlPYBrYsNhQv86iA5vQ
fO9CY8sjNBi77bv4yXHaoGjVA5s//9WgE85APFq69pA1O69r4NMpqFi0avmz/fmo
5x0QLJ/pCmwpa8m5lRWst7ehuouwAwYXDLrF6WWN432Zyj0GUgbH/JEKHt1uzrPU
ag0tCCrBFVcuveNGQ7vBHntmFocUssEd3ZdSquZkXZGNv2CGh/rDkouDFz4DZxGK
g7vE3HJn8CVHcQTskbwOfEvPECH0InJbnlrUpLKI1TkKRCPUjwkoTm9aYAc8jYBG
IkBz1caZTQt8u4Bwh53qFLhjJg2GXJB1Rddnvbr3MPC+GAf0NvbwMaXx/oZ/2MS4
o60zqQIr5YXdXHJ++hcxfjYpja6M9ejcExRj7j/gMYKO7v0nfm/lijiK5kpagJW+
Md2ERiOMB4XKvEu1Fil5UhI+BB/6KOVNpKteOBuukkGNpS01eVkHAjWL2IV4IlUQ
jUPjjUM7hDEbAKlPcWZNbCfgowHOmgrjqfw0w75a2xwXip0eaPXftL5pOVvoCj/8
73xnIlj/UryT/cVOw6mKIOXhTL2JMryCE/76mC/yXS143ynhwXFgyT2H+5d9IQHS
rogLt+6l+MlxImx7M86udQs8B6D07UOLXw+tpW6TDwYUx4dveMjCss6JhDoyisyb
y6hG8mBt+pHK5uRPIpKrz34hRX7dycEVEirPKhCFIrfWYl0+U8sqOuSo4h3Zo9Zt
/lt9odtz1R736nkYqzU9Q6UYWZBkskFsCr/pEpHDWi/vAXf50JGXed2ZvHaTsX3m
++F5uWxfcE6IdkNYTrc7Iu3+y4oNCAi2WwzGFnDE6As5GieDN/Ci/GuJjcyMqpEJ
Pnroy02LYXHP0mzJYBsgHVOUbQcPjJ9MOzK0PBoeoToo3Z3ktp7ZJ5vXbj5hK9m3
/3p+pb3q/V0V4uq8VnyEv/yzta9YSV4cGrzFrMYSanz/JlnwJ7n5F0En+FvFYha6
J4RS5M83iK/zSjFr49Oh+Gws/dOp7dwuW7rlYclcYRJb3r3a511fGrAEB6dUaxU2
WQwLKIMzYT6mXZ2rlEYAnYCdD/iVXO2RyLUdECKc+qYmWqXKvJpbE+22AXwkv+S/
troThD2NeZUUPWgi8XCT01k2JqSb0Nf0eZvkQuYwYdMT5FXpeqipz7LfAzmMVRUw
j7E9Ab8m/eza0r3hC+M1sIBWJzMi8mS8WsDArhVNQSrYXcL5NZfvrTjLCsqFNpxl
mu4xnZeloblvB/V590aLymvFGmrE/0lCc9hyX0Ijc6kNCPCWLuNKEgWbErmIGebs
OKne5UKy8KNxYuaSTpFpwt8EUG+QUygVnDdy4lnbsYFl0cA4peWjFdsPoahQ8gdS
9HJ1ryRMUWD4Er1S2n3tqHVX0GL7l4eXzjyNKN/9SqZx/64V3prc6eiSdUuLeDmg
l1Hqic5KDDpTMeWOiPeXbcGvPmI78WCdRXek8+goaFVCxYM/3Gnc0/eOdDK11lcq
U6pcSWJjBhuGRrXLBd6gVi9HLnta2r36btHjqjni9BR+L0Bkg69SvTEzrnipje46
ePFSzrEkmkeFkxX6ZmjmNAdJDY7t51L7KTqIRep17qpGawAt88PifztYBYDBba99
lKs1uJ1zVJP9wXacAncbBdI+K+mpk5aKubiDx4N3OSb7TT53x3wtLbc+fn77oxnw
8WBaQ2w4FfMCMZ84N/AXL/Yj81t5nPlNBwfH9gwKDKMkjcnLEbzHUD6LVZsMDS91
6EVahNy2GqXaCTRIOgI9eOYUeya9UaRCUJ/kH3NLe8xxlISge/dosy8Uz0z8k0Oc
orGfgisfin8fBB8w3tOKkWyu0xhj+rY6pDThzu0VYd0aV6tWtu3Thr5VRWqkfNF1
M/H+m5fNlN8hQAdU94Ulv3hH0nUgd3l2/yX5VU8Dg2Q=
`pragma protect end_protected
