��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(|����	t!�2IbL186PA�`�n/5_db�����~�DϨE��v�R��4`˵}�<*B,��ye�ɵ[��X�O�R̽��p^��b���#��{{1��HX��?ų$���=��wO	��eUMs��Ҥ_��_�c	:���<<���O����v�M���h�'j]���8ǖ�2t�H�=U��� ���'��k�(�%aG�V��:����@���D��@�(񽒦�a��mu���Re �+������5]�9d�ʻ�M
�c�����]�F��U�
ЃT�{`�*����܁�?��©L�N�1��D����8���R{�H�2Tک��
IqYJV�a/�P��O6HnPY���q��q?% �fO��-
�����S-� y"����σNM����-ܲ������$�C˽�L�ɥ�p*/W(&�]��Q�a�Y|5�0u��Nw2g�Z�W����
�5��"���is 0��pf�Z.�,���M�oy���@��	�l#�[�U.���;��T��Q�ݭ{�Y��8k��~�!��/D%��H},w�&H�2}�Ή���-OC����q������8�ߐ�yd�9�>�K0**
��P�i�Rb��g��20Ԣ��Z2�":Nqcǫ	U�3U�=��~�4�c���jj	�ﵧ�Kix�j=���x,��H�к	?��\с�ԭ��*h�d6���t�xE�X��� �G��a\[)����?�06��&`�栱��hxc-��-�<�f���K���`���B�r����/������:�ǰ�Q��gpS���\صY�(Qkc�� fޑ�>6�!1H�C�1;�E���I���ACU���l�<s�|y�ka��0���uo�⽴��V�9��Br�����CcY���ESw��"Xy��7V73��3���m�5�b�[��o�B�,!��K׭>��f�xL�(�!�p��7���HD��<���M{�ԅ6��	�`^i��zk��3슉zһ�1O��չ^��̄0��
;̻`�h��sȜA�Qd^f8y��c��6�s٢�����2����闃l�P꽆vW����᫸`�,���s�O������Mm3���4�ZH�
C�ԟ.O��Q�e�z�:~Y��'v����]ߢ�Zvx|��L9dk/ོ�vvbr�ڜ���rJ�7l��Զ����Z�@n�yN�0g���C�+�yQhL06l�����ݼW�����<;J;L��}*�k=��fA�]O��?r��n�՟�J n�Zt�W��y�Kk91�ќ���n�]��'`縱���m��DB�:���?_���N���g��r�d]���J�<����7���Ir��А�{�A/� �i���ʹ��O�Ga�5P����ҧ���6ͮV��� ,Re�pO��c��V�����ޚ���t�U��Ͳ�\�o"u䃓}F��=VB�`Lg��@guf�bT�m�JZY�J:�8�U�$�a���=Q�n7)[d��s�P�0�jy���@䪛�؛����-@r�`�.h�aE$ïׂ��?�!NRA��+#�Uns��7Mu�Q#��d�	�B��7�cM0� 3^��y���Ƨrm�J��Xr�v8�B���8/�G��D�@��^��xC�����I0)ZM�����JG��������9���Y�Ӓ�
B�Q�g�v��麩�����W���W=H=]�%�y��"J��Hڿ^
$yK���3�Ͱ�4(�_��^-;���)ٙ�lS�J��%���9�=�Yt��"�PY�6��X��c��up��weo<�ٱ��aӵ�rT_a���%,���BiMفW�xN�y!��7�S����U��\�6�4�m�w׾�NS8g[j�J�\�J���B E��^�2�K�� W'�~ڡ�P�i�r�
��~yD����T_��������Մ�D�Tq���N�����u��ԉ�*c�L ő�|�n��
��,ȗ`���_���w�.�%e0�"����gǦԍ�T��[��/����,�0���nu+�D�4��.Ӷ�wK�*bq��7��,�C�n�C��@/�p���I���KXW�dFI�	�︜��4Ed��zQ	-��s}k�9�]�\Xܕ�n�W/0�>~�(��#�l2PK���姨mx�6�?W�Q\L��X�0]Ȭ�(6.����G���Sh1��n���c�˓���GJ����g� p�D����N0ưz��!T�r�\�ms�q\�M�P�]�Ի	�9�5bq�@P�b@O7�� �S�!����Q��J�5V��ۻ"X5�k�o5Ѣ�S��y� .l��Q�U��^���j��mo�n�"��h��$�+�M��aM��w��ļ2������o�4N�C&\�]����A���*�kgz��|3�9nKv��VJ*��;���Na�\��i����Q��"��}=O o�r��D:+R99a�����VT��q~}���_���S���=��)֯e�[�wR�����^��N���@{eN,��:6������}X���O����� �ɹ����
���m���r�)�Wԫ���_�F��@��xJU��א˜�}���m�f}�R|<,��@^)]hg&�@-���A�	�r�n�"ݤr�qm��5v��s�����-UE+a�|�E->���u��g�&�V)�Ίi��'���r�����A�L������V�jb%�QB1ur%��/��I{�&v����tI�k
J-wBr��j8ӗ�i���䡎��%Ș�dZ� :C���:6�Y��/�1��S�G�{3ϟќ�Z���
?�+�Q�e-�i��hz�ܹU�Bֆ�ɶO�c~mF�A�cK&�=#Hvx�đJًx�	9�r߉�]+�M�:�8t�B��<�P�*R���>�����^�-q|��ʷ`�����o'��o:�`v�E���=Xlz5oӤ��l���ֲ�ќH��x�PΛ?Be�"��ISڑ<L)<��:�~5�� ���]lU:�)�^��v�-�h!�L�庾�7I7@i��i�D�^.��!�z��|�7�a���e�����EOiVC2�4�(��1y�׽�V�
\;����6�j(�6F>�!pY�MV��Vp����"5��c�K�".Po�����sx��H��<�2�ۭ�.�\���V�v��ꅦ���]�V�9��0���@P�/ε�V� 0���/�h0p��wY.��2-�'AK��x��'q�6��^ 0K*P��hȻ�ܨ�"�07A��q�Z$XH��$��"c|��2uq�v�\����;�o$�I���n͸ L�C�� ]����M����6ư�G��hzy����#~��\R9�d�͔�#�� �;1�����|\}����Y�
�{�>��7�i��(�����]LO<�(q���m��U����Ƿk����bJJֺ����A{��&���,�{8"��s1$�B�Dm��?���rFyIWB�m_.�Dy(�(軮�K�0�%lVR���,j����\LԀ�{�#+b��y'�z�ދ/���5 Bqa�~��!�m1�����t�����r�;�Px�n����!�p���0��"u%aq�����Ѥ�󝆤$x���l���*��=^�	?Ή:3�\:л͙=4fp�{��R��P�f�]@L�{��F���6����0�g2�(��Zyik�ڤ�\��)�~�5�0�S8�,�_Ψ��T��G��L�W<4�֭ug�0��o'�ֲ`�����E}�#=�dCW�r컇{�_�m
����yJG��^QV��G��BR,Z��-hy�|�(*'Ԝ�����7IC
4�������˞�c�u@��$ҵ� Y{6D;ߚ�l�Q����B��Gd.����~��������)���wa �
�Z`�z���r��.?��L9�b�ݙ\?��ڨy,�n�p�ϵ���1h�L���D��5�:=C���� �D���ԢԣG�k�A�g�r�#�����x�ö�2�p���ą���Q��cC�_iN���Q!#�pO�Q�BZ���X�)���f~0T����я��~i�ŚЯ�$ޚ��iδ��� ���?g��U���i�K����r4���Ҫ0������	L�~��������
��-�Ғˑd:����t�|@� �0�n�h��Ă�x�W�v��znB���;c�ZӦ�Ǒ��#1�<i"�4XA�2Cs�w�r�������X�~r���n�v@������p�f�<�a{�f�,��>3�5��1����jU`v��!��=I���w��o���#5����h2⒥"m��c�Uy,�3f�q��]��b*6�}�[��6��<��S���F�x��~��>�s�L�Cݯ��4u��������ڪjP�xAԔ�2c��A<��qE�G��v5�������Dض�o.���B[�DXZ�J{Nv��<cSY�i�Q�I����ODZ��	�2h�Z��B�����v����:\?y�'��%�v�
%�^уg2$��r.Z��q;�j�V-^"��d��";�`m9�ݶ�`m#� ��>Q�Z��H�#R������v��-΍�sy��S�S��cN�T?O5�?mA�=B�M�<���4����o����lcBL�X�GT������=2@A�v���C�P��+�c:
�ۡ"y&�����W]PC��F�Q�N1I-+L	K+o����ǽ����8�T�{x��D$�!PɽF��0����H������ݠ�����V23���ų_��[��
6�:�c�4ݹ���[+<��>���8G����*뫄~V���Q
I$���v�c)K)�G�j�;��Ϩh/H�=��f��C_n9��P�y�C��"e܍U��k�����8>!T�����W��b��L��jH�M��ݒ��Y���dw?X�����[Ml��b�?W�^�+��&_��H�� ���K�RX�ƕ���XY�9��=*��Ň�/�7`r�+�9��-˕v;#p��90����d��
���~�(�Ϭ�-R�f��M%� �驈[�$�ި�)�[�O�>�]��j��>�¾�	Pգ�;yY�e�mݼ�L���ZD�J5!�ߊ�޶Y����?���#_^�K�:�0��*�pe�����C�fƏ��]�JXp��9Ǡ
�~o�med����G�w��UG��	��.V�c����o���2��(_�������W��6�k�;�Pp���>l��S�i�)���!%����&�+�����]��H�嗨WvQR�[Zi5_TM�uR&Ԍ�w��H����'Q�D&�1�q>+O���_�R�XN��}��u�CX�����y l,߿�&|� �����0��f��p��򙎊�At��>��h	�1�*БV!��!�cy�:8��%�:~�C�(�C�4��R�x��kc�ѝbΏ��1�ׇI�K���~֥,u�B(�@�~ե���P6y��c>�o�ɖ�,�����[��6��˳qC��ߴ(��@�>�ƣ`�[F����&�4��K�K �~bKg_���soY��^p��ʀH|����܍��-���ge><n�`߈s�q�*��s���E��y "�`�e ���D��%:sPP�3MHf�&G�x�C(,��9�h��IͰ_��7v��w��u҄D�&S�8�� �����mUr�5z�P���y���e�Ni!�-��R� V�d������DK�	a&����bC���-�B�Ak�������	����'��������h$_�ݽ d�8I睻��D׹i�R���1k��0Q�rsEi����}~�9�4deAυ��0�e؊�E���[ Z�g�bƃ�2�Oc"A��v3:b�/н�$��w�*jx��8+�[gd;g���86/�JH3�ugk2��&�}g$��K���|_��e?�.k�O���s�'YZ�w�5 �=�� �	���W�V��Q۳-X��ܛ$�3Db ��G�)��&��|W�]�t���$=*�l���w��C���=�,B[#��B�W7B� ��[K�������o�<,B!�C>4�J�ί�e��zu�����f�XʽQB�\C�C��L���3����/M'�4=B�����O	+�h����bAbK�����d>]��Q_�ʋ�Z=�h뤮D2�|@G�)���v	�7����,YH\�?�#�7"e�!�z܁�.��w4&��;�Zi?/��0<חF����B|F|���)��WR�����A]}�,�5�#�N?Oմ����������,0�X���d�\ԛ����Xd�|ϗ��q�Y��9�v�ěU�欄g���0"��k8��FK��-�A�K����<��y^�����l�`W��	���P����K�tֲ�������h����`ӭ� �/'i�֧����͟geP���[��[${�T��ˮRؽ��DG�LZ?�+��cg�;��[��V�f���X���I��_o��ҁ\�1.�啛�xAP{oK�!C�Ponq��d1o�0�oy袗�y�<�f��0E��yԐ��x&-E�ej���w�v
�u�B�_T�,��	u8�	���l2�p.�EL}Mv+��f� �d�R����*$��*K�؃�wUK���2��	�j?���E����໳sr��Q3�\��'�|���������8��FJBӪ� ��ˤL��WM���N4_�h��2�[��6��|�Gʻ����*�@��F��+�E�h�����I����ZI�)�t%0�ԠJ�f� =�
3�!�qR+ZZ%����n�/�:�a��Y�����t�齼��RJ�q�S��.��:n��3D�Ԅ&)�*_#�^� ���'Ȥ��J4�th7F���#���:z�"�q�3奖~���5I[Xh����}�M��eD�퀘P�p(�;�Ɍ���@�F@�W�n���0XE�¥[G$�?1���`{�&$0��#����"�w��'j
k�9���}�͜�ą�D1�_����/ޏ�~�+�z �K�ύbp����#Zf�반��QjRO*SDhgT�+@�i�KZ3j��]���zg�ed5�xm�`xkPɝ�2��wmYǒH5�+#�}�Q��hk����U�K����5��H�ct�?ɜ$���iDxq���M�K�눭Z3:��i}_+��<f�g�*|�v��ey]蹨�~k���myX|���:�h4����ns4�@8|T�����Ta$	���2��_-�Ҷc<�y���g�w�a��œ�'X:�u�[�I��h��$��9+)6��Fi��g+PC!��*I(p��%>N�/�hNڿ�q&��6D`1��:�v�)�ᔖ�i�I�d��⚸���z�.��,N��Ҵ�y�5&D$oe�hۨ�J/�B�\4AX�;h����R�� �
\�X��pz�������.!p��)UG�1Nl��n�<HZz�I��gA??�Y�#?��U)���*�,��n�7�,�g��;�4��<ǲ��י`���a�~I=��� ҿ�YsGt[`ߖ\ߴ������s�n��=��LB`}3ҋ6�&�	c �_Z�-�\��7_P0�M�Țrŧ�����L��*B���q2�|m��]���.�3�{�k���z���p��Jl��r�"�8�6�+{v�)CLXDk�BG�.-[y|��/�w��;����Sd��f&o�Rp�Zk��c!�B&#�ǜL��/v���w���jTh�g��]7���g�Q(�e���$+��L�K�C�qX����%]����$��R�f��x-.C�G%���V�RhGKt��Dz�Վ���_U�گ+H�?��̀ơiMc����
Mb(Hn9GO:7J���kS���(3��X2��j�>�d	��ʵ�wkS\���ԩ�gBx7�A����y[R�O�0zj�[~��T3hS�����E&bq�`��A%�,0h��E˺'΀܃����(�N�coOq#A֕�e-��i�́��En&d���A]���x��u+����dvZ
_�m���%�=�X�g�*u��������
)�Ca�P�PZ���0��^n<7���շ��;Ü��x_lOk��t�6��]T�#]�� ��$�v��z�t�]�tE��D#�0�oς6<�:��#�ŔD4!���\��p������pW��ڞj[�㕦��c!L��w0ʵ�xo�,��o��@����ު	�nӅ�r�:�Q��E��v5���S#c���tU�г&���6���L���C<���EP�xi��D���o�������&����!���μ��\Qa�����!=�H44Y���w��>�3�I�rF�#���]w���D���OI�\��jDH�Ym<n���<^��6,yS����8�6������Ǣ��A󙾓��}J[�ʨ�t�ܫ~�G&z4&2�y���)�	��]u\RgRa���c�VRַ}�gf��7Ʋ>!ޥ�\%n�!��_X�����y�P�eꓧ������^zų�:ōPm� ������P�S��<L�E��3ņl��<�e=<W�$���܍�A�稁�u:�!�Osb����H��V&@�nF��P�O�?����񂙬$�����|!�?��D�S]�]�ڲ�BB����L�����~�~^�J:h�.��R�pdJE<PM�����#Ѡ���^���mC�P<z`�L���!�e��]�wL6��`�����n���4}&��&e���Ʒl�h/��X��������B���}
]@��5m!�V��,;,�x�W���RT c��0[�J7�N��C�r�E*w��g\�
���墷$��as�j�/ �=>"����i��ۗ9=bOY���)����P1��On�2�3!����D�T�f���HJII*O͋sgm���k��^�@��W��?��$�Z��qV�j3j�� z��^Q�;3�|wM�gPg\�Q�	����G�9�"E�P'�D<r�2�����U\�ַ�OIϷ=T�́q�C�^d��hA��"���r��x���n�ի+X�Uä{B���z|WW�G�����1��="�2������ [�=	\�#c��E	�[��`2����1Pޭ&<fL;d�ᵌ��l���;��J*Ʃ0���Q��c[�XȨt��KK��,��D��UF�m,o�܉�+��1�L�r���j�)	? '����G��j�u�X��f�]�!k��9�xg��J�����p�S�����:(��{ S��;zn ��ܙ���Q���f�d���y��q�ú�8Å��BB��	^�nr~�!){X1���\�g+�'K"�)� �a�uA+�Qm�3�6oN�F����+&6uX�+��D������"�������H�L����O^���KXm��=&��7�y�
u�x�Ү��K'͞�-�]q��a�/�C*��]��4�jQ��T٪�Ԋ8�Cmm��!��ַ���e���Y8�9�z~�WGy~r@����cW��΅��[O�����	}�o�'Y[T�9�Bך�|���T�<9����0D*9�a�K͎�R�U�3���'��70�34}��УO�*�[/��u�t�wv��iY![����w_e���8L�|Ř�7��i?��J��!�8i�o%U���~�!d��ëA��%,��0/!�k/��8�;1� ��6�BZtE��|��@���1�@܍5�h�;�����Gb��3eܶ8�[~�*��&ޤ��u	2:$Y��!�������-*��`�6H��Ņ�B����O����HD	t6�T%�r�棣�er^�}��O���� �%��]�֜�~���T.�pֿ�C���`֘�7o�k�Y�7�
����:��x����4{��"�*�V��Ϭ=�7x-k���u��	o��q�zO�>OL��&��^�$l��װ�20Q���C�!0kx��b�Y�s�P�����1�[s- L|v�a�b��)~1��h^�m2�B�P�*���"@���r�W�n)ni���o��C9�P^�. �$Na�ee�/���z�(�0�*�����/��x+ 8Quu�z��%=�dR�+�}�ȯMH�e��(��8x�V2c�s6*=db�ܩE�Ѭ�	<��TT�`]�����o!�^χZ�Kr��X~���P<�R윤�e�5-��{M�	�8�o��T��g�ǥ*�٥���8�B��ִ�ֳȮ�o�;�W�n�|dv��yv��7�^�l]�ف�#P.YB�����f���Mda�y�ǡ[W�9�7�fw*�-�F�Hg3T��lxs�g�(bM�(�ڪn�KQ�+��m�$�ЌY�Ęp�	�15��t/�(��,���p���,$�I��d��]��i���ʾre��4�!h�䖏m����i* F�|$ܥ�j���
�*����4�E��~���U��eJ�~s��4B�O�h�ԪQ>WMB�3�A�� ۻ.�mY� &��z�\0�o����8�ڏ$��򘉌����|dhu��ZU��������q+ ��.�4��>�o�u>��t*�i� �2�J�g���(�0���o�����`�,�N�{��c�0r�}97FcR��o�=Ń��H�"�+�*w���2��ii}y �T&�Oo�W���\Hc|�� ;�6t-9�/i*���c��1\N�����wn#M��::m]��lv����oEO��}A��-U�&,ݶSһн�vM�t���G���4��E�X*"�`���MLFwH���TsU*��8	V��r�$;��� �w��x�UtF��7 �~�o����5L?HK�T֎����衢Q-dȄ�@�ܾ�ebU9���0��!K����6Cr#�?��d����,�'�7K���;��A��w݌��⒛_'mvJ!���ǫrZ5��oׇ�
y�M��8)�mg�'��������X�Gj@�����7��[��ȗ7�Ўd5[�o
��4.��v��,y��H 0���z�`�	O���-�gk����M�l��Җ�X?�����_\�H�4V>�w�i�C��DW�T�c�F�Wp#��Z��A	��XZ��F.�S)w#�b@L�;<�'��ŭ��Ar�H�TV�f�}Ø�X`�0w$��,�X�.��WBw��Iջ�4�?50�d��Zk����	'�(�筆�ӿ�Իe�3�`0aW)�������Ӧ�.�T�)�0lbA:��Wwu�mqȌ;������ݡ{�\�=�?�ȁ� ��ؚM��d�	�Ҽ�1�j�Q��v@6~
	��ĆƗ��K}#�8��Ft�{=/��	ש_����v���#|e��ھ2D���"�5�\�c�7�����	:-�̣����<���!0ݚ�@�; F����f4���FTq���S�r�e)ts0ă����-wP��E�y���h���C�~I�Uv[��,�r����_-��8�Öus����2ao �t�X�<jV�Z�%�g��d%�-)>�y��r�Bnd�+"�	K�6im>t��\�N�����Ty����mQ �9Rj�T��Sk���}�Ɲ<(��k@�i=����]p�.DiQ��r���SL��\X�K�љ�EA�J���_S������W��%ln$|7���a�
�p8:�({L@�FD��h��'>���k6Â�_b[�[�B�ȫ��������F?_T��ò
i2�O0=��U桸�F�/ߒ��%I:�K��"�խ��T�%>���(7���6h76��҇A��7�>0��ut��U�V���q�8�S��g}F`��><���<�?X����|�����KP�M	�~'��o.ҿ�У�rV��OƳ�[z��pjt͗�8F�-�2b_6�:`a�F��`�t�4j��#���)��Ρ��*ۑ4{�	끆����!a�m����꽞�'���Sx�`�x�Լ�� ��G��6��Tլ�U�JK>B�->�2UDy��i��e�d��r��R\�
�"4v_	d�ы�2���+}��S+E�Hɹ�np֗%���:� Qו���Q��(��$�9��Ƒc�V�
�'j+:PM4�$h�Y�g��U.�Da��g�ګu�gӨr
���Zܮ	,�˫����� /���t�{�Jr�4��oi�$��wԂ���Z�7UU��IRvSY�VҪ�n�ί�߾[������ ��:�;�ɨP���{1�)�w�AOCe��tOA��ЇKk��F�֯�	j[����-`JL�A��3�4�HT����lcC��M]SUI�Aݞ�#�� �h��v�9��`�1���K`w�[�w�J$_CWS~a���~*.hBw�/<x�G�SL��$�c���id�y�)F�=o���!�^y�,���A���u��������#�y|�g�h�|��8'ҵ�)���%-�l��~{xz��wAbFo󲱊�Z#�a=��KFʆ�3�
��H!?Ux�A��Ϛ���D������t���ln���&��uNÄ́9��`��sw�'R�p���t�	�ǰ3UU�w8�5δ�?I��R}����@������(��L/_�6�,M��*����F����L���J!TȔ�B��jg����N�@��Y��'�\�*�F$hI	UZ�.���^%C�x��'g���Q�|й[f}���}$cZ3F��:A��N��=x��I�ڨ|Hr�^v��|북�5�d�*b�e+��II��i�i��8��E�f����T�jnZ=V,ɡ#�����!9����#]V����>��HK�s�@K�?��2Z	���z$Yt=Ua����-cy&d��\ʋ6O�뭈R�)_h<���1r�3U���JQB�.��]�P��d�ߩ�ڇ�~��H�W��*��"��,�\ ��@ɰ�`E�� hbS ��BȄ}�P{����e�,�G�{|��J��!�R) �ھ�0��^�j~�4�S�a�<aX�{��c��-��4( �Ԍg=A��5�Dl�ߢ1�X�~�lܟ���O�ޜr���s��*�Ƣ�K�2>p=�6/U	a��B˙ �{��PS�I�as@��!(V&��x���7��1t 5SMm� ��vv
�z)!�������!���|ޣs J�f�NMVD$-�Q�O�G֫�	v��i�-��UL��{�'���T��(��qn|I��
	1bMrW⇣�}d�Ϡ_DB��Y6��5�ޛ�fA$Ab��E*���s~т*?�{�������u�� `]�ϲ`Caկ�\/�7�YI�����=�����nSc�N伂�!2>O��Gp	�8&���Y;�у�dv�Y�#���0�L����qGY�����u��L�K��6��=�W$��yu��������*uE,�Xvm�2��pʽ�n4ft��[G�.���#�8x������oA��Pؼ��� �����8z�$�p���ڲYu�I\�s�~�y���п�.bWE�4�F�eF�
h��^�`�#<���tJ}^� �ORtF��oճ�Z�	f�_�?��hw���NA�:F�M�����{gq��� VsW�gT�f��"撚�0��N��E���.H�e��>���d�VJ�N:�4q��n@>���о���� qn���I%�y��_�ViM�fr��[ sXU��m��t��L�}z���?�Մ1utߊ1O�]�����'�j
z�]�l�f�f�+���&�B6U�CPZ|N��G�$��l��(J��@v��78�}��i4۴��F3�S�(�/r�qй�LY;�w&�3M��s\�)�W��X�DeR*q�������f 2V�Jƶ�+�D�}��эԪ���oL�:e���^�Ռ&����RX������s�Օ�]������D���<e�'XGҝ4��J�G`O����脿�ߠ��ݱ��8�^���?�v���-&��ҥ�^��$m�R(D$@�
Ü��t=�����3�V��އ�:D�6^=��QT�߳�/��֡
O��/�K�k��С�x�;{}�|1�h!M2��!)YT-�?��+>�w��x���5��� �G*��]�Oo1ؑ�u��C�5>�&�h���"�'���*LM��-D�d��E�s���fl�P���Td�������qN�5d���o�����{��Z����P�V�+����
�ˠ��3�`d���XcKc�5�S:�������L�K�DcF�y_-5����Fd�����d,�gf7S���S��N����_�(��8zݢ<��w���Q���t�u��Ѫ�!�j��w/�|��O�>�/QySA�ʂ�v��H��y��.�Y��yADR|7�v�H��F�__�v��¯�ߌ0�p�!���%(y���?�)q�)f\���/�<���w��F�� �vf�`"������֣au�|�]qԿ��9z�u���kΔu*�t��Hz�C�yK&�Xd���-�A������*RQpoEc���wS�¨�/�{s��!��5Dŋ������5Cጨ4�2�A��b+�J/b?�e(�֨�U ��U�H'�imu����+n��\���N2��ou'�D�|����5��>CT� ��P��%�ð�"M��sGur]�6 �bA*d��[�ҳp#�Wz����3D��R ��e_��1F���=�.[���y���W�X��+2��O$���X��/7��k�iq͓�MSZl���e-GH_O�阱|:{��0��#h�oߪ�e�w�\-����Y+��. �����ڹ&��6�K$}�	�8)��020�Ωa�Ǝ�)�U{g��F.�Y|" ���-�**	�U��nnӣ�t�O���#��n/��F �=����*|���00�l�����%������� _�x` H;&^�2�%Zh	ᤔ��˧�:�.r��Nq����C�*�ajbk�/����L�_+L���Gߖ��d�5'iE]7����Y�Zy����"}U�b�,[Z�7���O��>I��DbaRMy�;�$
Į�2����M��إ*��	F��R/���Ұ���1�2ߜ��i��o�}Dєa��6��P>�,���h7�͟a2�=���i�����,9l9����DժE�k�	`W|��T.(�\��ۉ>}����B��v5q��pm�D׼ru�.��?ߠ�i2�S�E�����ATr�kC�qi ��^l��J�J|Dit��<	`�������K� ip�-�V�eK�)^��fSſ�N�=��ĳ�D�[��� ���I�ppL�4iA�(/���g�p���־���B{�А��x��,� ��	kn�H�ڗ�q���|�<�z�K&�YrY��W��|~�5"���*�²�-�w�HiFBځ����@I/'� ��>��Ӽe���>���L�3��\�~
�$�)UM�4�����c��	(^f���	(m�!Ϲ=MZl4g�ѮF1��AY�	� UÏ��1Y�
l�F��-`��N��;�'�,\rg.�Z�Iwɤ��wH���}���G����·��	;[���pB�'�w�FGH�2s���鞇�"F����#�	��&YS�d����n��f�U���)�����<�$!2C-B�$�<���e�B�O��M���l�`Ld��Rس����Э����\odS���1-������朱�&�A#�o��8{�Y5*,èrN��.$q�5l#6"��������z�I�0�%C>��1�s;1��m������P��Xp�-�c~8P�!ab�۲�YB�d?;��QjL�t��\1�AE�Bt.Md�)0����鲬%ʦN�;o�={fcN�������Z�ePKrxl�#Bt!�9�����1���nI��9���op���WN�i�a|:�h�3��G2칙s��$���״���U*<J4�^�qY���)�4��K���;#;_'#"=�JDP`�~�݄����P�xx B��R��r�5 ���?�n�4S���0?��n���,����}Ǣd!�Q�-�������[Hk�%�X���)�ܷ��.�5��1&/�G/��7x���`W��z�5�3iÒ�~!���%����9�?�iUT�T�|�\=5��|�\�I|ޏE�1s���O{�^ԾoD�Gh�[<�
��29�S]���׫��������(k���@�u%�,j�XiKgI�Ծ8�����*�-��
�~r�G�"���%La�����d�߻zB3j!��5����a�"Ȩ-�椏ٷ���1��D�<��B� M��A�r�b�UV��1��}l�����a���"�ec�Qg5`/�1L�/��3k3]��Z��e�{��/���9�b=����n��X��eA;(�U��p�~iП���p�u�0�Y���X�����I�N�O�����o�����T��4k�g�K�t�od���PEGW��},}���q�bk����PR�_�I�!}H� �Ap��;��@!�f#�L��/���E$�A]�%p??�敮��h����7�L���e2	&@v���-�R�`\�įƜ2�4𓦴2X.e�6����`9F��f�_^{(��	X�b$�v����q͜*��s�����s
����He��݅䗽A���͐^өZ]��0����@���Ry� <�V�4��>3��ёhYjҤ8@�v�N���{v�����D�O�K��~���Ք
�.*����7�u��w�N�	������9�b��A@�EG���_^p�����AWeC}�d6���GM���G��2����6s�n����7ʌM��cz�k�<e%q��e����p�� *�%`��w��*����J�(�1&5�MΩ
Q���E|W��!��nn����U�4y���=��>���D6¹�-�lMg�b ��:Ф1
@Ϭ	���R�Ok� �8ŨJ�dּ�w�81
?�{��2`H?����e��nڱ�s��)1���z%�3��-����[-YӪ��F��Qp��L���-�3S�kTϳD�ȵ�`k��[�ěF�!���w2�Ey]�0��V�1���s^o}N¼ӏd�ِȍ�S3�"A�%ۻz6�-���'	��|�&.�������UV���6��V���}	3#`F婜��	�ES��;�]�Pn4~�����`�f�Y���u���}����TV��AK4v�����!e�nvX~ǵk��^&��wW��Ò)\ֳc��*H|��vJ+D�@FB��e�"����L�0^'|�%�!�a�KH�7�i�P%��7��_���I�+C�l��~�z��>���X�3��M��;��F�¿Q���q�e��Gʏ;E�D�Y�)��;dr�`�p�dZI%�8e�U��`I�+!���\Q�c߮�E�����Fb�Zom���~��J}��G-��Yܾ�	2e�+�h@԰�{]�Y@ax8�v�Ȃk��yQ0\��H>�0�]�uE����9�[�Ŷ�8��_dU���M*x�ݲu>1�o���}|�6�$D<��1-��>k8op����]�X2�ߘm�n6c"�t�߾-�i��t:��(Ĝ��l�«�O�B$�K~zZ�4��=j�xy���SR�wqPX܉U���yk�[��-�0o7�?������6�(P�bʠf_Gc���c.vcf���L�m�tI�s˭[��2WL��f��d�eK��)h���}����VtM�0[�Q*���q���!���6���`Q;�����yE�̙1��- ��>�)�9����-u���4�\���77��"X�s�a�0zv�^m*�9=S�q �ة7��VV�U��+4H��ڥ�P��
���L�66E~�p�o�閧�t�Z������t�(�CC��Z�W�5t��S�t~������aZ��a4^<Ц"�������&l��/_�S=�������Z��|�d�I��re�xk�&a��ċU+���[uh~y���rm��g�5�{i[����Z���?����bGH�4��m�s���Z�/�(9ZGͯuՊ̼�T0�f�d@�&�d8��8���t���o���k����]�۬������ç �A�.~��5�J��IQ,/�/f���rf�������ϖ�NSEQ��BU_�p|?���į�5S�hl�f���[ZrF>���S7Fe�8j�bG�>ڿƍ�3�L�ώ'�Ɏ���ؔde�^��z��������Z�~$J�\@��:1_��b�U-����L����*�f��	��:�mR)/�I�ғ��E�|ڀz#�{T3\�Yz;��s铹�Ɉmٝ=4#��7RTl�h�J���?q !��A�BK��BD����]p?8��ϛ\/؈a��ra�E�p�����W�>�XF8� 飹0��eI0�=?~$lܒ��Y�5ϟD"YH����� ���R�����n�lE�U�P�<M��7�|��F�g~
P8}�E<rfL���X#�v7�浐i�f�2����� �i-~�?�f_C�e��=�`X���$�hu�j��K�;,"n�|4fp�F�þ��t|��H~��_C,��Q�z�?C���_B���4W�W���w��Q�ҫ6���~u@��������F%`$)���"���n���}�"d�a�)���� �b�Fr�5���9��f;/�qa�^��U�;�.&0z�Mb�2�i�=F�ze��k9q�s�ڊ�LEE7h��}5Xw�'O������ ���D���OЍ�9*/O��k�U��eW\G�|n ]��؛�����6
z�?h�_"0�؎��to��ivxBx�y�,U��^8�#�q#K:DK�4�A 4>�#E�r�)˺���a���*@�7_�+��н�^Lm{�-j�E���*��Vk���m�� �K7)� W�*��XLK���#����6��|�e�α����\`��ݹ�# ����rTB���@m�s�2S�2z58
Ɔ���!������}�s�SV�:�5��g�fM�G�O2Q��e܇���j#� ��4Q|3�����_����b���Sà�H��H�\���nga�'��+����6�9}Ϣ�P����l�<RXhO��m.m��,�D0�P}A/�v��|jׇ�|2�J7���T�mߨJ�O谤zje7�Ҹ�%uv]N�f�2͹��Ƶ8�J�K{��8�b�˘�M�_Y2�3,]2�� ���Je��]W��ug��ȉ��3�	X��M-�n�}����!���$�-q�s�$t�Tq��(�#mE���1P�u������lm<5�߅�S����($W�������ȩ�&����!�'�`��g����f����*<�����n��hw�?M�gi|''*�r=�U$�!�h�b H�e�_�k���v��`�lA1Ju���[�:�c�u[�����6}A4:	"����x|8 d=�VZR������c�f7cdy�[�	Ly�ۋ�(�n	�8U�ĕw;߱���jR-1[��2�� %�OI@˭�r�?�\��4�7�Dg
�K��2�/U5�Og�E3���ꈚO"0ok���giX��`P�8����addE�%N���P����G�~0E?Ч��:���2��I,�\��F�S_�!�|P(i�S��{&f46������Vfzo+Hu�B%�KNC��߱	vZa�Mz&٨��Yw���1����j��I?�rўL���j��*��ᵮ�眖R�j��_B�m��Y�1�s�������"��������7+r(�u���!�pW����,���(��F�JqVS�Ȑ��Fp]	�u�eשn.w�.�l����0�8��
i�����Wu՘'��QF���7�MgKASl�F㺟�ߖY3ԧ�Y!)t� ��.�a��"��i�/���F;�$.�\n#�A����#�
�P�KT/�˧���i��_�H@$�|w*e�G:9���e�zv�R9?u�Xp�[��U��>E��q'�BRDp�� �F5�]bY�Q�WI]MtV#w�l��O|����v�A��&g}�T*덄!����Q�3?�Z��?����0�����lˊ�*\̩��ש(4�	_�-&�~��$��|n�-�d`Olo^ɥ9���@���*�h/��ĳ�zW��T��L�ʴ�R��<f��*t�f�N�m�%�lw ��(,��?����}�lb��E�*�+����T1����99�8d��_�0�.zLZ���o'��[�=
1���C���F?�B= �aEH&J@;f
y��������^mwU̱E?�ɛhz��6D��}s�F��%�4��K�f9+A]�`;�x7����>��	���8>Re���zsΛ�< l=�T�=
��1z� }��r\�pt����¨FK}������,S������S���Υ}�i�I�~/Un4�3�]��	���үk�w����;��ѕg�2o�h+geѓR�@�li`mU<G��)w��#�W@�4�a��	�A��*�c&׽�@"0`����P���WH�'p5�3l���)�#b:��3~�ַ��7!3+�r��c��I�{�F���T�����V��jO���[w��C
v?�l��$YqFC�*�ZD$�ག'�^��/��\G>Z�U[��-Uf?Dj˻�n�d���ʭ���D���&8q���T�I�~A
ar��z�����*�z�������ۀ;�;h�(l�
�Qo�(r�t c֗��@4����72��|`(N����t�f�����>�((G>�~s�n����\�v��̹C��wׅ&�>�J^�b�K�n��_�U���/�_�/��E��T�mZqI���x4/�{��ܦ"��ru�=���TO�S��1��~�F���c� �j�{��$nh�K��>���L�E�汗�ev�:���7jA�EN��~+��'�،��=S~�O<�����g~4a�Q��8z�_$��W��F��{�贞t1�������o���p�2l�it"HD]9�>)5����3�'z_����4T���6���Q��#��hTMt�';���#�$��F�s�/aԋM˦���6őX��ۘ�)������x}A�r�`�	@��T�!�2
'�['(�#��Db�%�ce��n87�ES�G�	Xؖ��W�-;2���cs �!+n��ʲ�DvZ��S~نSCd��͙>>*�~��w@56�����c���Vy��62Y	���\@��Xi':u��-��q����|����ڵ/���ϸ���!%Dai�
�M�ЂjO���p�m��c�dr.�sc3���#�.=ь�F��S�������h��|���WYY��nC�$�Jm�f&l��ToB�*����7����L�`7�k�C���K�J�`ՎڝG��o�\�@���%��ҳ�a���̏Ƿ(��_���d��Ӛ���]p|Y'5�uz�#kP�o�[�pr zդK��Z��C�V@�D�f��ئ/�z��P��	�&���0I�G���V(AWW�䧂u�g�������p��Q�a\1���6	S��<D��2xv)���H�sN�H�Öb�%�5��� 4j!s8':(��13ؐp!�M��m�X���H�ĲiM�CԲ�r�N�����]#�~#��~����=wj8�f��k9Ī4��{UT��?�pJ�Y+�K���~o5��1�y��î{�"�Y�묤��S�g�0�=��,�e`���Ox;��»=��1���>q x��,U������?��Vu��A��n��o���A0�ә]�|'��ȧ zG_��Ѹ��ypU	�G~-J�_� g�k@���=�l[$'�S���MW.F���b��q��-�ՠ�q�6��h�9VJ�Ed�U˼�A����˰\��k�V�6�)n K�#P~��i7rs�nM��;Ò�Fi/����v�7Sa~��3y}����L��a��,O�}]�'̯�d"T:;�v�Z��Ü/DXp�4w��n��?t��G�P�:2}&q8���S�rs�A�(����t�-n4��D�L'j�v�%��y4-� 4P*�_�	�,��;"-�����iR�aV�Gc6T�V�w)T� "mE�)����d�u(�0W�R3�e��#�_[	�|� PX���o��z)%Զ�)ӪYZ�p��3�L��O�ep�@��ι�U�YE�z"(
w��®� ��ẔH6���S{
�N���`�c��A@!�4}"J4v�UL��k~_����b�w_���:��E�k�m|C�o�
S5��
1�L�`,[gl��3�?���0i~5k�������tI$��32iJ������v8�u"�	yZ��)�=�L����!��p��p��բ@���B��;Y�ԧ橢�ӆm>�k��~�qY3m\��"fCr~)A�=5���=(��)F̮�>�O�s#*��h��lG� �L���`#^S#f.�#����"�s-��r\"G����)�T����@�
`�8b������C._�6���de)L�)��6�:{)[�g><dS�'�H��|N*��D�S�@��a��ա�?U��R�p5�覻����x<.��c<��=o�
�:�v2wR)����+��]\����!ؤ�3��6�p���ݲ���7xr±����t�r8�!�R���oV`2o�R�*��G)�ד�~QJ�v[C>=G5\���A-��OƮ�i�2���,�0C�0�xA%ս@��6T�9��m
@7�l�AJȤ-e{}�'u �����U����.j1H���(<���}47��y@c�L���i�>��D��:�"�*�Hu�/r3�
��ڦ �.3�qŦ]����?�^�e�n8��z���LczOA{�pNr5�=��h�U"1#h�N<?szC�s�K���S��2V�M�#Ќ �._�#˲0�py�7c'oHGث�cSy�g��F�$Qw��ĐK����WP��̊�ye�4'=A&�jy��vW��"�	��*�#Z�N��UV����CO\����Fu��՗������j��.*�J�/Du�|?(D:��}�u3�焥�̪gjO ހ���)��R'����8�Ot�!�����!N]`*X��v�@"��#��'~Pg����2 �?&^!�Au�ȣ�Q�f["gp���?ŶƐp���E�dC�Lq�êe*�#��i��g��-W�fک[p�6�ؽ�����O�̕3��3��sY,��{4 ���_d�?���iv�����|����s�1�ًH�C�Za���^��MΪ$7����gp*�A�Q�çw)����W����\�O��l��_n�t3�3����	;_w����]4�v8��gu�Sf7��eC�AGa	���GP���{_5x��D�&��Ɇ\0V�f<�٘��H�]��}c��Hrs�y�&�R]#��n����\R�d�n��Y��JOޤ�H:"FDF�'M}���.W�.T荌�$o��#N��s��/�+�Y�	=�?��U�Nh�zǓR�y�����ӵ �;����Rh��~)\���	�I�Ȑ�5������&�Wx��u�����BBRP��x�l-q�u�}�P�?��V����Z���^��0���j��ʐ��"���5����d�4n����JN��@}5aA��	K��75�8_�";�����i*;��6���f�Y��Rz~���;L��YS�9�;k���g�p�#.Sq���f4�?-���3���ش�,8'��j� {�o��|J@4�?���z"��] Va"��Wc�g��z}�m�e�9�=�G�gq8]
n�?xo����3��#�&��L���Ncm��E0 �ϐ�1yA�����ҟ�.�of���@��kp�2��v�2�t�h��W\+����M�w�%�V�i���Y��Fr�����.iʗ�2�a]H�_��(ؾS+��hP u�M��ۚ��z��@K-�M���˄�
C�-?��6Ո�s�� �W!�������73���?�0�0'~\��Ă3fA�Q,e��B���/���GB$J������w��P�f�<���P�\�Π�qd�5�@�v����	���D׬�Re�B4�N-�r���L����Kc�����^��gj	X^�\w��ᮒ������� i-����R[@K�T.���qa汔��7�~�=�Z�e*�r͵�s��
�248'8O���>3����N
������0��?Ƞ&N��kQI�%�h-�Rm;�ɫT�
�̦$F=<��x�q�|��,��f�dӣ��^�?��k�yhϜ�ۢ+*��� ����h~�����v�Vo3�Lo̗1_IYsb�i���j��	41�B���vQ�3MN9�l�O��7���
_I�e�ݽQ�g�L�y�b��
���9aG���R-���=��l��*�9c���Ca�޼Z���=H�C��+��r�
(?��(R�hG-bk��{2H�e]�)nQ�W�.R�b-j�P���b�/��Ar�Z����8�Vc.�D��6@=�w'2�&�r)y���yUH����(�c�ean?��GT>-��C���"�}l�؆���A5D�AL�����;?5Ly�׷\� ңN����I
��hL��y�S!��6�@������╷��MXvЇ�_���dc�rg^��ݝ�!�1F��?�ی6(���m�tEf���i�$evV�Yu����5�	�lU��������F[ xL���������	j�]/�O��wu�wX�i¨��Gǈ�C�Ƕ	�6�n�n͈>�I#����B�8Vzۜ�ϋ[ܕ{ս��q�D�xwW���R֚)
W�L�r�b0F�ZjF�BC*7��=���r}z--T,�E o��K
�����b�����Ŧ]<L	~�7�����vro�P���;�M�߀���DT�@0����(��:��l�/"��L���"�
-�r>�i�-�#;���qؾ�Z���f�Iʼf�fp�J��Uh�Zd[�p��	�ǞK��Y�RCS���}�h�4X����z�L�2e׌u�r �V���9��Hc@]���c{3���/���CFGe��0G��L�ԝ�[|{�@��2`�lz�VU��m0:	�5�X���^k�=��M�=3�L�S�5�Q�
�'Ae�Өɣ�]��m�A�!T�����!?{3)A�X=�90��I���6tg<�	�?�0����Ϛ^~����uJ�G������(j�(��C�"%��w�3�Sԟ�s��
�����s�����zĠ?�/��ٻGmB�+X��nP�G�m�>i���uĮ��d!�>�̝�9�w��%>�����(�*Gn��I��3)i���㽴SS9�1rhjENC�Ы`󡟗*���ᰯp��+:�������7Nyl�'���U�
6���G���	�$v�՜5U\��_m��?��� ����jP�U��Ï{�`f�y�z5�:�t��XًI�����[%�׈!�j/F����Q��5��8;O����5R��R;�;JV���|1���j�Z���qپ�Gz}`HQR����O�s���ɪev��1�!(�z����%Ul�q��WR���HKD�%��i�>���|:,�o��/�}�Sr�������w�;�K�O��.)�Ga4ZmQ� �\H�W��Hm5I	ԧY��=b��u��jW/�R!���9D�v?lQ�ޣ��n�VR�l䃐�(O\�6c$�a���8��fx�Fx==ݎ(L(�FӺ��R�4<�P��Ɉ[lt�X�U�F���؄G��97�#�X�;����[ˆ$�P䂽~~X[Ώ��;��x�ۃ�v�mNMj��A��-���9ך5������;�={���ox:�w��G������cT
����Mv_�i �M�U[�WIά��8v��Bc������R��l�)��.ҳ�
��Xy�C����C Ǽ=�k�)�;�;�P�Ξ����<�&�Bë��0� E��^L{��B�(i�+��|Sݾ0��1�R�8=�a<iG����O^"=1*�5�Z�D��� j��e�\�K��ip�����i���������ZP%>Q=]OMY_\��r�����?�ؚ%�����l34���+�b⼄s�Џ�q����k,]��4h,Q���#�K�z"��<�J}�,���>U��ƥ̮]\d{�5�PT�L�����Y�D�?:Sa�5�t�� ��(�b���/0F�G�_ Z�����5�G�b[8`6��Uk�[K�o8�~Wޟ��Ul�I2��U�/~+�z���~�#S)��Xu��)�¹I��׿����m M�i��Ao���L�i���Qmw�5fj����m�y_��	�3jTPN�J��v�'�\X~��4 �A�A�~���Ӳ���F7e�?D>e[5"�t/Y�L��ʂ�������IZGPg�vt��.!�W��7
	�^�vH
BP���:R�!�8(0��BH'�,nW���}Jŭ�Й~�K@H�b� ���0e�������� �Z�n�!֎X3إ��B�_��#�'��[���$~	J5�,ml"E�xP�KVO���"�؄)cB$F�~�V��|9��~�L����x%�Z�]��#[�5�2��`�T��g��glf�5�NZ� <����O�j���	j����O�l�A&�'#P�6^!����Ӟ������H��ׁ��bI!���6inX � }Y�;�g��Hf&�.���Kƶ�R�G���{���)�`�I������%!��X/�ǀ�T�"^��$��2_�� �o�n�x�❔jɷY���v���*����b_�}�
�ӏC�?���'��q`R?K	I�V���7l����.j�ü�P�sA-�`�^���
s*�����Q�5t%S���U�vɉ���1�Q��|�Q���0�rrq=y��i򬒽�;_�K�0+���p~1=qՅ�W�ˑ�����m�I��}�\�{��b���T�S��/#��= �Yk'��v@,�C��6��������O���=���
&���MzՌcoD)Z�ѭy����Lw��/M��և�E�Qcg�) ���9 ;R����u�r���U֑gT��~����$�֣@/�aGx�\�b�֞�G'G�Ơn󸿷����k	?�����->�a����pl/����5�PD�aϙ�\vR�l�+mK%�~�~�E�����q��	�jQ@E�-��r6TL̦��ʰ����f7��� �um�g�[��9�y��v2�uO�e!m��~v�{�X�Gw_t�Cro��Q�^��8�����}��x0+?X�b�!0�R*q=|���j_M����ָp��ט�s���b��~��x�ͼ=3���/Nٱ%��?لJ��w�Z����i�����[^�'��FK�Uxy����a�[��ـ���M�{���Zz� 0��.��~��0ֻ���x��/�������uE��'� �mֆ砭�"iZ��ӕ�������r,�{æs&&9�ݤ�e|�]|Q��ʟ��&�Ƴc�拀y����1-�=�׃0mr%i9��5������Ab�x�f�4�QR��T�BScy�*�Tz��ゅx�K���`������w3��kR3dv�o'�r�6 ��7�Sh�ly$� @�uً%k�ӳTG��]���1Tc΀ց�g����r�Hz�z�ȇ�z|8�]oo�a��tE���:�{^��<�8���y�f���*�A�8�k��8�]*��^����B�G*qN�$����s=�l���ڽ)#�r��]Yj�f�8To�B����y���?)�ɿ}������	��? ��,�N�	�D� UzZ?��z灓[���ҷ�HUf@!��Mz���/r��;�>�08`b��ڝ�s�(��؜��~n�H�}���*Ճ��,�<A�T��*�W��h�^E��p�{��K��1C��I�3�#�t��\s�)ƣ�z��ޣv3�	��Z�:��P`���=^_wj��P�*f��rx�ْ���2Q�ILC��*��7���mY��f�����U��e�w�1���"v��	2J�n��:<*�ю�'����,������eY.lʔ�X�V�sVQ�Ӝ�}}Q�I�1�@:���F|�3����� u	)������ܜ�ْ�A���oz�)�i����x��"{L|؀���M�FQ]��3=��xm�X�Q�YX�5%�����K��>^h��Y���q^������TFڵkƇ>297��B	 ���vW�]:$�$�7����P���iX0��Ip2#�k���h2T��qVTFV���Cz	�	z$��N��������\�1b=�慛"F(�U[xʊ �����3:h]!��W=q|����'��ŗZ)���VO��Ɂ�!�Ti������e��	�Y[�����_0R���v�e��$!�@6m���	W@���uG��E��{��բ�]ho�ˤ����6��g�B����i^�	�9J���
\�`���8�lS-�K(���ږ:������+n��I-�B/���Sq
f\�rj��p/gWI�I��[UH��ԛfo���ƜX��_cY:n[�	��8�@��ս3��ɛ�O\��Z��]�W�SyS&�!b����W�+����fU��&W�F��.��
�qp��P��Ƨ�Kv<#/)���o��ɳ�@A���! ����EIYxo4�޻�O��I9�!V��=���_��1JdUjةE����	��2?-��e�ۊic����+��&�O�Nϝ��b6m��������8E��i��,$m��-aN['s&Ma�Ljqڇ�1�������\�B[%j��B��B쀄�!�xw��*�'g֒�#���N�_�6��r�~�j�� ;d�T���!~����#[](~�A�}�a�7�=ut.�(YS��D�m��NcTG�MF���I��V�C�Mg�BT� �n���C�3e֎��n���1�t�h�X[Y��Z?�{�����$�FK��z��r��뻜u�ȕ�{֖�U������o&Ҋ('�3�f�p�4[!t���Ӎx��uޚo\xF�S�I�Q�K���T`�Jͽ�&��a�i�]?��Ҹڲ _��{�r꺑K�z~���	A�A9���B�'wt��������g�����9w�>���HR=��L"&$�b:�I����SR���g��#���f�-t(r�Hڌ���/o1���B � �jT�H�+�L�M3%�E9�Zs+�e��[B�e��w�H�i�<X�6;�g�bSB׳pg�e��Cho��� L��{�8@U�)����;�[c�~s\����!�(�x��P��tO�79q�џf��
ej]#��ӣN��T�`�y
.T��?%�����Շ�V獜���4���K}��-�� ����E[���/x­��"�[����a.����r��)t��wI�q�`�)�|���f�|�<i�v�� ��ؼ1M��W�o�h.#��^��q�YE��܆��,��9��+Q���U9��gc�G% ���`��(���w{����vI/�3S#��&�)/��Oi��>�ѭ��z�2?���x�Wp����`�E#�#8K�{�N|؋\��g��f6D�:�SE�7EV�Ril�xk0U�R]�]>�o$bE�V4w�Ĥ����g~�C��Ep�]5�R��_$���b�l�E��^ݴ[w� $*�}�w���� ��5>z֐��nS�b�b�s��ϒ��9��0즖,,�G���J�Z��*$����OkO��l� $$�Y(|k��͑XD8�yK�)�]���l�Z�H���}d�{��b�dؿvO?]_8J�c�{�Y�HO�+����$I4�35u]�)���s���S�=�
���7�/^'��}T�c�D�)�^�I�:l�����yp"�֗�@�<Qw���Ų�- 1i����q����*�:���eДh�>�DC���KT����@l�hi�4�8/oI�I�W�3�	��#��̦+x'��4�2R����\*v���լĖ�!%cBT�%�Y�ؑZrj����y�9���7r*ێ�(bOd1��2�������q?,��W[�D�Z����Ə#vӫv�����'(���@h�G�Q���_\{��u{G.e��ǯa�k!�+I"��M���A��g���6�C�-�@q/10�W�t�gpi$��gf�ɮ�<�@mk(�@�q����2��^�i��sL+����e��*�I9_�XY�iEԙ(dJ��(�cd�MW��Zėӱ�	�Ln
}I��]�z�?�7�埊��G�����ܗ�;������z1 b��;���b�~qp�h�C�?����4��zz՜.F2��q�zU�/�\[�ߕc�Պ��>��~"�Ⱦ�,�6ƕ`l>���+N��Ն�f��J����/�sE8�G����2y�)�������	�Y��;',�1v�P]d�Z�vd%G�X:XT�l�Zz�6�����"O����-,�0�����Έ�cec���p���^�G�x6�#%⾉�p�rJL�z�E�q������$e~��;��+Ɣ��Ǎ���DD�ݰ� �7��I��A�ǫ�w˙����"���������,:�?��#AS
6�c)78�����t��	G�k��?��=dCDzG�%n(���g�yo:�����m�̦�S���vj�/t����{�G �p�"���Yh�G%�c��tB/M����^3��^��E���j��xp�BP� �i���ͬ���1�,#����{#ށ�'�����?4��d��f�����n�f�btb�i���1���1�CFgD�7	.��H�4���o�9^�k�<1&c�}��^��_��p90�@8$4
U?b�,�8T�8FK���aQ]�ԴBH;)CX�|{�L�5�r��b�`>X�V��J�(!<�g�&�M�4H����
�.�;�*]�����B�u@�Y]��z���2�<Z��"�\���I{
��:}m�	S�$����%BE��w)0�L3��tp�o����S�_ƺ��(�I&�=#i�f��� ,�y��5� ��:Ļ��܆L�ޯ�V���^��r:s_E�s��Q�p��	s�����pu��p#�{��Z�Uƭ���V=5pM瀣��Zi�L�#m�b)�]K_G�r��e�)��=�ĥ�;���a�%�m�
�I*�� ��-<KY��^؇��0x���5zUT�{�"���7%���f��7��6�J��ޢ�59���y�Nu�b��@�d^��`8�\0j���#N�ZL���B�|���)0��P}�
�H���~ѥ��zK(�~LN�N���P��C�T�	�SD��h���������dw�2���!��:�f���9g��Ǩ�YU��7�Ť���T$����F��o�n��^���p�~�c� e�m�&'|6~���V+���p��X9HH����l �&��3�G�&�zU��0��L�O����6ⴍ�J*���;��*D{�}a�7|��)�۠y�UΎB~�.�w4s����8�m}43(%	n3�E_߆uSm��(-��Z�yk���EL�O*G�7�$#�
(��^��ק�Oh�6����=�>��j�h+�0b,�;d����=�cP����ٕd}���/��#���ҽ[ǩv��0�����Bdqպ�}*�/I�����7S�y�0���?M=d2&�e5�&��lҨ�A�P���|�$�ۨ��h7HOW�	����9g�+kh���ˏ�N�]�a�̫��e���}r��տ���!I�p��Dh��b
�I���W�g��t��@��r��8�$�l�����o\��6sٟV3���ީ�\0z���[!l��cy�<���{KT��Q?�����?ϐ���/��7�����z@C��M^a�>~k�|�K��?�<��M I�8��Z�����>��W���=J�+U�g�#Je��H��2I���y��Q�@J頀]f�C:u��qeO<�޼���������H��n�̍ Nψq�$p9�f�K�b��gح�����>�x��f��f^I��7��������Օ���b���]r��/S�l<�b��!XY�Axb�������&
ۃ���$�������Dc�f�K	\�^ӏڲ �m�w*A�Щ@�*���τ�Ջv_D$M&��Beb�㻙x+�b4��a���2��N61o�ѭ�b(�G�QP�0fK���Q���qne�4Q`�&h������g|QS|����a�{�����p���ۡE#B�rw��gZ�L�Y�uo�Ѽ�����{�c7*��+7�������N�OŠ���X/݋������'�wc�Ɲy0��	�n������<*'�^���~P��բh�_%F�����^�����k�Z��j<.j�Ǵ�t�r��1��T��7d��3��]UA�%l�#��m-�=_� ���[���֯np�P�O�w��T$+/�v��Ξ��˿8oQڈ�Y.�V�?l��66\��^���j�,_�&=�QF2�h��l���W���_�-���F]���n�j���"|�z�_� Mٝ��v%��
�8���܃��R�iN7*����Dň�teo�
o��!�� B�E)�D���l�P\!C�ڞ=!��J�I�j"��{����>�(R�t��8�%=}o��HT��9��oځQ���*�_:�F��r��kqj�u��@��{�9x�d�Y(���v��8]ch��9�L�Wđ�-Ck�?�:wq�7�>6�9_$��b��wYDy �h2<�|J���*��v82XMV����
nvD`���Շ���]V��Ky\t� �)ADB�AOj}޵�����n����s���yz��s�l��p �/���[�:�ݥ�J[�>ҫk�Sz�_ ✚�Az�G<M�H뉇�CR����SH:��4[���mZ򀭅ƞ�j���ݶZ.c�4_[��^�����q�D:�7s�؍TVu���*��5p!"��P����й���u����h9S&4����zl�"��4j��Q3�����������<�2|!�A9Wd=)h�������!A��v�r�Hvb�v�E�0��vK��
.�뎮�o�>��\���P���#p8�� ��r��׮	�?�G���v����9��8�?rgh����,�F�p�r��{�*��&�0�vt��xޕ�A=��r��Ni�:��/`��*J�L�h�����ET����,�#�Wf�(�#�&I��$��2E�T{de2�MC ��$�#{�HJNct/s�7���+�Z.)������F�KhFjd�VeϦ�u� ����a�;�F�.�(�v�?�,��sH`��D$2N���4��❺#Mqh�z�To�fڊ�ph��� G��v`��2��	[� 	�t$H�r�Uu|_����&�G
Cz�<��כ#���Hbk2���>՘kX��xJy9.�HN�[��ӝwV�Ax�m|НǍI͎���	��U�}��`�'�a��r��%�ȕ#G�PHL�Ue�D>Ȏ8eY��`�$��U���W5��_NupKQz)�N/3�;v��bx���a�"�̉!���!�- |X���z��OOu��	9��y�w���@�d��l���")��r&���!P�f��뉌����mR�>�����gy=!��g@G�/d�L��}�u8����2�� ���rL 9j�X��utP��2����5��]�`tS)���9f��&�W
�%���4'�Z�t�������թ:*���`wL���\��{��	��ʄ�kE��'+g����'�6�إn%6&i�	-����
���Ow׈�������=��x�A��ǎ� A���#�P�j�h���/�Lʿ���04ƙs�ϝr���( P�����x� ��S�s�����6����A,sr�-�
���g���W�_��V�5�V��0°u���A������C\J��)��t��7�d��N`���ڊ-Pɹi���S���՚"���ky�P|�������4�ԪУ�w� �̟�7m]|��qі��l}�\F��^���66&�9f��o��/�����w�B���fK� ��M�c+���)��PG��<�ucT���óW A��y�:�B=xvS T|�ƛ	��9�Q;�+��kQ�љ�挀��V�ȔMl0��l/�)�-l�4ʘ>��@s���Rv8�p>ƿZf��C��Ƀܽ�c�'����i���v7�������L��P�O��SP�n�h�ڕֹSo�<d�%�8��zmvx�^��1/g��r�#�t}�? �r)��x|���q	)?p�|N�8�H�gK���c4��{y�8�	KJ�+��D�Zj��M����Y�mwX�_R@��F,,�i">Af��ư��}aDӟyO��L����f�,���^���ұ��U�������_�u����?HSo�ͭ�!���Y��2aGu�hӹ:m��^��e������8�]E�y/VAv�:l)5;<\���<�>˯xRO7�S���%*�e���6���*���\��� �B����~MD|�$�nz�E�+9G�o��$P���w���~�lhPȞ�!� ��S�juL`ŭ1�Z�=v߽t�э�`���`M�*^ۧM6uy�'u����@e��������ɛ9:�1kT�e���4nf4uÛ������ܠT�B�tg
��pbG�L[�C�Y�΋�\�m�o��Ys���	��2q����m:éL`~#�#Is7'ZnGk�mB��
��y������c��ERӫ@�%AW���W���o��nf�q�����kxkg
�y�_�pG��i-:�@�]�A�y��o�K�����]n�򃷗׎���6�㨠��@����)��+���ܐgq:�v[/��'��͸�S��N�TP�yV�t��‏�0J�}k\�˓��YS���C��ٳY� ���(���-������j�9�D����AB�X'�ݬ�{U�v�X�����5B�$x�1�|�>+�7}�z�w��W}#fv��A�������"�T����O�D$Y�s?�%wp��ﷰCK�H��M�c���=Jtڷ�+�r_%�ZS`@�j��

�F/QQ���!�f�((�U��B�%L����l�Co�ZoJ�)�C��Cq�6r�˳�f��̞��1W&�>�~����QʔP�K9cP:�&eϥܭ1���k(G��(��Ԃ��/*�����,���;z��n8�*��;�-{$�Ry.�.��8xkSB�T�3/-�mY��N�:�_q����f.F�\�6��T�v�*��ď���'�s���&����4�m7W�Q�����5H�A�=�v����q���&by2#i�<�.�+��]B�sy