��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B����R����l�JxM%�$$���E`�����o)lh
6[#V&L�.2�%���1��(|6����"o���F�Q�,���-eQZ��m4�`�b(�I���w2�Λn�J�~������%@��~��� `aG<l~�tG&9��!���Щ� �;գc]���6`�AO鞱����r���D_?���0�����a/��3oE�p�:>�]������+��M�Q�'̌�����{	%�92�L�,ԋvm]�"3�F��Lr򱗼ݣ�65�R�?�}5Jj�%0Š������'�P$f~Ad
ң<Be�7Z��4U`oHj��3���܅K@��6��	����u��//���Z��ŉY�3�[37jV葝��;�[�˟h�ą�x-5��aDX�:�/�)���@F��+W�Z42a����G�>�mr��ʢ	kmǨ�����x>��!���y0c~}P��?��&�"G��n��E����oBjP������x'��*Zx��H&�LjϢ�A�Wg�3|�y)-�&{Om4X��Nn�N{:ӲH�wL�Op0��� ��9�ξ2cXHOmۢȕ��ʵ���ֹr��}�t��y��ܰ�y��bG��-� ��]3��ȁ3�&���$X6Hs�@��[6���g��lc�\y��6�U�z�:���H/�"h�T�d֟��Ʊ�C.ߩ���_��	*`ۑLj�'����X �K&d��>��Lc�L�h�٦���y�$]�� ��24 �R��!��Bn�~�!��O��>Uz�J�n�0��E/��."᯳?�`�LB@WF~<�HǿA��;���?�>G,D�0`�l�ګ%��(��ѹŘ&�U23G�B�Ihٮ-��5"?��~r�������"BW
���΂~�����eH��Y|�XPp�5+�뫂���c��B�B .��Ow+G��5�[��n��َ���d��H�����D"U�U�Ρ:d�Q�ݖ��E�� u���ݺs��Tǡ�iR	���;F��k�yODå�� P�_Z�Q��ܞ�nܖ�_N�F)��VnO��\)�����L�X�L��r\�-��&çrÜw�y��W�&l�m��r�:�_�����ĥ�5:73�t�R	�&�N�ȁ��t����t߭���6b0�nLh�SrXV�����F�Ǯ0�yy�TAP0��W�l�:Bk��i����"Ȗ��IV�J&�*�kW�H��C�w���o��x�sV�v�NO��]�JOrx�������I���G�0p(�]���2�/����a� ʍ�\y˅�0�}X����sA�&�@2C{���b۞�kU;��Aq��ζQ{���� |E�Y�F���{���C�AJ�D�0�(�-����Ü�iZ�������0��yC{��Ol3���vp'7�3��Ca�����I�9���1j��U�l��z���Nn�#�WI�{O�����1���h*�d��ӡb�����{�q��@������]�wH��)B��R�:6e[�О\4����đ�]Du��y�\+�~���/!3"2�!L��g���%���w�{�5��˲[ތ&:Ҥ�u��&4o��1�z�ow�{��߉Eg8��=���J0WXHB����D��\'
��1�
@E�֤:ך7�.�W��ȍ����CDEZ�݈;`�1�~Ô�k�L�(�K{&��6H��j�����O(a�[y??�l���Ұ�[ʰ�C��|j=�/�`��L���t��n\����-F���@§��_�C����CN�{���M�ĭ�ދ� �����!�S}}Ɨ�t��q�O�C��mp#�U]�_7)�	��>	Ho���w#2�V0��:�p����엝R揃���%h?'�v؈�b�Rg��٢�����������$���ojf��VV���g��!2���!Uy�4��z���)M>u�c�#_d�z������g��$�2w��TkZk�-U���p�g�_;/R�Hc��dQ��K��x75[��Zr�m�
�{����BݗY;��T�%��/�y
��Q��k���b��~� �u`�gtoH�.=X�d/N�r"s#����b<����nw�`��m[,���R����*�����?����ԩfu]�h�u�O�u�������Ok�	���J����hi\&��%�v�ַ�&��"����k.@΃���?)��K��?�;��"D������Y�0V[��I,?]mg5<K��ٝZ�A��(���j&��Ȅy�C�s�a�P��ugx+q�ғU��b�o���o>�U�=�
��t��LO�����i�e���Ц�p~?�XP��x�,�h�i@��>��4J�Q�M[m�L�6��=ՙ��z��:ٍ#:�Q�6Q�-~�bb������sD駮�KD������:��!���t}OX���m0ZcQ@�Y���"s]�*��֖L'R�����ż���@l��pz��q>P,g�p���pgV��5��z�㫀��$�z'�Ռ�*0	@gI���اAR�lq�!����1�9D鵢_uwץ�&>�1���rя6�ta�N+[1��?�ӂK��Q�8>i7�0�n���C����n��|t�e���P�����9�&��a�zVCSW�N����Akk�-o�|��v�(���@�b �R���E$�l/�禐W%\��)G����b��Aa���L�N�J�r�\oΈp��趤�T�%�~�W��:"��<t3i(gp�X�D_��L�U�{z �ICK32�����p(�[�(i�l迕Q����v��<<��'�yz)�X$�qS�3�"m;��m��$|ťR�E����1�3d��!������	r͉?���\��|u�K �/�dId�:���]f/�PIOpUuk-z�u�J�����x.r�lێl�?7�/���d-�]\Sa�2J�ৃ.���!F:B[Z]C�G���|"vV��s.��3�qa"�w�L_,�q�&'<���[O�e��<\���8���L����G�3B�9Ŷ��x�M��̫���6�6S-Y5��r��O
PL��+���Ё&/��?��l�����=wֽq�v�a�Ij:F�	-o��K �]ļ����͋Ų����]f���סp�0��\���s!����[�_����!�5�'' �L�`���M�Nz���FO�ٴ���|\���>�dhc5�Pc��ߎ]%8�Eu{�f�"�Q)���� ��4�5��N���V��Й�D(|{}�\�Y�;�<�x�O�۶%�����?4�Ʊ��h�x��l�:�M�¿,�7�$_F�tg���e/�
Q��l��g?���_��{gՊ�q���1%V��n�#��������݌��rh2O(�Ȏ ���_�,b�s����@�~�1���Wӣ�PI+��
��ځ'������p��C\�j���s�A2�xwv��-p��F�����f���z!�R.x$uT�ϒů�4m��0I�ъ�܎������5[	@��kqo��1�����/���Nhyq�o��I�C���A�V#ɾ8ƺH�6Җ��7یku��d�M�to^�0���2����_��ka��g A栩"�z���$5��.�n�����5S�!��_	<�Я��նdA���ќ���)/��/fO4&��Va?�e�"�BRֿ�]�wg��4�n/`nj���du���[L��?�`���uR���*���١@Y����N�
�\��1�k�q���U��dd2S"�ӳ����|�g!ذ>e�w����z�����M���x��~gp�^����'�f����ǣm��)��qQ���i\����R�]���cy9	j^�7��B8��P�2�@GXA/*�d�덦�u)����3�f�>�3���{�9磀,G$V��!��Y����"���/���=�1aۚ���aJg�;P��i��Q}���X���>��@�,�-lo�(ӛ��gH�� p��N����ڒ��q:��uK?��5?.����=��#q�4�?�X'�v���G/Ȧ�ʤ� 9��g"�V>���F��w�6�p������������,��nڤ�dM��O?�;};�ow�Y~�
oC�zLҋ#��G)���$��ewu
ا.��>f&�����2�Ei��@׳��Bݴ2�o݁"a�O�]x�ԙ��F_'0�&������u��\5���o¼h��R��s��,Ğ�2�9e%��	��PM9[�M�'TE�75��Ļ�W��H"��O���a��0���)��-Ӯܷ��u��5���
5��L��nN��0�\�!kߘTcaT;39�-�͸q}��f���Je|������+��cwB��T�H�h���9<DS����Q}x�;��X���e�t��[��ڸ�@�*�8|T>�B��ӲՃ�~_0gr�X�l𯑷��m%���`Q�tP��s�8Pz�0ht��8Eh:*��f��`}˨&��f5�2����="k9m�ͺ�������1�$�.��rwd�E���:�Tk�t�&pW�b�ȽuRI_80��a��d�Z���g/���6g�e5Ln��um�Ԉ�-�<�w��cx=�`�g����]\��8���Q�����B��D��Ɣp�Rۣ�;Yk���ZB��j�ʞ��z�4{9G��ߵ����R�U݇$] �]r>7��Iy�	dxm��ҹ`4��C���'���ߩ��T�ߖ�>4p��.ڼ��S(���v9s#Ο�`��>��0� 隣��~��m�%��S�\ZƮ��P�PX����I�ү1f�j]WF�<0K����Q���=4N���0�ð�I+�X���"e��B����ڋ�n�+�8~H+������O)��0:�lKÑb1�m�;�?���v��!? Zg9�ќ�J�o�����e��#m�f�o��S܆�\t$��'� ����p�n���_��[�;!E��^z��Q��s����r��(mK�lmU������5�}	i@@���T�
lF�n]�o�����ȉ��EN�~����<�⚹?���n6!8F(8��_zl$�ծ����$�h���R9�����xv��z�<ΜS4�,yٍxrA](���D����DD(,y�9p)�V� �8@����Lh�M��&������Bw�&J]J��t3���I�� j��a���R�\���>�Mm
 ���E�K��
f�3��%I&9
�;�ze���wRnU�f,�Og�ͳ�\ը<p��U����ePl@�@�H$��%�����")��j{So_���^5ۇ������Vw�����9W��f�^d�Tό����곐�Ȗm2���,*����r�#��h�����kdl��)̜A&XDx�j���{P6�qYq�C�8 �קi�zDc�ɼr2���dCz�B����j��4���?�=8.4�Ʀ�۝��_ѥ�-�*f�k��`��,"��Y�{���/#����&�M�̎�!	��oK@D<�C*���_�*��:��(�ۀH���̂����@��xB'�=7�s�dyߋ�˅[(h}� C+Oe���XM���c�mNՠ���}�ۆ O�J������H�e�E�XNҪi�1�����5�[���D�2FC�\نe��af2gG��'��4"��È�W붹V�ñ?�D�sfOn�S5��[��[kM 
��Q}�]U���||�ӪJwN�9��z1%,��'�����w>x��F�0�>�m�w���+CO���XT��
di�ͤ���Wwf'��9����7�6o)Q�Xͥ/�&�t�7ˉ�e[N{�v<���%�Ald��YEoZ��tY�-3�h�Ż�LE0ϱ<�	B>��:�ޥ����Y̴R���J%���y_�q��i�A���Y�xA񔓪�ȍ�0m�C����d;��;�^��ؽu&X�3��#U�/8�[D%>����s��� 3d��\>�:d\�u��-��^8ʍh�(��^Mx�]�;c�-u�e�-1���#���y͇J�!gd��o��bw��a5��_�����-d򪖶�9��XE�R��BeA�<K���ԅ���C��QZ��^⣇�q�#�w.�@����
��x�f��#݂� ��7% �խK��^�Y��F!NH���p���#Z�;(� �UOwA�!S�h��)f#V.Ɵ�,{j�U����8�����
��t6Q�#Ɠ�7���� ̹�)�c!���x^3�H8(�=����K	T|���s��S���O��Ҡ������X�(_� �Gg�����	��¹�\�'6��\L ��S[i(���^����K�����B[p��/L��%t��6�L��nT�*��l~��G��j�\���<QT�A4'�8��j� 5���-5�����Hޔ=t���A=";퓭��R*�L�_��nV�JY��"�3lv�B1��{��M��j��9��6N���]0.M0bn�Rp.�ӦAsdӯ��a�h^�>�&�P�1ɇE��G.�8�<k�a�s��F"��W������ �X�L�����Cj02����<k_����J�*8Kc��0:��1�,��ۓ�r��Z�G]�]ZE��>�#�mB^���~~�ܝ'�8�k������7P8�?PD�v�e �"��#r���'�"�/�Z���b���E.*�'�)��=T�$:�¹���䶹���ڍc	1T����wU�"�%��% ���S���[I���wNCae>���Uij�C�P�on� k1{.���������~]3hE���	�.����5V�MEN�$�#�cŢa�v\�<%o�{  \��T��ǋ�����a���K%���+4�iˏ�>5�T$��ڧ����5�ܗp9mO�[���#SX���E��;�4+�(�qX�'ܝ<�o� G�jd�/�\d��M�&t͟~:$ !,�7>���^J�_��O�5�wW�v���E�S-��i˹R�Op���ߛJvm�A�/�H�y]�P���T��Ｑ�3֥4����^��'�Y@��� J���m��\�C	�^�.��Z��W?`ճ��q���T�kК�THW��Z�Y;�
� �?3�F�a%�%-	����#,f��ԟ�l3H3K�^��'a:�)�x��7�[kY�@� ��¼q���"&��)�Ŝ����)�vy�j�S���p@6Ć��=��$�և�:j/��Kx�һA�b�,��b��bS��uHG:<����ڽ�e�
|N��4�[A@��Y�R����pa+C�^ad��;���tJ_ZJ�-]��dĘ�G�U^�÷�#=�m�z �)M���c���i�9�^˒H_O��^�ܯ@�Bz�0Ic~~��MyW><�V%��
.۪��g��Ц�b����Ƶ ���_#w.��"ZQ&��;��{�S�Ճ����lG���F�^�"��4�������)/���Q�h��r��LN-�,���`���!��ź��������kiZ��LB���M�~�]�I3$*�k9��=m��ʆ��A龍p�K�v�I�4������]��j�"�g2�{����܈�g螫d;�#_�60#�^����i�P\�D�^�{#�g�2��ptݔ�b&C]����6{a��sJ��f���:�N�z���<Py�c�;��w�i��H�t�!B�O�`���r$��ʵ���ͮ�!�)��`hq���X"q ��A�ݦ��)������T�{5i��uJ�pTr���Or�v�q�Z�h��p�Ts�龳��e������ʊ�Js[2�@��>!p4����a�4��B~aE'�	=a�T2F�����nSw0�#���.pހ���0��Rc���|��P������'QNX�U�h�!�;�����Cлj�d��nR�����(Ky��of�-�Pa�E�o�FD�Mf�rp<�:�z�����]��}�M���D���$�5?�z��:�)8�p��\�^���S�hA��z��\��c"p���k>B�d���?޴ �7��8:��PY,�}��!�?�<���B.O�f�?���;�4��p�M��d�A��	mIh	��c����J�͉��	��r{Rs�BC�1 ۪�h�?�u-��D<�����'~���?f)("��a�VG��!�އ���&Q)Nqo���zi~Ŀ���35�T 0�`e��,&sA�-�Ӏى'�7��M_|jm�O����\�![l��i������~�����f����t�˘�K�eZ����$7A�@ �Ǣ���t	X����O��YX�B�"�P��*-�Y��dc4��1��4��樋�7���r Fia��.��S91���l�h�Z���)E�*���.t��u���Sʙ֟���st�Bp9�985����r����#����f�t��j�#,���\Ud����#q��iH��g\>�Ԭ����i�G�t�?��{�����U��ūcYM����X��ϚtR��u�O�b�I�Ӝ�O-������f�&�`츪Ss%E#�n��&�jƭOQꥏ�Q�4�Ow�ц.{ے�e������0��(5ԿR����G�3�E�'�v�ѱ���=~���� ��i\ k
80:F
K{r��70��5�o�nU������`���Jh �����i�Q[
ZG�zM�bdqW��_�!l��{�[
_�M��5LZ��~�ci���cb����*!7Z��I�w�+ۉb��s+�ܠ�j �>���̰�9� 4�3~�)M6:�.p�EH�Nz�A�%�%@j�ݵ]�m�ǹtAvz�\�l^k²�o�=k(�tw�Aus��b�s$�Z���8U�p�/4_(E:`�or� �+g
ZO�ʲ󰅜�<�5U$&����ƻ	^o���m�z\�7����sk݁�.hӞ��P8������ha���g�Z�[&3�<r��\�d��d����ֶ?�[�N�X��v7(�R��'���[�<(Vi�����?��:���Pw��4텄�O�Z����^�ug0�����-�e9�U���6Z�Zڪ3`��;�M�4Ю��5;�z5i�\��6��oxD���ӥ�Kb���2%[Lҕr`������$87N�lB�������/�1a9;'���Zu��/� �mf_i�Y�J	+�1�-�YP��0�I�m���k��$ݸ� ���)c�H���v�hò9�^�f������h�A=��4���v�>D�E��]T�{���_y+��{���mޝɣFѓ�{%`��T�:��br]}[���HuD4)-9e��Yl��N�`�{%�W�lV��x�[�3�80��Yzb�g��h���u�0�� 	�`Tq ¶��⼑Psk>���=%q����#��"_Y�Y�@�G#�\�z���RL׷�tև9�֘w��Z��V/w�l��$8��-�ys��]��I�
D��h簅|֡�-�;�I�d̦V��`+.S�r[;=�t����*{��3*�J'�L����2��:tks���c��,8 ���ոt����M�-l�Ά�����}6��p��|���4^j��S�[��m�s���"�c�ObWX=7k]�)4S��E��tz��o+�Y%��ʒ
/;	�����p���
'�~�~f����,Z�j��K�#L,gщ]��˶�^�C��R�/�_!����j�G���Hh�e��3U�)�/��bO�e.���kغzO]�	�VHj�"�	�PR�}��=�mv+��v�N�hWP��Ltko���_���H̩U;~�&��q���g��G~�X�G�	=î9�x��&�"�c�R�[Ȼl!�9"�t�ɂ}^��&���xO�dU���u�$��+���C}���-�Mh`�9_R�	��C�~��d�Ad4���3LPp�E�g��5I�r���k����~\��\��oVfzG9xkKb5���a�W}H�11$�&�3���Y\r��6)i���P��S�Ft�����a�S�`5���`���X,��!��9ka���`]v#QB�΃��?6"%)Y��Nl������t��_�����i�YL�,sEku�i��Nk�z܋d7(N+]���������Y�{D�M,�\.���DW���ud �<Z�����d�'`9��0���@��tP��̷0T��9��v�X�Ř�,fG��Z([S��-ý�d�FF�#����:��P�o7"���2���y��'p�����#�+(��JFg��*�QɃ=ɪ[��΁t�f���$�A�N�[�t%6$��,�������o*D�*�	c���_����z!j��n����q��ıL��5�joR<<X�';��5	�򄈞�_AQ|׏�a |s\'���\�t,7������M!�RX�	�*O��OK�C�(��d��?ъ�k�1�Q��$�K��^�8�m��g����u2�sڃ$xa��t�3%7�^�P�a0��wg�bCa��2���xKp�4C�fG�V/�7�$�<���9�4�g��puH��).D�H�o9<+#��ȂpMZe/�dzW�����_�iAm��/Hj�Ym��,#����x�XYmF��X0��Zj�m{��\_��;���k��Bq:B��R͘JN����e���"�l��b	�O7�m�Ap�IA����U;�-Dmn'��/;c`�yޥq��>����Y�����:H�84��X�V���W�LI���`��A{��Ux �X��^���F9��<\�]�C�Ù��\��[1�W!�ζ�Z�M2��l�}	&b,���T��9�,]�����I��\G&,|67��q��%�+)j�<��n���/Y^���7fhM� ��,�WK�����g^��,ߝ�<�m��VQJp~gL2;���i�)���8�B�/H�+�6D ��Д�V&Ipb��J����`������mJ.��|�,� y�F���0ą�rlp6qhP��[
d���	e9	\�68R �XzŞ+.��ϭ�~)4�>�}c<EI3� %�O���&P�`?���t��9��\U�DH?�U���E������ Q���p� -$+]j�I҆�O���\��^-��d�����8߽ΛQ��go�d�.;b��?���,�ab�%�.�ْ.%z��V<�w��I2��[\��rǁ�z��4J�D����i���`��Φ�R�d��������?�f	4f��7�JkgM�5�E�K�1B�lF>�ݰ����p��p�����uO���X��Ca��ɲ��Z~��f+�\~{�8J.R[�);(BQ�od*k���[�ֶw�ac�U5Ue����O�,�2�%�+��QNA�Z�h��*\d�F�J�w{�L�W��:Q�����<��&������2���w�Щ�\��#
����=��c�����G�wemb�B�n|�E�D=����$O\W�ޯX��}h�����`D��RaY6��y=�@���eL���w
�9���M�-��Y���Ӈ���kR�Z�U"	�O�v�6���S�P��8�`�Y$�/��`%o�4*�z���`0A�h(δ��)֗'�vD��*[�.W�V��c��b%�Q�2�L�1.sj:�n��TT�˿C����G��ٴ-�pg�"��b����I�5; �Y,���Ck�W���,ff�.2dӷZM�b�S#oos,Ok��p C/_B�/	����T`����H���Rx}?2��~�C� ��(O��Hɥ�׽�]qEU���ړ �ԁ퓠�8�^�������Rt,�\X��c=˽��wߒ��Xl$$AX��9��|�Fg���g�{cf���\vCWZ
�:uQ]�����"�'j�i�w��c�*v��>>�2��
��W^�>н���|aj�O�;�>�͎���D��qb��{�^R�2^��c�2��w\_|ő���F�$�@}�zU�^����<��='����=O>ꌠ42�):駲ܫe�����b�9�=�)c,�ʸ�|��X���xլ��^�d+��/��桩q���: �[�W. К���슛�����b���ꚏ�dj�=��Fs�+�Sk��*1�?���xOqd� ��U���D���l��K�e�Xj7i���҇�r�=FZ�aw�/�{\^&����	�Ӽ���E9��)痤���*,A�|�i#��z	~0;1j��qA3a�1��\�[��[��w��Y��C�'�7ms�→�9_R
U>�f��&_Qj=ed:G�k#	o���k|ma��v��7"�����2L�g7~�X���J�t/=���)��d��ݣ� �4o/٨�ޢ���vT�E{�����v�;����S�;��>���&*�%�Wg3�ZV�.k�v���u,-{56C/���"��ek�.� g���ć[��Ȍq�vb�[.�+|d�:~e@k�_x9���_���jLt�v�%6w儚��0����DeU��mI�ex2a��Gsِ �z�$�!�	#�ᆺz~��F9Ƥo������C8"Md�Jwo�id�a�\��׃"5	�q,��#��@e��G?��*d�(��W�o���^�?.#	$�P�R��Df���	@J�S��&�-�$rL3�{[�N��2�/�rݓJU�x81���%eY	��b�:����9�TaA�`N�r7D6���[J�`j3m�!�4	��K��\���w3p�uY��d������PN��d�7�U����y�)�.��N�A��==��Td!�s"������
.P� �˂Zr߁��ՌV��9����\���[M���c���4��E+�����j^G#�-���Rn�7U ���3Y��0���^/1%x&�"�3( ��2����Ck!��s��Zq���3�\�01#��䎪5h��v��n�B�-�S7�6�y�ٿ9�51�lS.��<fT�����4�s@�R�1���>Ъ^Z��V�.#i7}P��{� N�qX�����TJ���W,}T�ȷ�1Es�[���9!�_���[��2C4[�L���γ.�o!e��q�l*�~��;~��*�I��wf���ap�W�RȰ���-�o�K�n��
I��E9�gm���Jd�Q�L�m$���U��W�p�Q)�dE�jL �M˙d�,�>�Ql�j�I�@�os/+�p��>=m��#4D&�*�+�{vX�䴴��i=by�c���k���3�9�;]\Re�J�tn��W�㧸�z�4��t���E[v67��_W��2�߰�|b��\ɹ���m.k92YU�:��ߺ��]I��+�k�'C)����ႉ����_��j����x����oJ�_`�@K�0�PrJ�&FJz��)[�P��,��溊5�=]�s{,�_��P*K0��x��SM�A����+}|�.���8|�S\�\5}��!2��e�Q�|�ē����c�I��m����
V� P-'���	.��(�6y[�����1#h:j��1���h��p�6r���:qa߸�%6�
��Fbك��L(��	ӛ|�u���������Z^@�t���N�?̔�n�%�R�2B*o�W^чn<�����g�p���Te`�1֙޽�S�h��џ�]�XuG|��Յ��Կd�ȏ� 0~�ޠM3 nO��_���_�d����}Ш�`-l�Q[�����\�&�^��xv�J,��]�7�ٮߩ�l�Z��A��z�)?FG��a�0FUK�5�U OH{�������a�T�~v`l��� ����;ܠ�$�-x-�u*�ω�`%u2���'@M����O/S3Ʃ��q�˩{��e�w�V.��)��Tw�9[`%	':����\M�_Ѩ�_��{zi{w$7*zЊX�9��j�"���c1w��ۓ����4Tmy�o9���cf\,�|����	zjF�����VC<wf�JnY�]��ƀR@Y�@j�{�1[���K�CG�Yb�3�Ç��L�B��_y�������ױ�']@�>{H�e�m�oc�����j��m"5��1z��p�i�Y'����1'%�4UO�q�$	�Mص"�(�(.��l��H��Y, A`S�-���1���%��_����{�����]:�[ߪ"G��>�m{$�q�5׽.z�U!Т,p	%@ .2�T��m�X�y[�d(@��4�J$�sβH�OT�b�����3t�R�Ñn�9W�(�|��9W�F�N������|
0G݆���H�g��ע�E�ݖ��7IA�{�ol�`��^�Q1��@N�B�F@^w�ެ�V��o;?d�8P>�n�u��'<W'}fy\G��������!z��B��gL���=��t�gvxut�CX*��wB4��f��*_Y�P$Pں"6����
kI2�@Q:�P��Ɏ�NB6��e7p���K�P��M��tqVP4�3m13�<g=����r����d=��u"�io��[ف�oj�&ۿ4�tY�8����d�Y��8ʡ<����2MPa�Y�a��c�"��
^��c���,70x�a��~?vő���&y�dx
�u���7ÒD*�ʎ�g�IyUG�x�� 5S�oT9g�̠�q=�UR�������a]����vu5��4�]ڄ�H%��_���	P��t/(1�M&+���F~��E���4�DK��ى����Pu(l���0	��k"��QBG�^�_���!�@�2�$�:�/gb9�71��sg< ��箏�sU*����h|�Q�:L
0dd2�>��<^�@#��~Y�7��9�4��3����)�����jg��Q)���u=L�æޮ��ˮ��7P?m���S�u�n�Ҋ���M���
��NqRM@^Ld��ˋ�=.�~@7Zr�a6������u3��$�����K�Ri�(N�X�d�Y,�j�"�<®��P�e��i�Ŷ�Na�C�I��k�pr�ϧ?|�|vvb���_�N��J\ϡ�i��m�YW%�_�*lѾ�Dp��߃��=�*�Đ�^@�[�j�����^;(��H�n9f/�$ft�^ڗ�����)R�7r	����}�U��h��������՘5S���_,����j�l�f  �o8��r�� ��Nx�H(*C���?��D��؆;MD�;ѸRZ#����J�L˪�^�<k����nR"xdEF������ކ��C���{\�Ȝ�H�f�(��XP̒��D߶�wÌx��-�8!~X�����q{3� <	n�1M('[�����%�8�����,Q*p�_�`��^����q�X���\����lM��`T���B���f���c(�:���T�.��]�2:E��N��o���)�2�� ���!ʦXB�������?�]âi�H�ΖS�
�|*�VùG�r�.<�rOevR�5~��~�J�j/t�P���� �l��X��ݨۈ�d� m�P����� T�!j��3a�b�Rkeq.+���@�Cэ3eL��fR6؟:yÖLv4Kx���l���1o��>����[}�ި9. F�Q	��^��٘M{�슊;�� ��>Z��\C��!��yM".�mq��dn�?�(�՛�K�$�'�>�?H�$�92㽽���8\g�u�] :��Ҙ�k�|L)�O
���/�KK؟�Q�����������B�܀V�%-+�v?8�JՀwܞ��{;!��߱�s���4�A������8��*���1lB�45��뱯t.\�~�z�e�6����f�W�m	��!�)T+еc�2�[�K���q�Q�+B�w�(�ۋF{��h� ���&.5|���8��X�\�D1��!��C@�U8X�h�BǸ:�e�f�e�*�R,�u�K���~�*I*KJqSl BI�!=
���}�y�� i�,��t�E`��S�,����i �	8�M�BVk9��5�ƿ4��W��O���/�m�q�<���v%l���9�(��x(�q�H�B%���Z/�]rg��\�ƆC�K�:/6!y�� ��+0����>CDt�_�n��w��(���!S">�[.,�k�O����E9�D�g<��Ǆ&ˉ{��)z ���6���ٵ%��zh1m/7���ա�3�\L�ݝƌ�Uk�:g]�8D��Pł��\G3ʘW�U�����������ud}�y���,8�*�L)օ�`ٟ���{�0xu����]��C����To�L͊��(;������Phf���b<rs5�aPs;[�!�*t�|�͌�?ŀ�L��\�P�a�On��+��j3�>�rz�	�=�d�H��%0}����e;�d�Wo�Ùs��-���3[6�.俲o0Pz�?�����/䭷k��ysެ��g�t��\�sW4�h�u ���z���o �p��wk��w�V�LyB�16��Q�Bqzz��K*ʑN�O�%�C�K�>_��,�Xh�DX�6J�O6[^���$���y��V�p�v����ŦD��yS�n@�b󣴍3e�HCD���I��t��U��[ׁ ؄!���fl���ma%����iA�x�	��=�?���*�<Չ�k�φٲ�:����.p/"������A�3ݜ�ќ���3�RJ�m����ěܰé�ڛϨ4y���\��p����n�i}2o�o�<e<�>��-�TXQ���Jo���%Uo�m�	(���R�ø2�*�`��{$_A#I꜇�&%x�T�#e��	�k#ĖQ)<�B3/1A��Zl��i)�N��e�ȑ��e�
�,l�c�T����TLr����U�ܹ��D�M����P��8�-��{Ɣ"���=F���PC�sld�G_&���1�ib<�{	9��)Қw��^�7�{Qj.�uЮ��7��e��Y���t������Ñ�@��O��p2�~UST�^�M�ۡ���ū���.�I�֖�ڨH�j1
t��[�Y�Y�;;���kÊ�����*�$ N�UnSИ#��B��tK�+ ���}�³�ڂ�	yJA |+�Q�4JIQ�>$��B��;�|�B�3o�]�k�0�h�P���M�4�[ (�!�Ÿ��TK�&$&B	U��dzv�YL���~ëa8l�hb�Tز�Z�]�#7���p������b�2��Ht4�W}�W?vPOo��V]U�-�����3�Q��O�r��1 �F��~���;o={�G'�_;�7����Vƅt�Z�A�)���]�me�H��Ă����#gmOӪM��v�K���6��v����U���=�(���e��Զ��t0�w"��*��"7�;�I��iΥ9|��� a�NP���P!4ٝ�JVfҪ\GB�����xX�=c�Uý�M��W��F�ghv�^�9y������ܢ]:�J_���cB,��0�\��
xΏ;N�=~V�تK�%q����'�f)#�#��P��e>�ho@��t���^15���P��H���Z�"���r�*��d1fI�7�9bh�Ύ��x-d~dtG��J�^���_��/Px��K�X ��{"�7_�#�D�y����ڠ�6��8�U���.y;��'�ׂK�@
����;+��1*�����
�}���#�j/�T��U)��2����YS�P��e�x��Z)$'��`��Z�n��O4����XY�D�ۨsFf�9G�������'�,����Nӹm�
�f����2�D��������Q��.D���~�u�],KY��uOtOB|���O�.�?�x��tI��u쵭?��e�R9}��f��="`|g�D���RA�Y1E�r #�4-�AM�>E��%h��@�ˮH�RV���w �C�;�Ws�#�,z�έ�X�a[�pLGP��7�D;37=&�y�+p�N5�Jv�c�\��HqXY��o�?��ֈ%�5n:S���m|wEuA�	��M8����M����.o%|�ٵR�����|Trw1�4�?p 8�JM箣/���x�B�x�*�r	��`$(���b�Xi	�yy�����$c�Z�L  |Ϧ|9����tY_���uo��o���,�-~EE���&n��]�=�v�Ȣk1�O��yGŘ��n���:��D�3gR���Z����Q��_��N�&�זz?���'�P���+�D��)7޾��ʕ�39������^�Gl�}�M	Z���خ<ܮ|���R�v����f�@�0����^7M�*�5�'���R2�i���ݘ�N�>̅e�����n��M8>&^
]X6��"H^r*��UGN���P*E�O�ǹ_G��y�A���g<�Ǒ��'���5ւ�^�.�e�~i˻���;��k ��xޒ�����9+�O��AV��I�4��S)��^�W��۲v^$��0���
]A�C�ĺ^���gipiO��{��RJr�A���
��V�S�w�5���9��?�(�+�����N5@���qҁK�<^��LT�1������A+!�mI��$�N���r��.-&:W,�k�)8mXfu>�8�"��4M��Oe����|��B�J��	�v(�c
WS�)H��k�Y���U&�����fR�WC�A�����-�!M�#���WΰP�jl�J���MV��T�i�0Ҕ���נ�Dw�?(F'��\#�	|����ͅk�\��&��8Z�1x\��SDc�v�Cb����䢉�^,U@��I���w�z���L�������t�m���0+�j;�֗���������Q��|�^���.�B��+W��
r��Ct"c�tzr5��#7kaɛ���Y������){�w�Ɓ�dٗ�m:�?�7o;�� A�˃�"E���6\|#c�Cזs?�`^�_����"��*�ak2r�l�W.�m`�E�C����:�v��Y[���NT�2Z���wi�q~V���'dJ[y�n0|�d�ְ��D��e��#�>L�T�!U��� �s��R2���k8	��Ӱ��uV�hT�]������Z�F���z�O�J��`:ک� ��߸�G�2b�O�[25�jI�I���v�I#�V"o�l�{�R��ʆ�|B31Ul6��֍��
 7��.�����F�Ѧ)&!{�@�ۋ��\�N�U��m@��;��!
��gƶN �W�}(�&��p1�ht9fi��j��ח�Jʖ�v����e�� Ԥ�÷$*L]���~�:3Þ�~3n��S��(�y��6����}$L�j9�{I8�4|����ǪH��7.==j�NΑ��:O"e��t��o8��S �I) ��E���|s=���&	�y��v���E����wL֞�ʣ�Z��&��Hq'O%��
�.O�*#ɋQH��CdvQ�9n&���R[�j��9�g�ᒥ�<CJ���AU)���Sv��ap#hQ�s1��>�2t���&�z��2�܎X���QŶ8B/fE��	�Z,�*�/8?|.�?���Ҧ�p�L��o�V�b��33�.z�v�b�C6�Ps�"g�kվ!lIg^S�4���Ws���\C�X�G��Z�B�(�`���h	��M�I[�U��o���6�@p��7�4�Z�n�+�����~�H�_4��"�Dv#�ұ��SS�.q�y�ʞR�-������u���<yс��4�]>����(�h��6��'k�<��tܳ@�J���Z$����w�15l�o���'k�a4D�m�42��]�h0AA�B�"t��"�� �Դ,رv�;�m}Y��+u,�Y�l�w�v�dni����t	�+>���#����
1���k4��]�vt�K�k�uU�-��E�n�3��S�<*��ޡ��&���\z�3��_"����<��b,Q�'|q�Րi3�4�����e�^=?>E�ȳ-�������R��O5V4~e{o�L��
(A�`*�*�����5D9�}�H1p]���.ʵlZ3Ǭ�U�"���IϰD��#�=�"T��K������ZsHU�	�7�s@���k�M�<�4��IGngp����p7��a���k�&V� V�C���B�u�&�ZB����E�����ޖ�+�F�VKQ��Zi��h;Je�Kz���`�l݌���4� ����m��1H�A��r/�}К�J���8�~-��}2c+\%,L;�..�3���ۮ6�֒�i�
�?�
��$�nZ�������!����������P���z���vb}J/ˏ�J�]G[�L; ] 
s�E�������@0P]ʌ�&i�3���(8��q����fz8W�@@o�6��Ms���Xe�`�9��ލ�̟��%�BC�u�oS��d���A�+�S�����}G*D��jv>�Uhp}1���{��be��G����d�f��~O%Q�:,7��I�4b�L��B[U�<��-w�O����ѩ�Ar@}]p��EZ�o���̣��e���	��=�ƪ�����~�������ٲ�BX��ͫF�c��я`#�FYi}�_�Q������VD��"��ޟU��Xԗ�_�S���)���j��+����a��0���އtmƆ߉�Z�؍�J�f~�`wy��w�ҳ�3�,U&���+� E#��2���2���@K+j̽Q���h�t~[�t�x�i� ����}C�Z6ZB�����C�QJ�\>��G^����)�0�s�Ay�8_X���9Q0<�\V�S:/�Nug�.c��; w����5��I���6O۟�Z�|g� x�8��?�G�0T�E��@x9ŬnX�]P�v�<���X-��e��(�H6��g`ʃ�����eN'+�~w��$̦�������/$e堗�t�����׃���#	4RдZ\�&�/�8���߹ܪ�5:�u�MƭAn~�K`@`�{�����N@��f�H���$y�T���Q�H��fӓ�j�8���>�jKv.�Q��s��|�W����CD8`nj���Q�n�(���PZ�n�PJ����s>�Or	!�7���������1���"��D|��U��$`}X�P�����c4�#-e������~����w1U��vLD �?ZJ��b%��Q$��<0J�p
�C/u�����ׂ���� Q�)NBw�5���P�z�7�3�
|���)}qXXg�钓��`~�T:�$#ʬ�Ç��NW���u�����~�Ը4�m)�ƶ�ߴO�����������u����"�����7�&�~���B
c�~����0��=��x)���<�Z�� ��˿��3��U�;�]|J`svP�l��,��Τ�'yR��a�����A綊x��]ˆd�{�V�2��Wμ����`hP�˨�7�Ἓ[E�	�Y_���
�͹$(m�m{�	��r/3l�$�Z܃�2Y�(<3_�����̠dQ���;���n���u�Y�B"II+$���ņR����-O��~- ~��*�+��۽�RQ�b�"�
��&9וi[T��p6�*�@�4F��TU��o�a'x�!)ʶP��	�/�Kp=��_����n�i�{�c큡d����!�琢fAә/5�7�����(�hȯ���<K;:���pI{�N;;���q��`<*�d"8N(�������*O�D����c�$�t��
@�H^�o$���L��6'�S�dЖ&/@�BG��F@	��Mvjš� �Xf���a���g�A�A��5� �VI���ª�}�3�ʀ��K~Cx�����U�jZ
�~ P�J"���G�OF\��>S.]��lb*���H���k⒬V]fC���Q�C�)�gkCrQ�R��i��g��/��5����$���)8M1X��$���O Sa��׾��vK9��, L�9�%F}���ؒ��`�S@U��"1��z}����b� �����\~8����������w��oM�՞W�&���g�H�OA	L��;���I>��-�X��{������4�91YGYҨ���I)@��8!NB������j`9%�`t�8ŔN��7l���aW�*2�,˱l��%	ᎂ���l�!���{io�a/caq�N_i����~�*
�,$����
��y�A�G�sw�3V��Q�Q+G
)�Uc��=� DM	�3��=������tǻ��
�2�D[����<0��ȯ�:-�"_��ƭhyC*N��2��%������iS,�#���bP�5�]�����zogO�v��О����t���#���%��9�7{<@�)���gkf�Z�9�����yF�����~�#cy1<�ٔ4d��ȝ��$(U���5� 㓟�ޥ�$�t�֎L\x�yP��kDUtQ�gFrzc]I%NtA�Y�s���
����|}~��X`�&����#�<�����ll)�m��Bb����(x�Y���ؗǅ��J�N'�=�;ˆ�Sh��;�K)��fj⃈6e����$(\���v��"�ȟ��OH��3K�ez5Z���NUȀ2�ږ�nY��R�j��9��#�!���'��h\4�4t��#�����
�**� ��j��9��wX��`.)Mf&M�7��Pǆ�]b��m�	]���n$F��!y��5��s��b/�*��cX B%ƷJ��S�g����Q���B�<��5R�,��u���B�����8�5a]��Y�0�g� �Y�����6�w�w��`G�@ƽmS����;�H��9�2bh�F��`@d�8�LD�J��B���V*�k�z�L��
n��~�U�`KS)gӎq�<>=�Z m�׏Gd���P��bFE396�bEZ����6ܐJ6��#�<�0��"1C]�Q$���x���f�+�@���@�=B�aV�T��A��A?�Wc+�x�K��x���yNf���SLo���|B�|�����M8*���v!���HA'�6�ə6r�-��zIE�4�S�24���iV�U4#�(��[�َb ��r�\	~��o�c���v�����G3N,O^V��9�B;��l���O���T���^r�(����?��'g��1*�ٺi"�^}������8�B+6"`������#4�~̆ߡ�-E����4��a�>ro�rF���O;�v�p�'jIBd�t1Q-����R�
����S2k�tk��y���=x_`�$�+j․<�a���=R���_*�^0ˢk!Z��W����@����._�8�"	��� �u���w��O���<	;Kŵ͞/�i/�{�*ĝ�	Z �z���}�Y�Z��8e���C�+5Oj�rB�o��צ��D���b%bX/�塱b:ہ�k�/�1ǩ]s)����W��!.�}�اd���qߝ�՛݂�����T�i`߆v�~��x�0��s���q���*�M��'����g�_o��ޖC�Ȉe9��iKO�� ��:���eX���-]�8�7k���ѳ���=Ǐm��,��Ȧ����J���E��,g��H�J�s�\� �⠔ꧢ!.��_��Օ��v��A\Cw�c�NG�,��*��X��ਤ���81;o�w��Ǭ|�צs���"�.���W��P���Ϝ!�J#/�?�@�N��������(F���o���ۤey{jf��,5�lh�q�?j�@�Ϙ��D���[%A��)�$`��W�S�رW�����W)�:C5Y���ѡ�.=�4�.��H�䌚	
?����6��{I�d�����{A���[�Kl�y���n��.�$ɕuؘ�����g���-d��\�H��΄@�����W�Y�޸�R��K+=�����ġ�����y%LM��e�u����8>���f0p6	+�yZ+�̓Y��(N�B(�W�;+����L'2�׋�b�/�E֛��C+�Ԗ�+m�|�ī}�c=
1���>�
X|����������~�8i�AU����6�IT��9�!��A\v���(S�i�IA���`Ô���=��	y�iz}R�;�\��hm'+݂�o1e#^�&�g?��7A���	w��z-.A�e1r}���5���p�)�Gp9Z?�q���1S`�rqћ�F�`�P��u�*g�ó�g��$T�.d�ڊ��Ro��	C�}��+���` ċ|�*B-��R?^]`n8�\%�Hq#��lA��B��CL�Q�k͜q�st��c��JSu�ד�y����ᆬ]����s�<��9�4��$[����%�@��ނ5���|'$��_P�[����~�Ķ2TƠғQ ���IV�^?����%�~W�k�V�WM�#i�d�k�2�΁h����R� �P1$��Z�:l0ŪxSN��iQ�;�%�;�2����~�W�m=�=U/7�QZ�
ri8�.2��N��~�|��.y���[0���3����d2�"7�Ei�9��7�p�hU�(=0�E���ņ���C�QuD|�.�#����g����T��-�'��xU�����-�+���w������:�~'d�=
���S^?��HS+Us�ց)榿V�G��VO�% �UCf@Nn�pU�r��*�,3%�!�v��b��ybۖ�bøhmڂ�[��������]4�k2e�<Ϝ'��[x����f6ۭO����G�pd�з@�(��!- ChJ+b��̀8��+~U�nE�~E�w��x�&��0zc�k��U�f1�|ogY���Jg�8j�]b� o�fZ��'V�dT+V�QNkH� C_����ܽ���Ĉ�A�E^^�A	�Wr^�׆@8�!Z���eR�����;Yw �bx�2-z���I��v�p���W�ʴ`��y�[_�l�WH/_Bl�lmL��
9I�Fr�+3{O�b���XC�e��}}� 5����?:��W\�*0l�yڮ���Y�${�%Nve�Z�q ��(��3��
ʂ\���e��<�=�+��}�J\�#�$pB�Z��l̲���7�O@A2S�;7b5x�s W!TMj���l��i9��C�m�4�I��+�h]�U�_�`�[������s�)!�vf�6�8��j{�<u�	װ�z��p@�F�uH�̫��N�Ӵ4���^�"���H|4#w��7Ѹ`ސ�WN[;�&�S�UY{���[^���&v�2kٸGI��-���X@B]�����#0 �ws��m5����Gϧ��p�K(���\���"\��?�j���ʑ�m� GV��ʒ�w{����]g�<N�6�w�=��h�[C�A��1��+fP�d���үf�S�����Jt����K��E��o��Pc�V�a�++�3�����`�^1���u	���{J6�y����'����C�A���gu�'x�\R��g��;AL��OM������p2~��� ������1�~ɞm�����*vb�[뮑�3�U���R�8"M�?	��o�&�]��ε�������Ϸ^;�}�m߈M���-����d�*_����؊��k.��b�����ufPJ�扊S�eb�!P�x�[��bE��H��j �Ew[\7�������h��y�Q1�-GH�C�f��y����R�L��T�;��������m�ބ��ex�;i%d�2F������z�y{�iL)v��iદ��X��t`8�0�(s�^ �|,A�g\F�)ge�zܴꛑ�r�C��C��Nx >���16>"ӓ]J^�^^�M�VNS-m� ����4r�n�lޚ!��<Ԛ��1�T<�
R�lҦ!��_.�*�o�2��4=�FY
�,Vg{g+­9�3��-�-�䔒�y~��i��}=��o��5W��BB�+�%;�X)�It���vo&�}���;�s��f"6I��3�������(��uqp��#���z˘�P�3~�c����y�0mpç��2���_�,���:p��ez7�������r�Q/��i�RȪ��(%lM�]��E�lu��|V1:�g���Am�g�������v�s(չ˲O��"/���3�c?�0��CS�lA]qD���H[]��/�H�g���m�5"iK�=tv7J]�zح���D�����7�ബ��:��W�4�͑/D��#�a{xS_X�#���ʜ|���tT�i��ϊ�`��߈Ѥa�(���=hKi< �y&�YL����(p�mh&4�1���;�>��Y�
���ON��1��?� �nf:�DOb��!%��`�K�.m�-ђ+8�7H�T��?Wr�f�3�@27u1�~��<���ԛ�#��K�y������G��Qțsӫ�+����x�C�YަcW��qSd�6���om���e��+��r��G���K�M˃#Z�/4P� _�j3=N6A�}k�����/�G��)��hD�:��09ʩ6��*,ZG�A��V�zd�sT��j����b�X�1��npt"bȋ�o�<pzZ��O���oB��ń�#�!�Pܠ�*�����ꕟ�r� c��AW��Z3����Pl�y �����g���r����0�܎��!���}�<_צ�'w�~�Y!��|�Cw�@B&���{��'G	�N��6�n&�d���n�{Z�jJ̾]�dOl�:ν�>�,�Q��V�-�#E�ؚ̩����KbD{�ϓk_��|�0��b���|��rv���Dm��[iI�s��+����fTK�r�2�	����?v�C�
�;���#�=��=5+'�i�p<K�TV[����j��Z�M��s͞��#v�Y_��Ogꐇxp��I(��8S��b�f�UԺA}BVx%#� �p���eH���(�Q��Q�+������H���#QqR��q��1��@����I��B2��L%Z+�+dj d�&�ΞٔF��j);P{k��.�����t�wdW��^�˃�X�綹׵,2=�˺¤�V[{�V7Uz�P�z� �����fQd�?�Ⱇ"�L���)����lŘn�H}�1s΍��M�cI8�^�!c�����Ou��Iz2,f��W#�w�T������0N�d��%p���v��za�	�|���e�j�3�[����y���eY��ہ�8��O���s���n�x�D��p=t-�U8�vc�/�[����z��C���;�]�`��<�B��-�����OM�4�7���f�˟z=�m"-0�W�+ZKH5�೮Xz�o֯vf����*Zg��yy[>�z?-�v	9�1Z-��������d���#L,��;"��YV��D���V98���j��׀׭� ���(�KՔ|D�5{�펢�bH>���xM䗩��B�9�ǒ�����I酂r��'"�:bmW�X��hf��C�����A�'���|��QX&ṽ�>X�YZR?���AS�
Mz����H!�3��N��ЂQ^JR	(�Z���Ӕ��u�C��s��d(��J{��	2h�)����w�*�S�V��v�R��^��~R�JS7�l�
{ y��ɻ�R��F�
��O=���(����	S�N�>[����t���b_����-���"qu��h��0�'9z�r�U�'Q��+J�8 I���C	�>��0#��w��-���"�]
qn�ϯ�8=<�|ZT�xy4KkJ�j���Ĝ���T�>Aw����(	