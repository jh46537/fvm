// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:34 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tCULMCvhssbmiRZj7fYU/E5p8FOG1Cng5Lz05sd8+HTGLXV0ED5o7foNRAG8Ptff
7szsB4Ok5QL3FdJc84a1CRRglfzOqVqqko/aCqHpOSSbRUISiEORiGj2Gjo6r1fv
wAqiN95QSlkYQACGLnXOxBeiHE7fdrtc8L9liCgy+/0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11680)
Mv9vrylipPP6gIXleQKd1MI22WSebmWlCR3EhqkfQRFAneU0ljitme98CWRTfmf6
Hc031azy1onKlbjChhJoKlv2w0vL1LP5zXO90jfkCZ7spVee8EDylZscj3GRcJQr
UY0YWyKsVbQeTZ+JWOVQIQuHTWW9Us8wNx06zxXJVO0P9bhKR7MRrYrxbiIp6ij2
lp/HN0GYDN9nyaTIXzITdFiHgivx06/UFvEstXJsiFATfOJ99yJr41dk36S/+LgJ
twbzRuJJNUuVQx/igTUFdsGPknphjDuNqf0S1icN72rfeUX5cnDkbTbu5MHv6Cpf
FSMlveei04u5Dxy7U4PNZwU1ugP+AJKZ7Yvuya3UMFna+3ktDWgJoMqQRffQQRrU
sbDAG+bo9PXZrFKyLjHA0GgnqYjeMQmkIkN0uPEdTyp6q1ijLVSPB8iSnfg63jjQ
ta/0TQG48x9x3fplc3CuxC8GSOJqwmbul1MeGVykKUuU1tDm2kdz4yFsKI3owXhD
1TzAW10pGB4SPr4MvpJtsWPhXYy0nJdcIBWeQcBpAVHbPAdntdqFkXdS5umzam3W
TCsH/ddXIXgCSLc8LhzkT1twhec9flnObKl2sRbWE7SwieQzPZET9mJbrp7qFmcl
s9AauniAfNTgjczapLrxZPCmS4PtjzBOY2Pg8wMzAE9C35QKeQvxEQNWdGhMbRRX
GAiBS+1aN9g0LmPgpZ0eNij4ntNWNo2HxgeEAPXDs/py8/2LrRINVCeHYtp0Zc6k
wWreNf0CwSlHddgbCbJArEuvZHs9coA4zqCWrO5YBwYESWaYMzkmjHtOWOf8QLXu
OT38ehwlFJ6r8cxkbhhJRxv8w1dEGZuA1vXwUDpxQG8u3iffUVWhm0j5qhLoLJpg
P0FW3P6Qd6t0vAy2OxPcCtUVCIdvduJ5DiCtoZUlm2zTjkHCmGRYdee8FdeSz4z5
tfHMgs5IdLrSZK1W+M518UThnms5Vz23Rr9oeA6DNW2s+wkINwFmoyPUH+F5kZD/
g5eryoMjpaYhqW4/Ep2lIhr7oZO2s/5C50WReFdcGVC15cFUJGiSQzVjmwYwk5aD
icHTfVr5dNUfsaDIl/v2CrCKE7iP9aO8lbGxIvYIYwSP77A38fHvIRK45oikLh0p
P04MckYWwWN5kce2nF9NpnkodGJf6czAhuvnWhcAo3DyCz778cAMM0qjXOqKN57C
GiR2689cDNGjV4JwE47SR4w2/JX+UQrIREXmmP2L2pP1W/Sawy5TmxlHVpef2kIB
rLOvR4VqnS0AVX/au2BJz8Fl+eh78dar2Pb5PXtKioItetIq2b5lWo6LNTGngiYj
6rINJ/JxGTCKzJRePK044Vy4oGoHzTE9EPbk1bswSWmeJUPvj4D1Gk1IUs4P5GL5
JmeKRROcGzyZoqw3PkYRJMdS9oOd/oy1v1z4hcHX+N1w9mwu8md5F1Qv+MeVF4co
Eov+PnptZAsmgBzBNYe/84ONe6/b75gzrhWJevnF/ykRTnP3Dm5HsQIpNtGPk1pR
lDpgPB6L8Jy6Du7U+ZVJXp9CiJNmk9aGxiLuqHw/cLwIjBIYbcWToZ9jmqfL+Hxv
b6Zx/uaPhpOdHxHhiVyqnDAEFOdpOpS3+KcIqDBGQMKR9XedPaHyW1Qcy6B9IUox
41apZi13De8rnNBOsdTF2ZABhWbmOq/zWzqbO5hr9ViaYX58gG2vdcv5tYOgcSFS
EJHHUMHAP5svP1PavoGeDK6VgnSHtpNZOsIkniPHFSJiqDjFWvige+WAYcZ0Mj0D
GAfPfd0Q3pryOdFq7Um9NaSxjdMnrXBIDMOeyUsHxiYGwBxXjdww3S8Wk0Xw0pa/
p3lt/lH+tUDD6CV81C6xVRgqL/zBeYHiNgfbjgRYaR1DpaBp7kDiqEnER+RveCux
ijMrWjwb7GWEdfdui3smYj8vEWayM7qILDDvhHRNwa7nHiNnhsEo07bjb5/hU2PO
mHkHgetkuor+4uirOgZkiuJMx7/dCiW4WwQROeX0icljB/drlNLzYYu/Yi3Czzax
wSQKKlwt6JFGHQ9U8HD6rnxrakVcgBngZuQuVDwv1psi7ENG5F/cFVD6z2cYNR7v
Fo22XKypCWCM57OpZXJnr56pwCQ+eJc4mUlVL/pcrKAekoBQsdOZOu6rM+ZB3IGR
j9pqzr5XNlfXBGba+0pF/D0XVrwAV+5bs2+9wazQoGDh6hS3hSLrPUilI3lwZzf7
PiLpqrYj3Ewm1sI8b8wj49C8BaJdktJJP5QRbzUb4X2xrHmue4rlaGsGbzyPcpBI
p206jB4yoQan6iJFQxO6C/ENKj1RZvSwOH2IMZeV7ez98uNm9Zfx0qFHDk32IuyE
/zrYJ87C7QTCFoBEtV766iN1fVTSNnfQBvxMUAGXTKEepprtD1daWUf2QTDFHVRs
/RRodo9kmiQ+wAZ9IujStMfpakf9PKsuUKxbN2ip/mKXb1nxj6rir2eJDWAhUzSq
2WmDcXm55Wb4ka133SL1GzSfwjnBjEu0WReoctxRFj3UuWoQnOrmINZsy8lvSBWg
tmNhuf5uT9cF72NRvIPuZsOqDCYIuRietOubiJlrcUb6xSJQ7Sf3wYGS++n5ENsS
y36qLbqscx0aKRLzFAUTUdWYKmSv4aQujnLoI4rFLq/ur9/BVsOkIO1Dl4A58E3l
6zO3PGd4wFv7d2WxIsVwQde1suVLMYPF2Igup0p8trf+rREJ9uQAenEjV+yA1pfz
Y7uGl8HNtuo/pSONdlr74AOaH/inrtGbRJ8RRoyAo/gxHAZKvLzW8y9IptnIGYNt
IBJN1WsI0VqA+kOLzPlTMRAN0AkbTIq8w8qPBrAXCGKyC0R3T509IDDSDGB7Nasn
NJ1Aimp9GrK5wdP6ogafNNQ/kcn8Kpgj3ID1LzTWowceTouqJZ/e6UqyiLRawhMs
8aDyNXIsEFKBibFmdESiqmFfDiOdfwXF7b7sshLHCJXxSjL9seQ9pNf0o+h1eRZm
bAzg3H5YF9P/Dy5msthvrbUat2WAQgKKClv7nfRh0TwqtLDphBS4m7LbrCBOfBdZ
v/AXsMnnBO1/FNKbxtgHsZ1iJc57MZCnJea2C3pfsStByEAcpEcNCawrc4Awg0Hs
SpeKb1dmka+w0nmwqbrMfdpWHHqVFDt1u79x/cq3ca6+l8LKIf3Q/85FIg2kGCm/
iXcndhg65B2YL6mWtFy2uya8MiCZs4r+Y18/p8+ocdD1eqGndM9E7yBfMqE1Pbx7
81Zw4TrmK8VgqcBddxpIqLBb2+DnotWgRJd6Dfm9HPXeq3rHhj5q+Lu7TF0g8ndP
9kX+3PUWz4Nav8Yfme5ZyPklol66K9dXlVJGfr47RastIfm1QuCUAdSwBSKjIppk
cJMa+UC7NKgk0i5prUuafSTa4fV2iBua7SQyRCe/ka73GcLru8Sx7PUFTxWRlrYh
mc7UWqy8HcBRXUmBBHzySEfo+5nZmd0gNtk4iwwlf2z6po9C5YnGqnooVQHVq5WN
NHbFk7O+r2f4Gds0b0M0fdx48AszOPeBbMbb4IONoW0Hemwxu/0jjs+rvgnUb+CY
tOIs3SFe4MQkYd6L1nJuxO4JZBSVgokJ8mQRYMLrvrNAFJwjq/fqk6HMs48lGbfM
JijV3dZNv9fFEhTEcWG0JVMfzUxod43EdDRaMVJLw0GnldGF3zJBgUWINFG9NNYO
1O19mlVwpnca3VakWRe/nwDtuG6VcYfOGIZe+gtkfAKfjKv1EySqGiGX7ZR+d6TU
wx64r071rDZAi7nGUgCxYDnJKKIfV1eOP4njEgia5nd2CMuo4mUwUGtfWZmbPtG6
y5Hey06EjQXpjs4Mqsa+aF5LM1d0g0Tu2iYmPMF9ij9F1lOrWRwvWOX56BE9VqAX
sjFnWQkmPXdYiOpbRbtFk791dGZo60IbxgUfqa9BROL5xFOJJ7qK89fAH6Fbgkhw
eo4DJaeDQh0HNmGdGQRzvgNOqfAKBH6t5dz6elgLeTcySMdnOHRpvGbLMK5C7ln3
GGPzkvnuNZNydGZhlBzFDiadpSISu4vCNI43FvGEyITwy3KBNwgX+t06+rkiKgPN
rkodLUG32cT7C1l5wBLcR9Qpb8lKsMAMmmRpc44eRheIdadyDafEpDAeRWujzWfI
DTnPyfas6Rbexn0gOEQlZrafl8E0CsFFEB6fYrSLblSgF2VoDv9eCuwh6wgDVuVB
nylksJ65bfiDACNcwPc0sAPE8rxeaf8l7JnJpehY0UpyzIrzSk1llXiRBL75G2fi
bzDcprtWoxXaXYoIfOwDwixn29yMZjfVhxWNPQcEJES6MmHK/cknP4eYcRN+QP9s
U5/h8R71YX9ber4Ym+pp7GkJOEPH28QD0HgXTliXmvd6kjQtPX9fMCwViOnx9SDD
d766qr/om6Q1tDOh0mqlKc5T45fAnmgCIYdjMbplt0RHN/in/MnV3D21Gt82xWrO
YW5JP8fCGOTiAbqDcuU6gjMzDqmlxXarDDdnacWvdxmrc+eT+FEsRIvD9Gj2oEcZ
+xFti2ywhD1Oe+5GJ7jDLC7TKw3toOYcMC6LZuYA7zNd7k93HYHMCCDb8VgMgOvv
mFmKnLw3d1bEOd5l6WDFO5WXl9Ya8wSFMAzTfZvefcBHX45WLU4gNF1JMreEjOTY
SPpJrh0v5j056b+J2WLeYPjb5Z0F8w+MbVSAznDnx5r/upKdam7An/vB4+Eg+i8Z
J4M884KeULaj2S3Di/TyhqMP+KyJpfpA4ZY/uOYVStQyKQfERlqibwKcMx+jtGk/
Je1X9OM7QUP73YIdtLJhy9ydkn70XTZRVqGM5WqsDNtOP525Oj98lRFik5mMGTpH
EAwS85FYFUNeyIB5eqVqbCFfqkQGNU67KtRQid8wBxKCNyz1W694pBtR5hcfrekJ
36atp8yW9JxumVMmhvrF4A+7N/r6q5/1lx4+g2IqxjhG4b7DTOT8UTqkUU4ZjgKe
mPg+ghSsf/O8h6hSFz9GBtI2334dYJaGbLlUYU1nt5HKrke2JGZmdAeGovDbwo5b
mwHFyfkmxalBPdmgirdYVWv0ZjyAUGI6luCVtkw09g6Rh85WQp9dRlVgYHkMxT0N
g4Icflostq7UVFQCNwg8vdyAY4YsnBZt+On1Nt74F6NJXUny92XT33hM/LUDLtuU
Y+gGa77e7+ryB1ALbXNFG/LA9534CaTmoSpM+vJXSIHnk4I09O07NIqLbhK2NH09
Wa8ylUut6XeXh3gJiAkXpwVRnTO8nu2z7wQacoH9swFoUbVXw7vPKm5jE0KL7yAa
ne5C8sje6pbsQjx93xl1/m3NJPGwZQGvd2ezP1JmYKuBXuCxb/cOWgfpMkldRZCU
g3ZYENvj1KZgEEdmVkcmFiCcQPFNshGivuroko90ITWlOZ6ZIRgXuyXdU4g2FwJS
lumAftr/FP4SqtgWYXu3L3UNwJwN7zvn9kTe0q/koOJ7oRPw52XvDFL95P0WC/mr
zEWgjNkQKM6BMqzCj6/IzZmKAUKMSbin0MgXmCzXGyMBRh2dH3Y9IwILXmeENd0c
snyWhwdV77qCRm0ju+BkMqmE2zJ/stu3aDIRtmQj3cCn/CjdPKYRRhP53SAKwVVW
0awZrOutaLJcNGtmdiQRg6omy8KvhwQb5517uNa7XNMmOVHv0mj0HVeCtooAlPKC
gRLB761XbtycKnd6qtpJOaNHpj+gUTPpyxD9jUwaeGjgPq9N7s2ydjl7lMa7D2xo
6BIq0xfbYlkdG49+bOaevM1JpL4pXBfjUo/CB1Mwy1FMePXYvXRMlaS29QSjp6Af
/tvv2c0/Ty/PX1yBJcSLQlLLas6ftDZHIoUFOD7Dmt88P4Wf5+76cSH7ScgDTdYV
1lwLZvSWitfiNJs3qN5JmpZeKWfuY0mlgO6+3fLRztdFNJEvku7qSFsEdVU/2zsH
akmOhspME/h3jHiBzc2/gL4kw0EaEnNvQ1qorn8kEbOz8qPOv7fFKnaPyWHvKnba
1liFhDsmwwgbsq/T/2rxw/eE6KuN3Drq1819GKxyF/oYISb4sc9Itd/RHddQpM04
6NGt3zJqEtTa9+zIfXF/wHprHSXcFIQJcGwSTm9rwl+7/I5qzC18LGIR1DbhH4Dm
oy31klE2ew6cE+4OFbFeJbQO3wXlam0n+wEjLxvIJYKlVpSZvElM/w2/YYgLxYWh
jwO3hK8QWFbUpAlv6ARs5EwE5MKF6TgcMmCn0AJLDHLUN2hZjguJmNyeIyxv1jrc
ZZBB52fKj45BcPdRli54BnTCVCHPKnA6femVPy7NwtF0Vta49u0zl3OoTPezD0ka
2H3rvSh9Hlu0OirSbE41iPd+8R93fh2cCZ+5lUHij/k9b9sSGIHjLAKHPhGRaJBl
ExOHLEsCK5B/41CdsRbH2UQRi7Xbo7lJ8/l3AZsLaRyTkPFb7EzQ1f7SDARzPuzt
c1OvqATEe7QM3wKtqkE3wy7wzlkeRECVPo9IpLUy2LIPXt6fH629qsjb5k2us/S+
0WjURIZppP6By0eSkqoyhB0NCktJqwhKnDVXeMhSg8BWits5/WP1DV5t2k1b+XzU
QzvW/2SP414TW1dZVdm5QvXyl6LDNGQkv13OZNZtMMhFYLMNZcQa6orgFw8TctzD
ZN3GwAdv125XMYXJ478mLSa5KogbmeU3Kt6iywVA8oiv2ZKl6pw/sAK0Fh0KobRK
KzgKHIcD/6LFzb5nwUAvleiV1H9yTaKNAVn35lHNkDQ6BkPYIKj8sfAyioV2c8cs
VGLJrnbBnym+i6yl4cjWLGIMTJy9q/bUbOdkAYLJpbRuMfYxXWwlUVMwgv+UXgBU
6WsJZkea4eMhBmdRfSnOdxJKz9PUs6fYJMoCJiz2LlGv0odovCkVwp7P/f/oXmYg
Q1ta0U5yOh+NEC/TFBKKGE/aLa+UDo/HNgRyfJAQoEM8rHdKurlaEPNiuTVL62bx
9eNR+oj51d7hS+Q1e1sD/5t77+PXdiBpU1hkcuwosIbnquLvKkK5AvtSgnBs2Jrc
pDTvGdR0M7DT5DKfwBTQjZBsN1nbStjE3L7YO2ior0s2sBDzh3+OoV2VnJSxZn+B
2hknmi8GTqDWZX51GaayWXRIIZP1oiGv9QR9tJoCM9cVt2UdSpdZOGQiXrQGM4V8
zXG4LasYfyDXAQXbkIo2x+lOtTayF84k+0wFaBI7esTIdJmiO6WEYs52HXnImW1v
srizctmgpDQzs99/cFr45EPTTBDxPk0Ot3CSjmCLCNf7bU/NSvxFuLqZ17UlS6sv
b6BsjTU8y5kv/fvnQabyWDrnWSFOGf2ARHD2QKrJYQ9RnmVCsKWpG0sa4CriCnMO
+MMUYOvIYq2m8/Yw//jqLsRtgCcYiSuwNZNSf53rntZa4lSS5HqrAevdHMz4IH5B
/9bGVNnU7HaIq1nKmM9F3VETAEsZSjGwVK5F5sX6RQ1ahR+8CRV0VeEfQ9frhfEt
5MwUSp3shsISxWeZGpfrcW75ew0sIpBs7RHlvz5dmYcvFQ2naIPglDyJwPkk9uYt
IleKN2bQDhsDGZmdIwwfcGa/f2yOn9NTz1+MR6J2mAlvnRiUTvDKqAf3rqr6x3hZ
sD+pN14rGl5lg5nbFr48sw7l2HSmG2eP8o2VIzNmKaLAKPPqGZ27wJSpuyTa9/MO
FbjjLl2xi2IDuxfVVrPLlPTcUyVgI9jru92YJsquLO1AARgSoY3GuaEhVQqU4FJU
Vdo5w7FFzBvM4GdNI4OFHtSiOoeY4npkvHGqI6xzPm3pJTNdW4yO77j7yDVmMX+p
Y+OrHgly839DfyrfmZRH43MiwXQXpuf3UW6TlGSqP9JHlZJAM0xSWT+y9HwDfujz
9Dh1mPhJo0IHx7pjOSCDPUYi2sKgNPKa/TEAQvSvAg+es5StozsGaXUdlCU9zpdF
BkbNhcRJh7LvwkBrCLUGj1gds5h5lin9XOaz0UISqnG+Fxx2iZPw9PTAvWqIEGPr
5fJw011iAFDLMeSv8l1gfOXWgbp8eYUPunY8RNJLvw8ZyJFtiLiLSK6C4gmf9hBO
/ehclyF36axeskSjxDjR7ZylFjRbXT5lae0UHMlAVqOSyS6xDZow9wySzDjrJ634
zifyAZwBsUak42G7Ot/LvBz6YGaN52leq5kQi/FZkk0AoG+vBWcO9DiAmCg41Eai
v/Xko3dgBeG6XUqymbhn5TRRmImCVjcdX49I14JOWYZHEaEU/ozxZyHkax1zRDB9
Yts2tvA0cn03eNk5bnCpjlZmaAsjwgP0DM1Chu/UyDO/ijkBjj3ULW7ZqHwLm0JW
Ht4mFd+A6s6dFcGl8Y0p4h0e/L13MgA6s6ImS+NO15OJJ2mJEwiVaPGvdo1nXh7s
CjtFp8Zy8rukLAQFOazbAPme0OzGUdC6ydzaejf5AyDviP2S3rbBd65yLdRiSRTd
j02ux0hKYSFLMm8/RCM0A7pYgEQ9qMnttFwkJUPVg551XowHy/x2L1MDdMoXQj1H
cxd7l3oPABN4J966oIDFcDZgh8LHX9pML7HC6RcxgalpJn9VAkbdsbqugutBuCy1
sx/SspgRZ4OyoG6VdtTVtXQ4ydqLdzgl6hN2NjABRbsm/ieb8Ot/E+sashGYo45t
ppQKdFQMvsOu2FIXG1XM5q3zD09cjMQVczc1oSYtkjZt0wJpj9e4iB3ZtwxVblHj
pkEovj1gOwgZj4aajr0FijawP3BriTL3iD1O6kJBfPRUJlsbq+9TnEEN3BL1nkBz
D2wYUHULc3f6xBB49bux7pbav9E63yXjlAU9z0lmzHZfQy6Y45kKw+bo/9VBa+GX
VOqMwr2nzT/BOqK8JNHm9b5bj2vFC/7knpBpjf9548/PXzAc/9IoUdecH+n+kxeZ
/ROgE+b0jyk7j6neu65iBdbhLd+YGHZKC+4mzDpZOzIcMsGCkhm5CcHr9LvFpM5p
NfR8+yEdEJ2NmNePFBHZQNJtPjnzwV4N/Q3x2Mu4f28tObG6Gtcn4/vKNjioNkqL
tXcRQmtO7GTe3q/fslnS0jAB+1BV5ewz/VBY7nrIPw/W5Wyhb1Qy27uatzQQzWC5
4ODbdo9hImVexSERAe3AiLk4dNwmfJOy0f04FN+OlIB+Qtast/Pv753WG7m5+p+7
8qoT0z4/zsnxjKpbF7fCqlIdMX35kjLRyqgAdsMgbxDVN1WyZ7bJhsqo+uWV7Cxa
52er6rUW7GocFIp7gPetQeYrDASaZxS97QyjM/OVQXpLPSKORMkwUE3vjadEiUic
NKVihfdOXGHDbmYX1/etNrS01oeFS5cp7PSW0qyLIY86P2aYMaIdlnjcWp9Zz/Cr
rLN9nGv/x27NEF14yuQLmlqhtwb1QMRklxUKeESxxpvIVhP7Mq79eIfUADe3FvVj
pE6iYTkoBM+zVnWYW6WC1std9w/9GtlfGIxE9J8jhjNE4Tzp++fYMYINmiyXq7+N
QEfrJjx97xFxtQD9QkFd/ZvAgdVTBPYUIJ/mFMB378xeDswqWl9FQA7rUKXVLdsL
n6cxX4BCxUzawYKIEdEOhqaaCv7s+T/q0whqNV5YC2ysgku2Otry/T7DTB0O0AbW
L2q0HugSCm92CUXod/xqp28gKkQqH+OSHJOzQzA3QgOYSh4sZkZhdmH4FjGmFCwX
eHHorjXt3OoV2eLdvOfRDRRBBnp7sLHHZQ8qqmcYGpG8HOkkZCGyGJU/rNgYjGnU
pNh+N0TwMZpdibjG3HsAVWGuOdB3PXWrgKNbsFAO7AXfV8OxuMLHeLrZ9fX4wxvU
0tBpbE69S1+Hd7crEAt82fwQ9AK1sKcBZS82wpRxMdPBPPFtn38dFpLGv8ncAhYd
qwbgJKJgps9SEZK/nGHv/NCqfGpQFUjePmrKno+sN7sfuaA5LyihznYMi31Iin0q
eDB+lzKWdB3sMWFwK3o9SSyRvV5AbayWrw5J7GWE/3fA5AYx/1FMqddPOISiYEcH
trwLqNbweb7B37W3rnpW/duF+2aBqDdHa3rYSBN1Nci+c1V9fOms1ZxDOA5WPZEO
fxlNIcURT8VAox3cBqVdwMef371IreNEaAvYKP6UbwzbJApGPxNQ235In2Gnp5UN
uKnSaHQksV0nMuNrFt3+1U2/7aG4QEFSAn4A7FP2BH1xIRp1jf/fzJIapcvoMfPf
keU1EJiGiW6jextK8ENw6WFLZ3mGVIiN3gFrPHPPvkbzDB9vqvDFrlIG0cLc70iW
sRw1ZJc6iDKn65ng06eE1pOCzoE5tCXBHPCgzg4v1or0tJfpZnHz94KtG22/R/WH
xvI4yV//PoTYRqn6QaUe64o7xZ4XL7uHknvmzjoVM7AWEFVG6+TImAKzZqW87+C8
KP/ibz7paVWY/2XuNLfK8JDcAwgUUeqvYFw875wO5hO4PTrkj9SAwF8nIwzlwjzq
uwYtNI99hgWOCvil4W/TfUf3SN5tch+CUZn4aK3BxdP1//wD8RU+K9oRridJ7NG/
jYqXoAn8FNoMe+MU/etyujHgtxiL90HF2obFGQY/GbyIO2dZaoZCgHY9IAGzzEVw
L9FRv1oSB1f70lGYz7g5kAEp5Z9NLT5NMXVWAEGIrL313Jhcjl6osF8UzKy9K6KD
inpSRyb1yA7vGrXd9z7aRR9FFVTWXLc9RxBRXDpVaMX4VDMtPnrvuYMaE/PGI5Qc
0KMBp/3plnDGwPdWULnpKNOF/tfj0bg0JRofB9RsWPYLlS+kg++HdR1BsN+qah3B
k7zPvldR4XpIkrZqoAgLs+B/kCnm2YKDIvHS4tuzyVyOYt1NtG69p7j/1gzHa7Sb
ABJsDe8gRqVABQnOPS3srpl7OOlcieFdNDrpZ8lXIh9g165PxWdQEfjntTnymVcp
JeGOCRpymAPOzrXsSC258CT4pfFHAfyttC/v/7oRSHGJnmGY9I7kd7bLUzKSS66U
/J3fLmjkX8SuW8b90sYdJcrC9X7IfHxcAB+vHiPp8AzBH4HUfVsqsTQ6Sycx8HK4
4mSHSM2i3s07SgYPqfHAS4TeB5Sw06sLrarTevBZjXfw3uJfRZn6t4lBmPtvcadp
6+II7UlFkxcvYhGgR9XaTHcC5/z3I7czwYRyh+pxnlQokQ/DRxujenFeKINhKFRK
mOg0xiNVR9NBDrUsdpPWf1WHbPDV01IJ/11z4W8s/TBxTZKtwPHVzaA9hG7/sb6W
DDwq/HX+LZviyhr6nMyJl10EfGtn1mkwVC8YeAlM+c6pat0cTcWamf0Xmz57XLI0
REBCVt7fZr67QLGhE31hxpgTe4Ep/45pXRj/TgXi9jGV1elfslgCdOJslUCqQrYZ
d9DzmCfhmel8TyA9zM4d2hOGlmisOHgAsb7o4ivlbAF2f6b93IItTzBoHDAexlWB
RjKAchcYkN6FXoPKoejoIipECqL1QRiJHWhLXnz26I9szY5xBbLNCUD9TKfgPAqZ
pAd/U7cNqHrdIotGXptSTIr0ciu/ygzbCoIOAWmC2cQcGjcQkO1abQ/e/+XD23H+
ipOuGkG6mEuBRUmCcfNR1Lc76dPVHo3m+0aafERZ+KmdKYgffRtaJR7buOsgzErn
EqYo5hVSGAYpu/EPElqe1Xg1VajwUdhvYFR9B+aWwZ1ccJQgNwZvQ1b0YFFhmrK5
B3hQLvqbgfY2A24g2APpwcu7S/OsqCaQbhpKgi2FX2nhE2Xd1Q1locPMMKhhOPHt
3aCvv1kD4TEnTDe5rDT2T8WfZyOiZWo0JwEoIZLbFxTNVWcyCAcmcbyjDGZkK+TZ
H5LKmkqclfOV7wWBHTT4/n3oXRavyPcimMeThHuef3hOaobKzE7bbl4POlStLu55
FxA1paYWWfCXt9Lqs5M1CLnjM0VNKDtlqXTi8odLgyJmgjx55jDhnZTl43FUgmj/
ncP/gqZSMtBLllowveojUnhpFH3k2DLWu693/dNy1wfmQRjKP/CnBClAzF/59hXe
5KHSPoOvl2PaeBsGCeRk4a987jVvO9BJJPX3tmhtlvhkg9KUqpzkoxK/hKiswdhT
13Uzywg5JMx92Xb5Jdu5X45oBOXh79BIDRWPblPXpSEnkERPIx2aM0XabcgOW4bo
76Cj36PaQ64jy6Ggn6TX66Hfg8shdlZt2H5rOBYs8N8Gz0T5c+AVMWq6VLcPkgxg
XOaSLIfqVqvTU7z8w9cu37WRFOtDBGrBkrGhN3Xz9arMpAWrSqGUhe5jwNvn3mKp
FFuFqHXysI2gPsFAtq24a7DzGEro0hGA8xcvbH1AyysYe9YrtaKVBvUWChB5HidZ
AgNfGjyKxyf+1yta4TKmrmB3Manr4wZw+4+adwgAVr2pl2nbW+q5UTZ/uE6JHkUV
U8WHyJiTVOfCigPnpWqf9KoxOPbtbILHZEjAvqXZ+vyjwPmHWHGg3OQyd68ChWkD
0kXJMMvR7ggTlzNmiLzA5BaTUkda8v5neYXcJstaSwvMKYWi4MLyf7u8QnYXBp8s
OfWF794CqDre57XHXiDZUPB+nHP4eWLT1oYUnj+EgtXIVweLSfSi1BDGc+L1sdKa
hb9MX+cy2U8KFvW3Q4VqSH9n4G26Z7hSsQ5oPmuv7wn5DWswhntI9RleDORYQ2X8
PmScQlkkhX4AH1ZFVRzJVWroR0mGWNq4layAjRW+zTpCu7l6h6id3AaW8LTaC7Rz
snRjpEexovsC4nqAgLkFj3EgXurc4oEiHYvCfcroYbWajqTMtqtcpTGYfaxxuQff
un4gTj5f+FzryJNQCDhdrSKglmUJCpOYC/YVcbCFokQ3TWJO0lcZskT4IjnORFwc
/hm+4wQq8vOvwMypx3ZmSWVSx/1mRPO47QpeE6jFmH5AiiAlzyj8v1QpQK4+ulUJ
czw/+VAev8SDISMhB9G3Uck7+usxt6CvNZ7Xwx6YMBRqy4qsfSwRmBc9mNVof/JQ
wspDYmguLj/QT0oYyMHG1atmQE5eLsM019HOjKGB1mzGAIIkGOeBIfFREC+RqLdW
DRCHVbbAzM/tye2UNa7AKpDIID1WpKaqnK3EbA5BxI5uqem8q2elWUlVx7xtlhm2
vFquBOVBcHDIFeCIeKfisVRJCBUOvOEOmH4QbUuu3ZBR7qhfyDuqSp5NK1XmVLdQ
v3mkXBWR+gfFkjJ4qlYCjeRhx50GxHaKZiLQRCAiIq2vGT2UuyWdB18QxmaGfA2P
vH6qZFBur1nxPOpdMkj7R2TfsVY414CuiiduuCsoY8W48nUMy4H8eDmswm0Kzip1
sr0/HdoFav/eXHP6rw0Dh/+wEJ4hOFP8RRQ/ZaW2HFPbPXW/Ct7bkmD/DfZFbejg
fzVOQLRsh6xMohknY+k8L5Rlg4E9CQvQWfwzPxYJs3YjCHmrtnKmMP37j8pAIjGs
erv3nVoAeg+Gv84cS50aK+0DVzkp2kuL2iCA7dDfJjxWSmqlNWwziynwUpJ2bjGB
JOWbUPIu8I637NDnvREx/W2Y0kTbhrOtDRa2d91KaezVWCU16TgAaHuJh3jKTPtr
MVLWlLc3F/ok5xRiPZ8op3SzbstFlMoFx83y0FxLR1P02Q0+niF9C4uaQXSXICXn
T46oJIXbRfEMdmtX/zJ7F1NZ9FYFFHg3mMviqzPuwVBzzJo2MVtHP/RPgHtZ+W7G
aKZ62VWgFQWruG/AxBiwFtXy8jTWr0pbuMbAgr2MnikhEr8nGGYW/jY1vAQwBXFj
ccBxBmRkanKtfiSAMckDPCqodQys6TETHncsn4XOW39vjT42ZgbxRsEZRhJugOD+
Jy+zEkHTzvDEui9JPExkIQ3glG9RDYSylsEYLObWQ4FKNcApeBZYcGFXiF5fNdHu
uE/f2tlQ492pp5RlCs6/xinwGrgZNtGxRARs1PnxiqglwYoOJM7qKAwiG0Z/+6ID
+xo6NWjrv6YUgzQ3oqaTHHp2WBzl6pgY8L2Pm5C5FInG7+f3GqRYo5/+5sZiTgIe
ktKy811K2cLmc3hlCtMMhK5TW5B/9wdG7tiXYW7YRXROY7hHlpZjKTWEM+sc9ZOA
WUe6lRuVh2wOtMIctlDniD+/Mc/7mMnSglJsWrxeibI1eiKoPo71M7/1BOsr+Ams
sXseg0B76G4pDzsZfXPAvuEey5f2roSNzsspsZSWQYJPVqvkg1dsa2IfJ1pikhpt
6/AkdxRNegktHp2vM5MJP3usikaO6s528ePP+X3WKEJSHIvCRaxSVz/ssiz+Uk/Q
woGq77Ts1qNEPWaFXpwbElhAgSw/92FE3cPyqoCQT/UdvRmSf6nuYl/5RWuGMXzt
GCZgTGG5aQUCz4U6A86Df9drOjK8uVXpov/kUnAA3wtGh45SvJzShudtrvMiQRzx
USdJQas8xciQ6ZYyXju+eVcKldbYdng1jkPvvLe4nOGcLpHHlBFcJsrMD6Ce+X75
tOYyPwYIzioIKHybQOmazqV1nJCAgBRTOIRyrfRGBpL8nu9vZVZ/XHzI0ZVKSlmV
YLA8FYrZfFcnFbWDJOsOfO0eLUooME7VMbv0AMlfNQwkRb6JgfZDMgAzX5PqPVLJ
94TPdcj2haGIJpjfVKmC1DJQEeauid8qMcUl2rLpecwuxvvFTy4e+rIAc6PFkDXa
nm0n8FUw+JRstr13CWQtAuoFfQ/o//eP3d1uu7defodIjmvT9if6nBHUqCMHvhEw
6U9Jm5q7Stk9SbyGmPddkv5+hnetWyuAX68XwSyMb5Z3PcBbPVD2ztUTs1sJkzg8
I8RZSdcKFYpNV33c88chXk21w1tXmSk+W4l8cdxMI3edoe4P4D6xIc8BzqjFesab
dT8sLjVegpLEsZrj0TFYyVIhUsQe2Pk6ZycXpV8OCEuhz7OnLguUbm4DaF+dOO4D
eIPbNAZS8IsU0orgwMAryNVAtaQfGyh1LmEnoyAxq/lorXIGHy1/YWcodrlp4k01
oWC7h1ujK7fnyT4DyQ1vL1oFS8AVCSu1txblNuAsoxu1NNbhR9d1A6UCJt4u3UUH
cLBlFPyA93DMsf3odeoiGFu+t3iYe7u9/D3ztpbqgM8Pcoyr9EyFj94zTBh62sc9
MiEG/so2tX0wUmo+kbgZxvlFNUnW03mz51R/RtAxrpZFocjReQSbSq+fBIa4GFPy
uPixy0kOj+vKzZBSTZNwt+mrxz/iKqGjvr6mBTcgHILIRbrFXVeDuVCZV7k3CWvy
TJ4WdzRLHUN8cW2om/c6sDu5OdncQ/BMSYjrHvFoUyONhOCpguuPA1+i0rlj85om
UYycOp4Gb3W6rLn0t3eD9HxTEegN9Tt+ZwsIL4k4SxpS8eOWl3/51sJSM4NWOu41
bTT4DlUTN1z7yHbMqF1MzixgPRQG4iOQlLuvMPI9KGBBZnxghkIsZpRocEP7D/W1
QsSfqUpN3bvbnhGqOQaMcehNzHHm7jZotpcRig9HHQupRf8MEIDM5ntxDjIAvNfR
RpTMXdsYOR7JeDEL/GWeE+cZ+Tj7end6zngpVLtt1PyW9IaSPIyjO1BX3GzINdIM
Z0JKc19rVS2Dl1liHYZ9FEkAP7rMwsEN2QudG+euzpU5WnfEfSVog2QF7aVXbdVq
OxpPx3zh1iDVSPJEnEynHw==
`pragma protect end_protected
