��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�u㎺��`�R؋l�)D95F0d"��HɖR�C��lq84Wͩ�!�_.���� B��G��Mq��������'����(�16$q�Y����o|Րױ�0��4����<���ٰ���:� ��aB�Xe;�x�C���aKy��4o���n���������]�~�lƊ��YK�$���Y�X�/���C�&2�7�Υ����#lu���Te�H1���ρ�LS렮a��Юэ��c-\ e0;J��w�����i����x�=���~�yD����Ĭ����;�����#��E������0������J]�:TD��GUL@a����:	dLڨz?��D;?�����!�C[�գ���뒹a��w�=����a8$!]�=�a�;��yj�%$uv��ew���Z��#�k�e�Py�[t/�* �/�b�x��(�#'���f{�1�
%��z�>h�$�F��"�W�i�Xk�����1�>�����ҚWi}�����p��W9&e�]�J���C�<q��4�Ts��G�h3S���Ƃ��X� 3��vK';o%8���?jx�,�ڏ� ���_G�/9K`9��T%���lc~}�>������)9��n���YiIZ��UN��O��J�Qo�����V>���v�ʑ�3�d�ŻP��.�UTО�,�[��pG
/��'{9����^~�V���2�n�r�>��7�:�Ǐ:�D��)d�N��3R�$�~15���6�}@˞>���]�k��a��V�8�4�m��
�6V�=*� @	�1xѽ`s5K���J��y ����:�5�FZ�iy`��\�%Vg�a��L9��D7���GO�P� D�U�%��t+n�������v3p�8�UPwV!ˇw$0��^���(\�)Ż@Ik]H}:�R�Kq8SɸS.㓉��:a���S١�0fU)��)�Ȱ�c�}b	Q��ω)a�iJ��L��6:d�י:�Q��ұիr#�?�$��0�R��kQ�:|���$O9\]�T����Q���� Z�,?���v���JCy>��߭�����E�䦲\juC�U������G���O2��A��؍o~�u�k�Ӡ��> 3�1&�5"��'N%�Z��&p��<G�.��i
y�,}��2�ZX�Y�%�=�j�{�o}eT2l�6�IOy�wce�w.h�Ư/��Ћє��r3L�;̵mD��$^�~��r��2�8�,Z��N�3�e�'�B��$3�&o��"�#�a�Y]�]�	�R3��-�+�:��,�]gf|ͺ�Q֌:Z6/#.�	��;��Bp[%�{�3F�dq�ZgF�{��� f���m}cA�����#�vi��Z�a@�d_�+�_���!��9��0ab��OMC�ҫ��a.����8N��i*��G����3x(h�ja�	�b0�mP�<$)@�mg9!���2&xĿZbh��]�0���Xr�	(��oM���/.�G�-;���c��ŇWP������Л���c\��0uz�2��j{��AY!�	�^��(ՐHO��34TC��n�&X1������d����~U��O�Ӫs)���d��kJ����#]��~|����=F��hv-�Xʭ�Y��� �t�����)�!�u��K��@\�lr���+8��~�U�ZV�E��]�x7Ȩ��HRٵ�G�hő\���G��.
1��oM�9��(����NP"N��Rtإ�������X_�lԹ�'�6,`��fч-�7!?؀�����|�z�	E�Z�`0g 9����e����RjoaÉ��$��}!1B�}�M"�>gM�ܗ����=���Ҁ0����O�F	�Ǒ�#�׵�����O�w�Ѿ�p���0�p�Kp�0V\���u�i�'m�eq��O�qT�OU��Ejn*R��V��+���_UN�Hh��M,b}!%3mn����
�\�晿�&1�C#��7�OPV$#DHk^oo����=�����
�ST��#����	�:�ٳ�9�|W���� ����5>�
�R�h���Ê�u�A�xޒٜ�1�N>��1Rpi�*d�����&�������Px�>��H��z̼���������d���J1�[����z�"��i�(R�8�zl��曙���zL��jV�ۿ�p�N�b���T�ή���@5�oY�e���D���5�?R�
'lq������8?!X\v�z�N���nK��2��ߙ,�ɞ��8�|G5!E&�dlt��A���b&ʉ$֖������y�\��!����}�&�.�,dHؖ�0��g�܎�m����0�fIF=İ<m��v�w��1�?|��P?��9�H���:$��ǢrѸ���V�9;[�dYx�]W�����J��[1�_�EVUܟ?�����`��a�������W��gf��ej�B���@:�� ,棐՞���zh�^c$����CϜ�x�FS��E_]�̙�;�c��'�S&���H����3> �V9�l�x������"�CX���GJ�&	Dt�>)H^��L���~d�[*�������s�/�LL�ji�	�%x�o�ij4��8*b��UY��*0�e�������U�&���A�ڟ���ALv���~�w����;��YW0��5	���}��v��xjf�p2��/X,O?>?�jF�v��'sK+����������������qi���vkc;���*2Dc�\N~+&iuT�����S/fo�|����� ":�(���1�+�_T'�i�:{;�Ƭ����6��������e�B!Y���v-��-]�1�4oF7߻�{ۊSBQ�i�V���ϊ\,.ߐ"�
��\�Ń�wdMJ�JOI���%����b���~C]�l1d#�]�t�����j�<=7}�HqG�z�vLx(�O�e�B�(pG
�.B��q�������ŝ��'�x*��M�%AY�>0.�7k��'�):�<��2uQ:M�-��:lg�_�Y�y���)3�mRv�3�hE/Dg��e\9'�ȽR��QfD���eҝtR��	s�	����yӉI͊��}���eH�7�3)?��N�K�FMÅ�;l�!��&SΤ�L��keg���UB-D��w�����z����۝�9T�y�.J~��s�]k�����m4?��;5�	��֫��F�X!+�{�	�� �T���E�&��}Kyܸ�U��:��QY_sW*��Z��NS�a��6+�Jf�CmA#�?�0���oP�&L��`9^�I�e��S $��t�$tV�)P�jD�ϖ ���a�Ў���Z�,�]��F�XO/T�#߫dm�ñ7���p2���JB�YS�!�9+޹��/op�2UG�Q�k���`���V���%<��/B�Gy��2/�`�M1)�bnC�wۉ���o�?�_� �qѸ퐲�9�O��Q�=�4�q���(b;~HO�4�8/qA������$�M��������( ���D�Ύ3%���U׺���;�_#ED��t�aG֦�iu��S�&���H-گ�V�c�h �*Y~_�8�UR��ͨ��Ȑ!���ܪPP�2�1�fN���Y�M�++�N,�#2ǋQ4�jv�=�ձS#ʻ ��,���N��q�a����2�ԥ���>��:��UҰ��c�T�(�{/�\3
{&
��mQ��]�1��Xy���5xQ�mAb��q���5 D@ʺ��"�B:2fb;���5����y4Kk�����s�����@��bN�$��{7%5��}ƉO}1�{	�)�����#�<��M��{��hu�V"�Ɩ�'���&7�?���j"7��_S��XX7l4�:�W��Ow-ZH��d,KT'ԙ%i]|�3���P�D�>6R�����C��zB��:^˚��`��N�!Q5��S�ps|�`��"����D�6�b5$l�zp~�]��6��vA��B6"ᐜlѶꭤ�5�Y���HYN¥̆��LJOb�s�g�F��	U������׹]�<C읖�5�u�BFߊ���=+��5$�jF(��F� e�K/�)��=����������ɀp�K˓�m���������S$HC,\�w��c&ȡ��`��7�M�l��75��_��,0Y<�9Cǻ���g�6�f|#<bvY����x���� �!�焣Q^v���ǻ��@�=w�e����8����s���O��ю?�A��l�J�Zg�:�z���	l���<�`Z��8�'!N�7	hM�7�Q�~���˂���c�o�� �#�5�6u.vUD�h��1��r��T�p		 1�{i�E֧���KGz8�?7�T(n	�9}��5�{dG�EcT�E�+� ll$��fx�z�O���b�gex�h)=����K�2������ȹYvhD;#�̰o�b��j�1��y/#n�#���vg�Ij6�^8��_�I�+!׷I��=9�`�Y�=ƺhYc:s��a.K�s	2�&�A��WoA�nN��`5�<f��bx�o�b>N����I��V��� �r2�92|�9�Ad�g\���J�S2�8��(�OP�S����D$��sӞ�z���i��9�:���&Gx΢PϨv���A��?��S`�����E�+[ةm��'*5�l��ݮ�=�@�\���K�����h/RL~)�i�q5g/�2�>�QƷ�c�`�+�!��[��9�/ħP��Z僐��6�%�h��I��Ӎ�4���Ah��."�Of�O�<Ҟ��
�.qAQ*)..��-�j���O�o(-r��"3���@��%.G��G�=�κ7�Ol�+F�&w�=���G��!�Fd�$��Rm	���<4�ࠦ�&�|J����6⹵�1d��z����

���2�̰G\�~8<(���CV��X���h�g���y��������X����r���ߥg�ߞΩ
�M	Xxܬ��S��E�5�����06"n7.��(0��w���'�w�(�!�e5���R<�N���:�E�ij�0�uk�lzӋ̃Zy݌e��-��7�Y"C��'�2�'�����/+���TJ�(��F��n@�:?��ίĀ2��p�D�g�Cv~*m<��C���_]0��'�y&!�p"��(�|���.�`7^����r_X�p#��Ko.�'d$�̬h��T��(����¢F��|����`^r��bl.QE��7 �"��/��=}U"���{�0� �Zl��`��5LvnȆ`��u�ޘ��)��>��d���?�=��<&�c���+�q�JW���gsY�u���,�Zu#��3Q���9E���s	�Y��P�*鴔���?����{}$��l��䒿�4�hB�6����nħ=w�j�2Wp}�=�VLd��:�g��қ���
�2���)�%�;ks�����p�$�Ѝ��Ce�*cʆ�9V\��jm��d4�g&�b$*��X?�8d^�\En4}tX�vی�4t�J�hw?��ݞ�.�e�p���O�N@�8�ˊj*���>F�CȜ��|h&�#Lz���ۡ�ɕG��+/���_��ɯdu"*V�m�H�PO�Ztia�8�n���C�٧Ͷ{��g���)81������_"��b���!���
W��t�<(��?�j�p��O�d�3��c!�t���A�XO»b�Z6���<�?#��7w����j��N��Y�~{X��p�
_�唊�C�����$����k,[u����kM4>y�����7}���,#��]�b�V}n���]{������(dNjͯ��/o���k�{o�
>�V�]
m`�����\Y�F�E�F��*n�PQ�������l%5�V0�bDC�3�'.��*�-�A�t��Q4�ܲ���d��lbw�� 4(�n��M�m�u�x�m̪X�x�Gہ�F*�Q`:��y�?�Z����&@�H�S��j�rO2��h�Zo�c�
��1l���Ӝ"91/���~�;^[6���D!�7����O��ϭ+�j���rA��PiE�0=%D�z�O:(k��ę���������TN��-9R��.OJAD�E���ü�C�.��Q6&���Yڹա�yq�Zt��'��u�1�C��Y�ؤt��I����s]��V%_�2>xM��P���vx�^fQ5�*��3?}���~����X���t�Z��&�j`#���F����z�,�e��*[��\�n��ɬXU����q�>MDЈg�hQX�<B����k(�y�?�C�
�U�4B ��*o1�����2��o�M'�gw+`��մ�1�y�͗� ̪��G�i�Es����6�-�ъ,���I_���q��p!W����4������4bgK���*��`�If;�9�M�	��Jee�|w\鴩�J��x�!C�m�;ydf����6?<�2fb�,Ms�^���>%�3O_ߙ��0z�!/ܓY"噏$�X,хs��;*�J&��̬N���js�(�,I|�ࠑÆOBC��/4J�Ȍr|c·�M���~jm��=A��:�/E�/��� ���!}�7|�N�E���A䀝59D�6��:�Of�7�wV:a\�b�/�x�v1�N�ݣ�l���:��4YDZ����Ji��,�}�����?p#1^�H��B���AS݊���S){�'ٕ�O:M��º�C�q�?�oZ��Pq�gp�`v�}�)$j�� ��kJ��6��w��&g����_��`�J,}:L��F��^���+�j=�P*�@����o��y�)T7;�]g-Wp�D6�i���4/�B9�f�䚧��Tk��.0-!�$���)Y�F#�QDm�:N��ryr�D������X���~�݇T��|	M�V��BȯȣRD���FG�ڇ�K�
C��i�8�e����֜�)��~��Q�K�`��h�����J�)����v�~%KR�ʙe�\�v���:m�ޛ4���u�I ���%&O_�ut��F�H_8���l�?&���G��sp�#/�?,���Փ(v�6�OR!_��`r9��{E�ˆ<��6�BR���c���*�w�1����ÒSP#3�������ޘ�Wu�n.�;bx��;��_��v�gn|<H�]A*��=�YуE��e�@���Q�
V��TK���+������r�W}s��gI��Ё�[�E��8�:ܰ���(�Q`�C�l<L������p/Ҫ�F;KN?�J��w���Q�<Ym)㓫Am�H.���
��zC6d3�P�^�ѐ�^�<@Ŭ{�5��.��i$�p����'�)�����Q��K���ݕ�㸯]��0��f$�
�|��T��(���r��\��(��v���N�P%�D�W��,Y3��Y3�.��]�o_Ӣ7;x"�i��#��b7,�F%$.�v�q���V!j��pj�!�h�?�>�|�q�)��_F���կm���		;�/�Q��X��ݔ�y�~��y'�T}b��<m� ���"������ɾ�[l����񸆳����s-�q�Hi(�@���p��ʞ��+!s�T'9�So#v���y	�#��=pa��Nc�:�'����qě����E��Lp��[�,Gp�u�1L��T��D?�B�3��Y��s���.B�?MN�<��I�9�El���9���9MA	�ʲ��������?�����L/������ܫ<\��
M��\�i"W��#k�{iLL��c�k��@Y�̥\��z�$�<����n�D��
a_���~d4�U�`:��\eC�	w�f�I�h-@jo`�b� � ֪[*�h�!���>4�ޡ��I3��n�3j�L]�����曖7l5�v5�\�JAT�2�ű6�������T����9�,S��u��=�̑Ӵ;���l��a��*������;�r�5g��i(�����{��iS�2�ވ�����+.C��l�j�D�8�	�"���z����\|Z鋪�I��$��1ފFq�O�ס+�7	�h݌�g�'����!���A�gUF"/�Σ�I�	�/��@o����*^~7^ e%�ȿ0YbBc��|����$*��"ѱٱŁ�юB���$*�V���/��i�( x�|ԇ���Q̑�G^誑�(O�u���O1�2a�~l<H��������䢞���Û[����7�aP���kY9��W���vH��s6A��4ds��hlU���k�n���Xm�E�{G��<Q����V(#�CC��P��?
���fk����Y�qNƊ�h���B��70c��'�2�0r���a�h�"�R�+,7r��=Z1�ጋħ�6�Y����OD��&C_���LԲ%f��=y�wM��T������4Ǳ��P�[)���N�dI��ۋ��k���U����gϺ�(����.
��y���oj|��75��V�ġ��fk�=~�(�G�r�"���O���'�����b������D� T[��7��@R�M�MS��� ���gg�]'#_/����=_��/O)�NY*
A#�8�O�Ω��ƍ��6���w3�m͔��� ��"'ҭNҕ�Z/�i�(��i�y����z�M>���eݽD�ر���ֿ�hW�vz�����ܤ�&� �Ϣ!C�'W[���ϴ��%�#ǂ��@(]�Q�����a`�	a�I=Z-&����[��7BW�ɑ�8�`� ����g�l�ˉ�`گ�>��运��p�M�ʼ��cr�'�j�pYxSc�0��f���S��#��EU���e���W��W6��u��G��55��	�*�/�3�3�gh2�xrݚ;ޅӊ��*os���ǳg8#�U�d��A�(a篚iP���+�/ɝJF��6n\������n����
�O�]���l��$�E'��H	o����RC
�����(t�d���6�v�ʠL4���oDp���N�;5��I��N}r��	��9}�Jif�|i �1���/�ۨ]O_�[���X����M��\L�X�z�?�AA6(����+�\���Ε[0/[��I�>�>f-�Li<��a-�`6g~���oj����fK��>�,x��7����$�������m��T�D���E=��
�)����$ҽ�2{�x3
�IZO2ci���#�I0��+�n9�b��W6�D����k<F`�yD��vlx�z�Le���=F�UgC�%�L����Ѱ�y��a����~���j�� P�z�#��N^K���i<�7�]pg��'��_�E��ư�7�PK҆����=*V�C��%߁����)3с�Z\��~ԈA3JD��ޣ�#����)��܃�w�䎳dc��X�Ct�W$���(��9n��gZ�mZ>䑧�(Ghվ�K`��h#��&�w�A��;~9�+"v̏>��/��	��h��JwA�ܿ斏��U����������$e�gKc��Q�j�R�ҙl�l]�	C�`��B����br�w*`t&�7,�:L�~���/'�kϴ�e]��zk����}�tt8���������P��cc����3fˠ%	g�31�9y.��Q'Saw} I�sT;ZhN{BY��0�!��)ɘ�r��G�w����8,���n��	�!��=G�@����=�Kt�ի!Y
^����<��hl� B�˜���-�W�2|����D��� ����Y�na!DB���rp�ΰ֔F+�����ިd��V;�.�Ih�d�{`t��S��v�-��n#a�W�� �PL)l��m�;gI�M�W�����/TZ�"�T�`ǿ�ba|����=X��tD}�s�_�;�6_���A�����i�@B9�I���m���ٵ�#���H_���X��C�o������qR[�W�c��U �X��-�,vQ�� �KNT��5 g�ο�miT	�X���óR�K7��7g�kK��%'!p�����d-�U�D1�铚��c����p�-+M���y�9��k���c���V�jͲC���j�`q+�˛���5����ov+J��ظf����ls���z�8^_?����r
��1mT��b�I\":=~pw=0k�~�r;N)��)]��PV>-vF�x��@��N�[v���x1� �@���T7����p�D�ӟg��G�i}���� ��¹1[�mI}P��fdC���1��@"�"7��R���7�`�-��/�r����DC(�%�F,�%�EA��l�����Ü��w��,�IE��}I�x�{�+[� "i�h·K�R�����O=��2��0����D��������>�33}���y�B�V��gsA���H���NA�c�'oH�m�M9ǂ��K������3]�K�%x�k�8��n�ew�V����	�>-,�gY��jmCӃQ*���ND��8�q�M;Z4��ǨH��LX��a��I���ƾc�<d����S������9�&�rn�����bR��YN++^��B���͈=b���I?�A��߿�r�3�m��q-�;"�
f�����qg���R�2j�]0�k<��?v2?ʏ��u(F��F�޼�v
CI�TU�ԶXA[�T|� ��"����a��]�7�L�֪��ݢ~ت�ݣ�OY����5���{>�EX�e�ҁZ��jaa���%De��Z��������-F�+pˡ1�)�
���	m���ʎG�m(�SM&6�-k�}Y�U��<c�h���]�ًrwG�Q��K����.I�'�d�?�����g�)�b�_3�������
`�V� p����B�n㸐W0U�nN[�M���l�F���s[��8��+TX�5��u;�X��OA]kS��+��ܳI�3<O^A$(}y���m���>k��� n7��ֺ���z��	p�D���7BWe�3����k��Xy��/���{?�D9=w�m��o��51�;o~�pe��	8f��}��u^W�,�t7��������RK2����P�����ִŞ�e\�z��"���[��������y���
Q�����F�� �¢�����{Un4��S�f���&=�^�jHB7v������ˇk�f�V M��&��t 3�gB������)d0�]E�\C5�:{����G�H���n��dw���\���i��	�q�
�g��K��cJ�b&��zo��+d���t5��!�RL7.k�G>T�V