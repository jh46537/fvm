��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�k��&��Bvx�s�!2����-	�C�o$���%��e]YC����td���bQTTn5��r���]��ו������`��r	��ڈ^�5Ng$�]��� ��ڷ$@��VEbs,��v��a1����UiYAY�֮�}"�ɛAJ����Լ�N�$��Q�Z�����I����\�9Z
zd7���<$�
4;���/xLUd���\�נ����{��?ҿ����8Iј8^�6Z�,z�7]��Uj|dӣ�����vE�����{�M>	�V���_~v���ܡYQ|{s�a(�lK����,�>T��3\���,e�US���c`b�()��+!�H�q�]����CV���F��^�~F1� ��+F�H7�IT�!�S�K�-��cW����=��8!EM;�X�ß�Z5���71��a:�CȻe�(�;N1;�Bi��[)�{��c�;�:&�{8��p�w�^�\G���su��|�]��	'����4oo' �p�e�/j�Gf�ل֘�#�L����Ys����L[Z��Q�(p����J��Mw_-u�w�M�,%�$fG9.�|\D�%*	�2�^}i����3��ʲs�t�`��A�f�ǂt0��q���J�ǖf�T���5��9i4�.�6
��+��S���X/t�Un�n����"�׹�U������*��@;����RituO��pF�$W�G+~}[_�MZ��� ��=é���Ӓ'-�kr��̰*�h�P���?�xG�\�� 4��acf"�M
������qp��};�U$�\����m�"�1�8��4�$4����
�9y&�彧�XDyjdvL�$��ƥzz6����]�Gl�t����|g��X �sб�8�V���8�q�5�l!Za���G0�L��3̺!���1�+����F�L)��lʵ����x�,�̕��|���j����`�����ȴ�~R��v�IIL5~�i��Xl��{�O8�D�5�^�زՔZ������ K�rf�� �W��O����3��{^�Gr�릈�|�&H-�~��ǃ[�h�
���/&��u)^g�au�/�9�"νem��W����&��~�:�5�--"�����!���;ʄFO�a�����,L��enG%�rt0�R� ��bRǉ��Qk((�Y�8A��E�:���s-��?�Ff�'&I����������Yz�d�un�<�"Eq�/��|�t�}��nɤr�|���=R�/�3�[���Xu"����%2
*�1�+�ˌ!���X��D���9JU,��e�]Ksm�yQ#�� C���rx�T���j���v��G���v:0yB�,�\���BcBYZ���L�sjyS���)��:�;��3��)֭�7j�^#���҉Mj�Q��T���\%���z�n��|�mI�f������&\Q�bH����
����e�A��4.�˹\,�hޥ���#�f��=f�����vM��+�����繁E���	�Tqn��h*̀-���I{�8-���.������2�Q"@M �Y���fBRHH��Vfl�>F螒;$cۺ�4ߧgR�#���l�����η���B§������/i�)Ϝop*a>З�	��j�v�ڕ>e��q�ρtn�7b.:m��Tݢ,F�(,xl�?w��N�K
��H�8����J=lK�1�!�%��Sjsp[ݻ�2���K1��	�/�'���u*�h�"������,ݓMFg8���e�Mm��ntˏ�w�s���ӓ祬䈘�2�i\�v���Aq�NS� ���@��wp�Q�Fҗ�m��н��6k�Fm��
ڂ����l�w�H�A�)��b���\H6�Y��)��7�D�����^����qY�_�]x�Dyj�ژ�d�>4��47Z�)%�j��[EQ9��+��"Z4���~ެ�La��/�Z�cƒ���5�\N�M�{�_���Ϫx�W��G_e��
������ﺑ��XN�><��N�����N:�"�u���e�\��-QìK�N� ��/wTB��8��2>�@֭Mt��h�m+J�-�|��J�����gN������oR
Uts9���Jơ_q��d��|��SP�BD�hx�F>#��/A�y�1��q��q��wcl�|7c��ԡ�,@�=���_�R0�����NPu�+�C*�����c��`�[�yC���J�^LD�����Q�l�L �ߕD6�� �Qء{�' ηX�Ʃ@j=��M��']�Yt�`�Ҟ�4�Ҕ�o�U5lRI�BI��C�5��cJ��v�G�r_�/� y ��	?�wPZ���i̅���vF/����6��&�Ē+\ OX�0�Q$�{t;���D�@X<�@�ޙm,�Ĭ��u-�R�b2l�[���7#޻nzJ�,9<�&�~Gӭ�YL
�ƙ���Ն3݀p6_Zn;*M-\l��S\f�B�F��}�r�T���ɴ@R��X��hY8�oQ�|c�lMi��g;���#"i���C��7���VU�a�{<��˃�\:�s�p�ň �ǿ��f���+([�9-��,k���/�I�_U��aF�)	-��2���"Oџ<R����ъ�H��5�JI7�%���D�S�`���05%	��YEez�����hWͼI]
�r��CH���-�E��Aប�C�T5���C6�`&܊��\+��ڙ۞�_�.ox u~c��!�b���Ǖl܊��I��v��;�����L'�Z�WKH�y�?�$ґC������$[��'�Niď��&nN��ި���������~o��E�P�=��HOв���L+�5��}�sՍ�R��5/{g%�yqɄ��[����n��\�+(�z�i�b2p�N���>Om^�)��N[��˃"j��S���(�)f"p�
b��V����\��q�!Q��&im�$�`�v��"�~�I��.�K�@�d	�`�RSA°Ҿ�*[́�(�0Jבg��>8�il��!������}E��d"��X�3$���"y0"���O�:Ă�5��%���|m�A,L�����v. ��`�� M�b�h<��ј�ǋ�|���4���kύ�_������L�^���o��?
rP��Q������Nr���q�iB'�� �y`QA��䴚�r������Y���͝Ք������8��^I����Q�N|�={�hr��HU���X�w�m0�����:=q�n��j�(�/酃V��\�\|�Z�ok��@���EI���j3i9��.�OD�z�q�~�|*l�'
��^�T��������V㠘���9
���2Ƕ��<G�?f�����o�$�G_�W��3�]�<8����a0�Д{{2��[���6�[���V�@`��SF+.�S�,��&����{����Le,15e$(!�����.��"V�U��26>j���K�kzw���c@61���t�\y(���tl�1졻��b��s�H����{"w�r���]�0&�o���JY��&����F]J���c"q��	{_k1h^*E�{B~R�;��C�ſ�;׺�_�o�\E�E��Td�����Y^0��<���@ҏ�Q�S����[�b������'�d*�`j$7�]I��FJ�r9���}�;�V`;���.�!V�ʷ(��$�W�f�F[����=/�;$���@ku������"t9}ق��YPvuZ�~��rG�5Ӯ�� ��H������=|��1��Z���p�\��:�[bvW<#�$!����Q]A]1Ԝڜ�H�z)/7K��AL�j�[�WHUҖ��̺��T@�L��v�F��p����,qJ�S|5�O�u���6}*��p%��i�wʎ���r�a�U���U�Rc����*��M����0q���E��.�,�f�o��|&:��~ߤ�� �C,�'V$R	�����翇v*�v2��#:����Ψ/�!9����:?f�POq���
��o�.{�� t���QKO�OW�b��K��ag�݂�O�xM�k��	�y'V�i���偫����c���.�U�Qu�F��Щ�cPg*�]6K.+�A?����xʅևOrzP�H�\��V]Q���x�py0i�1{8�c�a�"+�g�ٓ N�>����//��آ�&�/��.���A�Un!p|0ok��x��t/���1ӑu�5AEg���a�a/�3+J����zM��X'��a�Ւ!<c����NR��5�.�3�9љ�FN�qfv>�*��Q����&�+�F�|y��� �/-�(x��# �o|��R���63�=v�텅{Q��>�/3���%5��iɬ�`�\
��^T�S��j���n�<��3�ˋ��ĝ�5��>�#���YT�uI��oy�51��Eċ�'����,s&��:���-@s�x1Ͱ�\�?��+�*��h����DZQfӿv�èCɒ��1�X���Jd&L��LN�xQښ�-~�A����;�B& ް�dʣ��R��Գ����W���5�}��{gH�u.�	ΊF�]C��W�ץ�F��.@9����J,�O@ȭ�������'�͖k���s�!f�e�w�^�lqk)P1j�y+&꾄d�t���[�[O����&�/ll����{�2[ҖhN�X�Y6�FSz�
����S����Mu���U��tu��tԬ'���2�['�8��U�w�hFN�OYJ��o�&�6���o~��D~����ѯ7l��}�']�w˔w��qwB�g�A����P�m��Gi$9�Wp��r�L���v���ì_-���{�~��[푑�aH���l͌Ԗ�c��:���Y�n�~��i���������;�d��0rL^!;L�'c�},)I�:o��D�=(HA�D����e
���V�}?�rB��B��%�HI�cLYӽ��ضՂ[d@H���g�o���C�\��ɢ�2ba�k#�����v7��e^[�+�Nґs*�d��@���kTվ8���_���4��ʱ�^�vU���dD�kUQO���Al�n��U^"äБs�F����B`A��-�I��u����s��0�{A ��!*����� ��m�#�*��Gh���vcnV4W�;ۜU�v��e~�X��F��0�s��b��оN�/���f��Ūv.�Ԑ%k��sH|l-Ʊ˶���ı~f�	=�u��/A:S�1����	��T�_ �Ta��U��Z�_��L��}i�u���W��韠����oz(μUd��7ʣ���=�dK��`3B<�_�w��n̲���4�fR�v�jn����J�]���j���,Ŕ���wK�٨��lL�����n����'�A3ϓw���J䩃2c6rWy㺞�b���ꦲ�������䁾��)�Ԍ���񅇇���m
-�����d�M�̣�?C�\����y}
�k�X�\��(�����MSQ9Y�,�/����~ys��,.�Z��X`D�@����Q({gec�>iҨ�2��6i>ѩ`G#dXs�#������o��.�2,���B�9�����뺻Y��~K	�5��f��ۦM������U�"G5%V�1q��..�i�=\�1�!%�ػ�m�]MQ�T�7'��=���_ֳ3�l8;f��^Ȱg�V����g�{~�5w����ni1Y�����Kfΐ��B�u���wp��c�Ɩc����t{q팑�B\.���ܦi:SdZ���/2�m�bPZE����o[��ރC}f��1]��Tm����E�NO��9-�~�ޔ�5��36���G�ƿ������EXm��� x�2����+^k��^�������@��o�ʸ�^ʹ� #������D�G�rA�ͻ��$R�����Jň)f�J̮�'jc��!��_p��&��}*�#��,l��҄7�s��@�'M����ʴE�n<������/��w��_�F�Z�\4_UW5��+�ҷ�tQ�7ګ�d>�ɤ��~j\z��x�S���,��!-b�������	h���=e�8��Cy����f%��x����1��unl�D/�����n�'����!(��("ߕ� �g�h<�ϟIW�ֆ���ΰ��0Q$��d�9�b-H���j��0*òtyz����vr�Im\���4Q��ü��l6��N�_��i8��e��������$�k��sԪ��,���#�L�9ko_3�gf����
�s}���yQ&�d6���, e�����8�h���vu���2Xbfؑ�T����@���ʵ<9dBtE�4�o\��B{o�*߂�gC���PS3�{]U)�;8Zt�����oߩ�� KƠ�H�$�|��E�]�Tӡ�b�2�tpL8(BU�u ��5�|�bg�:��ǅ�<�9��7�Y\>8��4 %{���ꙫ!��Ȟ" C�jt�z9��ȟ<r�'6Z�� P�F�W���aΦ�%S�Y߶��?d:�y�$b��Df-���YiG�w�k_���B�)��, 7&����DQ 2lM2�-��k웸��E���=�@�1�4r��J�����1%s�5�S%u�n"��[&у��b�@��8�+h�o��?�x��}�0�!�e���h�.5(�Fj�a�$}ΦP�1@��	�����|�g?��Q�wA>�.폰��X�e"&x�#���:���$��_hr)4�#�eқ���V��
��ǕZ��쿕� @��m1��JmPچ�<�Bi��x-�e�ӽq�F�q��D7�&b��!!�t?�b���7� d������\O�a�MOg+91��9�]�4��!C1�:v1�w�n~�D�Ɩ<�y���LA�P���މn&<|>~X��:(�,\N�gn8�o�L��v�U��ɭ��,w��k͙j�tՎ5����g��n�Sc��� ���ng��u_]��3!���i`Go[��XZ�e�䐳D�'�iP_�I����!,��e�-�F���8��9��A~}�=oC(��z.=�N*���z��A�}��Q��I��+����AR�L��	=i�>���j�J�_mqr��a�	�ڣD���<��\��H7r��V�wD�B}��9mRؚ�ٵ��ΧC?(� �~̱s7`_�����H�A��w���8�tɱ�(	���ɑI0i�-��j?b�'��>x�!���53�O��-[��OA�z�C$r�ln�tq�и��yCt�\pP,<ÒS���]��ot!����G�{��7W6�Dt�
[h}�P��f�q���dS v�&��6
��#�CC��FP���� l�C��y�C�de����	���q{`65�
5T���LMĥ���{[�ѝ��xy���gRCk�z�_;'��m4�@���v���-�����P 饣Ifqp�� �2J�N��ݫ<���.�(:�H�����j ��/颃�m]���I΁�.0m$;�[�N/��(��f�=�)m���9V�4�#0��
+:��.�	�'-X?j���J#����z�3p�w��-�j˾�p���F���M�.����G�z��}���O��u�ޗ�{���9
���h>5����̶�C՞��0�UZ���
��˟�V��`O��2;�AK��F��Ţ#������KB#��x�[G�*�qŸ}n׻�:����Ho��P�����5�R���O���������v`�3SW�U�&1f�,d����9zt�rڪj��?��4�䧜Ŗ�gT��R�ߛ)�	�lъ�_��2C��Z|ՙ�Ʊ�hh�7�az��"��$//.�fo�)��()���)�m�P5P��s�ks_�;����18��>���k�V҂1΀�����Ə�ߟ[����x"�+����ԏ��I$b�:o�+�d�%*ŃRiFZ-�>��8��p+QV�۪�0��}��Wʊ�������Vv���z�64=jRR!=a���*����:=gH1�[BHU��N>U�xqU�(/��L���A��ه�=��LM�!�z\p�X/m���u���7�U���]�ı��8Y!Ơf��E��[s�i;B*v���1��h�X�-K$< D�%{n������nY�7����[�hr��R�wL���:�}/����L��o�ܕiT�xƞ�[t�ǹ�;�p&��m��Ţ|=C���逽�.V@Ҧ�ˬ�?7�H��u/��rd��ES��C�O�.eW��P��^YBb�/�­�9���o���m����}^���μex�1��#��� <�{X�k�R+�:h}��m)��%o}���d�6�Q�a��ju�7=�⒲_�#�xbP^1��lׄ�k��
 dQ�ʳG�^?w)�tU��B���rRGi��J	�����s:�(C��m��&뎜aA����M;Ǐ�>CK��|;tȵ�S��%���v:l��q+�+�q]B�E��D�ʫ��u����/PG����m��mc���)�-�q�]��HIyPn7Uq��9*�Z�[>�d�`<Au��L
�'��$V*�b_�nk�(>�V�����.�=_K���H��u,�emN�؃_�qo�/gP��	~=SX��ڙw�3�$Ѕ���T`)<$��D�c�Nʧu|�<G����_�i���h٩kYV�&�ݻ`TN��!l�����i��kTo���9��� �Kqf44�-0ۧdC[;�J'B����ǒ:r��b�����W,��أ({vq�������nT[{�Id�h	�fN��_�2 ���D?/S)�q,���wz���Ks�A�~�H����YE��0V�o��^�t�z�+�L
A�4�P| ��.�ZΔt��r}׬����o�)wK콝[�D`��>���.�Q���M-�y]N���X!����s�V!i��qq��Eu�6��pc�f�k�\:��ӗ+h���'��~�NJ�m��#_:kuP��2�r�b�YN�^h>3��~���_~��*	�D�s�N��	T���3\g/�D�'���;��Ql�a���c�(8���y�܇k��6h�������� 3�}����x�� ,���X��-�9F���r�M�́�MC�#�T�{0#S��/q�wC4���Q�}�M�Y��½�?ܧ��ݸZ�_d�&J�������l���DS�H���h���a�P�q�_��E�tZj��0IS�{ѯy��*'\����d @ o� ζV�j�M|xG^5"�ā�q)5�Ni�Z?�sn���?;��u7C)�?@<R��B$����+(_�qD���浩Ŏ����5�o`�m_3�P�~w9x�V}'��D8��U��E8��i���	��ˌ���a3�-Y�����:J�j�#'��W����J���bR� ��AX� ՃH׊V�~��^�Us#'�)�vTء��z�cט4$j3F1��_�$������1E�]����U���2Y�B֞��!��C5i�Zp;՟����SmLǴhW���zt�>7*rw�l( %ځ� ��J1��pf��\�
F���V���  ވV���Z�i&�s������?!i�=�y���X�_L9�@�8h�dq?�|>KM��T��T^�[Щ16lsFڟ���u�ǄW�
oJt7?���G|�/@%�1�v���ކ��#�����ͽI���׎�S�"�S��}���T���6�
�ϻCS�|g��^��H~�n�Z"��Gw{N����݆����Q;�r�WdZ�Z =w.�]���zSMtD����V�!�'��?
���5���@<��)���-۸y�9wB7r\�a(v�l��f�|
�g �\�[�٣w�5�_�r uBJ��FT�7a͠�_���bA�[�_k����J
��/� �Ȕk�Mw)�y�������;&��+4�oxc����m�}�N8��'�7�����@^J>a!��җ�#�����V�@e�Hl̪�\�Ϟ�k1�4GX�Q��]Vq��	M9&�S�U��'#»XG��	K�����s��,q7���6����˭�gk��vӻ�/����Vy�knr��]K	�'�h�m�|^��`aBr�'h�O���nVL	�E<���*D�d3���թY��Z�Z��&��@H:t����f���g���L�ѡ����]����l��!���9�䬮��Ū�1I�H[��_f�*�t%E�R����̌R��q�@Xv=x�c��ݸ�ļ�Gい��a��ek�=r� O�|�C	f�5(.�Rڂ��ʒ����c�]�ZQ�{�D�$gq��,�m�IX����Q�y�v6Xb�4�t��������G��Vv"�V�(��o(d}px�O��#9U"�Mȷ�nb��+�2� t3�,G/�Љ��D�i��C*th�����烥脞h�!��P��˝��h>��0֬4W?A�R�&GD���z����z	�Iyz|VG�[��ms��9���&��ۋX���HOQ�$��QMW:V�zCf�PDz���铧��9j��l1��N=���j�'/��┭��*֕��A��\A% !�:�>r��Vv���5���[�X�RZ/�\��:���A�8ToP�̛�r�����m/��g	R��{����ߠ~�ȇ��E뱡2���@q�&܊�α��a��������sw�4$6� �?���=��w��]��UL>p9���+�����o���>J`#�����["�]l�uUgb����"7	++��^M��I��ĐDg�COa��w}bJ���׸�N��e-j]�0��~�
H�M��%�NEր�E�]����{VS��*�U�����9��`C��d��|b�P/\T�?8���'u�騦)}��������ϙYH:x��\o
Z��s#M�De�;��}�~1h4��[.H�>�~����&#O��:vqM���`��oaU�!�U�45w6��������k��^�󣢐� ��q���p?�w�/��u�"ᮗ�x}^��
���	�JE�Šh�{X�20��^%~�`D5���mpS� ��HIi��� N\j;��ݻ|�_��x'y5�E��W�S<2�+PD�q+��#�)��Mz;Q}j g{nԚ��������Ce��<=�&��)��*
DCl#mM������3���^�u�ȯ|�V}d��]HŖ�H�(���4)��Q{�#�o���#N�=#����p�j8���ә���ߒ< -K�	&$M�L�<�E
H�M7�cI(m�������e�PmA���&FB$$MkZ�?>�o2���4��j�!x�Ux� 3�R�]gݪ�¨bV�ZG��!A�P
��큏]���T"-����Ou׳��Y��
�Ⱦ�ջ��dK3�k��3�̝��^�k��E�vb�Fi �"�=Z%8cf� V���<ӂx�w�o �3%C�kjtX�/�����\�d ���m���,��*��V>R
�/Mu9��z�S�]1^W��<�4d}�!�v�6D�XX����uj�M�d�[�C������lh�����6��-Jԥ�Z��*ܽ?N���W��%�p���1��a�'C����2M	��i��W�u!?3j��Xp���Y�b��߬j�l{XԽX�p5S3�_x���"�L%�psf� ��v������7�����K߱N�k=�sǷ_�qH�<9��
�!j'��.Ƿ��m�z�r����u٫H��*=$�7^@�uM���k��݅d^}�7|.>d��z�Ӓ������-��{ڤhp�k��(�O�x�ϥ���(�X��z��W�=id�&�N
 ��0� ���g�_TA��K������J��99@����G���z���{�ݙt�OJ6c�v���# ��ⷔ���P_7��u��6K|"�,Y"@�f�_T��5/ʓ�oCQ�����d٧��������E�����Zd
����NN�(ܦ�7��G?d�m`,9����[�Wz*tA���]Npm����e.��$�[��q�ʊ�<��K��f��n�Q-�i�?:��qN����}�x7Fꁪ�'��o۾�ۛ<�k'Zæ[�Y�4?Hճ�\r�T��Q��{�ݴF|7Ĝ�Y�����T���S�"d��M�Hy�N&�x���z����4��H~�cU>ɻ�Z����JG�祴�g�ZF��S���x�N_gԊ�OE9R;��
�<A>�)]���p�!�
"�4e|G���cɾiҭ�oQ��˲��0$��N���b�����q�D�K���8��!Ǡ�N�:��hʙ�p����-=��i���F"(�! '��!Z���E�m�v5���֐��
�{�;,Lh�U��������NF����C7N��a��M�mMaV���D�n8�J�o@��8g�ձ!AK�S+�`|��ӈ�=���l�׈л��k	x��a�+�=�ur��K����){��R��F��>��[��s-+a�a�@�.�I��ǜ���1��8bR_zu�@��|}�|vg���ǭ�]�z����ukg�f��Q�3(T|?a�Ĵ����E��&�_��"g��5ˊ_E���2�Z1RL?����mWP�{M�hi5{SN��癭��7V����a <�g��C�c�~�}�}A8����%�M˩��t��	Kw_���;	�q�����Gϸ/ ���|��ua�{A>�����8��7�;�eZ����2AA(6�_�n�jݶ�E|�xm),��_|��y��!��dt��ם<'�kw=f�:�Db�� �^дb`@�luL�tMB<؂��MA9Q�?�"?���l��(���yXvA�^���}�W���O���Cj2h����F���f�͏d�G}4���Q���[�<u��aSI�1aV�����`�6k�HN.�<`��� �0L�W�3I5��'��HC�Kw���Q:Q�����b�ռY"�xwk��t��̗fV�S.�I{�}�ӿcU���F�^�f.�5�'�>��ʵ�� '�c۬�>L2��1�1ѕ` ~aN�"����ͼJ㭓�����S:V��-;:C�Dd]��ak��p��-o��	�S����/\}"��tl����x�D����{d����Y�,������t����QI�T9��ubI�o���[��Ԍ	z!e2���]�O�1.���W�_�"d��~�jZ�������9�C�Y�c��Vx����0���'Sde}�*��eA�w��GԈ�R����?~7��9-Z�ohZOam�0^�B������q�G�@nR\�)�N�	�0��0��Ɠ �'y�oa����JZg�#��0������VRo��ǧ�4���ے������0z��!xP��y��u��4�;��~��/˚Å��W��05i�:�<AE�Ƞ����Q�K�B�5��[��s�Ӎ��K�V��l%����,GL���Ϛ�_�g ���\�C|_*�b�ū�Rg�	�:,�ǡ�4iҕ����H��_G�^��[�T�8����R�/տ�����fw��&�v�Y��p((�������5�ƣżm�!�Ř�&lɌ$*p 5�å@�d?_8Q���$�:(�>�����.y��W.��� ��������Hy��������kˁ����Y���>Z�����U�U���d3,��7�V���[��n������.��$ٷ(�W�@Z�Eš���.&�P�蟜(g�2��T�x�'��ȧ�;�o�����i�[� ��?~_�'��܈E|ǫ5����Z��O��HSmZ��d��A3\�#5\T8��A	���[�)��h�~���Y��R^e���5x�:����5��k=���bS��+�	�B�pֶ�?V֝m���ސ�d�����`����ó��5s,���ď�Ԫ�J�B�O�@V1�##>bm+��kZ����2�w M��F�6��kpvG\O�C0
�����匇����
�7n�9�(�5��;2����,0"�����[�����/n6�$[����xY�������Ma`�-�"�����zO���O
;DYD��Ŝ�?ɱ�7Gf�9/�Q���N.E�#�Y�[t���ɶ�ER�}�?�K�"%�Q0s2.m��j���;�U�rةK�8Pz#�{�����{��Q�ھh�+�bx��Ps�#Y�gpA_WӋdl觥	�jj��6q���Q�EΜoTW���ز�6��H��9��c=�����|�9xE� +Y�o���SC�mp�(#j�D�C���M�X֌a����U~��hXob��ˍ����C\~�"�٤%�®�`�����&4�T��Q���`%kDlD�
 f�}��4�vr�=�:d���������@��ń`h��m�[RJ���7]�:o&�fĆCafD���Ah�����|~cB�%��̡A��d�z^<8H�i�=T�|�c�1��]��|h��Ce,Wc[����ǥj�剷�F�����j�?P҃���|y;��:n���|y�T�== �VJg�=�h��kٶ��qQ+0EB9e���t���v�����پ�ŔJ�S�}P[�J��p�"Mo6;����^�	&Q���8�ՠ��Yk���u�NP�ꭲm�h��o�PK4� ���R�Э�b�d1�J�,�-�P]_4�հ/�o�ӪX�>7�u7�k�>���;J�����\V����Ū�GM�5�g�v}
��@�'o�m�e�},R��WcBF,������
�D���	Yo���̱'s*��&�^�Y���VXh��U^�#�����=1o�ҙ]�/ ����͉�f��Tw׆��[U3_�jo�+85�imh����,T̼m=�b��x�$堾<\�Ƈ<�>
8@Y-��sw$��*�H�����Y��:0L�4:��h;����\�����o���<qR�6Xѯ���G�n�+���Qb^��O:)cyp�PT� z��#�!E�o�׸��e����?Q�(K���P�`⣊���_���"�qg̾Xe��x�W0�ֺP���5Ã�l��Ф�BUS�(�C�<�V�B��u8�M�2i:+0f�"n��ЙP�7�[�Y?�+�,9?�燇��%��ɕ���ր�S��NkP���6h�1�S�̌�nw���>�3\D�,�����$n��WP����-`��p�J��]a!𩌆��"�����i0��&��v�fe�~&��|M=F^��]��(\��k�!��&�L��bu%vh��m�y�����-�c�o �JJ���\I��tx����S0�~��"Q�k�0�џ�uE�n���[����&���F����_��z4�_J[��P�aj��b���#��<P�.7�3�l#D}p!��T�W*W6`���J�1Yd�y��Z�2��AδM�-�X���bNw�[C�
m���yEk�V8�,�"���P%��.{@_�AdC%�a��ɤm��d�F�g��z�'���8��5 �U�e^��]�>w߹�����?�8�ϗ_>ߡQ$�0� ��I�M% ��/t�Kj$�i K��΍<�UD�'+�:�o�%,/I��Z�������<�@7�Q$)%��M{�Ȩ���p�k��o������εڤU�մ��#c�'��l?}�������\C��K
v�t�azqR�"�/hj���Fg=m]�:ᵸ��l49K��n��YF����q���m�7p�m� Oԛ�d��8)M��Ҫ`�K���x�4�!�z���G��9���w�^m!�v���<F�5I��]~�����_v�&���6h4p1%0�|}��] `Q�/�=�|�Z%�����B���?��l��4�gf ]�8̨K��|�KZ����v�Ϥ�l��	��,�vOc��X�q�{�C�UB�0�*ڔ��T�]��M*�(����Q�Nƨo������6�Z�|�t�8��џ�V����:�\����
!��F:v>�	�K��ˆZ�*���=s�,ӱ��t�@��2��L�k�M(!�?�"(,���C�&���;m�g�K}	n-�z�v�6��ߩ��O�
���Un"�\�@)�`u�L(l2���k�*�9��:�iSw��&9��YB(������IZ��/��t�ۂ�}s���o��~5�9dΤ��^=��sWռ�f�P���<wt9���
����g	ֶ�p��M��FM�S"��p���ޒ�:�˿�:��%�s�Vqz'N�Ý��O9�C�hW��P�U��>sy�ZB��-�퓣�[t�iw���{�6~�,���EG�)�ҹ��*>�9f��䌇�o�~ae�w��$B�El�#A�����Bp���^�?l�� ���@�7X>uh��,:���yl��(|Ș��y����W�m�C���I?%��X;.�A{#�1!R��ܜ>ft"�ⅺ�kZ5eoPm�Som#�>�Dkܮ�o4&����|X�R��R����wg�O�#���@M�Hٔ��` �!zНkz4�������^�Ө�mz�K�#�!�����Kxk_��O~�o�bT&��Fr�X�43�j�n�a��iYc�.�£�������h>Y�S'�FYX�����lܙ��@d����sQ�]�M�i�?�E�0+.�T"�o"� �E�`\6+�j���I�C���m�ue�Y�Gca���Q����m댢s�O��h�>U�YY��������صA���rc`�'d��?i�@C�wZ2��9�����3��AtI�f��
���/��[�y0FZ��c��B������fp�XII���
��;X��U�޲ͨe9�(8������n�}Y�5HD��湥�ֹ�j+H�%O�����l�Bhv_r��U2�S���9�Bv0A���D�/�$��@����p��w($GR�"����!���*B�nk��OM_ݕJ�.W�q�Sr]z���b���N��2�`BP��}��!�fk�g�@����kt�	�脌����'sQ\�֖D@�����.�\l��,	o�H�����Y�'����)ǔ����S:^>�[=������c�;��P{�G��|�oy�� �C���R�Q�9Q�	U["lկP^(U;4�HX3P�`��To��2{x�r�╛:lbN��%�`^�d�>٤]=��M�Qt�z�Ju�F��b� 4:���PV�!������7>>iͰeʁ�����z��MkI�,�T�i<r��7��N���6N1$:���x-�'��~�h��<�Vܜ$'�	���T�Y�?� ~�jhÙ��������"6��`"�ӈ���˃f?���
uHk�g8�ZC3+��ڌ[-���RZ����Vh�s{��|.��[�A�1?LwNM��<,��In��t�Rq�E�?l���ۉ�(2��i�`)z<���0	P	3|P�h޴�9��TU�N�B^����H���̬\n�����ƶty� r,�߫��ȃ�y#_�ȅ<��.��r�I	��^�UK��0T>	XMN	�h��p
K���u��b�)�Y�{y��(w�Ew�f���SX��V��s)�pzoH�7���>Bl.�,}�w�&�ׁ��f�?*�6*�sDJO�'�3q���:�Zr ���Ԍ�Qqps���X�э�,���~�a���_`�
a���<{��%e�7�x-2���zW('Y��-{��A�1�z[�@?&C'i0������i����c��{Tzu�b�0�z8d���3��b��U1�Qo��)=�^���J_�՗�4�׊���e�����<���pF�{���c�k#9��,\PH�/[��ц�Q�i��!0Z#/��
C`C5�&C�yv�
���]_�D���:��h�T%�q7�I��M��U�b7���-˻&B?2��7��À�{���o�8eԮ��y�}4J�݇�ut��	��E��;x8�V������wM�f��H�H����"�<��R�5������f^`�����Ug�x�ջVo�8�#�]���1�
�[���KpXX�wF���l4�����Q�Y�6�Kٔ����J����o}my��E|"�o���̓o8�U�UYÃ��PܫO���9���?@ط�h�%����1�&���&�M�5څE�%/#�$��0_.�3Zfh�o��H��@�E'b˦l��Cw+y��}$FNn��5�j�`d@jߋ{�Ŕ�ߢ�g��ͭ?��BHI�����r���S���Nvq�㚻��=�ug��] ��@����?³d��m��ѨO���[�����X�/t*�73��Z5��HNd��;s�|�6�p�Ԥ�	�����j����Uv@i�AqA@�^�m_�5�����kboq�}VPu��yp��%]X���	E�^<�4)Q/�����ȫ�X��E��@�w�b#q=���aj*h��mF���Y��>h4������v����_[� q�����Nw��	b*����h[dMH\1�b8%0��L.BT���=� �{�ou�c���]��U�<�IF�
���6�ۊ�z�,���^B��,SxB���"�TK��h�]�kpj5�cಧ���ŀ�'�_=��[��<�xb�=�-��-+�`�P�4��n<)yZt��@�;�V�V�����4� �<�p�G��?s?s"�?�î��p�{L�Do�e�@��^�c�c�B=��vB����<߼��+�L�G}�|��f�R�}��br��(#Sl�"c�c�x,QE�ws�x���i�77�4ʤƌ���(���'y���P@W�����⭂{$-�QK�W�Bib�}ZKf�|����-)tj�o	����ڶ���9.MĢp�=�S�t3�rx�&(�D�2�={���^����o:F��`�J�-~�y&��=e/�����_m��R�$��H�a�y��;C�"�&�cBBh���b�[m�z�}��S)�5��	,���,�#����S�>�T��o��_�ݫ�t�n7Ԃ)���ָ��;\t���g#i-�����o/8�;ꐢ���uW�TN����p� i�8�(*�A��5kt�Յ)����<�->����I:���0t��b���K)~6\���W�5�q9�N�	�ӫ�Ym��kV�y����w�YtE��jg�u�!����Ƕ G�G�gt(�J(�ӿP�$7Z�lX�M�󡇣�ܽ`�#�i���ٮ���fb؈�Y�N|ѽ5��J�F�HGC����4aw{q�t˄��ӟMFS��w����N�:����X�;�o��i�<=��\��!�D�oH����P[��d��-Rq���ѫ�*����&yc��ح��!��q��A��������KRiE���B�
�%��-�~}T��)"�o@'2�(���Hsv<�IK�1�G��x=��H5���L�(�Z��J'�X��2�b��/@#�S�X~h�׿���𴟁����=͑���]��;�C�v�e�#m���������]��o�#oޕ��	%wBl��j��;0�p�oH�>�"�CR�Ԋ���5z���x��6�L�_�bS���XZ�.��HʢD~�3Ű`%�ww�۔�T|�:�����D(�m��j�иA�x�Dܞy��)���m/f�nY�Z�SY3�v�C0���Bw��$&������xb���s�n6ߜ�/��
��B��DES���	򯌖��xeg@�O�/o�|]��li����˗���}�<������lg1�M�p��s��X1�A���O)7+�K�ƭ<��z�=��=AN7��?ZBnQ���9rF����8���xヽ�w\�|���p�gÉK���}�.�E���b�^�?}j}���ČY�l���ʠ��@��~�N��"\@���94���w��UnZFg.����CZ_�~��SK1��v�~h�	l{fDg��j�6�f1O �z� �e�Jd��������E`fc
�܀M|u�L�NA��z֥��ڃ=H^�P�ȟ�;��G�����.�4��P�$)��A�8��TǼN��I��_J^��#E�N6�H�w��K�kΟ+�ϼ\�ʻ��bӸ� ���^��e��4G����*!E����Sl����8�����M���*@���K�Bݕ�Oc��x�J[}���m���Y�3�k�B�6����:�E$�C����dw���X���C�⻲#YP�L��jǣl�����'gr6D`k�-_���٩�V��6�SxUw��z�7d �����zѴ��R�V���9���J���"��ƂR�k	Vs�⯛��5�j�)�Y#|Sj�E��T�X˼)RO��!���2��`���;���J}&�	�(��F���b~�y���tM*o���$���Č7̮��+=�S7V���q�G0&	\�G��qTǇ��pg�)��
�����>H$h2�9�?�wm(}&jT�N0BwF:��ަ���@7L�5�'���<3��γ�6�Q��;
Oh��[�@?�m�?S�B�;!���;և1�ϙ �߯��Ľ�`aE�2(�@���>�6A:��Y��ȗϒ/�Uǈm���L@���Ï֕�u�+%��,����ú���&����(�p<�3:������=�v���j���R���(į�,3�IW2�S����Ũc�f�Ć<zZ��ܐ�~�!?%Թ]{d�Q�;O,1U�Bj��i���{������,v�Njh���W�`h^T�Vv����Ut�B��H�,aͪ��5�aHc�����9NXf��,��ۜ� �]ϰ8A|O���#�ź)�M"�U��/�ao_�����j]B��e��=�çg�&�h�r6{���{YheU�Ͱ3�h���s&�L��!�o>�M� t����3�'�/���<�[g ̅�;���Y���у6_/��+E�*B�Z����Ϻ�wSi�n���9���Si[?-�*3BZ\�쑾]�DM�6V�?��Ţ6ٻ�@���~�K��?�8���F�͈n�O�k�pS_B�4�P�����x�WP�e>�3�[:Rd���>��d%�@�m�,�s�Pe��~0B6}�%ir����lE�ip�'�"��]�5$��ou�j;�PTcx��$%%Ο����żX�����x��9�Q�;��� (���`�f4�xԦ}�ӹ�mD�Q�X�^����kP"�?hk���i�M���d�o�GjH�N�sKm�p|�oz�V�=��M�oݩ����`
��j����S��+,��b��Y��h���=/}�xK�PG�(P�+�ޝ#��� o��+�I��?4ÖN�A�Z�'�P�^��F$�2��s�Ka�wL ��V����� N����oG/tc�����ʖ������H\}`�X�rW�����Z���1�*�D�D��Oo���n-b��z)%ޤ�P��!'���6�r��č�>��L{�����!5{� ��c�"Ԍu`�<.,�R�ݣ���uqJ.pMV?�m�Ix+�;ӹw�e[�ͷ���[*�z��nv�S
��Ү��rb��'7�4�U�0�I�nܾn,LAH���iG�w�m�:0�D�aA�`ɘeY���g�hعx���[��b�֞]l9@���vZfI~<\���'�'K�RkT}��Nh���g�Ҍv��zE,�8���>��D��<�U��d(i�"��Ǵ���C4��G��M���n���P��c|���^�@H�E�wj���^)����?E�@U�ґ����Pr�j<(r�a�c����!�c���.� 4h��bnt�fL��Z�z�Aɢ|>`�	�������%.撹�J�;`�nQ=#v�+�_c��6y��z��>e Q�*n�Qם�o2�w�d"Ё9%���t$�P�A-b5{��]5V�3e=�[���F�G�I" ��'vv�tqcK����2QԻc,��S�_�c�G<���N�E��Qߤx�*���Xr9;�R�p��.��e}��0q�P&��w!$Ph�&�R�g���Zs^�1��-Czeku8��~�x*��CM��n#�w-��/��~2�ܖ�sZ�%�H�LM��~i� �êۓT	N��}i�HG�Ud�ql��6��XJ1P�wǧ[1i��5f��j��FLN쌜N�b����e��n��Xz�Vr�FX��{��+42��*�m��K288-d��b���5�mX��v�j��`;{Ej�ϧ^���:2�$�� ��.��7�� k���N�Q�<8f�~�� ��d�q���I����0�Q���8߮E����VΒ!�i�Z'C%����@)��V�KjҌ`��	������T)��(�\�����+���m	�i�)�տCC�^��N�)eU��<wјY�Y��uIzZ�$�,ȢlK5���:�	��������4����d�!"�Q#�C�Q1�v�fqɝ��"��RY�fQ<��
�wT�|lL<���ƨ|f=�h$9��bb�CC��®�㟾ME�C�?�6��2d���45��tHЦ�sv2q	�m�����@�R�Z=Z���0�N�l���6l�|��������L�n���q[�,JR/?�.(0����婨z���}�:i����6X�ɠD���h��T�Z��{�\��Ht�8&������=fw 1���5K���]���0����a���M=T��}���	Y��[��?�̇-�<���S�9	T*�'>f҅�<w������#a���*����@�I;Y[�''G	���ҷPL*]a�l�����r�����5PT�Is�����n�������S�4�,J��y�}j<S������Z�"��ٽ/y�Ζ�R��b�:� ��.���v;|B��C���}X$�Uu�Lo\Tp���1t�?�f���bUG�%)3iõ����B~�Z3�f~9!�A��e�-��xٶ��W+ b����٧��.'���¹�oU�(�P�����҆t��9�DD�㎕��,�$���.Ur�迃�aI%,�4�G�0�<'Qi�(��q��c��{(��Epv%�ī0�_z��8\�tz����V���E��Rۃ�A��ER+X��W&��)�N�9�lRt+u�lߏ��S�07�gS�d"%�����pyO˵����V��d_�uw�GQ�p�}kǉ%{�sJ�Z��G/yLڱ�v�6�>�6�"��Krc��%�y�o�����֡������"�����lU�F��1��B�z�m��U�{�8�J�Y�4U��U'ы+����g˵;bZ-�TW��=��.WS]���_�
o��D���`�e/�ښ�<����؊̞���́o	���NaI ����nrN�?ڨ��Ld��w�WD*$�Jc��n���D;M�ҙ"�q�&�rw2��s�G�Jn�ߍH}?�r��!���_���$;��bF��b����������S��V�(^P,ڎ~c�gyуN�}��X<�"�:VZR��7���9�HVI-��<A�D�e�\�/�kF��j�ۙp��Q�G���� ���m`�8)_͘IwLQ��]m�s�m,D��[L���H�d�@�@+���0d��jC���&�3\�.K�
]5�%<륛r��;�'pjU^ �pg�m��۾xN^�����n�*�ӦM�U�M�d��װ?l7d�9��u!�A�1��y\�هt�A���2J'�u��$(� Y)̤��/��YN�w�QℿW/�G���K��v��*�&:�/�z��-�����&�R?$%�e��qHɓW�1P%_��APA6�L�.J_��R`?�	�?�`G�Q�C�-Y�T�N��݆�~���"p{� į�Q��>�9��ɟ�D�+�x��})MgO��#����1�;G�iOT�+��_q�cg��7W�oڽ�l�4&���;N�ؑϷ���m��g�Pv��ʍ4�i���1�� S��uXl�������a�@ۏ����o/��Ѽ-���*�>�G;F�,�,ˆ���8j_�SՏP�>��`p���Ԓ�@
����9}��h��c�� �{��O2M�%C�f�D�z�E�a@��p��F&w8P�k,���v#�~�6-�u����� �B�gY��t�GR~�e�_�o(p�K�;�A�g({T��J���Y��¸K�>ѭ(���=mɔ]�g�p�W�J{]Ptz�x<P����u�k@?�{�ئ����=����L�y!�:޻�
e!�a�������~��NS����&��0 �ksfq%v�Ԙ3�&g&2��-��,�|��A_;-z��NV����k+HRM^��������a^��)R�f�d��*s6'�T��Ŧ�e�t�&�ۄ�-B���o������`���a�^�#��J���,��F9��7b��9�/՞|��k��9�J�G(R�(u���l����X��0kNP�.`҉�۴�=}�S[�D���Zp8�;x�ݲ=
�QI2�B�WOd�+�("�{���|�Sy�y%p��]m�K�:]^���d�~J�����]g����u
y����b-����7�d�K���A�s�0*a<H�m�Xp���ޡ��RJkBL��Π�<��_2P�^䪆i��/Ur��8��8Kˤ"�zDB`�8��-v�WU5Iu�)>V�趙�02�U֩�f"McUN�T�T�JP��V�΢��i���s�>+
�;^��#�0�Q�RRV���}*����	�S�E;�zA�<;ml�:�A$�X���C��m�i����E1R��]��`Č��oE)���>\���N��*?)��-���Z*���0��f��a�@�iw�D��T԰����E�� d�� wC�F�.�f8'/C�c,7(��S�C'�ql�Ǝ�|����V�A���.�Q?Rs�;�Rw;�bj�#�4���,(�E��A�zp#�e����	�*U� ���>���cs�[d�ϊ}�S�߃�(���W��r�R�8v�^�6W���Q52h�Ǻ�b�03E+g���i!s��o%����ߴ�? h�Z�n���ã��"?s	]`�~b�,:�Ä	_��"w�]`� ����cz��!� ]Tp�i�f�F������8rO�M���*�o/܍�g]Ʌz�����-�AB�dt�q>?�^��D��r��Bo!��A��햃���5�RG�)/�l�
aѱ�X��4�!�Է���][�����+���(Y��>Ԙ�|�^�a��
�!��L�C��	���'W���n	�ECIl f��+��;܈M��%����T�)��hs�SQ�V�X7�����/�V��f;-��ս4��:��*��
��,֡�S<�k����O;����K;"�36�u�1�i*H����B�)���L��s�DC�ɏ 
9S+�ܖ�9� �x�Û&���}W<[� �iV���1���r)P��L���Be$����ǖ75W�ȑ#���LI���^m�k/��@Q~
 �-)W���ˊ�R��oY���ٰ
��jE��kc���MD�1-�pJ�ϋNȨue2��yd�iJ������^h�6�x`�"�R��9�/6�k���� ��r0�--��}��t��܀�ICjS=��*}p�:�Y�j���P��R������Ǿ8��^�a�y�B0\�@'2��
ұ���wq��9c�Y�I�^dP���0�p�"���p�4|�'�����O��n�&���	����{;�lR��]`���maD0�*�2���C�ک!� �Ď@*`GR�DU练*��){7�a*g�kВ������L�7G�?��.M7�e	%�0M͉�K�j��]�\��/�,����ċ����c��&�C+5Ț�o-�����8�{L�{9J��)��e��گ�O��πN*��[am�s���j[�f�٤b�H��O ���#n�;�`y���;���a����X��!�M:wj��΁�4���_����D�T���$	�N�,ӵ��U�a�����H��4��̮s̼17Hx��Q�UnJHb�b��9�{���ӥ�j�@�x�I_V0�)s���TZB�j��=vM�
o?-\+/<�>� ���������a��Ȍ=�@ ��-�Y_��e��h���?Ś���G"=�9��܋�Ԑ41�#��0F`�C�M���B�a�;A�E@X{�R���o��|��Gӽ}EG"����r����8	J�-�w�fd������B+�|Á��p!9s7��h��v�t�(U�ӗ�a�q��V%W�����f�R���;y�Ds��)�)���1/�N��dm-��ER8�G^��R�u4��H���sٖ���e9���;y�s�!��_j��������a"�gT�$+��'òjj5���`���k^�R�D8w	h�AJ�M$X�>�?��G/�+j��<ý^M\�^wX���Hn~�8��h�������YxJ|�姿��5R���P��es�@!�U�ہ����E�����G���Ё9;ں$8�{��=�%��)�Y�&[6��\��d���0���Tw�:�"{�;�l)�@�(-��7�$��L�f߇ZQ�V�wWn/?�0WG���m���A��U�h���M^�<ɂ�u<|���bvwsu����>q�uA�e�2��+h��۳w�#
#&��cZ)�DΟ�ϩ
~���%�8Fݥ1=��#�T�E;�Ʀ	>���ZE:�R|�W.iQYDK)�Y�(
$�^��KM	���6�Т���	��F㨕��7�<z����>��Z%}zN���`'H����x�l��7{�x�zh�jBtR���H_�+�_�mJX�Q�(��{�(�_�/MT�����p>����}fmq\�$VK��H�["��A�҈o�k��Cok��itVe~(������J(������´9å�)	Z���J�����8��(jUG!�T���R�X�;�l���IA�Ì�#���3}�S�ZqtHn��	}+!R��<R����ly杸uS�,=�}��>ŉ���2:T���~o�=��I>�̮�.�{pSx�~P�7Z`W#�e�Z|Jcă��^[�ďߖ=���wU�F>4�VK)��\��`�ݹ����)Dr���TV�D�k��w�Ǜ̝��Rb��2 ��� <_$, �	��3�A��}L`d�W�K��>K�}�q��w]uw�E�����epZtG��b��zm�@`�-����O�Oj�,w(�ӇM�L|�F�-��m��e�E��.�5�s����d	�x/|��)^����X�
u<ˋ��f�_7�]�:�o�9k�N!��q�XeTps#A����VD��R�6:�wYl��M���nR�j��1����(����u>�!���	�[��P��`�+'#-ea2�{�V��ʑ�m�~\��sq��a)���N��{�+T� �э���w�"6�� �6���E��`폼.��jե0���*̀��$O�Ȫ�L���Pf��T�<���ڴ�J���lݯ�n���6>���O�'Y+Jt�6�B�ĹJ 0HΆ�9dmS���`%��`AdT�x���^U�&$mx�l9yn+&A,~���D�Kذh��z�A�`�5�X}=����ש�7�ꌝ8�"��pD#�%���4�����YJ�\1�+����xh*�i�t����U��\��ݍ���*�_uҐ)�/��:��a�;u�h7e�T��8k[�d�;�t��w�����A[�:��yR5�v�߁wS�T5���uca��M�f �	RDv"[�?��$Z7�Vъ@]����g��-�,&�*,�N|��I:�a��:S&B>���׺#�8�,�����\'��)>� �S��{ 1�v�a]���r�ev�P�t���W2ߙ�q/i���I�U��`[# ���Eϵ�Jn�}�y��0��Q�`���ݞ0�����-<�6��`#��e��(�H*2��{�.3��tAj�AK���v�aofSڟ7ITغ��}��¹�ɡ! \ f����{~Q�uE�AR��*O�s3�q2Q��<;�?���6� �W��XI��,G%��ROS��0����&.>����#��dC��3z��p��������ޓ'�5���q�S}���Q���A3�4¿���ب���#�����gCs�^\��C�w�6%{��)�C$r="��B�ɁL�CR�t��Tr?�2�b:�� HLC�rd�~3��]�$x<.��tt��,��,��n u�x"B������������2�zVڄ�����j��<,�ɩ.���,����F�vA���T�5��7��b���\c�����_?�,B���B�8�"1;�j	�"�v���2ύ��;aA��5HP�N�i�D����MȲ��_mc,�.�<\6&�v� �-�j<���8&�ok|�=���^����F�d]T������/��%Y��Xc2���o�juD2��	Iw���"-pB���l-��<���^�v������("Y�ypXu J�"x�X#h�/��YDZ����r^꿸��R���f"�%V)4���<�!�6l�V_eN��H[v��Q��hG����W���`����$u�w<����dy�Z���5ܘ҈���l��𫑾�������ƨ=�6=��Q�[��8�L���<*�ME�j�ad���Ѩ��Q� �o|p��Xx����r��HD��4��,���"%���-�h���%��4��l�u�GqX�J���ِ���!q�8�:K��Z���.}Ug�N�=�*7셑E�]VY,����gr"g�48i��z��E���$�p����b���/��Z��@:�A;����S,lW��[�^x��8�
"B�r����
9�����0�y����E�^��+�-BiH��[#��O'���K�8��$w$~��RZ�V�sj�)�GD�`�Z/<�X��b��K���2,)�������:y��HH�<V�/(Y�R�aІ�Nv�aN��-���$
�s����jG,�d�{6��]b�&�}Sf�e�Wĩh�kʌUW6��g8+D6�m=���P�>��'Ī:KDyb�˴N�n�!�+ҿ��,�Db�C15���C X����CI�s����������]�$1��}��"O>�n� �%賂x�f�~�U�K�G�2��U��ra��D��҂k���Y:��jEh6i0��AM�%�Hmx�W��Wή|�e�J[�8jzǦ��mwu8 E�1����sB]$(N
�M��oq�B�Y���#��:턓F�����J��sK!#��S�C��rG �
˾(��cW�Jsm(Ny���?1�,���fdy��-Ta����< ���� �Vx��j���|���ňH+��Mr�Q�]��9��h��߽�	^J�g�R^�F0I�[a@�[%��i�/�;s�~�!60wˢ�V�1�ώ�7����B @Q�]�ہ�S�
���ne�*2���^\9��WaGԺE����{=tQaI�4�?�q�[�paXȉ��5�}T=�A���n���R�
��o�ƍ! �c�;Å��ߎ>�	W,��(Kk�E�Aj�܂�ĝ'���ƤI�n?���Ӝ.L}�Co^+u6G�����ͺ&<����uV/aRT���3����6�,w.��ig�M�t	|.q+���Cٿ��t��4��|�`�D�㢇�
+�!C,��<zTB�;��4��?��X�+��f����E�m�Y�E�N%)����,e�ؼ��"�����K����	�Qp�3�+�R���vrI��i��n5Y+��m�;{6|2���β����هI,d RV�����Z�����,ܩF�7���IDb�i����mp[ �W�U�������[���u�r��贓?ԅ��fh&I�!��b_���t�����k�(��&i.���l`nD�/ט1���2m'kt�m<MgN�f�����0&�ӵ�������O�m>�θ�~҈��0�����fI�,4Z�{�b:���<�蝈n�|�Gɼn�j�C��*��ڠ�L���v4VJ����!��qk��^������rC�0�j���M���%�����(�K��<c�+M�+�����%P�������BKb{�Z:J~��%PL�1t�z�{�R�ԋ�k��� y�4�`	�g֜d�(����b��M���
�4i����٦��k*d��aec��ƫ1����G��d)"St3!}.�IXsT�4�$F=�fZ��U�B[8��4���+ !��b��%.%y����y������������-~�y�%��8�*S-*5�P~O#��|��Z�X�&L�2g�����ĩ���&�Rd>��~��}�����Qu{;	����:����,D����~��8 ��#jܓ���J֤j�!��O���x�ż�k'B?�x"���_'+�X�Ac`�g����ܻ����f�U������,��+��d���Y��F�K��kbl��Kf��*]�q�e
e�d�0�	��ꫳ8&�&A�0]���Ǵ42�pr��\���|f�t_�wK��l�f�a �	�1%�����E��
��P�dJ/�����r���r�̀Y����+��$ą�е��8���,�z�t[~1"%�_j��[��5z��w(T�׫��.���
>���ә*�M�B1�r�8E#�D� ?���z���B���n����,8�-���������l�x���:=f����}\k%S8s"O*eXN�����)�`Go?�����T�~�ƿ���c��*B�,�K��P`&v�٫!bb$Ϲ@��O?������V�1�9Ù� �Ϣ�F�Y״-��V��m�^j��`��k��*йm{�U�Z 
iM�2׽C��a�3׋�6S'I��P2�+�r�H�z {/�D�@8a��u�i�u����T�j�����B��h�k����h���n��9�2݇�����!dMF��������β�
۬uTm� dïӎ��Ȏ������˒v�2)c��F�KY�[s��%�kbm{������ƿ#'a���KeD��^o@�� �|Q��woU�g�vd�d1}�#w7��*%�������_�WT��.m�@βY.u��j�1� ��#��w�g��!�#����~�M^K3%X�q�Z�f��U�.B�a,69߬�+L�{�xC�J�2���r��Q���=��=��Mm3�X.�D���iG/������TH���{Ng|ye�I�, ��D��r�����d�"p*j���"�t&K�'�>�%�����mKrZ�ƀ8�� E���\hK��������_Ҵ��¦���Q�r�6��n�3���zs>(��p�Z��t�%��g%��s5�u�?^��$�G����Kӡ���n���([b+�eYnEc^��W���4yi�W��"��;~u ��
� �ꚍw�c��2���T�Ik;;2��l�i��w��fM7`kuDpݬ(����B3d��sncћ!�����a�}LN��P]\��򏭾'�g�u��[UQ�q��i�cy���~S[��Z}�:�N$i�O�|�-P�
�t����JǪa���"���8���v��u�J � �l�bs�'�F{l@�W��gvy`Z�@�1�^�B�ۗ$4��ʒ�=�]�7@�R�q�Ԙ0d��B� #���a��!�#�Q��a+�l��yݲ<:��g�Үq�D��N|%��������W��-���hw�AȇR��7,~�Mw�^��i��!ۣ�) i�tt��c�/����(d�{�Q���xw�J����.�q~��!VK嘞�:��N��D�F������di]�� ��ԇc���T,����g��vCЍ�8�J���q�v���`�sQ�<�_��6��.�̫m��D�r<������&��V�B�h��
*�H�Pm@U"�ҏ��h��Cpdqw�;�����;U�3� ]e�;v���6ܸ�����K��w[��߾Tͮv��������U�y�-���(G��a �0�"h2f���$)����%�'�cn$�'�x��k3�D�|��fd��d�����R'�nY�6;׮? ����e�H�L�5����v*�^)q���<e�7�Ŋ����R� \��}�N����+4OlM��B���ݸ[��V���n��8���⬶��@~�����9���+�J4�����������0��iC��We�<���4B@z�^!j(��rJG�1���׎�UM��}?zؠmO�e����o�	Bn��ڕ E8��z�Yg�֣GD��]�?"8�fH�����c���kT������`�ｉ�Aw��8i|!kŔ^q:>�`���俠te�D,��&��)��ڪi�0]���w����J���ob�Wl��+I)E�`���2�@�t'�`ږidfQ�N���z�,�.v�o{��L�aZ ��#��Y5�MZ�_�j����Sՠ�����t��H�^��m�����u�9X[��.����ʗjө"m�J���~-���:�b���]�B��S|9j�C�7?:wbޝk�N
���'�F *����U�Ǉ�,��.Xj_P*�9��vL�|7�p��.�.G�Id�c7�Q���EV�O�b��4��921�"S�����E�?[��}8���f�����VMd����FB_g���ܲ�U=J4�Yd�r���fB���#&��7s/%��Ћ�X�h^�������pi��������!n=P����|ϊv1�\���_ib�SeHO�=d�v�Z�e�y�B������8)⌱9el�o3��ǟ�w-���Q����0\B���V?����e�k�����kaH����*���W0RO���.w����Z������	�'�m����v����x�x5Q��Mg	������B��@<�Gt.���,N�ˢqc����4.*M���U���r^`u�Uy���V��1����v�{Z�o�o���9y�V����3��X�i�&:C�R���gY�f�����1sy���`�ɋn9�z��]��4T�.��.��I�v�g�;6�2*
%L
�4�B�I�`���c�ٓM/�yd�|i��cC�����g 7N���`d=������2�\�`^�3��x�@���>�J�O���7��(Q�R�<��lO���Ӣܵ�H�nI������@!�r���Wl/'��~U0KW��p���ix��]�^W�΋��鏰�,� �1��2H�c���q��!O�	[����G��=��io�F�ߓ���E>l@±p�%��[+��2�?�s�%�ic.4�5q���W��P3TSt�o�R=�+�E`<��~X�XrS��۶.>8͠��.Y�{��c��?��� O� k�$5��vj�xW�%������}3�9�0>ޓ��F���0�w�UX}b�غOj���.���l�C]�H�O�$��kz�u�ܴiѪ`�]���>w�B�
�Y��ѽ�JQ_�� �HC'��L�Qu�g(��յ�t�DK�
�����Gb��Q߇��nӎ<(̝�ٶY�D'ָ�%���0�����R#\�yv��Ƙ����C��q~M����~%�h�uh(qmb��N?D���5T�`Zen��S)o+�~�J,�jݕ��m���7�����8���
�y��i��ӻ����%�Dg�<�0NVH�عQ!g[7D`F'u�ĵ��������9�PƢ2�t=�e���I#NH:�*߂SR��T�b�x������O?�
���FY�s~Ҟ=:ݜ���@z���.&(���B(@����br>��2�O��0��y?��D!X���4F���gm��!�� ���Bעo�d��m*�L�LȢEQ�2�G#�?����:����׸��d�I#���(ţ�%��$�%jE�h���Hf�=�{zG`+
/�Ý<�M0�p�B�m9��V@ܧ��#��b�1�ї�2����7�?��uOH���ӫ���ȵ�� �y*H����˓ΕYX_��֞O��Ɏ�R���A勀�:��j����p�L�u��U�x������<��!��5F�g������Q���)v�Q1Sx_nעj��#�Zb��h����I��Ӎ��uH�M}�J�(}ɇ'F��d���u�-/��탊���{c|�mJ�a��x���#����K���ts�6p� u�4[�#N�L��O�O���iB4]� y{L�� U���G�c��|��_���K	�ЬL;���A�n��F3E��HK�kmo�$Z)���0F���7X�,02����t9"��F�M�ud	l�鉝N^<�q�k6R#��ݝ�MX�)���"D��
f4��\4V��ֶ�5o!Q���;j�<�:n�Ҡ��x�U����9$���?C:b�z���-�����OG�����:�u��Ĳ\^��������Ze�Y����4bD�փK;7�V'�CUs��l0�P8$�g����f�aG�Z!�s��U{����X�d�>��5���s�̴K�4��Hh���F:2$t�4���n/�؋�¬�!A^�~OG�L$iC�����zQ�Y��%�_��3��՗��K�5��k�ԩ3e?��^+�Ҥ��k�Y���z��X�f�����C��#0���Y&*���D6�2xg���	l��4�p.Sʻ��\OT�R�ނ0s�ڮ��h���$��+�ѿp�����N���$E�rv�������L/1	\��"���}��SܩdX��g�p�:X,�[�����H�wZ��o��ΐ}�{�}�<����2�1�������_�A��j��Q��W쁠#/_����U7���зԲZ{1E����`�8�S�n_ˮ�I�˄pwHz��
"_���G��q�˱NR��7��o�/�p���n�G��B�e?j*���5Q�?"��T��n�jk.�[Y���牦�"��7�5i�|j������^_衞"��m>wm��/"l|�t�{��Qe EU�F�o�j���{�*�gP����
�eŹ1��u����}2�����F��I�lu*J<n֔�U����ol1�0�9�q@`�5��ҨʸƐ��Z��� (���U>�+���p=��H��u�T39���|I��q���t�$�!��Xy_(7����HiJ��W;�{�ֿ-���s�r���KAsj���\R{��Tؠ!I�J3]>�&�Hq��ж�s�-#O4}�Lz(���d4d]�S������w�]Ŋ�貈�g;�]�z7/�w����"�TKk�*�傢�uf #���믦sH���9�6��F��;�i�W���k�_�{�,��
h�J���JvfdU�s�TN~%��fm�؇��ti�@kM(�k� �s��ъ�9����B��4�	VU8N�1��[j��o�{p�p�+_�͖��b��b��Ŋ��]$y��:뾡�����Q���z� g#�P��L]�O�K6���%��N,h�'�q4��PJ����]�v-�>m��א"�|y�v�خ��5��kN�V�+F�Sp����D��T�%u^^(,bHŎ�?��=��Ǚ6���5ݘ {z����	ܓ��w�}Ш�X�Dki����}��8�B�R�cn�mya��lO�IJXԹ|ې�
,rN��,�D�%��l4B����.�8,��8�طؠ�%��v+�H$�lM�#lN� ��#���Aa��pQ�^�4~��SI�p]�O��*s�uL���/����He��.�׃�8���<�1�C6��ŌǗ�����m-�7P@W��@˵�����߇�Mҝ�@��!\�����Lgֿ��C��Mv�v7%�K��͢���D$�7�G�&��N�z�o��	�7)��~���d��A�P˙c!�����F_���ϫ|����&4HN�@@oki�&qM&;��s �x��̼ 
^+��#6
a��Ǉ��X(vN/$_ȉ���+���ߺb6I��M'rN��j2{�c�=�����@��Wj���;Y6�_��R�h�������Jm��x��Ciν���\��S�"�*8o�pk���
�uU�n.@CM���<���ʤ�'9�T��'��������GYJ�,��Jp�����r�/,�8��x"���D��ݹʾv��Z��"ʱ�ӗ�`Bbz�Xw�̫������q���ǖɝdoqj!�M(��j��9/6a}��\{�yxNϺ��f���)C��"TP���P0[�ݪ<�����F��{����.n�FOØ[���j�e	������F��^сF[�j����E.t�Su}��"�':x��@[�󽔡�ɿ�0����E�n/�_d�=�n�N���"�E��H�� �9C��#�����|D��ʣ}y!ʢ�
rr6��V5�:�'��Sݒ1wZJCknZ(�O�X��j����Ѥ�	��ڑQ������������u�L�Ws����m�%�☛0b���sZ�8�;NΏ����E

����%JN�8&�6u�_t%_����-���o�!;� ]}HJ&��[ʣH`Qŀ��9���+�9i0+�	}���^��7"�m�n~ZO`C��bSoe�#>�Ȉq�<���vv�����/"��&6qJ�$�[%h���(�*/A��L�����L�^?�@Gz��ST>�p��2�N��Y�GV�>�K��/j�dCPB|�}���2�)��o��$�&���!�^N�,�����W�w�C�[�+�o�(�V���\w�og��y�Ŗ���8G�;;DcA�Z�O
�p��E!~���2���n76�Ɲ8�&߯lA���XL͐?,�U�v�Yj��W����Q��%<m�X���\7*��22ͪ1m;���p���tcK/[	zO���wAdH�Z��$�i�w�
UPn����g�o������39����O����j!xQx�a�l�C���A�����H�s�_ham\p�O@��cI�k��VH��rQ�&�`��@q閾,����ߒ�UR�n�IH~-D�,u�$7|�n��-����+��r��	�;c��p�ܸ���;J����W����� %��?})���/y�K��D�A�8���T�[ ���
��9�Y6��<OJ�ƊP�*�	�^3kxWv���+��l.RC��t�!&�(��ǹb�>od"<O�Ze"��I�<�����̑v�.��^u�#�r`��?B��R�!(���مT�gn)�>3�q�I��:6ݐ]�/?%;V&�h:9x�tA��c]���\+Z���iB��ҧY�Jږ`�W�����*��c	Rk0F����J��N���d�����,��W��8<sj�$���|:'���z]�E�f�j�
�"��Ē�1ƫ��`C�v2&�X�=0-֫xՙ4���ׁ{!0O,?�,|�SP�x� Xu�~2C��Dm�Z��h�Aɺ�ߚ
%q�]�=0�鄴�lь�Q��|�K����������]�Nx��*�A�P(x>�)��}��)ˣ�y�5���(|�r���h�m\�!�[��lם@N~W��6�͍b����va���^ SF+������h!ӧ��(�;��U�%E���`[���~A1$��M�_�b����W����<��N@M��V��]��pу�O��/UaFyC�2���~�@vf�C��d��c��������Z��R�w��xB\<��e̾�Q������Z��s��2Q�[N5\\�C���!��q�>���b�m�sV��eo%����xy�{*7P}�l9 �+w�e�����(|�Lǅ�3�����U56n�$�����3Q{=��$�Pp(��#B��j�v�/iRd_?�bi4XT!p��(����F9XM,=J�V��_�	Y�>�W��3 ��tlt]���蜇'Y�3��	=*�Ɂ�V;�B���Id��` � �(�GM3q�	1>�_�.���B��25G ���=u��9�tG�Xj���#H Yj">�LO{#*�>��CG��CxK���W�]����`Cd��Z����[|?[Rvˠ2J�j��m��P�v��-�8F��aF�˹K����R�d7����I�Ov('����i�y� s���fL���*ɇ�%��Q��a�JX�������3+@��P��]���ʈ^7��ސԑ^	�̦�]ǣ���u��9�3+x���EaX�����N&)!�'�F�'x{��̣Q5}N��=�h6ݹ���h��>*��:%k�'���`7 �f���d�˻ϟݨ���|�3�r�cOM(mo�%�o#��Ӛ��H���H��������-6-���?ibU�i0.4Մ�g���}<G͠�%Tm����WBb�I9z��g)\��}�?�i��2m�����,�K�'ˎ�(�2�~N�j�+�Ӳ<���T�����`�"��o�Mf��ǮH�����)`35���8=�{���.̽�m���n��V2��rw�!�cU 9(Yx\"�P���.��'�l��ֳ�c
��w�-q�~i�9%�,��ZȤ�s�����ۜ�&Z������p�fm9^ Ҭ�H;�Q�. L�.fz�=2�(����Piy~r���B����#��f����i��ry!ҵ���Ϥϣ5c�w>"z�$�j�#R��"��-��Ə�^8�J��]�vQ�h�HA��{H�Tݯ�h����Z���s%\ҡ��=��H$���V�z.�#���c��@�����r���H��g���
%�>0}�F�ſ-����o�x�дĥ@�f�����G87�R�z�ۿY_�M�a@�n�U�h�rE�HXI�z~�,]�6��B��� ��_���p*���G�kV�����\���ĵA������]�ȁ��;
����M�t���� p�k�qp�vӿԥ������*�u�>������zYC�x��t�J2'P|s�L�7�ooۛi���ֺ������I�ʰ&ꄰnm+Qz_`���!n���1���v)>yC���M1�Q*ǲ�gፄ{&nO��}��ւK�X��͓��0Y"8��(�J�gL��!#�»UQ�:u�G)��{rLLW���ۜ��7v괶�,����h�:(����5�X����&)6A(J��y;,L:���&h�sB�0;�Ǖs�V7��-�����뷘۪-��l���%m��W�ѥ�;gR�Y�hW� /�Q^��34��	��T����Η@���[>�
@)Dm0�TOm�ts�*���6�������W����#����S� RM���'�fru��^W$�J�m�<N2A�(���S�z=tڙu�9lP홐���օ]~��6����H���yL4bI��Ԓ)O�8����`7IB��P���:)w�� �Y�_�����F�aav�h���*�?X��dG2�����6�]��2' ʠ�>�8�M*R��{nu��O.�v�C-y�����N��&o�BF{���'x8O%\��L)_/
6���?�7�0s��nPA��Q��*���r#�(�Y�Z#'/��>������H�B�r��_�Y-��#�~�.���ه�u�S�H�d�t����z9�kd|V�)���t��r@��έ��8վQ�m�ܰf�� *�,�Ӄb�/>wij��S��3��`tZ4�1{��ЎL��{�����7�c3�V�I�Y�!SHn58;��5��u�t��o��h��Y����O�p%(�1g����/���f9�MK|I�#��|�S�۞S�Ƃ����Y��H�q\6�ED��pf�M(�Gj�>��I��Iե�Z�ظa8�YK������lT�K|!��9�ڀo%3�3�4��
x\��_^-��[ùt|b� �p���3T����
}l��|K���dp�K)��f_W��`h/�J%:W����U�f���3�D܉8J>���"�����t2��mC��Йμ��X<��HQ@��&/h��m
gF��L�
���
�����1���*��r��]c�a����Q6��0Zj��k���t����%v�{i{�q+mn4��G��H:�#X�cb[��q^�����[��l������sF�+a�u��9i�DP��B�Qf<CC�4W�A0�lg�D�N�
D�����s�����]���I>�B����<{\V,����]^qG�:8G��o��U�H��A�)�Vi��x>���1|�#/�
���9/�K{H9�_�M"�t�a����FeX� ��@�a�i@Y��W�Sy+V_�9b����I�a�8u�ˏ��L&w2^l��[�>�%g�[sFN�s�\���o'u"�ϛ����Y�G4!��s1��������E��7b����[�Ev�\*:y��KW��}�7�	����Ou�%�'?K��2����Iչ	�Y�a�L���$�=mɞl߂�����k����(#�����b�{�\gӟ��.|���e��v��� 2(o��9���o�C�ld�%�&_�v�4�O�e6%�I`ݟ�������
�@f��YJ�|c�~����n��^�y��׵	t{�!���TC��8��(B�y�`Ԓg��{	�?���Ί�
��%��X���j� ��Y�dt�cj(��(�8�N��6�n����ы����_pU1����W6�h�S���[����L5�����bJo}��7&�CPw�^��0����LY?{GQ����ĴFI�4;T��$O��T ,��D�q�vc>���%=�^q�n��2[W�� .7f�}��pM�N�ǆ����ǹ͍ 2P\��^�eT-c9d���z3}�<h��zgQ��w��
�`������*P�g}jK��k	*�E�v���(����M��r��*#�����-E�-J�@�~	V˵Q�S`)E��=��B�d��p0��ӈ�E����y�"UN$��c깜�N��(�-�Z�2d���h��uZM�1�A����dYOBlj�}��p��Ɔc��o�@�7��)@�#���N��~ϹGҾG� �M8���.pmT�#'��D�=WGܸRRg�)l�\���?}�8�eC��S��Y�_�P@_���?2��Nu���|���`;�zy�R�C�b=AM�Pr���X�?6�yf�='��\/�aT�ّy��"������
0Vв�����7��X�I�h��X2�7Z�2�qڹ����g����i���w�;	Q�eH�v+ݤ��O������؛�{��`iyU'F̞֨�l��5`�8�(�ė1����8wv��E�����l �QE/b��i}�?6c�h���0�!C�;h=�;���BP�ę��u��Չod�x��~���d��0��C�=x�8x6����r��� �.���V��
	�,��a%^���l=���&��Ȱ�})t� �y��	��;�c�b���ԅ�v�k�����s�Ǉ[7.�Xc4�:����>_��j�P78 x�h��`� wh܋3o��L=-��A��#1��F ���Է(���d��~v���<:"?xn��P:4-|��N94^��ԃ�.�^��!*�����1jv��X�p��;�-�\���7��4��$3�=9�	�XP=��Q��r�(��j�ɑE������I�\�"�u\q�~�=�fD=�p:2�BG�j�������1�ܰh�e! Y�C�C���ž�4u��|�%��_?�˪�>�WP`\��8�Nt�L��7�-q8�k�L/gO���Uf?�#�2�Q�[6I�w�&i԰��.[��w�CC���r�5����NT]��	r�4&����`/��g�:��Q��}��Zݪ�|��~f-�&��/XG�?�0���̛g�E�}���!�G7!�rV5��=�/>Ⱦk/R>Eݴ�\,C�K��R�bC�Cg|N�Y�����ӵ�0=�h.֥�7���zJ`S�x����S�'�6߈���ڡD)���B� 匯��Q7�?����	�~Twm��ҋ��[P�iA� 6^|{�0ɯ"f�'���%0�7ox�����v���H��I�*A�V:,=*v7e@�(���k���i�֎����KF^�c�Ij��祉]9�����$=�/����rY�{�[ʁ�s2���9AM-����-�)d�V�Ԗ�웆P������R�N��N�wݵ�T���#�u���:�9��HE�}�aH�)6�u�L������'���.�j��Zy Ux%�'�P6�B�ݒ�Qمj�q=J�1X�����>2̒�&����������������\CV
���5;0�D'6��AT�(n4�S>�i�2�#��{1٥��!L�5%W��j&G��VV��|�X�ܮ�Uu��aP�4�g]�St)T,>�
ld����IE���MRk��"v�3XYy�i�z$���r�%��r������¬���JM��4e��d,���zy{V?-�!ST}��jtk��~S�;�T�!�)�u,.���;/���ӑ�Y �AB5��S/��J���ab �s1��\HZmo�/����EG$��tt������e?��Y(��L��f�"ï��!���#�&�}��UV���&�o�A  �D�3�T1��Oٌ��?Z�c 8�V�%�S���-�l?�.&"ra���m��#��N��`�g!����!?TYQ*���53H|ֻTҟUwj҃EF ���a�Xq��Ћ��;����Wt�nKj�Í_+�����IB���:Po<�c!���}��[�d�;�p�烿+�v�D�R�<x89����>����6{�>�d�oxBwXۢE'�Ek��wܞ�K> ��ٙ��Ⱥ�����L�݇q����}���Ϭ����ȷ��=�ijqn�9���]�o@���P�$Xܗ�ČX{�� w���S��U�e�,�^-n�ȴ�*z�;<xV�V{ER��.ʠ;�*�Y�oWT��$����f6|���
�������xh�`��o'Y�.\��fd�Ate�X���֢E\�o�q����Dh����p|0L�`�L[����o/{t�������\�����h�3y��C��x*�5��Jzj

��S�⧛T�A1`v`bM���b/Pg���?��u��5�Ż�昡=�/ ��Ք?���V3nZ��ls�񽝉�p�Ȉv���;�r�ϸ�Q^��Mf�Nu,�ʓ������Hoi�o�;�U�aD?�\�(ևju�3�ϧ�V���{���R�?>��y�|�P��y��.c�;z��dSE-�qE��_�ZB+�y�ld�{�!&���|��`�l��N��	D9ض��\3�ji�"=x���b�&4F���p��9��:mIw�r�A<�
M+9�(������/xc�����.�� �KF#O��jS.d�=FR�`ŵS\# A+�
���T����s����*��0K+qa��q^ͽ�_	�g�.�&��_I@!�dNAE���>GYQ S�>ы`Cq���^9��&���ߥ*����<K�u�����wyr:��v']�@X&�p��eb@F�@�s��~��̷U������d��I��f�x�)�l��f&`Vw��X����(�'�D�Y��	Zb�eל�`$^�����4�A�����a�HW����V��i��O-YpD�1�b�����7�hm֓�����趛����VP�Bk�����S@M-h�����'s5k�������SQ[/��ah� {3���a�MZK��N���M�2
b%�T	�bW ��>#4Y#:[q���"�X�KAȎL�
�$�W��Ĭ��XS�?�O�M��-����ԡM�R�����6�����u�k��`ܢզ7�3K��y�~Ƌ�|�L+��q�Lĝjfk<�
���q8w��-{mJi"Q�ʮxI.}2$�(�����#��]:�:�|��ܵ=8a#s���]0�S��Vc%ԥD%��/yg$�9Ê�s[�T���A�$�S�� $�CS(m ��e�Ҝ�H���qu��цX��L�>f!+��)��f~�K��:��4*`�X�5̣D�Kiu8���9
n�h���gZ�16�� P�K������><\�k5�C�&�.�+"��K��k�B%e�n+�ў�I���&��q�~�p� DO�|Fg�'}{�R{m�C����ݢ�qFT]�ɡ������.	F��T�|�����m���}uŭ��f��p�nk5��\�@��+��}[�j�@��LL�I�q
>g�w�7��mř���HT{T�@�X�/���:k�c'=�| ��m]�	�_�o3[Yj��A�p��� ���t~�u�@է���F����G�k��!u�6�D�D����>�դ�t������e�S�ႀ�}��[��0�Ej��������"��t�A<�7�%(���F6��4=�p���Jq���"��	�/�&�B���Z	�{����ã�u/K��q�3&F�O�7�̷��IP���$���<�fx ���X!ed�:������������.��I0��P�N*�T�q�f���𲔱�.65��ESze�pt����ɢ2�,͈Y�sw���?�� W�e�PE27R����Z�Q��(`1%��O"����ڶ^Ӈ�����-/y����!K1��`$����̞���sw@%_����f_H�kJ"��L<;B��!��U�>����٬L�"��OȈc����-��#�*)^n����o���� /���q�:qۇm��_�T�h��@;�=����]o�(�� ���r�`�zxpz�ϑS�NwTR�8^!�Շ򱰘��&L�ʬh�K#�n49ʿ#��U�yH�=�G�4�C�'hn��?��\�9ż�C���=�����Z��&�N�����#��=�Ĩ��Ù���� Mmr�8=�b3��k�ޡ6�Q4��CR��5�.S���@%�
2�|6���
�y<γC&���� 
��JXZ�?����B�D�؅,�ID>J,�ɤ�����-�4�Q.a��?�_>K�H���t������?��5	�wC��8?z��r,��x�=���@�(jH�n/��E����
��G������W�}���Z��UJ +쩍U�VH��%�����'��|����b�B�H05+�˨{�T���	v��K��z��1j��.6ڱ��<|G/�y�^��~,�h�UI�����ԒCqr,���j x�8��n��"P� db�Z�!e'������@8 Q�������ŵL`h�?�^�B��BN�X*����
�N�?�U� vCS%7=�@���#PmZ����(�$��z��75`�:�ߦ��a��67���k^G�%��:\d�V<o��d�?Z?���Fn�<?*N�l�ńi	���k�@�p#�$ȼ)n���t�uwp�qu{�
��9�n�ń,mUm���
"'N��'.@�tI&�A�ʕ�����)�biG��{�����g�Z��W,x�7 ��X�Y,Yc>|3��ǟ���,���n
.҇���Ѫ���
��]GJjZb֡X����Fz���>����'�W��g�]fjp�^A���5T
>V�B��Ѳ\p#���i0>|M{G-k��9,2�-���ۚ��N�tfA)(�	A3}��ΫC��|&��5p�o i)w�*=��M��b���9�T�|�#Ŏ�*Ͼ�����"��Y3s/�`�r��-���k��Z��k����ࡈ�4T�=?��Rb��g
�R�u��F�lsr�DC��W#W�UY���<l�v$ԋ���g��f)�]�,��ϟ�iڱ�]�LR�1�3�G�V��?�<�]D�]���uۆF�Y��%���DVn��\ �=��r*!��f�8'Ej�`C�a`�ݴ�:f�
^
혝Rq�^׌��gM�����@�����7�}W�x9�L�����K�G*#8x�{�,�𣇼�����ڌ�+�IUgv�pv��=��0��ǾUx�^�^��`F�;;(�&�������m���?��!�ᡟ���'�����W�P���w��W�J��'c[���џ�5�-5��u�-g��@����:FC�g3i
��'�'�(<�6�x�J���|��1!}�m�=L���~Sl;�����������y�~�tT�	˵��?TnzB缾���� *W�3�a�%�����X�H��Q7���s���+����e'�)p�S+O����}9ĕk�1"8m�xa	�y�f���Cs9oÊR'%B&7�;탅���蟍<lb&Z����O�m�}>��9�k�%�5��1��$���S����Lh@����Y�1s��ti�H4l�i,�w��O�:�C�j5FiJ2�ub�u�!�kl��Iѕ�%������P���-e-���EylX�)a�Գ^jů�0KN�1��
z�#�δ����E�;`��:?��*&W<�\K�Z&*�;I��\�JҤ��&D��ᵮ-�'_�u�5nf5�!��~��r��Ol˩�?�h��2[\����t�~�ы�����Tla��1�_w�_{"`J�+��ܽ��0F�f�wr{~e:�۩���j4����I=f3�I���V���]�P4G���\��DqK��z�^(�N�m���-l��>C�L��&�
����<����DJ���
)��
:��Uԣ�Oo((�sa�����mD5�W�!�X�U�L�)|���-+��eW��j'������(�9[�Ň�^�sq��u��6u�*_oT�|Z��&�d�f��+ܲ�?	Z峄J����ܕߑ�J:�gu��V�ϯ�Dۍŉ�(�Z,�59�:
���s�����.��!q����yb��A��l�=��i�$Q�T�Ȱ���9m�J -���O��6��~�� �ys����ر�!�-��A)���`�2�=p51��h�t�
�h�x�����9��|G�0��]~)�����]��
4�E�,]1�N��A�V�IN�"P1,�|��D�+@i��%#�5Ƣ)x�y�q��g6O�-c3'�(�w�*���s&����AE-s?���Fb̸ x��η�a[�o�[��� ���ڨ��ƫUՈs�i.���LܛT�b%5IUwN�	�$�x�i��K0t:R7ˈX��8�a+��O�<0^/�ّ)���Q3�B[�g�a��] �9o��HT�&��W��=jԥ~���V����ʃ$��R��{1�&AUk���;dk+��z�6�Y3�4F�\��F�>}!fu�e*����R���_����q��z7�R��NQ`�U��c��&��Y�ڍ��S	�z����%�#<���^>h�ib���C匃5Ԛ�l��sL�+�u��".0��fI�sgtwX�%�TQRd�'���K�e�aKL��$}�W�T������R������=G�l2��%�e-,�ZN}\N\4��*�kbDu�+SHR*5l|��;�����!�qt���,��A�RJV@���˻*%��H�Ъd���#��ʗ@F�>�
�����G��O������[/<3���	M����-�:9�9~zv)�0��<+�����4f`����E!/������	t]/�����c�Q����|���EN�UV�8��L�`�nk�[��A�eq��ن>��K��uةk�%��:D�&8���af����8���~��/NTT�ܩ&���r�I�HW}�s�3��G�� \M���'c>���%\���ә�l���r,�mxi�O�մ-���ys�pvZ;<Փ�qe�x�(0�M��ov�M��!��c�h��}�1�g��}��vk�ꜝC�K�4��қK��ƈTcV�sP��3�X�?c��m̶�s$��>)�v_���SSq�V6G���&� ,��i%uC�*�O'J��s�ڽ�#6���ck�S���R���V0���3��j�EMEM��n/��9rI�ʭS�=������J�'~U#��^���m�v{y_���=�L�ᖼ�2i$�5&(��1Җ~_����.L��"���Qkm��+���_=�+m��9Ya0k��E���y�Vn�.�1�Yุ��9b�ٳټ�����`�޿h�J�=�������w�gx�g��j�4P<\
�/�A���j���k��Y��z�L��y\�^_r�(~�:-cT���"�
ӑP2ڳ�:Chq���I�7�36PDo=x��HU���Da��\6ΔgV��L�h��J+��g˅��:>�pJ�'@��)�dsp�*6U?<�:O[Q@L+=�q�֠�:��N�|��Gӊ'%�fbh�@�9�p)�KDX�������e��i��9��<��1�Q�4~ �m�}�F͘�%Y�r6�x~i{�U}`:{�L�S���E՛4��:��4B�n���Ҿfy|ٟ<����6aN�Cл�w�_�&��3��!\�wYȷ�&�	�%�zO�χي�*]h�׌�FV`��=���(���R�f��bg9u�[��fj��a�oo���������&�I��窲5�-�{W���C�q{#vu��o�Ct|Hcίw0�_��~ӂK�Ł�A��>����.��ࣼ���� O�7�h�����4��n�e�m� ������ιY�W�[����s��}����r�P�C^�-��t8�ݮ�2/P�%�Z�~�sY[~#C)7!u�.<��k��=�@��m�@m����yj�K�d���r�!*I�g�gȭӼ -�c�Q�ɒ���ʿ��T\���j�ZK���9Mp�fB���>Al|�R����ބ� ;.�I���1���h��<��<9��S�J����2-�S��KOyT��V��ݧ.����ُB���gg�������/� �E|���R��8�4{� {p��^�PǗ�xu����3(�.���U�?u(����v�_�4D$��I���347C�a{��,�I1��ԫD��Y�॰������+5c�}��>Z�����Đ\*�܌XoæE�9%�=B���n�n��!2�{���eA�����=�e�+�����\*"t���-5b�;N��U:;H� ��%7x���:�8��4/u��F�W��[t��j%H�l���ma$��s��Ԋqr�N�I彾y	�Q�|-�@��LLn��&\Ȯ�@P�;����u�uT�i��|	:�a�dt�)�mv��A.<�C[N�,�I�%�2ް����υIK�d,=�����-�q.*��?�#qcu�
�9��b�d�%�8��Z���u� ?{�h=W=@��%�CX��6�p�>Vj����3��k�]0�C"Mw��lr�V�#�V8�]�{$X-Ub!�$M���"!��C�U�4����/�B���)��o�bd϶\�G
�WH �	d�ٳ��R��I��]1�܆���z���,��؎s�	��^��K|�u�}��I)y���{X�o�C]	8b��q��½c� ����R�@d�N������*b����*w��*��܌/�K���(`�iV�\���ꚱ�"E�����.�I�����)�n0�+�E�4w��$!�Rh��;�f�7 ����[��Ws�9�����3��O`3fv�2]�tL�%F*r�� .�~�C���n��2��RF�����`���ç��I $��Hg�1��cnΤ1����R�cE*
����˧����u0�aiz'�/�-4Kp/����?���|�B�Eõ�J!�ok�{�A��{F]%�bU
���c\uQ��_���*ֺV�8�śwaωyT��:tꮸG	"�ܽ�,�a��| ��|\
�v>������`��LY�-���4���{Em/ֆ��>�it�(=�o-(�0���R�t)���{��=˭"ˤ@E�c��!Z��&p���K7r��U��5�*��9�H���~��5�9]�ɺ��^�lYbf�F������-�JP���}/��^���j�������yd��b{^�Se>@�{o���ƍhG�NS�6c��},�y�I���d�z�$���e1��	Ql��!��[`�����;Qv��ȈW&�o��z�5Dmp%Q�o��_�F�a}D&���,#�j@���k��Ig��;t-�������U{���&Y��z�DN�5<��[{o�P߽���{GwP.�@4�>=�H}�<��;ᨤ'�ĵ��78�Z{�5���ZJ}�����"_�􀂣bف��k2�Р�d�����4H�P�J�d�T	E����ͦ�3�!6z<.�dYv����4S9�M,�gc�ۭ�iֺ�+�7�Lbc�U'��Gv�(�ȉ�2�����Q�1�wx�IJn��I���������/��AG��f��(z��Y�Ɗ��'Dr�k^��+���t�)QCo����x���� �̘V��d���c���ۜ��1��Z]̪�vXx_���9RJ(����$�t�ԧ쓁O�(�j����01���L�b�	M� )�-���������#�wf*tw��%��X�������kK�~��Y�j����#��Bi��
����(�����������jH�i��ߌC�7��b`p��#pܟa!*�I8�^�����鲎ycY�!!봅�tY��na��@�Ay~J��'g_�c$&�[�xG�+�2}95�H�b��� �B��;��k�,��`J��-�b���e�%H����	�_���k\��FdJ��9g�0����k��F�͌���t�O�H�8Y6`ѿy����(�R��^y��
7��!n`���	������=���R�v�&I��.r�I�[8Ӧ"3�� �m��!^v~�M�����7��U7�F�1�^{�����.1�w�Z�>�cl�c���.۫AH��M��Y����Ve�}/i�����9Sǐ�U����G|c���B�AU5�Ռ�]���V�ׂ�b����r�CG����^����"t�"g"U۪�↹h��:�Lw96\��X��~9��'�J�C+��L~����f9]q���vG��l�e� a����9k�!u�7� �Z�e^\4����5[��s(*�Zy�����_��y�@�4�R;�F�����K�r4�`�(�&�s�QQ�D4o����>�D��z�4o�y�%2�\15'a�u`_��+#�ưG��a��˱�<)5I0��,x�2A$$���jM��~�; �9L7:]z�$�� ��}͠D��A$�v��lg�)/r �@�F�*�I[��x�=��6�����#�$�GJ�Mv����ʹg��n��4z+���Sf������ ���b���hg�������ϙ�\|י�s}s�|=�[ķz?i�_��7(��R$�]�3�*5=M���T�k���aq����D���o7�v�[H�O���e'�V��<�\�I���Sy���i�Hʥ)��EnHO������%�޸�`�V����vQ�Q�V��lΧh�i(H)�"���D3Eg�4��4��h�F7��լ��J��]�l5%��=4�W�d�AG�x�p�k�l+>?�L�[����v���	4�"�)\.I�1�I�}���y ���/*!�ꇐ��@`K��>�aQ&{?��DV��D$�(6��-������:���R� ~��/�'��J!ݖ�G�5�}L����Yh�ns��g#�E��e�=����_������_6�{��\$�j����ӕ�J�&��ֱn
(��%��au��I@L����
�����_V_�h��Q�ۦF��.�7l�$PÛ�M0��
����@^=�H��D���-�k�� <	Q@�8���s�h+3O�������"�rY;��G�Ac'8Trϴ_ Gh�J�7$q3Q Ov��.�"Ƿ��_w#��s�g)���9�=��
@�Y��L�h��;����dj��CH�"ݝ;y��٤��ØөK�t"	��^e�!��/���E�on�#H;{ ����-3�h�#�cw�c��u�#H~}�IZ9j�֭CoɊ�'��e�g ��ɖ�S�q<�~�萫D��c>#ᚏZ�Ɯ�.MXe���(�/�Qp䪐G`9�O�<��˘��;�&��N�ur}[e�҈���YC�����H�a�p/gJZ]��1�kak!��e_C���@1��"������ˀ�f~ˤ�O����{o��a\@"�(�T�� �H�V����Ir��G�.ՅV�G��b��7�����nP����8y��Z~�O��c �ý����̐Z[ Ş}y��\$�/���hW��"a.�Λ�UX��N�.\�Ny���8�B ��.=̅J$�'h�T�5�vE*^A �4���>���/�]��{Π���^�� �`��}1:���%������ar��b�b�m��Q�\�?9�BbKq���FgX�N�!m���K?H�+��h+p`/��P�mt�Ҥ��TV��Е�>���N��R�Ȯ־b�����h��D|z�)!H顭���Uf��>�R���ƔQ��Q�Y(�̐��\��ߍ�������A-m�)g��s�MW��b䉩vP,���7
� ���H���/�� fɤ�Wǥ�?����YC��:�c�kQ{�j�<���ѐ��ט�ٮ�A�Eϱ���4��Z0Z�	��K�E���tRU ����.3euc�D� ��?O��uҢ{;Z/��4cՔ��J�(��X���t@�|g���3ڀK�s�&�y��"_.O��B��?s������zm�r{��HȾ�7x�+1��ڼ�3{��h��	ߓ&PS�.�Q�K]쐵�L��}�}cW��E�ro��]k�mp�<�Y�5^�GТ71Hc%Q\���}`�1�L�lp��DW+s�'f�+�4'	n���*��0a�9� ��ΝQ/�Đ�5�u��(Kj.�\m�"9U�ؤ����'c� ��6���r�ƌ"��c���}�����hNz��d���{�Nq�q�z��z�Gb(������X����<򆨤e����� WM�"����g
e��G�K	ײ����Z��t�N2�,���	E���P�ݎ�r�r�l5�_qt����d�4����Fq�Z�Ϫ�0�a��<�>���1�($�3(E��Y_�,�zx�=!w��bIε6��#�S8z"{������dݯa������n�h�5W\��?O�/��7��p�)ם���w��u2k���s�%|�CCcl�y
�
�F^B�@҉�筜j3��<xC���vq�mo�S__5r�b�c�k~{Z��%�^_���䁦i{#n�%\z�=h����6�r��K�6;�r��R�,�liKRxn�E��x�7S���<_}�0K=N�����1sP����xl���ϔ>����G��	��{t���23n�>���T]��Ы�o�=5U�tnMV��[�
�>���������m�%w�@��5���bx���@�u�����oJR6L3(��`jV��(��c��R�E�K?)�'{�Հ���4{��sJ��t���9�CT�)w�YCN��xyϦB*&+2�����i*<�$*�F����G,�����_?�K� �^��g"k��K�3E^!Z�5�E���=R�H������m`^�tv�VEg|V]�3�eD[�Xۀ�#�4򆌭D�u��k���ְ
<�@�=��C�C��2a�h`�ֹ	GO@�*�cQ��W����/�?��RX��(RW�n@�@�+� �q`+yXĕь���-�~+9L�Շ(����G	�:������0#��(鮑2QFw��Wm��H��1�4jx8�?)?7�Ջ(C�Z���N`�4m����y�D��+"�n� �����*�߿oe�
��Eac�H#^��!�Ų=y�8��7*	�~O�?c��Lj����K�d��#
�� MF0���J�7.��0R����ouD�dR!�j���i'��\\�f'��	s߰G/z<
��
s*��G^#�7���1s�X���u���24�&�g�f�<r����a�G��g٭@�Q�)�!I{L�OJ�UQͣЦ�)��%�L�P�.ڈ�J}y�?���F���O��2j�7#n;��	�����wm~6�7L);�Nya�~�y�U2�� Z��V
T?�N�=}	�m����d�j<�n�3��H�t\*�H�6ښo:�Ig��R��E�3�y���O)���g����y�$i $�'}y9T�M�fZI��� ��o�1b�xFq$�ϴi��/}W�6s�4���6O9q\�������&���$�J�	��U��u!�d���38%wT鏕��Gkꮳ��9���O3��e߸��N�����v�ݰ�}�[ơťX�bz(Pf����Ȕ->�e�G!L��/;�Sj�Di�J83r���L$�.$ ���*1�q[1݀�1~$�)����=�#��]��z܆����X�MC���7 b������3jw>��賳����Z5o� }�7�F�`��q=�s�c��rH05��aJ��.���.S[��ez��x�ݺ�/ԅ����L
�V���s�9�h��Fi2Mɖ;�BM��w�����m�c��'�8����~�f Z��x��I�1U&^�#�ƤFw�*5^ e���,�����D�C�w)`�-�?���d^�.�~Y��}Y>%�X�BIÂ�:�5��V��t��G�2�Q��M��h�����B�lӑ[��%��(�kvc��d��f�ɼ .s�0�j��c&�@�IB����RQ ��o� ��)�ԓ�jA7�HC[&B�e'��6���{���9�a¥�\�a�;l2�m���Ϣ܊Q�I| ��
����$�̐�!�Dn�I#ahu��r���/��5\���w���7~m��nP�Q�sDp��VsA	��43x�C����O�+�G��DG��4���j.������O��Lu��)Q�l�셺t�j4i�a��aͨN��MY/b�{�&�k�<��H�ot�/'����if}sL�X�]ޓw	A>���(J3P=�iN�;P�v>��d���<K
��iΚW�E�#��W;C�u�߶�*_9ŷ�^���Y��w�|Ը�j�sY$T_JU_<hp8t:	�{�u�7%�T�v����]�X���w��PO�����Y�}E�[��s�V����6>T1;7�A�?
}�AE�P���9X�w\/[�T؅m�{����w4t���h��e����2uk#g[�ѝ��,�W�RV�d~!b�#���ea�z�ݳ�c
c�]���-6f�dػ��5�}�
�	���/�m����͝����2��_Y����j�3W�y��w�@6�k;-]��B<Nk��㷝�_`������
9D�PU��a�J�EF����h�`�
��憫8��x��ղD<Bּ2�Z�Ǧ-�V ^Pzs�k�_� /.x�+WIΏc1�{��2B�����48���;fk:�g��N����X��}AZ�X���	l���}[�=:��p�|�Ǥ%��w��~���2r��>��rB]�=o7�R0�˵	&)�o|sG�BC\��������эG0���k@��԰G7R���ZV!��'X*K�"�b�<"6	��g%��z��{ʲi���@r�?��sx�Q
����t��	��q�5�Hsu��U� �n4C�t�l�9;��>��5l���\l�5�7��E�w�s+B`��1��ǌt񜐣}��(�E��酷�ֵ&o �p�"��^����ab~�q��P0r�9|.���ו3�L9����-�Yn\��lń@��pӦ���$�╚�ʟ7��$2L�w��2A;�$��G2w�Si�C��êJ���K�rm֊%5vZk:��_��2T̮�`���"5.��F��R0�ya��C�Ӝw� ��h.��G�V}���2���m��H)k��S�Oo���L�v���� ��"RpX��o���p{�Y���E\�Q5TD�����?xx)tm����1�#�����]���r7	�Do���j@�m<��<���JF�e���Y\��΀�f1����>m�����Y>����ax�ݨ�H���U=�0�f��H��7ﰮ���ְ��/��+A���ed=r�V�b���ǇH�:[�CL�@��VvIo,��+�XM�
�6,F��I�	��R��m�� xǂbů4J���yj2+&�=�zMʯ)Y{G񛃐������7&�#e�l�R��;�4ʅꨄ=A0�ch5�����T��־*�^����b��=���%�a�'G�#��E�b8y�dڴ
Z��Ǣ�D����i���]�2f2���3���QM@Fӷ+���?ֿ�b֔P-e�}��ڱ�b��M�V #]��TjR��۩mX�J�b�hI�eh2\�O�#+2�������כ޳�d�=x���U�\-������|�i��*"�l���fā�C'}����~Į�����/M�.�N�&������}�!Y�ɏ9��Z�𘟱ުۈ�w�Bd�����7*�5x�Oϼ��4��1�ꏢ��Nk5���!k�ˣVz��'��m�^��8�/+&���	�-k��Jk{w�AF(w���m���O�=|�;Lv>4Lb@��Sr�b������w����6*�
��>/ٟE��:��7��`IIp����Cp�k�^�L����?�7c�,�l�KV�vV>U�QR�1�&p�ֶ3N�H#P?Ap���"���g4e���!����9+��.�Xr��ܤȦ��J�q����_�t�=�1��p��0�J��X�R��÷g�ȯO������!j��[��{��1��N��o��PY��B`��5�/|�آ4��
e����\7����#mAl���ju���/d};K՗H8�[�{�^�c%>o�q����KjQ�2Q�5
/3� �i�x���ȡcכ��:�s��F���<O��ӆ��Qz��M
�[g?���������Iq35:����`��E'����nUP���LBz߱ۊe�+6햠u��)��]ՠҘI�E$6��M�G⳰e[�?9���������o_f�H������jh�S#A�,'�މ-���CF����G���Wi�}������g�M**Y���x�U�7����VʇA�e�G�e��Zw�ĶD/Jӵ�� 8����+ω1V���^�M�*�E��T�-z�?z��Y��Av>e��	�� ��D��sv�����àV��]���!a�*������w�?�v�u5�~���J�|�%���f5>r<&f*֑�&��һ�����Q�XR���E�/�3^?�\�F',�8�QR�V(3纣$��U�
ʠ:�^�|�'o��Ggz'ˮ��~�L��.NN֑!x���9��;�۬���/�Lk���B�����5��Y� �D��5Ȥ��SۦY4ƽ��.��@�dδ4XQy�U*���ą���c\w��-��S��pݜ��W� _xZ�z OBbbk�����)R����?��M$����}��������T�#!~�|��� ��y�.�H�x:W8��';$x���41/bٔ��gf���� ߰��K�5L�1��d�uU�Y�70��]�ʑ�%�{e7 ��`_.�D�<Jz���dz}��{��J�4(<	�gR��K���0H�^(�����E��P�1F�Ͽb��}��g��뫹6"��$��0���xO����v�W�5��:t�v�ֆ�nѹ��hw�F\*�x 
��ywP�70Ie��=pq3z��������_�EFt���y3ǅ�V\�jPx���^�>��ޒG ~���j
L�L���o��J�KO� MC/���5�rD�I#�_)�v_\����`�������?��� sx�a�x�4bӉ��+ ������	eb��{�NR\!F)M���T[��9�LSc����0�BF�[x�]1�#o��D�ȏ�t�-2h���8YR��� ��Gw����
�jqf�d�6�}�A2��8�{��K�c��T5�vb�Rk�/��^��r��|j�&�?D9���Ø�A_k�`e�{�	�Ɋ?O{jm���Q}�\Z�5<�Mt�x)n�I ��A�^pw ��S�a�A�"B�>�=�.S0���7T�����8�,J��(���	g*#q����Gd �}�pf�@m�n��ddeOفM�p�sr���=��!�[~ۗ"l9�o͎�idj!R�/�:���y�U��.�%I�� `!_z�D�ә���o_sNH��Ȋ�������Xgh��j�!f����{u��w��I�(F��l������TJ��]��j�aHA�c}��2޹4���[�.�1�7Ȩ'>�nM*�6��̦� �MV��寏1;�+��P���[n!#�G�\P�)���ab,t����N�t`��h����3��
����J������S� ��A��9ؑXW|�e��#�nט�@�^�]��g��Qo��(�8=����|�DjM�� ���2\%㢘xa��ҳ��\�Ms|X�*$��F(mH�t�b��(�jwZ1*�q~�w�_�Z�q�Jy��¨��<NU6�ؗb��8]����K(��A5��f���<���zD�%R%ɑ���nA��( Vy�$�c�d��ʎΗ�R��ʆզ��aO�㑅/	J듽AU+ک��V�$�Y����]8���U�?T�E�u�F����z��^��-�fA�x�yh���s@uh4H�;Q����.�N~��-��˼%��[n���e��%�9�8�%A*�v��*���t�r��g{6#��Ͷ���\��;.���.&��v���m�Z��1��*���E�CM3Ρ��K�o�D�b�gg焉d�#YaS��7E珙�V�A�5�M�+��P�\�V��6RJ⎊�1K�:��x댙�%u�U�j�^�o�������h
 !�d@�PpK��i9�8�}��?��^W]Yu���?��v�o�D|���T�)�-b��|�H�ͽ���N$x�[.�
�Y.�*yu�k��4�$���Z�~$�Q*�E~�ߘ�U�l�2,�91�XZ��;7���{��A*yÒ����:���j?���$y�/�T%�8A+pt����VGy���;��eα��Bx˔�M��TN��"�	�d�V�kF�o�f�!.*H��ʟ���0�����=�@�p�4W�"��/2usi3C;'�������z�~�H�v��	'q`ۻ}
.���7%Q O�r	K�{�%��{�M���k��L{�ǯ'T��M�HZ
T���,����vK��L]8k�����P- �QbB��ȳk4�-ۚP�����7����]M��b2yOt��u�2�W\xQ��;Ney6B�2����P�#9Z?Th�B���Y�@��������qY��	
t�=���ߔ����m���l(`�Z0 O<I��1k �ςҎ�.�����v`D��Ir0��g)C1;l�Cw�{x�/P⹉�Օ^�N�^k("jIkYӗ���b�)��Z�K�B6���(�p�D���S[$B�=�
��N����~/V�<��3�x�:zKJ!z����5t��I���!Wk�m��"��]��ǡHi%�*����*����>���mY.R�7��o#��6L�����ARɧ,��$Q��Ё��~�g�x���#V�~��`^^���7�縃y%zU�[{�h9��iw5�r��lI��O��)��XS�wJ�o�i>[j��������t�����@q~F!@Am]c�D�}O`���a�����2�����R�X��+i-�LH�.�0sJ`���h�x�&�8
�-d���N�#�:JD���Hf/4/y������]+)8�T��E���G���=�O��@�A�	��a�=�-��fxZA�����v_�6�{_�����U�_�ӆj�iЪ�zry����(�U��WD��]���D�\��Xx'$oUȟ}]���m@��촓7�)�z_�)ج[S'.��k�&Z8ba�!���`[ �
��/�߈��)���_G��^�
}�a0y����lwo�\��������?���K �X�B��J	�����#�-[�^��Xv]S�ǖo�-�Tw8}��?9��Pb�ZT��L���A���a�Ok[X�I��1��v{�y��L���5����f(:�|/�MaRf&Fӵ����WЪ���Cͻ��o�^�L�u1v�'��R�3��8n[�r�	��o�(��ލ�d)Z[�c�֣\��a�B˱ܖ �bj���˲�0�ͺc�8B�Z7e��W"e��3u����:v;��$��_X����9��?_�2ƨ��c��P�؋���w��������"
`�0_���3�k8�֮O.�U�7��D��E,��Y]��@�;.�9iK�i@n( �|�h�0��X��T�-X�o�y����*��=a��!���*��uԐ1�j���nY�/��m2��.����6Q-�O8�<?9{�H��)>�T�E�B��w����a:.%�C� ��W5�֝��oF��f�i_���1m�D�\Fz7'����8Ɠ\�w�X�p��$�br�I�שB_���=	H�����h�uWe]t�6c�v-ev�~���]\�X�l�����&4�+�*y�}�Q���,!�^<��9��>�3��Y �ޠ��N�K\��KԄJ�F��.��]5��W MD�c�>��Poџ�iL� �Օ�0�dT֤�@T�݁�Ť�@��T�J.�g�r9�v�9�d���G5�HM	���H�6֭jy�1	)�;�.���Ks��h�$�t�8��v��JcHa���FA	�$�:�LL2����0X_j�Bp�?4SH��#7�=5�������=�������{�U������ق+�=���Ee����<f[��{.C��N¥|���"�#�=S��[��)�X�r�l�F��:D����y����u׍Pѹ&��ޖ�����v�NO�ͼ��CK���B��h�����n�6��f�Η򡧝vE�g�xŌ=��YI��~��XE��/�BTF��ݚ�d��#�;ۗ�bY�p�/�Р�`�Bf1$��`%��>�u��[���U�&�1��@C����?^�U���~*�6��⫉+0Z��{`2O���ud����8�@�dj)�����?�M~rh�ؐ��g\�x^K2�e�> -�6�v�L��JmF��"�ᓲ��~���S���!2�?�:dp�?Y8��J�WME�)ߋ*�dV�R�*��NϞ�ZQ�M��Iw�	�	�XP!ΰIN/�K�g�O���*UA�CM�,�6i졷s�F�1��F��tˍd��a��F�T
�څ-����Uˮ���[���f�f;L�j;�h�x>��(b�u��ֺ�ɦ��t�V��s|�UY��������ޠȥ�}�!��_S7sD�U����jv���j�`�a�s�t��C�
˨���"��\sN�	���?�Ů%$j�J�R�����v��y�f�a���2/[$������9��f��)__8�_�]&
�_�sg�ʖ�*�/��dV��(K�n������E[l��j� N8������?�% ����J)�9�<L��]���V�-=���Ċ�9P�
�J���䶢��ƴ��M�<���m}#�0Ks�&��x�>�v�+܃۵և�X��U=����}s�:R@˯v�U���^�uh&i��DE�����$q�Z�H2���^q���]�QTn<�u쿸�ɨ�V,�um���!���������@���p�k�f������� �f���卫)�7�,� Gh��ɐVD��ǡ�He�����<3ګ6�ɶ4�?Pf�;�!����-�
v���%�W�X�� �F!�MJ�$rh�䬒�F��&��Y1��#�{'b2X7%U^�l��%G��m�&�8��"���b8�vl��P6�l����[O��7gv��WXJ��_�)�n��3p�Z����)9�Y?l-T��f��>6W�򙿕.`� n�^N~��	�
�(e,7Ȳ�_��#:!-j	��I���Q�n�'|��@S��Q��}\�}�O��pF@f'}
�Sag �9osA��b+Z�7��H�#z]�t�̿X\D���w��-��N�qޓaӫ�������M�R;�K�g]x���MKSD_��gCA�Idʡ�+` �M|���?d��{˽M�Ǆo�����'/�c��ݿ��Hə���.�ū����79�ۦ�C͐�����ܤ9f�˗͚�Rzr7����^M�������`��&{��Ս�o��6���ۈA�9�� ��b�R�� p%[�J^�ZuZ�a�>����"J���az��6�z�V5��7��RH��Y��q�)�N�ks���W>�"� �^2
��d���FRS�r|M���3˰U��BcgB�&���(3��R� y�];��t��-�V�h���s�V?�|j��B\8�@�.4��������Q%
ʀ1�sUfQ�*��!�$�3y�_����$L�M;�p�)r g�Q�ϯ�_���)��fm6��Q���_�0~��z�Ah9�o�c �^,%�-a��E�@hG��cb�����W��8q�ͪ7���;�L1Q_�.��OH�bH����QC�%��#��2���,y!Κ�|�o,aq����6���GDRS�o�I4�T�����:@�m�-���⧝z�X�����?��-X|�����f/
z�
%ӈgD��~	M�3�@�J_�&�RMw�V먳������L����mc��ʎ�L�Ɨ�/)��7TNy�P	�$ܫ-�2:��]7l�_y(��R���RV����ʍ�vm1�l-�f��q��d��PMد��$t�>ڀr;�����ϕwl��;��H��?��^��HJ1R'��Ł�{�&�b�|9�r���D��[u0��Ə Q��屿z�#�Ԁ>B(j%�(I���
00G����Ģ�&+m'�A�A�Y����F�K-��r�\5JJ�� zm��=�V�|�G8�_DBΗޔ	�z>e�p�/�mDP��|bC�C�����!�3�"}M�V�6 ����������]��Q	.=&�B7��|pc~�}��=`|���oD��>�������m�F%U��zp�����Wˊ|.}���烙�iBr��#�S������"����!�.���us]�n�K�k+.����2�7R�B�=�	�5ݤ��:�$~���5H�0�bfY�ƀZ�N̪��㠸!�Ᏸ�˸=�o��hG:��R]\9\LZ/�*7�<����(D|�Z��E����R��1�(���:b��aa�|��������m�?�A�G;�ݭ�Wg��6~m]ᚳ��1���bU�UDt-���*���&_O>Z�Z �X���q+��:m�q̑$�#�n�h J6�� iB��*��ؿ�lm����.�ϋ"��G���'����9���@��ofo^T�1[��% �ZIH�ws�s�š�0s�d��hi\��gz_2@��L������T&��Kr� V��*�bF�g�9T3�LE�J��g�Jk������(�}��FAV�8�����}����>
�F��\C��T�w�?�7F�h�rBz)�-���YI4^��}٩1���v��{B�G�ͧ�4�3��I-R� \��C��-�VBo�(&>�؎V,�����Iz���Zx�X�|P<O�shJ�C��8l�Q}�+�.#�}�R"��f�?g�+���{¦9{['0�38Ip!D���.����/�gƔ�\���j<v,8Ur+�}R4�gCjW����ؘ��-O3���l�to�Y��>���S��׿@b0�C�|I�ū1]�;/��u����ǚdu�s^-��,8�$�_��P�ś�����h�1i��M����7r�V_f������Ǳ�j��{ø��^S�UN�U��0o��c��q������[���WY����jdi��Vg��:d��bI���)�#��Ɲ��K94P�����Ufq�JA����m��mY�G���u�(k�b�k���HQ�1�4�v�Mܠ,���.o���2�ݭ������3 ]0�d �~eĬ���uo;�<:ߥa,M�B7�'��U��-�h�pɦo�T�A	g���7�Ԯ��q��rH~���G����*K�g>�AZp�J���	O���r�M�����fE]�0}�Y3l��6��mK���w���#�����j�ڷ+�����58 ϭz�0@����H$l�Z$t��Q�|��8�4/HW�>���D�sy�7D5��<�$�������lE;BA|����t�x �Wh&&�f@�v
&4��'�p�+i
�����L��"g ���9����;��#��d*�5�]�H�62��q�G�q3Q�V}f�:Fr!4���;�I���T`dd%��Uݢ���j����F�i��QL��|��x�eX�gO�}�k��w��l�S��щ���"�۾�ф=��s���_���(�+��W>ݳ79y=�_ @E��Fҿ��7��>�^N%ь�C��^�,#��k�|�(Mv�i�q�u����٧Q||�/����&� �vm;?�K���a�,�p�B*#�ת��L� ���+,Z4#�k���%T�@��%�4Ϯ����P�ܾ�U�}rK��Xt�;Ƥ��m�v�]�%��N�pd;9�t}�OЂ�3Da�Yo�
4:ؕs�����A��s+ߌuƝY��?~�yN�i�s�Q*���Q�� c{°��S��7�#1�u����R��4�қ��g�0�4K{�
�����ȅ?V`*����/)$c�Ub�����h���T1���VAДLK�(W��{�w='È3�s���|D<8��s$n&5��i�=���=l��L�oS-�p����%�O*�#�,�Ɣ"I[{��k�#�˞T�s$� �8�3�m��.��V�A㋜IL���l�	�/!k����p�L�bMF>d��N�a'(}�>��]>���Z �~��j	�����f�h5�04T����?��j�D��х��YcVMw�����T|���.�4���zE�w:�S,1�-�F��Z8��X��e����5d��x��f��w[;��#��份^�X�h3�i�p�4������@l~ql*���^Q���i�K{�î��xտ���}-&���>ct��
����]�nAŝ٦���Z�*��D���_SD�S��L��3�V����2p�[��v���T$�l�R����.�b俻��q���_�;�ɣK.j����.��O-]��}83�|�y/���_��38Pʝ���g}��:�WeAfH�79����T}���ӆ1^%��	���?SM�9Ư���&���tR�g�گ���>�ދ���qԄ���
$�C������#���)�`�W���4"�a��\�#�^wlN�p��2�`�߭vT	t>��q"�۳}="L�=)d���@1Ew���|��!`M�)�.��±4��9�@7[�lEo�Ț�L�G��<��t��ӂd�ɦ���Z��³Z-�4�&���
�bhG�R�=L{<�G��`�9��ח��a��ʟ�2[�C-8����1��L"E�}��	�:�S6��nA$m��=�r{�"B�J%-�-�Y����&���T?78�A�	ؼj�r�<z����9)�1��Pv���*�2���қ	��Ѽ�z�����;��y�X*>��?������ma�#s��T�ǫ�]��U��RЈD�[�Z22���s3�ZbH(GV��Xp��@Nn�Ϝ�XΎ�pM�#�ab�H�jY'���������=n���+�����嵓�9=�2�u��IE-uM ���Ó<�����= ��m J!��fQ�B�o���0�X3G�`��P*^4N� ���sg»o�N��rx��$�j������j�o�=��� �po�"�YF_)���wU�ݜ�R�-��*�7Oe�l��:��F~�g7���'��2�B1�qZ�����Z��lg��H�7P��V�O7���|� �,3~@f���/��Ŕ�8��+��7*��Muŏ��������(8��X�;�iΙ1V��b
������`�@�ý2�ُ#Pf��r_@`=��v�{�w�Vý��1���QJ�bB�Jҭ�3�4j�������z7Y�Y�Y"�6�S ��������;]�G���P� �x϶|�P�J"����©�{���+xY�Z��jcH6i2w�u���F[b�qs��.� f�t��%��h�r��e�c/־]GH*M�8t�O
��i���3B�wG�n�ۓ���6m����r���f���۸�.�u?�P��ԻN���+�1��,�$�/db�O�@�|� 'nhΫ�{]!�D��N>�0�\�q�H.;����*~@�7�N��H����j��F�JE��F�ީm���/!v�ϱ�e�[����l�I7�F�b�*U@p˺��#Z����mG��F��R*�蓔��"���a�+�wN5��'��ps�Z��&�-�>�r��ϭ$��	�|T�`�xO!�Cj#�ad����#pX8��/C�	�NB6h�0��بe��r'˭q@"��fi�R�YuOP<�}�,��4��ȜJ:�s�߿*���T�DQX[e[TX��I$`�KM
�9]v��&FyTo��r�mrky�ʔ/�1S;���Z�Z�+��-H�8�8���8L�S[%->8�I�h?-;,����!�"�QA�m����n~� *i���/0��۞�`;n�3�Jͺ�N�u����������]� �(�1.�S��qų�=&�j��	@p�n�GÜ�����{�u����c系_�NO����}�fR5;�k�`�ykшHB(��\��,(1񨄙L.�� �RHӪ5���{��*'L�Gŏ��pzӅUF�g�����qv����^���l���u�ޏ�S�]Ќ?8�7}�4~���0�Cm��E��j�dz��'<����+�(JþۮBM��ƿ�Ͱc���FT� Ճ�L�>���G=���o�4���c�7�4c>�K<Ƭ�i4X��qf��M���n�#'1
��I7��Gv2�?LoA�
���d�ݛE���E�MJZ>;�X6�n�Ao��wӀ�_?����}�gx��R���F�_�t
�0�>�+pvlE�1�RA�3o\��<Ҍp�w .'/K}�uG[��w�#������q�d����61;xV�ޒ��.YC3�Lh�_��+�)������-y���H�>S6'�9�Rkg��)�{�Y�&�N=d�c��WS�a�)��p��>�i�J�K�IJ{�ŕ��V��f<���&b]�O9�}b7O,X��b<Gq�c7�O ���x��@�gkޝ��D���j��X}dy�l����kK=��\\:I�Y�R����	W�4�^��]DIuR�%���1,dV��ŇԜ�w����{��*?���W#��+�-"�h�G*�M�'I���������!?n�+����(w瞰0#r51��!+;T:o�_΃u?	�;��������J����R�J��zn"ٸ+O�eZ�IX��4I'q�fXH2�u��ݲ���8��Bjɮ��4�*�C�Fҧ�ʷ��t�'d���6<�ؒXuE�C�ٵ��M]a��k���:���`Q�[E8�>��6qE��#g",5Xv�)A)�Z���P��5�=3�x��:�Щ䯩�.���w�(�q���h���"�����6ߜv3����ͣ���O���$ �;G�Uh>������|^�tncD�%+<�H�e��3&�R;C'e�ٖ���c�»
�w��*0���C��wY4�Y�ɰ�w�6�ҚR4�W�����M�К��,�?�*�%���s�!�`��.X�A!�|��~����;H4��	������0�A�^��}z����U��0�o��]��Q)B��:A��Q�֯\���UM�z�NX���}I����{ycze<'D����if��7�ZNɳ����#b+��õ�a�V�z��%�!��_i*`��Y�<�&>,I(ZW�O�^��:kyʐi [=�f@�E��Vp5�6:�j����4�ؿ�Vi��WdL9�2��1fMH|�+��Im�_�+������￪ݴ��ş����5߲G���o�"�Ii�RsQ��Uw��h�ٍ��4�l<�}V^���ʰ^KyĞרl8؏v���-_���.�0���Y'���%�C����k����cqC ��b��8�ǘ�Ԧ�]\T�|���]n�`X	Oj�����z^�,����\����'I_������U#��Z����d��pu�/}������0���f2���Ky%��F�[KH��w�&/����Fo����i�y#K�:�h�}�
O����W"z�Ȅ:�p�a<���9��LZP�
��4@m�X)��xi�a2xmx� ���"�N�
�z�~�R�t(�P=��?��]���MM��l��0�'T7����++���:�}?_�(��}�#`�X�{ڵ�����#��=�9|�#rV"XtX!5�]���0m��@S��>��V�5�>��3R�����{����Ȟ�/�t��a]��Cr3��pG���U{�Oh2��)��������C������a\�]�tD��`I}���s�N�n*�����T==Qr��J��\���B7;K�δ9�W�E�X����?��1rM_9��"J�C�cyJ���]���?��^6"p���M7GT���?�zV�F�w�u�y���&��6��\��6��d�,�%Kt�Ȁ��}�_��6�}����^��ஜ��֩(�ԩ8�k�|���X���{4�z'Os8��)�zO�	+����$z��0����P�(��U�{�K^*�&�]�ӍV����+��� ��O9Ka.Uґ���P0Nw'��{
%��d��7�Q�ӭN�5\jE��ݹ�4��|��Hb_h+q�*�\�`MҰ�>�t��o=�A��%��ҾE�r�_LL_!g�u�Wز�A�SF���r:`9ɉ�����8��ue�_HΊh]�:�<� LH�ɇ�Q�[��\|+��,�*Js� �����I�]��9&i`P��nL����Z�:v���VLn4��s���%ŋ��Nӂ�Ai_ž�a�(�A���nn�##`>�fօ�&AP��Â�����ݴ(~�y�W�2��u&'_��9[(�Ϫe�v�e�
�X��f8Ӕ"�����R)��3 ˠ��[�}�j���-��[|%�����ȡ:p��#�"�-�%�Ī��YWw�i��߈��ڦ����I=��w<D��g%���$��"��\`�)i��Z�'@`�55���v��j���ukb婃w�:�_�;�L�`�K~YQc�����ݮ�X�
T����ͫJI�t-B��Zynř��A6�$��5�����}��I5ֳf@����.X��+/	��c��6�_��=*���ul���u0��g� ӛ<�`���� ����ϪE�K��rw�QRR��ǯ�!���}����$Y���N,#��}�����t	��z�Z\�V]��EŹ.������"V�6��; ��f����߲ԊV5��m����lex�ꕜ~%o���ҫh\qo�E��a�	p�M#��5���O��A�J�A�1������1�l�4��t���SÃ��~+E(.�P�r^^LI�e�x73*a$��{��\�y̢(��Z�lfj?AC�,W�{�ޅ��.��]���[�Of���MV��2ZB�g�r`wogf5�:7��h)���K�db����^� 5S�r�&�6�����k��)�G�C%��U�]p#$����'m�ݫR4�4$��H���j�AX�O2-]�ڝ Z�voμ�W	ʏ�_~}P(fi~�{=��� :$uA�Ťh˟]��Y�\��̆�C����v�~&�� ���D�+䱈.3�Sǆ�F�x�ą�P�4$JA+�29`>������g#?i8�dg�dV�!�5b*�%�Bx��Coh!�������7���Hb�d
�
9 �r?!�1v2�r��ڱ�UĎ)�e�gړ�J	Gt�YBvu�إ�����RN;�4�y�_[
�U`�S�.[ Z�l���eE����񡄉��{����z�]��NR��R��+��Q'�$��ݥ�G6ѷ����r��۠�X\?Ѡx-��Sl��C!��B�`#���|�@�zY2��J�Au��O�}>G���n}]�幝�C����3}�E����@8��H(���?�hQ�K�������k�ż_H�7-3�il����Tx�s���m>�k{:����.j��g��d���Jכ�&CG{�#݆��źF��-M��uY0]�J��֐8c�����
v2=���B�{�.�y����&:A�@Ҟ�@fB4�	ϰP'�'�e(��l����E��]й�h@�j��K��l��"ƬǓǗ�_S���m�y�}�_�%���gj�&�M(%�݌�D�z�����t�'^WJ������&4�G���IӦ����b�R1��R�o�Pe�5{�E�Q C�n~Yb��}Q6�/0(���(iQ_!h����s ~sm8�-�M���Xd"�e.��U�H�D�|��b��aJ6�3���~~XA�l@�:N�`F��ymFV���y�����m4���ֵq����4�~�J�M�����h�~��F���u'�9��^8�Riv�jR		�'��'g�-N������z�)�j�����So0�!)`b��#[�:�Ll�A�>ȱ���vt܂�=S^wG�d�w�n;�`�gv÷�]���]�+���	�z�5;�^E!��Rӟ��]&�!�ɖ���bm����{��SX��>�A�Ji��p .��8����.�D�|ۈ��g�,v��[��.ղ]��Ũ�&�JPם�M��g�!>n��25���=���`��\�t4����ě�.W�<�.�ĪAK�]�Z�yUN� |$��٣y=2����#�����:�IQ��BՎ�R���3�\F��9Um",�pqZe��H�[�L�-�����L��F4�z�#��p}��3eJ�Y<���^�EA.]��OE���_�TV�4t�\�x��n�I��Pؼ���´�@������F�nM�7��g�#J���!>v\
�Bw̓�|�0��0�|/p�:�,�U`0 ���$��#���A��2��:p�{�n$��d*�%��5�n��+�K�A�	���l鰤��1>��GX�G��n�Sc�/��!)�(��I�EJVQT�/�E����a7�s�F�k��1�*��'��ht2an)�[�����97�l����	R"����n���a|�봎�?w�z^V�Gk�%��s~C{�*������c��mlAC6�RY穰-e:,�!�_�i0D4r����Y$�'�tCKl��H��/Z�������o����ڕc��m=�w�$x8�D1���j�[�,燡6�Ƅՙ[�ວm�0�挂���v��-5��Y�!=�|�q�i��,*�Mj�c�smJ���<J�;�|=�dp�D��Ү�;@�����X?=�٩k	�k�m���V~����f��yݫ��4���=c3��
���N�@{y<%����6J��" #^T��%,�B(�H=gRUi^����Z�%H��`�X�0j���:�6�//��A�����ͼ���Jd���߉� v�3PO�%.b�H���u#f�J�+ _�m>����gp�}�:�΁�仝����A!P@a!Ѩ�?TƄ���+Jl4/����K�sH$��P���wT�:����l�#v��*���7��(����F���䝞BZgҮ8��U��Zf�����������w��\�.���ʔ��f���M�� ����Ɲ�\7�+f��R��2(+箛l.SvFؖx���,���rX�;��b��wW�I�b�TEn��M�#��+���(�j�XH�=a��-I�) ��:�E�jv���KM�?��[���=ߡ����<�f+��ZY-�sI:EF?��*į��o�)=�4-$x9p����mqP����s/�sDJ�jf)��S���y\����H�'7���#׸=�mz�^��9#��3���7���R�)�9�a�O��;0�>�L8�Q�4r�xC� ��n���7�!Fi;�W��&�7 �;M�n��z�+nJ?�ݧ0B�����n��P��y��2}����i=����ۂ:����D�3�B9\�.��,(�~�D�����e���+_�;֪b̌�D/��PE�))pf� 9�Ɨ�$G�)��y"�=���1 n*��  �qS6��1��6<'������j䆆/���j$�M;��QI��M}�V���1��8"k�-sR�O�pO���:!܁"�k4g���@��`��X�p=�g�d�g˿P8�;����Y�p����s�0�j=o ��}6��Q"�U�`�VH����P�g�?��ׁq�בz?z�[��&��F���J�L�����O~��8������Z!�D3[��1�q��ս�A'��ؔ��[���>�~��C�C=s
���� ����`�;w{� �J���-�����O��b�q�#����p�0�Nl51GƼBrL2��k�L���4`[R��1}ْ�S�$S8A�5�����1��Yy��E*ZV��&��`�Tsn����F6BW06�{es�F��Wm�Dj���aDiN��\�����=N�i o{'��+y��%ƕq��<�� ��^//��2T����Yd�H��je��Y���YH@"���Y��N�BޛY/Y��/+sK���S�`@���<N�^�+��֚`!�Y�k���
6�רb��h�l��5��r�U$v��Cu<���1��O�7-Hu�i�^2���2 ��q$j1�
!��v���N,��籩�`wA&<V�U�\��D�>4�Vѝ�͙�Ď��h|��AЍ��Jq��4���^�X}%L�Ti���s��@1���Є�J���B^�7��O���F�T���"��4\K���=&�.��^- ��5� ���$f�ߜ��[�P�:��L�$T�7>}� �c!dn�6����H��vm�kV���i�<-K1�PZ��|�R\��	Y��{dd��v�Ct�8�W��fn��D�	d`\h�/"�ɝ���h؃n�-:��^Έ�o����ѵ�`�Tn t5-��!�L�h��(�n2�aL6=��k7�L��I�m:~G�:����k��5Ǆ 	8'э��Ey,��6 oG�m�V8��L)%�a,��|f���9�b�J��C%����.��V�Z�6��"�?P͘�CT����A�e�j���hi �2��_�	�3a	�,ew��$.���� �Sѭ��"�k��ˡД:��sO�� �8腁h -�4x���D-$?�tד��j����O��J11�4v�G�s~!�6��R�\�A���<�����cJ=Ŗ+*���&/���q�R���g�Q(�p�yc���\��-�_z���S��f��_g��U�۝�c�|�r����	���H�y׸�|zVL�����':�j��	*G#e
 ���wg5���#��wB$β�cwX�c�K���>�G�?l�DJ2r�[�/�{k黝d�c�Y��>�����P��-�1��QB-.�9Q�d�`�K%/ E�2R�J����ڎ3�,<��E��,�B��Y����"��L��v�`p�
d�ڥ���pο%�w����Kgf��Q��c~����� �n��ѹhG��Iѳ�_Ѯ��>�88kuQ'0aA&>A}M�1J:��R�=I��)����'�1�ɨZ�(!��+��7Ed�L&��D>>O��܊oKC����n�~�nM:�Y��i	���
���iԹ-�
���h��2-ь��5K�?<.N0�P����;]QfƆS�鼶jrx��Jhv�.����I��E��dwD����T�4,/�GX8w�}��B��ʑr��� 
�Nhpjo��k�.���v֝�w�-_��vδ��{3�����o��Lf�������P��Q��%x6e��$�ߒc%ܡ����Z_Z}� ���&dܚ���{�+�y(��[g}冩�RՔU�(��\c��tL�������ii�����0H�NiF��`�4���c��#�?�;�_��.�˵���-�%��2%�&��o7��ln�ُ��gևF�UM�gփ��y�-y��stW�<�4Fv.��3���)x��F9`�s����JO����1�p�����;�%�{3���ht�Q\-^�Ol�<�z��5��] ���Y�i�-�� �rե��Z�����>�#���ו��`0��X^���혨y���iB��D17ǀ,�C9�<A�t����2k�K&���QM�q��.rZ���L6T7h\�~����>a����_����L,���7�	2D?��Z�=�z��ҡw�$�G�~<�Cd�f�3�W��{b��B)]���L�i\ʖj����,��qJ�oh�~��2.L&�	D�N=�:{ (X�軅��K��e��_�/1֗�5AG�lL����;���pg�G*�Gw7�u3*�'�����̮�Y��)�#�7�|$<�JpH�p���9�-��"��*��힎[�X\�G]�eg�:����X�L3�����W>ɘ�+��a�V��ٻwa�_��*|�m"*q��6���&�G%��b�L�l��,�r�¯�Rb�b��'���	��q� P�N0G3�H�����nT�ot?�,W�vV@�+Y좻�?��D�B��ip�\A�dsd$ƞé:�r���:T�`�vS�[N0�M�ar�� ��n��R��I�-��#��年�V�o��5m���?����U{�\mYO�p���ڪ��6�kdsn����+��Rā�(�&K�+���K�`zV����W�S�?�F}���U��m=�Q��w_`[��a7�;9��3��Բ�{|E��I�C*o�q3�g�tQ�5dw��외��F�vaU���۩50�(�Ȁ��k���ǈl ~<�8B�&�F��:Ck(��&ݤ=(��$x$�&/[��n��Zҋ����'��;O�<ݴm~!jI}�1��sz�؋-�Y�
v�sT���(����ҩ���O|%���~���Y���`�9�F���n�7��;��0�8q:��#\9s2B�Q�q�o���"\܀y�0���0����I��%�%�z��-�=�\����L��H`�ݽl[C�nbY�������{_	�{Q�I�ۃKy�t�w�㷮��4��@4�6(Z����ߏH��l��j �~�5�̺�;Z(��zf~��� ��,�������4R�}��|<��d�	��^�.ϋ�r�>�oO�ܯ��{^ߎ�Ț�����j�Ȣ�����%�$|��^Olo�J���~���99�k	�$��,*W�M����;��l�GX�����wl���5��[��pX�o�XP�@��/l;[N��R%��1����+J��Dz��W�ˁT�������M���Rڦ ����y5�e�B8�U,�t�f�"����z-��h ���R��OG7k�Tqz��D9w�0��/C^��[�Q�χ��p�sJo�P���oO��׆����$Z�)�%a�Stʙ6����Sa���Ô����̔(��E\��%�`7��T����_��5�H��j�3�C`e�UG�r�ːV&����$Jё�LL��W,l�s�*�����7��+��L�����T4dh1�ލ�X��Y��F�Zc�ъ�9�z�>�^'J���5�â���x�Ӂ`j������;W�ɑӄ;�	�E�����&
�����Y}¿;��zy�T1֟1x�)����`s0���M��L���'vNb��	3��(�f��J�����S�J�_����8k��&���.c��GI��R��3�Ϫ�*Q��4�˴�k�V�����PB�Ʈ��f��Yf��ٜ��i����v,s۝��u]r���-t�w��Yۇ>tG��vS��R�WR�z�̵�TZe�c���2p�n�:Fv@rp�{S����D!�cSv�ҳ�⩝�g�[�I����M�%�����А
��u�n�8�[|r7P�{�*�Y�.].��/7�I2V�;�<`���ux�3qۍ&�K��Dg�[nM�OsK
��K¾[����^j%o��~{�A�uγ�Z���{L�#�R}T��~o�(k~W���N��?�v�8���3��Ϩ7�<���0����Z���1\��E~�Z[o�A�ȧ�F��	9�%�j
5�
����k���DW64dM���1��[�'��SI̜X�T-2��>B��1��Эo����=!��~�����>9+Uv%h�^v=���[H�qY�(�7VB>pBH�s��<a�Wܺe&��#)���E�~�ob3��k�uG���?�<ǳ������,��'�147�矚�0�[��w~�Af�Lh��h��SY�ub�+!��P�n�)���S5=?�?�o��m�+rq�꼗bg q7C'm��:gL�	O|����u8rq��@��?�����]�!��Ck[�g#����d�z��t�N#Y��t�@~����	����9<f�]�H?�[#)���a�����Ӏcp�PY��-Թ�j�=jH[L[I1Y���C�diTl~Ρ'�8$5�����Y���&go�VSfU?�����IP%o��G�j%���4�+�L�9c�(&cI��a��7W,�*g-Q�u@�3̈�4��n�G=!G�[B����������w!c�m��TynIAl%�����}�h����)q����i��֤�0};�c�D�X���~n�m0����Xp���LK��^~x"��igA�>Đ7��Ƽ��}{��7^7&��ד)ލh��4�)Q�f�=>�<m���T]j��kF /�R�#Ǭ�K�Az#*\#4'��:{�����D��mu\_���������[f$�+�}`e����A�:�[R�9��\�>�$pQbB��p'�I@�y��x�c�IS��"���˨2��NL�F/����h���y#tm���S���Q�Y�Q�Q��aH-�t�>+�8M,vyJ�|�������w�|��s�m����WNE�b���c��a����z�GLs���+0��cKB���f�/;m�B�"���δ#�؋�f�yh��X�]��+2j�]w��B/�{����Z����T�e�6Ģ��l�����u@�Z�6`���?�7k6�Q���5��TZ�e�T�0k�YoH��K���Օʕ�:���a5׼�W�L��U��؃<�"�j9r�,�/N��ӧ� ᳑��D�>0aH:��.˩ �ۣ�N\���|p�Bo=�Q��A6~H���$���A�:3=au?�\�$Kw����{�%M���I��;���P�'�Tl���Mo���|��k��em����N*�f����W?����}�Ħ<��ݢ1�2m�=�YU��2�@�a��|�6Ю�7���j���"mh1���=M�KW�Ǧ�y��Ch��6�C����ʙP{:,n[s���9ҁ/h��I[ҳ�n^Y�����M��v�a��0���gm�^*1�a�� �Z깣y�1y�:ي�i�����O�	�ߠ��o�"�� "�V`6YV�h�#BO�����p�֌G�1Z\ �����l�N4�b$��#O�"Q.M$3�5/��ǣ������yF�	^�q�ٕxW|��D��`aŘ8n��@N\�͠˳�J���=]����91�He�f��E�|8=1��I�
���3�P�nX��u=��pRl��ԓ�E�{)1z���D��Q��C�����A���-~����9)h�x�筁g|z"`7��/����n�^�V����j��'B����ʩQy��5�0Ӆ*����U �)#���e�n�`ߴ&�0������N8E�r���@J���pI��Ih&�t�`�֠ow�0e:|bC�5c>ȱ�{�LB�|�j�?�
r��q�hH�́���QȎtǩ� �*��}X�8SD�h>�'r����ё��UR*iJf�QDɝ|������8��b���+,���̍r.�4@g�i�Ѐ�?�*6Q�N�v]����ł|��w Y�¾����q�>�[��=$gP�:���~�����)wY���e�C�5T%_Z�v��0�eߘ?Mta����j%~���B�f�y|����~��$z���&<<4r4iIe)�t98�n��,�� f���,������h
��O�ýv����Xm�"���q����Z���5t��5Z����j�s�>�Qds�?��&1���6��c��A�ŭHgJn���>8.=ހ���qZ�����*�����]�
2��J�-���e���}�_���+�P���H	<�����'!mPU�+��[t��
e5^�_�
����[C�T�Ij���Z��K����H�HB���ւ�������V%F���7�L~��Z_���3l��c�%2���o)�芨��~�hD�����$������eׅ�|T�<f�L�)��h���k��%����J]��Ar�U2 k7lZj ���7
���0�iY�����V���&��5�Pk���S�k]A�\�J���HO �5��\W�L�݅�)��@�?'�c׳, ݪCաiI�_IG���d��0�֤��jaJ�!���G<��+����uOI\�� ֏�!�"�SR#��e=!�+�9T_�leɵ/����YyA4�%���Ɉ+*};���p��Y^�������dܗ�A$��]�!?Yk���dl�bYE`�\�N�H����Ӯ�(v�������.3��}��:�ݿj��ʤ���lv��P0�%6��M!�$ƝC�rj��Av�
����W��V<ўk�n}��bM��ߗ�q���`!)k��"D�,|sx��&�����&p�O��5�"�(�:ɏ�:.��L|l ��[{Sq1R[��}�AܺOxX�~�c���M.z��k���	.A��� 5�%F����
ϻ�	��C�L���e7��N�gvKJ��+�#�9R�V9:�GF�ң�_���r� �a@��Y�C.��Jw��}<��נ_GäF�*t�׍,��L�Ml�$\%OO4�h�<�o]��6om�u�j�-2����Ɂ��ȷ��ɰ�cs�Ӆw=�FS��x���8�b�`^P/�#� �u�M�л���-d��{p��j�A���y�rϽ�4�9!���8��;��L��lZL'Gt �14�S �،y�����8��䨊�`�Ӻ���r5��������)a�1����]�w�}�ǈB������m��S�d���b5i�ֶ��z�8s
y�c��u�>�O^�����2�پ�4�b�ރ]���֠:�yN�z���/�4�s�#���N�Hԩ��֞Zr9���x��q©]�݊��,� �Ï�E���[K3"��gƵ��JV]�����Z��,��qS��p"C@�HV�;E��d�]y��_Myy�������zV��;I�a\	��L�?����kF�������d��C��ʹlcl�/r�[��%�A�i�T�ge��'b�h�	���K!@��U_�������*�6Wv�u����ݑ�h"A�:��ە�^/�q�M��d,Y,?����%�aO�TXdc݈A9����K;C��?)3Z�[9u��n=��S*�i���iU��6�,�&H~�@��}W�k� �W0wY;<�$�t.k�@���������M8�-�1��>?�< �ϺIѨr��\��Q}�\o�g�����$x�q��0��$H�]���zD��f]K}N%K�|è����xR���uX�22����H���a�BaW�VzYh��l {x����Qe�Tfq�I�^q{�s����"��hJu�%�wz�WdbZU/jޭSn���G�)ʨ��J,�dfjC����)���;��$wܚV,aA�fb3W�N]�6�9KV�<eg���κ\_�p�
ӥþo�����&B�Am|R��d�ʍ�2���e��pUR��[=�Nj
�E-�����~���*#��x�̃��?�������k�(��f��8�Ins�����7_R�<����$��1��������K.I�ȯ�ԯpי�D��-��Hw�/Nٽ´�s]`����?/����w�{�s���M<m�Ts4��3r��Ȯ�)�������4~>��_�7iE>ƅs���\������U%T����A)K#5(���D�g��3����ˎ��S<Y��J�/���Y"��&Σ��Bc�O?�L :1.�OPN���͇?�!#X
�)�ߝp�|-&���kB��CW7w���Uҟ�ֽI�]��qQ�K�h`ڄ8R{�,_�+�i�F^���[5���}2$fz�75�60�o�������⢫��baDj�⏢d�����(��ۺ���ƲϢTc ��Q��'��$�+5�"��T�,�����b~��)0�9eF_p$��UCkX�V��=��b@��
���8֝O8zwE�r]^�'�@)�ԅK��b.>�©�J��Y���v\)`�M���V�>�LPÛB���C��ݹ�Jlĳ�&�6��8��o7	���S�
�3�J-R�nu���e(6��@�muU Y*���]�A�DH�� �,����$1@Y��/�ᮐ�1�8��"���F��ݬv�<\�|T����ht
��c��hIP���8:]�9�2�S���p��Q���"���u���I̾�p�Æu \q�;6�s�	�{��w�h���̄�����U Z��8P��9H�7�3�٘���K�UQP��/�4%S���j�j��S�Fg�(��`�s��%o�l���~�h����Kض�q�[	0����c$�>Ce
�!��x	�YI�1Lo�70'�'2sH"��t5fm�)R�	�}SW�0���u�_��R��@��3б�#Uk׼VN֢��6��4�	F�����?֯)ZW�n��O5�ƽ,�/71������1�Kw�����dj��C�ڣw��JZ�'>@�'����
2��ŉs��v�gvp ��b�����!�V��
�g��6��;d4W��2{Ī�&��K	MBTsvϊ��ꯖ2�S	��.�4 �nf�]W&	���ű�"�NT�_DM�[���5��_|i?�Y��Z�=~/�#XQG�����)���f侕������g�Z7�P��i�~�� �/�"�v~�)�,7���Z��[v�ك>JGȈH��M��qx�l�)2����Q�hڢi
(W��Fj�af��̲Ӄ�.��*I>k� [�m�� �5aM��R���"߹�92�9;yN�c}������拰cRҫ�xV#M�b,��z�{�5:�O0�6'%=t dB�Y�]�),��ھ$LN=|)���x%���-#b��e&��j���a1P=v��hۋZaA.�(������>���O�vD ������x��-N��&a�^�L��MK�l�A���>(�7����yEfo�<:�{p3��ïj��S������q _�Vظ���W�~�vz0�<ԏ��� /-(��Մa�/bՃ�{^��	
��5�c��QΧ����A��Oe��}���:�dvs� �������P����վߝ7�ƕ"׆ت+<�FMcp7u�Gq�lt�yb]�ǡ�_��-����9M�}~s�����mq�8��]�̯�b�x82K\^��*w�ھ������Ex?�Mh����uId�X9M,��R��sh�Bf%�� �!/-Y0v%��C���^��R�|y����	�:�l4z�>&�"�yi��9�2d[�?'dқ����\/�����&�X����U�͔G�����Cw��O�/��g��,J�)��.Nn~���5��Q����[�Z���g$�I�|��I1� =�R��D�ա��[�U�p�Q�[�.fYb�iR�F&��S��|���V{47����^��v��"p�0?�7�S$�]�ϊS���bj�v������Fr�s���:�G��u$�}˧�G��rO���;�.�8�lC�k���З�c��KH�l�rӳ}9t��9�E�ވF�p�l���6�ljR��
�IL���r�v�4ľ����3�� �^S��` �i�D&��1��V }���F.�?l	A���K/�x���Ђyn!���@wt����s)�X�HQ�q^���縿�r9\9���M�"~��tY�R��wH&�&()#E��ܾMH�t��,�2��lwR}�2����W�˱���t��(F鏧!k>l�q�\�DZ��v��nq�G�6e��Z���3�y`���lR�*ui��6���~Gѳ?�Zrm���L�]U++1��l��gl�����J��:�l�Q����@�S�Wm3U��a���|���X�<?"�B���/<cA�/b���I�qt�ǁio�Ax8_�3��k�:��X�����Im�j�n\/�M�3��$88��m=%��+��B��v���xm.�X�T��S���4o�����ox��
�ߴ��� �����}vP�R"�Xn���-���S1��̶U�qρ�9ي	��Z�ڿ����Z�mA�����Ǣ9��[&��@�X���{(N�L��r4�w�wu_�4hPג��70%*:�,0�P�[s"�tNyo�]8�u���\ϒb�Mw����эJ�����K|��
k`sMj��k��C�ͪA>��p��N��h0Q�(�b9�Jc;r#!��"��w|TH>D{'2B��uH���j��q�"p|��_V7\�jA���Ep���u;b�d��Y�te�s�I�C� �'���3/d��7��tK\+����tԡ����[K*�3���zt��[4荽F��UM��ݺ��M��Xیא��slQ8t�PƢ����6�&sJݓ���%�Dя1��~i�S�&�kx���Q�q��f0�ߥ<�Vܘ�m��u�Ք+�e2��N�,�03k��"KU��p캠p�N���Kxؒ�\WO�Q��s�Ez����,3SM�Lxj��N!%itdp�%�Vd䃣��0"=�'ݥW~,.6�7�- H4��e���0Ǒ�7��nb�/>�S6+���G,şŻ���)OPᗦY�{���1��	�c_G������E0j��H��/���U��]�dȃi�wW��Z�3��1\'�)�G�pBW>���E2a~�9�i�� ��T�|)"-��΍����st �3O���9Qn��	�I#4�flF��\>|����؞Fa��tֳ��o��ɮTX��5�Y�C�[pԝ����K1[]N'f^ڑטC�\�b�<cy��^�eOL�B�Iql�g��Y)}&v6��� yn�|�D&e=��ب9Gҫ;�VS|Ro���
q2��ϒ�EN�p���9t�v�Ѿ%�ћ�j^�&j+)#�K���-�û᫔�Y���P�ȣ����$dp�ipJ��=g���h���C���`��L]Y������e�N��e1�x�1
K��r�]h5�UB��T��X����C�	�Y�E�)�N�LJ&����D8��l���P=@Y*y�?��R���;}�O�ǯ��X�j�O��X�P�0����2�4��wQ�x!�_��T��g�J�R?̨Ce���4c|	���*+Kꅷd?h�=]�\t�SG%��^�U��\�[��}�~��˝�/�}�qԮ�q�C+jj繕T�,����:s������ '��] N��B?��Q
�Ӗ8so���������m��vaS�7]��I�M��� ^fZ.h�p1�f��PҰ�ٲ�>7)ޤ���]<�V:KPl#wR����DpD?0h�x�$�¼��̻�h&�72
��9E^Ѡ��<�V��[�z(���|����� x\����f��!d�hX|uwGDt<j���KK�?�f��r�fe�L�ٽ�6�A�\>���|��Uh��:�M*�lc�x BG|�JQ�cɔ�JЦr��!7�z�?^��Bo��6!�y�p����hz�xV�œL8Qb��Ԯ��.������`j�2L֭ڄ$��-�fm��"���t��D_^��xŎ0W0�آӽW�C��q}����h7z�u�����I?p�e�f��KQ�?�<�w�ۗD���}�L����O�,`�b޴"b���ǓcT�)�2���Nm^��;P��2rpLņ��Hu��}�|q6���T�S󲵬����TFq�Bf1��F�t�2���|uI������������Y��)ʩ7q�P����䀪u`ќp�� H�w�;�H�P��O�q#|<�9Gy�"$�Plq���Cp�-�΃�9(܁b#�H���d�lc��?�L��og·�8���(�A�F6;��	���+�fSk�?��5��t�=��n"�ˏ�
�Ó���q���Fl��h;Q���9�F�x��Ϥ��ZᏐ*����,}x�r ��-��'�)<����c#	>����i��3�E��XEը�@����d+��IR�.����$(+a��MX��[;�I2�n{(���J��;�ކ���=êѓ}=ٓE�����@+z��0 I MM�C��!�C��T �nJ���B��GT���"9��EΟ�аҠ����<�n���fЪ���ȷ�� �u�A�UJ����R�Go��䒕�VǊ�Ԧw���f���l���M��5˨څ �z*%��, ��;>��ە��y�#�	�>��q��1Ę�s�뫋W&H��LkS�07�p­�0��ґ65���-��&�1#�5�	��������a���[N��l�U� mjə����Rghv���X$|pïj�C�C,�_��o��̍
=������{&v�֙�F��	�T�tI���L�J����_��A���w\B��P�ЎO��U��� ���Du"����}cٙ@U���Y��Z+ᩊ����ù�a&���}�I-]y/���8�H�-��6su��6�b�ߵ_��d�6ڽZ^��a�<ϟ�@� �f�GPoO:�n ��\��͹��6�~�p��ִ��-?�s��h��ko��A�Par�_'e���{��K3��>S5��CgS�[���R�!����H0�#ٜ��ė+z0ʥ	���ɹ���tH�Opw���pX(���i���g��o��H��A�����v�L��$`��ƴo�f����F�W�d��EV��; ��k8���y!�f"Yf3Sn�Ox�%)�>�o����Ϙm����R��yH�o�g�����>Yq��aG<��4c��ኼ`[�4�w�R�-��gw�����~q�%RF���i������=EB�b�L�'�,�(�F]�a,X)��՚y��H���,�ܼ�Q��z1P��vl<��n�o��a{��E[n�"V�y�m��y��fV��/�چ�G=�K�R���YV�ZWs b����ph��N讠A\P�?0�� ���O	Em������&r�Х:�AAs�~�ؒ�ߞ��J�pfiֹ�=.�+���uaF9~� ��M�r��+�{��B�2��^�Z��<*�C+���s�^e;���+M�2����3�v*A�h�{R^��*Zĝ�0�ƥD��4�M5��AP#�|6C1j���V��{�X)x�`�Z�%�&E��o+:��
ո��?<O�<)6�� l�5L�� ,,�[�_��h��"v|cG�ǝ�j{I�'ʩ��}Q�˃�y�-�K�~˃�XkǸ%a�{,�G4�#��<5�'&����f���d�#'F��Ɠ3S�$],˿�8�-�z���j��-�|�!�{�mv��S)�o�=ؤa�<,^�s&�9���Z�Ҙ����SZ˙4����q/aܐ���1�[�H� �;�cprm�D	�1���'���r : $qh8{�+wN��Ƕ�,g�.��k*������Z��zyC�;���{_!�J4D}e�DP����dC���A��}�
�kK�D�%%K�$E\��vw�Ӌ�-�HC�7��y�8+T��y
�M.�Xf@ࡺ�N���M��=0l���g��<A����l��ŗ��\)�ݙ4�f����N}75��3�&��)���kia��Oǡ�?�f����[;�J:�i����s� /��ژ:\1ē���9ݩ���lK��T���RiN�_�-����Lk�\u�O���.�3>dRR�m=<�hf)2_ށ�vt��q�L�{?%�% ��d|6
��Տ
*����j�ۭ��4�Ώ��:��:�׿#��wURH49��7��	OW<M�Jb ܫ��QG�0,�W��&H��#�ʬ�@�Br�Ġ���P(��W�--��NP���:����G��n�}����#u�vc��(]am�&���ߪjef"%��(�Ǣw���/�h�Sa}0Tb�F6t��K
(��F*�������Rz��̘�I�o�̂�	+�<L"�Rג���sm�xIz�nyrw'�6��\^׶-�tb�{o��\��K�+��f�fJ�Q��yi����S��j����xN֊�ǽ��r�0gSf�<I��M~5%_����Ä��/����KF�k�S��AS�b� �Ղ�����I� �=�d�;F��A��L�H�~ НS-~I@ڻiM�����\I��?�	���E�2[s"i���:1�^O����~��`�}$�99����ԟ1��k��0��¹�(�J/;7�q^*�@�ӊ�������(��O����2�I���-{١t����#\q�z8{v&X�_v�ᩁqt��_B��'6��'��Ԙٱ����6Y�6��>�5 �Ō{�<�wy�^��y���|h������nT�kӗ��9řM ľ�	��ot4�o�cR{\1�q��
	o0S�Ш!4�L�<��{���q��Kl遠OR�Zp\��+�UzdSq���9�^�'-$��'�3.�� 6�)`dએ`�EfӚRP��.K?a(�J�M�*�ϑ�a��;r	� ��=n�Z!>q֥�ӵ��f$��6��FB�x�`�C�]�B*QȦ>�z�)��s�1�M����2&�Mխ�t��o�v����Hbޥ$��p��A$y�~�[��Z��,%�@��!��2�<� Z���9�	���U�����($���\ea�Y{i1�v�w�'�i@B���8�ˣ��f����E*|4|w��߾~>^�jkҋ��b�������U$ԍ�qu{��6����$ӽ�H4	�U^� �*�K����s-�X]�R!�f�Q�]
����%���h�l�2�l�U/����!�%;B�f�ܸ&C���; (C���.�
W���;����g�**�^�0���g�N (NJ��u���ƍ�h-��N�X�T���?g�r9�ҹ�]=���c�������F�C?ii��0>�����E)�,K.�rJ�hHi[��{�r��K=h�[�נ(i�����b>�S�hx�Ŕl��syX�,��Ώ<�)�+�D�J�z�S��2�
p&��!8�8ۘIM�5e����E��Ы]k $����`nІnv�1z�I�K.�^�l�J/�g�{Z
���Y�k�/-'!�#��e��)_ ���a-F�8%�t��|݃Ek`�3W-ԕ�ކ0�-$/�lL	D����t&��*�:*� ��Wƻ����3��w'�b�{KJu�_��~��PfR$ҥ�7��I�-eȐ@8�^x2���ݤ�}�u���>�g�͉�qB�A�CE���$�"����ذ��ꍲ���09[������;�E�,�,83q2p;;#Q)B�f�·٭L}�U.���4
D¯�2C��h��<�p�!HjҶ�c�rv^0(���"L�0X��/�7�dkE*�����bM��-�:ׇj�4����MC�"���ǭ�P�=۔S3m�ң�όn�H BY*ez"��1�~LSӾا���P��\7_���G�v�e�k�9��J�^$X�t*A:'v��35^2 y�[�-�����ӒU^v$W�#���wm7��������[��p��L�x�p	��$!�=�'�� ����Qf�� ��C��#-+�D�Ķd���P>���/�K* 0��D�� a[ҡ97/-�W>�X�<�R�(��-t!\Ѓ�2"C��xW�~kf<���r��p0������/F��j{:)%5X1��u�e�xy���#7�|s���9�9�~|l�㈬�D�ܓf�T�3*s�¾��jB1e��䓯��"��
�r��çAf'$�DHL���FW��k� C�3!�c܊�m���Y+��ݘ�י�}���.'�3��տ!gEm�.���k6���Q$����ٹ�s���?K�	�3$\l-�����.�X[�=����3p�YdϮ�����:�&�ڗ����_� Tv�`��*�0�m���?Nb��I�$�#�]B�b���}b
w�<kò�i�BvӬD+Ԑ%#�9�� F�H�GG��6�� �׆�c�����xU��
���#F͏�f����.DĈd'6�t,Ec��'� ��w������l2i�I�X9ų��g���A����&y]�Q��g�4��9o0:!�n��%�=+ق�3ӽ�P�M�Pn���4���䨪�֒���+q��b��sT&#�O3�ӗ�e���7ǧ	cfL|���0�-Cʐ�{�!G�q[���,�'~F#/@��x�@��c2,�3��bW�gPqO]�������#�G㨄51[t�и�b��BW�Z�N�%,�Y�ծ�$�i��lw��azЖ���_7 ����X�Sý��ғ6E��e�_+ u��ru6����\�#����;��G��Vo����ᅷ�cyE3��FN����-X�4�Y��bv��.�gx��]˒0zL�^�D��iX�K���	Xk/30��?�K�Q1���ue!X������F0��y�
e	�fU�lݖ�%�+��d��Rw�$5��I�����Bx��2Ͽq'��򫟴�'��7�B8o�Ӈ<Q��,7���$�����wvة���k',':�D:��[及a��̈�7ފ#��*�9����ī�%v �p�uݒC�K�����4L�۬�'�F��c���AJ������7T8�C��{@hē�.�o���D �
g��߼�p�
�@|�^�h��(�zA�o֍#��[I�;,���k��#�d��W�!�,i��c�����H>b��Z���x�}�C�S;vD��Dm�ހ��S�7�/�@���fU:��*4#��	N�#�H/���b'�Tp�0S�:�QT���B������ߒ*~�^X��XP�b�c?�W	n:�����4��k�"YǼ�@ٴ��J��F�S�:�'��9|���71Xn�6��&╙�Wa�8>U�ݓC���R %g��vLY��%ߘ�(n�ɣ`=<O�vC��JY�e|.ܰ�k�so%y�����K{���4��p�����s��s��x�9^��j��tB�-��?/���<R(����@�����!WhjM��4nm��Y����cTx?�*v	�;R���pj�\,yU�3&u�yl�bЩ��,;f���E�	<�JF�Z�x5o(H@�._���l��=^�}���Ӭ���-�â�b��.�J���9�!s��ш�u4�LM��*4����9�%&'-�&���֙�
7e�����s���rK�URN��Fu�P�Q�z����F��iSV�+v����a� O��-��"z��a�)�E%�����a�{���x���A�tp�Mӡ{��Ս#��O�r{���O��2�rѭ�1�9���voӇ�]NY����ipƨ�j\��7����0���:"��fū��0ڡ�'(��8�&H�U,3{���e�b�����ҧ�V��Tb�a(������n�R��C|@�u�}|��8�� �ڮ�t%M74ּ�����aV��l=U%�_��߂�`k�m��w@9�^��������z�5�~�4e|E���.���k5s����$^�1�1�#��w�ё��~�5��[1��A+E�9�+ͮ���A	���+l�n�V*M�D筷��M��t��j�K�q�e�]?��xLl���-������^�١-��sc)���I�ZK�d|��[�t���9�z�h������� �ׯ^�&HTg��X��\�:T(�n{���[��=w��V��!z�p@�����ݹW5%�Ƴ톆�Ae����ֻ�'@I�m�ʢ�L�7�'zLZ����\*:20x[ؠSx��]�~��gϦ�	�k�,NT�\��n�{{:�*�)ѭ!�[r��:��o�v��L<#yU��랖���A3�*B.��">	1�kjȘR����
������B,s�m�h2ɷ+Kz�z�7_��a$����O�c6�7z�fJ���Cؾ׋����:fd�d�~�@���tA�1��~k6	��\�՝��F����k�t������I����P�W��"ܘ�Me"~2Qn�l'u�S���%�캹�����ނv0�r�������2�)/WH�s*T=/������t���?��o��0G���zx�͒$ >4�|H`#P�H�3�o��_Kv��и+j'��)�̈�� �f����=� ��ށ?�<�"Ր�O�<�"5�h%0��w�@�E4�4 �	қ�⒉��=P�<�ǅ��A��@��>����	�wFuzu��R�*��q�n�J]��~y�yٳ<������֥/��(��F�q�o�H^�P��g�2���ǅ���2�� �r| �� +Ϩ�]�׍w��x|ф@/��'��┤ݨ�s8���e2ۚ����"5�9��!8Tg�N��<�k�H�W�{V��O��_0ɧ�`���X��?�QPħ'�� �k�5���y�S���!z�k�a�<�v:Z��}
�,����nA���ӸC�������{^SE/�	���u�곏�Ka.G��-�/�xt�F�x�5�c��rs9�MC���We�2�s����,Q�;�^I�F�/5�[�����[�g<���
�����1D�3�B���ȐV݌l�ҍz8X�ax��bO�v�2d>&"b��lE��zN�	��������֟���LN���)B!��g�̖A.�(̺<~�H@�Q&����c�qY�;�k����*&����ۀΎ!�J�O�������hvm��Զr�/��=�@gV8'߱2��^��We'j��W�KB�	Dz
�U��ߡj�pE��o�`;>6mݐ
�V�ٻ�Q:I����T�)����ŒA��r��<�����L��G�H�u?cŪ�¯�sQ��OA-���h��G*�Hd /?W��.)c��n��r��#�nK��]�3��SJo!r����'&1����kQA�n���fX;t0H�g#]�}�C&��(l:5:u�� aC;ږ*�"�k;2���p�^h��
(]$V������9o�`�e�Ϳ*�`�V�TAn�8���OV���Q��6e���S&mo}�|�h�h*^B��rj�m�3]���w�ԛ3�ގ�J�%��=kՆfȝ��5 �FC~s�q7r�_�?���6�|���n�J�u�����4	��O�9�<}�:�J�14l'�W��sfP�sɸv���~��Nƍ����,� ���{�Y�0�1���5�1�9��ک�%x�~��m���2�۟��x{�c���)j�ǰ�J̌��ʒ��dü��K�Y��0k�[n��l�B�o�Lt|k֝3G2�	9�w��z' ���1����$��cΫ��ʋb�Eo�'�Ey'���Q娿�ebUE���1�?�ʙ�̵��A���@�9�#� ��}><��-��X�!�R�I��45�&f[�'T��-����l*�X�f_g���z�����S
}seÔ�n�ڸ�cc
��OL^��E���Çu�9��m�V��8�>y5��΂��HYT�}�"��OO�j�N�*�&=��q����|Jw"@fJ�e���4$2$��ri�!��n��"#�?�Y�beU�D�:�)o��n_�`�/���ak�ӑ->���o�=�	Xg�l�`�����BPRѯ�Ӂ� ��Bހ�׫b�I�=��5��&�g���Ca��k��.Igd�yrpo�$AQ.�M��̿W����YW�h"���x\q��7�/����N�H? �j��wfVhd�s�N-���a���4���\�Rc�l��	��ZH_>%����w�$�6# �@��⪅�����ȫ
*��̽�f�.E�L4R�N �$ooj���$Fa5|�xƢ����h�	�}E�\Q�xʕ���K�>7�,�O�����������lӓ&�Z��u'����K�\���ƽ��� �P���~�0.O�`�bT�v��|�zV�%"d�x�FL����-d���$�O�xx��O�.��LSĿ��$������wJB�P����
I~h�	���-�M�����Oa�
;�2\��m�)��A�,�~)ޓ{��vم_�5v�m�ڲ�X��aٓU7!��X�']���d�t�Ě�tMԖ��^=v�R��M{�u9h�kk��2��V��*�
�A!n�E��b��HB�R�9���G�b�u��&����ˡ3�v�Y���`�aƸ6���3�K��d�\��,�*�.�����25�AS�9��D;���O�T�`���rx�&���<�4�v�{�>ߙM�o�ȣ�)=�}�]*4X�%�\pw�d��ے�mTI��FgQ�Ŗ�k��p"�h^[�G"]Tu~�v�N>���IK�����m�X�SL�Gd�,� �Z���^:����M�q�YPy�?35L\�"�|���yuy����A}
ꦼ&n�$�>����Ɗ���5�#�(y��:�35�L�ޗ4]FD�!�c3�?�����vB�$��R�+���b���E�!�F��eM�'N�I��20�@sE�h�v:"ŗ��$���ٌ]�eXp��[���j��S�!^sK�K��8���F�m<���)ȝҤ���)���@ٜ͗�#����A[�K:Uy�~d"v�ڞ�D�YXhW_F��jHJ9ά�ĵտ\�`�$���Dų/C�0����\I3��G�2U��QX�xPU��C��z��%��+Or/�z~�v<�uޏs���VdI^�3��H�T���J��%΁U3DX�m���[`��Z�>#nî�� ���	:=5�*8�5RvmCm�JCӘf��.�����r��9ii�9y*L]�b�$:�J͑6�6��~p��($b�R��8�O�,�3x�s��g�sTF�F$�/ϒ{��7��y%��Դ�L��2��.���kg5�yQA�G^�j�*�$c��*�}X:�	�(��	<@F�EVMiia��	a��Ϧ1kH ��F�u/�[̮O���"�^{kM��"$��ܳ�&�{�)��T�q�S�&�����>����� A�<�P�:���_�>� ��3U~uY�>��gb'���"�_vWA���,�*-�^��U��@�P�n]䙋�����L�w��u���r��g׆�a�Y*�%���W?��KIuS�A�m���~E��L�5Tc��EΌ/T@��L�b�����a�|i�#i�l�/!�,��q�( ��I�U�*�k�3!R��K�z����?a�	�t����x��N#��q�h<��c �C�j|�1�k�]�Yq`�����\�>��ۅ�C�`k��j�Ñ��o�m8)ą��[Kq��'��$�f�<��l�����(��.C}_�T�\j�l���.A��̥��G�4X�Fw���C����2<���zN�踺.�E��#��:d�T��?ʼ��{6���oo�]�ӓ�_\ϟ��m����$xy׼�{R�����AxgZ��;\��z�g�*75L�J�o$4A?x�U��_Z�fB(�H�^��)���	*$��Rт=���xG��:�J�:�LO7�p`������J�5ð^��?E?\��huk���M�л��oQ��wo�wo��m\�Q-'�[^�-�^|�	���MW�key��AU>�����ѹ; ×�أF�	|?㈕�b�_���}r���P2&�w�ԓ=ڤ�SBMDO	o�K$�.���ϩ���~���p����{�* c1���z��K�qW&�&}S.�:j��T�f�KٮB���A5�PV!�68	#W��G,�h����A-��i��%��E�O�j�[��Y]���9��q���B�mify��=��6�?�#A�  aD�f; �V����mnn�t{p�!��c��|n;�Z��n�`0+_=�9��|����%�
:�ÒY��~���ÉM�,e���� 6��) ��zO!z�,}�q�7���HE�zV�~J�} ��)ʹ��N͎��t�U�p��y��I������@;8D�mr�P��z�-��d�K��+U'$]F�]� ���	��9�B���<t�U���C��  ���?�ˤ��1�$��q�G~��-KA:�-�cg�Ӷ���/vN�B�y�P�)���n)j����\���W����{�P�L6����&��l�mA��煼,�I�<��O"��`���{5S�WnC��RXsh<P�<ޓ=m{�ymb����g+�Ov��x��c�pM�2{ڶd`q��::	��am���z}2�:W..ݞc�.���w��<cB|�5�#��2;e&*�-n�i/�'�A*�.���h9���^����^4�q��o�7D�ʾ�jO:��&�"�<0�^�3�b�v��(ӠqЪ�S�U�i%p�<RY��\IК`v� �~՗�e�l,�zl��k���{t�q�=�C��p�;d�۸���x׹$�}�DbQ
7�.x���A�%He���|(�d���F{�܉1of��A���V<��9/����O~����*SA�l� r��'��}�� -8���-�5��>�n#T���
W	\J��ۺ�u��f���8ПK�ɤq�[,A���Q ���C�����:8���f4�`�>_\CPݞ��n�-��Z�U {�n�ʛ��>+�f�a��4����_���6�=��>ዊ9~ -�'����#㒸}`�9�
�j�H���m7� �Qs���)��� .(��69Hr�ܷ���Z���� $"����(�~&��1�yb� q��q5�Zr�`,���`��S��L:$v���+�}E��г���f84$��ˌ\�>�`�)�f����@�a�+�⧪����ō�_E0&�
��J���cF
�z!�%�Ʊ<-㢸��\-�������Q:�E����
�S�wE6'��rQ�ѐ���*W��"�4{���5h��A��o��o7�#����f
��*q�?�����]��2�|*@��n;�)z.5H�)���i�����YF��;H,,X�*����C6��ӨS���j�\��q/ �w%���d>����ߟm�v"�5\1�<�Ñ/Cl>��R�Lk* ����=��]�Y�U�~,���yCb�)m��HO�A���W츩eݣ�m����}�V�h@�G����k�)Xb�ש�m�ujũ4I�����`�k1����bJ���`⬍bړ9�mN��:�v
y��^�)䈞#�q����bvf������;��;��v���s���R@E_L�A$��q@�K�������|0��I���o�bAy̢/���;5����fG-k���U�p�� �ճa��EF�R?�q=�m|A�j�a�/�>z�sL���+�B�,��vNi��t�Y����>O�?�|��UXI��d�5�h��Qx@�2pI �_��ӟ��zYяU�
�W>~��ݳI��2چ����r�����0>U������ԊX�EH�%�A?iɉ��}�@D�םgx�>� ��}2��"��_��`���y�Xf'IRN����Bc�*�0
�/���������[9��W��kTS _�+ˑ3�\�|�*X��ط��'�p�`��(�L���;�/Ѷ1���>/鱟�)�_�규ɣ���7�ܑ�iJ���eG݌y�_/49kE���E��FK���ݚ�m`4w)ā��V��d�T�����ͦhP�Xh�2�X�� ����0��-�ࣨ�f�w�f�d������
�7��1��ED��@9�sAr7t�V�S`�� �SCՖe����c���(�e���g�=�Z%�Jp�Fp��ľ������)�c���Vݴ�t05D&?������d����!�S8���&D{&UFӇ¤Ms�q��j�ols$�Z����W8�><[_T����r+B~?�!4$b��O-@K*��5�l$�"���'nn4����l���H�k�i�U��rGB�.��s��c�	����.�ۥ����UΕ���bL�1�3���oD��Ӏ�̮oK͎�}j����˿��|.İG�jز�qƛgY�k���m>�PĊ޺#~� ��)� ߰��#"�_��ٺ��W�Uuh&��Lp(ԣ��\ǒ+x�3��-�5+h
kN�e�^�I_���K�	���¯G'�O����U9;�J	*K�ӎ�	�����Ǡ��{:��˸	H�7�`l����; �{�F��8�>6�@����~���'	`L�J1�x��ޭ l�c�LB Yym1BQ5F���Ha4P��#B�ƀ���R	�T3l�ym��~ �6xuN�c��c6_��b6	�[�k��_��K\;���o��]��0L�Z�Ɵ6��s�2lw۷j����o'��4OY����{@�C��<�u����j����%ڦd i�q���o��Zi�x܆sԬ 7���u	�������b+V�S��2fZ�E��m������2C�f��2�a`ҫH�g��1�����~���-��9e�J���f;#��S���~)�[o�S��w{���\A��j��d�U+������"+�,F�o���G�C�*��M�?�%w;������&<h��X+k�E�n��<�1Q�A��c"�r���3��vM-�kE������Z�-���l��f�e��u!p�e�v�/�
S��}y���63�7S�w9:9����d��:m�<HUt23̺��N%����&��ZE<����ָ��:ש���F�#�*~�5U�7�:�8b�熵QgtyGJ@:D�d�[�QDU��z3�k���?Q��-��Rښ�6|���s�A��N�\"�=���2��������c�)pc[����m�א�k�.��� ��B:%�N�$k�(��P�ct�|�U8�%�6����O��m^���@����{��nM=��q�n�Z�araQW@��h#���xo��������d�����:��Fg{�^�x쉫�=Q�[<gт�{�#�rс�6�U�2�qr�n�"�|�l�ڬ��[.����H�0^[l�K<�}O8����"B��6��.!�I9����U;���K#�#DZQ"9�H�Qb3[���ۡ�[�L�u����"&��W�n�O�M#e���UÕ���j��`]!Sć�릗�6(�<��l���x,�3K�`c�^_o�_0~G�����-���T��.g|��ף�d|�sL�c��%��o�������[D( _?�!#��h�&�6�3��!8���%хZ���x[�ڔ��-�%�Zrq��
� zRXrû������Z(�+<惭�R�z�G@a9Ǩ��b�V�4����IVQ�}ۜa�8^�:�Kj@�e��<ɩ�~�����d$n���":pD��t�Q��px�@$H�<le;�x��.��!*<(�p�L��!Y�FJn�Rʥ�Y��Fm��~Q�J!MG{*\�g0l�"��w8��ZK�L�l�%4ۍ둮�kI�s+�5�C�h3f�&��Q2�ӊ��w�V�ꘅ���ȍ�����4<'h\ӏ����D�2P>_[��wG����b��{쾽�%=@��>�G�#�R�CJ/L������Ը��|30^�3aMU$d8���I}�O��6B� l|WPDb}��S0��-���p����L�?GrB��b]#7��IDN=�q�"��)Q`�Mt�3�t��-�v&])	�lM��yk+�������N#�Oo��LN6�	9�o��W�|- ���֙HK�B��#VN�^��]v��ZoԄرg��P$�������1޹�� p�����(��A�K���*z�,�ko&��.�OY��i����`����i1`��jlhsR$��J�:�M{���3��w�	Y���M�R�p�%�H�[��������s�ok?Q��j����3��	��p�dsдC3��h8\��`e|�$��D�w��/4�F�r���m|���'H[��5?��\���JU���W6���n��`�k!��>Ʃ!?�Ti�rӐJ��&c��bC�6E�{Ǝ��M�;7�0g�~��v��æ;�b��/~�x1�����$3������ڞ]җ	��[��3)ȿYG�\mWG�M��4����)����]��9w�3�߬�5�mގ��(��"[�hHY��]r]d��lH����r���	�wEL,�l���yU?�k�Eq찱LB
����$�]h8+.�����]Q�-Z2XlՃ���i<*���f��hkN����q*qsx���n�cn�ے����W�������_�HF�
ふI��W�+6q�:dX�L$����D��tkʒ$JT.e���1��BO��V&��� �D�5��U���9��^n-P�b�u�K��`�/n�l�,U�+ER���Q��_��Ó�r�w�*\������yn�)�8d"̇së"�m�ӯ ����j�P�U��ݜ�����M�/:O�#����b�AZc���L�{o !85��H!��ua��	�Fw6Oҭ��e\���^Ż�H��(��K@�G{`���<LM���?�U��7��!�j�3w*�B��}ժ�u��m��`��7�םm��t�86���N���<� C1�?;
ֳAEa>�F'3�T;F�� 9D��� �%�TqɆ��\krW$/�I\�����3�N� ��t}tST��\}���e�a�� �n�h:$��U�<���G.�D��E�)�		zP�Y�һ�Y��r�l�h��Z�<U������F�|���U��f�E�%�~[��o�|�Z<��
��ᮉfh{>l�S��HV����y(���#眹�# ���-�IX��Q�v{��<�z�܆�EzP��������@�-�Q��b	��IA��~���j�����s����v�t.t�����G��"V*v'�5�����)d��l�B�	��|���.�RT�s�ٹ��_���	|B<��Ĺ��٤��>�ZM ,���$��f0�@/Љ�<R
gh��>��m�u�{�&��z�R4	��>U��Głc��#�*��.��x�e3�T�>�/����%�z��}%FmOv���S7�Ĥ�o���2��A#楡���8/�L_�<�đ��dj�^��mR�F����\2��D��� �|RTeG�G�f���v�;9��X����P,><�9�
��^gFW$���͑��������+��n���s�뉌���aߟ+�f �q,��E;�"��o��=�T�U
I#b���5Ư��Ȁ�v��/dn�/����iR���	T�7�7�U�Krm����xѥ�l��lZE�y�_����0[~���ק��L�����ȳ�w����;�|+�N�7@��痼�b:�ծ9(�*�ם3��a�.7&�d}~��Pr0�OcZ���!��H@��R /��]���yFJN�E��DM�<{M%���i/N���]b��R ��٣=�P/�Xu�.�#T������ז�M�'!�n�&�&8���6N: TGx �o	��x�'P����2I�Ft�=���^a�j/�DA�"��)��U�!�q�+��o ��_䡨A���mԅ�ؕ��S���7�"h)��3E�K�kQ�D+�A��
O���7�e�A|�K*
"�*�#��K�.Q#^S)G�����Gbq݆\ثA�Q�-�Q�Ĩ�q�(x޸�d����$��#���:�x�������J�8���j��P�+�_.�����& n���es��A����FkԴ���B[���%����,�t�̎�����8�+�ɱW��Rp�Q/��L�Rp�~G�).�2����7{F_m,@"������r���*��2����z��%Um�<l��E�I�+Ib�֚���SM' 3f����{ì� H��M��,��}������ȧ�;1��`������uZ�J��K�v��j=u�#�m�Q4J�"����)9ˏ`t̘`��L�)�BD+ϣ�>��]��`�>u��A�/^�f(%���'}�þ��
��K��ͣ%��ښ ̚P�c�_y��� P�� �0��vL�L���s��ԠbM4{�����-�PwDAwSU0	�]`�n]� T-�F*�}�J{�� �ҋ��T�ndX�%.2 �$�Ş�^RGo����
;l�����cЧ�#f]Q'��A�|�w���?�"�˵�7".��kC;J�u����bIH������������#:��MB@��j�e��	v�Z��>8�wC�h9���澒
@�� ����P.im ���~E���K�C����v�+��kHs�0�UTW�jr���5zٸg0v��&�r��_V4��&���zBj|6��y��h~6�N��R2 -�lss��l�#�u�	�4�� �F�@�"U(Y\o��4#��7>�`�/��j��?l�׳�N����b@��nłӏ��b��_l2VJD�B����B���R�� �*��PEz�3h]="���y�(�����NL����h��{�|·eӢg?�ZS��O�u=�*��K����H��VC�d��;�?M�(�S�>`��Ǎ�0P�\��="[j��j�(���ɨ�%R�k�X����	�ɚ�ȼ�V,���/vB�K�	�����S��k��d�F������g^CY|���H�j-|en�Q����0#m�hph�KPU�y(���;X�څl��}N/I/j�#�>��k賘:�:���$g�<J]%=�D����&` ���s��w$�3�)ڢ��5)�~�>$�՚�~�I<�����������'T�=��5���뺴�7
�!��QD�㦪�Aj���{}3X�\�xjEK+"r���v|Ĳ�ݲ�������{#`S��A��̖w*3�]%n9F������#�T�ab�odPd�X��|n:$�i+Y�a�����$��y��2*$�|(�;��j�W���;��I���F�E&�q�'�c���OR��PkV��QD�x��BUm㵫΍�����Z��:7����@/�dt�f�(�}��1 ��m�]����o��w>&d���}�0���Mq������tz}}�����'nL��$����ƾ�RSC�ūY�Oߌ��jB+eg�F��/fr���%]=5
8�X�f��Hc��0���e���{f��,)1D������{��^�7���]o%7q��=�;����7(Aa�=��DGbI|�IqS�K����CJ`C%�󲈏3�0���W��Њi[re����&�p���IY�hec����8[�!���8">-U~T�=2ڝ�5.����������(dŘ����X�H��&��b��n�����7�gՙ.S	�M�D.M�B��t΃�=��o�Nת�"_�'���R�Y_ea��ؿ~t�]�7;���;T��Mn΍��l�E�f�/?�3��|��
hHc�&G���;���"~����.B���5���&n������5�-n���C=	�h8��2��մ{�f`��Tmi90uR�Ҳ(!?��s"�e<+ъ�,�cZ���%ńr�3��FF��W\ڊ�ê:F��\��jy��8Ph���(��o�l5=`�}@U�]v>\�B���w̓b�?������Z�Q�%�Yj
��V�aJA�O�O�#��e���eKX��݀1�/3��U�H�a�s��h�*` @�߻E�P�&��>��`dj��Ϣ����%0�T{�u�V���)ed��V���U�B��������n)ް�8S�9ܘ�CY�����s���1�ӌJ&Jp]No�y9(�[ι�麩�E�Q
���$�q;Ⱥ��O��*!���"Zѧ��W�~s��C�+.��\������)߾�d/-�)~k^�Ar��?<qsw)0�),w�e)��/�Y��T?��FL �eR��+Up���{�:~�~�������h��j��������: ��Wtu�A�����&������:O+S�gV�.���|e3gtr �v���&Ys&2�
�kh�5i������ZD�|�,\��	)�����݀�ݒ�N:�k�ǎ4K}*���h'����F6E�q5ؿ��O��6;�fl�c|�8�?r�c' �h���u�����+l�w��ꥵ̝�N��GX]T���J;�o4�a��nbď%%��6D�'pv��y�����Q0.㭆�rkQ��וb�c�K���&bk�|�=ԩ��xrEB��L�׸%��C^�5�v��85v;�dԵ��x�UE��?���*]�����g`j�Ky�<�_#��_r��T��#0c�nEGΈ ��dɃ�H�7���iY��WC��`]���*X#2��E�n�q+'c܁��Ϸ7��=���e�t����$2t�N����KB��oC�w�"	<@��M�&���R7VR� |e�CZ �oH�J����ayF�U+�Ӂ�}n�����BeUY��Mz�E�G�`�bQ}��gEU��������$�PEba�%������	j�0���PN'�Ϩ.�(a��u�]��ʤ�&��g�s�p�>�	������:�>���%/�cp�,�iI,&L[i)�N�8�k��b�)��3Dj����+����P����]���:w"s(|��P�R�j�i�p��hӔI�:��e��v�Vm����1�eK�A�F�ok_O�5�jc��t�0N6��������~<�����#])Js���E�+B}�Z�.���e�?��;�F� ?##�N�J�RM[��׬@f�f{�!�\1�9n���v3L�/�+��&��xֹ�k��ElhC �u����m1�k�j�Q+��0
������o�7�0ݏ�r�-�ʭ�B�h��tj��/�2+7��`�gR�;;���&nѕ���g����t�g��u[�=��߰|_f7��p�>�L2:�>yr8�+_����1�f��ZG��I'���\��@_���}�r�r�q�I��gwg��"��������56ۀ^�Y�ʒ��GT����[m��4�B��-n04*�K�1F�M1_��h��>��
M��HP�1!�A�N���{/q:O,�yLd��ŧ:~��л��b�Qǧ>=-����,�G�Q ��qX���
*e~G駁�FߚQ� �+ A�Oֻ"Y�:�-,�a��
�:�6 aDC��u	�A�ê��Q��f����>��/͐i�4�v�7�������H����T���"s��Yְ_��G��!�w��B=Jy�ƭ,0�R�V��k`�`��ťݚ<Zvs.e��f"�8AH���#�L��h�g�ߌ��r��?���K�Ʌ���bD�|�����>�gn �C��m� �^u��;��h�^��p>���K�⧦�6.���˧j�pܧ����S�鵾ڕ�s1w�̴���A�m����$�a�|ЕW%=��B
	��*���a�PÏ7� �����X/E<�]0
Kc������[\K �;��Ս+o	�N?��Jr����	C��X���[��Q_t>����[���m�H��������@�t=�c��o
5U�z��6�)���_.�z���4Lf�p%�x�W�gW[N���_Wp�lEڅ�aC�o����C�ږ�oc��6�hN!&�M�I���1�����ux�#�E�e��$�\�~��a��}e�d��'�K�?5��{CU��\�#��@촹��>�/c�.|���	s�s�L˦.�7��,�?�8��/�z���	�g��w��?i�=dGP����	PR��3��WO��n��E����ؙAH�DI�H����GrP�5��9[�ҧ�(i�틹6��T�8��_��P�e	�2;]IkI��M�G{�A����P=��eN.�w}%���l8V!d�4HS�~�,����Q��2m��`hτ��]Gx��/���8����^WO̒�ت���	(V�wm��\�ngb�L����8�SZ'��ݵ.	��j�[oi���|��`(�6��	ʎ�[͌����)U6�\&��*����^��(B��V�0�f��,���5����l@{�!�� ��iU�T�J|�vG�=TS�j=�{U)t��x齮���I0;e�L�Ν��oe#��Kr�!a�$Xw���/��R$S32�)ng@�f ��'�kY������hf���0ue��"���&K���t��elֆ�UږeI��0-�ڙWt�7����ON�}��?N�����c�~M�y
�ޢ�c�kՎ*�#�(]��O�`#�;Aj�@3}6VM�����f�}M�5�|��̒��f���T�
r���۝�D R�I�e�����S�71,�+����E��pH�o�b��k�Y<1}��'b�U�2!�E$�0��v���2��0�:&��o�tj�NE�Aڽ=\�?��P����"8^S$k%�r��z�!6"u�1;p ث����Q" ��QD��F9��0�h[	�,l��c˙���n�(O��7�j#
�ݫ��fӲ��NvG^�ħ	�7d���TV7�o�!bf=��0�#��O�8�S�&t�|��:��:�<?(�[(��u4�uLm}d��l����_��C!����ǝນj��RyX��6*��3G�����ܺ՟5��-G��F��h-���)���9���Y�R<9�qu�Xe)�,�o��]N"ک����ҼO|����I�s�ju�2T�֞t�bM���3XOxo9�sb�S�
���T6�-b���<�6�܇�H�8'�4k^Z�a�yx��w��zN/[b�n��e�q��9�k�m��[g�"CGO�>BQ�2>�7�J���p�N�%:X�e�h|��3�]�[X�.��,�Z	4S�pp�O�j	U?�]���yH�Q˯���"�*�x���H<,ˊ�x��y>�E%�5XУ<���Y���8n���]@b?�SnmH�buln���o����?N�z�Q~>�	�����I��2�g��� Ο�u7>����Σ������8|��P�3 �Q,�)�c[��g�)k�X��~^c�  epЩ�!����ܜj<�wG^��1ҟ'{N+���j�Ԉ�xa��5�����x�)0�[��B� [VJ���֩�� i��R��p��8��J�>ʻ����z�9u��|��_���Ukr%	?�gqD�n�,��n��[��lt�"�f��ߎK���2���̩8J���+�Z����R�j�Ƥ;���rN��9���� �.K�4�L<�V���%앬m��^3��}�������y���i�ϱğ��=�%�!���e���x��Ԅm�r�d����sT�Wɬ��a�~���n���GC�j�(M
���;fϲx����n���	E�(�	����8�4�<4C����>#j�+�y��,[Fa��;]So�jdQ$pGİ����?v����9�w7C"���D�滋�	�T�NtU��L;���RW�iF^��Ù�1ֲ�c*�A������/o"*��aOޯ_>!�چm��Py�a�Ӿ�{�	�&g�^D�ODM�a==AT��b4ó`67c����s���17���k\��ɮ�cn�Utq�۝����<��/1����y�TO�� �ր?B�]8"e�1868�~�X�E�jC���_�u��,�ۋAU��%˞o��1bМm���!*xC�������R�h��T_fH�(��~�+�L6�˚t�bu�"Zy�M]2GI+w����S�.�O��l�8�)-!o�=0�3Ӧ�������:/
��8Vr �jV��~��)�I��| �!�y��N�Ȱ��'�y�z���*��ַ�7�.XO����[���xPA'�|��`ye��N����uCV1�Iw��w�
 C��?���St�[ -b��2�����ݎ�g8����Z+��F��qr7hA��}��Z��D%�[6�M̥�4nH�]��T��T�ۄA�bߓ�F�N!3��$i��D��E�/L
�zk���ڀ��}�A~�,W�#�V��'G�zRC:�٘�Q~[R�vk��F��f��d��"ћ��e�0ƨ�:)��@����zcEZ�d}e����<HS��q-�_,\{�[ˬƐ�&<���1@j]N|�^�E���ʑhv���*�J�܎>��kR��	�6mm���<T ���Y��U,f����4�mXO���s�˺xJ��ְ.�̫KP=�0��o���{(���Ҏ�$���n�tM���A[]&�Y������O����R|�&YG�Q�P��k|�iJ�zr�8�+�7�_�jN�ñ!o��&�`P<M�M4@0
�LF�7D(�w1:�V�o*�+�G+L~Ů��pJĦ�j����	����T�q1��ڃ�F�c����k!�j��+�����n����\�$����h����wuU_2�'j`i�>��i�^f��R���u<��~w�G�S����5��/��t�����m�\��18�L�8 ��%�+߻wՀ\�:�\��}�¡�ᗩ��Q������ޓ�G�_q�(��d=n4ź��-�6.��4;�-�v�٧��g���i�)w��w�n8��'���!xn�Bsϻnpc��l�uj���pB�{�C����>���]���N�o�"�H��-kB �׼��*���GE��#֩��Zn���� 韼�P2+�A�x�`a��<z�p^�_����z7[֛=�t��5#q�AB�7R��"��N[rI�6l�Hoc��d�loA)��%=���~�%�� �lGrKm�2q����s^��	
�Rk�	�����%h�b`�Y�$U��p�e���m���HBM�����?�r�N��� h���bH���g�ڼs�?%B���8���T��0~����v�m-;������çqS(}�)-Q�n�x��" �w��gȚ�(Ʉ��#�I�e�q�S��ǟ��A�d�UAMu�	�C���/R%&�!���Gq4S^:�>�C�� �8��U�vqu�p2}�-�ޟ+�g!��@��\���zu��"���%Q4���J���
=B����),U���:^�0tM{���,��� L���v���f�U�)���2������4MFvf!���8�Fඔ+Z�6��N�-M`9�,o�>τ��_E��K'������.�G�4F ��`��<�Oac&�!f�A5�2��/=RI4��y������FPV��5m�!��NObo�oXc'"YS���0�<U (W AN�T�c{l<��/�O��b�۴p���vrU�Jx�G<x��T�M�kf��^`�1�^J NMG���yP1��A/w�I�1�s8�����AF#�Yҡ�(�ZJ��i�<�`p��!cyg̼�Y����cF�ar*C0��Y�)J H�E�Pݡb6�޻�*B�W^���ay��rX���J��sq-�2M�E*�Z�Ce�Qٹ�L�$��5���| �[J��.y�P3hkb���Bz��cQ��/1�f���4ݤ�Yﹸ2J7V�|EZ7�|��Q�
�nR�d���uą��6�E�xc|� =;�'�MO.�C(R�z�7+DX��5�n��f�i?�p�Le������ �Ű��j�9!PGZ��>�ˬ�eln�rzg17�X�J���/�Kǹ�	��/�B�6�v�/���FO�L�]����Ї���,'LI��]�et���uV[XS�u4�'�̐0�
�ܱ�U�YE�+�x7�V!����5Ρ�Z/�C끛�=��13���3�,�,(��s���?�0�@I{���E܁��a�/G>+��8ܺ�;�)��ꪤx���jE"������b	��`n/��1���
b-��oGg�N؋����k@Ok�a;B����x@,�i�[�e�>�jL Dј��?�Y���`K`cD���'+���&Z��iF?�nN�w|Ғ|��� �u�U[���5&�:q��]��A�Y�����JG��&�Q��7��J�3h;��,�2
�5�[���N�w5�].�+���Hc���k���`p林��ۭ�<�Jm"�4ry����1���v��ÌJ����S�^�I����*�����,mz��Ϳ����6�?)I�%$�ĕ	�}>���5��MĠY��B��v�J��
�|M� d��c/����%]��+��h�IY,[�Pb���`J,?C��P�^ָPv�@��wQl�#������a|��'�.`�?�2��[
&W�hQ�G�Am^�S�A({��*�W���:�]��������~܊KK�[l��,X�t&}���٦%��FcX-K��R�*��s���Z��8�m�'��;x���I`�̧k��Q�	�#�{<�v��6�Q���e4���z5"ɡ�	��\Mq 	8�����C��~jhC�FI�tm��8^QhI�����-9�T%�G�����>1D��'~+��� Y��Q��<�;�I��1��Q���I��@v�x��/i��Ce�څ(BݥQ�#,.���!�q�������.8���\����%3���}������T�ڰ�_s�Z���BA!��2�',��1!%�<I��m��QvЫ��:mI'�� �9x�u;{&�� ���|6�ĸ�r�i$��h�+��1��]Q�i�/_-�Iѐ�7�A&�x�>�-=�qC��~K�dd��^LbA��C��/M�EE�t�ek2xeE������]��ḁm�7ɞ�"�jL̡�X1�����H�y���y`�%�Xu�!�ik�o=uz�pm�[�?�^��[�)-��BE�3s�Xy�K���@���̯a�|,���2��1i� ?Xd����pkȹ���?�ͥt���F�	,�"���*�rܠ[��욋���b?���b��'qBl�l `�m�aP7X��P��&]���7q�0N%@�M����e���I+�x��sy��0Z3� )׹�����IT:CF��vh('�(�S�9�(ZaY �a�7�'c�_�2���.��A�墓x�g�Z�s�T6�E�GܑKdR
tv�/m'���i��jl�\��-`��ŋ*�D��xY��(���@���lI6^�8���A�9��I!,d�&x��M�@�$��:��In#ޜ��܀�;l �4�MI�������_;5�i���`l����ׄ�"A����Tz�;�2�k�/�D�{���m\�����J����MY�ʕ�D�&��ia��0�ӳم���OZ�$�r�~���=H}��5�}��Zk�+�M��1s<8}$F��bsf{�����n�b#, ��$�ʡ��惿\j>��?��)��&�kwaX��A�>ʞ&�W'A
����5�#�1��oEb	m���Ckݝ��C��@bW�߬�ћB��Z�V>39B�_�cb=��at�j���8���:S�Үcj��]rSJR�1p�LM�xG�v��$��NM�3��sl&���3]?�`�i�߰z�A8�X�#�{�h����E��${��T)�f��PƱL���^���z����M^ڳ�7����`�h�u�5�F����f�8?��+Rc3nې���ڔ�z3=��-�+!*ע$�r�'I�2WD(!�[��:��� l�ň~��
� b%W@r����qq�K��g��'���)�5���	��K6�k�QGqI.{}f1+���Q��J�B+�ghX�R2�m{d�͢\��LA"-�fX���!���K�\�)��՘�Z��������T�W��E0@V��E��FW#�)�˪��l�2ϓN���ȼ�WБ^I���G�d
����W���R��F�m����]��^@��ک������0��������.����	$L�&`��/V�:X+�n�mi�yV=�L�)�d�����&7��h�s�e���yP����[mF0����&�C
ٻs�aѓ!Ѷ��_�@yޮr���(��f�.�8�4���d����B	�2^��+v�o�c,�]�d?ue��ߟ�n��������w�Vf��#�2qyx��X=��t�)ԎY��х�w��;�새;5�hJ�)�A��*���v�A!"�h�$��O'ń|{���j+6�1#H�N0'�F,G�0+,��.�?졥��XX�i�*����ͪt���tO���0?C�vJ�zUZsL�0/��϶R~,���ð��R�գ>�K�� {=�3��I[��?}p�en0���U��i����;�$|;��A��#U%�_�,��)
���h���� .�_���n`�^�T���`(�����|O�cX��P���e���)TX�܏J1��V.��1mh+�u:ռ@$:�O�c�4�G]x̣��Z�C�dI�ۣͣ[�\:߄@ؘ;�Rc�SYJ�IB�����@�>��V�/k����'�HI�v@
�ǭ���$���2<�Y��Q�����,7>�/��ɒ�)�@���pb��c� {���lw���*�0�;� 1-G�o�<(le�Ҽ?����ȍ�+�������*gFS9w3W���Z�$�{1R�u��py���J��DU@_�R/�g�}�05��k���}0�lب`�&˥���@A�vC�E&��W��}��zq)i�*��'�R�,W�>��t���`�}Q����hv$��i$�Z�8-P�&���'��Dr�J\q�٧l4�v�Ou�T��n{���è�Ō��9�U&�n-V*M�᷿�7���a��Xؼ������g%O��x�j�6%a�e��r!���N�mL�C�7~��{�Z�z�m`�ٚ%���ݾ@�@�����u&���$<(z��ԩ�q�s������9}әx�
x�]�HؕÙ0Ͻ��BI/D��#��b�dQ�*ߵ>~�Pd2�k�5����m�LD���V���iV��;'����&E�R��Y�2{�����٫)-�ރ�?�����|�E(���s�8Z�'��Y.�-W�E�.�z"%�CC{�S�Ǔv�y�2Q}�ҁ|_�#2}��
�{Z�	��8��j�yd��e��>�:[�`�p|$�uΤ@T��	X��Y���r%\O?Ef�[ׯ�O:o�2��&M�*9�G�}9���.��n�ܡx���;އ�Fw�(�N>p���d��s�NUY]�׸��Q��V�G�=H�}��V�g�RN.�k�š����<�I �f[~y���:��O��k�Ի�Y�o�߼TT�z�o�׼�cI��4DH�>����lk�=r�=T�{���-Z�@�Z��l?аP�ȺYqw!�0 3{Aί�2��DE%�GM�(����;�e=�W�j�9i��\X�!���k�/6�,���l'�B�[�V7�I�׳��f��Ŷ�aaݰq����!�ڍ�G����NOeW�-3�TU�V��ݢ�B�rA��8���>i�4�]�������+��?.��k�j�4�d<L�h�շ��>s���,��H?�%)n�rO_*+�n �p���Y����"ӓ&�fXVXF�(���$������������D�=1�{���Dѱ��n�S�n�"��[L����S�ZTp$�_"�84��'����yb��.~+��،��Z�n�;^l,�7ǣ�!���Ϟ��.������|Zx=,,�j���ۤ����Nh�0*�^�`���t�dˑ�zP�zS��H��o��`TIzʾI�1�/��R�,��ݒd䞀@�%N>G�j��h�1�S�DNq��#nk~mؾHi�]؇��>�"N^�Ӿ�K�Aվ_��:h�}������~�����"�j�k3�=m��6�}8v[�K;�P�񅿦@V�T�dG��:qh�D�_����f���W�e�e���MC��z�w�̶���t8d�뜊� V���×�  ���|2��%5�V�g�I�wU?`%{�����qzP����
�:�
2K��B�6N�3�x��H�4ZD��/����ew1����t��i��iK�wDi߄f8�3����Lx��_1[�S�)g��=����Y�4�A��'T�	!�fi:��d�U�)�,z_�gywd�]&{��{�hl�7.������$��R�
4��!h�"�O�D��$�y��?n��;�a�֖���hk�4����69�o
��#�aM�N����7�N��W���A����.k�^``��4!:4b���/7����_Y�<	Ѿ�a���o�D�]j��IK�tC�Gn�#G`E�]�ڙ��S��j�h��P��a)<�{FK�h���]^�XC��W\�����Z���7:j�7��~]����kf��,)�]���y����N�.\kHUZ��O��}*bCD%7%�<��X^1��Vj1|؆��^�Q�(?nYRo�����
@�MR����89�OAl���Q���~k���W=�·�L����#��X~�#Q����7��u{+c-����kV��K~����E믵!ٺ]�d>��@�sB�p̫뽃kl}�^$�o�������E����u�XnM�y._��E��Ȩ��W7�n�p�_=���,���]���`Ӹ|�Q�����MS]�<E��H�������u�o�{�&�&�]���6��4�+247t��*��:�K��f+]�|�����]P��`7K��~d��fT��s��6�����L���$�B2y!`Y5�q�x��F���hq[�=�$���������2����E��3�/��(;�=�i ���6���9sg?�A��uÅ��w����&�%��Qi�Z����a�%���5��M�2b^�ޯ��['v�kw�
+,c����``�k34u �+��A��۫P8�\.	�"�����ai�]�_45��f������g�t& H�)~�E��6-�_:B5� �=�:ym�V�Z�r���qǧ�ċc��A��Vž���:(�jÆij�	�^�K%ܺc�	���N�������L]l</�;C�L���O4�^��nL}m���R�.�!ϕ��M��-�ic���\^ap ?��D��C�  :��y6o��i���T�d�����1���µ@#��	���!�z'��79H%<�+�k�Z�[��0Z����	��S����9o)�I�ԇ?̠�Գ큀�c'a���*�^��y��UW���@��P�t~>u:R��/{������Ӻ!�x����Dש����\1��6U��,BG�s_u�c�DT/�S�"�&kW��j�3��^�:�G�x �F�@�&�����5�Yi	��t.]"`^�se�9<YEyj��u�2��F{�ԭ�q*�>��1�r���	�U��3��V;ۧ߯34���(̠�Ps�_[��FFr=�����W��ːP=�%��:�W�s�O$q�y ���2a�R��J��k�OaV	���)à'��zR��O�'ļ|���t��X������ك>'�K	�L�O}XE J�,��gi��>�Ш�����|"2Z�{��q�du����� u��!ZV�WQ�	H��.��In�w�C*ѕ�|�)!%.�0�4�,�R�0��1}t(�=O�k0Sx�.� xcҩ��	�9�):��إ,4�����9m�d<�DL�+1��JW�B�JU�0��.D^HTHKT�ǩ�)?�"9�:�WV
��@��;"^��Ł��!�^t��z\*��e�!��=습��J����	�#/��Ѡ�奘�!�cޗ~	.ӂ�!_�LS.������EK��|`|t>E~�yI'�pd����	�-/������7"��(�WK�I�˃q�'q�X�<`_>!̍ץ�L�/�vlQ��.���n}ZC��KRJ���mu-k�ʬTh �
���j�W�Е6$�.��wޙ���5+/ (� �,wG���?9� ��'D����[�R�JR�sn$�g	�	�ԗV��X?׵�(y@��.?��L5�~M$)�>^��1��b��K��Pj�_j`Z82��d��)m7x�x��u�L'3 :풛H�g��⼞dM�D�������R�CҶ�\5(��{FLk-u����L�̻�m,�Ɔ^�ZO�+��hu"Ԃo/��,�=94m~W�(�m޽�vQ��աp��mؗڍ�j��_�����V?LH$ʶ{{}c�0P����ʝ%H�O�\P{�B�����'����{\�UQ�e�#�G�����e��pƼ�gֶ.�M�#�[�j,3d�!���ȏi�li]O��)=_n]�������}��2�^��K[׸ǊS�����o����Yӗ��:�`��rWn=��,QX��2��:o&Ѐf�U�ȍ�g���jI`Nv�36���F-Jq�V�]��w�§Z��w?K X��q�>9��R c�+O���+�!|�D"��<K�M�� $��6 r����l�e����4���0l_dѸ�%c/]l:�7��[ y�h�8�e<�u�;:�Ҥk��e&wѦΑ�Q��3�
k~ڒy�e5�Ж��L����q'D��%�	܇�`-�k~��jR�5��Bo��]]?z\F������f��~R�uu��t2kؑ:Y�l��$���c*׎����:'�me�k��O� u߰ɕg�Q�4������U2�8� g���Κ%��
h��&�}��Yv��g�e��WW�����'���|���%�Y������N������pHN�U�+Јk����>E��!	�'�i���9��"'3	)��e�+�j_�ƥ=��5�4v�����*Hj�!@S'��|����}�!��Dw+��J�)=:&E�3FjAG.P&�ac�M�Vk�'�&p�6�L-�����n���:�������7���{�Ԝ�e�l*�4��n��֑�me����j��9��m�����@�I� 2((����v]Q��\��h����n�9e�>�+i��	���Ʒ�v�h�<�68 !-���BO���f}sS����=�3�ް\w�P⚛��opr��lĴfK7������ʹ$� ���6b�2[�Y��.J��w?�߃�P�R0<!|\��chHsT�&�9��76�B���o���[G���?�������j�,/+�fn�C��V�f<ΐ��˘4U�
�� [O��]�]�z�ld|1�V.�Cj��=~��P@*A|rR�����=������b먍�w�@�2Ju��u�&��{b;�@�Y�_�� ^�i�l�K�F��=>���d�ҹ���6�4�Ƶ")^$�'�9����u8�r�t&�y�T�J��F��|#�KC��U���V�"��[U�$m*�M~�*��(����<	I�ͶՁ�^�>�j9R,3VP�$�Zݘ�$C⣷����h�������0�1�H�Z�ރ.�=@L�{o�sđ��.N�_10�^G�1h��յt��xq�	�6p{���?���y�_�@�"da�q�KMF���T�f�f�L�$'�K\������f$3��xJ�,��:=��8[-�oy���ˤ+4�P���?�k�X��౺�/����4�札:�ն`�!W�@t'���ߠ�׾��~�t�낪�3��5���>';��v����%dk���a�&f�fs�x�]ٮggJ�z���^�OpU�:�ĸ�l�����> z��P�׾�O�-R8�w3��fd�%��|�uI�q��4�������R��bQ��*�E:9`N6{�ץ�+T��$+�,����P���("�lh��D$���	
F�7��S���'E)�!�Q�8��Q���t�^&'�*�3�qb����1F�Ta��ҙ��
l���8��։M�z�!ٚ~��	N2�����OP!j�G���ҿz9n���?-�Wo,�8h``��m [~���	�E1�[;���*��
�g��E�U��^�����ӎ4�m%l����)*�$d�x=-�WQ�e�5 ��P���3q�>=�q& ��D55z�oA`�����v�rT(p�:��L��V2��*�����7�@�����M"-�b	\o�V-�08��cW�� �X�۵Fˉ?��KC4��h�9y{��5W�v.:
�GN+֒qc7��RG�c\���[���7�zł�O:�)�!�ao�4�_����W�Y�풋�3	��]W�)�;}��f�?�F*�1�����!?_P ��_����~�zG�}����ɥ%��SDf��_��S�nO�xk�)pWͦ���5�T�0�1�_�2�=��(KYX ���f�Y���_��ѮSR|�D/��)�5-q���v5�=D<����M�x��4������t)t��H�* �<J>�e9��_q�#9�Ht�|�8�ح����2u4��N��V磾߮sGj�y���G�=�D�Rl� -_��y��]���jew�X-���������t�M�ݪ=}��f���#��N���Ļ�A��}�(��
��h�}l7  ����(��&SÓe�� ap S���#�����˷�㛳י;f͏ +�c��|X���OQ�|���o�]�xV,;��k�h���L9���]�vW��<�A��||�]Y7nN?�N<�%LQ�F�ĥ`�xb����|ӣ�z �ޑN^�z�&kɑw*�ws������p:r�����g�@�V%���X$6m�)���/#	<��m��E�?Sd�Y�`��?�6���!u�h\#���}�"�-�tL:�!r��ၰT��L�	7��h�L�}b}4�ވ��?�'Us������ 0�3��fȥh���B��_��mVz�B˙��]��=:@�&���^�e5d���F��-'������H,���ԍ_��Ӱ�J������NWo��+��|.���X-�B&��Q�I9�Í�w�2�^t8�v��ߐ��n=�P�d�x��&D���B����{�6t`���������Î��t\jy��)��Yp��R�V�z9��A�jr�����"��s��GϷ��XQH��-���)r�	�(����tvH��*�[8P<đ���i����t��C�
ku��CC=��V��"[  R%F���88("佭Y[�Q��4�r=�C�[p�j{�Eu��b�4��U63����^������E�\=w���ە��e�p�[�M.��'�U@����w���tΆ����#����m�"�:�����������*&E�wz���8���t�4y�	`b�Ҏ�,����&Զ �?�w�YQ�h�<׳d�1�������}~��Z>��W����IЀS�m�A2�
�QcrS�D��z{҉s�~H*�i>D�E&��;*��_�2��:�:I��P�U����/����)#x>��ٴ��`ӊ\�j��xρ��
T�{.3pPj�V�g��ZY;�j���!�[��6=��.��� |ҋB����b��/\�Z��é6�)��V�����E-NQ-�Ν$�|�2ϝdL0喖�J�.v���K��wH}�Y0N̐�L��A�*�_�:�d+�PX�Q{�4d�$���W���Ҹ�Ტ7(|5}�*ϤH�;�f&1%f�ْq��J'�+�}69�E�	`�V�5�А�����8����z��0���\ϓ�k�P�M:��m����6#nՂtm0�$�}m�PLMA����8�z�'���a`�;mx?�h01f9��6w�yۚMH7o�{��4����LJ�3l2n�2��ܝ����j\˂B�����I���P���rI��4�[Ճ�]�O�ΈC��9��I��"6g��TY���	Y���:�y�����\pk�f~�*�DkS��;��8��x��!�7����	}X_v%�,�)�\M�r?�\.�q�Lc,�L�o�ېˠ�|P$����st�JO�dH��=��v�T��@�d�j��񿪚TK� ������6���&X�e�"�+ޜ��L�Wa�P��S�F��������MD��U�9[, ӛs�1���{5��I������+�_�)�\0wQ*_��{���l&O���4��rmd�ˡ����RA�a.8*��k�dy2`̫s�����/�9���0������:�v��k�ɽq�HN��Jh���
�=.g�٬8OU���S}뵺^�ϡM�ʭ>-��G���d3J������F�p��eٸ:��v��Zj����|6p�G��;,��0	I��Z��
a�-�S�~�6���X�x
Z�4uN!�}
�"��*gj�O������?�&A��μ�ۼ��i[���u*�&��!9�Y5���T$27�A�vҧ@�p��ʏ_S�:b�j��: Hͥs���Mĵ���HR��f�{wJYK��:ia�j~M�ZŚkM��0���=Q�?�'�PL��h&r�)(+H9�c�3�$*� �j��SG�Dt̻��\=&�u�u��g�Z~�bwo�X�(&:���T�$^q?�����Y�`��Nlτ	��	�d��T�%�DT ���CN/��
�{BK
iGw Jb|��?h�A��O����b �� �V���	Uޫ�7�M&@���W�P��Zd�Y�/���dKp�oVH#� d��!����Z��g+g�^� ��� �x��_A޽7Msj~ �uf�N�I�S�'�����V���|ƶ�
+�shheX��z�V}k# WK+�k-h$���\?X����;�r�66�b!E�՟�ؙ�"���u�� p"��;�L�d��Q�pEӭ��-�3����g�ˑjm�~+jݜ\}�&��Pg�6�kpL��"Ա�2���4$��z��F�[�*y���F�C%;4��!,���0��1:\���<���y���~!\�J�mU�A�3Y�FҸ�i��A���-�h��5�������D����^���bӷ#��Z�B(��:���bֻȩ��J�@%9Ġ❻|��ߏ���������R��Qc������CfmҪ�#�������/@�E�Шh~����ױEQ~���_@�����2��ؐd0}|h�d?��Ѯ(2��gmWq(]B�H-˒�>vկ4F�@����:�!D[h��;��av�;zgE�l'q�TC���m���L�yi#��R��U�.6b����/�/�ۋ�1�3�[|2���O7X�s	߹O�ʯ3�rw���8r�R�V��>�mgt�/�Գj�]�T������5d�㸕n���I[B[���	wB���Q�7�]2��>����J:\I
G� ��2u�����ҝ��D;-�2����
�V2o�ѫ���ۈ�g�d��ĥ���Ʃ�J�-"A�d���E�~��wƔ��t}�
���p�_b�!�N��ڻ��d����$e��U-
�����9�9gK�E �nNb"�`8�D,�0���$�	��PZv�f�i�0ky�\��ŏ_�ӠX��+�N'.>r"YC#�x�\]t���#����Qw�d(�J�3�-� `*&��w�k�{6����
++��@3����h�D���D��(��|8��T]�2"Aˍޖ��`:�ې�>s���%4e�DW�auE �2JE	�|�\��(6�+)��x���7 ��	����Q��t�v�zY�͚>-E���8H��"�<O >���z�B�@�����C�`@ b��xG���u��� �?��{�1�<�C�v�i^����Q-V`�<.l�E��X׈$�%��TQ�{2T�����3~T�8$ArFe���_պ�:�Ӵ+�N�<v�)ں��7���|)��A��&4�Zk��E�z�<�U�t#�V�_teB^�4���fǶ��֌�dHm���/���t͹Q�*��n�"u��۾��T����}.�������L�T�VG�'�+���x��颎(��Uw�z����zzHn\�b�(�Hg�UG t�v��g-�{B3�d���*D��<�ZF1�M��C�As�[(���!���'Ve �"�S ��(�&���]�	$'�HFQ�M4��/o�|"ɮ]5=K�Ad�ጣ'���������ޥ�>z����u�G�[���)Y�}ٟ���ci�x,�J�7!2݋�i	U=�5ť��{��6�����.N�W~ۨY��k�c$ɦ�p�<��t�^�
6�7.��a���d��r rf��0�3>�\A�0p� �'��<��B�u�)�lâW)"�ax'Kph	6|�	�t�h�'(r�2�-t�g�5������������ԥ������'��W�b�P�ž]��T�W������� ���:]����/�F���j����B'�V>�UX_�|-����J��=�;�w)๮�b�s�KZ=��z.w*���}�R����I	�N5��
F%4�]�u[��
d���ğq�s�^\�E��l|�hBޏ�����lk�V�4ռ�o�!:E<�-�3јDU܉��؞���+�@���GPC�8:����ݛHE��'a��Tu�0<�hJ��N��;fQK��Ec�}�4��]��l,��T�+�>�=Jx�+]�fYK�0� Hl�S�),���2U�u���f$q������ˉHv	!��xg��t�&����z%%L"mP%��K���n�H�P���?17`kY7/�Y���+x%�H���"y�v�c^�S�?�
j�k�*1]����7׊����1��h�<�&U�*�NB�����%sOm�!�Pv`态��ގ�>���w8Rд�!���#,�f���\�����	I����o��ɵwSMJG�*{�M	 ��)�2¶���;6�pd^�����P����}�ۯ�)��w���骐�Nfm+�,b
�[��J��-�̎���bC/����m�s���VnḖk��R�=�n��z�{'ؿ�M�1va3Li��s����Xq���J/��S8��o���ǵ�{k�9o-�����vz�.�Gi��e���j����_��2�����V\�I��8:[�ߕ[�0���m[qVC�M�<����������A3IpKau��:4:�:���8�����ETC��5��]MP�ÅETq�����E6��W�lT�g�Q2w�5�#lA>�v���!��A�N�w#`Lp���i�o��'a�i�">�����Q=�Oʼ+řJ^%��[.�b� ����䝑���y8(�S���~@:�с��x����=�ԡ�Sd��X$��u��5_b�c<��~���j�JU���*�se�N�6{��͓˾�����-Gň�R��1�'Ѷ?�{�xO<���Lf�C��><���<#1q��Y4{�61�ҵH,j޻^eXџ�����$����B�k����"8��gCY�ڢ.�tH�u��Y.cŤƧ��2�K� C�Y1е<U�C�]8Z�fv
�Y����� ���i狮���
lCg�T-y���i0�)q}�I7v#;�
f�U+��եMKxٷ�naOz����U/b�"�d�9�2�!���2W%��hF�q����^��rF�'Vt���ù����V���UOҫ@>b`�od����1��bT��Ƽr>O�Oe�����	���4b�OA�8�S��M�����5G�z�Ѧ�!a�����y}d1xu}֦�ֳE'�Vh�:kG��X	�
MA�r�v<l�/��OÇ&2�OO&�P�38!.��r�
$B���|�<?W�*�s����L�H��*󏅸|Uu=����������Q�scG�Ov�b�DT�Ǹ{�փ�iD� �Tn!Г��T�������VlC%T��ծ.�
�*`���c�Բ���W�JX��C2���՟F�ğ)��p��Q�tr)TC๮g�o~�In���R�[8&j�oٵ��69Ob�j�����ͪwa������3���rn�dⳆ���gz�[fq��Ad5R��k�a�t4�D�k��Q!�c�AZ�r$��v0���$y;ě�eV�m���{���oV��_�]3Օ\�[9���&>�mv)��n��1t��1y'x��[�+[Tgp�h��̏Ca"�gb��� Ǳ>or�4��bέ��ҊgWm y�7*8�5mUx��D����w�&ڼ���_��1P�%Nu=��7�ߏ��D4�!�ύqI;kwa�"��������F�:�Za2ga��n����|��D�)�A���e�9�4L�r\U���$sS*��V?��	 ޓp`TV�Vɩ�?��5���~�˗�W���hἮ�3�=�e�
�t�aQx��H�IS�n���_x	ߚ�=gޣ���`#�W���F�i��؇3Ƨ���\0(�I=GRkl)�T���۫��Z��j(Iǉ՝&���5d���㗨�^���Ai�?N�Zm�oT�^�7�E����h��yd6g��Hp��x=���r{a�����F�D	8lW*z�x0 n���������T+)$�(�}��m���J})���7n@N��ʌ��h�m+�-�����=��ǽ����</���<_������脿��}�F�i��Z�2��=
�/Z�x](����k��*������FXD��ҡ�D�p_f�"�;88;�c�[�9�9��b�᜽IW�o���O�|{�~X̿$�����Ic�M�g���v��Yy�!�D�RV�1�f~�6����0xO2���:�)��P�:��Z���q�9����U���~�\�,W����.5�w~y[�|��5ᢶ逨�ӾҳS�/7��S~Sp�!z4�z�m�ym�{��a��V����̈́
����R&��'�N�t���g�Ra��v�TX{�,�'����3/������%W�<�p�Iʎ��X��>e��6�����N!֐uwI�b�˱�7p�U�m;>A���ꞓ��4L�X�Y\�WZz}Q��n��쟹!�:�$�o�ĕ�HuO�	=�w�oUkT�3����	D����	�OF$Y5�E<<9N�Y�]W_P{h1���u����{��cH�W����?�5�F�"�w$�4i8��8���b�yIJ�{T%`�&�O&�kJ��|Sa�c�Dk���n3�4La�MS)7)F��E@�H���P@ �?���h��;�$i%է���]����	=��o�`m����e��_����t�d�}s�Y��J���(>��î�ꩴ�l�:���9�([�qO�m��~D�ӽU��Д$�y�K$E��&�t��H�1Ìo�-��'Ֆ���ጷכ|	cx�������2�z���tGg���f�H���f*H�T-uΨ�L��ޜ,�S4���{�00~L��JmN�(��N_J2мS��0A<+�4����z.{hlS7%h繧����_�tc^��ڸ�Pe����q�/��>�e�'�[K�o����m���"Q>yW��,W�Cc@�g�'���9�Ue����J >�����"����}aJ�r�ߏ�	�*���l5��~�%c>�f~�HD0���4Jj�y j����3��%�r}g�^z��)Տ� t��s�s5���U������
!��~_�
���a��P���d�}m;k������I!=v��E>(�0��{]�N�� ��q�0FM��c�lʅE"Q�i���Ţ}~�>�$��vݢ�1�R��Q��/��B���1?%�e�宷y�P�*5E 7\v��� ;ơ��,��(�_*_"X�D��76;=A]V�q�t_���0���Od��X_���%��ޔ��BZ���]5W��/\��$!O�'���p2 �|L EW� ���nE]/��ۺ�c��+�����폯��ģ�Kb?c��*,\+G��`j�^g����;�Wh�C��GV�����(��j]5M��'�8F\]��
��\�Ծ�i��pI�y2�����5���퓨�[�)=��%y\����z!�','�g �9q���� YoTi�~m�A�P.�G�{��;��G��0m��v�&8v�=�qRٖ-�©���R�&@g��1�5���ߓP�>�RL�o������!�0�������+�o��\G1�Cok-�ħA{���6�T��V����B���m��l��	�ox�{�Q�Kٕ{�[����0�;���q��ޗ7�:����w�S?aT�\��7tZ�����)�h��,���f��.�\[��[�������|���f0��lh��~��e��v�)�`����D�h���]�[A}�*������V!L7���
���7��9Ù�{��: ��g/�w1��u