��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&Y�%�ddؐ������&F퓬�`��ׯ���+�e:Q6W��$�I�Q�	?G���}��h��E���8%/�_��wc����7I�T=L4Qŗ�?)�3'��P�8
����V�N6t��G�CW��W��SjK���b���������b�(��sQ��/P�z��}������'�4/%i��ɤ����f݇��(Kx�]ZM�����]*"�����,��23x���c����Ʒ}��<�6(���*@J/�ӷɨ���9�'���$��TO����/cD4��D�����|(�{����üQ�w��%ϖ{ٛFd�18�9���M"��(����	&l-,�?w�	�i�q�#W�n�a�-�������	x6���,�q jT��A����N$�vl���jĂ5�Ө���{���z��q3j���aV㈒^#�H��H��#�_4��&�td:z��r�,�^͚,�9�� ɻ��1'��:Q�n%Oܭ�?� ��l9��+6�A]��H�ܼ�[.~;�d�8A�z`��]:Ӱ�(wSht�����ce�0���gSO/P����҂�b����\4��K�X9�w�kt��_�fz�����Ɲ����hM�H��t���ۊߡ��sR�g�f~�b'I�P�>
����YbA�a3����Ž�Nh��� �����v��k4�l�@3+�vA��l>%z5
�J�4T�w�$��2[����=w3���?t��@d��=_S��w��z�&�l䖆*6d�9��L숗��#��Β����g�m�/��/i���H@@N*#Ȣ��!�1TJ�R@���&6��l�9����l�dOKD���t\6U�ڢ~���:�c=#w�"�d0EF�X��Uښ:�Q�a�s�ZVʨ�3�Aho����b���y�9`����xI !1;~�Kd^{���ͽ`�������U	�����bQ�?r�U��ãa^�C=���V� rd��g�!�R�I�ơ� �ǔ�{��O�k-�͆E7� �:\=�QѲ�Gx�C�g�n��ݿ��:`"��F�fC;�{J^uź�p`��]��:X�6�(�.������v�;�C��#6��H��/[�|�;̜��Y��i�oC&|�	5R~b�x�l����5���*CJA���j��Ǖ@=Ap�!�MY�_._�DS񁿜�Q�8��Y��/������P滺VֱORL��}A�`~�aj���)��&��qYy���+������c��HV'Ml@s&G��n�t#�Wa�+/�&�o�V�@/��.]i0Vʑu�a͵���SO�@�~H����"
�ޯm6�x?:�"��t��>I��[�k���6\����=���c�[с�7�o	����"��㹨!Ic�k'\�zHQ�������^�"����Ut�pk��|��	����t�e����K>���֏8�$�zh�۱_����G��3����9�#�==?��wV�ߞd�-�+��ʜN"�<I�V�!r=�3� �n�����+���OY]Ȣ	��;g���SE��ܧ>&)p��i��}h����6�<R:�L>�b�ͭ�J��\mH��D�Z�I����M��-uY�����9�?�R��1v/�.������>
��N�r�4�n� Ќ����suB���:�`e����8�]7��90$�۟��&Dv/������n3����㇅d]�%���r��9=e�!���Ȋ-�#�'D��/�tZ��co��-gi�ĴQ�rƉ�1��J�Qf��� ���?�h�k�\��U���=<Ht�qD��be���l�N���N/.�g��܀]^~T�O�L����\
=z,g�0 v9�K�ĆD����F�}���	@z]<A�-탆)�.ȰŐ��Kr�vG� �.^d��1�%O�"#l�"�t:�L~Q+������4V��Z�����J�*4�r�]���4m�L}CxĪ�S{e� �yԪ�w?[�7A�s�"F+%$62��P�쵼�AHl8 �����o����a��C{>j�˾�'k٠��F�g�Pj�!��;����Y�	��W�����7	;>�<�,"�kܱ�B_i)��&���m�5�^D�����|�8��drX1����"�x3ɱ�lV3�Eeo�������].�ڷF�T���n�9�\��%+�DX>j�?S_�+SpBx�[T�\�Z����XL����S�;ig���I�4�4�����x �0!�J�����"��:������0u�t���.+"zۤi�u�G���������끠_H>2���*a\8������&=��fl�������ی9���sC�=l>�*,Ux��)\\mc�1�5()�1̴�6-RM�k�]5A�=��+�i#s���w�7�gd�4�:�@U/u.��lB��d)f�j���Tu~�� 5�_�pt�L54T�Ǣ4��R�N�ų_��2j�l�������
����W�P[R\�=~g��iM 嘳yIB̲츂�i�P�̹p��8Gp��h�ې�´NMT<5��13��NK�_�V/>���q��#PQ@�k���l�e�� i�m&��{ޛ��)��9��ar����1)��P��Q���aF_��.���7H��Q��:k�A=ɉ���#t���.,�d���u�
>��p�H�/Q���)}޺<�}�\�0��D�w�����tN�� �c��H"'�'���5�����iXX]�e����(��?g�۩]����ᰅ+�6��邲����������Ԫ�s�Kkd��P�tוֹ���b��H�	�	e��dpa B�C����?��N����8��C߲�r�?A����ÝUK:��9�!cm�S#����=�_6���l�$l��|�=���FDʗW:']:�����穓���w�9�~>6���)r;�x1R&�L����*��)�0cc�!�ͧ+^ae��e*v׮'������0p� ��;�q��hJ擞�z��g�����$X���~Z����.��nH,+Eһ��c�����ִg�&k��o$������������܃�����'?��+�g7� +�E�<�Ul
)W3N��� XҊ)f��ohe�Jn��쐅t�� Y�A���W*����&�������9q,(w4���Q�'�!E
A�w6>
.�6�d�(�x��7E������`�ɗ7W�A�J���f�R�+? ����i��k<΂�%�56B���%��Ȅ-J�/j�.�@ycp͞��5K�F��L���3�/vN���q�U�>l�G�@x��K�5�Y�z4�e�p4Qޅ	�bQ�$�q���`f�
�`<�4*y����"fc37��C@��i��I᡿��k7d�)\Q�� o��ήY��Dz���h^g�,�=q�Ђ(�/�c����?�fQR�-Q�1�����j�g2$� ���/�Y�"�G(N��#��Dj����(�1��ٟ�:�iz�G(�A1�F�"!Pe�g��{lj���l@��ܙ���wa��uAZ?�Phg}�n���iw(_���ad
6G����,^����쓋��h�erI����|Iz�jB��0a�h��pБ���̂���*���J!�n���)���j�r��+A/T
��R:|�,�3$1i���v��Gq�A�u�zU� ��	͚Hܞ��,����l`r�Y��a�K���qT��S��Kf�ğ�O�C1�toOd�^2ݾ��F��=AbT7%4*�ʈwј'=�������oC��T����$8���ܯT~��Va��s�14JL=���
:�:�.����c�dKMS�g�}�`���Nʣe����=B4�'���碢��s�^�|g��-�,G4��>�\n�۔������x�d
�?<�3+�z� ��=��SJP�ӊ�U�!����\�)8:g>�g��2����C}�n.&!�M!Ђ4�_ԓ��������{D�3�O�XA�*?+��	�