��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{���b�e��_�@�*��Ht�'�>��j��vm�s���ӯ&1�)�z�DhK:��������j!�I��(�+2q��}>�̘v��0��;t�/��[b��9;U�n#֛s2�R���6�8�(����G>ҽm���h'F!se�P����p��y��{�2�����T�	AS���}J�X�=�l����^y�� �.��S�(�˯���<`��"dX�h�}�����L➐�S�f=���Q�~����t���g.+D%Уb �ّo��͟��ԑ�~]�p�`�;�=��j����!	�� ���L�Ew��`E�&���U��K�M�Y��&�f�&������1�$9��s{�QJ�|�:6W��(�8I(��jV�Ј�X��H��Z������Ky-���g�$��
n��aJ�4��;O�~�k�='�N����ȥ�\�Y%H"fW�S'1	B�I]x�HF�B��Y��Ym�^��E�IZs��iv_�V�h����0���g����6��js���m��ӌ�*�,C�,$?D"�+f����`��C��2�����K?ljH}Z4r�5���	B��wB�i�h�&�f�S��8#��>4��g��|Vn֋��M��ݞ�ĳKJ�G���y���Q4-�lZ������!��y�S�)m��3����t�=N���XW��a����8�b�m�cV!w}���k��#���� �G��o������g��5�Uq�ݟ��p��<i���Ɗ�C��+� ���)ɸ�����T2���)}�F�(ނlg4��"s�\�2qJ)��ܶ�,�r1�_�9�.�s���Ҁu_�.��r��$�/l
�tRj(+1�~���� ן<wW���#�̔�h;O���L �69J�d��u�#u(|Ev��H,`�Y�����H���=,�D�2�0�NISY�*�����\� ǝY��������}�+�=	k��T�.���2�Б>.Ǚ��@\=�9A}T�6p��fh%V��Ϲ|�<�C�`@�%�td1~$�R������4)�X߾�Op/���D"�g6#.��:���c�u�F��A �a��\��������f�YpӋ�ˉ�)RjH���uv��8#���(�;�����,��Yeq�l)qn��%0��I<~��ߚ�cP��̇��U�m�X�^�DDt��o[�G���j������ix�s��6�j�w_�$,�^HEr	\�
MT�ߊ̎���/BU\�Fn�c�9i_ %�V�}k�je���YaBqr�nUT��b{gHa�
�=QI�_��Z6R��@���`Z������&�k����r¢;�u)��ʞLNKC6ՐPtOd\vu]κ��K��� '�$��օ��͍~�#c� ߫��׿��?&nmٿĜx8r�;���"��$KO��v�s��\q�Mrђ~{t��<W��h�RG:���.-���"1�LV�y|�Bi�QnS��l�Q�\+�oJ�i�a��g��U�i�`|=Y.�┝�.Q^��5�Un%�|��f�$�Z�=� N�z?˰�ї�N*�L��$3|@�v-��>rf%�r��] �^t�_�:�������6�ah��Sb���������k:��&t\i7,������6�mT��\�)��[@��9��Vȹ��=���}lǄ1��Ce��SIN����˽��e���hQ���9�-����j�	��$�2td��f� �i��LٻS4Ƃ�D;) �BJz�@����x��b4.�LlY����W�XseJ����1������.�_0WBqK��jow*Z��]�Ѝ��8�`eyI�
��/��Ht�G-�-Ֆ:���>�c�!� �Ke���C���u-���y�Ci���ʢ)Lv�R�,%8�vDN�KJ.����� ؾݿ��
&*��i��:���Q:B2��`r�vↂ�Q�d���CC�/rg��#Dt��c<���[��_EU��zw%>ά����LkC큂�=�Zr�3C�O�&q�Y�[���1aX�!^y�CS-�?�������,U4�8T.�T�Ląʵ��@�NE��G��윚Aym��|�h}Ƶ`�>��@H�}�_���FV��	�Ju�?�Q�cEo=}���_�W�:fgy̤:6+Ǖ(��`Z�