��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,�������_^�6�3�@�RU:(�3�у���aL� }5l����X&2��\�+�<��`D��0|C�b.0����,��L2���\͸�~��V;��_�	��e�TaAF�,}wN�aue��̖T�1�d��gY�j����#l@�j�C\��2z�a�!���>��Qpo�Lc �)6"�N�x�
��YY������ߥ�?���/��H��L��f�i��0���x��Q�ǅ��ޚ��!��3!��*a5�����!�6ݛ���˳X�Ycyl0{"�V�gp�;�^�"%��{p�sA�-0���۸ƹ���'*�o���o�y4E����mά^��*����P��0-뫝�( ��2���iq��F����vM��s%��3m��Ӝ?�^�pckN��L�҆�Z{�s��	I�^?��hf�����j�+��_�1�S�슲�]�D&��[����/����Re�W���JyY{�dpHG��6�I���ؐF�ǜw|<�q���f����<��JBb�k'�S���	v��R�C#o�4�EL�ba��X�*�r�>�Y�����I��kۨ���^+H��5u峈�'���bR���1V=d@��1����CS�XxyX[?�6P��@����5���];ѱR����ޅ��9U�>w�qy	\��&��QO'2��
m�k_��A�\����/=	o{�G�]^��"Y�s�eN���.��%���I"���\3��`1'={e��>Uc�Y�b�ܤ���G]���̣�Yγ9+�|��C�@wg�J�z���z��'�J��`s�p�a
!q���N�Չ�����Ǒ�Ґ��c&N�x�0����ӥ[���C.i)f%� �6+&�ɝ�c- ☰g�U6��N��/������{�/��].Q���Y,�!���؅A�3u��A>Xq;q%���E^��$�t�a�{�<4l]S�b�R{<b>R��-f��1�����H� ���O6���'d��?e������0ϦX��� ��
�}G2����7/<w���(�.���U�}�+*r�['���ӛ\����2\�N�@��|�`�� �T.;�������>u:�B�<��TL�t��/k��[�$�B"ee�;�Y��S9Ŧ\�-gPk�����-��G��F��>>�v�&v[����"n������L"��}�����~�pp���ُ�	�{H��qH��?��$ ����pfJ1�̘����r�(���8�E�_��wSS����S�,�>�=��~K9����=ThE�l������^�=��I��< ����x4A�8�[��3#��q]Yݸ�P�dd��Ё��{��:Dp#��ﱷ~l����TN̸3��������q���N�����S!�p�/�<�+齄_�$l@kqV�B���~m�� �;xU>�Sa�l~<;�{6$����i�����h���'O������0������S��<ۙ�c��ց{���3���{lb�|�� �1e�����'��Ȩ���>��w�.����VkH��ђ7�E�d���b<���edi5�h��+���x\�֊���ͻ+�Ȧ�wB��},a�"�	&�M�vʧ��<߿Yȋ�?}m�,28I�����~�����"�= �Ũ.