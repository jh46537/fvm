// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:33 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZhA8TqX1c6PXSadP108yEy4XgaLYSviPTzypcP/fVR3zoyXGZmZEshiB4vGiUjjX
Wul2ihyrXvvc2+k7wK5wUNda6iU/9louWFv6Zhn6NihNMcdL3FRWOIlLpBIpsOgf
HM6Cvv0UwWlEcqW3FCeDnd34NbiQWQmVjxliHbNqBac=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16768)
I9HjdPUJGeybdwjwoZ4BlVkewcGkDCIRX8zGPJhi0rnMe7lxwXQcUhpZTEIBMmYF
zCvFnr6WrAkJ4+HnXgSoxn6VwWqjQtrtw+TYaDiZu0AKEAelPueb1mkaRtigvYwb
i0w86EgEhwjlXY0N388tZ75V/inHskwWBNV9HNQT0A52pifwnM1+ElNc8C2Rgtpf
y5O1PUo6TfghUZl4Yxs729GMYbx460masDABbgfSUwov5qsiIwopEYEzm71Tvki4
OQ73eS/wnxDkATD1y7FQOc/FB3MDrMwwONJaidQOZ/WKi2RhpUhUTra7aCW3SIG1
FW0MRVvwzavBA53ta0EPV+/k5B60GCI3Hz9xiGaVDCMMTJirtaCCgPiKa/cM+2Hq
7c5TQ/V13QGAztrDiI/SNkgcIxiR9/PwSWcQTGVwkOJXbVobfNNKWc8biWdMIDdH
JxsIX759b7jM+X38coGIMgJE8hBpbpSgG7P4H4NgSsp6+BoWajSkV5G1CylFiGgn
w/JRCewmTkd4YghmcYW/g8VvqELPDQn8uwAxI5q58hCIj68joXBMHrCtNnGWyAKT
wprLzhDrq88rm5hhuurFuCsPl1WCqUq39W46WHUnxXev1qSm/fG5YAjZR8DzlEsj
jbPCGiaUftT+8+cFrpPrxWCP/9Ls7urRns7v1a2FHr0umzNnu8EHmWNEUnBKrh4o
N3usnMbTbTdPVrD6qbzj2syTB7OTiwfc17hD9D1phpo1gvwVQg9gWuaHkGh4q1Z1
dcSjj7H2wshprzhsME8syBgIWbryRd0N9S/pQgulOgkAqpjyGflYj4WTtnbOTih9
zvpk3N6EayRDifMnQFs6ZN6mvCs6vm9VrS2LsPx0Mqt0I+UMFWIwLBmYSDFnxQ/W
bhkgi2J39USbRHtFEh6onJf1NwZ3cPLbyuhYkmooRXP3K52m9+DcYU5AMoJQES8y
lVWwJKQN0UjZ1KXRa3qGMWXub1aUt37/gjLVlgCj98TkJbNnEvy8QhRoceCcDAWW
Ciy9be7LC6Rbn9ef7HripUJ0C62z6uT47QRR4FQUZHfmIIWvaQ7DI5DfmUquqnJW
bnKMyO0RY35YNY69W25OkuQuobilNQIh5D12V+cqeT1NfK98IJ+UKFp9bMDEsDmY
wUwVMD0H9Xz2DjiiTkb5EkT2fhVQZdv/yLe47vMBlAFUK3Dr7mPQRUQqJv7w5OkA
coP4MBMTEBUTUpbw2/HMsuBvV76OWxYa7rahQJRVnsf6waZ5mWXpUnqledT8MDfJ
yYVTeof47eu4zzuHVHJ2CNvOtEIBG3Zmm7cmjJFLv9OrRqN1Aj8buN+ffTLB4yS0
0AapUr1P+CBkI0RCf293ArMMAuCj0rJhE6vlJXuE0NayBrEIbzTdkNYNdYNDPPMN
8+KcTNQkLpWz41A2fWXG4oPjj+9dYY8PfrUOgWUTWa9McdV3vp27bnY/eYzTZvEX
/KHiey37E5g3f/bOfayi4Q4/HevsvZj0LRm11kZzutTXAO0KPyCueozo7SICaJ6G
mau+r66ZMjoxj776DNG72LvbDCaBKUctHiR1lu/o/ZUxvlw0tS+8AZHGXL71MtG8
/MgEHR2JHZxsjXwAaxQBfGXPODrQfbtTwoLXLXZ9ScAOfPngguyIEPj6zBblMsq9
n64YTinzVqA8vnNq+eADSNMNKcIAOrS05ioSawrdCZaHfNV3iEUZUnafPbtwfhSn
t3Nt7gnfJ3RQQqSOFmac1thyghek/nXAWdEofMCoV3GGZm5AFkW0MtM7lfvNYWmU
+BnOdwvtS+Al5eJ/2bG/KKqNG63/Tr2Y1PVX8EH5u3Q+2fz5KKX21K4T6+2RzPao
ph615GkIH13FuhnJjte/jRyeDWrjTmBq18k3UcKyV+dd+TbOW+7oudMe67MO/GTd
M35plvyzY+zaOvtbD6tyqU7iPbP/NRn01PAW4HROJidn8cDEmxHyd3M8Q/QYr72b
qSkXhJL+KjcoXoiJGHqEBw9B6M/oU23FHXEMN0ETkFzl0jETDPe+FbK2LWFIJkW6
odUvXdlXWDb8cgdPI9+rqDt1FHCpD9y1NiWyE2Al+zwFtws5zfwE+srLVre6xHbH
A2MNmrb2W2nvDDFuW7Yv6RZs0QJlw/FAE+Ko/GkZMwUe3Sbt5ZNCGWLQtG1NRZt1
o/i1d7eRBsSi9RFW3dSid4LEjH+Mi8CIgvhpz7HNuFqL273y+yPAPKeNw8WRq3Qv
6FXV02uH+VNBUyyRNc6uItppvHoT4cFexlFTgolUXz4g+cGH612I4fYBuhNkSrtV
fAyut6Gn9EM/87CrlBtzvKka6/4jmLArG0WYao9OB3rscNW9cmNxEjWM3WA23OdW
trVVNsLSvR2F4D6yMxaUFdJlhzKUyFyMOI7ZHPtKE+excrM1EZ5LLjubGZbTK1gR
F+EkoUXZQpaAxGbE+4pjSZsYuEp6bg5DgKETJ/wbZCEAqZu4RUlo/ZDWA3vSXgZu
v/tRLLmkosF79gKWirWFgqrsYT+vnrPLdF2vs3FWKguyA/joeQwUK7PVGCCPi9y6
SBW69iteCHxKotIH2+Qd5wQ0jA1o0IEsgLiEcPttCSqeMCrxKLh3YL0p/GhadH8b
b15jZfvGi1H0Lxzprg7/E6NrLYooSFkin/U6drOFomU6DIn+uCpne2Ia29RDMoXv
/IJwucyVZcKTjscOjgxUeY96IjIhEjHevG6xItGXuev5UJt99O06AEdPbCPkKQ1K
JbtpNHCoVWw2LUxP24wv5rlJ/WdRFjSRSWL9u67QHBGaZI56TNswVTfLvUzL0Op5
zvc+PM9QhuqE68kUPQ3222hy6kCTwz6xWOSkQujWSu7V1kOvTZepVuFOv1fq4JKw
qxJ8CCzmis4AcpCrpcjgPINbTdbbdDFiUATcIQ7Ax8oYEjku20bxiPh3azPuDJ9n
M1YFydoCQ3LFwXdlUVJLUPPlLtobVWrX/0l+RCGR3HcgleAN9e5iDv7h7N7qkGna
EdBHiBxvbnSpAPi6GJXGjFxr+frMurW9ffWOTCf6Mpw2ttwQwOdSCxc3XvHsfmm1
Z4f1BrYn5NSn5BFId/V8YxFUUzmnMybnd//kxfw3b2C1sEgT0TslUnBdx32nVG1c
jKQpGwxEbYs4c/RZ7xD+S/+KRy8pPDCsoKiz0XEzl7LophdGeuOMVRWwngNjyoCu
ogckeKexz1MdrH7FXOi1cIHsSJBgK8+83lEIS9lxzVivZ1KnTEOU8AL1Js7izBWU
WGfObmKXRj2MXcLhwDgFypDe0mvevXtzGTYD+a3N65/WmT3L8pqPv991qVFECSMW
zy8sEm/k0c3Inh1pKRC7pzDTtGWjV1eN5XR/pgAHe1a+pvC2wUjpeyYknuVq7kgd
iLJA5M6hLOr05TYrAcHZXpvzTsZJI4f+VjeJjUphdjGeS5bBiLj8Lauloumi9x7c
O1P4+u21O2tnR5OKgL0VoUeyFPY0uQUo0kzIPaOavy4T+pGRRNI001aVVPucKrpJ
gxAgt4JN59E7bMYxhwKj2wWSkKZbWHBaxwv64eyS2utKjEnJtHVuBEjOdL5vU5CR
5EudYZhNJ02vH02XK7E80KJu2NLgikntyUHLTYyOQifXBRmRoSz2hPfiqsB3WVgC
CbDTZ0lro6PMTJ3OJYmN16WX+jJZxug1QHhPhNRGnulSUHsbhKEHqTMn4EyM6X2J
KxKJoylK/Y8cJnNNT9jB6IAyXhaoIB6SnqXMl8hHtoKMWwF9Aik9mki4HIEbP3ON
d0D5FQJhHbSTJB/IDoxxOkD8zHLUX2Db3Uhf13pyAgVdqUfDghUb3n8/8kAFFVoj
NUiXJpsNQsYzZgLEaZmwCD3+kOMQolteE2kuYLoWt5uvq3t1m1S1NnpBWESzQn0G
oKRMWttlgyGlOo8p02oYsNqb9ggWNjY4n7VhrzGsRPysXztSJ77/ldkLfTFwOOB9
T6SlCw6FyxMsutuskt2Yf3ZGS9+f78qcgaLHRr/fsr4Vz5iGnqc3FimFmCSEeAg8
t2E6UVnEL4nyZK+YLK88BhLQkZDsj/43lsV4cQiOAeZZBh19uumenugSU/bGxyQ4
wsqSPGIYr3HN1oQ5zihbF/4la0Z93M2nFMD4YK2qZmq/NahFNW8GiECUorHQOgRV
UXUlhCWVPTi4jJ/4mEM9PXsPpADNqkkQipQ83tlmCElNjRiF/1PL87dgYgyGYSau
jcEN+VFUv/Gc8Kr/B79NZrrDZOTjLbbXrIEowr0oMjqK9J0gVEM9VhgCUa+bvnDC
oBtvahGsf6VvNXwqnAPe6A3sd/E6Wx+F2QylsTH/EhJ62QD1swsxcJe+the1pt4n
vc0hz0Sh52shVPX4salOv5oTWUB7Uq6MXc35ipCbSjQ6sVbKCWxmg9OvsjNY8LVj
v+iKSf3IC4rYFBxdySsWYKO5afknsy/HI/njP6J8OFrrRniaRaW1fbOj79HsW9oO
MkupKpXQU+bQEjtYrJtnW2RU4AbQuYjHoALRFfHMKo6sEgxFVjOcjcGkXYcYt89Z
a8+gk9B2Ghs90APvy1JecNsfbpW5kIKHjEwGLVdMVyFH7M5TvODpvtRvvYwErTZZ
CO6FcCJExggvrz7Fh61Vau9tXRJYKoJuxHpqpnzKvwbHp90GuwTRF40O9j1M4BaJ
/+WgqjPK0g4GEnr+uyyWVCt9tyb0Oc7bRr5UFHzOZzkZ+fonmLyeFAdxYOQ+DECW
DMWXnCD0AP4OJLivD5fOHrbN5kYw2R0BIyVWifOGHAm4ykmatwsUJOXgiwvC7GDF
my7G8Zw1XnYFE4chxovYx860d9l7bsxotj0z91Zl36uWhIxezEd7vDmHJ24OQNrx
rvy+wg7Dj/puRJvb7R6ppBV8pKdQOo/LsAXgtpcCuSg7Pyfm3cSF7ui8rXBx1VUc
fOfb99/9/WPVoc029q1PU/Jghm/K3ROTPN3p5HoVTE88+DCd2Wiid8suVK+a0uZS
qhtkfCmG6AsioNBocaB1sQOBnz152TzjJTuz5RUjgLVS8rS0dXwrEuY/DJhBzj4n
m7qOKnIXLOhx2YbFtTYkQ6LmJ6/4LwTKSREZJZW1+HVStyUYVBZ4eVXPJ6aJfX+i
HZ9V+QZb3o63+UmQDGWsi1oftuYWPBzWfL8HdUoEX4/puoxendah+tVCdWgvzLA5
8NA3nRQIbvpQEMiw/u8wMGAv0/XLwxEXVJvnM7Rd5QAjsh1StJhdDRurcdhDbnt/
/6TmEMrVSpXt6SvGOuC2orw8hrR4KKto0LRl8JsQx8/jzDj9EFr8a1rl4WvMQJgG
GksTooxnHw+qq8OVeKsDSZsqJlUFd9T43pbDGjF/08dRO5m762wQkI+OfbLX/C9V
1cR5t28dzDZGbhKe22fP+Ch7uAt824NwgV2kXDVf6LHWQCfr3y3Mjnki4i6VVJHD
kmvn6Ax0kDtj+k4j3uDuJdE/ZDnAI/4iaYC+LErUTLu0jPNmIvv0gk6NTiYxBjfh
2ZZnsLNTBcv7uwLKReDsJHgyWc8de639zXHIEdMLb/Rua9VZ4MIJwtkDFUkPELBc
QAjT2r5on6aUqQ9zIe/XnKiAJInSRSN3mSIl+pP0ay4rRtHvTVjyXLeLiSSBU4a8
46kfEz28a1VGfICUi8AkKDspXFKcGV5JTYUTmUwbwYAfk0b23fux6p2ZfUhhr/O7
BTuAvmW4CG1CVunKQ7DYiqjHgvXpngCqMdF4vtUBveB5olnxu7e/AngCuZXv3Frw
9sBRUkkfu83ClBAfnLJXf0R5ZgywtapUjs7nto9j/fMMI7bkOr9HeViFHEMr7Xiv
1e+TfOmzA9xvNAIOvXCAjl+h8R5bdxcAwhD9cNXVyh6q+SEgJdhkSwW4Ml3BuTON
rab/6KaN6cidXDhAG00nTXwOotutmbckk6fp8pQdxYNyDL7AAqHBV3hnuqO95h0P
fuejY8qtKY0fkOX9FFWufEKTgP6O34S7ea02urlvJTG6qzLNNAS0svz1DVCHdZiQ
cruwlXxWYgFZgALOypM8sM+LKm8rdN5VqHni9TfyW1QcmbPQxhXANlcpN9WT8N6H
feLyGra2viYmiIuorvh/AZu6k8wG+hqCNwpvtwjS+lWs/ua+Y7HUYCjPMNTQ7vAn
IEf5i9/7UwPfx9mg8uFD5xmDgvTkUMn8x99Wi9C2dZ8wjC9lK+oox2Rp6bujnga7
vHfopMH4HTFmAoAIug3YpF2i0QZkMf4suNpZXmCcWSCK+V4FLDZJDn6By7YWhq9O
ho2qSpqwXQBllWkMBDH4XX1r9ZdvG6mOCukQnjwctDP5MjtRIGknQ4jW72mX8ryX
UdE9PNWWa0hPp8ZQza7s8RUdQ79D6zMPfcvH711ClYoqtjJLdfgLKdD3EAgsBLos
q9UoaKsQY7v4b3GtNaRsl4+02GR+nu2XrDeyXXRZxSWlxV4eW8qQqd0xOHPKJ89I
vuX0OUJdFudq6l1604VY48lhxOWiPUdDsrhnZAx/uicOOSkftPma6oSFyKFB0fEg
1QCWGYoBRJZG+AHJWgOiE8YytE8cuW++eK76rH1Ab79wIcfD4Y+JRLHSwogpUV5Y
IMYPpVF5bOfsD5jO2ggGxkC29h0/xvzouDyao47wmml+DtwRKdY9rXgnhBHC7Ac2
a7goZHMN6MLGC8M1xoWBOg872mDBa7Xc4R+SmmI7/UVdWWDJ5Ejrw4XWrjsaap8R
AWzJCy1bjaUUtl7KEYkFprrQhbCont57p7ShNnZcFqibqDU7pzAhW0XbK+8Z9nhd
BPP9wIyIzj1alh4+gUsJEz5j2GLoFVpEnzGIDjwoPIyo42nSAv15t3OqKeBGR4CY
7GMo8XMTLiXdb/Lu5NM/IyOvk4UMfUWHf9h9hPH3bYarZR1oytIiR2v6iCZCtpsC
W41+2TE9ClLdRL7gggIK5rUy6gIUcdsqyOJVSOl76dOsAxa03Nt+PVcgg5HldnS9
KPxRBrg38b0UEMYubJIhbH5xlDOP47PvwRLRhIW1qRTrZUCVloHGGZoPwx8CJpAC
6FJ15PU0ZTEJ9me85zL1k4wSquAj8pDbssOFxtJGDa3HlEotdn1ZxzX/INqRUyi5
RQkXhGrzeVW0sFViqN7giMmg4BrdaCSnPqvQJG+AxQpe3nHeAUkojYb3SsyU+BWs
QeQ+s73u2hHnOjEl9R9voTMZKS8Euobxf7SbVgXMT39lbk7Io7HaffKJ6qlyPLrr
AdlXi8qX4dTW4PyQW480aXPeVZgH9lC3ibayWR2GrGFx6WQsXO23lQIWe5Ql8l9j
WpR15J1yEt6aedOa6Divpzn7gq7e6UPTg5CwvoGZFCPjItSbr+tKdeRvoGsEOSDc
Ru9kVFlPvrD5WHTfSJFuoQnq0Tnn0Nt4ROa3uVelm97f4z0PcSYhQBrhStCRhAOw
jYxKs8d3qF4mCVfKUpeby2C1JVlVv2tuA4Y/1fXf6vvDjVne/ZhVkcmO3Pooelsz
9FuNPWDarxzukqTq7nBjUSpDymLQBEqEA2BpCLwUC8SEw7NtYafGNwyskpL7Tca8
b3ESoTuLnoL+nYf6sQ2ZEnMXrAyehwr8+2Vy0UuSjQxgOix+bG68YjzmWsPq6U8l
++UW3kgWpE2g50HU3irUzkP4zMb5+1s+DHjKYxFC9NFu1/8Pa25BKlu3/Nnff39R
FNZ1+RwKv8oMBu/+NgB9yk8WjGIBraKlUi34UbY2VtsiWecs9PP6pcPUrJ4LU624
zkLK5CL/3izlIzBEk4aAohKn5pGe9QV0Tt31RStP/Cgw7b74gG7VNZa86p4a9mnA
84RK6d2yB077N4vhG3bChjlhRAVMrm9LFMalEtT/AdqQSmBd8+M+O2sbUwwUi85U
tWEBvW68A7y0vVLN/z7YRsP1EKWZ78yK7L63pm9xZzHOqMQhwI87uhERS8mpXZXm
6MfDH8lbKHlrlcchPt+bklb/r+fTNw9lPvTZqS+nrL4WDUBiu6szR7kxcFzveYQR
miFQUW8FIFGhbE3hJ/dKfxdL7i7gfLgpZ3Z6jAq8adOuQAS/bbhHMelsnhUAJDRW
w7XZhVsuuRYzD1Lj5gM0Cztgu+FLewEZSgeQxzi1MSnhdIzxT/YrEchBeqoqEMXM
dHzX+WZTRm2g//s7z5SCL0nUescbphK7kzl2N5yfv8U98oWd/vG8ETGndDvqi1fI
Ryq1kpW8fO5eBfKtyHuanSkjgez+I8avcSQPtQJflDYcF/bTJ9X5oK6icRYy8e3g
/cgDPx8Np6V7C30Hsd202lV6HXov7GDe6Iqs6G9W0MmfVOg3bYtT9Dhdg4ZU7eci
SXAVsVL8n3CrZwabi50k5AMxBwZktNE8nm0DfsxQKRpWEJkRsZHNOa0ZBnSDBF+W
TicP8c2JASIaSb0NXR0lQtj5Nqn18bwpRzcMfvJ4VXhBVseuAee9JJ0dsNJjg0Rj
2yHoq9qOxzEBNFnILb1g1YbPWKUc0tfJibKGASLCsY3e5Xu7G32lUiJYfsJRCbpq
2j84sz+BzFSKlPvXV0XPY848DQCH+nQdcyKUk6wzThAZfUfhjyZibShLDvRYn12+
2rvOrOQ0GtXf6k5S7Ad1ctqugPzaYS3mj42NSAL1LCE1TCy7+7f5CPacDOl9pU2n
d5w1f9whkV9WOzrJ+eyjF74sli4T/FUak5kxGNI6VcKhns1STuta5GXSl0Hul2vC
f5FopzrRGFWUGO7Xd9x/43+rQEGpqiv4pS5TVh0zAiAi+3IpTeji2hfebQRx3piW
xCjVq1xCHq5df0R+DvY1TtALUEqudFYSgX+q8Vx+6wHM8XzCqBr50CUm++NIOoBn
R7bwxs7sfLyPdJ9FjhZQKfh1sMjvLp/7Z0k5nyujBronnMUBg8O0XorcNV9PJQf4
kUPIvMbsIxbuZAjxRHg2HGClqdg34D5Pqe6pNh7BHmppiLQwwR3pAzNf4l0c+QP/
UTRaTm+/l4V+TYJ3oILm58NeYFwrCd6mspbTh3JhwHaikMIDHh9r/OlPXAmW+Mct
9XteyQbf08ntSi/Fr0DRbD54g9nWpBG2uS0pjrZELMh8ByqxGaeo0HF7V+3tzekg
iynlZ2WjD3mlKh1E0Ui/55eo536XlKOb9wZUNW/hRFSP5RVZIO8x+znCYjELMqm0
8FRYf5xySXD0FjaHos8PpH8yY6qX50SOU++eKgplPsgOfyrjFjhrGeBNfodo91fo
F04IqGkSIy9RX6JhLbSmwFJg7x07gyLsaio0BlQjTjXMNEsxvHIovygJvFVthQjK
w4/treI6cSWeQPg6KDxjpkDYbV0Y2O5sRS8Q44CmaJk+V6EWEBfIxR8mJRlmBaKT
u6KXHaSElWHGZqpn8N4BRUVWhqOhjTHK4FCiqp1mIFA1H0i9ofP3e9D5fQfaMIxF
gMyUxrTQRa7RUA3DILyPdSoAr8mhPlzALAH2hRGOsgWQWgPiB0Nn2TljSbxijWaD
wveTuF6eJGhVqA9wOdFoIS47qL/nJDiXGjzLx2wIBh9oi+2HnDFCsO6KabQgC4oc
oFNizOetWka3UBE4BAZiMNUFA9xYukjz69WVLgdX9DBiHA06c3kLuiIt7OHlLG5d
GvsflyHwT+WK4GisxGY8ZO1EoOeSuJtKyng+a2UiWLEe6b/oRqqFqov5lFLIVr6u
6zOhMq4sxxhiHohZF9RMBOOX8mBMo+J/DFhtpBZsG/bgni2QuVW549ac3CI2w50h
KrpkJaPYPwDOVZkcQsjE9fqMB//DTKTnRCKA2g7+fQ8BuE8M+OAHcRDlPuzvAuC5
vQvmqAqT3pF32uFdfur6B63IBd47OptCcWVmCLmHgVzV3Pu1naLOTKVCyejZ4Qle
1wmHtGqNQqke78l0mNqPJeKBWkUMEwzbW7kHLfjT8D+CHw9QtZOz1IMgdpUsJcEL
dNs02rkUIFnVoZyweQSrQUbIaTovXoYliQMOj2QXGh/7v7TAhRnuP00YONMOQcMw
A68pKxYq6h68wxnv/QsLwdcvkFkkcmy/Z94AxFZJ26TH3RBt/4JjPk06Eq7FzoiO
ms9hxTo4avoCYSwvIpTTG1e4P9/w37K1pxG8tkWmBAX6mryrhsp2ZvQ3+MeyL/J4
ZuEyzHhZw17X6MD7MiIr9q7M+BZx5Ur6Q0jV8AaMo+o7gKPEYSfdJ2xZr2wePncQ
NGD2PPh0SiyiMEsoRJnkxYK7ztdzanbY0cqDomo+Moxk8pvrozwJID6xRwQwU9VB
EoBa90DE4a+/0WGhxCz/ulRTFIVqL6UV+5jpIvrIj2bAyQb+9vL6LNMwvGXb1RH8
6fZEdo+cX8Oz4aNa1O/g96E2Wezzw8ypLxIKJALqZbWb9Or1ujZBbWqnmAlZ3k3s
3KgZvQPaxkAnURrA5plBjOBOkjPiutMGqbgpSY16em19in9dhJiv9WTR4ZEw3Aw3
s2pvwAVsMa0LowLGnCTyxEhGF7DBWkmtFp6cTkSI+5dIJdjjmeFInl+cPGNLuTrP
3EnfnqzXbS6z5nP1lgOWzzjvQ65zmFqBZRSo28W/syRkNsibDniHTgkPPSIe3GDM
jK0KX9rXkUedRKapKjzzJhbOFzirRBe/cJOtX8oBQwAyoNTCmuGyPseM2PaEJLev
HEjmp0Uug/7v+/0/z5HwbNFLSbFcC7GRdHVm3rSdA9l9r+XO12S7vyuw0asFz9nJ
2SmZobFXf0t48j8Nz1NEOU5umAZ9PvIBCVQXX5g6kCUpF6f/UWFvUOLDYkfB0pXt
l19vEQhiPTV2Jr1dzF4w2FcZvD/UpjYIS+SdT+rQdjrhsnUw9tnfL/g4u3A6CJ+y
fOq8FMw5fMFq7RgWQKX9PGUWgfkrQTdm4f6yFUXWTEHK/XsdLmCKjmNIYKzLqOJB
kjmas8JbBtFNQy0HO4l7oJR6e3k8dNzyFNbOsCClStX7zcARABMcdaOaKsmRNuqV
aj5mFeDTksLqZNX2StFKWO6EBQID1lRhWbvZ5LARqn+Cj9eW3V1L0ft2oVcj2K+d
FUfyPwxO7YpwAUYwWL/KJQu9cjHb0x85FhabRypjF/8deq3J2zQQ4fjlWqFBKU6d
9SzmT7lvD/tqByT3Y8IjxhLH8zhcMBzSrFG0lmbT5If+6B0AvsNvD22k1JYypK9m
gGUR+Jnaw1P9e2LgccrxhcfTt+MfEbDT8xcm++RGddLy3PLY5Hyps1Oo+JaUm3dL
953RNwayG0hRJG64PVyBxF6rqk9SQFdTlvMQYmDg3VtidklsE59LHvY5N4DiUxUJ
DtltUfyLyn3bpDW46RABnXJRyzDhAgtEWrt3MKVFCwJxSMIjbg9zjTJpWjNwOmH/
F9qv39bxDzMGZENp3aD8hgnvSEIkFjLexrhJzWsB7NcLGSe0qBa4r/9LW6t59f6r
lv8FzXQyrv5wqhUijZqz6VFv1NYwbq1axWDHjJQpT6dY5f5Cu8RUTvbWG69BXXif
qJcbIH+Ve539bBfP103AlbkVKsIxuP1Lv+ukTs9mFcMDWTy0SnHzHAB/XnO0RL6N
oTpkvnyGlT6POUaU/n4KYLWFagBRfVUOfTpdZuNhYQ+MLf/eUqiMmRc7tkEXqKp2
xdKHUdQndjgVA6ZkWvDXkUb9cmiElSX3RDpjTQRbgWs3BB3JB19n+zpXOUSeDda9
kKBRrshvx5DQcrjPp98BM6TxgGOetVsXj9dvbY5A+ezeomSfkKd0mZgjoCGS2Wym
CeZdHeJCnSVzwlvrB4hVfa+neXFyG68brVtRhjCeN48MrRCN+leP8+sRcFnVZrmh
R1wB+VkUxh7n4LXWldgNYrk4UOcPLgnpS3Zxkx+OmZaii63Hf0dq6f9j6+2SRO3K
+Z/luqKzh3WxKIBlkmw1oPmNpPZ4aPbnjVez5bM42u3zgMO4oBk2rthuJdY0NXHN
/qXVutk5JcjS94qsONBM1F3epjR8yVo/E1EUJEgtWCYF4sb7VdIURGVFat8ZNnqZ
LVRqmj5XA8C5AYhcfJn99/DtFcNUxI9tffwCadku9VkKgNZL+8Liu4AWlsWXKwOa
uWEVKRt3OtiCTFKRSEbsE6ImYBe4zfMSFPIvDaYxyzw6PoCwWkjegGPG53oErvsg
gjcC9BHnlVVQ9SraD3d6dEAcRJKIXcaUPi0l+THpy71Yqh2Ys+PJ+M3Vwb3lBzYr
L1BX4a6yxiieJrps5Fkj42LOwBhKt+LkWxsp3bDUdIdC2TdfXj37uVCaIC3d0/w7
CY5W8+Mp+Ogu9zCRBBOPUAMfSQEC71/akmT8ZqvPOD/VNXZtdvwhn/1BOb41JNko
VPH8UJamjJLwKh+a4uJzbhdvj4zpAwG1GVhZ97xrH34cxA3DU0pUWqox9SxkfOq7
9kGdwJUUfldPEk5N0wyGqJMoY3Iqcemve2bWvp4qR+1amZmxC739Hq2jtjxgh5tf
qBFNf1I1ybd+1aEZNani0sgQjYBOiTE63MWPrbmSwILvYRk7XY+JM6p2Ol+V8Cug
KiIg0U/wU2x/Tt5j0ccJGY37NXqmVoco7vYaipH0liqslppORMQoe7+p92VZ60yu
zmyzsmiVBvYsj5U41m8CEZ2ba4TEvQuhiF8qPHRJl/5EEY4RqxadUR2MshH5tXFn
qdCWY7JTuadvjdYnR0Ra03SVDh2jDLgfjHdb7MRYzeBtEmXk4T+ngjHFRCKeh7BM
QcdDgfraBFgyhPNijHepFpVnrQ+nzfWuZgPLhM1/Jho/ghKMaZXjVqNnt3dbviXF
/X4kaB24m7l99/PM1ZaAvJ8yTrpevPbV8Q+5BMWZDzfsW9BHcn1RRQ5dcQvf7YSX
wma8u/7KBUH79PGUoiNJAYW8Gn5EfcoNsND3ioIpgMcuxeYikGEvviYA0oNL0k2X
n5sAcr7vJg3OcUQoOG5ZLFtMeI/jDl2RFe5U/7CSdjaY/rH3HArN2Tz+gqhTkKdU
BdzFtbqb5A7YrlSIQsBsnzE5QAUequqBoQyumSKK4N6+vd/aD6uf3HCvnp1n9njo
4lK8g09o4v+kUEXwkB1jmwkeVCxaEtzdJEMfj7IsH+RkBJtCKVs3yvkzg2Ju89jU
wRdUM9GF8IKoBhJvcLOgC9u5wFrJX+rkAQmr7BbW8KXMBaO5hOtoqPY2EuNAm+D/
gLCJrc/9EMYvd1lk5ihXiAZswTxlBP68PDZz8wzLPpGlavRi4c4QUQ0Igs6OE/oo
tCKSk3YdUcv3rqUa7HAvnoVomIdvH3DaPMJe6O3SLufgA3n29I80u0V8wuk87ZtX
dxfT0vpyLxKqE+uNKslGjnp7QIkU0PaEAqA1HbCcqlGKera/bfkJcpB8BGOZFBI9
zWu4uXGE6j+fey3r+lOI7Qt3Zoez3BhQeqsITotluvuzMopV9UEMBBpYI2o1OWrt
8RwQ+v5sSpxrz4XP3hwMXAMQUoObmtS3b/zFHVfZ+9NdHySgWOFh/MIL9T6+qgPz
JBM4E4095CEKDr9S76uhTlE+4DPXj97FeVt9xNzvkHAj+kFpNEJu/296bF1kVCQy
HN77qYfgVZUXK0uXn15ZX6TTZuGCvd/ljCj2Xe9CApSg1nJjqOOSYMhBF13x9vJf
6T1c/Iq3e771uW6PmFCTwI3ThZp7REiXntqUIHx5Q/A6LHtoBY12SFzMLAwRHgol
FYQvA/O0yoArtF4bsxfsNW8bjyo4FQhgYW+1c9oKNgSVTOB4E9rAxLO4nHqnYC3e
fHqQFpc32gzAp0XVPk1DJ+ljnH9zrPnNh61c/1fCIt2Re5QCxrryk96n+hXxsCfG
r0ysBr/nQsx0X3FUezBSoMmg5pMD2RA3AAFtb+JauJaf5fYXniFGm5z4hvPhTJEE
rpOoD+ihtGiyfFqgIS+a0DMRFzA7JhJqm1wWPUmp2M8rEFONt+x9HWgfrDeIDpGw
M+bvMkIUAMO9NHoGaGiGaq6KTuEh1lloSdmhpbnxd6nl7v6MujVbFrlq/9YFQq/c
EVrQj15aPBAHIxX3S2I0b7YVQ727N3Ad+cl1WbuMszgtEDzYepi+eM1/91PcF+ta
FgHveIkH4DM4mBXeJvpxlJ6+oMkHhSQNQ/4ohj8bmlzffZ4eLeRSZlpXjeoxopfx
LR+enRay6YrWqPCRkh6d8YQgUqsgSAIc8PR/mDLLd0VA0/5QZFyZa/t6FsACi0sS
kNm4Z7Zt9tB390AoTktjcDnVrGbPo8vNn8VPJH8F4IATqYkb46yIzTtsqNtVaQnQ
aZkmxlNwe5+IjXBxG6OUBgNqpIbi1+yooM/a9KrQykb1kTXIH4JwBHxQzg17zsni
7RJORn54Tuw67smhzqWSDsPQUqrlnKaBK6vh4XrDahBQ2kWSCeKL6YE8IFlHxgM1
akbphgjCaW3GxVBHHCtB5QMmOsRH0vCGub274FdjvptmIZVLmDQwBWq3mQQAbhDT
6yrn0fq8iFsQa7GuPWBpeGKzuaimTGAfomOj+71ypjt72+xnfJYw0dDP0K+yqvZ2
7ba1VeBVoUlRkDP/mJBbeMJnKxMA31GySxJD0UA3EwBvxwm5vjiytQ3AyDl3uVSJ
Aqg0d2i2DIOqzPwhmf/p5WtV1a++CmcsLjyzdup6uvjV97V85g8kn8hg2/S5VW5V
6oixlGXGsS/yzS23GeO2AVGjsn44IoCsc4mQKnWwb6XIGTRMKeOBHYfIeMDPFm3d
Y7XWuAKs+QD2c8u3FnlEUiaZc5IdFfS7rLsuSEROU9LGxSu/yK+lmuQFM5d8eRaa
U9dyqSbhSYxAngxaAQ0OyO4uu/aT9iqUoNARdLwtCDGPevF+w6pJq/5apxCAGkHa
vhSy8tLsxnR2qNz44LrNiC5I9KzCncTC3w4oVtn91OCJppO/hLg3Z2GCCfUauqPw
F9OzFzfUgBgP3/NOU0hiWLESrFAp2mqAG0CXPh+ZZmIK4XHQo6E2tEjlG2VkPTtC
pX3yspgM+5L03/Z3xgjJ9gN3B1G0tZSZmT9UsC78VhbPg8dcXRJpCxlUdVB5X5L+
frHGyZghHR/UkazNu/jFh7Svlxq3yYi8t6h3Db/T0o3p6ALaM5ccxfKHk8q7jVLA
lbKe+uX+IPZQEyvkpTZu8cLS7xHUXqJ6iymUHrXWdEaP5qyCJru8gB3Xm1/Dmu5x
Zk+yYmGtFz7hdVE/fF4/xH3L9KO5rmEqK6t2IKKe7PrP5oGmS16qnJHpVQDjMZhN
BNfS3CYS/2l68hxhn+WLT231rdGaBBkFkdAVUFoiloJCO9qzxQqRqUDxsmtiee85
FDJkmm8deQCz+FWCsYQu8GM9i4owx+b6kGcZu+jndaLJgMyTWixCCN4VCLADSL3j
uTSeWoHmWxFxfqS5EWwxfmI2fXFvORft8ql2ynpWdxRdNDzUUaKwFmGcxg3i3QCZ
SY7oVY95Tda38iXBSleNrZKZDQcKJaa5zMgOzd8Ur7YbUyRVHKx1THspAdOxJHMY
Bt3l6NMvWY242yc4N39+EI+yOT3OO1hlLDMhUYaSpIQsuV8M31Q1z3mPv/CrZDXZ
qied+kuTj5MLhab8bWalKZQ9RMEuaGDEkbFb8/sJW0elx7MYhutGDh1rPUBWg/nb
XLzAzarvqnDeh8oV8x5DvmijobhaaQ6xrHsPYKhUXHWjboF6Ft0epEd7fM9JCnWo
9ueUwLVqaR2ER4ykZ6OwbzJeBj25L4kR87pqlJP7zjnLFUJfllX1wJqj2pouHUFD
DPxWZx2+c88lM2oBdLzbZSKCDX0fMN+76tG9CI4jWlAd44KHjr/TZc4yW1Y7lGOJ
myIEUg5UAXYBBlB8JybauEO3GI5Yyulmg7o9VbfSLFb0Z9As1mzUCQhltzIwI9sn
8makLb6+8/KUH8xryRyBQt22z66pPePPpK9m1+Vb0BYbPeZ/zaWhYeuhoJhdDyS1
6erOVq3KZUM5AwaJ5nBPDD9aWz+13n7tlciX4N5X6OMCOIjWF9wzidQYMhKTwY5Q
Egxv8eaMkZLisdt453Dp2GmS6ZiaRIpkxMkbJrmdWJKAKxu+loDa0KZ4lNYmVt6u
py48Clt3vmLiyfOVfImdMy9sQh9AK/Iy29dcg3sd9yLoucsShqr8BzJSrrlkwL42
bNaXacWWk2utRMdEVXLKJu5Z1A4dmW6m+B0UagDGjZUvuPDYpz/GlEbc6z66YPXh
PVIap/iuF4PSj1RAXoZtFE7ZLri3C1MrEm/wQwfw0PXBkO2MIPgAAybU7jY7X/Ow
pGfineYkGa/c8tUSfwudm/41+IXMVmbZDH2CnM4z+/R9sMVuOPsL0N6R+xoTmqLJ
n5Vuv6H/H/kkrwIw5RXWUXs8OgvU5rRpSqApN/4GqUUxvkTtYRpuEsZBHAVV7DWe
lWIlhbYAbDrOGozsgCo+FfRaKYCWwTI9lphDCHU0809CsrCN+OJStODM9o5lwJ7n
0Hhm3yCq5wrEJ++EeY1frGRvBuiI4aP401YjJC6KCv3MSLks7czUcGTJGi0OVZ++
3vVz9T43vg/rWhI7HFGtUPh+mJAf6Yz6F0utTelMNubkvbzrLaEBxaF0Cp8W3as8
MJGOUvFIqjoxw533GQ94yeq8rbn58UTNlAnx8xYApmsPZ5eOnlLbA1Cw0ErNSAiW
DB3Nos0cmf/r4PMx5nWnUl5NDs6R9IwHT7XTIqOlOcLPaZ0ZHWcgdIXAnd2EamdN
1H88qxRxoW+iABMd4gGbLVb5BnW7Xtg0MRs7XWU+u1Nlrkje/gFnKgZWwuza51EX
2H4fM+yyPJwqlnl/7LKeAl2qzRvLxCU5fWlxwHD7qQmJHb5xC91uNlUiHb7BEsp5
VAYvR5s2oCHPYdMzefCpZEF4i4V8GToSI1VYW1Q28im5MrnLX+FnLkVGPV3ZS06K
lzYV7sWGmQv8/t0+akYn3lvPRv2sX6a61UHAJg5hMolrBACRiQUoGNZYQBRFWc22
HCeU6YLSLvTSzkrpBJaYBq4t99t+MA2plAv4vW3Lu7YSDKbx+/uTE3zIOigvJWfa
HJ3AKcZsu3q8j+gvV2UFfYB2TRsZwU3+BujxfTLKiXTjc94QNd4Xu7Chuoy3/a6W
my4m6aayBatb06/ZxD0TQSg7cZm5mg+Hkdvcq7SjboM93SG79E6SI6UlJ4WpWka2
cJNXVXXJ0ZtQiuC7yyniyaoUHo3nPHG169vUuGnsAtSYg4wwS+v9FNnEnYcZUJ8d
AsuSWbKHa9mFmUBSGb76kZTDCNNFzLtHqle+C/D2DCwd5DoreFowCuqGiQ/Kot5r
m5Dg5pE4pSFjPIdvIVipE1Snm+0qI52RvHoThgCdg8/koc54lhebU+CxBfxWL90v
a5KumCh2mWgnMKdnJlQQ7/bS/8dRCAmcKebtiuAEZg4sPzu2UA/XdaSqBe/hW/1t
s4qQ85gQUD6tCGrqfun+tdDgM8T1jbI+qfEHrWhnzjJqXbNc4l5lZQJC+AdvN/lp
u/SjfWYsNiwY1PbGGGt7wSJU2OkfGaUowOZ/a9MsfVHI1cm5WX8KZNIh3oFGOTcO
mcyBIjUAneslmZhkw4k04Fq0mGKr2Wxl0xNUN1SERH2qked+MU+9mskJZPPHHlFW
qPQz+ZoMjA8AOxfY4zFKh6sOZ2ykKKCfr4e3d6V6Ix3r3BZpd+tte6J5DzuYFeUa
4Adv4MGSFjS5Wn2AgwnG48K29ZxbeQyHPYy6z9z5BA6cdbWL+c58rZfRnsnXyA6f
KuJZKK+RgyUiAcFm5HiGxAihesti2h/1bVOBjO5TeMoKSVFBnO3SxnL8zCY4CDtf
HfM8hHC1CYcV66bNesQ0uarUyy9fU3ZISuk13075w8MbXEk+Msm8TqZtkCIfJEdp
RL7BjvTpA6recfWFJeSnuP+V16fYlJKV/dA9TyXhVy/FhohSeFbeRlfbmXT1BgFo
VJKKpLb2+ahlB7abw2oNeWv+nGngv/LphezlF7r1rbCXtCTsaJ7AHbn6G/uCaKv/
XCriYEl4pDqkUG6rUyL+BG/ZIA5qM3iZMmtrcSNFyLbdrltaShRjVjG+6Ihcxs0p
Zhiftg8iKsF6T/TuaIWvCmsC+OqhhdkaondIqkLt5xhXbgiRxUHxTC05Du42f4ND
Mm/19RJVNlkrnbIhlyZhWw2E1x1xPSiBsXLfW+9dT08NrpCkhXnr+7q+Ca5/IVnK
xKBllZ3Z4xe0nzYzyWW3Upz90Qu95yJ3NzWtv/ro1mZOqqDw86lyzPBPm1mLsUdF
B72cDecsYxVyh1b0vReQl6qPd75rjot1rHx6FOP1yMrBWtKCo0kAS+A828QdEbFG
/8c14qbgdSfmcYzHs1cp5rXvBTqdO7ZA+luQR40M5zHdsSd49c/hFNijfgvQj8Qv
vwfdZ1wSGOTBDAi46LA8pbLFTb7jJY52h+4Q+iF8zdtXunk+E8NA/ZShPwwEqh/G
eqK5at9J5U7MADJUXu124UVFJ/r66uMHsgk80drcnJbnDFDHOvV3gZts8PFwKQU4
6hvj0irBebPa0mZIZZ2hOA5RDrWftK1lP8q6tffbb+9hy8CQHsEjYHAMXdhT7qce
Ur4onGIarX5q8XGI5OFxVq/Cd/2dGOrofWoGz9OwiD5G+NRpeTKp5aRyBpTZ0cY0
fqwi7bktsfUStNUsmIcek3Fi+g/DEhkEOWvOM7D1AtRkhKvxb7YbGjYGkMev6qwN
WYhwGlQrW5qlSgljy2KXiYbLFoGhsJP4DacE/dk8iUN2ND8WYoR6C7vxG+tt4Y8z
3FTx89nqgHZFny5AKGxawGPF5P93VMm4PKuru1WeXotN2Lbo7sD4H0dQWQxvS2za
/QRJeMMubkUEaSqPwo8QaSwNUgfOPx8IA3O6C/dl0ZOnDNLfPZEX9ub5X/NJD0ah
kTsgeo2w7ZHSlw1b1Eo42WH1Rq6GSfCybmJTd71Tv8GcxPFXnD2b2GReGKy/bh3a
p7czWvg9jhhWQFPBjJ88vL2lfMNGAnFefYr3oPuMUS661F3CysgGBD/8VOrvIjKr
LsU/PlDDvXw3CY4rFfXJG0Km05Kn5JNC5aXYp2Eu+cA4N7O+0466tlhyoYLy09sV
kFFf6FWnFLiHF+dT1ZKx5n5lQ80Ybl1lxyW6+1qbCUlCOMxFX3nXm+ts+PVaPttS
LodhF3iAlL5AmpPit78RwidaKmAhvZWWpRxAtRWRz98Pt3ep5wmn5V3gr0Pm3gbb
er/F94Sdp/SISI3DpVmBUTmuhYTFX+su1LgMCOTiO9RQVigRk8ADIdU9/xMQDeuO
ccmMWdypDKo1WFq4Vx4orwYMzY0OkehHDUPf6DHAjTpq5LN2sqe/uYKvuzP3qwsV
FrpHT3IxPJMDy1ltgKs2/GsmsPbmtTXvyu2Co8thDRMWaH0tSkwt7BDR+rjEvibP
AsdlycqeK4j1MNgfzLUrs8nln+iv9PYANXK1o5AcN5fVFzM5iX5x+g18xOZmnZXD
P5DFBn/4PyGpz2Oc9MH6dWMOAQTMANFcCnXrulyDNP7sYSa0ESO4y0EAxXXBkxrZ
AQQaPQusa63TJInJhhoOe4fJOXBaOwHXGOMW6rUluuDf+QxOfPbb/jMtcw9vPn67
Du3K0PmkFBEi3Ce+aEC/bynvzVHYwPhELV5sYS9W+NqjJuguyQz/Chxm8thDgwwD
ho+HkdGW9/1tLGqhO6vSCywfrGMduK+ia+0zQkNrdboSICWaqL97RDP0xFSDk9gP
fQNi51TYvp5dIR6+G7ohEtfqaI4/nPC+9e0Md+9eDGawuNnN648fW4zmsaXpI3lb
xzkERFouONVMOcSD5A+bgz8gwAGXH1bcHMNAc82fduThFi7SEz4ahB53JcC6gmOX
wsxDflueYl0Qss3fHHeN29hu6C47qto32GL/DfR+jd4Om4iDwDAX8yky7jkE0Mmv
sYJU4XEw4x7bTQF1w7wxoos7OuA8J2AUULFaoIDjpN/3mWdqkQNRUOhxFegizdOL
Mt3GurnTEoS28m+rmrVsSlTQ7JWCC5GrxE4CCMOFdkjOD9Ru8KJGVomDe1IFj0zF
lPJoK+Yyj37+/SbqspDKeLCk7GoKARAQqvHS9a4o/CHjSdYUlgjzehdNAggARDPj
97RttxVkA66K/rvVVpq2ASyxSitRwPtD7vzbKkvxWFcwWskLSkgIpHdiCOLef5ci
mv68KNL/wTKfRuIL3YCkhTRSOlu1UgK8/dvJtVr7+a54PmdhYpPB42/oW3qleNua
NlOqgsJXTtlJHaxGYJC2UU5uBVFucw8eO8aQVoBY17Y6Uaszh/8XAmZa9XdlVlcp
iOz4eZCvSltdV3fpjNtEdbhYO0Hf03zfIEg8ktHnX231mhvVk1rTVaLUUs5cdTnp
rD/BVmoN3+b3f+HJvpd6ogL3lW883tToIJTHtk19DcILgvYHpd/JKj+a+N0qQeet
1xhVaZ/QlbpbL/+nq/+ttjGSRZ1diA2WnhDPqyTMs53FFI+QrbFHBqWsUljB30YE
LgdciWx1+cwEuHQIPAHUKY2K62ohOeA9RLz3+CSMLN7U2sJtThNeihLX4CYztOTC
6Vdfa6bjV05BwSAxSR0aHTRpHCUoUzzsbF86LFhsfMBeMq5Lgg3gk7RO91ZTI9p7
zLa1WnzaEwRS5o+XAE537R7Wl4yBUATagLTDryPGlDWmPwbAslWqdR8wokPlKw6k
oYiiGdEuXHSc2IjjPJ90vFRIVz+pE9DTglJrdHPAEtwVdlbNyalrAWvbWcmvkjtP
9bBHwYz3c2bcwr9F9ndfzw2nyl6zUNl5Qsgz0EAZIZSg0wSGxUj+Q07WM0AxX9mf
EHF0/v7aW8EqhuqSL46Z7ZKEfFA+SVAQmoszJFErsWAxusaGKBOTsMEEeDZ02zS6
2LoLwkmJmFI6ID060IlyxFxeeGdp2fdwUP/K+XFCaLv2GrvdRiQ6MqH7bKkIFRpK
t7AXJi3sisp7OLFe7B36qBBmz9LbC3ELlMM9rbLZbKaAj0wfsePZgUmQOonllvgU
/5hEgkkBzQemnq9uRDUG9+9X65cAAnKLXhcEWvAxmdg2xfMLKYa0IeQEsYVKJo13
1Apb/G/5M5GFSMkpbpT96hHqg1VcjTAbhETLKzHTNsjzVMgm9RAVhvR9H5yjv0O4
MDCt4gBqZmpsWUBMssmkMy/2yrQGI1a+2p2E9XkW4NCwQL4UcmvKOUYxQ01vPVQ6
GXWC13MQ5XZUeyaxOPd+Op3FUNPYhZPOmQF5c9bNL9/r/TkoP2+mKpv/uq6YB3zy
vPzFLsNtc4r78q8iVJgvBTaDhbtr6YP/zaLjWMBHVsDZt0G8X2gbNt86b2QvmnlK
NPKvmuR4r3o/m4EZ9+sI3NoLV83vWT2b2VHKNN+p0LxAldv/A03hLmj579Gza+MS
OZ1vh5RAw9urn8UQEbYxExYXh9PGf3+OZiunV684VCb7JGa7S1sljMC1SHCgfv1Z
DBk5+skq+O3DtIxJsMeqQqwP7ZapKOMYFHmsU8L2V8kN5BBKrKJUgNiO1gwOfC9q
gQLeB8Xt+0ZgYqKtRpKoewAP/O3oaZVHpNKJ8NLk70X1KVmTvzlBqXekRql/Ri0v
9u4nWU5HmEu/vx4viYRUfNoJ9LWxpP0bd7qJPceu52HaWMROALpnfWIHP6B5TPOZ
cn3M+2XEbonIcOJlfjQE4+P/MIcb++cdEDngOqyi312TgYTMYi9l70c6hhnr3IEu
P1v9JuGh2oMk5vl5/SbuPOIObMrCGhnbGnaviOA9ExWl7KKGeBA7UP7NOk/1iAci
+lmc2ybfXKwr9eewpbAvnH9o1ugT8GRTdSZSjLJRhOqi2udxV6Cv2lfXQosWB/w6
zwWBIed24Vw2Pihpsu51P6/0gQEsOpi9WPrsGWTC2zc0OrjOO2EbVntWhLJHfpF7
XHOdUXw2VVvSS1QlNWjTHQzq0X/dV7X82VRj/6wdXW/O44urBQbTn61SjE3IEe61
ivjWXdDdGoMLqs4AK7oIBw+5yjm7Kl8V9NeWkef9d+5fa5RYa5Wa4NmaFysDpZHD
JKtwiNDr5WEr+ZVFylSF7MQ8mSQxxKlP/LJud78fomaAMyW8gN7mRCBqfQldhiO/
x+xfXzTL3s5V3qWj8s2xlgiK8ZxJVehQaXFl8TPbE29ILsgqSLbgKI6smP4KOxmU
7XR84dxa59lDCYnuIVAbG2JCCwkX/2jEuHbjiPPXnKCV+MKCPkX6bJeYTa0TFV16
vbawtSoS2qXNpCQwE+uafyGqajTLp4XM2SK/FEiKzD+GvWNElSYnTY1eyviyHlLJ
VvWAMzIYfCts2dHG64Xcpe4HhN2rJSY4Dr+DCIUyjV4AQ8990FzTdjuLxM2zt0UT
tQlK7noGMWsr0HqE/WEBiMDGBEpDzwodlfTjdo4gUV90dXXFzZjmI66K+nvdU8Eo
/dNqWPU1WBDOgJIdaaMDew==
`pragma protect end_protected
