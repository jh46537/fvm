��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&���2r�7^�(
b������G�����e.�� ��/�?�,:;ј+�9�����
�ɘk��<�Gs����q��D���3Q�z	+�)���2nl!
Xee�����7O���r���Cx������(U�]��lv��L���'�,�h�b� SG,Z��C>aϨ�����R�[&w����#��E�Z�[)PLҗ4���[\~���n��w������R�D�l��#`�}(=��ɈY�g6�zCCе��d	�I���n۰�`e7Q��k���'v�0���d�P��Ʀ�ʁV�P�.�
]�����V@�m�E��	]�ݖ���|)����*&Ӱ6�ܒU��o5雭j����)�L�H2B�ވ-v����~������&�G�'
\�8�����Q�U!��t_��qr�-�tq@��瞫��&?Q�lʥ��4�	���h��y:�#]�����<:w�(!�-J��M�em�;��1]//��L��V>Ǫd� 8�Z7��A� G����dG�i�@u	�0=ϊ��h�ӴLk�����!gb#�p�YVlp��%cޥu��ZhK��9�ɂm2���+��:���QM�������͇�䰋,MT�Y��'���ONY?���~����<j��r����d��ڸjF���	�@�	�2UgB�!�I<���)fz��U���'i%pF�@`�ƌf�
����W?���D=�FZ4�R�eu�j�c�S�֚ԓ�]*\q��@6H��K$֦_o�*u��[�\����&k�SP�C/�cHڜ���ᛡ��z>�S���%}�^yc��Z�Y�b �Y�H�B|��lt�3T�������س�;+t�9K���r�ܲ��A� $&V/�z�%��\�z�Jz) |ļ5��k[�$ˡ}�
��dž��z�{M�(��l�\��Aʏ����C���؄j}O�d�^��+�6���'ֵ_!"�0�$��YCbBa"2,k�WX��?�b�}�jU��RNH�}D����dK>m���wb  ��ܥ����\���]u��܊���;/w8��ܕ��'��
ۯ��z�	�ZnW>��Y�7)�O�/���7�e&$�8�_��Bu����C\�ݞL%��.��LU� �U�&RI�DY6����|VOġ����N�f�G�:`�I	�!��h�w�ӳ4�F#�\5��F��jH�چ �lb��ȒϚ�ĳz6�3���k\!�QD�|��=�D��D�Z�D|�J��je�ueѓ�����R[nȞI?0����[�p�����^�»�k��gs��plG>�����ܟ�$���5�O���~'ETT��e��~-�����bJl������R�S��g�x�l�N3d;Ɋe(��O�=b	 B^���An�Y4�_�05倣z8z�'e1�$)X:^h�Qg������!�_<���	O�vD��լ����J�fw��Y�c�:�� �[�۝cJӭ:�������ί�p���Q2���g3�C�bbv3sIt�=ޱ�s|(�!�5�Ek�ϣ��-:6�t?*����j�5��`��A&�FáС��ZVW2�T1�Mj�%I�ޒ�>�����A����M��f�h�!�*������umC��N\B�%w�M같��)�����.(��+멄��I�It��/��+f�t�K15�_���)T+w���cYY$��X-W��>�m?@��P�AW1�釓Q�rϻ]���w�̼U�0�W�l��8aC��g���×��Tp[��EF��MN*@e�~�-�ɹ�A�"�40,c����*V.�"w�jԆO�:\ʹ@"�@SMξ1zu~���>0f�
��n��pI�T�m��Aک��<���mXAf�`a���H�cI���y9o�t�<m#����������'���T宍��{N��0�Ho�yUT8���XzyM?u����_����qmN�V~zEA�>�����U��K7��,If��O1��4����Z_
����2��	�� �����ɾ��W��1�����`��(��\��U����IUؤS�Jn ^�
����a̠x������R�K�$��G�?�
���҅a�0��ٔ/�yg(���K\{9]\�"ؑ��V�n=�E5��r��L
j/'���[>���A�0���	��KQ��g5$�Gp�7�ϱ�HA���d���2d>��'����Msڼ:���i�i"���dl{8ۘ�f&����ÈΔ�q��n�u�X=\ʣ",�+�����z�Lr(�VK����p�(��7+x]a/N��i��	jH�+U$H�)H� D!ͭ� `O��
�^7��	Ƴ/��c	�7�՜~�PƩ����GMmmM�5	�|"���Ȫ�\�'��y�F��K�1W#bN���Y4�ؽ
+s��2	5
��E2Sg�[�`b��.I�r���$ȣg��z�,sQ���onց�������b��ϡ��w ��C�v�p ������Sc��|���"��14�O3��B!DR�=#�G�ٯ=���%�?���'�:X���+���4�})D2 �'�;�����tf����0�G*��(��:}�R���%��'��	��%Մ�n\�L,�<�l
m/����#��u�=���:����!򱢬)!x���+��@Л���/����m�<C$��N%��n�uke��L
7ا�`�К�l����	�_[��H��O�<_DU� �M�T�ɤ7�MbY�t��Նgj�������T�64�$�k����Px��;'ƥc�r2$~����~��2�т��t�����R� M���5�~�܃d�6Ͼ�pK�������-�m'�N�,�e�=�¶�Ζ*ܙ��B��p�r���ke4kخ��HXx�k�}�4�xȫ�U����62}�,��Qua�\�'I��ΜP��L@�1�5���N7��{�a0��=p�'*Ѕ'p�����V�NT�Nu<��<hX쬢�\�3>�����w���ѣfCWZ�ឺY�6����p*Q��\�q�Ï�Pb�7h�|L��ܠh�4��Q�v;>}5ƞ�k��;����bх�}o���M�+�_K�\)����}2�iN]����g5�X&��,�+�Pb#�F�Γ�a:�����f.0��^�Ѓs����^�I����O�Ӣ����96z�c)7��~65e~� �o��E�i[�y��RT���Ʒ��U&	@Ž�k���Nz9ר�N(^�����5��X͸�˷����gˌ�ܳzm[���[����5���6s��Z�6���!���0�f�63A�uѕ6�/P��� 6�[,���˳�/�ci6��(#�7�H��3�S�� x&��Z���J �	ǩK�㿈�5�Ć���z1����ي'�R�"y�y���zʹ���.��2���X"�k�dY����TD��g]VQ�q}!��q�{�dM%�
|ƾ,���&q����Y�%�q��X��^����:���,��S�Q6�*	�iԍ [�+��rEN�\B�u,��:����2����? �#��,��m��""*M�,�����P-<��΍��@������G*�_$�
nk�Fy�G�e��=���u

����ܩڌ�o�'	�����ohm�(r�nY~ s�!c��?e�K��Vi��م�R5����N"_�vg7�� ��g(j{jD;��_a��'_4�t�>9VJ�6����j5.�2%$D9�WL~(���j�����Y)ۃ��E��sC� �D ӌ��ꏣv2SO���6�@ �l���ԗf��ib�Y���&t�d��lsP�t�L��a���ݱ�'���Zy�bO�|�6�d�ϯ$��ᥙ�%-�A�$l�?���@���@�fv\��'���E��c�5��6R}�f=���h]����A2��ʺa�BA�ngWO:�dN��*�YAp����`��!��6Մf�1����=�ݸ��y ���AÚ�j�Qn�Ѥ�V�c�J`"��@D��]���ԥ�d"FIqxBH���؟��as`��*n��g}zF}Z^���lWC}��]j��f�k��~%Dח�Q��r�P �i�����,��p'ΐBf4��Ѵ����B��@с}q����Ꚑ���߬���Yr�0�Ģs6��!�]�O~�'X�䕂Wy�w��4J�!yEvH[�s3cbi�r�/|�� X9�l�].�ˠm�bxVO�eO��3���]�"�0d��wݷ�g�bP��l� M0U���V�%[�)C�s[J�f0Aѻ=�*���W�y�"��+���p$���{������e+lU�r�K�m�G��; �P���^���!F����L��?�z3nkH�2f�biolaY.{���3E
���ڢP��};���NE��x#�Ț�.72��U�rE"Cq`P�E��=u�3T��N Ru�F$�� �>��R�U��I��\�Cz0��0d����{7"V�W�ě^��8 y]i�G��D�x����_��Y��f�&[�<�H�R���U�'����>��;�����:���(��>��� {r�����`52��k����;�.FE�����kCkj�Y��3c;|ɥoN�����tksg��K��E吊�y�ε�W�"� y�H�焤g��8���[Ļ�5d�η".����T%��і�K4^G�x��Yc ����O/�D̭&t�i������Z�U:g���2- '�z�ҭ��1����{��v�c{�L+\�d� �mid/��x�W�h�`�z��o��"��qy���<eo+�HoN���=�ƾTZo����!��˗��L��?め�s�6�n�\i���:�V9se�"�
�@�\��ϧ�ԗg�+KkbF��+�tb����0՚%�P ����qRͯ��ur8�-3^ÓӾP`"(V����/@�?���%l?K�SB2��]��4h����:�f*T�'���L��lO���/d{x��}W�h3&Pȝ	94	�ھ�������<��%��7�=��&��)�n>#�c^7ʍ��aԴ`С��`��i��Hs��n{y��b� �!�t՛�T���Pc]������b����U�lO&��z�$$W���ڠ�
�+���j�AH`�����d�IǟQl�����ß\��*jMZ���}���j����a���P{��j���q�V�]t�����U [��i�����ݑ��:�o�����ED8�i:C�z}�I��{?�V������A��`�G�Ȫ�#��Ur&���lb9S���l*nP����7���S	���a�IM��ە2{�Z� �5��l(1��|l^=�δQ�N�Ypj��#@3�3�lWȺŬ T)Ja�
�lQL:����#uKƚ������%=����͊tV��-���g�fdK�����\Z
��c��"�Ua��N�ܭB@���U׍�o��l��v|���ry�K�\"��.
��Κ��C�5�n+j���T��B�4�6�{7�!��8��劌�b����8&|�|���T�S5՘wT�mA���ם�:����@�9x��`[��k�{;=ǿ����^�2��+���'H����d��m��߿��/�}��Z�ĽM���^Y�����d�g	��#v�5X�Τӄ��`ؽ�Ty�<�����ſ\�b��@%����2)':���Y��&�=U�]��3�l�����ɘ��Rc�O�%��û3MZݖ� ��A����+2�0yNU���A��<��0��0�����<���v���Y)��&��h�'���]Ux>�un-2�8�Vس�W��K���i6���n�6��XY�c�qN����ו3NP�����|�s�u�;�0��|����{{jMw��bX��m�g���K�p�hO�N
�`�<�Q�--��G@��m�#��r����vNĭ��[�h{�$M��R�Bh1���}��������X�6&vj�N���=��}�ߠ�H4=0�zB����7�J�L�	}?j���4R���cS	N�*�1�gS�̪�g��/��p��&�X���?���Q/��8�Ї��L',i�iFu��8a)�������ė �2��F���e��բ�ߧ�9��"�K���gVZ�?�p,)i�GXV���W�u�Mp]!�:fNY���R|�vnG0��_���<1�߷���G1�~>���T��Hpch���N�,Cա��R���ގ�
����.L�L����P10���Cx+�α{_����[�
�5u0�|�{B��4\|������H���"B���gn��c�0�Ť���oœzhi�5�O�bDe`��8���;�u�%d���K��&����~{�9��4�x z���5m	�i~����*�N���SL�^����6N�'��6���C�vA���:��+�v�Yy��yϨ��Yv�*�&�m����g��n���P᳝/�z��B��	���=	�A��lA}]�qi�/����w�E)��@�ԌI�>uk6mo=c��3�\3�>�ҝ�~cHi@+�0�)��K<�u�`�B��ûď��-CڅZ�\��U�BΏ�6򍬧����21�k�D>��hdN�R��=��ifr���ϻ/����d���!օaH�`�Z|��1�$�������S�"*�]pD<��(�rN��3`b .Uˉ�e����y�֙]t��āC�=_�f�BL�\�o=d)q���]��.r����n%k�����W�4*�#SM"y���	���J+���
��M�K�P��d��㥹ʢ�&ڱ�ɇ�N�����D��K�ҳ���g�<����dw,}���h����5�6�!�,oe�Q
�b?�y��4ɾ	�Lo��*�*��gu濻o�����C��c���'(b=����%=&&EO��];#M�1�/T}��*�##$�J�j������f�fF���ɤ�2
�l��fc[�[�*�slC���q"��Y4Wl��Ę�G�9[o�.ο�m��Br�1l�U��{���_{���݄/
�q�����yA���~BKmJW��l\�{�Rl��:r�ȨuWz��佝ٹ�+/����CNu�L/�S��j���tA>" �1 �7.3��St��_k H��F�[�b�ǲm�����cq���:��;�f-b��ܿ��b:^6���"���+���\�@�Hw����� �S�k2y�L��U�d��n��v�⃪�HS�(fgy�#<��i#l⮝��-d=�%7�HR����.�v\�bI~�
��<� �]�tΔ�i�
��]82�*��:k��q/6�kë4B�����zCk~`���wJ�����G�_1c�ȁ�Kp>c�E�������c�M��e�ڐN��1���%�TU��qlu�Go�/S�Q{�p������_ /���߄|wT��a���-�#��j~�$ס[{���l��Bw����D+�Ř/�贋I+�9͋?��R���g����K��?*+a��*T�ga�������rq;{f_���/�8Z �d��:$
��W�!1���$��a����e<_���31�?jF$���]4�zMK�j����S��OG���Ro<�:�\�����~jV��$	�7[�Ķ:��BŻ�� ���rp��)�*~"7;�I�me�8������%���J�K��-}�F�i��G֗���C[���d
�Y����jV���J���;�T�;���Ϟ	=$�1D��\������rx�:lnm\�*�V2�V�w�P[�3���޵����6��w`�T��殖>���.Z��`�W6Ϛ�B[&�g�XӇ#�
�ҹ��bh�3����L�=�[�xV��TY�!���
���eb��|_}�-���Ļ�]�4�{o �{�D1�\;���E�|�MW
R�e�{�9?����Ee�f�L)�Iq���Н\��S���i���7�����^����95sZ� =��"�k����Tq��TK!	*n����7��Kj߅�l;,���0����o*������a��u����!�j�OO�ذҖ`�W�˵���}���_C���P�/��`%�Zln-Va@,�x�J`*cwx�65�l힌���i�M�ِ̻8��r�o�+R���B�_���������H��gy��V16u�J������DsQ��| ]o�mQ���U�M���	r H��O.���Q��;�wV���$�}G-�����|H���4���gUe�����}��,`��Ic$�Z�H/�n�(X94�׍�*�/���V_
�	�o�ĝ�� H�~�شk��}hh �u%*�Y#	�-��i���FT���E���n��������E]^�����e|Vl�Y?�ƣ?�E����]�bM����W��Eɧ�ԑ���Ѷ*�6��R�����8" ѷ}��~��*j��f ��^����,�E��%?}?������рv��W�ܐ&8�~����}��L��='���=t��M^�M#�A�ΆL��ݭ"UM
�Ko� f��Xt���W��{� |�亄��9�0mg��%�h�h���1Gŝ�ݜ�Vۀ�P����Z�*]�P��2dvӉVRq�/���s�F�t&*w�6��Cx��|����]͡�K�W-�Rg�{�
�JM�K$4�>�f/(g�-%ĖX@O���603L?�X<������s/�;�>�]^\�運�:��K�����Z��'jű���B�U�c��~؈����[+�<Ą�OAJ�{��UC+
��e�R���]\׮���*@[+��Ζn�����a�.\N�72Nر�
`d��,U2팺��#�O3���ԨÈ~���J_��m��`�����!��J���k_;쌛�^���m��q6��ǃ����d��w��>ś�����:3XT���ѽ�p)��+���ZV��Rt����D�lM}�'>�iM~�n�;+�q+C�Q��e���F���FTd�Q��Jo�Xn�~�B<7x̵�i�kD���l�!�Ƃqp�X�6l�)/��2Zt��|5�����^�� ��蚤R�"�a}���fC<<����m�hӑ3YQ�c��F��C�*��!�z�����p����� �k�y�˅�G7��U�Ce/D&�z��͡���4�p��<ZS�%cP�J��z���B�E���"�S�ܬG���n�y�l�~"�P�bdT�9�K�7���D}���$v��ʾ�>�X��x�4�I"�����߽7�NVW�K\�>�ՍA\l<u�^��:3Ej~+K���	+��xb;�0�26�u��Ʌ\�D^T4����j+	��C���/���-����@�7W����E�;�eζڨ^_�|��2I����r#?-�j#A��������̨dʫ��l�&��o�/�B�r͌in�0���Ð%5F:���(Zݶ��S��B�c�X-)Ã�\�;(r���OtO��7�,���B�)����%x���V�[��l7�%��L�|E�t�m@���E�p����T�I�8^d"�R�Z#�5�R�Z��������s=�Ź3��ϗ��戎�p	ym�Ì��HFU(S���G	>"�~����Δ��I�ռ6F�p�ϫ��c�A`HԎ=)�g�8��ly�Ph�+Lͥ�l�+�L�mt��C�c�B�	ԠC~a��I�kbeOh
��}X��'�*��41�J�C�nS�,g�G�n��|dW�cI@]}�ε�IdA�G�f����u��n�S�;���l�ev����H�M�����5��z.�(�Y�9��ˠ��H�X�8aqM[w$�j%:'�+�`+#�� �u�&{��c�@@+��^�#��j��SC{��H��83_�&;��PS'��Gx�e]�.VO�>{���S�I*��%y��T��@�]�x�B�S��<��|4���)�h6��&u6&��Eyt����픏�%�/�{�s�#e1!�ͅ�`�1��L��`.��4�	`�m呷w��#7��ꭍ����!C6/̊Pr�z!���xa��\���� ���[��?(:!�2�Ỗ�����sI��B�%`xP�T�+)�qK�Snd�5]�g�6����K�3�XU�|i��o�}A�P���N]+�/�G��T8ٮ�EKf�^6H�ynҴ;�	�ʓ[����*Vj�w�"\/!��*��^�o~��2�6-�Ң�HߴaǓ�r��iCu�s�fݦ��1�*��!�r�d�u�^<�b����I_Pz�=�E�f!�e�F��7"���`�F~,dޱ��S~�^�֊l<>��%V��L�ED���o�ؿ�/(ʈ Wn����Xi%~!�<�_~��?�b)�3����.aRY�X�)�}��9	9����|/_������p9�qD�)}}Vd�3���T*�+s��F�"*�����2��+0���r
�����ûQ; �;��T)��|����6~ϓ�& �ƇS�.�\��E*��9�����u�U���dP
������f����Ji���1;7֞����u�|�K�L�R���T}��J���f�1�b���8�<��k�W�;mv�ܖ!�H	'$�CKz�Y���R���GU{v���^��`ʨ�D�U/��ӽ�@��o,Cn��1	�(V�A
�?�����ԕ�|i֤��1��D~��>�`;�|�?^K[�ѓ(�/]r�Q�&C$�w&n��V~9���1d�K�KҌ�^�4Ǜ+��-f�v�ʗ)�]jt��5 m!ԥ��,4��r	S����y�˺�:GY3�*�CX)�^`>�팿p�]�#���G3��#.�f{T��Eb̍'t�R�!Lo�u=�lq?$��A���_�ɵ�R
	���7�8�"x��z���p��9��4b�B���g}OL]�#��d<������p������a�e��G��{B_��ߎ�.x5<e��;f���`.#��i*��i�}����5�I����C�!p���;H�����P�Ÿs	B���ͦ�Z�F.��J(�(еQ��"�CPO&��L�;��=���ʞeA ��0��n�Vth�gJ�v
vG�'�wcl������O�4��-\��qc��~<�9]p��s%|ə�0;���D��fqY�Ws�w��H�2T�ovG
Jd�?8r�a�![4���j �6ú�P;�I�������I3�:m�ř
J����cF�TJ��KuQF��Q\���L�d�|�tԋ|)�f��/J���!E��B�I��"�	H�u�L˲��׼�*ֻ�������K!kB�^>�Q���fs�ڎ��	����_X[伛
��&i��"�*�%��`8S���й]��[�Ӹ�s��8��D��F~��H�vl�r��� ���=�m�h��~����i�Z�5@h���Hh�#���2e=�woDalǨ�4�Q��?p��:���T���N�4�̨K�B���ޙ$����>:�ϩ<�X��f%\�Qs��"*���Sf�eur�X��Z�p8Pa,�"��s��b�Y��ӽW���D����y�ơF���"1k����~���s<�kv+m"��ng�:���ג>�����ㄪ�������8I$�'a22��%�b�ݡJ�C7���?>ߡ �p�������^���ŜGu�1���t���=	
��Ҥ� ��w�% ���B�#���e�?��D<ݰ焭�R�|E�z�i���p>^�,b���ϛ�{��4e 6D�:�����A����{�n`>1��s��zS@K��#n�	p����Dh���h&�ݸ����^���ڹ-��9P ��.�`������d�p���F��B�!t1���h��I*Go�Fñ,IW�ˬ�2�e�	����������E�J�y4z;f��������2;�\ ȠW��\�{�P	��;Y�.�C���ߩ��KA�ۊ�]��bR���F߼9J�(9	^X�.��&L���zpb�vnT!$�Opu���Vۆ�P��=����<~�L�B(2��jI3��}������G�[�ɗ�.�W�h<-uF0b�-[�M���g89��LC��D�;R�7�LU��d���=��_�ʋ�&D��Pv����=n�2K�ҧ����2�d+�:�c��q6(~;����R|o<�TR\�y��8�x��?2digr�r�/�}du��=B>i� ��E��*�q*�}8����z|���u���tT�<�{c�Xr��9�K)���QMT�<�rOh�?��z*�eq�p#_s��̜C�e�K-���ePhӂ&i��q��m|t3Z�+��ޯ[W�v�)�@|��S�unX`�1N�>"�E��3'fƩ�ґM��ڼ���I�:�5H�"h^l�1Qm^���\�wu�a%�h��I�+�lVI�V���zU �+�uBW0gupA�B:1�$�o�c��� X��wxÔ�!p���_󘷈�G�ܱ�0�~��:�mݖ���"��l<�g ,R�0�l��q�w��+D����"X��:��:%[>�v�6�٤��Y
f��n��{������j"/�r/�SĉXɵ�}t��`0U�����x��p���>�5O9���L�"�Td�ZKj9�!�>�^"�P���7�}܄���1������m+P�{D����Z�������޿/5�hAWHzʆ�4���ċuJUX��K�`�yȅ�;
���x��5�~zf�A��zs�k���bU}�Z�v�%AP�Q�k���~���\.��s�mf[қ\�r�c��=�o�C����[�J�~�=x�s�lp%��(+�1�@:h�5�}w��
ꁶo����G@���TI1-�G���,4(n���ZW����4T�}):�,d4Us՚���Zz�ZP�5�ȖiH��,��.��)�[1�u-)˴K�3��x��V���x���FS�����M�x�Ŭ�iT�i����Q����ց�M�a�����b�6�4N�C���A2y-�d2�
��b�nu�3.P��J�oǩ؅�t>�Hp]�D�	]}x�=#�&OL���B�\���m���1Q]����B��W4���Q�$�T ��%Cd2~�˪�n�)��M�Z4S!e��|F`�O��P*��bB�����X�T�-T�����C�e��KC��-�h>c#l�)��Td��~����{�>I.�)� �Y��<��}%\���4��҅k���0gB�w�������/���bAI���R勐N���gª�A���yDE�g�K�~��n���]��ZN�u�Ͽ.��T�
=H)�t��-�p;�]����wt�2W_��ojE@���ݙ���SV�N��B�+��Y�և.z�AGI�\�`)Q/��R�<��J)���]�iZ���^$���mO���Ф�P�N�Һᫌ���z�1U\�B.�=����=�N-״�
�s�=��pAG����;�d�X�*mز��p>v���b��'�v���j�W����]Á��@i ��g�Y�O����d����0R���G�;ڂzb7�L.��'����z+�Ȟ 	ؽ9]ÍP�9�mJ�
C��ʢ�[���'ע~�7z�g�(�D��-�=8�9j�U��\�u�9�l����&�Vz��-��]��Vi���լ�3��I��F���!yʳv�"@\!Ih��@"1��oR��>��R��4�=J�s�<`T��.�9{���2H�tQ�EP@��z�ߦ6�Y�j����1U�����	"�nO�����4h��M/&�{HEX�N0u�*t �_Fz'���_�;˙�-P���wB�{d���Z+.���e4�tB�V�i�5I�;c�+��U�v�#=h|Ě)`���%4Ad�Ča_�����ENVD/ ���uS�2nRڭ�Y�(H�����:�V2T�"�	g���;3[	�O\���y/$kX0M�R�->%ۙ����Q�-�f�"9�R>@?A�:����=LKul�$,`��W�9̲^f~��K/���B�q<fG��+z�a��U�v�`	�%����"�5��˿-	/�Uo�IT���%�Ni��.�H�a��>��\+ڻ'�7�=?�uk�~��dB4�>�����`iQtO1H�6���]�S�?z-�3�1�Ɯ�RY��t�Jh	�MU��@�\�&�@e5N��E<��<Ⲡɘ�)��cf`!*������8��+K�`��هH(x����nެ�Ʒܬt��u�XG� �ڰrB���fِ��Z{�S����(;�Ϣ���(�3�)�O٫���r�YB��]A��nSB���YLAji�
�٘N�8��?
�!�D���q���T�Ϻ0Fg�C���
}�l�ȏNa��NL���>�%�������M���lZ��"��UN�CMb�E�sv�Ӈ�ւ�Λ�ˊ��t�0�%��i�v���B���sK��"����B0T���%T��uŮN�� ���,f|�?�Ba�?ruа��%E�w����݀��0�}v'�a�ݤF���3�}(�0:=��%X���v4�x����buF9E��;����~����U�$�ֿ�S4b5{�I���1�֬0ݗ�E�˟�t���n݀����~�Ϟ�����R6&�l`��
^��<���c��I������cg�6���DZ��R�"A��}V�kJ���8.�fd0[^�|�]{3cf��\�s�B}h���`��[
k�6K�K���O��F��V쒙�������������w��'���7RX,�ۻо�=��ϑR9~5]�uw���;�iԽ�=uA��l[0�1�����'Y6�=�B��14�@Y��T�%�" r�݂�����	��u�����Kqf�8Y��0r7��hEŨ����
���O�M���#]CB7o�e,nm�3�]
��KUf��N\����`&!�$F��lf9Bi�`�k={>��)�ݺ�������3�F�I�^���ݰ��׷�Q���}�rZ6�x65n��Ϭ���e�ʜ��<��+��1X�(�ǂ$�!D4<�, ��#X���ũ�q�s�R���xo@U��%��:=�������}�����l2��1����(o�֏�X���?U�����ff�f�����e��|v,��`Ś�S���V3'��d��f����/�v���x���R����L҇6��,��8U=�~A�P��,��_%00鍺�ظg���N�28��1��ֆZg��gU˟�����m��a>�!!�¼=���L�Z�my��rK���	64�N�E�2F�Pz��	��oj�v�����Ά	�+�5��TQN��ߗ��/�*���2����%	8&Pmd���X��G�4c;բ��`;�����E?Y+\�l�نA�挸��5�O*��<�N�,���GӉ'M��gM�j�>�t��|�@�4_x�T�9�x���;0)"�_j�!ܧH����۬C���F绵�W��ȹg74v!���
���{>('V�c?���<�\���(a.��:�$�_H��q"G�\�n�o��A��!���0��\d؜A����"$��Dp��(��iK�Dw0����q/�����j�e/�o���yJL��ʑ��2�m*��)�Njb�01�N�c,�+7���]O]4��JMꮊ�\�E&0��OSS	��/��"jp�ów�D`eA��ި��;Y�)p��P�|��#c�8���ǈஹ6!��I1�^x�󰟳%������*w� �Z�����"��� ����O{א)/|�P�tE��?,��������d��Qr6�v[�2���9*v�	�eFy��3A�)�I����g�Ɔ��'V/9�@B��&��M@��=	�XΒ�|;���ϟ��Q�����&��Ռ��R汊��H�nw6��Fa�-��i
���q�b���P���pO�sη%�H>���-=�%����YR���[*�+Y������3�5��m�f�:��H9G2I!�#XC2%�8z 3�b����B1[jG~6[�S�ePr�|�mzI݆�L�5V+�$�7@���)�%�z^�=��K��ko"PԮ���'>���&/#��b�.�R��u8��@>=����n��D���)oq�����b*���Z�]�T'd����R5�:��^ps?��6x���v�8�>z��	$?��r^���loI{|$[cޓV��Tp�J���d�����Q.����e�'�tbk�� t�[�Db�q��9r�,�� �9 ��|����L�):���>Z�w;�}���4���֓�Y��I�l]Wp~�4�|#<���@����+6?���`��EYB�r���\?@��'���{��� �@:T҇k��2Nãѩ�F�Ӭ�vd��6�kwR�٢P�xly�p��4{�Mc6�q�HV�M�X���y�HޅH�b����ik����Y�NŠ�D_�i."���#CB�?�(��A��	�)���@"�f�Ǔ�P�+����S%�bu�h��J��e��g�xs3/Y�z���������I@��b����_�>\�~�E�B,ƣeh+�H���.
U�i-����^�݊��0`��ܬ�e��˥��&b�0��΋���3���/��UI�:Z� ��=$��}��)�~J��Q��3��	C��ZK{��O����ux9̉jFOz�9TaK��S2QG�oÁ��l+��׉3����Յ�� FpV�#�%A:�����)�'��(Ya�����솵�1�y�N�� �>� ?���1��ǚ�$�]UZn=��ﲸ�A��r 8pP��l1�p�d��z��u�	u��(�)�ZI�� ��K�c��:}���]xtan���=l�D���X���.n�d�xQ�S<u��`a�Ŷ��nCn�
�K)�'�D��%c���V�Ժ48V/@�h����l��}�)q�:w�i��f��W�^���U!%[��1"���8��+��!b=��M	f�rߑݙsI|��|vJ[&�,*&7N�<:��AC�i���я�Z����>8=�S�Pb�"��d��NqF9-��	���[| ��O>���������@{�G��eP�/IO�qXdi1g�}���F���)�g'�H���`F����hA�ݒ���u��2	��J�)[%�z�wI�?���-�� <�
?��b��I��U�]����2!M?ܺNW�|y�+�x'��h�m]e�k)�vki��%D��daoo�ِS5dPݰXLI��Y-1a��H�Cu��#��ͥ�Y:������Dτ�L�
�nj����4% ��H��1�_X�{]�g��G�w!�%|�1�̹4�`"���i7�>\�Aӝ�*}���Z�r�6����#uT�|w!JNT�>�H-MeW���R��ni�X2�'[�EI%�7���֡Z�z�o8�&[kԾ'�,�NZ�F��0�Qn��|gns�95��e�19>������cA�#���E��)�9�V�(�� g�O���8By����愀�ϯ�ݲ
V��]1pn��4�vk��4�� W=�I��~���d;�!���Uv+��PEl������"���^q���٢h)�WH���̃���4y�X�n�@�B���\]\̓Kg��tVr����t����?V)�o=�� �J�9a�S�#b�?0q�#��>�QJ2f�!I?-�ľ;�u��p�'D$���9��q�,ǖ��^/h��������H�އǷ�C�=���a�pA?���`ٞP��@��o�G�MQ�G��4�NZg��n�-W7o�HfS���(S'~M�3Y�}�O��%�Vy��J|9ۧ�7�3 ����7����b�s\-42���A��������띁=O�R9��o;�������e��_�����<�.p��[� Ktv�A��r-r��NKܧ��Yx�O>G�/���bT#-�����c�I��Λ{4����W[���2�����V�@����GìB�)-�f�43�?XE �ۓ������~����BO�r���U�p2�<hY��|&���p���v��ĵx�dV�G���in�$���^��pnW���6w�{PXK�`�����ig&1�Е%E_J��mh�c����w�%�+�o+�逋�=���a.Fy��}�q���&��Q{j�iN�[��%�:V��| {��|��jW��=b�{-D�W�s���m�<��^����}��bҰ�z���J���HVgR�Q�mrFm�5Jp����ޢy9�²��T�R!�X8gь��k�'���#�	�״Y],&�͇rE<A\a��F��ֵ�z(���R(
}�"�?��w�ZJ���hd��}��{^K�溟.�#�#񣘁����D�N�A�A������c�hf��Q��E�"�C|%]FK^��%~�Z仃BYԽl<�<�G�~�/�2��z!�_= [h��&M�c���]ҴXn��ޓ�L#M���s�YmgF(�|�ۍ����<_�$��K���>���7��b	��Z�t܋�)�n\����W����|>ǉûZ&MO�#�'���/n��u�tJT��t��'��G��Gc�����+H��{5Ŧ�z"S�B�9P�Dm�)k(_6����X9�.���0�ӄ�\�m��"-Y�_�Dc�P4J��i��r�2P�'�T3ؤ�W���	�fp�署ƕe|ǠY�ߤ����湇��:���~����S��K��F4Q�5�\F�æ�	��r��l�.�{J��I!�	��iw��������)^�T�|�����]v��J�-rVZ`.������J��6��v~VE��|��(`�y��8*iϭ�M��x4 �6�7;(�P�l6�{�͔��qh�����n\$ ����!.4w�2L�T�|��y�T�h�)}�a�c�4����r⁂��`�� �tXPJ^�i֥��D�Kt�Uф��ք�Y��1˥��7���6�;}꘿�.�*?�F��Z��7ߍB��z*E�ł�q���#�w�WО�7�ml�>���l͂Jr�F���[7��4��o}ɽe��
�EѨ�hY�ڥ�9o�<�s��J$��7���7�����"����:���1��W��i��m�vQ&�.D���X��p��ZI�1���Vz`�q��_�_9ԝk�I'�1���R����n8�sL+ɖyo�M��6������:	+��J���j���Ա}����@��^qŮ�3�-�۱��le��Ϡ�))���C��0���pXc��ͯ���Wφ�T���"Y�.@X�.ф;��qtju�'�R��"� r�	sC��u1�����a��t��|2{W�0����c��
C����Ɉ�E�� J�H�!6����r�sH���hIL��>=f�i���":זCV�p�v>�-�N����vD -1)]����έ�+����K���/�&�;�4 \��d��Ͻ!��\�M������3i4�u?Q�_��F�SR��i`\��xE:/�(�j�k��Ž$e�34YF�z����!�B;p�"	Q���Wp�� �u�}�y�yq_=���t7�g}x� �0>K�Lnu�h���d����	[�-V���킀.���e��>/*��h_�L���J��N&���õڭ�k�L�|��Ag��cJ���`��rsy4v ��2��M�ݵz�.:�l2�Pl`�':�8����t,@�r�ֆ7��y�S[��ٴ���7Q9:�}%�Vc�������hԈ�"�+9���nTW���6�A��ʢ��m`A1#{��΀zq�f����%��"lUsˈD^cGt�m,�����U�V>iEwr�p��
�6��Cf�9��PǄ�.p2������b 5�^0���6����&�`:b=�@�~b<�nLMTK���ژ)�M<[$�n�3C�@�|���G,��/�Y�R����S�\��WNŊE�%��ՠ �x�z����W��|��P