��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����,��f9t���3>��Ձ�A�7M ��uj��M�0��{�ơ�Wa=Kg��!洭D�2�&�6����2�����X܋��x� ����G1���w�S��3�C�1�9��1+CH�<3�vwN��F�T�\#[�'I���ҒO*K��V�6�k%���D��Sn�&$Y�au��Q�/���OO .�XS}���9��k,[=0�hj��V���w��:g�!,;�(���1��+�\�dn�/x�o�+HWh�c$�f�!��e����o��do�d�_��X-s"�M��b�"��0mI.�r����~ד[%n^�X�ɉ�&�e��XC9�2"��E�w9s�c�������fڤa��Xoj����qy���ܸأR���5_3+�����փ�K�_�Uj��ȸ�D��N~�VG��Iu���f{"���U��H�`�%�bM����k�J��ԧ�6���b�x�4���ڭ��!��Q��y�~�9$���,\q�x��jSQ�g�;C�����k�x�^ϳ�T`����z�(��A�aM�$*�ם��s+��ǀ�e��RV��L%bE�n9�=�@B�h'��˶!�\��	å��������"�KݜCE\���#8`�O�ZO�[�;��P����ǹ7�ǟ&���ǳ��֬N:��[����cYw2(�o���P���*2�ε���5��R�������Z���F��^WE�X�o����	Vf�)5��~��/3�����)t�2N��ry&��܉��xD�G{�'	&l;%�D܍7V�+����M���n�֢:�+:�vUڹ�����0
���[�p&?0I�N/�������<a��r;�r���ÄR�c�fwvI�o+�Ż(��a�^o ��N�	F�|�1֮����"����l�o	0Ko�|�2T,�K���2�\�v?��lf����"=,�**a�R��޹	���V��j�6g�*�<��ow��I}���<�ĭ߷4׭�L[�B��+��������=xG�"��UɢWt�4�s���'������k�Jr��AQvM9C�{a�{�:��(]���}xJ�H2R�p�q��(�I�Tc�eG~�u��p�����>��l�sG���]��u�FS�_@3�˟q|��A�Ҧ�6�ı��<��}��7�c3��`p�V5�g锧�(-�S�K�����$V.��T�]�8ߛ�m0�����,;p��ʑ1��ed�Է���jM^R��H��)
B$a����d��
�f^�|N����m�]������r�"e�\TDA�8�a���$�i�~�(��o1�*�uɸ���*� �2�rB�\��AJ�Ypk2���-1'l��݉�!7��{�sB��:�_��ȥ���%^��%��?jP�k0����:,=XoT�E�����-��;�t�����"%KD��(�qG؃��'J�����Q����fV��� '�������~)s�φV�w�@�3~�kԕ�� ��B5�P©���С��d��,�&��1Tv*#e��l��?��v�l�����4}J����4JA�aoN+���������	[�qְ���ۙ+#&	[��s���X̦n��5խZIFb�3}��_'i�ze<�ĞP�{�˧t�Q<gZ=B�������%�$yt��5)l���r\gǅ��c*�Yp=<�a����M&�#����x�٬���/4����s�/��J�����j��Aw�hq�+DD;�_�xL6�x\e��'O?��ɧ0-��켾M!	,���kj(�~@+t�ۤ��y�< ܙ���"��p(�^��[^hG�y|����F=c6��H�
��X��c�4�G/V�x|{�Ҏ������E���[�ԓ��W�?�f��4
��.���g�Hr��&�Me�z9�œ�*u����4�O��t�!���;��x���X�ľ~X��\��SiX1����q�DRYqd�|xUk�^�r-���=���٨;�=G���Y�k_)���]S��ߝe1�E����K�Ib�z�U��?��L�d$�ke]�I����;Q�ȏ���rJ��	�e�Fw��j%�q�袷 ܶ�:0ʄ�ǦKS���<P#��_�:�����\�̎�g���ä���߻1�^�J�M��2Il͔�U�m��42�Lf>�!���<�QbDt=��:�f�d��Sj*��#��g��i�K�]	�c^�sd�6ژf|SQ��X,���ڔ�y��Id�tp�����>�5a?����L�	W	c��"}L>z����� d�HC���ӲI��5Iea��rf ��߷����`{Aң�`QX�t
E�����F�/m\{�ۛVb��+��CP�Kf��Y%�&Ⱃ(���Jm�/-.m��A�K��."��/Sh�s���r��?������~�\�(ٌ֋jr.���<��hG�/��#��㣺��?�bXΆ��o�\/}s"f�UQ���+��v˵���_-�����K�a�=��u�w*4I���z�0N��ʨ�Ѱ��b+����-�b!�~��I%W��M/ߠ���[阸�}*��wp_^w��ea������u�>��"�����Հ�&����aj.�����s���~���ڂ|fg����7�	��}��f��d3ki�S*��֫�-�y��7�馜p����Fz��ĸ$�����r�˝C��(�>�*9R\f�p�}[X�4�&= �%�#*��# ���jq
�~��e�44�vݗΨ��Xx���WQ-��Ysm�.v�����usׇHX[wÉi�"h�Y�!����hآR�R���WnK�ė�=��Nl�n%��ɋ.���c�U��zHU����A�b��gy�kj;�M�Æ�ʕ�L�g�:��nk]�P���鏜�x����|�����/d� ��d�'��M�4�om�.�N��<��`�;�5�S����.�s����ժ엖���x��ء�lfQ z���F&zR
���e�����
��ی/a�AgZ:p|	�91�&~S��l=t�;Q#X4Wp�t�˭m�u�6N��T^�H�<9�w� ���(���̒9m�Ʉu�5�n��u��d���N+�i�b�xl��-�e�t�d#�.�[ܱ���={�el���Y��7�x��X �r-�IF=�t����NԿ>L3&L}���y��*xL{�,�z.�wc�w���5�pY_<��-;}C��c����d5��}!�J�a����aH�M��S�{'�C0I�\�}�u�}���O��z�bz"�V����5H�뻨�v�~�G8%P����h��y	O�����Ak"��Ԅ;gW�I���o*_MR����Sոp���C��>�0��ƴ2V�.]N���bս|<���F46�T��Z���b���^�K��-	�Z	���ؐ��_;�B֜�em���~���J�!oڿ4s'�%��On@! 4�#7u�yw12Q3���#����n�~�� *��b"8�NUʾ�`�0cXE8�9��m����R?�K,1H��Q��2w�P�00}K0�۳P>��=˛�y�vOӆ��ε_���?�Z�؉Yu�\�FB��Qk�@�S|���t`g�@�`�j؋\�.E��������W��-��>�l�J���o?|�u~�G_s��gb(RT�=�[���H��!Z�[8,�Zs@;~6�ESX��]�R!e�R�v��� 0n��({��b�C�3*N����L^G҂���o,U�"�U1����MO���D,�C�a/�FQ��P�H��/U��^������ߟ;��y�:��T{�AZ�qlg�@O)ҬP��C�I�-t�ہ_���`��9'���T �p��Ӕ�O��\���^�R8�J^�4�+b�`Ն�w�UkڵnG����Ӛs��]��2J�k8��Z�:Sj�g��m?�����2I���ߤ��p�pD��X�"RD��g"c2�#}�'Nb`�k�J�ŋ!��Y�^�Xr�dJ~���?Uc@y��q��Q�IHL�E
ͺ�����;Q�)�[���-�����'g������MDt�!
ٷ��+��v�z�r<�g��@O�XK��{��Q���3Ί<g�]C;��a����e��it�1(z͝�}�E�%�W�2����+�$2�J��P�F�4�[4��@�h3���0�y�@(pHs�ؒ�?N�x���{<���=6�����_��B�Py�fQ f�F

����O�<7@��s��������}[@��%���սť���m�K�g��Jx�Ј[U�{�Ƭ�vL�a[����.���JH�ް���-c͗Va��j�v�1A�"��u��YO�����]�(�bYl)��0رK�a��!C�%���Y�����l�-x���&h����ֹ���net����%Ciиq�=t��������wU|�X��UG�ř/I�@�\K���k���-�]u�*�Ҿɋ+0�cy���ʟ��������l�k����9������عbs�١�<�j@�ȘQ�p��2�!欲`��!A�\���t�S���}��U�C}x@�A�U:v�Uu"��~ ����S��!Oi�Q�B�y����H�˗������E�%�	oJ�����WBt8&�TBQ�lR-���o%ƍr�#8�غΈmBt��JǇ�����p������(AV��GS�X��g�J�	8�&�l^"�O;�hp\�?�-�-qz�Ȧ�T�Ѵ�hx�~�
��9g>�<��\~��epÁ*i��5�� {�@��(L��;,�ч�dTab���@���
߫��W�/��d�˖�'I ���e��3�ǃ	p��b�0I�eώb�Ad����m �>�gg$�y��Ȼ����<��n䙯�m[m`�R��QO��MO]�/��.D�b7��S[�Z�lt��{��2s�Eh�z�3�m�+vd�g�.�j�l�~���������t��J]Z�&虇�*��p��8��󲠝Z���c2*��0a��Ѭ���6aӟS�3Oc :5�VZ6\���(�G�ds<������X���`T~#Z}#a�=����Z�fl31�K�I����o���k0�'pMĻϪ֦��$�"RT���l�U2{Y_y�.�Davo��+�]��*�������k���γQf�l)u��L[��<W��ؙK�_C"H!4����H*�mK��k�yX{VTu8��27.��g:��V�S����E>[��`�����ol�v�">%�!����G��w"���o�Q)���@�&:�~K�24��@��������8:����m����P��y������}��+o�e�`ܟ ��l���$B1���,�@��gl8�X�X؀��K��0oU)ߴ����o��ǷC��"+��I�G��[q�.�X���~�\_�K�]�:7{��������[u�=K]Z)��-�X'G4�u譏�Q����K�
g`_z	���nb�s��?3GRͤؽW��v�`�F�
ڐ�UU�R7d�rJq�nϙD�� �;3$ΟB+Ǘ�MX(|Z$���'�i��<��9}wn�%C�x`�[��^D�i��Q�������n0�r�g~�6��u�Py/���k��!�"�D�%L_�j�+�����_dwڦ���n���L�.}�u�ϛ���.��O��V��u81���f0�*��4���:5]��!�~�kb��E\��h�FL��9���k��?&x����!�`���+�Ó����X����h��#�+�kN�)���~ᑀ&s
�^1���5�k�*2���g�[CȤ$��N01a�yZ�+nS�h��F`����!D�T�Pbb�5	����ۄ0�Z�$r��b�gۺS|�b�Lۿw��P��	\و���q����/�_8��Q�R�@j݅�./�ɶ��!p.Wxv!:G6;�Go�E(�񗂇li��Y�����M��+�	�0����ޑy �@��+��� -�ʆ�b6 \y�_�u���[�Ɯ�w��������!vjo"��D�]���zc+�WzX)��nM6-�Գ�a�g|��X|g�)���}����j]�D�$�����t�n9��6� 	$h�z�I�n�$�f�v�6��#ª*��zN���*:j�D�w����_�_y�g7�7!�����QԵ�K�E�����Y][c��D�Z��kX��l� 4)���?��Է0n��w�]<� ���ې]+4��f8ud.�so�,z&����"/�d��ՕϢ��K�}&�d�<v�>M���r�y�h�6�с�x<��-r:���L���L������%��](`�|Qv����R��*�GZ@�F��&�a���T��|���<n���k�A�Ty�o�󵖅ƿ|/L��@G�{�λ���/41��%L^�Q	5���6`�;}YZ��J\�_�x4*2�/����q��!��	Y�H��W��O�� ���|m�^R��tJS����h��0��`���7jP3"���`J�~w�o�?� e$T���x��2/��>J������c6!l)��ҵ�[՝K�����F�Z�O
��R}m{{)�`^8���J�P������d<�{��i'B���ZϨ���e ś��X)�=2"w���C�ŧ��mr1˨r>x}ˋ�����Y�?����je�fr���}��G6Pz��A^� 
&\ ǲap*D7M���7�wU:��=rҦW� L@��t|oXN4�lC�������rш�R���z��)���(uĹ�%�6Ii^s@}Q����P�W�y���u��m���Yrn��f�~�cȿ���g[��nڰ^�-��J]��������>|/_�~A�xx<�^���_c%R��#�CD�~��0������Ax����!`��cmn�.���:hF������Ñ��T�b�ƚ�
o�q�{��MBB����*���֘�zn�� uϧZ8�� ,��:J�n�{�W�����jNMp�5�-��G��<d� 1��;�A��n{qJ��y��/d]�w^;0W|���A�w�rB�ʹfk�(������ p� y���)
�Ђ��r��O�J�8��L�uEv&D�=zc��]�>"f�o�����Ⱥ����I������s�V6��N�5��$�kҤt;�ƮG�͓�3�dde=ςC��w����&c��o!�ۈ�:���@8�U�$yF�⩃<h#��G3�����[ ��l�Oam�OZ����m,�\�b��8���B�7	�hW!����*0�odݫ}=����E� :#�ÎwEe��.7��J9��}u��
Ê�E�|j]#��	�o��k��%�
EO��gpecY-�G����@se�j� �2H����eɘ�i�?�o��F�ɞ����ҕK3Ҍ_'l�{�:I�:k=u�BGI$V�OlDa!��D�%}pjՄ��F(x7h�"����*5�b�j"�ZyJ3w<4Z��$���ԜJ$N�M��2��a���>H��܈L���w�щLC��m�[���τ��2��p���J�Z�y���_۱�ZX�p/Y��Q����:�9���~���(�8�����&�N~y�v��H�J'��c�H�q.�{�
I�v�שA��\�(�(�QQ�v�YQ�9����-�Q1�P���$'�&��8�0�n �*�F��!�L:���+F�PCˆſ"[C�LO�
�Ra�F��d�V I��2;ǰaSR�K�񇔜�([����뽓:�G�w�cjZ�\�	���Ӏ����~�$A����:�(�h��2�T��xʁO�e��
_/�.(�L q�d�窮�X_� �V,Q����f"r8&,�����F��uz���F_�*Tc�A���
4D���Ϳ #�S�:gV�"�Z�� 1	, 84�A�[q��hC�4u���8r�ľ�m^��G�$�һ�����s��F��!6B{�DDP}���c	3f�_a��N�ÂF���V8�G[��/�ֈV{{#����a7J�*�^�0���,���l21*
��@�U�Ss:�r`_Jo3η���Ǳ.���P�!E��V��u�޾��� }�ϊ�poVf#	��'I<�fr�b��T���@Q�Q����2~� �"�?e__@���E%�v����ʘwt�����'�X��]�U�/Z�P�����4�� tfv�΋/�������7����Q�+��p���O����6.�猨�f�Q
�\�S�}E�Q�0G$�|b��|����]�*�{|C(���\�G�Bu��_���O� �3J����+UN �O�!��XBOz�_S�n��w��hQa��-E���.e#z%_R���\�%��5�Y �(�Ŵ˸6쵮�"k��?�ѿX#�E�ʳ�:�Qtd%߲�vO�W�i�����{��A4��9S�?"�a�{D��s㤃�`K�p�X��I�y�p�`p?�y|6y��u�0�D���b.�@�7�6�u���PX�q�:��1f9"�)�b��H
���=E,���� y�M� 4�cԼ�����
3�G��6��ڪǴ�/>C�;�L�[��d�vjJa���˗e�v	'�w�<���2)z�z�_�\�#�E+V���d7|ʍ3����]$9�z�V���9�*��[@r9"�_�.�KE�ud��E� C���z{�e5���fng�ېiT�lS	&�&D�J�X�_?Dk��4��n��n����Jn;KI�y��u�˂=A�>FBܪ�~�<����?��_s�z��|X�����D�^f;��&���o`�D+��j�o϶}E�ý}d��i�|2��:��7���0s�h��#�l��^�y4ǢeL����RrY
v���J�$�b�m"�>����S����m�
rlm��/AG7�?��q*���1�ݵ�.Kͻ�j���ʶ*��hmlM��-�E=�,���Qv?�,�{.OK�~�	w�7Vm� JU��R!�sAg1�ӭ��jжAx������EOt��y뎷�e@�;�xy��M)~
2����4�A�2�]����S
N�8��ge�5:U�bN�N;���c��Q�-o���8W��P��9 #��l�D�����H*2ڒ̩��΄;�s+,jEu��^�kh�>�%�TQ�q�kJ�G�l��	42���d!�=�_PrLs�[ m6�A���Zզ�h��1�"VG��qYȋ?2�X㓦�����ɽ����Bf#��%�{+��e&a7r�OVQ�:�>3�B�]��V���]Xi�_�/8]d�G� �O�^[x6�P����׃�!�}�h�0ɀ� Ս�v�X���e�^*$4���֥�#��L��[�m��iX�[���;%��W�=g�ν�SŲ�V��p[<��Ω��n&��n{f:�\ � W!���m�V˂>���9��GԤ���>��!��&Sfއ�Z1��^"<��٠<�A�F]���7x_�@K��4z����p�q�:C�� �z�'g[�8�Z�Z�&=������wֿ���Uc��(����U�N�+��&T�5EZ�;x<�,{eR�� �_�;�Hv�(dE���-L�����1��;����ý嶺M)�X�t�򺖄�4�h�oL�E����t�#m53�
x.����7�WĻ�j ���� MP�̠E�%��/C*�B���*�$);sQ�	������~�]��d���� %�\�H夺kzwf�ҿ�z����@8���� .W;��R#˅Y�}�(�<fat`eg3$���=ogyq�oɻ��y�Fef���ߛ�������2�D2."�a�; �R<�X�U�b8ɻ����
V�6>�9Q�9L:�*�f��y�dQ-q7v�S�*�N��-��響�h����ea�Ì9Э
�ͭ����4C�'�NI|-_>X݌jkK������'��Q�,����+&�X�lp()���o��K��d� ��T�G5�����xE������$��nf~�-S��[:�3�6+���]���c�mG��Np#P{��p0#�BtL+�Ԝ9��-'g���I��QWwn�q����ț���_�p�~�����j.���ћ��i�Z�i���<�N��?�v%�{T��K���Z(5���T���VAd�c1�Il�<F뒼�ɸ�Q�6m{]oهE/�%�=�����i	���x>���m4�; \	��q��_	�����S}��.A
	Wb`]`ʛ0��7O�)l��=A�>w]F�yb~��}���j�����ZX3OOf]�{&��qy<p�f���ad�G^�+�X;�
��{��u����J~o`�d8!��<��@<�:�V� ���{���9���i~��,��"�ָF��6!�D�T%G�>�>��zՆ�y#ERpE����[F[=��~Hm��rJq��F?Ԋ���;̎h��ؠgc)yf� �=���9�jLr.*� w��@t�����ɱ�*��
��TvK��h�Q��A������l�~��B!
} ����!#��'���ى�Q�t���$�WVvio*����ی�+{���;�[ �'ߘ���P��"��m�L�,o���M��aT#��Ҏl��&��6��%������_����:�cDy�l$��D![�E��]����`�ƹ@�w��Q���*�7�6�,��f���\��j��k ���	�,�E���e�/*��T��5?����6��"T,xbg���i���߽wqɅN-EQ�=fk��A�8��
��7�L�b����?"zذc7&�#mÜ#~�{�﫸82v����]�ʹ�8��Y�Hk�j:���uU%�)��kq�j6^w��3
xU9��V����BK�q�@��Qj�����_���!�'TNk��h{3�*�ƈa�6:��w���&^��w��}�}�ѭ�,%@@\~{fkLU�z�6�̥��ޜӘO�Qs���Ef�>Ъ2A�
.����J�W�&2���m� m�����`�\��V��7�63�z)(��}J��ݡc�%�k����?�z#�h_Ƣ�R�������*G�ZY��k�L������Iύ��Y����C�<���/(\Ʃ{"���A]���K�D���L|�
�C9#	$i�ɸn���y��z>�|����^�*��m���8|�w�ɤ�co��s|f�E3�m�����sEܻ��ZZļ��sX���d����[��f�����5�JLe	{ȣr���v.�*z�N��遝x4FOyn.�U��h2k��Z �l�Q��x��G��Jqo�^a��Z�ǻ�k�y	�x4kz��Zٽ� '��A�j,�ы���)���r
����Q�����{u��9�.I�8;��gJ����{Tnʅ|��Ứ98��&^�J�d~+��$��.�Z��j�?�Fݽ����&���$�Z]Z͝�5��`5
	�	�\y�u~ʒ� �����v���VE��$�3Nm��P�y��?5evSxj��Xل�͎W(B��������m7.���ϛbdDwO�A�
kH#���8@~q��'���m��^�|�	b�ͪ�����*[���ƬO&�gP	ew!��1���;�e�Ѭę$�t+���dsT9�&�_~Y
�˼�}Xy���8��'u��n����^-���F)���b����ّ��8$\\+:E�{O|�-�W(G�����ߡ F�a������_{������v���AJ���*�� �+�}xk�"�ؾ�+ǉ�����(�O�����@���h����&�}Bo��0����ݰ����zDelX��Mͳc[����:�jN�7�qHʹ��G�W�$�ұH�a�A:��u�<mt����,�~��ù�Kxuݛ��?�����A.٭�2�zH�z��MxEϰ�c�y����.�	@^��}F*��7'S��8��-�!Fn�7?;H��|IN����E�����0f�7y-NI�?�!?�(B'�5F�m!��\$2'�������U$��㸧��|�u���4Nq�ʣ=~�	kG
�א]^͑�C���e��b���rN=*�.yn�E�����H���Z�ZC��LO���$�`l�e*wp6��kh�%��ݡk���� �r������.�p�u��'>@ys�u}�ϟ�;j����N��z�C�X2b�=�u��k/���ΕȚ������2�'�&�0��A ���[s56�ץ���̋R���Ȋ�\�c���?�Q�b�3"0�Pa���+u�,�{p�C�����P�:
�]P�6$/F{�ʠ�7�7@���� ,lRvepQ�0tn�p~���26��Ht�#�8w"�(��0i��QLo���r���(g9<��P/�aJ�9�tgb6��p�Ƥ��%�>�)�m��.@�����$�O �!���_B �z�/x��������8�0��@a��T�ڰ��������i^���u��E�K�oHHY�Z�GX��^V�m����R�p(9�}(�=_��XOv
xC����N�'�����N�������/p�.3$W1��9I�A�>��P'���u�*p󐨩���X�8וj�����	{S�IE׿�`+���`��GrL�JK�?ٖ�x�h���5��P84�4W\$��%U.����}��
�Yٶ_J!N)���Ey��r��ce�5R���vҼS���v�S���R;�Z@�Z�����q9b�2>�VU]�쨴���*-g:�T){h'��)�R��ϓK���a���c�>�����bKA:�d}1��XVB����SN�\�!W���aP���J�)��=��~	����ߐ� \��XRd�WdJ7���W�۠�P}q����R�-�/-��K��GH�� +O�9&�-R�򘅖�0U�A�����s8#^�8���nO���!J:�QH�Q��e���+�]�ˊ��rv��oK�Ng_d��U�tx�`�Z|*�޾o�s2Nh���u����W�ӀFuǞ�7���&���53�Ha���`���g[�.��<S��ޮx�S1%�ޱ��H�i�4�J��w�C���ֹVf!�8�1���KOIZ������s^ܮl�����1��T[����Sd_�X �T���X,D��V�qT�~�f��4tR}�� pvK-�ZK����Ry��_d0ֲ��q��H�BU�z"9�o�:��� �Ô����v���(��f=�H!���ZH?�pj�q�����+�����f]͟�������~��q���#\��x˩�@V��מ��<��8�&�\�Td�����H�sM��a$i%�+��uZJ��5B���:rq�����I���Isل��~o�$��j�����K�[�����Tg	��
�0�@��y�g�p���ܞ@v��i�ȵ�2�ٹ(���P_S�~o���ןH�P�V[+�Ĕ�`tc&��o�X�w�U���3#9��J�i��QAT�Ŷ�<�Ȫdȁϥt%�A#̹`9p�tu;J�����C�K3D\E�r������� �hŕ6D#݅kQo���BJ{tE*�+���KZ��m����,�&L��3'�᛼NEh�2��x���,:����+H!��p�mg}֭P�I,�pۇ&�d:�},y,Ѳ��-�2q��}'���NfQP�<-��N�(xd;��^Wϕ� ɌJ�[�������{y��)�M,���,_K�a[��jw�x�}o��ȅ�d4�F8�"�V~x�w�ۭg�"	s}K�`��>"'��6s�br7�����}*#_:���N�$�����4���ÈB����4�.�f���R����w�ڊ(��6Z������i�:�5�F��^�~�����Ҿb�4]I� (�w���"���&5O�>m�:K�NYZ�����غ~����Sm�H��>G�aB�}�Z�\Ֆ����U���r���#n�J-�V��R�s|�(�P�ob&k��9�ܡꌵ�Bt']����E�(�G-'B�VO,;�D�vf��1�06���Y�`?R/��9yO�	�%��r��k믭uND�*��רm�&l�h�I�ޛHbWA���K�<Z{7w��e��Aw!����rP�K��?K/1�F����eL���Wx5��O�mMA�V"Ly�(�_)0 ��B|�v�Q�0im�@wʀ`W��exH�F\!��i����h���[e���ݕ\�LdD�~�R�_��(t�,�ܸمg6f�����*�59U����3���[Α�S(��i0�����VO�HP�d�9LV�E\���ԝg���l$�'�����7���KIm���K�E.�tM�W~��%�eN�5AY:�W�hZ���+�JP_q7�����K��������D5��Ss{�E�a�7D>���8��؛���jH��Z6�P�Gn��4i o�H���Sx�+�V78��S�f����7��2X�ɼ`lr�����r��e/����!H�z�����+���d9��vu�t��0Z_�O�L�ߗz��L���#�W���>��u��V�13C�[��J�[Us� 6�<��p����q�fw�V��~y�b3�$�u40w /P�g��� (Cq�\>��W!�R?{����_��]�yMQ�J[tmQ+�k-��� .e���7-��Xb[��{
��@�D�.��R���T��/��s�=,����sl垍3�]߲I�3IwK�_V?D��`Tosg���,ϯOA
��@ӶbOY}�5^���^W3��C��8� �?�[�	�o��k�d��6��0���:;�`^��I�k�������~�bb�� �c�+O|̢��Q�3'�]N|W%;2����O˵A
\@Yf������j{J�G�qƬ8�3�g72c.|
��5�o#�C��u�I��'`�[&18�-���[[°-Y�����3�{p�q(�a�#w�~ϼrS��Ƅ���P�ዽN	�DoS5��=�/F�~T�A���*�H��o�3�G��/�ο?�^�o?i���T��mL����G�0V"���� ��ZBI��C�ä�V��k*{k�ur�h�� ��\^�[�j��5�O�Tm�op��*ߕP[���>?�{�����]��鉵4D���W���7�>��sD*�j"��2�>��R-x��A����y�H�,��hX�ۇ�nϫ�i�������s}��1�>Q�{j�BiM��|�k ����J�?�V^u��MU5/G���BY8;�ߘ7���z�5vx�9~u������mXv�S��h� ͳ�_l*e"x�\�Xς��N
��	�㘏�&���d�7��8'�T��:թ���Һ��M�7�|�c"�8�c����k�/&��L�;��=&�[u�9��{~^�_/�ב_���XA�y�����븂�ִc�H���<:��}og�kˑ�-?��M"��eA�+�:��dޅ��~�4� ��MT����hrǱ0�W����.��u�S�i��?sa��"��0��3���n��p�1���l�{󉣏md��'w��q��v.-��[˼�(�B��Q�>E#�����( ����e,��H��a�X���![���S�`̄C=a��x�l�k6c5����-W�:�M;�^�%�7�y�BĪJYy�̸D�W�|=߂VJ,�(�8�Zp��.���y�uKE���8 �:O��O�h;�c�-�`^��g���_[��7cn���E/�S�HXI�����Q�k�w �s���K�u��W������ě� ��f��lv}��y�,��y�Ps�~���i[+H�U�����C?j��E��$�<�$��n!3��XZ�kT��t���]텮D�ze"����Θ�o	��&S�?|&ke"�G6����?o���3�1,�g��h|zP�����ZY�M��)��10�1!�
��$û)&�NJ5�t�_��[�~���9��_R����X����{ 7�3_ޘ'#�~�)�<O�%�+2�~7-�$X����Vs7L����T�) �������#�i3�%�掉pG��Z����-�e�j���� �c�3������ewlğ�AӐ�������\���	�c�̃P����>�9�d������u��d�W�1og]���ǧ�"��*Wm�Y�^�K��@Vs3}���߁�|���TYYY�uP�5AQ3D�:��i5y�үl�+��ȵ8�F���ъX���,g���/�Bя-�ia?E������!}��o�Dg�2|QB6s��0g�!��[}6������j���h��F�g%~��u��M��hu�ZC�k2̓}غ,fm�*6��i\��9�6��#�=��9��L!a���P(��n�啰Ŏ�2!�H`_!4\B�Ov}r%U֞Y�U�ߍ��͟�Rwe��f����̜��lY��&�TKL�{�t¡��nE|Z4��`s�e��:Zķ`D)Sz���?���t���C�JS���Q� �C�����TW' �Bgs��X��F��	�d���Cfd��3>遚���?�:��<�~�gu�y"ೋ+�=�_�d��!CYV3u!�!�Y�F�<�����e����E
�!XQ��[��4Ը�4��sl������[��M���MM$=�	��L�y�k�_jE*x;� �E"ipp�JeV�q�HL�+66�d˝	>[�(�k$;�|g}a��Cd��;N޶og�gЃ���L��O�θ9����= �n��|��%�;�e�O���0S4����w��3q�4]��!$���������1��~��Fʒ�P̙}��]QK��R^6�[?�ur�XuY3��1[z3Y���D�0�N�t�ȜZh��R,�,6�6���Nrs���9�Q�S�=�h�E�_O)U��nk����A:d���?o���U��&:�S���R�0h���x�D�Y/9���V��S��f�Ғ�'īzW����I�:lW���G/Z&�K�'	1�P�*��bN)�?3��f�VwihT�G}T��IU���^*P�<��ð�8D(���	vWt&)��T�Q��9����e���|l�3� B�����cQf���9
݁���T#Үْ��g��huهh�V���b��l�`|=B"}��;��0)T�P�]f[F>�RB%�8A�H=�'0"`EW���9��p�~��m�Zֆ�~@���n��.����bM���<�ԙ����aq�յ�	%���.�3�XޠE�v.�R�����s���j$q� �38�/F�wk�j>�Uҙ�%E�� �]L�H�Fl��Ӹ:щ�g�_m�ѩ������M�Y6z��@\W��(��^ukS��F)���2i#��Ƹ:�n���[�kP�TL�T�j���1eoe�]�+�hZ�ĺ�v���������RܢR��3���h(,����&�-�5=yA�^�M3~��D�=���$��zU�:���4�4�,�%������� �	\������}C�6��s�-�q[j�$t���V{d8�A�Z{6}�/����H�?�OA�%��q�A����Z���pU�b��`<;�H�o/�@G΀�`L>���5��رi7�߃���5�f�T�ϼ}�F���H~��)k��`4_s�"���(\cԸ�w����?vZl�`zIU��e��o)�%O׏6��ˀ�-K�ˁP�Np��c�ó�J9��tz)d�9$Y;"Cd_�92	����(0b����$~=��4O�y`
�����${~���k���C�[�V�f}��i86�EA�#�>u�H���C�:�l�	�0�-��#U)C���!߀X��k��E��(�kR?�7D�<3���74t���їIh=t^$�Si�K>���='�$�剡3�)���d�VAj�D�f[��mgf�����1�#�
�L�$��Z6Ϣ�Lx��^��Lj�A>h���]���~e�eRc�	�M/��asA^/�,(}S�΋8�K���R��a�;|����q���2E�h�k��j�c-�o\�䥋�a�_/�������X�L���9���lmW�,Gqs�䒊�~̲?��p�T��1��sP0y4�@8���ވs���#��k�Ooq鳲Z�:��U�����TS
mC	�y�V�XVKVC��xG��(��%�����4ecg���xb�0��x(�k���gj������{��0�5�7%��<08L�V������O�|�s��?z�t����͍�1��Ԏ��X9i�D�Π�"�e��%���G��Z�]�f��w>�ݓF"'��:������X{"[�{�kEk��
�	o�k)���� �Iɽ-=��
��ɻ�u[�8�ێ��0�x�U��j���f�s�;�ar�,�	nBFY���n�+܆�v��j�;)*�%����t��;Vу�4G�/vJaa�?睩��⚸}�,uԎ=�Z�'^��-$U�O�*�"WE��R���'�^1�֟��� (C�ƪnb�P�*іN�UW�<�P�9/�G�(
����`.�e��Z__�!y����g��$��pɓ,�sͮ�I;�ZA��N���X����J�U���-�b������,E� W���9 �S���uAXdǟ|��q3m0K�IơkA�����ڭ4���u�\j���v��l�1]#���G����s�c$m�[�*$(Mr+�� 	�d+b����~1����㊍�h��4�;�Ԑ��q���l�}"8Ň�Nq��g�ifeKR�kY�NR3�Z�$�n���i:,�Oɛ�z������@�&�)��'~/L��{���A{3ܾ�p���m����O�ސ̐�㿞�E�Bw�Ӡ?'�_�u��eI���
���iW{s�?��,��%��ՋsK��sőS�)>	���$X� }��Q� �ʑ	C������Q�?@&E&:�zR��A��(�Á�/Gp��9ֈ��g�γn��������=�L.]ĺM���!!*�t�q&����K��f�����T��w�*70k��Y�]#�Ps��q��U���F�v�* �uV��.A��؄���|e2���o �S��/1܋G�������UPa� o�$�P�o{8�_	���,x�)ż(W�V@}�wV���T�ͽ�u��Cn%��o�@���kܗI�/(�e�%�fV0C5��F�z'^��l5Y}�X��#y}Y;�����c���ғgYG��HDn�l�$����5M�=�)���Ћb�|��FrW����h9k�A����
��O�sDcE}����4*5|ɅQZ>t����8��+��{0-�N.�_�+�CD�Ա �#V���6� �������X*I���#!�L�Al[����s��\/�g�2��R��q�z�m�ޭ�BӐ@Z�r�6YM�ʼ��W�&U�s.^_գ?X�[P��E_�u���*οھ�Hy�tŴ�Y.�\i� ��S��xcy�ȵ�~,�'��^^SL�W;Bjl4Ŋ����9��ؓ�;�-��U�VdM:�7wL��*��9c���z�j"��2̹�"V��		8x�(I'�߅d�{e,�#��ь��Ke­��¶ܖ���o�L�
��� �z��]��فj�w��U.F[�����FX��Y"������M�h��~�b����vz{LV~�it�GS�lv�V����7�+�؁&q�"~���5��.x�v�&�8Y#�͜V~@˥n;�i�����OY��Ox�-2x�P΃J���]^�Ŧ�%���!��|9VkT����S$��ҕ`�$��j�z��Q�E��R���w�����@�(�t>�1����#=Â�=v0��lRx��#V�2m"���B� eL�2y���"o'0q!콣s� 5	\��xDT��'P���.��I�ڳ�ў����0e``�X�����hrO�`6pᴧKk8��%��濽�_҅��~Vy��ĐNX:�y 4�|�	%��U��AB�ǜ�z3��8Z�鬹�D�z9��0�̄x�N��zY�F�ɋ��ٱ��6sb����K7d��*��frs�K��<����1ڔ{k��Ve��WR2���i�i��J�7Fh�b&�1���� ��m��;F��sRA#����9�jȕ��t��T��7��E
LvU�{��r�kT`����G��%���Į��:���Jd�	����6�=�վ���!P%���>����r}?��~9o�K�o�j�iD�i�h��њ�#�DT/tNNO)�	Q�ߨ*̣'
���L��¬C���~�/
�<
�L����G�,����b� �˝@V�m�=#��s�K�/)�9�v�>�l��Z��52V�Q��&a�7���p�����xH4�+�BgnX�ŕ|�c�*V���YR���!� L;SIس�"����͓��w%����;]��o�8K��OK���e��͇��GM*9���=i�� 5�6��*��d�΅),;/@t��$�RE�U�4&DMt=V.��b�J��C����H%|�zK����*�7�2���H�iw�.g��m�h������H��~jL��,Z�#V�Z�C�v�t������ߓM����|�i�1w%�F޽7�w7����	&~[,��Ԉy�a�XD�Z-��\-��=�Ҕ�d�s����k��ʫc�����ԣg��^]�T��7�Â����`�~������#���;S���f"�ڬ���~�R#�����K�*�	�}	}�s���$󎣄ұJ�D`��׎l�g��wC�T�$����Z�*��WKO���)}l��\z�j�l�"��NҬ��<�g��f�-�ݓ͋�^��h���1�q�
lv�j�Q��4��3������*��+�S�(
�����м4�����8Ϳ[#����)Z�&A^�8�C#K�p5u)���@	,Ř�"<��L/F��g9�X��^�@�y�X2������6���=��w\A�Ij"����[�s�"CBeg��� -J�R\�
�{u9���:v�R�D�1�n.P<섡#UH�~pg�a��魾D�O�WwdUR��@}��r.���ǂ�$��_n(hXk�f����V��G�#�~�����v�7ֱ�V�	�9���1
�56?��zWJ����!Q6�Hz	���.}���������]s���-��*���"yy��tVy�Q>^��iU�;�'4�L��a�}@���y�T��W��Z�g[��}Њ�U*%��GwSb!�ݲ���c6_�\-�����}���T<�/�"���+�v����n5�'ke����S�Od�@�����k��j�al�7 z�9m�z�ߕ_���"V+�?��$�G���� �z���)N�F]�06�[�-o���"�ݫDhV�nR7�H����y�202>M�F��vmy�%�I��̬E��P�����N�0>y��b�K��		1�thEp�8��ϰ2>����"���N��@᩸'%�z*q���}�`������d�Y�=��p����y%y��I=q��أK�'���e�(� R|۱1��l!���ʻ(��>�v�
��F�)�v}�=w�s8�ԃ�N�.�xN���ppa�g��g���>V���wX�X��ِpN|�_�,���F���}�G����f�X5uiw���VW	����s9H�怋X�q�O������B�Ҫ<�Pz1 �p���g�E�������۞��\�
��FYP��t-F��zS�AI�1�S�ͨ�����B)��1��[� W}�>�M��e��р�7���糔E9B|ALh5��e�q����ga�#~�IYo&o�b�!�4w�g���Y%�b/iX�Ȟ�~���6��B�����Z��_��������?1هi�z:��r|��:Ot*KƇ����B�.μpva;:�w�j���Qw�}�]��?!oJ�-�A�Fψ�������'�0jᬣ��k�]	!�A"�[���~��@h_�HbM��t4T�TӪiZ�.�H%�74`{�|C��V]�(��vZG�(�I|����f!(-���8����">t&vϼ�:QQ��*W"�7&}6G��v5/̈́�ł��z�Ѭ�N�s��d277��w��-�V{�~���T�O�����L��y�\ �3$)B[�4e����8���-1K��C�o!h4�	F+��At��H�m�)n[�~�@
�P���E/������nt(?4\�SE�G�8�������J<�z��f�z�0��Q�}����C��Q�-/�=Ӟ!�?,7ίe��v���(��MOz��դ�������Q�Gvf��A��̉�Tu*h.g�Q>b�kh������_���+V�g��)C̸U���⿙�n�9O`���4g��co�d�/��q$���Ǎ��Ʒ�¡������
��E��]����V��Vb�t+G���O�>�w�hs��a�R��=h"��� ���s7%���!H۷U�����ϝ��1��N�өL����t{��
��4��w<��+^ �<��J�?�/�TX�<?��
&dA�d�� �Zilv�}O`9M1�b��ct�o�2�R�^����g�2-�04*)aZ>$X���?�ޒ�� ?K���|���*�YJ�U7]��T�`����ȉ=�Ĝ��*ۧ0��E3���f>B Y���7�����m���h�y���VM7�ftC���Kz�#�6x��}t��س1��&�c سS�{>�3��d�&]F
��m�$�摿��se*���������G�-ͤ*��ZuP�;�E� �I/Q۬�7����h��(o3%9�훀��A��w�{��V�c��l��hf�gC�A6AkZ��6��y�a��0�!��~��5CbD�@�r��!c�b��JH�a�H��m�k��Nɰ��k�1#ː'U������M
*	�+�/���	ׯ�W52{�E�&��ի��w@�%Ƿf�� ��Zׇʎ渪A5��Bry�X8@H�A(�%�8H�[M�Jw�y��:���R�c���(��?e�����G7���8��R������,[���S�;���~���7e<,�ro�}Ə4q���`�죣��xQ�/F�0�s�kru���5!���@���\u�(��bx�w�,{C�cRv?Y���i��h/(a��qƮ�k/*Re��UX
���4{ ��t��0Y��8��5D7�'}0׻6��BKc_?>��b���4'x/��du��d�w���F�6uyq&�Q���|�m��-l�[^?�����+SzwVC��:7,3��s�f^���\�9+f<��9��X�:F���tT��h�l*�\�[�(N*�F.l���5i�,���>��O$���E
d< ��.i��@����셦����SI����Ql]F�?�V/�O�� �5��|�����S�&+`l�P.gi�r���Y]�&���=��f<�)���6����� :�^�8��Xr� ����쬖0���JS /j���V�%yj2�:����C����xٮl�U&��,�|1�=>�V��5-R��>,�\_�15[�O�-I�B��{�xtOUA�_���$�1"������
B3'K����9�W�s��/�##��y/<���%���QaЂ�>t��2W���"�0��3e7je�6������qH%�}�z."r	��f"Uz}���hj$k��i�DO@�q��Vy�OW=R~=fJ-�-^�'�eQ��&�����Z�:����}��ĩa*S��7��CQ^~�	�����r����g���uQ69O+V8��lR����N�>�u�n7�0�oUD-��*o��~�M@���g�u�ڊ���}#6��%ú��jY��d�5�	C�tP��$4t��l�>��Y 1��oRi��EQęc�_�<�:]�s}�\�2ۖ�5e�8��/$Ly�R=i���L�������.8K�'���]T��=�H�e"0A�2*���W�*���h�/�O��F�ȶ�����j�T��Hd 7�s=gv)*C��"o�mcP=��p=�G]��YwMs��?�M_F��(D4�&U&�l���,�N�[Oɯ�/=��!O���T
h�C�6H�r4x���À����G��Lu[	�-w�e%���yt��8-s]�7�|���%�\�� ��xp>fP�=�|��K22l��X�`�v�^���wot�#rr�-�Vs[�����*ć��볉��.Ǘ�b���N���ȵԵcp�����6�ܮy�={�L5r�9������;
r+�?�M Yw˲����y�@Pp?� �"e1�I�#Yէ���!�'�H�UyU�|�JC�;�{v�B��z��Jџw�i�islL>��Pe3t��N.���ԩA�m¬�_A�,iH�&1���xo9{�
�k{ n�H�^]���G/�rr*�DLX��%	�GF
6HJ�ł�[v�D3���
���.qR-���������
'q�������2�(2qtqsz�
)?�Խ"��rP�"G�>��#�s� ���ޟ�ve��:��=uHә�U�����@��Ri2r�1����0¢naQ`�~��'X�b0�M�ڍ�`�~�1>��y�ޓ�蜛G��Z�J|[�þ0:fL|�}�(-<_smk�(yo[����Mvj��>��8�N}|�7�4�څ߃qo��H�e�	���}�}���M���t|7�P�e�� ��o.����a^�h������8LD#``��S��ӊڸذ����۸��+���4)yE�2S���,�?�k�!�6|y����p���o���ќ��?�&Q��-0��/��<\���1fH�<�Q���D�����$C (%�IY�C�E�i�r�$'�ǖ��_���&(۽A�9�r"��{���j��e$� Dzß���"|�q���$4o6�ud	���S_�|>��K����/�i�Fd�%ru��i�B�2�޸g�Rc������'����R1R�s�,�6g9&T�q���",}��.�sr/3�Vn�x8nY'=J*��N>��Ϊ� �t�ܙ�r��cJy�`&Y��T��0C{BKB�i8f��͕����z�o|C�L���h���EA̔�қ���+_6�/d���ƔQ���{�ܨ.�G\�Z��7��g�Z8r�����2nj�aTW�^�9�DɃ��ZPr 7���y�v;S��HU�JW�'��&	�GL�H�"`�� ��U(R%��Q��Ħ���9x���1;|�� q���mx�n\�9�����[~�+�Lid-ʟ
�m�ȕN·Ah+ʋ	a�Ȩϕ���]� tKs��"���ȸ����+{cj�c��T�ۄ�s^�^�h�������9��#U!ȭ�J(o]m:�E~+.	K\hUN�v�PB4�_����u��o���oy{�P]#F���5���Rb�+���Qئ��J�ZQ�
��y�w-H�������y�=��v�#�>�+5
�N���EA��s��L�� �+��9
@�ud��X��tE��9���A,JS�QC�,kC�׎���F���Y,�A��2O���̬�:fIm���"Jx�m8g��v%޶��7xWQi�}�Vg%`!����.�>9��:���;��xf��3
�4�3pc�h��<靰9U�;�b��ju��a�5@;��uwco���G����2�"s��]=1�N�٬p��)W��(o�"�~<3��I�a��NV-�5:M`v�,k�Ѻu������O c	��\�	�?P���.	�÷� ����%#�
�*?�.���������~� ��i�X�2+�L����N��#
á��!^1�@ ���X���9��4���fH7��
w�����i�'�T�Y2�2��n�H�Z0�υ���y�b�H��8��i����FB&@4q���h^ZX� -�>���م'N�"^�)Y��V�-S9�������8mA)7r��g����]�<�m�],� 7���]�-�EI_��o5���Bo�x�}�<��Db�5M/�Y;����2��.<�����V`[wa4��~ע<>/<y�z�}LH/��1���eŲ���9(}%#�����!������*�ǂZ��G,1���E�L��}�v|�}�#=�[rs���N��A��P��FEH5u��6��V�iC�E�����`O?G�����e��ou��])�eE��N����}TW�v����c��{�;B�"v�_���8��:���*�J`<�j��p�f77@���W�� 6E��G��	C��dn^�VS�}�����������׵� �x���,EfD�GTcH;��A~u{��+C��y����������q0!��_2m��v�7V�����F5���-��D�Υ�����=Wg�9B�	Q6#5�`C]%m�^	�v7$�\~�sTb(���2P�c����.�aGHxOB&��ٶi[������~(�>⌘��ľ�����n��\iFe���4K2i��I�Yξö׬u�W �pާ�#�W��x�),��q��������	L�ퟳ�����1%��c-X0�g���
3��M)���YnX��􆛡��K䓗zdM1~{�b�����Y���F+A[�<�leC��H��Z���ڕ��N�y`�bA�� ˩+����4���]�����;���r�\����ߪ�ӑ�ظ��������}���G�a�bo��@R��u��,���IJ$ssxh�L�2�]��Xe��I�����¸�`��`x_u|j�vE��;%0�}dw?���-a��Gf�Y�a	|�Եv�_K�8���
H��W[�8�!b�����'�,�� 2�_�B>[��"�;�Υl�籛���#���D��F���Xt���|p��Y�e�,��C}�ȕg�x��9��x��4�pw1�êed��r�a���ci8����„��Hc��'��]Z+5���ux�G��?�����_�d�����Å���z�d�j� �%�[���C>�O�ժ���m�W�+��~�bc`j���W��<��T�.-a�ܹ�1��s�L�U�jv��%Qo��A�O�ʋ�����6$��W78�I�l֭�8^����+�I��dˈ�j[B�֫�����n_�	�E�rP�C�lY�s��f�wV�)�P0���B�11�㰠nY�� ������$�D�^�@��We"ј��gPl�=!0!����TIy���c��fn`�H<q���W.#�p�S�S@����䂖Dɠ4aǥ�դqe�&u�~��I�]��o)�޾�`�?� U:[5���@����TS��1*��^�^�lC��C��eO�-��6��X,��yM�f?NහZV�Ʌ��:Y���+�G�a���9�_������U̐����-�q`�qYoV<�.0���w.��[ܥ�<W�.[�c�5j�Dp9�W/���:y�U4x��4����M�����7'|N��j:���5�	��60���_b�����+]FyӾ�Ҙ��ξr*���(��Xo�_W$���l��?$��8p'�~����8��F��2"����+��Q��X�0((=^��O���Ӻ{a�9�j�/a�����{��3A���),F��`�J� �������@�l;v-��ZJ\P;n?<gm�~2�+�<��h�g�kǳ��+DZTr�����h��'�rC��	Je��[G�:����D�W*��\gЊ�o	��y���%J�]���+��S�Z���;\ڡS�(o����ܖ����Pd������^�~�J!D'�CxZ�D�E�9l:�R�db��.?�M�[�wދB�="�V�l��S�V-�F���R<�)Ƴ�:�	T��{��r4��s������w�X��k�a����Q�t5�Fd6>VoQ�o<Жp{tRf�I��ǣ�0F�IC�Nn:�G/7:����&����
K� �5��-�&��&g��f�nf�)��Ρ\o 6݈�O+O����({5�t$/A7������#��H��M�.�*�Y�2�=�9�`����Y�K���vQt����nTJ.g������Q�K���q�#~�������)$����ܧ�^�i
����&70��+P�Mrܟǃ���V�XAW�X&���>2s���/ExO$Y��h���I��[�8"�Vp�����Sa�~Y�1A��9	CC���U�2�粛�@׏�Ii8y.7ؗ{5�'�$��*�v�d���i«�����vRO��v�Y�4/�!�T�z�
�h��}��Ƴ^59%��r�>��T{"5�����G~Y~&��Ħ�����z��]�U�X��f4Q� �C l��@����]���jP�%}ӻ��%�,8�O﨓����D�'6[��ڐ "N7���" ��J��]ς~h�{���┛-f���\�l�ͮ��cB�bb�T�.�i�E<&�#�mL�?^�t[�G�77���ݵC�4^A�!�bz����������"�W�z$�G� ����8d��n�h�<����8�ɲ$rߟG���e��.�O�Qz���ȹ�oe�/��&j򎃷E��S�Rq��\���l��p7�3�up΋xD1�!����]�u	Y�<�_��!7��7Q���W3B��&f��f2e��I<O���ȸ�'�$��B�kfj��J������ѭa~_$d�S�'� ����V�I��5M�#�]F1fW�����b���Ą�d��R��dD�:b�r@�ґ�0��\�i;6c��y%�\����aߴ��3)�`�F��L4+��B�s���+�-
\6Z���y�+Б��g]����|ιG�[����)f���]�!�?]��*�Av�%����ct��@x:�pqn�S}�[v�j���GtAYЀ�"9�ݐ��6����8Ѹȉ���Jh��J�[��
��ݮ����*��C ��y�<)��/H�2b xT_�0���]I�Eapp�5m��ڡ���O&
�}\�~w���r��&���u�zY`=V��xw��+7�c����a�s��jd��J�k�Qk�ɦK;qI1Jb?O{X͘ʾ�*t=RX�(��GC�ǁ�m��''.%]̑E��R!�qb�;?����▒(p�^��r�,hV>��208
s��G
S�9>-H�|i��A�Wڥ�^��!z81*1��������}�i�=�H�<���Wœim����o�M�n�@W�[eR�Lࠡ]�-&�\g鬒Jz�cV����'�j〙��i#�df��0D�O���h �1NP��S̻��e]<�N!i��r1R�[`��9�����	Ir�J�z7��ݻ���T���!D��R���ri0t�rF֏D(��� ��}�[|�ذfj�r��� ]���ї� *��u{jʭ~�O��.���ȴ ��}60I}���Q%3�f$���h�`����K�:n76k]��F���V��l��(�6�h�Vl"��	��oN6��ZDq�8�%�3��D {����	<�2:�G�7r-�3<4I�ep0�G=$�T�u-l� Q�b�/6k(�\RH2SAb?7�^1��81���ޠ
�����`1p�H�^��;�|R6U�I�,��v���=�u4be1φғ��]�j��FtVt��M�	y
�4�5���%�۰,[�J���8�W�_sy�2��޾�9�JH�{���v$�g�+��{��y�0&R4ˆ�̭�O���aɛ&hK!b&���9bp# �q2��e�~"j�Pf�"�f��z����m �*a�#�O`��L�
�1^�	�;�l\�_�!A=��D�kJ0�T�4�L�k�S�����?�G�\��o��Vrl{Z�o�+˘�Q�O�	M���1���Y8��z)���0D��x�u[��?��0�+��V���L���[9 D�s��j��a��rB?�b���{��H�I!��F�)��E>(d���M����67h��Lm�ߛ|Mx1��E�?=[gXY��ܻ��ϟ���N�߇?�˵Ӿ�o���� :��u�|B{Ƌ�ƃ޸��K5X���N����-��mmWy�;<��{X��L��`\�>Ɩul�mV�Yf���"�����*�j����>�@�N9�tLt��ζ�N��5�����n���5_�c�R�R�1�͹&��Yr�TkXf��R@*��H��c�9��Aa�/�]c���h��>�2�RY�L*F �!�@�^G_����^�7�?�X�(�J���*�
�~�9)`��z�oD��QZ&^aQ�ے2<��K��*�������m0�Ҹ!�DƏ'&����i�A��붟-&u��n����ӝy��ʵ��?r��Ե�s�&wi���mVo�����V��>q?���i?��o�Z��Ҧ�Ukt{eY��E%`g񼜮B U�x��(�ku��3	��&��#^�������,(�9�^��&�p+�E�[-hn"�بt;G�~��59̄TI�G�H2MH����m�h��3r���\Z>	�U
f��P�v	�۩NԿ|����/�%U�'8W��$��n8�@Q���r�L������\���kڶ>��*����-t�'bu�{O@^s��q`�d+r�/D���20dU���{��ޖe��x�|k������0��|)OPe�?m͠�������Quu�<�O޹��XO��^�]��,%��/Uލ8�<D$��sl�0W̄��q�['�z����:ιc(�=~�{�e~x��P����@B�� ���rA�=��o��]X['Kv6y��k@��[?f	��<�����/�_*(�����$w�}Y�����z�a'ۡ��������1R9O~6�w��{��T0sdm�# w�p�����b��Ҕ�bf�7NLVQ4Υ�<G�3�m�gg��,E��`��%����з���a�:W�l*����ZH[$�g�������i�`^s�->W=�1��,7Fbo5U���qi$���>s�I�in�y=u�ލ�L�w���a�?�>H�����"* �����2x�	n��y{0�h�_@Z��J�2����Ά{p
*�|(q��.ۇ���M/+��o0��O��i��������{�Xv�d��{	����w�w�Y�2 �V�{]�Y�d�;5sT���h;�r�F��+�����X�}�-�P�ۑND����T�T,�"�^�߆so���J������x�@l���S��Ǡ�4h̪�ՉD��v����{�t��
���̱�ssK6=�njN�jI����e�����S�C��1E)�&km�f���s�g���6��-�cd�z����¬ =�G�'*�����Q������Sh�ۼ��leo��{U������Xe�:��hP �C�yqg�|wƫA�p�|v��߼� V��<Q���L����C�D?�[�����}ԩ1
�Y n�S���.k�6��S��������0��1�.�d�QGݕ��g��R����m��
����n�K@�Ux6��]�Ʌ�e"G/i3���'��y��X/@���Q쳁���TZHX��<
L<����ln��L�/���(��懩 �l�6�d���HH"֕���c��� �4Jfu����2���/4�ʱ{�9�$��_	_���U[S=ʲ�燛(�����T2�5
���P���P?�oFw�lM偋��-C�̼쏉t �LC�_˔�l9�û��<�|L���<�1S��(|���S�l(8GM�]U����>x��7Bn�:(USv�	��c ��h<Fu�q��J�q���Q���?�ox�����pWL�X�w��G<��[�����q� �apBՕ�VrU�"�qLc�%��2�)̀s��,TS���_���*[��k�W>�4��IML=��k�Vܝ��p�2����.L��`b6���#�D�����2n�D��~�͓?z�԰�(^K���U�@���ϡ�08��]�Հ�y8��G��4�\�X�o���ݵ��%��`d.����R����˺�jGE:���{7-�3[����Fw���;�u��5�l��T篘���9�B���6�Q���o�QWXx���л)�d3�j��]0�>3�3��)N������h�ʱ�D�����9���x+,i╾	�\ڃ_���yh��q�!���3#���C� )�Uz�mV[�2�
����������Տ�*(ѐ=�d�ǴMa��s��Ҍ��=5|��|�󙣬���G���5�>��񑈠�6��G��5��uJzF�90JO��9�����8tۃ���W��3���!��6��6�F%���\1�,�1%�d�̆��N������@J ���r��ɠ=��>p?�h�� �P��&�*��gcll�N���E�+�\f�g�#S�eпl�4�; }#�s�؄W�|�|z�����.���EF�2��ܡp���c���P�-Rc��S	!V�����?���w���X��6I��_��`�C�P��1zrp���>�l���Ztm/8�n����K��Q+�Y�~�_G�	�#&����S�Z2�V"r4Qz�[�p��خ����Pj��Q-�1� Pzn �"��~�h��^d2Yw�p��*�8��Ky\�Pj�}�xv�v���ܫ��X��t�{F���\��7*S��=���''��K\��|#��h}˵]�Px��L���`X��.�~�:�yYM�MD�1�.'����r6�V�g�6uJ�e/�?�'�+[�;*b���4�1+2�N<^<�.?����5Ts@��L��"�����f�n��?��Sx���C��d�+���ӭ6�#�B #��Y΢a�ě0*vD��n^�wsb���-�� ����]M_#8k��a)��^T�s�њONY2�,L��&�R�D9or�<v�u]�C��&��$�[��B�dEŵ���;C��:N��g|�����(*f��G�����C`�|;K�G@���Q�a��/����2t	&��k@ �t��1��s��{'V�f�QX�\ɾ�yz聄�t�F��Jz'�2�ۮL��m�5�C��A��%���Y񾐤LDR�>Jg]>�8~�c��gb�z���]}�31ju	�^��w��V���Ic��X�q� ���:���~�߄����M���S?��؜�/�0�->WZ>�H�ej����\�bwa��w����:�-�ƍj�Q/�"��;���9�e~M�O�r�$�����{�P�1��C�pUQxr��r���s2B�/�X�Pb@�%ؾSd���D,�;-��w؋@� KaE��������=;Vl��c�<��c�Fjn��P�?���}�-g<~��r�!��i�&��!��XCD�mV��8#�\�A���Jl��~��ק&�y�˜�['��8]\�_��0|k�]Z�/��Bv��d� �B��{Ҹ��S��f�<M9���YgeZ��]Aҿ|A��@���0�_ Z���a�KB�H�-�����7;� �*�DJ2<P�B���~t��6d׶�x�(%^�U$9p�у�!��ih@M�*Tv�\T&��&�r���$:������lX���t�3���"����9+''R������qѱC�n����E�Zz2�12���+CԹ%��,񍗠q�e���|(����)��#��`Lsk�u>Hd+]vr�Q������N�����J{�S�ü����h���r�Wk�0�)	���8�fx�g�D~�7����]z����q#�D���YV�qO(�x��xD?�[��,���B��Q<)�(�wT��x�5�[f�/�Q0� ��v�vZ�X9��'���W�N�����XFP�]��8��mkZ��8�B����q��S�6�ӆB�9Y��$�<C3.�a-~�om`��w���1g��~���H��9�s]	��J���-���*�M=m��5�m�?�WOR��GQv,�!�}��\F]]��h�GAd%�wL��T^}�����"ҔK��%�i��<U�}?���pP"2�r��[���}p����6�"[�Ɖ���~S{���fm��g��7����Q9�s�,����]���e�1���S�Q��,Jn��,��v����P�W���_�� D��`��E
xK����.c<�+A�3���2!uZA����e1F	�e���]�Qs��ꡮE*Q�錦Y֚>���D)MV=�o�r�������r�����(�#赹��jV��?�a��[��՛���ʻ�Nx�qF����h~B"�4�2}��Ŧ�������+1�Ũc��n�
q6���G>ޭC��KR ��ԅ��BǐRÆj���x�ܵS0�x��\�cw=SN�f`ط�����W	����N ������jd�b���V`�� �]��bsL�1m/h*�^O���у�@c"E����6�>^s?�w�?E������`5��k��+q�\��y�����3�ۓ�r�DQ���e���5ݺ���%6}�MK&�����-hS0�\WxO-��Uú������WS)�����`0�kw���]�f���r]�� ���i5"!̻�Yi�� 3Rq�����ԯ��4�L%�V�V=N����!�w=� Զ!}u���o>��C��F�Q�^�L&�c�:���/�,*v�F�큉]��&�"� ]Җ�����*���!1S@�s�3@��QX���\_�Ӎ�;�b�fBw��+%��7h��.��٬�4�jȭ�*亴a�����,y����t�Cۆ6i5)y�{h��1�]�f�%[q`$�`���`o6"���Wjﮋ�u�
d�r������_���8�ĥ�_��
�b����\�ϘR����[�g�PЗe��[q���l��4������AF�s�@����_Ș~���od7���J;�n����砼\�EJʴ_�sx6S�����)��i�(E9������0����O-��d㹓�#�P�|� c�F������ɻO�/�w��F�[�P�o�e���1�?���V���JP�:�v�Hj��v�ƍn(R��|�m�4���VzwD}��֋Ą���l�/�(�(/��r���/�N��-��/�"��DXU�"ů�&�Jbݟ����l� ��*˾��`{�D����m�9�WM}J���X��*�o^�F�YɎ�I�0{�
��q(����}�U"��" .w__���"9D���?����1�y������l>�qg9��ڥ44�a�n�������>��#pܖa��p���1��v�J�r�o)�/��?;��XG����S�P�3(h�DO�����/F!���ܝ����~�؜ږ���hS��g�U\K�P�T�`b2'�7(��p9�+pc9�D]��#_|�������m�&�����
�K�[�*o����L�Q�5���n!<�tc&A��I|�b�� =*��ܽ,��r��,��a�s~�,��n<��"��]L��_�S\�+��
�1)� =�R���+ E�'�?6���S��`���J���6M�}��O�sU��IV��
������ǸF"��o��q���S��Ͷ�(kO֤kp^0b�k�EX��j���(�U�j��iZ��	��MKʧ!����&"Y^P����e��N�6�0�\K��Ǵ��ə\K��箚�p��׍�T��I���?��c���#�!��H�ŷۮpM!�OW�^�um�%�r�\u��R�?��h��y�χ��&�ƴ�
��ԡ_��H�M<a��P���[���<2.�.6��C:1f�o�[N�D�J'��V���b��+�"͠��r0�,�Gz�u�f`�rn�"��g���E��q<ݵ�ד����(`o]Ō߹LF�*,"��~V}hw�rO*I@b��o�Em&�" ]���^U�J��G��J��If�(����(]j�ek���F� r��*�X�ג���R���e��?}�f��8W��ެ����O�߭�Ϲ����+�����p�+P�ߢ~�Z�e�qTk�� ���V��-%��.�v�8�G>]�~ߙ�r�"*B�&�fo�;#3V��!x�Ƀjӓ�����B7�D�S�h����6�/�vZ�<�t�)�Ҵ@��/�6�x�=z����+�XqNF��{��B\g�����;a��d0�>�pq�H���rkm�ȇT�u�^ �!n�e'��;'{�^�&=)T���6\W�^�q��5��Z��_��Ү8�~�i۾×k�vˇ���@s=p\��4��T��__�P1�H���]c5���⛲�C;��ς������(���
����,���w�jĚ�T���<L.j7�ӆI35v��Fi5�t�����z�Xc}���\�ǣ��m	�	��Ŝ� ��<B�b���'�����Z�E��=C����g�Z�OG�W�t˗^n�\8<poo��VV�dFHw�����:�K6�5����z��W�"���=�)E���X�Fּ1��G���9���C��
ᩧ����qN�L�x����E�%�u�u��D,�����k�7f�{��4���	@��8�e�0����1����I�j])���3�>��+�N�����e���$��*��>d6����k>�L T�uN���"��(�}�򠖌u�tJ{��+`d"��ƽ
HQ[���K�BX+D%�3j������?X�1C�,H��\h��Pc�'����k�Ca�8`[ 3M:���� �Ѻj��Q��?sB?�U��;ۓ