// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JVpIb/YM8FtoYXDBxJWG7RRyP7Eian3piqSdse0WSYlMa1253FPissKcZbWI4cjB
VCiHYj2rnoosgqCOM5hMBlMcxOaRHf//Yf8N6weE0KntqsItBj8tysQDbO616JG9
Z95O0mfR4HguTzEOKgYDGqL+JTW76WOq8KbV5oq5h2Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31440)
bOOkoUtXWu+fR2QLpXH/JWBvObyvatf7LG46Bc5kybzTLefu/O57WcRYZcVY4CxN
o3g675h1RqvUTNGIP+Z/uokYi792AWsptyIyZctA4StKVX3G6JdWOOyz1euyd91u
97wQL3Wc+DLsZaP8muqxbOmN+T5Q8yPWFhNPGC0QgyddXWR9YOBNS6wo/3h9ANhr
syEiWGXXnoLKyloXvagBnKnPFrARtZ/RE8tP6ZxCYZhl/+Lotu3ZY9TWeoQS7Rrq
aeu4EuusAn+nN45QjiJT9gD2NIqMTwCW3l9J00zsUnmRvQy/Uc5FHtEogPuF8BdF
MAZe8i8cxC2TbHLhlRfbSd/AZB/wjCOP9vQo/Qm8WuZwN2YVGkmIHMyV8FYkRECf
q6gz28mkLivpWhEfi7+faLi3m5QCzqS0VEQhQHoia2lzxNKJb1X2nCQjuCNJosig
a3B/7QzwGnn53DqEinlHNb8jdMtBTG0KM4MTQ0lASiFjOCml/70z5aN3SkZIb0Ya
kSrvVtPDKmahbH4B/a6vJjiarjlwVtPBl3hpGC5pKFRmsk6c3n4s/8wtIvUoLpb+
eP3gRkuM/K60HqNToTFdgSbGBhT7ruZNTzuQa9iNgXZAmWRigo4oeV+fJiwAu+jP
1h06fDFDiCvFAo/D6yxtFqyrh+bNDwbYhBVh0qHjfeX0mjz3gw7ar6riZLxJenIM
xyW8kavRDAAQjm49+tMjfTUw8Uq9Tr25D8FAOzO1ScTgHxbwMyNCi7PpvvHF6jtL
4sA4BZ51XZRii6Qd0QsLYXhwjwsP6/bRClDrEWMlxXXI1QXZmfqw1oDuddSWbRmw
ZhUZet3z05wc3eVaNt9cq+PPeWbEsXj/JofKKAG0ZkvX5EKEd1o0uts+bpRe+rZY
zL/ycb6VfbFpmpasx6slbBVeLCESaMdFEquKJWxKqeIyVWyFD+XNMpIEGssg82QN
VEqbiTb8cWqqAGeRAy4iMd0VEcrkdsbLCGamYn36dNDQj0PycDjs2X3lQ3Ipwzik
l+CWmUci22dslrSkOjx7auTVwvP5UceOFoesEu6XH8P9S2ULXFdjFXAjOyYVNNeH
SggIHxgOo0GhR5DQB40AyEFWh3fyXttvyFW3HgyItmiLsFN6+uNp1CLzB/5qWFXP
EiFQI9SMsx+IiXyP6/sxklz0f66RPDTwYS2DgnDDse/cLRmqbhKDsWaGz66vDQq6
mxZed2ra5u50GW7qYGnjax19kqF6sXELCcr0EsYTf+feLiyYM3KR3A1hdxt5GHBG
TwyiECGVLx9Cir40KIqR3t7nddAvryrVbgfq/F5qRBTJoztBrRqRkXZtGeI4TB18
BdguJNFCu9HHImwSdHaBa10zG1wWNkJ4QRsjolHnO1m3cnwKi9fluSeVWa03xTNd
YUF2PWnqx0TK47MdhTxUFkWyv6SdxYcpOg83dZ+LqFDsmfdbVe6O/Yty2NnC+1xr
9FTGNmqc/eKrBoIztv9Ok4gCKPhKEFMIuZRneY8mYCy06mXgjoO3tTDH4CAfQTEf
/FAhERwuXUbB5iUwtwzsqpK6ZPtIC3tyLImf+vSIbA+/kdOSUjx6BdpJdTs8PXKq
WZBwiq02adhccBlFJQryfEADU7eNSc8prxYpQccJaA1zJ6jWub+Nau+BvVrGgeTy
ke1h/FnMnluzerGyoZb8KY+GLcPEESryQQkO7NgNCwsuthPO90nsyHaiDeC3HckG
HAYKpySllaKus/ahcFgC98rLgFcK2IshRx4966IVLE/HK8ZMulUznI/sYCkvDudH
AlmpDBW8cxbj3/ra37QtBJOi5BzyvAFQC0sF7oHBB8fQ3X+q0TV+W5q5r83XPfWW
SduJ46/irzJNWTLOUC7nxvUJJNsHZeJzhTy4Lr5q9RUPZAfwsPyaIPTBnHrRvpy1
/hi8tIYFnxymVTarC5e2HRZipQnN+7rrBSg63AYjn6On7b21fJNVJyEUD4V4gcfs
sVT1/HCLHwSeK2GSqYB3Kw8rHZcw9u27kHH1r2gWAZCM67Wm5Wc5hRQQFTzoc9xP
T54NAfy/vGJj+RTJEWBZKvzV78L1ycBPp6Dc/BWss8HUvFfGoSD5D3K3/s3I24um
TMKnMKgf54OE69H6KwdTs+d/P0BYRnUlcGzhuRN6IbsV6R7bz+ToUXOECIjtj8P+
yVod41djAJYkg9vhV/ZH3iWwOP3hVHddV55MeKitTGd6v0yWiHdtVFHGHQ0LrsL/
x3z/IQjbGsap5rP6cGxi8RsxVWPQ+eJ1zMmCPzpavMHssTreDiB5MdUB4S8K2Tox
rMsga0Cf7gasTtSL4BUadqzvHBmSqW5u3iUsHm4+If8QrmlJHVmrdhLICHexq7nR
JZmOZ3oHNOOOua3KNY0gUfXc6wluW7Oku1qmqIgzy5iCw2/NdX5mND+Ptf6sNF0k
LUJCLV3/lXOS7YefrX6y9jtOm2KRkGJU+KIvhTiTBmSB3J9lsuPvPVSTyS2foAhw
SpkLxZIAxFseoNnV+wiWNBTTcGDy/pBrGWqLBkT2EFbXy9DddpibnV+eZ9Dgjcck
YtzQHoMQdHj+7ZIFlIFTzGgMJ84t1PWlYYgTyX1S0uMy3vRusTM3mVa6kiwg/jpQ
qqn5QDSnCBs++QnfoIlv+haLsjmKxYsK19CUnq5XC3aP/OSWuGF4CORXyucT2LVw
2/MGyyKN4Et65WslP9OVYkd+c3DWF9QWogNzOes4/lKDgHcByMIBCAZo8S0emIT+
smDCEu7WhVBKibJSfLu0td7a9BgGH9tlBBO1bsz0qlaO8jY/Q54Ay0h0wQImKXh9
qD3e7ofgAHfZH3w85DglcLTVbiJRWTH9DUrxhtvaB9Hk5+JsXOUb9MtkkYwBikOS
Tccdd1366rMofd+wWbd24ymJCgOZ4sF6c42Bj4XaClFbOveb/gaWLI3PIXMDLU0U
/OpQU88dU83VXx7K0EouczSoOnra6upqEHIfHK+RKuZc5IPFSeFCeUImujeByiQ4
knF9rGFdULH9i/3EysvDcfiTYaH+zA3e+fwFwAERjvBUv+qvYyaVC6Rq8IBxTfKo
glj9X2aswSQjYp3XXM0gbVm8/bOyww7A6iNbTHw8Li0oiowxqJc0nW/qRaDGsQHE
hs8+bDdVHjFm0PFE7sbNPAX3Qxvol7eJvBBhvrKNZaRj8VC+/g4nS6b7HnirVoJe
Jb8Bz2x3EtRRaZ0A2zymxavd8e91DuYQtz44PSFIvFIduAbKEPu47YqEEs0/04E3
0VoQA9wsRbHs1uYOPCAkcESLf5e5kbffNBA8faMeP4vAhb9hepSqGjwVYFh6j20u
fo+EV8cVVldmWO16J5+JKGoBUM7h1X1oC2X7g3vSEzNFt4o+EtB9sAr27WQTS3T4
Uoa7uJe93nSUeHlFP/T7B3VLbfYTBcZy8LSPgAk+6EiZIvghrye29Eko5YByncqy
blrzo36CZ1zkbwleEsIF2399YUyC+DW2w/CEqe8iGFLoLz1E13NXWskspXh1R7gW
AmGfS329av+lCdbxquwnTH1U3RJFqtSn1SwYJQstRdIJX9F2Av53tPHFMV49s1e2
/Q0/Nh/jS/8I9chbIZKKXoMHFPs3PgJAQ563uJrdmmRISq65M6hqzk1nrwgEkjNo
VRjelH+bE2+8KAErfCTV2J7+kc/w9nSsaiopWHDi0yx7HtY0AJuyIl4kfiY8xeet
plDnVeG4k8yh8/wpknFgvKtqk0XP6KZ5uM5HiH0KdzjYmxXY65eZSLtAcRjITabj
Ofqw4eaela9EU18w6lQc+hy3K4Y/YRRyuCyV5PiT8nyIGeVxsjlIgCz7NyIjjdnu
oOyCXT5YrBqrvQ41anVYc1BVgPtESVxAF92N4FZ0S9KgMRV0UMKdSeGKrexmc1wj
NczsYNr0b6ara5jnKBF0O+v1tPkjvU8k9WUSnz+UpYM5TKkVJJ0vveFrBBkiX9Sh
pjb4ORayWQz1fcIJngB4BZWaH64sMnZPLXc9f7CtQRu4tVZ/8Rz2NMgEqEX9xOjr
uRnLNK/HD8pa2m4p5eUsCcujqCUstbjlCM071fRXawvRs0K+zuF8a9I+eYiSuT8C
w/Yo+61xQEqUdjAG8PmHqqizdh1SdDaNXEsZvtD5jy/ZdXfBmh5QKghU5xBlQhah
NSHIOqr4gtAkXfAgWyWxXRpcdPy/kh8MvgjzCRfc3G2tteCh3tnoeJEqgtVqHkHV
eoDRd2v52j35CXlbw/e3bUHYPuC6RPdvXY6ugbAfn1SqQDNWtxFBgHy3AWlmby1D
++76AaDdX5sKiMilBgiuacwAyOvZjg9yAG+BwrSBAQh5/R1olgj8l6KaOA0CeS/X
Wz8F5LZmrgV4lojcI6Yu964Jr/j4I/cCGGebopz0M5o9Qf8DeTRMy8CtD6l+TWDi
Qo+lQit+yJlXcSl6fv9paQuanzOXs4FkthDw8t+HETnoFUnfvEo9axSwLLM78Bch
RHmw5ui5zgSLsA7Zf0SiQF4Bn43SXryYrzQu4QtZJMnJ77vZOnV0tf38C9Wy6nNs
lQ2b/VNTyKcNSSyooKSxLfj4anbEyIEZY0SmoLAHwZdrmjD1tmWhkCEkUh297ps5
O+bB8bLFZTmGWJwkHIVai5y998ix2Gc/rBjlnEcwdAJ4ehAuwY5cM3HikxOM1p0q
xV6ACwhXieyITOLb7ioWmroYdnYj4dGF6Zag1/K8ajjKo+XVYvfqOBXd321JSrcl
Qr+qT0w6qA7Ly7Nr4kmQXluBGc/F/z8ejLQHiipRSTbsYsg0IsKnm/qwubjwqNOw
DH+8My3i4pBLRHBt/Sa30qzSRUEy1nefweU+16OE9GPh4yFqFDHfbMz+L7Sfk2Ci
d177tym+7D1RW3MyyLXu9YuToDC9W0G6HPUK9o16jmV07Xr871ZO+W8hxPviqgzo
8noGxoUsQHjZO1ODnIVJCGVjmbhvb+uqfbp1NwWbAOZPFkcq/Rl3lCU7mwNAItKz
aaMpP4sfbtBeRebyuf0ahQakujRvge/cm2gl3NX6xtqpcHLoDxu23hChbS/0pw5G
hO564vRVoSwYlm11Gvi8r9C0wtJgn4U730nADOSuqPrBfEAntg+1taacjSY02Hlk
h3cOp6ZVuuA6LmQC1b5uRE0EHJjMFNRs70LPfHHwPXh8SxKID2C9+1avK7l1SOaS
8utXdrqPGKsCEbn5uH8uXu786y2n6S0l9TZ0+5QJ5bxliLibOBjUscDiEaNz04r7
wNBSbRxIg7r6J3gsj6WJUZv4Vy335Ki/2Mpr3DQtkyW9BNW8ouiUcsinHzH6wM7k
xjQyzMW20lxninL4mBdaU5DJjn3AbK/mOfzHqVuV4X4Fcwb8HbFdBH/dm8tfnq7V
sPRW5NqjGexPKWdbVVtBJBMEDLXzti6G0RyTtQ8p1L8qZhfopjJz7Q5+UMntIUvr
3CyZDF+91lutWuIz07f/4Ub2lSSSRpMYcsdacYG/OkYpBrte4sqqMQVz3ndQ21Di
BT9wF+RdsshaKCYeu59UaDRLC5EJ1qzhig0Me9ITAg629KdqvzXn3lM2MEGznsM6
0UmkVnPKc0JuHTyKaUotqA27lFO4qcqQNMKobjJ9v8JimSgOiqgtAOnkpT4GdX64
66m0Vz5C7ufCyst61l4u4feqcTgv9rDCUS1zNQS6zk8YbjAk3hrFidzwTqSrhOu5
hNEBe85s9vYZ+ploJmo/GJBUnPmQTOP/3YUYzdMueEd+q9UD7o2yedS7vBMAFOO9
RNyrylrzwoTLGHh6+RPqngHedagi9fv3vwDJ26asx76SUeLSpaOQnDR4uubN/fdc
WTYJqPusBNyKGZerz4oRe8QOBlka4bj+zFcZJrWDTLrFlD+9q1E9QLLE5sXvwTvK
ljj7vIerAPw0U11Qif5JWClmMopw7KWuKUrM63FOLlPo5TYdSY3RCxCKmabV9cev
fob2t2BciMji9o/sMn4qH9Mu3ScZBDYmlFlDzQKfzM2IQcpsz+DFHt7+VNLrJf6R
p5vzMgL4328KyR0T4sHgdREEs14AsOcGOWSpA+C2lMsWAqE9g0URjvJ57EAsPbRs
hpmdcB4UKC5K7bpliyHuGhTTEqyHCcLYPCIXEd4KCP2e8zjalQOzdLvtPJX3vkMB
vHMeFlJnr4aBOslmfnPOf8a625vVr0LLqb6XuAbV1KVrt/zO8kCPDi2aeIwagihn
MSmiUoiQk1c1SOxlVGurJ277cjGjJ/Gww1mVtwV+GZO4UN5Fllx9VVdSGTySyRYm
5b0QDMKmAffS+/lxi3mlff34LCDfhFqVAO3IZ9o1PUpbQ3C+dX0yzezP35rsWwGd
ioI2eYNTplugKcjQvMQpSHIELeQghwjYCMaznMqVNYyfbAur1LQdhIGA4s7HmZQt
Z04rNP2Xg70HyI7DTQzMNCrQMb3R3NvTKt8nQoGeFnxRkm+QAh0+eZP8u3hJw1wo
Mf3D+fV4exZi8P9TSY7xedb1M5Ef8ng/D8NJt1kyZF+0pvd9tE8GrNgCr/FJD5dU
mC2IuhX7quF6zN5NIBssrfYYefSzKItSS0A5tTOGZZ6YCMtqr32m+IQLnXtW/fWv
0FVJAVTMzs7EF4ahojKonQP6JLrD0HYFY34jpDC4Z+FMLASBhjSeIqdUAKSBhy4K
+LxhcW38BmEzl5ddmrwafkOZHTAxSyxtth47wiReL2kz0IWDK38ltkbe5//kIS8a
hzKU5Y+CvLZrXdnwvnUv8b2+VOqrza3u+pvjSj5qz7gjwuxJ2wQtg2cS6Ny8k/yl
m/VILdacZAt2gBcrYZkYp8G8FWxfQ8majBb1JHoHvjxkdVPJd/rHhMKzsZqOMmho
sKMetZR0bT8F0Uc4l/OZ78GHuPEM0hyYJE+HoXTzuXP2ybE8xveFB4nDhXYmhWH0
uTQQgPMoZmn7X1UI/ObmgUrzfeVN69vAymfUnHdS88iKDtt+YbjNPrLne1LrasPR
zUlPQgg0ZYxQ5Cf+Tu9DCwaQvLe0hkMpWp9gDKF7ja08/fexgmod+SL8Qx8MH1m5
Cq3jbtxJh940Ar9XIDw9oZXwOlyKcGL33zyI5wmuPLA6Tg7NqjZqlXaTdnhfyB9v
CAOeCWY68Nj0dEMW6r9ZkjjsJ9+gtTM10kV7eq9gPMtR4gwufgB40ukfBL5zBKLR
hABYkVpMlndqF4wTt5De4To3pRcgwQgdSQjhM8Z0abYe1vJ8lA7NVcObxLmaUKI/
LXGh47vS2ww3gGuux7xGQAekxnb3+zg3izFipys8+NJSDtw5qTPWgEWhpyNqzBMD
uI/tSyT9Hgn0lfxOnHl5SBUzwyE5ubbwMmCsKaYv4EJ3CPjBdKze3IR1ICz2uAnM
3WUTisse+xPNTkmhnCZqsIfOjhjU/z+gVrqQ05MZSTPjk9lbiZal8Nsrys6zQWH/
JSJQr8aw72i6aqlTnhsmUQwCCsEvrwcsQ3XWtaU1ZggQqJwqGMlA9IdSobZF6d9K
BQGHsVZ822x4RISlFJ0OHZJmhM2oIXq4ZreUJZaKHlFNutuSkB4Pkc+uPQNF+jak
9/XKU7gZfm4ndfsfpU7e/+kvErBnMWOTeHlof/q70F5SP7b+akLolvLuwL6+sVe/
UwVkhZsxnOttkBfWYCYXhRJZuWax3BLqbhxlNd+wSBvl/ratfRWxf1PWAy0fKyos
WD+8y7bbhUKbzlElnHMSXjQcRIR2bf2mFdJACL83g50z6S+NEoTiNPjkeUop+IDB
T8EdF0lek8G2jqQktscDRUKVBNepM6gatvBZrGX9Nr9Ltaq/wa57fmIP1RZKVm0J
uV9UllwP+4HYws9PT/jDZttydP7atI0xDUjiFZLsYZPoB6KfOQLGtT2CfaqCd9Zg
A5x5xo2IkMdYaxnQ7lwff7gVswvApCtGmaXuKfDGzJnDDM741b+ZwMMnt0lEnO18
Na9tbdaSsG3a6HIAcgQ17iZlY6in8aqc8Fo8lH/4OSw+sWEvcnN8zCAZfGK4Nyaf
y0Ixp+8sEcOYXchACTPeWKXt2gi1Ica1Oy9mZKWAFL3gkdavcMzUKga7ivIZ/flq
eikHjVokFXfV3E8Gk9pMqa+N++XKFAl/1A+Eyo/fJDAKVkRP5ZpByp1oyV2/jNSW
kywGb3UWehwh3+E90JJQh3Vl0b6nSIoKJ4A3K+59JA7EYy1/tSZX+2HMADw4poKA
2oTVcxc+L5tV9a13v1XeQPe0Cin0W7D0nBONWB/k5GN48s1uSZLGWQpBsLq1bPfb
T0TGqZhZUtEG0BM2lbMjPn4O+zYqWiYl+A2R8SgqE2hWFQcM1QIWNJUgJWJ9QYMs
o+gzFVmpvSovj+kIIIvffZtOnb1Uu18DXd+SacUZj+BoXA7stsf//ubY3jXyjefY
VRwSW7f7yVV6jk7vv5vLuYTqLmABkfj3pmXmMijQmk9jTaDDgxwnmU03Ol0uMPXk
FJnYL0nTqMRa7Hd0OJVk4hb3E4WTATctrDdvvUz/FRM3obl5qZgxjVfeL0YxzJDT
uy5aku4hieix3qCv2/k4pFr9I0JjMoI34fvT3fvD4N2+uB/se8Xyv1JTIG8mqBhS
YRzWAjIvOvw5MCE6mDrt4qeebj3fT61iRxfbmO6qVB2c2tUVxyj50bcMKc2PjZl+
04ZATXdyKc2SEMY9nLtwSLjrUrENZVK3SVFTBuTz3179yH+pTNcHjTOX7M7uVnkX
tUX4Uh8SHjJ+EEU2H+LIhvmRU5b1SwRuqumzvSrsZ0cwSGl3ydhoSwp9CNqElbWZ
ecZo6Z8t6bfoy7ZR0aFt7AcvAN9wBdbkJZ2jvidsLv/9lvLVEdq+q3dcbUF/Ssyg
3f/Lc+7EM4Slr9PdFs4hddPc2dvDt1gLq61anCQ5Uh8Uit/+FNZuQFTwqEwSAGhg
383eY0Zdne43EjjfMqFNcZOxOWgpvEugnwBfNKJgAZ+Xe73DrB/+I1PSqYf+MwNZ
Wwk95E5dz5TXya07+qyNdGWCDJV/w5gBouP5KPxnCKTnYFY9/b2ckLetyhoN55+L
slbDGcH5K9rH70Sk6lbzSUExnjmY8wU78IQUdDvdHgSLa04jZq/BRtsLP/0P5Igb
By8KuPW6MTfHl4QrGi8ySnqkMUVBUrh4y83CnEZK2S/GKbGO7402EypvIRNWmd12
Rp8GOesrVbEz4/0kjeM6fXNNSRRhASa3r6dY5QUR0RemsDzORObjAnRbSCGCBLOS
8eLUhrHjIeJhKh0dXm+HIRA7mY6nHC+mG2RhovMhKKCn1lxEoHKOaZlz2HicIx7n
drdSvmfMJ2XNZCV3zHadKqKpJWdYfGCJAJ6kmqAmT6EVU7oaJWWfU2mXUvpaMyiS
NYYUCwsIhJgIEjgffXi0Cv5DlnhJrkG3PQKg6kFwAHJ39xZSV4vc93q9HWmR97c9
ZnEiPHqgIFXbA56scqlzNJD1eluBwCIVVXOy/oj1w/rslcZ6WHBW8psWiNlaHhJT
Ei/zodfUpwd/dEuiUWaF9FjOYNjC4Y8D3ELjTex36MMW+a9QZyybzn3HS3s9mDdJ
1PSv6tHiW7u63rIIGlGaM3wK0F1AsAUAf5ooPTA4MInwNCCkOV8R2YjrYqloIHG6
egLaYhxglG2sR5kPPDiNbuZEkFnwOzjTznn35gdRBw2/7WEYa1Gf6/CoVNsDrn4D
KkOec6S0ow6Qed+IL9h6Hrz8fQmJL8iQhxc8ErfxXcVSQriBxBPX1gvAW7suRqwd
8eh9n4Jr1iX/+zJCFnDWIBWswgC8+OD8s+vBKPJx6Hr2TYtj4ZQvGjTxLdqe1Wzv
mGW2TZAE9GlUkN0Y1hDyX8HxDqqpbJS6v3Gl20/n57vOULjqPypxNyiRH6w1OgEu
r2CDGgt+Febq+TrH8rYFaVCQ6urIgrwgRRB63egn4z4OEGPR7YkfD2ZykoZtIaqu
L8FR84Z98cVlll6IM2lDdQBaVFAFaX6CUCsNOIKlrD5JG0CDbvxi9O+BCUplclXg
tChy8M7O24F9q1vfGAxWK8HReVpfR2GzWjndRU7V2NGQHBkeIWdj4MjFrtErD5YV
sQx66cTIl6XZYzFNBGmgaIK/WB7FD6oJ+B+LVJBSrYgY+IaZpn6J2nm8G5wr28V2
ZPmSkJdPIqBJpwx3wCxl/rNWgFvC0gKtbrh83FvaHWd0qynhUhGlcQv3mRsqu9Uu
vGyS3AXYUmNLYvedLMYabmTuniLNwrA2/aHd8JLoBknvu4i6TkXvSGN2hw1wUeml
lU2Fuigrwl6VbYHyPie8A7QnnggcMmvxYlP76cyVixK+mdqo2BRgtqq3Q8fK2MYO
k5Y3wZAxzRsneQoNR7V1E+5BQmSDWMOtnVG9go7WAJ9FoRKjZAY2sv5L29K9BreJ
z4Sfti7mkjVJ6Dkh58jofRGHXZrzhjL2xmbQyRNoYZF1QWIfQM4dbyJy/0Zf/kGi
zsCZ11wBDHBk/zJXJulSsmGRZJZp5BjdfGVFe++q5mVoVTSNYBzCN7S28jYElbcy
ju7IdPs2Vj/io1Kc/vGAwZ+tE54EkBgHXWNoQQYtQLA7ChmribYX1xfif/pLhmad
weuAxsZpXD6HZ0YH7Nuytr7lhrFw8nOJe3vqgLAr6S5iiLvBmkRnAFqjNJsXAS4D
pgsIERCtfeLyw/J5SLQfRzsVUvbxx3RBuaJReXtNIGs9S4U21xLff2Fi9Nd+hGPR
lNz6W1bZKpAMiur1B0jUVgCugLpi0mY86lwWTzEYoubrFsAgsUjYgJGrWjbKyOSi
cuevcUUn5WMrIIwq/LrdtQtiHWZ1wSncCplgbz1AF15dMvvunTRJbR5uVOIFGAx4
GenPyUSS6lcBfT2PxN4xitbsglFnIc6XgnzjoqPwZqsrsuMfz7YYp5nxlvyAv0Kt
Pkmm0EyRLE30pwpm2/9SY+j5QdRyAumz2+GGRKg6wzn3BKBoP3IDYzpaf4zJ/v51
yKze8ALmLh6obMMMTv9IN75fKc1u/FoQoMolvJIzo13r5eUGJ8qZM77WKPRM+0mr
SVEZJwg+WYLElpC+R7L8P8jirosSHhDURBE2wxwCBQak2CujktotMZGIPVT+5LfN
j60IQos01Kr66xaLgECgtQpPvQDFu7E4IGd5iOTMyc9EBBdE+Pkz3wwx6NfeGfuU
TVovizjMb2joG77nLHZ4nQbOk/bYPq7eIUpYbTqPtUCosZQ+DTlX86rOFD5I1agf
8wIz4D8kybYog/gwhtrpISyzPuVnQxQS95mvaj2lofPzzX84euhBZFdWngx3Y3SZ
x9cD2KM7nUBynvQGxGm6ilDGpy58CWaAoDS17ueyBqz2waYEI8md++LhLzLe8ZT5
zkvyDTuk5dECt4GfeCuykpv8yU4ByTVpyhICw7/My3WQPvaIYQgLR4Rqy6Uf1uI1
GrZGTkkw89tzcWkM8KPYz5IvKW0GCkEYlq6MuDNtW67r15JEcFkmdAP/cEKQP8Mj
Fn9utNDHwqfjcsU4Y7oM6EcSoA/lQGjNkLCEF6deabGcbN8fzYoDHmwsM5gxFrZa
zQYtALGWdzdLs/mzfW2QtcTvTNEb06yJwFZ+7RqGfehvVFA7XaGvDKqinU/1uAF1
6i1EMiZ4tK5CDFESo4f5EATEqJx9ip0gqieT2Ur7bNGlUjmofdYxrDVGgG2RvIBM
j7UIxkLWwA4BRCq9nocRzktgYhrgqdDJKnpooqqCa5vuKI2QOQxCZbi9xEvxjAOu
gOOjMxgVqpZUFeagnwuvdNwFDp4x/m0vMz4bD5PNeMrsIB85xn1lHCKzt4lluQSK
rcpqpoAkQ0jzeHu1K4iuct2GTMegxqqrJhkWM10y95xqboKoCbiSW9YOToEbaFoD
BpGLAK8yX3+g2hrGS7XKwCywcsL4t5CsjTesC6Xu2fF3INB94wQyGWnO6C/YfIO9
r5FuvSt3MNua/7UHxgC7k05/ONvairuwzIJYePrmB8kPvItBQZTXml2o8nqhtk3t
yYgpf0ua/pmmNeBElpxrqytF3/wGJVvJCMiihlweRb8qjmBOGUsGIkmr6KMU8UiD
MIMCQTI8GqZeqj+Wr8UcZyoa+ge7fGA3GSlVvamSa9UWl3a68J0IVz9cm4PnZELw
LO/FO8AtllsJzr23SeQPpLnGseFeDUhruWdLj9E0KTLHq3L7agA2HSeo9wjcmrEt
bST7apsBhzIpGH6mR14uawsZu4ZWv0O5ESDAO3DlHCxqqx3OKEp1aQl418wTsQBA
ZECOPlvm9GVIaJ9DKkQA0Ly/7IhwnVuqbLa99PKOKtcI8mEreNJO0Vp9ypK872lo
tGM8g16E+6/u6E/xllewdCCZn5xOeAEAx7RaWFn9w1aEIOxN6OFgCI8JO+6xyK/W
7XOksekWB6VW/A6GSGb2fAirU9lHzXPQsKCCIsM8SOHZ/HbRJGTRUMa0mNI62aH7
e+wdSwhUEa/gVy6PC84ZVX/02C4b3zG9CS4BesvhlcjTK4kdbnzNElhEVqJq+YqC
VNV0lNN8opnWIKqIMNX8RMEz1qssktsfWsh18bDwvToc3zZDmyTZWoyVliUTkmZf
bFsBYTgXfmT4qVroVrnWyH5xIhkU0i4JtKAKzfn8gUhCOqcNI6/m0BKuim21P+Mm
efR95Lv3+phWRWd1gpcnJSNE/d4Wua3OevdcvmtTgDAK9TNTP1V520MOYgYJIUpB
56DO+NHS0P/d4fFyWbhsPiVSQMmsxpgZOBj7ep3njx1kcLyi/4KDPiIRjaQr3tJR
DC8tgVGAstHq6VDqKaZzBHubTSaHTFcKNU/isVBmSfi8wEjYYzqXZmRQZVQsu/uD
jtL2vSgIF5FCHuQTM5OphlVjEGxlf8x1wNK45jZrtfONkhoxqXRRmNFOmSjynGXh
Vu/Prmn5q+0XnAucUjsK+bUSXRD0fA2EF1tsSaf7tCo0pIQiOBMww9mCELDK0QWj
tDm2/Gjs/ImGmgpOFxz05wh2/0KvUmCqpN4+0YPhPrMEJyjNBxhJZfjjhEOXWyrw
9cyjjhLforM/p8eSINUNKV7U5lYrxsvmCwpTcmftDjcSVc3fgFhiwxePYazc5UFI
zf147n1Tth2B0thC2VMNthw4ez8AJx6FJp++kO4j9ZLBZwpjl9QwDeKoUL6zqJa5
9xmmZe46PGKBGEyqjQpzuRm9KdgUN7JC1GxHtLmqx+XLj2IkqdzctDGNtuNnJfbl
Hv+QLIW3pehggKwy4XF8cSV7fzLbcuCm8CRpf6kFq/hMpjvOkryEBWjJ9Qnuk9JN
/auYw5sVsCm4OViC6VNtbYBzL6FM3gNlBX7p+PVDeiJRoamSPDs0F6VHvESezt5w
F1aa4XLo7Nt2p5wKJ7VSsyYS0COzFyYz1/bPk+GTHu83JFyyZFlhyC2DUx9g2JY1
iL0he3K1qOBsisKXTsm/3X83/Zaxg2OMlhjS/IUSxa1O12cea0ZX89Kb0d4dJyWS
fm6XuQ3TLzgX01hLcc+XBJAQSenTVDd/EeZH9aAM/uSYg9wvm5BaxQw5n5iRJ5j3
lo9bGLvwlUs5scrPwEwKoIZttKXbTK6d/I7SKzPijO+2OOzX9OeosAYfZNHzcGcR
MmCrEvQEqcjvQSF5MtPQFl3BlkwojMfk5W2Hfn6Fi7yAqE9UEGSYXfYTRllDWmKx
GNlxZWxAwLhOmFxv5HTS5iQ81Qjj264YXL3kLvgZtsc1HkPQ41ZUcbQgoYE89SWx
+MAEYwXCNyc5m3saEJdAIzx+8npAeo/RAal41rdkOgO7//Pz53n6HgsQFkn48sjH
q9+r2u5RtdusHyZn6IqQFE5j9hxGSzQSWreTEs8nASuzc/ZVU/qVSa0jSzAQdCA9
5NPi05Co154j8Sv3dY+yOHGON5DLbHKtIRl7qFFIWph/NwOGHv53cE6HvA2h5vtd
5Dq4L+BKMYDWHVipHpp64vRBm8/6Met9+OBVtxl+GCf5OutmAleVfU3wqClyg/fc
xkIB+gsNJveAzQiaXUQLufvSUqObjuPvXlNBzOb6cxo1NKnImX9bXl1RIQswRSdn
GuyGYlbisVWX9U2l8l3w7OxKlehbtbkQHat6caG4KKx8tozygbnpo6EU5BmAmzzw
9LhvYUfhy6YEKRn1GVEFGVo3GAh1Q75ooaS9lTdvdJAhruYRbXpvvW311P3TuLNI
0M5SyuZtRu9uHHjSeihshN6XuqkY+4cNqnI/u2yk5Y6xHleG0UDIKYBZmGJjvfXY
bka3VCOFLpRELFflaKr3CTouN8Xq7XZGukCUVtn7hbMYia3z5BzkCpjG0s4Q3QDh
XcjUKIMehdGx81LuclZ/mFhsipfGOjodGWSSJLhpa+gkLPrCSrKzXPOZep6DJVet
chu8dF1sapXsUDJWqWnGaTNc4mKzfP/Jx+MqNk8m7UEPqxC+/SFAqJWfIeldNybE
RAim/m6l1estGEmtiBrYymaoLcw9kmQQVuaE1EddNDg/oLoSEDqK1jvH+OwXAQSL
aA/KvO44bdqko0WApKe+bnxK0zK70sKq5nJ0QxZ6L/bygSk1dzRENH5F5V/173LW
MbAea74UGDDs0rKE8q1YmPZLlpF27Ovi/P06veeoG9Dr1/qdrK3PclMELaJ7ZQsa
NS4akiB1fQK2LeMWTlpHXRbMWTzmWYD6rUxl6Gg6hKgagLa+YPMfKNy5Gk/kGRv2
9KHthfyO7XY/dLBmDDfV2N4jZk9Tm3ZiBOLZsmHDeiKfPYe6/R/gJmUuFexR8Dij
+FWnGGx0QsfrgQJeQXYTPFAiIhw2LndJ2xLj2goaB5piWhAQQBSoTk2aXCYdMIVy
QbaR1HIxKLjD0RVPkbt64ia3VVUUa3e+kYOfuBZ2F84+rD/PZLgV+6iogc72CKsd
EMmaIJObiJPdwEfPJNNKdKwusaMllaSPhe7ez5RV2i2e5wg4ggGodVxh4FC/TIVj
1JgdUdW6JrzwvYpGmvl7xByxQgR9Co2H9ETjt+nVZbczAGrN5Y3kVqMIsP6SXw2N
O5cF2efHPHo7W0URjNoYsnjfl9QN36h3o3KtrJ3K+lhUn99HZIcfeTX4/wKEKQaL
ZDJfRtDrE/SYy0IaHqju7YK/SacHedoidSY0WVezf6Pv6I5e+0XQTr6RuDSpklkK
3uhvSF057oruRpWqyshIDqqHsZkvUknt7GZ1rzkCkO9OgTeuySnghg9xjjrUVfP9
MmDv52g/9OtTDyUvKAMDvCq+RUo6qL4gWowwJfrwGezj70rhemBkQ7Yo7PA9enpZ
UCEKr01JIoIzn0XFCKqP782uleTOyXlPLFBCJj9w/vdii63jqO2GVadGigAy3JEH
BBskfuceg79BGE3QLDI0zlVvmBsIkGGHz65e+w5PMVM2QeGfRcTk+7ZZwjj6oPQV
HflJKseXbef8pk174F1Kf5O0rvzXyBpKwhqwqVlOqAdFXqJM6znZaE42MKW/Gzu5
FMl0W6KWo2P1eSC3Efcw+/t5G5IuW4eEH6lXdS0Yob9m6fxiraF62QogmME8aayE
KNZRmsjgnb9kvLZaxpcyYR/CGw38PAQxtr0OxfKKRRnRMxzA0b7dL4F+Jf86RgkB
3OzNfYDWkb4cg9jCGgscpv2w2M7PKaCCCtFqxYrgmx7TMXMvgeJk+fugperGYckX
z671lAPDA439cvhEm86sC8Qpg1tPoAxZdrRDbYaG3a7V63AFT2cAPFPU7wurOpEp
PXWv/hV9aZ7H1nGXn4bpyA236i8K8m12jiBtSCgQdKs19sRj4n2EgtPwTw7N4eU1
29pUmkbHDYzDVx6M02i+cb3/9ikoZ0ndGNGuHQOKouznVfCdPGUvJOLtkEjE3Y9q
gJMpQDeFvcBG3xjPA5jLCdOyGsl4f4dx9LFMD1Wg0iu//Qh+n0/ME/EfERucirZD
FhqgVJ3/Xl2d2F7LYrR5dnMjqdzvP0CmPesNv37sW2hSLcwXCKXJJ1RGK5QyizHH
jXFhiCCF79Fy+T7DbKGHJeDpTISVKb7B8XpsXRr8bfLNSxq0vQTc/pii8fnrl1xm
i/yGSigEbXFSmPAsw8espYpxYU+VxlkElMtrdPQ4RC5gmEmbooXJ51izV1G8PYhP
YrI+bvd4ihLqduMtrYKXrPcxmmccNBMYbxHyBtTbdb4PutuKdhZvVh85w2Y48I/w
E8YohQFVmbVi/B5U5h23akCfl2ysmR2GMn9cAOWn7aTU1xnr+9aSSNIGDX31Xd4k
SCxQu0Kpkzys/ulqbcZneGdV6qlEhmsbBLGmX+lqTUZuc7cj4+H1J9IrOhhXXwR5
3pis/F9l9c2RB05wMwPPDueWUH+DbHKCpt+AT8fOdLwJaz0opfHFKnu3tVpEAFXU
5KDJc0tVIEfD5eUMqVtHp1D+BVAUHBFZ+L43n4IkEx5C8JfUXLqkONXxWwD/KNLK
a+V/GA0/v15r0XOqOdSvX4w51PcysqVhvisPvybe8ltSyr0vAS3g04dDDxEyMr+b
fIfeZsMgCwnJhnVvPrfzK4j4UM+C5rbyi4/yZW2TPP9JYPqSR994Ou8Q5WJroZYv
SfqFFtBt+1yOICYXCB/LLE21B/mE3cByuXmOfbVf3E4Y5/Aznh1aX+XGj4jqZJoR
01oX+TaPfWkxrY7di3iDFgH9daiMsJsxWP7FTXXHtMHASDHZgUVDTYuBzb6GGdJh
yA6Ep9F/MGCb1ZXlI4hdIInkNEvStpLbz5YBUvd4lMXNu6o8JKQPiFR74mDVNgny
9l+9s2N1ByhUohlag8G20DiAdckMGPXIDY6+6LAI+yFiAiqcjuJ9cFQZQoWHIWrq
9xUjymKlp4itgN1ObkzIBMQLuiTbNsw9mWlRA+1IvW0xaUr/CM/TUDFLWhr3OfBA
GeyFhmERvaVW1WF7JH4uj0tu7VxuCGGqak69+mXCS+hmThHdOaQ8v6DdG2d12+2s
fZfSjVhZxV2Y/fzQG23f+9CuC9AG35SaDJh0RuECikQvXk/n8qi2TVG2MfP3RE8e
HJmVUkpDKS1mrbkhgV+aJxqjPVDCSk6hlpJgPC3efcsSbVbcIfllI/5DqdBQPxZY
zK3FMlYgaDpXtAY0U4YjKiBkMu2q9XM4zp2h8ojQzvq+LdeL8TJWy3cgFA6CHV2E
M/QFqU8+miZ2BVdxn9YvJEX8rCKdap9c/5ZoYvn0Q/QeZGZOlsrKi3iOwBSpF/Nn
nW40Qvdk3alVntB6G84TAEchSp7yKo3DYllLOYRVqLjQz9hVu+3zix0Iq01ytupf
eTlqZ27sTE4qUjNAKPsEczmP8JfeHYaJZGEyFWIm6sdSlT247E8chYn0V3BIfQ1j
o518IsjWs0WZB0EF0n5X5bE8mxlQkKkW8M1KsB0PMcuNNPZlmrnXoV+Ew0J2mwf5
YOaRacqlKFL/SPnoIEBbfgTT4j8yvgMjApLOaXTIawEp9XAWsxmBML8qf2pdWGgW
CllYrw338kMAYhZgVSTUdamoyq/AZXPkbxPWlfDd4ZHGDTEQXvFaKt3u7uP1rX5O
5uKmfXAmslAZJGB+k1TRCKiVgaeEet1Nfqb25gNoHEyzEwMkfqTgXXIsfUFqNH35
gpBBjQKwJigpIPEym0ndRRANGY1CadIhw/RrKCXJ3Woily2bFVBMb7Cew1j5n4KA
c75Lw87CLss/F8sGl6mOGYvIeom4xylwy559RxCvC5HbharNJ4Jxz+ckEu5AbZlg
5A3KpwmdnZypo/UWb/IiyjPpXZuBm79rkdcBy3FKZ6EFzGMLoV0VW7YvE4iTq21a
M+Hf1l2Xz0ZZlmmh80WLdSpS5gwvAxHVl4g7eXtvfAynGiFEz8lIR58wHgsmGYJm
NiwC4vLd++dDCjayZaxeINVmyJVObwnsY9fqfuIarmKNTDMuO1F/tj+lUGeKtQjw
CqbWJuDK11hU9/40k+nc01RkukjGsj17JIzlIJ3IhHKKrhb4MCQDTnRxxgmSP1l+
l22OxOnyUe7D9k3U1l9xejPhZUXpjf8NveYAcaxxCmBD2pMZyhmK2iq5imd2rEv8
Eqrqb5hZMMQhMU+Zo+RlkWnw7O46saAJzR3Vh4fL2JAWf1c0ecgywzRC8FKwQCU5
5Cd6sqyAmbMbkEq+kzvFEUQwLrQo8tTmBAc6KhOxX8zUk7D/6lXUdoF6BKTihVpI
V0yNnvphcyvKgFWwSjM7gHpPs0LzGuzia+UgeiF7LJSxcKWcSSzzUBTZB0OHINyw
V/CWceW9b5OoeWmIfwhC2xuSWnvjVJ0fPyYZRF5mPIGCn35pOQGF4T5Pm2hLQOoa
UAdP3lNERFilLL5qsz+BGVRE5S3UI/apt83c8Nd3yDYNSi+68jf6TbPvY4IMZvKC
jIDEKUZb5oM2BicyqPavteZP9UI3P05sgpvL4cZ0UfS+L+MHrimtUYgX6gS6Xrxd
rdsAkziG7apqFm6/Qs6cKhH/zQEepQ35/QhVFh16Ppop5CtN5V7NaDWo3uqB5/bM
F7Di9zTg9m/uC9tdCOvTpNEX3jLi+i/xd+rPFVjt5+pcx6KpP1KYXyCKwXZ89YOd
ReUT/FnFhINeuHgKoDvXiQp5GfM6+1VIwr/W3R/XClGvGc7yEozTXraVn/jVi0Vq
UgrTSn0PBBcwqvuaVr1mLQDW0l5ZcAXrGJpzhSgPBO8Pmmc/omLgXXqAhXcxPX50
J/bztgd3vcuKQT0LF5zds1a8EjLvHQFDgWPRff/meeamNcgQUMRkVWgFr3ZF+pma
b1FlC1fu6REc62HWceBxyBsrUoAtwM6MntiIXKihDEQhzDCqmp0xob3WnIpiZdTn
IiJAURx0/D9VVSSyWi4VwlMLWss4gYocvQh1TAbJqBQvMnSscXQ3a7Kv0525rG4f
oFqUxKLdIcJew/g5iqCh/QmIgz9opVeX8sYhFdIH97VnE9vb0xfEpL7EXXZF2aA5
IFLI5asUap7VPFP8ELxe29Rf8MAA/9oAxTU57QQQrqVGrrbLL6cIygX4sW9Q6phE
Ty9XJ89WEpTX1S/W6jEm29cZ9ol0Ss+irn1i1aNjJREzQpXaUrt0pNKSqbNh0wzc
6b6zOC9qyZ6NbdxjGPj8Xk4CfCQeQ21iQt+lVjDtpKd2b/YhPFM3Jv7QA+mg4sCW
qDj1vVhmIKshorWtggpwaXbNEsvk+PI+DT4AMQRTBeuoylt8VcK32EFYkx3qz+Ff
vzt84y60Un3XtaxcBoLOQ/d8xHKfFXUiepdpvACV+5cY/2kpbhJ+blTZnE4P3ciH
3rsTeAteviz2VbCPXIZaZ+W0TnRFAc3Rq+6iKjpLDjuDuIlj8eRjGr0ql72yvPL4
HmjImb1pIeJrYFxCuUiGkZiaqg9EYZSnHXHo6tkfj4K0GxY4A0U7hetQoi1hDgjw
V4eV7c2PO3+2dlKVnLC/0mRQROk79KU2968GnHmB0McEQmhFS1muldAqFG8LGKSA
IlkdrCfKu6quOFj0JvhID23cYPWhmFEU9ALD7YTHPpZqaWC2wpi+lIAGCkfdaPiZ
vCZOjIVtH0aSThhFP28NISzCEvOhMDT6N4TLhDrr42RzYtlRWyviLlHCLUL7pJGM
+54GKm3nRN8haVyJpQl/zxaDBbKRH5gOt9M5uZDCsc5Q6p4aw77i8y0vvz3QMIxN
5cYWxqrxZ65hJ89p5gCWkUrZmmrWev9pSLXmcbzsIDQq2suj0/kA7EGSUpAqayTG
0n7oa1iBjxPl0T4ay7djyRcodZE/MdDf7r+WZ9298wiXxhkw7x3xbE5fops5Bh5n
sleH6hlPL3zHzeWhfke4LslJQoiRB5smbG1FNqVa0BG3j+Bwha4I6GTiUrEIjZZ8
vvSo/L0modijf/WP3NXssi7152qQTDePge6NCnhL0U8Wo4sBIkHAjEFl7EkyqQsE
F7/AS7W3y/REq3W6IH0w0QW6n/PD5tWsyrpfYxqfK3+0uMuo02Wry149dRdGkgOL
d6/KvSgc0EBaA3SvRltLAO4PjZRNuCAIbRrjFpdCgdJriIAena354Sd4SZv/dnvb
M36gWqn2siTyEtW8/iyqyr1lxSxu1+jakbI/4Jx7OuQz1KH/ytcdt0De2IjLV8f0
2zFYM1jNwb6oyV4EygApkLASppwqTVhwS8r4StUaUaRFmYupCtvQGTzdWTCfIfcl
GyUcVmy5BVPpfhNgYO7Q+gQ6UXsF63BVj4pxOglTCk+6yhzGfYegj+AsJEpn+8i3
uiUAQKJS8WA7RmuYXyEjKFXCllPCox9MsTLLMYSEu0aRibyEK6qbdELVI+jw6p9p
g5j339tL4zlPiyEcGAn4qVox3BxYKvbMRqIy1y6RWTS03Ke72SDfLv6IQYpCg7E0
vNqUmQI7ATPcJsfO33Nn2XdexGjAwQ9mwMhNdc07XCqv9oSJ5PJo7hnU1vRwlVXU
dm0YNiJewi8duxmduuFlYsjFmIWx8qfgB39YvtKOAU4rNgYds2KPhfF1mdbg7wpY
DSvEXqaK0OA+y+QIWMnlzHiHujkNQeYKyf8aWV9PHDgeuYClmW43wNApFRbE6i8u
lxd9IhFQrr6Oq6aPt4j6UQDyWRhagPuH6/Q7Kw3ziUQ/O981T2wg5iEyWXBIGYao
qohnWQW8bH9yNxY4JyobmW5IQYBCryALFD21o2u305sm4y4ikmHxqhFOnTJHmZJw
VkNFnLamiORP6N3UmZu2+3XwvUx6j/2QrgWk4JePXFwkn/zf0UVlvz1Q/wxIKxA+
RaqIeLxfzli8OzhWTjiXku/yK7V8z8A0pT5Q4Se9zo8i418tCmo6lhO+qXHDfH84
3d2hiVoOpYLNxRf7MGYZX1G7zP/bKBWiPmRSOFJ83Vpt2pWejqNWhRo5TU4XwuAW
fIf5t5A90Yyow0Fehvl6vHp8dXUWPXK6H1rlF1zUz6vJNVpQbt1exyo5RC1IZD71
i7PdhWbMalTvUkZdr0OigxXS63BNvgeabII9jeL3tidD8/tsFoW4FShJh1Poqyk7
duRXl9Iq5WfKibhAMOi4WyN1KTa7NJ7A7g9DHfFQQ6WzEDDbc4eY6sm6l1/AMgwf
tEn59kv0C1cTbCcYaDTq6VxCIT5aoH/2Da3MVWrFwuM13SW/Az2sGiKU6oDtYv1c
5hOgN+eS/oKJCocuVT0G/8lB8Tgo0/fvIltre1XG/UWOe4cRsMzQt1tcDa0t+ur/
7YMC0bDyl0TF2X8q8DC27EEtIQZrlctKrtaju6y8PhQdtATZPFLxNplHqq4C0nLC
+v/Ccc9zr9ze3AXBRF0omD5bBPYlHNQVwcl+zbyhVQLhld/r15OzkJxsD0dmpsxP
ejQwCcB+pHgGMYDF37bDqXx8OBIJMjns5NaW1cb372ZnpO+rtnNTVvCXjmrl0oNG
q5v9fHOMfJmBfRtunVInNSUsLihTlEL8ZAGrc/GvHKV8xp8YsxS9RQbWweGG2j+y
EKe/wAscQMhcbv2I5qpo7vp/WkBj8vhlHgYmarCeB3iIrKWdOpi8M4wvBULXtP0X
RTGrHTW6kE0wqppz3d/2ZGnEMcosamnw5ImuodjZ08qhxyNZiyOLH/CmMVjoSmzD
5LTldaMA2dzEIUJwNxofsmDxGwesgOTfthbc2f4TvGMo5hf1KYVFQzTleAb6dvVb
e3wbAu1o6GZHXLKfICrnMpqhHXdMQYgdAL+IvyIFnt9vjsQWWZeuBXJ7mIy5g5Se
rrFBcDfPVrS9ufea2SwVqQfvSKzZzp2pXFhKejo+UySnrG76glS0F2t1zAG5rx91
2ai+IMI8i2ySs7SGU7Bp3OU4kXFqVgH50XbPHL2cMougscAFLNBDAb0LI7s1C2Rw
RrePsvEQC0nSFauf63AMFezRaJnwsn3ztG8BszXx1m04zDmgvMS6kNQjbwLtZ9pA
KNjGZORg9oG0m7msGQnEBQmHbd+irQNCoa4MctSh4vJ7vIjiiFNOMAyz0v8CRSW/
SdyzetKlv1s0FerTIghz+e71fbcZfJGaRT/okpGjN3gACWHC8G2o4ImePN/d6VZZ
5D/UEmZ3mqRZf1610/YTSExuBedMvlNjaprLkBNDqzjhkomDD6VZo7zmiy5l0DSB
/D9R4Grm7umn2tl1zYdPUM6vPdE2tOgnkvU20U3xyVHpi8vqi5+u5iXkk/Do8AEf
HTbd/Pdyiu4FVV/p1Kfnaz1uUibOuaq6tVGY7jGIwNgDTHQ/2SGw2CNyz433K4XU
LwV8VNAFTbxrDBg8op/n6uew37yBu0iluQH+GrxR5uhLrX8W4fVrG9n4qXkn++X8
VNk0G16mi/9GCD/Lr90AD6MZ7HS0jTKYuxAuvf2W/eFrIK7g3A0hf3Sl9THvTrz3
D/ZZr3JOekMZz94+3CNTLWXgRTAK0uWv20lkKz9oqS5yrJIxpls6fpYDrXgEBLzm
tzF1T2fc+F5VYkoC5ZXWrExreUmNavJBjxinSOBcoGW9OTkGx5zhQhqMfXjrKy0O
JgON2HjLYrIXnmCAJgAhl7D61K3Va0YdBG9dFC7oLy4Em+Ewvxqvdd9thDoli517
a7xHDILT1vx01JbmkH9wwYI02NcLvb0OX1kd0msBQ5e5xwjpcFmG+si30SLparNT
6WVhgtkxdzR83THMosxcudNZtnZWcqd7eQJSGGbyMavBF/NYR5l6/9Xdxm2kb4V9
H0GI+WhDiMwmbps/qJ+X4XasLNCxTYA0JHZIjMMpcS9KD1uKDCn8yK3t0StKtdUC
2bLCdZXnnCqjoY8YZyg7uArCxRP3vYOGJoyjmqWRgoWtw4C9rEMAtxirJ1+LaT0J
W1qD7eS6A5aGZij1ttbyzTLTYhzT21w/Z/osfsrP2DNLrTUAafMcW7mgQMYTxYbN
/g7j7gMm8oEXjpk4aEIoVkxjOaoRABCdPfbMPzvoIew6rwCv0sc07oypFW7VjoHy
dh0L1dvkldGQo6Gp6TCaud7VcNU+honfERL4R+DcK6ndSz0YUyvumxKoMivYE3RU
ytqj4/5eqGc4RljkMeqAMGA/EUFa7WbwgLiQfkREePzdMJ8EmddQYZOQH4JOy9RI
tz88fNh9RgbjtRO3HzpfQY32FF0zyuw71KC7mgYOyoyXBN58o/PRU4f8mhFUqupK
eX1I2t8Mq20MjhQ12ShuuGteDl96td14b6OreifzoZKewy+37h/CUbm0Oa4mYWZA
9BV7+WyOdKFxXxCi7l1zVCM9/H9WOsI/vHhIwP3oTLwISMhQxGycdqoe/mqZW/HX
2IutB68Ai4cyXUAGnEUUkKj4laFTKWopvYdDMPV+SNyWtuT7Y7pvN75oK6Ze2BQT
ZZAQuxNvc/2X4p1D5QaIafSMPjoLZ+Quegpeb74IsLkC4R+q3dbTnyHYaGXKH/Kq
V9lWSgPRLm+WkGvXBeahf4EbX9FW7/JnyoFnq7tr2D7BkrxhOn70pQkwCvsCV3Ql
LV1ikSQws5keXGpmRZsqpWI1S9OVVgnKfLttYoHPTBZhBXt/FqDedJO8yAi3Z3/Z
cCoJG8W81o9hPvJ1biH7Jk0NGrV+h3W2qgfayGK2Ljz65YfKW166cmKrInn929xu
2XZdJV7RDN/N+C5rjxywWTMFJ1xQoi4hoSQBYF0hqkSRRFLGf+fHe8D1UFNTx2/9
RFuUhO8Styu917nnEgh42W6sphzNhErVvWD2mABPOOJEb9X8Gt4LtyhPy1QArVbW
t7rncEaL0qEaMrU/ZR8SpR/pXA0vS/6Pjpcg1QtTvJcKJV4O7FalLY7FMPgOzJnl
MAzXfZHMUL6d/GDHphtEJSxweAwjTyKNdjjWJuR6P4XBWVMUsjzUAzen1uojol+V
xzEWS8ep/NjQ6/fi/W6WYkK+kI0DR+eFz9873gw4GxzlTaeMDjSmTh8trGojD1or
pCsx4pm39j1E+qH9evhNZyBWDp5wo+QsTO/Kz6xDaG2+8pIms0RTtQ+BFWUfDYY2
xRgz4/WNyC2NA2JwwiGpWUkPZCUsKZdArQlGWtRRt2qKIKPfVeZVAEg9vLRZ2kIq
H1SctDd7CNAY7PaFjdHTxWvXANxodAJnMFNxl/pKaSMEMqC6t6hKKz8c86lvyVlZ
hk+uRUjK6L8DaYCowSHOCHwXxWFT4YtQSPlCBjytHZhpU+gVbUQL1KWQKy3VAz1h
WxmONlYNdST4BGq4QOfh9UT8PIewMGwUwSa7BNMcLoQFSbfCqBUwg5NvwmbRfltm
Jx0U3WwWwtbT3N2L5zm2ixwXnk/bJVyP7lNqJp5QLx8L9u/ur/LBd97L4xTTOafx
MKQ+TVtROXj+tQQpmFW26zhjxKpeCkv1noj5hidSHBLLjlSLqYN3ns5SULj8LvzO
4QOzWYs1G5CgWWH5iHTJCR9HbiUg8i/loOD7+TG+J91c1NHDn4xDgqPsFtUJntec
IfdV1nhOJkuJfVd228TTx8VI6K8cCdDX7fnhRprw2016MdO6W5p1M2G3S6kBTIij
rT7dC09XuPhwH8fLxfgMxGRzmPn6l1uVQlp99Gzsv6yAXXW4YNFDIeZLhSPFLgOT
SQBeyDGAFxEPEFEYo8QBE5kYNQhk11lHvYk+HjvUmfbc3nFbMrxbZEW0zH5Cut5L
d0o4YHII3GYS4Woi0eRFlxe7wB2VgAvs35WAQzTytpY24ldhdtLG2ek8LSw32IqH
MKrbzMy9Lrq78p9bxWn5Fngc6BJJilB9Doh34Iwueam6OxdYGIlUMfQEPWlaIUdP
2HBJfy5UT446jWb7bMCn5iHn3nN19FhjcrwPJsTz0dGL0ggOxpE0fBHG277pGtyH
NKN2IidMGDifrhP0Qt8VDMTFTsv7RCS6NFV5kO0EEPDY2VWQQ/W9AgEIeJIvBOzB
mhd+98ze8OgywoFBBC1nsWMutgnnYYR5/QXhYVe2cMWQhq4NqUJR/tvtm8v+HpsC
KGY2AIl4vJnGP129trKCKHiMdlUiu5/J18bnnUJ8XWJhyHmx4Yqll4V3c3NIA28q
x6t31LsSdYChRa/FCRNwyP+4vD+9fpMYNaFq4Yk7c8KJQBRroq1X4vUitUBoy5by
WXmeqnFGgjwEnAsJh4WrO+R0YcdbwFr/1KkauFrNYVd7nDV6TZV4wHIa1AmfSyEs
WXQmoiK2OWumbC/0dR9JS25AIiBdOwQshIQxZQZj2pYGWeOd6IAs/xPRtlF0KPNx
2I3V7c/LTXw/qcbEZb5AnSBMnhsfyyafNs2nDyPm1+63dg3BOQEowatksvt4zKJx
e0w8vzeL1eEtt+Ofdpg7avmbnD8/3IFIKMkWL81hPldnBVEqJekSl752Sb+PVli/
rQGDkFsEa6tZPRqtYgzy22yKPifK1xETfHqIqA8pg8/bMzqnhW1RziBzN03qor6c
nsjrIMWmYatGba+/L+5dOZKaHZLIe2rUfLJMvPO/8wk0GrsdzyFugYrDMJHfMH0K
7GUmztKKbOJw0AjDWZv44HKz5Mj9F4b+Cjr84pUEVSiYsPp0d2qUQDchBQ9tRsjx
F4DSpJo+1aYkC9tL3C+9ztyvrDL2pIqL7Uhb23cvRBboalg0PxE1v5JRGKqq4hJk
ItjpdebefBTBFwFCMAUn0yhULl3yAgAPlhD2hj8q1gScGqH8V0b3XJQUSXWVnr2h
P78YaCTWnq5XkD6FTA/q8IWr3Oyxg4p0ffkjFSLNlviKbNrcsD4ZxhIMmgvFAMRN
D7d1XRx5xFLoJsxk5PIfFQoVUISfvvb2fskjoWruc3Pf7JHHz76fJuU9Rg6D6/cq
wJxcao0wo9wON2gNTcwgjxztAKlNoCdqE8Pfzh7HmS07xZeOsBZXyuP4nIDgyUvn
4vnIo5hwO/zV2OtBrTTr4BabcelNLB6S1MqivnMpyzyKewTvZ08QxDhYUYsmNH2R
nBUSZpoIQoIDHBTLzx5YCdT2fcZvF5BJjOi1fjSt1034hR8wD2/rado+YEiV48o8
lYbF/Hp9wcF0zCS4Et+X25SizLzGUJetiqmv7+33TCh7+Md14oKugUTJk8ronYn4
XDP0ZqNTYJ9HYJm2rII7ZrMHpX80YOP3OGbcZwamxzotoNJLZdelTXSATdaoPUvD
ezILqJO9RJ1Oqrl/BL+eMUvtX6aoxM3L9W8TnUrzFMcW8vXU4e4QCepQsVYh0UxY
RNr0XRxnE3MDcrDgMN3hjDvfR5UiwrKh7F0l/Tp2HtK05KlkgANEz1k6kqiU+0Vn
25qE7Div2Iu3hA5e5f7HvE6dkwf030bBS4VOX1yTd0Rf747hsNXBEWWM6E0UGQEe
0nUNDaY4tT/Q8Lr4Y7eAfxCzPdxCRRhava6Yv7AE2GOEbxBtK9mSAud0qLY47Fnv
4tyUpeG0FzPo8OXfWlMgWu4bmwZ+OXQmaPd6F1UfjvUprDBixmTfcCJoQo9N/Z+o
PTLzu1WZdAVNG8sXxpv1PnCEETk9tM1a4z4Crxcl1DAqa2q+ZaOZx1h8IjVu/4F7
O+xyX0q0HcyFR1p5igE1Yu1KkGxUEuQUQ6LKGPVEU56l3Ok7z17kgiZNrzc34MWY
uPwlykSgxYY1ABs/DvLwsAvrK+9K8daXRdmnNlnnUhkW8rXDAb2eBloPyRHkSdgs
XCizwBOQkvFj9hNe8g7rvbFhrsJl5nhCY/Ds3plNl8/Cf2Zm/Ll/U5u29FiUZ7DG
dFSJypW+sJxv02r8peDBGvTzVOlHyGRbA3NFpBfn1uLEy7907U95QIybg/b8AiET
/ZJJoMgUo2LFcBIK7dIMJ32JI8qtAoY+UYzTJHgJuE8ZsctLCff4xJY7unMgQThH
RPJJV/L/UIYWHf+BHUjEsIly6YBcau8zxAvh81pNjt+m7dnGzcCIPYq2jXZC5UYf
ctnkaCczDkFKCTK9VCq+9HGScCiwbHA9AamsJ7sHGHVhPySWFt7lpOBcEpDJIuwl
6zCwz8oKXwof0Gr0h6uxuCi0t268cR6YlaNVorW0DBmhJk63dRs3O/ADCqKTGRSZ
yv1+XcPdw9Oh5i3i8zFYeG4QrwQ2w7XHd4b/QrryVT02ciUFUmEmxNenaQ4Z08dq
Yp321/crcMjHjjsFZDhczG7up56qYYb9Bj5OKh8FMheuBekFhkCaOyqZl6ggPuxV
bJUeLQH8yOu2eguZWhWZ/gySAQv2dRrKRB4etuneXdu8OLY96jGisQDUJ2U5CPHp
aQCZzEbTFL+AG/i4MsGUJvf6yMH9hu/TyaLUE65W4gELffHwftc+1OS6XdNNhZyn
xMNXEMfG2LidH8LsJxCMLv8jtwy0TH19AQ8JaWCCToZHRcDa49Vci1FVnOGNvxok
V5Lyrhh737Ury4j9MjnrC3QjrPXqL79DJNT/EaENN5p1aBt8p6hSLHhe7LFyOOBg
P2+IL5hrZJ8KqJdxEXes9DkhDWoL3uwqXj5f0w7Fj2+FvA2nssD7VklnM647y0ib
nBzVabyshD/zDo4D+0/zQJ1mn2Od/+emStIn8qeuM1fyKKLAYBO8yku1jkCCHwwb
Om/9oqEAR8ZIsORkIdvMoET0FPtOtFZ+oafUL8lSBbBC+kdW+606w5X3eGugEDRl
BQKtVasHUWv1Qv0loMa79QL4gAW4a8M08gbWp+Di/vPHtLGP2klz0ObbNBgh+pO1
d9B8cJ5D5/THFV8IKDP9RftDzFRc1GQyCrsOqW0jf1oTyUWQCigY9dwEQhRz2J8p
hjEVzo/h1C2Z2dRIf2sj4etN1cS7O6XvavWMcrXAxB/Pyg3HimP8Xg9Naa1ggfgd
8Kfdnwd7KFeIdPmB2fUwBVTJ6zFdxOo3cWRX+wVV7tod3OULUUZImfIusqJnNDOe
OGPVhZAGKKFpjBfJeMdZx/zWm0K9Rxa3W+gdsEWssA6OvaTx3MyVp5CFrWMpUYU4
taZJqWBnQ2WDgJ4FqBq5iuYokVUvaFmDGMvin2GeFH+GlJJLvy8uH0cgp7yh0/FG
q2jUKhxuB8IRCW5v+F9/XNP3o2D67z78g7PcWrkyB/bXEjIPxGi68gJiEBRbeYy+
yFu3kT8Faxpcyu03D2EAMjeLD9uQC81M73ssZTLszc+DCweWF4QGFb+ktD2Q45R1
nhdui24eYuNB8K41vql7ipeH5yL9Qa/Xk1L+h3t5FE7iUJ0bcbU8YaPII4h7lgaq
Ahum4wqFKQRGCGoVWrB0COnuzsvJ0QfrRqN/R/1HHR1XrJYz+nioqNQFBag0PfiX
b4ix0uS0gB7W9DS9uM3QJONvv//QpJwLlo5u5u3JIO3Tzk+5DbNLYgFrjymjBZXL
EpqaDb79KavvcpLPZsIRpFbCxy660ATC2hWw0iO0a+CDHR/bDVnJOc3SBwmIuCCO
/gaFrS0yC3kW0LCB2bltc3fsrYNGEocnM/n2qbbWBITuuKXlJpHYvZ7GiqS8uPfq
UzCghxcL9LyG63FfNIzYnSfNFcAJ8nHTTCquxvZ/EwF2z8iMsWJTB1xBWwSKczsT
xsRQEz0fuW64ATrsQ5VEVgwyTVtViPsEjzu0kEPZmKTIsjxi7W8ALTURuNtoOjOQ
rK6kthLZ92IIT1G8rx0WaB8gaOs3DP0ZUrRW+Vsv7nhvGUYRqRzDmEgRstnllOY9
epOwPdfNvMnMC3asPyza7MzsJ02C67ZjqE4WAR7gSzey0k1j1M+upjMX5xCYctU8
9HDr0l85ItGIArnycQ+H2899J4e+2BGWoCLVbHk7vy7eDbz3CtQ8mqKqI7OYmseD
n08au2flDkrwgDW6YpBKvCJTyrCUAJLUC3F4tfPl47SLnHdUgqy6jZq3EM9p1E5B
/rV6X2yoBlVI+0N47+PzMr/dt6BvdYZCgAO967GRfuxNjPN04XcC91c/l/hDfl4c
U8UXoAbHRWtqUtfN9+LYWI8vlkVPn98Oo5kIBoN2Pr22ZZIc3CSI4qgfBH4o1lCD
RURD/7BPchjLOzPoa2a+zoBEWPLQPIHkVUof55NlyKMWRxGQoQlBdkKTT7JJPOki
6p83RJEBDY0C3UOzdXX5oGGJpkZ80zBOeDe6mK4pOo0NdFsC4a5atEgRi+GVlPn8
MN5R0Y/b9f9jpnM+eZLtUOMBQxUwmGjIO3USOr1IKAzxJU69ymfjHWfCZXwqmS1U
bnv568R0mnhxLzj2KbF18nV53zVpFN+oybU4iI0Yjg9Js3i1x2It7JEbWZABcXNI
dsNzbg013tAY2GcjT9isFT1Me7Qh7dMsPWBJ6BmWs5Cla8eYU0X1qmXJItxDfzpB
jses/WKqtRWNKHJgFX0cP2cParKwhM45K4x7G74mX6xTQvKquzCjYeUAtNKQNtGh
GyHEPvuyAMFO0mfzKreG+i2j2TPqfH5VbmTQGF+6f05nIqyPNcna+wZRpyiRp+cu
0PtT0MuG+7MgsfTeg2lMmxlvJcZC9L+bXm6XCE+y9VpnapZfPmWrhMhXgff/oZTL
RlhCKwO7jS0/5AAtGVYRv3uyuK3Hgz7HUGnh5uTs1nj/FLam8bKAG4cuS/MSTuJs
9gIdgEHYxjpQbf0Q0H8Y+m/F52X7set9QrAGpl9mh/llfP/XOIxV6VzOWzuxQVag
Vo8WLvxYB1xOiwj7YihWVR/mfBzBflzFLYGRFQNhYvwHEHNJJTm4UpWl70B1UnZx
Kqb8V8p6kefOcgLEAw45DbiFWb+2IiCPI0zkWeFDgR0rkF66nmlu0uTcguXHoWud
dZXFccF59KqSjo3L5iMPdVTKcTjuOcruOqzKrWVRPC7YvS90oZRElGDnQtiOLhmu
SGu3lvMs6BRFIw/p6Z2sDDg6vM7lV9rTEuq4HF6fCYPugyTtewvePD8/nV4tbqn3
9iwp0WPUi7Pjs9ZNX85HEk1VU+aTLc1QKRry6GQBTf5ErLPsS5dtYgLRUMEAViJt
Nt2+tZI1hzzujjV/prd/YjMhoZYtIZp2Ba57lMd82qAVoihwHyiYKM7XNVdqZkvn
VLwDhGVrV/v9n0j2aG0Coil56z0b6JPt7dSi6yfp1Qv9eltrHYbvmVSD6CKIAoks
6j4f5YFARCWI/G4z7Yqjpg15lOsTWfbPyvPsSOgLBCd6w2pI05x1h/O+BEqsTdQa
aTsiseKDKoiXhH6ras/PO3nJORKdIkKGBPlpY47drcTsmUIQ/Lu6LleIKzuWjMkP
JKwEP+5UO3jVggjzoeaiA8pVRTiSmc5sFq4ranQjw3o/PrBcvo/eAeQiKyy7lcMz
8XpxqcIfoAuQPXepKr9udJLyUBVMNvxtw27rRYWIlsvWrDcgRSFKdatrNgzJX2Eg
s0S1dg431bSYF0MQaZ0zhLWEDbOwCBimVsgN6UKrL+tGLe2QdhSd4R93pstUvyVN
1pz7IEfAl6k7EMoNi1Y5LNDNn3JuOW6W2pTXHXl7v3dwseRstb35Ai+a0uS7w2Px
8HNsYwSGVOu+Ri6T7amOauzWO7sEK/iMrqEFUtAwA0qqAzRd8lpCnHwTXGnlyrQM
XmmluBktLV5Xnrm6R6jrOUSwoboSKVESUXC/w/BMAqfQIFTuQSGDx+0a+A5Fr3zt
+uMMPf0a2pdYNkGN1zB2OuR7xi5YeVUn5fnp+YRgKYuCgomy5wArsPqeOg+cFqP3
l7jdWQLOFrIhBs8yJYuznBlhqvm/BBq1SK1ZvHcAL2v+gNmj/wuJlE0aCc3BZpEj
SUe7tRFDjWx3wVR8h+zZd7aTRlV0lJJeNGMclgLnDzGqJaKFMKhc8L0ky1XQDvZq
NgwFdOXgU9lCjODhYTDgLi4yFwxe/J2OIkYgnDumkjit4WDdDk2ufA/vcB8fnK1+
+pygieHunIgFbiuw8Lv6MDqIR9OII5vfy6CZ9PUmESnB794WbwApjUHXp02R04tS
8ApmNm4+mo/QxRuw9PsZnwOyk3tFhQkU22eb7JnNdKp9QFe5KXLJ4n+A6agQNOl9
AeNc/mOzCJ4HOSgeUaUgH+oJQ0M5JVyJB85bchMowRsBCfalvEKzfL3qZ8BMRojF
TsLHnH0cMcaO/qFV1Zov+G9kJC+KekBMR7rGPYnJG+zKU7SbQK2TFvwyieDIwG45
LRXKlISBotSmN2XXcRkmwpnVYZFd0OzCfHmIvJ0SQ9KNQAlpOKUKXlFU9Eex5aUP
xzlo7b3XDOSQ/8Js52kK6vFRt9ENTQCx1l0Q35H3XAlp+ORJzmLHaJpsj/oH7Eyq
BVrr+us+4PBOEkCaXUkAHRE/iA1HhhON5KblQB6RoTfLoCaRk/KcmsbZehsACFJZ
AxBPHVAy6vGwzO3lRT+BUgPVvJmBKNYAJun3mlmrbAig88BHXvCm9sbAmLU+HZgF
LQY0o0oiykpZ6o7Z3LGkSOFPIEZA+3pHCEjRNG13i3s5PvtdWTouS4o7EwtWJsWP
srcVZ+/kx5U9HnVqVQsxrttTjPJBMK359s2g+AoQvh5maRtVj3AAo8tOam1vKRpE
fb4YW1N93lRzVSsNtOPL3yydXgqyjygIOpdgLkKC1IfqrYkdJkf5AjBHE00l6hKC
4eJycWTXU480veZ6N0QT1Kis9+3a1zwjScYIn6G+4G7RNRTff8+b3xMToYTze2DX
2U/71eZyLWSkRVUo5RKHjCfmyf+pJO3aK3LyN/FoPy3/4aIy4WD6H/VdqJ+B1gHH
roi1MRcFb+v1yd6GB0won5zV7XRE6MupmayRgOM0sS/nazbPpwtbuIAEKo1293M7
CtNmt7OkOLk/ojQS4MK+MdetKX66Ju66TtofiVN6HCcSW3LbKJWIr+iHhp8CFBWY
J8r9M5HPY1uqaQz+qN6TC4/f8rta+3B3Wv+3wl2t0tY3pyoO4fS4ZNiYbWm8nQrm
7cAnzfC8khNKBSVrDfjsyouzAqSwY7QMm/Z9soH8QZ/VtlMsjCAkWUXcermk2eqE
L7ULBUwOKjXv0uY/gWj+fE21DPC0zWF6Fqozd/DXJFl+xpkw/WVL2gWpW2MwncU/
rkA30O4MKUUqg1lPlrZkdt7OlJ4cG5QG6RsGtvFO36GwQCJ08yO9e0n0Y+CnjGaN
sgWNbBNg8jzK9ILbMqJBq62gnXN5VC1hJg1vlByJqoCsyQ2YRLTWUZuRLNSflGG5
He3ub9ZmDpMWf6LSQpI9vhKO5yDsRAPc0ArVRePTrJG+VxNe40TSIjey4IqzrR2+
JOzx/9J8HWXTpJfcTJQTB1rJVV7ynv4Fs7rZe1usiUvUB8t1F1w9O7OAyXZ/ne+C
xvo8tdehfLIK1LhkN9KhE/cf8cNw0oaoAqwZNww1KA/c5iMGzZew2wtaIxI0ngXB
w6XaTMSWeBoubuUkz8Zbaf3vFuYNtoAHkYulhRPpcQ2vOF6TXdLriIgntx0Jo3JQ
RdFVv8C+NuK1VkMI3KN1fbd5llaXcCPAJyYYkLECM7mZz7fewk6Gh3EqsIo/aA4a
z7rhRwVaBIrPnaRnSKiGjRi4JaI61E2+pTtK4E1KqPZ+2AqrnqaXh7mdeRM5U1cX
yShK+7U6Gy/+NGgmfSvzgN/wIeRhvSZbm2tzz4OmDxQC+32U1pxHqPKfnh9qABbV
RLrw3VTvYUkjhlbKMNB1ikhg0liLpvoY8+8YXZ/dj+C3cYYd+cm8AYfodQUZnXMV
lu8wGN9zCutKlkowuDfpdGr0nE/pzQfer1byCt1wJ/iQtOzs8KR6W14D/GwZUAj4
5h5TVfjZ6kYruvdhttJILMgWRebazak0ZYLiegvWz92e6lBhk2uGEl/0qt5u4c7m
Ojt7kDo735P8jxaCX7enhLusST45kgSu9WR7M8UubGw2kbKODf2/uKwfTM/f3aiT
nseXgOEctTT+8nA2IwyRTOHbRPETmlLZJqwfNzlMC101rGoXhEOjUJUh/01HWN2l
gLTWCx94GeeNaAyQpHk+IgE5DyA/G5Ubg7WLG5AZ2TQtg7n2O028PJdUyjaExhs/
7bU1xXJOKfuXy3xurYe/4NmH29J2cXp4RNMU3MxIUw/KPzaSU9HCpDi4HqbnXTyz
49UPF0kf3+62MfTWydKal71nLYV7p7TVPhRmdwiqZ31On4Bqe1VQLrBK/9MoQqw7
0UK2eOoGD3BtzG37SMtYPEXwXqZfhSweiaegxJmBev4Tq3dsJt2DVdeg8DaKy8dH
a1iA3ADGW1fdjQSzs32eW31C2NLTFaUkoag+cLN81+f4Y7WZZaJ83FVLwFiwur6r
y5Dpf86CKmVmJelTIl15pxVFxhp16BM50aVBquLIsTbFmsrYjoQYtNjpHWyxEaWD
8ScXtYGEMAS20okScqW53Ci3w+FvoYOQnIUY59VfBvTAOcJ8FBDxAcWmVBtKmr1q
oAdUfz3MatzDB5iPk+elB6gpFxLscGfAIAs7Tn+rl5Mu3foKBMNkxCoDrADmm90y
FrNAQyZnkjNXrlmMAKmVnZCn35GLYRIEAgcQsN2ObWz8I3ISt7yzvC0aT68KoK4B
KciZeKsduZYuV3j0GRYhkI+0kE9rLDaeon/9YgIJYOEvbWwewKwpRr4S/9lyxvbK
0TcpMVcnAo7s34/qh2dV4zfdR326mgYVR8/RMseQHzgnRxD9pt8NDu71RLaNawlg
5zSq9vpRnjaPMOZ6yOzZBap31iJkSO353vvlnYSygOuyxvce0V9TeW7Vx/N6l3RG
uS8kN68YT9IiOjDvWbU8Xho38N10Jr6CHBdICgqnWEaeJ/wMF6a1Yw3AP2Y3SR0K
PbwiV/oRh7sFkEXFza8TsJg34F1THENvUqS/HYAdu/szo/eVQYPCjjS4pcOqPfmu
Yy4jfIUZrt+LPaY6De16rRPvK014eoNKjr64XCHPpWgTa2VnkJZUKVsg5/6FEO3H
fBMpR4Vyd9nIK6NmiG4YcnosnPKLuvmtpqyyiHPL8WuTwJZ+EYosLhAHJNtOz9Uh
3HzDs6BswFOotvg/VMskFSXw+D2Ld6HYv/B64tGotgrG0E2cq1IxjkIdFIuEjCYe
9EPhTg4xrJS6T0ym0FQ6LTin2M3GGs8rKFVTF9Bo4BZvn3WWnkZcTJXzwodYmLrU
KaQ6Aqrao9YV/r7JcA3lcyq1c+2sVuGBLRpIjASAm31HSwYcpnNKCD04p6OE6rDA
QVJA7hJFvezyj0GrCD+p6q3jkRpdfPSbLs96zkL7Uv3b2G43e0PV7EUY9GBXfehX
NqdfdbUqXFvu7lFjMDcSuz+RjJkzwOrUp54hDYLaxvCqW6CeMdiNQ1lv0iy8sUIg
6GULYzuPPnmIJ3lAMsLth5huc7ZIBnZXDyGckAl2mwwmfRCOyhXIFvx8cq2RRPbF
dfyCo2sgO/Z3PH01Df8+DCvp6ByhvRJ+XJTaKdKPbm7mPv6oLaiVBFvS8L6P9aKT
nBEOJoOSjFQerQb4o+3EfNJ+KJPigGa5pOyrca/LyePjXlaPdOW6Xe5gOIxb8Rqx
H3bweFsKW8Cy0im/R6P8MaOHoEqQdvwEowsvTvOtduH9XgPmj6FK8+s8bKnYMk5f
DLkbCjZAyeI9floP9Sw2Mg9KE/xF5ZpiKpN0hmeX5v7bUZ1OEosV9NuG0K4QaPEv
1ujggKGn9xVCcfGtsEZITarG2mmGG0p6VPcUQuZlCdTQlWY3gn/XOOh/21zxFC2A
qAF/5llcDnx6wj4mHjfAZHa4R2fgHT66jbtd+g6cuSF4JgtMBDVbJq8XN8bjhGuo
53XE30RdIWHTm+O6zYVWAUHzCyZaKDANRuo6Y1bkAw4tv/TFgNfz59E7e9nXkoPj
SoEHmBO4GQY6X/J7ODu+6RGW9YL3Y+dRtIQ/kDn9y3TNuyqsEOcMio5If1CfXfyh
KRamwgWBDkG4sPgvpKwSyJAk5umsg/hBy5Gy6Ml8leta63IBY++FZ9vX/5Ybowb0
xZcAPZ8oE3oaJJcKWDgbYq6VE4VnBoPQ23qzvscIwBKrDCly8a+7xJq+7RpEv63J
e/nOFiDEWtDpHT2IzJd19/y91hk2gm0fPycRNtrGr8QTnF4VntNV+SuFwbKyjsxs
wvgxOi+I1tl4z6/sd8tXHgfUKzRb0b07j88oCC09h7tSWMin6HkZAMM+ZAEHk7Mb
HiXCOUKE0x9iX856GvEHA8fy/3Em56Ku5xF6HPre0U/iW7vwnjytFvo5E1fkY+iJ
I45sIiZhD34rSH9G1KU1/G9NcuFaGT5p+Ta3bZwDLuv+KKPEiZIBsjQR+V2cTPFd
rhLikxWmO6XjculjZFC+JE6Ihjw8gZHwcspXy+Hqd84rQGzUcVEQoPBivmt5YeAo
AL3Tq7J/Jt9kvV18yFeJeojBsK9OLXjWebmIuOXXm+KVdA172fhzNutTXqHlweAO
ZwXzU5ilcFxLGUer0E6gSu1NlfNTaThTwSIbrepwtFl5l3ezSNBIQLRXNQBPH5u7
z7y3XRM7LgLrw5oLtCBV45M/DvuUwHLQps/rIxVVKuuKEdBk4GAhOG+7j0xXeXUS
e1tprMYo6v4wpzmT9slBBt358o/aovMMmD8iWTd441YWylUrC9VwJjCBbliGK7vs
JXHpfr0SX61c6hsj2jcrq9L+sBx0hDmcK6eHNOQqJ2zosBf9r0K51BuwTBXrgEcJ
KZDnIY7nH+Ye1tOXrBIYQXFpCrbBDg9TFr0Ecy9vme0HhIlFlIM568bOlTLZr2m/
rdw1rGWcBhHaCPErAMH+HM2izIrrmwOgmxLAfJYWRNMVl+1qSSDwejW+OAWWCuQm
Lu3xqMnfeGaev2RkojhJRlECva0QA8joVq8jFhkNfsi8PkbyZnmt2GrhAYBmdmBM
B78y8IafSYMMQnnWwCBT6nmCvY5Bu0j9bq1q9cRyBTSUtatj5LV0SqmriWPQbvgz
dUlZf/glejeErRWT0RzLOiTJFqMTnRcJ1ywy1zKnFbsE9tGAXolrQj98JAkE1KuA
CCkYjkcg7EB1fPVbOP8n/EcGXddifchIZqKPiEx9ptdM0dZpdIZNjAu8af0YZ1qZ
jUeq+o2wJjNUCvREwx9Ik2nWLEEYYBC8PqsqtUfFgFTRYdXF6HsXOHAfv5ueVSih
4EY6AW2nsuvaoVDQ3AXa9IIEWcjtbqcV0aj82iXgV6XD6H5truITQR41ehhlNrTz
UiU3ds6/YF6e+qC1NKxOz0YdxhdbVSN8pi3rTmL9XFBJMAkjGJMdMao9m07+JgnV
nLCstHPSvkZCgVPD291DM00qG+LBFniDKQ3ULtSrBhTiI0XQBKphmdFk8p7uwty5
7XXVuGL7hFQ65/sBT1KjGKOH4co+DyyTe8Nxakbj1bnMN+OyF+Yc2zPVYfeWVHZF
AZuspNPjIGGwmheWFDw9lw0E7mKrbCRrvnOwsF7RV/QKRkCTAZFydnuPIK9ka92q
mX+px6Gx/SrWmbmN2lZlR4N0HWcJjZLlN8TKsu9BQcscjcwvlsy49q1+pH6QOhxJ
UjGR5GB3jpMx0uS6C7XjCMgsouA3gxaUlMZ+9wFPBYZDABKrQpLk2IBVt316iBiU
otqLJerJdMoEys9iq12spGbyAbWYvDcd6XSBchCdHtXxnehmJZxOhT//rGosXPj7
hLtN81NOMucikDCLkhbq/NtbBO0hH0HAjb+c/GVrqQm19niE9Z8cO7thpVqnTle2
WnJTzfz3ana9PQ26GiicojJCqpjUd0AX68JygxMuVnd0oqjZfFlF+LqkKGi/Abdw
1RIUrUrsDDuiFOaaCPwaJiwumDsq0zbpDlNIusNnceTy8G5QwpknmYSuoQHqnXhz
Q9u8Dzct69bVWzjRXJzBVc6nkRip0ek4p8heSxxwveQZy+46lq/uRZuyqJxqg+Yh
spsMnZJ+trCJl56RkFLKkSdhCTQiUcR5uMbOGtGNSBk+qTGmFQFx9Qgz0UYwZSgk
eMpShjHC5NF1paC9NIC8MNgQduMruIfD61KTtaHvRQHFJE86hRlz2wlIvjLLqLTK
FY0h4Dmk+SSEBL/nnjsAz6k7Dg5zYeHPYWjfx8kmUCzpj951Vbi8Cd0gHtyfaVYm
FxBvVcCXxo9EswmVcFv6evLVQUMg6acw/K/UIcolbcMIxnIsqxcNMMpEst1RIkJV
Dw+g0ZWQ6pPwzBvPruxd/88aO5Nn4eZ0mYHMtbR0xaKF8I7FcK79JEZ9tqjAx+YC
acbTB0+8JCGi3Ge1qaDeQMh733TerjH9i7pWQ4kmyQyjuaIaQmBXewvUGcwamjzY
MshAAFDM/5m4uOec5C3KLwQipr4mryAoXYBOVTOZOUIfoj21p0repmEqDs88z5Ya
A+1UzwIdx41NVWyy20BNSjtyNUnek4+G77yB8xlW1YqOQtcIt5AGIQaSSnInuWhT
RPsM5I6ry8c8G8qclkzcMv2Lbz8Nw5zF0Frd4kk/xt3IJBGznRMdBokd7glHJBJZ
XFEugRGiJiyMbMT+8695K8G8Rhmq/8UMuq4SGNbIOdVX/RXHFVNB+o0mJry7zie0
LIsL1oJtZTbF1SH3PjJsyaVOvCs9Wgsl7dkN2qjYhbuxj1XiE7zVj5A0VvEocDmN
zyIe80n+KILYrse9mZ7vfU2OhvjHu1VAfvbrCmfFWrvK83FspJpE1JWHxwirJEkz
Hw/psBhU2x7Am/Jpy4JOIA+q0M9Wnm92zUMBRg5GlW22H++dqBTh9nilSOlhNIhm
rYWs9oX3B28udS4lvHBRuMDvwh2nOerbQBihrdwgWb/Hz8EZj2ckd9+VyyMKjWXT
hslU+JrxdstUJ6h/A2j1z8AULkR6qRvGjqf3rvWGoKcADcvET1wMaCnBIg3O0+2F
5dHoIypdJeZwU/P2NGW8eBl6vgjeBFVbdmF3XVvtaw9DV9/T64LK7Rdo9s7cIyzq
8lUHA2tQykr2RT0R0FThO+XJGTaoFI/kxj5IBEg3AsAQ8EljES2tauzX5D20TgbH
YHd8ASMG6T8y9aIvhO6lfyDExISJH4NFJ6HrlgbCs4JFwvL2FuyFo7zcctAlMkZw
T/Uz/GDhv3H5UbmOWxp4dcN2HUHq+2DswGvUKdzJa4mgbjlar4HC79cZ0ENFUV3b
Cjf+dmqCWkASE/9p0HLD0FUdJwUE0r5RCR5MyA4FJg2FwbAOU5Fu15JBhytGtue6
dJFBoPOyiPtmVP+0wkEvRcbKnNRWXWC59KP4274EmDVVgGVHH6OwuI6/wvt07c5Q
lAoa/MAUesGd4Vk5GT3/1wXh51Faq9KL6XYhL3JrKrwIlbJElJdIQn2JYu06gGii
yhI236vS7qf7VxkleSfVLfSjIQNEsl0OZypkWsNKym5f5ZY+DeH1BQqDuRGoqdR1
otqgqlln/Y8yrkiYreLnAL+F2sFQbxlKUfRMlWeCEvpP0NqHeO/QOw1aDj8KzSmX
SOfLTyGT1/jU0yaHnzm6m0HCC/Pozfsp4crW8ueUOq6MZztjgrYrs42OOQ/U4Q1x
ijS8+K+lLmFSlWsMU45kz5vUSAD8B5a48W/yzHvBOgPSEQ7jNrisI/Mk1MbR0am+
pX9QVHYNEK+lHlUd/Y4hUYOUY2+mda5+Rb2KqJwx3uQlmD2XyWsl4SY67e1fgI75
xEFqDfdoLllc30y3sIFGZozbKod5rjMpU2bFRHtQH9Eb6xtUdeZlFTDmszXtORL3
o6t46LOqBw0p/eDEq7Hn+vABBef/eNrQuswGxs1q3XrhWPF4Mjng+g+Yd28/PmXA
DFNl2KvT7m1MYn/z5VlPl13l5N/RfMsBcI1YCid59S+Avq2kwxgO7iCHZdXMSPKm
fim8Yq5TxwLQPVk8Q6D6Ap1SpGbSkY+BJR7JIlG5mXPbDM5YKz33VfZ++aNP8zQY
NXkXVc8/t8TnULuTJbAGI2+DOknHgagEqNJiF8Kwv60TAwgB5pEXyy1ZOHGE63QR
rJDPxtxOLMZoBRVjFSVk8nQY/Rgyb98UUhHi/PZyq6VZPb41ZeGx9zIDj+7Ptdmo
L8zI8PCaQWEgqLPP56Q0lbUW6pYgYciE7Mbw7ZZs7CBp37HEhnHm364cz8gzJ0W6
j7vJPuDJbxaoV4fY6qHKwilc2tcu/WpusbzjTyX5Ug5hNr6xe5Pr1AN7cjmww22y
seuNw2RjvexpEk4XRJNWbwOoXJ29n244zLuYIgBD3RyenRNSWVC7yR6/BVDPBYT5
RR4vfsS0As431LJiyxTMb2O3moqqs0Gd2uRnkLaAlxODIy9dokbeBie9fGpnNin/
s8pNR28MdfRuKYBYOfd3bREYNQIcwvFZ9WTGUefBBR47hsE8RA9QZtdHHf/tKdPN
gqABC7phsx40qXqwqJUNfbE1M35YfZJ1Fosl5c5yKQ2iGBo1PuFRcYg+5XA7idm8
JfezJwXh22WL/gQc2VuiDlMObgzRpwpvC9UMjtoeATQjfNA83+26VMcP8k0cGbMG
+JlPI3vSJEAG3/ui2k2oHpFc3RbFhE8NX1mF+o/jaChydTDutdOHVST71EB91ilZ
HIr2C6F64flQzppTQsyGrGankfjYyRuW5LiMEZiBpEydV1Whj1my6VZogG81cnzE
3z0dFNyHf0pFFqdoGtLHyXpeXH7XgrugeurUxsrvvj/ryF4LZp3sllDy99WPzJpy
1dmSi8pRz5c8SMLStHmVD/lz8kPOntwX2oJQKIcb+tm6dLfwfq4Un2UUFpewmRyc
XKwjaGkd8xEZJkV84l0pa0JjIKyFTNN0euK+czp44gabYoEn42owKKPKtxNJAtSw
uLVssFZHDkqwtpQ2Gxu0LECXkymjZtWBCoptQLqbgMNY6iWVKcSPGBI5z9EtiPfI
r1XUBO04Ygksmah7hYQhv7U3wOwCmefNvzyPCRDIh8berO04r1PYlSiYRCYlV8bq
ouS/PuOuSvlG6Au6JBZorV9/t+JRlTOXztbxu//+t7+ptIb3ZlxfOJiEG/7JyX2Z
eK+xYmKomUPMDpmSd3/K1BRwNxVD0SWt4Uix0FsqqOGtaU7PouT7mjcSwVODVHh7
h3TThczRgPifGxH67huAPRzL7dQcXrOLxwNHN0SNqzl2D308QdpdBqwZQQdY/oXv
Lg1l1PdewKJ+jabk99xW2jfCJwmMkVKGQe4Epsvjw2q4XTY65W2pykD35X3ihCCx
qPqDpjHqAS6rCe4QT73Y05tDxXIHzGdP+VYjIyLf2plio5hf5hPundpxxXh+vwUL
zObuygzIIroD0nnoJzXViOLS7CNpwuVFqYfV27OOls5vTDZy+e9JWUL2gqxW/xYq
1BzEb16fuebyQhYqzOsQxR1xeJWrswEsZJCirwoNoUZNqhR0g51gifW+oiOx2Pbc
2siSvQqh/Z/xUyg9YGTV/YVf2fPB0IViC+MDp5v/L8KcnRcakHSmhH7Sj+kVZPtF
hU6qaYaHd4udVB/YwQo6ymnZzKL8hE5/eimiSlnM23RnQTKdRUBUBrUidIYlSau5
HLrXs/IF31rUJx3hjKnwu2a7emPL4CIK++zQTa8STrtVkLFyM/VUnAyEsOViHvFB
RkBXKeT4C52RmoktaNpdlPscBwIOq9X2dNVPx8RePzaIkkWKONURZ8Mbl8BCT9dI
f2SypoBH7W3Ow5iIrwCVp3oK+m0v9UaKqcj6nQJp3bhSZy/f4IedVN4de1sh84on
ei4FVgaLj6JdQWCZ/zEkETx88P9WGze+Gd7oTKD7W5IV0PXW9ALBv1E1SztCxz70
JweuHFpMA2189rryWh+V1p0ni5hmAitNaBqg1QdD2jYgExsgP0YMEkIdK+GAHNQY
vNBpBvxjt942vQq5GO8cxvfypNCBK0RTFKqHFbfvXsCfdr5C0r1B4SFXVSC3tvCe
V86UNyElt23s1SY2TRTlAxektelC8aQbmFqA7OVreAWA2CEwcTbU7I1IBWlGI6FF
jMzncZPxP6cUWZCqduSqKQfx+ukQh7u0BMfFh6Qe17vdcFPiPYmCu5oSp3hdsKHt
u1yfTbmIpNhuOaJmrWqert16ZonGyYTFLhqmHgB2VXSU9mBusKNPs+AKvPf82qDs
fOs4LmGOWzzIepMzy3Rhjx+4VkAvF1hntgcK7iG/8loQWHJ4CdJeSkUupv6oWIc/
4z62kBE1/VNvGnJdJBzBckYPQQ1oIGi4AZvmaB/fFJULfK/HTrG0PuaJ62Aq3Da1
cFvAiBI0NUISUjSUZZVox9o2yQUYMnw/cfstxgKaobsvsh5uZK71jR75DU6cv4yG
MKC6ujaWBmMt3+w97JNqN5MdEDREzw3wWzF92X0qGswNVisFpYXup2yLxKcrdxqw
3jd3j2WO+19gBaTLJS6X5szJ8Rkm0Wukvl7hEf1idProCxWRZoFRE0Jn/1cv99fB
VXg+qbobCnIdvWrGdLuAL1f/4uS6ULli1tLfS9i99hqr26qU1TlM3EXLFMBoP2ZZ
8iL1iwJnacuItcUOXlrvzZUXU4g1ogXGcJSUyZEk97eZQBVsQoStjDBmaZwF7xMh
htss+tNDC+x3n62ezPue4FAiHWtQFhKcSV8O0WFbHLejgpFXlb99l7WE3CYzjjwa
VGMhpdfFl4nZAdwax0mJLEgltBMWfZFsJYJV3G32wbwluiUPOQSujVvjj/OX7myM
i4OufxxGghhkZ9ECnwvNU7HPMmdMzSV+8m5iouuPiXY1JRPdLpPYjjvwDA9DCP29
gNUI9bcYKW6O8IEhu6QPakemHr7pJhzKi49xMXEASY0EZkHcRAnH9cNBsPMK5M3T
yeXmWusIKeAGZa74r7B7t/92zS2ecfjTLsbzPdKfn5kGPcJuWnvMi5XvNjFT3pKu
Ea6VJ2/7NFStwrjdtIAhp3ZyUh2dDUtNuJqLsccWR+Z705+PGJLpVhU6otSRJXPp
J152hWFT7fheRFdLSCy9maB/RDgS7tGyGIGUuopEs3s4uKf8HvakIj6doj3lJ6LJ
AciDnhRcuReXZFbg2AVe1WuSD6DUIFpIXTA1+W/JYFgdPJ9u4EA0twNp3VdrvxvX
OYagDqQCYG7CZVLukla0pNC7xA7OIenWuaka00MsqsOo2Ks3JeBQfGQtKnteXIiU
B/ZsuPgmv2Vih2V9kPJa4c5iAa+uhtti4zV564UFiTS+NOR3dti1exk22J/YgNro
9gYLepyMLZ180dPkj3egnkkCS18Yr6Y+n8r9zF6UhyEIgPAr4Tqm6MHbUHLUaIsv
`pragma protect end_protected
