// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CbFBpq4QHPTVjMvgoCurjMHVCt/MfJfPCbQ+0U4xbywWz4aGSXO6bKkQFAt0RXw5
m270dqPM0DFMJPre9K+nNGD/BoybcwLWkUDxsRm6p56vDnlCQ2Se/c2r8Zjt0s5+
A0SAbzyaoBCFQ7awQ9tBhRCtBQvs9E39NhNY5iq6Suw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22688)
k5oUCNa+p5DMY7gApS/bNIBvsIruJQ18sV4kAvcy0MFp0qEWLplJ81ybnfkXCnwi
4jFyaE662ULBWUL2vaITmyHTLexf24klMjp+latRtJLrnZHjbx9WYVbx6haLUCDO
UL2nBqJwNIZpawk+MUbS51Q14uTdjSPO4giwuzlQ4C+KExE2E7kQslgbqzSYSIBi
8w4jMBlsqbWewZtT+UC7LNMXeQ8yDr3lvL1EVBUNVm4Dawi8mq74d47Hp5laopoB
Jt6OHTQ+2Ca4OWkHfVnVFsCVgrkUqV+eNJFE10wGcNmyPan/XN9J602ase8ZnCMj
KzPZQjv2trM9GEURRN48DOdB+IQkOHuIk132QqXN7GTThY+ie2L1GKRHk8ELoWHP
cEDyJmc2WxZEzQiYBjIUDFZbtG7S6aZ+O4bxMwBfdZzfenddRXpLKJFYAAYVSMCG
6lxsiGjddycKUIxhsgN3gmkLdoTn9E08KLuMECM7oNnrTjQ1KIPyDrJVtkxCcnlm
NNQ/dk+SRBFsPvPNh9yLK6q0IEExk38oKkaiBJ4julesM/43a4x3iwIg3TGiAHeL
YpeC5GyC56TNwXb724ptVMSL+LVm9DoKIwSbdF24bNhLQW8JruufpEhPTF24a3w7
RhuH9UkMQHcyuHR8tnvpGiDpdoLqtrZzwW9gAXqu4yJH0tmZCySaBuBb7fp5+L4R
0qXBVG9YBGl39O9SP7p0JzGi+xaRvltALKIARh2SHAJBV8kCPnKieX2pFYjSzBal
CdyvDQYic6Sv83pmWj/BEW203kuBHyk4z02VlbD1/szUVObZd1ndxemajN/uUvAN
xLj5W5hYrOI5GBtRJrQlHIHV4xCLX5KftR9oNFuUOeyy+SGW0W5bj7Vj7NrWZkDq
mwaA9CQCJo3VUjR27UMkquam1rT5GSsmHvnJIy+xYxuA6RaTzhMWpu+r0cNGdkS1
PAM20gwOqc4GvK13qQ2ZMhr7xSxRMSURTA2cwc6V3cOrdnK+0tsbKK/Plqa/ao9I
VksoaNfoUty8E1fVY23Nht00I7J+jSl+4DlCYvPQXWoCLF8eqSkwG3Jubdmu6aJB
gKvVCL24x5FCcsE90RgmKmIaUKAia0X7hntJC5nmvKeLFV6lxF7OSd0nAhAeunwQ
A3bM/6CEZv0JKvyTqa7bE9AmqcfD7BKBPnNwmRji3r+lDnWusVws+r/EeoLuKES1
F1uTMegBrJ0jqZk8qiexAcokeQThG494gZ7A0wIeSoa3pOFPV522lDy80JOHN6Wu
y5eCG57i8CUE2lsEnBRU5srCyvx62hrS9rtGwfRfoih8lWuqi08zRm/s6vXbx3tc
jNEQk47uWMoKk1ksqhOA69xuwuud8iGK/VgATnYegWcj6vc81XmQLjz9srj1JB6X
t/mjsU7A7ZReToq1Q6LSozsWyJI477Qb9SsW23gmKqT20p0Xz8xtwmjb5nirL8qm
kr5asCGFTPcdAMy79pLz8QUIWGdZvwqgw+LYjkNpiipt/6i23QyBWf1ulNX5Mv0x
bqq3Sckg9bbISfDTbnII30SFrfatMPAZidfG1+zag/ZU0p1ypHhXzQPC6p6ineJ9
CDmXhP9ViXZxyAsHEhAEa1OP+Vtex/Jo+xAsZa/5KL52G+FQzIkMD07d/8nxlqzC
9vB4z+zXFU0YlP6Cb48XSfZpZHMxnu1wqDCE/gNb0rkoqTXEktIWx5c1Zt/+zhWT
9026368v1DqbjIYSNrlxzs5h2alCC39SKqeAf6jFXPPvvr/gcRrGpH/KdgzIWiQ5
B0EP0gkKhbkP02EASntevsfkyKTxK7smHUJ8MLulbjSbXCp54Pl1FpAKPDwyMnQw
Makr9EBcPUuHXFcpzgbBsadt7VMOYM+jjbiJ1PGY4b8xU/iw4lpN5gZsFXz3maNK
2+SsM+rcKi8qcl/SeLllsHZDITx3prapLB4MGb+lTRSjFOq80rLzxmtqebOYf2NW
7HPCGrL2kolYhUzh9pZHqbMyZgZvW7zcBpwM6ZRobcu7v8JVQYE8W72wEKOD0yey
kDDe5ZUHPlNWObuEotGi+vzX7409sJzFwJZZkeK4Ad/m0Mnwf1qQYmkqyl9zmQEQ
jb7QTn/mpS0Fibn5e4TLOnCyX9wLbMlsWFKkrJOO9/E7xrw8dkrExaO8sCVCGFlZ
jNxk11s3pK6NNiptr8txX0IbDw1lmOLNg77vwv2Q+0Bhb8AY4R6ldOLK/tj53gK2
XDLLraRSruQUvi9lA9TTA0iiiD5XPr5B0kE0CAbwl0GuDGZ56UXg1fbO1nQFuxKW
L1HZ82ZwMoE+M3dRL6Z3f81a1wzNLsLbDlnbbK/RHRh9BbSVEyGJKxWN3DCzgmaH
boXScX9flOVkWeFHlMSj3AtVKSpi4swJhhF5B4QaeBVa6388WgTBKAp7mR7Rat4T
0NmhIDF51mX7CdXY5J5OW+CjM8RDY/5huxHvB40yUpW+xt2tLsIn4S3poz7bwL+Y
dxaPsX6G5eQuhoFYKJhwtYjG9lo3xrPmFEpfuuXQMSnmGi+CEXkV7+Pav4EE5KSu
oYt43+rQeKMWqrlMpDm0huGbixJ3Iu6RRwLXtyx523w+EXxh1f2jwneuuh/qA0FB
KvrD0z7L2KnlBa0DaRkEJfglS3+/KX7VktmFQxUyO57FG6vGjVA1XZGoeJ0pDBM4
fRSQXyr4rx5vmK5+Xn135rE2lMprlfPDI7XLJCYgYrdSLcZ6W3b45+qurS4nXZ+r
vBmxjm3FwunnI7WM6aebeW8KMVhQxg5IjVQEp7glapxy2LymOyYBNeHxPdz20n0f
NEuDKOgxM4WhCBXVKv9i6EIoQOmGZYoiU5i3rNAs3iPVKsklS/FEsXd21MEtC7Jr
rzuYTm7S8t2xakepwywEUuBee0eYjETnjnTjjeiebkEy2umypR8bM7kocCWLmBug
Pe+lfsCf+og+YgEjrpRgpX2s6yTHpWbMniUKUZFfxKkSoaKwpVuxoi4qCtKC9KuQ
9R35344sa356WTaAJVYuRqApx5Wt9qTY+z0YZlUTFtNu9agHyEGodBo+lkD3oh1z
3MkUS+jBg1dwU1tUQGLPSQNe09OqZnX3KG55k93whkd8AMovtiB3tE3p84jst7s2
wyunccZedFi4eSp8XgaF9++xCKRivc0CEt8gKeGcVssj7QEwr60Tw1PE7jc2JlkQ
QcuLrvdsgE443zbg9QfQceu8JCgiHs2BtUp9Sja5BBmCykix2CGPksV+6cHinXoS
2xN1d7Ami3a64SVXV60YOSFQcNYiBQwgAGzijuOkvltBCxuqbu4txbOujcDB0zuM
twkzWfFZTwqTDMOHsgSNufUd6kv++ePKwl1HDsJc4jOwWI6VaRdXY52pXP3jJeY2
YiLUSrYG2DFBVEx+BbNIqcP3KKAyZgNvxQ737M+L0sK0Pg/eL73Ku45ORERG9dsd
xSZamkZ+W1GFatwyIeYpUrMsC3t3PN0PfZlceOYpMEX9N1oibjgj4ZSdThAYF4mS
e1vG5zHFCzZTkBAADKI2q909BsE3FsE7vsK1P5k11ABSjBOiLmFrO5F9ul9rtv6/
4Jim2xZW7VSpOT1qz3fzEZSNVMx4FEt/H4P2SEGu9PiSk0LaUz8+/RDTVTuilskX
4TXeqlunew1fBFYNkMLJp6kesZ/zHhlSckzA4ElJdCTG/38ucErRCkPs+Mq84CVl
ZkJLuhIM06xUUIN5xlwiT+FbQe7ttWljo3JOlHyfKrbAiYy+6ZwnKuctTWDUyPa7
FpY3GqmHKJXnjToFzWyDySu+d+71vzx96/yArv26xKNV+DIv9JXKIlt4G4XHxX9h
uZ87aL/GLajUUZFgTOp4uIBcOIADd36Lfw5wnAYk3W/P2E190XIR7pkgQ7UZgDcT
v4iZkjrZVCkso1hO2PhEFpXW0OgT/B56X1fumpjdNqf4UbBaKvrAeRyQKTic9S6O
ApGlhcYsqg/y4t6jKWYOV5qntWTqB3aAWFW7EkmJJ3Jp9JQ6KMXUrcTUtaVGsDyg
9Uca9JCBcectS5sKYRuJ4B6HU3kyCLn2N1xqWqEPkZCukBb3p/VDYdxrOHCZBLqe
vDhJgSjzZI47HTwQrzMpEnglby34riQ9oAdT1nV9oNLwlPVI9CcLGsbzPtQfBzrw
KRpiiXoj/94sckwiULzUXArE+FP99Lttx/mbnexHw+TIoH40/DFREwNiiCDwxU30
ABT/ETTJ8kCfjlDM9wJ6lcEovG5+viIxcOSmls+PtNqEWu/+z5yQ/uh6ZcSv+VOl
RIadD84xUoteKx56NNhoSFqTKiy7OxH2eEjK+SZ/Y0PvGfe5+LCCRXbw6wFfJFW4
r1o1lJWrYMEloTlsOKrT5w9Js5vtga6vRCaqUUivhYU5SMkka+WnFzmhhWJj1BkN
prQ8U/4Eyhd+zngOu4MBeVl1TceBqmzHepPDCpJEhe7sh8mp5/N5RJqO/nYf4KGN
gqZUcrw0WpOx0iiHikBNfl1dxsK2Q2f/EtlNrFqTL+AsSqbLIH7VjC5LEr3VYIQV
X4lrv++x1ha9R7opok2T4fkhHWAZDgHqmTb5iacW09T1oMYeWHV7RGHMNT+DQjck
C1elewI3NGKzc3Qo/t/VNhWdU5cKB3kJnAtjbqzvE3/okd9LhURufsyQnLLMF/HV
cS+7Qq5a53shUFNrnC9Np86x93mtC2AK6nfsYq59pMwU4Lw9aQqFHXS35OOavPJU
O8RQe1w0IYUVCb9JBB7cQS48YdjlgvGRfPCbVmvwGei+o0SGgT/sCVniKNdG3wh2
buvSfBe4wl5Te30ISSyJhS65+4deATZ3ydxlNbXiykB2C7S6VG/HFE5eKmu33E+S
NWE//2NtB5e+qXMwYiIIRVDS3aIvYaCp8uFLiIVMoyJJv3N0ComfJdsONnhnKDGr
fI6dSo6a4A2PXUPZ7uxklREWcqf12aptnbcJzoa/oRfRvZeWZ6hMFmRgjzmlAWlN
N43pk5Q6BnbKDvBQ5vzYZY7T7sUjISud/7DXR4eJgTUwnei09kk0vGCB54/TkD2v
qD8qCcqTNAe/A77LCHoOXaqsoWMUHC3nLzFdf6GiqR2HxMVTn+60KlOVnPpLwLUk
LV6kZPC//zUCpuPjD49qR8A7WZArndu7rCEQtLC/s6/t31vWx/LNzhtNWEjzh+C4
u75tBQiyHORW+g/9gFiUcq22UrFSga0uGYTwcXRIhRUybMnAuZyzuWkXTA8FduHX
TwErjuuf7GAAtSuSEGG5CdNL3DxOC8X1h0AyBGwjRU7VWHz53nBLse0qFuoBPBfy
HWKgSIZXLeW8Dsl1bbg5YQCODN3yaNxSoydnCluqg3UaDjlAPScDa4xZhs0758O6
sTP6alVW5kylpeQKgoHsdsnKKrEdgLByPG24jVZYE2uG0HHLgtjCZAdP4FI6vOcs
j2bsmDGXU7nB6VHb/l/1FLx5v+jmZ1QTVjniU+2lN9MQYX2n/7UD6fLc+eoH8TTd
qLMtQEtQ3PqlqlsYYdSB5HOLnhlfUjuyBOT7hOIKXqDN8RPPD2ySHu9xNwUQ1oAM
/dwat8+UpB4Th4Ub7BBiNiKFGr2brQrg66K9Ifet2idcZOupyiTjPxcqN40eMwQK
nFxnr1cw8p1LOWYn2eVoNJcDoD1JQAXst1K+dwpNrqMbFqSPGvvlLufnjj2QUpfH
bE5gHsPeklj4lFJZiRntRjABlogLB2hacUKC1vphgd4zP8c/isfX7eRqf9B5O/z5
FYlivenexTIZMspTzi6TMyIRHvT/JoU41qd35+bAUXuE86THqjAwTvmywyZEeCcs
68c7yONi1bsw/IZ8TFjKKHlC/JNDgBvDTW5BSRHOnuGityOfzmKAkR7KY2oxTgc9
KHX7v0PicC+f2psnyb1E9OLYTBscqWLDBj3ejt8jRhdRZBH/V1vLOHEOLwJ9TfEJ
s8MPF+bdc+/Gcc5vKn2Stocov8m2WHR3urR6RdVejNegaEy0+kegNn7DblrzDsZm
bxKfsVkGMqgtoJ/ektlyHaQ4nR8aDo0cOkBuH2mcShI4Oji4/uLAr7W3Fxp7PIPx
fMIiwk6HicTASfL8a9Ut28PZ+EbTNV4CyDSkn9rC0FYZMXcB8N9H/b4fxY3Oo9mG
17CSlQbEOw4yp2tmWjw5dcnDZkZkfWA1Uou0oBcncqMWHNY7mkcMAwHlRRWVu0MN
nvRoyGB00WipZ2KTiU2h6ajHQpDlzKIc6gtpYWqUGnJpHHiFY6RpodiqNtqxb0UZ
Gkqo+cOxOEXBWjSL2ySbEu9q1otdTSKDrKKkPWkIQrixr8Ds22tdj2OGXyK48i4G
Kkxq7z4RYsQitVlaF21vTivj3Wah+khYhh0EajCFoq+tVP+gFyDmWNvE7HXdrIYg
CzpecC532voOy9sZ+kjunfGuSxIcMxHJjd+KZC5r+VP0FJtPIOIKi+3EzZx7kA1G
7703tIq85vDZnG38webrVQy9Zq4HtRDoia1ix1aEQwjQzNA3IOZWl+oCzHJ/61e/
p5MeFNFltj38Ic9pH2NnUA0h34KjwWMgARBaVtbuDFri4ymrPtszjCGIn8jUVaWv
9kzZNN1MOG24bVXzZvWFyjr4DIfZ7mPqY+Gnxzw1R3yJEOQSzAcgqPLMvPN+W8hq
9Q9R2LUDdOA596rMN8pjd+v+dh7PvBjXRGaowLpXVtsUBY1ZKTnH79cljh49hRUU
AVQTlQpQH83mWnk04XLtWgciTMAGypX+u2B3siUYF0wIiKLmbr/YJrUqRJlX2Lrq
ZPBDzKCKweE8u5Oe67gnfGH5Czq8CEwX5WduNkXxufGOPToFhQOhDoVJeCMVTVL1
FZqNfRoOOkIVmk3x6x3XO3w5GSWUAy/BcXae302Wh0kSbgyIzotulYl+b3L2AXbq
PpYM8F8kGkuidqfl2cqSOMUn51NMc7trKIY1qRtXTYZTaSNmCXTfMON9dzBpREe3
ThRHByj9RqwfN+FHjv2SsT82o8B39sKfOk8T793efBLWF8L8NvGqHXhXh1bWxzfk
wc5QOWqxgMt6vhSGuoV9UaPnjJd7xnsl7/U7qtW6SUT2V1BkPq+xHKRn2RgxvJut
BLVKfePzP8VsxLvy6ziPQjfqRrmYmI/3caTLXIi8x0qoG80wseqwIFFRy3yw4rCc
iXMuyzMGxIr9ArAppZibm80+C7txtbqmgn5MhhLSfFkcVhNZcrBF3k13G5Glbk0w
uhslYeQEAXIskmBkzAGBQZkyXs/sXU/u0o9YzZwJeXF5GHMKIljc4WeEvIlh9j9p
Fq+k0ERQQqLiP2BKtLdAA0an9TuemZWhjwjTXp3eCzYXA6kRXWGOpMjUa00c9+s6
L3Gk9g10TcWaDu98ZJ8/tqIRm+Qe976nV2BBRLVzl5KsN9A/RShc2sT38vKbRojf
l8Tjd+5jlqxSCsN/PsZL6weo7DNtg8LusbJi9xUqIg1kCPyNAfTd+YKxb+2S9HIe
zR/g6/bS9Vcnb36F9695yEaOaFmejQJIlXjtKER/CxIDnZDqONymjgJyLlKw/NtR
aReyuc1ry+dGayp+/7yYw+h6aGBclfBr7SuOU4rowMjCrp59f6BhvN8qz27zpMlX
A3PUp3uUbCxVOBuC8ABohAYUVsczV77JL2HCXu2cO4li66uzx/tMIdh2dtdW4Y9v
4XF/vfUeXtStFWxefHGg3goN3B8ZF4YZVNPgs+ngyDKwpDOomMSBXqX7Wfiki1is
cD0PNWrhTqnQGrvqSPZX0GVM0+ZdWpeYr9WQGfasJ1wX3G9h6Igga0COx4MPdxQi
guvkCu9L54/1AJr/g6o/d+1sRAf59uo596gl7Jkpm5M1hHos3ohWkQ9NqusT0dYj
RDtkyMpEZH3K+wYlKjtcKZCeFpRYpvIbpkDZLUvOzh0+2vSpLCSLoXApU66SxAz3
cTgD3HQiK9xAZavEpu788P3MEUu7sBfIR+MFM+ynYlaSLwtzZWB4aSs1UFKl1ZJB
0d4AVgHZKLQHF2GfVKG2Hhjw8bbGhgXwTEMvHpt6ZkpLRm9IzxgwoOt42bFCWQA7
d7QbBTf+ZlomG2p2khyytKBha7YuOBCbeSzvbgEFQrG/0XZiGNUqR+X93cwLN1Tw
c6E5Hq9u9uEz/tNhSZoFUd3m09d79SsEr2OndQGbeA8jLn50dm77Sf2rV5KxWR2Z
HoSntykq2mzJIyXPVefs0sl04jp5j9nuMJgbNR0lCtqLxolEcb4ihMNcMTtxXDKG
0xjIAdXHzXr4gdM9Fr07IdFyG5PyvRS7ej3pvCEyETuxIZjVZBC/ukAsGKNEn/nf
H/lt6BKfKBNgCK9Gl3bnsWJSCfrD58pyZmlSZn9rzDJtsb3NJwqtmp5leQdRxqdk
jZfoehZBxMOvgzbpvMe4Yb3cyYS8GKW0UFp93k2ZZ0jdqZlA9BOu5lfBw/o4CfR9
p5r4nEKdOpiFbS1nivPnjA2nGg4CqsiMEDDU3uRjQ2vcXY4XcjCrBcRIV+F5JlmL
IqeIKGHiXbpkNz8UXV59zwScoIn4smyJfY2v4A+7DnBFXLzAizuaL/tR7IWz+wvI
2zdeNT9+p4iWJmX+rg8U6WaiV9FZVNBVoWdu1bBoIXpmFrn60MVTCiwypNHuxm3a
GFK3wypF7yBXYbZ0Lv2PceCGnng0BlBdehdYQK/8WCNSE/HUKS/uiPPnRTsuSwiT
MhE22Jz/LSwB9Hr+TZ4pWMlV2M1MkqkFyX/mD+8qlXWDTjbZyRUjWLtMrAjLxZgB
Fc/PDBU0oyArB8yiQ9UTQp3NhKNlXuK64h8O80RaNJJyDjP6GwdFKIE/pLF6pPZm
JjkvSF5xECQ9WDUsZx+u/9nDV1o9Uk6QoFRVFFtmwnLOa+ofo2v+Gr/GdB4bMIRj
+OaP4Gm46vr7OxhoWDkRvDDq4ou0lDKC4S7byB6DRvyHTx/aRfm10Lr0sO5cqrRS
UsBytsmnXD4tzPoo6tSDgWl9vrRSf2oWEjpkax66fkS4Ym4gEBoC1cQN82B6mDty
loQApAZrP2DoZS9iFGhMO1KBIxb0NF5TJl0Bqmc47BDshN7rkKT2rf3H307bqKQj
7DIhsJEqQEeDCyBzppoqf8M26iaKuTU6UOBRXxNTAEI6Ia1qUPeVArrYzbsRjXsd
AUvOk80YZq0cElu79IihBcsDxad1lyqSlRwCyFE1kiAff3yja8GmrT9n90seFnn+
IjBALHPBJrKBDmzeKZ7UrLczKJdqYh4dfQl8GGpMIOg5KVZUaueZdrpJhW3o7Iz0
l+ugHJlrvzUUAk976D9EnVJNneyB8YcwvHIOCcoOAJJvUtHkRM8gGAjzPje7O3qt
LuNVUMZUi4q9RcxJ4q7HVta9eB/8Tr07wlQUgY3+5yId9Ifs7LYTcm9njQddOGGK
BnDW0cz+1wVoWMf3qOP/uteqyuSlAahJ7yQjK8JDkXC6L9U4oNW2VwiYSFklMhq2
geXrOj521oeLNwNLwfL7TyaR+bWBegQIX/AgksvkWdAzXSmlPZNwurwLrtc5i5GN
tAhGfIiKdCZwQrx08EtAu2wJAqyvr6o1R5PTfii+JOvxjNMSI0ZxEDm5nT2P3DUZ
4KePVnWgCZBQI+PD257O6YAgxP2I5b2uh+c/KtDLD79nvXxglBDwq+SXlcm58La5
8F3cqJ6W2p2HWqHuCcXNpFg5UlTbodzcJz+PKFZs7NWSydHv9xBOhodFuz639orw
DYknEtRv7OU+L/oPg9wtL8xTn28Ci05Bniv4fXZ68KSNB6F2Fw4nI3/DThBpoSgN
T0PPhuEgJduvHk81n08P+q//1aMjhNo5L2RwvkXW6yus9g3nwvgCPN72SFzWgWah
b7mIK5BbCxgZMNsgicyxywFVOPkfWVInVvp6exbH0alKFVelaw5FHw5RYtexqwHe
tFuFgAIPgim5LUW6K6TID6+GExnV1UMOw0zahPyo41JRdzpru8cuqb2oof15DE7P
OPab4/jPRw5pm0fGdR8dvEf+ej5LP8ZxM72fseTWuCv7frllcdA0PWAISC98QCiu
ZyZflWp2JBhfVq4x9wmsVH96z83+BUkDtAnR1ZbBTbf4hes/m5qS65DOsTrD4nc6
kduNr1sdHXwg3k5aNHwIf9E4yERGgEeZMx7neJMprYtn6CexVArzMsaIZztT1bkg
oVJdLcT2bacEg6M0bBrOXu73VxJdXNlygbIySom9hx97AtXTdlwBIYBSuSmTpwU7
MFd6IJcePKMroq2bVqRmWYGxJIBkB3Yo2RO1U6SJTX7owtunSyi801VSn7QvudPm
cZOLZy5VkLoiieq/TZQjURHhbjXbE5bDh2ilQ5sGgN/XIqzFFxTGbAV8a6RV5wk+
bqqjyHgZMRvXnRiqG04fmDBiCOfXLhLYTIGS9Rwi9rchN5thGWG1Ph5UQwDfUvFm
1JmnMba/9ggqrzsd6L382fnQrmwhrwbwK3lu2PvDpd7J0+GOOfdnsqe7BsLloxWv
8LCwU78MYhQRaMOcSBX4cQ27LGJ4IajNH5iIVTs57W700ulAsuSZ5ea2P7UQh6Xm
YOj0rb5pHscSahIDAqR0Xhfr5Iv37NbGN9DRC1XPbHHnHyknfD/R8+SU5D0G6SSI
jUHLW4mQrG3qTt64H0y57W5EXLsisQpQYPa37U9ty/R3piHCWoKf+WKpG2oX60Ez
YOlNXKDwPON15j4kJ7hKRD8+1meJBR24sV+hs7Q4/HT2xLnE0WuSM/Mwfv54ZRmP
BYWP4maKCMZa3B8EXQk0HTzjtuP16r9L2vl3cn566Tq1dwb4TD/84XtwlQ3bLIen
c3DQXIZS2PQP+Lnax/coz0J7XQCuwYbEGa1d9rlkP8FoXUdrThBnx9C3eFuywFtO
zJdYY2Lu7PkYiCIgFzOhPwpdC5YD5rb8/gSi6ieChNxNjFBAtRhfYqAFFdc2Oj2C
D29vQskSNqZwceHpwba+pDHqB/FX3MPZiPgJS6QpS+QbvkhTy6aN7hFNHE3fib+1
wfPQqS17XS+mDNuYtnysZeNolNZSQ5m02BJ35zCaKKVPdMIMuZMZsNR+tNUCGOf2
24U3fPMR7Qtsd/IBvS1yV0vYdWTVbL1Fchdu0Gh8GOlhJPT3+JlMAVwVT7gZBqHt
URVOYarrkAOka9RQIOdmd4+SOoeT67VAurO/aVgKx+GUA2c4ni18NiJNFK/axxbR
/CTr6TT+l4Y03IJdUD36bOgtUIim+s6ageEZ3dV6M2qbV2rxfT9kZNMNUgYLWfFk
1s184EsBz9GzqhBKMwvlyt0uZxRHllUmt06ZljTeXQLUgI7twOJSypTjcJPazKkz
JQSTMcWFwqKDS4uMvNxYHspxUemu3RdbvRcBBpIlVktiAurZeeG5TzkYRjwI0fSs
KVUpDNOxqFocMMOwtLSF9G3AVKgeKX7YE2VC4DdOJlJ+atyu4aZpcqr+2GwPpzz0
Zmh4n+l8DHHEQVUG5/cS884hKOcaCX43O24CDTYhuQodsS8U889GGcAPN6uTeYVq
nXQ0QKF00id5KT4+Zi3aIBEUicz8G7fTFynpZTCZN8vytnB7Nx+HWy6HrukiKpg0
Yf6FK0PwAbbF3RSlOsREUMZb8Z01Anu447ejqE859B3LSEGxqYA3WoSOUJyq81pd
itX0dfgqf/Awx0MQo9C8Yd70lHdsRSvcSvwaLkCl0bC3T/T/tIa+973htFjgQshh
Hi5MiL/oQ2qDxsfE0l05AshNU/y6D12eQ5cU0TvKwDrrOmIO+AbRlESoHLDv/YDM
HUjYoZI8hr4jvka7PH54MKACoyc38fFhkqb96VDe2pFyHd9563ovVxrN83Pu/Ejv
Tw+ayoISZnk16NrEDNYUGZdprSlYC7KpNLSKO/l46LN/kJfT4PbaD+ueXGtsh7h/
yTzRh/pUxtGQtlei5nb/4sztfcrlA1e6HrCr/9f8xnR0wKgZUf37EjcX/a83rM1y
bTeGCY6j6Ay2I+j2++DVq9SkyOo/WSf4bIrHU/CsIVz5mXZ8zWtxdqNYa/rfjlBX
ymt0ZvMzWnudDUTNtlH7rU6VAzbtvz1D4Pl80LC7bRyMU45PaHH3QDpoNxWA7ySH
4rStKciB0eLbQPf8fU8yJlKqfhWnDfz8N6XQr81XOex4ZHFZH0frgbFHox1nQ7aI
RjNZX8/Jg0puWTEm8toHy93S9qtIibXVabeRr/uK3KpMJI0uPNhzuUK4WVpY7G1B
fP8/Mn8kTbMVIa1wkRN8sBiQQ4F6D0rK/ti10q4BfFtAGoaIefaSeT9+URvBFIQo
WEj/OEcb2ujcUs/TQsMtpk366I9b/swEfMvfQ0Wdo8JGZgJxx4dlgNwyg2S3cnMl
JtCf11jLw+vZNPhrBbd+bLtJePhPy1iA5Pnsmtks1Gx5ed9j8+XL3Q8WqF0AN6GM
dkSvNnz7TKCt8o9y/lI8Gj8Uo6a/RlGfPj0o83fSDjvJlVkNeKoNIOCrcVtY98L2
0EllHosO8nG2tVzhxM6c3/EiQCOb9p/IdkGuLeEPPZprywKtydbclYS+8tfLbw+f
SuuWmD7SE3VajsTk8xSpnn5GFJmi7+EpFVRUlhbDRhZ4aHHtPZemyHVmV7fJ/0L5
CkLYkWijS9fC/QQMh/9NFo1TG7/yjDIoGZfzt/3QDQqdB2PqFGSgYb9z+nPJONLU
P3Iu0ak5ULQzds6E36/iutMpn+1Nlp+28MNpIu/7vrMaYFbjOG1SwISIXnMT8zeG
2l4FXTPKkVirmLF746HLdtGH18X3X5AhCp5ERg26UbGRP1EUo3I9kRlrJ/FNtsFu
mickDMd4lnh3wk0GdJhwwPVbJ85y5ybtvLWl2p53nTDYy9fQw7K+R4DVGk7yGYe+
kTMkA7IHXVlr6oS+rMOAITrGevKJqKWoeU0HI1ANqfFPPO4abffq6eK/tZGOQ/Gs
MPkAXQUreJNLX+hGSMis2mouy2YW+qlEmjAg2n2mET3PbcKD3yCGADBTDE6S+vyf
vIR9jab5EZVRIWwBqiM9zkJtq64dx1OMJXp7QJeISqbRe7YV5cgAm4n/4WqsDBOI
oT/cgzjaJJCIYs7v3SfrSm+32DGiSs8cHD0U8Nbl3sEgi7o2PO1u8YPncj7kPE5Z
H3ijgMVGRVCdjFs6QDSky8LDxEuKYpucSULtDyI7AI3aFpW++7vDhYdZPkVR2eyy
ehoPoX/PbU1g+0szY+h54OFACI0pxWlX1pSJ9wmN7K5h7iaOuJctglqA14FQi+HF
cR2PLiArZbwo8ZUDPXkljPUV6Z5Vvy0zZQ5Kic7et+TV1M+L677p2rm5aq1Zo2Lt
DZVmrH6GbE2I15X6VAZabfkBejSsGTujgxH5pJTLjA/fgxAJFtpswi86hMoNMQvN
PhtJTiCEn6jZB/L3qL4PCBsrVTrSZboDekm5kJ0V5EBwTtYtGXzofHudKEyK956x
vLXwOPoHR68VBgmAYs/YP3v7SSNzOXbMkio6dUjbgpbGv6A6g4fWknwm0z5U8F9Y
yrt1FPJoOK+mIhTURbepu60znQJwnB6s1RGz5JrtFxkeFy7rSiANiO6JkxGrlMny
CG18HQKy/86yyv9kBY4v/3dHxEoZ4yoDmJPL/ihdIZA0X4r8m+3YRKu0wNkQ3WWd
Oq6ZGytHXZMAyOVjWxBw4s3K4+EOtkEHzFSULtNDfmeiRiiHBnWe8UCyKthvg477
MgeS56ujM/FB/jQa2Qou3Fn9iB3JU0hdngO0xSZMhzrld8CE68h7EFtJGmHQcUuV
OEKQEfS5bKNCxrs4Cf+vqtEMKFBVHfEqMlHAyF3Lzkmd59aGza8yZo0BZR03HKJH
r8lrudUWJkI6CQRbYyfRAxHA/5ZYpddA4GK8W7TnX3COQMPAhhhbccDSeTx4AFRK
KNfSTJfxNUDg5dGI0JUSj6UTVQRZgp5wuISvaE7VIeOBHQmrCaps3FCfGK4NS0Ro
Me0/ruFaXbBk4OD/LNa7qEEkrqFYXiSbgznpOcZiUewctXPlAHxRr38b0dFgkPqs
BStIxT+gRcKt5wNpnRjIl0V1HA3/O8yHv73jdP9PxPWAzryIn5hUp1rSeZVzx53I
KZHZlC1wp0dKXrZaw+WDiKYi7B476MRTzQuKowSlqjhAcis0So0BlwX9SafIGAyQ
Mfd0D++ZKaQus96Bn+Nmq8RhK96hj76dR5tUHBnTf1x/ac5Lc0h5542iZo/JOMTJ
jKdNG6StZ+fUQucBy0QwMAuUf20JZLKHuEKecehpVZNhd3H8flCUZBDFta9w/SDJ
BBPMqJxM+o53pWGActU+d8pzomnc1e6Ejqneh7+JL/MFjGw4ohSW/QLQfR2rFrDr
qUrdYujK19MVYS/LOMz0rjQkeyPsrN7lWwrnUxPYv/DQVBNuQcfTX1X91tCRjdIC
W5m48fvC51fiXFEV9cjAP7x8NWhHmbFnETwTqLJLwGTkEcB8m92ti8DuOdFzvicU
4TEZPOKkbp8LiIMoO+V5VSJcYHxf4iQUCaE82E5enZafYIRK4hEPnNJzXCE5jlhY
5yNZLQ2lPqvoJChWz+r+kQKon390t/+MDKTjBhIE8HMct2l5hkPcAzGbQagCnd8l
xaxyy6LYRZyW60MJz1xja4dRobz/6B4sd8g9SvRTnDpsl9D/NDviQ4hcbYGACIXX
ZHc9RroY0rjYzLbZwTEhZZNMTli+rTCZIiwWo3hV+jgvMZsASsdl5hmp0fN/LmyU
X4Ljc4XUPihsGSWE2AcYRZfqd3Gc0qAfa/q1SO84XzoF7U7DHWoJXHwcCyblCzup
pFbHfAnZ0wskCi+Bpf6D/lCeCtEuL1nUFk754utxz+wVUHFBRGAujYWglX/4YXfT
5WEdl8W+JoBR61yUJNxRL2B77APUjfp+Yw72jBHDqtzoXO/lTOPIMkHtrj4Dma+a
sC5NKNeHPNMOB/QrzPoCsA447JGEJOP+zrGFsH1T8B61fD3egtvMdxuHvHBw9dpz
He7tkPS1aq5LbIYRSs5tJzMjpdt/G1rkHM2VNZy7ZcnijTBai+KKlcyKACh1MOj4
0jfg6TyL2iKdxRm+6U8lTPopICjiSw3Jb5XLdDJc0ladRTjDc5JJ8rImEn5SXRGe
f1U045uUb+aMqMHpQmk/08I7PQ/fpdw9T3WKi96km1boV5lBDfWiH/vBXJ6GtQf8
i2E8ZvJkAVxjKe7PZGz0wAafUgsoQugGO7MCrHZMndqvkVVqIy3NIUx3LbqrKYiL
fVcGhWi5bPi/8OBSLUT7IlzoAeoAOOTtl3WgcBCDO5shYnbwBcOQZgQr02hJf5GQ
DNpvWAOMItQl/PVhm+S1pIOWtCOnfunQSWcpffJxuVwigEe5lQZ7ufquvVW1sKPI
RUs1PGtZFcLE/Qc2kS+furZkRqnCo5g0VibSuvURIgeFMvofUP0m+MmrVbOOtw/F
h5WuM67HBJBQhHnj3ojFC55GBg95KzAlj5MGHLDmgtWDfYje+hQllsga1F618Deg
xyeklEY46P333pwZJxuECqtuL4ZSGk8K7dmXZE5kTyc08Czj1+eSadgpciO3xa1V
jj17GJt/zYLshM5aqnJl6B7LsmI0T+F0FUbmPV5k6Nd3yhjMeqAUUd56477S9wxF
Fs9GXF+OBwStxk9LA55fjIdUv+TGu3UzUrICtXRSpKrEXbjlP8hnH8Idfb2AODVC
rue61US2jy6sSBdJ9z+rXBaoApHnkWVUByURf+QhOAocdEfc5J5mIq7stlZSlDXL
euqNgti8ezSSCQewCuyD4X8wmd0dpJOucd6QEm5n/v46DNEPgtCu8qd0rUG+59DD
+eOrHkfMrZcK3UyuLV2wtYV/AW5ZD0Vc2EUItam1KlX0c8tRH8IMlyiaUbGiTm0y
CLYHZ2hOY0hw44KRCL9LplZJqoirMpVrcGfXv4b0EKo5bz5rB6/+x/HGuKIb08v2
e2E+/kzcPQjwViKKuoVoJEK15af1/tJaEEyRZGIMq9z517EfV+5fMl0eARBfdOqy
Q9mcwwYH7ae1VS8mT2LpsFXbmOI4Q1OXFMmt2UHEJeejh7vaEDJofxulMMNm1De2
IfezEKzfFrwdm6oNXWNYNiAcggF2rYeykdZ0xD319XiRrFL8rh/90J9EVN13zIkd
xurIZEYjgopU/omTa18TYulIxv74Mgg0A8uBXEOiE4XKlpZ3A1J3XbNuc0s2jqvZ
L87uyBJ1+21gNo+7kMKp8ZREfVdRtyHhiJfQ2pR/r0mKOkZOTGyzuHqInc256s65
sL2yaZ9TZxFGy9dKTyMfJCdhDJXN3UwnXpc1PLI2OnIu1jXW6Lxyv92b2RJ97xeF
JopFAPaTky2b7/Ctn2tliZW80mFE5jkduV7ds6vUGiCXUtNE6Hm8qnwZQ6BoJHWI
lWOvuBFFEmmmhLMwY8ktUTmuVngAGJ9qGJlOr8llNw4xfIa++x7rIUfd+G8HWPWb
lwwZLOvSEcVwvG+c2sZ4NLOtpP7mWxxsoAR7/eAWAD/2h4Gsk7QuqYO4NxjW3EqE
c/dycYDeAMmVboyPmcUcTF5QnCbOTFQWvowrn7m8TjgsPCOULwvN+LUM6F7GaxVe
rl7asLspiDolFIeidyh1JQ4RntfwzrW7RrxL5uHTl8kWz5zYlsawp20bxPQVROuR
e7a8Q2vULN7FTqTAuHKcq1Zjo3IN6uvObazP6tLpb3HG2zFmXv+C2uY5tEt7VRSb
W9JdlzKgEoz8NozS5XsKj0pKwaFAlz250lknHnWM5zcFsvo2XiYuEHr5lWsoDAb/
nNxMrRNIpP5bhFBux4PX/n09MFCBrGoXay1U9IvTzhhByAx6Bh69p8yYiOqQ4FPF
+8aKGW+jlujwre6PO0JcomFw/GNEJmpKE3IIpbEijmlU6wdmUYskWp/mtFoNTu7x
v5umepwmNTi2CCsgcTGEeSJNChP2mlrUqsBINg4cwk1L+UJ75CHszwqsduFrOPbK
RprJTlBn/O+8r6ngWWydfo9MnDhtdfI8WrW2dmPwHsnd7T2NMJj1zwW3CJHkEWpn
qLyy9zdL5XI0vDALXsuo9XstZVOxOcdaFtGkTEYLWJbni3lEWgJU6CQNFDMdM55R
S3oTCxhdGy0eqbfSSdwAhiwrnoGlxOlmiNKBtqvCGK3kdCL/BdzICm5gr6X+nGOC
4Lnt7YgfXexvxwdT0asUCL7/Lx61jmehQEvjyUJLxRr3DfvlWOSJ8nwfSHXnJZvb
BgAGoRCjj3RgfdxFpCjiNvzp+fTliaE6FCCgSVmQS/PJd6U9jtMf7zR/gsPh5y65
NXVfvXVrleMIjAsyX7ZzBgTsErpxLu0ObaacMKp7cRbjN2qskZ2OSjHK+9u1MmTC
m4i51qLA+nv2hHIKSlKKcm1Wa3z0fy9ehhsAP+b9W0ocEgfL84wOJEdiD3yRpHuJ
hzsGb5csl+4ZVrMg3nQ+01WRF9D0mqCxmR8Xr7kiN51FEJDLdQv4xECbM/kgBSH/
aLunJYBuQmiddfU33HZJrxAvazCrAFdp33Vt3Cf/FJZDQXM4xCkChKtBrHe9rfHV
pp4g0yhUGmpzZrItV1gQ0i6HWc7LDZNaGLO00VyFmcAgwxkAjRzreQKaD/VJHi/U
Pg8oP23GZYEb078Dogs2TIkHRNOmajg6odjhvg5oGN+5bLUpXvakkCC9DNlA0uHu
AVC4lwSlaFftLUwDKRpnMF4V0CXPOW+o86Riux1tfVuJi2CbF+SEApwNAVpZtqkI
zswu66LCiX+qIEU4UbbLJSXv9pGLY2lCnY0b8j1VoW/uZWJ5UZYWbvQmJdhjKjpu
bdhtcBsguveCZxda40//EzjvEYbHLSiMFuyB7Z3es4uMwsrzS2TCh6vP2ybF1aWH
jJ8IKTrWwUJIT5e7Dxj76CnTMO4trqv8N+Q2riI6J++488gUb+dwpjd/qUJ0SKyc
lkdJt1Jp0C2ptu0D5wI32hl8wb9Hs+miAp0jV0BH5dteaGqZg5QW+Ggj+jjnbbMP
UXMXLKFbrvLL8yh8pIOIDFqbnH85KnAcsjxzpnBR+3PKvridl6UD9ASeftmsSoop
fO6G4J/o3x04SlD38jJ1SOKUmnyXvPR8St+zPNW71bLvZFd5GmHB9MxeUIkKxRrt
kisB+acwuBNB0zsV0I1wGbK1z22C7l81bbnYce+1uomVMPBjDDxEARVxsSjpuUKO
5GUaaPE84ElsQj4rAmv20QvO5j5U0JinLodsEv1lJ/Lm8VMwjYuLBO0BcQz+eHAN
k6mlSi6mfl6ctZpifXzqCyYUMGdfdgYqR0xTxaif33DxWNal0esZDWxkajSy1Y/N
dZr+ISaGHbKwZKQCtxeSHPLVPwC7ODfultTK99sy4fKFTvs3Br+irvQgDPdLfA5+
W06ilgvA4e3TehG6Vk2TtQIXtTqvvVIExpWQOxV4QfvY/8MY6QF0QdoVXwaTAEDS
ZL5WAtUmGzF/SCYWOvC8TrRdXnIVgxd0S/s/nYwJ739CJIuG9czUYPAA8dNCcpbL
IIaCHZig+wtljlyTR0hKeVRi1cyy44Lp4kwi/Pd9J/s+PUkE5KBB+OyDcaZA4KO/
AffSwSM0l4tC21uF17C0Dkjl6egPrtAH9Aw8bPyDJHOF/aHyLB8KmvEa7XGuy2id
loeK7xPDwE0GKrTPkwFYlCXJ1+YiB4PVDTZl4BtPzYiLk3WGHP/GDrFlH3FB6FDS
FB013ddywpty0QSLApHjigWGbJFirpwwYGneB0pvPmVRxlfAJwIReBbVjyWQTQjK
YsTcziqpIHDpknPKfEwl52ylD0+Gn8YtQFxfGry9fpuUcl4Iqfr+0fvULpcqXJtD
sqgpFYDvmMvSavEZ5nQ0yLzEU4yRD6iOhWPsPzGWjbJvUEacsP0RnfLvNf+lORvP
Ms/1mFbwBFa2t6LD8GpOFKafmZYjUYp/Cj4sawo997U7jDQA7XckXEsqFn3lRisN
jFcsQPoxMkEWQ0jOdap45/Xc9lyTb+Q2K0u5B6MBB767dskcxh6xCgZ8OO56IRd9
4k1QWSnu5+O53O/b7utlNoEzPq97liQHEQHFX8S9sa/AYW3RE/4qsEibJMir0KE0
NFFpW58p2QoBfTDwkaponlh3b1aHmNhnb4iJCbu1HAg34xCs6bL3eTWX6d9Pxepk
qaKRR8kiQEvo3Qqd9wHd7hbbDIDSnWTWBP6P5Gl2xChC7HpL35Ksn28BNpr8JaX9
31tROc1k3UEsxklswxpuKq8fU6Jqwwcgr3fB5gnVyn/4h0u+z2Gv+SJjM4GzBDZv
PS0fiec9bsrySvFu7o3u45mLuINqadrTQ8P3516Ch9zG/53TcgIm4lyIQbGQN2Ys
sc4DOn3+qrHLBFxGBEK8gcRTNyD0x66FW+DvMnULpHq3XncEScUtyBzbVxU3GHRr
eH7a+NCiNKJDWa5eXJW+VNTka5sz8eE+GiSJ6X/GD1YUF1SEENviOGbPCZzX5vdt
2+67JIRxw5cd+9pLdRk3N3WEjW1kzgfATg5uqCrcBs+UD2NEM9Q5/wuAJSF6Z2+C
C8Xc7k7y7s8L9mtWHErdbS3Nfw/FTth5o5eRqbAQYjjIV18zRbw1JxEJiU44MN5D
usqs/bDXyKe+pvswlahLaGg37YFBs73DFXmwt/QjhamINXQLzaUx6Sz7LmhqB1pg
hudqkdk4XgKJ0YG6Hd6O2Mg5E0KgEcvS1gFt6knOSDjgmciB9eOnCGPZHsiRGR9r
Ni+xA/4BZUBVINRBuIpmjqfHPd2o89EUx7iCLDRcDmTNhHHluq5iPF69o2FJH7gn
CG91C7KZoxS0qZ31dql6dcp5Rc3rTQMcK8A0AJIlv7O0zfLXZXUXPMriitC/PCIr
q2OQ9S3NIGJuqsc7TK/Ps7f3w4wWZP2Wh0aaf5TWzcSHxw2rvzTzHA08qYzBAJ7u
PjMnlz0ClnKgtCOhSugT9IC9UC90vUGH80RnbmfYeIUslIIFFFoe+BM5qByj7eOf
7XfUosLfQAiTLZ7rIGsPjkI3n6H4D4nVQrA0/NeRXvofJBdjFASI1CxANfe6F81S
2zr/JXrshUCdl1LmAmIlAN2/H4crn3+NR9o4sRSvsPw4Rx/NjOjFKcTjNa3MEFrp
k3rkZ64Qd5LwheyU0ZOSk3C/KhhZzNCVscQoO5I7bekFRJJ36ONYlRhRHnp9YPOb
4TaXptAxCkO7DEj/dpQuRL2SRPmuFSOCs5bSsWa7AkHdMye/fsrwfoJZEdTJ1LTE
rriev9pcUbbPfCfjAXUDP7nXWRAQ4j/8RzXPLCPCZQpjYI8g2HBQPpYqEoRGtTQz
J+25XkkmFOZOhRf8XfZiT12H+7KNYDoTNuhW2Hbk0LXGb0qkg7MPOSjlVIvZeceG
sFtALsfM3sepLrWy/MKqEl2m4Vw8V7eCuRjayPU85Yxb4x0LKMO7M9TyvJfu82YB
drdbHA5f3U5sDv5pngsHsfX3mXXh6NKuSl2jh7mowth6BKzG5s/cPb3eqCyKSxMb
+/F0v2tR8bLyIsxUGAyD2QxkSzsM37n8xeTFbGWmdF8hb2oxlHAfCkdYPtnaqVjw
fNsua3vM8ABGuJ80JnLQ6xnzCeVnAxPWuhz7TwHarsCjO5Pca8UkMkcQNNgTuCqI
K2M+xlJgUksbJYiEfkAH6XKXTxYqUa0YI0RLCooukusKlsggi41fy0w9KF7fNpzc
F9eN903eRi0hu08B5xPwZ8DYFVmrc2pvBiW90s6vFYta8dSXMerpkbJpYiUMED5y
2Io3QJysebMnmlZxrdNHnssFfSZEw9TW/BB7FGERIk8MvT6SB/ovMeODBb173l5f
dWwoHZV2s0Ab16QJnBKl/Rq00kqZzyfZXwuoQFL0XVWb1OrlB0cHJh29WotGDduv
1mZYy2ncqBJaHu73QMhcjIIA/Clwet/yK8Tk5kblhVdRmSRtGqyQREpCsUxQ07OE
hWMCdFUNjN1ANLlkwDlS18FS4puBc/30LO0CyNo1FWOYlkGUefSUkXb0CM4Bvnj8
0WInVC+pdM1h3omOVn08k9/GfpESz/CXEjpDXgqAgAW3WjMDwDBxWtdCASYyo+qy
OGqbP1xqX/gqEs2Ii7dBr8KdbGLgRTTTQZklx/l0cFUSLZzBYAMmngfg/tna9TXP
Udtau1/D6TdW6KpdrIpecFKljbP2VVp8JHDsHkGZYRfRlioujUaMbyAVpmPyWjfB
E82WAwKB9XKRbhioCr1wTcNsdm0IUt9mLaRgwuP+Duf5rvlmchG92EIgVG3TGVpV
vfOjTlNRlGQU80Zrfhxro3bbDxvI9q4lEjw53rZ4ZPx3d0aE0ROtldJ3BA6FtLzE
M+w2OxAwh3K4U9/xyCs413eFxPihA3snQ8kK8nafFWZsBQDImba0put4IPE1ajoW
WbUqo7YSJPGhkaEyKp4+Zj0eSILeJvmY+lB/2n03JV9BKv5l+SNbAP1vl/GNyVFw
VVLmckFU2rXfOsYmb+2KJzldjh6ZyLzBaCv8IAeDw7cxpawxD4U6c7NJEvVwyvXh
hQ/uAfYXv3kxITywW5oCRRGpxh3Ya0f4htUzVVENnJQZmNpDVCkUQuVHNvufcPsU
diQKYjuKJf8xDXVJg85YPXHIZ0bUZpBVyj7zO5Mf/IE1btwfcKpFvu4s8A7dkG/k
Ru9OR3vNW3OCAdbKzzDd2N1v8AvT2QYySfTZrVhz32buBaUND0TJtidw9uVhwWAp
mwiyVuJvz4xlHAiM65kclJKreoPdZFo8tgvVVEJ+0DYPbnNk39dwc+lvPE2VdTtX
ZB0f3NTL+fbe3gB+LnTj5FZJDUmrQsRmos+lnVjQ5D/8V0euiEJw2EPhpjh1ab8H
W2YjrU1a6jhW7s7bCIphAjI31/VCSqcfGyXnta7+zdUTjaXwj1rtLZX4bnUuaTen
Sg9r6aECqEL1gNbi2H5zZqfvo6NrrPYdSinNUmD6126tfpdQx0rPZM5yChAmOn0Q
RD4+034t70gqoEboiQF49Yx6wFou57G0I5Bm2nSBLQWyat9r0IbgTmqZX3k1Z56a
YPfXBrpqFf68KGuoniyAPCeb4misIR9Vteh9tOpIjM6SzFQIZs70jIC9p6T2iDps
82jPJah8oppDTIgcax4hg8aMZRLzzipBm3huhyYi7GZOwCkiQ4QFuQHBCuAuYydI
PqnZaE/vfwZAqPQxf2MpBpFUF5wdiYPTp+9+J2Rt2Gch1+voTAFQpIvMsdiZp7k6
Vm22KQUPOR5sf2INJLhh9WvzsfJZt74ZaWSTFdQufn13ai1Bg5yOQvEyy+NYOc5Z
TL0fptgCXjv6I6pAkdp0FuzvWBqEBOrWoYAHIfubQj5nRFxPbQYAG25TPt/j7R9Y
HOwVyzsOofbhxIMmrvVNPbdlgSX3Kq6Hq9+XTWcGrPBjCmKufPLJaTJl2dRfA4AQ
/Q5D/pZY6ip46BF1zsKJXvjyBwvNIKVSnA19zMc/SozRyP8Bff9PAEQyk0Yzjtz1
YmGACGS/2f2vWD0raxhnMNHLv9FjULxKzWfWYs7MkJQSrUIbW1spLCZ1bvuUkshu
uxMfGl7gS5H+gAgRE7nRIEj2YpXMFfrwPGN6SBr61m4UugEIAZ7AcKFnkT7PuWtw
n+AZgJD3QVJnrFxUF/M/OB8OH5ed99sLFUEamCeSMXuxJqzU82FMsSYFza7ehdYB
twxITMDdn3bDikSQjPQgGk2qb3JZmu5vULmY5KR+tPeUQLPnXY3a+qQq7WeK+z9M
wQzbwvxUg12mlDb9ZBxn1GYqGui9p6/UXNULajJMqvzJB2PTaicv6ztlYdf1VeFB
k9XKmBmXPReUd5kvHjy8Zi2uRsV2fXLxEvBwX9u4yPNgOcY5HM/G7P8HJvPAW3JB
HrKANuPFuzSF/LHX5fTPg33rNKxKUL7wwwDbJUlRIVvdEaE20YtZCxQJYyFjvfuq
KXB6cyicFMlz4J5oUeTkBOPB0WUG+ZfjihHs7bFz0/uCWfUClPS7W+XAEKK4Y2JU
E1orytYCZf2/zppnPE3l//sAqPf1n3Kf4ymB088tBgy3a4idIUtBvGh7LqFYyQz8
4eEClZ0w3zDpZhnwNpc6CN7ixm2hlWGGsNnR9dXeRAlKgBgchGo2S6eDYhLsnR4a
nJrHs12NuOscg2m/+mDYxWmIyA5lSqa8Npfg9x64aYUSHveQaoSURFIRRwTWO3Ed
8Es8gL8HKS3Eiw4WtgJil04VKMLDrnfT3/Ogm6BkXyYmdBChhihZUdA7N5QRmw8C
xrx4oGoEka0GZJ7JeenhXMeQobN62iEnwBP3UkUVMBv/QNRjSt4OIcXzECvUO9Ip
NURFnULs5f1+chUwIlft5dVz9SU0aKvtO15Bx9zLJk/PDoBuY+QqN7ZgIXv7PJVc
jtqLxltQVtXMH7oylkUAKnJ0Tz869vVQ2d9G18SlHEFaU+RQVtt/oDzO50ccaGrX
YOjZlFrqXSxtZLNFribnX8HuB2xk9ToTx28FPnUijyw/DDI+2/EpUwiMPSuI8CXW
0x0nz/eXUA3LJkxdYKFGXOM3us2Gj/fLwuMvbw2fBH+p8KvLtc8xvcFV+fJ3CSc+
6nDYJPzSkCz5y5BoYa0h3LLbFX8n+HUO0uxqI20Ur1AxZMFTobbqu9HOAIwMAjyn
HTt+yGMO5/pNpIis8uWvctgU8NUcA5Ii4qLkQ1rs2rXYIv3FAT/t94UAJbq/fU4z
RZcsBeH9WwsiQafb1a6ovoC1ekWHCw7uY1NZItUOdGkgJe+wrjK3FS8+Z9JyQaEX
28VakHG0Sa6l4Ra+6KAdPDZboCmk29WT31CfTCPYV3Ntf31+1HrW3p1LDi55loXB
aE8dCOboboZIMiJSkxlvCabLEsjh73grttyonAds7dEE72uMRPLD2baXb54MOktf
mm0RAbS+X/J1Ds445h8GDMuZfDIx50q7zF2u8BU285xsTIzG+GOHWLctlTtkbwAh
TFrttU8VW0If7p+8DiNIli3zPIWkkelYIf5q2ueujP6fE313Wq3oGF9UrIdeTtJc
JyK+cKs+a7jOEkRqKtdSy1ql0SwtDm52lMQzUTmrDeTAC+mmfudZM2EY8gOmwBlx
0WCJTRFennZFQ+qyD6UGQAj0gCLTBWBEoWNhihhfQ8FUE2Dn5Jsrc7m++8SM29TI
lu9/b3kWnDicSaq2e090ozTp+aTDKeQDTS13Az5oqEHOKqt5Dlr6EeS7PmvYnF5z
ybFwGDzDdqps50GRG2RrQ8ZaCn7r1Uv8RKKjMMnFzyvUEgVfCuw7J33qoSKGa8kp
MclXwm/7rzf99AguXxHX6gjvJcXoYbmL5/nhOOxVi7xxjPhq/E/VtzR7dEJkIO/Q
9M6LTMxJzFIud6pVYX3eflvA5hU8gTZTqGPU6exDFeNrf/JLifjCt81RcVc+fwUP
XnAiGJdZU7IK3QseZGb9iAQYOErwngI36pLKjY03mLGvHf8VkP1jXqYq/om1VkmQ
pAayzHCqlFn3MzIMNSynlfneEUSdQcAMcqwdfBr5NCVmUvUJLuDX5EprjkHZn0Lt
1EQizawiRd6jlrKSKof+Ltar7OaAO7x+EcHnDIc2gimuSVeSpzCNFletKwwiPiSk
87U46ncr0Yhm0b1po0MKpfJU13mAs5zwM2QwuwOC3ELGLbYdv3BcTBgnKLAE5gQj
UG/k9kU8eo1Rw6Dn4c6Dmkr/atrCIWvHk+jXxddj88qhBc/r+yDGoGg6wz+th+ER
KyZoIBvZomNAkP1I7QtmNFS0+BkjVLeARD/6lCNj5GPLn4ZoGkggb2R/bjQhmkNc
5UL/yzDuK5CLTkKVITKPcHjZ9nfzElFICFhqjmeekbEKPk9vo58d32C3+L6SjiN1
rYdutXSXxpZjNGj3O9CAyrD8S1AqWou5C53YzmtqJ/U22dlAxntbbeS45OvPbWeO
dPo51U0cKJIfRSXVgkp0y3bo4s1FEt3yJmZdlDUrU06Rxmvx797SS9yrmj4TdG0V
rqQlIs7e2w6wH/U3WmJJoTncrogwk9Hq1hSJ5RfZvlKzlAKSgvi2qJLEueVhBw2X
lmF2bGRy21HprUsRJzr646kfd+pgtT6S0rC4iq3MMkeb47FQKctJtNT1QR6QZDCV
1je1oXeRUyLHjtz+3fWKWPoWTkV+ineTheG6OBI143wUd2y8uTjgy+8vGlNxmC4B
zaq1yIBiIcTjSUvqUcgxPVOcmG+BLAGkJ7VrbJd0ryu0YhAceMi6BX7QOTDyehJu
W9YYybbi7Sfxi0WKtVcPtCq85TxmTr/YaVBZD1B0MI+LTPuqpf+9cv8xzoNx15hJ
zELXc2DyIQ3Kx5GeCDizCa6bTfqnKuig2MQI+viYbojXTXlmkVBl8AfOah0bSZea
WlCnxS1m/OLL5H7YBOFnwYaFUwVBcQOMU6fRQM3LAb39fRJY2N7uhcOmhmuGjfhV
ehE1evHeLW4f8DfGZ3QZqOarrWGdKGgxL2OBSjUySUF4X17lQM8fG3YQqrw6ow8v
3Fnu7YeiHzMhPCtoRhbBkx7AzUuj34m2GZdBZkuq+zggVE21ARb5zZpm3p7N/358
m7Tyz4WM3tqTwx9Q1bk0yufQYiO6ZY0fRk/8MjSOEyUECUAXr9QBsDU5pCCkhvXI
sxVRX4bFABtDfy/TgahO/DjRfur8rvIcSZ7s8Tn0jxIjLrGQrG+VuSbXzDGxt0DH
CQGu7h1Ideyp1VLo2hpKeqG+lSAYKHIcdkm5yCFSMocbvgLS5w67JukXGNEoXu3X
rMaTwafx4VbmucTmxDaPSntsfsMdmjHDwZSf0QLeLOgtbaZ+6ilGW8M7/KvMOgaB
S9AXYfEEkeEvVlQfL6bvO4GxUGfDBppkJwNBJ2DvGstfzEbi0X5lNdtJY14pd6px
LtfYFiORAVEk4yNMZSj3gVJwF9XBXB0lxpvl1T24hQmeCrC2zONiZaEywOCdQkut
zByUdSh1AzPCKq4azUUhpvJS80Rq1sA4fHT6k1FZDOF0SHjsxPVBEHfuu3BwmYHY
uqqfp6q4I+q2FYgVqvdIYMeU39VpyTCvv8GaqsgjqUufiN1yIa8CEkNE5u6DLfLW
y+Itpb5lAwurHiXpx7ObQsw+eQQ8BplXSWNZzA3AQLOaUb95fIZaLmnQdaxYq5rO
iwQjVG1ioEZTdN3L2rJ2DtHcMwhOQ434RQoN43gq/2QGYIrH9B3KQS/dN4lsI6na
byXEhAPooYwmopVWBvFNrL7mRUDsISIASeQy3YPogqX0uLl5hNTlMj6uBf6ag/sE
XAXKmRKBnMDteffq1c6YVZoJd/9o7BOdCVZKEDc3mJP6BrakE+cY23yuDfj1rXsO
puJtFU6OHNBmboQJ+5p4+9uFIveSdxggDaanvwiJzN212/ARXziTx6wU5VVebJT5
RDxLHbW3QdaJizVEWhVwmhhWWcALp5JiyYArp+biXD9zNmlECZtuU0oXKu5uS0Tf
S8OKun1ETMGDsg4+QcP6Ek450COCOd65eBZi066n6FoCS9GjcbXm1SUpCNP1Mfbs
iT9eqo74Nwc6YsTdRNgERrUn4bJ4WoukMemw+V7llRLHnMMMh831Z2auTenBhbwW
J6ciaqOTgdjmNM5tli8mvc/B/8t9Zwo3cCTs2xFbd9KsqIjJx42nFg9YrATwRi8t
IySqYZGhKNkyqxw6NY62d0DRO8j8VFYL1S5JgLC48dJmELv4BwaiWYj3zXurmUxQ
gtl+/pwij/t9buqICnZzB/n82FrJHUSNGQswDtxnTYl9F2vYzGDqaNrT8yNq8xut
F8JEyonmet+NXJmkOy7DKR/mfiOUzSOMrrI03j0eaWNjxxLlQA7BLkLtxe00Y5zd
yyaLTdLF95IedEv9/eSmQmNQQl1GGtMTxzIln/O6wbW6Rm/kkpqT8Ew9Ncl0LwMx
T5uSAn6SEGAsnHZvbPJFBjrrAfUBSumRyCi17Vv7AM5ZDPcR/QsdeFtD0NcFDRjv
qBN21dG7LYtrHaJo8ttNfjEQ8OVpTfDz8wExeVwDrOKFHyG+Vl7jNrE0Tghv7WXX
1Hbzv9h0BJtNU5ncyu8skiO+k7qVH2af11rIRTrdJGacSMYNWGtK+ono4qVWii5n
oBo6PKg5Ad24GmkH6MBxA9YI/7ymSXGpz0ppGutTLMLjJbgZsHklChPBg3lzCaSH
/sN5rsWXgFKcIO9+cqRsqqHhCnwHpzAD2omqgAJcJbineM7g8U7Nv/4+rTeTHgV5
v2zacR1ektNt8W/hAhPt4VybEppj5bETUz26wy1XDTwmBZ/Qx1AIFsXRE0d6u8mU
GlfYFeDdwIeN8VMKGkq3WrzcwCSMW1eek3ioKPrmXOCX33Csu9+KgOEv6m368xdl
zi4Jg3iSAdnG7HpWSz7D70+7X9PcW2ifT8mLqk7G9SmCSZ8PPqktWMAxq8ouxWMt
+3RjWhCakvgA7fS78k81H/6x4jXZX6rYd8zq2/GoNeuvHf4Q6KGQqps/8n68JZ05
LpRDHD0BTZi+/aSRcLnoUUNnxEuGWshJxBy86H0tu0ZC4xDjRRSPyIDMCNoWAHAL
sMtMs+1mI5N+Mih3EbcKIZXUCN1NW99btqMHWr8Hi92ft8LO5j1pIag6XpJym+vm
B9j+i4q+oGDxU09RLhy8XOhkgEyqC7U9D1xOiszVLltFFFtoLz1M1bi93V8CEaue
uDt42kXhoS41eC8ss9qAoLcwUoXq1Q0bzUkhj1U65RhvKxrwwO+FFfGnBo6FhJxR
CP54KQhFnGSNSrew4HyICUiJc3MeEtRRVR7NdBoWjqNGfZ6vJSMbcXUBsM6eMrpF
3te7vWbd+QcjsQ8EOdaXSmqKpMdPPGYzrtY5qNDee02n1XqD/2E2TDHDlZR4zNZ4
3d4MZkiATkNnLMb90MsifYu9FzqIaDrQbMyQnkCANSZsagdZMWriLKmvVctmduk8
J+fumxaA96zkoP5DKbZMn58MoEycaIgYh++AAkGrlhspbqBw3i2+xEDMhGT+EA7b
pVZ9+Pgo93Kb6gUw/C2J+kXiN7hUfhG+20HwNnenxRg0IURl6gdrC1vWmOThPggs
Gpan/eKVAK0kCErShkM99JISVmVNjuieBFQnAxztC+PDQhsSm1vJwvEZRNgOnP7m
saA89KoEy/tVP65gkA3BSSoHWOm5aI5d4VP4z6KJo033Qlv6hp9O4JXZvLRP3ev7
nnlcB9XyN60m5nZRuZCamrKN/BxDbCUSlyNXCdgTeoTbBopBOz5iAjKq5n4WTUJV
5uXQ+gyn5/WTaownpW+b5CWYD7pbwPMJvnQumoFT6+6zvXPzSR2Ozsuy3fGjl4Bp
/n9COr0WVyYXON1KxZV0vV/XQ6Dl9qSMm53EZB+MWkxxvwuJ7pwt0l7maG2MGt0T
G8G3tlDDM3UPav2Q5aW4e3BiNIfjTWCEDNt3kNS1Ea56ZGxCPOzN+8yRbRjxKSEh
moOWj2fYQf3RGhQbRcRdsEfagwPjMcntK5vJxT1qxbmUsBN5JLrW68OqbOcjwD76
4VqWjxOhV7ZkXpRJZPjJLkWjQSwlzTSBMGlvi3Yv890iAuhlpoTUr6AZD2NuN5Eh
RddgFE88ZhfHW8sBA64pvmRbvAisskrZaBqVktZP4I0o4LJr2+5sg3ptrSvy2cin
C4fvrsGZ1LbmSmUKYSkxVgrGU7DBbsOQb83o1lM3L35LWwRmochHNeUjld+uvfAm
/+HJHdHiYPBh5BiOjzlEhxfFDVwQBA5QkJD2sqgjBsJ6vcqqSqecFtuXXPs9NZet
V+4qTfR9F+nWuoJYXzxK1m9ybiWqmWBXgBpa5oHBLqd09UOxeWardPI85toH8gRN
O8QERKawKrxEIaL7CuYAArL1ReuIbr/xI1HB2QJLVB8uSm/+LYpCjZcEZPUsEY8r
6fBmoDwIrOEw6QiphNZ7ebyAzBGg6FHRWJplQTkRRb4Z9RI4sF1c6jyzZ7Jn103a
maPUFxLmBR7XAcXs0WpMm1sNZeKM4BFFrxtUwqAqlKk1jEduX/PLkbOmyawEBJR9
iwoTPBNyOv3kg6zeYzCfDs2A9IwH/p5DQVoH/cZFn3kopU0PB6KwyFDZJabwxFxq
SfuXpDax/ygaWke/Z4VV4gTdbJvLikgug9g/AyiCvOZiaQyEQiKzz/dPWBWmrDV7
OAWvI8Uhem4zCEiVp4ZfyMknakfsaQ1RcDVfHM18elW+UTzcboI4OWuIHhGOHfOp
Juq1nm1uLaPLc6NOvXMVf8hsY7ZybXduSguhkVGIAUMZng59NXmrqiTGWu1H4nmR
w55aaI/gldxifQznk9VIcieEQ4vrYPvqMq4DTWGsFSKYnxX7ugFQVnUA4m554kb4
BXyYGE5fyJ1hZOhkskFMI10HfSG8A0dDls0tv9BlohB5RTNmWxqRiXtO3eSZB53R
CCeDRoENTy76fxEZiLC4fTRXYiBQN3uHb/O16XIpRJyp01kJw4zbhw7igSHIfgrf
yDuXWr4b4sTciMnYSgPUwRDIGo2Q/3xYy06NAYvPgoswU2H8vSVXztaa/WsD7JTb
pB5kb3Ao4+DkCiOPPoUZNhjRvgYEFE8kfqr/evtSLEFQkSNAK7ae3wLi+LvaOTr8
NYV5h/4kJnno2NUPQeoWwp3b3kBajDL1tHf0hAsZ+phwLVbSCgpDVhZcXD6KPL5D
VCgBKnzXvmm3Oalhai1cbCac0uSvMaN+CJSuXlrhrGeRXNAehtE5DpFc+HPxLn+b
3hhn+YFEkAivkt6ifAvP7pC4LblBUAaN85COfvdS9ywCx4KxNFygahQX5AGi2l0S
QndngzgiEt16zXQZ6vopjmC6djuoHL3QFDX74+AA9/Gxb3TpmL9gHjW0Q52OGAcf
9UPVi+qDK8bIlsG2sBAUdxxXTCyw5tZEhGnaDCkrtcP7s8N7/nCM0jMETBnAIhwB
Z37B/VriwQXThQpSArLE4JGV5FFVIoVHvK2+Ri+ZxkIs8EPMg5wo64Ls3N5f3UAE
MKObFKnmrnJOszZ2DnxcvaVEP6Ocg9jz6Ui+1kcOTrMfXJuARdGwuzjJbNNnR6cB
ca86T9XnrNl7aC84C023f3qf4xzu9JTyQhZHzzBy3oQZ7IBUCwsueFXJ//ezfdPB
UaruUym5GR+DW8i+TcrZ/rnYvljrgSiJLcFCh7frRQMorxgtkIj2LyZHVUzM5/24
VunAPFTyeKBO0/lV6BUAVV9wQ/rvsulU/kVad6/bi9iStSjqY5ISuzt1Ikt4wngl
tgaXM76se8bezKfYtgqaLwmsAs1UVPl5Axmz9XYAWYA=
`pragma protect end_protected
