��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�؆���o��9_��ʵ�Fꙣ>��IG�;�bHύ]+�;��� �O�5�=L��*םiJ���B��V"�������Oc1]���?�-��7CI�M�*�-&�i���x�)p��$���i�%��2Pߣ��K�Ptx��u���������V��],��yo�k��?������8�G�I�_iঢ়����; �̅B�K�oa����p/���a��*�koH �~܅�u�����v�&S3'��&��m� �]`��	xP����n�����^�"�'.��0oNw��B���ƕ&k��Y�+�d��^��*Y���~����c�> ���K<���cs����T�Ԃ��4��9�Sq����^��ffQN�;�������
�<*U��d�xx`�yM��ŗ�ɠ��� !%ϓ�:��  �A�B�ߍu'��@�.��{�F�����e�STـ�'f��t�fF#�-Q~���Z��'���-f��-mb���J+�sQ�v�7uT�5�4��5G�H���h�w4�b[��]�t�f�
Y:P���VW/Ȼ{�W�Q2` q��^�y��%�����A]�e(CbT(��V�F���Y��Wx8���'��q�j�u�/���>�.��ք W%��uOrJ*-��3l=u���0�E�j��m��9�Pk�����`c
��<�Q_��L@�"��y	��so�P�J#����N����Q��Qj]arUz�����Q��[1 B_�"�J
dIM��wo�SJVk��aR��^DȐ۳���]7�9��x"ٓ���5Y�!�j��C3�N0X4^�p��ia,(K���]����6�y-�^�D���`���u�P!�%j��otnԞ�&�>�D����4qY�7��p;n���S��ӉMG�L/ިc�1!�TҨ�}]�@��� ��<��1�OE����J�m�+�tq
�f^\�0���e�L3�`�<��6���H�[���ݵlVP�v�|Y<�|�l�R�b4�jq�� ��
	�<m���u
v��;�P�3y�U��k9�j#�rں��r"X����Ȣ���@���G���w�&6.��s�ae��U��-k'���!Ϋ8��0T؅�Cpk��X��/�O�&�v�龨�O>ӧ�|8P.rn�b+�ε���~esc{^0Ů�Z�3+j�LZ�}��oyX�J�������\��)Oe�y�V-f�A!H%̬�]��.�6�@t@~���V�k�^,��[Z���8�5��{U9���ѳU6q-1s0Ԋ!{ :��c�֨Y�X:8�2?���f{
M�j�>�dZ4��Ja�Z�q-nk���5rDVR�w�%G�b�
h-�f[���U������T�ԩ��pC�B������[ꉑ�~��Z1WM���:��0��ע�����n+Wd�[�v�FL�ȋ��?gN����S��B�]���!��8�fbo�3��B�SJ7��H�<yx��8'�8����]���3C�9c(���2i 쒊��`�����Al� ;�9dI�&���)z�YC�?3�k�%�Jܩ�$��2�a�ȿXZ\�Y;Q�q`�%#�s�-!Q҉�UL�2��`�����n�3=�E����6N5������5���&� ��cC����� �m�W�5ը���{��X��%���v��j�,�Ehn��G��D�;[���3߽�B{�c����(�d���1	=��X㐖W��s�����PJD���J$5a!'rt�#ړ��9$-C`�U�t�_�[`SmF��|6g4�'g��y-�����$~}�`e�{�ێ��5�?A�Q�^-���s�dt�������܂\-������״N]��B���R/�����+U!|�˾x�|��
�R�ʇ���PN����9�[4���B7�_!��aP��]J�y( 9�]���%�E���Jh�D\����`X$(�Ȃ�3��rD�!m��gh�TL�h�f ݑ�x���L�z��Q���v���v�VѼ��rY&�
"^�%b[����SO(T���wnb�󩺭(�� �-��j�=�P�>����G�"��$���/$����'
��<wo�h#!	̖��&�4��Zl�pԕjP?H��y��v�y��a����E�xڲS34��[�����ٵq�H0�#��k`�j�3lg82~.�ǈ�8����Iz��;��>�;㧺�Q�?R���L�$�zK�p)q%��rZ~�mO���}�v�@���o�w���}�!1��L�Fl�/��m�3���ؤ�۷�s�k��LMi>�S�LoQiI4��Ǎb�$M�/�S���B��������6BKt���p��5K��h�Ol�"J�3'�g[H�f��C�4���放	�p8�X�0������^�X�/�w׬�(��\��Ư]�Nl.�h�R�S�%C��~�V�Y*�9���ϭ�'%%x�B���V�@��o���)n	A�`���Y�S��@8IQAx������ą7e �b�� -&קK��������b�(Vo�FRJ{	��H�:�`�Q"��S�s�W�U`����0�9�_Z��8k�͉��]~��7��_9��jI�$Bt�/u�K*��ֽ�ǵI���'�� �B����������\N�+����wb~���g��+��ݱ+�����
��eWm2u�|����ltJ��>������f�m��W��|�꼇���,��CJ�|Ca���I�� �a���Jw>�'A�qP5�9D�߰#C`�(Ww����#A4,��Y[ՙ��a<;:G�ѱ��43`���z�vj�����fV�4,r��œ�۬{+q:��+3`t+ʑ~���=�;�n9 �=pt�1�F
Q*|�1��B^ڲQa�0�o�8+���>AZ���G�L�� �x�̯2��7S��qm���~E=[D�9Lϟ�C��*s�:l��Q1��3�����_uמWFV}�e�_��}�8�"*6�������p���)'˅����ȡ�rok=�m����}F"}��#N_~���c<��f�)ޱ'HA��ْ_�+����lҿ�E���P��Ǣ�~E�8����[ryl�1w���$�N��4-�칙�_i��fz������0C����Ɣe���2.h���2�-,H=�e���]\�fiU4S�s�X�Y�%���%#+a����O�&���aC��y�M:ӝ�&��}�u�e�Uj:���kTRt���w?7M��Cq�F���a����6E�}�&��}��I�/��Ƚ����S��ˤ����9eFquݷ����%��0���n���qp�I	*����w�B�ȑ�YՔ�pÈFS��3���L�pq�õ/�ŋ`��A=X�r�9�'�`'"���Gλ��Q? &w<�X:#qalT:����7Dܽ�f{�J�������;Cjd�Ľ�+�c�%��M���^���ur>���&΋R/��5lҕ�ʌ�J�=�f.>���[�3�~��zr���`���L���������b'�3F���dY!@�?�vd?�]�71|�pK��'����#~v061����oU=�;&����R��g�[�d��X7���,�9�����Ҥa)��I���pK�_ez=���sҌ�ps��5�9.����]W���<�q�6˅������w^,�QC+MI���� �"�L�(�"	b���T�-��h����K�<]/������ �8Te��Gl!3^����Zg�k٤��Z�Uٴ�b-�/��#L7"�������i���n��Sʳ��:obӨ�C�Ϊ=��y��>5dNs��T��Z_*�k�M�����Ǥ���#��ĔۜI���8�	�۰���
�0�S����]�*���Q#�Lf����oӓ�P��aw��j괽��,��s�J�aBH;���9��	K�N��2P��>�0�,;h��)�U�P�L�8���q ���p}L[R��E
�j.��J6���R�]<�xq$�P� 3���C���~:j[:��9�m/	泰"'�(�3���q��b��.JX�2��RWb02+&
���We���:�輤�7/�@TϠm7p����ٳ�A Y��[A��
`��1�4а���7��TW�������N�����F�p���4�b�!q�/>D�[]U�s �$�&*娉�spc��5�t��+�������Q��o�Z�?�7;$M�o~Ʃ��Z���.3��e�Mr����f`�4�|x����
����S��mv@m_���wW�䋖��EIRna|=k�9�;<D;��k݆S2�l��RPogf�sFu�~����Ճ�(ǳ�����d��S-[@O5�����7f�����wQ=�0��ej�c����(y�Ĥ��?��A<��S��YR��d���{�SB �f"+,p~֏w��G��U�:eF��e�)c@^3�=�g�f�����b$��E,_����3;��E(������ez��<)����*�yNa"���(������WC�<���T�{���!�0:7�<z)Ͼ�{gR��<.�F�2�-Wo�AoU%¤$�m�C��Y��c�l�>�v`�y��S�g��Ҧ�?]W�*z�pb%��T+�g��	�e󘄌���vd ����
,E�� 'ؽY,�I�nI
N�z��6���[&�O�&��ʎ"�[�T�����4���HQZ��R\�'댟8cpO�v�Î׷~s���@Szvde,dI�O���.�WRD�m����m)YHP
�\UjȥY�8�א���sm��q���>|o�yu\Q��r����I�"6iFyrl��!����Y���0J"������SdhF����5+�i(����)9KN�>�k��]��+�hRL1����,��8�4D�TX:y�O��)KL����x����"
��=^s�}�9��<�8M/D�Du�f�|��_�t���ʬ��*���L'ul�{39�UN&O�hum���H���r^���_���Ʈ�s�8�ù^ԋ~�p�����2���"	��*ۜ4