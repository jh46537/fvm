��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<s��.�V5JK,���z���$S��r�OT4��:�Ї%F��o2����6+A\Ag;�{9d�\�H��YQ��l�
�q��q�������	
�ߚ��!f�z�_�8�!.8羿#@ /R˅��C�΢�� l�
"c��ś���-���D7@��]�����'%�@��H�X�;�gsR���o�0���Jf��q�pN%os�^��;ˀ�m�8�_yh}�b0��1���L��zvv�O�d��멫^أ����;�λk�L��8}�E��V=죏�V��(�%���AV����Z��uI1�������E֓��E`mO^�<L��� P���e셿�*:�o���<iF2A 4��6�=����i�M�M�=�Զ!��/����<��\��l����L��b�zd�����կ,K��}nH��j���O�� �xR��c W��XA��0~�5����,�����m����!m�No��R�	��u�E� ݩ%��],t�R��T�f���+�:UXV�,D9�ֲꏢf��Vؼ������� ��Uk�PT&K��9*�	!�5&
=���}nH��y��Jz�
��2\'@fU�?t�� ^�u���C��Rᇐ����!Ȍ?��L��}[��~PK2��7॥)ELEf[B�g��bea�U��4�2���t�+	t��Қ�L�L2Aޒ�#�� ����l\���:!*����r�pR	(��
Y�F����Y�Θ6�R|Z���VL�d3�}�̭z��8KR���nE�OIP�<�y2��tL�[�rr0U�cY�'ڤ&���$�KJ��RӺ��;��vxf4���5%�FR3�S*�f�k�6�;�d�%g(!`WUB&��k���>�N��*��1"d��W[�i��V��YM�+�7 �`UY@��!P܇|�V�:�u��BU����Ю��3lS6�����T	�mcgW�.��X��i�����!��_���n�2����V��%f%�i��f�ZN�Ă�bU�y���&�b����&I|�@���ۛf�(?F��F}�!׬Hu���?���*'�Iʢ�<>�������i)1��Л�sn��+�O�Ǩ��$;Ʃ7v�6���;a�
���lZ�A��wa�WY�!��I�������_��-r����߄:"r�I]ޯ6����%�)����y�P�Q��?B�=�����4#l#���/ԾD�����|g\�P?���t�)���W`~~�~b�e�5���P9�Y��`�C����c9��GJ��z$�����  �����0�-}Y	ի�SӤ��/��k:\��� Gj,�:1�~O"YQ�m@&?�S���A4��-2�xa��0�*��*2
�[����b�&dO����E�GU͚2��ːyx�T� ͤ��i}��֖Ӡ�sT!�"���^�~�I� s��,L=��\.|0�o9�d�kN�5K�;��'_���sn�����k=�����"���W�*$�z��@�\���UvК�^)-a/��1ҷ�Az=����X�Z�-v8�p�"?�y�vp���k=��9"/P"U�Mg�Ks@u������ A�W������R�ЩHK��s��<�����u��,��KE$Kd*�-��=3G��iݨ�mʹ��["��,���iv3�����ףA s`p�m�F��{���΢禆Y�'rP�_�td�
�m��y݇�����%�2xV.^�(�S^�o	6	���x�DY���1�*��]:���a
?�Ȧ;j�]�!9h���1���@�R�����X���Gc�^x���}�(Yb�Po�����a��Y'�)E<6��K�HӉ#����<�d�6��(_�ĭ@�|��nd,�p�@,D4���[��
�2B��@ݏXQ�#�1V�%�+�������7e�5�HXDJQTv9����(�OD�w�ӎa���]�I�Cv�p�h��3`f����YxM-_dd՝�F��|ê�8k<�{�ݞ"��8eTD�����]�ώ̺k:}��_u��7+��l�	���,�)*���M��Z�<���
%iލWε��9����*�QT���ei�������$����d���8˺k�Fwï�r󭭮s��}wK�Äx.J�P�_��6�(���`�.��T�.!������|u����*/Ȯ�2�'U��m�p���o#�f�̦e�U�Ih�<1�v��}p�N��qCP&A���(�[47}��w�A7y�{���{�^mb�cj� ����:��GL�i:�J!�rx�Hh����:8:upY+X���3rYw���I��H

��$�Z��؍�/�r�25ٲzˊ8΢o˩�@�Y��Q���}ӣ�2�b�Ơ�g�[#�GK;s8�Uw�z��6Bc�����!>։����V�%J��Ȕ����<�D^��pW�ҽgbS��z ͹��;Z���I������
�}q@��*�:�C��?>C�f�l��<�=Ìf�����M���k�p����b3>M�׿;q䚟��E������_�g�t;�*���6o3�Zd^>��'�)p�8O"���!�(�?Z�%���n`cRu_pC�H�F����K	���m�g�t��>^@��l�9���wp�r�-���}�5���8͢PT����� ��A�Km>��A�{}Z�%�=N���;A��'X���A'�L�S���R�NX|8ND��Ā��@5�k�cE������ ��;/Vf�����:H����.L���ډ��S������M3:��@J*SZ���=�P��&���>��H���}X�ռF������V���?����|ZX��+�Q�|V �[I�|�{44.�E���o�7brݲ�&S�����l�����Fz�C���\_2��uE,���!�#`��&	C�Sk^U��u�Y��ls�}d��^<���07����F: t�G&X'-��*��t@.ѲE���SB(jY~����a��m�]tg�g�/](�'bi'��$��∇�JH�h�R�����n�^�|�(*��t��E&�����;V��XdrȎ�d����Yo�E�p7Ԡ�-�3�#!�&	� �Yn���8�"T�J� GR5�\Ѳ�/�FsK)�;,������Kx�J�V:�j�����*�CQ�t�+�"`�4�_��WAح�G[R�Ժ�o;��%�a%�t0R!$����r�Z�6�C���W���9��o���)�_�.YO��B,�e�Ts��J�r��j�gf����c�4�\v�ՆY��R���3�I��댞�(h�(�U�Q�J�Z��b�V�PyQ#���PP�� 7a]׶#A���?�R~Qa�y�û�qK}#��Ut?�i�����W����-kv��(J�𽦯\�S`Ng{Ct�F�7��6�XAn($������'m�z@�3t1�'�U�B�ǒ������&x ��[���F�S�s��C�*J���b�]��$�%�f��]�˘�e���V�a�;�Z۴rў�M�ě��H�$ߴ�%�k�.�O�q��-��PR�-9	g'�2��<�A����iN�1�o�hW���&`�]֓���p(�O��^�Fl�����YpQ�r�xVm���.�|P.\�*T��.��/�i���b�\��]���R��8���0�\��D�$��6 cZq�
���|=�m��s�=�O#M} �G�D��P�h3?�j'��x��8�sjI�Z��u��v�Mj�LAT��N"�N��ά�M:8\�gpŌ+h�9e׹bEFO�3�3n��6�'~��x��vV�i���������P�`��Ӂ�|���藘����I�I9_��x[�BR�Sc�m��t�H%d�}v��)�[�����WЎy��yo5~�IG/��|ڍ/��&O��7�����c��Eٿ��8$��{�����XHp��S����z�x�}�j���z���x_B]�(ీ+��r�js��R)�o�mxq{�p.ߙ$p{�ɕ@�3a�^`o�zk�5�'�Փ���p�H,��
�L��ӸI�5��h�1��I���X\�j`����*�Xݥ� �/:G�>�~��]X}�7{5���kV �۹8��+��QL`�΃���b���D7�dk(�X��	�t`�}���v����iޫw���auY҉�@���x��s�G2���3|I��R�ܞw∴���'t�s�XČ��e�vcV��h����NQ����+�M�*P�4��mIU��(�Z�x��v��"3�25{��k�\+I�X=[�&�������C�r�I�voe�m�i!I�A�"AK��>IzQ�c�/|���ъ2�1�$�yJ��g��iD�54���l6T�<�q�Np��qt��&K��(��ܖͱL��*$;����>�,��X2�EH�ޏ]�&�s�$�́�
]��g{���U��_��:�� ��*���= "�_����5�UX���؄q��m��i\�jU�?���3��/��~p[򙛩ҫ=lV-�g�~�	`�[ϲ5���9��J�5?�-2���S��p���vf�C6L���n6�����y	a8J�R�.�b����v�m3J�1/���^R�2)��L+p�
0h2(�����J1<�U=H��l���Paz���/�;�! �J�����'�ǂ�
}��J�N|������ �M���觻�`��b.�*{�ҲK��SS���f~�|��Ε���Wּf��W�sk�h�!��)�C�)�*��`lo.�\���U��'�z�D9�z�����2}��U9�S��x���U��#L�W�D�roҫ����!{��H��"��