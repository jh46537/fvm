��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,V):��5�P���!�gPQ��B#�.&�I����͂)K-�-M�5�<���i�ô~dS��l�U��6��ʮg���w�!;X�r���u�DÐ�N�x�@��^T�(Aj��Y�9K�s��I�v�b"��c�k&/U����t$������!�h�<l�8$���k�Lc2M���9��γw�� ��-D�dPoѡPˆ��_������o{��l�a�~���W[�s���[E��:���]��e��J/��֛��Eki�C;���$�T��0lT��N=�V����7R��P�u�ӥ��
@��u�L���}�f�3�\ vΗL�D+��bU��ʉ�4j�`�ia���s��i�:q_x�ң2\���_�z�
��te��A�Fqȶ.%*�(�S��hW�#���L2"Zů!0�U����K�J��������(�r�������c�M���� \ߐ@A�E�Q#=�]\[��7wE���f�W'����;����~��Q��kM���L�p#$��>����T��|=��fag�w�M.u�mY�u��p�Qu!q�*�e�vB�QG��\�"c:��zﻰF|�L�_aY#Bʰ����U���f�SN��ر�
�y���Z]U9x�M�/��Ը��`�3h1c��A��1ǋ��{��"v���/��C��2l����SY��La�I��P���BSR��ߌo~�]���N���o�L��Ka�`���r-RU��1=����"s�R�<�YR��Ԍ���65�}��`SW�t�˄��s�a�{�o��rtx,0R%u��&���z�C�������յ���L�5�!l�C(�N{������j$�\#���`���-|�5�I��mI�<WO�+	����M�NX�Ơ��ؤX�B�Q5m0%'�K���џ;m�����e�r���n�d��:�Y+e��<�<aUw�t^�>(�E�S�!�� y���ڞY��6��V��!]@��ɔ����@J�\�`:ׂjXR!gO���[�.�&:n��I�G�ω'�T�{=����=�"�a����2�`P��	O��F�
(�Cs�}>�r���B���{(�-y�$yldM r ��xqr�][�>qq�����$�_X럻Wp�k4�*p��S8�i����}��knXv�>3������ ��p����뫓^����)_V����>ߝx�Ϡz�n�)#s��_���C<�j?�����Ur:�!jq�A�&T.~��1^��_$L�/4��oك,�{�M;�����z�w����]���d