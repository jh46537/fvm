��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb0(����	zik�0��ܴ�/�O:u�9��Yn�Y2�w@�恲�ۿ��FV'g��k
�e]���"��(F�[�;��H��zL0�u��L�2,��sv�EN��i&}���Ks]��(�;���m�N�Q;]�[�'2�57��.S��U�_c���kz��lPjt�>���T���e�O�a���E���E}��|��kba�>�S�p��[�>k���Fv8�{����`-��g� ����	�k .�%����%�6޹�!_��<�X�V3N�o1������I�e�tU0+�dJk�lG�Mʦ}��}&Nя�������AO��R BTXJ}��]l����m��y}軡{�#t����ײ�𺪵G"�����K1:#�Z��	�@�Joj%N�>z�?�h�i�̊z�g����OW
�|��q��>X�>��`��ҧ��95n �IS�+����~ ��9M���ݭ��>���%	�֘��&oK����|��u j��9�{�4QW/�_�n�ʫ99�p�b����k�ߝ�p��S�r����V��]�����$(K�o��:�sZ>n�`R���vb�K���6����[qz="b��q�2�m-�1A��>�$(��̫�6�g2�(0�����!n��~�Vͬ�%.��7BFٮ��⧤�fZ��v�>�Q���T�ް,���h����Bἕ�R(�ok�&BU��� ��&V
�I�5q~Ms̟�SD����(zJ�b���^�C(�x=��^��vzP ����j��Ʀ� 䅜���� 3���o{O�?{iP//=���\�I���7��7�B�$
.ND�;����ޯ &�M$�h�OOG!Z�X����Qh�5��6exUS���P������߅{W�n݃s&٪�(D�g��ϺB&�қT�e��y�2sآ=Uʾ��3뫑�(�U� ���x�&��x��{1�N�2��\�)���B'��a��:X��n��pN�$0颤�/�Х��X�[�ʡ��u���A�E��TtZX�P���;�}�:}j�D-�4���Ie�)��w}R���b*N�
n�Sa�� ��[߱�[�SEC|s��̲��x�ltQ����)�N#��>>%�*�����N���f��݁!��t�"�<ݚ��M�
S�� ��T3<�U"@QN�[����6Np�ҋH++e�g���b&Q� ����Ԅ��p���So`�U:�a4�/���:E�}�f������si"��Sז�ǚ��5�5=����!eF{�hgn��`݆I��`� �?۲��2 �:-�%�"��q.rs�����N��JpO���	�Dj�VU#�es��+f>�I���73Tg:Vq���􋟫� Y�82I�N�7�����iOu��qjϦ�����m5{&����l��h���%ȇ��J��<�!gb��(�s�c�e�!�*�7,E��f�"���i�|�uq
�8��ɒ<�W�f6��b�K�� ��(	K6#C�����e!$C�&1%�-!�(����D��6�',�=�+h�-�˂*A��-�*�(U�3&m5��|�1�����W���ۧ���N�c,Q6�'�׳Qk����D��k�(l�p&��&Դ,���Sc�@q�fW�<K�e-�w�Ht��S^���m\撏�4&��2)��@ur�����)(]E� 腾5��9C��d0`��>�l�M�u��R[d�Y���d ���:l�(�џ~Y��fו��K5��`z!U��#bSP�͌�ר��V�1�� nU鿊���aS��ڠ�ҕ�O�<��<J�Շ{s���<:�Ǳ������P�.12�Gԕ ����q�U�� �f�I A_�&�a�uj�E�3I�gc��g.Im���:�zKh�n�ؘ�`�/��v�}n$��ͮn��*��)m��%0°�Ձ��t;C����`=o�/:�"��F��[���|Ao��Q�Ќ��A�!�Ui�#M�N�ڌfq�=i�_t���V�f�-�_b�'3�氿�����~�j+��X�����	nx�k�hi��\�~�̽�!7@O1
�cĞߛ�}�c�b�&�|���*cy"Ԁ������z�>�
Q44��{ǳ�oi�b��fGl2n�%>3<��xB�wܸ(�S���D�w8�t�+C��!�>�gj0�ju#~�D�eFi9�R���������/�r��DH2 �Mzh�i�o�DmBXT�����Z$qZw�ωx!��VyBO��~��;7����T�\����`S|(n�ͦ�{ Nx���54K���Q`�������&У����4o�6�XG��CE�����ặ��f��4E�f�����X��$��
6��v�
�i7��2�co�:�C��'Z	���l�ȴ3���;)~��\���w̳���ZJ�vA�k����7���>�tu���İt�M��\]���!l��T@�z�U�z�܈��35�ri4�Z�����+�=�k����ZeX
暳+�10�  g����K`aj�F~5��5��S�����7K�y��<oM�����f��F�䄕��q8�F��>r�M�Z;�z�I,�C�QJ��HL��i�ߟ���ݩLVBd��Y�o�05?����=�u�jH$;���J߀�G\γ��\D���s�w��c���eU ��!�Fݣ�	��Ҷuj��(���b_ª��j�L�H��E4�n����yI�`g�vjX�^p�f��6#��4پ��ƶ�� Lh�>��y9�Wb�I�U����	 (�?>�����WiY%@��E�0&�M~��{�>b#��^(q�Y��4p�"���z��ň��)�@V���bҘ�R HԶ��SUm� ���^D+�(��g�p#߼�����&�Aƞ
��`���O��4���)aEJ��*1�3(��$5�%��[Ƈ7����y �eF�ڸ\S5z8�����[�s���jO3�ji$Ä��_?�y>�#.���`��Bm�j�e:�I�뫲"�Q@aK�
��d�ʱY���72W�b儔}�xbǞ�����gP��6��`���E���ip���o[�z�E���p�!գ��on�F6��w�y�&��k'Q�Za��1v��
��%����v��F�/}���˧��t�~��![wG���H�/DQ�����pX��w*]+	�b �{�'<{�F��9�H�k���c�	�9�yC@^�8h`l�yn�Ps���{]���� ��R�U��� �2=�Ң]4��,� ���X{�b��^��@xP-5b�7�_�w@gU`A���4&��\����Ç��m|��\�z�������is��S�B66f�M�Ώ�I�3BA<$���j&#��1P���`�/�}!�bו�Y�z�y��3Du7I���V��}�\�i1� 9�d]h�`M�W�\�.�z*Q�	%ݽ B��hni��j�nA��%Lcۚ����/j�~�4����Q��T����e!��n�y�8��B�#=��.^�rT)
�sͮ�0i�u��txy.[tB~��K��`+d��0���k�U��ȑ=d��~�IJ5ЈIe.l�%���ى��
z���\i�-o�|�'_��7��Ӭ�m��9��B���
���9�z��f�g�jK��K[MH��ͱ6�i�)~�E�S�-�G}
Def�V 7\^���o�������5�Ӽ��p�%]����]p(ŗ�����3+r��䈪7��@c֭(��<�Nm%���z�3f��}���"�U��3����{-��׾�<s�n[7�ueP�t鐋��LC1'�*�->X}������D+y��^o��	"�]
MI��XT���JԸ���s��*k�:����m��:s'v��WP��T�h�Df���[�^7a�@c�v�U=t�bT�r���T���w��B� �����Y��lKg�,���P�qM;�:��l�!��>s�8)��-�	Ƴ߈AQ�բ��R��(�?�Բ�n��W����yR/��_�yIx��A�T�ey�ݾ����c� e8�]�؅[| 4�d@&	����lEbz�ֈb���q�ti���xe]�%�:R~9�lU�C}��pje�M���D�ˑ�@SB�i�^��Z04���n�,Ot��$jS�_�b�L0�	B� �+	�}�c��y,� [�K��?c|+�6{�9���y_l�"$R,�Ȅ�����%�X��r����tCVe��(��#utX(�*]}�!���M$$�~EtH� �= �����(�=<ւ������G��E��,��oR6k�ߑF�f-�p���P2*p�r��t��"�"�6N/��.�ۀ��@���L���&(��wztlV�J3GG�V I�E����:���� ejx���NZM��9/�����{"@�'�ݡ2���Y���'"�e���۟޼�
������龘�yrl����~�EN�3[<&���A��ICL>�@BxW#�	K<�����F|a%��<�5&��Nt�L��5@��gp
c;�aW�ֳ`��\�_ת��i� Q��d��C�B�-۵�������>
a����˫�P�X��ubG/w�%4�R�S!�v�(�X����m�Հ���!��ZZ�;��u���]G��(rS�
9ӟ����i��Űg��%��h�K�b�3�Mk���4GĨ�ī���+vt�汑b�Sa������T2��jx��L$swL�ey�Y��e��Ot"����aNEu@��Z�:7m�cw3�+�zd VH#�B�	���a��s�˗�Ʊ�\��Wd���iѕ�ܕ������.�N��beTB\T)�t_�{���i��w�|9r�F�˛��&eOA:����Jj�j-h�t�=藥�� [���F73�C;>o�I��ݴ����?�v6�a�c�9Կ��t�D4��(5y����	I=k�q�هHCw�Z8gÅ1�j�G�H������v���E��H�(�Q%�����.��D��P*7 �� �'hDͨ2<������S��z�y'<���xh�����NO�Mkid���p�< O2��o}�br�=?2�:c6�<�������IiPfJ[iqjo���&��@t䚁���,a���j�AJ��{�)%����ԁX�x�?I�7�h�4�3����c{�(��1�h@�����Rܐ[�"�[׍�kRۀ��U�)����>!�~[|<�U?}�3��'4`GB���
�S��V���5KI��k�-n��<@�Ǎd�1��_��,��)�H��{�j��Z6 �O��.���*��!�l�{�oC��y��(wN+������%[|N#�tc�o6m/&��#3�*3t}$[cB��:o;�%Pf�a!���R�0r��@��?v{�7��������)�u��_��o����=z������V�Q!5E�"���%����2�"�ϥ�$h��H���ޟwr?5�9r�_<A�̅e�m�e�����̩��|�3�4Q�kSI�83x�W��� x��S���̪�W2֮.㎸�0hG�������Ӈ�p���@b(n�, �w����z��f�=�wu����v����4�z�ߠRy��̳�B��ךE;8/5�-)�����Kƍeb��.]��� ���Tٔu�!~�Z͞�W�Є��4�d�!��}~�It��L.>P���s*d��[ɧ���;I�6 v��(O�rRԐR� orj�Ҵ��2��@8e$��t�^G�h�i�b_�z�?>�~U���*-�J1���y���ʄc�.9��P}k�晴2f�^�iOB�l%T�z�D	�Q���֮��U%��Z�d�n���T��f�\��,c�_�du�_!9�P\Df)_z�?��@��J6t�L��/8O���Ket�^�8Vgy)&�j�8B��[���\>��zLNM����gji.R�����uT=�������:\�
�%A����@��%H�\�ĵ�u b^���«���q�'3'����nX� �v����I�WR�G����������>��톢��r9.S� �䟠��=t3��YiA��du��#:��X�h�����0B��cxDe�7���Ѓ���V�w��w��	t*��*�!i;^�<�oR��D�O������A��CY��?�����-�qkq��a�FÐf��1˰K�_f���=�G��4���I�j�S*.�KE���BP�bƩ$��{�33��V����m��X��V�v܅�f(lۇ����"�Jn�Q�Fo�?����s�}��yY�b�m$�9BU� ������� ���c�P��vr.�N)1.;��am����{����bJ
�Y7C�H�o1�6��/ N}$�#و��֡�T^�V��+'�� ��GM��v�.�R;@��X||PO�v��-	豒ߪ�r�,��Hc5�2&�I�\˃��WᏀ�Z�˵~��%��5��'v.����;��S��i~<F���ե���[_T��~1G8	_�z�n��	v����-�'V�ɡx�v�����3U�i�f���'ɣ�=~o4��e0���b�t����ڕ��>��^�ŏz7�ǽ�<���kv�H�A/���	4�M��B^�	M�;�!\slpH
�@,��Ղ�{A��y�b�Tn^�K?����*�X�L�m�T]�͑C�|=�?��FW��s�5W{�p�i$[-��\��� <��=i��Q�&f���x'Ekx�r�il9�4���m"P�y@��U7{t"L�^��Q��)��t���3%���Y�ɪ�M�)��eF�_�C<ex��#���	 .��E�I�v�n>u)=�
�}��]̓�T^��w�AX�F�X��$�D>�yY�8�'��y-�\#F���=Xղ�{["��i�d	�(�L#�8U@G�wF?��`�������*`6;���1��-�,��U�μ��w�-r���������*��F41ԑ���@��#~�6 Џ�D�����e���qʔ�<��h}�*���]�j��Vrv����p`�%�Ԗ��i�L�W��g*Q|�t�џ#�O����=K��ʾ�US�n���LT�]r �)>��(6a-���iw;l<SL�&��n��cf�O9�XU=����hiz�J�M��^U��\�d��+���(���Dȣ㦅�x�#�	�)�Dd�M����/����)J��������h�����UZԛ���@t?l�t�<y]'���8M�U͍��4�����Wގ�ж8971���7&c��rwyD��aW	�Mk�(�Z_�������a�ST�^��5G�q�~��$t;wc�,�Ԑq2JC?y0�Yԣذ"I)�ك���|�2����G�z�o`�߽�8��MAU��e���/Nb��%C��P�vK8�Z�zY�M���fA�q�%��f'��������摎���ד����4�G6/-���3��a�$�~j8W��˶R"J9*���*�9�#�Is���%-�b`����T�!2p!�ư���}m4)����:4A&�Pf��������n�dX�b��\Oy�]caK��_���w׳qy��B�v���vY��՝��<E��,�G1z����:�3�u%ͫ���1Z�A�aQ�y�d��	�T_�m&�ۯ��=�L*��G�=�����L�����_���@}��<�J%���7L��p��T�R	r�ݬ���D�K��-!�[����