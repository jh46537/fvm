��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�ֶ�3�4q����}��{x~�� s{��TFҫ��J�^���n�AH��k���s��#_�;�b�O�u�|�������֨��#�:�b�\77���}T�I���kX�ի@�6���12()�|{J�4�&"�}M3���_���mD�ی�`[�K1=%"�T�3����j�;&���%l�`��:��zAjG�����.{��X%Q�Ͳ|)�K=N|�lw���XP�4�@]��D�����2b��"u��eg���J�u�%�4�^��2V|�]j^���
,�9�O�1�`.�2B��9��5?r��7����։rmf��퍱��CP�m]��}���&Cw9Z]����u0J UO��t�i����i�O۱/g��@iJ���2[�LC�(�$sZƌ i�jw�ҡ���[�c�"�Qjw�cK�َ.�$�]ɒ�\N{?��/|��X��_��(���-*r�{�{��R��PB����m��Q�i�W�q�~�.){���/�^<�� MgZ����f��� { <��6�I��}�pc>�=F�1�jG���-�R�Xԯ���fS�6�1޶V@$��Z���M;��M�`�0�d��u��#9U8�reX����N����6��DF��A��|3�Ӵ/ˆ8���ZP�u�Ħ��ܣ=�&����G�(����<���nP�a
�ƴ
��|W@�Ыw0J}�s�W�3a�{�,�O���9JfD�4�	���|�H��[N۔)������<�ֹ��N������F�Q��]N���J�}/<mX��ZS�؎Jŷ��x{�/��r��Z��<��PɄ�no��R��ɡ����\��`���J�D{�ٸ�������b&�����1@!c(�چ�e`�� �"H��/�N�[���Y)���ơ�z�*��"���QRT��
N�+e�fd�_�;��z[�C�$P|d���Kks���G˘��U�����R��-��\٥y]P�ݟ��^�;�&�`���� . |8Q�Eu�{)�aY߻��H)�۹���̶��f�ӍA��A�XfQ�fF\Y���ie>��m�������]���x�6��Q�8n�����}��2��c�&�ֹS�j�\�_-�*�<�e[mTq�@����X�>�7Ot:�,7i��ȑ+�Xk�>�4�z����cW#��2-p<Y2�a�2�zs|4]��K93TfYN�~���@�2a´�@RYq��^�e��ǁow��l�.�۸[^Ň+e�겓���}�w5ڪ��/y��f�PuO�U�߃F�.W	;c�7
*�½�9����]����>�M�q@OLb3�)DC��l@<E��hZ"�ql��4�N.FF_�k������X�Ә�H�\�L�1xje%)#�=޵΋�h�ΆO�`8X�8���Bw�����9im���[��� t���@�@J���p2
��2&��O�#�X��S�	��<G��2�V�����3&��@�Q��m�qc0�Yv�*���[ۘ��Q�~���)Hc�N����F`f  ��rs�>���E�	��_rH���Y�OV��h����Bݩ>���uJ�AV�B�ᔽo���0]�vcJ,��a+x��,I�u�4�\��̜f��V�����%�m#)'�*�L�@�:��DL=�TC^��?��}�)�Tm:�t��A�W�����gU���MG������'!����> �HEy1B�0!�2�Wu�.�;��K0a�e��9M�(&��Ų�P�͟��Q�ش��eD�V$9���cC�[���Y�� ńЛ�'9�A����eƍ��R�a�!;}�3\ ���f��Y Zo�	��q*��%0ʖ�n�+1����Z��ņ���`�OTp{qs���Qm����"gs�&?f��	-evygF�!�k��(5��4B�x(���3>�=6��-W����\w��`��U��ǃ@��@��=�ɡ��S��I>O��UB�)5�|��N["���?I�}v�!H��=i�g�7z/?_ޙ�O*�D��U�#�*�_g�$�&�m��>�=��4�,%K$Ɵ]ؕE���R��|��M�������@O@x2�e13GnF*�U��B��Q�K��+ͻ�����m����ۍx���a c^��l��5X�!lZ���?@�{�̣��0h�q4N1�l�?����7����=�E1�
f[��)J�|��7|+e�S$@�O�NO��h}��XRy��쎾7����fI\1�u�W��~-p8��/?��3�sֳ�.>��S���� �=M(��/��m��̈�V��#K�ш=;�p�%2x��GзJhE�I|�ʎa-F�"�^gBP��z�`u�ΥJ��M�Ԍf���l���}8���`9y(��ޮ�3�`���\�
��D����h����s�5x�6#���|X>������]+��}�:�m�%v�e7�eك���B�m,;H��@� �c#x¢�1��,T����ذ۝�I"I�'�3�k�m��t3�����1�dc�P� �h�.V�Q�nഺ�QVL'�>�Nx?P�"ONR���$�kcD��:Y	-��e�O2�l�W|ܞ2/D�5�U�\D��(�K��eH��]���;
(I�_f������UZ�Ѡ���{���Ə=}6)B٥�]�_�<u]��jL��$00�)'�_�����x��_�]>^��%�2.�`�,�@ly�1j���&C�1��Csǝ��J�/����}�v��@'FȜIG�{j� 1�op����>a�� Kxil�k��l/�X۬0(�	x$ی=�h��������1�/���;A6��ߙ��}q�A}o��>����O������o�O/8`2�,Nͤ*�r�|�1U����ã���c҂0��U)�5�5N[d�-��9�ɪq2뢯�ݣ��������E�'�rIQ=;�\��ft�h�nt
	@��}��Xd���3�2?7f��0�JG�88�G�׍ Y��,�7L��FpE+l�\���k��H�/^��V"i�$M����u�c��;�㵽�4���#���-��Z�\C�.������>{����Zpggܑ/�4��%S˦Uk�Î�:G�gόC���R��h���;E�� �9H�I������TB�#	���ދ��W�Z*���x��8�+�z]U�u�$�i���I���,$�L,���:0G�h�1��šي�Fz��L��P��(m��#�6�$x���,g̅���I��<IW�S��HfoDX��'�Ä	�]�r�$WX�$��:̇2����7����X��?`�y/�?m��r�0۲�N!����>���� ��?�b���7K'_dm��2��BF$��P,N����Ĺ��T�1F�Yey�p���6�ѪM�	w��HĜ��@�QsàP�͋���*��m�}��v�A����M�AD�f|�b��x�c ���N9�� 
��ߟ�R>�_��a���Ͻ���*t�>����&�wy/�����r��1�[p��\[;�99�_Eo�� \"x��u�I~�*W�NH��*� ���{��$���C�-N EC� ��d�a�1mַ���ϭn*̴m��=G �(a%{�G��b�Q��� A�X�nڬ�g�&ap�j$I�4[LS��J|�h���ѣ�`��il�sܭ}W@>$f"E8�quS""�0�0Z-�����W�� ]�AGd*]�"T�;֢�C	��`��2s#��{��GIe]}&�bk�9����#�
Z�xKn���m{5Ƈ��%��A\IQ�Z��p�� *�˕*��FL�����ף��ʬ�?���~{;󩶭���>���Q��ϔ���-;+�(�Se�kd�#�LV�X1�;O�vJZ�e��;�rp��r6�
��X�٫iJ�b?&��������f-��L���A�6MK�!��"�T�	\�6Fկ
�3Y���&K��X{�>M�E�h�.�1�⪉�`$��n�a��!�BU.��jD��{u'��R���*�֭<�0J. �ٷ?�k�n���3�g��Y����u?k�3ND���V�6�AqhY���0)V	�̍��S��OD�%�Hxܛ�Em� ��Q[�}���,#�^YGn�K��q�g��b��o�cZ�WZ�d��y�N�u6�wI�"��j\�5yq�ѳ`�(?e�vbU��ۈ��oǥ���c�u���wݏ�;�6\Mm�>L�p�"A�=���ұM;�i&�F�gn�\ؔ���2�r���a��	��|�?[�K��g��"q�q���mW0�&m�w�����%��\3[�.��L�}5�i�H4M��C���xҙk�^�B��A����:wݾ�����#����'���N�<��ڶ���R��:M�7&��NC��P|8ْ�r��r��T�����o�P\�I�.�)a��ysX[�SP!ζ^���֔�m��Ɍ�v{t���0�EfT?���N��-�����ė`�*]:3��_T9[�z�y�g�w�YmP���~����"t�#J,��*��\L���5L�����T�{;�"���>�&|g\�8-�p6�K���co��,Z�@���ifĭ7p�C��3u"�.��Fa��q�k�8�B��p����S��>�O[�l9��+�;���q����h�:���kUx�r��:��o-gmJ�{6|���	üs��#=3�����!t��0S=_Æ�هs	�����e`��VZa$Y(�����zX$V��Eq�Y��̒Vl5�5��:��U�gY����~Ef!a�gN@�<db����	$�%f����;��@���]�ԏ3@����V�L��3"gC=�,k�$���$2ŋ�����Z�q��Ȅ���~&����!�˦��ß,Ż~_\�e:J
����on�'���r�Cě�B�������Z 9�T�0}������A>�z��8T�Ж��aG�sj���z����P��Ԗ��Ԗ�{��6�mN�w=��\Q�IBÚ���_m��� EG���ckw�
��u^��y�^0�K8�=�5�c�l9G�Q���	%?���P�v�n�lD�f�#��u].�IO�Ȍ{�Ih6wsTK���6�JZDV竻�%�*��E��Qm-zn>p��>gIR���.�QB��B`n��]���
㔉C%���nF��JycY� \�V���~��/�u��"���כ7g=�{��$H)�(�3f_��IòB���:#c��"ə���Ͼ��(���������0��T`_�)���R(�Q�ƚ�ཀྵ�}� ���X�����{�m�mx��������7������(~~��D�ęb���M�;��B*'����]�
H�7f$
�F��\���F�8��[W���Li�`�c�
��u�O_�A�V�{�I�1������tY�Z�%ҝ���=�p��壻=Zp�A��v�	1��kR;mA�~`��p n�ߵ�^�r�Q�An�2!V_��cI	f*�pR��u���(.b]�5���Y�;&��v���:Qx|�8d����{P��̽P��M�Q��	r�b�TU�t��HV��ݸ�����u��hS
��6�\�,�w޽:0������6��W鞸ʄcpy/w?�.�4��p:�N9�F��~�aEe�r�©.����Ϧ`��F���p-��6%���f�#�!�����RZCL�/M��%
�,Q��q�2��$�Q�%w����Lg=�>��+O��|���*����c!�U���?�!��W4��n�_a������2+�1�ӫ2����|��K�-:zNVN�=��ɘ6�����[�@uN��Zn+�����{����!�
���C��*�e*�/�1k�����N�j�������;��_��얝�&�t��Ih��s��=��xΟ�����y<6�~ͳ�Ȅ>�HO����h��#��p��ў����O�7�^/�R��ZW��*��&��ۤ�]��~�$I���^�r^S ���X��.1\fq���M�d�C^ d�W{/��|���
N]\�ٝ�U���)��>Z�l
"����^fإ���;��6 M�UI�L�?�:nR�X;��~���7T��1�#S��Ѹ�Dޓ{fZY�����u�p�:��dov|+�r!Zۮ��§���^�n_Wa6�Wep���|�a��i6��i�p�w���NH�WM��iU�nB��N��i-!��Rz�H�&F(r���5)�J��n�>�6�"$�,�	#4&i�;E�)�Č�uk7�{i%�h`+l�}��� ��	���$����ر���C�$ص?���7���1����������N^NӍ0pp�ڬ�.y,�y�\&m�H�St�@���+"k뼅a� ��i�=�x(�J	���tXB�*_¼�E�u�;�p'/��A2�V��K�� �Da�]�2N5Ɖ?͎��c4��T�c�C���:�AW�DF^_I��SJ��������5J�Hq2I<�l�:��]����F��|��'��;';�^��� �y�+2gJ��O�����K�
����C���I�Q����k�%&O$k��2Y�1#W���V��.�1kQ=*̊���!�t�P�+ɎsB�0��!��O�p�����	n�{��ç��V�h���q�C�C�qD�|%q/Abm���>d�ea��\Ŭ���v+C��'��5Q�.�&�QU��S0xdON�$R�/#�>���5?(�Wi��t
��ڨ��"��t����j�Զ�݌�cfkAUJ�dK������^��u�>�7��+��ze9����iNC�ro�(I�L�c���<rb���G�����:��P�z�Q���[9�I2�K3
�rm���7�̄�Be�QB��퐻����2�n ߙ���PxsT�[���m"�d�l��T���˧����[���ߝ���-7�Z\Ҙ*9F$DY��@~nS�ӽ�s�I�y�**�lP$�qv"	\����c�,�����F��mV���E�Z�8�#�d��L@3�hU�q�[
�G�̜#���յ���O8�6 �a�Ddf>��Ջ��/u��gp]�	GH�L�~�^\[1�D����������KB������WPJT@���Imۍ�9�-���;+�Pc�<�@ڮ�)/�
�[��Z����4�λ�� �s�O�,VS$��>x�+��^�gA����B(��ϻ��-<Ypp���!Ng�*H�c���5uĆޥ�G�6w��wa7,�Յ�fUc�F�rq�Ҩ-��T�����jh��pt�jR�C{���Pl��+�Ж=�M�x<�\ ��W0�ٟ?�*���Q.�t��Y)VL��$��:M� إU�
��6�p#$ݥ*�5F��2����Ѽ\<�Q]%fI��L
�b��%��xO�6s�b.��,���n����cħ/V�r@|�B>_^B�z�j,���s�0$y�뜀er}����c�yg�wl�g��`|�7b��'���j}fX��Ώ~|~غ�����e���Q5�}/��O����c��!��j�&"l6������y$�ԚՁ��p�y���g�`5�c.�p~�a
�PXѴ��8A��@�a�r�/e��Ee;u4�*Ml�ˌh�
�+Z|;q�`8M��C�c�����jjJ�bn畦��һ��w@م�,'����|']\�E]�jƶ(.z��
�sYA�aIjӞ�wYk�����r�&y���	��i��7�����P.� ���J:~
��.�&/�EѦˌ�0�?��׼���*���Q�:;V|��o2�(Ϫ�a��׾��jr�/c����z��i]�9﹠�'FvG�v$���4l�|�>�;��v�ϰa��k0�k�Bt�����}|2[w��˟i��L_U\P��wb4 �n;I�'�C�J�z�Ң�\�w���VhW�s8�!�`�1��c-@W��{����3h����j���w}e�l��d̅C1O����X/��t �
�5�=�'73�%�%Z^Q{@�2m����9����WLM"��b��i>r��ڽu��f07F$�6-��Gh����{�AjG�W�[*�w|�h�f=k'{��jȉ�gR�
�0u8���.Ü*Lț��jGM�߀jo��DP��&���4ْ0��-n��Oz^s���	���9�P��Ƒ���-v"[���:��?*9Ϸ����E��C��zb~��۸c
�u�����<���d�"�\,�c�z[T��U�B��ǲ"��>a^�١��O�Z�}P��JR��4X�#��;B(�`�u��[��P̈Vԅ��р���J�f[���V�����W�������,�g��e
����c�z��k��G�°p���HӰ��l�șk\x�|��EרC�`��q��۵�)��r�a�Aꃋ�R<�����%)3�)o�C��`Q��\]P<,ZN����2Q�qB]&6Ǜ�w����Y���3z���a�
�����e#���?(iV�w7�<�5�;�<c�kH���2���֎ P-l8�Ԁ5F��AQ��; +�0Y��\ګg�C"��6�]h'X�MP���R�p'�6��nb�IQ��5�~Jr��EE_��(�:2}D�^����؟�MDd�'��?^������?+O ��;�ݏk������]U�º@՝���������"��9����߷]*��������+s���f�O��"ff�	�#X���D���������b���AB&�	��U�N�I:]���M���$�}�P�|*���B'�og2qx�!�+�xX㈽$v��J�NN ��7�;�� k�L�d;��Z^�m�Z�g8�ɃE���~�)ޤ�=j�#�^�]�7��wN��fv�)a.;�?G���֏��ХH�~yS����À�Mjg�A���N�E�Z�m���<�ԧf��j=��\�C���z����p�qQj�7u�J��2��[�?�?f})�B�gb7n��>v��kE�wږ{�6�z��8�����Qq�ܿD/��ܠ��i�Afj�.Y��mY���ŷ��2�a�++�K���w��=�8�|�[fV�X���͒z��b�B<�簔�a����b��5�p���YRX��K��ir7��Nm9.��&>M���/i��E?>�d2�\��d�n	�/��X"��ղn,����q?ڟ&��V~x�Ԍ� �p��A�X��Y��y6��ӊM�A��T߹9d���H����m���x�6J����[msb��Qm
�7p�
����_���F�4�J��/��+ˣ���{�ZIf�lHsEʖ��g��M��ܡ9.�}5=
��7�5ݓ	�>�m���$oZ*��'�Y�)���Υ�|a�&>#ʯr��O�����́�)ʄV��џd=��3sO��A��P���&�@�bG�K7������*ǔ��l���[�~����\�����!`�w��Z��	�m���ҁ�FHF��x$^���wΊ���4�)^M�Ѱ����OS��J=�t��a�8rJg��/���w�-�}{����kK���aϲf,��`�j�v���_��6����b��c���DgM�b6>��HC:6��s(ג^�B���Nq��3dF�����[$���}��/#Ǘ;�c�;�*O�Om�P�ke%��ħ��C�]A�9l�~�}3_�]V�C!�b]߉_�aT�����Ǔ�4��b�+VM�"-��vjVߺ�����'I�
���]�m� _-�^����]z�ۈ�s������x��4���?�&$ł&qȎ��*E��@g�G����T�'YQQ6b��&�V��� �-�����ȸ� ����ؽa��7�+\f��Q�j㋺H	��8Mi�۵�GZ�����>�.�Z�"��`O��I���Px��$�2流_"U��]w�2ϊ��<�ʻ/��� �+T��_��s�c��1#=�x0϶?��L� YG>ɢU|g�dA2虝��$�]6�8 wOiÝ���6�������n�N�!��sx��L4C.Z��h��������+��$ɎX��-��:wG��f�1W"9=�� -���՞L����-^0��<c��,�
���l����JU�4��`��q�����:�
	y}�j��3����ζ~7j������Yu��()�CnS�$�'�2j��g�/��(��@3iB0 5q$�ʱ٨��h�p��S06#����0G�}��;/G���7�G�,G2���v��z�3�y�}9�$f�e;_��7�a�|��C�� Ӝ(_�EP7��˞S:mN�N�>�

��t�Ca��Z�^Am��$��x��[b�g�!�����܈�E�|��a�&���=z��B
,�,���K4�3j��ZS�2�s�eA\[V���Yx��~��tO�z�+C���^���z� Rd�J���tc�>V^F`�r�hTF��8w���ک���$�"ߓ����h*�qmȶ4���T;��χf*��������CՆ��l��M����of��C����J��XL���H�R���au�2.
+��<S����F��*c�sQf¹=�%�L�)���̺�.�5&�!���?a�f���D�\�(�E6K��A�l
c�t�*44x��c��.*co�t����0�H�"�bƳX������"��rhy4{g�7�K���Ж��>��Z/�r���yS�-�0J!6چ�O����V�W��!@�V����Z3,߱�S�bυW^����(��@B�h9�w��b]�қ�z`zZd�����dv���H�:3��z���.�8�Q�5H�=�Q�ܹx���5Tw ���y�k9��V�yf#`2~�d�#Y���<�8�X���K{��I!b��/~s�(T��{��5�`��]��Ϧ+���#���q��kvw���)�Z<�����/>C)�@��G�����;>.���l�ѝ]�.&-s��0{W|.�=��dW ��6\���q�i%h^Z$)'����0�J� �c�LYf˻�F�Qr���(O%���yd��DH�Z`-�xJ!�v|ȴ7P.�ś�o啡&Z����G_��!��r�b�J	�uV]�B�x�����K�1�sc�+�2�B��z�~�
m�F��pl"?��h�Ϋ�;7�
{Bf�K�L$�<������m�i����W=c"��=:�\ 0�#0���D���:�֑�OYf��]�G��ʹ���)7*�,�yL�{�Fz�o��4�:�)�nK��
� I��*�n&ھ���)�#����@��&�&!�5[�n^�/�qڡ՜ʓ.1���������i?A1]�����eYe2ùFC�����"0�9yޱ����@�m��!n>5E���-�[�|H� �5W?6	W�M�}�9�~4~�,?]֍�eߐ2�;���3�i�fk�%m���\J�Ԕ򔑿(�R2�H { �����e��Ox���)Ws�������MY���g����W�1B�~4��>t����\�-����׳�[�Y0��:tyD�7�WY��cGZ$������.�s�c�:��?�z�	�kUd���l�_љf���=2pͶ�=NJY��jDW�j$�C����^�J�.��LP�þp��J�&��L���@ݩo)��F.N�N�\��{�c�S�\�J���8a��n�/���?t� ���H˨M�ƥ#���U��w#b����Y���f����V^Ġ��+����ډ2�\V��N	��\�	���܁��d*H�!s�-D�<�'Q�,ç�(�r�f�"���G�#�������b6��+��c3wG����td8.P�Ij�@r̙���W�qIE�V'�QdWl���c�}�Ѹ�`�i{�.}�ʣJ1&�?���F��7B$^�>^`����B��]��컓�-����6�S]#&��m��?[{K%O��?����4�u�]*��䭖�@��f���X:p�����(��>��yn�W|��Q���!�}z��1Z#�V5��!�w��f���f��]m���,M�n����x�f���\ �eY�&��$��0�B��ך��o�K"�|0b�{ki@�N�q�YĬ����?����0/g��Z|�GK�tƵ��!�{jc��s,��Y�q�^�ۼ��'�y�7C����4L	J��yu����11�,\SG��!�dBhsQ����z��Q����5��\�:&S�<yK̬�����d�R��a���c�(���H�`s-�{�?a����u�����n���)P����p�aL�1[�Ӌ+H&��c�I	|{
�o������t�m壹s�¨�m_�|E�B� ���T5�(=j�O�,c�U1WQ�8�F���!�<��|�QRI���.7_
'� o�_h���I���7	�h�ѧi��wfπ�e��'Eܚ�.3��L�� WR)g�Q�d�!pR5?N�W�΂P,��l�����y�G��rX��W|`��Sev�ˋ��t�PQLc-|����F���b.U�0J�l��ӱ����3s"ݭ�E'�H���(�Sy��(���m�f(/ ����A�g�`ӣC/%��]!�fO�����������O�Ι-��t�ӎ}g*N���h��s ����QB.�� �8u(�{�m7 q����t$+;�pH�0�Y�`�)ڝ���r��X�b:��u��P�Ed�˲�(�@�py���T�.�6Q����u*�AdNJ�C��]�֖YO��
��$4��N�-�+g�_~*�Ay޷����A��$Q*�YQ�D4Tznh$B-���|;��W����1�K-�BEF�h�h��N�Vu�.�dK.*Ǣ�<�cIa��Ά0"+���fL��ADR�gufAi8�^]Jj�*��o|��@�h��*��]2���={�I����C�Y��,��}5���3Y��V#o�lU�D/F~�?�C��CBR����"�0�pf��(��^�8`��-Ѷ����W����"O�<�6]8d�'l��NB�g4r<�q�|Yo�Rl��>�����F	�$@l��O���5<�Ϳza�,��U5����w��[bL�H�Z��(��J
�g��й����:�B���^���ŕ����8z��/���3��B�A0p�X=�vw
�>"�p7Z�8,X�oA�T�u��"�>>���.i���[� ςK��Q�;B����.��!$x�J����>���ݠ@	���5��x�!)I������0:�wOP�4m�Di>�_î���baG�T�%�a8�`:A��O�O�͊#N:�ī� 塶]�<{9#[lϪ"<���{j)O�h�p2b�yw�H�n!H}��y#b<�ڸDA+Q�GmD����r��p��t]@�e�ĐN/�| z�����M�`i '�k 8(�=脿#b_�|Y�M� (Y�Dފ}����g��芭S��L���M���$&�mz��M�]6$�Ӽ@�����$U��2�8�+�/���4�WlG� ���\ϗU*�V�U"��W�ґ����ڍQHt!�ݫ�\5�..����1X�O��N����P���y����f�<!�ΰ��U3Z���lʎq�p�L���(fGŌU������r����;�3��/s�nX����59��d���6
�ߑ�w�>���G�/VwV�=Q�y��g�z�hu���Gl�����:.�F���`f�)@�o���cװ������4��'�ޘ=J�Q�n���&���i���"�
ĵ̎Ͻ���:�
un!I�U�(φ������H�ȟ����im����f �] ����CZ�D[gTq�o�:6�����kŸsj���5���)���$�F��;����*�ݻC���C����
/�6;�H)U\)���b �BqWQ�&\���c&s�S���Fz�����2s��Ŕ��#����9�����*����J^\�[!�'�xt����g'�+�mA�f%	��\��N����7A�O
���y���`b'"�h�z������\�����H��-�pk��c�3�n t�
�_(�+W.���{���#%��)fd?<~p�t�(s���֩!*�U�ch�C�JFa­dz�����	�ws��dp����ȍ�"Y�~S�Z�m״�����r���Õ2�zb�k.&ۅ�c�q��SO}�S�g������Ʋ���^�S��=�-L
 ���O���w�hC���%"��D��F��hT�h�BW{�8�����φ�a8W j�*�^F����[g���嬗�Ů�c|[ �Еo`�C�[��)������Tm�zu]��Td�v�X���*F*��@ɛ.M���x���~.� �Ϡ�����`w3��^lITCe�_ ��&v�Obx-W�W/�l"]�@��VH��R����>��$����ϊ�֢-W+j���T�XՁ���0�
�%l�1>��Yb��T�4	�A���M�^�z&��[�9�	�Jjऩ�0fق/E�ZqR!���M[�B��l��s3n�����_�U�L�m�7,R.�\x.0��x�u^�Έ������@y�"�ʏp;Yx[��_���ѯ��d�^\|2�	�Yy�L��zH����'�gzj��{�F�9�4S�dȹ�WчV����|����c���G<�ָ�%W�p*�89�q>��LVp"��`��S�<,*��i��R�X�J��l�_��x��`X�HF��&�$as�YvmT���zp���R��-^��d*?H~�;�_�S���Nf������o� =�Ѹ�
"<��p�d�q�G(����	y�؋<����τo[���S��z�t��R~\���g���3Ѥ�>Ϯv�ȶ���G�$Wg�����쬺nCJ�{oH�wr�w�7C�(H�mF0�=�۔���b�E0��!�4�ID)�7u& 2߲Z�Gj'�Uʂ`E@�X2Y�}곷$LR;�1jt����$�I|�Z�4�y٪��P�پ�a#�A���>ޙ[s8�a��n���-�]BXMU�p&�c��6�/mϖ����W�>-��Q1u���R�IWN��B�"2��V��j�l-4��s�{���5�6^�(%�V�y١Q?��Sl5�z���X���M�m��'���^ķ��4���
L��"?� �BɄ�j|�}ғ�4��~�{�.e�fNja��";:��D�C�c��7�JҋD�&�w\�B�h�6���[6(��[���!h��n�^�pu�d�*���G��˧��ԁ%{k݋��eM�ZXA�S�ؒ�%g<��Nً�e��}i��+X]F,�5��D�JJ$f�BT���G7[�*���g\$ԥ���,S�����^{�@�(��O���/1�5&����/7�<��ʏ@��6���nY�\
st�;�e���-��N)�f+b��1sTAĔ+���4��c��x�O͔�R�~��(�R�F'(2;4u�v�o�z� �#GzA�95�@3��I~LJ��6���Ec�������S�Es���w����'�Ň^�9�U`����� �N\ad܍:T�g�H�=һ��k�}a��3���*'rq�yd� �������N�X!�����@2^�C)��;�+i���q�~��?�A� 鰌K!v"jw=���"��!��u��;x`��6��h.�tk=�F�t7t�B�Ԑ�L��%��ʅ����5bKHr$�yhcC5��þ��u߆��orY/�i�x�ss�fJ\���8��:Q}�j톅�`0I#H$�b��ח�M�!���{]���1n�~�-XB�N�=W��ꝳ6s�2�h�P��o�������3���?4�t�������ş�/)��U>� ���(&�j�J���=��7��/�!��!�	��	�,�&8���+a�sGkb��0�	𪷷^���8th�v��z,	�g,���Ź���L��,�x�D0�7T0-���S�AX�NGM`ot`

��tx#�ı\cdĹ/6o�QO4�� ��Y�h
��zE<ŭqGRa��E����.�'�)ة����6���3CV��#��B�1�,������ln�{���*�iF��D|PM+'J�%"�KA�hMSl4���Y�ة�&u#���c��r��8��R���<_N�F�� ��q�l�ժ�!>�K���B�DK��N�Ti�^���:�yW�C��*�%���	~�^)�Ģ'�=����f�x�2���t�j:Vy�N'iT*i#3�+���i����F����|�m�G�nA�|��MЁ�=F�����8���7v<F�-� �\�β��(�����^�σ;L�P�)6DA�B$^�Z�1��y��~z-�����7���.ќ�D�?��(.�1#�sm�	��D4�+h!(x}���=q������Ki+�!���x}��.�Ə$�����1�ܣ���Ӻ-R��F�{)�Uݱ\����t����vG�g2�+�23��AK �X]� $ⴣ�hǌ�&s�&gԶ��J�F9���|�g
�xZ-�<� l=�}W����/��J<�cC��Ch�w��
�倗�c!;�!B���R��������Ħ���<��ؙ������2?���p��K�Ի pC7�.�GޚV��3[ ��g�/^h�<g�"0�h\�L�֗7d�Py��y��A7N>ey"U�:˝7҇EO��t�[2.��ӳ~f;w��?�AE��5 8�d�ߔ�2ۄ�w>�钳sGZ��2L�}ݻ��*��h�S`��q��ZQ��涇�]܃=带HWv�yyd�VUӲ"W7X�F_��w�q�+r+3�
E=3�r�v�mo��d��"�Us�2��LU0R-'�|�FdC���
QYl���u����8W��>a�������A�V��q�k;����u4���LHs���1�w�,���H;�]·��{�j͎�]�k��I�p����%���g5��p�D��(ݙ�%ܢs����Ō��הV��4���c)l��te���y���@���]6�4É/rK�Z�(Q����ASZ!�>�SB���>�@��w���r[Z!�=��y�乭�6#!����X�-s�7�&1_���'�?�1�|���l���j�C�q�x����,]�ڥ�A�F'��W��:�I�f��0��K]��e�7���O�[��}��T�{)ʩ
n`�,�g��PtQ���޵��n��]�ǔFm}-Q���o~�[̀�I@W�pN\7@l,�D���G��aXb�Z����� d�6S	3MeQ2�l�d6!��8�0�������B��~�_zo�Y�	TF���L�d�M�[v�٠�L���_L���b�j% 6J1J;��,0�k&�#9��S&��olMs��������j�Ega�� �;��mNO�]f�AP�_
Y4��ylIW�$�]˅�7�˶�y݁c�1�D�DL"�:@�a+fEDN�X;]��x��ؘG6<1�%�;R�;�*a:.9IxѸo�� ��c+����<8fѤ�x�i��q_�KC�F 9&�C�i�r��Z�J���(ig��'�A���n=C�ۥ 6�dy\l���$T�6GVF)�.^�M8VxK��ߞrM��RܥΌ�K�D���f���#~&`����u��AzEx2.�A��0��/�"�p\vM���v!� #$�z2��  %��&A�<��=����n��U�.qv�[~���b��:I�<��oy������ B�b�-�Qţ�׀�A�����FJ�p�ڍ�v��v;kE*jWFws��Ѐ�������e҆��6�NFW8K�H[��tM��0#'�ˠ��)o��K��f=�ס��a�w�xO W-�\�uZ�BwR[w�TA�4�aQٔ���+���X��.��tW���|�[�.��	,���	�Fw'���t�5�(Ӕ7�(���i�{���]�X0�(��@����_��`�P�76P|��.��	[~���/�t��M���������K�u�e��B��|�����'�v�b��e���NZ��9Q7ō�+lb�h/
�����F0o���{� ���
V��f�mn��U�K���y4�OH�ݬE���i�UEHvU�8ql�eb��~������(��Ǣ0Y���V�˭3��� 0ġ�)�(9�Χ7����o�:���0k<�ٲz�����C�����2b��?+ac�Mv<���:�V>�gom��(��!��9��P�ћ���EU� M�0+���N�I��8�G> #��ѣ�W���Ѡ�p�5�p��lƈ�� �j�/�m��0��}]c�4�M��QF6�TW�W�:.�ұN�ݕ%|"G~�8�Oc��=|�Ri�+�!�L�bG-.� ��x��e6��oϪ��5M��D��i�޳��hܰ��}�AE��<Ed��u�D&�K\ڡ�n
r����?���v���F$�cy8�9��yD����?g+|��.&�xzJW}�	8��$���8�� U��$�v�Iu��Ҹ7q�@~w�m��wN�i,�xާJp��tW�K?�E�lM�>#�.8ofu�۝�)�u6&4�r��Ht��Z!٠��}�VO����8|6�yȝ����1� ?��d�c`ʲ�'�O�f��aG�0i�����U�{C/�?p�������L��a��ٲ~E\�aF���"�猤V�h[2DF�"�����J�$�Tcl:���W��w�ܽ�8�r�6 BHmxQp�S>�PF1�Z�ιw�m�Sv����k�{�?6$Q��խ���i(�*W���Gɨ)#��穈.g�DKŅ=�9��p�.��4#��E/��G�y��gs=�
�⸝LTIz���Ϣ$�c����4��r�4���h��.g;D��0?1"H
���wk.�`2Wa'󚚰�ky�ސP2?x4l�F������=�"Nw�Ԯ�hu�M�b�Z��KR7ze߲�22�p�\�Oa�y�{ƣ�����k����,a3�m�X�| ��`��*PF��ure�o#�,zQ ��=��/���䚎���qB0���\=�W"
�|x\G>��idq>���#sR�R�����eW{����8M�yw[�ݠѪ��1���:1��9��SNs��
o���FcV��%}R���EaO���a�
2 �)�������C;��y���}�+�n{J�W1Lf����Ak�
ӹ��3����5F�Z}u��c��ۻ-[�:3@�/�<�۴�u������-��A�o��(:D�Ȏ�D�������}~%�ҏ�b�)QΟK.���1mDI�"��Ț�r�f1M�q˳u2��>�<���B�7H7�AN�۬���\�SR��~a&�^G�>/ OYs{��Y��s#5d�yaꙓ�N�g�M8aoUƼ ���sR�s��qяo
g�"'�me/W"��3�JD�za���t;�JG`�iY�6R$�u�+�7a���9����
�
bt��_���"�s�Z��Փ�AŌ��ZHSH�1?�Mc{�ags5KE�Z���%��Lh���;;:�d<A��l��;E���{Sr$��gi̔	_v���W,�N��.�n���{$����Y)|�������:.Q��dU�g���.;��<���9����0��{���z�z��>Ʈ�V��
H����Τ�����W��K�f�`���#�u�fg��S���-}�eW:!���J߱��Cg�v��(��C���/�x�j9��d���:f5
UL'��@�}E��'��i�� ���X��PCau,�-�r�x���^E�X�����
�p/�9����K��������p�6l�.�4�Ʊ�=|!s�q���~_}�%����'~����3-��V�Y
����� �n�,J��`�X���|�m�6�	�>yd�w ��l��w����K�/I�a�⭇x̜'�"H4�狪3���t�c�S¬J)��{BI���k�p�6	}���q�/m�_nT�kVDi�δ,��g�C�h��>�<e�_�m�:�g쨪���	�>B&���?}��;����R
7U���}]�x��[p�p���ͅ 6<D�g�������Vn=��FɃ��L�����K���N!yJ$�-e.s�I��U����f�QW����c���D���68�O�h��p�R?��HT��j&��5?�(C��U�u�J`a�gw5|��F%�3���oF�tA�1���_����wc�y�[q�Lr��~� �ߺfy�r��|]��΅���v����gʓ�~������ց`�'��s��CQ�*A����`��Z:�<����񈲝��f��ʺt4�G�l�.�vɂW���SND>Qy�2��[[&�Y.�'A�e�:��ˊ,�q�u��k]#~��Q]g�2R-�� ����wD�ML�`.���1���3N�Y�i`ğEA�W�P܌}%ѡ���4� ��@Sv3��X����U�@�� ��yx�:�.�� ����\D�4��?��s�(��G�8���j�b�B����/n,g���½�����R�t��1)	؅��{ìhAmu�U�a4L��=U1Gh�dI�/����?�&�.�c���!��*��|f�Y�K��d��=��|���3����Q��4]��U��IJ�����%��?^�ӳ�����i8i3��Zj��)ӲS��)d����!���
��=����j��4�-����@���qG��O=�����Ժ9� ��z2��I["���FC��]�%��.aAYTp⊑��a��3I�B��ZK��ܨ�� O���u!tȍ��B΍"7N��$]��Qu��|iH�S�o��??�*�>��%I����4���$�wY���q��\_��
%`��]�_V7�y�Ϻf���a�`�ҝ)�8[�|���daP
��;��}u^Y,3l��ϐ��3G��cy��^%Mޝ�Ggт�U����h&L�5�0�����&
�"�q�R�ڒz�A���f��%�I�1o�|�b�34c@�>����ii�c�����3('�#sg_�jц�DkIaܢf�:�~�h��|�����SR}�o�*�/[ʱ�;�Oy=c�L9�̧�)a�ao��0@o������nXQqѭ̳L��%y��$A��3���n��}	}\",��;h��z�2Qd���h U�	�7�F�r�_I��{"ߟ��*����?�����VM*�\��B�dб�ș
����4��TPݱ�=����� �P��J	�O:��-is�~ �`��y��%��(��}9��k�f�Dm��b��3������1��K�6�r@�Γ�<��ތt��^^�9��G�ͮ���d��J7��>)?�?���U�GW�/���ʉb�,�~X�"�^<�>�Ն�x��@�еז��+U�#��n`�"���g!��ٓ�#�%�,RZ�]�e1�C@�`g�ry���0	��M$�~xF�݈��<sk��V��.��f�|�:�s�!st�t�& ����*��6���*�gC��g]:�};/�?����8���#x��,��(ti�o�J�x}�i�
S�D�a�H�OO�X׎u�"7-���̥��툟�5����&"b>�3�O�20��_S�~��Ti'�;G��lt+Y�Cg�r�ރ����U��o��u�e��Rֽ��Z�M�C�4	=�'�Rv�<9_�\�\z��a�rND��uUv�v>~3�����D�`�½tCxs�l�Z��lu'���g�75�1�)9$���"�G33y#��fs'�:�퉹Y��{���0��"#Hju�d�]�0o@j�7Y�E��KY�#H�^1��0��AKrAmH� \��_/��l���HY��y�St�c�?J�=��ֶ�W87l� K�[sr�>�`D~�UK��O��R�yrc����>���������T�֦巙=��/U!o4��Z�Po!0�����.�7?�r�SVᯌ��N(�^}v�����	��@\1Y4�>t�Hvd��;�^�����!?an��ݕ����%�#�5L�v�t�C�rv���`bӎN�V��b�������E����7��Q�N	�w��i�;77�L��ou����b@��k�����S�/	Ε6`��e>�̇Z��N����|�b*6��Pg�~'PN\:���������\��0̩�$�F8�}�60 F�����H�z.>E�	��NAK���G&:���M�z���� M��!yۚǍ�h\8~�E�1�T�T�ˣ�H/��d��`[^��Y?5�KL+���k� r����$f��E~G�3��lf�͑F����;y[�[��������(#�
�F��a!��Vy�G�x�xi�����y#+�M��MR�)}R$'�:�]]����k�����_���?"|�:5G%p������D��ZZ�^�<�k�2J��"�kM���K�|����~��/�6^�{0�-9�V�F�#���>�4aj�����DQ�74&�$84�b�Lm ��
mN��s?�s/0r��9����A)�"�fF��I�E1oO̵�}Oy���f�O��!v�����>h�����`(s`�1�RIq��IXn�Úƕ���r�AV�����mk��l�-/I� �<��c�R�xJ�z��@�P ���e*Pٷ'7�8Fd�sHV�W���.�4C�3�f��-T��z��g�����3���Qu��K�� �i�7ؐ�p�7{�f�� �ga���_/!�%�*�Ώ��zf��8] �z���`��(�;,tq��o��q]g��E�Z0e3��z�����i�v%�w�$���nR3���NG�g�?k�����+6~J6��V��e���nW��LX�(��>�#]<Ъ�����^�ll�V-�o�]�b��OW�}�V؍pu����8QgiRH�.;q�}A	��������fүQ�A�^.0s*�W��"�E�W;����\A [��F��*��=�H:�XsB_:vl����l6Y�~ز��h��2w6�,�0�v�*�]����꺼%��G.0І*��W͟u���"n�w�W���	@P��h�	#�oP*-R_����J��G�ŏ�N�9���ކ{�F����:h�;"�"%k��4z���C�s�f-БP�WaIs�F�m�����AOY�U$PƖ�@��E|E՚7�lUд���K��� �ip�gϚP�x3	� b�<q�Ҳ���騝%�b�(92�13�Gՠ~3|t�zrpVr
Օ�
�$��.!���z�Vd@�mFj׋�3�c���b<e�%g�! )!~��so�pW[���O��W��G��Q�Tp�"ۊU��o��y����DgB�w��y8~�y��Bx��Ndͤn�}���y�Q>&��6l����?pCcǉ��>