��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�×M��������`�X⯰�]<h��� U���o`7Ɋx�!�g���I{H���f�����&1�+)��ڷ����m�/��(�+u@��K
"��?A���yt�tn��@<n>e�q'J1B$\�xG$Pp��(�n�����k���6��[�ھ���K7>wCHYܨY2�d9����\&���~
��z�0�P�`F�����lȭ����>s�jO�aߐ-��>h�Y�x?�p����m�$��l�|�,��*0�J)��$�PC)͜7Wߦ�K�"��i��j/��
�[���IKT&�B��rN��,��<3�FI��;�
�B��Nj�tO.�һ����s\-����3v�l�����Qc�+Q1r�0eP�Z���O���J��c���4�#�bO۟��3�!t��-�j
�~A�̀��e����wo�fͤ��U��P����X*LL`ɝK��4ˌ�s8Ļ)M����W3�*1��lSU�Pj9Uz)�؃���c@�,�2����WDAro�/>R@S��|g��b	v+B�ff �c���~,��ۆ'�?�5���.�yk8�k�IYݢF�x3�vW����g��a\�f'{���跋3'3���ô�� 1	a��fL��&3*"i�x�N�Xӡb�r)]!���Y��T=XQ��s�KUE�h̓��I&��N@R~&����W��ت� �Ä��[W(���p��B~���k���.$YO�H�;�LZ+��l�"�7���G�=v9"�X�/g�j豏H�	,�/�!�p�����	���?�'I����ƅ\�r4K�dB�������Ūa3Dp*3��+�3�Xly!��;��� ��|#H	�}"�y��Y*
�M����&�-��q�Q�^�L���vN��) �] ���B��Eѕ(�<����R�����z���dJQ"���EX�y={�}s0G��n>��1��<���x�4�[^�����)q�#Nn�[�GB~GS���Eu��^�~��p#�`a�>Y�D�B�Ǩ�[����]0?w����~`��m��@?fn%�7�bk_��"�����:ы]��گ;&i���c,�q�l<F[�F��w8"��X���p�a'�!T?d	3�0�)�\UB�^�$�#<޻��*�n������ep��K��h������z
�_r	5T��!�x��nqr)b����6.}P��$'K@E�����;��1�T���C�����s��4��6�g x� ��3�+��}��J��c���O�>�z�I.�	d� �mx��og��p.P�I D�-� ��*�u"�����}�I�Z�ʷ�7��չF��[�� b�i�Ʒ`�V!/"�� ��![�i��2ѣ	ݫ����V���Y���j%Ĩ𲟹�A-�zo�	�����7uaS�4�^�M��,�e>�@z<����7��ߋ����\i�+��B�:�O>(�z�|��Y�7�K�P��ng�ݝ����-�eL~.	�f�g��O���Ҡ�#K
�[��K12t�;�ӹ?��x�/y-��($��S#�1D���dJsO��w�ي3fDĲ	�$r���[�N���|x�>���p["��!����c������ʐ�CW�k��m��I�
ܫ��@�S�����r��3t�E�t��������IF�$J�E��\M�خ�
�P�>@(��ni9�e� �>�V�
��Ãc��S�M����YӬ܄ɹI�T��S����&KH��ş��3��keC���-=^z��m�AB�qf��vp�ez�&熻�rj��Ux�b�#T��a�z���,�sԞb�9�c����BZ��@�u�7���<����#rBP(�<{)Y�#����Q �RN�a�gKpr/���'�G���a0�/D�i�@��%�H=y.��/�9��KPw��5�M7��T��j
���
�[Z,����e`,��s�����K�)Pԍ�rp�%�`�I�j��v��,���,I����4U��橴��7<)S�sG�.U�]貕���\�t=��D��^��{H�0�V�}͂ϮN!k�+]�0SPI�#6ێ�>p�DZտ��z��ׯb-e�c���$Tj������VVǱCu]��]^�8^'[۹<�B���	�,�9D7��
^46�O<�Ar�7>�'��߸�Q�}���jEB�'�99��α��DeJ;�K&?0�bP$^�|�7�*���UILM.pQ���x~����*`�t�����4�Glх�Ub���HҤ����!y�{����GZ�xЛ�8�^�+3IQ������<��������љ��z��Kԓ3j~g�%_g�L2�N��2ft��^�bpf|�N�`Uf�bbbF�ۺ�V/�0�)tm��#U. �hQ��W��c(�:�C�n	��n7�-����2�\�D��:tn�n��/�w�(>�Á�y��k`�N�7V��F�3a�Jx�ȋ����^)�`��t)E���<	x3[�ю��G��J0���}Q�mZ�̻�-�����}��y��C��Z?{*oNZ���v�dQ��?Ab�Y@V������3�R��rpHǸP�cn��gФ����}��?{�ˎ9hX��: �����Għ�p{kf��l�)��|��������E�$�z.�3�Kd�p���v�Y'y���_g2�]ɠl�_呫C�	��^��F�0Y2�{+��)
1Hj�/���.,� V�Kix<rj"�섣e,\j]ɣ^�ύNp��3��M�qG�E��ݐ���`G����߾��QS%�V~���F�?:�@	��C�(�������PJʶ��c�i�W���~�
@�_���RR�X�G30fy\�7�KRh�����:�zS���̦�j�	�4D���2'/g��:`6�}k��:�猵�}��ߨ���@)p\���-rř���*�'�r���˼&f J��7���*dG(�>O�^Ӎ��[�o�΍�${�i�&�'�*��$#�@�2W�a�i��leӢf�F���hl)	eK���4�T�*񋡱WW�h���֡����Ӕx�R��{����Y�S�Q ����r}
 �%�Dף(Es�&�Ϣd��F�\�ϐ�j{;�ͼ���$R�x�Gv@/���r0_�|�Fha�Vq��6�ɨ@����=����J��e�?�Β��D��{7Zc5ޗ�
��e@/�P��-9����\�l\,�Bm�v	�V����- &ҕe�0ZX���+_�=ՙt��a��BgS��%#l�b�~���2X+��W:CO��u���_@D:�0��(�xNF1�L�3�Ѱ;8��쥃��9V䩏��,Syd��zW�����j+��̣�2��^YJ�K�W��C��:o�ϥo��	O�Ǝ~�jX��t��=3�����@���`#��,pK{�ҧ�w�|�0�\������rX�W�K���I2���k��s�����A��w�{�o���f|��M.?�n�tr�n����-ϣ�M����H!�Tb��
C+�+1�@���A�;jd^캬����,���'MM'��n������(�UVϩa��<�8_��~�o�kH'AYA4kU�|��!��u����.I-	7����/൵�z[$��~b�<�}�	��M��# ��]ų$���,I��wTN/�,25�F���F��T�y�= n3��!��q9K�%��]T�T���xQ��Z.u��ͨV}�|�-)���x(�O
��[��A ���Au���mA]�p_���=8�_��=�������5K?߹�8�Y�����h�3Q_�����gP��h,W�G�N��2��/1U�� ��5��0'<$����Ul�A���hNp�=���z8ys�L]Ov�*��K����aOh�$y��pY!2v�W��zC��I+���X7�drO�"�Pi��܁��1<TS���h
.%:EҲ���x�N��Yۃ��9��C�3���X? ��_|�x�%ď�Q2����*��^6��}�e[�V�!�nm��
`P�sx��"/���Q#ӖD���9�D� �*b`32��N1�,֭�l�<�$�}\n��F����p�����Pa#K�G�"��4�ʙe�!@�kh�`�X�r�{n_n̴���1s��G�t���)�K�Ŷ�lڃs(���y�u�Z��S�A8��
Շ��$�ƜtH�C]�������G!!��(lPҡ�����Tf�l��e��Io�̐���4`t�s)��_��h��䢔�/���é�$\���m����|'R����WesM.����c���_��˗<�\m��]P�g�}�3e��a�e�<`Nc�1��Kg*��e�\ľ�X).����<?:q�赿�2��Ae�U�1�72�({ޗ\6���z�3��HD���y	�n��~A]:���t��*��3�v����d��QLC��#��H��F���ѯ���!�Nn�Bq�%Rv.X~��2�����x�^,m��L[\����Z@L�J�K˰�l������gX96hi�>/Ho}�oG�R�b�׏�0�P���#e~���5V��R�[W�άL���8��r.ж�h�>c�ͭ�!���Ir��)�����T]箺���i��cP����z�,8���z�M�׭G�E����<��T�� �y�1�{�z?��GJ+�"���|�h�C5���sU%�:��|)A]n�&W�dE7�6bX�_�,�y9�l���F��|D�H�����Pt�ޕ}dy��f)���6��zb_���$���5Q\u2�?��PlԬx6,�9C�p�Qw�6�X/��j9�T	.~�1N;2k*��y�ODS�)K�טu��n�/�".�"x?# ��n�q0Wf\D&�ㄽ-9�	�C�n�e�O�P|Ű��TC��I����wUY��ĺ3V� ]n���q�6� �=G��vlaҙ�Y����o�vO[nP�f[�k��>���	��9�`����j0�y�2�Mhx��4tbo����K@�2��X"V;�7�^e�HN�ކ��Y�<l$y"{�L��0�k��!�y�~�B�򇻕y�U+W%|-�_�L|B�a@R z:;��͟+ �Yi��"�/s�Yʲ͒�t����<)S7;�FKUz��C��,��箘{z`NC}�U�(�b��s��	:iA�1��������v^B~j}��͗�n��#�ρE��G y��)_J+.h� ��~� ���>�/��Q`���"��:���2^�)�< 6yh���4�k�"���.
�@!2Fj>�)�a��o6'X\izm�+5�l)�����Y�Qm���.�NX�(@��B�G�C vJ�q�$�k��^H���hf#bf��~[�8w<g|�f~�Y��%�}�%�ę��`tj�^�V��X+�5&V��<���?�D��(�K�.��sI-L}N���)B��U^�*OE/�\�>��BW���� ֪R3/
U���ɑ�q�D��n�^�R�O�w�
� �P�]7jދ���r??�v_�(XH���%K�3	1��\��� %I�g�M_���߰mۣ�<���?
 =	���\�X�_l�$�.�6�����_G.��<U.o�zb�ꦩ�&���z}��2(�l]�h�
7�(�ߤɅ��@Lj�0z��*؏`�&9��Z�c�ߺ�7!����P�j2���;���O����yQ��tB��M3^���D�>��t��.�h}d�)|W_��yXnE�C���d�ik���#'�|�FE�]���	���Oד�Z��UA�;P<��иW?��~�@�#3�Ҩ9F@z�����u�*,E����ͅ��O*T��2ez��G��-��ݍn�f������P#�#A�-�����4㡘?��#��ڔ=��� ��%�#�uA�|0�	nd�v�P��pn-�&�p̱�<��6�Ȃ�'7�A׃T�(����,��Z���eu���j�^��L�:b�=�>9u�F ����f�[���7x�o��5��ˣ�B���';���gWC�'3	�"r��8���=����yb�S���hp<q}���f�dcVD��8Qys��T��6H]*hQf����J��lg�-�w [X���,=��~���hIЃؤ;3��/	M\͇�ܕ"i<Bؿ'$������Gdv�,A������^��6�:�|f��瑀#��U��O+�_X��9���?�
��%`j*W����?w:������7����i�EB�g0���ߦ���M<�/��t[��%�c45B�M~�HfI�|��sWQ��|"��H_���ۥ�#�TѝE#�5��!m-���x`�E���jG���/5��H���x���:��wv7�;�M��ImU�OffzSO�Ͷ��RL
C�T�Ƈ��.��@�"f�ʀ?.5��߱G��=w@gP���]�) �s���8�K{yZ���I`�����k���ɬ��ㄶ�����ٍ��{��L~��![F�i{�c6���w�J>BM5�����^��94cO��V��H�;���7)�����>�5)��BNHYX�&ib�7~��������˜{�G�µ*��i��fC�&���A���™+��������T�u��[��sKq���	d�d�eZ�e/�\��ry���V��e�*��VE1n�Ms<����J/�%���?h:M��W)LF-��U/�f��߄M%����W��p�u���`�n����RCR6}3��	2�ߜ��ׂ�¸ui;�֎e�h��U!�<����n�F��:��������`OЪ�����7$�"�+�e��~&r�@@���y\��w�u��Dյ�>1���?g���`W�f�