��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw���Q5��x#PcJk�� � ��Z�Sb:5�,0����b��ԉ���S�
�����GM��T�aM0��R3)Ö��w.��:��� �0m����<_L:%��;:ڒ�uCD��yY/���J=�ՠ�9t��Ր�ƒ�-�"��t��R-א�_hE�Ɍ�X3�F⿀KC�{�	�բ�Kn/+܄��@��=cs�� ��<O86�K�҆58
�n��|�/� b�9`L��R�dh��ۍV����P��s��fA�B��t����5n�.b�Յ��F�,8������
 #��>�
�6�1r��kP��t���`����Sz�rK�B��/ک�Z�X��Fsc�N�hj=4��x�����;��]N�q�޲�����5-���~��C���e[~�f��G��[
v�*�?�5$�:��2�[�?���5.�� qfz�Lw�/;&�]���^i��Ѡ��^ņh� �+�d���z�"4e9L��L�x8$� BoʖP_hOz���V ���N�:�-[������;݅5�>�C6#p��?����W��3!",>Q�N�m�@\�9�Z����Ԃ����բX�K�v4�H��]Hd�:�K�|pϵ2��Wˊ�L:�=��rt�K���:� 7e�E8��k7�~�������ԴJg}8�bSR�@(�}x�V�����[��~H���X��hR�z���?�l� 1Up7����eK0�T��>�xH>�,+�vEޱ<vH�H�@?�{����+K��( g��u/���l�Q=4?:4�]�@9�<O�/������<@sF>�te �#JUA��q:ݶ��4n�#܌T#;�M`��5�U��4�֌[c-���P���?`W�e���%��]FUu��}��53��n��	$�(]&v��:hh��m��-�D�Fvϊ�$�C�����Dhe�:�q����"���zy��\v�� =UT�_w�ߵ�����U�,g���Q��T"���ͥt2V�𘆅`\��/.̀o�'|�����V�����}elck�gG�d�5k���x,�{���*š2�t�뤥qO�6Ɖ�B�`�W�q۝���6x��hY�O*yIs	����N�}]�ٴ�$�汗2p��)u�������Mʰ�c���ï97�Ϻ)�	Cpv�.:�Q�ߔ�H��0��y�pĨf䖟��]�����D�Pw=q�uS@��=�&�L�p�˘"|Ԏ�=H�Q�.��dN
�L�Q��_�!H�T~��u��2�ć�_�]��PR�bԓ�f��a/Sl��fמ���nl?�� e�V�1A�JRަJ��x� ��;FWPr