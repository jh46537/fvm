��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQG�.�����=����A�\�r�|Q� F�ׄh��)����b"���!O@��-k#�W�/K>0�>cc�|��B��+u�ˤ�DM����7���C7 w��ݳA�����AN=�&�A����/���]T"ʼ�N���B>��L3ʃ2��g �9Zh%��q pUs�2>�W�N+�B Bm@!d���GT���`W}<���y�5���U���!���2���A����l�#���cXh�ݬ��5�E!4�^��R��2�CF_����WH��*��t2�Y����أ�����x`��|/������ N���c,���qّ5����%*���&���]�d���5|���uH�6��SCa�ӳ룢���B���Q'*��6P�7�{���;�;�.+P5�8��P�H�
�z�Q6����?9	��
e�S�hC0۾�Hgæ¤��*��H}�<�?�\�{}��2�a�6�/[U���Hcqp�v�/����?�{t]K�=�|_�!���Ա4}���U2�]^J
�PO	�!��`>�"�@n0�v����)Y���=	�h:�q����TH��WM�h�^O[���HBh2�%j��6��5�����u�:�����$����gƎ��ي����͓���n�"^�l`5�~��� [O�u]��gz.soF �;#�I�{��)������Vc���g��U�}��ؓ�e�Bc�3�62�8Y�M�?4�ܘ�8�=9�Rג�~�T��nmk���?���F���f;6�F��w�І=���/�
u�J0��l�����ZJ�7Ӳ�ўF��?$��K��}�~�<��B?�a5����'�# ʮzar�zܤ���aڈ��^Un: �=�J@��|�k����L���Z�(­��7�4��Y`�ݧ�r��l{�������-{��7o�fe_��J����Q�&��v�ӭ��Na#&|�zB�/rҙYW�R�}��2M�R��Z	�H?+}��!�<�<�v9Z��?��Y')���Jь�K�]2�:$PݍP�8����q��^����+Fz�7���2Ҕ��#Ɩ�L�	`c�gzl�����~
�K�\�=� V�qY�Y�j���7�W�Ee�-�BGL��;ނ���$5����*;�$��+��M����#�&�r�]��Ot5����軭B弻��<��Ⱦ�f�ڦ%���GsE�Rd��p���=� L>LeDQ^ܞ����G.�6�DT�-�]�Z�%��e���6лD��5U�������_��'PQ-5�%;�a�o�1�֋~�b�p�V�j�I���@u!/0V���O��S�������i�~�ݽZ�cxt�O�P2�b��9�wA���J�9��F�3��%¦	�O҈��c�x+Ǥ����%j�K#�\|�SA���\�XtX���� ��K�+-\�����ohh-.���,3P�9�š؎G�`:����j%Mi���"w&�F�;�)/kͣ~�^����D(E�/�ױ�F�dib��7w\w�b[���Ko]��n�[ceF#�n��'��¬w�����\}yճG3> e�X8I�����m��0����k�Eע �B�W�ke["��}N\І�o��iچ��+-DM�Yi����g�{�;cBqi��`0k�5���{s�|S�/ؤ7����{!
#����&�f6F�R_�Z��;����O	�L��� !��Y q�/�΀mi��U�И?���������������KD|܍���w�a�I<���0����fcio�g|��%|�:=o$���:$;��x2��®����|�T���ܢ��r�P��9l�#!���N��?7�$M���5���>�ޫ����
���s�M�6Y	�%�_7��V�/{X��'��y���>v�Y���:e���H�E�/g��8W1����a���WM2���%@��g�)}��N[��j�>zC��Q���ʙK�3׺׵�d�i�C���!3(R�c��GL�����Y������` vB�+���+�XE{�����p�%~٧s{��j����
�!<S�֏��eW�M)QU�G���n���y��L��p?C��!~�C)1���)<���ۿ�QC�"G��>����J�bT뙆�C��i���;��`�b'�Yd�?�}��P���];p�2�AQpg�_&��H$�#H2�Fܡ���ȑ,O$Sx��D��Q W�=ؒ��8lvD�#t�ʢ�����}����R�9o�LgQaH��j�*O]<���I"��O�������0�*?��7�g�����r]ϝߪ�J��j�E�fū��d������xqʫ��<"��xD?:
@mo�h�c��@�������բ:�p~�N���~�K����a86�0`���E���N���t����=�Nab|1�*)��[��L��5�f�t����I���WFݑQ��ʙ����b_�(��~>��l �v?�Ny��;��䎞yt����C���[,ڜ�j����9j��s���͂m]��q��H�=�L�a@U+�ȡܙ'=fx��м��%�l������c�ҮGɣԽ�r���`�2�GqI�������0*2��iP=�W�LTt< 7*��p���9}
����@���٢B�?����D\(���gKp�7� ��L��8�x�_��_'`3Q��ot���k=�I�ц���lH�g�g�\�L ����lE��&�Ŋ.M���u��:ވ�(s��驠2��J!
!+��ND�2��~��3��^��a��K�9�?�f�D3	��צWO�)�B��#�V�uI�.����(}���}ȽGm"�.x�g�z�7�N�u����05=�+�x9��ܥ'��5*W� �Gk�y�E�,+�ԵҶY��.xw�Z��W�k4e�k6/DtUm�7�1��J��D��DoU�x�Al���������2��^0ު0��i�� !,�C�,B��#P�x�Ng#���(&�t������$w�2� �:����66�T����RCwh@PO]C�Ѫ*���$^�V�����{-[��
�N��R�>��y����������0��РB�{6=�h�����?�\A �<����%DOA��0��Ǯ;CiSw}�z�1#F������K��Fë;�(�y�L��\OZ��H� �NJJ�;�y\�0����h,G��V����d�`�a0	��U8�֠q�F.p���*TwNq�o2�r�!½n��,�[�!�:�r��<�eM�9Id�?	�Ҭ�� �6�m>Rm*�=�>a���@*f��_<��?�X3g���	Ϯ�;x�'�4�Bw[c1������h���O��bܿ�-lm�<��
�6�}�X��Z�G5�s���,��^�Ð�zsК���Ë���!�)�ȷZ�ފ��/��!S~�J���|Yk����v�⻟<��pj�0�N�ن�K�Y����R?@�8���0���XB��e�v����(h:m�p�FA|��7�Mw�%��Zʠ��Q\�+�lU���:�H�L����Z��:�Mx������Ή�b��?���3�.T&��C����<���Y���">V�R�� �;j��N�r�9Ψ��a�ޛB���Cî�0)S���1�$���U�Z^AD�L4W�`�"�J1�؅���*��d����A�ذSu�h��h� q&^E�X��9DH ��̊v/�1���HZ*�㝵T��<��Ϧ��n����ڶ���q��r=�����6b-��O��~�/'p�p��Ր@t����.�ʫ��E�'�m�ۨ���V*�:lG���nD4燔����N0�DZ�ldu�đ�T9��� �	^^}h+%Rܽ|�S�����JAc�m��N&ܐW���.�"�YS�W�$�EA��{�%���9�����
�F��D(t�(%P�L�y���W"��Ł�A�;��s#��M~��Ybd�>�n:�&$�d#�;��R��6^<y���]ܘ虏c�#���X��]�]s�1X�� ,��<�����+p�{�����\'��;M`#^��S5V�v��|N������5j�D��Z���=.9L#7ύ!�N��=Ka��񉪘Ki"�BuNj�^hR`dׇ.��l�cZh�\���{6�JX$'0Z���t���=����3O��K�Fz�Uk%��I"��B����؏���!Ľ�}��B�6u�5zR?X̀�A�5�jW�~.�}��hA#��'��-�׽�ݨ���|�����$��A-�vӭ��n;���.�G�fSl�_�⳦�2ik�g��m�<�[-n�]n˿{��q1��~0-!�_�c�8�\��}�}�𽡝��2/�}�2wL���M�%���IL�{�[b�Nc8B9&ta1�=T��w���7q��t�M��`�;�;	;�^���(�0[���fXԣ��i�8H;�6��6(&�yk���`K���ޑw�&)��꫍�Q$��3�c"�K	yܞQZm��0M���R��;�$q%���\�Fʑޖ.����H�,�BK�c�E(ZX�mgfyN�뤴ʦr�o�E��tp7�_*ċd���s��m6�\�s6&��G|��r}��G3�~g-���9R��e]��tJ�c���EZ#�<d�� T��q$m�"���G���׏xo 3��Jk��K���;NP(�<1y���.�9�k���(��5�K���͸U5�җ��٨�Gq�p�ӧ.ӱ�q������a;��/��!�g$u����t���˷���:��7�2O�;E&�����c�Zjmݛ��36���7xl[��A��F=
����ݺ��u�Y�� z�,��8����{��`Yٶ�������'DTR����q�?m��w���kA�R��t����Ql��D��'R�H��?�|<�e�kܜ�ܠz�>�O�\�^�&�t+h��@`�FxX�f����y>�o;K�> |<q|m*�P�~Aq�Bc�^Hu��ݪ�����ɕ��ĵ>f�d������*�l����ɹa��L4�Tky6�,����#h�I'n���N��� ���n>X�v�G�����	�=��h>uFߞ	k_P轺��E�!1L*e�-�gơ��3�^���7�h'R5n�h�'�y7�0�H�=[On�A��߰�u�D����O�9�r�1