��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B� �⡐*��D�k�(ʸ;+.~/jը6���1�@�P.kZ��笩� �hC�צ�'� �.��%�x�WOL�^p^��L���Iv�shI ��>�{5u�����9!cDn^D�9�b�mp�r�|~f�l��j�5��od95�� б��P�a�f��>�l'�w?5!^il@^+�>L�a��*r��w�Ś�М�0�P�c�͏�B:�I$ZtE�Cd�T<�	!3JCǮ�8Գ�1��t��>o�<��������vY�s��R 諚�̪T����fo���)�a6��l�Y�A���toq8�rݢ�$:+�~�P��# ����dAe/���A��ӳf���|�K�F�!ϵC@w؊��)��ZG����Ǣ[M�iS���Er�S�����§md���k�sR��C�����u��촒�7%&�	�uD+Y�h�|ٻmz(O�:[,3�Sq�$��U �-�+@��֙���^���}����CUV�+�*��s��~bj4�|���yr���t�}1}P(*�lO�L�OY+�Jt�bR��L�qn��4���c�멏�?����#B�s}��ժ6k"2���qpGBI�	��a ~�'<��?��wMdT�	�{���\D���%�q@�]����v�$b�\`鸃�ͽ�����?	X-��b��%b2Ҧ�U�o���`P���@uޯ3VX\�H�)##5&�Q7�Q�џ�.h�	j�yI��Qq*s
!ϟ`��'j����`VQ���ˌ<Gr�c����J�{���t���Z��ƞ��.���͗ (�_#��}�,����L�maV���1�ȅ�C�E�ME�Gj����x�?�����2fOȥd%S:еα�=���:/�k/{%��A��Ƿ�=����G�bS��,&2�C�t�������L@�����'l�S��a|I��|�b���)z\�&���D���!�?kV5 ��{Z�5����-}>k�0 e���r���P����Cȅ�ƭ�m!��g�8�jNoK�l ��y4�R"2�d��7�x�C�U;"�X�6 ��]@�뙯q;b=� Uk5��L�C��q71yc���	�)_�YR��9G�(w���3O�?��2Z����(QA$+��CVqM�꼊uqCA����}eu�O~Y�4%�-�R���-275\��\���80�b/O�NZ�6|���N�L:� ����z�Z�!���&]Q! n�1�o'�%�Y �!���j�-�����w���!��:�BF�=��X��}�����'��z8���m����;�Ԇ�( i������O����O9��;����8������s���-fP�[�`��ȃ��;+nWmDS��c�T �1+�F>�WK>w[����B��dTt�J~�g�<
�Z������A��I�q�����f40����u�o&N�>�Y��В%-v@p�WZ �$���{�]�a�Q�a4�X�˸��T�ki����D{)b�.Z
A�8��v /�ދ�\��%
v���p�c5{�©'��� �n���}}vC����A�7��ߚg�Q�l�O�olڴ�U0�b�;)�2v~�/4����$y�'>�ӯ���)D����p(hH1GvR�r��2�uhB)u�!*] ��b@��îKo��{�=7J�}y/��k�����&݉}lr��K���<{��#�g�%�z��iO��m��*����2�M`�D�Li#�x4�4�����R}�[���4�R���8�j�^���)o�V�����O3�>��ڼ��j�\9���J�l�Kֳ	��9S����ɝ�"��|$Cz�.������a]�?H�ƇJP��DH�R�7��<��v�6}m�G��K%��'�H��/T©�xX����Ι����dn�R\�%��]\��2���X�����ͭ����V�nS1�A��PJ� L�0Z|V7x7 gt	j(�m�!%�y>�����l\���d������|2� 2�i���fTh�����b���
��P^�,@�
<�/�ozFN�u������Z���D޹�9��J���S�a
t�$��9]�uu���x�Ž��\H�}$jge�� �L���	l�*�3Q^q�haM���HM#���u!�-��u)'� ��a��Z*�N�Z��ڇ�eX�j*�`��f��K8g6X��V�{v�)R��Nb��P�A`�$;�����Syn
z�k��7���r���������m4��Λ���wb�Z��=��5]B
}�!��<���j^
l\I�6����
�;�3�Y%l��H�U `���U�ɤ�Y[�*[VխSqm�K���Hþ��z��!��&/e�-i�������y�D{�.P�k�nG쀔(�����X�h����*��CM�����7�>��N�XHy'�`%�~H��ߦ���D��R�e
��3gؤ�p)Zs{�}�B�� R���h�,���$x�m?��?=�h@u����!T��<����/	�c�:��5n�Pn-���qdy��X������i�ݞ:�kh�ֽ��ԭ�����[�@�DC���'ӏ�����_��T'�M=�t��yd/6� ס����A�1�;D#��s͒��"�a���{i�W��;l��gh]���n���{�e,*���'
�o)b��戼��d����}W�bi���C��Q�O�:��́�o`v��:�b�����'�E*2�M������E<͈�� Tu��H�\� �˗x(�ܩD��^uK�9C���'�(w�pYqm�P:�LiV����)�\��ٍi+�L�Y��ʒ��N�p�{8W���l��ȉ:h��A�X&X�em�6`��[�J���f2���������j5g���A؄�߭	s�p���uJ�l{��s�3����сCB?����Z���|����}|Y�`ǌ�Xv��\��Rs�mmv���w��y1]��c��I����`�9�
�w:�eH�_+�WѝT�Ku�U(=F-:�� �����I��=S�q� �tCjyT���U���)-��8�����!|��5q�N'��**b��t������*�_�4X	,�t��Z�S��ޤ{)/��$5T�	�	`E�6�w�����1+l"L�i��_�0@�v46�)j�+DI]�p����y�BY)�6;X7k���\v�������w��rE4����h��L��2Q�OUc|�*Ŗ�d��C��u��g�55�Dj	�mjl�=T�d�y�y��c\�+�Rf��jCm1,�Z����#U�����SO��p5hV~0�:n}�� _Hu,�w�<PЉ���o��5��鹫�@�ͽ\��S�wj�����:hpG�-�F;�'Fg��7Y?ÖvҲ�UJ|	��؈$�}q��5{^�|yM$�R�Oo~˃��S�#����#�x��m���gZ�8"�x�ۯ#V3�>V�R	�,׳���51���9�٫l)�0��z�0�^�zΗ�;n��b���ӿ��4(�Vb-�?{�o@�@��㦻{�p�s�O�r�X	��e=/��N7ײm�f�.����?����=�`�>�n�-�|�'�M���*��mT���*�qN����џک��8��+���T?KG���O6W�M/�i��ۋX
�ʂ5 ��M�ym����Z
�~���ǹ�?E'���%���� -��h�`�I� 7Zڦ��{�-�Y�X� _!bT�R�x��$x�5��b������@;:$ �G��Qa���+�~+�F���)O���y,���g8gۏ�mO����wj�^��Ot."�%1T_^�AΛ�M�Z�����m����F>�a��'��ˁ�ͮ�^����+KDm�0�m%�=�a�%��ȐGEj��>*�;H>�$ޛ�/��Ÿw�ҡ˖U��ANL,Ӕ_��BH�j�����պ��ˆ6��afCj�`�7ˑԠկxnJx�.t��o:!'d?����,����4�6*0������-�U�I�D�L���,�-����-a�&K@u.Q�BP>?0�߷}Z����8<|<&��Th���5?E���g��H���U3�n�*2iϴ��ӭ�W��@�x
�,ʄ��`T�ZE0��x��|�3�K ���p̶�ihz����Ⱦ�3�\D��j��ŷ3,��{j�˷9w;�OG���4T�2��9�y��=">�n͔��dv�ߛ��w~L���Mn8�ff�ٝ���NT�:��)Y�
U�5ZFV6�	<8��%�k&m[��+P;�㐺�����}�@�(t��?��4����W.���s������${���t��sи[�T��N]��8�j�����i��YJ��9k�S,�U�*6��;�ω]2��K��g����<������e�I����?^�B������P��!ϸ�f�'��9*�Ws�R�����kN��^IﷅP���2�~K�9��{B�ų���J�μUܱ��ڭ�����Q��hDf�&�}v�P/�,�ѵ�`��T�F��V$��UĮ&�wm����]�#P!B	�Q+2�9�~���Di�#)'\፻^�ֵ1�9�j�����=��Y6�<�A�?�j���jD��%[�0��xf6S:W��Ic	���tSr����<�v��	T���Y��Է�HLݍ@�u�,1C���!�%��%!����8$}O��X�� ��4����0�H�*{dPm���.�m�\�s����t�m��C���E��Q5��7`z>�աc�~�lX����7���j���
�5��&���K�	��R�`���7J���'dQV
��X�B沺hy�,�d[��~��[���T���"As��9��4`@�n_kv��t)���f���E1]i|�=��!+U���4���x�>��U�6�zfY���e+��`�Y��
A�DJ*6#)j�i��s@�~�X<�E��k��H~�{o;���ѡ�� �ͅ2M����!;\��6�hJq ���U�.��&N"�I��š�ǘ���Q��ːB�*���<�Z���AQ����jT����B8O ���g�=����#��1������ �\�Y�֊꒭Ǭ��fiɾc`qz�ۄ�?�I�;4�t��=�v�4?WOK���6:���<��ɲ��?Ϋ��tw�!��Wg2�Q��I-1Ϟ4,���H���v�kH�0F��o�(�������.��	hb�����Ԍ<k})��F]8�ӳ)+��`��i�>&��A�3Y�_���
~F�[�~�B =�\����<?�J��?��IaU�i�|�G���7׋A��fɺK�L�̓IR�.�Nmz-6��E�������Y�.����\�C�d�O��BUW��� �����7��0�%��9WoAsp9g�C��J���aYU�r�_��tb�`O#~�(H�����wQ<tr�2\#~��tpZ�ߤ	�oD�r��a$�S�F����rp���De��Aэ��D��2f7�l�xhy�s���V�T��������