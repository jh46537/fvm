��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�Y�э+�`"lQS7���8���:��"�_؏b�H�\d<x���S�EMo�^�\��f��ش����r�aB隵oPB�=�Ž������}� �9�K�g���[Sm���&9-�)J��4����+Z������Cx��WgN7}��Jm�1�FB��.իV.X��,�6��m�qRD��� xJ:��=A$$x�0�GΒ����$-��i5p��xw��D't�A.�s3!}�
$zk�*R�p�b�c �q���V{Nθǆd>�azd8��Z��q{I.��~L @�}l�BI��&zS�su�),ecc����=�uL0b���E�W����nB����i�{�I�NT��9Ff\�m½�I���+=���я�=��^�!@��[�GAD>���uO�����5?���&�]u�M�F�R��Z�z�&kH���4��d���,�w��Ĩ�D��f@����J��+�C�4r��MwM��燭"~l����]g�zZ��}�gȩ�+.|K!A;"�c 	�!AqN�9��az��S=��Be�̕nymw	e)S"߃PK�9�n��k���5E|h�C�/=$1�lm`����ߖ�Gl�G�s:U����ʆ�g�NJ�I�k����"���z�H���/�m���DU�?X-h�?����^!�͑f�1��4;�,�~�{&�"���YLHp@���ǂ�j��/�["�rv7� V{��Z�K5��r�f�%֟����Ҏ���dN�7+�6������*ZX>�%����S����F0��;a��t`��r	���a��_��%��[m������x��#�i���`��ч��f�.:���(��E;9�F�I�i\"���ӛE�?_��6|.��,z��r�d��w�w]�Ƭ��zj�)&43���x�p��&��uN9�*-��a�.�z�֕(x����`8�`m#>�����d��uM�$a+0Q��t�]��3�Z_�_�W\�gך��c�a��������f��=��C�H*�>}#=��ܫ�}��
���I�B��E"d�!�+c=��B/K���7��A����̴ �yX��]4[tDE�%"��l7꽐O�,�	�?�������)Aݿഌ�ل��$�nf.Ҡ��̉Q9PD��GW��q�(���4���o�B��PQ�z�]<6xA��o7���C��w�s�/[?tO�C�̵hq(�]���@�d�<��� �*��M���W�\��6�����v�w@{<��.�N 0�}V,-�)-���ѦM�񩭮����f�beS�2�&����N=>#D�3���g~��N�f*-M�9P�!Q&��kAp�!�pC`�9��F�5��r]v@�<h�fjm�n��%?��i�B�/�G(u����}҈ {J@zd7a����{�l��7#�Gi���B2�t(,Z�.`wwM&<I};J�R-��v��7k	,,�τ�qYBi�,�<X<��}�bLO����ͱ+/������a�����[?��@N�`;p���(E+^���DI�?���q-h�6��r��|�_���LZ�ZX6h�α�$����;�y��ԓ�H�5���U�S��Gi ��V�ښO�4t�ET�|;ˮ��]oE�n~��������	��s�-�Sf@�~L0�Z�nv��S-��ey�e=LI-i�E�ٳY�71S�Bg�HZ�<�\��ǮI�ɶ�F��l�E�M��+'�{��{	��fI����}#b��Ɨ7Mm��<'J�Mt,|[��D	�����uy�s�7�#����gX�ߑsl�s����W�~U�=�[G����6����V�N��v�`���U��2�7�4]��J�W=�^7�t�?��kP�/^��^bR�	����I���,4�rX���	��)��I-�U���R�g������?rعRq;��v�2S������GZG����dݩL
����G���s2!���'*�j(�1!^AV����B��㈽I*�yd%�l=�����@���{��gDG�P[Eb)=���Z �l�w�)�pl�~��;���esX�rJ�ʪO=��8��Fhф'���u�{Ŝȴ�mΔYG�RR���+,S�����ϲ�ͩ>lZ���!�9t�R�Al��(:�j>��@鞗�XRR`x*�F�@o��(��` ��Ǥ�kb�'�9�-�`����ɑ ��P��G��p�*�vu�@Nd�k}ߚa��y$�'�Q �WU�pЏfĚ�>�q��(t!޴i���sK��t���,>KR��
恐�3������h��:�Y�k>ro����Zo�}�^TӲt���WK�GAA��=�B&6��}���G�YךvG3��i`��gA�H���
��~.1�i�Z1���с����{:`-e��k�K�HՍj��p�,,�����{��F�ZG��W:(��堀v�-�M� +�d� ������n�4P�1�n�a���T}��-5_�u���]��D�Q���ƞ4G6�%V��73Y���?FW������	�T�y�����u>����:�;𒥡U�/N�A�MS���V���D�\�C��&P��)p��$by�Y3�	�����.4�?-:�|�� R�N�B�%����bʂ��&�	�`��P��EJ��>j|���rYԜe#r ��`�B̜�4��OHt�@Y�O�u�����h���\f�����HrZ�
����Q\�og�dB�u�N�����v�ڗ�E7=����H`>m`.M~MWI�..l4
�Ԝ]o2�t3�s �W�� �^V�<�n��� \���*xF�5Z|����\�#����h��޺��x�~��t��,m�Lm�,olJ��־�8�|�j��Myl$�c�at5����_4�$���7]E�vᵲ�ej���D�+a�,�4�Ș��-hV��F-ߜ?�uU/y-!3�`�aي-�`�3�kG���-��.�n5��I�aQ�����a^lG�W� ��A,?�R��J��T�K�٦�>3Lb�wf�S
.����l�"$���Jm!�q���bR��=��03rc�sw�����)u۪����úԒ���9����gLW,��*L"�7�M1\.a�g�5|^v�[���̠5(7�'4� pѦ���}]M}����ǉsW�R��	�<�6��6#�S���M�v_��B��,R/	Q��D$��������y|