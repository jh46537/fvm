��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���a�%�sK��h���/a�y���v��=��w�����:�y$f�*,�RA\��S����ћW;�U���T�Ǔ�q�0`�eѓ^����8YU?to�Pb�I�����9���������:����l	�~�Y���)���L8�|m[P��Z�ј�79Ӄ���e<���_�����^�2�����
v��;�{a�<Vx3�-�����ٍ��/�[�mg������o2����@�m�e�?ኂ��l:g(Ozl8S
�-�CW�gF�5�դ����>��'K�:���ϵA��8�l��X�0S����b&�7�%)����!�h/Sq�㾴.��"��w[�Xe2�.ƿm�?�g0ۉ.�*9D��>[ˬ�?]#��m�g+��;��Lb�W%��"�����n�F�`��VW��th��Y*�1 ��a�|�!D�+�iN��C��͖�?]b��ukƻ��P�ԛ>��ngq���GK�����,RO]���J,jE���bj6M�L�Gf	J���H�wv����Ƞ6�s�$�$���z�2L12R�=��9��e�O���2�V۠E�|�;���?%(օ�J���m\�B�L�>�
��nq���vz���[��}�o�#>8?\E1ƪhi)��o��`=�	sgl�+�����B<5L{L�gڬ��z�o52������'�ֳ$@5N
�y{���ᚃQ�ݐ鸭���ϓ�?�I����U�z��k,sU�(��C�o䟩$�sHf,������ٱ^Z��`�%�B�!�tv�%���ӡ�yĎ�o|Ϡ���	�6Lՙ#�"����.���/���shl��Ͳ Αw��((���٪H�4w4*�o�%����q
����Y�?�f֟�x�:�(3�N�����S�/W�5AF�@�M��V_�+X������OG7�����}i�O�>���&f��bv�k��`܇��׋��$�>T���-����ց�@g]bi������D\cbhKq��p�@*�ځ3�jU�y�>д��L�#GͶZ����O/TJA�Ԧ��9���bj�:�������O{,��a��g�EA���wퟲewO¦��CG�\�s�g9HX��h}LL��TV_�żK�I���U�|+-�q0߇(�'|t�K��D,�b�p]��<��C��N�v�q%����{yE�u�Ky�h8���",*;�(���;{	��T��{a�O�:�V;�dF�*�m�-u�-�X�!`9��x�<�c!��ѱ�c��Oà�<�>��B�Ir�?`Q���RM�h����C_3�X�rM����DE��7!?��׋8V�����ݳ�Sꪁ������і\�P�z�N�mοA7	�jAI�n3�H��$��K�`�#���\� �]����W{˩�B����L}���r�e��z+y�#Y���i�ej�����܇��	`�oKKvB��Y_~�F"�Gf�����c�.GF�	b�b�С����ӰR@�����>�01E;�4�^'��=�|��� ����u4�����W�3>.MpU��?D��v��4:+�N���%�|�Z^��Ss�΂k�MR��~֦�8FP��6=E̜��|*�����]d�D��>�S��r��D	�jl�<���!��EB���rY�8.)YF@�e�>Jf���]>�ƙvRm�9C�K �����n���N��H�/M^�E�P���z�!KU�J�����)Up�G^&�d��ǂ���\�շ��վl�N��E�j3|��%Sh�_W�y�}�N_��U)���"^�ؕ�ú���2�ߓOԪ�� �j�o~�d]Ch援���|:p�R)�B��VGlgBH3��ƏN4X���J�R���;��pW�� М4syG^�g�bdO�vzy ������E���'{����~�Ԕ�@$,w�}��̀��e�����S�g�;8����ɥ_ٌ�Q��w�s�˓"�ya�z�E��0򟞓`�s��mH�l������0ǻ��|*� �e��|��'3KR�^��2<tv�зI���$ �K�H�Ð-�X��dNu��V)�����A���\�����[M@՗�|QΓ�Ũd*R��~f7�����.c����뻎�~)��/R�fMۃ ��]d�]�W-C6��}�C�@4'*���E��ق�5�"Y��,0T.5�Lr�d���*}J��؛�Y$����� ���9��f��%��g�geZxS'kͨ�k�rԧ�2�Sz����[ ��4���ĝ����&����|�y�wn��&@�� �#淕�wݣ �x���z��ڤ�O�-�fM��$Z\Le�Ѝ��'Q�o�L7y-+��c�;�O[�ԭ F/���8�����9ȔS�p3����+W�O�@�k������"�'ѕЙ��N��|u��=��4��gH���dq!qwz�����{�J��+�D���#�{��"̵�=�2�ER��YCs�ot}�8巙+X�����51A��C�j���W���KV�Nn5#�� ��VS�zv�|�8�qO?��@��	��B g��9ւ_.C��Q��&;Q�����Qw*�D̻"�C !�V0�8�"I��rXAсF�.�WL�w]�=����tE���P�?�߈$�Ӵ�]��β�bT�}��x�B�� t=�ɟ'6��;�< D�II�9E�K���b���x-�p��͚��>�-�CB��w��t,ie=E��Ɔ��O���Zp��x��cȝ��;�\��ꭖߏ��0�~g�~�Y���ܶ}��jJ��>�!��wL��KI$��_{޹Ӥ����N()D����~�� 9�x�6��q�w�""�בz!��ݩ�|E�n�<��9�a;���k�k[/�4My&�N�I�@E�C�@�ty���=���5�Y��ѠF
e)�%���'�{|�3�Q�J})7k,[�������?���&�B���c�V�`Q�x|yD�$PA�Y}M�1j�"4LU��!��]y��P�U"o��^5��:S�:��-�.�V���U��
��f�%{��Z�cL�J7��U�s)|�G�vE��HY����;�TI@[O%���(�R¸
(k����bJy�;�Y�����=h�,>]c�~�8�;���_�Y�/��~�;�̀f<�����z�rٺ�#O���"F��ĎM�Z�Gs��,}N���S���`�D��O�S�_�g���Y}�{%�MɁ��3�;�k������c4GP[l
�"�MY��t<��}�3�B����h������X��"R����0��}�N� ��O�F��d���Q�g�m�̾��.C�r[�y�s���çY�����
S�G�r'$��h)���[k1*+.���\T�1�S-�3����#�2��Y�������|D��4���W��$q�i��4ӌJ�>.��[ZNj=$���?�Y���c�mx�E6,��V�z����8��͠N�`�wsr&�v��ݭTpr����:Hg�{���!�:w�@�`�(��?�C4O�h�� �u�F�	���#O�8w,��;�?�E��3���$�d�M�"�Nhϻ=�#���c9B�D�Mšc)S!"�6D�1'��鷰0c��jX��Oؿ������Ml(����ݴ�{E�R��J<f@ue]��}��X��c+9����@T��=l�����(-����S�[��1$���}鉥��(�h��HfcgO�8W�e�-�L4�C�?�j]��19j07���:8Ħi_)^8��.�.�̏l��j���wh���:e�R� ���$�(g�t��Q�p�q���ި��o�����*(0�����s?�v�k���	���	Ox)�&�	O����C%��$�B|n/y�,��[���Ș�p���Wes�O?|g<2�l^�AC]�>���N|��I��������ʢ��4R�i�)/zE=r�N��h#��
��{��[6�ʳh��A�[�%D^�u:�b��7�O��o����Zf߯��l�i�����B_�ޗ4~ٯ0Ŗi����e�����Ԯ��3��k��|�[O��vn�^�Cԉ����T7*�j�A�ۘ�Ԣ���J&��F�d��]���H�qpL�/\��9o�=�#M�t[��L�L�[�Tp�߼
5ɤ��N(�[���5�� �Γ0u������b�O��s%�7�����įq��-��𼞄�e0(��L���6㷉��ЖU�L��E���Y����Һ\�K�8�yb��)e�B&�2��3�i��jc�������Ņ��2K}���M�?(=G�w눝>���G�O�A"D�svRGPኁM��e�e_E�{���^�6͍��f�|�;�:a���MT�*�\F��C���K:���ƶ��aj�i0���A��e��ܴ�NL��i�+evQً6B�s^��s�W�y|�^��������ٲ���Eh&�J��8K pd�k��i��?LQ����K=�S��H�-��V��7gm�6�t�j���aLpz�*��h�e8����wdo���U~>��d���,��l�WVR��TI9����Nv�黓�u��>�p���Kv[j0���
��j�n���K��6�!&M�Y$��}�b\���.���'��:7��9�վғ�7�~������u�El��� �@�wq�pI�0#>1v+hևJ��n�����o�j�v4���c�a6��$9*�^�������Ź����vݹ\"o�<���xëdo���VV��H!�x0�4Y���gۚ�O5�
.?J`!��v8>��Y��M�,y����2�����=�2���dԢY��W}A�\��3��d�c�5����Ed���ό~���v��Y)�22����9%���V�=����_��n4���Ç�	���Dq$ /�}�&3�&���xc[���8`��1rd
G����W�rbM ���J��uO��~�E[Ƚp�$k2��Z�n�{�Z�9c]U�wLoJ�= �i�I�>1k�e����v�?���pn��>��Z&iD�1������g���c�܍^�H!����e>c?,��?-\��n��/:eEGY8S e���0�6�}Nd~H�&_��%Qd�M^o��0o�ߤ=������� 5.R,��u�9�ؙ��*�:�47hA�/��xSn�2U���]�Ʊ�S�2��cR���dk�6��~������Ñ���� }*�\4�����M3���%�KE@vM�;��L7����LV��X����s[�O�N��-��6�N�lG���ŜS�j�fcQť�@X�|�Ȃ})Ӭd<�'��E�#��d��Q�X��@Z�.[>��m�/a�t��,�X�
i���%��a��t
E�ϯ��yyRk
B����+�Ǟu��v��a�g�@a�A����7Gh���/9>S�t�hg���U���U��w��&�p�:]��K�ʖ����Z�j�㠢�_m$9�k����Pb���Rd��>v���`�?�J!�R���j@�lģ�#�V�PC2�~;mT�����t;"K}�.�fV��
�$�vP�R�WA7�.pŢ+3�mc��P깿�;";��uڅ�A��V~�b߷g�����#n�Lx�~�
�!Dy�~�:i(�^-hj*j ���l��U�YtÇ@��������Z�'��o忝�#�:�+���;�̷��9�G�wR��>��$S�$M���G�+��t�ݖ�U��B*1f�-��5��}�:�Q�� -z���1b
;�U�3�	�F�a~1JvS9�^�B%����v,�5H@1UZO8ͬa9��&��;��d�q�ξj��3��oe��[o ya/na� %�S~�|����~�����v�uͰ�d�������yy�p��|�6������: �:�b���KxY�&ߣP������"s1�͉��z(x8��W\x��\��}U&��Xi��#��0�@��F|3Ai��B;Y��rc�e����A����|p�v�}8�0�x��=z�֊�L����!�]�� ��VI--�H���������1c��K��4Y�w�|^�*�ND��fd� ��a�4�u�w� �F)��E�,E�[�w�����_jh��Z��G��y�
�0d�~AyW�R��΋B
G1�1��Td:�(9������!~Wb�Q(�O�9�XL�93-��f��%y��*.���<���[�
�3�_��jf��}=/���&���v�>b��0S�\5]�U=��=�Ƃ�f_�7"�ٮ`4�.ſUt�=�0ܩL:<{&d���(���vd٠3�tb�7��"�j�l,ѯ_�5�{��,d��lޟ\6��T�Q�"~����8��d�#ܳ�͑�)��iQ�b�4�%x��*9�e��}���m�����f��&=��	�a�P�z1}
q�yt����fF���,��<����҂4Uʝ\��/�Ɖ{�t��B��S���˸�%�̃�;���?�fD���&6��uF����}'6��&����1bΑ�0+>p�g�k�&�f��Qꪌ��-Q�	W�۹]����Fz9i+crp��c�۳�7����r(楝�4�'�I�}����]���|Ffu�X��	U�~�nMs���4իX�W�c8.�����AQ�*g��H\4���J�Z#@�~�@��);/+,4 ����TT���CxQ祿�N%�͝6E�p�)�P����� ��c�C`g����^�=��΋�@H�$�zGH��q�I� x�P�lq�7�x
q>K��Mu+���b�2o?��S�{����CR�4{�d�'�Ͼm~$a�gOL�Q3W�5P�!K��	�tԳ!��h��ke�M! ���o�1f�������([�,cֿ��#��P�\�jѹ�B�>O-��ל5���6��/~� 9th�^c"���O^��5/"���k��&��	�k�1]��YM�{����]�ꪑ7O�
x��>(�t�~G���y�p�{+�#IE�2�� �d��5�Q���T���f�rw�0ܬ�z����x�j�3{#J�#wВ���H��Q)3%�O���*zQ�L~E`���1�-�Q����ᴫ��S�)��qn�b$X���C����9Έ*i~Vu(,��)�&�G(BYl�����n���"f��p0U�=�`�qKY���QX(sUdY�{�t�OJ�l��Wޠ�ٍ|)��冯�k����C���:_]��� �T+�9pp�f��D���C�Q�bl<�Z��l��'�G1�qش���̏o��m}e�o4]��~GF?G--��|@�Y�)���H�N��bk�t�+C����ݥ�k _���� pπ�؅(��w�F!�M̋w[��G��o/��}[\�MIT��z���=�#'5:S�@������qas/�D$��(�Sp���aN�:S�G���%g��*FY���P�G}������w�bLH@o�5�-�v'8����8L�j�0�r`�,�8�(��6g)� ]�Cjv�/WV�m�Ի�x���9�ȀpJ&�q�<u^�����,L��%}� c�V�[�r�:��* w�V-�t/�Bs�^GC�dq.K=&޻3�̵	z�F��Sz��=�o^	nPǶ8�y	|���?�F���pj ���V��"A�)�����~V�Q`m+^͖�9���Ѻh�0yg3������8�^���Ԧ�