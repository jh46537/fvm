��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�/�CZ�08Kh�� ry�z���������Y�e=�͔��/t�������kUO��9(�?jw��RZ;��NU���[>��1����ș<^S���m�>�%=1��<����)Hcފ�=N�و�[y�j=��ڭ��k�)2Hᚮ�5�@�7����fb�G��@�%3?V��z��;�*&q��jo�P ������O��cj1*��FU8��Y�73���DP��E�_UO2����i�9�N�控ewp>��`�ϩ�~o�H �6�y��'��r�P�s���ʆ9["�a��D6[�Nc� ~�7B��^� ��zS��O4Y<CM:��\ŚED���K;$�QQ��YU6t�4{��݄|���58��Z���������֚��:f�g�����C �8"-_I	ج�u�K֩�}����q��$�TRX�?���[~�U�,Z�"�z��Ė�4cDP�#�����l���� ��>9��`�7T��7C8�]ב�V7�)���	)��
5nU��N1aݦ\��$��n�P9��	H�	F�f�Ȟ:7Ū�;�������1�dc1�7���{9����E�4��˘��Qh�Y-7�d&�g�!��R��Q�_�o6�/xk2˙� SH�;��_��B���L3����7p�kz�p��/�h.�s�E�����k/�K��L)�7Q�Y�]*�Hͱw�,
�k�w>�^'
�*C�����g��"���Zr��$R�	�U����HX X�i�=`���������y�E|H��!,�L��J�� K��#�)A2z�����N����܅UX��YL<���<zR���V����8�C�5�~-�l���Z%i�iu�1l�9���H����w;�7G2^�^d�q�N�P"��N������r�(�-睶�)l�s�16{Os�xŨ�.l���ϲ1�]=�'�xk>��]�����5q�1V1�PK��9[sk���q=��jʴ�v��-�:�N��K�����T5�����ӢrUI���>�$LL�Ǉl~Q69��B��i�/ �9]��Gޏ%a���R�d.��Z����U��D_M~��^(B{}AT�i�R�f�)]��H�e��A�2�}��u�,��a�r����Q���m!I���eO���
��[ҋ�T/����X��m�!?[�E�{\|�*`�"a�q	���S���K�%o
�
@F[6�;�R͟-�.9���ٽ�����zs`�7�Jw^C�ZI�d�8yk�����:�3$�y ���+�ѫ�Pn���3
E�A}� ��9ְ�k������儒�e��������{C��E�hW��{�ZA}���I �엮4�~��w�׉ٲ���m�� Dcy��1�ѮE 2�'��<_��c�s��o;50�<�>)C��a�[P,�:kW����$��qi��%�����\,X%EŨ����&\~�k�aE`���&��"����d���e�T~:ä@�O��48*e�b�����z�w�J�L'z���EzX���bT&�n�m2h�����Iy}L����Y���%�
�&O�Jb�I�ծ�&���<�@��sl������#���O7����GR�[>y�~�u���Ìr��ݓ@��l��9�)�R�sB�?��!�W!�j=���vI"�,`����H��'F����h|tձfB��)�iwJ=���Ȕ.�Z�s��J^<%����m�,Xz�(�4D�b3*%�*
�������U�N7�2.�#-{��/��5^��t`\���<_ r���C��e�N<q�o�ӝ����-�x ���r���Y�K��^�s�w #*���JQ�/�+uO���4�o�#�7���JaS�����j':A�cL���Ƀ�'�T�x���Xc;���Z@�
�]fa��Xn �)�~��}C�7`.D��%pT}1��S`��VQ�R��e�Ď	�aWZJ���U
?$����!+����Z�@��(|P��~�Z�B �؉�}��ъ)v�k�W��!��j���� b^��25S��`��7y�e�}Ģ��1��=ӥ2�.7�h]֋��qI{�Hj���6r� �[?PD{n�Ir���q���L�^�io�~���� ��<Y�4�MpFdA�H�޺�R-$��P�g�3�h������*�����K�[����^x\��M>��u}x &���8�1��<vD�a�?��|{J7�q�t�ʡ:�z/��"��3Fq8�u١�D�q�K�kz:3��=DPނ ���2M%ML	��'�.-!�^ŷ���l�=�A�v:��fv�X��N����,R(��K�����M�Iͣ|���Y�i����~q�O�<1����J���EW�0O��:�r�a�[�a=���>��7������_x����b���m� g��� ƤGT���0*D0\���vQGnU�,���S~S.��7�_����;��ǅ�!�z�9�0Oȸ���M�#�����C��tۡp�[�b/����0ߣ,���^fH1W�k�%Z�J�f�N�������a��]��	�,��li��k�q�����EA(]�{�k+�E�
��d�7����y&	�e�$|�o �t������x�'Y�|+�J�/���'��[j���K�EF/�`�g��Ԕ��
iF!���{�h�mA�]�݂[hBJ;sͤ>��̴��m�P�K잋��c?�I����9��<���