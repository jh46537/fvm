��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,��F�X|�ע��R$�O���Lev�O��#�t�wG�45�������j��{�&[�o`�Lnq��v�4G&pr�[����p�r�N�NHd��`�� ��p��Н���Bq뼐Qӆ6zg����ED?0ê�%��C+�60�Lu�}f�C���e�ԭ��	9p��H��lR��5I!ntm�� R���C�g8~��>�Q-.1��!h(�B�-�#�u�X�qtX0��!��ήS��Q���yA�p_�� �C��t-ܑ�~�R_�I���[�觑�Թ<��,ۋ44{�'b�H6b"" ��/�)F���pt5$Ŕ�%k�~�H�w!v�)y�������l�<[#�t�����|�-����T���|\��F�,O�~���h-�(�Mf�� �՝�ن����rԳVtv���*�P7�B�W?���BG[3ŋ���bA��+y�,h�q�ޭ�9&����F���<a�P	�5Hx��x�)�`n�����ë&D��	�Fr�� &`# �y}`L釪�w҆P�a��K�3��9���%�5�d�@)}�I!Ƕs9�"�E��]�%�����U�>��5�b����i5H�]�Q[����2��Q��j�p���o�_<0}���0!7Z�Mt�S D���Ť�Z��_B���2^�<�j�x8�h��"G�lc-���&*��𠃻���*�\a���^U��(_��p����aq���8���t���q��t6&���������ʚV���oH��b׼��6�@������Jz��^�.�����wL���V�>a2+7P�C�yX{X�Zh�k�@�������tm!�}��`��<^�Y�Ա��eƳ���%z@�k9t�������ʻ�^:�i��Jx3�
�jI�`�fG��#T{���*(D�ڿ�� �� �@*B68��Q1�U��xczj���jFt}j��]�
-�ܹ|�X��O(�C+ҍ���JC׵�δ}��Ԑ���(g#�p���Q�oo�!�hx�#����@�F�����!Y��_>��� �]Yr��G�/�m���xTC ��`gu�i۰B�.GS������ c�p�.��[9�Z�����gS�ZB�"ʲ׋�$�) K�jدKΝ�iT%����1��y.&�uָ?��w31\Y���3A��f�_#�I4y�L@��*̜���Du|��̩Ҳ�EJ!�0�Ng.Y�(Wk��7�ߜ�5��7�|�WJ���m�����t�.�uh�U
�t�6;��_Lz4.LU�V�8�����h�r]K�Cj_I��[U��y
��e�@���[6\�B��MZ3���b�Yݴ�TN�Je-0�0�W���[WK7ď@J���5/��rH�`C�Z�����L{�t�� +x(ž�DDf������y��B���I��u�#)�nx�[���$�y#]|9�a&,�������r�T�I�����;s�*B�,w�N�R�/�2��+�����U|�GS0{�J��i�؅�S�EM��6�tjć3��d��f<�*.['�tQ�WfeM&�\$�X�{o<�+=_W����t	lD�~.�$q +o����L�rz:v��Ӵ��:z%�9���QOw�g:�pHp�x��`λ�@ü�ۛw?.���0��4qL����"ہNF(b�nAL�g�	���-�s̤[�Z<��Z�>�y�D�ԑ3x�!�V��Y� �$'�a����W�P��,`�1g��p�Ph��|��1[,�'{n��YH�B޲�������C9�q�;-��&K�� 2ُ漀>�`Vd\cqP��#̣z���ޫ{1��GA�	��ک&o��]����j��Ai!����J"~`Qя����Ԡu��l��ư����s]{,��9��Pľ�nE��r��/��M��rS�Pc�o�՞�*Y4g,U�6R}�d���%�M��h�c�k#C]���o�o�+��աb�qTEw�^wg�ǂ1C�V�͂���?B��F?c�ો%��] m���|�G�7�3�C-F�P
���\�i��^��?�T9iQ:�n
�ܰ)�Y���x�a��Pp�,+�c�m�:�������w`n9��$���r\�qc�_�Rˬi���F>�k_n�F�A��g�0 V=