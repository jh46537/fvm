��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw���Q5��x���A�E��T���߇:�zoU��z\׍���8�t3�I����U"�̗�e�t���V�>&,'����e!Z�{��g��j�i��1���"�I���y��D5(7�N|_��kNI�e�ƌ�����]��ȓ�W-��p�ZC�Zt�Db�Ƕ]�o54;��'��_�,�����!�K.�}�H�x�2:���M�Ӧ�87XK1��k������W-!�S�e��Ӈ:�E�"���;4�i�ˤl���5��>2����Ǡ�ȸ�]}`�K|Ov��nt.ֿ	�CW
b���|΋7��d�saS�a��KU�#���ߧo�`���G���Gl����
W?�/\�S���<#�!�~e��uwW�жtՄH����l+�WJòJZ��<���p�pv�E�~Y}z��6H�����pDK���^�����U�apz�~H�s�;͙Y���y4�� �.M�cyP=�E��\]�D���Sŵ)j��9%����g0֨>-��_<��v:�N H�0��O�'^_���[�^�+q��7�W�^etA������;�)$����X	=��2]�Mr�d���c�^}*@L�h�0�8�Y+Y��y���!+>'b�LJ�`j�Z��^K��p�(N`��B'd�6EA��bZ�&��sR��y��4P6�a��9ZX�Yv��뮁pb��MFґ��ۋs~���ٌsfH�C���V.jFdV~�,�rp���*۶H��U�,4{g�9��0l����q���X,���~����PM��-8^��E��6�/!̇�·x.��S��c=o�zlG���Fp�v��Z�t�,��뻾ď"�g���-���:06���?��d/DQA��n���`�3�vs���\��	�d-b�/�_�c��4O2]�M������R�XTD���@�p���5�:ݒ`sf�?���OPz�����u��/��:�}ƫ�����W�_��L������Uz��cDN������yߖ�1�s�����nX���fYU�9X.�Hb:��,$}�����T7�23�k~�y�Az�O���h���p��M�fū|o���A�
����$=�D,�{�{t�Q�H�c���)@$�I��>����L:��u���)�J-H��JJP�����]E#��J�$"�nP�ej#EY����&DKn|{�]�gy���`T3�Lo>,� c@``S0��	��g��0fYRF��H��%|=.�"�u||���E2��š����s�.n]���4eSB5��[���84F9��H-��Hʋ����%<*Q�#2Y�("�f���*+�lh��ꊭ`�+���F~� 2u�ԇ}�eP�0�-_$��(�K{v�������:���z/��eVSX���*����n�V:���������m5>b� �f�g&�!��d��"�|۬���M��w�+�P�I����?!�Fح$�P�>pT� ��x*�I��6rs��)r(V��V�쪸�6��d�"���+�����3�y�E�z��Or,�8Zc�����Os�p�xx5��Џ����I�~�	]_v���ɪ"#|+�t���Fϔn��	gWӨ����_a[��KF�2�Eb2oʿ�O�Ҵ8��^@�x���ڭ:{3B@(��M��`(x�0��z���`	܍��|���������u�in���~|��>�4�}�v�y^"�1HL��
�O�e.��G(%�^�[<�:B�tZ'YL���u<&�o-*��$bLuru�7�0bo��K����+��?��1�X}s++�S�N\�s���Y&&�b.�Y�=�'��c�qF�u��
{F��ç{���4 �Cz$�T��Q'dю����̼����0)����u� �R�y���/���ѽY����b�Ip'h�NGP>z�P��X�`糴\&�q�1���*���_~�x���s��ŮA����4,>kX�W2�����Bؕ�@�&��	W[&�{I{܌a��fsNC��%�Ш�9�!��WpO���׀�쎺�Z� 4��\�y�Z:,1W�le�6̸Qpo��$�I��M%vU�%���A�����Y(𞼲�(�z9�@[ ����];e�Ɂy-`���`]��,�}mfk��mS����L~q�mA�� .䢗�k���W~R-�2�I�e�[�6N�N�aH�Xws����iL�>������'S�����h*C O]'����m}�����~�n��iA^~����J���=R�z?��PYs�C�f#�a�����_Zf��p����!/����l�K��#+�6w�Ե�#!%�}�����]}��Žx|���H��0��"}�3u]�8
f��崬��"��X�Py�vZ�4�N0+-�s}��DI��Hup���4uKʲ8ţ_h�k̿ZE�'j]vM8t7���)j�1�@��B)P΅m�=!��m����w�b�bq��D�I��:��_�����rT���S�]�߳�< �"lF!.���p4�	��^�)�����UYNt�=�6*\����9UT�騵��J����z���5�p��;.7�>�D���wTO��-2D���j)ǋU��*!dҜ�:Nc_9�T�1�95Q��^��(J�h�;%���:�	X?1w�r7��P�-c�'�,�~����,ڰ�tG!l�b��p���	���Rڋ{3��S��{g���b�Z�y% >���U�����ݒ�\'��*�f�p���E�Ly�5��eu�9h�'�Y/7��9h�˞v��8���D@;��j}@\c�ί��B&I=�sMk�Dbi@��JF�@�G�7�Ђ�U<#���xg�+pyΥ�;*֏V>�b�y��3�'�����;/ʒ1����X݋����I� �5 Q�=��o��B��=Rɖx7�P�s)��..-b������o9���'��yϳ��@L�V����	�}�-��s���!l�r��Ջ����S9G�6J�}���r��@H?� �縵�2z��4��f
_J%y:&�n��	��,D0Ƈ�FpU��v�z n��=5TP�脇���dtR:jL����y�%۸�=)�;�a37�z��\�� G�c�`�2t	�7X��a�Jy�O��0�U�Ҽ3`J
��*�Oɉ�:r�u,���t�T��M�Y-wv��N��!��$�O���h�/����Z9w�������7��*��W�r"��O�kH��F�{����'Ǆhv�|����� 7���ANI��K[�x��"�Uea.�|$��X]�\h�|Q�N)�qߍ
#S$����J�w�si�i��|���۫Z�����2&-�����
�¾�3�-k=��嗥��(�
p'����Gy�z�I�Hi�n%�����mqt�q��-��He�=l�c��we��[	��o	_F�ܯ8�+�d�:TnU,�=+D<jrޠ�+���[N�3�����ZJ����'��R[��Pȶse�}��Ѱ�e��DH���U�mI;V��Z�g�~�H;g���������k<h����r��ό��Ֆ���b�����^�5�,S�W"���w���!��˿��xb�P'-�/�H�Y�����;�&�h��1��9?̾(�V}%�R��\d���Q{>�.�2L_).�
&$)v�b�s&�"�8.�ir��J�ݱG"����p:�kߒ�ŝAmA�P��3L��G�k��>q[˕P���Kb�X�E�2���	1"b�s�j7����Fr�F���%�����?�w�`ԁ�Z?}���i��fO�Uq�ה�dN�vgX@�~�Vy�]!����V�H�����,��������Kӝ�����s���#���Ջ��U�Xd�:��vR��@һʈV����cm[׃=U��<�|���v��az/;)�t�s7pJ�ȓP'����o+���
5��".&�\���y ���$cL�b�#@��Caa�?'~�|���%����#���%��X����nL��)��T̴T[^�?�� +���B�\54׋!�����ڀ���ظ]���RkGŢ�h��X(�x����v�b�IU��?�^Xy��'�:�X������|�Y���\���Hnw�I��z�x��>�鎑f&��ǧ��5^�cټ���C�!O;�D!^2z*�dg��>�c� T�SMmt�����>�>>����Qg���.�E�`�}B>��T%ZȲ���
ƑZXP}٨z��m¶�O�����C�`S�3{�1:��/kv�M��y$��C��z�
���pp�c=y��9RB���{�eFҗ}8��pѣ|�ķ��&�\^�_䊌tP�b�h���PE�gU�'}n�'�Pf�K�ʀvZ��W�����p�cl�U��}b]+�v�������F�%��a��u��'X���Osh�N4��m?wxEe��e�s��aW,�Y]�N��k%Z�lO~�H}��>���
�M�|�]Z}�Y������7Cd�����
�.�b��ּ��eS�N2n��'+�i����9����������'���Z��c�TL|�M?bud��$��28�Q�KQ!��rro)�s��O���[Üt}���nƽ�����?1K2�Rd��d���/���	�C�l��°��]�G\ w�7o6����A��.v�pg#1��Ϯ����n�T1�i�,�e�;Ml���V�k�h��l;]n0[qy�XBy=Dib��=,�&�����]��I��j{
 ���|=�w��a8���˴���ω��`��tB&���� NiI��W-�w�6Ճ�5�$Tgc�w����ˇ�%m� U$���U�A�WC�����q�F��/��<���ʮ�y�@Yj'U�R��\z}P.
G�n*���GP�t�w��[�=��v�b�F�76Y+�����Q��e�Gw�w�O�[]���gwr���p�)�K�V`�EB#=ˎzF!�[���SϦ�� ��y}O�/kc<��<�v�ƻ^;}�ݠ�
1��#�Q���Q��ΊKQ���V@��SQ�l�Z4���Y��p@�^�C�?���x�Iv_�Q"�:�O����I�=r�� #$y�����O�i_u:I4��@Ӝ�UQ�A%����`��!��&e��O�0�{��KY���-C8��#������>��ub���*�����hB ��.p�q�c��� �#�YLՆ���r�'ξ��pb���e�,�_%e>n�m�`�;�JP�'n�ܝ�O0�j~n�#�� �r� �6���/?S�;�/`��Xi}<��V��<Ɛ
^��56p{��a�gG�eU�t�! 0��Aƹ���yb/Fq�9�S�n����kã7WѠl�Yt�<!R�����I�cA�D�捋Xm���� @qG��ݒ��~�Iwg����+k�+� b%����I\�Ы�ZQ$�=+���aah�Ń.KɊk�8�S��(��
EqM����i��K\n]M��tA���@�Ϝ�	�S9���Yl���4yb�)���y>,̹�6�VB��꾍��
==���b��#*O�Z	��n�u��N��0,q�J�M��LzZX��)��z��Sa���Q�ؒ�c�^�1	,pt�B�����r�ȕHW뉽P7 ��E���ϖ�^�7��Y�F���Q���x�����e{�,a:��mV�����i�C^�O�p|���������*��;D�<O��ޖ߃J�u@�U���Kћ#bNx���QUj2Ӳ
o���_+L^c�@���.L�Ei�C2�*c����S~c+��v� �׼y9ޝ�eÁ*���@�nm��-�Z��s^�7��A�=�or�r���k��@%!�3ZE#>�<U����"ŞՅj�r!��Ĭ>]y��tTJ�5�n��w1i��b�O���|��՛T8�o$R��!�v���A�{Ȁ��t�\!�V��n&��3ӽ�5pX�`�k�b��ϔ��=����z)���GH����_�E]�Ҙk5�m/a��a��5I�ǡOS|���E�@<�x��*f��K:t�R+�B��҄����ǝ���Sv��%��������ҭ�q�0+�(��dq��K�1:d^QO�xQ
�q���:ÃԮs�`�cAB+���_uz��c| ^�k�����]��d֭�\�y��bK�<�M�gr� 2w���%��\��֏�l����f͖�q���sRO2���D�0�΁�Z�<��{��}9+�Am�Z��;��5>\��7�6Դ���Bw�%�� ח���i�e���tQ�`"h�t���XO����&�x�es,&��z��;��6{�D�r�
.?�i�����z䪆C8��&/��J:5K��LT�L�1�H�>���SC%X{�pP�����"Ɣ�E<�_�|����7|=㬐���{&��
�U��l��gL۽uV ��_٘��Ah�/���U*o��:??�/���^�x�{�W���͗H?�0������s-<1W'6�Հ��'�ˠ!,����F�qp�+2�������T� �e��|Ssv�U	�l���dz�����-v�i+�O�nr�6�����9K�ܟ���t����t�0����O�TJUT�m&r����/�ęp30����	�\��"���Al������(`7`��Z-{Ŷխb����
�E��'�G��)x�E�C@6d�݄��=��ܙR���o)�\m8��Ns�HGw��G�q�g��������F�O�3�2�*z�Qt��z�@�(�R�a�j��I	h�V�X�������J� ���W��/)C!٤���\HƁ�$����j��̙�v��#$%h<����%f2�0y��%��	l�T�'%? 4�@����_��y�8�Q�k:��C�޹��eer��o	N�#��m 4��>%�t�O�=X��L�p�e՘w�e	�^e�P�Hb��|3�����i�FN���a|��_�r
�<[�;�JI��K�P\�ZO�-�}��Z��]p�އX0H�;2ˇ*�d����ߣ����=;T�Y^�$�2ʏ��b!tA)7~�0���>�a¼����S,|5�nY`<���>�׺ ͫ�}��
Q҉'|<�{sIWĞ�4O{I�]��i���D�P�/'�-%�4p��ǖ��q��?�B���p�1�����VC�������}V��(/��	�ӣъ�_"v5�h��!��~�k*C]r*`����KoYuz���2��􉄹
�L��A��߼��'h3N��؁ ��E,c�F��`d��w"dBv�T �L�w���U�%�)}�͡$k�����duv=~@�
��^,/[4��� ��
�f'!���c�؁��#3S��1����9<�n��hl&�0�k��