��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O!) ���Y�Q΄�O��*Ȣy�dsuQ���`�Q}SA[�.���(��<
vɼ��;4���͋s1D[
�f�T�[��h�K�"HO�¤�TwƜ|�J�tR:����p�#��;������A&�K��HȮ�!!@<Ȍ��VV ��k��ko窿ae����ZS(�F�FO��2�;Z=��t�)W�{yo��r��(�K�StcN.�����s{P�8��AN�C�/��~Y����[#�z�bEB97�'���?�$'�����ِ��ǰ[�'�d�X�������%��`r��`���8D�]�At���w	V�򴴌���R����F8[4Nj7�-���ιFUEp�]c��$W��9P�|�Ԝ��L�?�9�8	^rA�Ƿ���.�He���n0�u�+}@I�2��P%p���-���6��f�8Џb̝h����喥e n/&ρ�1��ue��Fw�����s���Sܿq󀷀�	�~��ݒ�-i�Ȳ�G���S1	�g��<�ד��f�t0-I���:oۼQ gD1M隬it�;y����4_���TB�چ���thh�bL0���]q~�����4�Pw��Du,��8n�,�045��u�3`G��볮��"�W����`�hR�u��yI&n��xc���&����7���W>=���Ű��T��+�ς7
�73�ȥP#�lm��"8:�K4�j��c��<��d�eA����
���&c.�nP�	�hy�Q� ��l54ꓭ��ٶ���j'bz~�������,��������&l$� �+��D}�4j̢�0��)z���#ef �2)AuO�3�ۉ��p���s�l,��p�J\W?��sk\���k��}�a�.�.i]�q��W���o��9�����^+@���T�ӷ1m�$�X��<�j更�UGk�y��b��}���8uw�h�R�b"㕑I`}�0B���B��v��u0ۇ���A@��D����N�Zۊ5&] ����I��-�K���_å��HҚlL#��^�p�wo�O!�`'����^6y1^��m��7���s�5���"����BM�&+��#��_����'k.�A�$ʎ����ąI�4Nj�^��Ⱦ��4�e�zg�J �Ty�hL�%� 桐e�L��ɏ3�jyBh��ߕtͼA+�)Y-��Ż��/�xf4����[�����2WUP+�ಁ���m��0�L�O�j+�^-v�Wש��9������F	������X��#�U��@�1/�g�cL�	YC���s��M��P�=҇q��̈�? ����@޺LN���g������tX�{��R3f�w�2�}��d�1�����'Y�'��}a��&���֛�)�	Bw�.O�x/�]���]�Qͣ��~<Sz�M9w�n *�^,�С�ƀC�u>ʽ8��6?�;�݆dq�t�r3�*��Eav�~'NJ�R$�D��3�Ւ�R��h[�����,~��`�ąI�!x�6 f����H��k-�B�]�Rc� ��f�Vh�L��|f�໵���������M�U9#V�?����&]�aã��![�g/3���W���YZc���jX.ؒ�֠�[�Y�֯A,��?p�S�a@ss�;��j�~Sz��ol�s��7](p�����E��E�Y�H�Tg��E�h�3�T����	(���
}��؉Z&ʬ��M�z���ZQw��Qs��+�0z;ș��:k��ǲ�|3�v^֢�=�d��! 7���ߕ��%�a�p�NXj'P0W_(�1(\� �X�yp:N	�1<��ܗ![=�CPMd�\�����Y=�YeI�/OVH���(�nW�F����34���¯F�+�!��,A��(-��`xx���#\��?֩Q�y����@U��� pzD��Ԙ��̄���gfIL�7�-P4涙�=:B*�隸S2�,�W��N�FO#���F�MQ������
ny�x)g���i��|O=�[��50N��#�H]�)DJ�X|%9�H;���y�9����w6S�KpJS��7�r:h���K�^�:J��.O�BO����}�9S;�(�{��-��$Z��s��7�qS���%6�j��$�%$���1��~�
����7��J2�t��G��QNL�p��꘢Zr�ib��ڗ��%R	و,-���g�v�e[h)O
-Siѳ@ a�2���gײ��+���̹����%R��&6���s��@��E`���Y��j2q�o�9���0���C
��C������9�
���|�ƒ�:���s��߰/�"�H��q}���u����O7�}��ܳ�M��[���t�i~5�Tv�"�J�qFFMtχ`bW��N�&���&i}��m�"b�
����/��_���A�Sb �Yw�\aύ��`|5�.��#�Zbm�	�-DB4{^�����u`S��˭UP���S�C��	~r=tg�v��/?\>fj����,�+7��O��
��������`���
F��I�.eV�n�����O2���POBrv�U�gM�����D%K�ج��ί�xxp��Xm8�s @�)�
z��_�C��IcjbPS�л#�Pp�
%�dť�T�w&IK��s��A��j)sj��p�&��:Z��$E9K�rR,'�3�3��5�cX����=}�<]3�u��I�'ɓ��|z���U ��IN��2D�xǵ�n�CB�T9 ��m�����
��
�r���{��f��BYd�#5&x�Qn�.��͕l�-4@�,��?{�P,�B��P*��E�d%�,Ԗ]���{��o+�;᫜��Oz3;��k�O0zR@<	���a��V���� vv=����}x7�.x���U