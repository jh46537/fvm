��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<����d3��i��:��@:$���;��U��zV>���=c��Pz�z0�.�٤#N��v��A�󅺱P�p��Q��9���G���p�z�.]��8(�zj��U6����8�~tRi�C����`x�7�+�O�F��J�0馆kgĶ�+��d���}�ܟ��˰#��L�F�f.St�k'�cD�/n��F}������}�u�e$&ޗ�S:�č]��b�9|�e��Z�D����-��������E%%�o�_�Xz��
�?<��Wyv���f�ohHo%-�C?�Ÿ�3Հ2KP������,��B�'�^.;D�����OP���!|�|?)9;��K
J'��յ(【����v4���V���):9p��I�-@n�]B'�M�/����_�=e�9xY��E�;K�� �*�rTs�+]���f莇� �&��&<�h���~�=�u��K���"�C�v�	x%�-qV��F	��m�&�@X-G��dy'�S3T���%�9�)^/E�u������ӄ�?���p՞T"i��c�����Va��o�	��J�L��㮇
�7ةv�'S�c��Z��uhG�mPY�����R���`������ĩ���� c���9�ddQ)o�����u�=�l��5��-{o�A0��Oqx�j����|f�q�@qX�+l::��U�m`�RF��y><�5����]��}^�6�e���q��2mU�s�������Y�b�����ԻE~��F�׿����3���G��-������iVݖ������6(�+��(��c��q1㶢-�<N�x-��cz?��TտD�-X_�zf_�_&�Z#XM�dM���U����Կ=`h��ҬO&9{�ݼ�ـ�t`K�گ�V!��,HLv�w�; �bHED��/���F�@C��Oh�SP����?��1�]�}��Je�5�!;��,��D�S ��9}p���*�⚃�x��He�I�*�/�I�g�]Y`%	2�F�{�ģ�����������2������#�=?9R�73��������zk�bx�Ċ�g^^X��+�T�.q�;f)��6Ř9���^Г�rL���6���œ�ht��7끕���&��%P@�T�׃��O�u+�e�&��
���s	�jj�&/pA@ED-�>2�Dw�2�Q�9<(B���'����W���X���y\�U�a7�tS�l tS���nO>)p��6ڤ�&2A7�w�GP�lLܬ��@�f���W��ۭƤ��
R ��*�
Є�i� ���<*!>M��5�� �۠��jZ����u�M�C��3BV�C�����Q�$b{mu*%8uM�!�������2o�i�W��(s�|I-W������G�:�Z�#�۳L_r���K�X�R&� >!ȴ�"=�����I��%H��!WpY�����d�VvJ��\Z����U�Ɉm�bA�X̲�ȸ��X��({	�s��1����*���N�iz�/��Vڗav��b�l�����-�w��*�}�Ct 7��݅��`���1��DXty/����T��@�Z0{h���fx
,���Z� C���>K�I��_Y�k��agMPE]����G�)ުhi����X�\�p �%��zK<��/{��F�-R7��#���(�\Y����Ԭ������x�^�֬!��k����1_���E�c��J	�h�
�e�@��ů�e��<XJ�RW���6�XCP"��T�~`�Dý�b�JF�W�0�����&F"+���R߷�_���R��b��?a~̌W!�B.�9rLi���}�\���WX"Ovk�"z�ߤ�^Z@9~0��Kef���!x��s)J���h赎!_&Œ���`�&�#a]��?szCf�KWC�g"K�h���#�q��J� `�[�=�~�.�V;e#LS1�J0�1Ԧ,vQLL�I���C��ZlG��|�^�2F Yڎ�85������G�s�+����<��;����p��Ǆ��U����-�r(({4�x벻���`.�Z����0����<�����t�\�$u�����"a&	�\-0|aa����k� �xqc! �!i��r�۬na�芞$��o&Iz���}�J7C�-��C\1J��@bCnd�f��c��^�&�s�Nig(W#�)=ҟ��Ws�.����i�аl�-��܅�D��ה{��H
�*II�{�p���<�����m����+�/�o� ��[A���ea8�7P*$��Gٱ鉍�	*uN�y�^,�)��1��	��3+����Y�+`��4�Q�0]B�J�.��?�
�>[���v��=�kN'y|��:o^6}�hN��b����\�~����S��	����%ྖ�hhX#<Q{����S=K�lݘ>Qv�0N.���]�c�U5}����U@jMT�l(6v��<�q`�/x�'\l?��i{�OD�n5����?��\��'�b��(�A{�Ň�|BW�
z�Ǭ�8�\�,�A<ݒc�nIz�n,�3-],H��!}��N���@�A�m�<4�Y�ۢ)�v�?w�_�㑣;~s��@-D������J���5V�h��:�;��k�R�~�#�����)ٽ�pm�������T��ጙ(���S�㘀B��K�2�t�j'b����ND�ʗI=��r�i
m�+�?x��	>��