��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ����|-��L���S�u�c�>׹y��d�ۍx��+�!7�3:K������+O �zb�K�̖�N����C��:O��ѻ�rؓ�
�3�D6|[ȶ?�����Qǜm���F~�Q����C罹��7�ɞC>80��� ��z������11���ݓ������Kq��Qy���Wuaoq�azW��n�C���I울
C-(�e>�,S/�U%�&��	��Ch�nry��	^D�e����5��z��l!���-���X	������N���ml5�2v��)&�G�k7��2`�͆��M\��9<d6�]��lh.�*���p�������S��hI��I�F�:5ss��$89���㶤c�[�sa�;)��ʰ�Y#�*|=���Z(tNP��,n�����9gHw2����>����U�B�A�s��o��r��� 7qPB{�͔{��ko"8��B�i�o��ː?}Ҩ���T	���l2�	K	���հ>��[,%��7ޗB�f������Yp���݉%�ƪe�1�Gn��hK{{am্~J'qI��_$�	�~Л-^�xmï��k�'���]-G�G!�g���n���>)0�MP+�ƴ�F��'1ƅ^ڡ�iy��0� �i�8̾,�}'po҉�M����Q3�$ri�X훴�b����" 4���d��#�L�?���~�M����$���'���o�M�:��e��nK_�	we���տ�M�y
�џ�buBSv���XN��=g�����X�=J�� ���@�U�3��l�#ajq*� �Jb��j�/��'�X�s&a|�KCfH�"f��!���#/�;����O�ˡ��>��I������j�[�����O9O�i=s����՟���Xͬ�i.A�<��H�.&�~��bҜrY���y7#�+�;صS(33�wQ;��E���Y�"��A������㿢7e`�{#�1@�;�i�T �`N6�2�x��3�K��f-��C�;�s׿���P�j8��8�)�ǯ1��v7¥�Q�!g�뚋�P���N`Z�U9	���9��&�di���D;���&��x;�Zl�i:�v�5�|��7���\�7���.xu�d_���`[z���;l6�w�o�GA);!
Kx%����ޡ
��3AjHh��'x�/�Ua2��#(�ѷ,��R��̒r�;i�ۙ���3�i�4��[�)��t�	��-�s�ɉ�%	\�T�i�Y盍ƃ�J$п�ݲ�7�-�?�c�L�-^v�5e�l:�n�T`xb�1��H �**����)Xp�5�ꄵ�5
����Tc �p^-���Y��âm����!:$���G3��I�V��-.V����$רA�.�d��Sv���g�^J��>9�{�m�Xq#q��i|>GW�2]���β���m7_�fy���f��q_�7���N���	�'�c{oF����u'��q2#5T��2-l�4�t�d٬f��̟���^��m���iW�E�dMǅ�\��n~��v
�Nu[:�����V]�ĝ'w�m��6"�wH��JFy���:1�B�����R�.�������Ҝ��>[���C�r�r_r��_�ՙ�����;%'��3M�8�UR,Y�v��L����j�����渌��fע��n�b�n�wb�t��@������Q�ޤ0�WH� "KK�J����8������r瀥ѯ����r���u�����?�}`�L�s��d7������1�h��TW�ç+3������Ts��iT�SS_�5t4JFg􎒟{�]�K�Q1��;�u�n�m}a����m�Пr�i!�R@bI���9��!+7;Q��69���S�R@�V���BhA��LV6y��6َ���쳋!���k6�I	�h�v`*�������`��3=���X�[�[�C[UW���(�.�]�t��+^t�������ƀDE~B��'�������d��*���y=�%˹r7?o��֓�(��B�� �����Xw���u�W�`�������'�2����;CCN����
ϊ�+i�Q�;��$Q����O;Н�{�RL[��u�~I� �Wy���j�ȏ�<�Z!w��f��|Z�d�\KI�DUM�DȎJ��C����ɗ@~������+��}8��p� �m�18�j1	�뙟voq��� �q��vKV��y|�2�fp!�*�j$V�����GG�ǡZ�����=w�9�XF��	E�z�0,����T���mO�?���v7Dz���S����s&K7�X���.�*/1�����t�I8���A%�kV���G;�af�N����]f��x�y!������q2����g~Rr�%t�s���,���j���D�l�{ūC���m�cz�١���B~���K���k��)VN#��9;���3�F}�� (~l���C��2�!�ОoUZ��Ɯẁ&$a�a�N,����n�s��/�1X�<Ry��kc�{� Z�	��Q���>Fo`}�1���Ӏ(�h������3ru�{'� T���rY��e܂���YF����D�o�
���t�yJUe;�#����jF$Ɩ��詴Q����gc�������R0�r}9���M��B�欺���L�'zzd�TL�"v�+t���qN�2��p9wx΄�/v	4r��K�f��8��B5��,*F�����Ue	��ߺe���,r��s�LFhI�7�I�Vj�R�o�5 ���J��}Q��#9�"�;�>g�'��:���C9��}������*o�7b�2��?a��fC�iUv�4�m$�Х`k��� ��g���.xX'�3c�������Y)�v�b�Թ�е���u�����)y�<Q?�4��N-�|aRFCp���ca�<��*��é���+���y'7�tb���ƭ=���^�(#ۆ��F��z	����Ȋ(�r�f=�t���P��*X�1���`~A��#b���r%�j��M���*m|##���|y1ߒm]��~ؚn"&��H�G���T��{�jWG��6
R�f �#�~&9<�k�i4�� v'3@���w�;6'5�UviV/����!�I���##��ߚ|#8�S�����mBC�i�e]���b���t~a׮����1o?rp;����!�f��ΎNd�<��z��u>)>�j�uװ.Fg�u����w8��xq�!�6�c���d�x�(��Ճ�W�$��-/ )�3����C�#1n����2��l��<��M�EDC�W���#�p;��)"�De2 ˾Ԝᨄ�ǎOZ,��bҌ@	�2~�_���H�rE��w�9>?���ie�mX>�-��e��뭱ϑ�*&�@6h�+���jE�ħr�"@�rTٲ�5Jn�e$5_>���r0�c�4��*M|U6T�=��G� |�v��[P�zv��j�j�^-<��[Q_��>��=�0�7q�M��>`��0.b��4e�"c�9�qAxd`�Tu+���=T�?�1\�H����(��.��<d����P��иt1��)�u[���1X�`�XU�C���fZK��
=/'����0cl����'o�4g-��l�a�����Uq\�faUI�ѥ&+K(��J4of�"f�pB���d�5��XC=�������ro�Jh?��c"�(���ro�&n�����P��*Os�$a9��+�}@х��&*Ҍ4�7P���ϒu�,	�0���f���A�⡊2�cmU1����fuX�j�_#ˠTmj�7{�j�_�;����*{r�o���z 4Z=��0_����2su�5oD����	�w�0_�gC|�g	1�B�p�{�Sw�2x��}C�I�l�V%"8P W���k��(���j�'�����|0�!��(��-�-%y[U�@��:~�>�B���� 9��:�w+�U���L<O�2T,����jY\�d���7"��5*���f�9��*l1U9���-�G���Ó�_�̡7����7�;f�~�KQt1j<=p�gTFr$�`�]} ?(���SU���O�
x�2,��hJ��<_�Z��b#�b��T��P5��5�C�~�Rϐ��֣nC������y��(渳�N�7��uD���Q�%KL]�D'@�TΝ?�U��R�x�\���\~�g+�RF<?�^�Twm���p@�+{�
�u^wODi������
5�c{�/ ���ҫ!	�3(�p�<,"(��Vٸ�$���~ �����9�����4��tʠ�� ���l ,2�����r�	XL����(�ɴ����G.�ef��b 'u؉cX�6B3�@P4?�U�.�
�l�i�n3�N�h'U��wP)�([��E�}K1�v�!���Q�t��z~'Փ\��~��;6�U�1q o>������+�`��pk4�үL�&�/�Lx%����x�!l��E��ml�Ϯ�	�8j��0�G�K2�q�3�a\�rgQ/�.�@��k�P��m�����B���ԌR+\�.)|Tj5A���$,�-?��qB�tAs��.�u|�gl�8D4Tt��iQ�`��J=��K"LT����+��%���Œ�����s�uNAʬs0 ct���%�U@�}v�t|�?���{�@D�sh���}a����QtF ������G��������ؓڹv ��,J��I�����m��!��!�����=g'�ϑ''�8"s�&����{ƭ@K4df`�Ќ�8,U��a�c���}����=�Z�J^̅?�KQ�P�����!�Q������9���:����������Kq��Y�ы�����w�nɷ'䣌w��6��t\�`^��!f���Z�Є���k}���q��������NKD�h�HG��D�x�� �4sC��-V���U���wld��[���=��]�}��������'rh�@��0*�N{F�3�X��� x���� �}��1�Ó��w�ۋ5^F�����Қ�`�a��I
W�i _[���	