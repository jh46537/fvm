��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<@��݃VQ������k�w�
��T ���6Y92;�R�3�C��7$���]
�	��ݓj��t_M0�+ob�N�VT�Ϩ�m1�8qV ���$ۅ��|>� "컃���=}���$�]Q�t
H��ip���J��k�,����/?!B�=T�zmȮ�p��9z�(�,�%��f���`�k��x<~Ц��Z���Tk5n���y	Y�E$� -�M���Q�"6;���=]�n/H$%nL8Jg�RXphOAC�b�ᲈ��H鬟���e�ǟ!�ק
O�J+�i!RlQ�\��`j3�/ņ#<�G��$��:����9�n�L6F�i�a�9['�ͮ�e��4�ȴ���M�V�?9�� �? S���(� u��`�M���<Ʈ�"�{�C��¡P���B�m[���*�7ǟ!B!�8�?�!h
�_,���_������Q|~�le��a��C���,K6�!�"�aBb�aw��ڹE��Ҏ�8�����~�哔�x#�*��I(:O]��k�*B�������y$ƻ�[h�P����~W',ƞ�z5�	������Y{=�RN��k���̕�KFI^�'g$`�:�GW��zv�Z#��E�S|{@�I8�._\����y������5ʸe6⫾�[�����כ���@4����'��^nnc5N:.��1�4Ͳ$2�Ԣ|��w�:��B�T(������f�]c��o��z�����$ ��y䧱��{�ڮ���ľ��n�O������'b�ީ���6_���O̔����(�:`������V�� �!�?��y2"IO{�B����C���M��Bѹ���+������᠑�]��(�~���h-@�B��W1�Ŏ�~$��mk|��/���ھ.r��^�Sq�0� ׁ�`{�%)�b� ���u���pQD����sV�x�d+�� �G~��}���ZZ�nЅ�s&Ba����)�(�⭋���^��C�[c��s�JZ���8������Q��*��#�osIt��[1�����*eRW+B����.bdV��]�\ϫK �o�DvS*?Y�7�o�g��c�#j���Y���se�2�/5��2�K�����`� jYɦ#1��y$����%�*�$Üm͙��$�M�F»�i�����-�e+;S�o�}�8�|�L\�����_,H���B�Jo]6h|@�0���r>T��4#�+h�<�h�q�evk,/Sb-�d5�N�x@����j� �ٟ��@�]�8U��7g�����C5H$(���J��j���E�0!έK���V��gpD^U�Ie9�U��`Q�Ge����-��(����t{ZRL�2�Ƙ���^��}\�p4�v)�"D
�7㥮,	is��T�/�JeWiS��Ùn��u�ר��`Ψ=�	�P���w�I#�ڻ6���
&� j�.-�7���Q\���TSDj�04�i��\�3��Fd��t�B�6���c�����n�iRv�p�8�d;�?���v@;�! ?��)��:�?��1��!^�\w��>�9cX�B��?@�m'�B�-4�t�������GB7I.�!���a������G��t��T�h���=�����^@@�M�w��c���a岲��7���RZ�a�x��]��K�DE����l�bk>(2̕�1;dvA��pc�⿃W��ik3�G�+7��/b�=��d���șv%��i��~T�^[ձW\�.��)Kc���K�f���(���f��	S`�a�rl�|ߟ����
�v�t>m���
=]����_��B}3��e|���囷ֹ�:e�q�!3�Ϧ�Y3V�F�#�l`��
ʩ�&d7'�R�v(hB���W&z���I��D���V���#�p��ˇ�݅�	����4�3jf��ɟ�5w�0��.�0�[DK�@�`ti��J��;�C�N�����Z���=0�<�{f1L���%�xN����0�� f�AϠ���=�f��b�Vt�^�b�b�b7��4�x��	�o��E�I���N��/]�?.�Zm~�9v@l/�K~��42$0IA\���VFUb�\D�v���ϥ�_F\6R��[\�؀K{\������e�/�b�j��R�;�(;��ܪ��(�E��\��iF�n��_W�ż;oPH�as\�[=�Mp{E	1F�H�#;vԿ.I*ӆU�U~����hc�:�{:�(t��tO�������������8�
��$N\R��躒�l�����I�l!G�T��<��0f~���i����d6�㲳�r9��a;�*�p2عVo#�W|m���97c9/�L�<b�"�_��^#�8�d~#���2�4�����f�O�TD�'��{��D��,�n���lR=��2g��ɯK� !�V��^Ѧz�*P��C䜄G��a�<�f劆At��}<h���v��B�jҰ�@�*+f�Qͬ�g��D��6������ӕ���!�( C�X��I^
&��x�R+uP���^/B1,�S�q��fj�)-��]H���������f���d�j�b]�^HhQ��0C�h��w�����78e����|Z�3E��S��h�dP���6�y>�q���Kؠ�x��CNPNY�9��x>i�d#g�3�=���sF��}���ǹ8�]�áݽb=�Cg)����)nvR;�s�I��m�g��Q�3��hb� ��D��������%+��� �����ʟy:8���RĲɶS�=QW������57+!����ш.��i~�'A�a�n���LPl�0�ލia�_/>pO	�d� )|-��F������7"gaF�\.R[k��E����r��k�"��X]ɔy�(8p�tEh7y�Q����<u�,�Ts�6=C�z�}(��k5���wd�~/�g����W�����~�v�F/�~#]=�20z�N�'W]Fn�T��\�5�߈5�K~�A��:K
���w�2=̻{����-���đG��F�AM@�8d��]���k��v�\mR�)�B�h(���\�S�6CI �}~���$F%oq���}^��-,.Y,$�r|�!�f�!��r}b��.v�V�h�7�1�(��@�����-4�s��0�����eA$��������},9|i�}ۯ:e##7qś\zc�h�pH�}"�s��0�
��п�f%�r�/�[q/�~������U>��q#ЛpN��!�� ��Q�ĵ����u��w�̩�V�m�[kW�sV�ѕ�v����⪢k�k�z�^:_D�"�1p��-�2I���D8��u��@���q"�X����x)Q�z�O�1��g���t؉�A�ə k�BQU�6�p��bqA��8�:�6b�qD��e�?��yJ�#�hūѣ5z,\�%X�1Uڀ�c`5��?3#��D��Ug�Ǳ̰�n`�'��C�y�{��܋�L�y��H������gq����M$d��n\Ѳ@��E��"�tH(·�)�j�V�I`��B��qnKs��ℂ/K����yi��f�4�ϓӼ��ԕ!́�l��r���9[���{��v�층$��;� ��j��� I�'�V��<���sP�����Y1�;�b����D9�#.�d��"I���!��ب:%��P�)<�?�v�+�Bܧ����k9,V��Z��8�5���K?� ��(;����Ζ�:����W��cLEˁ.�s�"�?LF��]�G(�U&*N���O��y�=g�'S��w�3���^�U� �IMf�y7_�|�q��j���Dշ���9BW 6	C���m��n����KҘ�b:rR�^v�"�@/<�q4C�I��VT���q�I�_�%��g��-!h�N,HEM�6?9;kz��%����ZYJ[��SkϮ�E/
�]aN���;��V��!6�����ǝn��X.�c��iD��,)%Kn��?:e})g��'+	%_W�]��[����P�cj=�aHӴ_��\��]?d��S���0��Q5��H��$��N$$[��Y��';�ż��il
��+-��|N�׏v�Rf�G����(����{R���*:;FM-V+��,���xQ��*z�	�)��s�������M#��4ڀ�
=�
�x��c ��&��5w�O�[�\�b��Z��5�	->򽤜v�V��Xy�>0�}I��[�y���R���I6�|dR��l�/�Y��V�>ʿ�����O�*�Şbg1
r�3�:_�����
f{��K�ɯ���Cʨ
���0l�:�59�l�v�~���G���
�7�тN«�I��ģD���E)ڊ-�ϳa��
��_��]n�?�܀�CY�Aپ&�u�17�Q�mb�����@��	1:�s�$-��;�:��^�Jǽ<J���X4�T�f7M���c=����Դ�^�]�8)BhSCl	�?��I�!�xLX`O�/��Y�s6�ByȾ��Im��W6aPħ7�d/ͥ�ȁ�>�����T��c5{�	i�4�S�������Il�$/�F;�v�#�@�7=��ȱ�2��z(,RT���l�YM�~<F���*�px�)����ʥ0<��������a,3t��l��=�����䧼@ƅ*��V�[���d�5�kK���u��X^��ߨ�?��H�~I��q�5��H1���:����?�-��2���ю���6lY�왉(f)Tf��u4���*Y��-�Q�V��&\�ǒ=6`XS�a�@,`� ��I�� �d���z}R��!�I(��-Z������p��]R��?��bX�j�y�Wӂ���F)8Ь=S-��ߧ�\�{A�S��d_%zo<
��w={��<\�]�˿���[�x�E���:6s+dn4��_�X� -���F�M���v]}2YvT��סڔ����7|�Ƙ�X��j�{�v?�==����M�跔mҏ/��0?6����IY	�L�*�@w���Q���tC UeO����2��@�qKݜ>���|��0`Ք�ċpߵᮿn��zE�$p�~�e�g�3�� ��O���fǥu�K�����~o~������x���� ?L�.�q����2�� N�>��jx˲v���B�"?�O���3y�� ����#�h��u�/m�!Ƒξ���o�.�K�Bb���u�n�\�\�-������@�h}�;@�jU<�;'Z���kG��yo=v��8d�h�h�0H-��i�E�K]���;�M5R��ü�q�O��{��C�jT$H'5|�/���&H���n�+z�%���F�����D5��{��	+�	�����\˻�/�z�}��������L��:���ԦsW�K��C�k�9]�VġXn\Я����+-A1�~�4Зe يL�V���'Yb�{���Rg�A�7ˇ����/L��UX��e�7mk�Ei��/Z.�2�2�4����dgX��>_���Sb�ӹ���8U+� ��-+�D�F��;#�^�ڡ���;���H9�7��D�s�S���&Xg��\@h ƌ�����Ց�':���ړ~�g�mÏ�ݞ�!؋ɽ	ol���U2�`����Ĭ6��H<�z�Q�e4	_�X�t�h9��*x�ϓ�i	l^�����<+V���М�ANXݜ�&)� ��e�	zG�v���>P�d�{��_l�)��_>k��d��%J���m�-�G��
�{��w~� ����/u�;y%'(�Yj4�L�ss�^��MK(p}?��8����a
<^=��\D���h��e��T���=��]�>=e%nt��e^�	����Qk�41+	�LU��k gY6OH�Ϥ��������"�M�/�S��dIkU�d����⹺��W�͊w 2��EQ9PFu�X��pퟘ�vd����{��d����cEb�W�B��ٵ�Q~P`��,�i��J�CN1�6E�\��|$����.n����^�8�y��S�{_Z����Y�M�b�+L<%����I"��B1.Uf^�r9�fgA6���J;I�7��K�Q���fn4P�#1�y���d'P�e]^��X�\�`IkJ�Z'?cԕj��4�:�n�����a��p��tQ�nPR9{�!�O�����D��[��D������H�����X4�+Ѧr�æK{�#o'��Bi�|�X��	<�I��/͐0���Ex2"�h���vQ�7X��N����ُ��_��I>n�K���eHBpl:�7c�/�z�ѩ�&G�D�+Ļ�1
%�i1����1��l!r�z^U+	���h.8��ғ7}[�'i�mS����l���C��m@�w�u��A�j�[��*,��4jKe&}�c%i�<N>dT҉�*G���f�?޶II((�c[Kp��&�d� ,c���:.�xsoWv��[���gbyH�����*����Tr�t@��(rJ�QO�d������LzKaD��b�Q&��1c��hq��疚pq�1��X�i����[V��wuK/��N���=�Vc�Ut4;e�S�;
P��^4��;𕁈󶄰�y2�&��µ�@�;������}�՗�p�_j�l)� Hdt������a��"P�'O���Gm� �dAUN��׹ځo�m��7fgZo3��Y�7fj
�V�cI0+'�X���YE���#������j�,��k�
pΖ��}WS=$�cs�/h���M���s�����A��K��Q��譅���V�i����E���Sl��Hh�0//����
�*r��0[�%�yJ.x�����̇+�x���0�#t�E��G[�8Wc#�p�;��x�S ����|F%stv\R�~��dy�����A O�y0��%XcF��W3�kU�R	�8fy�{y]Վ܇�t�Ŷg�{/���]b���&V����R��G�Z7��r,���y�%*�yR!�� ��8e~��ݵ8z~�+�,�e]�/�T��5���cծ^z��ق��9����f��g�9�p���\�>ì�<GQ�L%ΰT�ЄvQr
+�Z���Ξ"�q��pKe}��n &b%4�e�iPG_�l:�Ed�)G�W���rᭀ�֜a��NY��\�F�"��Ҳ���#9���A��Mm�0Ȁ��f�����1���/���X���̒�q0��z< ��l���Ш�s�H<��#M�8�>�@P�i�o1��琱��Y���/��n@��2*�Xsw7�;��.��愐ՠ��d� �X���pm��� ;A1�ɺ��AV�w?*�\���m���5��{sZ/�(R8�������iq��Fr��U˫�-3�y����nL���S��z-�VF��(&h���gidB��Eշ�B����W�GlK�TL���Xw1�uZ�t_�8>��dq�����>���"���~����BeNݶ�r@KȡC�.�䮗G)d;�~�rF8w�m�A^C_3@����W)��BBS���<�8���3�(�6Ú�����>���=��1����g*�K�����2@�xi�� A�������-�X6��nC�لޞ���n�-���C��H"8o��םjB�������ܕwsdS���f�Z9�����`�=%�!NH�t���䞪E^]·L �E�N=R{�!�{�����r�q��H�K�?.�ਗ��.�:��-?���d��!���A3:RBH�Uք暤�{$?�a�^�d�ǲG�*l/2_�T���]?�����j�vj�S�x��}��u��A�ba�X�����/����aZX7wa$�GI%��7�]�Z�)�M���M��������B�$��D��vBwpuS��2�5Q��C;JB�snN/����F�����(<��,��] ׸&����M�W*?��
eD6��cc�?^���sh�m��n�"����<�R�O��M���A5�'�v��20���D�бߘ�6���ɴ'��Җ�K����,."y� ;�2����]�{~��[���<ZՓX���nU�[�ڬw1�_q�+�1}�pyۤ��0#w�94����~Rk�E4�
V���j�?���[*�G^�qDVS���9pЋ��ul"�St�Hhr��N:����h+˱.䳨]G VD�������'�eZSC�V�q?M�v;�i�%�:�¡]Fb�=������D��o�هc_�C�qU2]~���#����X�5&��Z��3���L�.��OM�
�/��^���� ��=E]dk������_��dp!� k7���9Ek��ɉk���RI���O�������'���<i$uXs�;�f&�|�����!�W����&b֌vyE����ƶqG���Y4M�äfM�+f����'����-] ᑸ�{�Q��%t��J$Su�&�AҤ{�Kn_�"_��{6�#�R���S.V��TG����T�mC9���M}��-����.e��/��AZ8o�J���B�VU���;�"���H���������⒝��;�*tFz�	��?Z{��w���E�|�v?���n�no��[�$����g���_{���h]h��삚�g�w���^�F0L���(�N�D��"Ē�>�V%�;t����}�VL�$`yd��p@�v>Z˔��fNS�`�O�A,�ZeNF��~f�G%�{y������`�E��#�(��查*��J�Nh���7,E�s?{9���=Ҡ�G�@�Nw�?lkԨ���O/��x]@��P�`,i{7'�������D�Azz�& �?L	�����D�����f��gtr��q�?��Y�$l�Z)�d;O�l{�ޭ.�`���`g��ө{d(9������rL���PT��a��g��vw��L&r�������x��i��U�l,?�n��z���')�b�MEp�?����m�H\�����4¤�vJ��69�U�Ȃ8�Z�?���-�ϝ��� �NfZ��Q�s�.�By�u���?��H��;m����#�u�����p�D�ìޅ�P�A��/B7*�Byy��NB*�Ϭ���/Thյo����(=�{,�>*p���=��?j�u��n~p1�Mc�w;e̳���F��c�oD�Od`O�Nh	ϋ�#��pW�̧r�YE��$��~v�!��]w��
�������mȻ���#D��rtTR����&���J=�@	.��
j�~�A�1��N�H�|Z�|o�� ��D=i�N��6��ll�N�;�����x$��?y$󝣊�(wR��+W5��Z֧�E�8��_i�[�i��A�J1�*?����~��Rd@�L�������_QQ��fB���1p���8֢�0�θ嫻ƻ�O�X��n:1:*�f�;7���[��&�(��ᴢ*#�֘s�K���X��2x�`�h�~'3��P����SبU�i�g��rH�Cl�O?롪�s�� �����<bHr�Y+��h��n��B�>�-lη^��\u'~����o<�6:�	RII��zC�P��S,�N�y�a����)�捊��Dv=c����b���Ϧ?*�m��S�p]FT���A[�BJ���_j��x5�����3��J���R��V:_�����)�5��b��uq��?�K�>������hA��_��%H�٪�*څ�%pҦ�B�Zk2O�o�Jea%��S,֋o��V4�¾}����!��]�C��USF2�'l�� �sGe��vi�=�/mʬ���=8IHA��&��ߑJ(c�ҁ��[(���Km%Q��׌`��A�YC��ؾ�![��!�^f�h�x$eQ_X��G��`�`0Ct~���EE��������8���=��W�G��,P:RL{�ҹ�驳zڭ�@�$McR�^�8Q!I�;ڣ	*R
a~�,���zm@
�K-1\D?W�?|�qX8�:rU=�8�F�LYQ[�P�"�w���^3���%n���W�r�]2�,�~O�4�es���꫰p��?{q�C����3n7��c�kQ�6��?>/W���ƣm����F�_�p��x�C+Q�r�WD!��hw�pd�|Pu�M��B�;��l�W�-�eB�w��?i<�K$6�'�!qg�Q�^ ������s��0
u�H�ΐ0�~�+y�4Cf+�;g���!g}
?�b���=e����=x$a�F9�@´�Yx.�97�A4��*#�qA]���Q��� G�bLW�dD���)��Z��g	Yi���6����m�ϧ�8bT��Xчm+}~�g�<����B+V0]a��u�5�����ye��Pwp�� ���DX��	Y��'wO9�6�Gr��$2��~0o1.ܤ*�S����J���D��J���|�jL����)$b�N��p�дf�RAa��4�	\��4��ߐ�e*DpS41�@]��eL���(.Ϟ��H�¿��'\y�H0�m��}���ư�]�^p�sv?M���k��Uђ>�����
G���v�/5���}���rf�csp���^��F�S=��6 �����ۦ� �Uw��o�Ʈ��«3�/�7����(0)u����K�v�oq��͉P~m�ɘ���w��l�~�x�1"6^���㺁HsR��m�cE��wf��$��$.���=����2Y�Y�ҧ�a�_ڝ,�����9��$>���J�oos�jv�P���-;���ķ�&@��Ȉh��Sx�}; NP[�P�C���0%�72����D^Zy�\ŶWD%[l��^�Ƶ�������T��T�6~�� �H��<�������mA>�s��l���g8��T>V#�f}�����-V�5r�H�R��y�侎9��u���%Ƕ5�͜�������z����|~���9 �(d���Z�c'�Q����xx;wn��Qj{W_��:fy�����U1?o���n��ҷ:��SBܓ)�g�W�����We/����9 �i�{�Z�B?{�285x΍��')��1�D�Ȗt W��׀������v?���{�s21��,r��h~�x{������9`�A`?/�C���f���L%���X�_(��Xɰ�۪�ą�)2^6� �?!�Ȥ� �f�����{�i}�o �<4,�8�K�x"ц!n~U��r�T��(>��!J�ي�{m���#��p���HB̅��$Nl�s�d��5�}����t�'�(�����K%��7+������։KVe���Z�d� �r��h��R3%���A�������~ӓ�C�y/�)�2�Z���}i�i����r͇����O�D@�������n7T�k/������o��0��hs��(ˮr�_s��@=hkB7�V����?%�<5ڣIrhì�Mb�r��� |h�#Az�̕T�{��=w���yJ'�A��vP��Bb@�U�RY浢Daf��!��$�WNc��2z�dR.�"�7D��ʋ��C�W�������v�coZr����\T�ܹR�]�����D��x��4)8���.R:�[d���x&�
W0f�)�?��9�t� �nA�)0�h�r��:x�ē�7�
Uߵ��X* LbR�����˂��%.?�s��&M���Z�8����Yt~�%A��,zj�����iz�\Ú�Sq�a{�P��7O����@.7���ޘ�~�ԼZm� ��'��^��* B�e�ʁ�f��>�8B $����p��o!�5��Ӕ�=T{��[�V/���VuZFy�7�3�'����5��m℀?%���+����W$�W��i��!X�n#}���F���'�H�}�8�՜];5�R��&)]q�R�XsS���,����m��|#�oZf�F}{/�Ŀ����R�=��V@��W���1MNb�e��J����u�E��n�Y��eǉ�Law�@i�!C�e���3�w)�c]�����\KUwR
ܦWRD�ľ/NN����@(��b�>�)����O��*�;������'?�����급dZ�Nu�Jǳ�vI��4-�U���liU\�\��O�Fi�W��m7'o����԰k-����5���``���K��
(��o:���r��dr�=5in�	wz��[��pU��H��u�C�V{� "6>�����ql9'e��l�m�s�r��T{