��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^�.GJ��-��?f�b��(��ҥ��Y�����!���نϊp��=׈�kS(�?D� Y�S���#��f�����V8?�_���Mg�\��gѵ����s=�B_M�E�B%z1�����U����\�����ZI^C'���d�_ ��-[b�DU�Vյ��*�0��/�^�]ݚ�Z���r �Ї-�l�h� n��ࣁLR�5���e��G\"�JZ�z�!���0�.f ^w ϴ� I�L�J�ȷP>���ө�,5�%%�bK���>�͇_|'xƈ�&8�.�7�ԯ[����!�X��fŷsIE�~O�l�d�O!*�W,��H�����;}"���9��k�CD`Y���r|��# 媑6�x��31�_y����ъMd����<y �߱o��)a˘Q7���{;L��:�:�6�w�K<�&W�u��wK�M���b�[���h��������HC�δ�;ի'�(�����Ӥ�@��$ �V]z	u���#���ځ��2G�#�B	�}x��G��߳~��Yi�y+�����(r��ꕛߥOy?���B���W�uuB�d@�Z�ܩv��x= �ap��X��(O�vNleJӣZy�D�o��/�?t ��0��犢�?�T�*0��Z��}N�YE�1`>�	r�D*�>���NqxVJd� S�3459��]n��H�Dﻅ"��7w�a�t^|�p�v�5U->���^� �}�c��@T2��)6V豓�"S����Uf9�g�$j��j����{?��S�X_�H�_\��ݞ�D��.V�H��BF©�;)B��PX������ϒ:A�%#�#�����=r�Pvv��a���)E�yQ�r爗|
]6�HY�:XPK���(m(��4�~�y����m;z�x�sQ�4�YV�|�B|q"(DU~תK<C�v�m�s�O�|W1b���/s~�I�:�l�u�Y��.����]@B2��A����� ����K��l�Xx�ew�L�����C��re�7z)ϣ�3�VjC�=�朓i��5E�I��Ņ����>��>�D�,[�  ��p>k	��2=��K;:ɉң?����p�_�}��=�˝gL~'/���c:d�1�)���8�t�V �X�"����=p�9�˗��I_������
��&ёP��)5綢�(A�3���}�J����M㉳6/��{�揁��k����>�+jr
r�4 � ,�q2����jG.�p��<��2�N���jУ��5&C��Zk�)}l�p6N�K�L�{��49M�%�l�e0�
gss5���.��W ��%(A1�H���g�ں?|�6��|K�:��;K�64��� �9� I?�GJ���>Q�qCbŠ�Y�����X~C�J��C��v-d��U�@�#^|˽f��\�#;���i�^�Z��'��k�+�.���@O������8�qXG ���@�E
��P�BocX��+!�4�o�mNO������d��0j@�T�]�����}�ƓDq;R�n(ܡ�.p�e��P���Vi]�=.3�\G;��wb�9���mq�fe�]&x�yȕD�e��!���M��� D���bzJ.��б������t��_Pu�BdVx�љ\F�I�Ɠ�)R���Ӛ!�m��r�u�%�B��"u�/Ș���	���(S!������F�c3l��w���2��O�p�gNZj��� �TV���F{Ȏ�*�̂���堕s��J�:�^_k{|����:��H�ra�*Y���V����`�Q�JW3望�)�3��@4����+�xR��U;��l����<�|lc���_�0�,~��� 62S!=��b6��K���S�{z�5͏@E��߯K�{ȿ��ܻ�E�g��ۉI2Ov�鑧���� �P� �>�?'����	o������#l�+読8��KcC�����L�8s?���F��0����X��`*
;� &�g�vH����Hu0b���}Q����ZB&�r��U��N����Rm�<6�lp9+��'��J\�^����:Qr[��|���ט������?=�n���m�Q���y�o����:%'U�@н�����5�.UP��f�a!��r��H.x�-��b{�'���s��5�:���σ�^3�2o��*�*U F�`�!A�j�k�쳕Aά`0�Y31�8��%u�'`�Zk0��`m��F|�]�s$�+o�d]O��_J �ﯤ ��O�J���3_5ԊA����g��=���%&��ˏ`���-�K-8������͂Z�9V)_5�1-�R�Z%<S�-E�����[��$��	��\����aiI&��/d}���_�lJ�R�a�k�j�~����O�0j�d�H�T!����^�p�;�G%B�Z�J����B�x�;�	ʼ3eE�����o�,�J��Vr��k)�1��]����R;s~Mnvfy���l�#�����ME��E����T���7I�a��+��5^eRQO��,�|�]�9.8�i]�TYU�.R�	��'���pOǷm ]=vU�r���'��&΀��@�^���H��՞]�,��O@�<'�@��ֽ�}*,2�^Rv���kĳ5j3v�#ھ�����������'�7��g��k QΦ�cP�P�����p�a���>>|�%�r��1��Jyإm۟�I���ߕ��nm�E�u=��9b�g!��@e8�]R=>RA
7�wGRB�������-��NW+�']DT�z2��o�$zr�G�g��X�z$n��~
�?�� �w�^����{�.M�,#i�+M[�E�p�*���6�����Tq�Ȓ�!���f�S��J��𕡞z��Q,C�G˯C$wh���|b��qZ�5��i]L=:�*�	a����B�6Gߘ�Iǘ��|b���â*+c8�3�Ȯ�C����i�/zB�S4�~��_ἰ���ȅ�z{X���QpK������� @Eː)�f�F�����duO�A�x=�>O0S����a��M��c�[��,�ѱ"x84Yo�쪕9��ſl�J1�u� �J�;������4⫭�m�H�j�T�5�a�����:���ӰY���46���>?�$�*�^���{��`Z�E���v8�<:x�1\棊��~G��B�g) 6 6����2��t�n��KӃ�6ǺO�Sͮ�1�����w�`,�P�!ko���ܑ�>��@E.��t�-B�i��8 �1�v�4�Q�q�����3����%3���t�f��$�%1�0�pg࿕+����q♏�vF˗#���?�Cҷ�)���8��3�`�{�6�e>&&W��.�o�����w�[(�a�Qo�x+6Lĝ����a?u@�jAb���y�Tm���f�:C#% rz(+�a�H�fl�:�<rf��J�D��ݢ���}�ͬ�Jd���[3�#}z��ݜw!�9[ٴ�a���g�F�� ��!/�7�7�
_�Y��H���f2���{�>j`��#�upjΏeOtR�{�;%�`׭ȠTH�͑|IϿ�K�ދ���G�z��ݕw�Ci�\�@}�3rH�Ǝ�2.��2?�l��D�2FwU�C���F[4���ǘ*��5:n-���o�� �4�v|��	!w��Mhk��U|����[p���ˇ���*)���h`b����  ���LLܡ��r8ј5�ED?�g$�8CâZ!*Y�L�Ӕ�hV��z��_����~v�u�	��vi�uBݔG�F��ρCVZ�,u�y�8�:��¬�y��*~Ma8��O����������4����zx�v;H��M��GS�kpV�ŵ#�.B�>[r6����Q;l˳�93c�B�^�$r��ڊ�r�����Ҕ�bbw����kM��u
��E�e|%�\����s 	�5{QF�ğoX�N��l��1+�=[�NG�i!��JJc������{`�J�u$��D`�
 �J����m0f�c{hE(x��$8��ёl?ޭ���Dq�ӈ�����TS�߫�,s��������\`ʭ���w{��_�I�A�e�||6�P�"��ݠȄo"�o>l��8o]I\�d��G�W;�)���G��3�e.�ZAa��y�ANf���ڕ�2u�}&��  �m�Do�u6l�����CYV�S�����R3'C��c���IV�P�Tj)\&�����I�GQ���$յ�+&�?���?���A֘]��Rh����vb�յ��4��߁�sV�����J!���YAKI��t� �}6w���d`\q���T�5�m��M�b�U�nhߓ�����(��+��(��y_�Ͷ�(�c����O����f����ٳZ>�wF��Y4N3l�<,�����V��bKM��]a2��o���h�N���q.�����P/	���r&.��r��B����m�zJ�z�̏��O���NyA�*@A� ��l��j���/C1'W���Gu;��l�y��x���|����,)�xY�w�p�����i��*�6�/Y<s� z���	�V��4��Pb��|��x}�bH�F ����S1�s�g�Z3�����M&�А..�Kor(C�MT����H��.xn:xz�_�P`�$��ܗ�_~O�Hg�� �2A������gI@5���O��3�ў���qS�p�--�rf5��+�.862��l�'���{�:��^�j	.O]������ty�=ǿU�㨃��$��wVۉ���K^��k�w��̽��yl~|a&	3��1jP&'�u����P6����;q+�+���r����n�Z�K�4 �b�#z��^���p��e��͌S�Ё�:e��u��k��.>>_L��<�ANp�7/���w��G,ޟ�|��;�;؟1	<kI2n�بڠS��oo�iϹ5��O%����7�ި�Q�����R4\#�t]��O�[����	�6}=aS�o�� �������9:�����A^J�j�D%Ȗ��}�c�Vߛ�+��8��2�8Sy���k8��Rw�������D&���Z�����*��r���m;�3��M�www��Z��� ���8��x�8H�1R4.�a�����т"\$�����a�aay٣�Z�o��V��jK�A8��Gi�F��e�[`����m�qo2� ��*�[�t�.-`�ۆc��'�ȳum����h�M|?UxN�\Ҋf"��L(��o_�o%!�y�҂b�Ê�~��Ʀ��[�so�..� �pun	�߮s������OȮf-����V�9ݖ�&��O'���V����[mʸ�(Im7����e�r������e�p}g�][�᪳?���&��<��[V��H�L&h��t�j�ۏ3�X�u!EИH�C��?W�-������?m$s+�Ba�/"ɞ�d7�o�U�@�U^#lL2���qZ�D���A'a��)�`�Qz�<r_B�zq�t&�36�+��ա�q�k���ѥc��;�J�2ɭp[����A�n��<:�&`d�\t���0m4:�9MJ�������^�Ս�H�TE�-u��U������P'����g?o�V��.��������'��('��t�v栗[>3Xzg:��j����'�)�C/�W�g�eFM�㐴�(e�H�o�i>�J��j	�N�%�;|1�F���PR��� q�	���#mh��Kކ�z�� ���论=�}EK�����9�a���PGuxV~_cq�y��\=G�f�g�|�e2i��*�k�q�T�V��
�;�jB�t/�(�؛�f�C�������i����g�o�I�dzљ��P�f0�_���Gp��le�'��w�DS�x�5$m���IGmj(w7]���\I,gE.�h��'�3�3��Y	��Ɲ\@��rE:2�\�����雇�bԍq/8M��o���j���+�C�p���=ν����,��􋽌M���xڳz�Q�6Ek��r�go#e��Y�r��-�	x$�	T�������]{�Ph;��	���H���#���������}��a�"�@l����%�~.� �O�c
�����]h>05.ȿ!w�lo^��7���8\�Z�Կf������l||,.�}c�6(����(��i�I��~�{�n����7������^<����W��z��zn�~9؍Md�GbN=]��UP�����S`��W�l�g�[��y�TK�XS%��c��Ͻ�@>�R+�<�!]OH�Ԓ]�%~
�1i����c��5�]��N�����^���W���wF���yB�a�П�����_�W�l9�ʁ�U��T[���T���e���!٨�RUg4B�%�Ge� $��׼��c�{8��9�Us��wʑ��6G���0��H����)��^�EJ���<��w��Icb�@�_[1Z&\<�*A��������ӈ��DE~�N��ݟ��P�t�Z�9M����yJ`Km��ى+
/�;o�8n�)A�n;��8�R�:��#&i}����[�&`����WI_-�ieʌ��6���R�n��"�s�</�n"��OD|�}j�q�qN���*w��X�Ǣ0�+���.��-�3i��m�^�|p�01�#�#��/�?n98���ѱ�R�ƟC7�P��f$J��BH���]o�0�a;�!�{��Q<ҷՔ��H�zڗ*mR)}��'��'���N'"�����(�#m];Qa���d�{)bWѶn>��:��{��Bוї�e����U�/��*�z,n�yU�"���x~��OހԤ�w�!�3�����iR6H��T[M뵢u��W�b�j��*�#4�8pO�|>0�⢳����~.����h��>���e���Y��q.3M*VDT�V��양�>�^?����Pw#2�=#��J�������%�C;�k���m?���=T3F�zD�QTeBM��5O���j�-c�l2	��.s���:w���7����D���N_�!X���Nǎj�㳑6vS���i�.�
�%n�Gb��a��0�= H����*��%��B|�#	Ǽ�]�