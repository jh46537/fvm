��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�'�I������9�d�:���"��ApuiI
⶚���Z�M�� 䯨L+8����f�L�c��(|d���%��q�g�N��d<x$V�/[&�WiAq�D�d}�kF���Vp+���GO��0�a#�!���E�^�!Pqf6�Ӣ9^m �|4%ӂ0M����`�
M�r��,p&�:�p�����H]2�l�"g���d./L��_�C [[7�ݫ��
�I.�Ȣf�0��{{WXI��!M�1
%!���΅}���b�Ȯ�^)q�i.���3�ݪ�;�mC~�~=I���wm-�3.��䈭��w�N���ɻd�'m0ٝ���KO�i�����6+{pOLJ���7��]t�"��� @� �W������s�����}�఺�.�������E��1:})B��^�:���8a�t�i� �0�F����N	��K,7'=}������2�¾�xB�'2~K�}�,��n�3�*������S�W�Gc9�!�%攻d%Q�s��6�=�	��t�+${L�r�s�W@.�ve{�Rkk�Z�/��Un_�MNt�@¿[�3��j���sΥ���p�&%tSC�I*q�q
��X]B@��
�.7b��������%���o�|6k��|�lG�+���&X��)�f6�#�[��D̝��A<K�;��a���U.|������l���u��K�`ac��l�ɋI����{]4��G�`3�ͱĝ�rfx�T��aS6�</��VI�+Ix�k<*�½���G�0�֟X[�`���ˉ��K�@������ߍB�$���I�m�v��R})��x����T������3y�� �T�����e*4�b$��34� ��ΟY߁w������oCRfi8��^
?�=�ā�CG
<�gd�����Uљ���Ǭ���`��=hv��ƶ���mv�76�i$�LW�X��?��	��)��v��J==7@���������^��؍?�(�4��E5�{0����o�m5�Q�I� n�я����l�3�u�9��"N�J�TZ7J�G4��k�9U|�
�H��b��
��aM_CY�L,�^��Υr�	�I�/Zɮ�N���Z|](��|��4uRkj�Ա��u������������H���m���QbG����qf�#�eO�u	H��kg-��^�Ĵ���C;cD���o9Sѭ+P�g��?�b؄�A}��-�8ɒ[�	�c�-#y�Z%�t$�~]�%,0��Y�dl����(�fG���0v�K�yX16?��7^AC��R�E�C��=L,����ܺ!���F�Og���TQ�8#��ǃ[Tʈ�e��<ן`0������ܲ�y�qry&�
HB����iį��*�U�L��'�����(+����6�81�*;BE�j���Nfg��I˻c�t�rc��9E7��;�;Qz|>~9��n�x!�szNXp���vX�$�l�o�4��9��9�U̺'ӣ��	l��:j�/�"j�f�[�Y>��QE��K5��x��1JϷ����	����n�ͺ�X��)�M�B,)\P{'�M�H�Yf�B�`�y�I�?�������V�J�t��͠�>���Mj���8}Z�Մ�d8��s�5�RqŖ���>\y�z9���QA�X�ֱ�}��;$%Z"��գǓ���k~��ޮ�E͡��3/�r�@�t�)��B""@A1jB��6 �1J��[$��2��?'��)���5��r�	 �&�����#������fA�Oi=�v�=-�1V/��W{F}��O,�ڍ��ֶ�8L7gt�����!��ףjE��|Op��4�{*�2��!��|*:\�I���*��i����"�1��'Y���Z8o����}�T%"A\K����z�tWͅb.$ۤ�Z�>M#��S1��Æ�yDt���3��`X�e䈱+�G0�]3J���ڕHyyoJb5Cv�waxIQ�\�d�����mIbB�oR/,�j������(�pU8�����Mڱ��u�0"g�v�xb_���2_�c���l'��q�馐7r��X�U��"��'�i���jL&�����]]��[��e��^�eeW������Ǖ?�(w%�[��Vh�݃��"���T�B�Иk9:�l0Z^d<�
&�������6N��AO8�*V��{��ds�M�Q��B5���V�V}��S�Vޘ�d��i�Yk��gE2�V�
�9e����x����lL>0)~�0�*�'u(s���j�}�A�ᨑ���y<�mη�F�1U�^Wo"�< J0)*b#e~�]�}����E����[OR�e�/'���f�-ƴT0�j�3��~(�����n�Wy��0�Bx*C�j�d����X�
q.����)L��?z�������o0�צЪ:U���JQ,B�N��_�B��I�^AόRm�92/f��s5��Ux��N�#G=삵�Ր1M�xY�/"t��6巚��v�R�tlcf����FATZ��B�R+=j(�}���G��റ�H�u:�-zY
�,=T���l7���]��a����86Nլ�x�I䔹�y�lm�0�*r�N~�z��~<9�N�����QʯBA��͓G��������n��W<J{�����|��Cʉ^�tn&W����6�3h;�E@K��ͱj=/X�,�Pԣ=�O9��E.�-^֝�W��F��|!�ub�����Ƕ�]�U��nN$���c���ZD��a!�M' ���t�R�F�8��МwP#��Z3�� �[+����H��nE����w��3Q�ͫ�+,R[%$���X:+"Z�� ��d˓2�Z��3���,��
����4=Vя������K��oU#M�u���=$!�2��SZ����l'I��/�U�P� \�h�����[|��e7�lۊ�c���B�*��j�n