��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�U�6��v�����(@�da��Ku�������bF�\ou�e-p9t.�e0��z�>v��V��;>��0TǠu��{!e�3�=MR#E-��l�l̼9��T/��y\_살��p���ՄL�B;�⸩>����
'��VY�쏚n�i��{|�C��@|Ύ� qTH`����ԕ*��%OF�tbp_�@	R����ny`//\��у�%��ǋ�䏙�UFG�v��!��GD/�K�t�H���fT;�q�Cx��ޢo�t�$�`S1L�j�V#�Wiv�?�4�Hð�dʌ������;���ꌨt������G�ڳa���	��?�D_���=Q��J�6���.�W����[�	��z�(%ѱ�a��5d�Bſ��Ǳ E��R�З�&l����TȌ���l��bÊ�6�`��x(b���)'�νV��i���_��l&햜�4�����F�&���E��u���N����_aY4ˉ��@�+��=�M��iSY����T�֍�W#���ON"�S�Zz��US�d+z��æ��*f�2P��Ur� ����������	\�o~s��jB�.gM�1R� B�#�����<AϞ�,:T(�JmVd&%\Bd�<��pc��O<	.��(z���&�A�Xoefp����ޢ��9�D���<�L��ʷxV�tR��q��Y,����B^�k�b�fH�'���=�G��\��5H��m%���>�R�D�j,~;�ƙ
�J�Q teb#Ρ�piT/�j��:o���\����R�n� ��}��|x@�{`G�_��*�n�[Ց�Z�a�(��ӡ�Ҝ���s��y�9YcCj�jnT<�CH�X�����<'�t)<aO�(�H֓fa#������,q�Y���`�i^zgx��X�5u��m^�˧�2(/2-����{ܦ⬕�'���le�0&.5��$�4hY�c&&2�ձ�& �za���h�y�?���L���=$|y_Ww�F���b'�� � $��~ݓ�ߝ�ؼp�����0i/ˣU3)=.a�)���]���5�8j�RiA�r�u	�j���� ����r���d�h�\/��.g�3SO[��c1�AG�xA?�l2o&N��WR�%KS�>\���{��C�s�X�ё%�y:9�hx�g��|���כ��A5�0�jo1���Tˣi�A���i�{��u��
Nr$^��L&����"�jG�膃��X�$����,����j�|�7��ms(s��#\rcc�L.��J�$
��䝵sa&�M��1���l�s��Zü辸���F�ϑvJ5�M]��x�~@�I&�C���j+�1U��@�o�i4���Ȩ����ȧgR���Lȋ�?�,�I�/O~Ñ�h�[����Y�4��"�+�w1ba����q�d�t�(l!��1k�:,Z����C��d�%ד�&E&��N�l��_�ie.$�lKە��8�l��E����J��I5G ��M�̻��qS���b�9�z�b9�%�,�8�œ���/�&PF�`3>%U��tI߹������]��o���Ĭc�-Cs0�.�?���2���[�Q�}�%/3�v�Ό����<\��?�WՆ-s�?D�t=���1v�}�� ݨ|MH���� RO
�Pl�0j�"RN��.7j-O��)����0�̳��;5�9�7�{���r�*�O����	x2���c7�y�bS}߿�E�<��v����;/5w��n��V�｀<�r3�����0!���I��=-�ڢ��>�<)��8�oI�� �w+�,'�m� ��0�̠d��� �>�[��r:��o���{ɿ=5�JZ����¤'%����z�/@��:�;:$��~�z�Ra�KG���4�#�*����v�5��dL���a�d��q�op�Y��4�#�Sx��K�s]^X{
ga�t0^�߆����n�!�����!���s�]ࡘ^�L'�9��v{�?&)��SF��y�Yl34dU�r.�ʙc�Յ��$�"��ڭ����P�h:���7Y�Zo���������[V�:�U߰��Ʈ���D:��lg�"�!�vO��k��k��a�!{fl��L�U�,osQvrU"yH���.U�ls��.C-'��%�r@M6X�dT?��$�npo�je�<��	R�,Sf*6���3����~! ;���fA�u����&{�Dcl�Q�TY�>x�V��n*�p:�����rC!�0}�\n����7@�W��K�|	xb3�O=nRv{�v��mO$&*�F:`��V;�{R]���ЀB�0��V?zEr�
�,QOlT�f�� 5����<���zŎ�?���+[�!���7_�%�%o[�U�qR�A蕩��A�G��QOu�2K��uC2$/�xq����_{Mb��6�=Խ��	�6Lju&�N���=` Z�m�_�3��=l��	�.�3���vW� �N��2��#�^�r���2�[�f�	�r�I��}#�)���w ���!�9��A�7�Az��0���^Լ��8��9YĖ#X`;˔RI\�Ml�sBg8Һ�V�-ͮ#-҄���0@�m5�[���X
,��tb���7�F'���G�[d��ltR^���ƺ��Kf�R-2��P|0%�LN]��KV͑�>�,y]z�j���R�!$��Ko�k��(�g�Q��d�)H�K�s��|:ч���q�cŧi���h�J�{`��tI:d����ءT��P���|[�w�i�Y+� #�&͜��)�0���zt_DH�)�#㆓x�1�˰�^4�A�����!���^l��Qe��P�@�����1_����4���A��m�]Wz�{�t�O���q's:�fb@ߛAPNL����V�+Ό���qX<��Vk/S�+9AZ֮���A�-V��@��}us2!�	���|��}5o�'��ԋ����j���7+�Q�l�=���'{�*�?�0��NmY�R�G�$�O��&�K����bo���	�a���L�8z��\O��lr��:�X�c��n�5N��o����OY��c/*#.���#��kD � F�"h5E1A������P�7������:��
��e����r7_������j6�9�����}_�����?�h��+���W��)ڋe��̬Gx�S�ͤ�f90.�P�XKH�ǂT6�KTT��Ɛ�����%3�]�q����-�ݐ�VRf[�8�.��y�������zb}/��*bX���L�e}:�JZ� I4~��������|�*�P�G@��ĥ+���ˍ挷�����z܇&C��s]n��=b�?���]1��4ȗ��`l[ْ' G"9��Xޯ���R���r��Us1h6��\��So�2�ձ0�|��Q�h��C{fB���j6cߤ2��Gc�SkbqP`�C3�����A5\�P�Iߧ�a��8]�����$QN\����Nk���q�,��<�Ƕ��ЁR�rZgǓ9��T�s0���(�e#H����-�nl��������^��F�ATU�����li�>�|�쉃�)�M��,�eF_�yUc�E�e	o$���'�U�WFa>|�c�F�������■k-���`�k��׆`����R��؝mCq�uu{
�B �x��2�f�B;�n"��X��<�����-̵���%rˉ{�Ad�<�	�%~L��vl,.�:���Z=�4y�$U8�F���4�x�y���7h�5�Ó7I����Vb��Zb�ɏ).��U�� ����D��� ����L���zf��֝
�Zld2����-���5�XP����w���Mn3S�N�K��d��Ɩ9�,���Zt�V������l,��wَ��X��Ҍ���pp����.�V/ lEx%!D�t��A���H0ꖰ��hu��Ԓԑ��1�p���O����[�P�{{�����\/��it6Dq�����
� ��a���c ";l�>�2$�*��ӊ�� m7�Ag%�:1�?{b��e�����H��� �D���ix�:/�Q�W�:�Ր�&Z�ʕ�\Lm�I��i1��t�d5U߱��X�OK�2	�s�&8����vT�z�}E�P>/4��%m�l[H"a�E�����S��i���e.,���"/�y��� /��3	2��]�j�+�ln8R%�g��B�OV�
�Ƈ��=佱է.��ƀ��eI�Ս�ýC�#rگ!+�N"ӷT�s3��Q�R���<#/+;嵱�f�Ϩ4���)�|h�Qg^x�T�Θ�-aܚmR�Y!N��VOd����(��/�����	OW�P'�֜�a��y�|��c,���;�n��؏��4}��}�%�	0�E�$L;6���V����Q�v�ד������&�:�%Aؼ�!�.�{�-�~;���=\�xI
�b�+��+�MV�'�~Y6�����
"�ܚ���eUd���/2>�s�x�_g0\_�r�`,*���cۖ�V�jv�_�hƒ���W�V��W	6$]��=�?�/}�1�4�|��!mwrMX8�it}��*���<��e��!L��󏱭q#8	�,�گA���yS��ݕ|��չX���Ķ�o"3�5y)��jK�e� &x��\цfzE\iV�H��� �-h��oW^R�q����L� �Y'*U�0�]�A�Ug�	�e�/%�0d�h]��zO��1���C-	��LȜ��/� 4;�T���F4W�pF�^;��/ۖ �`+�A�e���X�A��u
����^�v0�D�{UƳ��6���շ~?x ��;څF���� -g�.cq=/�n/'l �e�:�<�T�	���5�3��m���F8���B�^u�y�߇��d���ځ���rQ� lrA�I_�=ky$$�2�vY��-w��d����Y]�4�u4,�6'f���PjQ��aQL��=멉*0O��)(�C4��s��+v3�U��>v6 �i��62�/�ٚ����(ndp�dp'�()D@����&�Ƙ��'7��{��uɅ�������	���W���7"
�K��{3=��t�F�ܬ�~V����X�L��kt����LP.�Ұ*�$^f@\5t��C���H�u�9}9�ԟ1~긠�P��Y��U���U��يO[sʤ{�]�G�bwH�����۞$b�<��.?jX���WA+Bc��wnQCF���6�`�#�,���돴��d��� Nj'��S� �sc��B��J�8�"o�
I&nx���i������v<�{0w�B�I��+���\�c���H���ef|PG���!��o�qN�Gy{�OU��?�PON��| ii�����S�L�@�\��i��ۻ9E(^hk
@�RR���2��`s��>��Q�3MJ/%#w�/�$�1�M�ۅ)�)��� �3 �)���]~w��5�o��?��+���V�i�����_�L���N��(T��6�"�" MmX�zO�+�X��7N�O�����&N$�h�r����'�k��h�\�`�%k)LG���ﺿ(^��}o=XV������6�x�	sL�
)�g>zReR��a����*3{0�k�_�X�v�T������:�}���V��(�3��oe���<�"\F��+}�	A��u|Є��*���#ǙB�$h�O�W91�+n���D>��=�2�g�G�0�nT�_xX��a���b�-4N���=r��6�P��}�ϸ��J1&Y��(茪�Y,����,� ��(;q�3��?�t.W�Pd*�K��XM�/:xk�zGht��8ZK��&��m��Ƭ74@S
o*�i.�ֆJ2�*�P�94pOlU��(.
|%��r����N�l�g7������;�L']י�X$���0�o��,���T)�q.#���SvitW��a2`���OИ;㯱"iP9��&HK-��5x��F��E�=��bכ��
�����A|;=n����e4�FN����f�B�}�zWC=��xϢ�Hʚ�ج�M�SV������z9d�n�Î)h���p�&Ⱥ��Ǳ�)�U�6��Dy���7E�5`���
��Wq��,�����9�w?�M݊@ۤU�ZK�´Ƈz���/�bwH.�rƓb�s3�Ku�=Q+P<�m��9i6|��lh�w�=���*Y݌�q-�7��c�4��)H��tPlt��bCg����s�`��xU����j�mWxY'���s��?��\����I�v�\k��5�����1���<l�����Q(���k=3��S��d��L\k[a5TR��4��N���fHVa�J�ED�/hƷ����
OB����l<ɕ�;[4�a��m`8 |��,�6H��ܼ�QbPuSK�8��R^�ƭ	�h\'ߌ�rC��X ��	�Cjᴎ���6�.y�"�ǘ�H���sq͗^��������f�7��P��lh?wY�{��*�aס�ϑ��;��v��%~W��sh�ִ]�5���⸮�L�l`P w�T�Y
s����X��if=��i���� �y��l �/p�-�M%\h�
�['�:�J�ʍ��DOl]�u_��`2��Z%����*k��R��:�a�N�rp!B��ό��*�@�Ha�9��H�Cˁ���&�ew�5��5�oz������".1�a�"�����}e.Z��2�t�篳�N	GQ2�,�����w�w顆�7*V$?�;8��_	���N��~g����ծ��va����m�}��Ӛ���F:�j�^΁�Zi�׎��g�0?��ƇR]~�ϊU�+��JB�;�2���!��\�u�1�U�|ع��6�r���[VC���j�&�X�b�B�.B�y�ΘNxoCK�lA�?���
�\��p�ؾ���%��h'b��Z�\,�c��B���r(���U܇n����<�)��-�zq�׾ x��8��&
5��t��2�d���?`+A�-U�O}��Cֻ�P���0���$�����=@oVU��Kv��Ph��8�`��ehX��$�UZyX0�t������K~9�gy��j�_�bW)!�Z�Ʃ5�I�;�nեj&rl��|K�u�f'�z���b#�~)~A�R����R�@��Z,�B����OU�Կ���Ɩ�[<��v��UD�Z��%o�C9��g����J�g���}�U��r��P��pqimC�P9�:4OWN��؋���F���K���^X����	�i����T�֑0��r��s�}T�_�B��v#[�$������%��8�uk��e`w:�@���xN��8Q�m�Kx�$��0��u��e�ʋ_b� {��z�ֺa��dm�Rp)��J{$ �<!;�zu�O��t�����)=��A��ܝ�=:0�.�=�~��+P몲@���|(,�]���%��{F�thd�&�z�XZ�a1� x��w�NG��n�K���A��:��ѮY���X��C$�����20��<�5�5�0��XIl�!xO��[�b�4�i!�_��l� �0����Y�����_�þٍ8����j�9��Vl�l.���diS�V��#tg��m�������s����6���	v
ğ(�����d��-:ҵ�țe��O���ۛ�T�Ѿ��
ͥ�ro�Y`�F��	qbY�n�v�j1u�/�B��
�b��&ōΖ�����'����D8skՁ,=�����$�����S��x����;�:3 X-s�N�ǌm����wz9X1���h<
��-c�oY�~�N8q�O�Qp�%��^^�YX�%[��l�D�Ȑ5� �u�8���Y6�;nf�R41@8�xΖ虍���B�!�<s�E�0I{�"A<�pL�>nV\>td:G	�Bv�m�8��0�΢�1��%����=�?U����.E�r7 �]l?&��VR����fu�Y�L�Ug�
�$N�v.�	C�;�3F�P���xf��
{��#mB3�G�h��G�c�C��E��fqSe����!m�!w����(��p85n�����:�i,���H���V%ˈڲ�*�