// reco_4ln.v

// Generated using ACDS version 14.0 200 at 2014.11.13.10:18:27

`timescale 1 ps / 1 ps
module reco_4ln (
		output wire         reconfig_busy,             //   reconfig_busy.reconfig_busy
		output wire         tx_cal_busy,               //     tx_cal_busy.tx_cal_busy
		output wire         rx_cal_busy,               //     rx_cal_busy.tx_cal_busy
		input  wire         mgmt_clk_clk,              //    mgmt_clk_clk.clk
		input  wire         mgmt_rst_reset,            //  mgmt_rst_reset.reset
		input  wire [6:0]   reconfig_mgmt_address,     //   reconfig_mgmt.address
		input  wire         reconfig_mgmt_read,        //                .read
		output wire [31:0]  reconfig_mgmt_readdata,    //                .readdata
		output wire         reconfig_mgmt_waitrequest, //                .waitrequest
		input  wire         reconfig_mgmt_write,       //                .write
		input  wire [31:0]  reconfig_mgmt_writedata,   //                .writedata
		output wire [349:0] ch0_4_to_xcvr,             //   ch0_4_to_xcvr.reconfig_to_xcvr
		input  wire [229:0] ch0_4_from_xcvr,           // ch0_4_from_xcvr.reconfig_from_xcvr
		output wire [349:0] ch5_9_to_xcvr,             //   ch5_9_to_xcvr.reconfig_to_xcvr
		input  wire [229:0] ch5_9_from_xcvr            // ch5_9_from_xcvr.reconfig_from_xcvr
	);

	wire  [699:0] reco_4ln_inst_reconfig_to_xcvr; // port fragment

	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (10),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (1),
		.enable_adce                   (0),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) reco_4ln_inst (
		.reconfig_busy             (reconfig_busy),                                   //   reconfig_busy.reconfig_busy
		.tx_cal_busy               (tx_cal_busy),                                     //     tx_cal_busy.tx_cal_busy
		.rx_cal_busy               (rx_cal_busy),                                     //     rx_cal_busy.tx_cal_busy
		.mgmt_clk_clk              (mgmt_clk_clk),                                    //    mgmt_clk_clk.clk
		.mgmt_rst_reset            (mgmt_rst_reset),                                  //  mgmt_rst_reset.reset
		.reconfig_mgmt_address     (reconfig_mgmt_address),                           //   reconfig_mgmt.address
		.reconfig_mgmt_read        (reconfig_mgmt_read),                              //                .read
		.reconfig_mgmt_readdata    (reconfig_mgmt_readdata),                          //                .readdata
		.reconfig_mgmt_waitrequest (reconfig_mgmt_waitrequest),                       //                .waitrequest
		.reconfig_mgmt_write       (reconfig_mgmt_write),                             //                .write
		.reconfig_mgmt_writedata   (reconfig_mgmt_writedata),                         //                .writedata
		.reconfig_to_xcvr          (reco_4ln_inst_reconfig_to_xcvr),                  //   ch0_4_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        ({ch5_9_from_xcvr[229:0],ch0_4_from_xcvr[229:0]}), // ch0_4_from_xcvr.reconfig_from_xcvr
		.cal_busy_in               (1'b0),                                            //     (terminated)
		.reconfig_mif_address      (),                                                //     (terminated)
		.reconfig_mif_read         (),                                                //     (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                            //     (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                             //     (terminated)
	);

	assign ch0_4_to_xcvr = { reco_4ln_inst_reconfig_to_xcvr[349:0] };

	assign ch5_9_to_xcvr = { reco_4ln_inst_reconfig_to_xcvr[699:350] };

endmodule
