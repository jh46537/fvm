��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C���P~�û��2�pn*��J@?�f�f�(�V~�Ts!h���P��(���hP���%+ÿ���j��`�O��V�4%���z�4�rC��Dk��;��HsJ�6�txVO�A�1��2�R��\��,�d�Bm�>4 N��q; IvDVKl�+\8(�e�u�����.nך�
�ZV٨��A
.[�'�Z�dg���r�;�b&/k#eo���;ssTeot���O:�U���O����s��8�c�v�Â"��6��`�ڪ�I瓮�=D�H�y6�e�P�&�#��E��5������2G	06I���,�L�Q�P�LwػY�i���Įٔ����:W�^�f6ф�ߩ4�dZ�d��F��jy91=�É��eا[�Þ9�*��:ʅ~ŧ���k�Z�=����E��#k
�Ҡ���X#�
}5^�J�9��b�N��?㲅6]����J���~�9z�u/��֎u�z�P�CK�`!�����><�𲷨����:
�S�J��z��)�d|��ך��{��|��`��fm��m4�����(}}#���)ծB�s}��C�%��s�!!�$s[	}z�o���M�Î�Md-�ޑjZTNOLyA�?T�{����_����C!D�w�@�OYC�S����t!��lh�����2��^~E�B���]w���M��ܸ�x���a����O�[o_�.͘r�����p�s�>���ǣ)R!r��������O���$�� O}�V(h�J��ZT����Gf�h�ڪ�\V�HsGls2(o��fV7�Io
 *Dو�Ӝ:�p:�1��)��W�tk؀���im8�����
�5��;�3H�[���by;���-V8x$B��V�N)�u�b�E
�2'22J9`6)c [�jj"�E�Wt0��.���G��aI�G��V8�����鈥�׼R��j�!ɭw<W�J4��b�f�F;t3��gmll�lP�Nw�'e�.D��*FgQ*�C����o��� �%(��>�X͹��l>�}�i��1�J��}�஢�-`�Cq�s)}賧��Q������!^)��53�$D��|o�N��=�K�f��d�7��du�H<	�lsH�`� �=��%�y1��n��
�/ĝP͓�
����8~e�,9����?�,.4/M�� �D�41�k� O�H���-�j��ZI3�l17���٭���k�륙���6B���W����GX��*�U~K�[��[,���gP'��$���s�aLԸ�����{qm���������^�;qr-�� �Hu�=��u@�@$̮�5v�'-	�e��_q�{I��]����^x#�۫��� ����pk6#5�kX�xɄn���˃�΂0�?mB����O$j����I����S|�Z���-�o�*�!ފI��j@��gо��Fn_�ݓ� �����.=)�u%���o�\���)R@N>�������*}�8�r<�{�<��v�r��UtL�s�����PC_R8��(��xa�'Qn��s�����c;����2M�������ha��N'�ĺ�o��T��*�z{3ngX}`����X�����|v9�Iw5)�[S�� ���R����������ĒK��?