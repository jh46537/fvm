��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,��&VSA����U�i'� 5ևYg~�D-93ۈ�&ߺ��u7�Z�;^�\�¸w��h g~��
ܜ��æ�A��6�O��S��=F���lO��L�Vp�����?G��;�O݁�H�9�mm�a2يdO^p߬�GNc�������Aج�Al�1*$lS]Q�Xƞ\�?��r��Ɋ��g.�x�E��5~���Aa�_:�� �������m�)c�N0(�KHO�B)o����qPW�0�L�AT��1��$���*"��T<���I����/fyU�|��C|�����Q5I���U�^ �g�����/����gd�W`|�faZ.��z50��x����N�k�*��QϏ��vb��1�MĊl�A6���hOa�Ô�H��ā+RTR�V�t��
��x�S)�����{�t����L,FA��+(w�q���*Rߝ;{z��onq�:9�-�gll�*���w��]-{�	(�3����SVl;��"��0n�G�n��ƕ"S�F����2tK d�M
fϙg��+R��$��6�� =l�\>��Տ˦�]_UoY�+���Xl
�J�`��_z�N$�$f�S�e-X����3�T;}�^ �~h�Nx���ͷ��%AUVc����
�K�-���7~�@��Az�e��s�a�G��?��ٺ�AFC�M�Q�>�YA�o5=ɴ��vp$��8֦�n��#N�0X����?Vk|HU5�W�M��]]����	�%~\��(IHڨ�m"5�%�:��y~�YK��o����p�ōp"bP��)��ð�2C���0�)X�y�%�՛E�|*0��;��s)g����u8v��������.�=���}�ǰ��'U�i����v��x�82���+.M����U��?��3�Ck��p�Ō������+	� c\Hå,A�j�Ep�D�%tF&��W�L�U� �f�s�M��#q�:�o�2�<3L��$l����<Ū��t�������x4K�I���]�X�1�/�I�b��R��~���C������@���D��5�jS�=��ę
|Z�}�l���wh� l<u׬�r�5���*%IL�rA^hy@5)��L#�q:��09��L��@�_���1�̚C^Ö
�U5Ҿ�O�) �C6H;�\3�y�<���b����Ǫ�l �7�ʟ*:��h(y�Y���87�����j�q�jTl���a�D�a�e7)o��4E�������� T�������X��t�/Gg(5�7˖�[Z��_���M�6����U�(`P�4#��F�XC�iB��ri�Y5�	�LȒ. Q$�t�Ie�e�l;X$�>�� X�zB��W�ϙ9S��&�h��ȑН�4�؍��K�6�^�u>8����'�NVV;Gp/��=�,Y>�ŏg�dV�N�h*!t}~�&'�#=�,�{b{���S��!e&a,�w�F�(�d�#HRs�l��t㞎K})`��p�)�(d-ϸ�t���DS���[��F#�[�Ѩ���ڭ[���9ŵT�#��EkK  �`8�Y/�jj��tx�m���ޤ��i���B���8���V/��B]6X�{&Ι�隟v��(�]M�iNPk��{�Ϙ�?��~ ��1�H�E5�ЈV��3"������L�e��Ab%&*E6�W�( #f�j@b����x��;`x�u�4OE5�����Kʃ
�CϨ
W�xy�s�r��p׊Ҋ�⼈�];�)�����(�)����Ok��:
F��SU�X���1/��p�: S�s�λ`U�P}J�)a�ykGR�]meNwD45]m���>b��<�� ��-��ܲ7�;$�U��Ҷ�n�~0����@lt�_X�m�m�������O�K�q�&}�H��5`�3�w��FѰ�:Ѵ���I�-n��X�ĭ�_���㯍9 f�7�p��S!���T��d-̌ˏ���k�j؈r��v��U^1�}�{Q��oP�T����������#�%�\E)㐑d��m�ayC�y4�8<"5��l����3�^���}��䲶��BKN�u���{8���5H����3@���GzFm�����w��aT���s-Y��Ҟ�-i;�W��w;�˥�A-�l#��e=ꖬ\����)������C_Rkc����K_����rp����Gq���r�����'�Αl���I��M"�G|�x/1����.x)b�^땴�$}���h�����^��U�L�UG������c̂=��R�	.}fɖ ��2��ʂ�CO��X4�ت�Q���P�`�=dXRv߿BōfD����P�ޅ4�?/���mg��r)�������KB���e�9���ʯC)?�V�
�"���������7^K�)"g�+BF�@�����+������.ؾC�X�K��a|S?�V�l�������y�qe�te���X$aJ��Eo� ��"�3�	ō@AJg���U|؊S�����Z�'fh�=�^�#h11P8�ف�M��K05��F'��ȉ�����i!x�|��ȝ�#�C3�lc]s{U ���9�4�H~���������k %m_�"dU.�<{�Ka�80� X�.�O� ��E�U�>�]��4):n-rY��S+6��
<<�/k��y�o$Z�c�U���Q��l����|�F�{]���!�O]	LP��,�t�