��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^�.GJ��-��?f�b��(��ҥ��Y�����!���نϊp��=׈�kS(�?D� Y�S���#��f�����V8?�_���Mg�\��gѵ����s=�B_M�E�B%z1�����U����\�����ZI^C'���d�_ ��-[b�DU�Vյ��*�0��/�^�]ݚ�Z���r �Ї-�l�h� n��ࣁLR�5���e��G\"�JZ�z�!���0�.f ^w ϴ� I�L�J�ȷP>���ө�,5�%%�bK���>�͇_|'xƈ�&8�.�7�ԯ[����!�X��fŷsIE�~O�l�d�O!*�W,��H�����;}"���9��k�CD`Y���r|��# 媑6�x��31�_y����ъMd����<y �߱o��)a˘Q7���{;L��:�:�6�w�K<�&W�u��wK�M���b�[���h��������HC�δ�;ի'�(�����Ӥ�@��$ �V]z	u���#���ځ��2G�#�B	�}x��G��߳~��Yi�y+�����(r��ꕛߥOy?���B���W�uuB�d@�Z�ܩv��x= �ap��X��(O�vNleJӣZy�D�o��/�?t ��0��犢�?�T�*0��Z��}N�YE�1`>�	r�D*�>���NqxVJd� S�3459��]n��H�Dﻅ"��7w�a�t^|�p�v�5U->���^� �}�c��@T2��)6V豓�"S����Uf9�g�$j��j����{?��S�X_�H�_\��ݞ�D��.V�H��BF©�;)B�6ƨ��J��>@&O���Ӯ��~:9����9�$ �H�J��s�W�i�S�����A��G�	6¶D��������g��HS��C��'�,6�Y�"!{u�|d������9�"�Hj\��*�Լ�����(��O���aZ�`R]�G+A�&��L<���>�K��(�	"|j��Y�,J�����r�~�Z�gC,��X� YD���L)�?�͏��Թ�_c�S��6����t����W�h/7�Օ�^o���qYX�-V���+M�4Z���^���-�(�[i>��Ͻ��X���~���2WC���}ğP~���DX�<'�&J�@3� �,ʉV�,��q�,7�Q���Pe)-�n�!J�(_�ʦ�F�E�������r~	Tq���#��RS�(d��kP��&��Z�6�<�kz��,��ۂ"4�򒄲#���J�za�������MCg�#��^���"������,��`bY��8Of���f�u��jP�@� R���>F&e:�7�<^�}��P���	��8��H��$�����$q4~S�'�"G��dJ���N�K�:Y\�L+��9�N�#�Q�� ��%����h�T��0\l�����zI��g��q� N�Qh��N��P��������@N������`}(�ox�'����f\)3�����A�UY���ڋʃ���z�;6�V��Cӵ��g��f����XD�;= �;��?U�#�(x���m[�jm�f��T=�o�F ]k.y}M0VD�cЖ4%�����]��08JA���Y:�B��lв���q�a�a���ДS��ɽ�X�&ӽb���!�y�����p_ޤE	���g��qC�KC]��.�Q�!W����]b�S�|��c�����k��툷��|%��:c��}��z<���Q3��Zx�XuCh��ՒT���9��~�>kމ9�%���(1��}Vt)J���[���J�#���h��8߆�]*�����
��6,h7�,��S��1ĥ@C�%��+`��2�H[�F�O�Ji�Ũc 4�Tg�rU�j_XM����<6�;�)b���6W��%�5V���m4������R�o*�fA�ϬT'���6+��_�/�
=DN�����gd9��Q��6붷�qU^�*+6�i1�1���3d��X۫MNWxmcB)+q�"�'.��bȺz����ޗ�{�d�\)H�<&���~����X^�h��1��C7�@�f��Z�n�)�$H�B� ����F���hg08t��Ť����"��|�QӋ=�	.ߺ)B�M�J����6���6��5V���sɅ\�~a��C@!����`�u�}��s�Y�<H9wb*Q�j�߰mD�T�v������à���~�()	�TEUtF��#�ʃb����K�6h��}��9����e9]���|ȑ�mo���3�iz�g�꡷!����h���[��A|�Z��S��o�]�#���.�)9P��ous�ݡ�:��ͭ���D��Uv�*�fK?Kj��'� T#�j��!J������d��HN�aPS�j�j������a���T�]��e�-��9�@�����3�{��o4�rΣh�����#���8��o�^�_���+$GK���?=Kj'GR�לC���FXA�0��S�X����ʶ[E�2�N\����`�x��9@�����;��|�S���Z��ѧ��8��V�z �ȯ���'��4Z�.[H�S�E �|@��'���(j����b�aEWۈ�e�;�,�n*�$֜�e�~4?6�S�Q���n�!�y�w���]v��Y�`^�Rp�J�xU���������g�~�	���
{)�&����S��e4V[�8��+$��;�����t�dD��p:	>��	��=0C�[Lq�j%u?m�k�=���5�( FR�>e:H��@XIjau<�s�_|�>��M������	�|�!�O�igD���h�.Tp�52��jG�R܁�'�6�V�(I�9�d�ѽ���-!uGO*�-z�sD�&E�w�s�^����� ��.
�����u+d�\,ARRE���όʋ����EQ����8�RUi�ᛤx��0��Oլ��
�Z	��jI���ǎ�x��1�Y�]z�5_.6h�XA��� =��z�e���1fs9Z�5�ȫ���uc��ce��9Q����e�` �j��8��䒹Q��ݵ�۸>������7|�=��Ў�p��iF��S���Hn��6�C���V��pn-�+æɁ%��ټ � z�,��]�Y��T��zSo	%� 4��WS~�h���*����l4�J��>��(�
��k��9��[�2)�.G/�W�0�`j�{5����pS����:{���h����O,�L��0�����Y>`��
ڋK�sD����3� 6�i��S�}A���ӟ�8\ /��+=1NM����ר|�*�9�I|�)����6����(��Zx�c?f��[����!O9/�^( �s�,՛U��<q������5͟��^�$cY�%e�[���t����Q"{��̓��1S��_.EI�&ɧ@U�m�bA���3#ʛUέ<������J{;y�۲x7Es/��G�;s�X)!�t�;�`�p>�Ú05�"���#��%�����F���i{P��`�y��Ƌl�*���뵧G[�E�eQo��id<[��XB��Ϝ��!�QK��R �H_�s�Ba�B�$�~P�a��#B�e;̑����;�B��f�s��#��gX����0(ԥ{zÊ�.�!��4'(α�@�Mw@�M�>�,�u��^X�*��m$K�-[���.���`f7�	�u�T���|���6ת[�<��αF��y�^�'R�x��;��|�t�*9�a�>�������J��Ղc����#�v��\D�zU#uq���+#�<1�Ve��ύ����a��9��	��"�0twA��K�rc�#R�5���,������J�0��w����Kw���D����D����u;���s������;�1��t(�H�̒�� �(���^�U�Á����`�L���ܮMZ5�vI7���[�֋~S!t�n���܏^�Q&��X�

�m�2t�4ͰMR
�GE��n;�p�%/V��bWB7ꥬ�П-�c��X���;S8���֬
}~��@JC`����E���Z�!���u8���n��Jj}��E�xV���N���0��I��#.|�_����5���f��?E�WC��JcF�x�fl��#.u���s�������t���ȡ���8o��r���Z��Y���%�a�*���=A�6�+C�cM\�k�oB�+G��	w9���X��H�eNBV�Xn<����i�Pd4�{EJ:ҍ�L2m-A3'�1�ڷ�����+���j�W���Y/K�=^�G�J7�f���,�J�^�X�֊�Օ8�EU�LC���r�R��J�M�=���v�>�@M|�w�N��B'���=�O���N�7� ���R��Ȯ�f�m�a�^�B�7��L��](ݨF�y~a7YƂ5�-V���������w�ߺ6�Zp���f͂���R�ץn�!H��}��^3&��I����ay^�}��.��x���̌ė����6Xd�@W�5%\��p�'��6�(���n`˩���GN����Ł+�H�z�hŁ�<}��S%�
� � � �H����N��^�-\ �0y��Zw��<8Db8��QW���k�6��
�a��o�׷ſ{���'��9]mm��. ���{�����ڥ-N�v�9�a.`��M}".��J�W��"y7v��,}*�2����	�_��u���Y4 \n/ZzӢacL�������s|x ��a�OUi�#��.����3�u �Ź���&S!Q���t�F�u3��;���O���ĉ�
�㬝�6{{{��n:"������!y(f��&�ހ������޷�L� �T�����s*�[��v߆�j?b�c�H�1��wX��~
�9�f7/3�A����������V��uČq�'����}��,!r�ϗ�2��.�r��6ׁ�� �ڷ��Y[x�I����x��]6:_O7UF���,&h_���/zOe���Ƹ����)Y��Eћ�L?Z����	ql�5�L3��q�Xj�2ܛ~� �㌔Z��Y	,������_�騻�A������5�1�!�D%8�N)C��V������&"��p�d܀��<�$q��Ru�!C3�����"ɏƬ�v�5?�4+u��d�#HvfY�&�ȮJ�G�<x�����%��%~�Ϧ�z(��*��&t���s��2�x��	��ɄR ��N��|�4Y/9��Ze`"1��%�B�+�łi����ZB�y���@��*�l$gT*[�"�T)b٣l�)�@����s�@咤Vn0�z�kp�)�6R���t~W�#����W2�疃�`�X�1 V6锑aK}��ms���,U�p6�c!��]��gxq��foN������ӄ��%�y���P{�y·���S�n�� ��[��7���Q����J;		@����0�u�Z7lfn
�O5�G�}����4���gD���V���֔us}�\����:� O߂@�E�P�7%���f��Quz�\J:G>.'��$H�Vo#<zG��]$Ʈ��_���GL�	��*]Jӯ@[���k1������AYR2Y�+���!�''WU�WT2���B�n�1��8������DgGƠ��g"�܂:ɼ8�ONwY!��N����j�6A��E}��;0nAK��.&rk�2b����8�vi��2�����I�T�x�� �痫bx	�`GW�P�ZN����a�0Pq��İ 0�\"S��9�'Hnt�+����d瞧�7�M�;�p�[W���v1D6�\� 㴪q��se��]�5�8\�KL=��\2$~��W�yQ?�����n�7�3��emg�-�C�����	�q�&�j�G��xz5��5FO�)�=���E�/���G���Tx�PNv��Ko�8�5w�݆�6W��PA�V�S%3n@F���.$`��8��