��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<����d3��i��:��@:$���;��U��zV>���=c��Pz�zް���5#L��I%C2!:	v��H�?kG�<��_����ǻJ�I�JiUK�Kfƶ"�&}Iƈ���[̭3����(������Rr��<F��0B� �r:[��	Ԑ�pA3�R���}(N��1*2����Es����bt*�x�5㗔���W�\I��?�C�$!q�`�����J�)PXf�z�9��D�����I7�l�~�J�R�4}/��|�oO�>1q��P���@��֝`�!�g���3n��h���4K��Erd2��I7��,u�(B��Wqu7�y�Q=3�:�q��ߏt�"9,��"��^���ಉĜ){!�╁�*���af���⣳�Sk��BDq�^4����]�"$���Y�*y��B+�j�Q��|�vϠ�1G|���dbl!����R]�	��q�m(sڋZl�l��Y�U\Y� ��ԛ�ޟ!��Ӆ�y86#y��[����wd:ĥ�C g�9Hv���>oJ����v�s�*�|��=d�6m5� �O��������E}�.�{$��>Q24�n�P?»�b,	&wYhY/��C��>t��,���/��D ��nQ���3zi���>+�ےϸIrHy�[��n-IG�Ϗ�^L5�8�3���Dh�R�����p��2l�,O]�8���5O�%]����L%8g�Vlex���ms�l�XZi�	�����R���mxXa�z�\"%��[�����F�nG��t�e��-"h�:�:ɯ���osYsl�8@�)�ZK}�ų��-"ݓ�ߑ�7��Nk\AC�w���O�*6+����A����cN�U=@�m�].���]�*^B�}A$׬ֶ����:�p�m<ݶ=3������]�����Ҭ��Pu�z1)\4�L�%t�Pk�pUжGa�D
	���p�ۢ��������&i_K98�F�����sdG��x����Ņ��9����qZ?W�����`���P_>�?"�vԗ����df��~H��_�C�N(���vs�tR��F/�W��6�s�J�:����H:�ӭZt=�JlZ��nO�nz@���R���R����z�$ī�KJ��yhf?�D�dm΄?���f���M���O�v\��CmP眻�LT��2T�z���X4&֦�;5؊�`ʯ.]��utlI��,\��%fήn��y.bX��13Iz��z��Gᰓ)��f�䩏T�3{�:�����:���yٍ,g�x_��#	�NSk>��D�9��f"����͓�;�ρ��s�xo��Q��W 3()�o+7ڗ/?e�%V[�F�%��m::HZ���Y�`� ^!!-)�(�6 G����$���r]ߩ}.�"]X���\5�������Gzn��`��/3�l��	Q4$]��M�_tk���v5��P�t6�"c��J���ZNՕ��y���>�g]����֋���.�_��1��u&��oč��*��V���@[�1[�Y�ݓ6E/Ϳ���p$�3�5{s4�[�v�rZ^��$����ƨ��ƫ�ws�x��~��ņ�m&�:������o��s�̍���>�P͚���DʿDj��m�:����2�iK}^�=�ǋa�ҶiX��qL���b8|�I=~|5��+M�c1�~��/x��?��i��=6	F]>�r�}줔o�����m�{�-���E�s�D�j�iڊ�ЦE᧯����3�x� 	�(W�jL��
n���Mn,<rk?��(^rD�'�5
U�ݲ��DƑ���(B�Pن�V���Q{0I�c��O���N�a�չ�כ'AV(RJ���x�=?�"NS���~���鷟�Յ�\��{��8k�8��~k����hŏ[	
z��;)6�E%,|~� �XB�'=NTL���ʽ}�s�5hw����b\�~,BƖ�*qC��^�U�O�N^>�5���%�Um�k�p�l7=��q��x�	��=l�D�.��� 9-hXCA]ܨvݟ��T��$;�����k��ȹð�le��Ud%�
a��Y�K�]X�1�Q��Xa���)5���/���>��8����@]��a��ٳ�X\Zَ惴ï�D�֓�EbK�(���3�&:�P����$��|G���ë�C����<�Pc��cˊlUon�̀��fV���S�G$9�� 쟯R&�{��=���D�<0�E��>Ԏ������Qwv7���S�K]H�W��%/��9��c�C<�z<Fk~�)�7FL�#%��?���G�	$+�o�bϓ���k6O.G��j�EV�m��Tu�#��ɡ����Щ��ti�Tע�,Y	ؤ#�����m1E�qP�ޡ�!�h+��y8 }{ �E���}��;}"&*��IwTZ�z�Y�Q��n�O��qu�@��qRi���w?]�CS8�7�����ʩ��})_�T��˹���6�x��U��cĢ)˅p8)�>��j/z�ߜ�ͥ��㓌zL���F��M�Q=�%ͺ]nəy��%��8_B��X%����_A%��?��7�=֥�f�]D��b�&��I�I;}�5��η���#�^��f�,F��X���Dd�ߺ5��|�(	�3m�VpMJ��|y1[�����å���?%�7�������L`%�H�X U+\<~�dk��Le
p��U�Ű}� 9v$-��ҵZ������K�#!�h<�,�7�\]��d,�?��YP�O��R9m�{	}_���)���(�[�r��&�)�{l�K~	��_*-��=C/g�l��dD_iZ��W�oS�@8��1�B�S���#������M�q`������2|T�<!�|���
\Ů)�.}�(	A0�����5O�߾/��V�d	�$�T"�k��������*���W��_��Y� ��_o�v�7}�l�Gu������=%KVW��E[�CzBTۚ�(k���;�o���n0�C�OqdΫ#}�	P�V��'5��S
��r� -�4p�E�lLn�~ң�Ϸ����olB���>�ŰM�k��Lj���p�����+����μ�!Y6P�
�[>���ǽ@�P�H;��5�Y���惠@(��bQ���?嬙ȻE��C t��m��������C'.D�-<��[�*��߇�?G���������$��'��6�?8D_��l�?� ����qkg
C	�R;L��¶��J�����p��Ŋ>��x�T� F��t$Q�W���\�x_�R�ᓕ��b�<���o���!�)�=¥�z�t�d�*WC�dx�p���Ƿ�72��<�]�B.,��W��D�iz�c��d�m��	y��p�=
8�Z���+�A#H�+��|^V�m4��7����݇/+�_FWzkJ�M�r����l(O󬧥p��������I#�Ӑ��a����ag��s&Ȧ�dV�2�(��t�dSع
x3e�S���a�8Pu0ݽc5p���)��6�i^�GE��"8� Ƽ�M�y�=oi�/�����E�G ������x�31���o��=�ނ��(��w�S����}%|L4+�(~aT�B���yT�dMk1�|4��Bl�h��j�],�M��$|�Bg��Q���i�2�����M�Q3���%A��lQ�Ջ+�a��������6}P�B��,�=Bǅ$Ϧ�Hc�3m TAEk��F�(t�u-ue�xH��L�(���m*<��-������ 1�n
��6��m@%H|ʟ�l5��4nN�y:
Χ��Dq��``oe�ճ���]����6>�|k��|�wv��G9�f^��1��8�Lc$�5�.N�靥�M㇁�ݵ�/5��m=��!�Ft��n�k��|��$�c���gW�/xs7�<� Z+�ɲ��$-�̣Ԏ���S������>�����zLä�!��{'���U_"�d����v�o��.'�A�0���������{��𥉉٭7�kI�j0 CN�G�v���Q��0�15w� �f�*G6=�¾��XN��{�s,��-@����\��)x��Z�:�< ^ =Ys��׈��CH:����
��~�Y�]� �o��6������܆'lWHu�ɢr#I�v�j�f�y�j|#���`����t<�~.��3�����y�����6�E�a�Ύ���lUa$A����V1��R�ݱ*���5����9d$�Ce�_��Q��%�g��G���7�NcJ�x�@���&���1_8��Wr�u�!����+>�~`�ܿ$�&F�~aB��܏6e�
z�J� ���7��B��/`̗�)b�������-^�7�O�d{Yq/n�<������'7*Ź���>U��Kd"��k��t���Z�$2s=Y��?�}�)���p��� k�^2)���f6�8�f�C�<��x���6L�݃Ӟ�v/�>S�iX�8�U�>3Ϙ��
��<���ܞ/?W�B�
D.T�ߩa�6�&W�(��r�Zzp�a]����9�l���^ꠞ�~6�t���3)�K��-�ElQ��~<Z���?����lh���3j\":[yI�������&�@��i���ީm%�9�!�x�5[�O��\��8�A���jK��^-�_�`�9�+�B��9M����P�x׋�����^��r�"e���N9�2ObF3�e��\&ψ7�B�����9����H���ׄ�m>�bUj���3�`��u���B��r�_O����Ǘ��8�1T�8����S��9#t;�^Wj$�uŋ�(�6E���i6<R~'Җ��z���o��.
)o���&˗�,��\�̞�[�K*R�@���v�d��օ}"\͏���l���S���>��V�?�0[8��" <O�0�*B���LW���z2��50�|��ɜ�t�턏�&�����g��4A0k�9S_1!S[W>.3lgQ�@��$���ǜ ��=��J^�iO)���d[a�LN�3��M��* 1��b0)�|�k�
���G
Mg>Mv���&H���%&�|�����́���9��|ʄ�οN
����S��捫~�U�aܷ�#�״�r�~���`NOi:$,�fK��vF�
��F`�c�	W�J��-�f�Hع-���]�'��k�`ԩ�S���}Y��P,�2/�ݘq����^����>�/�H	��	��)<J��/�y����8~+�����hj�&���w�]�4u�z�VSp$RP�-�ԓa��/�4J�zÛ��.t9d�Y��IK{�׵}
��f�e�9`�L��b��s�Z�VM^�gz���½)�@ﺢZfTI�	�����ަ�ϧ%�������e�_A�����/^ wK~H� �d'��t�V$�@��C\�{a?����Hɯbt�$��Y������w�M=0��zl޵ah�|s�J�!���a���Z���x�y-ypߎ�����ͨ�J����."g���Edjv�2}Ө���
��Rt�]�K�8����F�����O��.b�����>��q�&CpR�O8����
�Jq~6�]�A�i�$�z��1�{�(����TBZ^8�r�j�CZ����Mqu���?���,�y?z�iw���yjҏ�r}��7����ֹ�XS]�9����O��Ҳ��D��2s�+�S2���i��Tд�dG��2���O,����	���]�])�`=Q!'���GZAZRD�n1h�����~R��i(�cO�N8xHwzxBI�b�b!�]3ָ�{^U8j4�Egf���%��i�g��XPi���`�|{�ʲ��d3��Tm+����re�_�>��]���bz2:i}kZ�QK���fƓ9�S���Z�T���7BW�o���ߥ�]C���T_iM�A��"�����W����KW�i�	����l�w�����#����5\T�y��3��q(̊6�%%Bx W�&����������ڋ��='b�CT����Aךg�}�E��X�.s��C����{�i56~a�����z]<o��$�*Yo�-�kX��zV#n��tM#F|�.�n�n��y%n2lշ�c��jCn��ӕ܋}^j�7�6���A���h�{)�C��I��2�d�0�52+�zt *�S�})&��e'���5Z��`H���S7�;�tq�Y���ӋYυ�JJ����O�n�5�0��"�"���S{��)Ĳ�O_�+B��Bp�vP��⭀l
�9�I0�{��t=��"^�mQ�ވF��!���1	�9�����fhV𽣡�{J`�k(�A)��D	P�pT8���\}3�RFK��AJ�1W�񭵮X#q��p�`"&yU��%�Q���	rz��6���nݸ�S�����S렶����C����$M�v?�#�>I4�z�V�4�BB��D%�oOF|3.h��8Tҙ��`��0K����(S�́$H�H�)oR;|j�)r�?��yU���(Ւ?Ͼ4�C�n-����0�jB���E}�yc7;F����&�*�"�V��l_i��+>J�����.H!-�#�q��ޕ;�ٛ�-����c+V�*����@E%�#e�u�X;OeՌ� ��Ay2�WS�h"$� *}
��\I�;wC�����Ú��?O;6H���l�5"��>�͢CBC�*�o�*U��/S��i 
�|Gp�چt�!hD\�h˪1q/��X���3���<3����y\���?"����bm98�f�i��ۉkC��jD�!�:���+K�p-T�ۆ���� ]���5���P��+.al_�;4�yԤ3q����*�v��V�m��f<��4)�
s;�����V�Ϸ:��� c�d%����]!�������9����WC��U�;bZ)��������H��o��ȡ"�P�)�����t�q����e�7�}%W���lr}㪘԰��U;u�����ފ�Z`R|dr3?]���+���0�Sȥ���r���x����H��h��h~�_��_���� >�Jz	7���\r�
KU�<7��/~��R@yx���e���7�E�~v�k'T
[8�C������v�Mo����x`E��}`�24�%(�����e�2�x
Z����ݦ*�7��1�""�G�NϵGz���.�U>ܬ(��	�e5�}QS�n(	��.��N	�̯����k���['k�,"{�� �Y��I�J{O�tϥjH�L�k��I������E�W����X����K����㐱�x�sVj�H�YX*y���w�l�%{�����8�̨��TY�lZ]ժ.����:�l��=ؽ�q���x��a��/����yJK���3\V�QDٽ���|`VZ��3B"k�������RP^������j���L�ܢ�����;�F�[\ռ�Q0-+�W��rϵ0
��#̥��@�U��݃�v����ibN�Zi�gI`����4���'�~bKȰ�J��[7~�قp�ǖ/N3@"#G�r�핑��]�BB���d�%}�a�8䆛��~��O�ʂ����{��@lE��=���o�:��t,F}����{���<�V��ز�X�;��gt�Uuc�nn&� ��$k0�<��y�=�m�:��J�3h�N��L��O��2O�Q��k�E<�z�,,!�F�pR�5���{�<�(;��|UQō�Ʈ�h-�����3�J�u�k��)��E)3R��S�|I���rY�sT�E:���R��������lf�Yϧ��)ȍ�L�]�y���F²�|w`���FYϱ�[&���/4~HE�W��8"rO��FͿ��p{�z��9ĝr5����f�A��� M~`��?����&rP���{���Ǫ����� �@=���(��p��/SW54F�Sw�ϡ�Q=7�G	��Y�}�(��pt*Vߡ�2�7�Q(Jɠ��/u���Y�8�C�J"����Mc�+��+	�Qk�l�um�"3P���2?B��m�o�o�j͔�=�B?��#�.2M�$�3�
.�
��Pvğ>�To�7Ӯ�6	G����z����g"vJe[yAF�,\	<�e�:ikF�W��e���4E�=�?#��������v��AJ}F�!��Z4&S��X��:	����d�3��YH�g�W�v�=Ш��U�\�u�u�L�ޓ���YNx.ij��B��̈dˌ�[o���	�9�r��f�z�Ӭ/��� .c�^�����.١Eߥ0�c�r#���� K?Ȩ�щϱ�H�Ђ�2˨�Xp��8�ѮhM�f�A��
pܘ�#�*�U�$�p���&l�N����E%�<�pk.�w�g@�Tx������?������m�sԍ���1��X�*�=�x�N��狜Ɍl�M�Lz��-��P�۴]$U����"����$Q!���N�֯§c
\YDaA�e�ۤ]'ݣ�#��?��0c���I��˂!�d�+�#gy���n<:O�q���F�r��[�����0�7E1sC�l&*,���k�r?��O�tG-����WJ�K~$|Z�҃0~�)!d�sW�*1�O��C��9\V��Ҷ�1���;�{&���>�%QvR�\�;�u\����kt�J