��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S�VJ���ɾ GK�rA�!��}�x�E}ݨk�fի�u�(���L K߲w�.L}x1F2�#5H�:�'))�6_��\j�S��W��w�.㆔�[NQ�6��iM�@��9��eh��L�@�Fb�%FZ�"e��R���W��@�s3a�����膂Y�:�D���!G��j	�E����}��Ui����kh稯ka�"������e�^��6�ɠ�Ij��-���jW}e�@,��=��\�`�Ǩ��:>_2�)����������t*�� *��%/��X_0�2�KwS9�ڪaԟ�	�踷Q����Z�@Z|�歊�)���ܰ�K���"F�"�;�ŰS�d&>�،4j�o�9���xD��h[JH)���m�tS����\�ɑ� �n�{ƒ;PM�����>"s��R��m(ɠԉؔ�W��6���ߜ=�5�%�_��+*�o/�Wv/�nW�S������50�u#�����=�O�3b�w��Z,L+F=5�'�?y{��yN�2���D2�m� �p)*�CW��F�7�Ye�ȼW�xs	p���-0Gnނ���Q��	��q՜o
����D+�g��!!|VeG*�s�1� y��!��FXV/ao�
Z�#o �xE5�_�=��جƒ�K����#������\?xi`i(d����#���&S����$��a%�o5�H��}\�����?�ՒI�W��+|Vz/:�2�T�K���f?�k��A9���d�̺}���6���K�����T�ʫ�n?�塲������*}�Y�9�{��S���c�{ҩ����H���qn����qh��W�"�&sL'4Z����B��,8��w��BFd�8M�Y�b�oe�Wl� }�$�ՇD�O����r,���1�υ�\\v��<Ɗ��h�L]@�'�Z{�e5��w~��t�qJsP�X�q)��"ˀ�-׍����������@�(� ��bx������O�3�Ӓ[O[	�Q�����c���x������_��˸)��+��hNۚ�-�4�G�[��T ����r�͸���6�GY����G��E<Cn'C@>^=0�DFj_�hEň�
����6Yv��ݚ�n��r�'U�d/"�OS����<�N[�-��������O�oH�Xd�K�qF����mʞ淛�vKBDݽ��F*m��W0��iH*�SM�-s��a�fո�5/?�ز�yw����Ʊ�^3�T�%��ޮ�~�N'kK�u��M;�&8&������0a��B��{B�t����@ֺ?n~`š݀۱�
���
��ާ���2o��E1��*?�X ��1֐��g�0� Z�(ӖrA6��r|�5���"M��� �zrU�Y����A��-���Ӂ�Q����Z/*rl8g���1tFC�c���$	�����K�?������5w�"����xG��i�&�k}�k�*|}Ӣ�#K̉|u�_&�o@&.�
�\��w���ߌ��L�S[ {��3J��2���F�م��%���}~t�:���]�;�q.~��j�+i��L�_|D�s���Qa�!�_l����=->݅�����()�L��̾��94�ċ�2C4�N%�*J��&�+N�,'/0�^,a��]S����;�A�H�Ȍ�6ua�=����F��%T\�4���K�I�2Ӡ��R�D�-nt^4�P��y���ڹ,]�j� <;�f�I���\JY�Y�����Hu���RK�C��p�2k�a�M�Ǭ�uR c�H��(1����" >��[:�
�⬿�(���r<3Ku��K���{�/�6���w �z��݆�����-�u� R��o1O�[~�����?�b��)�9��L�	l�vh�/��?�g]be�*N���)N�W�ZK��x�)`�*R����6@ID`����vFګ7��*�^�ck��/�عx��Q�
>�]I}�b�&D%YD�E=�-������m�c"+�d�'i�,R[��a�p�O�2	6��c���~CÈd�BRAڬk���t]VKĕ[�ρ~o��������1��>�t����c��x�X,�F �h��������ő�s�֓ 
N/�m�y�VC�����B�������e��ѱ�nBx�P˿����H)�������p��W�Ϳw��"���4�Z���?��m���
Z�a�&5�=���Ԩw9�����j�����5mM�׻-�z��EN�C{>�@/�Gd�:%xə:�9,���̀C6t� K�Iγ�.�����d�LX]9B8T�R�����l�^��V�ӆ�i��4��g�s?AtH;?�Lw-U�yg���ủ��k�0� �"����<���o�dƗ�pBg��#��r�a(��ho���V,�b3�u@2dk��'<�t���GcV0�]��,��-������iY	u<��F���D(�𥛞ޏ9�H�ƚ!�H�}@�Ԏ%T%uǽ�=I�Z�P���VC�Z���?F�����*�h�6���T�x2�va�8� ��KRgi�W�L�*vN̚��gY�WU�
�|vq{����b���2
>�-��
:�!�%��o�է�1��k8�:�"����7���K�b~����$���IatiМ�w�9��H��G�iӼ:T��]�@VS��]	�Ԙ����\P�����VǮ|��R˞�����'�{{ӣk����sD����m(g\Ner'����kLhhΰJr�AO�J� n+���rIm��r��p�.ܛ�m�W�`���.�q,�&얡ڎ�u��UIQ�UR ��y��+�2��h�O��o�f��md_��s+�31�q��csB�����L���t�i����1�����'��yބ%�eI�%�Ό&u�K���9�oY,��Ir#���n#hh�̬(�S�"ƻ4�~5t{��^9|C9���T�ך����'�F�ekmŖw����������:��4!DP��l���9i<��乥o�!�h]�������N��,�Jέ	��l����;�M�g�z{�mY���}�� ~!���k�K�6��,)�?'�sn��G�p�jXݴ��t�8҈5..[�?͸;^�C��F�_B��b�E�����&�c��ηB:��l������=�j��u�s�I�q=\����mރQ�fr�1�5e�D�	L�xl�E|@��KM'9n�CiL�`FyN!Q�u����4�qhk�|�	e���f'9�\����x�l@qVWxsAq ��H\�����5�`��fl}r?v9��0LcSt����R����(af�[$�e���w�I�,=�1�aɮ\���t��¯��3
n��m�����3Fx��S$t?�� ���yt�y�6�,��^��bz�"����ṾGmo36�R�B�ڶ�2��_*KCޔ��<Yyi�/?q��aBob��R�D/�#�d�n�;��0���W֫lo;!{|o�N��m-
�= #�/��~2u����z�V����^4��7�+m�D�X[��QcH@yCO�Ք`�o������Ӫ���(�l@��Q�+��G4�E�-#$��j�=T�e@�����k(n�b��'�l��h�w������4���»���߽��S7z�%�5�z�9��E´�#�ow]g�^��xpLF,X�S̗���T���,�6�'�yv��")��#"S!��/��_I�f��(�?d�¾ ����LYijl\y�J�U���,���~������B��)º����*�?�Բ]&��#�`%�M�����Q�uW�~�qH��]7d$96�B6��W6c,�A�dq����s�lу�Ol�꾌E;�"�	����;��굴Vv�r�[� ���G0U1�e�D�.s"��+Oƣ!����͹?���� ם�[ԩ�5��C���fsBR�x ��_+�l��>���=�2k�Y2���1H_�/��=j���P�m�c$�VDȺ�¶�.b`˶}�e�:G�%����u]"��0=�g�ΐ/\��kܫ"�s;zz�n�Qڅ�e��Xys�l�\�t7�z�D�uC�q,�����K��3R��0�1g0��QlPQ�ldV�(��̓D\��,l���ʈ)�0�����c�i��'���>��h�'vj��9��.+��^�`��) lf�Cj��n.d�!]�_\nٯ��s�I��n�g���B���X��ဠ�6�A�Y��	��.w�4
�K4�q/�'�CM~�g���(�O_b3>RQ|��\���Tw�R�� ~��'TFc39�T0�8*�NN�[��	�!����I� �5:@�uN���ʤ2D�;KA�U�wۇ��$�6�s9

��n���X#3:�����L��nd�# ���&	��+`[�4�p*���)Fl�]�C�X}Όq�����e���b��Sp��ȓ[lp������&���ǌCl�'���6�Q�ip��a�Q>;72�O�^�4ăFSw@�t��B��<U;�Du	�tVl�tvWuT|ݓ�Y�>~�OGF$�Z�a#=eW�%��0Z�K=��)�D���+x%�{i<�97A���L�I9W�L?r�@�D�ۈ���� tvnp��c�8��ؾ�^�v�K�;e��(�% �~E*�;��;ia�E�1ǽ��i�Qi�@&݊��  o��{��$r�4�Yk
���k-�"y�7��/���z���F��g�`_��3��R�A/!vẁ�]	�7Gs�7�M�ΑI*@`�P��hl�u�_�#II����r=|מ�&^Ξ:.���/@�?>��8%ϓ���)�9U�"F(��1��I&���C�P�B��/Փ���և�M���9�)����
?�\b]����١5A���r���Y�w�������X�T�D���@u��$Tp'�����ic>Jf�^M������0'|F�:)UF�� �Yi���Y
�`������o�
嘆w�Ru����
Ej����y�]H*0]����
��۳JݞN�~tj��d�m�ܤi�M�I�˴
lqa|�Kv{"u@��n6ȭ��n���:�����+D�WPB��GDQRb��j����UW��V�L�oK�$�JǜD.gqD����L���T,���m�.[ є�i�ng�V���`�����.�F������Jt��Ӵ\�Ed�~M��+���%o�#�	�ϖ�k��*�~��K�0-G�� �0�6��v�L�{K>���,00.�,��s&�i9z��!��JYlx%�P�^�(3da$׸W�s��41y �te�:�U�T�&/�P*+��gD?��iN�2�R�z7K�i*��[s:
y���Q. �3�J�7��|�>�K�q[��>��Uf"
Gi�0Q��_)@+�f{��؂��0��h�Sh}Ey��,k���V1޴�����vR���Ɖ�i�'TJ~�CJb�aX�A{�m�~����J�c'S��>z.��8��<g��:�ΜPe�Eo�N��%��N�[��1!$��uF���n]r��`aȂ�H�٬ӝ�-�&�������Ę2�;�Z�5���i��r߅��AN���^����u@+�w�޼x�;�%��5����\���b.�����f4wN�_���	�T���*��MLr
M"��:X��D`�CJ�`�o�K���mb�+GE�sr�G���z�*���������c�*Nİ�aڵ��Q�I�s�~�G$��;0�%aW�{s��Ǜ�6[T�y?��s�3�^�ȼ�
{08!Xh�8�h��y���"���g }
�'�mѸW"����-K��(��XH��rF��j@��X<;�E�̐w���ZxV��i&rd�'V�ۍ�
ü���u �Ȳ=omk�J��~����,���c�Hq�<њ�Ut�n�6#�,���)��i�s�́S��Stk�Wm�m���/���i@��,�s�G{�+k���xa�Ů��V�PC@�{��2S/��C�^�[�C"��G�D7����[�q��ۖ�DC0BPnu8�0�ڱ�qt���&{�{o�l�;��Sj4����G���h�P�#p��v��']�ps��D�D����r�peVF�Hc��G��L�T3t�,[�ãX"yI����N�Xq����|Y��41�7��S�/����[��6�繇✪ �0�=�]���/�|���jŨ���x�_+�U���A-a�+�Έ�ӷ���R�O�Y���R�M�Y��ͯ��-g�2�|�ߦ��$�1A�?T�:O�@i���-�	;�:�\kS�nB@;�E_�@U3�DMt�`�88�P�]�C/�x V<���ni�[�Q��I�m�b`�I��$, 
�vZP�J`~:�[�t	���}U9E��(ٵ�>���C׫���'b��u��zhf�&Ԟg�������܌΋a��	��/�׸��[ׁ��P�%}��a��L(pÏ=�J��[�f5����K�o:K%�N�?��e>�,�3�Q��� �����'.B�*>�y4UI(G�|m�8���ZU���=F�P���:3��=`.U	0%�t��1���2d���>�D�α��ƾ��{k���P��#؊GDJ���D��'oK�S�ۣ���[a,d�+كǍ���[���$�B�������]�����$� �O��2sP9�;2rM�{LЗ�^�MR`(&g���t7�4(�����S�+s�y!�練/2������R��u.�������P؃$�9R�|QM���#�Nv�3�ɸ�qU4J�PN}[G|*�P������	�xk)�b��S ��p��]�9y�y��K/�����B5��V����`�]C�r����괭~����h>Ɖ�Lq�o�@.��y�P�C���n�qq�����P5�J2J2W���<\��ʇ�nj��g�����Ll��Z��(#>̾�u2�f��r+P�P�ԕ���@�K�U�ma�4hr��,�g�l>����LnbE�0��A�
c�Ī�
�|ӎ�� �O:��C	��Ex�W)�q�F�l�F�_��k�+ ��FN�R/�wIhp/5��.���� �@f��&�b�c���k��@��%��M5., �R[{����Pd�Q�e'��g�&�ᄥ����TE#�X��q5EƁؗ9���K_`|�hD���㧪�0�W�P��m���BO||��T8�V�_�M�-�X6US�(�ڥN�bY���.�W���Bz�L�����GFu�s�$V��$