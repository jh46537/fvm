��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��)Y� �1�c�{�C�9	��܈Y!����lJF/C$d,�V�<�.
Ւ�-!S�h��n����X��ѢS�R#`�ǗG�ݠE^�^HQ�JDbs��:��y��I����@�1��'�1�Б�4۔�K�s�~�Y.3�L���G��6���<\�.�
�m�܇��Q�o�j�>�o���L0��8_����M5ZN阮(貹��.+z�9�Y�]}"t�(&{?���s3�!�ii�ߎ�u�+��S�,�mI�=G�/I� -�Ez���xp�󴽏�i7s�[��9���?�i���m:eT�!��W�T�Ì%P�Y�M7?(�V��ē7�=�@	��$����ֽD�(S٤�����|>
LmC�r}��?]c���r%����D=�����h֎�	)C��k���ˑ�;�,E8��5�'��竣sC������O�X�Ur��W����q�N$�8�$I�a�J۶�J{�O�~�ϥ����AB������8�6-�]9�w��H�,��'c�b	m��F��A��6�r�i,�S�EPpJ��X�&0U�9*��;�B�k���Z<eD)�DH��Fj���h_��
�z�<�?/����_���
`qaw,���(��wh��k~��2���٤䧩c�3������]�F�b��Χ۪���r��L[�A��|��o���.����P�����,}��)��JL�����$js��J�@��W��φ9ÖQ�����	�\]h��J���F0bY�e�\{�)a-�������VNT�����A�Z��\.���/�P~
�$�5��J*�d��W�F߈��?j^8�:��Mj�%u	�!��z�Խm��_�ۧ)'u�)l�!l!<�Zc%!4]vO]����������-��5!!E�� Hq�Ҷ(z����^~8˹L]*w�F��u���TM��~	����!$z]���BDqDړ�I�ޒw�1����%R�%��5�|����� �bs�s���j{S�'�I{���=2Pl�*���S@���'9D[ja$��%����!\��o6m�"��m��K�7��嗻�z ��\��i\��!9��� n��~��T�;Z��8�������X����b� �3,���K�h��E��h�����o���dz䃭�&�̱�Gm�+N��ˬ�����݅��ì]5{�!6�O)�m�u��k��4o�Z�ŧ��<:�B����C�fQ\w�@�eı6�%i�d�oӘ��#A����`��WH���|�x ��
f'G�	�����*�!e$��}�TU�~����@�L:���m�^"��}��Aㅊ\���+&p�Z����t�!�P��Oh��q�71�Q����(����aۺA��ښ�k>ys!`��a����6f��_3�剶F��)7}>�˺�,Ad���-:Wqc��Aun���T3���᛾On�Ŀ�
�VD#ˊ�}e >���}p*��N�BSb� ����"ǚy�����S*ڮ���&-j�C��[[�}��y4�*�z�`LJ[�1�sQbϳ�l���=�U��J6e��#J!<w�SE����!�T�S 6�)ؠ����j�>�o�q�?�G��,� ^�cn?V#"Sx	I��H�G��\�ÊlB���,�3ȩ�Q#A�g�-��ᔋ�~!�Ko<�A~�R�F�,Er_����IjV�7�]��W��F�_J^޾WPqZZ�Dc�ɷ�sr�)���A)N�z�_k��Ȼ@ƿ~�r�S�T"�̛i����.�����,�>�
� v$��]��\��(��_��Mf�a�*Z�s����1��
;�pt����Nk�Y&P�x$X�U
k�Q�>Р�*_Q���5�s�"���6�E(�(J9{s�G���W����y�K?�����o:���c�צ�y-E�t�N[~\���p�a<v�UOMG�Op�[�1j��l��� D�B_������3����/�0��*N�%cc�'�PH���[<;2���5t��S��Έ�oaW[Dη����3�<(��m�eǭO{� ��2"Y�o��(ڻ�F�Ӡ����l�6��O���݆߇����!!�}ã�7q��2������� �}�V��s�Z*e��m��V�}�o��>2��a���>�dB���q�������.-��A�� V��IʴGk�A�g:Z��
���H��cB97��!��[)�]����ZH�9}�]����*�BcQȇR��$���C���$���!~���o����V�IP�]�(��Q�H�0�mf����BC�k_�n��Ń�,M]Gvzs/�]t.�Ȅ$�A���&]4���T�x�J���.��;@�}�IwK�!��~�O���Vf
A0i�?I���.��Hx�x"=���eX&����^,{�K��J�\�쾕�u�WT~;F�#�}h�o �O�����v�X�MW��y����^1H�&M#�ͱ���c<~�L=X�=;�w6怖v�v�K��*�id�ep�Y����,%�$�q�Auo�A'Dm��Fm�����S&P@fc
_Z��I�$�@��Jb@ڪ�Տ�x����sђ{Ν����|RA�0؂պc��֌;�.�͕.9�KbDqn��n�YM�"�a�����y��g���0�-����*�'�'�N�=�����}���R/�'�rYӣ�Ua��N��$��"�}h\�0�3?�w�����V����.�:t�����G�p�h�emՖ���7#S\Nn��Ŗ�Aɫ���3�,p��!Kr�E,ث�1��ܭZ�Qu?\-� B��0��x�y� ����Z������YB�Z���(��`����b�����lk8������� <��
_T���w ^:�P.Ѹ�Ĉ��mo[_�{?u�7��h�CP@S^���A#��@�~
�ݭ�	c������e�}1��[�Ɋ�J�����-��`|}D�����zC7O�¬2w��_�`����т2�[?C�*�% �̙�-���@�oS8lL����t�:���*{T�F}�-y
^�w�ܓ֍������3�mQ
#��ь����k����.ԉA��"�X�A��մ��!l1�T*���|"�K��fzݻ3պ�i�׀K��U�����>��i��j�2����1Ǹ��*��Uc�S&K�z����y�!�r'H-�/s��F�|E�#�yC�Ʈ���K�˓��0'K�L� ť��x�Nk/��Z~A��k�=:�ܴ~m�$7�^���и��HB�ނ�����_�������Y�6��8��c�[j���ʪ���S�]'����
{(t#�<Wf�h.B�t��x�a�B_����J��:VNuNtn]*ɛ�X�_�>_r�ޕ��>=�/�x϶�P�0�U���_�.��E���8�R/�͜� 3����0JI���-Bԣ�z>b�Ko�k�q�ӠG��dl^exH>^�	���ɣ��	廞K@&�ZI�n�1Ψ
�KFi�3�[���)�.�'BD7�Ӂ��76�b�_zdk$w�L� �+NH�t�D8$�H�>L�Xl����7Yr��>%41�������9����u���  �Oa~�����gN�p���Ŗ�����X�ދ�3��'(}���sqM`�Y�Իk4G����eM����Η�]hcA.0Otm�d���On�/��,Z�����$&oѤ��3^���]��9x�.ju0v�&�����[tH^$�a$��%R�_jܢe@�k�#�
̧�D^V4��v�ql�<p����l]��=bU��ni��n�M�9U�/7De �\���.�X9�́^*:�KRr-i���a��0��E]5���q��R���v\��w�a%?趰�z�h��얇�Yq��L�L�VAC$wZcǧ�!��I�. 9�M!����Fi௴�LF��2��g���a&WW��K{6������:�2U�"R�+s:��t�(΀�y�qZ�w�E�L�1��)I�/\g����"�h;�T-Ȼ�#Y�d�;:���=3X�����RhD�{J�H��0�+ɪo�i�r|xS����T�[���t^�j�¤�Ǻb��� K�R�n��C�*���x�6������Q�E�{f��ŀ^�&[��EG�B�|����:*j�-��LaNS�e|�f��+��lǟmy)�x6p2�#7�.��9EX�`lv`Z�9�K�S�!vcvN�2���S�V�NU��%"��
�W@�5�i��#�� ���NI��� 7 �K�U���?ȃݶEMF4�"[��	\�f��б�GTL�_X.���p��'c�P�rp2��֓��x��*�bD�����T���a���UO�3���H�+U���������&�%C`�䧍�an���Fw�ܝÍ 
 4o���P���Wmu��I`�p��~�5�,��c���1�����w2`r�z�D�f�$v�iS�����w����~ր�$�
�)�i����oE�}@��r�U�%f���+��u/�b��̍�8g&ˑ��KY��Wŋ��ѯ��*h�b�<����������2��
�*@��C+p�P� �q�Nws�DrKM��^pf��膊�l�=AO�ڒ�l�V�2{�����]v9�{�2}s�t�I�*��HAt�S��{�����Tw�Qև�m��_�9�߿�b�+k��U�x���q���O�V�sq�E�7�65X)�̤sz}hr�"�_�썣�u�c�ב��W��@$��n"sn���y�R��{CT4ۻ�� �F�9c�({E���+b&�	E�k@9�����w���������	�ϴ��2}A	
V���C�6q(�m���<dK�*R91U�H�l���}=�Ql�}!���Bdׄ��!���"��EYM�b�h��L�!Z�5��E���%���3����ۄ{��ş�š�h�ʆ��8�}�e���¦�s��<�n���}��i�S>ZA���ܘ�Y�9��L]��I��	���9|�o��m�܅�q�˫ =j����A��?Z�z�^�N�<���%-/}	Db君o�����ǵ�c����LX����6�:�|GQ�2`\ϲ��j5��a�����K���D�OS���s��6����WR��k&�/A��j�1z��7�?pM��J{��֋�j~����"m�?GᇑYZMJ�H���?U�
�i�9�`�Y��ْl֕*Y�K�;�h	5=r1j����ƏԸ����̡���������Z�����>�[�,�u�!|o2�e2���?�w���%iA�J�4{۵�a����!÷�vGrx҆����m���He�T�
���J4b�ہ��y�}����$JG�O��+T���g���c��U�'�2�?h,��:�T��*y�3�`B;���j/x�G$�q��p?�4�5�*l�ۖ0kF���huC��T�ݥ�i���Ҙ>�Nj�����6�I+:�(��͂
�q�[},f�i���3G=��w~숇��i#�h��ý�R�wΊFo�N3�1�t�D���xl������ϛ�{XI����E1
�+)N^-�6�2a��s +��r�f��dѷVQÀ���җP����	b�VC|�{�vי�L�DՑ��R���v���"f�����W�EkH��n���V�o��my�2a�4���.e�`M�oq����H�V���Sٻ��F�m�U?���������#���<�(/W2ŏ&��q�^q+�6����[2'FUyH��Z��SF�3}�D�����C��M�}|v�E���ٶ��y�Α-��?l݃� i ި��������>�^��,Ab��1&�5p�/�� �x�e]QkX�`y ʼ�o7`-��{Y1c�4Fʜj���#�����qCE�����;�K�/�Ơ�{�����p�p�&�!��d��c?���%��|�u�%~h`g��:�S��D�-Y�_�2�G~弸����G�ϰ�� �oh��9y ]�t;zA�;����|ʕ�_��c��5�3g@��9�_w�}M��<�C�"��#+��{E�ڊ*�yJ�6�C����td�M>	���`����մi�k��+ZY��'�,���@��6�S2F)d�z��ߨ�;��Ǻ@�d�"����-��Q�n$������͓̑�u�{��ðؿŢ�Xϥ�Z���v�z>���g��N���p��kS�RZt���b�]Q�k��ZǌDz���AS��}�ϊQ���Bv�Z��h�kl(����,�?���(����N�,���6�};q
��1��"
o�v����E�9�` �ݍ� ����{c���0�ƊԶ��xy���e��Q��0r�'�d�����5(��t@dX�>�;�JE�[+;����Ê'A�w;;�𼨤����n��p�3�j��'`v��}:�i�c�wȌI �He$4�������J~�5�y��fA� '�.�t7A�鳩�2ͣ�4*�Fd��4x�c���څ��)���v}�mC[�_�\8�+�J��Gj��$S�����?y�&���s<?�����6��gf�	�8Z�ޫLNr@��w�k�� �����A�.��m�?
e�<�J�ޚHB`_��Ņ�s�Aǳԃ�������P�?�� �wk��x��F�4&��k�ק]�4]������:�n3KE�q��:C����������7&��U�"�e�K��	x^�g��FUD ЎI�J3�V�B�*"s�s�6M��m��!t�:����˯&�˼�Q�b����l���+~H� �~���蔋F�����ysS������L=�v0Dq��}���5�"�T~�?��#�Q'��<�	/�d���P5��NͱJ�Y��0*:}�����wt��?c���P/����j��,N��%� ��D��rѩ �*]����1(��]�F�/F�N���T�(ޜO��A~���w��y3!��,�:����">1�OL�	�n0�ɪ���,j��U��@~�����@p��M~��ͿP8�؍.m����B{�*�X�h�Z�2��Z	��y�,�^_w�@��˨����x͑���g��z�|�A�,�X�c�}�'g�V�ȒϢw��� �3��6���[0W-���iN�e� ��;#�CBx=�4I	��2n��8��l�ېJ:�މ��#/EM�&�hFj�O���h���3�i^.y_�Q������1���ǿ,!5:��u["َ����9�ݞ�w͝<�i,8a4@��y�V���#g��Nu�s�th�#_��S���mF�o)��k~�9�#��t �j�e��A��k������s�G[И�/�A�x�Y��B�����z�j��6�薔*Ϻ�L!��*�$�}�㋣�+�G
"r��-%��[&~�F���u?b��?��Ǆa����r��Z�?R�����͐ub��c۳Il-0m��|݋���ƿК�<� M��m�Z,��� >�2lÏ�ꃴ�x8uiv�Q3�w�b��> ���I��w,j"�	:�x�T,��Ifa��T�g�G���j � }���=Y��'�V�4�󆐺�Aa�;ev�t��Һ����|ǆK.�b��ʼ�i�ʹ_���k�_�皰���n�J�:�2��uL~�u���h��e(��p1�v�ɡ�������UĔ��5�j�䄧�C$���0������G�g���P
y$A�}[[�����LruS,Se/Ě$����"2yR>F��SR����:���f��cd�`�B����~,VXB��o���R�l�M���?ȬP։۾��KU�@s��b�a�#�>��Y��X�G-W�vK�>��B!B��|��h�V�Rs��2o	&ܤ��<�hDu�J��UY�2�M����U!lx�@��R����Co�2^��F���yr�8�rr��"��6����{@"Z�
a�/��O���
�QW�t@�
���:[ k#��T��9��b5T��U��q�M~m��a;�ӊ���5�p%��do�.�] ��s�}��6f����#5���M�_�V�2-y���]Tں�42~�i��-�-?�[�?���T���{���b�1����A]�ۋ�%VTf��؄h�~|h�5�XQ�"nA�=�O!�F/�}(��ؓ%
S���"r�\��̾
��p-@P���%����|R����� �k�͡��(��SV
��N��A� /~+���G�κ؃&m4ܙ��ԏ.�R�_z�պ�Í��g��f_��|���vr�w���^!7��H��t��'�3��~�$�O�k�޺�謅U��Ay�ז�]�r�_��a��,e��N{�!vߛ"a|��3�&��Hƈ9�����x�
�3̃v�?'=��Xh�ɬlK������:��Y,��MϺm�lg�k6w��t�We���*<O��`G�l[��fg)�tV�kM�U�tL�
$�-��6�C~��RA����g�q��]���$3�]�)��-9���)�G�*O���A� �V���o���8D1�
�$�yV����� 遑���H�=��7���a���m�#:u��&�~_��M�p5��jԀ,,��:C����_C��<�x���2��u �m�X�!�@(��!>]���D��ߨۓ�֥��F�����xr�Tz�4*�tJW}����u����f$-���_yɑ����g��іU"��%k���Qe�1o0�����	�L�*�_��j<�����HX����C?86iR��*$�#�Z��^�`���#�	S��e�?[�M�*�X4���d\�G��[TrOG.���h��|�'Cd��.��s2�Gœߓ�����#�('�/�B>�
��� ���7gד�P�VWh��J��^�D�x���Y����#1?~�����+q����������q<?���W*�o=�ֺ��u�;���f�^+�ŏ��g�5I1������9��_��@��s���L�'�_Tg��� H��3'xGrAO�4!�����Ԋ�r6�ǞeqįtI�;܎�FSE`�˳�qT��b]����L�,��բ�=�D[�S��¦� �̐�pDW��7?y�f�G�����9�W�g�;<�xv�i��_��^�
+�Z?:@����۰�]��!
c�gm��f6-TIY`V����9�ąhV����cՇ��U<��5�:R^�n��yQh�6�\^��<+VNX�5!y�c��bV5S+t�M���*�u�?F!�}�Zt�2Zt������T��������[3y��n����絇��ԖG�;.6��b�;����`��p�	��(���=!�y(W�Z8[7x�Q�oד�.G-��m����M��4ᗠi�����$8��3z���9����#hi]��Q�
�%rt4��9��$o���ږ������7'�m��*Èi�ǖ ^�F>ș��y�.;�K�����]�/%uE~�3$~]�x�~�ٻ����,T��}R6�x��Ɋ+��%��^2T�Yɪz}�v�{WB�=>V���{���ˑZ�r���ӂ�����_R�IҬ���o����9�� �Q��i��i~������x"o9��Gwy�ȧ���8��-��v@,���d�Bۉ��юB�_�M)��/95��clpwɹ�bq�Ѳ�$ں��M���AR�K�o�r�D�Tɒ���wjn�e,�ub����l_@��i�/Uk��tx�����S:h���v�{+ ��JĖ�F^��B�dRxC����(�-s+�2k<���暑Y��fOrrj����	�LZ�L�mr+���pF ����	�fS/1�%<�^�yg��%5P2G�D� �@:d>j^�K#U"UF�8G�vވ.�p�G����6�Bݬ��)��C�Y|�����}y���M�tM�]pKD���m\ �@���?:b,�٘=��AR����E��{�{�|�L�^���h29��GFDEo6�
����z�]r�5=�d�8P@!��\M�b9JϨ��$���;�3.�Ţ49���Bx�E���V�wB���@�Mw6�1FI>ʦe�d��)�V�]��2O����O����gJ�'�C���9\�U�!�1:],:�d`��egb��h�r�o�=_��+Զ,�!�Ѥ�`:���a�q��4�q2�Ewz-�#!`��3V��M��9"y����Y �YftŊ������G��!M4�%|T���S�bU(w���Vڰ�A묌�T/eZW�!�r�d?v��!"NS=�/t)E��>p�	�ѱ���'�,�h���{����ZKI