��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw�a�[W;���(���=�+V0�[&�v/9-�ŷ�;��Ў�~t��W�W�n�I�T$�LR!� ��\��H���l���&�'Se +��>���6޹����-�2��6���EM�Q-[�4��mx{�7.���DI5%�\v�����B�t��r�E�fl���vO$�.����@��2�G��b9��`�=��邩y�<�����؅5��*t0���|��?y^����튥ӻ�7�tA6��[��Vm�d����w��J\��a�$c���VQ{JU�:�'6!zK��#���I��g�D�1�2���[����p�d%�]Un'�}�8�*�-�6���l�����KW� k/�.���@�F�d|��?��2U���9J�_(Y�Wx��$�k6?=ƣտ�7q<�*��)���6Y]��?\��WI|������.S��vG��|���h���֯hQj1Ht���<���ѝ��zR�̾��J�޽[�2��\��a��!��1�yU��$J=�J&��#1�L�Lx��$�$����A�����G���CA�.�kM�@�*u��B	<�(�E+�e\ܯ�P'�.��o�F����8wpQ�>,bJ@V+7TE�멖�+0�mknB��񔹛&���&d?�T	:�9bH�zqyC���a��k�W�u�p��.�^��,�k0�Bлi��L@�ؒ�m�no����,i�o��L�C�%�߰���R!*2HY��ʲ���ܞt7�(��T�� V#̒&�8�}��X���lL�S��CdS=�wΟ|�;I%2��D/H���,,��W�2RcV��E��s��h8Q#p�"{�:���G�dHmI̐��,��%u�x��}g�9���002�FZ�y/�^$/͸��*��-g��f�]57#}�XA��	�&�wPS0�fȯ�B==I<gXj�]�4���i�N"�a�w���Y��]�ھ�;����E������?��n��E<���:������m'Pv�� &�<TW��Z �7.ߪ�e�U??3����:�+�� ��@܇!��J�j����	=E��P�환���L�r�u��x�*]G�衊|��T׆Y7~���w��cx��7Ǣ��bd 4����������@���O���Y��ʴ	Ү����Z:�UC���-V�*jb���_���÷V9	������^� ;��%滩�q8K��k��f)�tc�|�l��O>n��g���]�6�U�m���U
�1�-�o�>Z�R~�O��t�����բ�%h�����ʐ	�&����;���E_P
��	���B�5 ��|�^�N����̠-}V��)1������ԭ:g�/�K���w,���H���!m]��%E�!b_��[ ï1�8I��8P8k::4��]qQ�rB�|��UE�@��P��	l,�@�NJE/�b�OG7٨���֣Y5�YzYކ�P����"�l$�kU2>6(uh�~IT%yCmdj���s�<ՠ�����1�*@[�zG �=>Z�H�DN�O�������^ƮKgaco(
��� D��%�V�69έN��ێI2�➻ӿn�X�ؠ8��UwP1
��u�
��%�� M�b��4%���)��Kl���5��_a��i��0��_]ZZ�-�p��4����J��=E����%p{�艅?h�4q�l���E�li�?g��Z!�L��ʏ��K[7��ӗ@ϙ���8��,K�,��Frdc�"�/(:@d�Y���a���0�0�)o@H=��)�6YM��jأD\�LH<VQ����BŊ�.œ[�<jb�ݨ	��x�~h��+�Ĝ2m��C���1��A�*���>��;bf�ޚ��Ha�oܜ�7d�X}�z.�,�l�����Ϟ��j~f��~$�I�p��f�J�C���
�1S�eUiU*�vߟ���{�6��m�`�w'7����,���#��O6ږeF�,M]��W�'X�S�'1M����(ܽ�^�A֜6���N͉�)�P��P�Gav���/>�v�0"g�s�ɚZL�C�p%A^��S5��H
������Dem�kcI�Lޮ�艳h�M*jmM��#:e�����e^���1�N
�Ԟ�ҐZ�%-Ai��f�c�;c���t,d�&��=ϔ$K$�~ܦ��[�V��m��������%3�mj������H-
����J�E������x�$�ad�Č]�-+�>���|�NA-aPM�O~K�}Y2}U�I$�M����b ss�K����*��\������_�	��+���1S�Dmg$��������!�b+��O��a:ڻ/�M�D
ǨO��(��q�R��Q煄�V��\����ݻV��� h�(+��dM����
�x����^5:�8Q�uW�P!^�H5�r��fI����'H����V<��aw�z����������/ԭ�����o
t+[{T�����7y]��Xv�h����JRrG�$�)�����e,[�2��_x��A��[�J��}����6�ޚW^�tm�<C>�:�4���0Nn�'�&���	F��F-R;�6���,�(?Q�
?�iLY!��4T�LSM����襖�0ǥ��8��zx>�]#A&�zel�vX�bEppD�<�A܍i�x�6Izw��Q��O]�d��1�\�>�!߆1N�oxq��wex���2J�#l�X=�
�I��AN`���>��"�~f�-F;w�u5-T毴��y���p��sٚ�Mm�/�|��X�K���j�8��>>D]��8C����P��~��U2q��e�RK��no�������a;�mm���y�(�Ӓ���x�FE�<���Hn(X!���P�e.�r����L/�O�뽵�Vjg��":�f��>
�K\�Q<�^	��`s��U��Sí'�>WG��%�| 8 ��Im=#N"�a��)֩N��H�FC=e	�[�s�.�D�H���������!����$�ohu�<h}�!%|��f~�����Ջ�����=#6���]_J�W�L���,���E�Kd-���3ے�nw�>��y����d@<k
s��/��:\��Ka����y��H-�ҥ?�D�RR�e6c����T(T��1�����|��3���K�k�!�`h؝ZS���jsr+zX4���	K��y�К�r�N�F���C	K(����G(D�+���;��U���r� �c���v:�~�k�DI+��"����1�g������2�ܐ����ʙs����VA���V��$?���w슢�������9y�N��O��m�v+�I�*[(�7�"<�Cf�@�3X��Iw�sO��,��kOtm:��t�K�˰{�)T��k�**�_D�8G�3���Fp���Q�Z�D2U�b���O��1��O�XO�_��~�� /������l�������(��I�&͘%���?�_�m�8C�:��Y�l�'�&c[3�mPA���ʎ8�s��\����������(֌n�%��;�e�PM��q�f1�X��1��s�+�����K:{r?�LBē/m���F(�;xc¯-��=~������[8��T��u�M�6"���T��.�}J�����L�íu��/ՙ{T�M߅��4�{���6s�I����v���~\� U��,��=��#��8��8ЭeR��4N��R�D�0+rr3��~�&��}z�hZ���
5w���S���3/�wG���!r-2Hkm���z�zz�V�;�J��D�� ���͜���S]A�ga����j;9�M��pY����ܶ1��"�X�{�^9��.��D/ސ���/1�Wc3����T-�l��x�����pm[6&U����q�:1J�j�}��gڎbӔ[4�c�V��M��2��	�� ?�us����(��ԅ`��FL��^-	��C�+����ߑ�N���H�����'y�:&�4���r̠v���٨�Ga��Z�>Ù֫�g���T��BͽDY��8�wX��+��ك2�}�Pߟ�:�m6�B���k�=I���eSK�]�g�[jb�&T"t�(S�;@��;�P��,��5�9��^�׵��9Ul�l�+zk�Ԯ5�W���Uw�#�����Y���;&����$K�F�%E���R+�ڣ��
f,M�ױ������i}Z,M��0�ߏ.]?V\��H_�
�b� �*d��b"��:�3��~U8Q^GE�Bi<����3�3A�Y��t���:��^��=�PDe�l�s�r-%�%�!Y��m�gޛ:��sn��G�˲K�H��c#ʭ��R�v���΋�������)��Y�I��(��q�?L�pE�q�1`F��_#-�͚t� ��~��E���ݍ���
(ؠ����eMf�;f�}:A^�Y��N0ƲG��n���ʳ�h�0�mBU��9w��ȸ'(r@�/���G���C��'=*Ԁ;�'��*����J�����M�J���kwkc��E��=��RP>�f�Y:g~���+��]ͥ��h]*�JC�Ar�y2B�j�?�fA"�s��}�jhY��O:JHS3x+S�g'0rc�����+�C�����~��x؎&�i�eR��r~�	b?Ў,��E����T�u�%��H�^#��qA�6�����>����\ov����O��Vpz�&����$��]��L���m(,!�V��~�!5��S��Ry�~{��9X�\�(}�4T�����V~���� @Ɲ7n[I�٭��=�l)�*Ɉ͠�oQ����n~����X��E>m�D�����.ց3�'=!�#`i�p"�G��RN�H�� <�<QRO>Ŋ1S �ɞ��6�!����:[��=��l���C�v�{���2�ް1���&���~�NW���ίWH=~T�t������_��儘�c�O��#���\����BYRq��X��skH���v�%���8�X�6O�o��>ٚ9�if= s�`���j$\�K�E�	.����T��o��~`ni`�L�YQ��=���#��)��̉��J��C�F�W9���B�b`KEk�}:�D��b��MTӅ8%�|@�wO��O6<|�4�x�te�`���)��9,�{��5����Pm>Sw�� ��X���^�{�^���൓���;Id��v����ê��q��&��țo��s]b#5����!E
S�v6�Ib>:ƴ�*�۽�z롡 ���V��{����S�6�{}��_�2�/�½Ġ�����y"��?5.&D$~`}��fbŊ��;2�w��s䳚ql������^ۃ�m����)��&�����#�# ��c�1�qK|�ڙ�z.����"����|l�c_0��E�DP���{+,AjX]}MB�	�d������F���6�)CZ�e����:��/�)��[.]�D��5��m��-��%)%w��h�ѳ��eE��n�E�w�	�q��˘�YZ���͠�7S/(	�h	���طڀ,����>�:`����sOF�	K�E6/���eB1iolS���n��<�2^���Ew/H�i<��=���A�ݞ�d��|dpJ�	���Li��9�z+w��f�g���]�e AG8�w �TbRɵ����F=H�6�lF�ȡ�[a��ЮT�)Fu�+����z��XM�� �BjP���e������\o�Gq#�8�c�d� ����?<�W�Tk��U(#:ҁ�z��LP�� ��=�@�
!�,mS.Z^rs��)�Y���JI���)}.�Պ!�Ϩ�J��V垙hIp��0�Mͱ���֦�BJ���Ĩt3�Z�����i
]��HI&װ�E��:N��o,"�V�f"YR-&չ���sʮ�*���oV �<�D���5N��{���4�"3��
��+�έ��"�tx��"a������R��zrlަ�c��?��O�傪�����q} �hQWH,�@�L�W!�R��"�l���΂�8ٰ�/}���r�O]ygC�f�]�_L?۩x�����5�����vH�o��;^����vO���]�d���j&�)�f� @�S���i�Xm
� ��e�B��-�����|
���Y/C�Mu�����fW��LD�)��EBpo�B� ��00�ŀ��Cef3�Y��GUJ� y4<}��׋1�O��(-�����|�1��.��=�f��N���(̄���>�TD�� $>j\}#�^SС>��h��0���?8�^ћ���eM���
&�R����d����}}B��~Mk�	F���g�m3J�y�y��lvJ!{(>��a ��_��z@�Y�%�6�P*��o*+��b�'B�K#�/�]q��V�\UT����i屼F��8���F�����Z{��HGj�X�C:ּ\�l��է}n��l�����Q��������(๔���w�J��;�~v��-��#�qp)Ͻc@$����b}�gD��IEHo�}R	�\��S���+��$�ɡ�Xx��dK���>��c`�XԐ���}��
&�1
[���'��;�,]�{��� �=�t` ���i!�U��(���'�t�F:\���S����PX���no�DX��sC����.dMDGK,ϴȪ�{^�l�����rN�B�l�'�������=�=�~tuӍ�pVOC�\։A��
	mP����y�TcGeI�EgM����>7i�m(���?#$jRr�*�&� Y�.�S�B5���Ʋ��b��2v�٧M�/�ӵ�.�p�h��X��I��p�������֨#��H:5�QN�\S�rɋ�7��٬G��-������z��S�F���O+C$+��y����m�