��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���;0���[��q�N/[85��1d�nޭ�!oX!�ذ��p�ޥ�4��^H��*��i�f�m����l��&�<�]\�8e�44���k�t�CЇ�+Y����^���($�?�`�\!��?>���l3�d%�	�]�_�J��^���׿G����y4����bI���Ѣ �4�L�:�,nmE��HHDJٰ��B��A/Y��́\MD{�+��<�Fb˖,�r�I �����$^�tL v�z�ڥ(������k4zV�%Vd\�l�̽��b6��C<�������2�	��ډ#�X���sYag�v	M�¥�.���9��䴘
0����m�}d������W�R�S<�V�j4I0ҙ�fd���K�]�іn��$]��z����}�7�O`��r\]1E%! ��)�)ua�(x�= :��i�(�1 \�ȁ��S�ر0暢f����0z%�d�r�3��i���N��o,4�E�BE;��I~�1�~3�����7���Eh:i�]�1]���d��Gܬ�o�x���P��+���Λ�)�f�fj�gI��C�_|`����igE���Xx?��\Y�M��]I��&!���]<b;	*��JKlcP��Θ��Z!F���d� ��d���Fw�-�ɾ��e��Z�Q��Bo9��]h�&3�Dΰ�rY���cNk���$�>��6�	�B_��K*��JΎ��t��aB����u	��];��26�Y���?��5�,��Y����������*,���n.<��'���m���� DVA�mX�G�"��\|ޠ�ᰬ��'c?�M�k�JO�@l��1�X�"��`���C�Y{0	j�k6��	,�܌�i�?g�f�����g1�L�ߒ lP-.�#�ِJ_�}������������r�v�-}�Z�>Q�м��#���k����篹�ǆ�Q�&g��
�'hJ�#��(�@:�/�kwJ�h2�h�{[���/�E4���o�@Y{Kj�Uo�c�<)�-P%-�&��"��[��p��wm�����&C4(��,����G]�F���6��]|N��N �T@���J;f�Ў����ɢ���>*v�DD��Ss�g�iu7\��j�d/�� �%�u�F��g4d�O�8��FT�����7���1�݇�Q��PW�l^��硉T�S�ˉ22�Y%L���_����)�I$�6��u�R������ ����̀lf�xl��c#Hx��+���Kꢝ�?�Nx)4q59ʋ��A�I����0pk�����@+ƍϧ�H�U�j��W�ܑ�b�&/��VJbs�Ulxw��`Z?5\.Ne�F|�V�>������_��m���_6N��w�����:d�}A��1�#���9�y|.��Y���Q漿��g|���MG�U�T{;�؍}�R�t���T�1J���V�F�%Q�l*mI���A�U[IRɃU�dxs�Z{[^�JW��� �Q�(xre�O��ț>��t������3�b;X�D38��У���r���-��?Ǝ�D���7@�u��G���F� �:%�n85����P[�_�JP�kj3a�0�����/vj$}Z�An�"�:A���4و��#��p%�-�kI��uf�ղ��%��P��,��<��J�06�	������K��Q C����}�/��=�Ӿ��K0����q_D�>TP����)��"�vO̝�}k<�`�V+��3�)�i����-F��(�'��?TSsBA
9��CU�[uN��BKz�"�G�g �Ķ�E��\��A ,����Y��yX%�M��\)�i��2�GW=�Q6+w�ӽ��O��:ǲ �<%ߒ��DM�@���x��_�:����p�K�-�U�M���W�����i���Zs"X��vڗu~�y<���٩���d� �vjX��[� ��yf$�3�?�g%{�Ge�i�UYg��g�e($̀L����*��UV��w���&
S ��I��x�'���ϸKk��6��ں(.]�{Vq&`j{F���W0L��4t���sr�b�dzt�|���U$-��E�a���rO>3�\ف!�H��Zy�8l������0v�46hΫм� ���e�!�g�*��z�R�8W?��A�M�t�C>Bߘ�Y���y�ĳ��>��<�R���
>��^��o؟��G�����u´	���������.��5U����2��t�"N:������K2{)G���l��t��,��8��(�.���x����л[3L�!��i�!
E���^V��wzS)�t��L�]�.޷B2�%9����y�����o���{�����7ԨX�B{�Z6:�,������k�5E�'�� �F�e'Qv}�z��i:�Dj�~c���(��`�D/��<D3�ٿC�%b԰ �t���4�,�;����7�k`�$�ǎ�1�+ ��2�3�;o��)�C��� �0s���1�j����j4�F�.�3!�C5��-:��l0�]^9M�C�J����.$H� ����E��J��X�bj��܆I��P���b�|b��<	v$Q拰?P�b��5����/3��	�"z�C��7o�1�:S����U-�9{C�`��Y=hj�p��K�2����yd��ǣPf��/�F<�>�͝r����x$���py츱Z ,��T/���v�*rx�.��dl�43�h�;	t��A�B��WFyYp]]� j��xnMv�ipLL�Ck!���gV��֐�|���-#ˡ�0��K[��<^V�T
Z{<�@�H9#	�9�-v0w�k��r�rP��������6g�yd:�l�ʀ�$[g��<�gz����Xؗ�'M�u�W���^#}�}��{�������rb��K�'�5��̂�<�!ݗV��Hv���L��ޗͮ���|�n%,�_�R�*ڍMLGg���8���uŻ���� m���H%:ŋ8^O�_,�/��RK�ǜ�3�1����ȷQ��NVOypo�Y3gI�����).A�;v�;\��,��҅���Z�@����7�l�����ZB��[��]R <�w���$ ���*(y�DD�N���.f?`�!"���H�iɛCgi�k��Gt�>��v�r��!�F2q̰�>��I49�|�F�f��kd+��>�^�qe4LBu!����x�j� ]������<�
;���kɃ8j�����"O��G���k�Y?�B��H}V�).}Z����a����E��釯"o$�^p�cU��Y���a�Z!�G$갋��va@Q�`8Sq��G�P)t���V(n,����.�_}/D�xB����l6����?Ս��������z���V�`t�J{V��U������{�CN����@�+�5�;د$�_a�;�'�����2K�< ׻��$�/Z�_S��X@y�1�}�3�����O�>����z�68�(=
C|��y�x�:�o>M�ԧ�A+K����$1���^
�\�3O�����8�]��.�T�Bp%����@Q�; ������f踗�4��M*c�������Qʿi/�Z�L"�_�İ(��oisɨ1ua"7�C}k�~)������1d���b!u*�� ��H�eGT\]��48�	�&n{�@5�����f��H�5i�A4��:�Y9�+���{zF.ox��"��`��U�ωq�!&���`k��7mʧ�	��C���B5���oПԳ��c1���u��s)H\ņ�!�E��!�(n���MX���'j(��Ӱba'�Kv����!����x,��P���y��l�5�H}׽�
C���%��Z��[f��3��5�����
O��C�l�W�k��y?d��8�p��68O2��m��L����q��T�ۉTq[�m��C�|Q{�Y��8�"�9fb�P4[�Mٙ;#�O���]¼�%w%�>t�����}l4zh`̯�mV�����l�l���|�v?���Z�T>��r[~�0�eӗ���G�\T/�2����c*�g�C�#:ӑ���2zZ�p�������B��v�Sx�@��޳��9ܛp�Ų�����3�]\�Ir8)�X}�T�-$�B��Ø�T��m����SN�}%ӊ�����ϵx��ݫZ@�ѧ��փ�G�d�i̜D		�\���b�E-ac�Q	���	9�2s�B�ԩp�����F��1��)�kV��/��1Ցz	��۾��f-�j
����Z���������8������/��&A�s	e�j�:B�K��ȸ^F��J�fE
9�͟S|�-�=�1�0��a82-y�$��);űa�!���-}"䏗K�\b0ϗ�O{�e����1p����Y�R�b�-E��TI���q�h̐����<ĊQa{Us��<�w��|'���L�0ʺ(�;|}�$�$�.�<{�8�=�Ȣ�,&V��Ii�x���Y�K*h�f=�@�����M�gd� 0��2��� 	��+�����B,�5�=�1�r;�p��/��˾S��^)4���%s˵i�WG��	��]j04�tڻwϨ�@�ĳ�n~Tm�4#2��),��tHX{�>��qFЙ�`�h���f�ڢ
G�����V��3N7F�InLU�L�^�&�k�O�������2�|���5|��k%��d�Q��p��ǫS�� �����PO���ш@2�Y�M���B�`�7�O���Y�� �
���	3���)�nBy���o�6��}P�E�������[NQ�ʟN�t_k�	�эT��@2T,Z�Lut�eE[_t^��aĖ)8�ژ�w�ڕ����g�[vZ&v��~�JF�dm-�w��af�n��Bp��r�vg��ۋ��ŉ��i�W�%���P<��^�A�}-TD�]�K�=S�F5�DU���k�Iud���}��7��g�k��脟��L�ZCZT�łYk�7V�	-C�wn	�PŃs-k%J�L��m$uIϡ�$��8Ċ}��T���l�5j�~�F� ���MzD�G�蘻~v���R:#�o�O�X�ǟ�����p�,� ?]~u�M܍xK�?�8�:!��,I^9�'��Y�����k�C�}�a-˗j�?����ɼ��R���t<�$Z�9�[r�a�D���%�E���C������4CT��Xz.�>N�-��
��_|"�[��.��4h	w�m/�20C���!��� �J�'<�����5ט��=os�9��?{����i�������|����M�����l"3���Fݍ��iG�G�F��R�6���J�k��1�a5�"����On�5C� �[.ƤA���(�+�8}f1HT�yȈ��O��@���M�Z�����&8��������\8��D7<"ڂ)�z�ܛ�[.G��&:z]�4�<�f6=�pU���Ë(�5��)�D��1����1��O�I�^��2>7g�L*�T1�L_g�vm�춧7\ Q? :0�&U���l@6���=���-i�x��/���%A� p��d*��gY�JU �X/Xb�(��O�wZ�^�?H��!6�ǜ���C��Vau 3d|U�p�V�]�KS��c�z��}�s��[�3.�[n�L��s�~��¿?D-ڿ#6��bU�mo�Ij�F���0�}S%m?[���L���="��+��̒%���!p����}��J	��J�� �m|���K��E0�M1·�&�ak��Xh�YLG8ן#�P��	��![@)PBJ`�ȎtԕE�P]�n����tNwc��?��C5#:��C�Y�����y�Q$%��N�~y��?��%��._E#�=�]��C.��9���I�(���nXv(A���W�d����6�0Ļ�<"]0kF�� u�a�RQ�#�z>�ަ��g�� I C�i���������ؿT�hY)�s<Y7���WeQŮ@w�H�*�=lؖ�h� �%���3� |Hd���=-_���zx�������)�c6g�T��j�g��g��	�L5;[V����=OCȪ��;K�e���i��Z��1�hh��+ +.$���� 1��+p����7�F1�w�g,»�������.�b�?��g�eN}V*�<T��ی(�1���{�4�A�����#c#�᯵��(�&����pȷ�S
��7�yv��)���5y��e�/���8bY�1�ã�1t�lXZE4N�9��'H�X 2�z�'z���^�O�M��jH(�r������(3���@=��mou�oL~wv�Ɇɦ�Z�~2����<r��%��]���-�9�'ٴ#HV*�j	�*dz'5���7v�"�)̈����Z�g�������X�}Ñ�Hь�)vK�$0�*��lLrL�9�r��Y�tiW����5���1���>�xRv��6D��Q <t;�3�����}��q�`-��F���+lӋ�j�����m���L�p	��j2|ݞ�`d�$�j-�{���ќ�wIc_Y����n	 �S�1t�,!�JY����K��2�:���6������\�]����#���;�W�$:�]`��C�TݖuU0�~Z�[���+hzX|�
`'/���g��[��Bf|,T�&Yv���%u�?
K���rM5"43h%�M�}1يn.�d�U��@eW�`�q�xF��vzDk��W� 	ˌ�C���e=:�+~����.od�O"1)격/���&�<�#o��;���(�����̥� m.��u�꫖,�lj@ߧ`�Ts#����lן��U?:�0˽/�Dۂ6����Ü*��6��|�?��ηI�9�c�f����>2M�Cl
�����b>ꤖ�)ޥi�U6�ΰL�d%��Y���k!z@�!'E��tAO�-j�4摹�aU�,9�v��ȅ�č���q���Q�`N�B4���OLO@l�HvD��<>��Q�K��+�B��@���xT;s�E�Q��&.�=u����@,��chv����i�	��S7L��O���E�� 汥V��Y�~�=�[1�7b}�L��bG����;2�s�䟜+����I�F��S*T*T�攊R�����$Y	�}�d���Q�
3(\�qǱ\n��R��K9A�݁�����_ۡ;�D3�?��ˡ9�
P�~��Ĕc������P�Y%G��r�rOq�-;���U��>��m�A�q���AR�p�=���N�������gcՠ�9ϴ�I�v���# ���"�b:s[���i_�B�=_B� `�ߺ���(��6p��e���Ժ% ��ҩ:�ׂ���AÂ��'�%�2s�V1�o�A�����"+ۆ��d[�����y�?XhF7`��2��1d�0}�2�)���׺ld1tK��g�q�n$�]�d�	�$�J�4]<����N� �޼#{�~��?\�E��[@j����`��!���Ѐ�I�[�\T�zY)�a��P�#7m��MhE���d����+����N����q&�vZ�݋0sMa�zO��?6ן���ћ��v��lGz���p�CL�3e�i8F���2*ч���Գْ=�u���'õFh'[]ś�Ң��4&����^�R.�"��b�\2�O�b��ju���b��Ѵ�5]A��3����G��yGt��d&�+z��OfŕI���~������v2D��C�u���d?���7������b�Қ�ϭ`!�Ʊ��N:����;��jέh]{�������`�h� ��Vu����ӏ�?����0�Q��2`U�7��wQ/NK��W�퐂����a� �n}�NGf��z5�i��(�º�8�3C}��M��)�?����.�Hk�O$)5��� �5w(_*��ä"a�������y���i�O7
���)��_cx"#
�#���A/�6��ȼ�7�������.��NV ��(����t�agM�5K��7޿���oJ�BE�(�PRjՄ���궁a�&�K��׍gr�$�A���/'4ؐSX��L�#��]�_��ya�4!���\ �����BI<j��($�D�P����X��Jߓ�b���o�����{�I��~��l.��_s���>��T���4;�S�KB�6>mZ�P�>I�N�j1��kx�y�3
áM �z�N��P��j�9�?�5X���Qs��n�cv�x˂x0N	r[��_#X�W^$���#T��b��;]+ɫҬ'�̿����<Ib�q��U�SJr{XNg�ƅ���oW�&���?a�O��F��O>2�T��
[�]��]�na-9����v�3+ҥ�����k����#�w��M��|
� ;I�Ǭךʗ�l�ɄF���ֿ^�i��V���4�[�!��W�a�m�!D}� �`�6�4��S�����Sۆ�nG��u��Q1j�t�w�Z.�ik��t����*�|U_e�$����7��:��KB�v��ڌ�
N����q,��� $�f�� �@��s���y�M�#���z�|Al�e��������������s�h<.Lȴf�;q�,=s����-�>�����%�{WT�2��%��:}+�<�OH�]{;K��{��)h���Q������Q�55)HA��T"K�M��F��s�9#�4�zw�k_[�V��rDp��O�����6�JQ�E)���#������q�."��`�7wh��@����⠿f�&Mt��GHk����uh���<8�%C��҉t�ܥa�z���#���,	p����$G�0Γ�n���Ƀ7)C|�05�.�bvK��J@����b�J��9Nџ��\8k��t~0")F���K0����N���GWB��V"FB�7'k�
��{�r��s�\<�8.L�L�-�?��q
����44y��ս�;�ZQ�[�U��΂���̠ΩC��T$`��+�i�����>�p5��L���1�43�_ �n�;�`�5<ö��w�f���ѯ%��^x%���j�x����%Cy����F9��Ш2f
�~s�TȐ/u�3I`u�1��g5.�� �T��<����:xO�q�������A=�Z��'\ȶqV�e9�O[�T�Y_��M��J������Z�0f��j*��s)���H�k���+1��7���\�&�;��/c��D>����L��h^�w5�Ɂ�����o�׭�tԁ u�˲��@�f�>M���m4Fb5(y�'[Q��#9ǽ*�tF�w3��
��BVR�nv=sƂLVh�١)�֑���3)�y�
��ȇf��<O_X0��!MW�+�K��q�����y?uoΛ"ŅI��D]�Y�"�ꮕd�B2$5;���c'���V�s%R�$�F~hP)pSd���Yv�{�B��}ݐꐀ�Y�V6��C����K�O�Z3g�m^q�H����j�j+�?E�������d5��e#�����Ds�0Q��}V���c���(��X�����Y4m�e�4��j�Y��WN�I'��dBpH�r&�S[����{�SfXZ��,x|��%�sm�:����m:�,}񭁍���M>�\3ӎ޷��U��)�I"�HH*1�y������� !H�<{��3͡U��"<�e~��D#Ṿ�x�O6��lC��'*ҟ��� u�_��8՞$J/`��.X�(&�ꦌ}"[Ky#0uzɑ�I��T�j�|)�r���������t�?a-����m�s��Ց�n���-K�Ck��9syϱ����ҰUD�"���tS�7�%T���f�Y�����?�V�Y'oO4�w�����_!SrS|�L�y̠��|���0X�<���VX`l[���.ip�.���J��KE߲�a.$�B\LcgF�M��5�x׋AG�b��q���'5@���.�ik]��ZQ2�<k^i����-'ZJM���ѻ h<����gwa2
>&��O˜ч�8�fI�)>��-UMt�v?�@B�3(2����zeh��Ǌ����N ��\qO��Gm��'���yEՙ�Cc�n�h��)�~>�����`��9�Bj:����F1{�[��H5~����G������T���&��Ԁ�N�l.���|��M��dAD���ӆ��A���ZFzd��5�8��0�t�y�\�6L��m\.���hX6	c�
x+3؜\Uс�����Y�V���,��L�s��@���G.��I����^WC�g���7k�>%�n?ֶ!�9�1JlC�s�/���d &��_�VN�}˟��g��yG)z�}�>�-���x/��0����ÁB?��'�aV�셎f��%�&zγvۀ��.�~�4+�WpAp��Ι�|D�J��w[_D��P[�:u\�nc���Z:���F�S%�[(W7�hRi��@3Z���+,uq��W���D��PM4.�?"AI�/Cc��!!^g+�l��9j�D��/W#��.�,wp��/�i;	'+�8���I	�����c��1�S`bu�:����8��E��U�9���3]4O�z�FGk�pڦ35F	��ʒ��0 � aw���fBJc�ȅ^����������h���{��`��i�V��D�\$���ЖW�h�����xk�w`�ӘJ��uc�W���,�if�s�|�4H����j˿�(/���=ά+����6z���ˏ��mh��&�	4l�d�s�k���8i�uLv�]	iґ�;Hb-�\��}���	��[������7�p`�9�Sd�톑A�pK�͖24�K�)�^$߰��MOe�p��k��4�j����)D芻i4xR����!,����i-w�����Tv���_�m�H����y<�u�������n�H�K��\K�M0�p�c����ۏhh ��lT�e����yը�·����z���t��'��ůr��0"�(Ua0�y��؝���=z�D9�z�#C���NS�l���bX�0�QN"��,�f1�I��s�)����pNzo�p�|P����W^ԿQ$�D��Q��0���9�b�=��?X��xlByP�,�D3;D�|��JSE�~�(2��?.��<�8�u��^���*H=�ԯ�-�9�?((����[ݶi������Ź0$eE�=UT͈n$L������*���qҽ����p}�L??��UEYC~��n4������ҒG���H���U�����㮈8���ED���r'6��3FWV!���=b�ɹ�����~���E�Ҫ�J�&B@�v��ZY�[W�-)x�MG 2�x��	R�@,.Χ �J�	k�"�s�a�K��`
g�QE�x���#1�f* ���M����if����<��?jȲ�>�����~���1�X����'�6&�Q�g��K���RűBBf�:�a��ܬ��-S�|sx�S-���c_ٜ�^�Ր3���ѯ4��s�`��h�"B�t݃��N{��4���]ҵ��e���؉��4 ��/���.�e�6ｏ���坂*vv�-t6��i�ɻD��8̼�8�=&����[�����z�5�H2�a�W&�ڳы9��T�E�^n�JäԽ�S���U��6p���5��8}*V�Y��&�G(A[-n��M��E�L�qu��_�eQ�9��1P�eO��B��s嬔���}���VV��7���k}P��R�%��|�ੜ#�X^�B>I++��5=|ųoj*�^g�׃�6:M�M���_�U[��^\�s�\k����)�?GXܲyA (�1[C����UB�9ԝ�\`���S�8
�����8@�j�~��h�L5hw��D�x�u���M�����bځ���I\.����Q�F��/�Z%����Բ06���Ҵ9��������G�AO�7<,�B���u���d