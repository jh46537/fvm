��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQl�E��*�����W51R�@0`�T���D{&l&W�s:�-�Cj\iZ���*G�W�T�,���*h��q�E�_j��v��n�����V��~Z!`�@�������Jo`����ح��禽�ufL&~�!:ubs�r�SF�Z��s�Ig��_N�i����
Uڧӫ��e�B�#��yAV]�ح�����q�j[ڀ;俁�и!����.'20�5���kpx�)Wѹ>s�qI�jt��?ϛ���I9�M6���|�����u�ްq���,�=��S^Ax�0*��C�*�Cq��j��=up/��l97��w��l��K(_7%�'��Sv=��V�VK+���#X�?,D�i�"PeR*=�\x�?KWȐP�>'��H��KO�q���|�o���p�l8Uf[AԂ����e���:I�����LFN��yF�����<�5�
�<L��%9
q����r��!�u��/�];��Q<:�������Ò���J\@�Z��Vb*)��PU�Q	=���q������z��=�85oW�`yJ���R�C,��Q��Qs�� Q%n�9�U��T�r��B���V�`G�?TE���	���(?�F��F�>XN�`�3NN���;���P���])'�<F�
Y/>-PBT4���S��<)J����p��=�W��m�@��ӗ�w�(>��/�>��X�P6	�G��s��bS������U��n���Jq�́�e}�>8M�$�[%kg�^�]?I��?��A!Q�Z����ߤ�'�0�`�T�j� �\[�X�9V��r�s}2?4���f�N��C�2k���l���a1���Ő+A�w�'`k:�A���zdd�"9�$��m��k�D��w�qSR �m��ڿ�]��y�E����d����7�^w	��XZ`�	6ALe]M��?�a��vZ���l
���n���ZlA�QvnN��d�6�i�F���>�2��$���v��Z�-��~Ӥ��p���U�Y�U�Y�'��d|�� 1[�.;>_nR\w)����I={���e1h���ˀM�>/�}D��-Ǹ��4��8S�2o1:�q���^�n��w��#�O���7�	����6����I�AI�����WDệ@�"�����ZD/ܕY�V���v?t��z�)�`�����[z�����Xys���6����[5��d�MH�z�!�YiрDn�m��8"t�]i]0^|��*e���XA*X�#��a��zq��&���mG�fwd6o#'f��͔�d���|i��I�g�Mpc4�Q����(p�	
d<���'�g��1�$Џ����Ї���v���
$y��֣O�[�����n)�'���������^��1N�n=�[Tu�>�3�Cto�K�Ǆ�d�n�"�3���K*S�P4�ַ���Ð��P�M/b��Ms��,��`������5�b��w6 ���s2xM;����R�t�+yS���R�W�� ?���qF�H ��Ȉ�C�̵��(굵g����ڤ�=��(>]���a����L�'SY~�$�uxd�Э��,�$��<>EX~�>��Y����Nn�4��G�8\A���Q��AU�j����R��'���Ѡ8���h����Uj>Nc�	��iBҁ��.;r2՘P?s�/�\�D�>�u"	�t�& q(g3W���$���X~���Ȅ.���;HR
��(�u�dn0+��D-~��P�0K<0�/<cl�)�6�r�Y�0a!A��� J�V��-�6��B����uP�f-��ǟO�BK`]&;F���+P�E}w�7e��O��e�F�9���8����)�;�0X�(�	��Ă��@9|X��D	$ës��_���6
��s.���<	�bq�㻢�$���e�Bh�5���J�x%~�[�%ث��ͮ�������9GЦ�q�]�6�����3���p�_�v �(CC�[K��4������B�uU�O��n.`�'q�O��'��(�{t�D�'S��T�=�f�'CI��	z�+���$,�2g}'$5��?p���b��3�̬�}��-��e��>z"q����s��O���F�Yׅ�Y3]&���F!^i�6�'7p�Z��\?���	�g;|���><'���)0��ݞQ���;������0|�����tX����b����p2���⇆��nȊ/z5`��pCBҩj�����׺���)���<��J_�UW��H��6�׸��;�Q��Y�z9 ��y�e�GV������mS����sZ��V�$L�'**͙NB��g�A�@�+,{]�m�)v.����ma熹�����.�_�FA�D� �G�IT���D�\@�<֏�v���I��6&s{ڞc)dao�����������r*�xm{�9U5 ��6婶�\�� ��qV�bA�������1
{�Ɗt1�_���K<2�7>D�������x��;]4�Bv�_Iǯ�"��JU7(�˟J?I	��!�|V&��|��@������6IEܵ���7�	#�H��ʕXc����܊�i�Ձg��*�ɠ�ͤ��n��hQaa6�|�ph�|H��č�i�VY�:=��zz/
I���wD�zE��摓6N�h�yO_�k~�&oz!\��#�wͨ�\�}�ujm$,;��^��̢�1���Gl�?>��n�4�2�4DU}������''KQ�A�R�5�!޹�6 ��|�v��,f��@	1RRLS��=XiWh�0�뤀���X���;)�8��(��M76w����G01��t�Ŀ����*��wL�ac��������ğ�㉞�JXV��E�����6|�/V�������u�Czobn�8�yZ��o��z��6�H鏥ɍ�֤@�޳H�f�=�Q�vp�Rl@3�	� @�Ƌ�v�N��Se(X��_�ӈo���`�<�eA�&}g�`�Q/;���^I)���w�`�NLS��H����j=]^���pv��	����RrFAwO��o��dFl���!�W��}��B��=������њ<�.8;T��/���]����j�ߚ���4Y�Q\N��0����e��ĬE����xu���X�n|T%E�֤��&DÁ��(�I�=�5Q�࿂~�r^�3�2[�|x����|Y����ɛ�%��&���Ń�H�I��lF�W�~^/e�?�G�{��t��M��hx�4�ƃ�T>�nݢv[���I?�)b 
fT�|��-0+�#>{]��,��<v\�>���E_e��[d�->�̵�?��I�6l��Z3\�]ټ������)ӣx���C���&Rq�ѯ,���Z�ڐ���O�T����X��HBÇ[�{;MF ����:��B/�jc��@���˵G�\��ySė9ܾ0��&#����*���.JP�����m\凭��a�*���?�I���
E��9i��z��z�	�&8.
Ϛ�T���3�d�A���ˑ�_g�?S�yB��g�8�qm��E��������1���$S=�B�X�i�J(�YFaFޛ���yX�d���S6�i-��J���?���������Y'����	N���3�,pg$Go>»@�tҾ��w�r�P��:�ۏ~�9�άM<r���?���)��~��&ϼ�V~&EN}����+�8
�1�t�C�U!������E҂p�I�u�� �! �װ���jA$`P��f�АN�[ef��%�o�;�j^0</���k*�KCZP�n�ߗC[�i�0�����ډ%�t �J�5a��A{�OZ�'��t���Q��>��;��F�q���u1�S��l=��#o���E4�����;�'r�#R��<9\����!��	�&6ҰTa�pN�*
G�۪2ﰂ�����IȖ9�QTW
���8f�C��dX)��:Ө�/Z���ߒ�o�N���w'�����Z��f�k�\�ki���!�r&42Rw������ځ0w��1?a���
J��d�t���8�}�h+���h�S�>��WI ��u\�o���Dv�s$6�c�>$�_�(F�13�8;��H(;Q����3*��}���N�Й"N�ej�H� 1��"�� � ���gT��C�%s��.�2�nX�x�=�y�Dv��C�c�O�oz_�W��1<`��|B�>89F�LҧGR����d��B,i4��ɪGOK�㴃�]!�6<�_����LG7�GNe�wŇL�o��jS� ��*�$ع��j����-Fg�	:ŏ�M�H��l�%���EM���-�^�8�"�!���4g;MIO�������9���<\�a��B��@�Ag6L����jn`���(ۉ��մ�)�V��q�l]2W�)�kQ���dB���8�����@�O����S��TU�f��g�_B�vx?-U�2<����g�͊1�t����b-u�d6����Tu{XY��f�V���b:fH���A��𗜞ic�'jk%�#��jW%�����0D�/�Mw�l=�����İ-�⡭[�eDw���0 W���/�iB���LM�@GHje�������Ʈ�Ω���g�f
#��a�-X��h+?/GJ�6.�e�,�=����	8]l̶e	��~����vJk:���a�����+����@sP��8	����j�{�r��m��K��a��"�Z� 7�?f�p���eS����D�4�-2���.��x�3@�
Dt4�9��z���i�
A�[�{q*�W�A��8/O�	�,�f;]�6�n��w�
��v��W#2>��qrt�<�>�HG�u�a�؞�s�F�5�9���(#�RZh��:�ϫ&���?���Sߵ���v[��Ǧ���F���ذH�I���_�x��1]���6�������Q���\Z�i�������+��k�J+�W$�[G�͗hű��j�I����L�sf�k*���4h'�$0!��'m�T`C�dw�W#̈�z�K��[韡w����+�a�eܹQ�'�6iQ��P�99��g�=l�q ��1L��)�4��zm���1��:�F��uy�+�ӏE���j����Ɔ�����N����
h�yd"�ì�z5�^+v+v@�\�Q��Ȅ ����&�
蔇�����+���3�wR��u?§Ȋ!��d�6|\�23�����T������֨���kT