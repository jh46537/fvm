��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�姫�gLk'y�ЎEM�AɬA<!p�o���s�+Y>:��h�p1	�A��KM�1��ف���1��B��SS��	n��^H���nP�ˆ���/�>hAx ��לP�9��>O�/:��dD{�����H���]�}�����aѰ�n�>��#"ۃ�!^��qZ��6m��:�̾p��B�/d*���)�Ǹ�y�kz�X��ڑ�Y���R��;���ꐞ�@̀�
M���c�JFU[s��^ؔ��@+�"B|a���a�e)F�$���ROZ���,�c����}��"����M�^�*�� yء�8ѤU9��Or�M_*���5�������h�K��c��#
�Y����ڑ�nJ�,�7�f�6�zD[��n��v��ݬ���	���I���U�wȤ9�:X鸂���X���2]x���B�}F�nP7��R��Rb��X�-��Q��hP�i�E�P�E�~Ss��8N�cZ�/�;�]X��dY��>t�A���#+1�T�an$*VuEy�G�� �H5ͤ�o����Sj�6#��]��X3&]��=�F%��>���,	o�exf#ԍ9?zN���'�=�7����!�P�m���1�}�\Col3��9~Z��Vӊ��mN�ֈ8��I����MdO��'V�:�k]S�"������R�R��A���)��*v� ~��N�&�c���V̨�K�����S!�E�k�ӂ&N*Y�0"��3)@�u5#X��&��&w(r�a��	#V��v��ak��X]�l,�\�J�m�WU2t.^�-L�Rh���m��C22R���c�4��-�d-��i�ժ��߾Ay��w[�1��W�X�Ա�/~�-  ���L�:r~/�:�.hY1"�|B\ܺz����>?M�?�B����͍Z�!�EL%hݏ�\�JU��5��^���_�������G� �d�����t�P�^9��u��HA�62�ۛD8��57���"��m��  �M-$���%2�x���t����� �:=Or���Nz��?�nFgJ�?�����$N�S^	'�GDҲ-���"X)%=i��X��E@�lZ[<�J'^�V[3��vh|�ϝ� V-(�{�i�JDSmG��5�u	f��_Ad�E
J��A���w[�Q�W�b�7%������O4��J�.���<�㎒Q���T�Ԟ�:+�t�HO��DH�T7TLՒ�G
Fچ��"y�=HI9�^�q��/~�?�tf�	��.�%%ɰ����?�m�'� �s8��ݹ%���&���6��Y/�[��rKBw?� ����-p��%�^�-H����E�R�.l�]��M�iU'�i�lAu���:�1�$�@���n�A�_��>-�Y�=�5P�IOv�$�wT7���t����ȸ�	�c"�e?ލC����\r�%��ܗw!�O��cR�qN�!d֝�ϩ2�ԁ��\�N��
&;���B���0_n~:;4M�BNx���P1?�K�G�-S���k���AoI�L��C�o���~�vnY���T�$�q�:�@�s�i���Y���������y���{��l5\��K�&�-=��%>�c-�0]Z�$��i�k���9?[T>:�(���h8�u���I���{�(1l3=·�-Y�˛��[X���>���K@L�꒼KO�o�.�Kr^2�_��c)�=��]�
�2ñlb��� �\�������f�x�������I7@D
u̬QнW>̺*�a��eUt{�.8J�/O�.��4CJ�E�s��(�:�Ĉ���D��	��y��UX��,�Q��@������_�Bڀ�aӈ��֧'���ו	��� d��L��t�&6WU�R�3��V��K��N/<b��	9�q|�#����)|	��k��%�UmF �v���rN�Ō�zw=��I��W�&?y��k$G �O�u@/�Y,iQM-��Ղ\��b�Z���L�j2�R�>�:���'��s�F�|zß+�P�IK<Ug�5��S����={Uf��if�?�Z�y��2�Sen4����y���(�h�7�(������������h!�n<X%���e��3	��f�w�af���0;�O�0�R��1�g<����X�d����۠�d��PS�=�ݚ3=���wKh ������^$Ǎ�}����e�2�D4�
��%6M.�M���He�V|1]�L��g,�Z�E�ϛ8�T�.@m�0슶���,�G<���1��ױ�obR�G@�hJ�\C����#���Uۡ���w��v�A8��,���^(�5b0<1{�!j#/M�ٕ�,�x1��&ԯGw�h��J���
� �ӿ,�D�4�:�`� 	���q��!�`Fz�-�!\z�_
e��Vf,�l�[2�	,ޤ)e�Ɯx��%cs7`�n4*���HP\�	��a/ϻ�׶������g�Ά��d�t��)�@\,S{>���]�#�Dz!�z"9�nFC��Y����ɚ^kax� �S�����m@&:�K(�U���4*nFg�'�X��j��P�d
�;l���l�$�c���9;i�/c�̝�B�'�R�h�����ɞ�Jz]j2GT6-�y�z���9�CúTNS0();MH��"U�K�,b>὏�O��\s��hH���sn�?��*[<ݔR!��h���1�Q,�o�:����JaD.7M�/���"FC�}��i��h4���e�Q�W���'�=]�b �~^fy��r�_<�s"Շ��$�S�|
U��˧�XɨK7^x=n���AѮ�����y4�W>��<`! �>�OM�^�\֫�4uߊ�3ld���n5'�j���S1RB3��v\#������`�ƽ��Sn�w�\�s$]Vء�(�7�^J�{�c�IF��)�O���?V�vs���pօ���YUOX-��ى^�۷��̢�֤0u^��@���b�����嚸I���osi��Ó�I���.�@)+,��(]�\qRECP���ԓ_�Z�x�ʡ]<���p�ì��샪ս��*3���q�a�R|R��Vk��@��¦vď����F�^H�:�u�{3���I^"!D���Ї�K>z��K�<�Y`�㒮cir�7AKb]��p���4��S���}��I��N�t7�Z��?��=1�VYG�}� �Ⴛ.��(`����L��8Wm�%���L��a�F��)^7��AD�[�lZD<缃.�����ʳ�N���F��QuT?7/��Y�����DI���Gћd=G��V�Ú�Q���! ����4�՞��&k���[���[��{P��r`��ۺn*�l��]y�l��RZW��:�h���\^3��� 	�K��I�|9D�:*q�y:������f�8����Q��C��>�w�'P��B�ˠ�`G�3-7׋��X��g[P���9��J�
j�@<�d�H���(���wL���-�*C������㛿��$Ǘ�w4�����ߨd��҄j�����˸�k�o�K|����;ކ�?�=5�����c`ʲ�>�L���C��Ϝ}�z�V��\��
�_��˜[�-�a89}@�o�"'��� ���Q�]�[ּ�Y/�P!d��4Ƹ"M?��_)�^Vy���iz��q>`
�Mg�ʒ\��8���}[������pdm��$�����0��fXt��%e)�|r��IK�<��aW"�qnd�n)������.=_�H��w�}�^�z��ʏخ�r�`��
�e���J3]�.�C�?V�>��_�W)��7�����9�.c{��	��f_���֐;|Z�b�
���5F�8!?�����n�;����l+�YF�b��C��/2����7�Q>]��
�i�et���Q�色L��ѕH:�X[�M�9{�:P�(AT9�����0g�Ђ%�rSw�р曖�鹁�]�'��J(:|/I�8��U���OuR�j�L�˶�DLJl�]P����2��?�Xr�c����e���<��/^&���3��{~�h/�&����e��{3�ٍ�;w[�����I���0U�Z0�$�lz��V��	��,��D݀dd�÷�锦uLb���W�+ D�+�#����Xgϙ�G�*��6iܺ�����w���mw'����z��^�U�ޠ�(��Zƛ@w�ٍ&�U[7�u��0�M����� 	�	�ҲS���h�kl�% P�L�jP�'7	�a�'J�?2�^��
{O�ߪji+�"XR�zۡڧD�������}"7�̂�`��QK���7��	�:r�;�$��NZsq����I烢OT4��
e ��r|������IS3Flf \e)J�x;7^4"��ѵ�iң3;��~2X�ƚ��ɒb��ه��\~�{�΄8��Jhٝ^(�x�Ґ3�� ��ۂ��l��R�4��~0"���'M�8t��٢��`0��X��R��H[0i4r%j�7�eg���i9�)�����MѨa�E�_c� �'a�����D�A(RP�����o"�T�hQ�'�ʢ1(�S�n�߷IC����;����8�M�90',R��a2U���ȧ��bOV�2�y��I�1��^����_�7�%7�R���vZ�dFg�l0�l0&��b$���hEa�9_=N]�3�K��;�\aͮ.�_Ǽ�<��)_|DO~�0Y�}�e���>M�Rs_<�&�nrn�3��**��c��Օ�1��	�Es�4�<$��9&�67��6@L`_t�@��/n.���<_��	��l�B1�2�q�mؑϡB��@6dx�M	��<\ǟTltփ��L�+b�$~��d��a/�U�q�Ǯq�)#C��8	�^px�^u�Yd�ů�١Z1�{:����f唱�Ѩh�4,^w#����ՖuD�|�/�N����J��K&,U���A+�1��8�<t���cwX����'Rl卟}�A��9Р����7۸����4Q	ΛX�7T���&{��%dk�����5%��c�o��p��l�����,ٖZs��i}�H$��kmӟ�3�׊���?�.7��g`�ýЗ����y��`;��BJ7d��3�Y��G� X֯=;��
�N^�7��:R�i���`3�Ɠ��4�F}w�KY6Мm���W�{?>("l%cM����!��f\�&(΍1n���a�r`je?R�wܚ��N c���kI:��p*�5�<yD��?�	4��O	��Gk�,y�.ܬ�wm�~��r+_�D�((^f.����n�
SN�N@ a��<��V�ᐨ/K-���O��B\��E%��ǿ�j����!���(��Y�o�/��m���5�'��nJ{�W)ET�ʘ
Uk�ב��t!��<��4s!]�"�9T:�{<�^��R>�{21/�ۘ���K��͎���;f���e��I��E@�k���\�'��mu��_s��ԅ�Ms�;_��S�Ǡ�u�6��t'spn�#�nB"�h/�=�4�"	�I�o)�jK2]�Q�*�Aϫb�~�Q��h����fUr�Y�p7���t� ;�m>�\zc�s��Y��?i?�~A2-~�z�S�������תP"����
��6�}�p�/�:�Z=n��X�~��;�O�����ߪ͖C˘�����M?7�'�-�Et h�ͽr��c�9 ��+ÙHi;��t�94��w�Y���sȞ%�%X�΋�u����SH,ϲE�����[7�W���˫ze�殺�5$6	)�*ۃi_2#��z���_�D� �����[%���D�n��ހ��pV�R�aF�Y���k,�l�o��]��v�Wq�i�H�J9Ѻ~��??�8��*�Wv2Y(���N��wŇ.uL�6{@�A�w�c<t@���ہ�f�L!$��V�B��]���mpɬ��x�I�z�h6�5�b`�rK��,Y�\�Bx�вf�s��~ѪsA���d��W�Xy8qG}�T�]{�>����V'"��M��%��y�s�j�d�m�W���קs|t5�ٱ>5��"��j���T_k��\��ԼtV�	�e��'�}s�?�Z䔷������M�"�`���2�Y���b�c���6�)p�0��tٰ�+�zGx	-5�")��|ߝ��R���d�E�i�f`�t�Ϟ�=~n֐�Ϩ�u?�@��$�����۟@-&������\
�H���Z�	p���L���_�䡪8p������5�}�/_��|�C�[u����ټ�aaG���р>_r�>�>M7?��x��
rC�� �Ę�C 22��~gWϏ�y�P��D�y��ez�K��O̓!Ǽ��>�MG8%�l��ܳ"sw����tP�5��W�?s�z.�
���<�K��u"��h�����[[�E�������`��6nwʨU��-�7�,�А+T&�}b
���۠s�ʽ:D�H���-���p^	�1&���S
�6�� ��ߓ�Wz�M�KYA��g�h5��ڋ�\_d��W�_�g�RF�4�/3!��]fX
P�F�KYf�b�g�����0�����m7�܄�i�0��ŰS_�Њ*R��d�3�����R�gB&��U���Kީ1�;%pR�oW�p�;�nQ��O1]�؝i���xԀ��v�`k/�4 h��a�k���C�n��#�"çG/�� '�M=b�m�D]��|����
^�r��yet�9��"���iEEԍ� %ՙ���lg���Q�K������_�(?r��!>^��
�:�rv�ai�͘��W@�f�d\��������j��_ՠ|L�vU}SjJw��w����gj�T�^1$T�wL�
��ө�^�>�'�8d��#a��v;+0�����ve�᝖��	��8L�d���̴ȋ�9,��d�Q`�����`��+�1	m�P�����Yu���K���T{�v���c,��㐕��%b���>b_����9cҀ�8�WV`Y*Gj�c9�3�޸Mep#�wk�%v׼�\�b`a5
�����AB�'�8m��`��~�Y���џ�5�+�����a=�c��'�Pwg�Y�A%�~25[l&��S���kwG�����^Hn�h���2|㌭�%#��H3'�������b��G
�wф4�ߜڤ�_J�iK~c*/�L�
�^�3d]��q]W����\�n쿛�����5T�D�V`��b���z1*��wA��� g���ZO8�������W�5ɥ���6�L;H��ʾ�pH��mYУ�ʔ[P��E�~��$��7Y�o�����N����9m�����O���~�����+�;nV��P�D4�ry=<΢�a��H�a*Q��$�
(#W�hTAJ��������)�x�ɍ
ٯpD����G۲�V�y��4���d"<�:�����*X�8�C]��}J�u�;U	�S�$,��2��(Ri�u��q���i`A����H���̈��XK7�炻����o�Ѥ��V�~0ߠR.��� FG��Ԇ�Ux���{_��I-l"��R����9�`|� ��)xÑ��d8�  ���?B��x�#l3`XW�X������ū�_�d��&��#�P �__�`����Cz��m���6�0�"�3W�w��ܹӵ�!E��.?�����A���.��6d#���<~��M�v�[���J���K�z ͣ!W�&Oh"�D���ӭ�J_��Rõ1���D1X��H������K����+.V����Gbx���/[ݾ����"J=l���W�D\	���8Mt/���1��s�ZJ@jE��"
�ui�1�4�(�[�Wc,�:�����ԊW��S�1��_$��Io��f��9�KH�Cن�Z~��x*�Ӗ���;{
�#�_��5�����|*��ǡS\M�^D�b�+�U���J�I�M��������J��f�Hl9/dm�K�.��"�á���
�Wɺ:���-�.D���y�,L��|o4��=�hUg�
��˵�4���qxD��}�!]e$��R#���-;TA:��.)�(��+��l;?�w54/u���		:�}g��=�W�΃L�YE�S9�?���	�byY�����5���*�n�5�^Q(|�m���4!�9��>������Ŏ���47l0*�+�*�c��CcX����o �g�](�"����_e��ʙ�Կ�t���Hu���>��}�R�G��,&��s��C�NH ��rtmbU;	�������C�K�iZ��U܏TFh��C��"'ak|�?!� ���4Î�*А~0c�3B�c���݂�i�iI���L�y㤳4��k"R4S}���c�w�O;P�n�#�yv<�Ѝ��{E���&�E�y�~�B:Bu ��bC��7̈́�zk�Ӝ���aca]�s�2�
\s�
�{��C�m�E�Vx��S���sڽ�I�](���K>#���%0d��K����6��/�0=z�~��^�����i������p�����B�}_�)/���}�$mcm�/+����"WI��Y/���1
c��M���0�Ȫ�E�~QpW��Қٮ!C#<���E�{r���@�9Z�A��;�<��:4�M�{��56o�ɔ�[�*�ϊ��jJY�!�ˢ�qa���]��P��j�U�1��Ň�������&�D���m�SV�u�� ����b�����)&�Q����^�@A�*�k�R�R.
l�����8��V�ń��l>��S�u��e'��"�Zw�n�[�zۻ���zi��}��d��ݱzy`~|9�"�|Ws�>g���~o��4+�N��M�EHX���(���4�_C��r���GI���
��8�v3��l2����@��!l7�K�:2����G�?��K=]���Q��("a������u�&<�U���c�i����I#K�p�d|���5)��`c$DT�Zy�5�m���by*v\9f{���%�[�"�o���S�0;�7e���?H��PLr3rV:'?5
�膑�[0�{Q$�7=I��1&�v�xf_�J)�L5i���NH���gf�8�U��a7�H�����D�@t�<�Q=�j�S�z�̋�x�ٌ��,�x��j,��Q���/��Z�����\��e�d�����x%�!���R�[!"@%��wk�,��i	y����ˤ��odR��X�9��!h��������A��!.)�u!����u��3���y�����Շ�����w/N0L��[��8L�^G1xP{�1��%�M�+ʧ!z�		xň�J�	q�@v����F����ߓ��o���p�a�}�8�).�\P:8������4�c����d��K���b[/%�7���AJ�z*�o0��H]�n����)��BC�h�E�c�A��q&�{����:�d:�L��_8W���� ��Y��r_tU�9�PdlL���(3�f_�7 �������vZ���m��J������E�x�n��;���A��Fà���G������|�8�3>�ӿz��
}�"���XH���T�'k:jB��Ƀ-fp�V��t�b}��?���||� �H4d`����5��#��K��"��x�T���j����ǭ��/{�g��5�����1*W�	$r��bWf<�r��Y�Ź�[�zs1= t��� _�\?���1�Xo�W Z��h �Jg-�XX�a�zx�]�Ԏ<9����ZQI��	J�j��7�>0w���F�b��3$�?��9�2�o��q3�W�&��D3"<ح���j��hgj?*(E��y���	+�#������S��>Ƭ�^M5��-'U���8�e���b�[)<�ȧBwi�~N�ZLq\e��܊`)��D~d�8 :X��4��X�n�I����\���`G:O7Fr�kU���R ���� b!�.��V��Q5<]V��3�;"�{��A.���~M*��4��3t>l9�-|ό�����Xobq���;��S�A,Z��Iد(�L�������8w������"�80G���S��?�����w!4R��3�Y �E]߮I����_�-	�K	<�Ii��PM En����'�{e����v�4l,�'#�]y�w0aUB)iLbd-�2;O�3��?L�ܛ�I���^vd�����;����8Xᓃ
d���-Z~9��G�a��N�O̚��+���u0���@�7# ��]g�n�)[���vBU�̂�����:�	K="�*����F����?�OU�\
�W�eE~Jb����N�'R7�;f����DE��&�X�s\��[��O߇Y1���K� b3�D��"(f����6��pl����6=�n��,��O�Z��K#��%�ps�B"7{�I[j���Η�G;�xaޥ@��O��V>ۭ�7Ú�ޕ�}8�@GH�(��^�����MЇ9���B �ǲR�HX3���bI���?c6f?��A-���.N�5����[��g��	��sO[z<}[t���8�ܡ	q���>��F-7C����s5U\�o��� �.�G�B�PGŨ�;J[E�+=��#?Į�H���%*��a�_f��!��)6���1ͦ�hȡ���w����[�N�M��.����I��Lr)���g_k���6��S���X�)�;���)4���j�@P�j�oxd�^�^Q=Q^EU[YI/W�e"R��J��G��t(J�vV��|^���ch#5����-���E�6ɴ�K��p����n�G���In��×(��;r�V�/;Ԗ�o^���ÕQK��7Q�&ćn׬�����rv��4ׯ;��q\� �	�ޖ�d��4?`�kϪ�ť�P'ѱZ?.���?��r�GO���[p,OC*��#mi<���<⩃�@X�5�[ z*阝Te�ǏqT1�t
��F��ť f��A� ��0�#��0$�I�)�A/�S� .��j�3z8E��ρ�k�qzx*쌚K�1ʠ;.�,��5�!o/;w&�m�Xu�ɚ�Z���z-�+a`�=>��d,��y�ly/?��ȊS��r(��k"Z�x4��u^�u�KW�8�q�)�~��^gt&UTi�����A}n#np�
OsEl%l5��G��[v��#��:�Ӓ&�>�NiN2h2 ���1ЩX5WQ�\,2+ �hw����	,ɹoÌ>.��zp�#��3�0� *�o0�͠�5�zJD��W 3@�ؤӰ��R�.
���7�]���۽02,���N$wOZH;�/Z���dK�+ӞZ�� #�����D�E�A
��/oNR��lz�>bd%|��Ǟُ��I8Qy�D�o�~��H~�c
�ȃ���nM��0�#��R>.�<�����طa���(��o��#�r�,x��cy�
%���۴�e�N7\8�1�R}|3��\�������v�m���Up��C�$������h�����>t���]n�i���n�v���ՄA�V6e��7�@���j&���!�)��Ӛ���P9�9��h�賌9�����A�;��i-.'1_ԃWA���f7}��ꋬ�E�>�9��;#�v�d�E�8J�;U����0^�
:�v�]�	>�9'�ܾ�Ov����A��joO�>po�w�+u�M֔eZ��ƍ2'����²!T:��#\cʬ��� ��߆|�Xe�^��Rdּ���qj���.�{D��w�XL��y@�b�v���\��l�Y�O�|�3����I�t� �~�� ��W�;~��}�؍Bz��')ؕ�Ή��$S��\6<#����ur��i�ށج�����*�c���#�����V�	8��V�����R��q$��+�{֍,ٴ����b��`���m���7`^wm~�Xp�B�"����Ç��`RṔ�/xIı�z
�-��ۧ��Ӆ�'8�Fs�@?��9��	��:�B��������U<���w��p<a�>�B��q�U�QP/�/�葭�S1F�ǐ1�P��U�^��$Pm���Y��ǁ�/�YJ��K��p��s�3�`.�tĉMg��"H�C�(�7�5�?��Ѝ��M�}o+.�j(ݾ!?�s���~��n��O,��yd�g� K���r҅�zB�����Ě�2�E�
�������-+4��#]Ѫ�uLsk��;EHَӴwÿS�cT�oǠ��y��e�I!�1�1iK������D��l�_p�?z���F�8�C�~�7��0��~0n��.����v+F"��D!���3����1�f�̇�S�Qq��[RN�oّ�R� �~@]X�QR�C�1@�J�,|���T7\1ǿK������H�b�S[��[�U���(Z��Edxm�$�~���K��s�D�:�v�"6��˔T���"�s���=K;(C�9�ƭO��r<bJ"��X�҅�&\̛9�W�y4��i79C�= �y˰3�8�����r�et�_�я�с2t�ʝ0��uw��si���_�{|��n�`)L����[��[7����G��o�6��L�Lđm����(��{�5ibeF���WE�Jp�[K��Ԑ�*d(�F�р��1x�W�O��w��_��͌��2F)���:B�"���1q�L��͒~c"q�L �6g��5��m�u@�_}��(e7c�Ӻ2e����i6�"��8��m泏�r�\l��Ũ94l0����ɠ*�jY8�����g�|`hU�K����Ҵt}?zl�f��x�TdOe�ݢ�Qk�����'Y�U�ǝ�6y��x����yV����e��=��2�LX�U@�#i8�J>sUF��I�UF����.mW1p�F�9���A|�����Ѐ��3w'�3���RN5��φG����厵�Fm�"���p�Q���(�̋�w!���I­5zH��k��M�͐'&s��7�ڳ�މ�L� �o��i���TT�W��ˣ�ֹ����m��Mμh��~=�=�?���A���~x��i��%�K�⨸?�>�Ϩ��Gt�?��	����^ 	W.	ɸAK�]*u
BZ��5��r�s�o�b	����)&��fr��kJ��?-��E�Vt�s5�K���wb�
��g�����'�y�1e`��="|�|�?�5C\?!� [��+7k�Y�+�i��#��=!��i�˸�c^@a�C�v��H�j*5��p��Y��r�B������&�$�t�-T ����gs�wap愇��;���RX�'M?�)�炠�5��s w�=+�����5�P͙�p����{r��n��"�#v�7���(������JR�a\�,������S�oG��:[�)�f2՞��W�w!u*L�_aɶcS=Hb���[���I2R1Lĵ�_z�61`-�D�_;b�1`	I[��x�ຳ��8�<m�,��o���/��6�E���ߜ�.��6ٰ�bn��x�>V�zucц8���[R Ķ���x�#�M�+��X"�����������n����}Cq��Lv��AX?Ɋ��Tx�V�r�w=�Q���;`@%�=}��_7.�DNBӃϨ���R�[t�r��K�U��=T���50���b�?#[��?��W_e�G�J��Y�W��)r��Qh�*��S�6�j��b9+��\�/�.T乞P��7����_��R-��3µPɃS�B��</�����d뗩YC�N8��"8�ಿ�5��[E���]�GiDx��\�햧�N��0�(�y���Mr(. �o�"}g���"v�I��wj^�
q�ԙ�n�c],�wv��F(�iB��ݥ�4��
I��؈�v[��@���"�'r�,���E��S���Ic�
�m�*���yw����*��J$�F��M�	?�Y>d=�]�rd�p�k��N�QPh�,[���j\�_�l��4�=�K�X��cH\�ǌ�0=�@����!��`Q��H�q��`����b��GP驍I���1�?�H���D�b҂��C����F��lK~����?WP|��9�5���fii�n�&Ѧ)Ӹ�љ�ɸ�B�{�KN����B����"� u}�Ju�F$]x>P{��?�jtR�a$�lе?�f�����2�FST,z�����y����H>c�B��7��`��M�%M�NW�]ŲΏM������ĳ�����|=q���
 ��)����H1�C�Ht��sD�R�Ē�n�E"��:�-�����*7��-C} *�,n�9us�2�#�q��ȱ'��o�6�m�K�P�չ9M(��lT.Zr^�"J�s�$�t�D�c:� y����Wp����X��$�2̐JM�n��V�o����1.�U\��g2<�M	��Y,�D��"��z禊.A{wi:S�}� (�*^be���v�12L�Yg���)����u�W��F�����k$����gݜ��A],:�)�"F�E�M�KZ8��5�C��Q�\��;)�Z�VH/��6d�����
�kSP�\�1[N����B�g �u���!��(q�}��#_QZ1A�~��2�d8��+r����T��qP�"����!�Ys!�	�6s�u�0����j��l6zQ �����`�\o�-D�P��Gpn><5r�� g��(	�|�ߎ4�>ſǁ��i���gq�v��{��Ruy&ސj��7���K��$�L��kfd,�`�