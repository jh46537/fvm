��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{�ףe��	�A`������I���;���a��5j3�LkW^|�y�]���tZ:�$]]�jvg�g^�`/@v��ֿX"����<��JfE���ɅJ��CΕ�H�����{�q�d?��ą9�KIYCc�0�C2�dl�$x�co�e�R��!��ӶU��-�ĉC
ͣ�2-��Ě�5ps
�ӣ�,.n��z��N���A�ç���ˍq�����o�.A�7��w>x2bW�)@�_1��[Wk��O����4i�������h�s��VV��<���$ �6-4#P����r�7�/�
�B�+�媉�{|K�ݴ5MQ%�1��֕�R�"�����tq0���{���ݜO)���}��D_��֍F�*jP�*��g��5M��N��jb������NE4q#��+'kb]d)��~�7CXJ00�{��1�F�M��!;-W��=���d�]w�/��dmg�ǩC��C����$��6��G���_�b��<i�?�~��M�U3Du!�K�.}HP���F��M%"�\)�4q�	���]�5���#sP��Yd)���� �łF]��͸���7�5 5���BEưz{	E5c�?��X1<��U\TL��	�F/��q㡧r=��'�y�{�����e8%|˺�^���>�9vȼ%���<7	�"a�q��.�>Ái�%�|�g,��iq��^��+ۑ��:�����������w"�9P~mIR�F��j�-�a5��֨t�!�R�e������uM}  �w����w����7�ʕ�&:�;ĭыʛ7��Fs�\#�|�~�$R:�:�x?R�1Q#E��fxS�I����hx�D*�.�q�ղ�"�j4�ϐK-ټ�ʥe��=J���[r�z}>v�|�����@��>OZ�b>��X�~�T�;��!��0x�k,���) �Z�@7>�o�.����s��{t���׊��lvx&�����z�/Y�p�]j���$��X!���9��\��Y���)P7Pvr�	�����*���	
�Iom?ǩ�����כv$k:�W����2��Ib;��'+yQ�*I�Md���֖�c9��1a+�OE��%��b��IN�������#�������8�>xh���z�D>[�b\�R|(MBg�߶�Nb�*)���s�Li"^`���́'�!oz����L�Sᨊ��~	2��ow��Ь8�/6h�Sb��ϱ#�C�׵6/�+��S�|@�ae����q���4��!�v�oꭊ��$r���:�?���o�Y��cy��ˑ��k�(���?c��%�s�4����:�'����|����4�xq�[�#��;����=uW+�㧻ߘCPb����7Ul��M7�*��A�V$�1�bJ��ݧ���g�s��+"��	�?�<�̸��_i�'M�lrr���5l0ތ��d���׸��,>W+g�u�gvn�c�_�g��R쉙��W,׶h��ЮQ���D����3���+L`����͜��5�o����,��zߋ,��!�o�'[�NC��Z�z�'���`�7	i�?l-��#U]�0�-� �ݤ��Mb%CȒ��`�: !e�Z�PMl3���^�N�g�B��;m���"5���C�p�����v9\�?�nQ7�4�i�F�J4��]ܳ��Nj��L:���_u���F@� �QV�w(�&�=5�[S�^��<nM��#c��JO�4��5@����͚�(J�f�T�9:)�7g�`�V�l>�6+CB��]��@*Ǉ6@�W����P�4�sրa]}ph[/��/�a�0F�qJ�������+nIM%�kh��9���#@D��\��O�t�bo��j�8����VD���-Ӭ��D��"P#~����?�D{����2ΘK������HI5w吅�N\O�̐���>4XvF�q'L���\ʾ`�>��jZ@iCN<�*P���+�wf��b�z_"^�4����s�~�ڎ�<���"�;K���6
���#�Je;�
b���Z@�o<�s|�7�(G��Og����Y%H��n��D��Ya'�s�K�P2������ޠ��@���a.��f9(B��9/�F,