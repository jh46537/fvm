��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<?';S2s"|������,M6�L�C=�d"�a�NP�f�l�͕��a�!*�M)\_��d���kC!��-L�1X1-����7�L3	o�h�:ϑ}+��Gv$Gi
�T6�;��f�V%'����0�I��9�ߓ���:�f~�k#��8��j�+;x�wlc�z�v�k<D�c[k�����S��oX<��-�m���ӱ!l%����!"g#�i�������I����K�u��D��@�&�Dr?Z���t�}���#�&K��.�X=>X��Sf�E�\�v%�L�B�BlMLY��,�dr09Z�X�̳�ɧ��\�KOAYP�O��:)������N���.��b��=v5�sjsg�ػ�]\���c�2h�8#NE
!*�P \�'����v|��d_�y���o��y�e4�Q��S&s�.|�t���?��Ŕ����Bc���g�P�qb��,����qy�����$�������P��������R���؎�2e�=���:Ĭ�;��
]�!���OV_�JcO�瑡�=��w�{������s��<�������fd�뾉t��"M��ú.�����g
E�8uc�,��e��!�nu7n��o�i�j�ܨ#�K01z#��9�a��c��q([��k��j>St��o�E o��S*�r~Q����AE��V�������Чh�)�i��l|�pܽ�wJl+p�@��$>k�<�A������z��k�V�VO�����Iq��R )D}T�^v}AG�8�߅y��4���qLϠh�
�:��i't�5�
;��?��T�]����$3F<&�۪���W�B��	r��oŞ�������������s�op��7d|m��|,	v�\��I����4�8;��%�`�l�r���1��}>Y�|�?��I{��Th��dd6$���ތrU�}W�,��V�wh[����B�.���%����� ��;�3rk:��͋D/�D*Z��0
�b�	�
g'W��i����:���H��M��b[�Q�r̨b:Ǽ��+�Y����wW�ME��0�U�)�A����*���XX�Y2��������[h�l��jT�*$� SSՑN�fm��#7�6��s���b�9�ʲ��C�BM�S㧀��M��:3-X�FX�(Й�^j�,����ƞ��Y�'_�-���kd�w�������Q�nu�a����=tfJ� d�>S!�����lʡwZr��H��+bp&�ŉޮ�4pѬ�Ψ7Q��`�`��rT�%'}��hw�ʨ ����'`]K�e�.[����1:��eɉO+���3�-�V���
����-����������q�(��Y)�fhD�+D� �Q�D���Y�:�l�ZSly>|XΥC�Yj��&܈��W�M#{���&,`�;����{;��~�+���-W���KZ��K�h�2eHn�N�r"�3Z�
��%"�ש��zoP����k!�[D��	��O�Cuy[��A�q?��^�~��mn�y81���� ��q.lW`�_X�nX��;V�~�v��sukH4Tȣ�O�Gj8Y5����b��.�]��ۀ��u]G�:�M5��j�O��0{�"Hl�Zv9��Q���%H&�5�q�e��e�A��J�B-=��uF���z)hb�%�����ܲ��4/�$r
wr�F�����}V�\�ήT�ܚ������]m�m6�sgy��s��) �&`���bO@�8�Π֩\��k� � �Y�B�j��eI�u�4s=�����;�������e!>��VE�9 Ē�\�٫�s��1���>�����*�xB�̚)����Q�����<����_�Q�+��z��C��Ԏ��.,�?T�КZ�����ܾ�߸w��ܖ�<sU�@	o�]�_x Nt䏅��ѧt��yI	�,d�I��^HyB&���}�Z/�1�V�U�H�t`��Ob^�nK�w~`��t��i6��JƏ�ja{N
���;���p�nR�A�c�PI��:G��&�U7���X�-�2ꊢ��t�+a-�fK�.Ϋ�QO''i�pP0���Ŵ]X�G6��o��5�=��X�X��-@L��j/萺&o����I�����
9�XZ�+����$'�
��KΉ�M�t��!y\Ę�z� �b��!��o%�\'>����ٵ7MTt0O�r�@���rpCi�/�xǃ6>�Bk{i)~�� ��>'�VM(AX�%�	����^si�ķ�F�Q���hR#!���Z��� ��N���8���Sm3k�M�'��/-���^�T����j�kFj�� s�tR��k�Z0m'~�'
��G�H)�^�����^)�UH�vs~�,P��x�a�Ƽ�N�r)�
]9Y���,�1ry`��Y�K>7�Nu��Nq�s� ��Qc:��h�\��j�:�P��.a�g	B�7I���a��f���!a���~���&ſ�����na�ê�uy<�|��it�^�����5�N��v���|ԟ�^��b�CZ!�IO,i�hM�W,.��ZϷxIm	6�ehsE���OY��d�^��+dv�6�{�G���i�Ǉ`�ūC}w����@[���o��"f( ��z��3���𣠤8f���'�C� �ho��!*tM�RX��b��$�,_�h&�O
�#���Y�1�Q8A+�k���9�7�*��j���+tFK0"������GqpO'��y��I��c�kn�>sI���~�XYrv5,Hl�%�Xi�o�LC>w�}�Zi�g�{ij�}5X���K{\yrؔ�t��u`)W��>�
��oՁ�W�\��_u��fE�^W�uP�;�2�JՔ��w�,�Z��)�7Ig<ɳ�>$ǀmQqax�i���/L=[d��>��-r�����~�L�.�e�t�����]S�3�7Vg��n��Mk�x���$�v?6���L8{����DԢtSo�J�H�#�%l�F����ޏH׻�gK͌�����]���"�<�=�3h�^al@�-6�%u��뛦8�@�:b&,�����oz
0t��#��t��kO�s{pQ��"��D�k$��!w궬u�D�PЎR&���޾�>W�B�`�q�xJ