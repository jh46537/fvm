��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xMMh0n��f���X�h�ʨ���H�P�e�Iܷ �>Z{�&���|�w 0B9�ԙ��w�'���,[��?�3��,5��~��1o&��VR�6�Dμ�)��Si/�#�LrK6�҉c.ĺ,�2�z�=�:0Bߟc�1^['N�8��,H���S�|���^`���p�y� �1��j�2��j�!N�҂�(�m�*�cU��,�l�MR��� ��a��#$�����)C6��^��N��T�"JQ�;wt��H�q�'��z5�6��__8d��B߮�Ę�Y,�Aq��Mc8���!�B����u��G����]5����Ċ��^�u�D�>�"
2;P���3�,Sy��r�j4�־�1e����>Ga�-9�`��b�1U���+o��¢Y&ͬ��`�X��B�U��w��h9�+=��|G&G���l1C��H����iA����b"��5T�DS �L\Uc��|h��96	~��s�RlE��ᦢ��𢕴��n
���#���Mۗ5:��3A�R�A/ۨC?/F�X�Ճ"_2� Z�5���&{	����,G�νHVs�"JG��y������&�ń� �X�B�\��AN8bk��a�����Y_JXИQ0G�?��6_;�s����\�-+6�}s�o�z�����K~P�����
��{���UMb�ҘαY����H�%��"��~i�l��[|�wI� T���/���rs��u�V&�h�ߥM/J�}�bޗk�=@CX�@	��J%����F?_n�A���tt���ZƠ�[�vGg��À�w-��R���/��x@ �0�Hg#U�*����c�L�U�Vi<q�ŰFA���xX�j���.hUs����5�zVk���7+�deㆶ���pg��2l|P�1�����G�XXX�:�G���
�W
���	�aS@�V��=��Т`�ݞö�U�b�ID�>��'!h�݇�~���Z+�w��c�A׫��)�����M���[S���Zk�c_~�c�g�������+�ƫ'S��*ܨ&��2렿xG�	e��H5J�JJW5��S8??��b3������"�O�W<R!�u�1��Q�V�aq�?I�h*uuBP�JuO>���?�@�B�K��B�Kpa���$?Ƴ��	�� ��䦲�O��7�*~����-? �ѕ{v�YRc�řa�9ϦU)*�O\�:��t�8���G:�'�	I5R�^QVg���&@3m��������b2A����$�k퀍
�?�1	�"� �ڛO"� ����Q�?���Y����e+@���H@tp�X��I��*:��a]%3t&����*������E<��I��Mv����o�W�_��u��Nh��2�GR�v\Q}`A���6�(��:ȷ�u�5�k�'�K9[`��-}��@v?_/y&g[1����ΨЦ~b �P�qS��H���&����]K�����z^�K�?M;��3
L"E=�����Ų���3��G>٠X���|[i]~rw��?�پI��M��й*U�hb���H��ԻCmx؟�/Z�"i�"�<�IӪxf�Q>==+�S3qy��ME�b���e-���e��/��H�4���e\�e�~ļ9�3=7��#5Á�k������T(�"�r)3��Q_����5w�{��1�m