��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>����rhhm���%�ñ��\X}"y�GM8�,�eP��:h�Z�{|��L�~�t ,������DN�F�	�:j-��u*�zn���{�h^���C��zlC�Wg1MH����{[�rx&R�+0,@Q:/��ц�?yU��g_b��1���C��M����훅�[�>F�?X�	��ϟ�]w&A���E t��/y[�x�b���튟Y}
�]�w3cGTe�����F;;�A���|-�¤��^�{�w\e�+����"-�v�E�`iӆH��n1��Z���Z"9߸���֦�}Q^�t%��$w��=6�e�C�?'G;n�F� O�9�Y�,Q���X^��"�p�񔺖�3ЄQ���W*�'0J��kq���>|6d$j���V�+�{��Yf[�( ���_��qd�pY�o�4�8h� 
��ɴ884�|�?�f�j�T���� �=��m�?5�y���=Ք)&��=�8m����,c^���N�f���~D0�	_�W2�� :��o�$��&t⫘TV�jXN�ߓ�.��G~��E�� �h��0�Oٍ+���<�aV+!����	D���5�N5a�L�y�<�H0�݇(�X3�����=�y*~ƞ��o�Dj�uxSVӲI:ot�?Ԭi;D��9�uԛC@�$�����ٔ��o(�
a����5�bu��N8�^�M��Y�b�սU��d��5q��խXݑ��ni�r�%./�|s�T5?�-�b�F迗s��(�L9�O)��d���TM���9��2ı�4�a y� b	A5�$T�%�E�[��6��^u_N�H��e���ګs�4�n \��Y|�%�˫b��`(��!���C�8��Cy��4k���n��c�I�d:���P��JM�O��Ss���@!���p�A�ZfK	M������[3��/���}Ğ�mI4�>;�XT���G�8%Ih�@<-):GWb���F3:<� �����{��Y��'�>T� �V��b��r�=�j�t�Dq?(��d;Ec�y��5�#��c�d���n|�|�^�6�E�x���b���Ѧ����]o6���^Up՜����Nq�ɘ��-�����e]���O���Z�>o8�R�'��[�(\U����͂89��fkw�E���13���<��1qx�����:Rfz�u���@�g�΀�wV"[Z���`�~^�������	j]>w���Bf���E�#�fk�ض�U�*||��'�q!JZ"�n>�^�s~k�W���C�HO�h���d��(5���o���<ن��DU*�˥�q�q���qvk�M�U�se�2L|�U�ϐ���|!��
`�"ð޼ۚ�iM��\����M�o������8_�h�FaX0	�X�o�wP ܆��#����2�J���Q�����ZcA�.�1u+{A&/UM)�詆�Q�̦�pnִB��h�-"k�2.���/��j�G�ޏ�zra2�?d{iΨmc/Aw':���jR�{��!w
��~����~@G�7L�:޵���^(�4O1�5�l�<y���9�&��++��k�:��s~���z�RJ�z-�_|��?�37⯭��.��]��k=�! ?���}R5BFH5E����
J �HfH�?��r:-UM��.��=�`$��sB?��������PrW�.I.��rJ���Ŭ�.�⠝؁\^2���H��7���7�H�'繒��DƜצxzZ����8!E�I�3��k���Hy�\��<å�/:a��1E�s�\7��i�/�a�ؽ�<bqH�b��鋔�%��t㢼<$�vW{��^s�����IDd��m�9>�ق���d��U=J{)��'y��bf���*r�j+�A��BIx�܎xE?H;����&1-Ub,o��!�^�h�|0�ڹ�(�v�B�`�s(�K�;v��������O��Ǹ�����
��O���r�og�$��fK���V�h]c��#��4_qT��J�_�k[�˵�f��R:i��� '0��n�ķmv�������D��/*�hQ�6?��|�0�,�"�f���^GE�*#H���`/�������Ùrơ����ɭ���a4u|?տ���&{�
�j
&I�,��
^W��zɲi�@:̤����*<� �Ëi�t����/�;N��Q$�LR��0D˚�Z˴T�$,�k<ǯYIW�uN��!�����F[��Ms�	_��5[J�h��&1�n�Xm:���K�8L'\Q��j��=��0uLPR�G��B;�R���/7#�������s��[	���$d�hY���(~�������H�6k�o�4���JI&cX����p2�%��i��:=@@xꐧ��Q0�B��v	
�J�9�o�;v�8Zsғi�n'�{]�;�S�X����α �6�:B�]�+v"��kͯ�z��\�l�D̒@Y�U$T�>xZ�|�lP�u�X�P�WT���'\S��+�#F�4����v�}q���h�F��ݤ��Ɨw�\��%��ŠTsC4�q���N����Z�^��]M��Q�i��T�����CZm���IRs�Ŏ;ՠ��	->��]
[����I��#*uj��Ns7�����AkQ� �=�><��=��vU�3>�F���c�@�j�M�ٰqp��9p��!I�e=�XK#��q!0��N�$'V|J�_k6�@y��ݾ�9���1�Ŏ�")B��_��cܷЄ��ϫ���U��|���~>X}���Ʉq\��yn�9�Y�����\�N!��dv'Đn�[U¿���on�����-H�#�{�eV"��u'�4�w��g0Ȓ�Q��9�Ÿ��W�մ<w�
���~ø���?�pyX�?���-"�Pz�����cR�1����E�Q��d���=P�P��|a-�������A1�;:U�E��
�}�4��҃"1�e;un���I��(����zh��V��񯥴I�\ZUծ��io�å,V�Dw��F��o�Fk��3�nGS�eʻ��������t�PZ�W�����8�߼�֯X�ʟ�ݿx��"G�-�l�Dg�9��⊸.C��n�`�{�Ak�]���:ci(*BQGv:r��Wz�Iw�La��s��xn�h�SO4EE��Ba)qM�-9��Y�K�63�c	~R���1�4��3�kWf3��W���{���j;�]�w���l$E٪�{t�ĳ��1�}Iˤ����Ӷ�t����FU�u�Y�}�����.V*�{��­��ke�RG&(�� �����8j�Z�-�RT*V^{��_�DV`�v2��G�n��2�=�(3T�"�M`?����`�?�0�i�o���z�ufS�.E���l���e���w�Jg�뤄��8ˌ�j1@l[�����gۄrt7.�h%q��eʸ��z���Ж��*�"�_aM�P�E��M��R�9�?�`R�`��{��+���J�h6�T����Lm�u����>e��>�	��m3�"Ő6������K�ۡ� �> �q5H�"�����礢�DrV?-�rz� )o�����U��1��櫤#�GQ��N*��==.Y��W����{��9�_v��!&��Mw�M�IU{�&�A �/G��eP�Ρd�bp���g�(�0��������ÄuU:��2a��"?"=�`%�֍��y�sa����#���6�P�.��\�����JZ��tt�w_�c�W�ۑ=N���Yܰk�9ڮ�ˏz5�LJ�d{Һ�x��m���ဈ�ӒzR��++z:�E��~���*�!���h���a���znNM�z�p���D��4�r��iAk����,�~��&��|Ɂ�x��Kc�o�t�@�ٙ�jK���>G2��\�'�w���EA��5��%l��'n���hE�X#n�h��AR}����ɏ14i&U��-.U�'������#ݑ��7�J:n�/K�{���<K��h��5O�-�=a��I�O���4`fϋ�Rѱ[{#|w?	}P`27)�B��3
V��#L���UM�x0�iRCYI�b�%<,,:lWu��b\�&��Ҁ��axף�7,=�5A��Y�v�#��G�T�]�[��5�7�ۗ��׾q�F:I�K��c�l�M����.!�ḳ�'��\3Xy��V�q�p�'���<I"fl���> �3x�o©�}�<��������Բ�sؼ��M���iQ�e��.�;}�$�^�J�]��P��s	�P�����$�d6m�=��n�Ux��V��Kj�N�e�m��q����"�#�X��*�<���D�<���G�tƺ��$bvn'��%"��l��Z~������)G|�*�i8���	#�8�i^LT�hJD��dp��m0=��p*�
U� ���{�{CY�V>S�����V�i����U���M�$货��اB���7e�	�W�׺��(��%UdvG-�

]�H쐤Y���/s�$�S����g	:��oԒA��r����="T��3�o��b��P](�Շ�4�����5�+X��՘k	MvY����)�ƅ��Z�зB�;��M�%?!�<�Κ?YN���6�i zv�=ʢ<"�q���Ec�VV�/Z$�}ӄpqAIQ��&�i��;��o�[	-5���B�3�sG�l�e�4�@n��w¤>�E��s�fG����r��
m[ʾ��6�%�`�x���9�\��ߢ1n�����[���L�A�,v<�CU�-k[�Ŋ)�=1t���5�����Q���������.�ݼ9��.ܹF���T�mߛͫz���$r��-�B��^=���v�)R%�n�D�\�R�B3�nzD�t��[Y��z�`���>�l�*���w;�5�6I?*�34�JfZ�����(�ޢ�	����: y��ac����� ��њ-��W �B�!jios�k��3����֧Eo�D�4��U�[��e���<���Jԓ��2&�6d�	��a�[�8�2�bøz����.�bj�4($b��=����O��3��FB٭�C�X����o����;!v�*% ���n	\ 3w���3?���+�4��P _Ʋ��y._D����V�����5@;��~hr�r�[�9k�}�Lǂkw��p�:<Z��	��t
Rd��-��W����r���
��_���[!�5�g�