��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	���uYC�т��dm��JP. S5&�Ac��<r�Դp������q���;�� �ґ�$Yl�JLd �9�����:���l�c��BL7�#\
*���~��rO"U�F=
R��/yF'N�t_b�u��]-R�"�;���j�q�&��i��.O�r���h��+�]��=�k�=�%�Q���6�crWNk��S.Q�RD<,T��|��"1�K���p�p���ш�Ǧ��}[��c�jw[�:a�zP �}F`Y�� �JP>���P��D:�V����R8)s��9�?��5M���?�*��a���$�*Z���1�0;cm�����st
]e�����n���;��h;-�����ف��F�+"�����c�v�,��U�F[:��A�&���
��\"��I��L���i���@kM���ۜ	]����ڣB~�S����%X���N�J�Ab�H���Y5���g��_�+���� �.�J��4Ri񛤙xO�:��q��{1r�Q�U� l%�1X�(f�n����D�״N=s����*�����]B>��f��?�fR�ZB�{1����J���1�ڭ��h�����a���1mլJPza�m��e���\e�:Gﮧ: ,����C4��"�M`Q��Y�Ƞl���K�r��帢�m9e<�bn&"��U@(��"NW��K^��[\���.�~	몷�8O��_��D3$G�V�z-�E�����T�tY�:V�7�8��̻~G�dd���e͝[���zTw��4��IS�޿ �<Y0k���l��(��}���	�WciqoM?�������NB��~�.���iT��G���=��&�?ۓ!w
snA�Ď抹�fl�Km֦xS>PW/�C!)qZc��2υ�~bC�בh�z�,���A/�S��S��������x�9]JX惡8+��6��Y�+�2(VO:>G�U��E%�9�/˲a� ��]#�A�:kÆ�cdv����GEP,�UH�Ō��2	��!W+&u+��%�����C���F�h���d�����}5[�ȁ_��L��f�� zN6��s�-&*%4x�T�6�D��Q��d�O�T������R�(�w�$x�me�/#gU�R������e�x�Ww�N��W���N~�Z��R}��x��*�/4�.���m�&�+X�B[����֚|q%r� �l�&���� �����H�S����"���M�>��P�@)8j�[�<"p=s�g*��pjQ��b;Ъn��	���ҧHF�L��N��i�=�
��#�|�.���du��\2�!a����~�+@}h�l��Ub:��߶�O�?�hu���\�����pŦ�$�A����DL_����w��(x�b��E���I����B����n�F��܉�X�Z�!wǙ�M����$N�r|�!ǆ�M?�����y�Tg��%�����K^���� �`^���(&��Q��'��ެ��pQ�h(@`�>˻?���qΰC5}{Rr�0��=�����s����:_Qm�
���}���2w��t�طݸ����7�JJF�^�Y��$�!�-#V�_�ΗUJ�HV�ՓC�����g'yN,O�O�u������I�n��Ņ[�ŏT(�� �k���L�B��;*���I��$3��	�{�߳����%����^�þ�j�-� Z.��{�1��k�.�zH:�N�yzt� ��1�����یw�m3���m�$��ľ�C��*E  .�0L�Z]�r����&�<��EH�ы�+拉��	7���Ad��m䢤���P�K7�,�0������^S���X--`u(!�W9IX��(�m�ss�H�$ݚȽ�?@�62�|B����Z�\�q0��s���{n�4M��!��*���ʕ�ǼC��P�g�3g^S<�0��yqʉ��e�ȪՍ��-��yMM��G�
��`0�g{\��uV�@
#�
�~�|B�0a�چ�$�1׬4��c[�Z�kPpS[�XP��=Pq���l`I�v�[�>=���.T���H�������Y;�����r{��숈lr^FA���գ�_ܾ[H�X�
B��ӗ�
R"7�´l��?���Z�|^EV�
� &�0(ᤝ�@\\�������������K9%*� �A�𠒪�_#�)�v:n�]�E�* ���W%�l��TH鷋;���}�_}����[᲼�Ӎ�_�옿ߵy����F�Pg����<y�K�� l-����}���UU@�.Z��M�� �Ls=��7�>=0��2}�zr�K�I�f�(H3�o�Ŧ���ȸ�ĴG/��J��DKF��Q�U5N
���J��߀�ܟX�[D����X�oWJ5��H�N�������eW���Z�=��v(˖�$���]�gB��=[%����g��i0B�m��{����v!��7m�N�+N^�䭯�N��9��ű	tս��F�q���ǘ.���E-*�r�j����<-l))ދ̎����������܂���c�L�tJq�0��_c7�'�*C�+�k,*��s����K��pO$��<��F�2Γ}h���Z��C���ʊ����W�|nE����s+x���jo���V2PP���W�(�p��vM�0ś�m��Á�M�� A�I���3�t�[�B�w���U��V�<_t���� ݣ�T"E".���1$ŸxaYk���E3��SM:�챥<���\�J��4��Q�h;*�����>D� �P5U//�C:�XJ!�c��5�6�T��{}������7��+/��[��۬������R�P��-[t&�4�/�'�1���}��}�x�^b�w7)�*�y9�������)�!�����F�yJ,4��p�w�$�)@�U�qx�ɜ�nۮi4�})���t��?��n�y�j�̾A$���1��j�w
`@�<�\e2\���Uqy�R�5\Jy��ft���ja
^o�A{�5��.�Q�{�C�fu�S�}<Z��{x��U� l���錰[�Sx~����7`�B��d � ozs�6��i��Ȫ�����Si8�E��u�/"G���/_��%��d��*��i3�%Ľ
�{��� 8K�6"]�%#E!Fʮ䉐0^Jue��h�:	j�B��?�wƛ����
Yz�����1.Ԫ��3@ԽL��ɜ�Kn�]�9P����!�P���*۰���+��2�=�C�O5�x�ӧ�(�E���֖b΅�of?�t�0U�TK&"�t<`�>{����2��lq�6�}(�HK�4�s�4���I����Ma�	d��E��zz�pB�����W������V;wьe~Pu��#��޶N2Z����?ΐbНR����iW����4�Q���}�Z��<�>�c�W��(B��y4�hUr��I��y�HZbrP{�3I����y�Z��ϴ����~��=k�wi���M�/��~0�wً�R�D�����We��$���7�i�����P���@��	�0��M���61Ҟ̋VdxJ�F����n�OU�W,���G�I����+�Ϲk�fh�K�<G�D�LI��9�2ol^T���������+�Y�`��iJp}n�xF�Ҽ*�^joE9���S�9��]1lS`��%h�`<f3��'�^V�4)�?�xw�J���+~�!�fE���Y�������|D�-*)����`+XLmEѺZ`���u �[x<i<�z�w��˖/��M�=[[Q���io�tG���q�I�	F�g��w�:+F�1����z�>��#뙧���(O�h5�{n-�����m�UxJ���cd���P�~�=��Q�����D��T�*L����,m�S����V��f����
Dt��aUCJ�s0 @=Y�,�K���,ԯb6d}�.�����D-l�" �ԡߋFe�e�:�9/s��v$��(ډ��G��[�����+�K	܁�V;����6(���_e�����ѿ�1�np����/��M{���ȓZ�T[|�n����2�['h:���o�)l�فK���B���2zg����������o�~��u����;ѯ��]��"˲�cn_�������'L�����Y(3lҽ���WE4� �� ]�|%q�h�Ԫ���F��!ZR�y@�r�*#�j,����v%�"e��=��p5K8f�x��c�
���N�d����J�`{���(�#�hxl�/n����W#��o;.�A�q�fE$uW�(���������";ē�2(���ӕ�OH}�?t�NCH)$%9@��<n�X�W�<iV���_�bq����	��i����|����h���}w}=ipm�Fߑ�5|a�����e�5�+�nX_H�((���p��^����O��Loεi��#���ڀR$���eZ'��	���C�^�7�Rb�2�b�z]�]4�"ߋS�	P� /3"�$���R58j
'�p"J��a�2�^^T��4�ǿY��%���W���u2��<�Dn��1KJO��/<8\pUPf��q���
��;ߺ�O��~v��(H��_�����,f�U��	�F_g��s��H�٤�����V��I7`h����z
��[��
>���1�iᮨ�`]�o]/�C�#&y���#�� ����������o˘y�dۏY��o"N���)~�����e��0q��Bs@�c�֏j��y��'J��Oa���zr��A��}����ϗ.ٌ���(��ո
7Lل��7� F��hZ�S��:`�Y#�J4{X.�Õ7L��9�*���\�eR}��X�.�RٞL�U��DZ7���jK.����%��?Q��α��E ��pP�4.t��i�L��WNs4� 17VYL��_z�x/����~����S5@����y��rũ������Ȼ.X�{d���``W:[�^��3��C�����>��3|��#��;�o0�*3a�-4��Z�@��RZ�:��Ϟ=PT�~��Kk�ڈ�Q�pm�(_�^X"э޾�[U!F�!�Q�c0z�޸�^�����Sg�@~�}��X�
��<y9�a� � �2�_�yx.���JH��u@����^���ЃQ��}��Z�O�n	FyJVa�	���Rdo����3���u؍-�͂(���HK������%g^s���nx{һy|��̕�2��S���(���Fr�%��ل�ڕ�N�+in3Lԯ�(���h�E��#�zT�?#�|��pf����B�*
��jVWH��;_�+T�,��]L�|/<B�oW0�LUz�V2<G�.)���s*�40_\i�f����b��8���M*�ٝ�������\g�Y �H�����������g |<|�z=]�s���ET�u���e�o�!\B�����"��C�q,��N����#�+�lD����+ Q����^^���͈Y���ӣ�X�����0V���O����С��p�dq��$аU�峃Gü{�j�b���ݾ��($6�VO�O&㻮Ně�0�t!�y�H��$�-1��El����E�;�@�R-}�DP	m�v�Yhft�q�^�n��P�����iغ
)5�Y�P��߯u?#�>�o����/M2W�Ƽȝ%֩s�A!��[�8/O��Ȱp�c�5
$�1S1�i�5�b��&֌���vk�:�JR��Y���{e�T]sI��е���2�Q�#��Q���Y�]m;�e*|8��9N�O!�u�L ��0~���F֘����wͱ��
��w~��/�M/�s4�\ɄFf���W(<W��-�GY��H��{4�0To ��MH�m*�M<��/�踳�	����/y_ ���l��������.�6���o�����ơ�f��$|7�����U`)�4�$���U���3;(��,��ӤbG�i�z�|��j�޽i;n|���Hk�,O:�� (��շ-9V�X��"���e��V�G���S2��f���.-����*,K��"B2��]�׎�JJ��Ѕ����.9�d��(����z��c���|�o�,��H�΢����6�r�A��������J��T~Q��-�����R�y��GX@Q�э���uX��-�2�	����p/�~�.\Z�ʳOw,�z�Q���!6��֮�m����|Cz�8J8�/��{NlJI��/u*�NШ��VZI����EXB5 ��`[�*��=h�5�����ժ��$� �n6k�iT�.u�;���S�g|���J��~�_�S���q��ݭp�B<PHwK���e��0��S �uS)��$:�&�,�J���I�:`�Kp����AA4i���$�U�?׸�����,�������G��[l��>���xU�����a�\c����v��%N�7���1�=��e۫"������Fh�!!��u3�p�BwXT��u�����l��+�_.�N�T-@|o������o<�H�@�b�-1l�@�ۘ�]�����4�Qp�p��Xr����v0��z�F�1S�C�WSh=|�XP��j�0��wJ!��x��>��3�����T:X ]ە��br
KT��J[̷܂�0�\Vm3�d���4�3�}w�@{�}�o�C1�:��*�P� �y��˛���~m݂���6l��#a�c�B�e}G�<{���k���3쏪m'�0�sA�������~��yG��6i�)�,��X"���k�^؏ȝͨ㢪�>��u�� O��j��5�B�DK��-�������RܦخƤ��3iv��i�."����V��qf� l����C��G���|����5�׵�Yn����kE��^� kuG[m�Nb��\۠��/c�����pRԥE�`�������n��,a�y���0���6���b��d�38��Yy]]��-,��/� ��EG���
����*��$g�k�9��-N|� rϔ5L3 �og.��W����yR]�r�����Ų��FlW��w�O��0�J�h���6y����pGQ�'>@��w�h"0m��6����±�P,K+��'ԛ%d�g[©��1[֎�?4��rf'�Yu]9%���L��O�52��E��4�zߖ>�&�dq&>D�,h�����H�s$��c�x��ZK�v���m�$�/���;��l}B���K/�ЬJ���uH����������&#-��@8<�H}x#+��U8�N��@!y{��c'LE�]�VS�����(^]�[���W�yI����9��o,4 S0��ln�ƅ|����P�bp����2��Z�ӏ��K�`ifW�Z���j�U����]sc}��1�-ϑ��$X�y����_�n���d�C�P��<E!�$�cS�V1�3�
�.U������_�*�x���Y2���JhY�����.w���2�"�iVQ�E���
�D��
���A�ˍt���r�C޹��j$4�|u�`x��8�s���)��^��{��ʛ=і�"����R��S���42�:1�( %�O��2����yŔ_P��,�Syu��U�lk�����ߘ.���6�C_���c�d�
��2���W{�F�H��X�\�����y�V�qH1Ϫح�._ �Cr�F��}���\�p|ȅ�ڎl!%��VZ;��n�g����:�¹�AO���$��:��)��ʫ�U-.es�m@iI��"C��@�+ �A������8���4RϧUߓ��S�6&�uw�&�$�
V!�=�����n|3���@d����o����Iw���f!��:���f8���ܗp�Ck����2���r�4S�{��_ݞ���C#YFE�����(ಁtڢ0m2�ݐ3D�Yo�FoE�VQ�^�8��l k��M��!����h�t��c��Mۗ���B*�2!�ú�9.mS
z@�w�L˵�3}�&ۋ<���h�^1t+���_0/>,z}�'[u+�8�cN+Nxٛ�e>�%�BF��H�[�?B������]m�9��u�w ����NN��M-�p�2��t�v���Չ�a��o"��!>zRB�oP�ةF|�����%i��`����E,���l�BRYj�9Xs\��A��8�}Z�J�:�j��p<�H�|��6�
_�@�?2�K&��<��8�Q4Q����8`~giv���N�:�	l��b��o��l�*��h��8��IՋ|�u�ʖ?�F�I��oz����W�7Q��}�w�I�}�9�?V�=�f^�TRH�Z�S��ږ+�$����*\e�H���3���_�s�
,����{�����8���js`��B}��O�,?��ϳ������\/����Z2����q4=��f��Hy�ү>B,���JW�Β[���8��ꖓ�R�Ƴ��7�w�#��L����Z"���@@���.W9��Z=�3Q;����}i"|f�]�j/��0�{$�dZi(�G��"�3�$�_Q"�}�u&����V��A�qV�WȠ�V�P��)ssK�A��O�x��C��|�M�t�(r�>�fA�K�d:�wRb��ع��,�t2�.+��)5��4�6k��� �g�觀Ro���gh���sz>�[�����ch4��&"��(t^�bCҼ��^,�R�L�~���e��������o�m[�-���_�zS&/E?�ʘ�z���צ��%9�����/kDEe"ܿ������k�B�f���2��אݦ+��A<[�����y��|e� ��z�g�?�e�f�z����l�E���;ś���Q�Lç����]���*��bEG�:�B�j-�!�E�j��(��X��ge�ʳ���-��Ij�-	L�&���f�?W>$F�AAt�d��t��4�P4Wtq�FjO=���]ʻ�G?F[�Gܒ���i=:�TW�?���u>���f؇�B��dF�\�h�I�aGnTT;�
�W_���s�)������G8�
ro�������H�� D���]�c�����#{;h\\�a��-����èO�S���J����{ Z � ���0"yu?��"��be��k�H#x���~)&s���={����ﳖ�N��h�Fj��x���"�/����,؟�{�3�s=�{��7�o@�6GA���ӝRqa�	q���%��ޜ�T�	��=">S�Z�g/[���ȤA ���x���}-�H,+�Yʘ�@���f����D�:�d<�*�
�B�<�ߴ�޾���[�c�L�(�fDM�l�����Xv�"���n��s`��Q<B7S�����\�>�D�yz�k�A�c�T �-l����g���� 8�~��!24E�e��s�v�m�$�MU�H;$�4��ɜ.��3�dۘQ&Ϯ����M�S�g�,��<^�-t��G���6��E�4b�}rx�PO���<_�#�qX�
4Z��PBȪ҉ 6����W�E�[�2S~��Ԧ�Ow�M�N�R#B[G��c��.�v�r���?�M͞f��N��3uwn�R%N! �*�~�
���͐�89�D�>��t�@�΄�r8�#	b?Q�q$���\�>k�tyԒ�p�nT�J�J5����`� 	��Ɖ�pʘt�O<!;rv�L8�����ĥ������)��N�?J�Pٱ)~4x�h�z�y:c?�������1��v1�i��,��p��P���cFN�ޙ�2Jq��㈕)�(��P7�����L
������8�Җ:�e�G��T �a���
�'�t>G����ȉ�֪Nf1{g�)��<1�]b!qRS�	�_�u���*�s�s�g��%<c��-���Uh��U���:��>��t��U93q���ЭyS+q��ʷ��XEL��9]�b*X�6|ވ�7��=�W�����0�㧼�Ԅ���#�.cINv@��v6��3��hn���q�J��U���:��;�k@qa��q�S���xyƔ�txF����g|��~1��gYr��T�ylw�9��E���#j7��O���j-]�N�`�W	Er]y$��������c�����+�#����@��t|=x�M��3���t�BPJ�M��v�*�- �h�!�2����� �� ��x��hzh�,8QIg�31wm,�O���6�v\)%��HﲓK��X�<4�5Z˳z?��-z;����fT�W"EEB�(GZ~��~�d�:O�5pȕ�6�0��w ��w7���!�<�tLVߤK��9�0,�eZ���,^У��$������|\�mK�S3<�v����O�q�4QQ	s��~.���,[�j�9�=��ܭ_-�d�Ԃl��x�6�<��kÂ����Ssw�v�!�pHw� ̯�hN�F��}s�wg/�/�C����4VR���A&'at��:�E�n1�,�jn�top3�ld�!i�vO��kN� !A<-m C�]�^*��y�	�8b/"�*�I�|C�DG�����^﹉�iuy�����E7x�x,�F�U�� r�W�+Z�E�x�!����Y58����?ҷm,�	Io=:5���5��Z�D[�Sc�:�Hy^0�+`W�s���`�e��E%0���f���-�g�Sﺧ�v����OE�u�����18�PԊ�Q��i��œ%IXe��~1�[Ԥ��-���Z�+;��M�4�Y��Z��oF<�(_���B�)	�D�'d�T�8����=7��`�ӓ�邜�}����Q��8�����rd�DLcxn�O�ș�w�q9�T�
�L�h����пW`mfi���#ԏU�X��m�7+g�J��)���1#2!P/ݥ��33�-�4�`�L���'1�]n]�Iѭ�b�9qo�c9���w�˭*ܪԹ��pJ't�_,`�(�l�\�J��͵PF�e��be�'xY�'i�AH��P����������e!Z��.D����i5��ɶ\3�ďd�^tm�O�����[�X����iV�/ʍ�6�~�>���c/Y����^S�y:�ՈŚ�ÿ�hd)P �w��/O�
��������Z�&���@�QY��f�B6;���AˎK{ݯu[?bm�g�)�=��#,Oi�>@����&+�`݄Q3Ü� ���$-�6<(2�[԰s&�jh�JŤ��'9�U��ʶ�����עW�f o
��_�|
�F�D�H�j�Sf�)l���&Av�+�w#�]>H�e��L���XZ�ѽ�</S^^��! 86���#7F���J��z�x̊/�����B���A^���Ac{��*r9&��*����}7�C��1���u�+\z�ޞE�ma���4��,�h2�JC�}�X��X��0�z�^���NNp�����^������u:��{Vvu���7�H�Ty�����l�e>�%��� ��p�Y�%�:z�1s�W�8�#m6z�/`�ް.}��w�:#��K8������Ĩ.Ǆ�#&�{�S�Y�=�xE���0��|d����r�\=�~��5�ԏX#��T�N�.��������s�#lq�Х��^��xE�w>3��&OԚ�B�/:I���2��d��u�]�	v� ϊcJ��H�2���1	$"�:A&'��d�����!#����x*�P�_d1�?k����di[b���U�|j����e�SK���p�Ygn�=߬{��C�M*]�&�'��	n /����L�
r�J}��tϟ9�=
s�a�4A ��0~?g�I'��7����i̡=q,�Md-��O@�R��K�F�£��9�
A�V=��ҡ�YK[�7OOvB'Q�9��s
�06�.�A���T=����n�M�Gx8r�	�X���-�=�xOV3��N��a���������<x+���O�G��8��ch͊�9ʬ�ؼ$�SܼW��v����s]ziy��`�9��+��l	@¡���/,����-�/l����m���
�Ncu��Ə�Nr�&����ZiP�zS�ߦ��Y�Y�!�G䟣��Z�K���$k#�mJ]�{f׿�g�{H��qӌ�<㇄��O���Vگ->7��4�qg=���!��8�b�Ab���|U��5��_��^Lf!25���s�d"���j���"������p���1�2��0+�Djy<�u�J�t�tˏ>ާ�����q��\
�tD$Kf��Xq���c9�"9%׋<&�܈�O%\9Q��i��Xj~���`1�"�S������H�!.�V:�W���`�/>��� �`�N�!@��U���ȼ|3����-�VpO�������p�`OXo���4!�)��glg.�F2و�􍘨���]Hɛ��ݔr�$�#��׭j4?�B�_OlJg����`cg��m���ә������[K2�́��D�k�t�nz����{���������t�13�rS�thr��s��!�Qϣ �]<�t7���+"Z�<���c�ŌVjၞ��9���#��"M���א��3��*�\�o�=d�a=�Z�u�P��!i�J������E@2O�{0�Ip>�� E��[;Rzx@
�dV,Uf���$�Ҟ�_���U6a��[lÂ:Hcq`,-7X�������Js�m8!S��T.�zE�%�s.{�!"@n��ԋ�0�+<
���]�"�ޢ���*LI�B7M�!ug׹��8��M��yWE�FL���������'&����&��6���l}�\��i�Ц�&tЌ�N��s�/�1m� �[7X�d�#ě� u�ۏdڅ;���v���k,R����g�BN.���+�ͱGv�G*�I���{�*I�͗�w���8Q�1]�֨�\2E��%Gr��+�$j>`{�>�в��-��ֻJ<��a�V�-,d�S420YS����!s[z�y�+"�˵۔� ���e!�ң-W>"M΄$��a.w)���$�ms%T���F����;�+|4f����!�jaE�f	йF<��ko+NRn��#�t�(H]�:���s�6zD�ZB��!��}o��))��m&[l��B�DC��C�A�u���Z�ct�M]V_ӡ���\�t�k�\��ȿb�|'F.ڴ���|0�6�mXNr;�A2����3. 1gGvS�WDS�۴R [��^���4d�:����	�L��$h��;hB+5�	E�~mn��z>�t�n'������`�K�.�qvYՋo���$��*�40=����h#=�	�eծ&6_%���N
F�u����`��BmC/�k�7����8P��.�u�
�꿶��/��dY(�q�뭄�X��z�X}�ƕ������[����zK��ۍ�	�{ޮ���6Ԯf ����Zi� �eI��sx���i�h����f�;�~9�l�0�˱(F0/׼n'�����h�UO%��;؟75���>�m���u��<�^c����Ka�w�|���^��w(k9�PYWW	KA��6�߿��P��0QH5Vb�@�f�kf�պN|�=G�=���f�i'�x�+�x�	��?ۊ��Q��E*9[�v8|���o��� �?C<�L�E���XV�ĺ�]��P�V�
�]��TG�����4�W Q��G�2]k1��K��c^��~��De���!�h~Oq�\ʿ�c��q��)se'@8����%el���6)a/f�s�ݷ����B�#���s�]���f� s�/�"g�id�����^�>����Ҵ����sBQ�k�. ���:bzH��Ğ}�Ww�v�=��x�MM��p�"t]����)�yS�-F����w��ƣ��p�j#��{�aن��v{�D��T+~��H����O��ay>�5խਐ�ع-��+`�͂z>�N���_����`i8\~�GJ����(��Y�$���"}������N�B|�]v�\*ã�*�fKz:�䪻����Qt�q������ؔ�(̜��3�!fE���X���8ώ�]7A�X��/ק5�4����L9�é�¢�c$��C��{[�3VY�����8���ޗ��3�b�մ^T|i�nF�����y�O���">a��X��B�k���i��<�q\�J2�S��U�dPfu���i%ؠ�񟳅��r���,�lZ�r`���s�p�x:�I\ɿ��W��-Q�S���n�'B6�K9>��|��s*��ܡ�`,4��(�R��SC�@t��k&��/����ZHx�aW� ��69�a�n���+��A򚚲e��-K�W\A��5iه=��e)��\��k�1����P\��%�ic�'��1��c{�9M���tJ��Z�8S��m;�#�j�z5���~��;(�/���lP�l�6({��g�$����\�yu�(`;�u��,Tl~>d�	���ԣk�Q�q��6�R��
(e��]g�J�7�P�R�@���0����w+�e�����)I�\+6�>٬�룲FM�0��m�=+}���r��&��C�����n9�~��d�4�UW�d)�I/�����H=h�}�����
3�y�]#�6�w���(z�sF���-K�сԫ��l�sߺt�kR�필B��M��V��p/GN9e�@L�o�Wx>�U��k�c���-J���,����j�`R�ճSc	��	�:��F��Q.����yv�K_�Q���^h��7nx��o&O���e�Rj���6R����>T��1-���]l�lzR��Q���Z�S+������~��q�"(�q�7��d�o�of��@�v���U�Y|J��7�6�D2��C��Z�\l�ՓlI"��+�h��Ҋm�V�eY��&���)�O��1�L��F\�3�s7C��. �p	*����HMߚ�.�$�~0����ξ5sJ��*_�]��b�\*h��$f��D�l�s1�u6��"�C�Y���E�9�ަ1���'ØZ`[�}�o�z�
#�k�zu�U�Uo������BrB��[���J�_���X�.�����#�+�4җ����v��b :���۫u$ݯC�
鱰Ә%�0!PV�u�,�|����7}�tw�'���6�"�{�B�E�RF��Y&���>}Ǯ�������G�T���+��T�~u��BN���1p=(<��B�����[TS�^�u^e�E�C���� �q	���^:�5�������"�7G$Ye��R��"���=�|pE\��{��!u��{�/�JZ���� �H�h��}m�w1/�{�0?l��~E�Ms�dr�*1Hp�sgӊs1�y��C7;��Â� ���,Y?�Tg�B���ߒV�D�ԭhw�2Y`�d���Z=���3�1NpkӴu���$����i����+���~�d�R]��t�̈́��M�R�5i\�l-�T3;sX�E����%o$�9���S�ja�:8�@�Hy�$i�i�!��.J2�N��f��2t_K pd��lْ�F��@b#�r���[�I�t���� �ۿ.6����jE.d笓�)ؤt��|��=�>��S�g�2��^�R�����4Z��*]�����#��qD�w-�c�3�{�-)�?�#��p�:D5^�������w�NJ��|1@��TV6d�Gw���MT��ݑ���lۦ���Bxީz�˦���C��)0[n�N�#����Fɥ\�$Ϙg�Hb��M���'A�5��][Hv���jJ���H��nbt�L ������E����Ә֑��=��ͯ�|qW|:ևC^��Hw����m�P��y�k�&��-R�-\�K�i�ȵ�pF�u��/��wP�D���L���2������I� ���
K�T\%��j*�H2|�=���hL��QY*:��IM�o3r�U��,�u�Z3��`����=�(a!!}�1��gr"�B��h	W&Y�oT1�O�lu0��0����m��$*�X��a{�)�2�Ӟ0*\я�c�w� Ͳ����ӧ[̮-�3�5�2�Y7X�񬴯��8���W��}��ǳ�P؄P�6N�~4�.^��	�l(���՛��K��@'����tD���{��^:��3�0��KP��G<3�8JoS�(ڛ7�5�r�� (fb�,�lb�9�����C<!˘0��]P%�QA":��\��C���|�y#��:9~�i�[�#����u(�p�1����2]_�R�" ��#��V˟�����((OW�C]��DH�A2����/Y};�6���B-����A�X9e�9�>DU	�N;t�/�U��4��5�2h{���lt:i�s#m�F�-Y��LnY
�b�-�Oc+�����z�}?�k;%�ޙͧsj�����}Q��I2�U���ixH�|/h��s]�q�H�-���I%a�.�'�x�w�>�D��/�qMN��H�%���h��Zwrq�Zq���5�BBq���T�S�=n�ui Ȳ���A�8xy"&��������:��M>�~�����Q7�L��妻�_�}Y��cLJ�q�l�HN�xS��@��r��ٕ>��O�L�Q���v�`ZƩ��{Nl����X�~Dr��p�}s��b7=u5	�p:�f����d����bYq>���K嗮]CЀ���s.K����a����#z�[c\ÿFS� �jd|m�_�G�u ��Y=��^?�LF'5��T��K�4aDpG�ǋ�m�-ӛLZ���{m\� ��q-S��_/�P���шL�Md��!��(��5o�k7NȾ���KB\N�r�X���t8�H��IR`@t��C��'�=��h�qg�L���CnJ�/��`zp�����Bv�cB�PFM�'�^�Ͱ����)Y]-'4��K�iZ��k���D���
��O.Kp��0�;ߏ�B�<3�3��*�''F6��>��Is_Y[/�o���H�V�	C���j�L Ďѻ�ݯM{"ٿ&h|���`
^-��y;�CB�����NzA�ٯy�W���6���c*r�ӧW�r)�� �Wy�o��^�$t���v[؂�#k��?����j ����*���硍���|�P�j�]�d}$]5�\V��0DO��9�m�qG���;Mc-�)J+AA��8���C
����8��X�.B����A�K��:��a[�H�o���������x��C�rT�<iB��i��.'մ=�1O.�wF����G9��l(u���x;ң�vs�Z1��}�����* �����������:=���b9Y
x�wO�����^�d(S$�� wN(�<t��wVB�e�X��xx�c��-�i������Ճ���;~�����Fʼ�!\Z?��'Ũ̌-d�/�� �m��@B��U��U�2Q��
QT���J���6N'�}�O�o�"��e��qh�i%hh���ɦ|!��{��)&�;y'�_(b�ţZ+�h��u�q\�������1a:!z�J�C�K	��D[�0  } Ҟh���$2�c6z��>OK�"��|�lk��Ʉ�F���JS�z���=���U�������C��E#Μ}��wwK.j`o>���+2��MT�S*�SV���H?S��Ca�:��2���:[i,sQ�����@��"�j������Ȋ���v��2)apo0���^`����{�|�=,S��/�3~�N�B�%U��Ʌnl�N$~^��Pnh�B�fk+��A/�,A��@Bka�uH��!�4�h̄:���[��E��򻸣��&�N�!�}z11j
d�P�۬��X��^B��<�v���-a��1 /����u�J��jQ���L�+�U Q�o����L!�8>��[Z�l��C�*
ڄ��/	C%�I*zU�� �����(g~��>�N�,�W\��m��U45{���� �T5��1nΫ�a����$"��A�93��\��(G*� �\A���GK���H9k�[F%�c�yV�	�d��d7O�#b�ǪU�� L%g���	���;q�s)�+$�L',��]�C�b�a��|�����|���ؘK���b��{XIa�ܹ�<�Vh����y���@(%9U�����Mi���n�+D*H0ll�@� q;2�}2.A�"�x���Wԏ�+��"9��m�lg_jr�<5�;.B�3��z�u^c!%󰒕��73)������@aY�#nH(ۗ�>p>c~�g��p5v��C��[�LTއR��D��'_ٿKB���}�%0�g��nP���X}��\,T��ɘ��`��+,,+(�W�b�ngwV�OC�v�0ԓ�}���Ņ\;�E&������p�fm��q��n��)@�n|9������S�F5�F���Ok��ص=�n'=�0i�r�Tk����Oa��������Tk�bC�] w?%C3`L�L��v������J�i]����bx�,��u>���=�H�"3�ӑѤ�o0�¶&��X�/�!�_�ɞ����o�������y_�q�2{�0o��^��md3�koP#^	��X��FAǧ�[�~^$9J������S�ϫԅ��U�w@��V�0��%"<
� ȅ�O�_����LD z��̕�d�H���9;�	��m�2Ѽqǩ�-D�'���bt
���W^��P����w��ק��1L�yZ/&�9'	=�S<�D�F*��Wj�]0��.d`$#nP򏛻oR�����4��+�6�8��v�C|�������$�5�:x�!7��~wgC%��������QR����w���CX��z|q8�u�(���"ݽ#bP����gF���!g�=�̼D�!���%fV?0��?Q��@�g5h�٨�ӪV�`�������0�U-�Nω��;�K<�<h�����e��-�O{=�~!�ؿD�Y��:��4�KA E�*:�_}�;��%dw��.)4ȨA��)�n>H"(����723.	�j�ғ�^���}�UTM��-Պ=ѝ�l:�z4�i������؁:M��-[;�L�+ڹ-X����aE&&<�z���t�Vˋ��-UY)���Y��E'�~B�ax��`��_>�ͣ��'�<�{��x|��chhIY6�����k:��-��aB+�XAٰ�'WY$;;y��`���D�i��(ȋ߂Pm�y�˭�4#3i�
pu݂�������Z�(Wu�,����"��򐑉��σ�R�<L�
��g�؎��~�q��/���z*�>�a*����������B�68��ſX�s�v�T�ğ���/��xeSF�ה�=n�Ԇ��T߲��{�fs�Im%� ��	~�ں�Bi<�k� U
S��Y��|u):=z!���WC]<GK�>ܘoz��4�A�i�I��
\�-m3���q�p��{��z��}]u�vK?��P��TS��x�$��E��b�(�9����|"�Z�J�}����hV���s���RV��*c�/�>�xQ����)�W��]�r�]��C<�Aő!�ZVRG����51i�Á���O/��;@GQ�8M6^�>��:ܢy��2r�Q19�&~Q$4�gՂ��P��
FZ6���Ɇ��/\��&�m�c��&]�����p���Ϧ�=$��Kʔ#�����C�>+[~���	�K�J�e���Bv�~4��Wc� ]���k+�'�1>�s��٨sKu�n1q�7���Nof��z`=�[K$�.&�D#?��;G�:�aF������6�92���Ia��K���X;���4���̋q�Et�C2�b�VS_C)mQ���]�	�($��Z��Y.7�R]E"��Lk�z}����*�����y"� }}%���|�+��C�ʹ[����h��5RC�i�����&��c�H��y�w#e��'�}z(�Ò�:S�"ЙBy'/��(̀.]uG���c�Ck�5�YG��ΐ���B�yg%� (��;PX� :O���k�t�t.�d��ْº|-���E�k�X����$l�d�� ��M;�
�p���Մ:=�gt��{o|îe�^�L�+��N,�Ǩ���.��r��]Fϲ2����@*�9��WH��	���'/ �V��EU����Bi�%�ѕ�oO� ��$�EO�Â-ֽ�L;�J$Q�$������Ȱ�x
�=4[� h �y9�M�.Zj5�I1��ɍ��m��?��p�V����ж��n�����G:��u��:��+5ٵ�tvW��X�S'����t6�ZI*��hȁ�i?�Z&�u�4��0�%ӱ�Y�~`0�77�'�	���^i ��'|�9L]��i�4���l��6�Oot�������e��4�x�tj�~�aep�Ĳ��M�+2B��Ú݁V����*��gܽ�U"�%݉��ц)b}�3
����Fc��cL(�����W�~�o ���wg�`
X���1��37��͛r�{_��+K�ʐ���CD�ڂZ���<���EZ�S��`nm��J��>h(���*M��8zy�2�Ȩ������l����;��y�b:J
�+\�||v%TQ���A4~��}�	��P(��J��� u��T�}��@.���œ��e� km�tr:�@w���@�R�+�G�d�S@N���)�P�.�n�U���L����%�E8Ӯ5��H����?.t>k\��풁��X1��$/M�x����Ut)4�g�_�N���sj�1�'301Q�ء'����8$��Ig$����>|�.�1K	?|�1v4�q�s���L|ӦBY��1w-��Д5�1�&��C����	��H�+"�(�bG�-ne�\,ĕ� �,����7},�s����CBxd���]�����oQ.~�`歹+!;�JgK���s+Ut7xθ^R�w7�&3���%/���o�Isү5��˷X#f��=R��ð@�@�y��VO��L��W/bޞ*�a��;��{��z#TĮP݉��xLE�k�A�΋g,2BQr���]B�Ϯk��XO��S�5`ܶ�Z����|���*�&��TY�.��~\�'���=VoBjM�(�k�]_���-���d�d�W����L��[;LןHOd/�;r!��WC���7J�Xt�|@�$� �tq�У�:��͹ ���%ϕ�%8t3��l�.��๚���^[9Aһ�I���6��,/f�3�2�������0-�3���k�9&y�d���B�� �@(��\�"f�yE�.Ye�c��׵��`�L/����>H�[���6*^��
B��M�eA�3,Ĝچ},t@���c���� �����ns,�hl.U�ڼ�]������~xەzؖЏY(Ag6A�Tr�hD��y���bk�B��=LJ� x�YasKуj���p`����+���|)UԦ�m�ͳ9�!`U7��g���ҿ�Q\]���F�߷n��ï�`WU����Ī�2xJތ,#�o����*J��!��W������$��
�9(A�*����AȎ<���̄��`���<4~�vL���:7͜�>$(�U���-ŇZ�:��o��c2b��=[�����xJ��o���3�tN<�s��(瞈��[�Jq�����<�G(���5�n���п���B$;��������Mi�tM�z�}&��8>�S���a����?�6�X�VyW�Q����f�Gaek+�$%t���s���]��E!3M�Œ�@Q��>������
�'����䶣�����U5'!�YP2>���0ΏC ��<�I��7y��bn5W��WG���@�$q��z�&�(YfY��S!���V�P�J4F1Ɂ�Ŋڮ��f��a=�"�I���m_K���F �43������{�~C��B��k[z��}��^��s	�]�3~Ǆ\1�����MσP��Q�θ�Z]�wa�؈%q�R 18��)�^��&������+���g��	d��b���.���f���͹�3�Mk0Xw3a�n�"�-z�g��r��}��ى	�r���]����J`�*�+�����Ó�K�tl^X���ՀE������j�63�|�q��i��7�iysH�l2(��N<�Ѫ /q��p�b�q���d��2��^M�L �i�]'��-D�洛g/�%���+!Dݢ4����w1������^��u�=d>#B�0��k�k��^gn�$�>�QV��(�a�Nb�\lG�e�z��qSs���7k��%�N�%f����/d���1��*�� �ؘ������t��h�S1��^�\7�|C  �EZ�px�m:�Mn��A�#�P@��4��̗oFu*�D(�ˈ�w���|gV�o�z]A=��ũ�ڍǱ���PXł���%Т�J_��"^���	���߱(=��j���`Cifw7Yf�<~�N��B��KO猯�+��j��RO��X��a��(��?�s&�ϜG������X�*0���oP�����{�H*����XN����Z�*���U��pt���^��dH�t��7͍��#��Z�It�C�����HN���<a����I�0n�V�t���ز5�y_����Q
�<�<��N��v@�ފ�xT�%1�s�곒��LW'�ÃbT5��0��-�S���.T�Ip�90�niQ���1.��׀uOu3F�������VZϳ���Ȱ��(V\����5�I��:)㗆	c�]3�C�����෭��<��QLϚ���_�5�
�M�����1�h݊��;��Vf��D'��-J7�\��H��Ȯ��$���X	d��s6��8 boŭ���E2%2!T%�)���*��p�-��Ŧ�`��jd�T��cHܮ����a�𓁓@G��H������)�/橻�u=��}��7��$撮\sޟ�Ӟ�3�� ���6��ӎw}�����2�ֶ;�x��������3���=	0?"��fm�f�_����{��탂roka��u\�$��Ig��@棏�^t�(�B&a�h'F�=7u�����?"�:�Uu��ɞ�9V�`���Y�E~�n[�IN.�@�<�WIG�Kg��e��_q�g���W���tykқ��\�f�������!+&/�ؐد��r�{��A�G,f�P���g�pQ���C{H��I|+�_7��KK�M#b.���g�A�dˉ]�i�!Bn�~��[�K�V��������	��`Y��<ʱ����&x0��mV���K����Ih'��]�=�Vϔ}Q�J�M(Z�^�U���ek}���(\�!?R�#=}S>��(6�b�����R�_>��N�N���
�Ku�k7%�e��j<�P��g��_(�+G�E5�P�6q�_Z��ܸ�_9�27�V��q���	O���uF?W�H8-̄l��ɗk3%D��6N޿�?���3/���J�7�q�hC������E;��8�J�1@2�����r]�uO����r��0J$g�P��i�d��z�CJ�d7Bk;m�v���~����G��i���(����L���3>Q����y`Ud?���T�����Ĕ���^_5�r:�1�N���M��1m�Z_��/�(|�r�������Z�b}TR���i)P�h����i��N���DY�V��`^�}�f�f�}�e_-����N���e	=>R��h�d
.ы,�ϒ/�}�0s��5���&�ܐ;Dit)���w ���q�1�)5k�	��ķ�F�;�0r�~�W{��rM�<^~������Χ�k�#���ۭ���;*��.�w�p�q��A^|��O�*��� -��6(s���'�2k^̙,�jY��t��j�8��R�2�\����9����Y� `�����C�un�9fN�0ĵ�ao�Ek�9�ȗ��S7�E$���x�ۉ�Q�r�h��Ŀ���>�s;�`Y+7���H �N�t�=� Ś��=s�b%��sFaV�\Q���\����Ub��\�U��(R�A�P="�X �����T�z�5a��%�?����\�P����Ӗ�`�/֍���,M�ζ̮L���b�(��O�u͞�k�8K�r����z~g��x�=�ﰓ�H-�x���U�Xs�?O��W����?Os�!@��>gNk��D��S�TuI����#���WݛV\�M\�(�lS٫7"ʧ�����v�V�� ��6��u����4�� /t�_/Iz0���x�w.�v!�nN����9$��s�2�LC5nc�P���򪠋i��2�Є[n������#�t��Q� !�Onuj�^�0���B��X$�$�%��Qe��P�Fu��?��ژ�R��f�a��c!I�n�l������w��O��V�?8�N���I��tsҐ����*��b�)IC�1:ex��Q��[���'g����J�qA��ݭ� ��-)�)�M�j��b���(�}�۵��u��D#��Bc�BW�((��I淚�wz��1�ݡC(!(�O$�T��|/�f}A��w@S�`ŷ���tͭ䇲�3��PLLH�<�U]V�Xi�rT��
?�\�f�;k�
�(��B"O�@l�#����KF�Hq)孄%g��|�aBO���Ӣ�.��?��BΊ�K�c^�Lu<�O��:;ixĪ؉O�;zh!1N?�'��Dh�����Gإ�UǰYѤ#���Np�])2P��'9�
/"�Y�L�z��*�p0y�G3����f��(Z����ð)|��[%R�ʃ3�N}��~*5���ت߂Ȁ�O8�W� ����u"ځ�A�לN�T�,:�\e��Xe�9�Z�G�'�[�fV���}j�#f������YJ�����X���$�q{7�z8M� ����ؤ(y�<��ΆR%��d��`��d#>ʹ�&9=w&_v�gЏ�b�`��c�1_�&�~|�B����W�Y��%�a�\~�3��BL�y�Bb;3ݛ�;%��9{�ߞ�Z�{��P��^L������z�/�5�;ۓ����ʀ�M�v���L,V?�E�;�d��w4�IR��;��Ki��+�I���K����T��s�3�a�L;�����HH�(F	������̷������2D�CV]��%�;��n�N5��G��YL�7o�)|�!���*�K�����hre@���]ν|H��We_a754�Q���A������˽�G&{r�M��oO�H�4��I���M�VCA����Ɩ~TVD�sB��d��17�ː�3rۏǯǇ#,������8k��(��YYw������u�X�� ��Y��V[2m��w���w��X�`���"d�Вءc"��5�8�B���>%',��n�-�����q�Def�H�`ڡB+����g������_z�ڤ
%�y���R����_B��k�ۗ#,��D���
��=�ʌ�U1#$��.��C(ɪ|o���;v�	\�>�����3k5�;Fz,�����ѝ��?\���J9��n9s�k�������<�3~mIمl�Z����4�鳅3��Eh"�����U���t��G�  ��m���!�n/��-��;��m�~wm겷+���A#�����."�>5�,,�}�����$f�7ON<AKU���v���Οh!a�V�!}~0����~j�����#�8k����錳�F�,%�t��ࣸ���<�nJ�g�N쓅`���]�=�v�WWE~� ��L���("pP��g=�"��eQkN��S 3Бm����!`�������j�`�āZ~>���p��4M�Xջ����o�YD���V.�z��^��������O�����,D,Ǵ�<�#}s��u���
�[=&ߎ�8,�&0�x�����]��g�&y��M�B� +�A�eP5�Ǩ͏P9���[��P���(u'�Uش��p�`D���Q��ȼd|
P&gG�&��M�`B]�b	J�u��n��p�<ܔ/��{ɗ�ǱK��j�x�:#&ېq�`�q8���.���O5��U'rZg�_i�4�Ã���C���/I�z�.�
�R���33Z�M���n]'�.T����v�e�{��^��
YLW�w�B;eN�w�S��ρu+)i?b�YRIH	��,dB���É�Dj�|ީ|����D���À"X��ߞ���|0���V��o�^q��j�"��ԉ����q�6Π���\�����9Rx�1=�����9ږ�7�]sٶ��n!�]�Ϩ��q�3�{nάK{i�,^Rf���& ����ߍ`�J�z���p�8O�LE�$L; L �CD��n�P��4�g�|H�(�Me�J�Db�ʘ5<�$��~���Y�[=VՀ �!���_ףF5lm�;xr ;w�,�=ݨ��L9�M^p~h�Hȱ�¶��$���2�H�}j�a�ԭ�"%�q�9�vG��� ��[�,�����i�������ĥS	��0�J�G'�\#>=e�����^N�ڭA��Ț� ��t4�V)i��G0�
�j	aJ�>�#NJ�q�]�u?kZ�9�K�����KS`H"�R��+}�J�^B����OEv�W=����a�㶺��s������P�ֲ���kH�Y-��m퐉�2��S P*��#*�������\2�<=�I/D	^b�S����BP��՞��\D0d���U�D���y���$�� kM��p��?����{�-Zd��$]7U�G�&`��/h��Ln��s�k�*�s��mt����Ӏ(7 ���i Zl�+{�ή���SoM��?�!G'��djI�F��p������.|$��D��2� �],�!;:s�Mr���=1P�O�L2U��!(�Vx,$,�E�P�ZmY�ˌ%^�׷�uQ���;:#nY���v�`��j�����T0�촔�~�xJ���&��N (R�RB�*�s�3�o8z�2]@��E�A4DE���cE��'���S�_5`L���'��1��mY~��6�������	Ln���א; �S�)� K�S�b��v�y�c�g����q��< $�Ȱ�6��=N�������1r,k<D��/,��ԇ�E����x��r���m�����vk��E�G��?���+�T�ej�~�H�?�U��O����`X��.w�E�\d)vg��2�0`���ςKt &�thnf:�ß��� ��[��f�N��T#������9rJѹ����R�<���G/��k�7�@�'�m���IK_~W��$������ ���{��D�8��x]��txn��6���˹2�^���ۖ�c�X�����>��h��:�>V^�����Kd V���F�+TZ�Wt��UR�A���s�6�WU~h{�R������e-]c2�^����f����I���h��ݓÆ���i� (R�ٌr/�㓵Qc���$!sF��'$G�b�ptΠ�E�yޓ��d�p�y�7�"����b�n�s(��E{R/D�~�ߥ^*�pK5���2��y�KR!	�[椢��,7�3)��r
�V���e~�o!���~��.-�즨��I<�fk�s���,����ƅ�쉭ņ���.���b�VS��7K%���o�u����6h�D����nRd�<�'Ƥ�g	Hq$��Κ�0�-Q1LW�7_�O�nm�����;�8v�-v�.�����9Y����}���l�g9�&�=yw��@�Ͻ^�g�G�;,e��'u�	�vc�<�Qx�K�����ӈ���a!�ny�/�pn��+��+��G��Y���^���A�gn�I�e���w�1�4��P��c�t���G!�c&.s�cbIYz�-��N���MAr41��gL�"�gI�*�WPBT��b{Qڳw���F�R>mjB�`��N