��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI���!qp�6ht����B;dv
�[�܈
�/���t�!HO;���;��.$?�'�-#ܨ��q�X `*Ƈ'�e,��Sg�Bno~����1���V�0HA�=/�c�����)7!/2�����&��������N��Қ	Z�G�i؈�7ХP��^��S�T���4a��I����Zp^�B���,��1�W�؂���K�U��=k{�LcF���)��Idᦿ�_�Jy�����d��iN"����#�,^F"��.P�P�����9���})��ւ}�?�T��;_O�@0�|&���7cgKD��PD��댜2�.��%`:N���n�@�8�ݘ55{�K�l��߆,��`QJ���ɘV��kF�B��+]�4E�`�8�`�-��a$�$$�.~T������n`-*k���_�il�
�J��j�E�@���tΰ�k�V9�ň���Ԙ=�H�ZE��x��>d�2:��@��|a:�쎠e��������`�AF ����Fg��#�t5̠��|�ȯ�;�K 6�����xbj��t��[�%���;�<h
"nY$�S-��P	P��V��VR�U�C[�2J������1_d$2K��6h��)!F�Z]�
R�Ԁ�a�A�f���#��cv�-K�ͬL#�� I���&�.+�䔨�m�eBt���0�L=YH�&��� ^�1>���	@M�~���3��ŜX��l�7��A��p؝���
 �Y��wRd�W%>w�c|��f@�d��қk�ӮlI�үC�s]�\���êf�	�f.(����1s��w�B����Xѓ�F�ޙת��p�jk̄����_?�(\2K��@����/6���#���X��AW��pbO���/C-k��S(�7����>8O%�ե��5�����agT\�j��^��Sb�j�wCm e�l��<� U��|��Y�1��_j&D̺v�4�� ��E}�5%4�~�B`����~���B��o*P��glɦ8�|ny�'6o���2e��B!̇��`��y	Ѷ��΂Y�tB<+�藃d�O�Pl�؉j����<W����ia�ZM�?��S������T��@a$�2X�5(�����H��9�I;�-�R�ǣI�ۧ죴�5,GΆ/�Wf�vK
k?�KG��sz��2JK7���>h1~�y�*:����|Y�E�>0wȺA���~�՘+uꆚwF��oo�#�^E�39D���â�E#편��-��*�G�*���^op%�A/��f ��Ց�S��t�+��,?�Rm�{ �"��
k}��[ �����;ʴ��&��RO���i�0�.�e�*<�Y�<�W�<�|2���_6˩-@��apM�Gm\�F�u�����4��Ȼ�@C��!E���M^2��.HV����e��U�Α��Y42JY�����[P6���F$��i1�_����h���ѹ��\�1�4���K�V5!��?���f1#�~���=��hR�!�ܷp�ѩ��	�3�������U �֓�+eNl�%g8N[�Aʨ���u�e����O�T�T̗wfk	��ǨN���A(������52!ť�JuB�þ{6P(Ȍ!*l�sh�f
m]�q7}튣e�jՏ����vPѸ���q��3�,\�"U�$6i��_�](kь�#�願��G�р@���O�br��?���eʮi�Ffa�`
Ԁ�\�Y�����
���$��0Z�|K�hR��iήkJ�֯'��!Y�=�(!���gMR�Nő[+k�I�����q��C���� �F6��_���ܶ���}F_.Zb�"�:<��k��ʡ���H��_�)I�t�{����t���q�ԛsF5�k�!W�C���m|۸��R�:�:�sS����Ϟ�
���M;�6����Yʳo�v1Jc���Ǖ�?�<��OvKNyr�i#�����ne�jY)m�O..��&�I�u0�Izuzҫ9%���
Q���P<��U
���qy9K�3&��:!'ߘ�%
G�S� k0�d'�\�W�,�B�.1�9W@LZ��>��J�L���*�-.�Q
�6�B����-fVi�J�!mq_[�N�0�Lh�Pe��7R�?�p��}��yab���@$�a#��V�H��,�������������k(������Q�d���S�[Z�Ur��٢�k�|�]�����H���Bh�� ��a��p�)j)ȿ��zB�Nj�q�v��t�ܛI/���x\�8��w�5._�3�1�]������@~�p�q���Tc�{
:��R���2t̰�	锾͕�9fڃ�����=�u)L
V
`+��T�V��A�p�g@f�����hrS&F*�C����X� �Z��Y�zn���Juz9����C���t5H�r7��4~�Yi����02Pe����\�B۲�{;���L��S(oi��|�r��