��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z�O����_�F��<�DBz�2g�Q�����%�Foͫ�����n	�C1j�y�̩�YJ� �R�恣�Q��'kj��.m�� Շ��n^�1����a$<KԺ}wEI +�&*�����j[�� 'E������Tz-�<LԮRz1���
r�s���F�V1��[/#�;� �p�����^;�3��F�I�1!��L�E�=�K	/��6����c�_��sBE�m����.�+ϑ����yQ�LS�°xZH�z0�*'Iօ1q�Sِ� j?yھa��d8b���ϒ՜�+��1=�r�?ۏ	 ��~Dp���Cb��X⥫+�eh���!��9�oH��?�-�J�)���x&ȽP���DWڥ�{����L�S�L.���Z�8���x��e�i����$;�� �Lp�\s����7�,�#���O�*�U��£(�qj�������Ah���C&��1��ƗfMHT�v����N��=$�~ك=�]�r[���m	y1�2���b]��8]4���Ѭ���.M 0�ce��`W�#վ��k�ZQDl�V�Ad����ܮ�������)2_�u�Ě]��ך��%Ր��������%���G�nO>���(I������?(Ҩ��|�Z��oT�7�4l�O��Y*����6ċ�>w���i�����b���E�2\m]a�%� ��-N����ڽ�N�6w-��`	��\u&�yE%0���5ڇ���0�,1��e6|lrA�p��J;DcRvp��B��i���Y��L�ʩ8	�jw�~)DM�=��9qp~�a�WA	���=�ׇ!�Ϻ.���F�Q��/|��XK@��u
c�>�?�p��!�:��5�*H��!�Ŀ�e��,y~,ca ���6��*Fbgm%�Q6sϽ_�������ɪ����I� L�G�/��ؔẌ́�J{3�Q��BX���jB��N1R�����X|�A��O�	�Z��F��ͭo�ɪ��S9{ �au�K�.<d\�;O��Ay�P�kxg�*�lҍ,��cQ��m�2�C�k���M-��<Gt�<�ׄs/�u�2�����lAS�9j	���@(\$�fݪQ�H��i���fM��w��GZn�`�f#mGv[�5yE�QD�2�;�^^]k�;�J) ��������5���T?r(�A7Ӱ)����i�Q�k�v)y��L�����߭�9�
�����Ne��p,�[�Fvr���Ņ�h'�Y������p��w� �4�Y9��ˁ�ɱF�������>��E\��g���h�Q3�Q����>�FRˈcE7�į�/)�"W}�����/ү7Ɨ���w�tbV�-\˩*y��Բ�.R��(��\8�ᗝ6QRL�.�y��Ֆ��5��.栟�\�:���1���}���,�)���|��N�F0HX���r&��/$o�/OG"�Ro!P]����J�%[�������Hq�|�2 8\L��6�����-�7�*X��ҧ���bj�=��mw�G�Ü8J�jͼ�$ Xb85Xu�f��S/wj>OA�("Hy�3���&�r��R@����%k��eQb4ܬ��\p{�-��g���j5^�As��S[
�X����}���c�_f�d���q{��H���
2G���E��5�Ѕ�;Mт��H�����*i^d��J'����PT��X$��B�Hn�b)� ��$BC�=�n8g�4��y5Z����L�I'�M�T�:�7�ֿ)K;�20��1��)~�	�,�sQP����zP�=��Qg����)`��4���2,	ź�|�)FW�C��Ɩ�4Q��ئ��w��23�Qb
Fگ9xm��Ehd���G�Վp��Ԗ&;j��M+�u{ R�X^/��ǒ�ݕ���Ȇ��@U�D+`�D�ܗSƔJg����IE���7�KI��Y)b�A2M ����H;ĉ�j��N�(��t�H��C�5$_�9"5�_j���#�LNr�v>}�ۨuh6|��?���`*5S!�H�l�1�ƛE��:�ۨ�Ð� �tr�<�z��E��w��%�Q���x��Nً]5�:�&b)��c/n^˱�y�9����g�.�y���fb�;I�Lj�b��k�(�W�j�O2n��F�k:��o|>��oˌ�a�~=[�2¦0<	�@���Yr���{L^<.�G��Q=S�(n��ܘ�^��ۧڳ��DT����6Sx�<�����<e���!�{<H=����c�1���'yuY�dW!޿>jk��Ta��(9y���<��3S�q�`��.�]���X}���zN|�>�
��YGꥧ�Vf�:�8�p�v�ޫ54T$�����a9�ǒ{S*�wY~2�?{����m�@v�UQ腿5y|S���j����֛���%�ga/WgTiH����}@��װw6H,�vM5\�M�4�6��*�ETb�u{Rѻ)N��?s�l�?�u�]���c["憨 �0{����g�Q��.E��rv�U��`4�� z�Gr[�B��ں�g�(ɿz���p���(k�n��&�Й�=-~�d�2�W��v��W���m�����5,��j����S�|w9�Z�������
D�v�|f��BWz����ҭ.،��b_[Jd�½�Vmd����y+�ļ��ޱ+��/p�Z��s��ޟVzF�l���X�b�/B�f�V�*ؠn���6ڭ��+�(��v�}�c�����v�T�W9ϰ��-�PT�(����/X߉�T6E�=T,�xH欩x�Vd��tZ��5������Ow�E�H���ɨ��[I�R�o�@�e�nR���Jh���xW�_��f����T�?"90�B<g�}U݃b�a�Qr��l���h�)=H�/>c9��ګ��yЯUk�g!���	��]?+����ߖ��&`H�t���:!������B��!�<��HB�5��-r�r�`y@+����-\�qoi�۠ c�{LI��I�}?wЍ՚{���bɌ&�Z�f���EJRj�1@�N��b֗@���¹tX�~O�_;H�%D4��ϐ�B0VSPO�P�(W6E�d�j��z�I�4���DV���Z>E���_�XX[�o�f��#Hd��w2A��S��2�NW�[�i�#%��Wr\�dh�K1>���g�P_�G�i����+���"����1��\�2�C'
ȗ�V8�VD+�iG԰Q��l����:>Lg����ב�;�*����[��D��r�_Y݉�5l��
�&�t�k��� �(��nƕ��G6��3�iW�b����%ݮ�D;d�A���A8�nnL����:�}����&8p����l��$�w�9�3�;��'ʭ����@�Y�̏��>$�AYtX����獴���2��K���:���ic�Tk���ʚi����E4��[���Q��b����f,���'=T`^�ۊ����������l9�}��KM=T��������\�*j���U��8$��k㒌��Š�10.O{��pu�.0���GY����&Vi�@[mG���'�Yù�Na�!����ĳ��蔚�ޗ3�G���8���p�]���o�S���j�v�o��g�L�{���o�e�x���{�\��,Z��#�|�a��E/��:���<��Fu ?Z���`�La(���t�5��m�T�\m�P4Womx^�5yB,6���=GgJ&W���uK��Y*�⌥2�\G,|�@0��S������9MJA�p�XP���RW~c����M?$6���п����&h�%��܋���5�����F]�L:�G���L�X�_X��bRW0E�n�F�J	� ��O�4}I��k�^��r��l�K����
K��k�# �s!��K6�k����\I�����nN$�GY����V�s.��� ��.�B��+��$saxir��۔`c�i¦���@��du=[�;�V��9�E��d~�(���6lwp�K�y8�B���P���O���m�!���RK7�v�|&C.�)Sq� p-,R�kS���>��C���V,ݙ&��>^]�K`㡋8v�'��I����nwsP�-�mfp���s?A�Q��4Z5B�%�wA��@SM�]gA��%��]pNp&ٯGЀ�70�����yÂM�̳d�x�a�<�i�>ۛ�f����Y�k8����/�\m�JAY��0���Wj�(���4�rLj_Y'@D�V���`��FX�ۨe�!E���H��"lZkd�%����z��ɘ��gʒ�'%�l�[�ͲZ�]�\�y�O��<�� ї� ���\�"�3oKlT�Z�꾍�� N����c��r�f���1!�	ԩ$鐊]�M�k���%'OPWT�m��C�m�-Ä�I���!�c��t.b�	s�CE:G�"O]U�}.gfuT佽���uv,k�a׬�$�$�́E8q/�'uh����cǰ"�ءȬ��[\i'���WyMu\�xc���M����O��k!8 �(PC=�4=Ƽ��s� Ӎ5�tWt;��ҳ��T�0�lr�
((�+B���"z�gU�����#(��XL�J$Q$;�.2�U�Dѵ������鵹��r�u�+M���!$a���F�F�v��$_"�4q/�"�!4�=�`��0���F�yN�u���u�[};>��9��i&�2��5p���k\���܌�TX���Ã�~t�7S�l�����W�/��T���	&�S���s�NQ���5�t���5��J���)�.7oP!��_�"��x��N��O�䅷d����,�.y�<3L9��DCð��괺���^2g�:k��N7��_N�R�l%�_��������X`�F�k���C��Vo�;`�KX�z���}-V���F_������˔"u�6e')�I=�ܼJDhB�� �(��|�є��a���F�%(��%
c'��9ڕ��
����U垈��	�b+n�\np�����m����b���H�2pPK��Hb��ۇ�w�&��l@���B�L���R0��Vg�� ^�E�	}�X�U~_��L��y���̲���ڝ#��'���m��;�	�B?@4�K�xveiWMv��!ܾ��h�#�a��a��F�v���|@_��r�MP�wq�k��S���Yk��n[���VUB�;�?����Ez��uh��dO�VY�67<�d�l�P� -����w��12����c��4~��E���.)�[���^��vs�Yr&=�}m`�Z�O��ɭ��VKA��*@G��}G�=\ T���3�Fn^E�	�Λ��{���P{�ZN�OϏ���*�P�6��f���*�ŀ3Y?�Ձn���S�\>@&�̝��xq���S���З�	b��6RLo���)��P�sɾ՘�N��;QE"��8��85��#�͍���� ���|r�5���	�n��@�	��^_��axi�{�y�?ko����޾�*��TI��1!��]*��a���)�����)-�F����
���S�vI�F�mӲ�{���I�$���]c���)Z�K�9}c�ۙ�yH��% i^)T__}�H��Z�����r�d�S�s�wϏ�e��d�����X�D�����t,W��;!� �.���|{�@hg`�����WP.�>ZI���ayI���޶����"
���Y/���W��O��ց�[0�r����6�u�-=9��q@�p\|e	���tF��Q��3��ˢ5������p-�c�#��7���m���R�{!�Et}^�ʴj�����ƆE�1l���:�?N$%�:�:LD���ȅ���I�?<��M����0�Лg�c���ɷ@����@I�k�*3�--��"gG<l�R]U��(Q+H�p#�����E��Dy���������dv�Y�P;��ܮ����R��ج�����A��2�9:)��ҾG��uE����|�f���7H�)ڪ�н�vs�@��V�Z�5�sJ�8�琒;�����I���U����=j�t�F;�;�nTkn�m_;�0+	a�G.R�l�+Z�qH5/x��� QboB�x������ӎK���QG�s�z��gn5�&]z�n�O����z��m�ـ�s��ѬW�ڀfW��#6D��W��z��<��vկ��K}�{��(��;��PU[�j=� �`ə�e�x�f:�'h<�Σ�K(Y��/���:���e1�-�uY��#�,�_P���D���
�����蜫۫M�I�k�9�r�|N��������ZO1��W�gg���?|v�E�0F����ʾY�d`^��j�ve_�(_��q
�V[G�� :��T�g3�T6�g�U`q���� RH��	(ɝ�$x�&uH�*'���g
�D�\���XO?���.��ۥF�������U�;$�����\3S���<�W&�hVM\�J�_�L2wt�A4+bvsߍ�Rq�G,T)!
@��c0�b�j$f�����ì�>����Ҕ�)�����f]·�
�{{���%��x���l��Q����Z�k�*�&;���ʚ�>�Ed�	���5�=ڡ��GI_;������ z�Q5�Z��Q�����ڔ�Kk'Vw\�w�8U��mT�����e��:UL�|3�J�rSBd&��U	
�x��0L��7�'�$~\�(P�FE���.$l����5�#�L��5�k��I&�d�%�::����'_�Y�]��D�������LI��v!��]��X.j���ƭ�;���1 L�W��<�����g�lG|�p[��˿0�P;	L���gǝ=��e�9�ɯ@4�?tu)�ڬ��C���!�䜌��_9��!��������s�{˼s\�s��2�4����-o��3r�*��I�k�]�Uy�/~)F���9/�D"_������{V:>o� dr�{�j�lo9x~�C�q��x-s{.�Zc�b�R�G�ߖ��G��`B����	��,ڽ|ѓ�5K��8ʮ�4���F׋i�mɅxR��:M�Ǒw��P����W��hv�ϧl�^��7��OPc�g��qp�S��PQ���U>9y�?�?/#�5�x=�a��^�s�X�ɢ^M\�r�x�xE���U%��*P��&
n��Vǐ����m�q�f���|N���<�&��<�|��7��D��؋��8�]�;��Yg�܋��E�ѯbp��KD�V��3�up��C�%�sAp�̭�:.��5j�+G��Ϣw�)1>�#��JR�kpZ��n�Β(�\$d@�k�����9M�bE���������8kV�߮"�R�s�h'Ѝ����'E�t�[^L�"��dEŻr�����*:�Ƅ�P=��T�Ь,p~��t9�5>����r�rr^��(�x��&R��@6��ߛ�k�6k�C�u��b�&�m�7�><g�u�Nb/ը��&#�ѣPhw�$�B%3���t��慒dÓaW���46*��S���#fQǡ?�v��JA�~���,��7��A����>]��Ѣ�u��'Z�H;ԅE:~�㲤RQEp,��sE����
�;ZG�MN�y}_�v>�?[�(���{�p�&3C4���5�);h{©�Ζ�d۫�]��j���e^�A�%�1�]�E��\�R{�[P�v�M��y�E�iҜu����1
��&�Th�[��;��mm�����2_<��6�W(�i��6.ǝf��Y]F�A�dE�ia�JDy�gi����xYf�&s�����v�a� 9[̞�F�V*�:Эu�X\���d�9��ⳬ�g�ϩ3���E4U���M7/�ނ�n�_�J�ZnJ9��(�f�{ ��4Г ��X�_�3��{4��43�V��-�l
��k*.�<2����lP�(�<��,�<s�*}�����}����B���ˀ	�~�[b�}��GX@H:u���t��YF��5���}�1�n�i�Tkt96�0�WI�`�RK�\���&��b�%ق�3�׸�ٲa����8�c���n����'Ӌ&Q?Xc�Oѵ3��o�4&)���ōi�
9CA��Xn���)��p��a*�>\�_���&��?�v`^��u֥�۫�����b�u5��]'������(Ӵ�1L� oS}`H��T�?dq=��n���vQ�3
~�<�5���S���rE����I�&�u qP��������u����8�H�>���5n6DhʯF<�{���i	��W�G8�q��,������&h�nk��4�n�����~��i�:'�&Z�(�ޢM�&~��<����cs=��|aLA��E��b�9�j��*qeub%\��H>!��تE���"��H�M����.!�-Y-/�N���(�Y�>it,BnK�o� "gZ����YQ��(��
���xw3�"����A��v������:0��)��>�S��G$��㦁l3QͰ���%$�|���;��6{�!�?��P�P��u�2$�5A>ZΛa��ln%F���CdR\�� Z�~,��]9Yq3o� ~�=��k���G�{��4�3�n���C7�B0���~��1t�<�;%�p.!�KF������8���-=ڒ��S��~��z26[+*/͇���C����`Y�.y�L�[E�ˁ)���>D��4B�.u�����Qw�ՊU-$�X#I���)3 <逸+�ȡ�#|�d�w�f���K>�bV(ɽ���ߵ���ӑv,z@�5ԭ���!�1S1�X�����X�
�餜*���5���!����V�[3)�%O����پT�'ǒ��*�n	8h�_\�W����sb9u�V�g����y��j�9K������f�+��`d)�F+��a��za��F�3�(q`�6���-|��@�	b��Ԙ�p�[c淥nm������㐁DE�s� �[5���r�hl�Џ!�|Q���������d� �`��p�)���Fpp>�*�J��W��%O�6	fS�~>m��,��FCRKk�)U�լ�H�}�|��c6	m����5��0��nJe�y{��6�M��(����w�ÐʂmI^�V �f���d��mg��|�����|��@�~�E5�7;eu�,��r��m�PEx�'c������f�VM����!�� �`��M��"+b��vREH&9o#��coBt��X�V�*�v�,� \1J�»H�#�D����~���
5�]6���_]Y�Hej<?@���#۟��1�:��K��9��Li�c��^��-=�/�{N@Hn�*� l@��ә �jl�A�D&��*AD? �'�W�&T'I#�Й��?8��>�f��3��ᰒ'����[������.�n�B�/{�/!B�čr�̡�ƥ��y�%; [��f�I�n;)�U�K|����X�6���L�7M2�h�&#ď�޳��4_�Sݵ�^E�%�N���']�!Ñ�c(CƧ��Q�}*�E�S�nh2T��8��끠k����@|�����Ў^�!ԘF^�M�AXktI�� �v"������CN7�v�ȱ��q�ϑQ�Wh��Ƈ�	c��b�9�� lҬ?p�H�l�XEZ)����*d�=aU�\)�/�H ���p���4�l��=�ߥ�M�E��M`x��/�sfe� ~5(�Z~����~�,&�x`>�瘏����-�/��#z�^�M��5��}\�K�gy5��8�m�x-�@�y܇Ӿ�L��L�GRrJKe�8,X�!4i�b���E���|y���K�wSX��4�*~HB�,_dp0���2�L:��j)5��G�e�܋[���Z$Xl�d�,9��V���3�:Xͅ?��0��}b�ͻU�^#|/���M�W�v2�Z�:�E �~�� C;p~��c*>iCzu_4�g�o�\���_9O����� �,�Gj"/�x{ë��O����D���:�uҎ��S��}��i��kܺ�̲7Si��'�ȾG����S?�%��r�"�rI��Y��Kcۗ��pgh��̕��4���T��s;�l����<������r�N(�OPEI Hj��l��#��,����Mb�0�K`L�r�ı_D��R�Փ䜊����+Ikз3�mf?la��)8�2P����[���?G=r1ܸtH��Ag"`p�h�75�˸�G�� s:�H[�IZ�w���E��)_�9q��G�\[x����u��H!M���t�"Q�P�{ܗǩa0+^�/�4�)�v�Z��O�i��RIf�z�2�??��Ez�,��@�;�Z[�=��(f�m����^�y�a�֫Ay� �1���)[����39�����k������
��b�w:�����QE���/AU��Ԭ|X:��D:�;L�%Z�jL�~^��Ժ���ή�1(���G\ ��)\b�����?�Aǔ+���C7��Nwq�K�3C��;J��g��S��a�';Q�9V�!ǳ��'U]<j�sŠ"E�Ľ�D�Ժ������NV�+�P:+���ċ��X���cqbX���p�Äd��g��BT7E�K���'�V)�Wޔ�!�	)1�m"�*����A!��%��P0�P�@�' �[�V0�Jc�	N��ц���+��z����q�'���L����e��/��S�sLȷ!�������U��f�����NI$o�_�l�!֗��b��}��qP�=W+FX][Rn*�u/t��7���6-����|.�a�АH�<�P���'G�(��P]J�(N ;�o��Ћ��S.A�s^*�]��`�}�7�O)8,�_����^�]D.	\3a^Hf��:�,���a��R�oϧ����:<� g ;kh�w	���g_��Ќ�	l#�V���M�3��i��\ۧ�>PݝemJ0_Z[��:T}a�F����u�Ү�#��Xą9��v���0Q���P�/:b��[E�� � UcԍE8�,ɫ.��,da��F�xP�v�U� �9a����w� ��wT'c����`���l.^�&mn�avsb��O�nƥ��P�A�N��ܻ���j��	���Љ2N����琇u�sO``��_�3_�?��G+�c	�e��1#��犮��	8 ^��r�Bs��~(��Ҫ�#�?ﳾsh�y�Ҭ�L�b���_�n������G��L�;�������1(�
��fes[6pS�P�����^z@�C#�錥�Ps��G��9'*�M���7'�l����Lv�W͓2����s��Ɛ㶶:���q���t�ćؿ��4�du8�+u� ��7� y���K���j���!8���5A;���hAȥ�ʟI�v1�q')��!v|yS���@G��븄c� �f.��EQ��ϰ��az��H^jR.��a���V��zZiMk�4l�Q��X��o�ax]��n:LǊr$�ϨI��$���PY	��z34���296���mG��If#�� CoϜ{��\ r�rO�o����4��/�('9$$������*\YD�����Ĕ.tx����0R�{����<hܫ*�yBR��/�ۣc����FY������Pn&'9��I���;hy;�ќ�GI:��Fn��}��*
qP v{L�l��zf�j��jy�^s�O,�� ��
vKx�-���2Xn#�=ތ��f*t5;�"{֍(��)��}��(;�3�)x(�le�|�FS�f��:�g�	T��ͅa������ɬ��P,+|����e5���
C�0́:���>�S��K-��ɍ����C�d�z�w�.`��L��t^��u�e�m����<�\s?�: �f�SfHn�~�]H��3 ���[#��@o����$�̛u��c��AK�d���h�^
�m/|HB	vw)������7�B�7����/��h^k�%�,�h
f�;�ѕh"�@��\�4]�.C��K��-���>�6��T0��X�y��l {Iy���X&�D������u���e�!�������e�{9!0��L1�	����m���������{J�Jz؆��k���h�����B�Q��/�.��c��o�?�艅&���p"�!�=���8*<�xO`����k���7o���o3>�6t�M��8��^v�	$�s��nw�^$$�B)��j�̚�{Ǯ�p�|�U�f��Q�E����q�g��#��F~`�!0�{1�sI���^\~]�b"��r筂�g#>�ڐR톚NΝVM
����{�+�$��w`�m=D��T��c*��	�F%��-�\D?�ޔ��gi�G��5�X���^:�s����ב��%;1�P���9�p�1j��S�&�z�B���3�y\�h�Ե�Kwkz�c��#/�f��W5,b"���pք���I���<T�GO��Z����^6�x�eǳL(�&����F�wĊ���5�M�N�tf�~@�MǙ�:�,��l�(��x�k��ȭ��g���	��5������\����JR)��Y��	|P��풞{�	w��O�c 427R/�B����ͤ�U�� !rL6�
�K��/���v��l<�e�)�|a��̳��o��9�T�O�kGh~'T:E+��С+^|=��������{5<���X��xU�̃%�=���zf5�Y�#�3D��^����d�Ҽ��2��x����]�0�%$�e��ZI�!�v\��,���Q�@� ��5�����
Z�.O���C�hay�?GM7�3S��byg1�5G�7�&C��=`�/�nk牄L�����T�W*GR��εx:_�4 g�TG%
��왼b��E�G7�]P�>������ޜS�ǃ>:�"�c�fp�%��z��υ�9�	�k-�� �����|{@Olݸ����Z��<�bJ��)n�����y/"6#Xh��+[?�$_Wkk��ž@�������j2"�$R�!lG�<J��*�!���{�o�,�s:����<}ʾ6�՟�Y������Eؔ��a,�sh�M����C��VqT�T�?E*��MA�����>�����a�+IM�qC�^{w'y�0>�8��õ���#]=��bh���(\�+2䨺⹭c:�O0薇Q�����'�W���s�o��%���?p%���(�h�d��k*D��n���F�/�Gny9Ћ�'V����������`~�K� �ji�[g00� L�+Y�@O3���n���7|�9j1IIoUDe�*�Q�?SFs�����ǆ{��;=-B#"y�Į0^�X�w!.��]Bm˱;���I�3���k�y��"��q���>{l�
�Ὺ؏���R�5��J-�:�o���L�<ZsG�=�"
Y��2�me�Rk�8A�&�=(a�YS)ّp����>�z�`k]8��5��Zk�_ކ��wg�ny|���9�6�fҠ�J�z��ӓӼ�bᣬB5�X�[��UD�nR��7RM;ϡ�-�&x0��0���jEpY6�����s�14e �e�+���&�����A���{�ę�R�NH�]��	M�ph�?̓2n���ė4�+:����^/i����|SY�Ƞ|�L��G2��.�6��s#�Kd4_��I��`.�J̶D�M|�P��n^�����S��8[L�(q�ò������c$�g�ABbNgw�ݱ�~�Mi��R^DrjN����
yGJ�v�lF� ���YE΅(�l&�X��\u)_����o,"E���%@�f�]	�U7�ԣq��Y�����C�8Ki#UXI���LCl���5>������DĨ��{^L=��k�bC
F�W#N�T�ͽ.�?�}�ElS�lH��9���v��baVP8�s�o#�S($�*�]�V�p����m��w0�nn��l��Fo�h�q<������r2UU��1ihj�n.��d}�6��͠-��Q������]����f��k�� q���_eH��L�{��+���$"{l�(��r�� "	QW|�/b(�61'���$54��Fp!�C#�Q�o�������qQ���>W�$���cl!����W�4��
�NàJ=��Aǹ�}�
-uٚń��I�@����	>X�BP��P?�tA��j۰ok�I;���9�D� \OP�?y~G+o�����c^ķ�K���3����$uK#�#s���dd���}��ƗR�mJyK*��t����&�A +��y�Ma���3G����Pb�"�f��TL��L�I|�+?Q����ʁ^Di~�&�+�#�?E�a˛I�2��q�F�0���/\m�ܕ��l���_�O��G���/g��<�p��[+��Q
3	�BT)H%$����V��h������9�Ij\���e�����L��aP�N���y���������0L�9
$u.�Ɛ%ʕ����d��hS:�(bY�w���;W(	,&��T��l�N��^�8ܬWX�����G-��T'#���C�)�^���^,�C��:>��d�>u<!��@䋻dk�Z0�*y�ix)�$�Џ[8�$�]��Lb�vVc�]�':�-yb�ހ��w��Z�A/�î�X�G-_��X<[�d�7�Q	CėƗO>�=�S��=w���:6��M����sΚ}�&:sύ6�y������i��N�(d	�i{T�@K|�l�XJb"�$��cZz�4Կrm��k��H�,��y�/L�%;��Z(����JHQki񺶽�F{(#Wkb8�T�FK��W���s�a]~��Z��o�˸��"�[��m�VQ��,І;U�Ŷ@���3"�ӭ��S�T��d�D�|�D8����Yr;��$���]�:e�Nu7�E%bTB{g$t��Ԡ&q`��n�h�����
b��*�3�W�ho��	CLj���ܳ["���`f�Z�G��2(_�nz�|ge����3N%-x�	��q��3N��9n	��_�d���Nۢyi��u#U�\�b�L�T�o�Jj���+IU@R濟c�0�t����)�7!���1=7[']u	��MD�#��:frV=E�X�!�����k%k�U�`@��`H%y�J<A=Q' )��K�
��dR�|����Os��2��&�I�W���{ L��.pm�4p����<��x�̐��A}�_p����o��3�ִ���a����tY��å�lM�����Q�R�Q�l%��ĕ%K�8���@4�R����еw|ۄ��k��������;�7�T�0�j)(3��~SZ7�
� y6N����n]A�x����\�eK��}<f!y�1w²���v�N?t���M�B<����W����Ǎ㺘�;��C���үQ�6�x�h�r"X䬰�;����B�E&=�V���<������Z#��vo�Ɗ��ڇ?;ê��:��=�����i�A��׼N��+H1Q�Q/�M���ߔ�`����#*�⢖���I�Z�2���)��)���.9�b���^O$^g��+.s��'�Gq/"TU�.���_z��,�q��3������  ����+�j_�u���8��&;��"�/*8�cr���o�⺄������Nj&fs�����dvӲdt��@r�����l��BT�8C�g��g�-3�����>�л��Ix��>BR�|y�x�2�����=�Z�c����:{
Wi�H��^�����Ҍ�O��	��ՁH��tg��Ed諹<��%�g��9v�����NȠ���4�_�&�(N6G"����_�(�[7���rjq����n��1ڕ����Ђ2�W%�^��!�,[I���TN ��U������'����������w��k���׈ ����G���++�S��X7� (�S��ۖ�ݾJ�����"pT�O2r�+�NՎ�ō�ׁ@D��o<p����t�V�&�ش:E����M�D�
��rhAҿ`⧓�y"P���o���AO@bv�D7:<����7&�I�hs���c��*oT�z���{�О��誺��f��+�i���30���K}H�L�4 ZS����/).OɼȇK?|c%k���)r`r!���IE�n㩀�]{�Tq�xޛ�\4XNC�k�Ŋc�'*�����)��L��(��Āɵ��C�	;��E���ɀ�%4��	N�y:���^�7<��*���[��,a�AT���="R�����&���t�}�2��!��.������W�*:��;��Y�[L&��DB�k��,��5���ҕ2-)�ԅEjK����rl�1zcܷ�$S8�;����T3�XĬ_6Bx ��z�m�F3S����=�e��;o�/��~U��(+Q��p��s�-ರ��%�򑘹�Kw�/�գ�${Ul�YQ�e�1z�L�~�"���ŸJV+�/���T�Kg��f-���q�rO�ZC,��$�;����;ScJ��n���:�K���5m�Q8�Mم�b�b�v���kP3¸	��%Y�ʈ��pwx�1��)-����ZE ,���꺼1��?�LP��;5���Z�X½b�г3�����0�=�=��J9��-agr�
7��J�M㜞�^9�㹬��wb�r���f��N��mRIu���5��5���8��E���.�`sE�0��Ұ�iK*9� &�Eu��*n�
�d�е<����I��4�JL����M�
X"��'��%Z������`U��1�Ò�H�Pk�N3�U�ǌ�h�a���laZ��ܬPe����dg���$4!9�����
9�1D%qx+᭖��ޅu��>6#�2�v��a���r�'��6��{,n�i>��N��E,��D?��Q&��s��j��ο�.P35��y˻�\��j������$X�mު�cR�UC����W5�5�hMS4{�	�����B� ~p�������-�?��F�-gRת��X����N[ƍ_�����2�T�K�����l�w�@̰��9��=W%������J��u&��CY?S��4xeg$��<��go�>"EȘ?���%�0�`f�A��O�Х[����}B������gn�NRF��<�*I��������� �k*�|��M�P�#���������nH�(��+����v��l?o>���ჰ��w�(���{�OyD��`�u�בֿ^!�F�Y�}��Ra��'�����~J�.�[���E9*�0�"o�C$�7S�Bң��.���x�bNg��=�����͌H�P[$��GhJ@�F�ʗ�/�F�-G����������[dS�4�FOY�����W�:k{��K!�ʻa��@���ӵ5�'�� 7kc�?E�gO��a	��Y�ͅ�h6�e�i�|�����.k��X�`�Rك�vǢ���wE&(>��D�*�M���h���B��Аs�G��X�pSZ�|o] 5p��� �Y�_PTd趆��&���A�g)�yCj��)L^y�$4��wmˁ��Z�C�"�Ϸ�y�H��Ro�5��`�Xěg�E�c䦹n�Q
��j,�*�7��L�-=�s�����U�|�d���ջr�anjc^^Y�����/�%݊�T\8��f{	�ƻ�{E9�:\����WE�51�4$he��զF'd�)�Y�O�UҸ��K��,���G` ��D����dGC���Ӎ�3�A��b&�i�}��dp?[yUC���e���j�	����v