��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&Y�%�ddؐ?t��5�O���Y�G�N�{����̀C�p���VSs�n��TV�j���eRV,HW�r��9 b�V3I�ˡ���`��`,��9������������H�L|�*���U�;�'hMC��ߘ1�J���i�{�0Җ��ʩ���
�����l�(+!P�C�K�|�$lxd��\.�۶/�b����y�XV퇻��X#P�k��em��LXv�*Vڰ�k���E�`�3��%l��E����C��8�k�_z���!� ���B����3eؤa�� #'���+`�$�+~����HR��.�JN1�N�����+�&x� g�a�0���b"˭V v��G���z�ܼ����P�Yl ��|��V߭HD
x&X�C.Oui���e��֒q�p�+�2i��O>�=����Q�6��=��(k��W������^���Z��ɴ��v�����(�BZ�KSGf�-m^Tc�P�{c�jS�cV��䰍	�
�V��i�e�x�`US��p�.�زZ=I(�V5���8��_��XC�{ ���e�n���e�K�Zm�Q�nL�hn�i��]xc�5��C�:���$��Q��H�ɿy!� Y�H���!5՟IóofM�.��,�^�xrގ�{Ў�	)v�_6*E�39noZ3c����aӬ���GcI�u����J�ǰ5wq�0z��8���N��Tæ�Ϳ��\��ǅn�	i�ޱ:ڗ��nГz{?6^Z����y�טy��Q�kD ����h��~o�"Օ��-��B����4�A�b�a&1_�Ҹ:�
`�j��i���l!<b�r��JÖrd� �`c��L��ߙʔ؈s�R��6�e�Gs3��LA{���A����4�&a�����Q��A�w�b�<��� 'Pش���q��x�	Nȷ��W�����#|�m��I��G�V���Ȉ���+*��m�ĕ��Hz+�,��?��0|��5S����_[!,8z-�dN 2<��2_����=6Y~��.#GzZ���<�5�d�k@��D�י�"�/1�a���տ��mH��ҕ�5�E���\M�<�ּ�����VWυ%�Z��/#�}�y��!�7ʫ��l�S<JZ`���lzP ��օ_[�	�?���=���M��k���S]H��8��1��(M�w�6��b�Ԉ@��@\�����[����O\)ެݡ����`/&(�b/�I�ә��7�t��a	/���+��z F�PlFȖ��^�@jW��T�j~AG��C����T#2z<�\��!���a�����EmM��S�Vr�F������-����e�k�#��P��1<rs�>�P@�F��4����(O���Z�2kJ�ia;x�����A�rM?v�Z�P�ϋ���F)j��4Pe%�[���cU+S��������I1���Z@���(Ɩ�%�P�+��S�9w�]\�"�����-�\����iRlx�txrO��=�[�>e�iH&�J�O�z��Qo�
�v%�%�nszb��.�,.��A��h��"�/1C��S�:�~�y��� �X4��rqX|d����}H��JM�
���$+B��g���3.��>�8�������>c$��3�� ���v�D�i��T�G�e�y$[JH܁����+��L����<��TS���@=LV���������iæ��K�3,c=
�~�I���q�ċD��t��v\��nĬ���; �X�&Ye�15����S+S��8���L���[�" ��~�T�.ѓ��[獥�T*�Fx�� aC8�E�1� �Jk�n�n�"+M���\3��n��9k<�g=��N݇�k�f�k7���>ޏ�-��A94?��>pծd����D�AT�v��`�d��:2L��@���l f�|G,4��)a� ��۔}_,��]�G�g�&,������p�v��rиȠ5s�L.�h�%*��I��d�L�{8�U�!�ߌ=�}(�Dq$$u��yh?$ȶ�����hL�ҡ���g�$ũӖ!M�5y�~�0 �C�?��i���FH?�bq���� �} ^b�&>���J���za�L��ܬJ�"?��d{�rl�%4��)�gj���� ���S:Lz넥�?�OĪ8ǾxH��w�+�Q�ݶ������m�H�����"��y�e� +x��;�;�~[S���K�ʌ�؉��q� �b��6 �ǹ�YKa��K�Ml�h�A�0���"Zh�?��#P����W{�N��N��Zc �s����X��1�������+m�������n�u(<{��G���Hӏ�[�y
��o&�X�Bk�p�4������gJ�?��6\b	˚�K/�v��f�0jn�Z�/��U�M�G��R'�i?�4�G#nv@-ȡ@��X����J�<c��'�3TeTu>�xF�!V�;���8�U�� ���^�S�$|�e$K�L�<x����h���&M�Ԫ7�O������#�uR�9�˯Ud$(�Z� �)jo<�*���,��o���$��C����衱
W)1��b���kF)'���]�|QH_���^G�1��ƋQ�,C��	\qfb�5~U��!Y\�-گ ��N�7��*1���w�'�����U��{m���0Gv&�S�}^��zvW>Y��P�Nd��{�����{���ܦM����xA:ߘ�c5�F6Dq�Z(�Ӯ��6V�s'����Asw���t�����H���Q�5
�7B�����ew���=Z���L��	�T�NS�[TY���G��Q�o�v��7�̇6�<Ø�nP�5T�Zg�jOy�E��K����;��x�+��n�bY_��0s�6$�F�O�2ɞB�}or�>�2�U�=��!X"���������C�ʼ�(�t=�к����v̢<�m񓷲��Nfv0DUf	ܲ����X�����O�����1�5������p��G@�^�c�R����O�A�����9oؓ��c�ҳ^t8`}�Ђ�����˃L���7�i�����B*�!/0� Y,U�è�T�C�3i��d�?��m��t�I�Ar��<k��e⋨��!���qG:��3�T���Ӥ��n0����O��� ��8Z+T�({ae�cq8�c{�ϣB!���KF��]��N���t5�ɘCp���Պ �{3�2t:��+�BӖ
�� «����8�5U����h�W�δ��Y!�$�>`U��
�i���s�%�� �pF��w��O�)����@Ҙ��%m������u�0��<H�P�]�]5'\�Ecw���=��@�<��_�P���SK�W(�p��`&\�M8L�O�q�SZ��]JA¸Vc{����?|�鐟Q��L7�6���q��`�����Ű�a��mzhQB��?O��=��Z��a�^*Mڛ��W���+�0ӗ�-�W���SUI�Γ�w�(,/54��J�Op廙���������Lı�qb>b��T.cK]}\��1,GL�H.��i*fR��>1���U�z_�G��jq�)��3=�
b�l�:�o�aT]�7��B�Y��K�J������p����ؚp�Q�C�>'�/0�s���vyl!+����Nn�����ݥ�}:?h_g�36B�>jN9ѩ��$a�c� s�H閄r�&h�P�7�x+Ưz�t�]���M�:&z��p�'����\��a�84Rs�*G��n)�ڵ��"��K"f"��W;���`��w��#�^ʵ{�t��TQdboZλWl����y?�z
��Ԟc��8������w�":cu�����j�i �9����l@x�Nj�z�	���D�J���^�bY��YY��7���8������O�6-2�F@�bc�����*��W�aw}�`�l���V�#ʏ;n��J�1��\Yt�� M����z�th�V�����`�Y�*�1�۬a�:�n{)V���!��i8�K�wm����9�wVjM��<���������%�s�G,���"5U�f�n[n��
_���K�eē��i�N�9�.�ڻ��j��.P�Yb\j~�#T)MN��j��pC�pu�l"�L]ba>�F.��}uE������>�J����w]&Ҩ����u��6�7\?��°���	�^R�⿩-t��n�?[�>��޸�^��1�����E���D�V�.vgNtքB!!�1ƞ]n��
<ց�D��}H�ߋ/�:�ӧ�TE�{A�L!��̖0�V9f?
ɘ�_M����H�RZF-f������<ο���luJ�Y4�X�R�w�)�Ag'�r	U��i)%�A`���ū*9�"��嵷V�U=�4#�e^9H��#	?����QI��-�Xݢ*:��}�r��I����"�g��Tz���`�M�rwwE���Q�!�8�HN�wͼ:R�%!��]ο���D�E�8:��������HP3�umQ�Ⱥ8ǘ�w�a�?��e�$��Hð�}f;�AfZ�� ظ:�wZbv��'����[����F�A4�Q�z��"Aw4\��/#��&A����D��?��r����YH�>Rl~�+�_�#���ޡ���è���#-L�	��APŢ��y��l<�k*��0�O1�����#�_ ?ӊ�&�Z���|{\6���@�#&,�;�}��ο����8�厣x� �]�=�ܶ0Y#z�>���Qb<���b���*Q����e<�~���(���������>ݲ�@�W�qG~�a�̻Q N��x�'vk	���&pM+�ӛK�~�cZFл��Ҟ�tP��x-�"��Ffq�`D����"���RU����TW�6xxL�2�J�w�h�:�X��k�^�![���Z̋��)6�_�x	]�.�^1"�"/����$���4�1��M�o���k����O>ۤ��6��[	sn��w�:�D���b�+FL�3�-�e|An�`7bcGm��v2�}�I���db�yy .P���S��B\�����4Vn�>��)dI/�슬�ՎӒ�a��5,K\�[�L�x2�7�la3ѝt0}�}e���_L��}Qq�}��/���`����!ѭ�!�&�u��-�4�G�w��&(����QY���9��"��d��� ;
{^$���7�~K7�~$��G�������z*eL�b�x���'fY�uW멒V�Ƃ��p��<�����D䠎gf;�2��+��>��?<�#��^����A�`��&���6x|+#녾��n!�U�=�
�ܤ��V�}��̓�bq6�@;��|�J���}�-�Z��Z�����8�u�����͹{�k6poUq{qi�_���d� D}a���u��W�uRZ�������W��C��d�x��S6��9�$���kB����-�`�tO��4����饸��M�P��܋���/����j�_}��Y�9�.` �u�R����D)6)�L���(�zB�e�/�m��W[��s�����6���u ��ȯf����2���Ņ�`:�3�W������S�E�¿ja@��?�ZeWU�~ DJ���W���^��9|;KM��<w�]rtX�|p�IJ���u�S� ��΀"B,����L)Bþ�l��zη	�b�'�����-�(�2Y'�� �hX�;V֗���2"s�1T����-85��0�RN��4�"�<�{o^x�dn��l�zG�u�Y1�f7�#Qn�����"6o��N�|�_V�.���)\I��j\f`y�M��}���A�w�� �Ӽ��\��Ԙ�F�f�mEq	_��ڽ1�D��M��Y��L�v�v=�Si�B]s��C!c�3C_�ҽI[L��R���+��i��c]�#�X8���
���I��|�KhM��c�z�헼�D��=����9^���2���_)j��8�L_�M�3�2Rǀ�(�m�-
O5*isxw^�.�>��x �CN�'TV	�"��V��9�I�`\�n]�i��v2�n��X�F�F��%}Y��[�N#b�$/��%�nWF�q ��5>�|��D�&��|L�b��\������P*X
^�w��cY i�� �:���s��v��U�r�-y ���Ϫ����ܱ���2�k�]�Q%kdr�Ո_��t��U/Y/u;=IZn��\u!�C��,?-g42��nM=�y,XR����D>f�F�O��.��Q���	o�`�[�C�f �+�?I��%tҝ$Һ.\v���p�.��G���)�4w�.��jhҙ��$�w,
;�B��?���ꭸ�D���A0���N�5:�Wc��џ����L���y7����̡����C:5Q��G�cs1�� :�ә�Y�v���^v��2tܱ���F�����]�(�rͤ%kA^+2sb!|s ?���K����L�It���"�5�����(E�'�i_��8��%?�Gt����zo�M�5>�����.��A�g�0����� Q�W���dd���۶�=������l��'��y��{|�X3�(�{��u��QE�͒nb�����:�s8�8Y����B!�q&�+�cB�H�!8��e�M���m�PcVu��ʒQ5� �'*�����`�*��mu�4K��4S�[iZ��
bE9*�9��Ӱ1§
�7ߘ��o���>D�0_��)n��OhmUl�Rl�[d_�7���~h��'Ѥ�����i�u�����#e�KU;�ة���f��F�$���4��C���c���\Z����ap4�Em��eX�53��5�wo楇Q�vd��B�^�T@��ɗU�A4�zy@���4����� Y,��jAP_�3�=0j���_>(dݝ{�=j�����Xg����s��>2ē���̍}Gs�U�e������Gh�G�V�$L<�#-��Z���yx�\m'��._OsGC����;܄9kz~8N���,,ލ�z�֕��|�����h1E��h����.]�]3�a�WLu�@��3A�cG�;����Ōv\�\A�HSY�-���������1���t���އ��3��R<k�0q7�mɶBTE�����92��}��c�pt����Mus����d�N�y�'���[�W�Ɋ�c'o?�	 �d
!�N��5�[�R�*��P9����ʳ���ǔ�'���t|�E@w#��Y�"�Qg(���@��s���E��#֮��KR���`.�s��<����D�T���O+���H��6'��p|V�����I4�<�,+����`�b��	{K��qz�� ڻeVm>�+��C+�!�����Ϯ��em���k�d���]2��ţD��o����k�����u%�H�sF(��P�L�R��H��c\r'J�_>�	A#�Q��,��F�2T��
���P+�B�4��
�h��GUN`�"%(}xp��?'��8���OJ3��10g�;�nM���q�����E�����%�mX|�,ń^�s����ǻ~%.?P�G�xA%_W����[�t�.��O�&ֱ2"�B^q�8�4({.�V�8x�����n�	j<=o�3���`��~�_����Q�8���[�{�����<��}�I��#LW�AA�m_��Ԁ»��ª3s�F��B]#��g-?T����qR9�lEӨkB���%X�KY'��(0�1C�C�j߯祈�)�j²��

 v���
�s�G��=�:_7R�����
w:����i��'�uI�E��ИmV�O1�*���{��7��阧�ds4ے.5WLR|���j��X�;!u�|.EM�����0��=���Ţ}Ā��'q��UE�EU�Z��Z{�	粑$�`F�V���r��[���f���:X��8�PM��'Zq����ɿ��ȶ������V;�փ�L��k�0Hz*ZʎڦLў����"[f�׌��I�<٩q�*EꝯoU������H
"�{��M��v�βX/��Af!EE������b*�;M}�̑q_r�샋I�$�M�;�ՕɄ��&�6,Q������3�w�
�W��%�j��l5r�L�O3�gn�|���[�9h�Q��[�}FGv��-��EJ��")
�|"�ˀ2m-���`��Eh�Ú��&�E�����c�o��L����ek�~���`�uR����j4�6��I�@��ｶ���|G��d����G���d�+�?ց%F�v<v/�y�����L���{,H�l�\e[����p��߬\duƅ���9r+��Gl;�2.�Z��(&x�2W�/=�'[����Ut3��0mg$u�b��?U�a1kY������.�W�����rJ=�4�t�D��X]&BϾ<?��j}jnX��	�ku�O����u�Ӏ8+L=7xM(��l�9��D�Ϭ�+��3
L��c�O����5��d]��+z��C[�1��ͫ�N�~�����_1-hɹ��f���2��XhV�Tk�P��Q'oW�=N�ʶ�U4���J�*k叉�&ަ:d���ͤ�[8{�Xn9��} b���=�0�긛V�?��
!Mu��G-�����!�ca���n6����k�m�\�+��n3�[��a.<��%u�"6ׁ���7������^�S�����y� ��E�de�w�b�O��A"���b�IwF�k��-��Q�[\�;ڞ����	��p�����	t:��z^v�o>��)�	��SI������+�~�r�V���ޝՉ&�"��k�_�����u��P��%N��/�򑌲:�?_��R������T�z��k� � ,�E��ΪȬT�\N�Fo�ƙ�0��"�V������"��4�YV�ovH��{����Ԏ\��X}��Fl;� �n�1G{��h�*��IBt.�x|�LF��9�^ D$j|a�fӯ�%u>3gL+j����J����a� ��f5���f�[�cXȦr��g��؂=	E75�<q��s����������Z����<��J��al{��5�<i�j�3�w+hP7�T�dS���^���P�>.7]����2D�;a6��d�vT�<9վ~� �E��0`��OV�7^��t�S�G��