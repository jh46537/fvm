��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���^�T-��!#��S��v˲B�Z�!Fz'����tP&.J��(�S���t���,�б;�n������I���х{g�25K��U	L�m�5=N�4/ԣP3�3}��ϝ��?=r2���nQ�tVu���3�1���AE�~�x�(d���/����'|�aTr`؍lT�e�L3cdB��e�US}��1y�R/��e�ë���L�`�MT��MG��l����q�@���Bx�nV �s/���Wv �gR����κF<�{%��Vot�y �yN3���X�-6w���|��ߖY�G�#3��)�M�3��ueHM�H`"zG.ͼ^ZG.���3ދ�>咒Y�Y�5���"�vաZ�� $���j������l5t��Y�"����(KC�pf�hUuM�����lcb�d�L��n)nJ��E�q̟����	S�*����k��~��Wsh
�����D-��W|�,	�:��k<(P���1	����1㶞_Ԇ��n��\����c`���沯L>���1�H���!Y�6��o�%����"�B�� ���Ii�2�+-�ͽ�iL�}�8E�?��7��ɑܽ��$����ړ�����$N��S������r����2K�J��|'ҿ�9�e�c�-,D��	������Q����_��#�HK[�u�0F�L��lI�q�xe-�J�bۅ�K3LO��h�G:^�@e���x]-�/S��3I͖��Z����@�tv	��x�
��Ҵ����g���m``�!䢪�}UXCץ�:�q�e�_�d��b#(Ճi[�˗ܜ*-1|S _��k����kX �ϦG8`G�m\D �F���~p.[jk	!֠�!И6d��L%�\{Ѵ��x��������R�:ħ=i\LI�EV���qa���R���p��*�}(i�����1A���u�xmB8��]��;����z���	���Um��O�%�f�D���H�a~���%�;�M������F�C���)G����L*�Te��84m��C�[2v��43�N��'6;��4<r�-��!��q���fz��
F�p:n���m��U�늭C�ri�A�j$+�(%��myl���J<��H<L�lU�j�G~��]���6Dgx�V7Uo�7�K0n���z���`�}�*t�7�2M�
5>��]&�gBa�i����iǊ��Ys��������h;��H�4��hŧZ���/l���N�C�F13����T"&	!2.��%d�G�k��w,�Δg�aw�X�baRɥ�{���*��7�M�q 3B	��q���q 7̭o��
�V`"�	[��
����؛���J�E?#�^�DC���|��^��C�qn�9u�����g��w;%���rw����T6
�a�0�(2�rm���M�pY y�:_�TK���P���w�!��� e�K�Y��]��Qի���Ѳۢ<x�>.�>���2�*�
>�j��wOc�1c�[�"��77O�s�e#{��yD�KE-,j����%���%���d�N\���G�*wF�DsF�3�rØHzO�97�N��w�>Z�TD�-͵\�p�q������ ���X�4:�����Q���۩Te���EH��g�j�҄:���2���I��Lc��*B.���w����