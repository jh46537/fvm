��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0����>�P@�:���{������^;{�N�9����xMZ�*�����B�������j��v�1�O��{��U�K,2�(��b
lG�m� ����e2h٠�������@�@��bSK���.��_B��^i��
�o����������ѸLY'Z:������%���<ܯČ�8;�e���>�b��*'�Z�f���F����}$�$+D,+2)Z�|��4\r"n��#��cB�yy]��K��a�,/�+m*�?}X;��x�'�m�oS�*Q�E7����??���[9�����P����n����Nݕ�:��b�]�Q��r?�:m�I���h9�vf�����+ˡ��(�M�3�;�s������5N|�B�]b	M�Kf��p���<m�����FC���������6'��7uJLc�'���Z��R�!Z�6�S�+,2���ʓ���H0��i	w%�ԍc���#n�sa�Eh�@�VQՕ�/;煟���\!��z�/*\���vE#�cz2�a?�K4/Y�D0�g~ˬ��:���l�����Ne��pxE݊&�E�.�E����Bk밑�/�f:�њD�2wF��vn\�i>~	�s�3�r̷�@s=V�xn�2��q���k���e�,�"��Z&�Md�q2� 4XG���׬��R=����������� g�݌�X�*�1�Q]�'�XkbF.xܿC�ue]��1�r>�����<~'��?��A+���ÒL��j�4J��g�'�v3��-
��HY�Rp����J�%�<_����9�����f)�=�b��ۻG\��)��T�.��j��wUG4��h����]��9��لf���ES��3�ݻ6�Rk�Cvj�2ux�ڗ�U�@�7e�z���*-�ۯ�Hl�ݑG6�w������RJ~R�X��A�h���
I9��<������ȨG���r5�Z`����%������Ҏ:�a�{̘(��d2aI!P��/�=F�>�;U[�I����U�\5�rT,�S�����Qb6D΃rxD�k�՞`s�|��1�͉�'z��>$���V��e�G�%�������u��']��Q����"�-9	��2	��?c�
U^GD� �C���A�0��a��bd����
���K���J4��B��8�ͤ���ܸ�����#��
�4�K��pR�Wf���"}����%$��8��q(6�4 �~JAj�3>�oN>(>�L��/uc���y����6����ss� ������6Vڎ��#C�+�y`At�
{qs�FG��6<��ɢ�%�����*��=cA�a���(շ�w�=���c�$��yZ}]�k����8�sJC����`�%
�9����x@}?�9�	�\7E[;p�b�9�/��Dy�9u��d3�[4�5O=C�Fnv�vۡVai��_<��-��K��]Ns����W=ꎃ���̚PҦ�K[f�IsDr�jҼ�-A� �A�fk�1������(�X��?�U�З���W��e��J4�2ě��f�c�1��1�L��=?Xt���� Q�
�o�GI����$@�#:]��	�:i�s9-�l��"��j]{x�BMd�%��}��5x7;,����d]�B!$�Ӕ��W7RQ��F�\Kɹ��҉40ZU����7������m׷
{]ϘK��g�������B�(�-�`循�	�휒ퟹF�]sgQ0VB��P擓�������;B���d�ww5�T:���f�R����BT5�ʦ�6뱑	5��b�_��=Me���KZE��+7H����*Tuc/B9��C�o?�R�W&G�  ������
�#��V\n��M�z*�����eH.�M� �f�Eq�C^��*�U0��y ?���2�K����;z�A>�Dkv�`��yZ�PJB���w?L*|ᵑ�q�VZu�@�R�Y~{/�
E��o�����T�YA��p�j��U������U���$Hj.q�EǢ��L'�����hqy����J�2F��P2�C�)�	[�ڵB�u�u�$�FD�8=PCF����� �sx��0J�x��N0a2�r�_n~ƞ��D��h�S�#T��R<	e��rS|��w>M