��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�k*b���f^��g�{u;��X�+�w�O�%�Z��0w$T����'籥�� ���xO�-�ՒL�z3�̚4�."�f����u@r���l�|h�`(<w<��+�s��[�n����m�1�Z@6L���e�D���J_�ݦ5�1�Ź��@����
��s�/�y[?�L�灂��v�<�i��E�}ԽX�U��P��n��b?�X����fP����� ���@�vͥȼΩv���I����L�!��7����	N�2�)�]:Z�0�p�p��E.��О>?2!�����U8��IԎ��K~���`�F�-���ٝ�GFxW����&3���'��0)�h{���?<�͡b�M�f�\�U�W����)�G�^YD���Vpў��\aw����A:k 07��;��Gh�_�v�fPL� ��`}O�ϖ�g?H[�C:������1]�p�ΰH�z��'Ӵ:6K�uÝOF�2(I����x�W1��7�N� ��u:Pަ�YqI�I�h��5c�I��4�$��L��:u��#�� ��'= �?g�ZQ�tV�v�Z|�1�r�![D
AŃl�)�҈qN�v3�.�����cN�C��l�&{���(
F0�t�� ��H���o��+e]�� ]e��ԣ�7��6��$��l# |($#�	tJ���Nq�����ɗ6�G����q��7���,^c��*R��*�;`�?���� K����%���F}�v��[Pv伂��_d9��H����2�TZ]�D�/������i�\�����ABA ����6I���fr��~˕9ڛ01�0��V�F~�v�cT���Â�Q�J��S����/
$Ҕu+��<�;N�!c�Y���F�kdvQ������_���v��ޛ�c�:�-�A,���ݤv�i�����Ń�F���DE�#�����U{U��W����خ1ќԨ�U{��]%ZJ��{��d:]�a�i�l������Y��g2O�&mPX��o]Y�qe��{��}�0��w;��R
�Q��u�5���
*�|W ҅jˌ����I�7DLYC�/^:Ȝ+��f~2�:��i[l���Ew����\p.0�}��5/���w
`�:�,ʮ<����c�c"�C�XAK{�\��ѳ8#:��=�*w��1,dꃍ+1QI=��'[���`	e�|-���r�+&ʲ��)ɫ����*R�a,
g&G�<:������f�ㇰ".-����E�����\Z����aQ�s'D[���Ͻ����s/���nص���`O����*����^O��H}�Ǐ|��l4	�f�K�H-�a)��:�»����Kp�q��0^R%^�5�զ܉Z�Ɯ3s�t�F��.�	r	��Z��i������~W���4s����]�W�f�2�YT�:����*X8e#e��-��i�8`�����)t$�����l?od��d�kZ�i�K24�L*��!҄��85��,�j�-�N\z�-����ؿ㈋{�KK��1$�a�R��4\�N����.�� JZ��&��K?m{�Ft��Hİ�KMH� �f+�'���{�w+�s{�:��;�$6bX̏,�FJ�<��ͅ]�m�s�w�N��D��˙��lJ��Z4M�[��]�`̵��J��