��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQl�E��*���7��ܽ�s[0�ab\�H�&  e�����7��]%A6�~��KJ
�T�Q	���}Ú+Y����V�ߗ�@n�����[���L^��[L�4ROm>FqF��Ļ�{b�P{�1��y⊮\�!k��b���%�4���~�Ӡ4��tφ�_��p��)޲�a�_��h��iX�D^`:\�T����(\ˁ2��-�x]ɾM�1��I���G����{����L۳h�נ��+�T|[�6�Z��x��q�#z�;[���T���ļ�eĪ�g�ۺϒ+h��5��$��0b����$L����I�yo����-���:MT�%���C{+�X=��w���O��ʒX@�0ԝB��b�4�M�E�~@
�6�a
~��R,v䙦(�,�,�|�uˌ���'�K�<�熿��'b�֛K�K'���UQ�2���Z~�u�;�zH�r�].��_���3_/F�^2�V�Ow� ݔ�_�z�f�`�M�SI�	��w�Pi�E�J#�'��"	�v� �z�0�w�ꭗi�x�#���ڀ��g��%��.��;��4�k%fkw��w�Ay����gu�|���9�Æ�{40d@����F���v[�A�DK�~��hK��A<e�<F���aw�M_����Q�G�u����z��(�R��=�����U��֫h����&x�hϯ#弪�Ƒf��ɸբ$�@�V�=D����~�¤�<rx�w���Z�8�͋ �������L����Vϭ����1S&V�fd�=�J�j�ks��٫䱖 �*�r��?��Ŏ��a�$t�B��~���d}�
 ���	� k��Y[���楦�������;�{,=�Bu���;r�1t3���}gX����[=�d��l�q��<\�m䫐92�bȖ�<�C���y���7����\��o�[[��;�@`�����e���G"'�yI� a��],";mH~NG��~�/d[,��G�UH�P��1p��Xy����a�41Ur��h�����4��3k�(vg�:;8�\�|�� 
�zCjc"�N����K�JB0�Ə��=6�jJsC��J�H�r�U�	.4���Q�w��ȱ��`�k�*,��Ch��b��ߋ�⬄�-�Ks]?�m���5ǆ�*~�rϠ�%1Y$?:E���e%������C�C4��s��oG�p`���`A2��$��kA�C8X-�m�s�%�x��n��ø�GJ~Y��vx9j���o�ǡ���rT��7>�i���S�Zy�Ί�RMf^ua%�͇I�Cȫ%?������@*/����u�r1o�ͦ�B���<$�J垜�� N�Gi��=�6(��*1P������v������E}�F��d�g ��\
�9e:�jځ���O
::���T���L8�.M�a�]y����</�!5����0��5P������>��
]bbB7��"d���E#tD�c���g4N�lX�48�K�Z�O�2l^�J���ˠ<�&�ES��񫒒�\�u�U��3���+��+�Ъ��p��bF�d3S,,�eYx9��P��8�\�`3��<�b���j�99�.�L��|Hœd.X:'ܪ1������Ǌ����w�3m9��AK�\����x%u�u��*� p�K7Ǩ��%�����U�K�^��]H�5�����]��.D���ԩzgɿD�[vnk�x��oE�nN�M���G�B2yi�Φ!��� ����ΛQ��v�
>�:�郶*Yu�������#�Z��Lh����r��-~Y��{�k���b �/�oS���Dbb�V6j��>�3��Ĩ�Em&&�
�c�p\��dw�-~�PQ�����()dӱ��6������������8������Laz�����8�BR4�_��3��ۢ �g��9�A2,����ͩ�<�y���Ճ��h,�]����m�߾�,���c��{f�A��&��AEPgk�#s�S�$e/�>�w\�������3�վb����*�M�H���ӠLȀ�e�Y�߼;$̈́��B�?Rg�4:w�r�1:�������#4 ���#���y�i.��fɭ�|#�6�K�v�1�4TtA���5W�g�+=����3��hI�7j�k��X�P[k����'{a%{�e��M�p�s�f����2���*�VI�����`YV�?�/m�
�����|�@���-���)�4Ό镀��f�7h	0		;����R�h�P���1���	p�T;ם��&����=�J�q�*R�F��x��jA�'�l(�zH4X734";�YS�0-�^����'+V�Qe�GU��˥���y��Y�Jk����=K*�@)�Y/%�u�C��S�:���'��h�>�1��&�=���� �us������B������M�3��)7�D:wr��ﵚͯ'��f4�c�9�T�tj��N#�ߞ CZǘ��Է�2��B>�*2�뫘�ܵ�x�y;	�~lP�栶w��� y��[�e��9	dDmWus6�-��.�߷�0�V��1�^���Ք��"����h���lk7Fj^m�-�� �����H�����K�7��	=�}yָDi���Ը���<V���A�qG����%��.p3����
c�tt�c^�ro�^�5�<
��6,�&�r��~�I5S�W�����k
�X�"����0���1��2��r��ך���)1��㩣{��J+��D�7��H`𽑩HZ��?	�� ��!��JZ�����i�O��E}r�׌P����Q�j�zh���2@f�T�g����^0n��}�`�g�j��F��*߸�S
/��)ۗ�d_��i,��a��H��&�G�����](�)8�*)�DQ:���,�n�,�q	����7tO)d}��5g�N����M��Z�F����ve���rWQL&!��=]�!o)b������.���F�?x	2�Y�bh(�HU����!��HEv~[�jf�Qu
E%�:h��pˊ��ef6mG�9.��E?��鬑��KKP	i`�����j=+����z�	�g-y#��h�J5�X�RTl^<��ܚ(� #3�.%|�d�6ի�e�d/�BG2���x:�U8k�B�� ���G���'��kV��.��
(��K����`[w��X�U$`WMJ
a���G���gӦ�ڎ��b����Url�L�t~����5�I�x�q�s��w�`�STj�~�|� �gN2��J��9-�d���v
O.�������+]@�fq�I��U)��׎��5a��>t���bD�����ׯX^[MX��X�Wg\턈a��-1��fA}�Է"���~��(.\�0	L�&!������I�:��o�^k�Kx)E��Cq7B!��.#�Ń@Ё��g9 ����1��ĐMO�X��!��S�!�&��:��R��6��go8C YV?cY��;f4���3��6����u�s;BR��E��HT�὿~�H�Da��sc�m٣ށ2ΜF�Dt�m���D�e�s��%��S�X�~��v�Rl��!e;S�t~�]�t*��V!�}��M�n�6khk0[�'��P7�D��yn�WpP�&.��G�#d���p�����İ����d����+��z�9t���c"J���ݳz���u��U�� ��uI��
��>E.�����i�=����W$�+voAP*�+�ro��zD.�Y��+�e<�*�:]����?�JIG��]�q��&�N�GB1��-݅^�sr�<Ge(���x��266���Z2��g���8�J^���c��g{G�1�#�x*�B�er�`�ǳ�EX]�I��h=tݭh-짒yђ�4��AK�4$J�u����e��)fdJ�!WZ$]��G4�_�7��T�8St4��&(�@�I^\t3N�{%�ש��o_Q{�{���L��	�����.����fÐ��X��/Ĩ��F�$1�7�>+A�e�R��C���� ��=i''�
0��~�� �u�S_?h+.o��n��������Q�����c*�6����BU�H�>�:�����k�̆Z2N��>k�Q0��C���L�^>vh��%�3�h�~��|�jVJ(`~s�ۚ0~R��Io�	����:�h��X�@d��/�0@�)dXͪ&�_�1�f6��-��F<K������iO�=I���f�F��_��
��V\>ڛ���+R^Ǫ*Bi�1]I��.�"[�@[mوR�6��y��O���+\ș�*Īl����u��9�+�̇�ѢN6�u�8���Zc����/hW�L2��.T����Xù ��d��Ѻ^NVN�uB�Mg*���w��ϋ'p��3o'���"u���H�r)��MnG_e�N�rgh�@��!�} �NX��%\�f���q�#,�xG��&6���&N�ߡ-�c�)��fR�;��{�ҹ�7�����882�캵B��B2s�Y:��@$��u�6����mrlѠ���Q�K��F��l�������3p��G%����,�b"ьmȳ'4?ؙ܏�۫�@f��N�#���ܐ��c�
vS�;�����a�^+��0��dQ�1|�;�5��Ǥm\��/B��U&�ToM&ணGVkc�ȴ�U�ڊ����u-���ڼ3�����QAD����#.��і�P������H�S�Sd����(]r���&�#|�p��g/�1ơ`yg�nw00N��x�`y�s-�W�d��{��[�D[$�u�1w�/h�[X��|~��Y~��A#)���O!	�����4?��`�ℑX�_8�� ?VU�Ur����A*�#֌�%՘�~su2���)_�q��n�'oSz��� jO%��@A����[C"�?a�t&�:|sqU��������1���F,;�bNx�S�ܩ�ȧĄ��q������"���8��Jﯝ{�|��(��랧5)O\��ǽ�:|7Lt�"���^W�8'�&*����,"��s��4"�