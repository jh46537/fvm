��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�y�Sy�;��>��&�MA�)Cʌtg���e�8~�����=H�9����.k������U��U�Xe���M�b�(	
'�m��_�S,(
>ɢ&T^5�[Kم~�WA��Mb�c#�<˃#:}��6͕��F��O�j�7���'AF�9��'�ƹrq�9�p�
o�'�w=��v��("�|��ӏ�I�\.�V�����)���cB�չ6�t3sꀚ u?�({��_x�W������!�`�e�H�H���|�-�YY�
ꆞ �Ӟ냨��e���S�kFd�v�e����y�*D���G�>����+�ᩜu�f�x�I���*��/1\1����r�2�*M_�4j�t�'{)ȳ:�A��!���ש��6�D`��Js�[�a�O[�G�O.�����}�9�����E���;I҄0"}̙�������@pi?%D;�4M�w)COD+�?�Q�ي��v���@�Yb����>��$��|�w�A}8���/���tv>��r{Q�ШRu!�Q�zL�;���H��?�"�@����Z���.�r��� q@^��Ea�\xҷBIT����l3b���R�0�3b_e��傪�5L<e7�aқ ����V���iԀ�I��7#?�l�,�SL��]9�g��|b�UB�yN`�T�c����Y(u2O���L��o���4�.�|����"ځ��	 ��h�1����ŧ�)�{�7��xw��6?x�� �<P���ܰG̛��E|�H���s�DT[mP_�� u��Ȱ����(�V��E�_�H7�
Gם'@���PU�����Փ��>�@��0۠��5��Jx�k��y��ieĂ:�o|�/q����2��k)�ڀ;��f?*w��Y�s9Mp�f��J@���xu��#]�n����YtO�`��1Tr��#I�D�>����M��-J�D��*�sW� :���R�V��w��
���u����+�L����v�Z�}?�����8	j��RSN��.���5�Lu�W�B�y�G��iK���B^s�X�XQ��I0���緇La��P��)C�6�ר��p���Mv��7Ȫ�!�p�$H~
2�7e{�A���K��;�����#�20�?�׆�~��G��\O���!l����	؉
.�3�|���<�B�0�)��dN0����"�ߟy�q\*].�W�E�:���s�C+7�d�����WY����Q'�2-�:nH��Wl�k��ƨG�fJ���;�HU��V�3�#�=�'K^��_�T��/E��(��_ ��ġ8P[��]-E
��͐�ʚ#7k�i�DDC^E��5v�s2o��W0e���`���s^�Ky��J�9/�OO������-��X��h��[�;ƚ4��5-[;��ͭ�  g6��[#�!�D��>���Ф@"����]��҂F�w~�Lt��;De�j�5�q4�}��f��<�8T�*ܥYm���O��[�)n��&K�FBw+N���nI�
�� ��-!tLtm�LFK�57��,�i0b�Ҕv��X!��y9�cç<s�[���Q�������F��`S�3՘"����x>�*ihbi+(�(���:�����&�Qú�Z����@�t���$b��䥥֎II�g�o��R���
{��2�A���7x��N�q�x�U��~	������z���;@lZ�쪽��ǙRFw'�'�y����N?�����\�@D�18��@4�̮T5����� ��P�r�ɖ,�,ͤǠ7�g����8~Xۨ�7� Q��N�5"؟�IӮ���l���j��uӿ������r��x1_�=� 2R�+(;C��lm�Y��'�ths��<O㇗mv�B�ղ{�\'Af:l���Z�25B�~Uk�����D�`��/ƍhʰ+�U����1����k���G��� 悅~���	�8O��ٶ�*�������G$#�̙�דN��k���Y�x���(/��d��eIR�1��s��� '�,��w� ��P���t��������ER�R.��;y|.�ˎL��?zYN6��$G|{�z"fh����=F�v�z�u�����uhB�f��V�}j�ҁ#X�#:��i3F���U��K"�jȎC(9&��k��Q[K<�������E�G-"�������u��`^��W�C�¨<-"Q4�S�p�AÑ=|p�E����3�b���D�)iF_��&��騡ĘK$h�94����)~��#5��p9
1���y��h��PL�r��-�sK۷�ӹ��ע���rh>� ������#�<:{t7['B���y��m��,3��K�I��,�g%����n�Z�. ʯC���jQ�cY��cs
�
7*!�_n����fmI��/�T3z w[2��'�4$�OR�"WF�c}��^cϽ�����'h��J�T�Bg(���
�	rHTg�?k^f�(����H4Vw+e�`�Y0�����8�^�7�0�\��7������:���S��2�=��/\��-�n�D�w�9Q��^��h�5�DP�T�?��)f_(���c�Z� ��2��_|F5����&e�&P[ޜ�Z���Z.N��� �V>�q$����"�����f����~j�"r��|�^Y$PNP��(���6�CTg������LD�-Χ�>ZX�>1H|��+\�Gn`�V�a��<�~g�O��z5H�������3Z����TZO���,ݭt;�V({, %p�]^?w=E��Sŋ���e5����}�gm�-���L`��L����Z�DN�����G�Ŵ/HW2*�w'�I��8�}lnf"���"�C�$y�G��V�9�'<���)	Ö@yc@���ڔ�j�c(��M�0�L[�F:�Y`����G9E_��[����֏i��b��'3\�f�PYx!F�����߽ew�� 7mz�ޫ�nʝ���w��/9ܠ���>}���>�%.�&0�|o�7��"SCt\���#}F���U��N�a��z����=f�?�)$�u�ރ;����~݋-�5:`�.}+� ��|ϭ���X��`��5wm�_%�"�_Ha�U�]�aL�R����B�b4��.��6�KB*tR�ט���8s�@x��а�CK�ߚ�j"�<��?*Q�$Nx�S:�W���
 V�z����Q���rkhñ(*|�/��qW-�Iط�z(��	g���m타����ڢS9[��GH�p���^�TZ�>�`�^Q�:���<|93�d��x��',Ö�')����n���0�-*�b� o�fZָh/7ݖ��+��_�OP�Ӗ�E�N��8{w��Pyg��j�͜@v�(j��`t��Ŕ�b�!��D�(~�~mS\�3�Xx���̐�*����1	A�3��i���Ĩ�Yߩ�|s�������ډ��a4	�E��5�P��E���ϓ;����� LBȡ9��д-OxZ�|
���we���۱��ٌ���Jd��3U�`9�³�]됉�lڣb���̢�Bf&��'FN����Ŕ��9<�ܑ
���y w��1�u@�;HݮnZ�+�09�Մ���q�n�v�ʐ
���7���#���a���1�ju�0��lny��	�h���e�{{�R�E�C��0�]rA�f�>����80��0����x�1�u���N��3�������b9�M(������CGz���F`���\6;�&{"�Fr�.J�q��<�e�1p����z���l��U9��(�k���3�?&��-|�Z��z(��� �,��ǅ��$3zB�Mc0�y��^�A���u��@��AD"�G��h�} �ⵉD�ۣv=��t\��fح�d��Ʋ�k����!MƉ��Ȫ\��md�Y���GP4͵�GH�����X�r��?���k��;��.PJ��\��9����̑*���&�g_R���BW��'�WO��������K�6C�)^�O���Obd�|�x#��_jF+n�x�O�7���_�B��䂑�����2�xN�B�|[�wF?��S7%�*�*�l�nΛu�Xrg?F��M�p6�+i��xO���r�@f� ����k$w�d��C
?��d%M�Jr U:�ԛ�n�C�_����=�5�R��`�g،}N<G�a�u�T����a[1�Q6�Ba?��]�����T|��[��mb������mV�t�C�1��*n�P���e�B�����0Q"��*ㄊ��S����@�?-�j}S>a@�!�ԯt��3�	ͮ��,`e��V��W�^|�W��PmVY��b�
��v�ھ�	��b֙ �o�2س��m�~Æ}��RS���d����㐨�OTA`f	�m��y�>����l]���Q��������Jk-V5���PNB��E<ND
��{]!���_���s�	�=[�'�=Y(��L������8�{����[&"��oc���2I��}E6�bk��[��Q�mRs��{��!OH�VXWj�T����K���0�Dl��%�[ߪ����l�ԧE`*��t<����<�2"~��;�ҷ�A�i{T�o���CHR�*f��L/v���fF���h�f�D�l��'c�}�6�m�s(�w���6̅+���ќ<�D�qb�.�!컇�ڴ� �T��,��?'}��&(�2��a����p݀�x�B�_�!�fF����'���DM�YR��14�B�����ۦ78� ��%�K�:������^Za�6�p�*����oSu_�%C�υ��� �IGٳ�e���6]���IH�a��|���ID�(����B��5��qI���caj� �hD�!�/�6xpJg�J8{�V�<�{�~�D�'��3��z���ZZ�4U��D���<%�2����"`i	)��قt(�c�N[><�Tt�%�ëDJ�1�N���5���ޯ��8�bAF�B���|��&U�M�U&��v���ֻo=y���^��*o/����;: (�;~x=6f6��LѸ`_�L1�35{���fs	A�l��t��sg/�Ti-�0=�@c���x����:��,����	0���	0�x�g�Ϡ��^1�I#��4��:���	���9oQڶմ�
H��,%�i�P��?"�@��A��V��݅�z�(��R�fկ�p@:8�>_��y6�[xyT�7ʨw4��o�.s�7SH��[9������iC8^�ײ��{=W8�~��3�d{�c��T�nt�8��GlFՔ��s/>���܍,�g��xdr`Z`��Sw%]��I��؃�)�ѹ~m�)��y
�߮�$.%��k0=�ݨ��:yh)ȷ�ax���2�[Mi����g��yF�NL��ZP(�����A��'��Ё�zQٱo_胮(��!�_����v("A��b�?�\��fB�@v �V\Bd�
��ç�oQ��1�'_X����]� ����Յ}y���:��V��z�ɿ�8��*�V�c��1}�r=5��9���k��U�T��m�:��q<�[ͼ-`��A;���'�PD�"�JF\�l�%�}iHY)<HpD�x��O���>9�S�w�~� �A��-yae�����}����臫�R�zYN�3��:�p�SN�l~�VAc>~�<��Gj6��_M�U!M��,\?�Ѷ��%��U�*�F�����]��M)眖��Od�W�@\�(,�v��d��X�X���&�\.U�� ��@'��{�M�-����xa�謱]�!������}��=Da��h2��,��b��g�گ=m9ݿ�k��G�T�LK�撜�N)��T��I��GR�ŌGr����5�R�rʓ�dS����b�p�;+��86���Xp�mHԌx_x-�Uh�����;�p��qF��������4�w��] _2�U���$�Fn���mG}���f_Ҝ@�E����cZ�%R��1h�0OJ���xKX|���ֶ����GW��*9�� �3����בß�����b;x�o&�k�WC C�\Ih�4�^ِ[�WG��΅�����u��p��z�חR�+��A#&m]8�6Z@��AF�D�z�Vhl��&�q�E�n�]c_��X��Iw+����X�̮�[:S,�:A8U�
usEYS��)(�k$������o콧��]=���RX���zؚ�ŋJ{�A;l��vB[ɞ���Ɩ!��5������Fʪ�r]����e��R�vF��Ì��j���љ�l�����(�a7�Y��`�>KA6����k��������r�D��}����O�D�&��ݨ";�9)�D�ΑC*����[�=�9�B��[�u��O�;t��ԿPuϻ.N��l����[�P���*[
�=K�cp� �~�?{��(����JY�Wt����jq�U.[^����m&��u{�	�U"PS >�``��2l��̺�Σ�<ydW/"-1HU�ġ�����@�{�r{"������ah�Q��7i+�������w��c`�\o+��Ҙ�����[���A����������%dT���B�'F�r݉�%�+/��beD'%���m�n$��� ��JK�8>?m�}V���{5�]Fʭ�v�6[S�A���f{�.k���,�>� <�2^��)��R�eq|�f�}��A�:J��늝�Ͱ�''�g�����t�+��T�xku5�[��fȱ��2�i�r~�/�6�X���LD�5%%�G���x�g	'$��nj��< e��Uɢ	B��V�>�����y-�����ɷ�Gɶ�g�a���pJ �P���{ˢ{��t�AGsǢ4jY@N	��Do���Γ�������n^�Љ��$̳���r�7�Q6�!���j>�q����I����<o��^������f��4���B��KD�M�C��0@D��%峞���S�Շ�X���~z$9t�)5���)���Z�Ҝr�����`��Z��TSw� ��yW�<�-�h�p�+���t��ĭ�N��}d�Q���W=�*����-4�U5k.����n�[�IKG��D���]���6^��zs��L�r���µz��,�	�Ym��@xJ�ʰ��lK�P�}�.�tB��d?�#���
,�W��˿e	�����x���%��^/f��Vd�-ta�l�8iL�g /�F�J.Y�u���a	ܦ-noRY�`�������I|�2}�L('_�9�ts�?
�=��(Kx��0H�+���?g��67�H3�ޓ�Skz��8��MU`h5!�2�:=�%��^��]9��_4FSSC��gu��	&�{Q��c=��HnI��U�l@��a���	�Oi�Qٵ�r�"�R��,g�JW��j�(�q3�s��1�Af9�`�¬�r�^a�G,Y�{���G>M��p\�`-�w%�ȋ���i���"6O��d�Х����*Gj���`fY�L.�<{+]�Z���.т4�Z�l���y��ֳ/H�T|�r}�׋{�v=\�Z��Y�� B�`����%�G�ew �Im�'xE��*�xt��2��2�����$�(���|Z:m8�t�%P��7�x�5�4uK��zm�߀��V��*@�k��2����-h��"P��j���ƭ^g=1�����G;�M��2� �6㲩�.����ͻ5���f�]�B��<�8EP�Y�\�ǃ��F��z�R-���;v�]�Z��{�3��Az�?�R���	w���Tfᆇd����i�@?����m��C�"��1�>�w�R����/�e��Q�i��$2����Ўq�\Ģ��K3�2@��3S���ɐ�=��������*i�x� ,����?*��`���)Y�Ē�j1;o�c�J�w�c�t��kI���7徿Ws ��fa!5�xݬ�_��\γ�è]���Ft%���
��ʛ��iʛ��
�ga�(�w�@X0b��0p�X���"~��?�dI�ں5n��ch
�EZ��S���{�A�{����c�C�c�W���&q<ĵ��x��Y\DB�����
�K�0�汭|3ʺ�v�o,�Ew}�.�UA����/k/`�\��`,�k� ����!���^t(����������".��驌)��!��mH�O@�ɭ�Á$sQ�����}����{�h��-�S�iU�v��	�l�>+XB�:	84����2�Q�\+\:��s�R�v
����u|31h�~��B����P�2���5K'zRL���ɿ��� 5�l�{}X6�󮦚�zl�9�nY1+�苖r::���?����(b��I�@�o�$��IϮ֌/!?=ߠ{�kKu�G;��x�B��w����W@��T �1?H=�@J�&�l���FLO�}�����e�����yy̌�.�){�#���{T�-��>�㡾5�'�Z�y��P�u� OR3��DT	��������y0{;�k�R���,������U5��B�x5�5&��%���?�9�$�<�[���o���%�X�5~5_?��H%Q���(ʹ�Ə��=�lڥi�2V2�,,xf;���V	�����=Z;eSK�a�7����+닝R��m�/����f�'��R�Z� ��z.i;62,�"g�h����Vi�ھx��ֈ��R ���d�T@�\�T96�p������e�8]_EQ`k�@ѵh�+���}U�:
	v�l4���#�`1/"]�hT���{'�~({B��R�9��By��	�y�<Wq[�g`_���vD$��A�'·_f�g�n,	̕-��4f����h�7�t�5��haa͗�]y66����|����p�hZ`��1T��ӱ���jd,j�7���x�O��An��ds8$3���4���15K��XΊ��y�i�r¾C)Y�t�c/�y�$�����b���̬WJT� ա��*�{�D�B\m����.�LPj�%�X&���	���luw��%�ѷ\q�ko�n}�lc��o��f0.N&��g4���tyW�^�{���Zg�ԣ��&�ג�И�0��aIBY�w�t���3-OXޓ�uV�S~Z�0V�3��A����|�o���4䄴�����ٴB��hE���H��k����]���>'4;��E<^�z�g���Q�l�M%���+-�S�}���ל��g�(�̶>�|��U��S�_��Ō��<�\�|�v?s	��c�4���7�H�������΢�I�m
�#T'=�{ .���b���>hv>����?����2M����Q���h��i��m�`��o<H�Ok����@)Q�n��5}�`��\�j�ik���>&5OU�����39x�0�t��7up̠8���O���Q~�&��>���Z�_,)�˨x�/w�E�a�w�ig��[���9{،[T�v�7Qy�v�-���sZ���D��6A���%Za��S�w�����M�g31���f�,��ng�.�VkA����t�k.���.f��[W���%����4�v�ZJ��&���u~%�jD?5��Rq�ܭ;j%�$E�yX�"r�a�'��D�%�?��?U�~&$`
@�΅756��n?���K�������W�;�M� ț�BEv<��:�\�W��Em��sr��E6Kx���b�c���-q1uOB�3NQ�Ȥ�O��>@��'>&�-�jNY���,$��3?�EY����wT�#zz��mk0o��BO��S]��^MK�okS�a*��G9R!�D�d&a�9��l# >s+���Lq�ϴ�F��{Y<���+\}�?Y	.s�\9��.��o�u�gK�P<�V�͟m�ؐ���*ڦ�P+�I����DÚ�ل+���1��@��	��
���rC���]���5����9���웤�ĵ�#�,����#�.?�}��S�j�,u�y��`�Tb/	�巯�J�i)��N���Rdp0���� ���d�z�b�G�]�e���Ա���X�����\k���[���2vM�c C�Z�W	2�i<\ͭ��~����:1�N!N1��̌�`�|$WoC_�� 0�����%%�T�{��#S�Q��oP�9��lAހ%�6>�'�rV��K�NGTٺ&#jD.�k�7��˕�j�l<NI@*���ځ*~p�����`�