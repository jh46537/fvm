��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb&�L�S��O�2�0�M9-H��*�����"'�ӛG�n��pR/�|PŇ��\�A�6j��N5�V�V�@�[:7B�޾�r��]:�.�����j�Y�(���u�Wd$���8�AƇc($�t��-xg4M��u]b>x@]6����_�y�h����E���"�ޡ���*ﮝ��w�O\���4ꂲݒǞ����*��]ah���; 3�*^3o͵��WZ�F��Q;Ǐxm]����A����b�T���O L��ݥ��Q]*V�o��yZLF9�Ưzd�V�J��?�����8��1;�-���� t����}"}ǡ9g��m��ymJ�_r�'��S�E��L���м�	����,�*���(~���(�B�I���V�H5Zx�Y�]I�L��B���X?V��̓�S����$��ӣL��0�d���+C�Eᴲy��>OMΟRÎY+/�jjc�	��M�6m���ޔ9�LB�X��섏إR�
�aM�)�{��_�t�J2�� ���8���6��SL; �F����Dl�]j+��u)�a������]����z���;�AI�Rh�����z}��a��Tf6��\pW�g�b�����?"���4EyN:D��eJ�n�)t��t�d��E;T��mxGԲ`jo�}�?bq�Xx}w�����n��^��@�z����V� ���)�&c���R.Q�>�&�>���41s�f��	�,��ͪ ���$^�1XVQ��I�%� �Vx+����
�XU�P)�Kr�IgT�#�SS�̴�	x���0�l0�E��5�e�&.G�V�z��]��g����k@?<��������M[��h���4��JlR��Dh&�]~2���ɴŢ~~܎^����'�O�s���f�N%�Gv�Pɾ+6!E_����s	`{ocQ��$_��Z1��F
���	��>ߓ+��U��z�\��Aq��Pm}��&k�W�~r$��o/�?�wB>��M�$�t��rcOo��G�{���h���?�����w��sz��El�aT�[�Plh���!��V6�zG��q�T*�]A���S ���9�X�yhКˎq�*Z�y�5@ ��k~6���I�r�_�!�Jp�ۓuףskЅV�7-2ݴ9y(��nƨ�o�}��1*��-�9�f�z�0W��WV� z5�!��"�<�AlX&T	����{� '�(�-Z{]��"Lj�]��tnT��i{&�S�Q3���tj�N�},���d��/m��u� ��uPU2y�C7��.��o�rZՓ�/�%�����'ŌM/�S���1���(���Oʨ��p
PwQ�~�.ĳ��+N�cS��'���X��K�7��[t'd�7h ćI�K��O �u��,��:���)�~�����k,�cA��@J/�]GߓB\8����rS�O�>И�$d�ܕ�6>��T-���� �:1����'#/��Ӎ,��؂�ɊmX*���ĳA�5�͔��?й�G$`�� ������'&�8T<j"�����(?s�8���CA4�j���ь�ۿ��h9'{�ϲ�"!��S��h���q�����|��'Δ�܈�� �r>�":!��l
F��!c��D��g�Fh
���������Z{�;=��X�C�M$B�/%���[���,�m3"�f��#���kfχL��.u]�������ak�{R
r�AE~�X��7[zd�y,?����H(xKDg�U���E�J^Ġ8�JF"�9[�R;��p�|!�������z���\�j���N_�~9�q����[|z�?��F+i>��r[:�]o[�
��{�f ��Y��}�4>�W0��\�`�f�qܯ���Ö�204?v�|�7�2qq��i��@|�ւU'��a�-��<��SN���LL,g�9�-,ZPr"A�����ї~<,��ެ/S!����e���X�S�T���7��^�
�1�2T2c���qZ����5,6�����
�AP.]�^�_�l�K��[�ԙV��m��^f�cb�B��*y�؏�
�e�w��u1�O�)�B��t�4��2��5��'�)�dբT_��(T
VY�T���-�rh���>v�;Y��4����q2���Wa�Y��1dW08��H����TrA��h��%E~E}�u���V�1������J�\0Ct�J��uC��v�_���j?��Ꚓ^��~</d����)K�,}��
�O����g%���&��-�W�{�	wf�U{`.}|.���C��t � ��İ�H��/� ���O�D�XR9��U���P�	 ��>�{0���_���6�k�k��R1v
prGo2�SW����C�GMb������*�'<8�6�o/��c�vA�E����m�V������ݠr�a�}�|�`�<!|�b�w숂srP�����X�-Gus�p��lC�T���!�X����� R'32ƪ�V�ؗyvhǌ��)x��_v!��dl��G��c@n���=��/�[ӻ��L��-�ҼgƂ�#���0d�ȋ�)$�c�5���l��*L� G?d/Ƕ�����AMZ�*�Y�NeH墳'B �y��M���-_ ��~�������h��QJ�-2~ZݺL3p�Im�C� �)b�w��#��9>�M����!��8{UI2K���V�l�Dp�����j�F�K�o��t��|ٜ|��O\�b��#?%c�&�%�uԃ�ͳJ��Qc�ؠ���y��ݡr.�C��e�ښ6�"�[o\�2����f>ԋ��=�f�����}۪S��(A>��P"ub;o�6�& dU��i��}���%��Oq�9)4�V��2���l�|ֱ�1 ��N`�S����V�n�8��\��sJ��#�^?�W���^�*9]yR�IdJ'�p�M���3܂_�,E���)��2Ak��w~���}�-cV�$*�����4M�}��<~�n�2���2�Ӻ��80|�=�C�_��Ou�rj�GEc{!#I]�N�mjJ�4���Hl#�A�\�Ad�#yadx�����Gk��/�dV@��>!�H<�x���	�ll�NHԬ=�TL���o\D�^��bc}U�`��ft졉/tR[ܻ�2V�5�u&O���9XV�[6W�b'�5�\r��	x�ӭ�!�T��d��-�IvJ���p��`��6���NՆ"�<V���ddHH�i�[$S4YXR�E*������4�zn��Ŀ��9 ����>vb���t�@����3ѸJ�o���
Zl�r��m�1�g�����~k�9�/A���8d�(��W�;�3�����Q/�G�y�s�>�4.��H��Й�dD�-*�q��-�J'�K'Pd�y��M�8j�h�y���j�r�N�)t+%xi��~�u R5��9B��1c�7�}׺	�yi�c��rI& �rj�S�{��[�Ī g���YU&�H� 9�Nl�4Y�^��!RP��$Y��b��x��a�@��̞�*�	���H�e���p�|�1��T�@�Ùc��9��ʸ��M��o�K����%Ȭ�K5�c���
�񥖈����S�,�i��:I�F�<���0�}���}N�k�Ă��Ĕͳy�E���s��IԪ|�������ڈ?�T�tm���8o��7���B���a���6y-�dݓ�Ј��U�q�_�O�.��H��\L���EQ�������I�?�{1����ѿ�f��E��6f����5�=�%���;��s(�b;Y�ʎ�`�bїX]���hP�w�׮��_��
�o�V~����Ȩ6��$�x�)(w�;� �T\l�G�뫞'��ԳP���I��c���@ē+0�?�̄0�HL�Pi�?��x_�[疯�i<
�:x?�*N'|_ZI2���xAZ(�llBb���Nk�h���Ϗ��tRyz˪��v�<��C���#�{8�d�Q�K��C�Y���5�;T��O��B�R���3ɦ��.J̳�X]6@�/S�:���/���u�zO���M�֍�����K$��E����N�$ƥ'� �@��9p��.�<��!-�qo���f����ٟ��w�KˋM	���Q�f�m���,�@�i��9�Q�.Yz�Tj�{�z<���d24	0���M����MޑK����ܟH����O-��x�r�^,��L��Y����t�r>]�f�H8�TC?^�����X��/��r���td@#~_�rA^3�l��ƘZW7'hy}R�@Q��/ũ0u������l������R��Y�U�0�|�%�$	_�g��B��B�g�T޵�Qw����ؔ���c�ֺ5�H�� t�����TB�㏉Is�(\��b' �?�f}��Q|$�aK�@��\(�m��
���{z?Q�Y���Ǚ�N�ĚU�l��4X�uUX��s�&NXs�_��\�y5?7��"UO[��ko�RV�D/X��J�v;
�3j3��/m���Zs��כ�%7ጞ�Q�W���]�cZ�H�c�W�:��:NE���������eAT���;��
9A^��6�m��0��tC�-�����Պi(�o�a��	�قؔ]�����v�V��h���E��	|�c~=O6�x�3�xG�d�y{�&r���<B�X��`�lE����v�$[q)��[BKz�o|4���or�xu���A��)����4G~B���j�8!��������Ҳ�j�B�+�!W�����A��WF�|<��ٴ�.����*P1�2����K�q�w���"O�P�������l�M_���� �)di?t�U|���}��ks��^�K�$�55����	t��;n^��G�.��Q��O*'h���`�m�j'O)}�����{�M�T�!Li�N�Oa���]��3�ԁݚ���Ze%t4�c� ���s��j���8|+�00)�)��RW�}"��Yִ��*p����@!�k�?<tv�z�mk���.��Ƃ���� �֒x�Ӄ�@ �S�Tk�[�/Ӎ���Ldb��kfsse�}H��h���D���C�T/Dgu�������M(����F��O ���Un���`'p=�����(�^e.i�3��SQ6Zڟ��~J~��jPt�+F��W�d��dN'[�$6�(����ǎ�^0#S7��2h�j
Y�Z�JH.�産�+5��ׄ�l:��d`e�S�ʠ۩�$���6���/��/ȕ��*K�[n�J�'�pC��МJeqw�̯�-D�2�Vx"U��vf�%����a-f̍��i^���B���"��c^��� �<��H͜V�����d@`�kȅ�!d��������H���W5��z� �l^
ki�a���:D�h
��e�s�!�����.�`S��$Y4�;*���Q���@�J���3�
�����"x���Rk_"�5�%B�^Ͳ�ǎ�#��lOռ���pR�jXvJ�l+�*j.M�xe/�яpVh��۵
TV]T���
����!�j߆�ܨ��A�4'6Zuoߤz4r=ER)$������µa��ײ�����fqt�����~O�-�_�sp����O6�]n��H�A�}���VE6����l��N��g�@٤$D2��B��k�d^]������x{#�R��}�f/��]����,�HA����P�񐷻o���Q�:��}O��=>!ҳ��C�!W�2G�_�ZT����B��.z�݇k����@���2��M���#~}?�_|���v�v��ߕ�$?�z�Pl��Z�y	����Eu����HWp��iS�lz�y #D	=�����wp�P���]����̢,K�+4IZ�Z~c@B5�c!	s���{�=��\Z�T�M��'�Y��8H?���.wJ��v�ҕ��l,�r���E<"�qY���Xy��w<����P�fVj8������-ߢ��l��aJD1n�z���(�1��K�"��9��?@���B�a̰��\F��W"����*GO	��^�ˠ�QvaT|����n;���%~@Hõrj�Y/�~7��
���B���/��i����VҒ4��4�B� ��(z耊f@�6������QP%��$���y,��DD9�`E."y*��j�{O��&|q	TV�ߎ	Y-��lA	�l(B��"��վKr��t�� @��)#��d.�g�Z����8G����p���_�8Z��p��~��i�7U�ѮKV�񳳮�\��U�þa���m/����bP�I��]�d�f��d=�q��wV�%W� �Gi�� ���q�[0�U�L%EuedͧL����*��c�]j�����5�F�F}A�.�dq�R9��1�Dr).����m�oJv������9[��Z � 8U+0E՞���4v�����8�Y��=����ӓz1P.���e2����k8�ǀ�0�	�0V.�(�����Z��*�'�k�z��(<�?�)��� U��g9��6��E����z�Wc��t��>�����vIz9, ⸻x<���ƭ����O�g%¢sڃ�Ȩ�1��Đ<�)o/�(�6H7 K�����i�GqZ[5���t�!\5��-Z}G�R��KT8��(n��3C}P��g
��
�\H$��pX�k!�O5��Ps������:��)�M�Q��6��Ĺ�RE:��2m�V��R´	���T].�9�imQf
�V�j�Cj�iV���Uj�1Rܨa�{퀾�h�I��탦T��FY�E���Щ��TG#�Z���D�^hH����m�%|� ��<��a� �����9)߷�G�-�=2��G�-Xye���� L�B�?AA��Y���Z6x�E��B�@�N4�}�V4�~�Zݙ����*Dq��]D;�=*�p���!��� ��(�q��2�B��A�~!�5��^X4tj$
��#j��F�pU����/ �:���#��_HU�bW�|��*�xˠ�z��d)ms	(����=U�r�[Ã�s�7�n"[�T&��i����Kc`�T�4���WL��γٶ��Ҋ,�4 \�\ǐuFO��A���P��fYs�Jq���p�����4¥E$L�q�	���x���Yg �9�2�S�/\J(�Z��.:�a��~g��,�x����b7p���;:�|_���l8 u�_HNSr��Hq�C�}�q, �O�j����i#�݋'0�~�j�)��
݁)Ym�5"�&]b�*������=i�������c�m����gG/ױ^�#S��h+.,9��S�\/(�}�쑐ҸE{*��$���rBN�닯�+r
���ł9Kf�
��e4gh�I�BN�j���_~��y�Q��2A�'�O5���;�����:�k+��cM�"��<���hP���wT/��"�ԓ�q���#$�X�c_TY��K������vS;>|��0/��J�+g�q�E�*�%U�v�ރ��G�n�Y���x�q��Ky3#�,����-�J�ģC�����)������8� ɵ.�}����C��!7��er��Ԩ3|����-�g��[L��I�4F��0�p �\������F�j �c.c�2؊���ܿ��B�Vy�$��T{ZD�Ş��=�l[.�w�᱙�+�����xua�Δ\P��uJ~�� ^�$~�'�Ta��6�m��u��>s�~��}k�0fݗ[��V����22�۳ ����)�y_�;������J�	`�i�y�D���;�f�G��t�ϔP�J�XKvI鎵P���E���R�c�k�X@�H�w��� ��Wr�7 �z�l,�K9����rK��,Z\�~���B��p�*��ˌ�5F���0T�l^�pT��|\ˣ��b�)W#5����l%n>K��g�dKBS�'2�����|+�}K�?��(��4<����K��w��/�o���Y0�+oY��n6YS؃�"4�XFT1L2�D�f��!o�V�&�xoB]�V#�N�3:�UAZ!T�)����p��J<�S�c����J��=��౗��e+:5m����e-�W\���9*�~e��d��W�aޣ�a�/�`&&�ƺ��-:r�|A�j�����'���'Χ�Գ���ki��zz��ۋgi�#��F��trY�1��N���~s�����:��J%�chb��N��5Q�"�Q���V�T�ØɈGeyb%-�%0�(�(���+�_�����x�k�ە<�p�%2�V�U��*l��M�.�,�!��j�?QQ��1�$�����qv��<��y���M�FS`����d��d���>
�B-�/�g�\@�yE�K�KE-r
�|�R�=�2_��p>s,�'d�Z�"��������^{��31��T~9�[�>H�F>	����"��D�+�6��_g�ݕBV����u���PaH���3$��=Ԫ�6c��>S�	):: ���}���y�W���B`u�iь����m-)jN�M��xةj���ҥ�i%�R�D�1���a���	W����	µdW��須����v=��b��r`��u��.�^��Ѿ���vgd��
����|�f�o+��i${n"��[M�����4_T��v�a�"8�>]l]�j<��-t{~�˺�~E�O�
�EA݌ԭ���G25��Aے"8�>F�c��b�?����g��$֚�����O��L��Bʇ\�h��7�k�$O$�)�v��"����:x}wڦ���C�7Ӄ$��U���QVp�`�R!F�g=�z��t���G�F듪�t�+~��<��a��(f챉��(��ag�/��K�~(\�eϤ��8ʫ�f2�|�%6o�׷2���!͉���P���c�D��c����}��3���Է��r�³� ���˼4 �z'l9���E�n�����k�����z[�_�*%�﯅��a:I{�5듫{��*�[�!�����jf�2Q�G�?ba/.�����k��a���s�m�=V�l]�0m"�!�m3�\��Խ����
_����S�8X
|��ph&�PY�]n]_j��
"��w�$�Wf$^Kx�j¥��X[�8ޒ���ub�%N���,
	z�!�D9I�����{_z��󧣮�	�� ��prVx�{O�����l+����U븮X�	��g:����9s�%��73���QZ��c����2Ve`�a#8Z)��V��=$?&�kv��#d�Tp
��׽��ۉ�l�2��u<�?�#�V��+���ŏO�_O�G:��K1J0�ˏի������+��E�Z�?�őVJrC�pz�Q�4�ӫ	�^�P4k���Z`ՏX�j �7ta��NjcQy����H��j�ZNyl��������&?�?�%0���X���ZJHqJgη�T�j�Lĭ�+�_�g9���	����R��(x:ЊM�6��$&Y�*�D�z9����,oʕ����
G��5QdX�u@����?�T��R%\��xĜë�@LF�Z��E=K�ٺ�R��k?m�w�b��ޑ����-_j:ہ�F�:��J�"�	{����;q۰\���59�v��E�R���E�����t%#ǃ��
��}5��9��n�H�7�yKa�!|/3��d"�s�Z�f5� �X�0�aC���3�R�1��� G����F3=�!�����q�E���[��'~fGl�v�hs��m~�/��Ƃ����D/_'ō�˒o�+�Un��J�/�g�<���dV�EB�<�q���af�e��j�9@I ܁P������pSJ�i� �v���O��u�}�(�D�Q��x�Q5�6X�ڎ7�E��mI�Y)ȑ-h�e@�������Q��B���������Z\/ϓ9T;���;�i�W�?4�1/���f����~�5V��.@ $��T�ϛk �"�{���bW��z/ �\e־R�`��Iw��~%ė~Ƞ_59�ʫ��n{s� ���Q������ �J��Y�`���*ΞR�ڑ�yڇ���*��^s�Z��̩��l��Qs\4g��WYf�W��9家/@�+�*��N���"O�p���ȕ�j�9��H���c��|� �9�-�������p���1�@Xt�%9}�?�Ug��x�2^q�(�^�4�`fm�'����L�%�g����\z�0�$�����@����D$$�� HEqr��Q}q����>�H�MߵܐS�c>/��x���9�j�3�I���eF4�#�(��;�+�l�{�ϟ��i/�(��&�4���� T�H�:�>��w�'>.� [�hp`%%	�����1v&lh�Q�̵���� 0�aX��69�6	�E[Z�����Di��x����奉]��f~'}��*֚�&������i��C�yJ��X��y[���.������PeD�p�w/hx�4�4bo6�ck$�Q�D��=|�Uʎ��w;#�*M={g/�!50F��^����/�R6Ǯ+�1J��pAC����W�h�Ǜ��1�e�y�~1eòt��k�H14���z!�@T�i�ؽ�	���!���ϦB>��'�ew� '�����ȼ]gJW��+�z�-��|'H��U�L^t.���������X�"=�}Y�5j�uGI�e1@ ���b�P��0n�u.t�7��A���1��w�DA������Ό�D��)2j&��@�2u�?(�RI���+�4��x�vd��|F��<����.�,CD_���[v��w	~�S�����*�0���5�l}��M��ӳ�)o���Ů{`q�Ȑ��ܒǜ�r�y��D�`I�y��;G�{c+���^f���â�t�W�5Omw���6���K����M��X��7����Pn_M	�U#V*�D(�� y�h�f@����ϮZ�6�a�x>��ih���T�.j��馑=g,~D� ��U�O��\�6k���t�W�*z{ ��'>�=s8�.��п��Q!uTpq��T��9�p{�{ʃƉ9S�-�	���u��;�=u�h��U�8�ID�� W��������,�F��C��2Ibk����$�͍�>�2�J3�S��ef�������ʠ�N�ˇ�j�s�_T���l-���:XZ�1�Pi�&"ĥ<��@��W�U�/"t��ҁ⑁�C/�/���f݃*�F��}��K�Geș�L#@�H�1Gg�O��+����D�"v�k��Ү3uy�L�v��6�8�W���^���]�l'��ؐA������2�YQװCɺ��d�O#m��\����������ϰ�<ӄӰ'5��oS[�9j�`�����'Y(��gdC|c�Y��IiU�5�ݜ�s�=�E�1�fW�*t�eiqN��`=�L�e-�Ҍn�Bnk�#�HL�2IJn��^27��a��G�F���h��s�9�`vs����S�@ݸ?��
�Urd��� �.�c�Ԡ�i�/��*w:�g#��n�GwCLR0)^l�7zn�|��[��g���k(�?%ŖEE��>��-�\UVX�&�P��S�63o&-W��&k,������0�_T�µ���>6�Ou�S3<Je�3�@��Ɋ��䪕�ɒ�p��7|�pL�2pf�P�e���I�?��a���N�9��I^�I�i��&�u���p�'e�Gv~�V��1�������qK�:�����/T?;v��/9p]�0�K�}8mk8h|��e�m��B1��I$�I�X6&������>���Z.��m�N����89�v{b7*.�z퀱��|?��W?~�����2G�����Q��\yߍ<Bx������<��E#���v�K>�`\�8�13C=�.��U'ٟ�1��çqecTJ'���hcG��Ǭ�M.��үNay��7ބ�KT?�%7��E��Jz��QY�g�'���ؙѦ-y���e8C��G�<��)�үc���ڹ[+�Y� �-g���Eg�Æ	�CN���W��Zpx�X�0ļ�L����j�Cѣ��D�)7
P){����g>UpW^/��yȩ!U����E��e;�����Of Z ��5]W��%-��ns�;!�(���h������(����-�ۡ#Tf���}�x�} ��0�5��Nxm#*�ޥT(�Z\sl�H-�X$w&����n��|��h�bW�~���_���vM�kk#��0��X�eKD*|�?a�@@�O�y�yt����+���~`�^�]��B4f��b8�|�6��br ���>���������Y�/���r!����i��r�گ�	��E�:%��>/��q���6���^T��i�N�Pb8�Q��9�a��5\n�Q��Dxo�(ӣ ��;�H{=�s����'�Y�(���rǲ!Ę
���G4�����<����W�~�'hb��{�e�����0�ɖ9���Zn����~(XsK�|�.M���`S�	E�	��ڤ7��䚷�0޾��:
 �|�R�F���q�~��&���`zs�Y�T�^��-�	����C��$��){JC	��m�{v+����ti�Jtr��rb8!����������<~��ϼ�	�K�����^����n��v����	�����U;*�09�)l}�9��4�� ��W@	�|;UH��2��;��Δ����6W�8�+ْQ}���Q4^dy�z�����Y ��V:k���]G[����x٧ާ��C��	�	<��VX,}76�&\C	f�l�tQ?�c���O����V��n}1Ȳ���qB�0�vLV��@9T�}���I,��u|�b3%zv:�:�p`J�e�E�v\N�����w5�`��>'�)��:6s�Aō��x�{�Ʊ|(dF8�R�7�#�1$j�"k�K�z)�Z��s2	��9�H���KƝ9�f~G�$���xR,�*Q>�]�`ĥ�D�iF��@�W����,�|2�U'D���������P:`A.���Z�s�w&]�ܙͯ��I��gl��H`(X�=��q�$���?BO�8Z=M�{��
�J��{�Fm;����	T�D�y���	���ׁ"�(L�9��	6d7z����<VںM�Ǡf���TuU� ����"&��_f�7#�r��.�\���7�;�/@﯇��"?ޅ�hQ/S������"�x��\�����S��\^���܍�B�9Ba����ǔR��+�磀аl_�/%�rV��	X;[_�7<i�F�aM�2����\L{�Z���+SV|����d�Yd�"<�u����cF��hb�~,y"đ\�S�_KI�D&�^c�Ab����kX����R��!>t��ruT�Q���U*����h�l���/� �7L��w϶���yr�EDʧ����sy�#�:W*��髅X4*"�E@z�R�z�ʃ�nrJ�]ǘ=�,MF7���/]�P���fQ
V��b���,�٬cs�yQ�!+�����{.�mi���S� �y<ʻ�=��Ri1��L^�0��`����ޥ��gJG�"����t3�LzjiM�h�d�F��$�'�[�F�m�C���sr� <ۗZ�u����6����
qց�R�YH�ʺk�5���C����%S���-e _NHDd����E�i/��E�Z�<��2=�����>��Č����E/?���	B�9P�iH ���HsOI���Q��D�� (^��O�J)��&�X���Ra�G����	�\mX���}4�!s��`i���s�;���������q�Y8sya�M����[J���������}D�+�mN��n5�y�G���ɜ�Vh�)~�2@^�ӆ�猏W�A����bIH��>�C~B��d���&��]���8���]+s�A�۠v��F�R����z'B�w,��`jT'
|��&��y��jxm]"��|�"�q/��`�h�ǜ�.B[S͹;�I���G��<���z)$��Q�/A#�;(2��|�ˑ�{]�^���L��Dڸ�4�:h��Q�w���0{o��#^#}��m��>�m����!v�#
�����������`�6��Jr��/QY��Z�٧}�HQ��Ӑs�?1 �q5���=��xg�W�Y8�I٠U�J�="�N�>t׃���k�b�Z�T�&�G.]f��Ba}���<����� ��&Ba��Qܼ��~��Dvoϛ����	��;����� |EA�I���'P�����B�{�c�-��x�7$��M��Ll#	�ؙ /"A�԰WG���c����L���Ŭ<u���H��A��<�n6r*�Rp?�kUQ�]�Ά�rqn��sM��B���iq��"�I����j��<�p�s�c{��xȅ|N�)Ō���0$�qVS�%����2ԟč!#ƫ�ζ��~`�|�\�)��F;�=���1��F��>���a�㢱�2�@�<�a���U� <#����IJ��8�cS�LX��"�V� @����}�u����4I�����D�aLcv�֜R�U/��T'��Z��,��߂9\�S�V0�jҰXKN$���:.~v�^�*T���3�L��k���B�B����N�w��h�)BX��,Է1���]��E��S�W����j��ڝ>�wv	Ռ�����~���GK��L�nj��*ȏ� ��˦M��@��Oӈ������=��M���?�YzLC�9c���TG�5���V��]6�~ʠ�p�y�&ᗀ�-��S���Y�m�O�(��=�'�u���634�9�l�֣M��`�aR�t��R(��
� �����"'�p�i�g�9R��B�Gz��.�jc���~^ة�1�yU�ҥ�¦
z=��O�$./���禆��qC�Gob��:�~�V��&�2NxD����Y��vF��VD�JH���=4�a��e�.����'eZ��	�*�Ҏ� �|/�XaTu�,��ܤ�S�p��t����٨������m�I��O�����>��<����\J��;���Q㢬]5^#%��O�KRu)�k��a 4�e6Ϯ5��=��x_Q'��<� s�p�G觏-���(��8S�*?	�&�P#2h�(r��u��vm3�^qDB��s}�8,4�a��������ܫw�ErC�o_��J;�z;�.��z?1PO��6�m��E�X���<G��N��*�"�(T��L܎�i��O�C;>�YO ������Mܴ���5㭴��xK����	�4,���,̿�ݛۇ���i�$[Ϫ�#�֝l��۸	�d�ϑ�"m2�&%"iYB��7J/�q��`��צ�8��Q��L�(����u��	>0�T!��R��m���*�E�BF�ٝ콎$F:�FW�d��t+a9��Č��_m���,���M������e��B� ���F��[�{�fEm) 9x��~&�D�U�8H���bz@Ŧr�c�c6����y�-�  �2a�Ξ�#�������7s`Q �"� ���&J�4{�NyNP�)F���@���A��ֱW��e�2(x�c�:%�EIh�������L���#��򌌲���N�Q:��R� ���\|�Z����-����,:�$@���D��<Ɛ��.��6��@�cn�'�R<��ǻݨ&N1nq�ÈWZg@��/5σ���2�	���q���S���I���j	6�i�g�x�O�g��<�?՛7���Q�e���2���_���3 ��H3����VI`)����I�k���D>�N�¢w�ăx��tN�h� �<���Gj(P��;��f�9��H�p��`*-k��Ĥ`���5��ê	�\mER�ؗk�R�b�@YI��"/D��W��ˆ���[��|��Mw7;^m��g�7��Q�-
d��p(V���c<+�v~�:
�K�l�&"������V$�.��j\��T�G�x .���zW.FO���{ �$�"ҁ�C�S�{r{�6,�6���xC��/����� ��}���؜�[���Hm4�E�^�+��8?��xJ���:ko�d��� ��\�Am�C҄5��h�Ү��i��3�[;�E	kB��w���.۳a�-�{���Yv�m�'њ-�YK�_uO�I|@κұ��W�>�K^9��V�HW���bËV��ꉬ�K��e���R�(r�=��mdJ��X�T��ȅ �ݼ��?~H
m�VxF���
V�H J�Yx�h�CWm�A�W�Rً$H�߲��fT~��*R}�v�f����|u9��r�A��x�n%�J��	�j: �uuo��)E��ت����k�%Ҋ��̹�8��qi�
q^
�[��w���ʩ��#g�Ϗh<H�2\�6�A^��}jD��Gv�^�B�p��4Q����
�\�#��̝~��R�,y=�uN�C�'>��n�w~*Fޅ���]��� ��t����_��%6p��z�[�|���0ɾ괢ˢ���]��ݶ&��B�&��'���%Qu�P�s�Kly�W��,�p�_�Z�J�|c_W�|���)~�$�k��0|�?�m���'|`�I��@6��1��ފ
[�����C���EG���N��>㐤��d���ҽ�3=×�P9i '�LU��
 �x����ߘ�_yZŦ�(�������@"���� ɝ�v!ޤ��b�俳K���_�8��J�3ǡ�΁Q+K �R�`4��C��;��I,�8Bp��W�:�3���&�i_m ���2M
Qq�t�rOI�O����2�*L�A|b�PvU�c������)�nݕ-q�48���Oˬ�\�_��56��J+. �<E�6���y�r	r�U�d<����?�KV��ժ�(k�>yp�C)���B��8�#?n��@��y���[IRls���z+
<�C�� ~_��N�,>��_�����_���w-,�])7|�:���m�-���Fo��DN�)"�9z��:�s%���S��Y��Nt�6�2DlDXgʬs¹]��m���Z��ewqf*�I���_���Z�>��G����{ꌹY$�wo�ڛ~��o?��aeͱ��ܿ漘"��C������'��[~'�@�J�С��<:|rC����ܗJ|�Q]���{E�|����g���^[F��gP��=���$�}�J�����~���1��5��Kl �:���������С��=�MS��7PM 3z�=Ô��#��r�,���㟬����g)���D�#�%}�%�S9���>�At��'�ǽ*(މ���.ђg����y�V]!%Y �o�A1�?�ʯ�s_�*�"&��P��zC�-��PP̗s��U@x�l�:_*�ne̔�������C9����L_)Lآ5<�{��n��l�+R�ٔ��eK���L��P<"2sa���n�D&A�W?���t�"2Ӓ h��^=>�C^�W�O��^�%��*q�s]I�PE%�9.��dӠ
�8�ɠ��z���x��Q�"�^��&ݧ����vsI�����v�X2�L1��W8Q�y��%��]e���=۴�S�X`/i��F輨�nwt�}�L�㽳��\�"!��1�)$}�'[�$�v�w
/�X��&�����^u��5Z�XAjqQ��z�wyϹ<�0c:������Of-�� �z���)q��[���'�ٱ��
Nnq7�`;��;�>b7K�6�%N��hX��%4���[ezdZ�]S��dNT���$����p~k��X�~F襠�W�e���_�E�7(��Ⱥsֆ	1���,z�kfl���u�܉s�I�a
y���#������Ku݊�ܝ��<���aj܉�Y�&ۏ�yq��;�'Gù`�C��,��=/���(��A5��XX,�2�4-��L�)�U'�2T�g���!0D�^�8���i��'�kn�� ���$��M%����2B�^g�H�i�.h�S'��*oAʻ�ؔ�WP_��62� �mS����zp���ߨ�����I���+Y��)d֠=��.�)�P���)1�
P���3H��"]�a,v���\ 0���kN�TB���aS��8X.b��0�+�9֠��|�}P"v�j�j��Ĉ���^���W/Z�d�z�z��5�L���iQ*~`JZHN�j>��Y����,��N�7��K��412ШU�2�+�k8(�-DR���S�_>�"[;a�R��X���0���(�'ލ�
�K�g��ޛW��ܳ����_��TS����SG���J�_Q=i5:�z_�L��2�u�X{]jv� ����YP����=V�H_I�v@d�n6�o�y��&�2��*����M��	�_��j�H[��3DD1dg�2���(�7]��@0�8�yӋ@�=r���[�D���n:6���ǳns�ƎW��*��� 9ݴ���G\�C5��δ��B>[�)eE�I��T��@2����s�{W���f�3�b*��&��wjŤ y��Z�f�+�����Te��̥}��h�^��ɹл,��cfc����LH�Z�����=>E}�a�"�[���rL!:P�#`$�CCq�_<�PP��]U�ꨑ��"D�0C�~�򮙺pd%7�,s�/��`�ϛ�'��H㇎�mќ�����[���3DU+�+,�iy��F�G�V�4�Vf�MKFF����x *[���F�.�#�c�T%��!���c��M��ur�ϰp�C�='�-'�~��5K��fG�>8pc��3����?t?�p׆賹ǐ	4�6����'�ռ;�Z6�,�I�%�<�(���%O&� 0�:?m=�MV��Z�_r���sj��^�n�S��>�QS����zl��G��G��,"U22����d;�U!1|���e����?c��rt�����o�v<�t-KY&Σ�.���ȝ�B����]p��uj=�N8�=�|��T鋸�Ve��dl�Ը�)��$.L�%�4-a<g�#!��U�ӈ�mU��e�<C�7x��b���^§T���I�ڹw�(GةsO('n����7"0;g!����� W�j63��i}bFL,I�}���M��%A���!�nB���z��P�jM�6��6�nϜ!uh�����g�R6ڝ0�K ;A�{���HQ@p{f��st�LrX�n�/�0co�4T>q�I�^�IA��LPk�AIQj���G���Q`W-�P��Xi�f�N�D���o���+�u��j��؉���*��ҁ��<em� �B� �݇G(-z��p�m\>E%�չ�pɧ��z�6U��:�L��8@�b�WjPYF�	�a&�Ó�� U�g.ң��2C�37�����`��⌙��A+�8��?%����*+v�C)���%���� �bhs����*���.J��k��O;��Ȓ���`L�Ǌ9|�n�,��O��"�rv�ڐ��|ln��E�῜Т���]0:�T��6|0��н���V�t`,E�h4-�A��fw�����G����~��'����{�gJ/�	������"\F��vd�n�S	����+��[��I>M�h
�˹�V|��u�j(�-H����q�~�%	����~����srp��2���%x��W���,�tC5H(a��z�%$�\�Ԫ�u��:EՃ2�g��˃�Ө��~�ݷ�9�C�A��-�P�^BB��Gd���S�5]@�E�GF�2eK��	{��-�;]�=0xH�0�NX���k�!�`����:�	ޘ1����"��Y+F"�c-��3݈�ŀV	C��M��J>'U�:sF�a=i��$�2T��H��I�i��F8�������v7��$���Lp����>䁊��Κ�_3�R1�\��#��V�Xݬ�c�m�o�?�q/H��{�4<M��3A�g���f���)|���9Ac��m,��s�+��4�1�3������7���K� �z��{�Kxl��٪r)�I�*Mn�-�{�sx(�y�K�\��~���(��R��.����',�M��p�J�Ћ�M�8:e�����8'�	E��Py�c���f�6#�&~�z��(}Dw�'��\H|�/8f���i�,ō.u���B��~�J�ٚ�Ev̜����sD�n�6�E�8����ՙ�䒈����Ƃ97QE�n1�+\���^UN���L�}��Pw��ְ��m(�Z�k(��l�j]��L	�%�� w�s�mP�F��J�CIw�A�}�1�UD��W�]�O�J(�1Bټ�=�Ər{^�1�kU�q���=�V�B��1�|�����2�GP^~���N����I�?>�΋�,.m�eZ�W>�Z���4oq��j��Z����j�7Kp�8�����w+dz�;�9Q�]Mst./a��H�'�u@��39���Hkg���j���;m�t�ON��o%,3" 3�b���y~��^�ǝ��h3���Up��A��RUg�c���.�Hjmܔ�:�
�u.AEP��U[y���6F;y��]�r�^�/���K���P�<U���Δ�(�����7��=�i�߁F���{:�1$�i�=}��J�l�=��@��1����,�����7�5M���!ED�� n���A,}�yWRo�ӆ4p�1m��"T���_�`//y����e����r%Nx�}G�Ã��r{zK�0�0�q����En�0�Y��Q��ăA@l����t*/z�S�`�5��IRf(�N�(���jQ|�9S� +�R���.�"�U���TZH�ɥI��v���y$�<�����&G�P��x��(G�J�ǉuJ�������5���l�t$7�m���㿛W��
OkB���ip�����&�;�x�ݲ���W��%$ǚ���.��c�w�_o^#;�M�ϲ��3���B�J���6�µ�_�ë�*g�Zށ��0	b��)�7�h�8�S��J7
�~ D�&��Aq�	D��w|a�kt�� �UK�(�{�z�5 �e��*u\J��	����ҿ�SEg\���@Z�߳���-Π�H�;�5v";��M~�D�F�!3�;�����=�ǃv[+���M�{!)t�;���Ʀ ����F���d܎�����F��
i���f�G-��Ȥ)C��|�I����(��$g��Kʮ�|阂�b�/�1?/8[zf���.%d��>(0ۙ��>C���]z�c#M+���<�Ҧw`�B�_q.'�j�L�=�������͐�A�ؙ��b0bP�Kgcd]��v��(�JX!dpo҂V#��,L��퇐5b��X��EZHu$i���~ZmuX1�q��o~��[�~�b�e�mlE R�8V�o��+4|�"WxVȁ��7=K���"4�lp@�[o��
�&K���VS�$E8dg��wԸ8/�I9eY�7�|T͢FC$�ѷ� H��з��/!�w|���4$�0�C@ $�bz��U�*���E��O[�p?_���_q/G�K���I��}��r��eG���(ݯ���io���������x?߽�������
�vސtM�.�K���֕��+��U�0�i��E�X�"�a48 ��
O��d�1����KVl�T�}��D�R��+ޜ�q����&���ΈUVrMA9�*�r�ӱ>�K�s1a�n�&If|��Pu�����x왦-D��z�
����O����Y�S��L�
�o"��8�\�����K��:�T�����Ĩ��:J�g
�6O���6�3C��"d
��F�{x"`��ӿ��������[�v��F��E��� ��!�iʻ���oJUz����\V���z��Ȥ46�����T��?,�\��*�hW�/t*�M��M&���x�FH�˦��#��z�d:�`�
�\4]�� ��v ��׊�Wr�i�����L�-����4���vf�XTh��`K{m��%�5��,���5PI)9���-��ײ��?���N��%��J�i�`c>�g�ml�
��K�ϼ�Y�y���K�[�?����P�8�pގe�xZ<�.wn�6��H��C��T)����ϑ����J���_3�Z��f}��b�Jї�y��u�"��?����U(�n���or���|�T�𧹇q�z�6g��?O������y�#	�
�1D�Բ�O�7���#e ¸� BBD�n��hb�>�H��D��%�bͧ�t�L4P��s3#;,^ru���|�<��ҽ�m���E��	�g��$K}�wY�K3iϬ�R�Nf�����q,���{�9���#�RI��e2���;��z�`5�����E�|/|bxl�J�����]���E�Ի5��q[!R�1���>꿧u�ԝ��	���Gs\���C=��`�N>#�yx�����c�8{8���ͣp �+!�̡?b����ݳ� �}���T��"x0��4}�fT?��4f�|�d_�0&r�����P(�	�p}��3{����'H��Pt�-6˝�U<4˻[{��� ��XNHyx�NЛE8MU��6i��W��;�8���gjBt#��3p��eS��D��-�Y��-/��F0ʝVM�uѷJjQ+����?�J+�%��v�����r]�Ӗ�����T�T�t1tTu=Σ�Gٜ��x�fk�Q�!*Y:�����Lq} a�Y"�a���?q��AuoA��ba�c9b=H��2�YRs6��{�:5�5:�2@L���7z�B� �/+��|>W8���i�4������\9��o?TF�.[)5�D�es�,����m� Lh u��$�指~ec���op�N�|z]�ֆϦ���C�Y]I��e�z��ڸ('bq� ��Z�A�Cy=�<
�`��NVD�%YDk���Ǻ�w�_o���[֫���f��oϢ����r��XXx!�8��5�r:�,-��'�����Rz�����1|0.-5��$+/fg'Kb�RH嗭��Q���_S*�ZCQ��^���tf����~���IP�ג������Y|�S��`�]�}��}%J�s��/�3��E�h�-k�uS� �g��6��'}�&Bڎ��a�f��|�@�{qy'��"PV��-v�1���8�u���Q���)���b�>�</�b^7��֞n�"��?�
��n����m�i�c�;�*t!��9觵���A{$k��b�ٴQ��kh%��t�G��8lS�(�,	淯p�;�s�(p��3�p�o�=<&�v��k�0�{�2�}u�k�2pk����~~���0��඄4��>���n��y/��f6��-O:H+��!3�y�XѤy�W�^����M5�7W!�7�B� h+0�@a����8A	ei�z�l�>�,v7���+��c�H�Lᾉ���K����Zzc(�H��j��*�f6�cR�QG��
����툰�bbε�()�� o�t`sg�j�=E��DR�71�p�<q0ж��kN�|o�7%/�E�-̫�C���(�0ҹ�����Rυ����]�5��f�V�fuy�֬h9��$�сi;!l��w�q�7��/['iA#3�i�P���\����I&`�V��Q��[���W������VDI���5;�r/��T�\��~���h2v[`����B�T4�Yn�h�m�|AD&������Ą
R>�M ��ԥ�ص�蟣{h4�
��z�˭�K�[�Ee�n>b�J���- }��p�@"�:6�F��ۧ�<Py~Y�����]����*��e�����|��kj&��j����"q�S�ul:�]���{��^n�K�'�k�7]8��i�q����߂~	̡��Gq�w�*v�����lfh\��Z�8�	%��΀�Ҙ���1S�-qs��W+G,_����͓L61�z���Ĳ��g� yTӐ�o/�P���[�ρ��""	{W�j,�uQ=X��@�.{���s���r�#g���?9�ŷP�Ũ�<��}Hy��QL!��HQ#(�����'�ߖx�֯	>���ſ��׼gs5�6���i�]�E��T�4 t��n$kɥ+,��%�y��XF�_��������#�؅�PŷjO�ε~�g����
��E�� �A���L��ZfX����/�/^�'�0������������m)k��I,I�|�Nt��lE�<u�	�Hht��g�)Hυ<s]���9�艽�-�Q챛��I�K�����/yi��[��狗Yu�Nׁ8f,N�Hz님ϱJ��[��o���(�	��8��L�}��s�f!V�Tk�O��B��gl�eX�ef��\�(U�qfz
3����J2�-e�)qT�/,Ih?������xQ�;_8�̫��B�BZoj�7���Ct�eJT�Q��"���l�6+6|h��
�z��i{��L���m¦���QI���(����D����D�3��װ8�n� �詪@..Cb8���ڬ���HÝ�J�d�4C�M�o�r�V�y��2�♖�k��b.����o�q��,ܐ}��'��I����c��Ӏ�[Y="ѩ�\A���}�I�Bز�yE!���t��sH,���!�6��6�#C6g$W�ܱ��P��@g�`r_횥���G���f��R��Y'f����/�{k3(2�^��M�iV߇RNΡ��s�I?��Q��D<�|5꿓I�)���\��6��i��g��]��E���?��l6u?7�yh�k,���ଆ��d�1k�*���4��~0���Y�9���$&А�A�D���9þ�ղ&z�Q=�\���1nC�|�wS�����(�=⋍�uF�Ϙ��9�F�/�(�
��� 0�t�$V�8�M�EV�X.`��r���K���f��v�\|2��p_�<s4��~���c~aZ��ؾH7�v��⍙ӒVAA{��<1�j6��O�����UV���m����]�/>����x>��+H� D�*���{�`ק����w��'��Y��=\��X�}i;�4�|��
$Y���c��ܓ��I{�Z��s�)�|����04��V;-炔�53�hs�6�O�+��Z��$��| �kN������9q�x?��j���3_nC�)d���Z���{f ��Y]�</)�=�g��c��׹X�
o�W��~Ue����R��;� V��﵋-�g��b��#�)��WsdO��Q�ZW�
�c63 � ��0���I����"�oD9}[�mz��M��|��q�����FZ�9�!�:��S����{�F''J�;����b|E)�;�� ]E-.;K��0�{EynF�݊S�ӸUkm�E��U2�Z�L���a���&�l�phC,���o�;ț�ɊȐ�xN��>oO��Q̿X��"�DAzbK������F�
^�t��=���<Fk���?%~X�º����{4�;���3��i{�Q���h�K��""9�����n7=���9W�sub�����C)mUvy� ��cL2�oǛ���f��e�T��f��;��]������[�4.w����9lX��.��l!�!�!넞�0L��؀�)�������>��/�K3�^��Kk�E|��<�Q��q�����Qv�H�2��㷙��E��M��zl�q8La��j��E!�q�����q�dD~m��I_�,��ִ1ʋӜ�q{���Qi�XU�c&T�m��*���@�� �^���>�^itMGXf℮�0x�� @�����=*���ľ~�o�|mM���&:هS�ϻq���n>Z��L�o^����]rlZ�("�=��Ft>�{��:�hD 1��~h���=O���Zž���ӈ"~��.�3g�<�U��:��,hR쫛�� Bv7�9C?��L�Q�����%MT=(�x���b�����@�3#���|n1��uG 
W/8<�P��^3��+���"��~==��R�6|&�7ޔtĤ�
>�L�	m�G�O�Ż;r���[��0q�7�MX�&��=RT�.,�����Ķ��8Ev��Ԩ0���~�O1.�Cs	�$�[0:���Ǧ��GMz���R[!D�cVK		{6�D�-��:%���0u,���>�mWǲ�{�wy���:j�}3o�.8b��[�Z?�ڭ� QX���dlrnj�c\$G�n�����Ɍ%�I��kL20�����h'�QN��T��!�R�
}0,&��e��	C@��W�&��R�0���B@���4?�����n:!�Y��C}���o?��KWH	P�D��Q��gj��S���jj���<�I��t~PsO �h!$���
.�/�����X=f*C���X2����:s��7.K������ބ�}��P
A,u�f���'�(�6u���N[�%�>ō%�����jW�yv�t l±훓��*	�ơ�",��7eʋ
�F*������~��ǯ}u�A�_M�g�c;&/�۠��EY[-U)�)�#�[�t¨L;�$�zVMj0���� Db�F���;�@	%6�	�ݣ����vwO�
��ĖVoT�g��MGRjQx<�H����4o�uu�j�G�7���G�Q���m��\=�9�,o��Ҩ�\��}�-�7��4���)�z+a)$���<S����ڮg��X�N,R�n%��2#5���FS��y��)���*��İm���Xi�Cl�I+�L7|`����Fr�g���ȳ��ז��|����QdJ�bH�X�l#D�O���d�V�w���rf�_�h��\��ôf|-*|��ǘoKw�?.�w��/T�ym�\H���ث����K�Bp��(���J6m\pNU��_�	 H�c4��v!݉�H9�w��"$��0ϊ�˗Ӓ��THą��h��cK���h@�l��[���:I�N�&��6Y���7��C�6��e��i��!��+P�<��=�5i�����gݏD�)�*'�TЂ`h�`EL���4���M:?r3B��'l�|�;g��p>/�;�酼��F&�.��렯�����U{Ȉ��{���h�gM0�T(�v�3�!=hfp��M�G0�9�\I�e���Pc��ж����cS��3u��kF���;�|��9p͔]\ň>Сy����w�*��U��d>�t
�B�^����(�w���?
�H��gz��IT�m�7�.����T~͓�����wT���`*�� (�Q�@S�m�F~l9��w��@{���Dw�
P�.6�~���B��{��:��*��:U�{������E��В�&���1���{j��8[�J��3q�Q�w��<�H�s`�\�˱*�L�Su+=�-f���\m�d�-!@��෦��;���X�����n��v�$	��Hlq�+�B�'@��*�sr(O�q�z�����|
Qy,<�pfPS*�=`V?*��쩣�Is죘?��'	�͢,�9�s.���:$(%G?�����L�f��:��er>:+�H���\�����c�t#�]��JD�;&3�	f����e���;8�j?�6�Z�W�_��K��ԡ��D�����m��7�d�r*�y'Y���+޷OŜ��U3й�~M;o�������L#���a�h=7t�7q}�T#RV�C�~M���/��KԒ���r�
���-V������;���"C��W��oT�nDO'�I�g)#ʂ8E�����r8�?�p�dY�}������DT�L)	}��K���o��U{k�m��nmo+���q{�W�$�����	�sn@��F��>�0Hr7ID%��G��]�Ϻ�����m|4��2;W����o�|�6	������%�L��k�;w=��w��e�ˈ0�+v�����\h�b��}6|W�%[��S ��O�^ܛ&1al�f�R��ݠ�l�~0����nw��PY�*CLћ�|�8���UR��0ˋ�)q����	�>�dS�s�s�dFio��R�������܍�����v4�l�k6x:i"����Q`*����
Ӛ�<�~	V�t=���j���x����~��yj[Z��%Z�㼷=�Gg�FIܬ��2�8��f^P2Hvw�=�5�4|���8��D��p��X�Y�v�<7o�aE�Q�T��N�?����[��.��3˵`�R���!�,�������@�1�|/2����Gd��Wu��
ȏА�n��>R�C��<�|B,�ҶbA����^�f�d�ܠe�g��O��lx��Q��}Yw�
zy�y|��������H�.Q��N�I@Q�C��� ��Ȗ!���R!�Yq�I�u�X��ާC[��k7��d��jVٰ狑������x�(���1".֑��:�+J�%?���;�nZ��hϧ�����r�Њ-5�ӅS}S�%Ժ8 $ꩦ��b�s�(�/��P�#�Z\�}p��`�b��"�
�(��>��+�)����f.�쥜�e��{E:1�K~=wpI�q�o�e�