��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw�a�[W;���(���=�0�Cm���!Y�h`J��^��5�Ư����|e<5�����RM�p�a�'e.���ҵsV\��K]��W��i�bR�~��Q�P�e��ڔ>��~f�[�v_s?2���D3�$���Ht��Ct��͢V��~q�6��7ˊe!��u�NK@\�F����hӕ�.#��|�1F�BL��(K�{Q娓���ɟ��K�5��M,oA���:�S���7oA�H2<��،�K�H
!�28��X�`�bUM�Ԡ�[I��N��ݔ�s2�5�pp�4��	���맚�Gw��A����EH���taV>LL�5����_�E8h�.����K$�j���^]��E������B��L�IK.S5�NKq8A?R#h9OS�9��D��S�y���#�6�
�2�����!��8"gb��8�m�#���\�!$'a;׵�s�����BT��I(�	;�a���mX�C����|Z��x1� �[|���b���`Xs�xYs�R�kg=�n��%����sf
%�!�ҫ?3�7��]�^%)�4����L�џU�����X�Yh�����,�.����)�r%��G���~sTa����Z����b��;�Tlǅ�!v~��gg�&}F�����
�xƪn���rq�g�:���@!�k����#�p+��0�ٕ@����E_���E?!y
��ٰ�l�]����h�2�|���,օQ��<?�]���T^G�	?�d��8��vs���
�k�(�!o�T�Z�H��.hh���U�����Oك1.]�ʣn�`0}�g�x�";>���i�z����-Sc�x����"��A�g���^\O�"s�k0whOpڈ����gSKF�Ё
�1$mP8�-��j�d�zU�+lr�-�jjӇ�~_|BF�G����ix'דT�(S%2,[���N=l�������!i�Y��עH��_��\ �2�������������#�5{r?�X	R�[���F�+��IdRnѦ��S2�[�"X�*�wm%7Rr��n)��X���+k�Rg�B]-@�Ի��q��T������T���3��l�:��B���ز$ŰspF<�gפ�����j�/��Ç<���Y�c3�*��>g
��-)���!�ab�{c�v�ȇ�Pe�簄�J`x/�e[�O��ѐ1ځ���?�QtCN(�{)����pd0�n:��1	�{��i��b��5��v:��XXZ�8Vӊ�XI5�C,֣V��a�Qu��)�s����`��4S}[O/R�Ag�y`}~�(�i^���_����]f qW|����b�S� �1����"j�pUUDR��ߺ�>��ׂ��{�$�7*�(�p���	�Q���}�1��ী�� ��ZQ���i�iRP�:��)&���w��q�+E�tp�� 7�p=v��S?�����>�9�=�-��d�n��Lޘ�	"j�U�Z,�^þb9�r�%@,�͛��W���׬A�Кv�|�*rF{��?�ȁΦ�|O�k4�Gq$p<�p��b2^�N����+֑��d�a�8RY�����#@*�����0P޵���x���-l����%!���}�6�	���)�O���(�
��w��<S�n3�DT�c��C�HvЈ),���>�T�z�����	�0bX��sy�KI�=Y`�Ѝ��|cɇ��BZ�~'��dm��o����j<���6�X��g%�� �����S��հ４I������*/՟1���ځ]&nR��l��?>�
L�聣gܡ62�R@�
{���H�}бu��Ef�T
vt����H��������q�g�;�|+l��5V"g�a]��}������?�Q���R�7Dr:��M��#�s,^(�YŞjB�PN�7]<���S�x��W��!K�ʚ&��R9B���)Uv��_=�<	��h��=��0�&�5�Q��겥�V�we�C��.����#���*J�l��r�&�,�N�	�
q�Ky��v�J��S��b�#�����1=(��fӟ�K��:��P����*�͖�'��"R��8v����n�t��Hd�Z�Q0���@�����̈y��V�$3���g����{�E�?�D�d��.��Q���h3���%��A�A���ꌽu���`�2*Gnao=_����X$1s�X܂VS�!
�C��<m�0�zBl'�����Ix������`��X�L��"�-���Ǻ��\�~��e��IsQ���ס4�o��5-�{5�������1���{�G�񒵸�Ma�*����;`8�÷��Ϝ�( ���93��o��hѻT_�!��-x��N�:�!ʳ�^�A/ӟ�ZQ6׃^�kX{�&���IYOs4�����B��b�0��Bh�r�Dg��[�cK�9oJ�(�<ki�zE	(d�b����"����S�_3�5��ߎ��OF���R��_Y*
mY�홭D���]T�R���8	&^N���6|�P����cQ5ȧ��95��j�-@���B���>Z��g�`�1��s�yLy��"�z8�0&b���t���(��3.Xeoc��=�q�Ɇ+�KN�;;���+J�9UJ�-WS�������$ 2�@��@��9P�*��[)G����ca"`��x����ВT�v@:�n;��Wh�{��?��U���Ͻ��'<^�N��<5�K�'=7:u`�����h�T��b���:�0�AT+0���T�i�&�#!�%x���'V��G�~�8i^tY�e��4��R/k$4�Rt�.���JB005dEۋ<�Ko�F�N[��:�
�8��j�G.r�G�����A��y����.�԰ǾQ<����M�S�$��J�@dBL��LG)3������i��bT�j��:��}�����ex���{ q��}(h�[��0H5` l�¸�;"�X�ж�z�Y�o&�AJ��ތ�v֝ E��V�nvQŀu� �.d��ph��'�ǐ�Q����݉G��q�k�U��|%�����ӛ��l�+�1����[���*����@X�J>�Z�n��zy��� e�,���O��b����'P	�;��<5
܅� Y[4<*VXA�OV����X9T�z��݃�ՠ�}�u߶�Ң,�� ������.y��Tg�p��۵���n1����
��%���ZpsA�Rxx���Nuv2����5V	l���v�׿O�Jy�#�u	�>+jn�a��2إ��h��]�e|3
�E��ב/s�쇘����	�W�8��vMW?�l�-�;C7�
��APk0yQ��|�8-����xI0�c�����*��h_�J!����A�����gK3Ezƀ��+;��4�,俾��\Z0#璙"�|G�ǰ=C�;�_�p�J�bR�S)����0��F�B���S����4�����(��5pB8q�������Mar�e,�L��t��p�?�����+�����W��p,d��Yaק���,e<Y��e��]M`�m��{u��cv��l���2jrM�������8;RI�Yxx�Z\c$킡���#����^���SW
0����4�& U�(K��Ag�fw�1-�]B�/�MwS}��=��}}}U��U��kG��n���L ��E�������5q�˶k�&�`X�<)�O2�ZD��4A��su0@���=J��授��<�ZY��O�{�i�x�*��td�ܠ��y����7Bnp�N4[�b=��ST$T.47�M^�/�VpUY���/��6d�$��
.,����b�]�j��VM���N�˿q_p�����m%�K�����Lxr���r����+%�1_D��F��bj	!O΀�э�$��#�;�\�NvN��fmе����ߴօ&qG�>�����2ӯ�G;s�������w{��>���£x��߇
6M[>���^�:wƣҒ\�$S�T���A��`�#�I�U@����2%P�g m�}F12�<��x�]4�^B�4^}ۖ��P�	E��ݑ��&���t1��%$�UzWh~��~�l8��KI=\It�8��;��Nv&��恀��)��ptL؋z`�*ݴ��dsۅ����Sγ -��$)KT��;L��Ʋ��Y�;�X!;��>�T��o�O��F�:���C9l�s�T��u�l�h71���2�����eg�^r�+�4g3BZW��5�PY���%���> �<Ps,_:e���K�R�,�Q�Y�/(V"TA]��.Pb������$ ڃ��A<���l��_o$�?S2Iu�L�jY�q��QPط�9�W �:��bX%|{P��V>=��)"�#�����]t���m�@�����u�$�݈�͒lw�V Y��eE_xwE����5��O�^��NY��V�<h���^8���ssUk�.Z/��"���������g�>��$f����/]���/����b\��W���k7
�
�~w/v袰$�c�GJO��	�u�+�vZ��H8�Ķ��ـm�5:�)��U����N�<��'_Y�fVD)4K4O��c���J�"�b�HÚv'*V-��#�~��?xY��;%Q `��cJ{�3'�`Ó���!�1��Y	���P��1q���}�"������o��Z4>�?�/�n�,p�k�e�R<����� C!q�er/C�_J����6�R��8�X�c�����B�g�2�I�e*u�ǚ������[��z�Õ�����?�+�U.V�xO���]���l^@���$Aw㥨o�J���p�9����\i�>�M�~�^�V�x�B��fC�7�Z���fm��_v���>�l���x8HKZ�C�C�����Ţ�`���S���!ZR1� fJ�/ҍRS�5���bx�?�_���$}���᚜^�G�׎��ͮ��C�/e���Fpz����(�3v3�eǿ@[ӫ�B�G�.�f�,�e$���<�fmŁS�zy��:vW6^N-*{E�tP������^�	D��F
�?�l�_���j�Ԟ����S��v���j��к�bas}�m���w�4�wd��ܱt/�mԒ�S?r�X�;(��M7���ur�_/~���� W�ji�@c|N�ۿ��'n<���w�V��Q�� �6�tE.<,G�'$o����H>j׾�2�e cT�O��O��b+>pL�*�4k��RM�o���DZ���e��S����WG,
��*L��.ȣ��Z4���X R��Y�s�%�M`�	�#{:���C��y_W��ؙd��U�M�/�j��}���B}���P�"���D�������\�პ�՞,4�L`F+Y� %�����gh&�B�n��,f�;.Ns]#����H���K���E�ŉj�� Z�g������̓�n�<T8u���$�+4�l)��HHL
��m�'�Ol.�`r��@�����"$���-��&�^D��B���zD�TE�|�	����4.]Ðy�Cc�9m��fӰ՘'����Z�w��z �Y%�b;mw�L�G�)���s$/���5��6�sV<hG_��ws#
ˬ�B|#q�x{�zR#.��=�q�ns�����cF��釼vbgxH/��7�-���D/v_�b��U$���zj����PL�4U�_Zss;{0'(F����;M�Ok�k5h�Vasw8��:����v�%�>TC�:/��&~{PB�B/xww�`M&{t����C^O��:(O�O�8�U� G��*��@�+߸���a���Mk}S)���)u�ܹ�95/�!�f&v��FMg�a5t
��sc���q�#�A�h�34�F�/6lH7>�J����/)�r�&��F��zXh�V��z���z�K���P���"�6�g�Z2@�����l�O�G�6js��Ue!*���v3��-��ʪ�.)W�ic��4�����3��^Z����5�y�KG��r����Y����z��Ͽ��Z ����U!�^Ĥ�N�!�H8(�q������L�jG\1<]�uG���:�/ �q��v