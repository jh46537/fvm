��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�Y֢�08)��k:�ث�1��=�1��cO<������9�5�^���W���.�����<��_�sP�x+v^�Y�+(���TOŐ�ܱ*R�8Fa�2*1��k+I�,��K/�$��[�h���Prg�1?S��x�7����yj���Ϊ$m">�i�1�o*L2Md~�(�)/9n�j�߹uԔ7�w�\�;����又�z���QJ�ou��p�1�rl���<�\��~u��}T�g�]m5�8JECU#�ř��B�����M���1�8�i�}U��YΔf�G��5��z_Oi�/��������G[�~�<�06�^�A�ք�U�9S.\A��-2�W��!k�ȱ��<W��JB��F(.G��օ�y���O�D�C~�W�ѥb�&uPmUt������S��9��V�C��M'���8�G���Pz�� mٹB�Q�(�';|���/'�;]�AwW�PN����%皋��a�HN�R���eFXB�x=e	�K�����~ ��o�nw+OS������l��w�}�@������rօq�(\.�v�Qbw�^�oA8yV�h?4��_st�Dq+-��?�����>S�!�$dvtu�qx��c^���;�L���y�Zf����g���Oʣn�Jm�D����ɥ^dbG����Ц��46ϵHQ���3Jmz�.�)F�&��⻫�SC�,����)��t����;��iadH�a'g�L��o��.�K_J�0���%�#�1Wr����ZGC� 3�fǇ����9I�$�&���Ub0:<H�����΃��*Y�F�tb�����۸�(<��pe�aX/�v�|4~�S}�Oo�s����6V�ʲT��2(��J`�;��,u[4��0��r)��X�Ĉp��%�B�6:y\�w�Ѥ����6>d[��" ��P�Ht�P�r����0����X��vO˗Xs���<���!��Ћ+h��6�=]~�9��7�Z0�\�@�C�oJ�x:��:8iS։ӪA����^�4�%�p��/�4��u'���3�H;&���>�Ɲ9�:=���Ϙ�����kz�����Z�b܈���� �fm��<1p�DV�_�^x��h��ڍ/���9� �1���"�}�2��q����S!�Mƾ<��f9 >��q���Ǭ�S'e�h.0Gu���֓xfr}n��L �̂�p׫R��(������)�I�*HԶ_��{}�4��n;���
�Μ�[��~�
������g�D���y�H�Q_��y��Y�O{ ��5��y����^���ZX���6�g���7�9׃ъT9`g9�xt�6 (����t����9�n��Z�n���p9M����o��'��5G���:È7ٙ�NG��*7ٴ���e ������!��"p�|;η%����}\*<����(4�y\1@�;LXQa�1����Se\�mf�֮ \���Ył]!��(0����٨s���e*�LR(l�9	Y�gm�L>h��j`E'0�W։u�%�I�gM��c10/ǫ��lN
I��7��&�l���9�ž�xᔕ��F>�Ah�hL�)�p����dJ�n���]�P�)��s߰+���g��fc��L0���B���?���/�Ga����'�S���nԸ�0�qǁ��﷐T�&�����z�t�\����,N��������x��qEK���U�8��N��b����l*;^�L�|�ZL�Ցi����-�=���W?�e�<f������Ah�4/�5��̄�4���x-��M���2�+�h�	�H`���aR�Gg�B���%�������mcI`�{7���۟�����b�d����w�0w.F�in,����h��o>�}8Z�O��y�/X� ��߆4DJ�����̝��1�5���҅�¬$o�́WL/�"�p=��9ފE٧��N�����">���C��?P*��޿/|B��o�9�z#��%�)��=����_�F@}��UA���X!��q%Ui3�;�G��fEl`r T���a5��Q
�9��c��Ru�קd �l&�'j~�@۩��a��EtC�"q9?���3�-Q82E�UI(;�q��(%q=0�Ս<�I;a�"�J������!�㉑@�d��z�{�>l��ī�0	Y�}`p�t/�^��?�O�e�6���ZQ�EB���/'h��ғB��
ۋ��n~�o��\�jq��v���@uY��X�c��V������Q7˄O�*�M���Vy�!ӹ"�C��C��bJ���%#c�e� 7͆���t5�+5��ER؃b  T"Y�d�xj~,CS���1�R��udD8k�lh�Gk�-���Vrd���z>YW g5�`��$`d���c ����᠘w�_�L0$lҠ�^W�T`�����>N��J��k�04�vQ�IJw͐���柡}�=�&=�>z��윮�� �5fP��TB���͗?�%����4���o$�x$�c��R�ɯn7�~�p��9������� �8�>Q�Օ�r�RuO�e����F3��ry��'o'���(�*)�jt��`^��}꾬�
��Z�kn���v��0���l߱�2��M�oH�0�59-<|.G<���H�8a����Rrn@���i����W��^јo��'C�t}�࠾� &���7;|�*b]��n�}��qa��̘�.k�[�-�B�R<&�A��W�O�}掻Ŭq�Ԃ�5")m���c,B�SWx�n���/G�YLzU �п��^�l`������'���_�KF��B
k"�rn��+�ʲ�� <�L��Ǎ��a�!��*W[1ak���]/F�@S����ؘ1��y������iK=���bNT��h�p,�h��K��0r�3���<�Ð
����(�3P���3�B�d�� �.��%�Ԑ���GI�����9�JDa���[�2lPc������8�D��A�S��K��x�Ki���Z�Ar���/�m���[��o��;&?��\N���Y6�x��SAÙ��1�Fʈ�@V��("g��;K�L�l~/��5b�vE��9��thK��@{A�v��_UY�ΗM1������G�)k�S�*y	E���X����֡�{\�r�� tۦ�YL�ϟ�G85��BKf������	8��%���n�Oe�D�Pݤe=2���-�ո�	7�n-F�3�JI)�d7JY�ZBȣ02g��O[��Ic�5�0�{۵���^���K����(`ØN�S'w��}Ή�ד�Y��9�I��`h��aT=�*v��={�M&��|Q�id��2��	��Fw��K`�_�T��Y�2$XO�=.S~�Cz䊩��v��i��2c�N����9h�k��_���t35���]�ͫ��`B41���H�m��b
J[�8L���2��j�-I赚#�[��39�V����Xj俢�bn@�
\kv2�V�����`�s�����ҙ��rqb�,���3e��@)$��޿S�w�CV�;z�_ˆ�GV?$��8��0�Mi׍�nTx�ڻ���<�Rŉ0D�^��Z��S:,��R?��
�$����@�<_��V�h�>�'����C;��dB#c5����a�@�����Qp��$,]������	6}���EW��N����qL�¢ �og��"a~3ӡ����㗪28��B�
�j�����p�F���ar1-����}���'����S��1T�q4�.X1��O𫺖�©��W�v��q]m�r�E��ނ�R�^J�}1��gg����M=���,#��j�(��;Dv����`xfs��2~y(�y��3�j�M"{���e&�o�{�Y�s-��&��G*a�ʾ�V�߻������[#ކY!��1
D�yb%@阗�r�X-���~�v�=aKV�B��}U_����Jq}sS�*J�Kw�A��S�e^Œ3��s޲���7��.��� ���Tw�	,��x�F<�|n���Ԩd��f���y�|^п[3�i3��i��lIX觔ƹm\�{����1n�\<��
���4ɝ{I.�GJX����;l�a��ʧ�?5����O�A*'�97�;��;��ҵ�m�J��n��"���5U�E�����cdkЗ�D�L�Q�r&�Q#�953�B�x�9"9�M�̪:��L�Di�`��܄h�A_�G���Ϥ-WY3׻��'ىz�U�}3qDo��+�y���r���HB�q��7�^p�{kV�R�1
���i�?���p�����#V�v �;�k���#�5�1Q4o;Y���c6t����391UՍ��IYjde'��[�0L;?Y:Q�}�n�wK@�K;&T>�i;��e������Vڍ����ő�O�?�m�-o֜�%u<�����=�"'﹈��E?q�V���>c:[�7׬[W�A�Dz��nv�{F���_�-r�Byu#�P�3ܙE�w�50O��5�U�\N������A�{�Q?�����k�/OqW!B7� Y&|�7�nTMA�T�,z�'uJ�;��:9ǋq-`￡�-",־6�r�+���-��ӱ��\z/�E��Np&�T�Q�S2�D�@�^ȃ'�8���tX�/3�^�e��c�)|>�$ a���*t:������[�� ��Tg�x@���{��wX���^����X�Vz,?H�-�]+Z.كيF���iHS&��&�&VRs�~��T����թ�>�\�z`���uw%g�1]����Ǣ���&�9G	V�<��2rGujߏxcTt./���
�B�L�F$:�BC���!�!|P��.������%�q�~ǚ�˿-'#�*���O���@!�Zg��JI6�̡���=��V"eY���x8��W)7��Mc�%�b���wF\�ZW��}��$�)�u��:-7_��i���S�@PoJ��똪a��]��
��f�,���ܵ�����[;<ryHe�j0�a�.{�i/��nc�m)P5�����Тc���HXf��ž(	Bhu�W˃�}Wy2�Fj�!����r�#��
Y���kz֘��|���6H��+.���׸g�[i�{YHo��� ���]�tA���jNu�=ٟ���-f�頓S'��H ���:�OV�	)#$O��g��&#�\n�����C
4F��n�3�����q��,��Ë!ks����@��&Y�DeVsw�x딋<�n���*�����v��/Qu�,dshCQDX�J�tJ��;��c�5��E�'YX��|��	k�wj�����)5P�U��1��9*�lG�%���>��^�C�h��i� y�o���#���O����<_΍��I�/m����ҋ�F�����4���8���ɹ����	�HC�p;8x�P��Ǎ�1Ҩ\9Џ���aQTgS�~q]ìC�k���Oe�{�<n��f