��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�Y֢�08)��k:�ث�*e�(AOg�X5����!��1��-Y���	�H����T�s��w�=���ٹf���aC��0�VO�JZ�ж��N{ɣqĐҡ���
 ���
.iT�4h�,e���b+t$�d����Q� W�^��b4����nI\g3��pE(�;�L𣐐����|��x-0}�ZE[�Q�v�]O��a���`k���,��_���e��3��;7��� �M�}�:RG���=,��G��ж��-�j��<D����H4�(t�!&��Џ�@WD�cJ+�g�7/U�HDLG�9�k�b��<tu��6k��1�!�*��P~�K ���l��)�J��A�^/T|?O��C���.����g��Yf�x7^�+�>x�P��F�-���w~�L���wЏy�'�f'�:�לW��,Ҿؙ3/��D��ߗ�����~���jڍC�79k�y��4�1��7��ϗ��1��J4X�����e�m^J4\�X#ƺvn6��&��X��g����[# ���ϯ�A|||�,pE���U�1��?���i��K���QS�R�!��Q�A`$ �.�=F �%j1XVc$�����
ގ�	 z֑���]�T9
��y�;���B�B(��\�*q�{��*�*�j�w/����vy��E**?ef7:	+�֪It��h��|ôΜ{~Q+��b�e��g��Qa�P�����=7�)�9B�'����%��0�ȵm���1t[����KlI��P7t	��b��w���yGٟR�Y�z�ʧ�=�i|7ί*x�y!�@=ӱ����xP�I�y/��$~wQ.S�K������{i-]����_�&T]�*���C��`�%vW�����4��@�=3����_A�!W��B͔��`�	�y� CT��D���)�$�>��6@��f�h���;�`96�$�B��UPm��C���˦��q�Z�*�#8nr�ٙ��p���~j�� lάa���ۺxG�$	�/��:����U�1"�k��`0�?=�^�j�q<�![��p��kC[
C^���K���>�ץ�k���`m%��,�>��&)��"�!�IW�_�x�x�sȶ0�̪mn4��_����+d���4�����=.}��	G#��8�"l���H]�j6�:�IHl�|��������fs�����t�mܔ1h�c_�P:��`/�
�j����7L�	Y�7�#��jȑ��_'���f6V~�{��	c�6�C}!'��mz^�s/�c���b3��ֺ�Z����,��G�&9�/��dU��y��S�զ�:��_����5��m!yq���q�2t�$̮ �qr�������ix��2>����<�>��q�}�7��K���a'[��3;pvq��:�p��l�ĕM�]ް�Z1H��~��C ��q�D��=r��j�֒�.��D�+(y�X���V�������l]Aq���_���2��I/�>�J�*�����fgA�Iݾc�UG����%�;:��<�_�����T)�H
��n}q�&{����ŝ�
�z�'2-�=�Վ��6=y�1e�ځ�v���t�p�h`Ȱ��.*�?4 ������sw��wLu���6���r��l� �4��c� B�je?�N�v���ޡ+'[��\����l��-	�N���A�(�NA9_��L���x�Y7k4�/�TwQ�(�ޗ3ɒ%��n�lE>�'�i[��O b�z���G4 ��`Z�E��=�q�C����;�6�h�Z$��N�Z�t��K��\�.>HP�W�[f�[��:�,-�tC��%)!MS����w�:4N�4�#V�/����>A8v�Y ���s�I	��4"ج?�șXA@^��B�{U��0
3�;��k�ȴ@	P�z$����F�Vә���Kd gpD�P�
Կ��I0��єI<(��4>M&��;tmn��u4il��w�&��F(�(ޞ�o��A���nX~�8�� n����l��=��o��Y��SOf�>���J���T(s槻=��s$3��8�}�o�̱~�xO1R0<�F��c��u�ok�X2Ն�������UYu7�;@���x\�';�,����Od�Ah� ��b�\���N/��5�!ļ�}>O�Rtn|!�"���B�֨P{r޸93K���T�t� 2Ⱥ:5U��)��sP���Q����׹z[:�J�_5����e<.F��D]�������q�f*{��DG���;�
}�R��-L;S�05 �р��$>?R�kק�P������U\�������'l���^������Y��dLP�i�$�XT��A����z9��sF�����r��:�P��;�0�C�POQ����Mٯ7�J�T,��4��5e�H�M�!��_E�[ B����\�I�j-�}5��X8��,�^f�gڷ�zbF�˴`��97~\����NRuH<c�n�s�%_.<s��j��?�Z�i���(ޯ�qc���q�t`7���+.�j��������#�|���V��b>�<���ͪ��~H��4Mz����3�~;�^[��o��|�?}mhY��^��oO]��!F϶k!���;j�}�W���V��!��e��,�Gå8\2v ϝ�^���H���f��o
�g��Ϧ��<�+���r�`*�S��dF3�č�g;��qKF�Y;ZJ���]�;���������{��X�C�8�&*��3��|H�����cΚ�O�o��lܛi�bOṱ�B%��x�����:�p��V��<��)
Վ���.���T�]�Ŝ2�./����<k���	'Ao5�}�wa�Kk�:%-��d��������ٔ;EȒ�K/�x�3�>�p�ɋ�wX.����]��|�y ұm\��9V.�ikc.îP�_��vж^�J��?�(۽��aB�[��~�tڌ���N)�U7�w&K%
�Z���S	:��9WW}�DHE��XE�{OO�{��l��j0�X��:��j��_�v*�.�/.�c8�d$81�m}������%� �e�B9��~��%Y���.��M�5"M!pmT*�9'A�����C�$�������|(�w�
H�������J�s5@g���h���b-��!�y�c�F�?�L�U��ߥ�>�~���	r���23�P*���Z�1s�����oZlغ���?��<6ҌO�RL踌'ypTD�����-�Q�R�G��y�H�D���"�����s�#�a�����tT�	U��垍RT�u4��,�Bk3%v�5G��/G�(��mJ4�@4+
��ͯ�.��k��E�x'pfQ�ߝ;�kc�g��-Rx�~���a^�^�A^//ˍ��d�^3F�	{:�{���g]y�}���D��8��W�P�f����?��|�$�&��5�!��ԍ�r�ʥj׽�4\���Zq5=�N��WdhB�{;��~�-��Y��XKS�u� �#�H�~�j��@m�	��;�n$}acs`�:��r�&��ŵ�E����(��"���g����tE�f�Q�J)�טC��z����a:B��{Q��!M��Y�ٕC)�â�!�<m�5ʓ�2g�89�TEV�I��[�v�#�{K�n����TTլf��>�¬mᵡC���K�|��X��Ie`v*:����9�sؼPT����sBc���,��4������+����!Rb���	��C�@�Q��P���!�ꄶ�����r�oH8�x��AV`m$#1�Y
%��9n�	�=,�X��f��J���B�FJ$?�T�멼u�S��t����%�\�f�Q�"� �"�)gQ��8XH���ŵ�w��{�(�Ҙ~������ˉƱ��R5�'bq-���l��0��K���s�-8�I���Q{��[�a�uĈ7�c�~�ұ�ڵ�W�?���揜	��@�9�3??��˯��V��V����y�B��ع �G�
~z{#P/Y��B��! b[6&��
��4�OF:A�'#�'9T$��M�/B�K1�Z���e;��k�?��K�7��7��h
pb�m]��mzqc0�/�tm-e@�&W�
7��=@8d�1���;�=�?R�$�fw�o�l�O�([,篡Fg�K`UP��2X��y����x�n	��)7�Sh��&�n��F8�;�Xg�0F�v�"J��7A��t��W�,��PK���:���SN�fD�h ��oM��D��,0�7�?�I(���_<1�����!:A*/�aH��T�P��9���o���#I��$B#_�\�~y�,�<mG�ܽG��ʦ�]�� (�[��*��]��B��
�]�43>9���U����m�3�w���{3G.3Qk�S �j� Q�iso�/k�����<�nm���
PCV:wѝ��s,�y��uZ_mɩ%��6�m��>�����p/��7��?��@�24+|I'�����hU9���g�UW:C����3�(��@Z��?hN3�v���S�uf�0"��W���_���ݧ�لj�"����<�lL��=��-� �,��JuF��)k��d��	���p�X;���"kfa��S�Y�����k������Z�s��^t�F�3(9�r���߽_���<�+��C�7�{H��ڊ�sE�ϒY;oVQa���M��D\��³���y*�&�JU7��mn��0�.~7Оd�1M@��R&�]&����GFl0�+��ξ��>�%���sG�Sb��%���jA�l;l�� `O�v�#�|�%�؟V�]{����jj_tۆ�R�BGz�64XLc�+М�;|��J��.c���,ȼKK'3�Q_~[��r4w/
��Zj83P)��o�u�0�>d��_! ��t`k������[8�»��F�C�䰶h��%�
�v�X�bW�i��e�%���,�S�� ��`I�s���(@|%��5��/�b�K
[}]��1����­@I�乄��.��1�ݘs�'J�B�`�W���<3<d~�'��,�m����{sNG1���z�Q��D���c���e�j��-�)7�\|�p�s�1m
��'�5��-_�|�����ۨ|�?䆗�X�j48� ��!&*N^�Q�