��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�~�������8U�� ��Lll,�3?�c����~#Rl���ю��Ba�ĥ�>Ҽ	��a��v����'��p��`9�?4`��6�&��Y�B�z%�,7��/�J/4�ǑCZ�-�5���z�y���Ɣ�k|Yџ��L��V�C��ґ������H���ϲځ���U�s�����g$��-Y����9Xr����`��+L����a��(�:Q�c�&��,�e'�B'���T�RAu�O��'���<t�7�T�L"�6����0P.V�5F�I�N�i�.��x�c�ًӌ��ߌ�˯��tbW b�
>�i����0�Rk�8v��b"��e�F{��$�qk,�%����'�)�'��Sԑ��u�˕���dV�ǍCa>3���6��C�J�����7 ��3����K\�� �܇AJ�	z��|,ŰS�a�'�C3�ǩ�ŭS��pmD�n?�� ��1;@�t!m�v%������qe��S_(����I�_��s8�Ց�=�O��<uQg�/��
�$�[����R`he�VL��p�8���G��څ|gs��$L�ϐ3�<��Q�Cm���o 6�Y:�\�҈���{�TBb��ES���`Ɂ���]e��0Vl�v��W���MLt4�'-���)x��փ`T������v�U���Ŋ?_����e]��
������NK��Jd�`����p0��5��gv;K��q�,�/ (Z{�1V-j����51��!�EA�n�H�j��Ȣ�f�D���������Ԣv`���\�U�l�.dI�1�Ԗ����В�C��` ����:t�ퟩ��'���;Y<ݯQln(�6�%��E�֬mF�e�ո�d��2S+j��j#��#���%s�nRۖ^5'�ހ�����iS�x�y�R��S�ĥg�<ߧ���įC��A�S��TٽG̛G�-TF�,��N��QU�?i�&kwt#c���Lr���`j�v�G�r\��Mƶ��.��D��y@��X�Y�O�TH�.P6�ܽ����蹍<oђ��:Y`|�hn
�)�׃^ҟ3��ذ�B��ѐF�e�N���"$�����]*�ҥ*Ԥ�\��җ�Υ%-S~i�� �������L����'嘚4��J3E�HS׫���G�ǯ��U%>��ߪ���%ɧ������?���|i�F�!l��2�xF�f#��3�7N�N�;�{��Qb���c�Z��������Q��e4�Dbz���ip�&��������%���tIFGY�ȗ�E-b�2�Db�J���,$]��E
���E\S�
�Z�ޡ�&���d� ��8O#�t�5�&�1B�
S�y���ޭ3]yI����s����Д����Ӧ�����V��L�pL�(���i��w���"����<�>��׎�8�^�E���g@�q8�g�-�y�ɿo<ɬ% ��}�'�\�q��1P�W�T������9�#\�]�	�������^=���g�0k.6�n�jΧ�i6��4���U#��nM��u�ȫ�3w������؂�sf;�����wR��>)�/�]e|�[4�W�� A5��i�I���(��i�Y��}>�B���@�0�Lw�4H�������|).��ᙋ4B�鷴	�VS]�E��]손�=�������
!{}Kͱ�T��h�p'~�(�y@��&�E]���kǺnP�ӟ�2�g��=��S��Q�/���JC=��Q �sۗ##���<��
�)#�/S��  �o@��L7?�������Z� ��&�J����Ù�݇4*B'R|����3E�� �5�փ�IM�A�QƑ 6����s�o�m�|#)(qc���`ǩ�=zy�,���e�|�%���0ZW�u`�kxD@�x�ɼ���m�~�~d�����If!GimW$^���yj�yF%�xF�9�+CG��S0 �L�>����	]d��}Ę�>�QZ�^|��� ����� �➱�e�/M�X����[;�d.�* ��q��*��r,�vT���X�;���`���,��mr��4]�n�i��1f�H�^�8U8�v�y�oi	�}�,�^�r!O�s�l�u����%�ᴣ+�N���4D��G���1�yVy%�6��ajB�H��eZ�����,5�&ˡ�uX�9���}��u�$��)7�#�vҭ�!�@��k9e����~ߢE-`���a�l,�K�@�0���ȳl��@"���C?������E�/л�e =�J���\w6����V��C�Q�XT�y�����Z�� yI���)p��n���Ȍ�`WVnhB8��F�h�.�^�h|X|p����"����,�| .���j:��t��1l��<f���Yoz�W0_c#�-��uGW�:Ax��~����h��j��k�ͦJдy���\~�:��v�N̯3����Y� �RY;_��hK��wo�i�~X^����65��^`�M/ Ȓ�7�>d$�~v	�~#u*�LnL���^l*�/N/xڢDr���X� �9�k�n'}D�\n��b��L��;���Ǚ%��RǹD�>AÑ/Ľ�g�Gu��X|���VB,<��Zc6�����P@�03yLў�>yM�ϧn�8~"�*u]n1��G[��Ht�=�>����"�4|T>/��*:KWϷ��d�9h���P�f%q\�$U?5v��{f`�F��b�K52w!X���#�'ߩIp����%���niՉ��&�{��Ķ����o�!�2� ��2A��JFK��W�]��D8��,����4��$�U�
�Л3ZO���!I��.�W�ڣQm�Y��i�@����=���CM�%���Hn6�r} �R�βkH���	"`IJaL���z"G*P<")s�SBi��q��K��q��.<͐	I�
���7-�P=��aZU�˳�N'r-)a#��4��W���3������/ST,��?K�}m��1O��8 %��͇�����s��~/|�E��E0Sh��m�������`�"T�?a��Z�kڷ���I�
���A����˟Y6��`�R�ݬ�kN�OU��, �dy͟�9C?�6Z��	{SI���e��Yz/�����"ʎ��b��Ny �6־�V��|���7��� ɚum��*��9ᔮFzcW��)^?Γ��(����r�B6���F˺��a�f�Vz4q7�%�$��~?p�����6=���J!�,q#�����	غ��3�r>��؋��Z�cf��ו���!Wn�ݣ�	��q�`؉�ΫsN;�W�L�}���$r�������t�(�~mbR	S|��λ��/�hR��JvwCU����.����5B�i/B��'��@#�W]D1�R���B;^���c_^�`;�j�������*m�I`���k���%o��eN$�&����D��8���#q��w�����_mj����˟�A¸T$��h\3z���@�͇ו#�x9/�l2��mNƥM�{|�,O�v[���)�!�1CV(L��e����*��7?��_�4r>�s����Eb}9��#�k���A�������{��G��%~���uP����2���'M ��RV�'�{������o>q�lɈ�m�����#H���������&M�y��א�K���ivI����W��-\�3�a7V�8����A�@�L�'$,�_A�n�~�'�_��1�X��xE0�j��1�B��L��vB�#��.É�{������
-g����#��N1{)���8�l�{�p��q��@��$Z���J�&�q�5)�(SizB+��06�{�'��!�Ki�o@|���V|�Ax�Qu{;��=F|?i���b�d�ڐ�
�����S^
�L��B�*���?�*~�LN� �%�9��u����#l���w0A;U���WÓ��#����f���X��P�8��H�@b2�G��;yߧ��K������x�2���n��
T̐�6]�
� |�E�5_~�ͪO}Y�~c�nN��9�����qM;(��4��\Em8ϩW�+�n?��J��w�kŶ�+w���X�]4cF����B_gY��P�6��w�`#iQ&�2���?@��~/TR�5_[�D�o�[�x�֊���s*!S,e5a6�7��w�;T���r���Z��S)�~�x�� 5F0o��76!ׅsa������{���I��':�c����˯Y�8L��dm�N��Dژ�-R�N`�V��pw#�h`�sv�+�mE,r�ڛ�$��X7��{�\�P�
��8V������10�dL�va/FS�' <]�(�]�q_`��
`�j2�p�$Kt�Yf��C;�&
�l��L���5�S�"*{�O`r��n��S�5���	^�O�'�F�� �Z��:|�j�d|�h{bC����a��G`ŉ��Qџ�ޥʸ@g���v�6z&:�ԺM'OC�)�[���7*���XWz���&�5�Yc��$�Ս<��,�:��� 8.��'�È�Ya�aЀ1�B(5�a�+W�h��&�iT;{�N2���b��=҅�Ue'
���r����[p�_���������!��+����A��j�<[���A�"��QFp�	�[@�0�w1$�/P��R��f�	+�����~�dmY%��QnE��j� i�?��&ZUʏ{�t��Mk�ʎ��Y�+l4��������D�}�O$�I����E*��u��94���7Ÿ�|�T�t!'����~f�[�\8��"� Uq�2,]����-�S��O�W��16��[���`c��f^9Lk�t���N�t�=�� ���^ �Q�~�Pl�[�M����q�L&�+�kBgBxZ�N�>�������?g�-ҋM��:�o���QY�˚n�ϑ>h���[�Ҵ�w�?�;����{�%)88�D���|��"�ƯJ�eLP����i�4pB�5�����b<6h��7?oc�{̔жͤ_1�b^������+�^���p��U�J���1 l��{ȅ�n�P;�gQ���ɹ4���pc�A��Ry��:gV�oKG鸟LZ���Y� )�j-I�}�����������N�0Y�U"J��5N�(<���1���v��e\(UI�ф���Q|�"��Ԏ��Z�X6����cm������q8;�c�=]U�+�K����Ѫg~&��C-�kT@�4gd��X)v9�b�/�T�*��{g�%�C���{1�����+�ǁ�|�-���1z��q�ZɄ������'ǭ��B��ޤ�U2��-5�ٱK�,	-�'cm3V{��t���� ��QĔ&�g���U�G����%�j��K)���Df��Q:B�e ~՚~ܛdj�TWW�.��,F��+$��B���UX�h���������|�d3�ؽ���F"��D�?���X�ጔf��\I�U%�}�GL�	<o��K}�+��
�F%΢��֏<î���o�$����uiߨ*i���s������I6I�\�d�k"�ԓވpz6⻭rf�t�?�w�ƙ�L��� �	�mn���%���/)1����2�R��j�-��/j�r��r�2���#��˦�����$�������HQ� �y��XO����`%���/P��
��^��,��ϼy����2�²򿙻HN~}#�����a��&g��C�O�� ���>�G��U�Q'h��C\�M��zרs$Ϸ��ɑSA�_X�R��X�!o6I��(�*"}ݦaѶU�@~ :N���){�E֌�B��+k�v�����A������#��ԧ9f���
J��éE�!G�K���##�p�hTrBF����Q�3#��4�"�{3m�s!4�±��,�!{f��"�ل���-�@_�5�9q�^ l�X�x�*,o"��e[���E���e��(�+,!���A]f��<��"��)I�����֪G�2���(mv|�G�`��l��+ɀ)�C�8/�
�Lgrlz.T�Ny�R�����uc��> ڤ%Ӓ��̐9 �пt��������3RU<Kv���]ӣXI뢁Y��gJ$����w�hHd|~�}JD�d��I%�n�E�'�t;{xt�'��gN�2I�t�cr�^�@vG9M�}��7�`�q���UA,خxy��2�|�o� �B�ڵ��Iz]��P)�1W6��$����/��\��{f�3?���Y	�`J�AyȘz���F���r��/x`v�?t�2#p���ZkMef0	˱O�k�*1z�oE�ڇ�u�4Z�yf2-+�1W�q�z�^�i����:�+�F�/R!�WH�P�ԣ0��Η5���т��~	P/,���(B��pn��Яu�U�B�]2rͨ��L��En*�d$�ܰ9�mIO�j;z��s�A��z�-�3pj��v�B���Ϻy�N޻�p�l��KL�U<1�~Cp�C�O��-����MX[�cb�#���\ջ'�Ծ�gF5N/usf���~�%���������n7��#6Kb⨗������5�yVBpi�e�J�U$���Hi̊T�(��Q�j_C����>���P9't���eA0!�J!iJ<�H��f���֚7�5꿑�P�P%�%�jW�eG~l[�Y4�EN�6#LĐ!E��#���Բ�����1�͑��<��V�k0ʟ��2�⎗�lq˚�fnW ���j��4U���mQP$p������$�&�N��S�ڎ���K�K�޹�￢��P�p!W'���K��^��0ۼ��|9[�r�5�
i�a�*+}�ɏ����˺�0aMp3#�`m�ut��-����� ����O�^¥79�u�>)9��;��z�	`�S����	�(������ّ��O�B�&��D�Iۃ��	G	uU%�f�y��Y�����2�ԛ����ہ�.U(*�#.�k���r^ѫ��4�������R�)�KW|U�7��PC꼓SF%��Ȳc͙�J����nQei��V���b�O�c�@�!,ݓ����i�y�}꺰(H	�8�5iUy�h�i�����+���	lJzTo��6CG��4����(�

��$I�"��U���0�\ܮ��.ͭNd��zt�j�?H!�kA��m|4)+��z��9��J\\�rB"/�Q���W&�f�;�x�籴	P�����'���"����A��� �&1a���=F�)���Q��)Z�Sa���Z��L_Y�#�0p_����}6p)�#����s�vi��s�6_Vc6�&�B���:����I�]	�b��_����>w���f��l��M?c����l�n�On�vI�K�/̎h�%9@�.p�J�l�l��G�>�;L b��i p�,�+j�����FǾ�:�L�ڻ!�;�{�-��"�/Z�ڣV�VfQ¶���<��ÎV"�H�X��0���oN�C0Z2sJ�?��t /���H�5�_-�͕9��ф��:�Y�J���������	��<��3?���=E%���|$�& �E$F�����������6������1^5Yp:ԓ�FW�A�
Ip����p���]oG\�̂�ˎW�5��WＡ�G�ʏ �B�`a(	�P{d�
C��cA-�~t�-�JS�}�ľSa�N�fe<T8u(��<�u�Kh*6i�۞W��OV�F^���N�n����QK�%��]�K(�'-ӫ��?@��E���
+`;��>������d@�?�J�`}ۃ�ߜٕX���jC�t*Ǆ:39l�|���''ʊ�1��އ�,7CI~��lGzKLErz�у�E�'>!={�2���.Yd됦����QH�ԋn.���%�����k�����(7J ���Gk��%����P5��g�X��sR
߀@{}�,�'Ӆ�96q_o�5P��X}��'��q�7�RN]��j�n�tU�ֿ(�MC�Z��՞m9}^�T<����׿����}�=���v�U��Y���u!�U*b�Y}��j�����j��b�\�>7@�G�;��������Ho8��+�.��$a7�����_Nste�<}`�AH�f��Y�O}�	������v����	-�~��y�7�5�2�Y<x����NV¢#o�0�G���Z��=�?[���)������Di��VLyG��N3��J��K�S��N�%KZ��|�\y�<R!��-|��{��+�����B���,���ֆ��o��"��xR���'׽�B��h��+J�5�����v �*s�8H-�M�Y�N\c�/��I�&+y������os��)�uGOjX�5���Q?`�*ULD*��W��Q/�*��2�?��a����\'�Tf.���b�f��@��Y���)�h"L�pk"<�^.h�0�z#�vh�31LUB��jX�_ɼ��{Pzm�^��uL0h��"�C�]Ǎ|Q~�0?�8��!�  V Q�=<QG#[���[�T�8م�����<�r�EB���-e����5��St�5DL�TንAA�-�=��Y���ʎv_�����b��P��TƩ�f9ކ��Yh���0����J��]#]��` ��b֚ǩ��X�R"��� �����&�@b�]%~�]I�7��j�q�����w�!o(e��X�?7	�/�VF�i
�N�E
}V���;2��?�h#��%vj�'�}j���dIa���K�#3n�{+;�k0Qrʜ
`���ԇl�&��d������U,�����PՎF��dG	Egx�)v�}�
t@�e#�6�tP���'.sl"�6S��^��|�lM�:�t{���@E.�
^&�\��e���e��~)�S	�
z�eZ%��l������C?
��Ybz����2F�ZY�'*�2���,��T���zՀ�U�U��e��7���U���8�op^�,oF��٩
���ܘ��䕧�i��y�q�j�#�����Gy͉(+�K�����p�b�'��)�F�,�-��4���M��^��s�[���Dr���@<+PpH��_2�U� y.vo@�W�DǬ͋J$���p��bۺ�Fcr�B���0C[��݋�S)R��ȵ($h�7SY�jË����Įcb�ڟ�(=�ҺߠΈQqa��R}��􅴝�� ��z��=���m����b��?@S��.�U�uә�L[�\wt���S�Y �YFH���_��ɥ��PG��ض����+	���3��	�Pb2T�I�'6N��:���㖕�������x��o������':��� S{��-�(�nA�wO�nY'$hIĒ$��,J{��8-�Gf���Zoz��O�xg�N�~P?F����k*��Y�$	��eJ��?Kh�y�JUu�T�#SJ�N��L�)�L�t�	��NVw/ܐ��u��ͬU<W�ud���<�M8��$ u�|&]�gΒ����3���ZM�����-e���������+�η�<7�����L��%���I��O�/)��=�%mJ��|�}*������M��{�.�tGG�;>��>YS����EO��=#�g}����c�>��s���!��o:�]��n$��96�zY��a�O�!�O�R���p1�zS �~N¬�ϠÝ�T��tK���Jy:#*�<W��N�1h�݄:>d����`���W��@���¦�a\��@�G��z��S��<W���x}�p}O �I�-�ޢ�S3I�ў·y��B��×�.�p�Q���+3������:�(i�����v�1:Kӫ�� �x�j��<� ¢�-+p�࢞*��X�r����2l}|���q� ���R���¥�:�/����;*zQ�����bY�R1_�{��|�n��!iu4���^��9��*�Kd���S�4�
y}yM��~R5P��G���޵�:���ɲ8Oa-;N���V�0�ǯ�@�z�էK_k
t�`���y���迀jF۬�n��9`�HI� ��"ϸ�x���@���>a�ZS@�ԙڀ��Z3����Qi���6F���h�)�/��7�@9����Չ��G�Y? �b���,�����W�����8�$���Ɩ��v�7$p�^��c�0;�~
~�W9BA��`x�EM��Ϭ�B
lu;>z�X&s�.��a���:Snt�`��h��p*�R��q�\� �p�!������c��u��OK�s+�$j�2���|>���Er=o5�1/��~�LL�b�c��<_s&�͟��^��A��(\[1�������� �e�?�U�*<.�ʂU��X4�c�ض�*6�&[���G�כ,MZ@�	c�#�2�^�x�i&���P<$�2'P�G������[����7�k����3�C���O���t%6o�f̃���g%�diN�����\��=헨� �z�l����u��\7󂦨a[��@�U��j�C���y����;|b�A��P[���}���k�~��6��Oɦ
�
���
����(m.�K���$"ބ�������jƸo)?��y}�o��؊W�a����$H�j�t��m;�2(n����>�*;�(����Sk�{�ze)=��g(pauX >O0j>e�o_��v���G��v��T=��Ĭ25��/��u���Egn�U���\</�˴�`�)��A��'�n8<`4gM�[YU���n6�,�C��w��^��xk�IC�W����8��b����C��xL�����C��� m���j^�! w�x1YK�f���8�Qɀ��,d���'�Ś#��Q^r���� K�bL��DN����;F!qP�<�(�s �]ߦY��n�6{���+���=-<��<�~�� ]�mP�-��v"{���+ɓޔ;��6��~�O���2�~uק̟�zͽJH�:��e8~�CD��dC��(ʭ�{Ь	�,9Vs�ʗ�o^��N�!���*�ȵ��!���ћUm�I�#?q�*uB�|�T�)Ś>s�
������b��N�]�kW�ލ��*~ڊDm�Y�l��>:ö��J��w��3ۚ|_�o{�:Aٴ�8�q�){��������^�A�B�^�R�O"V븛�lQ��-Mc{�!�E� n��U�ɗ�R �d;Ŭ�e�.g��3��*@��h8VM��y"L� $P%L�5���Rio��f�]�Q0�k&�=��m�����"�)�O�Ka8����?ʥ����i.�5��.	d��w��R@��u�MT.8����w�`�8�w�^J�����#S{��qc����%Z=����j�|(�@]7S�7F��������Ybk��U���O�RS��k�Q����f*j��ԟ=�����@<�1��q�Jҫ��f�1?T�T!��cq߮3����Z��� }l����z�.�/�)#�m5IJ�C�ؤ�^�:��%ѣQ����]r����tA�9dc*Z��Q�l�('W�,"#H���u������xd;]M�yX
����˫Ps��l��vY%����"���ͤKcf;�E�r-�^����m*6�C�X�y9�*�m��\S�r;^q�fȭ�	(��b���$��7�V_'7�㮏��c�2+�߱q��g)��f@|��o��O+�����u=�U%P:����Dy�i� \d���RΖj��Ul28am|̒�+��`��fL����h���7��'���TZOw����rdZ7�� �j��(�5Y�l����%s�*���kq����Z+�񐂜/�z��I��^.�su��v��DX-�Ɔ=J>y3���yc�ˤ.��%�q>���ܖ���r��@���K�W�e"L.��.-�E�;]Mi�B�j�.�0zK���1�|���=&<���Y�¯�H�ߑm�b�vZ�Exj�j����[�WA��E殮��=/ש��[\���[���X�Y�����bC���]1b��&ug\�|U�^1��'�*B��n��o#l�+����U������F������z��\�+�`�����焁Հ��孮�u���y��N!��*f�t��0�X�032��oϱѠ!��~A\��$H��m��x$5͚��ȕ��B%<�B/��&�5������#|��5=?W%�&�8�J�]wBT�K�)%
F ��t>iO)��|&|�{Yo���{�ā����uf ��$�D�6�au�NN���d�g��/g^�z�k�_3�M��R�E"dc��z�NP�j��}��0)�-���]��P	݂�a��x�0/I��Ehe[��iy�׈@��x<�����8o�,쿀�����`�YW7<iV|�s��"��|2�w�,�� �1�4YG
g��n�K�Q_%
��������86+4��*lkC�2j9ɛK֙s����i��i�D��>�+���s+>al&��^�ދ����9��Z;����Z�H	���zp?
Hᕷ�^�7�Vla�hq�Y�|�z"vL��L恦Pr�
`F׌��h�AL=��;\4>�y���;N�H�Oˍ�>un�z���`�u`�2^��Z`���}� x�Mvh�_�
�q?������g��uGP:��p�t�NQ�#C��R� A���i���JS�����,��#�����g��x����/r�N�����Q' ��K7��U4��.�&���L�P	��9���X�ٽ��1�8��!�������=1�e���U�GL�ss��,�^��-1����.~뿣����]��v
Z��,���6:f
�+������ ��U�I��^i����yo�Q~���k ����0By$����I��������A�j-�Vh����i��q�j�/Cl��ۈ������XR"m�fT�M|�5��C��,��N��_����77�]�/�]]Ի �5�fӿ�#�L�2~�\zp�����)��ۑ�D/�5ݭ=���/ժ)��5��Ƕ����xu����HD]�j:r�.�G6�;:�U�}h��;W�#���	�5X�D���Q�=݇��p!�C��#��5���(�B��M���󷿇�%Z���J�Uay���EV��!�Fnkr�a���t�'@�Q���U��Q�W�뀑��{�!�d�.�� چ�pq�&��h_҇�Cv+]5@s\�������J)%����)���d)�֛N��h��Z��5q��'Tx�����.uD�Dv*� \l�����f�c�[���p�=�X��]�"qD������kT�@A�Lq��l�N(8y���j=T�$� Us�ɗ6K��r:�{���?�Kӡ��E���_"���}��q�u�B��x�[O�x��o�ie���UU�c��7���+䘩ٴ�^c�<���UP�����s�`�l�~�@��˫����|�%54(�{,�x�Q�0�X����tc��8}/]u��{��O�3�� ��#%�?:I��p�@T1������K���9{�c�
�D������3b��XRՌ�-�eA�K��!�`Hb�a�	��&Q��/�A(��)q�D�&9T�p��Z t�[;�����PE���+��ٍq�o�X�� �|�n�Q���$��
.��R�C�o��,�/o���K]qhFN(�	�~a���t�i~�<��^ 	Yn��zz<�n�n�G��I��$��/h88�(�0'�Ͽ�>SIw��Go<c_S��bz���&���V	D�S�?�^i�/�n�>yf�%�������M���(Mu��M�i.=3OQ���2JG����W&qrx�d�V8EJ3���Z:��9.�{���/ۈhf9����|�j����'�`~V3
�%�rf=tbus	u��xU;]��5yeC# �<X�����T�;ׇ�RZ�|�>%��Ƶ
�]`�#�"[$�p���m���b��Mf������Y�����)$��=�Tp3�C�.K��h]]z���gԇA��ZZ�m�z�8 �[�|�J5�n<�J�����G��`~4.��Y�A0wٖ�� ̷꼯��UB��/^o�mI2@�&�>�f��;8L0v�q$o� ���n�dl�#L+�4�*�J�-��L?S�JG�p x���K���0
�����M`.�}�-����x['�y�G����.m|ƶ���y��/�]cV]/�/�n���95��y3��x���l$��`��_4� ���'�Lo�/�s�Y�5%A�M �' �_)�d1.��]��6�Ĭ�#�)�?�uO�AZEd:��R�T�G�6�H�|c��mNqaw 3f2~�og�˸de��XBږ�eh3��YQz@��1v���V�"M�9K�<�}��6c�#����tȱ	�k������%����2<�)�*�&"��o�A"T�L���H(]���z	��a�h�g*�H=5��_
?�#=�FwB ����yM1<
A���p¢��o���P�nt�0�B�UF��UA�)V�z���ĥ
||F�C!�D�o��o��o3��3ſ�]n���ȼVW�PUH�q]����f����"���(_m��x;Nf���bL*D�enGnvT<�|��%���X:
J�y}� ���䑮E6����+�%e�ac=8Β�z�<�ڄ&�<�Fu�� �=�ix7M�7�H ޸\�s��q������V.FG�Y��x���<o͔z篥�5�b*E%N�Wx�M�q+�W���=:�^}�Hqy����̂��'������(��2_q�C�Eğ9�I>��F��fy������z�rS2Q���t��6O"bg�$"۵�#Y�@6�Xx���_D����5jƐ�V����ո͡��D�s2��c�ܨ�\�A��X��3z�>W��~�1��|>|�L;)L�]b���������>Q��|w���}d>'$N���׎}BHXz^P��O���֒	V/3����Vl�5|c���Kn -�j��7�)vc���J��\�_C��p�b�?P1K��ǅ�g�4w���qa�f��H@`W��=�u�s��+��6t�^+A��Uv��k�![3��`�W�����F�gr�
v���U�ǫs�ܺ��Y>�mn�Qt��9�;����`��c���LDL���%E����p̟t�4`�k¡��L!�_���"�2�}�y)]�.�<�.�{�'��9���Č����^�#��Z���J6�uʷn�|A���
Ѐ���qV����Tyb�_-�J���kc���
{�jTz3 c&7��L��Q>	Ƨ���P������|_V�D)�આ1�F�+c�̫e����WD��,��0��&�#����iЇ�K���@���G�JL�%0V�HE�)uUz>m:�#��"
Ր:s��}��Nm+�m%���
�q�)�C(�\�g���~6�A�<���..
��K��<�;`g���,���c�xZR޾�g_�+	 �#����/5 �x�}���� ��}5^n�+�T�j
�L����o��X����T*�f����` �"�7�?yKNˆ�@P���4O��0���虘����s�i�����^���	�\�
x�MG"D|��2���2�EP�M������@`��⬸K�l����h���|S�-h�m���|;���.�H����o�J�ˎ+k�ڜ�ӎ��ntMq�C�6qU�����_`P
"'�/ݚ]�-�gC�s4=sQn<P�d�� ��⣙p�'�3�~��N�iiꭋ�$lw��z�p�`x�߭��J��)ue��eV����� \��p+��Cn�"lx��� %�jP�Bp�� ��|��[�sN�܅���֫��*�z�ۙ"�g�ܲ���R�q�y�X��#E�b&Tޔ�md�)����/�����$�߫�#�Jz�>fq	�c���1�9��A�*cv�C��[��=��9�f}6�"��B�ȩڒ��Iu6 �d0���:$$,(�44C����g����=a�5=�BY#!k��.�HzOEX��V�H����iFO^ Pb�V�J��S����}4�v���>��`>��U�&N ��`�o��������N�d��E�\ѫ���0����)%�:��������}��!��F�z�w���~� [a�/(�:M'c��MF���H�.Z9��Zp�Ĭ��+6����d�Q�� �ۜ�v~?��0�£y�qA!6������C���"�G�$����>�T91Q|M��J�ӥR!�,�oý)����-&Դ�����X�	p��A�yܓ�p��~b�w¹�,����$8^�8!����3�K�JP�VA�s�/�
bn%�|(��:��Ѣ�ՙx��%��[2��u\�o�]�G��0�+��[%�Zhh���4mA:�/<���z���9���*��{�����Q#�鞴h�0k�"f_��x��Yni�p�B�2�J?�$�4�0��+ ���Q$D�I@X1=Y�QR08q�V� ��3�+C��Lϳ[��a$?�"�reW� DNGG{	��0�Zac�C��ee3�\z�B�����/]+KF`�G�d��sօ[P�0��w�(;�-f��i���Rͳ\;�0:��hOW<�NmC̼yF�hjS|�����&\0�1c3ϟ���y��/�[�8�ܺax�����Ls&s�J���d���������������&?���<�ΚF����D������Q9�Ql�~?5[��4�n�_�Gѱ)ay�m�P3��թ����JɊL���;�����y�X���׊2�'�;%���������}@�!�,�yЕy��N(�g��E)��-�g��!m�4Qx�lB�g��n���m9����˭��*1�{A0����}�8K�s&nx{<��7�����c���fǼ��+�X����,�����bOe�Z�Tmr����p��3.@^�d��4�,�G�wM���H�Dv�k�S�Rˌ��}�'C�d���Y�I���Ǻx�w�p��&+4���?�5:ҽp{��`cUSO`��nAw��=�Q6�ɖ��d��Y�JNH�Ӿ�U���`P��7��D�1�Y��l�r�\�j���S��h���jp�sJ�+f �	&H�蹞�.!0��fw��sP�V�;?g�7Ɩ���e)j�Ǘ�$ �v�_�)��Gl�N�F���^m���K�MC����������ט�MF���h4���X���r�w�#��U� b���ِe�����3҃�U�/�9A�Fp�M&Z{�FV0D���R��W���~3;L�j_܊|������g�I�H�RL8�#/1l=_�{��͟m0�M|��5��1�8�PP>��ΆV�+����8O~�2(��~���uM�����_)Lj���kjp���~,Cx�C�|��`��U�OZ�%��V�-'�[�Qv ���~������'�OJo�����$��f��о�H���|j�{���V�'h_�c�h�$H���>u�b�N�z� �ӟ�y�\V�{/򼫓u��(�{N�L��n{�۹�gjr
�x]Pk��JN��h�� :;R�ɇ-n16��
j�R�"Mzt�ثe���M�!��&�lzn�_N�1�܂�ܼ�U�?do�y�Q?I�O�߃n�a��"^Zۆ_ �����]�+��Ҁș[1c��7. �SY���q���*2��4�c-�h�B0��I���r<2y��񕲶�� BI��I�܄�e=�A�?���N�M����(, ���Ƴ4�e�"9o���uwT{.�%UEv�&��1�
k��[9	�DB��i1�M�R᪂�>`y�ɡX�� H���CJ�	��up���PΟ���">tV	A��}D�i+�0c��L̍3 ����3N�T�k��?����qA�m��8l��O�t��_v���ӪW����cߌ�o�u������A^��F	h��/P=x�-�9Z�|��K;W�ݯ�-5�q#�Q�!}_h��.IQ�(��c��iw��w�-6敼ET�8 �������y�Ҵ�h��L�v^��|z_����O�޸rkE�����#��ԵH_��g|���cx��䲀�׉��)���m4��~o4���5M�dPw��w�.�aO:��i��=<l��2zk����Ӟj�5�+8-�:+Zp�����:4c���z���TVE룦�<�Z4H��Wж�$�'�L͆OP�+�p^و�I�!H}�7+k�'@Ɗ]��̄���u�h,��GÚ�L��5<$���ؙ�]T�ن�Wtٔ�:b,J�;����/z���^Z��jfC�>�eP���~��W��2��C�����*H?��4�"+
��^�}&?�"�\���UPE�h���F�'a�>b�[/+�5 �5�D���4�����+s������0D�� ����ϸ��F3Q������g��hZ������v�^��i315�SN6n���4_i� �����
���|9�����F�hT/%��ݫK��ws�n�@��D�}�3�)�+�Z���Җ�����1}X���q̰z	k�ё� r�&O�*
nU3W �=�(>�T�6x�SF ���� ����X�fk�gƻ���C��`�׏Z�NW�\GZ�8��&	:�z�+��y�7����~�p4�����|��^�X�#�D$ȴ1�Xp����> G��Iڲ��y�� �MVlcD�8r��:��R|�����*(�ݎ�W���M�����E�����8�)4]�D{�X�$R μ�M��	�iK�7��RAA\�T�t�PD�T����-����Ե#����j_�j:V�Ab��ٓ���U��B-#Ѥ�IU%�2��{����k��i#Xf�A�yh����� O���R1�����a8�S���>��rk\��U���g�;�W�GOc��P���=����
H�x�F��}�$yZi+-{��w?�IP}�Ρ.��`��̌��;���D��S��|萤����m/�t�O�!(p1���zT1��6(���s�5�[xŕ�����WB�}V�G3SY>QY.���}ҙ.I���cXڷ��i���mhi.��i󧩹�9C�ݥ`W��ٱ#ǲ�S�>Jqv�����Ya�A�pՏ�/�I=�D
~�e]�o
�����>5���BN�E�B^n���#C�V$�O�Ƒ�8b���q#�� pk������;\S"��Ӛ�G�Y�.5�j��}��{�3*oD.��쒓�������V('�µ�}�?5])c���gD��TP����B��!X�&�D�8l�:Ǳz�Q��/-B�����睞p�
Ҁ�c�ݔ�k�2-�T�X�@�8o*6@G����_��%�zA}�f9#W�/;����±�������(��=)��"}X�f.l����lf�mE2�W����C=�`��@�I��|c Vzĩ����d���U}ý$�oB�E:�Ѷ���� s%��?Z�6L��ŅB|�QY�ښµg͍�e��1�qUՙ��l�d�.xJ�J����Ȱ-=��# ̍��BS�On�_�B_t[�
6�\6���l)��:�/���b_�9�NyG��?�ǢkI&�+@� �Z��w��F�+ͷ�\�zՎ^F���6����=��^A�C+stTw�=��t���/�`��=;#�����>�팱i��Y���A2X��(����sG�󄬗��b�Z��v�%n�M�Lj��t1�m%��	5��dIdRU���i!-�?�8����iX�s��2OZ{rs�qE|6�!n�sa���'�����\�K��ζ��6��H��ݵ�їg�ejq��������׊������L2� y�6A�Xoi�`H�.*m�Q:�P�6'+(�7�ɖi�X�zg�e���Z;�dQtC�qb4��I�%冘b�u��ɓ����u$D�'4�t��~�I��Tʾ�T�k�T߅��ܴ̭ut_�J�1GD[��)gg��U\q�	� ��RG��Z1�@r�f ��G��ʀ-RA!'�:���2i��dBUQ�r8�@�A�����è)��d��}���]-�F��h�.hA�J��4�i��e+$�i�)���a�jf*0�L�'�_�b-p���!eO��kf�k{^�)
�:���I���N�%�PpD�D`�'���q���.<���lʨ����Ř�h$����Ζ����y����ީs���l0)o�l��F�#������ ,���)���_��d�y��JA��fp3QD�Ч6�RsQ����D�a�^x��Ud��j_P���eق���߃�Z��t��Y�K���ύA�J��% ���ע�\,������z`!�A�V	f���$�u���  ���9a��P%}x�!�W7�hN�&m�R�P�Z�6�Ph��7����a՛,���)�_�;�@xDȘ$�u�aO΢Q�#"
�����B��
d�ʮ��3 �x�m0~Q�������;��=.�'y>�9K�y�٤H�Z-�{W�O�����[&�i��ב������J[���ڕ5���Zj����ld4��e{^�ol��_�9�K>��3X�r%{r��0�s%��@�$��'���&�|�p+q��U�9��d.e��*t
/N=���f�[�g��]��*MQ�Dk[g�8���(������h<�@UPWK�����<�q��T[= ��n3�-Ts4��H�H���9 ��u�a��Թ��� 73���q'�w��ޏ�1M|�OiK�h/1����� ���?7
 ��^�m�h�N�ÉYX_SDE�hw�b����9�H���� �S=�L��Z�\oi��v��LB�Ք��t�R�jk��?����'[�����+��(Nz�?�ɐ�HB�I��2b���Q��m/���,�] e�ޅ��Η���$C��_1��� �k������Er��=�ǵ�\�)�"�����ϲ �,�u�i0KG���� e�Ӝ5֭���.42��� ����7�'͋�T��B�{Q}#�)?{
�e+t��������ӗ�ӣ��k���5.��H�9�x�3��S���h2l > �x&�.p�qt3�BS{�p�K���THQ�������W��A�l��Գ�����I��8��%��m�9����]�
�4�p�ґP8]���^s����+D��SKLw��Ǧ�����ӝ�6_w"���o�E�mu/C^$O��{�Z�����5~���L�Wf4n�{K��p�}k�JZm�I��Y��d��x���6�P�}�MY:���6!l`��f#�fOx;��Z̕��H|��{5��ܸ錏�����$&;G�a�KV�a�D��Kl�%c�s����.�ٛ���l�r�{�H}*�i~�Qs{���� ��{���mQ{�~������w��-?wn[�"������ޯ��?N�t앺��?���b|�:�#���j�~�?S��b����gs���Y�r�t��(�mH��F\|��Z�x�Ͱ"}���ǨQ�-��Ȝ%�Lo����d����o��`�!��rTh`��'�
�C1�����k*�0ޣE�'O+wn籵FA��Z
i�E�֚T)(.9��$p�Ã�j�}@"s���e/����X¨<ۡ����u�Ex�Q��Ƒ��$qfe'�*�9^ܬ%ظ���fo�G'�[a̝��W�s!(ͯ�gr���]�\0=�T���U����f� \� 0�ŵeH���v5�yT���M|�=jlKХ<�n����R��ϱ4>d�tSBj]H7>�0EB��i�VJ;�D���j7F�E?�.�l>����(d�wz��Xao��^�|�M�+�&`��@��n���S��v'Fn��US�������� ��q�at��;����&-�9܆KOƯB�Je�L����/9��%�O@ls"Ck<<}�{���"��_�2ik�]qĂ��0ʂ�QGb�i{����
���L�Moߘ��x�[gw���iX+=+��!8�Dl�:��F�,ԁ��X8.W��9�emg�-O P:�(�����9BX3
כ�a�����K�v+௵Q�䓨�jE����CǊ�F
���I�A6��W杯�|cMT�%y���v"/Z�q�2��x���}W*zX���V@�U�2�����TFth����������o�ե���>���4Z|����Vb�э=���blY-*7�?K�����R��z<���$<9���X���o������W��=��3�9��������Y1y.�\=ݔ�4ڱf�6�c1����)>�z�saS����N�����i*��Oa.�u.��0�,鹦�Z�#��9(��d'�m��D�<5$w�17Inq��S�T����_�K"�.Z��W L�L��_���錂����rez��>%[IN��҆N:�M%ӫ9�iMҙ�ds�D��JDOs�g8�Z;&B��~��I@x����; jП]�E�fI�P.2٘E��C��0pH�|��r��ۣVw?u��<Z^��3-�%ap�#�kv������ҍ:�H���pN����������$rÄ́%���~,�Vw˫N�I�����T�A�J�m�OH�˚W���$�d����U>��4�G
�G�}U�Qɐ:Я@���Ś��>)X���7���҇���c��?���{I���Дr�r���u�Q��xSxUq�dO��2c��l�qx��:��«�>�~w)
&��t2�,�(�G����VmedЕZ��T� �[��!�bQ��W� ?:����}P�m���	Y�}v=������ΉJ�c�/�*�����=�c}E�o���p.��@r�d�?��F�x+I���#6��b>����	*�"_����AM��7	X+�\�̞�^e���<}�����{�M]^%9U� �*����N���l:��?�W�����6k$�[*6�v�N�ds&%y&f��Fb�>&"s�N���{haܟCa�dB�ʯ��٘c�xK�[�mdcۺ�7k�m����M������ES�W�RX�(�`֜\�� S�Ճ������H�
�h�|���[���n��X���/�$�1�IP�A�`{ϐʶLpcQ��ױ��h�E�BFj&�D��u��U�UM�PE���?����䠂�@&@�e��!�b�d��'�
T�:�r>�cސm��y�n��w�ހ����}1f95��~@d��%0J6%�Z߆���@|
b��Yi޵�K���<.��k|��4��9�ogo-r�|�p����;SS�1m���Kh�y4s����]e��.���ț7��f�{|�J�7c�� ��<̂���aYHe$dSN��S�%ƛxK��۵��
l'�8�h��V;[����8MXԋ*��#�8v��Q>}��#Ҙl	+�x�� c�T� b_<�
.y�R�g/�(��Y�d�!$��	
,��hy�r�������Z���\�G{&� ���#�h�n�ň����5/��KǬ��3G/��Y�<�=�3冱�,&���n�'�a�3�E�JW��������ߠ7�wb�po�o[~��fKi��!�f�yF�9�$�?vkZ4T/u�R�l�2���x�����p��?8�*(��Cf$���i'��G^|irf�F���6���R���"��k�-�;�8��e��/V"e},�x%��T'��!+���}��&3r�R���p{�{�k���Nf��_w��L�/d������nl���Jy���=]6t9ϙV/��ki�;o]�+af�ʍ��~�x6>_/Ϝ��� .��^�"K��ʏ�3�?��xz�T9[�h�w� ����>���(�	�*�m����W��eI����،�`�i�'Q�Gu܋�)����1^����+��.zp�?�J�Kd��n�^栆�������b�Q� ���(@��$���<^����r��pR����݉JVc���4�a��T�z�B5�\�0�"���'L�:]Q�/��[m��ۋ_��h�$L�`ߗ��1�lI^N�P�ض�2E�����%�`=y�u���n_P/���{�)��z8�S~ �UJW�Yp���O�F*�9���ش^��V�;*B�}ᓍ �Ռ���ڼ�(�C��	�E���Ѩ&���V3ڙr�,�7�R���1l��͊�o��7.��)R3�8���_m����X�>��U{=@�;_㫥'3��Ƚ%�%Έ�Y@�xݽ� �� �����'^�i�)E� B�k��U)6�����:U�8)��$V��9�E����G"����U�Ơ�ϦAV�����j/Dho\AY=���ƀ� Y��97�2�$uA�)ɸe��-PJ��?�C4;�N�# ��L.�q[;�~<�����К*?�=3�tŵ�����p_/���g�;=bY�1܎Y�װ�Q5�˷�3�\ē��v�㏺������c8��'(��bQFjcP��� +U���;��#���sh�~W�>
�.�ʅ(-��H�%�:���^T?�k�k����z�R�i��3�OpВ��y��N������ ��C�9�~x�ܭ}�B�?��A��'��n7[d�^܎��ag14��J䲿}�o�5n@r��ު�,g�.��� ���\�g��ԍA�W���7.�����7)f�%�E%��0�b����]������VD&�$�ƚ�j����PG����tj����^J������Jjy%��Vvhi��U���S��w��j��WՈt�g���<�����b��@Aj�I��M�xr�­'�R� �;�8f|~e$�O���T�	6�SS�*e]a��`(�M0<��?܅��D�`}nVzϰ�+��[��	��ݮ�'���%��r��U�[Lk�꼇p�j�\sk�y#���T�p2-:eS!w�bxP��ak<=�ccj��^f}�<Q�'E	v�{Z�.�~�u��O��U�Ǝ�V}XDl)��#AR�?6��^P��6���N��l;w n�\ؘ:�����mN��fZ���U�p�8鴟N`��a�*��p?d)T��ގ�:�YC�=+�JpQTA���.�P e t��q�B|��yc��׃njtUHp��x���U�ܠ�U����hy{��m�^�V�H��?��x��{��+���]��I$�M)p��|*Bu�]j����ud��g\w��ܤ��AHDU��r)�vm�`��C_�4��$����B��x���-���/\2����l;�ȘڿqG���׼������]�կN�m/*������7{ �Ԇ�U(�]d�ax��L�a��3M�����&�X4Af���u��#�tl𚞻��G���b��咢��V[��JEp=)�$UJ��d:��ߒ�*�>�k[Ͱ�)7>��gS
�h�z2��������3iŠ��"�f�+<R�Ja���F]��i����1���ֿEp�	�sϸ� �/$��F�Ѻ�i�cfa�}��8�?d���/`C�!(�����D�tԙ`s:�,�	 0��1���_ʹ�,���;W��	���38DF&,-\n��JH'>Y�O��[������ܴG�H{1����|�w���=��4���wsA@������u��8
l:[!@|����,�!$[�E�wj��@{��N�$�,*d��s��J����/==<�O���Y \~H�FI�ą�b(Х���N,V�Ϗ�ņoi�$�4�����lڨ[Ň���q�x�d ����E�\��m�SV�3AJ����L'�.��k�3j�<1��"��s�B�������s������g���0���=������e��{I�&B�5�6���dy�xr6����R^8s�B�lDd�y�pbC���Š���fxj��,����M�V��0KO�+* &�}	:ͯ�xS��V:}���@�F;�������C?���V��"-bqy�&B���?Q�=MZ��]�ȝ�k��Y�t��V���{�Y庪�CW���(���jV9��ȩ�=�C�U�tCj!m�"}����x>�=��%��~���X�߸���&�}?P�Wo�y�j��6��l�~�B�-8���'jk�6�5�v�6�h�a�z:).Xפ.!j����y�"��5�L-����mj������p?�+��#�����I�������}��e�za���-�s��{�!U���Ɇ'�6�x��sc��&�pB��u5��jf���u��w�5���`�c�Ny��?{�p�Z���;�D�6ǜ+G#5���ո�&ɂ|^��	��\	����;U��5r�?��G���x��,��rK��cY��~�R��;9����u�h��2*c�^��c�����{��J�CS�fEκ�k�]��^�r�Ş�e���\bF��?���]!Sz������4iV:�Ht&����Tm��=��&_�߉�W��o׽e�k�},kM1G�7R�	�*,�3��~w����,SI�Z��a�y�Su}�67���Yd�Ј�(P�OMc��0�%]��T�ַ����<���}�I57"fmb(����z6��c���	�h��ZK/�I�}x4���(8��:߬^�;Q}p��p]pQ�@6I�����6鶻ݓQ�wT8%漗�iV�C����t�)���8���ᇼ�E\NX���!,T���^ū���	|x�<���&�8A���ͱ�	��#礏�"�TjYZK�T���N�6�;��H4��C��n�8�.&��G	���B8&������S",Rs�p��
,`_J����[����� �����rЁ��~TA,��I!q��?��i�4.j�\(� ��  u��~���28":@	�k,JùM1��YQڄJ�yl63�l��Ts/^�=����QK��#��p�)�4�r�+�ܦC�PRMj��V�s*� t�
]im�N��j�	�f��[��C#]�4q��
��h3рvi6)�G����+'�]��.���S�{�<��Z�u�~���K	g���|� ��.
m�ţuj��d�_���ZVԸ��T(TV�3ď|�B�@���M2�X��j�"ӥ�&���Sv�YFd �m(�o힣?M�=��c���6�Jp@��ϛR�q3⭅�o*�;I� �kSPO��r���X<g���/Ǐ�}S�����%�@Jq��(�P:2�sw�[ߘ/�)=z���nb�q	d,�����]4��x����9��e��Ҟ��u*b���k�@鹍K�E��O5j�p����ln����Ӑ�3M��_�p��������|ǻ �ّ��A��
�T{�V{(�!ne��
XDF��Q��|/F����G=��P~���D���u�{��u�`6�Z�*�xq�����[�[Y+p�i_`O��ehzG+���VWJg��p���ͩ��.R$o���m��f(�{�ζ�)��1j���Vh���D�v� ����,�K�V�ر%�J�ҏ��W�ߙ2>N�zN1��NE�B�}j���yt�b?�6��X̢Qa��p`�3�'��MِI"pJE]�c�zΫiD"��c��1���EF�����
�<��a^#Z6���d���ب����ػ��BK��/���ި��xy�S���4�q�O��^�:2y*S�nY�R�����"i�M�1���߷"$!�a�_�	��B0�738f��ɹ���*O��@;ٖ-��\��|�LM�6?",]ļ]��~O}lJBl��E̊�@[��ԡ�:�b�}���Ȫi�㦀��z�F`)��ﬗ؟��~	��}�� ��b��2K�2���8d;���:m;8�w�ϕr,.��
��I&�4|2�<�U_�Ҷ����S���8i�{zQ��q��zg�ߪ��SY�O5��j�D����������u�-��,AJ��X�����m~b
?i 6��'���A�>���]i�\�;P!Y������hS���>����z,q�9y8����j�mu<���/n Ar�5Nc���������� [\�$@�e��Dt��7�)1�����V�2^Pc�;��TS�ؕ��y�� �7EYt &d�Y@��n�N?t_�OW��h�3+�k"�;�G����W����q������p�A�4b������~�  �T�!P�C%�@�@�3��pO�r�?7��?���kMI�iNډ��xA=+s�������w�R�����Z�JyZi���@�OB�o�,�m�����:�q������ާ�(�6����s/�]�/ڍH$0�����Z�{�:�=�����E�s 7K�<�2Dd����J���]�P^��<�ȋ,��+���p����ƫ���$mkϠg�
4�M�Y���E5���I
���_
9o#�Z%�C��D�tx��.xz��t6������\��.:YU�B
Z�Nk�>�o����	�b��ro�);�3�ÂL��?�r�yT!�VW�	�R(�nG�Yqf'v��]��$�+]��V��� �\J<����S'��y6Rއ��Ô�&�� OID5�(��t=U�������Dy�$�,$*����*8"�d�_�\��q�;n�$�y[WJݧ|��=�LE=	��mV{�S����4�W�j��X��p�ބzP���r�*�w�7��M��w����(?J.b���:���=�ӊݵ���yF����U��^���L��*�1̍������p��6z#�5�lk��o���/�ʀS�k�7wŵ���mO�IGiڡG*�( �� Y�uJr�_1/3_"(e��#�JlͲ�V��<F��;�'/ï-�:sH;��f���,�@ۄ�?e���#ša+1k��xM':3� 0s��:���.y �x��+8v���K�YuY�Qxg�*9���6)�RW(Z�T�e�hf������U���Ɠ�T�ԇ:g���,�'�_�ć��ܦ����ƔI���9K"��.��X�J�|=l�OU�R�*��#k�k�>�vE5o�6�OF����ȳ�؇�Ƽ���uA%J0?�v���[fKxð��r��QPz�*�J;w��zϜڌ�2��q���A���N&0�� s��������c���i��K�'MP�ܰ\:� 11HX��y�4��~-b��M��F�!����.�<\�=��
�S��!\�~�B�GF��#|),w���c�Fِ?��W��5E�3����7����4�i�)����$�_!������dy��Q���F���W}Vt5Z1<.W6YΫ�.���3�QE�
�xx$��xb58T�W46-��c�B�1�f� ]�'�V8)qa��wi60X���t���p��]�ȄrzԘ��p�?IN�K}��q�y�d� �?^�~^��3���pZp2���7E�(�;���h��)���]:��>S�j��x 8X#έ:��;cێ���+m��{�\�� ^�[��?�fE�/��c���UzV_���6B-�V�bv��w�W�[��":>`KǀJ�mN�l>��\�#ݳo�ş��<��H�v�x����)&�BXQ��Kև~Cx�	����۶�����ģ�-Z~�'��3���v����@��]�󷇺����{��ݽd�6o�]%ӣ�Gy���_���*m�����;��'<%_�t�j�������,v{�8n44%�N�{�%&����4�W�6s6`�ED��F�������E�_޼��c��aԉK 4M���N���خP2�ힾ�i.�7�RpQJ�xpn)B��� ��{��*>�������Ce[�$c��Qδ�Df�!���P�l������)�PšDem(@�V�_�"v�Q�N� uR���=W���,b�սM����Mۧ�q�eI�
*��%	�:A�����R�r:���>�ߔ;x��T��Ĺ��g^�DzpàJ��W�!�/�b�ݣv	�<�D_x�s�F�W%��  R�>f�6��̂�M/Q��sV���P�.?;��r<{��|�.��Vs������*��cV��M�[j�V��x�>gx�(���K�^�aM���MPU����w/��s�߷9����iNd}31j��.�D��#A� �,U����i�wGS�|F��M�_�2K�s����K' o�H3��P9�B���6������ö����㹌r��K�r#3��e�g��s����܋�+�4˹'M�"�(��U+f�o�T�3;~В�N��<!�V��,���Z����lH@	���o�%�^>Z���[�,,����9�@�E���q�3�➮�s5"a��ޱ�&���f��7�ߏnP|���a�k/v[�QLIl�scF�l%���ɣ!Hi�5�G��JQ�9H���ЌX�ƈL����3�[�q��A�/��6��e���A�>��AĺZ�����lYv����Dk�T���_3�����P*v�|��cC:%��]��߶i�����bp1�<v�Z\#.���IV����LNi��f�;<Bl���H㳹��K������C<X�Wo���g®�h=]�Jr}ܩm�A�8Z�f�[�U���~�Ur�LҒ��9��`�f{��`��!z�X��k4����bD��G�f����@#v�v��_ڣC=XN.J�x #]�{�^�a�W������b�+��;4��=NeA�)���:r������>a"��x1"���TNH�3��,�#^#d��d,Uxp=	Ab����Tn��]�*�%�����	�
�O4�5���S5���y��;eq�,��T�E��#Yo�4�򍨷����$��S��M�\��s�(Io�d�֫��{�^hg޲~����b�z��RDp�[I�ƪ�_k+��1<C�c�|BC��Ќr���\�T���	�����@��0�~��*���5vڨ>��;e����=������P{���!�����qM��~�$?��i��G��)��'k�G|�is3��h�o��ts���T��j��a�4�T��w�,������6��X!b*t9��Exa��'+7������(�ײ%^��tψTH!��]`	��}0NBȲ�B�G?<��8N���#�(o�V�ViƜ(�8��Ŵ
s{\t�Fb��%3Jq?������e��ڤ�ErF��7hW�i�:�X�t�0-v0�g���s6�暜14I� <���ܸ2N.1�<lh��㟡J�d����0�jrDUƹ���~�%,x��f�X ��3��+��}�g�l��Y>&c[���,d�����{�����Ιk�d�9��OS8���7���HyL?<-tM⍛-���>zV�D<��7�S������?�J?>�E�P�f����s[ ��ch�,����v8)׌jC1)xL��:O�
����6F�����D�����[�IO)��V%��.|r��|����Dַ Ӆ�Xz}��l�g��}D��k�ݘ��jN�P��Q��3f4��̤�%��f���H�����	���� �Y��/��N{�:��hؔ��K� �<�`����#ip��o
� G�d���W���u	� �¦�Іϛ��"Z�)�cs�X*� `�E����4�Ba�&K�5�s.�Ou"�Y�u6q��ǆ�|��Fn]����@w�|j��J�T6y�sH�`�����T�y�u@�Ze�Ӯ���9�@�C8�c��mzd����Q&
;���,5^}��nPq�-��wISg����~���j��ռS!�9�5�U/��9��D�7!X�z�e�y>'��'��6�����Ex�l%M�'���n1�n�+�CZH���LD���Gm���!M:p������/7��F����W0d��Ѫi���sp���Ͱ`�E����m۴�9ה�Z�؏��g���Ə�!�����&�ߴ�Z)���i�J�����Y�L��I�3�4'�(���<�G�u_��
�|]�t��X��>������v�~�7�ub�N]�G$&:]^C��m�=C�-v�ߪ�� $�̷N��Fͥ��K�|�Tw�P��k����_�N���~��}���fM*��`Q*�}��I3d!��ڷp����(�.kk�X���Y8#A����T	������lï͟��У.�h�%:*V|d
|M:;3��n�PA�"	�8���������f�Z��ލ��Eÿ���t�<�(Kɟo��w6���֯�f�6Ĵԩ\��W���=��ÂԤVpM�(�+n���}r|	��s��A߷b�(��G ���	��� �3�\O)��-���癬������7���\D%��K�^I�oﰐ���fpI�)�FKc��+Ӈ��h*RL�v��N�
V�c��W20,�'ܧV*�������֡ r������)�A2���t�3��uc#��;�ڠ-6����y�x8���6.V�.�s��DODr��ڡ�z�B�|��@�*J0����_�1T:���_[�a����Z����8Z9�x<{��:x�4E��P�`Q�`\��ʘ��|-E���.��J��K#	��j�Όٌŉ~�54w�4���TG�B���5��.�ɉ��g���+פ�������T�b&/��M�~gc��,��N���aV�|f�a����#-lN��~��~:@�ߢ���j�1�$]�z���(r8�(	�i�.2U�7�D�;V鐗���U)o�6�d�~5��r���DX5����*���l��%�שd B��9}Bd��H�F��I$`�;9�pD�jzX�iD;Y�a;$1���m���RP*c$+L��D�x����kķ�oS��G/��%S5��*����t�=�ic����'HDH�B	5��`ye6K�vjO
=J�ߎ���<�3t3���*Ct1.�"4KA����������2W*N�*���V AEQ=S�%k}<�VAJ���,�zW������l���ܕ >[*O\�A�>��@�\�9���E�;j��x�מ<��ۑ �q' s�@�D[ݭ^�N/��
BX�� fvî+�0S�0�v�
Qg�Z�P��٧i��Cۋ�'��'��}��$��ҙ녙�-��k����%Fc�*c�&����^IC�F�4Z<�[�B��A��oV���&hAV'cȡV�h1.��[�99J#�r��R�=(A��>c�U��t�%D�b�uH��$x�Rz���0	QٰZ��3Wq�۱|
΅�*/�#�u{l�g��}�2ˎ��	���bL��M�#t�M�g5���E�5,�݌�Sf��ے��JJIjLWx��_Ŋ�������=��Gz�7�E��Dʘ���,"ʬ��V�+ȗeYg����:/ �Y�i���E��үV�	a���z���i!��B�V�r߫s|FrU�ӱ�<�I�H|�V��%&�ry���x�}Rjo�(P��%���L7�LJ��?�9������T��C{��l�^gvI�"����/|��}���Ϋ5�u]A���Ԑ	0!S�b�2�#�cB��;Fk��滦"Y�چ��t�c��X��3��,�� ���b�QL'B͞V�h���h=p��V��6�����(c7[�������1"�ܞP��wHoQ5��ƈ��Wq	�2t����*�iuSS��1X�{�7|���ӻ�_M�^ś
�(	أ�6�j�Se�[��w*y�Ύ����9Ra/�4�=Ru� ��}����G8��U�e�L�fQ��D���
d�0#�h��~��?;�O��O���Q� "'U����*��]��o���\�h7E�p������`�Ǉ���	���4��ӭ2i�lL��Md�W_9�X�Cd�j�m��gZS
iW/�I��jݧ<N�Rx}��.�����zߖE�W�����gYNߤ˾�㗆�x��Irɗ���|1`�MF��To��R�ާ�\��P�(D��U״��\��M�0���R��l�[�N"+��J ��E͜��Wj�q���{hA��H��
�ӳ
f�3�y�.W���XX�CG�54{{���3�(l"
��,$�MS?���U�X��[�X4�C�+Xd+@Si��=��ov]�������ii�T�I�#�m�W	֢魿�{PC��Vk3��8�$�4�P��Z�Dg���0��6�25���#��a��r���yC��B��vx��4�E��x�m1T��K5��H��{����u4[d۟	�h�5ږk�����GUOY֭��JW�y�M�����8�KEc^R��hـeP�v$ �Yu}a�r'l�IC����j�A��ZRA�p������'���d���|<r�`Bk�{���ϐ�6>6�X}���0F��F���Q#�� ����Y�*ʿX���<�ͮfe� +�CG�l˺��3K�8ST��S2 ���1�S�g�Zwlȴq|6��Y�Y�,� �Ϲ��d����s�E��)l�qJ߿`1�O6���7���ޑp�i��T�ʴ0O��sN�o`��D�����}\o-Da��d����p2���jA�7��H�A0����z���M��/cϵ��΅����:�lYH��;
���= jG��.��~�T:��N��?�������nЅI{_t�Ҕ����(d�b.��Rl����_\�J�t���t띺�� 3���$�i�ӧM�4w�����va-0���LK��i�Qʹ&'��]j��K�_��%'Ή��^>�`��m�Mw��^�"�&i��������!$����%��KV�ke.�w(���ה%od� �.R��+���<�~���ެ�Z%��A�d�z����}�;'k��	3�4�R=�Y���G�Z}O��4�$��وg�1�A���.�����U��T�����Z0=;t����s\�����H�|�/[�s�`��S�#���se���ٳu)�񉼕�zՈ�=��sT���xL4.��ɷ:!�=���#O���	����"�~�Z�ԗHu�?ｴ#�,�g�i�(z�W;il�l�]�v$q`"����Ɋ�e���%��W��֗�م�>8
8����(�\�n~?:�:��<��\�O���%C9�=-�Z<ˡ�N��BB�|e���������gR[�+�aF�Kd �	��?D�(��Z�/Boª�5葢cS}�-4K�0B�_glyojb[]�#�4�NT����v��;�� �)5�f܌��mtQ8�G��F��?Z�����55���T�y�U&1z�Gb�|ts�.������7��w���Ie�_F+��U��h"o	����(�<��nI�%V�%p�F%I,�1��84 ��Gܵ�J؂����/�������`���t䧇�7�������9��JY-�i~S��	6��+�;��־��{&� tr�LDz[�H9��[�ǂu��M؄s4#9ӟǠi:��ۧ�?f'��=\,�f�����$�d��¡����ZAǰG�u��?!��g~Gd/^ŗa��i)����o%�|n���"f雽G�ڀ��L����~�����*S�L,s��KĈ�C�>j��l/��:��g��s��p�S���Q_Q��>�)io��J�_�No~��Q�O�[��5)�i2���q�_��@FȾ9��PD�Q�Pa���s�n�ln�i�(J�@(:�46��T��Ph��p����zw�.�ȗ�E�/r�w� ���.�9/����?�&�eZ$�"S�� M��!.$w��M��	�*Z���ebX�t���� 	=��ק��؀,J��S�fl(��'P\�r�F����G�,�lȪ>"ޖ}0
R�>r�N�N�H�y��ځ�q^"7��<:����EF�<ϴnƝ�8���̑w�|ƭ�j��
��� ? SS�IAs��5�@�"R6�/�#?F���z�wW�[/��[�N|�fV�5�@�Sl�p�<�hP��a���D��ߑ�?�u�I�n�	vo�]����6��/G�G�)�K���=�{�Y���|���ǱhJs�e���R��#r;O�=��BJ�e���Ƽ7"؛�>��]8�uٺ�TҽT�3\��c{N� ƒ��p�Ԡ���^;�OXBXJ���k�.UO�#�u�G>6V�Rn��C{�#�*��� �U�h`>bD�����3�Up�3�@��B�����,���s2���5`FqA%��"gz]l(�L�/��b˸@)�e	�LK~�]F�
V��(9�8e�v;A�N�>��9��	���:J�~_]�n��+b*��]�1�0�_���aM���w;B;��w��}��?+�A]�.���b����H����?�v���=H�,��92yH�x}�gz�/�@�vN	9�7�o�z��;p�DG�D"}���C��v����h��Rיo2���"��©��0�Л���\C��c���A���j�_��Q�#7�Q�O2GÓ���n0@���85�oѦeq:�����B�*�v��UK�@#��M`Q�fS�:ؾ@_�*_���Ø�����5wyN��rN�[dÔ?�h&`�Uڍ�i/ ��tb@tc�	��y�J��J���߼�*�h�;�`+d�l@�l0�w#��e"n]3S��#�t��;1K�����*7��?���FB9R�_��m�Α!��>�!�s�K]R���^���iI���|+�O�����v��8"��n�.1>�S���g��G��>�l�ՇO�_�j�Z�����f�
�����F~�U?��|��.�]���`z[C��4���;*������g�S�85Z��rA����1�1�^�o�(f�~�,��*ؖ�|�8��Ǘn߲��'t�n��E�-�ЀwhH�>v)2����Q��\����� '�.���j����Gq5W�a[�wx��2<�C�K<g�@�?��H��k�������W����s0��1w�==�CWn/B��
���w�'�&h% ������+�
�>�~�(��qHމ]���"���&�� SX�����b/`��t��w`��m^���>���&�z��j������D��P�>8�$K�=�Mp2�b�L�A&�ۧ�r<��]ڵ��O�&�=�U&��$/b
�����#b1<���o���X(�^�ѴvPi_�}��=������|a�N�Z��*BDh���+@�z"�l�����{S{�iy�R�����Pc�ڮcf`$CD�X��j	w|�nŤ��6X�����
�_�=[W�����|�FF>'u%�a� �)?��w��f��{;�b�Տ˸�Ѯ'�],`g���QL����1�}�8�կ�����\�D�8�XO2"�fbv`��
Q�m�z2�a�"��q����Iues�(J�#_ѹ���af�/O{�_�%C��+M�P4�DD��7����-S�t)�;X��jIEps�< ��z�b����.Hf'|��4n/���Th�c��)E�T2]�f�6��R/���_|�pۺTZ�#�k�}������&�ho���ud�[-E�pJ�<�$	���V���O[��B!	=������@�h���T9:���]��[lZKt�c�Z���E��R��)h�Kfw]Mj����|�'�,j&F�����~yړ蒦�σ�X0U��2<��U���6�Ԙ��G���=i��;�$��1��ُ̞�j�[����'}�@�/�����F�U�y�'�&�W�Cw�D[ğMx��g�P�����bw��G���f[�?_[yYr��
;��4爿Gb�BH,V-bL���h��n�%�V׸.�V�E1�Д��a�W�y<D�G�`b�k�ua���`����~�wyE_�����X;�Ȫ���AS�o��lA��3�=��	-p$0A�w����-:gi;�[�����!H��Fb(�b�����Z�d��s�����SXr �C��LI��w	3��{p���g��&N�.l����&^ ����O�pE����:�՝4V�!~���>9����4�c�*5�G�}��� ^���S"(p�o��?��7p�TC�fI1'��6��O���L��̛�1�j��!DB�j߱�u�Т�L�/��{{�I�64X#�E��?Na�}��b�\ ��Q�pE�u����n&����U�*�l�P���b�7�:>��ߓ���N�X*��DW���N�v�^�V�4+saq��g�NIص.���\��~�L��Ȼ�[�3�Pճ���4�o��,$�Է�F;���ŁD[��YԞ�a�F1�������-����.��_t�f-I���*P���|-�����{e�[R��^f'o�����q-uI��������0~76�
��6h ��Y{�'j�b<����A
�#T���\��?����5���� G	�������O�ʟ�Ğ<�
*�X|֏_�AA��o���~ee�@�1xI�̈A0�fDm*dt�}�j��U�}�Ǿ�6� � 
>Λ9J��ֽ��@�랍_� )�;�X���
V�.>�V�u�� {* ��t��-� ,����/5Y����l9S���2�����
�m���X0_E,?HL�
)��ϸ
v<�E�TN���{F0+غȭ�������7�;9��"|;Ә�a�čF��	�"U�&�U�ܳ���_b>G��
�`kh`5J����G��M��	P��;X��VD�| IkuD��-���Nl�IH�v�WV���Q��:�K�}�|��4 's����+
e�-��̑����c�RG�y�Pz�����YX�a#ҩ�4�,�x��8U�+6&WC��#D?Ĩ�����|��0�1�+)��`�]��b;��X� o	g�B��y���j�J~K��x�n霞O�c�
��������U U_L�X�$�|�A��y1��9��t<��tp����^�PCGk6c�vW��r��J�E�T;K%��:�\ҀVhh��Q}2��'�ϣ����G�D�"V��)G҃��pM?1�sW4�rp����7����z��⢤U�O�+̍Q��:q���Fa�kE���bc�7q�O���1Jv�������A����K�w� ]`cDZ��ǥ��.sK41�Xڲ�İ;y���m'�5!d+OGԳp���G@4�ڌ�17R'�|���(f�Q7�Z�"��a�:��d��n&�%B��k���+�׎�<qqvnXl���3�iE!j.�٧EHEAE�Q��aE_H�Y�ـ��3Y;
DqgZg�0�/͓���A,�F	X���O#o��߲f9@P+���lt��y�qYA��"�A/�<E�:cG�:;��v&Š�a���[��Ų��$�����!�2n������O-���H��-4�V�qG�,V [���,��@�����Q��V�%Y�^��QM�r.����τ��;[��!��R%k%3��aR��{O���a�e������"�۾|����Wݵ��\�3I%�/t�^G����{��Es�A�n�ڗD�\�9������p��j�.�����9��3Y��;�Ɣ����-V>�.�d^{�{��R�?s0��5�x�W� G�?�kg�5>(b���0(�������W&����u�
h�oSz���'�:�A���HR�b	�����JD!P�;v�ųksR	�0��E�ƭ�!�� �D�V@�e
����t�y��b�n�uU��u_'��f6�U7�]�y���+��Arl`�鋨�Ӛ��hog�A>��@�fR�}��t��q@1�p��:�ŒF�,&�Q��A+���!�
%�+ �a�ǞM��j��0�y}Z9{~������Y��!Z$�����n"f�;����*��v�����1�s�GIǋ�0�YR��� x�T��z�zp��[kĪ��b�#���%��YA�?v-��΃��}`���?n��8ZxS���I�Z�3aV8� ;�]'���~���Ɩc����j_5/)!U���|��C�O<�"H	ڥC<b`�Φ�Ew#�Uk�=7I�=x��;����L��/�:07��g��5�O�`Շ���g�p��>Ѱa��0 \���k׷�dU�-
�)@9�JJ�-���t�\�&-l�߷A]\	��a��Չ����7�@
�}|�Gk�o�Ⱦ*� �/tU�I�����Z9�}���A%bI��#���X,h��m�`�z=��{a�{�J���.d�T���7e�l�_aR�`��"K#KS|<	P�~|ͅ��16YTzQO2���x�3Au~:b��	��w_=^�>6���d�[#O�Zr޺0�"��U��6��K�*�I畇$���s����bnVek�����9��Nﭢ�j�l��'8Ͼ��@Ķ��M��Z>�LS��N�yZ�ǣ���{tɑ�(#]�>u8���\IX��-���]F,�濋FhCfP������	�{�dJ!����+Wo� 'z9�Bx�
N^�9�+��7i�6u��U֕�v٫�h)�2�s߬�p����HQc�"'x�0���N���~�"����u��H���(=M:�-<�^{NiB�G̴�%��Z[����*��<��V�k��O����841�/f��%<
t4���;A������s��������)�Cڔ΃o���c���ZBwq<�2�H�n.쫢jj'���~:�x&����nz�ϤAL}K,�ZZ�4�T7)�H��
L#�T�K�Cz
a�����j�f��ѕ�� ��h��Ed��*\:��\���v���۩�p�W���"�z������T�{����&����mk��9�q�RDӢ3 ����d�d72����e.~� �>"hel�_���"/}�8;�h�������B{��5��?I$W�rm:��c;�IHBe���Ρ�i��㔦�c%x�EJ��_�