��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{T#�5~e ���J�	)��2Z�2p`�
/}�dg�ѽ�c^p��t7>�lh�$1�c����N�"ؿ�R�z/�d#럶6O����<G\��Y+��6?i�f1�M/��C�������Ǵ����-(\������O���w��E�*�(3�B���򗤒�|�-sp���.����6%�.Q�@6�Qt�=�t�a�)~CB܍�c�~s�4V ��u^���^=[���2�@�C�9oM̏��x��4������y��m�<VߥB�(\�c������w�*;E�hvT�����B��棬��>�xe��d�c�%Q�IeU:��WgKT�Yu-:T�8Х$@���Ɨ�\zq�i��`3�c��*�Y��|�;�z�U+�jg�-��vb<�|�(���X׆����EݍF�Њ�<�@��Uh����m��s\|	-�^�U�|����ł���7��>�L_T��=;5e�T]�ܡ�+��z�wU�m��1yס��������:���Ts ��AG	�1:��aa"ϹL�J��4@W�G� �Y(]'��u����E솇l��#���c��'GZ�~�l�Z>�Ыl�Cls��ŝ���8���WB�>>�"E�Gr�%�n��n���v���*���q7��� ��e|ў�ZIj�䌊}�Q���J��E�P3��L���g��v(L�s�,��Vr�T�UH�����Ld	�"���
��ڤ�����>2�*��ǯ��7�eԁ;�[L��V�u��.S�4R��̓I� ��p��/�q˚}�|�g��,&�P
-.��_����3�h��S�"d���|��tJL���#���h0���[ ��,D�|�z���.�]ýɟ��n��?������}��|�f��j�P�R(5Pm	��j%�u�]��@���zO����K��̌`��{nu�xT}��y%[+GR,C�!���� :�׵��69��'s꣖��u.�����H�('���)�؏��8�W;N '���L�FŠ�h^��P5H�bA�Y�ۯ8�.BT��2�ck�
�uJ�g*e-0���hbus����a��J�LV�9Y H���k��F[�ו�!#�li�=벍���P���JA;j�y�Z1 ��~b%NTF;~�B`���e�Xge<����� ��D���mP������r���U8)���\)k��q�t�*����)Zd��%Ő.^�ъu'v�.6�E��@9�L�F���W�n`O�6ς	�� �ꅇ��"�f�j�H��#�L�\�֘�~Q{�*�mk2@}���{�a;�me�<sc�O�T2ú��Ԙ��a�,��/ep[
�J�a��>q�U0$�+��J����M�7�7���\�8�|�h��;Q	_l�,�ͨ%���P��U���č���3q��6k`N��)$p��"m�/bGt5��"�<��r�����H;�����9��Q7b�D���5��60=ue�4�!�w�-�CX2�پ`� ��n�d�Z_n�m`��| �SNbV4Xwݸk=��� %�d-�y�%�X��d�E4��D�� fs@G�9H}j�Vg�7�����������i̆��-lut��B��zV����E�������,`5&M�>���8j</×��ڊC��=h������@Y@S3�n��a�v���+��@�^�+Jy(əB����G*H3Ø�_��|<
|����{��W�9��
��v�c"	�&�ɴǓ�,΅ڀ퉔`�*E��6aS�qL<̉�Q�L��0����p`�`lV��D��2�˥3���qrt�URcEs�9��yz�ҁ3F"��z}|���wn�F��O.��HU��A�*�)��5��ЭN�<�\\Ӵ�}E��f�("�f%ˮ�CD�y�v�����V�3��G��O�BD���^�;6�q��{�\�7qT( �n�m�>xg�s�e�;�ϓ�\x��|�&AQOғ#��
9�C�������,�ш~۝�����1�&�vY4Ly�� 2�\���!F�x��z_Ao�ڐX�-�+	c՘m���A����pK�rm;�|���֘-_Yv�9��	l��_R\�df��b&���?;�ǹa�}U�ld�[+d\s��s��?J:�z��<����Y23��S�l�w ���tO�&n��(�X*Q���ο^Fd�nu�
hg�&-�;:��
 C�k��U�t��sx|^����N^
�ۙc�O�8ii�	���BJx�[/��kMTe���!��/_�	6ǐr?��+�O	��R9\�t ��IUc�[������T�U� :��8z�p�^���ȯ[����~��t1�N[�$�M���_��%oAM�};�����$���/5���j}ծ���>Zo��#��/�&�DK�^����p�+�]�(:)��eF������چǐ� �n��65DC��Q���L�6�l�L��}�on~�+��n���j8�1_�}�k�gZe�����@P'4�0��Dha	����o�R^0�<v�Q�W��+����� ���M�Cf�e��w�}����8����L��uR�V�*��ۢ4��3�����������-�N�/g����4�4�I��u�ٍ�6��\�|t?p�*�IH���c,�9:7C����Nf0�!�KZǄN\q)�=�2�:�R��]���?X�1}��:�a�����z��aGMR9���b����ɋ