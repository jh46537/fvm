��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���� 6�:$���mQ�$��z��˙Y��ˍΣq��pg&����&݂�X�H9�!��dv]E[5l�"h���L2	M��ݬ Dȟ���f,��o�Uv��rof����8�J��n�I<D ,Ҁ��N���w�5/�
�$���͠G�E&#ܽ�,L�<RX/�5� Ժ|dԉ<`��CU�2�;{o�&"r_�h)�)q�U����X����J4����Ģ+,�T��<��Kҕ�o���ѹV��e�:ܘ�+�`��\j�����Y��K
��N���T�7M�A�3����EQ�VX��A���#/{˅�S�M1d��uDSu������иY�VO��V���s-/k˥���8.4��vj�v_)7yc2`����t�dJ5�2�)����v�XF]�TWϏ �A��Ưd�9*reo�4b��!et=JH��`��T��#=.�DG���u䱄Ny뀺wL��4:�퇜�,@��[��ߟJ�R-L���Y{��B�	������g��tq�qC�GF+�=`��BH��+q�H1h��{��7��b�K��U�սT��d�`������A@ו*�J�=[O�Cx���X#�y�k�Wcz�	�o�R��'�`�Ÿ�B�8����1�h�����F���l��� �P)�&�6L]��L��	�	\�r�;�Fc�о6q\���.H�ejȢM'��Q7�Zt1:�����rJc��F`,�U�f�'�F�J�G����p@��-J��4��a��c��]l���F�)D2�'1"�ݘ�C�l�(�����rHi\��(}�A���ۦ
�)xn��i6-�B��b�2;�j�;|3S�>�p5JG�j��&�`��&�g���N��iϨ�C���h�ݻ\5��>#�p�m>U[q����6�Y�c)�$I�8Qh�����g:	>8���9�CX*�8��fm�ۂ�<�$�҉�㾭���L��t�R�<�f��wzΘ�2����O�6����^7�p� �C�����)�mB�\� _�}���o+�$홿�$f!�k�k�;��J]Υ�K����1��<��Z�=�!m�)	���`3�IP�H{�K�nk���>�N: $���<s6�;�\r�����G�̇t�*}ʧ���!��p�/D���We����t���t�=��9L��&&X�O�~?S
oa�S�gC���C+؛����~Ԩ���l���Vh�O�t� [1�0V�G����~i��S�'{A�un��Ֆ��.���+��E4�}y|v�1ݹ�G���?x=4�u|zE�>�>���c��F5=�`��$?�����o��c�!P�CU�Qe:t�^�����u��c�q¶>�GM�L�� �%t��L�s�8!.�8�u��[	ћ��y�y
�ֶ6!\#�"=	�OEpi�X���{� �,kd&|.'~�e�$�Or�x�!o �ɀoW���Pi���Xjyƶ�� Mv/`��%�S�l�K�I儘�sy��X�61<俭��Ap��KL������7~�ߒ�A�<����Z���L-`R���w� �jhho��S����؆�d��/o� �KO�7빕�53���G�����
dH��*c��<��'zU/@f�QE����Ed(\FV�!�G�Fӗlݺ^���wwE��K�9�*c�JM�KtA�Às�����r)�6���H�E
�SR�Q�Ĳ��\s�
���~q�U)!Gx�����C��냸�.����7��}wQ�(�>�(O���|��3�}��ajo$���Sx���HW���N�<�����@%�W@��vq��Ę]�aS��7�_S�M;�\�$P�H@�
�V3��g��xܞ@֐0�,�
<�b����W��<2=C�K�����E���i�A�9�;x.d����~����󬐜8P����u�F�2��Ǻ=�A�q�0k|��M��l�2�9�-Ոu劻/�^@CS�1����t���q�Fd�
���5��ݼ>V��M�2��7��w�=���E���\�L�vs�-bO:�_h��쐀��G�b��Y�C��5cXx1_��ԝ ��m *�t��$����>et�%Z�C��o�k0`�+����ͯ���,��M	ALh�}���;�Q,�~�
﯀�]\sx_CB���v!˩��}	�>