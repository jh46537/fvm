��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�z吴�)b���ΡrϷ���	�J�`,��1�{d�����߰{/б��R̟�I��!�����٧g�� g�~�N]�e k�#w%�5^�w�;�T8v��D\񐬪��#�����%�K�M|Y�Y���a=��J�Y��Lu��`���4I]T��]jg�9��Ko�8��ן���8��(8;��ŏ����ۈ�0"�qE֭�^C�fy�?~���O�u�/9�}�D�m��j ާ�xF�}�"F��W����J=GH]��ݳ0'���;�ɵ��������G��Ӿ��6�]�����ɪ��+�p����OYβ�m��.�\鶐�#�O��4�r>��uc�x]�.X��D�ye���3�`�����ϛ���G�%��s^���wJ����X�)!��zX��$�h(J]��}.t�c�L����!�_�8T0E�ؿz��Er�sM��i��B����*�8�����ç/�M��0@>�o7+4��V��*�A0���\]�z�`�C�	W�|0GX7�V#�)ά�xB��쾺�c
����t�Edj��� �]Oa�0��~!����a9���>S��}h��'ލ��ϥOh#=^�� �t�C�~t~7}�������2�k[^J \zt�η���E_�#rtb�n�,Q<\���,l�CL�����Rs<C,�׏�g�d�Z�V�8���髷��7v*��e͹O(Tg�}�MB�
�e���uW�",!���,.���q��ܳ��g�E�,�����ۣh�e���T�0�w�5�w_� ���qWF[9rC�(����;^�DS?ܞJ� /ϴ�������ǉ*�Z�1$P�"g��]V%C��$y�N��s(8����v�s�u�y�0$m� Y;���)�4A�A����W-^�;G?�ź���Bpo��)�-F�Q�
]���N��M�j������� �Vo��hG��c��;ق�˳U���nS��L)��=v�6h�_���S��:�l���� ���VdM8��"rf���m2=~Jy�X��TT$�z�!2����Q^��Z�!�S��0�0��2f�$��[���g�"�����Lr�G@�4OJ!A�J�,�#0EC'=Sko��Ur�<��PM���8ev��?�}�h9�znp"��Ƕ%%!��#��CTi��l�ުȨ��2���4�8���'8�з,���� ����Wѿ(u珤�<��5�:/�N�|�Ӷ"!���'j�g����>D�5ƈ��!��0O-	�RAa�I5`��Q�-B���L�l�$*���Z���[e����l=����+����VzB\x�m!��l$R"f���!�(�[�PV�m��j�][VuK�[\�~ù�k�eE��]����)�Å�������q�e���v��ab�*�讠�� ,	�2o���%�l��V�b����F^,Bq���d�ڨ�4K��Yb6�[��f�{ۿfඦ$���jh���*k{����43u��:_��=>�`P<���]"�!�-_���'�00mѫ'�VA������`�B53�0ҳ�CO�S;jS��Xn7�Ze�`3��zg�`:����Y�̱��
��s�n��(�ɼ
�|��`��=3FIM4g޹�ÿ�Lsl}}h5Ⱥ�Ü}d��a������:�f�~,����>A� (cݠVIc���/����N��kvǦ�� ��c^����%�O�^��4;���m
�P��?d,�p+�D�����pȎI�_��K�������ɷ�s����#=�����@�B%�%����=�;��@l�z�θ��d�}�U���Mb���f�T��i�F�>>�1h�����ƺ�x�O�KA~A�ns 2��4�C#D�Ct&���'��:�&YEW\`�}��,_Tq�ɷ�?���r��ԍw%�:��͐f��jcR�*V_��.������¡�^���1�o�@e���V2�We��T�Gz�)��Lu�W�o2ĳޙ: m�,|���{�i/����ud#!*�ښg4T��@0]&�y��w	���kX�RִJ(��ՉQ�����~�V]�7�O��i���ӻ�UM[�L SP#\;&&�6�*J!�޺�.�����Y�]��aU�ї�f7p2~ �$���S��t�
�u��j�8�� 5�'�N���J� ����%l�ٳxY穮7�u���4�tڻk�=����� f��B�F}Ѧ5Q�Vz��0s��-�A�W�*�$]�fJ�J�q���Y�qƟ+�7���܆��e6w�ơ����1�h�}�$!#�I�����G�}���i�xGPx�Escv
x&(k�U���J�WP�����u�
�H�"	H�o$,��m4͏�D$�}]n����+�:�_ȏ����������v!����[�"{��1�[�a��y�Ӭa(�s�h�+>�Щ�px��:����1�tx�}eǘ����_�Rz��
����ԗ
т���4TN��8�i�,��h$�kCH|�&��33�k���~g���\�q�l���Xg�KIo��y�o�N�A���`љna*��S�P�Dk����d��L���_�"�{me�����>G�ٮ�ۂ
rp����:Y��=�X��iȠ_�O����E�i}���ғ|�-O��D!��J��HڇmO�P�v�|)�ۤ?sj|�k+{D�-0)���\��Ź������h�9T��Me����w����������I�[VU&������
��a��xU�� -nޣ��:�����zz5b�w��4R�d~ߔ�������:� B��.̫�#��HЊ��K��b��Z��H��Ka�vN��ye�݅dn���(w�k���*& Ek2-�˘VIkb����B����2K��6�b!�^~T�Oi�[>��Y�[r�gNS�(-��|=v��ï������> �ȪK��B���Ҡs��wS�exȖ
htx_8���sھ���?�����5ފM�_�iJ��h�ps�=�LMK,0}���t��B���u��z�(�5ͮ�
L$lv�֎�;j�Q�
T4"���R���Am��Pj�p�^ln�M�r�)���M׳d���&:�M�H��� ۡ�b-�h5�
n���^���Y_ER^��o���A܍!���}�������y(O��s:B"߷:-���&��>��j��7�~U$�
R	����<wuO��$ҚIQ�B���mZ���;h��!N�j���S.�@ѷ[:�������1`%<�ag�-i�H�_4�6��$�P�J|5�B�@��/��i1���?x[8Rb�e�-�q�X?i��zy�O��:p�^�^��֓���/rg�c�KМ`�o�L�ʩ=�s�U��#�Z�-bP-_@|��=�&�#vZ�
D��Z	kcm2O�ݍ�0�^�!�����ɢI!�n��:�d$�X�6���j�>�&���uf��lK�2Y?���Hw��^�u�-��Q�x�{xx�f���?��m�'�=�h��@+H�iJ����S{�{ e�)zn��\)�| Z�B�����o��F'�t����_x��� ��X�"'����1u�KۉMJo����a���y�A�m�ү���.�+��!��8��Z�X��G-��rd��g,.�ah�
�te�~�����M|�W�zcb��^Ċ�?���P���%�͏��1�����Ш����x�Ui92D��ҮasHD����`�5�^���5Y����e�i���=����],؟�e �l�/���Ne�W���NZD�(ҋ�A7�-�PV�a�뾹�z8�{�N�����['K'}ه���^�~���s����2\��=:�l��1���T�ᄳ1�ۡk,�#�]Ϸ�ړ��αϱ�u�
)�`��?��ư�A�h�g<ހ���m���*f��aN�ٌ�۱��(�������K�>�"}�M�w�{�	7[g�Նm�*i����".#���-������HOt�mw�{h��|a\QP�e+�������ӿr�%���o�O��$;�Nx���&�{^��*�S�P#��Ps-l'D ��@՞pb�ߗ1S>��E����~+o�uC�����2��i�z4������{ܷ��f<qD贍����W�윊ݜ�~4[zi����!#���6��x��Qav��l��f����1/e>�B������j`)`�2�I�+�T4��0���r��fv ۔��9>�[�WX�.i���!�T��G^�$���vS�U�� E@Rs|��q֌s��`gFa�P�/��]��Y�d�+Gi�)+j�Q��q���5t��8;`?(]$��v��?�X�|`�~W�d�+�*���k���+='�����<9���l��O��9y��V��)+�J>�g�Ѕhβ��<Q@���n��~l��c\vކo=�ڊ��|A�45�\�>M��\,���Շmd^E��^{� �v�l���N5v�V:�_��~��p3�	e�2]Tm��������K�9Lpsx>��Oݷ��7q(��@�Nj%Og�f禉2�E�4���A����F]g��^U"�^�9dZ_ۖ���A������x6����D�"�d� �6$"�|�Y���}�g�ܿM�m��$�?��/�j��j��vcbcŗ3įn�Ǆ���_!�cr�oK�3'�^��~G���f�M�%	dpy�V=Y��0Y=�]�b�m�1Y=���R�\2Mu9Q�M1����25!��:�� ����0��ż�PP��z-)�0��д�kjy0x�/ w�h�+�}4}^0*�+iw5�8�],����7|r��Iyz^������6@P ������Ĥ��uLlw?�����m�ap^
�e0xzvh$��BH,��0����s�s�	X��D�Eq+�Y�5�p�X�|P|1���	��{�ih��;ޣM�F��%�MV͟
aeqH,�
��+6���).��R14p��:���;�F9�Z�@���d�v�&
�Ph��~��s�P�bϗPtP�k��w�Wh+��4�k?����I�]��mhK'�z6A}�Q�K`A��$�
�N<ñ������>��������#XH9v���J�����~�u!�yM��yȳ�x��?J_g!L%�&E��N�˶N�ޭa�]4j�U���~	���9��6	e��\W�\����;������ŝ�b�&��I����Ӹ&��rDq�����9ܖ~�
�����S����Rg�Q�%����a�uStoH�!5I*H�*KX��۳'S�-��K���U�{� |E���<Z��y�s���Ae�ˑxn!�9�FRi��e\\�mX^A�)��`߬6���g�	�Ղ�}�p~ �0P^f.sA�Vh��
)�Z�t��I�`��4�
��OZ���1Us�LU��T�c l�pY�� �l�o�,C�Fp��O��
4>2�d��� I�qM&+��M���f:���O+���(�)��I�u���� $-������˩u��@�F^�g����{P�@}+ּ��\ņ�9f��
���2b��"�+k�u	�m��y�Re�y�ĘV�ʜU��&+֣k-mW��y	E:*J�N
#p��s>C�N+H{��d��x���0/�2�[Xﯞ�6�]/.�L���{ak��^���7&��T�'�4dQꭖDT
�Ozx{�ȥǺdV�_�"%9~�����ƥl����$�;�*���?7��W��f����|ȸR�P<�2G�bP�;O^p+=g�����i�$���~��g�n\��8N��-I�b$�4�f�r"zg�r��EHF>
#�%��_b}Z��~�I~�kMZ��lF�|6����z��1��٦��i����-�)uξ;���F���'�Д���T#x�?2c���!li�"є�-��\��*�Y�ʽ��x4�a��m�!?�i:���R(U�}���[������qyEm����M1[H'�Z�(�9��w�V�o�:}�����2���'�׶�G����ΐvW?c�d�Ob\�I��/�� �~��B�$�I��)���o���:=��֡z	CS�N����׾��#v����Hn���U�7���E!���`��>/���2�?��z�j��z�D�U�]�Q́�M;կ�X� �������!�-��|A�
�/w�z}r��3yG@"�0ى���8�g�&ï�c��_�aZN�$����W���6�Թ:dc|)�b���ُR��c�g���Q�R�Ճ_����2��~�덧��?�랾��/d���[�:�{��z�i�w��{�ӝ0���fN~~bJ��ǁ��d6��?�mtB�y��b4qmӝ�a��b�S���*�h��U�\ӼrAd��
d#��r2#��@ۊ^�#�6�%�t��]����P��H_яv���1EՃ�6�rd�j����pN��ӄj6_��Ο.�HZ9)e񋑳��A��@����lq�AX2����<�X�����x��R�|i�=�%���4$���#���0�7����4�<�C4BU�o{!-p�T�Y�aP�?{ �Ղ��e>*O�J�*MY��;�u����8[��픠Ϩ������zN���~��z�d�h2i���v��1��,�gv�~Kt����7U
5���7?-��Y{��'b�7T%�!*(��ŇW��0��Et 
k_��5���wΤI�C�i��9�9 *nt�� D5L'	��4���]%�Qu�|��i/���|�\�~>ի�ڍ�;���d>�|�0�3��u��\�q܇��(Rӻ,P���1��/f�e��S_5�]_ǡ���X�b�2�m���c<i"�t3��h^%1+��=��	Cj���˜6.�ZQ[�>s+<�3.����� �m4� ��.�72Z|?_�ǟߓ��'bGҳ�_�_ĸ���������y	Q�D*uf
���_G�Q�F���A,���� �>�_��΃�q.g{ݴ)�3?n=*������P��sJ�e��kQ�L�N�#g�N^�v�Xҡ{��ƻ���e;/�k�����S�n�4Xȝ`J��2�;T��?��/����{��c�#�,+g_j����}.z�FV�wKq��}O{,�O���y;�e.p k�s�WW�3�L��a�İW�;"�R/����yKgHw�$Mk�A���s�΢�U���>���hy(f�e�$N
Hf5��6?#��s�g��ھ����JE_��7�׶7X%���d��I���0����Y"�N�[�,n��Z5�T�����V^�'Pj�2�L��V0��pk�߹�y/�a20R��[h���ϪD���3����̲Lfk�Q�-��^յ5����`��j)l��8qT ��e&���&T���屼W����kO>l47����r<�w��5�$g��O3矰��f��9+d'i��vHpH�f�Ɵ���a����o'�s0t8!��x�T	ߠ�ԇ2"jl)ı��l��o>�H4��\�M`�<�l"��]�F����e�X�Bs�	�6�&sw^�h�ʜaLDJ��@�ӭľ�B*Y�ǕU�����u�����	���[D���aՋ�-�}(��n���eȎ�^^)�|�ŏSw���-^��ݫ�Fq��Ei�9����j��@e�[���$6����g�F�;�C����]܀�B�ɋ��V��Z����U�^�d��EԔK_Nv��w�la@*�S�Xbz��p&��P 㮗��U�F.*tg�6j�M������3�W��I �]+��*����p=&�	��զ�EBh������ف�l-w��{o���=Q,U'[=��,�8�h�������XA�;Gt��|;����ʇcU��	�tF=W��	�.<wb\���`�V���.�8�h*o���U�)�x�+����$޺��	�\���V�,���@��^G����?'q�<�Z~�[%���zE�s"�;�Z~�"�<��m0.���C}�
z�����m�~������%w)�iS���>�y�m�!��d�6�ڣ�!6r�}*�.pӍ�����z?�����24�FY�COu!U�_J_8n�.�\|Fw@���->���<��?���>����'�5>41s,.��̝pFUώ,�G���0Ԗ�ia�3��ߓ!t��d��7x4[��b-��-o1N��7�>/9��Bw�QqH1�s�Ny�PI*nQ���Y�*�y>K����j�$ni����"��r�y����
����|��9��I|K���C�qB7��k���Ŗ�;���z1��mH��-�y9ꗘ"�΢)]9e�DFy���呦o�S�aHr�x���c Q8��a &F�$�/�p���Z�k�����fP��޺�<k�V�Ui�wv���?�xzZ0�qn�j�d��U:¹j8����(�@I�:�S�2P�l28���ww9O~��`~����|�(\EJ)-�j"���6��p������Г������������Y�I�g?�{�����h:��k�{T���j�<?�
,�U:�C���`�ɿW+6�C���r�bY�,�[�a��a�q&����'��ʩ(���{13I��r�_@�'�w���#q�q�i���g�� ��N,[��P�ׯ6FsZ��|C��忳&{^~�H<�ĺ����Fb�+s���e%R_}"���Z�t�J�r�~�1)>M7;��G�Ox�6��4i׵�E�/�Op)����b� ���_\9��&t�z�i5o�����+�#�~�=.F����w쀓$����L+���-�W�JQԩ&� ����6sP�^׃�,�5g�~U1�d���^�n�(J˛�ŜGHൡcg���Xf���(t�d��P�|��-E��o�`]U������������t����q*�2&:4>p��#���4�ǒ2-��KPP�Ʀ������$�|C	
#=
!o-HmѶ�L��©�x�YW:K���)U��*{�1�RC�\u��_\�^�uX�]��%�3�)�����g'��:�?$�FU��knx� ��V�-�~�,�u�\߃�{��T�ӱ:�{�xp��F���ʒӹ�4&�0
h4�dS���0�J?o���"ߦm�h�ab�S��&R<��_�E�ǲ#���o���'&?t�c3,jc;�T��}�{&�K$�\�	[V�h���7:�2J֚�p��)�i�k��@g���'ް�)^�㡅�8=-�N��6(�04���o�6�
��I�D<��K�H)xe	�sax�,ڢ;�sCK�zUUw��3�F�I���q�a����g��$�JH���r�q�-�җj�obG�A�O9B���qː�x���{����n�޲(	�]n�=�OY��+f�1-�������zd�ӹ�7$��s@<���L|;�u]���Dw��B���y���U�$��v�\���w\Y]�Lm�@��]�"�W�{8G�������;�b�UBK�7w�q��u�9�q^n�A0Cg+>��*e	���f��m���8�U�_Hb�be4�B�^҈�1]����Wo� �򚳚૽ ��1�W�;�I�y�Zr�@���z���h�������tlH�&C�	D�6;a.w���s:��L�PB��/����4�'@$p� |Y�â�u��CN�M�	N!K�9��ڢ#b������MwN^Kp����f�g�T�öΦ[.��6��"`W�^ O*'����v�0�]&��F���}i��GH��[�.�|��&��}���:��	ˬ$�	QKR����&��	6_�ymY6
���d �P����ͣ��=}yE����mf�;�U��{��o���Ҳ9J��(&��V����;��Jz�z��JEq����g�s)�a�G�����������ne��W�c�����_�]�3Q�N�g��#����EC{�1�e��m�ufx�O�|`�%�)f���+e"��蘹&����&ݱ���b������&��ɕ��H�n�.����Z��T�C�P6������y����]W�9ԓg��̫e��OX�cɷ���Mv?$e|A�pL��y�R��rO5����V���Ǵ���AՊ��lpj�Oe7��q/�P3\]���C�ӗ��G@�f�
ą�����I�j(�O��!�����}B�4��&C�S��$i�a%̕j��++����
���U���a�������*eQ<1 8��uƶ��G��:4���I�R�����#�I (��8������w��v�[��_��Q~)��;�����=\�R��\�	u��|$�: �T*�
r��ڂh�� v�X-KB%��oIH��
��H��ʌ���!{ˎ݃����Dar�M3