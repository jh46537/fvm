��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�8� �vѢ��~ᮿ�G��.��B ��_��}��nJ
0l�,�n�:���=h�+ƅ�'� ��lh
U��֠� (���>X���yay}'�o3U�)H�po���Xa����.�R^��ܠҟD��z�	�M;�K!��Pyz�E�� �y��^)�9о� ��̀��_h�\x�z/a�(�BUe���ٮu�qn3nAF2Ҵ_�X�z�) Ҫ��d�>o�r��S�ׅ�b��Yw��l�'I�$(��4���ҟms��i��.�P�#ރ�fj�냦��᥺�=����g%dV��T��rI��S4�DB��6��#�^�ي�Vˈ�l�[��j[S�}J��O�m��,U�$�n�~խU*� 8 	���EQ��7Q��,�\�ƅ�Y�ʦح��a�IE2Ʀ��Yhf���Q�e�׶�����{ۓ.���ݩ3U��Ѭ�>��W��.p�a���[DJ�J&ˌ^���Q&<pS�"��4�+�2��
��t&�v�b1 
�n<����p�q�iL�~����$#�x�:{�QX=�>�\�GG�)3��׍\�U��wVT�ĆB��z��t��u�>��Xi�׉Ȫ�g7 ��6ꉻb�)kE�N�g� �XF�����<,��v�
�Ҥ�fS'��|s�6�W��*,�5�<v�{�⑂�Y-:b�Q�f�Q��vP�LY��u�G5��}|'M=� �a�-�O<�m^.�~0�g����!�
g��WI9��3 )�sx��r�(�08
��b\��%�b�4�X��*����"���GUnm�;���s�+���bE�|����k����N�#�~^�>�,��5vH�u<Z�mw��{{�69)�d�yr�j�8�#{Q����q�/f�q/t�8����D�o�׿Xͨ���I�W�r��1�Md=>�I�+d8 ���R��/���p� ��LbAj6��d(��Z�G߱�4Fe�oǻv`z�(Jt�`�с�,�O����9��j���5�f��g�@��M�Q�5)�N*�j>�`���R����[�wm �[���DV8i�0��h��Ǣ��N��ۨ
��S�:��IW�T�a�/Ip�{ �As;�	�<�Xr��R�sAHB�K�T:�N*�YM���(g\�o�4��b�7�t=�����B��L��?P�^v�t�'&I+�Ϯ�㠴O���_b��Ě�E��"=Դ²?8#�P�(����	���9da��"��t*˺�����<�g�!ƭ�� ET������+۵c��婆����@>����T�RA80���;��[��Y<��My�`S��$8���vSδ�}Ifl�;$����}^��	��*�������"L����wz�}��=9�t�K��q�	������Q�O��
1�V�fٹ����}���+t5�*�+���j]��-^$��p�T��k�o!_GCE���H�Q���<�@tD�]x�_͘\�e�k�Ĵr� �0�",Dz���#�<fwU:�"ۅWᑻbE}���uz�2t��#Z 
H��oLv�8x�R}0	�<���s[��?�����gx�U�eJ��C�:�al/�tC�HӦu,Qc-������0��h����n!�l ����=�̚�T
8Ū����gZ%U�1�s����Ba]��V�9*��!``l�G�ck���1��l�9кD���F�\��.�<z:g�m�����|�
�)����z^�������#���4~N��LjmJLTו�6r�m����KE@D5j�n��,)�G��-W�)<z`�h�s<�e����lP����X_�0��y�B�~/�@��ON�-�,q�8�o�Z�3�RK]��]���X�Z�����h �JzH�E� �eΣvĉ~�Z/�ٕИ�d5�Y�(@�ϥ�R�<F)��������jj6'������p�A�; n4��=�M�*L���.�w+�s��i���c�ĀX�V�;�q��A��q�`�=������G��>ec��l�T��A�b��e�ѹC�ܢ$��H�I�g
8BW�:N�o H��
�1�w��w{8��cC�K���$�]��N�;y��w�z��-�h�U�j�%RN�}5�3���=�"'�sp����qQv�[p�'����DzqY�	�<�������$�x�m󈙔0�7�+!'�Ɲ8�
���̒G���#�[�ucL���BMul���͵�ʦT�e�̆�w�����B lM$��-C`���*|PP�*�n|��_�뼍ݪ�:~�L&o䌫a�ώ�U�Mv�%���{�<�W�b9ֶ@�&`��H�j�4�@W�d|��.Ka��5y�إ�ҦJ��el
�"퓎���q����D��C%}�G����4�A|���j�����&��w�X��n�y}W�ӛv��a����(���Ov\W�}I�rJX3�YհC8�Z8=|�(?����0�����
�t�=p9^�0I,�S�J�2F̫2+��&�Ű�O����44S� ��꺂="�f�a�U\���,<�_'��i��6�랁&[��La�]Mb�Hz�h0����}<n?�ǈ�T��\am��yjH;Q�cD?%��'�/��G�jr�C����3K�7�q���$�Q�4�`��^8�(��$S��e���~(�#������l�#0AN��s2~}ݡx�Ѥ�C����m��Jՙ�| �H����`�c�Gu{rb����aQ�cV4��ٴQ ���O�l˶��huՎ��0�v���y ����+�V��$��|;� �Aq�a@�ѫWXp�B�ټ������}cG��lB�`��\�_W��t��0=& �����RP��]E�l5��5CNLu'�����jˡI�O��;��D����]�&�;~��(�M}���İ�!�^�	���,1C�����gv�h	��a���� E�¶֑�	q�����'���"�a�������<I��_1T���Jl��`����"\�?}�)�b���5鶁��������WZL#M�����q��)*\l�<6R�5�����4/�~�}K �s-,_�1�v�*�� �O!����w�"�Q�77X�(r��oQF�����wY�
J���؜kU�s���Hn�i�+ޥb;J��k��e�� z��qw��se�lN���T벾`d���M�t�uL�
�Z,�"�
ɥ��R�@H��ʟ��m�L�iܚ���g���M�=E�B4�-�4{٧)kmh(�ӵ��z請	��x���>�H�A�#�
C��י�.��n��6�|�G�����K��uNق�Si��wM>$��)�Io;���Ẹ;࿨7�F�-H��`� 6Z[���_�F�eX�aL���φ�iz��r7��/�)W���y�\�d'����揓U�b�U�'�?��-��M���m�ⓓ�"�ۆO�#�X����h�����B"bo����JR�ME�֭ć�����nvd`>*9p{+p�\H���;���C�����m�6���7�j(K�Qu��k��[
�YԬ=Mc�����Z��fl�5[�x���$	'�G���?�(�/�Dcr��k��Gu䱌6>˟ �����e^K�?N��*�o�쳱X���_9s-$"�1�1�?�+lk'/Cq�/�e'�4��}���sDt�y�{�I��J�LR�Zd���MzW7!/R)�{�ծP�*�k�L��芊��Y/��i�6]��> �y��Z�>*69-f��o��V�ۦ>S��rwM��U�} �R�O ��(c\o����M��x]JK��D�z>S8W\nZ��((��O,D�z�ϸN=��B���FD"��"щ<��W)G,��|�� .�`̌���"͚%zV���q�8���z�kV����ػ��v�۠jՐ^o�3=�~�\�(��k��LD��(��.��t�E��/I�b�a��K��O�م�/�O���:��[/:�C�!/��\��� )z��8��'��)�ϭ2%�'���.�ʈԭG�,�/u���H �Uzt
�$�1߯F��W��W���0>k�b�W�cxih�����8��L'���qŌ�`�=���uBe��]�l)�H;�W�ۑx�/�h��Z"�� �����߆QY�����w��X�z���y@?좹E+��$,x��#X7�i%$5Y�7-CN����tY7r��8�߲-���R<EK8��WH��К����U����<�~ގABf�����p�2R{Yz{����Bw�E	���G\�P�s�xy�E�Q��Pz73̇*���>�Op��r�"�h���/�_x��.=ޛl�q��3�6{ok�p�g���<5רSwPQU>��!ljY)b��-�jED���L�'�K�U�0�xZyE��5I.B�� �B�EuMDj�u���}����K��*��  N[�!��"?�-�+>(�nB��� ۍ����!�&���OT��n�ͱ�&�aqo)v��g{�C
��i��l�����+B�d�� �b���qQ�rK�#<E���W�R��l�Z�Ex�V:�K1kD����H��&���H���o�\�s��