��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw�a�[W;���(���=�+V0�[&���`�F�}S���5?�q
'�D���u�rFp�w�H�����H�<�hzUpH�Qinx�r��4��S��*���5�� �b���qޅ�,LAX!��X��e����D4��*^ZJ[8��k�D��5�2^�gL�DI+GbΆ����{n���?�W���J�, ��`��>���v ���U-�x�^���h�l�E��׫���W<~ ��7�&N~+�D�%�Ӳ�"�^ք᜝v�z��q�N�9����XM�޷~_yћ�Z�`��A�� �����.T�ttaX�!��0��$�w��6t,t9|F�� ��}�����gգA���g&���|��p&��M��A��O�����T�mԢqS���!�_���S�g�y$>�,i<��\�|�7��X�r��Ud<��mӽ~��:����m��;X~2��d	�۹��a�O���9�����V�r�NmOƅ'n�����]+2��n����Nt3��N�䂌�ERA˧t�X�ַ��3k�����jR�:��
ڦn+��&3�f��߹ˍ�SB��uM�2D����,���_�� ��'Ww�e0G4Ѕ�I ={��#=豗�]�J+��H�qK�]��	ʁ��{-B�tͶ�C���-A#���?K��p�lg�Dɻ$(�ųz>ج�i*��%�kh�lk�G�)X�_���x���fX6���8^��5c�o��P�>�-v��Ҷ y�������Ȃ��&��������,�̘�Տ@k��3]�~�3��$q�j��,0p+��\��$j�K��ڧ��b?ޱT+�e�.��G���-	U�Q&넑+N���Ч������ǚ�i�J���]�`�U��{��v�#VWz�Dƈ�ԬQ��b.��j������e���X�C&��B�O��l[��I$�id��; ��mٽ-H���p�嘾�?p'��X�+�G���¯�䫯�$��1w2��.�6���iͫ0�76���K�>Čc�Y��������q���j�KC�)��ӫ0������Di�x����/�N,�Ԟ�^�@��#!��`K89��E���[�}ϣ�b3���J�➕�9f�t�;@q�NO!vk&��r�=0��z��#���
\*ň�:�7�Z�����N/�Q��e6� ���(}t�����ߓ�̾���"���m��+ֻ����a�<m��[=�B��&�3,������c���#�P9
f��q�^��.��{|%wЙ�TP@K�ۢH~��_,8Z�w�v�y���\՛8���]��͈i� (i��[8w�&���G���`M�M�-�a}�������*3�z�(�gݙ��.0�b��>������e�IiZ(s�C�BU
�px��9!eRye�|Wh\|X.E������%c����5�S����ex�Z�I�)j
�D�Bnr����r��"���TrYk�|F�m9Ԋ�����m��o�;��d ��\�@�I,a�����D�����β��i- ��N����c-q��*L�XC���y�)� I]�z`%�~��ǹػ��P/1�[
��\�&��}������le�����K�t�O&7��޷&�{�B^�u劏�vr��0���ҏ>��0��v_�g#g��.VJ	��2q �$?�&Qd�y0���T�ۖ�=���-:p�cv!k��A��Q[��^�D
� D���[\0~B�#y��P+������-���0EM�7�9�r:$�S�'�{�c�P����^�H��9�CR&��hhT��C����Au>/b�'��s(��]��kl�B�'��4z+��\�|�^Y�Ґ{;���"�s)ի3?d{pw�Pr	���z�����sJܳ�������,����{�_��u�WA���Ѵ�z[G�"Y6iI2&w*KF�'z̸�1�˶��S��`�? h�����(�N��e�'^��A��Kߤ1��nW�
v�uv`�1:�w��4J��Ƈ�?���R��_����H��z|�T�?5����\��$)_���Y��5쫴��� ���V]nؒ��E�Tyv�@s��!u�����<��b�7e1OSQp|į�N��	�3Xn�l���.�f?48�_U�n�i��1�R2q�d#g���Jn���v�
��n/�1ChG̿<�=�'�~Y��g�Y��%�|�F�#C�&�ݾ�G�&�X�	7.�x��j�<�7�����QE��7�=r�>2��P�Ȱ�<�t��+��6��$�o�\�dRH�Se��h3Z�W�Rs��m<�n���NdFuG��H�7HW������J|�J��䁷"l��C�Ţ\sNE|����Zs����1%�F9a�6�i�ت腑��m��I#�\�A��ս2�R�ϊsT4��њ�9�Z��5�T����M��̪�[<��~.t����yGDBn�}ݚh��È�œw��T��*���{9)pC�ta[��\�J@vW-�����Pd�K������9�*�^�5[ό)v�M�"T�t�|�#�b�G�-x?/���M�l<���;KbZ��m� <Ε~h�$S�u�
��+3�����ݟ3g�������v5����7��p�Gkz�U*�c25]BΙ�_��J8��/�ه�)�G>o���l�:��E]���[_MrY�rLQ��0f�W��6L��1ZdEs�8��'��ܑ�'޳"q�mT	=k5��W�޻(�P�	���rzR�Y(�nO���O���>��O|�d^�ŉ��:���5{��b�Y�d�L�~6�I3����K�ϱ	��7�}�������<~�#��y5)'N��]��s1�M�"�e��[�����of�ϸrce��2���	�R �twS��`]DS�8�[}A��U@�ť�|b�h�;KRTsO�)�[�-�v�Z2��돔�E�N1v�DN����u�1>���h�pfnsj))�>R���mX��V}SL���ոu1�.EtG���)~-��s-}�k"��u�W��V���oQ�e�XFo�Տ�>8#S��i7�V�^���K"n�	l��cnDпIK�ͽ����j�j<{3M�Ɲ>�{����tZ2j)�j��������ۨ��5r/HxPGT�a��=E5Y	8��*+�o�J'9h��1�������9�iPF�w�{�W�F�;2޶��b+��nR��K�yW��GG9u�J!�w�T�� r��s�T��͆z����c���G-����$���jT�c�V�|ќ&R-� �axG�!~k��t���S}y�hљLcV�3(k�����7 `I"6TN�%]{�tߋ{2�z�<���H���^b��p�cJV�Bb��ĉ�i�2!��605\g�3��g+�{޵��i��<&`��a[�9��9 ,k�jn׭������$���ܴb� �v?�q�P0���Q+�����^i)^�\9��|��[K�"�1��~"��Ht�9�����X˄�X��Gz��K�VtґY-��n���b�B�C2�կ��eMU�4B͵ih�����C��c����t�=b�9����h��2�;٣ph!��k*�-bMS��x��Q�emtw�	5��%�	�a�����ȅɟ~��������@q�C,h���!�8ef޳c;}��%��#F������/>d٬0���w^��p��j��@}�O�G�{�J5A����F�ؿ��ܡh�/c�g�!�����^u���k��%�����`���0�D�F�G2�c���%�
R9��4cp��?�8<
�R4[foj��!�^�Ǣ%Ք�h��02�y�~��ɭ��"��os���2��[d�k�Y�`����.K������^걄�l��@�%]�vlV'�e1��|
Y-U_�F{V�wय़U�q�O���}�Y�^L�~��V�
VH�<����`XJ����r�"UE'�XM���J�Y8��T
�aȪ�?  D�IX���7dcb��tJ+IF�&D��j3G|�!�m&�e5��@7�	 ���/�5o��=업R�C�	f�$^�3iTTUf N�J��.Aԅ����*�(k�{{	`u5�%�