��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���|����*�%����[�"�nj�E��p�)=^F���gw��;&����L�P@���L��7�]3�Ť#�h��uu��v���u)u���t��O����>��*�c�)H��w=��>Ok�:s��5�x������.��<9I^ͱ�|�56�)��Z3@_�z|�����́���&�p��ǬZ��:/gC��ӕ�u�O9{<yvl
�������z��ޚpm���#_:kT"��F���R��Gn�21c3��^^a*/�<��#:;>�d�d�F�=�}�������O����eQ���3�$��JX�8��:��I�	�������pP֩�41�KY�ۖ$L1��\[e2͈cT�}��y�L!�:#�tG�^��j��tؗR�՟t�35��ts�b�O��
�Z���?YG=P����S��!��,ԣ�5�;�� B���*7��u�
�K�ڪW����#���h�`~�Ө�jj��;0\�+f�YLE���Ø�A�����$�d�Y����`�ǉA�ek�&���C��'��m�Ʀp��N�&��#�HR��4��&�hB�RL5�a������<���u�0�q09c�I�w��lE�Oh��.��?���؊�������Ը
|�<=rQ��_��!�I�\�e�Wf�� Qo�9ާ20Rğg���k����χ�@�}�=��� z�>��'#+��9a2΋B�g ��_���rT�"f�I���Aa&�ĸLyH��-����q.w�Z���jA\:�d���T&�S��z�v�#�rbz0��?����-�������Y#Hl+��w�VLn���>����NG�ttT̜�<�T���%�p\<vO�=(���;:�O��-@ŀx��#�ɵ�\��ѐp6�U4�^��3�#�!��ᕲ��>6�l=|�H�)J�x�h5�J�n2���~�z�y0�,�6���tMܪ ��q��T�}��E��^(}�m���w�i����e/-��Q��>s�M���Ρ�hbQ�\� <M��X,2��Kt�R��]/���NL�ܨ���M�㼃�'DM��GE��zc]��Z򄤡#~ΗY�HG�(��pH��Yh��GOY���A�'sA���)�/���m�?�j��܂����f(�hsG�yG�B���*I���M��&W�.�9��gZc4�H*�h�ʇ��i"&^'w���{.�5g>�w:�s�TC x�Ɔ�1q�(����ߢ�p�cRa����������h�@����=�QM��Z�%�8��m�Y���7߭��B�ׄS�wB�e��A	h�"�@����
9m�Ϗ��ˋ	���E ;�(l�e���Xj�!�r{CFr���u^g����͕*7�~H�7�t��A�M�����"�	�29� X��p�1��A���������������s�o�+��F_:�u�梐Ic����U�g�kP���o�Íq"�A�B�w/6�=ʣ휝�aɾ�����*����fmF��K�ܰ)^c�B�ⴡO�.R��ޥt�s�VG[,�,�]�z�¦�2�裠>�~��8 �.{�	Wм=�t\��</�w=@���#�P�۠�����˛�2�c}E���*rwmE�(Dl��DY� ( u�_��4��cu���Eoz��o� ��	���ؠt���|�&Z~�N�ޅ:t��d$.`�a�{�txl��g��e )q�?�2�:?��܀��=�t�y"i���3�i�VUY:�;Q�L�FJ�W����w��մ� �s ���}�Q$æ��R>Rw�O���$�V��cd�m��y�����3E.����`����섙�ڿ�L��~���w�w�aW�?|6���z7���JQ��}+,zf��3RY1�ￛ׸#�6^�HH�
L�Q�ě�4a���[P�n���j�[�Cx7�r��j??�Z�Ōu W�	�}�WA�׸OWa@��d�2֗Cfd�jU�t�*�w5pT���C�+Q���{?:'��ﶭ[/>�,=FO�U��dt��a�K�@��J�ӱE̹)]�@)�rC�2��qrт��D ��<y)�h�Rt"�'1��٭����^�b�-�'�,	�ː�w�	9��h�5v+�-㳖V8�:}�'�>��y3�]��)2����oЊ��8=\0%A8�u��g��$�H����6��U�{���kme6!���XD��/5�2m��IY}aHȮ|�����Zl�`�k�Ζ�F�1�I�c������rO[Aa��*������9H6�&>n��X��Vn��uc�*]������N��)rq"_K��{�h�0���4���ы
n��gb'�g/����T�vT�	�]�[o��_/���6���F�,����]J�#LP�0���0����� 0�������t# �|��!U=o���),�$��b�s� �1uX�5�9�#t.��zf���F�t]�y3`@�i4�yW��r,i��rid׸�C��V�E��p��7S���Ui��f%�x�� `|ӿB�Ϻ��>F0�¥�����$�����bI]���w;���X��<+]���D����y�(�V���ͬ#^eQ<ӧ�4�&/�\_Ͼ]������fUt)�l��g�I��~5j����H�QD3'=ˇc�/�̄l���>��+yBo6핾զx<D֭�!�~�9}t�ĠI//u�w����#��*�w0tǈ��S��1�4JO[r@���n�a���7�<���(��pBh�:�M,����	��V�\��.������n�Lj�,ҒF�?X����y�\�4)Qv^�ԋ��0�ݾ)�tHz��ρ�+�2�Ʈ��	1������{ �F��:���.q���p�Y���٠b0���Ʀ�����Ҫ,����)��k*:���&$�g�ڸÕ{����s�qf8�iյ�У#��&�� %�+ȸ�1�J��a$��@^Ĵ	�hۇ�׋�j��ȝ��]�Dh��<��Pް�	�� �C{�9�Q_ț��H��g#�=Y���ˀ	�ٟN�8����
�v2�nJvl)١8��'�.�K*�Z?�X(���>�Yf��T�/b�\�Y�s�}Idm�$z>f��E�2[R����12����?[�䂡qH̓϶�����xȷy��gjf�׸ �]=�\�C�3���(�&W���V�2ԟxC�1#yh+ {R�<~�B�s�Y�E�>��Hz������fKP0��s�2�[X(�wצ��@T6���s��_�Q^瀓;O��ݜ�I��lT����	8�%T1�z
b>�p��j�A�tk�����q�Ӳ�������?-�����m���h��e�$�����2��j۹QX�_�"ͱ8����e�|�Z� ���9�Ô�����捣/[���l	��َ������mh�vv/��߰�
dY�h�X?�O8ND_$��a{A�RNg9�t* (�
쀌Ʒ1�Sg>��\��>ZM礖OOL��R�'��V��q��.�G�Y��j$m7��3Z$Ŀk]q���)+A�݁�xsB����B��> �aQ: @V�6.1��%$�э}���M�e�M�x�lA�f�r��1�#ҕ�.N�\�1�NO�+� f$8mP!��IK(0׿���"b_�[�/��)���SF�s��w����C�h�C��J�lϥ������U/��B��v��()�1�\�p۲=��?RǷB*�3���ԯ��}��B����]kgd��Q�L��cX�nM��k��0��@���d�š�5�b���X�e���K��#L�$8���S�õ��f`.���˷�7��}-��^����?���d��,}/2<		2v�^|�����;�����9�[k�!Ǐ6�8�kg_�A��o�5�S�߁���yR���o�l�3�#⽉�M�:��`ȯS��A·n�u��[	�s&]>ֽO#�����h��O_	ǩ��u�]a��M��R
���+��j|������Z���ji�1�1!��2���S�h6hQl��v�O��&� ���� <.D���fG����E����۠3y*m�FF�tD*�-VK⏜���(���8��r��3p�#v����Z�[��@ߍp��_���nnP�8Yl�ƭ�t�������.jp���)a��{����O�>Q5���`ir$����,�5	�B���FY�ʇ����+$"�6��;w� �������n�����Q{E\��S�����|}���>l3���/k^����(��ۂ�pQ��W�+
�rn�/��`����^;:�8#�{C'��ၱ�7Ȟv7�b�x2;�#�oQ{qUܣj��?Z��f���w�l���S��������<�x���"�S��f�����[A
G�Z�]�(�EK����nCgmğa@C�~0+m��YMs���F�Wj5���P��sv����{���V	���vQɱ��n���I��+����q-��*-Pw��9�������l��4�F��Fyh�g�r�~�ˠScͥ\6o�?h��p�B�z�e��9�_�jݤ�e�unb��<q�d�?�'�]P�C�E��F��0�T>��:Mn���j�rˬ�@�"��_>���E�^�t�lq�F��u�K�B���P� 6��2=�[�V{�P(���M�F��?���ʌ��r=���J�N/ "�#�#��@h�c�����=���/b�F��Wz���z˒�QY�͌��u��*�}��U
�fIĸ<�I��V�tw���5ξH���؏v1ϥO��a�5T(�Lid���57y4���`4_#=�Łn=5X#������Ҝ�Z��pB$�DMͪ�lW�do#��y���C��w� �����ܳ�Σ�aB��u{|�F�����h� ����~��.ވAy\�r
I�`Ct�� :n�L��No�Y_D; T�#я[^Q��f?#aHS�͎���� �5UZ���r����Φ#���!�څau�8��=�5Bc��m=/"A�x�],x? ��"�۝��}�������d7)W���t���|�],����`.8_׸�Q\�����.�\7�â��Iy��B7��A�'"@{�y�X���!c��p��Sm��F�i�hb�6F�*�c�E��-BX-�2KӮ��^f��8�f
� !��q��Ji6��1�&$�2B��h�%\R�}^&����Y�Qw������$��}
���gJ>y�x��E��cݧ���_$ὼ�zj�ዕ�s��8ȷ/��+�w��^��[�贏���d\�n�[�7��X5���}��ȼ_0q�n8k�T��! ���hF�J��x�e����@�pM�,�˘����m���^�P6z� ���,D��?��'81�O�D�ž(�b�`���@��ܼ,��*��;��~����p%�r>z�쬤
�D��'�n�q��;�
D��"���c�shO/w����ZB=�X�dN�.��N�g":�(r��ۭ<@/1� �>?�B�����*�c�uW��t��(h=΋v �6�'�@�Ԋn�#<�Vs��u[6#����Z2O�Q��py^�ۺ����~�m&�	5!��P����:+��a�\���υ/I8�7��" �&k�y@�un�b����O?���^'b�cb=<@�!��F-�v��������@��:R��8b��ֿ�3���۔���_[\���-�蠋��4�Q�9�����!Un�Y����_���^:ufE���}s���`�U� �P���;��8�-�5�}r�\�M�IA�4�z�
���|�i#� mx89�p%82��Q����R���i|�7�U\�9�t����G9�M�w�`���#�%B���!c%-O�7�6�����E��"S�O�j�(�P+.3b�V6<pc�jxczx�
��K�[�E=�c������鰭��)K�_���+�z��(͓��0Q�=n�*��bx������(�!@eʶk#��O,r$��֙p� �=�R��p��mބ�d�r�>��0*"^q&}^��y�����~�}l}�����P����"����jc�#@!	`S��L���R���]w)���v3p�K� 9�ymo�UT�Q��ьIk,$_���ކr�29���p#���ɳ����D����V��^�8���<%!�2��&y2�K=���G�9�%����n}D�d��,j���!��;��><K$���;E��������M:�2 ��Ϣ���dE�:i+4��0S�hK�����-�{�txA�l�dį��<�D��q��'&�p�iJ7G8�UQo�ku���<����s-+����q�����3���r�064���Rl�Z���4C�xI�{��x��/H��SӦbY�y$ȓ��ych��N���F"��қ?��v#a`��ܵ�����n����D*RW.��,�vL�Ӏ޿��	�д`�*�A뮋�%��l3��0.!�Y�بy���e��G���܎J�#=X��fbW�G���v��p������(~t�26��sųN_P�=�"�����b��q=~����7=��	p�����ꋣ
�ԟ�3��נY[�9�~M�X��"\��Ak�h��lɗ)%�3_^�g���E�a�1�E��8Q�׸j(�[���*%m��N�xO�d>�¸�Gh>ڜ:�q�h��ŎY�G�]�+���%��)�E���{̹��d݋T|�8ߒB������3�>`e]����>w��(�;t��1�h������1��������qD�]��b�n���4���5�����%>[�X�s�T~�㰎�[��뭔�8���0{}:�cv�{�KEq5�WD	6 �ҡ�XR��xK{B��3��k"���CgW�o	��W^!D�(��ȩ�ُ�)=��!W���L+ְ�l�R��;��6m�W7M��@l
�ס[Ӧ�<t�װ�ɒ/��.15S�k*څ�|L]��V���6��蛔�aǕlCcn.��H}�x6a�5>��b;u�D�$&��c�2����;cls���dO-"6����Og{X��>,?���ǆ����h��l��jd���ttQ��$+ĸ���TU|�Y�������W��k�̀f�!&\�T��+�����gKk����*�R��f�ui���Ӓ5�<�Fs�o�=H+��LP��H7Ɛ�!�jL����6�E�E�
���Y	b�����]�>�d�$f�݈Fʇ֊LPE�����7��A5u��G~��L�)�T��|'4OHR�4�a�� ���|��&gJ���k�k�x3��n�	@�p��/:UeP�i��J�h� ~H��U�~�pi�����@HmY�	�@�.����m?�j/�k��a�T�P��8r����_��"�^����T�U�oP�4���l'Y��$�oP�RB�p��懄�V�vo��Wu0�sO�2.���:�hC_������j=lD��1�d�^�M¯>����H�e\����3Q�K�io���������_v�q��@�E{j�v�e+`B�"ZX��֨��r�F5����vA���RZ��嫴q�8�9��U6� ���������)f�:p�kҽ+�1W�W����L�^^G��g�2�| �G,�2�7�D�}�-#YTX�[������d�M]k�B�1	�^�uK�b���մ�#8�=�IJl߀;���a�@C0�־�r$Vvz�l@bX�N�X�͸��|�I�	����bY���_�a������Yx�-������͈����B�]S��]N�s�s�uZ���=�{7d������P�'|��?��{2�8��ЭN!ٔ��f΢���g̵(��(Հ>9�^�Y ��yª����Q=�+k-�0f���*Z�NkC/|���Yk��I;��'޷�\r7ݹ_�S\�������Z��J	��k_�y�Ⱦ��ꍧ1�{�F�u��+&��Ib���Bo��hD=�'U����C�b_��۔�;N��������o�^]EH@���?���4�=טl�V��b�Z,����w�t��G
��h����{��:�$��]�}D,�˛c	~+����8��^���~cx��N
�]�8F���0��Y�zx��U�ә]B�U�� r���v��f�`�5�)6����>�u%c�8��^�tq��ۃ��Ka=��h�l^��^�I.�q�"�'n�	wZg�&K���������ELL�O-0��#`7��i9��#�Ϯ�Ӓx�k]��e?�������9�ߧ/�����'����c���\}R�.<@`�$O�)2O}�����Q�e���!�p?�{� uA�{��Y�mG=>�b�4����k3l(�0��q�m�}�j&Ҁ�FE3Ơj�r0Z�ʇ>tV�t!�A�C1�ܪ�N ��,��n1�i�!��;�����":�Z�L~��W���2��g��ņ�67DԱ��,8��T���uJ�(.��۹|��܊���uPb�r�����MRx<vf���}��C+ V�[Ԝi.3��<�Է���i�1���Oyp����P����܉��=���w|[)o:5"Q�<��7�Y��ߌ�J4�����穀��CVg�@l�t �]�/��̘n�6��L�
�.t;$C;E�D�x-f���L�ۨ�gݒH<�ݝAgmܰ,��;���7�7����k�o�
�Ӫ�ٜN�����H�fkv�8sS����jbi���>�R� �+�9oĦ�?%�}C���<Kꌻ�hP�1�e��#��>��B���-]�	�^Hӧ�F:����}�,V��y��Rp~�*���E>,��e�m���ig��G䱇�1Y7�W��f�WheJZ#�ŹG�F���M�����7�F��i�3��~�K�b�����l��ihTa����kU� �x2�oj�|:!���SP�y]����oO0£�!��>�2���Be-u�`Ge� YQ�}�k\�S�>ѾE�IQ�2� ���)�
���G��	t�.���p����������.���P�G���`��8%ּ�R���Zd�Sӊ�G� GD&�t2ʁA���t�����$>f�L͏��I/�|��T�Av�
�@p/��~��X�ZpU��ԕ�� ���x���ɱWY��``p �	EK; �Xj~�vݲ�U�,�����7�,=��)9�aM�=�a���z$4!�9��k�?J$�P}G�4�*����G8j��"�ʻ�����u�D(.%�9ŔC���^Z 9���*VO;Yyu|e�u�a�\����/Ab�j�M�L��W�3��"[�_G�Dݻ�S����f��
�S1h�C�A-%
���a���g�0�2�zּIί
Q��0l�Ws#�v;_c��ǅ/��]uW���*�N1b��\�4�^�*�zj٠k�:jx�7����pPIE殍�ĥ��)$�`�׽f�ŀ�&_9���`�5��3�]�␽*"y�%�?���'�nW�������-��?�/��_���p ������	�|%잶�������T�s'�q�Fa��rS�%�UI�1-W<�a��[l��nS[���lZ~�ŚvJ����W_�UW6t��Q*�A{S���ￎ�hiS�j~����,��TWk�+��K�hF���Q���u���˄�]����EꄰՋ/�����W(	���ވ
�	y�U��u�����3��ǒ�+~���M��R��"Pk[���[E�1e��c>N�����<��9��=T�fy�аa����A�[�|��i�L��:T�c�q��% �m�塚-��M�8��'�M�$N>|�.���2��Lɍ�φ~�L�d��PPG�6 Z�xZ����y����j	�?x ��[�2~*��1�]"������sg�K��}d�U���l`���I�̪��'���k�3%0�����ka��֍6����'`*��"��
E�q"+���y�#ko�e�����gS��*�E�o��a�>8���>�����C��="<}�,�U��:J1���5G�T2�K��gg�OV���'a��\� �-*GO��	�dǂ�C��g�3��;fJ]F�J�?#�~���L{����@��J�Φ���L�J�.�H��q�h���VY;�yۜ����X�R��I�b��úP�I�QT�y��u��4׀�A�~�#��6`4N�w�l���i�S+_��1�[r)ә��A+f��'���F)��T��J%�y�<��;	m�d&�znTk�6�߳���P����d�%t��k�_2l��C���so���D��T������CK�?H9�����H��\ڝVR��d��(��^���l��|���:6��"�V��bcd]`��S%��c�<;��1!�ZV�.)���`5{Ft��K�՝@<�m�'�"��ܤ�����]Q�݀�u]
:�bJH7��/H�a���Z�Hx��C����^�f�ed@�`���� �pӍo���L{�&�$��A�.����C��TtΔn�Ϯ������r�������G����!Czk0�<Pal�_G�Y�%�E��K�m��uU�N�rH�w����D�hk���A�A��AɊ�3�*������4k�w��nt�<�"�v�YlX%z�r�*�S�*4#Q����8������1�$2���7�L�~�}F3�m M&a��tt֤a���܆;��Pg�� 3�J��z4���U��ݞ �	~�!ȑ���\�7�z!���� ���X5��&Q2��@�Z��뙟�\�Q#���52r��Q����T>�����UW�й?�*���hJl�.N�A_Uj�v	���rU�	PM�Z�)C<�T*勞888o<I�ƨ&d��Њgǰ��cw�;/���ŷ�oUC��~u�^� >�s
#-�����3�2����.}���;�$S!J��~[n�'��8�m1g^*w�*�K���n��uȊ��B9G�˜�yFs�4HI'�x�3*�&ܗ�������[�>�N�,����#YOA(ɴb�XD�~�'�^�3�|X���D��.��֮ 	������_N&%>��Dm�Q�	��z�X�g�
��!�k��5"Rd4��#׆R���S�������:k������@t�Aڕ�)SZ�tR���$� ô�8$�e�}�kz�Y=�L��7,WY2�Xޣ�bKW��TG0��Ռ!�4[��Po��[�Y�QӀ|�,]�%q��)���>F�4��뿉T(U�7r�C�bi�Fg��_����{�dQo�����M�_��v�?��	��������n�/�gk��(*�������z�x��ASXK�\�t�� u񊠍iSߩ�*��ek"Ǝ��u�M_ZG������Kz���F�'=
%�CM��}D�ɋ7��A������9́!"<�#0�4��c���7�Ӥ�>���F��M���H�m��E�%�����m[RHj���{��2Dh���DpL��p%a�\�8as��3��R���a����F��������o����jdhҖA�͇+(co� D�g�h��[%N	3���2�l�A���4�����_���ERF1Յ�Wl�}
�tg�gPj�/I�Z�U�G]H��No�H|�[�i���G�{�^��&o�WⱙAx�;�_��{}a�1ܣ���/����7�Z{]�eS�M�c��uX���ͭ��d��L��E�Qs�����h"r�9�ݰ �zYP*�eS�w
��\u<��<	R�@��������ψ�!W����Nv+|�mҠL�*j�f1e�4xHN�)�w��i, 3 �ע��;��QΞJ�(zv}�OB�,�>S\�_8�
(�s  �kUaXw䂮8r =8�5�r膯.F�[��1��=	���>*�����mƆ���J���v�|a�8�+lXwf]+�b�����gj۝��Q��&����a�ҷ	{������AǸ�8Y�^���F2��aX���2�Z��k4=���7t�?�Ɲ�>~0�):��H�'o�k�iRQ����Z��Dig�6�x(#Nz�'7��V!۝ȎJ��V��nt�S�ns���̦���<�&���b�k~�`���7s@�3�~(������v��@��P���SW��<ȵ��~v�^��}�U�/�+пqb��#��w�l*.�����7���^�`SKK	�k#��E��>0z�~A_B3����WE�]㿅��R^	��h)Q₯��{0˴i���L��z�����6f10���*tV��}�l�_\ڝ�P"���8�k���Ǣ��+������Mr��[��zl����e���,]cn$5{���L>��ީ�ǁ�W����y���Z]#�L�-q�ӳ�E��f#�[o���(��jS�	yڂ�I�۾S^c�w�)�����Ă9@X�%�S���M{A��iX*�q"�e���s �������]WCe���5&�h�0Q�%/xp:ˊa+��}�3���B8�%�����O��hߔkFԈPXPr���Ԫ�b�'�CB ��[J Y�焁|��w $?�p~B�)���z:l�u9�Q��m�k�Kc��H�� �ʞ��4N˼�4�����l��*lfb��ysA%�Q������T�)�`FU?��'����^E�E����\dY������b_�m�(�u�c&�b��I�ijl��4���1?]ea�����J��T<vN U�!����-z��������`�����/tG�گ�]�x��8��`����oI0��A̓��.}�s��V$&|�V�'wY����������a��ѭ0�@a���eN�!D�5�E�m&�A;��CՒX{�uo&�.�\�G��K^	
�B����w�7S�侨i�/qQe ZT�;hx�i�fYj�L-�wO�eri[�E�]L��<����Ц"|jFWP�����$�u�
�w�K�LQ[�L8�Rm��H�N�V�W�${�O����x'©�*l3��v�hO>_tFr`o���2��L?�r��OM�y��&����D(��.!�@#���;_/3�e����[7 h=U�d̃ə�G�c!N^QL�J$��j7�$��!�T�G-�����W�
ů��YM��\��b�D��Y[gԝx���jv�N_:�B���
�\t�I��z2���6����C������4S҈�U�l�˜�����hX��L��Sf��`y�M�}��n�oD��:�\�@p��;�rZA�P3�M�5'��\�/�>�	`���r�M�N��-���������}8p���ؤ��v�W�¿�G}����ܐg�
�Hи���D<�.~�A��$���71����/P<�I1l%b9��2�D5�_��3���Y�3���p|a�\	��_哭ج&��8��Ns�q1�V��#�cy�+4̍�޸)�!H�j���[ZP\�t �6a*a	1�� ��G+�5,7����k<Q��~��	xkēe�Z@�u��x�:hz�(\��q*2S���(̞���:tc<�|v��r�Q/�?�O1p���j��
-g��a'����d �
�A��>���et�D��JX�����Y%G���a01?<e� ;sݚF�D���$�>�1����)���;����"��P���J��L ���࣋,$�{�w�� D��6P�$?���8d��J0��Ci�Q���s>m���xǝ�/u��l�L�FRr1��c4�tTq������u�O���4���zQL�z�6_�Ž�3yD���q1�3m�w����VA��gB7�<@�Z$]F�7�t��ƻ6�c���.��E
}����$�����x�4���-�"k�e9�"Q��b�;k�~6L�9ߐU�>�X����h����Ϸ�"�����	qY���,L�O�I:���3܎l?y�'���,��5�h��jƩB�_���jćc��,��;��B�a'��Z������PÉ2S�[k�a��kVK�N���D/	`�σ�f����tT��v^�Hwe�h���s �o�^���/|�@o����_���KnYa���
�9m�K��-:�3Bb�n��[-ye�3��f�s��@�Z,-��\����0vNȋ��~��R=*q�u!F���`�U?��o�j-Y�]vR(�)8t��r�����J�
Nx��1/���x��\x��z����3 �G@\����?�r튋�@�Gt�)�6�N�8R;����5��9*�F�VAl���oЦ�rI;^u&h\��w+�2��>;7��Z��Y���|U	w�vx~Hǘ���뮊�7ޭ7I��W���|��B߮��p2S`(��2�'rۅoE".5A� q|�X�X�gM�Q��}�-�a}�%DZ٭���^Ӯ��]M*z��u���r(��A<�b�:�b��jjU�I��C��7�����g��B��X��+@7�=oe�Hɲ��~��}�
�I>Ms���3��[��.���C>g��V���q���/ڲ-B�_�=
�	p]���d��ٰa9N�uÆ����u�X�Ё=k�2x?��
/��l��������`<�Uqf o��ţc��\�W�]V`�,$ԍE�,����&���tf�c�_t2�3�`����WM�sSz�w����=�Q<u�S���D���V;^p�:�k�m���8�h����OΜ����n~�ԟY�1��ݣ�ہ�$@���Z}��3��:�����޳|t��lZ�מ$��{�d�E�e��#�9F�#pn�ƽS�,� ��ғ�r*H���1��6�ܺ̆Kڮ%�`����9��r6D��w�~`Iˮ'v�Y�ML6�"ا Ȍn�7!X{$����V�
W}
F�dU+�}LA��?&ǆ0��9�/B����^��Z-`����˱�wٺ�u&�H�6썮�Ϟ�2��b�y�i�H��C,��s6���<�zي�n�����k'	ׯ7���7���W�y��Ӈ}������C�,��}�������4X�#lͥ£��?	i��4���9:�
�/G�K�6�@EE�]ԧa��߅��!��p0N��VW�_�L\4�ܧF���_���2�49�s:�Z�K���hlgnG�1�T�J"P��� Q��{��W�_���n`�4I-ެA[T������NN>b?i'��M��\��%罿|�`K8�����������%�[m!�Ɗ]��:�������^��M�8F5x�E�=��>�Gs�:��I��϶��ZN�4\N�}���}�-�V��7Q�@US��
�xUu�5�+��"�V��XP[��|,53�y�����Ӕ�$-U��ȏ�����&(Ф��C�qu�'S�v,��̐z�4���dT_�G9�S��
	�9wG<�&X!�M�(C��^���*G'�����H	bGÓ{�˜���vPԮ'��,-����%ɖ�g���|��Zz&��;x��P�[vM�-�����z�U<Y�^�����H*A���Gv��.��1]����Y���k�s��*���Z��w��P����zn�A�8褖�%��j�|B���-��Qr�&}�%�P��D�s��U��qJ��TZ 4�l�%��'��$+-��W�1j�y���ӫ������٥�fqo+�&Or3�9�E�ug@��}"�>pE�m�e���hG~r=�q�7v���ådvѱͽ�v�|��*����$�5ۍU���Ϗ��*`m��&��Sw�th=t�w�'`��Yg�V���J��IV:�Z�&��Nk%B��ʹ��d��}rfM����9�	Ч��W@��.~z����l5�>`s)0���J,��B�|�A�9�&���<���K���ַ��o�h0��a�85����8��[9Gǥy����?�7�9��E�G�XJ&7�!�0��rEmL���H�b9���Rd����h�^�P�0J�k�QnnV�}�U(SOH�Ff���j����\��g�ͣYPj:�O���1�K��G���\$���!R�Z�����NN��ʥ�����墓�ЂW1�$
���2_ٻ_ļ��/kL��25!{��1s*O��̰�d�7�ý����6x����j�ڣ[��E~���c@�7��p�{����
��Qڠ���P�h�[�l�%%��q<*���I�gSJL�Y�#����c'By�k)�kzs|$��a.�O�� 1	-E~"����i��&2���FR{/�a:;�v?�0��[�=+�J���3�3��:�4��_�V��ކiu�Gjoh���Z+4bC3��f֤P#��!%��sr�������ɱ���I�i��O�e�W7t���"���.U�%R����+{����ߵ��g���k�J�/Z�=(&��T�����}�=�>�^nr���pT�R�{z�p y�
0�V�t��[��=�̸W_�d� Q�_����F��H�|�0Kla݃!�YɽZ��qS�����z�s����� ���a��:���EZ�=�]W�:S�:�җ���� c7w���ݔ�jJ��"���a���@x�A�oT0�%z��x��wg���XE��߫W���������8`��i@��80�(�f�wh�v�h�Vg��$y2��)I�js������6�k1��H5SE&� ���PGj/Q�Bv��Fb�w�E�5˙-5��h��~�a�e��M��
����U�NvJ��H9��.�t�����D������V�$/�8�W��ᚙ\��g�K�_�纳����[e����m��6|��<�ĩ���
A��(V'�rk%����z�g�UĜ���X�x?�>���"�)�N:ѭ�U�
��S �D+3��_&��FIvtLԅ�2�h��#v�c�6��� cAf�2M�c!��B�dst�G�����r{E8sőO��`���NK�Lr�{��b�D){Qxe.-PO�p�7���r���Y	(RD�<q�ҹ�(�C+�I@�WA	�oP͓��06-�# � Лw��g'7e|G{AT6[���ͤ����Be�*��#?a��E-+��q
���j�6�_r���2���C��c:0
\����<�K��`oヹ~nV׬��Dק�YA�\d�4�n���6�,O7M�S��Ƞ��ouJ�J>�a?��ۊ�[��}��K����S&X���3'`bH�����Ú�Ȣ��B�?� ����{�%�Cg����4T�[]"�c�p��?Nq��4���|�����OFĳ�Ȗ�+����ow��U�7�A���8���p��Bt�8�R�e��T��L��:!�Hm4��X,Kc���gJ��Z��ʖ?�kxF�#
�N��]}a�Z������g��:��!<Q����vk%nΔ�8�hmݱ)5��^�w��s����nk��ʉ���Bq�k�����]�z$��_��E..��t��K)	�Q����@&���k���C��zӭ��B���\D�~ ����MG�1�$~9�@>�����}�U6)&G�W7��xn -�$��1�@��L�����	g�l�H�b%���jh���)����]	�R�jLI�� +��nW�R'��'��y\D��)�!��&r�ce+�9�Kg�v�*e�n2`���rr K�Ȝ,^�z�*P�����)�i�2_���5�5��8]ߊۣ�X9Em����=�%'0�0�.uG�����Ԯ���I�4�G��t8Bd���?;{�&�W�m�b�9�+	E�S5S����X;�V�tM�Λ���ɂ~�UX�P���t�.J#�GY�c�s�/�5�Ry4-�u.�-cB��	�m�]���Pjr����^R㙹��0�D�a��^�ۇ��������/���R�X�W��2�7|��7}�l��Y5$�����6u��AM�r�`OB{6��
촛@KpF���}ֱ�"$�;L���ljTU��Փ����t�pp�V ?�U�K�B��g�����f��O�$A�J��)C�$e�D��|����z�3��11�/���"�����m���Q�/LT�b�_��yk�o��̊@��F���eL�Kۈ I�2]2.�)���Wj��)�O��S_$62*�ĬTX�V���L�ez2�E᱄:.�6W�����pp����b@������Et1�5�ζ��毛Tz���q:"��M3'OYM�9�J���?��Uk��p�L/D�T��֌�!m̠dD`*��%�����9����u˱s(vm��4��@~�G�5��n���oJ!����s�����"K�	3�x���"���k�eU_涞��r���Ձ ��5�C�IH͚�:�+��in�������9���eau�6�vM�E�uW	|�r�/39ڠ�U|���ӌ˛��怉Y<��A�H�7 �xV��'oBa�m�g�W�z��h�D��q+P��%u��v�ljY6m;�TF1��o:u�"R��@��HZ��4A^�H��#S��?�þ�s�'p���6� /�З� UԤ�Nԯe=�3.(A`����ݱ��jd�IVI�ol����X�X�0g��9\�G���G�IrSdAz����iC.6ĳ�ψ�+����	'�� �٥���s�sΘ���QPW�	��9���͕	�2'ݔd��5L9���ס+F�9 Xo�A���� ��&?]�ѽ}&
{uM���a�lK��KxfS�Խί�*$dׯ�s-�-��z��4�����	�菎>C�8���WZS�E�D ���f;uWw���;_�����X�=��3~97��ti~H�U�V�Dc��B1Sb�}��1�p��#,.��������0s��L�+/�>��|J�����$}ڗr�����s��Jj�Aթ&D�|w8N�2$�C�M1�,���<��[�$ �%��mZ�f�{��ؠ�S����&p�4IB<7�K	��X�^~S��#����#�Ƕ����|�x��g��e�3�R���A�ߪȔ�qs1���
�t��H�v�ټ��e#\���K".Z�#6Ԉ
�!����#}���I,/s<O�T
���`X���)��}#�B��N�c|1�������#9��$�z�����|�W.�'cy"�h���B�Kr���J�#($����:��?g�}W�`]���D��yKS�@`TV�
�|�Y��բ�ҿǦ�}H�`�Ax����#�5*�I
3>��c�vI�����:����S�=1����>�ʼ�nbQ.� �W����lv��)�<��^5��9ݱg���Q��B�b�X�i�M�����+��z��M�]P�2��� y���n�{�Q��L$��Û��右��U~l�=�q��OZ9P�:h���?�~����$w����+pc�XD6Q�Ξ4��w�tD;� _�v"��$���Z{��)����z'*|�p��͸3�	 ����6x����R���S�<c��*�B�߳�ʻ$P	�{�iv݇J����c��@�W�[X��6EO����ٿ�$���թ��qN���i��,s{��&�oʙ!o�I�B*	iD�Cτ [���7r}� !?���l���Npu�!¾�Ö���|v���LaR8�4l�����Y�H,9���W�N����"�0�E�Gn�l�r��]�Fu#�����0�RN�"!�Z��C�SG�6��80^)�JɎ���}���29�//�b�>�@��yQ;�m=�}H���+�hv(���!<Yc1գ>���o�HAr�23���"�k�F���l[�:9�,h� ���*���{px�j���'é�	~2���<����<^?���)���XL��#�1���Z�8�<�338Ȟ�7G��sS��E����y�nI�.1Iv.ݩ�'G�
pji�Sff�������Î�2m�
f�l��r4N��s���f�]1�NH{ZF�كs ��b)%WĹw���,8ώ�o�,0���}�w��T~2��	��n��K7���4P�^�2<y���� ��ƴ��b�2�gfr5�Nb'������y��]��{�o~��Y������$��]���l��^ᜇ�O+é��f@Z�R�`�k2�~q���E`K�slu^Qtc*p �yh-|_��$gB��P3�pi�I�r�IZ#VA1��P�Ɋ�߬G�-��O�����Y�%H�̰I�l�7�q97�MVp�my}R��`��ӺΫ���h��n�θ������9��󞁨�ɚ~j��qM"ւ�-�g�a�j`y �4T\��F�]�ǰt�LD����p����*t|Ey(|��o[q�t��F��G�P"��'|��le�	�!�����+�6��|��d�_'Yx��-3xN�<�L2�Mzv�\N:��y����>H���m�o>��)N�v��﫺h\�%y&j�bLIc�ϴNޖ�b�+�����O��ynw}��9�|�ifit�u�<�2����_�;_�7�E`d�1˸Ι[�}���!���O�
o�P���F8*�U٭�a��OQ��`$W�9N 6�V+�{��KXD���ρ�����Ux/�|Ѕ�9e){�3�`+dYanX��k̙�b²�k-���Kcl[͙�-'<4���{�'�_D-§w����Q��Y�ﺫ���-�>ʄ�<�!h0-}�u���y 3��@Nf�\ hX��6��a+�3�r����TA(�W��=,8�������RN�Ɓ�JL��Ni;)n�o<�vIW]������j��Ţ����tag8�U�������q��W���O�X��&��>q���Q둌�t�I��眪aB�Ѭ�Q���qL6�g����f��q�;�S=���X�/�?1 W_"Y����VCL�m1sPo�y�����gbي
���B��s�cxw�0y�2�!a͘J/��)�P�г����s���:�:�n<\�Wz�J�k�Ae�}b�8�����(��o�����<3LiKg��(�[w�肾#�+V�ew��������p_���u:��[B������)�#��(�M�M!z��(p)hV�7q"O���k'?�����#B'��$c��/ ') )����ey*I�}<��w�?�~a��"+�i����j��v7��YD;-(,�RM��P=<��z�u~1ڞ�W"DTM:�I�l��"Zs����5]�6q�R���:�`�d��<z�L5���Zx0�0U�8�F*���w���%HI��ϑ��"��c�P)�q6���m��}XG�=�e����&�e���E렑��n���q=�UßA��Vq���i^��v�_8��Fz�.��loBs��2\� d�A2B9�n����K�'j����oj"��i!�6a�I{�/i�� ��jo���H��:ơ}��r޷A;��0CI} �k�YI�0&}g���Iw�0O��![�����S{� ZD��s첱'�E�Dw��b�UM\A�eJPą����؞�˘!M�O"�wq��`�q�}�/n����˚I�s�[δK�$�O�0dn�Nx0ZX�>��t��f���[qw��瑪`������s�T��UU6IX5��)������}
��A?��F�w1�Zaդ���֜P��z���J9��qs�(�xB���4�uQ�Ĝ���-�X��+2�߂��{m%AD�^�&�o�����0b5�J���/�{���_R)���v�(��sƏt��^ߟ�����}���6+������{�A����q0Ⴃ��]�0!�4��z�8Ԑb�c��=g[h}�TFy7G�>�;��H:�UKCw��w�<&���8G��<����4�H~���>z�c��ILt0�uFލ���o(����0�Љ��5� ��q�I}��� mڙ��}$�)�y9<����^�)Գ{��%B���_�pz8^�?x@h��1��5khN���&�� �Ew�,�;��J`6dE��A��c�H���>F�sn����X�������i��a	�a�O�"�_�u��]^FAKz
�KqQz.Q��W9J�����zy��ҳk����:t��o<d�g]�CdCyD'y�����e�1C�akE��!P\�.R-Ǯ#c�un\@��k�|�b���ߌ��h
��;��mm@w�&H��}^b��d�X���"*��M5�Aq^��]Hx��p�#�ޛk�����g#e7�,��
%yՊ3�X��A[jx*ꪴ�`w٪���T�����{�������A*�<�1o���������[k�|[֥�eo�v:ơ���@<��)lF�����VJ��J�%���F���i�CF�m���1�m�.l�@�)ާ�Q(	�?����f�QS�&4��T2��������e������Y�wƿ���҂�R��l�#�7�E���E�����8F,9Zo������{iq[�G_�]��wy�A�Kb^ϕh9�����W�;�58s|�"	�Ý�z�AL3@Տ1f�mH�!7�;�����Ve�g�œ�t�-�)|Vr���m3bV0f�;����^v=�B��^}�
Ot�9�CsS~�:�@��e����A�'�_�r����ɞZYA�O\S�6��盃�y/I�����ۣϠ�S���b'l�T���d6<�����YT�5���V�Y�E%��g�i?��/���P��)@��o�vl:�(~A2Ѭ�"�'��D)��]��v�^�.)�4&�`�u�0��8W��\h�o�t���C'7k�G����N{)���S���k�85����>W�ls���Ѫl^�+"��M.B��C�A~�x>M��
��x���:!�f��`�p����I���~��Fl0��T>9c�Ckl�9n�qX�ƣB�d��d߭�H�0�R��1�J�����+��|��r$��]IU�7�B�r��f ����%|G|�����3��J��G>;.�@���R x�/!@)�w~�<K�m�����Np�.���uLŅҫGi���!F�h�F��S�Ȑs��ͥ���c��&�[����%�xj��w��5�w�F�#G��[��r��Y*6����I�����O���u��]>�ί-k����L�?�!�䵖���*���%��}�¥�m�v������R'�3���JEQk��ԉ�U>��ù.�5�
���,�;B�?\���@3��s3����/��O� Q6�H�9l�?���,ߛ�.fP,�0'�Z`���`q]�*:�O���D+s���rVg�jp��XngA��2���AT���>z8�?�>35j0 ��*�0+W� �_�m��wP�c���oV�y<A%�T��l�ݯ�e���)5U.�ɲ��^��[ɐ:��ki1�����l�������@c�Z�G��֌f�A������K�)d0��ȗ[�R���8~��Ucn�	�����M��F��S!��C�{��{Ɯ!R��3�����t��, ����芗�r�I0�
믡��������++7O�����JN�)�nZ�`q�G�k���m
F�{V~��Xy���yH�x�o��i��;�
�0��
�P��T�Eg/�	yq�Zn����r�9>=(�T̀9�u��_���������:3�6Ƚ��P�`G�!���rq�`�Z�q H>6h�u�Wa��Y��q �lR�x�p����.���S�E���ms�w���wr���7�:�q�7"�"�9%�� G�Gi��X�@����y��=Rq'�}�,.�B�U�0���,�2?'!G>���j�2���7q{�o9��`}3�MRB��S5�.�o��	�o�������h���Gz6T����"���/0jk���0��&~�H��=$�čfK�� 5���3.�Y����|��R�P�&C���Z�[v�n)"�~�;B��p(<ꭸ�Mߘ���+�H%����G��s��'�x���ҍ[�{�Ϣ�7.�*���5*��Q�W+�����m$1�.*)zk�ױ����&Ju�{�e����D�����A���T�5H�Qm�������ᚓ_+���n%4{��(�H�}R������ґƣ�KSm섅��c[����!t��aLW˧�y����9��S:�~�).��V=�}y�*Ð�tWpD RK�#���$�(�˺v'���p{èfI�v)��L�����~��s����ꔕ���O?���'��gA1뤎2[�@4;ς}��sV�;��	�ipQ5��\�H;�Ks@o�O�:3�24 �4�o�?�] z�f��$� �W�r�ހ�$i�5�Ӱ�ʷp6�}�N럠�,8�-v�7�'�E�a�v���Ly@�B�9�MlxSW��芻tvE2.�]�슬��3�/�iYB�����i������ݱ�����4��(#y���E�?�O�2��5(֩��յ)��z}&1��勞#��c�<m���LHs��Jz�=X�I�B�j��Nau;�p&
A�̒��7q�)�6�#�&"������S�1pѭ#�
�z��g��X���n��"����ײ3y&9ݡ��0xH�O*@��/���q͡ȥ'���jT"5�:Q�R�� j�}$��Z�VNڛ_U�w�搱�j�SWz�����ǖ��?1v�_�8�c�[��#���^j)A8�ikr��b�%��'��{\#��c�ST�dUH|9����/��٧���t�09����]!���l{�C�`g}���;�-��XJ���/�u^�۱_�3S6�l��F΍��|a v^���T!�V��*������LS�N|$o���aǗ���ʢ ���1R�g��a��1�S>ԛ�:Z�ZME鳺L�����l{,x,E~�i8I���x��o:2*B*[A8���K�|��x=V.�>Y�˅�5��K>]�?k��r�ƅ,�wST��$�H�TⰁi*��4u�e_p�ǿ��׶�;q1'Q��'J	w�;�uEoVH�3���R<Z�����R�L��̆��3����V��|��g��o�t"U>|Sޫ�(h>U�B��F�"N�i��,"�:�����8��eR7rI�g�N��4-��_Ĝ��(���s��Fs�_B��	-��Eހ��8��\�����Ϯ�'�:P_�@�Q�=�:J@
�p%� �||�s���z�/o�O�xzAޫ��S�<_����R0���o:�����q������C�h:����r^}"��:x^�<JC�P���w1g����)�0�����DN�6�tp�����&e%7��f��UAi2*�9b�M�S���1p�� 
Yq�YUڇӳ���Q9�gL�
>����Q�WO�FR	׶��@�,D-�0�h�������%�F�ZB�"|�Ғ�JA��ڧ��fIV�t�7z�}���Y��ג���
n"�/�eb�lg�R��tL>N\�ly�>�A�f��i��<��NšĚ�(I���-��gX�qY�c���X�ԩ����x�6���~=����"äճ���ʝ�� u �t��X�S ���Ć0���@�J-���~�t�p�8�?��Z3k4�4W�;��-��TN����W��\�}d�se6P��a���k���,�LGd{)s����PWq���g"nU����~�M�z�p��L�NZ��&�2�Y�x��J?�CY�yk�-8r��e��8љ�L=���a���*-z	��HU�u��.J��{�p��d�X�.x����IX�6�SS�O��04�K��ƾ\I�'|�|#/�Pb8�8k�Go��w�'��7���F󛯃�WAIW`��r�y��V�����[@v�]�BEr����ܽ�y���Z�ڛ0� �y����HB'�?m�FXF��9,S��"�uE��>�]y�=����4��`"#W�٩M}�=����-6��[<��n� ����iaG'����a4c���_k����&�d\6վ6*������"��p�K��hh�>�Z&�ш��u"���5�p�2*��u|�����V,/b��^�G���ܕ�F�w �.-#{�M`��W�(��K&��`3�Q��Ö��V�X�wi�?b%t��QT/�Ҕ%')�I���O��%�Qg�I1�x��Rn�ܬC��93.$sOz �6u�25B�&�hRpE&���0�}�q���.U2G۟��	 �W��/W�<F}ߋF�#���_/%+���_�Cˢ��h�>���:��;#<��D?��Rǟϴl$/"LV]��#�|����xm[��d��F��� �����co��8��%D�ݽ�|�J��'�<\�tB��i�aUqpK=Ժr�xI���b����c$�/@�}�|rO���M@��~H���Stӎs���1!�]��k�51���9��s�3௓�0+:{:��ih~dQ=�C�AA���PٝC������M���W�hAV���)��uQ�K|��Rex�W���kC0j1���>��b�_���';�q°숇�Ed=�$b
�,������n�i�ۑSuZ��9����7��><{�U�T`�z��wƭ��j+�SfG��G��f�'��U�ff�6��H�M����A]xk�v�������p��k�W�kBA_SaF>�-=�q+�;��_};a��򈙽t��'Н���H���WmV��L`�2���;"�@�
!N}-�p���$��5w���y��|�0�$/��_1!zH&H�	MY���9^�hN��N?�#B�~9]G^�T=G�M'��I�a��5&��)2�!���6��`���8!
�