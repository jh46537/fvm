��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B����d��:$�馈����Vj P�d�r���rO4�`O��A��4�k�Q��)k���E�Z_��r�Y��C[r2ҖUg(���`�S�L��Ȕ`�?"F^���w�r������m�6鿜�7��~} �(Ĥ�n�Pe��	 �cE/�ݭj]x{�s=�Q�BQ��T|��-.Q�p��.�o<��A��3���$���'9��	�"�.M����(s��?x� �'K�S����� �kfI�Ntd�J�G�1Y�Й���eRo��@�*5�g�!�M�l���f@�1�&fZ�S3˶凨�_����E�2q�YW|���"��,w�	L���J��N��H�m�rc�O��k�#���g�T	�@y���c��v�Vu;O��h�ʆ��gi�	[ƁLT}[,�i�,�a�WC�׸��Qf���S��/�����|�c������}'�P,Φ�D��J�+�rޗ� �w�%Y�ڇ��;�����J,{;�m�Y�.�/!���FGI܃�x����BVi/I�j6]��m7�x�_�w���^��Î�6r���T.�ȝ����=��=��.��v�9����벸G�%��bU1]Z�0co��V@I�Rz��{���}�p{Of�G�X�jf�����c���{�D�]��r�%�S��U.ll��pyJ)��5[�67��i���w[{�M���!k�b�B�I�L���j ��%0^8�E�he7!̔�
I(�xX�R9J���x�#?�|�(c�o��f�%ӘK��S�Ɂ.jz���X���9DX�HK�N:�w_ur9����C`�h�鰓����@�m�t￝�y�q�2���û
�T��`]��m�n��/< �Ch������,],uJ��:E���y�,��E�B��!N�g��ҍV��jZڴ}Nie��,��;K����B�6�O!���u]�
�6����^D+����b4݊�q�u���\a7��)fT�%��V�Ԥ�ƍ�zY�+���H�G��ġK�E��S��Q���Â�Y��h,W��A��m
��悬�n��~Ō�(�,�o����R5��qx�V�b٥>^�I3c;E.ƛ()��M<����Gz���CYԸIl/>Wk:����P�'�����W����>uG����#\�Z<�@
>ڻL<$�l�=x�~����V!���$���$�ȑ�M9��Y�#fNg��(�R�$̤Zŕ L��!�6K�m�S_�`��g��	�����UܸH�b�ˌv1�O��5h�������������B��B�&2�ǥm[��q>�2��+��~K*��fsP�E=G`����x	�	���F�����h4P�8`�W;�O֚��7��DY:/�@�JH�}� 7Ǣ
��i�➖&�b;�w��3���2�i��W��������NîJ����ɬ��g]���V�Gd(����~�O��;�nM�� 4�S���F��U`��8m�7��Y�z��K���(%�9,�B� �&����Ѳ�BU5�Su�|���.�m��(L��ht�F��
�����~���K�h���m�o��'��t�&�*T�|�D��W��K�xy��ô�h�}���nE�[Ζ�děB���¯�,;.3�f���س�Y�A��ۑDG�i� PN�KZ���w�;�~�|� �.6܎����Q�[pO�^�3<���>�F�̪��{9:U^W��<�-�"'&epc)�� ��~���J�v��)f�d���2��k���(��!X�A�V���F�􍨷�A?Pe�m�{p�_?Y��j���~�"[��0�B�'�/�wN�R"ě�p�&r� ܨ3��6�8[�4����NqFdD��@�DAf/������2��ɴ�bZ�bmC��
�G{R����><�	q��s�5��%*.�ud=�8�49����
�T81��"�ܢd?tO��1�=����P9745��L\@�!,K7gi~��s�yaM����L�8{;G���3����L9Ҍ��y?���4{��	f>I�<rd����_���$Ғ<Y�qk���bp.@ʶǷر!�����<mQ�m✇g�l��,�0ܿ�d��#D ��C�ס���3P��N\i�����r�WΈK�s_Q�1<��GE���dlGÏ?B���S��|���D�������@�f �K�
i��2��P��������߹榗��K'K�mc�%�n�G�&x��_��p�[�J:�آr�kӭ��9h�Ͳ�[�������-�W �Q���N�"�}����L��>w�0�9�sg��A�{0�J{�i�[�G�<��u��p�&8����cgw��3R���ߤ���LP�ǩ%0U����}�O��<)p���=��4����R����9��P����N'm�Y���U��EydR�[i��{��n���6�m���WT�u�]V�"�ݖd.��M$��i�0�]0�{d�<-	�~
��������<o6��0iNl�m�(Z,z�[V��c�-��|8E�;'{wtc�ʨ��-�_��h��>�[��b&;N�WΤ��8�������6�w.TC��!V��8�Dd����Af�-�b@�btJMK�|Fu�`����IWy-1P=A�l���wǈ�(�wm��uw'�$�]g�Pȵ��7)���(0���	o3-�*Z,�C(�H�ۃ�������h�����f�:��!���nƩ�1�7��u)cH��ͫ�Yׁx��B#��ޏP��z�F�Y)-��P��a?V�ѥ��:��N�zaG����OS���'����!�����N�#�[z��<��OV�H�P�r������ZH���E��sZ?ۮYvEM���<�����2j�m��y*���kٓ�3�[�V�Ҝs<���'-�'�� ��x�Ы�y;� �ؑ��V<~��԰U
�J"��WV:sT�F)�/��QO����g�O���*��ݝǿ G����&�)Й8���{�r��}9P�|5 ��%�"1T����cb����Ͼ:�/3�;`=��tA�U�Ҫ*8��,�����w��]h�P�S��S��P�/�_bYq&�{v�6t��:�a�/��ȳ�3XL7o)�T^�V�E0�3���6���bR�m��S����%2���y
�Y�>!C\j;�:eL�θ�X���O_�J�5:}v �V��Io��jn��5�8hD�
���W(b^���L/X���NΦ7�}���ENB������O�E���>a[(���I�A?}ݡ�C����د�i��m"���ߦCmX���{���|��Z�5w{CκE��ɘ|��9����Ü~���╼�1���DR��[�T�~kW���B�ܰO�}`�C��5���l5���zn�ax�m��0��_�:+�o�^k��>�lT��^n_��Iۿyf�����{�:d}A#YȊ� ��ɷ�A�t����PI�q��#YGCO{�&m��MU��"9�𣰼c
�&�0�wp5I�#=�}�r����*�<cP�W(���x���S���t� |��B�>S$�_�f%�bPI;�*�Ȯ�(7Ϩ[� ⍆[�$΂E������5���˦�|X 9v�Գ�{dݍ��PwlȶE�����߳�]�L�����]��D��9웡�ÊMC��t��C'S<Z�	itV�m;������~:�s���3!������[4��|®'�F-�"�_Y��C6�
 ���u�����z �f_*���M�[n��hQn�$����	봈�aE7���5��	��$0+��IB4
��1�8J����T�4�ei�&	Y��3í�>���� �u��"eUc��	6�:�hB� j�~AKIr�Ū��\Qx�08��&��	�$[����R���ś�0
��o2?Y
�H׋�)�xA�9B�$�� ��
�^�ǔ�}TiJ��^�A���-~G��N���7�к2�7�(3zKY�p�~'ĄT���A�ZtJ�����$����m��*!%�������/��j$}��T�Ǧf;�4ߤ�����$UCq��a:UuEUL]?�3ӻZ�#uZ.�,4��ʁdAV���StK�/�At��
�;�%7��5�4ܜ�Ҭg��o.hQ,��l�h��U�zM_-���gD?FyRYc��K��́bB�Ю�����}W���#�X�h�Xߺôc9ˉ�r�k�H��p%Ov�)A�K$����3��?�7�tM�Y{�&��m����!�Gi���HHs��O}X�t\�HD��R�'���>qt�vT�Y�p[T�8�m��.[�Ǽ��J�+ȀH�z�9рo����U�AXŃ/����,%ڼ�k���$�'��侨�ʍ(VLv�G���)n5)��\�q���@�ؖW|~�f�P��V$���<�������ś[���L�>^���1�E�h�!DHzWk�s���i��A��y�]�"�V4m�g�L� �菱i-�P/m�Ƙ��*{$i���m-�g���h{bY����&'L�Ԟ�)�i���.<4AO�����(��|������Y�)O�]�:UB � N��Z�p쨝ձ��^\���K���hُi4@��<�,�i�:��/5��A��x��Y�.���?h��x�h=<�}�����B<��S�_?aʛN�@��qv���i��c�@ 	4�.�y���R
:���eyY�=<�O:�G���|5/x��b�V�M��7V��`������J(�M���^;q`�r�ߺ9@���6ԥ��f��h�Q�>�׮�b�S7��K�W�s}�UF�zqN>yu�^��
R�$�J6����ѐǃ_!rZƉ�� V�P���[�HҘ&>}RHҸ'��.���</���
W;�|`�����A{n	�7�x5R�Б��r�ϑ�P�Z����Q�uSg��}S�u�yҧ=K ɟ����#�/W��N԰5��<�v��O�䫇Ov�b���JU��P2zr�wt�5�UӾ�S����s��=BT��wyv��9E�=�,9w'��u���.N���|���j�,�K�WG�R�><Ġ�l�<�H���}C��(�����yBH��~W��h�/��+��*q�p8<��E��O�-�:��	��j��š��#]e�0�!~�Aׯ構G4��E#A �OM0.2�M�Nts�&A��^ᗤ0Y�W���@��\����F4�J�q�Q[/[���0ű�M|6�&٤)�fZMY��Oe�I��J�mv�i�.�j	W�&�Vfx3�5ـ��}�S,k��9G4jh���$�al:��������^Hg�1`)^�����ԓQ�:��Խbl��yѓF�.��B#�$�� {��(�_��Ia���q�Qf�e����[�n��OF?��=����o�=�,g=`��n.[��ű�b�@tU?�Z���֪��;���]�f�{>���~�hq~�g���<�UL+|0���W6<�No֞��rg ��� �4�Ż��E�X9l��!/c�/L�~�����L(D�F�l��՛N�2�ôֿĞ��n�/�ݟ!���bbAq4n����P�q���v+bz��6����Y�ϴ����,����,�>���}�?d~6�j79��^m�EWku���BaJ�,9)�!���z�����F�%_]�ě�5^}�d�=Og�k�e��m��~�j.�6]��ݦ�qKEe�~�/������=�X)5�_�%��m\���#'�*�蕑	�ǓZ�Jzj�N�^X��uds�|�X2II_�N�g�/�訃�G��<�YPE�z�c��BڇKAs�.��KE�;7�N ���bsa=)�(i�D�����-Ӣ�����,�;��?���N��ި�pwA�o����{N�Q��.�R�s�#���8�@Xѵ�CW��.�3��q/�=x��Sd�m+c�m��
C��np#���$v������Q����^x�G���;-q�C`�}(A'���?���Jۍe_��3���f*�Z�'��*03C��w���`e�-�Ղ��m��T�tzȑ T��T�D���#���tZ&���(L��k���l��D�z��x��׽�i�\��� ��pQ�*>OnTn�;j��Y����a�~&ܝ�i����n��t���?���g��扃��]v��A���^��J��l�E�`p����P܊� �e�T�1^A��D5E*hLί9ڙ��p)���>�w�-�.��u��#@c^.Y��� �R-G��-�|��J-�k~��Ǭ���6�����^vh��A6~Oݓ���x�����!�:"�@AD&��O����Z30g{I�*�%NP�z��KqU��<
���̮��R"�^�ßs��+Y��T�)	�����< �f����C�r?�
i(��'�}~�������o���R}6p��! _쾺7v�:h���p��b��P:5����ů89��^g��F�8xT�E.�h,�rw���=R�{��]}���B��H�n�s0>Q��_�x�jK�Ul���Xi���I��UvV,��2���(�t{�u�a�NP�[��C)p��Ǆ��2�ul<���0�[��߇"[[�z�Q�Y[%c��F���P�I(���������6�(|����1Q���y��)^]�АMc�����P�f�+l�8�����d/���c5��R�-�Y��N4����u�l�M	��c��#������� h�[��!�;d�P���SQ��b��|�~M9����B�C��şP�ƃ���0���4l�ӑv��91#%�����ŷ��P�8�����ߴ�_�������Vi5_DÑp����$Ө�]�:���f9��ֿ<�np�+&��ᙙ�az�ƞz���GϨ������oܧ�b .�AS�V�2m�nj��<R��czb��@��'�'�.�g�V�!Z�@��V]%d�`��'�P+�#M,"\PYI���I9JD�y�t�5@��P�rx�Wx7�p�$�����+�qu�	��[����-�T����F-��U�u�c���ͷ׉��uQ��Qw��.1�ԍ���mLF�$8N����0�L�d������L�82Y���.�rM��s786_��B�c��݅�jw��CYS�Q���A8}���"^����'W���y⋳��] �]����,�a�WMJ�$YS^v���`F��9�l]Z8y�<��HS���By{�k���f<�Ā��kX���,�z��1�-��}?�m|�,h�9�/x��(Q�ΞmȦ��jo��R�hJ�zW��XS�$��5q��in���l��C��FZΫό}�x�����L�\���o�<%֟$�ԧ_�}��l���O���T`���L�?RL��:) A)B�>^�&w`��u]܎\����	P��!M���? �c>��|�e�W��LL0����R�4���i3�\�<4Y��Fm�H��RX%�i�Э�	H=\x�t�;�K?x�8�,�wf:ڠ?E �i{@���I���'h�& >���j��������1`��F���]����v��/�)��!P�'�Տ���e���B����`�1疫A�ٲ$�!9��B=��BvW��͗`xw�vo���w���/m��'#ȯXx�v�d�7;3���B����?��l�Z6��x�L%���P^��}���}�nA7�&~�	#��E|����o���$=_�mzx�ƪ�1s�^�E/�/��GA�M$�P��<8ɢ��sv�d��V��
Q���
G�������r/D�d��▏�/Ŕ������q���V/�!H�c����E�P�O�<�D�b>N��C��(c�9+(F�^����6:4[�Q�|/�S0�}�T��F�MF�I����#<�����g��e���+7�jG�?:�0�������{�g.��4$���Ć ��;'���� ���3f"&ùdn�+P��z{p�՚��E����]r�y��<�U�����	)�ú�͛gS��G.MBT#V"O���D�UR�C{�aY-�1eo�Ӫ���;���?B��S�f���l�h��=�_	��.�W�܄~�w<��F�o�޾$�D��"Ն_�`�Q8�E���t]{\�B�
�D}^vq~ᄒ\hS�!�	���/����d���n����������(~�a�L4�V�NHh�+�=��}��Í�2���fᗂJ�/HZG3�n��|�P���1!
S8%��NE����4E��1p���|��Ƴ,?~)!��c\�s'���6���_
���a&>�W�0~�V�69yk�&9gE��y}��B�&٩TW
����)*D���&iN����s���Wu
i-�h�:f@�|r���p��(��JP��6�;#�~F�bY�L��k�� �3���T�ԦK޺���Q�]�R�'�6Ǩ�� ���,Ӿ�W�
?��t1Q��!b~�f��s��!���H1���x���GԜr�����;��ɚ�"�������8~+�����a�M^2�a����� ����V��3]��X �.�@(�Gj�2�J	CG-p�S�t�Q��=7N�=���8��7�p��Z]�gc�i ���RR�f�h�h��
u8�݌���5Rw��G�2�HO���@K�l�r׽+�^iQ��o���f�_/b�3�yih�s_|�xlg�7�����T-��(�o%T�;���<��c	�ܦA�fr:a$�u�7]�{�`Z�������K��Ӹ	��k�����ML��_�][����1�	�� �R��b�s��`ך����h{�ݓ�񤨜�Pǹآ�[WE �b�<V7}������zQ���S�,Q���ׇj�n'io܃K�a1/91�G����f��ksiRy��@�(��R�TT��dj̜Ba��T<�?]�����A�\&RK�S�j@rp�ǥ��͡��؛�o�)<�$jT�o3X��lЂ=U���Zi�t�Uاb�Ā��隷o��ޤ���h���ӸK"�6Y�9���Bm$�W�lFI��þ�J�ۭ�ZӴ�R��񿥋��"c/�G�A%/��yt���Ҡ��F��O@1�^�׮�:�@@�ג�$o�(�4Uc�hY���E5*�$f��0����[l�A�����M׸k����j�|ѫ�66�:O�}u�&{\"n�<��\�d��q�t���ّ�ޟ�^d�F8Tes�yo�����hyӭŧ��vK��#�p���mʧ�����;����`��R��"fѦ�M��GƘ8JD���1Y�~BD�
��x�a� [`����X����iԯ<Y�Z42�p�5��`1��nP�ʲ�"8Op.+p�P<-��P��;Bh-Cs�U��#���mH������q ���"r=]�2�ݑbMÊ�3J �ы����4_�-��L��E&�PL�H��o)�q�cJ6v�����d�@���>�UbfD&>�E�㋍�*��h��O1�Vߵ_m��S�F��6�Ȥ��s�f;y�C+*I�d�@b[��`�Ƶ]=Jܸ|T��̯a����٬�R�`��`�u��!FS�,t+�����������$�e)p��;+��F�5T
�J�" ��WE��ډ1�����b����������N����
쥾�ω4��8'kh��E�%
�u?�4L)����������	@�p��<��֛DXy���P�(u�\b�-X*o���rՒ��7������3[U��RU5Os����lz��_���gpK��:L�ct�o�}�,�b�=h�0O��I���CXHw0��z��m���P�|Vi��R�C���ђ��1R.U��R��PTb5�S�g�S�� �e�0�Ә��C�x�F0�2�G�<�k�#GpA�6SZK,�ɨ�'��UX!�H�R�+�8��O�}|��Ҭ��	1��G�×h&��H"��k.��Jg	�+��2�3�
�Pr*�Y�e�x�ps���#�6�.�Y����Q4�x����	�����H�;�߉)?�M��I�'��(�!�H���N�6wj�S��KG�{�
`/ա[(3>�z��.�h�}5������n�9P�ݤ����hBL&B�ln���;�Хv�N��Bx�gg#���-�l��k�	z�$L�n��Q����&�g�)�E�;@a��Q��40�Kqg�N����F�q��;wI-KM����4QmKE�����.�[@5g�ҿ�F�v��JI�h��w��ϵ��u��F���Ć����}�+u�K^a�E�f�xf��N�摭Q�O���"?����Pk<�ɾUd��z�a��B���Ǳ���9���O��
-�={I�s8����2J!�H��G�W�C�*2�����H0j��#&��$��@{{�.���*�J �_�C��i�d���w���v���٨t������������S�5-t�F�Wg%��¹�-�tjy>�AP"�S�>�;cnf��m��q�'3�,���<������'���"�j���	�K�2p�\D5�.��:��V��Tح�A9D������K#a_R;�:������	Ar��	�\s�4�d�n��Wk�� _���$t��M��j�?)�U8_lY�w����F��T��N���xzC��Z`s#���/���T�"?}�K=�����J^�e@�O�9zM��u]�Aav�XrV��Ku���`���/
�LG���Ψ�,�Gb�44�+2��dHv`�����f�i�OV��{p>�>�|���ͅ:K|C�h���V'����-���1�A�*��k{%��{x�m���V~�F��� �!�ml)l�"�<������$bH�1�kS�T�8����ڼ�3�p��o�;/Jo�kq�����蠣�,�p9/�7�Gb�~��w��i�#��*4�v�?}��G�!�y�S����;�g'���E��� RB�)K�Q^��D�&�<�"��I��\�f��)X�qGh�����szE��%1·���>bϮ8��؏�G))��eI@���n�j�Ͷ�I�3=Jڔ�@Uo���XJ�:y^��$ 2�II'��Z�����F�P�%O������{[��P�X�6Cf���ț����hpK�1w�L���f+w�$��n�6�pJ
��'x��z޵������Y>�L͹�[z�uCM8yC��5����.��b���
��3[��A\��K0�~Sv�Q��_�>)��ω��B�N�ǬOqɣ4�¸լ�h��
���ǽ����)K:�g��y�}cg�50��1f�ZJ$Zs{��I�1���}w6T7��i���;� ��MeS�W@�!vp�HoC�����(���"4��~F����0����@���(X�,LЬh�?�-'oQ�{~6�ο��4����C�R]m!��&�xcId��|kx��n[��g;�TԄ��l�����H2�.2
���|:�&�/|x\I�GֽE�gȔ��T搓��h��5��.������F���..e+�w7�r�mó_:?GC#�_�d3Q�k�أ.H���@P�-���"�y���$�����WJhpSYyp��Կ�g���\Z!ތ��J�,�s�X"]�8*\I �o�ԕ]��G�&��@������A�jZ��0zn�ԟWo/)����t�Y�ԕ)�Z�}P�����7 �&^�.��]�y�@�h ��\>l̲/@NR�,S�#� a��*��2�W��:� �t���� �>��9#�U�pɥQEn�䐉L�M��7�PH3ѵ�`�激�Q�����s��b�v�q���D�z�32��˗���qh�	�piJKE�]x��@o\5~u�]��Tj�K���|�9����F^ ���$�}4I�:9C �~jk�V?�=�\ߞ3���VOmaϫ�')0��F��΍����tk���j4��п��K9��`����N����7���]�BСoY)޹zf!԰�_��b�<�������?gˎ���If��TX�%�����@��p����3[��Zz��cA�!�˺N��Z]T��H�$|���|gϻDDj��ڹqz���\��cɣ��OD�i��� K װ�����ا��",TKs���]%"��uYB�c�1}���w:�ϭ?!�C��*��B��oi�ٻWՋ�p��ԉ}ۮ4#����Z̗�^!�3��h.��٥0쬱&�������^3���8��! ���MC�rz�ær��I�	�9��i�4�Q�s�GPUIG�����7|�#; h��R�k�u�B�9M�WGS*@�̚"���:��L�<~A۶ : e�~�;~�$qa� xiU�"R�����ѫA<rߊ4�ٳV�,r0jS.7�������e�D0�������J_�]��r�+�4!$�������,�[)CC����&�!����[Pc�����!�{̝#{!����Q�o�3�2�+c}�+"_-�h��4D�/.�������!�,~��,H�n���7!G�-K�+Y�E1��|����"D��(�ezd����DHӞ��E��ў��>@y��FE?L.&��V	1��D]O/U%��1C�����J�/VB���*�&$k����A��4�n@fY�m7^���2�����>�E	�"	�٩6\�+�=�� 鉨�tײr�ƺ���,������O?�U����ZD�$��iHb%90���x_�2��|�� O�-ۮ[���p��B*�ϖ�����S�g�'	�A�xԆ�t���쯯��4��ÌFK���Bu�0[����'�����3���OGHD[���E���tw�>4F������y��O]��hdu�������}H�7��O&��'���}�!o����Xp"
�������P�c�qa��ʏ�6Y��A���̰	�Re�'_��5�!B��5�nwβJ��k�.���]p^옔b���Mk:"�쥡�]j������-�m�YM��!������Ds~d�\��>�{8�����I���O��M�+3VB����;�g���/�煎OVF�B�y {5i�t�3ֿ^�.Kuq�M[4�t̱�����hMZT�/%\��Y�r���|A�h�����z�]eo�-&��dJwÅ���؛O~�k��-�:z�.%ѾcY�u�g���T�R��?��Yi6	�\���2v/�X�O�� l"��#l���9��cM#%V����F	��L���g8����Jx����A��$��-�)��R"�c����+����*��֋&�T��=j'"ė�j^�}�7��~�<�h2!�F���7tܞW|s���߀������{ߑz���K������F��v����5���|���U�K��ժq�x����|�� ��$���?��f�s44o �F��u"	ʨ����k�cyCq�?�c]���R��6eQhF�)d�zY�kwT���-��j@AM�v�Ë��U\Kyu�a��T���A$�Q`ʔ�85߃9g�W�}��6��1ͷk-��&���|@~\�I��ߨ�۪k�4y�c�V�[@|�4��\`���(Ȭn!},� Xd %�d2�a�Ao�4v�׼�E~�H����rZ��	}�|�O�'^���ܮU��Sk��_*�!�ڱPi�?�`��/��T��ߖ�5f�b���AR��O���&*!�����g�g�OB�/I�:�I��%�[��!Z\ Z��� ���ڸq��"�EN}纫:=M�G����DnLئdtQ��!<��	�dF ��z�Y�F�x/�Ǯ�}��!)�ٕ�T���2�v�={V�,J��2�A@L��q�K��\�����~i�2��=P&�&v�� W+�户g.�V�v�<�q���o[}��o��щ܇x(�	J�:S�v�_��)��j!�}G�dT�sf��ɝ��WPlfծG/��k�S$�'W���̊ŏ��p��I�Y}����*�V�=W��e�JXɋ�hˁ�sz���G�|c���k��ްv�!�-���%n�]��eo���[�I��j�k�/_��a�Z?������=���J2�=`!jFsb���Q|����t�u��~^\�����w)L�*=�#�	S|�1�UEGaa!�����lU�����[/�ߕ��گ�mC�˙H�?Y��:p>��z"��4j�}����3� a�H	�Y��Q��um*kΕ�FK:��.��x/YRϊ%��������k�-GY������㋁�������\���H��V��H#�rMw�vT��6:C��"~b��f��G��F��5����m��P|S�=9��_���3¸d�Qj!�++0ַ[շ��Q��{d�Z����´����'�+1��s.�
��s'�Ja�=A4�R)#ozy��Ps%-x$�凮ܼyt�A������<���z'���ݑ ��>��d<�ο�
�i=p[��S Z��0���ՍF����RY�N������_�����l�Ʃ`�����m1]��[3��\���n���aJ= �E ���:����Ee�%�f&����G���d0$Cߍ�ʛ�u��ظ���UX��G��J�f_�{y�-���\v�F��?�&�?;$���򖳴!����J��@�N\������
��!���J��j�t��f{J�XE"]��A}�x�����X��	>���Ao��8�h����W|4��ɉ2Y@ڵ�2]f��M<i�
>vaN{\b��MA�&��b�>p�GH������ ��s\<d;��g�k��M���Y��p+�Њ�����T7�j	[bΐͽ�G�LFB��-`����;#q�8�����װ
��G_\����&Ű,�L�yt�Z����k�_�$xvg9� �Y���'m�~YA@ktα�U�0���8#���ZmiE_+g���$d���e�T���?��򾸙��H"��m>��� ���M��~����N�8.��Ewκ���Y�EW�G�'˦�=6 ������ֱ=�1����~�,s�0����s�<�0C)�q���mң�a|��5������>�@�[#Xj���I�'���B����?@}EL���3�Ű�'ǉ8��O ��U`�b|C���@����6�&�N�e�nO��2�K݃m@��#�@����VОv��O��0��7\�e�������w����<��"ɃWЪ�jɩ	=F�wt ��+:������5	a���}r�ayU[pf� �c��)ﵦl���%T�	BP-�$x�;�)a`����U3�O�o���^8Wr!V]K��#�%��]��̳�J�mJ����^���F�ikk�x�hE����v��c���x� �%�v��`V��D$�L �P������$"a�M�'0�l(
<=������?��!:�	qj�â�o{gkY��k64�2;cp������8����=�Y��Ez~{%�Yj{�hU�����J���H`�;�zA����-L��b$m�ׂ^L����U�7聋k�L� �q�� D`/8�W͢HR���R��ۥ����q�u���#�U��@e\�.e?����0�Rz�!�d�����i�H'���+V��^�wfe?�M�z�b]#�#��`�M��9ϒx��7�����"gv@��(����؂�e���D���.� Q��M�SE��ͨX.q�($+θ��k�M���y��K]dܭ~�ڕ5~a�Ii-�����[�嫅���o��C���9Ⱥ���͸}d!�F:�pa��h�_�vE����s�W�56�e��B����R\�ӆO,�=	%����|ǻ�]�CE����u���,��)�	2A?�p�g����fTU\xcs��I�R��Á¤W�ѪsaUIW��Ő�I���x?�X�qjγ�M����~��$�yK|G��>��� �ՇPv�tG�ۧ�5_����������L�ܔ�>�B�TVPgVIt�ߍ����}j� Q�~�¥��VS��ĥ2�,�)�l�O���b�+>L�y9=�֋����a|Lf���g�r7U��G�>��5���\I@ڼ��4���z�n����-V.R�&=X��͢�3}�c����R��<߭k�3t<��A_�g�{�<��4��������`D���=�=�R�[l�),�������\ 0�����Q�����
��|��-�ͺ>�`v�!�,[uV|"�bs���v������Dy3ct�W򿫶����R�-T�X
 ���e�A��K�hk]Ѿ[�4u�K#z��s�%:G״1�M��j�w�9��&�h3̑e�K��4$<x�K
@M2XZ�!�?=z�,�Bg�~�`F�����X�cv�C��R�]e
������o�ϧ�78������&�Ԋ%� �a� ,��e"_��\�|�ϒ�+o�J�KY�~B���wW1���y5���zFQ��M�$i����û������/�������f<[w��b�66Ⱥ��҄
��Z�z��"!��a�A:Ds�?F6���q�1�(�9jC8_�T�@�$��be5��90�m�����jd)�*��l��K�����El2/�3����{fA՞��%C���=�*���	5����$��_pR����i�i� 69���L�zO�9���S���`��ג��$��`^��
�aK�.۹bN�x�dv��#-��j�dm��Z�m<%�/�2Ǔ̆�f2s!�S�'�9�YGX�ڣY�%l���tA!0��B�T�a-J�X;yf�������$��s�5A#��� >��;yi����%�
�T ����q�n�+���1q�a!DHSz�5M���͞$ܜ�OX��	�4���H�hǲ�fH�q��dxa��o�o���7�^)�o�eFRP��K�*�B�hf�� ��a��'$�1!)�Q�Z�%W��n������b��W�C�-�p���.=oT����Z�O���\7��ȟ�#����n�cmq3P.\�a�LY���M\�|�}�ǵe�U�ZH":9PR�$�Ғ�$��L���":M�����Ku`r�f��8��_?Ny�mM�xЄ �>���um��YK��A(�@d��'��y���n�T�c�s���2��owx�1u��w���FG�&�%�W���q1��hE��3x��4���	�&�q4�����KF0s_I���a�?�: �U�t�{�ׅ�m� ?���u�^8�.�z�J7����8�9��u�)� ��[��)a��U|�{]:�G%n�:9�x�L�w��*�3�İ�XǢ��ŋb=s���I2���?���W��a�	�~�6Y^M�5(�R�Mk��o��f�WP88x*Q��,=?��9>��7&���J@Ĳ]����w�L/u巀�ͩ����~��ޮt1�ghr#�FH���qދ�F�b)G@�N��S��W�h'�"@��ز�V���9rql�s6��\����$���w8����2�ϥ�H�~x���7n�;a�D����H�S��J�%�x�LFl�"l������H�1Ӵ�z�1%���}kD?��i��ك�q{�OOt��[>�qև��`Ӻ}�Eː��d����� pH��'��2h���o���+�~ԥs�p�.?A(*z�VkQ�]o�y��f�Gv�Ü7)��u7ޞ�;������]r�\A5�õ���gfS��3��V�+7m�9���;�,�4_���0l��jh!b^t��k�lWM��;9�uU�pB���s>�=>��F�%�����p1@�X�����ԥ)Ъ�SR�Ȁ�9�0MA�}���	uw�Χ[;̒(��ݣ�?��`����v��$/�����J�\J��ߚ�ǵ��@��#I&K��=%��>�P�Ԉ��-���v������j�V͙A�2��Ì+��9�Ӧ8A8r>C�yބ�j�Ƨ_B�yn��e!M���38=�u�]�r�D�KA3Q� &�F81�s%�6�|~���j�L�'N�����
�򾾻����G�z�T�F}��t�������u(�\6��ʖv-�W8���8�]<ȍ���S���qBb��Ϙ-����H�X�;%�7�� ��g���qn��-;H|�7�&����8��м���R��/<B�c$���W�w6g��4%�.�7��r����L؊��V]j�9�9��3xPǅ2q^p�^Tߏ�0��Ͷi�I2U>���vk��89$Ԙ�%י+fN��Tݪ
N��v"��]��X�zi414�	����.5创K�N�FL��q�z��4м�8~�QS�M]p�`���S���7�Y��R��1�t)�#�5���^kD}���\�"�@��z����
F��1��@�9�a�׾�{������j��c[U�lH�W�(Œ��͑�ɳ}/R�gl�5��=�?���R��r��m��8N�]�\�AjW_5EV a�<4�@����0;�{�N�	XrH�^�e8-YRT��%!���-ݰ^��R3��C��+"��!p��g���|����(��1tS����=*��䚀@Փi��B:�?0F�aB�����n/V{X��w�u�+�R%ңڛ0�����P�����a��k~p큡�)ţ(�z�/d ���T���Z���ō��$�d�ԹFqF^k=0H"-������w|Ě ���g�\�ViK�J��F��[�'��:c��)��NC��6�����<_e�K��5'{H4*f`�X��"���O�|�]��|���$?(����o`��Q��!I�4#��J��a��x*d�$��0���S�QX���z���c|t���4e�w�s~�%��$���A)h������KK6Q�zd�߭e�� ;�.�N+
�8��*Sd^�1b�(�����O�C��5�R/��x欱��y�D�[Y�f�I?��F��qOVb\�f�N ���^l{:{��:��b�{U��,�|�C`1aJ2�B�.P����0�<w���"�d��J��J4Oy�!	3�j�/�� ���|#Y?�Rj��
������S��"���_%��Eu� �VN�>��ukb�`��;D�-UG��OA�H�� ���8n&���Vmcn孲���u4� )CF�,�$ð$�����@��ʹO�����-�}) �8�PB���ۗoBw��Ո�j�M��3�_Tk�Ƈe�DHj����_���2/0����D􋪍���Ab��J�;�YI7���%����TΫ��~AY�"7��U�b޾���H	߬�^�����X^Dc�(s{�a�ִ{�kB|�nU � 6l�X��Z��S~��Aٍ�ȭn.��4���h� �g�Xh)��5���5D=AC9��@�����[�q��gG�ng����!JSch6���.U��S���Ͳ��pq�X�T>Z
`�"<)�����q��Z���On�K��|��aZ$}��P��s|TLl�"��+�W�4�\��4�_�(; c���ޏ&��h}'>왲������G!�Z�a,Mj��Nu�[�sG�K_qn�ܗ,Q�'��ۖ�q����� ����X^tZ"�����/%����RM��}5"��^'��s[�f�N�<�@f��7�׷�٤Z�������������h7��R0"���	�>E���f0	b8'~[��6��?�,��_j�PB/���c�O4�ts��du�����J�T��u�)�>�Oc�2"��p�9q\yEc����ߠ��B�Y�6)}��R�#R,�ǌ�ר��W�=x���̌n�E�ʰ�8���X�z�C�}s�>(����ds��A�XU8�� ՙO&?��z��B0h/v1�d����]����G��_-�`����"�X��vl�$qIO��������z�<�Ȁ��!iFEJ�Ȩm }N��thC-�H���m����i�y��%}����q���[���5��ڗ�e���A=V;XK[SPk��Y՛d� �tY��J�A�WSNaD�Y!��g-��
58k�W�UNq�����V���k��d��/��� M��}�Kڗ�L:^N�Su�.�:�9��[l/�J�Sz�i*:D��Dz���t���~�1pUw����BM����C��/4t����Dڸ�u����^���c�h�)
�s�g#���P7�#L*#P؜�DʵZ@�^�pI�A�?۟����)!tx���'ǀ������c?E*��h ��������ńxf!�f�-\�\���z6.8ՖXe]?���R� ���W��U�κ�g���>#U+O���C�!œ�
���vQ �;���8��߲�Q����ބc�'��d�&ko���ء���Hј�	�3���kINǺ��E��H��Щ�Pp�j[I��s�D���"X�%��"@k�'�B�X��wE�k�(}۾d��K�Qo^�g
�+)�ԕ	���4�l��!�(�����B��[�
�:�r n����Ƌ�yZwY4��z:X�����7n
~d��/J/�T%/7Ǻ�I�{,0h�G{F����B��e��<�(�[�$s�Y+l;)�G�F�VUHdJ����%U��rq�;ׂ�����'}ti~�l�	�����TEc������S�+H�]$qv�·ܬ��C���*V��6fl��T�`6�Prʶ������#8�!�|x�G�ќr�����ky��k�b�HlY��Ѱ�+P-)�֖J���;��ΎW�m�����xT�n� W9.cQ�i5��Uj#պ��L�8s},c����{�a�ID S?�2[�b��cx�U�^o\��.���C���9���?%n����ė�,��*�k�_�vS����Oq%8E���؎.ޠ�aR��k����
��"��Z�7	\�K��E�`�s�j'��nB�/�f����"��}��M�ǰt�[G�K�ɭOӁB�#�U1��m�,�\�g�M�7��%;��������/����<~������ʁ�n7[�3���!b<�0�l��.(������#���`��:�u��q�pt���Hb�pjU�5 >e��d������T}��s�f��4��qeU=}���a�c�xtZ�Bs(u���R��SX�6�8	�2T�yx�m��1<|�qzSnz$���79$�+`�a�]�o0,>�p�ۘ0J7�-���wZ�!v¶�4}�f*�M�B[���J�M�g�.�+S~��~��(�֏(<�e@�psT��E�q��d�	���%�tH]9C��b6�,�:)��#5MI�c����4��邪x|��/��	?E_+60�
�?Om{:!i������!������쬖�����t�h%77�\n+��O 4hҔ%��I��<���J�](Sټ�t��%���fP=�F'���\+��3��G�gY�����g�F��[X_ޤk�+����?���#/)l�(
Yz2����=��l���c��6�e�_���{���=#�	�v��7�z��3+h|+��f�">\Qv� �٤J��?B5O�X='�&�)�qN?�iÇ-�e�a^�N���H"�g�W�� ?�^�I�hM`�:��tZ�����XQo�Eͻ��Y����[h��758?�Ω�+�⢿	4XD���[�)=;`H���Yyu�u%�~�2_�T�>e���N����'���%�1��CʴY��XH ��朽fG��ߔ;��83�I���V�u-�G��aD�h�D��~l5T���#[��ojX������2��Q�Aa�3ԃ�xǄ�ok��f�H�CB�
�(p.Xhyu�B�m�I;f�;T��N���i�b�h�`�F�Y0��+�Z�ϰ�>@����93����M}�=�?�B���o�1�-C��䚱F�&Vȳ�3G!k��{%�O��!%�/�Y�	�BP��y���˓��B�~�Jn�x���]�N-w�����~��䚡a�n4ut%HeW�O�%��ٴ����?�����Y���K�w/K[�黴҃��p�&��G}��MF�k<;u���l3:=v�>Q��Ń!!�BZ��sXB�V�N���*OJ�o��MIiz��Ns���f�S�<f�!���8`-�RoxZ
AҸ�ة�mz������O%MR�{�G��#�T>�J\�9P�P�U���۫�գl�i�(��\T�#q��{01E�R^iAIB���ͪ��U!���F����[�|&�w�����Wߌ����	)*>�:m�$iK�/H��=
j8�>��T�Ý���
�İV	-�v�3��ni�ת����2��F"�t�>� �B�b�b���Wo�����6�#�֨/d�X]�gָ�ao܀�z�h\���-����n��5aF�����&��<2�Dl3(^Y~8�x�38�{DIv�JB�b�94&S�Zdd�d�D�]�X6�ux�����E�A5�k�';�i;��5҃G�����̳�P �}�\=���
@N<:�a�r�Ӌ�U��@�z�������!'������G��:`\��|L�@��Ya?��Ipz�TM:{V���-��,[.5������"�@�:	����N�C�U�͡�����ã���)d��2�3w��hf�0�`�&��fF��4Ԋ��։$C\:���FE���j�ju�*�(�6��?D%��_%������� �GY 3���H��2��'��X�	�K�]Ǖ���y��ЧI�Ç�����S<�7.v�a9Y7�-���-RZ�>������6L��))�\�YP��-�H�{f��@s��	�8�
ś�2����6Q��ӟ!�	RM4xD�/+�U!�wI��c7��!��M�|F=d�Q���G�S,U���H(���
f���I67�e�_���؍KV�+�f��f`u}���y�)�-p�9�0�XRJ8�;�Udd8cdVZv8PAr�c&��AZQ_� ������`;����{��dg	�'���jB4A5m�W���?��k�r�oH�S-�޹��3*ҹ���=tf�vE���M�ʁ��g�V�F)F�'�E<����?��T&S;�v-'ER��gv�Y��ꄲm�V�f�X�X�:��<A���3�A�NfI�6?=�e,2xᄄK�E^A.{�U���W�u�
�Ti��#c�镨�>|[��eN����Υt��	[E.�*��v/h
��T{1��P6:�^�Cd�ʑ���/S���U �E��_����#3��|Gc���	$y]ي�z�3%XliL���?��u��㨢6d��HC�H�\N��b+i��3��:��m}��z���'��6������'@���b{	�@�U��U�;6yu���|-"�e�4�yL4���kI�g��ӣ��ϲҽ#X|���<�Sic��*?�x8J�	(�o�
@Z��<�d�6A��7 ���~H�2�����&P��-���̦��oφg�wɉZ��n}-	�e�'�R�����_�'f�#�Q��z�n�56�G�%$����ީ
��.F�+�3�=�J/�j�;t���w�o��0����ܛ�2�s*�W���~%�	A�<����a�=�ƌ�#3Ԭ������[�m�*8\�>+�6�C�:غ��r�J�J��C�t�^��
�� �� �=%S"�����#,�A�v���B�f4���\�������.��_��=���,��S���5��ޫ�g8gk��6�0������cX�n��� ���iʼYk��=���чw���kڵ�N�V$���S^�k��K�����b*���P��e���b7��9�b>*�\�p�IM<F��+kF-ߓ8\I鴩��sxJҦ��� A�	Hmc�t�`)�4��Ql�����N\�!�J�C6�t�p&$ZWs����	���n�}�؊:3E�l%Ȯd�{�_*Vy^t��\eR�����1��ه#��(�|�^-�����q*�!\�jA/N'���O�z���i�㒲GDk*��N����Yk�?�)�wދ���˫��brm�¾����)s�i8}+�5������h�VJ�㭧Xu�ц\7��"��u���8��G��Y��j�E��\܎�l���,�=�+Ɩ� ��IL褰+X�����a��ƽD��:��x�������~�G0�I���,�0N�������?��o�e�>�S�^ʫ�&�� )u������=X�N�5��tR��ɿ� ��U�������y�d�^V�m2A?���Qh{ɘ�*�N%��)�N��^��\X���&��f%�u1�Lb&�OXI��������]{�n����f a�n,����=���<��6��P�6�}�[���Yf���_Ka`�� ����`8o�ه�|4A^���j^�Ł�ݲ��Hd�q�M�C�Z����qa��U)�G�8v���R�U$z��
qg����g`��n#�i ��H��Jx���^�]��w�0����B�@��b��7M����d��_"{X�\p.MLdZ<�&i"Y�}��F
���5u�������	QK0��I����p0qU��Y�y$��Yb*8(t�dN�5�N/Z��FQrøjZ��@�"��r36t*��F�����n��@�R��#������;��X�gԖ�.�J����,#��@T����,���C���
�E@`�iW� %SG���3��:b@l$ֱ���
� ����3�� �g�N��R���R�C��i9
gE�Im�'���ǮR�V?�S#����E?��>�K�k��hq$�$���&! ra�+D^(,x�EL�jϮ����d���1.��}�G0��{^��Z�@��/��̥�{�L̂�<����3��r�ڸ���+�5#��m���sy?�+�z��0���)�������A���ml.��JW�o�7��Mn���	Ԡ$�ˢ�)�~�8���3��-���$W���'�]���k'\�H��POHk�ؿ����C�)��4@�p��f�.=�븂|�u1iW����/cD 36޴��h8�G�s<i+ʡK[��|Ρ	���nְ�/���Y�EГE?��8���G��rJW�#�t�+%b2Eƿs���K�qgvKٛ�����|��y������}�*Yc������K�H��� >'��6�UP^$Q
��4�O3��T�W��	���u9Ҹ���y]"�J�B���^��c�O�^��h���3'RQb;�N�%����fiT��~�Q� �x�l���Y�Dq)	1#���6��R`޼��R������W3�v�1�ڦ�AZj�Yk��{xJ��݇*�Ēεyj���*�����:⤏��No-d|Easa��i�-��v�tҧ�m�Y��Ʉ�tk���V~{`&��D�#�Bcgh�+�v�.���K<���x����+�8�i��D,րPg�Xnm3?_���`���j�`�{dI�� �܂��lMh�O��zž�L����߂���w% �s$��.�f����J�B3��hP�C���ܝ�n�� G�
eg1����ED�������:����]7t
e�E��S�ew`�R����'�>�WD�eC�"<mX6���At2�*6��9&u���	2c:��������G�}��HR��V��U�"+~3��˨��R�<Ę�J�ؕm�$���ؽ;��� k��2����"����U��ۊ�l�P��U���(���z9�<��Y��\g��Ap��9����H\��eE.�2��X��ט"����N>�^�������,��:r#zR�����������S�G��kQރe=j�7|�-C?L1�ۗ���d�w�3�pVX'zl��]PDA8�;�ػ="q��=����C̺���m����Nځ��(��X��z[��}?I��A1�ꗿ����]h�O?SI�vT�j��j\�����%l�TaP}jnC�������/)�W	�}���5�O����x����
�ʚ e��M��l��\�{贯�T'5��H������z"���b�ǇI��.^'�Bc���i�'���P���_	��;#S�����(��]����!�R�3׌o��N����m�O�!k�-�!�0(r�0�ɥ�*c��1��]h�L	D?�u�Rۂ�`�p��xZ�sKQ�]OYK��s��}*_�R��ITt(]�(VC� rJI�pA�$x��$��^\�O�c�6t<0���~����jG����Ry��� �9��edc�$������X��,f�ιs-��h*���-���q�*I�	SA� }���J�sцϒ��������*��aZ��3�����D7�ZA�<[��QGr��-]ߐ�ȟ�_�hTJ���:5 ?�c<ׇf7:U�d��J/ht\��-Fph�6R֌�!����7��R��*��V��+ʕ�Hmo�I���d��s�$��J��w���i�Q��,Q���?T6��u�E<��lR�B �w��g��F/�Wn&h12�ia�l��0jUZ��{��a�@������۵�ܴ������ً�K��������K����J�3 ��^h�/�א�
G�3Cnb�A0K��S8���r�φ����ݼ@�h ����y*C���W���'w9?�k>��LH�|�Pٙ(5��z�н�X��L�R��a�?
Bďj����X�qL��9��	7�����3���ê6?�nq:���;^=�>yL�� ZÓ��7P��3`��Y��������Pp_���Ұ���hR0\�?q�����@N�P�(����0�F�>�F�������ih7��p���7�x�'E�Z�G~P?ڜ)�����F� }�
�l!��c�I����{