��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�@V����B?:S���/��݀:6{�#rY����z���	N[��ѲA��rQ��H�I�-f�.s6��`��zv=QȔQ�}�?��O}��h��)���wV�ϲ�6h��-t&|0�x9�:���0�T��C�,K���5�$����|���nW:� #���p&x�/��
T,��Ɏ������2戹�M���lv{������r��:%���,�[`��^����,b��*�J�_m��/�p�/�б�ɍ>���4��+n�������*2}����wn@
��]z��@�:�HG�%�>$��L"a���T���'�|J��4SI�A�[oP����;f��)>�T�9R�y�8��O�T�S���g���LҬ<���G����;��V~�܅����R3�qO��M���w�ɻ�����U�]+kjLzɽ�	�M��Kw�"�-�Q����ob�4�+F�Q�/���7���^-!�ōI���4�l�*Ȧ0-��3�!΃_K�[q�;�mAwP&��=��֜�U��s� d8�/�R�L��B5�󳲏}�S�Z-0\�����q�k�K��6�����ȷ ~�&�ӝ����9F0����C?�%��<�{��z���׹A��%v.?��1�5+�K��������-��F	�S�<�0eG�cC�^C·G�
h�:����}Bc7��O������)9���{��c�5'_����+3-O�KTG=�@�J�Hi�˹j�`��H�2U�c��?ڠO�[%,�]�C��p��5��%:�(em�t�;�[�^�w���v�l��,�u	N}����Xw#<�~4S�n}��,IǄ�3���OjF��~Bte�A&5p�ٯH�lM�e]N/������or�$F�������2bz��Ş��+y-�d���;ȥr.���� �
�A.���/T-R���Cx�Y������-u�g�O�3;��!�g�y��zE���^g'���x���C(9 ���B�=�%�G��� ��� /�v|�:���3[�=����>u���̅�x��{�	
m@�K���<�1.}�U�X���L�]D���_��"US���M2ZЁFb\D�k�s\ܲQ�AP|�#�RVA�"|;�!�B,���>��"v������ �ʊ~��Q����<bp΅�Gi��~,ߦ��[$_�B�*�o�//�؂��A�Q!Tó�/؝�L w", ^�&�k�� ���ǩ���	�IrT��L�fl� �����`�Z����]��vz�9�T.�!�Z�Tr�Ɣ�R������~�#}�=m��m�j�l00�A����!3ܕ����fJ=�4��:�a��q4 H��;Q�^��f���j4'
iw*��``�����f��/��w�y=��BI��m��zðl��<�� H��ñꕏ�7�������s��>Ν������GY�ա|�|���:�?b)���(����4����5����c�sLO�3��0<��9:���kݛͱ}���_g�L�b�y]��c:4�Eq��A��� ��M�42_
��7�en*[���F�5$m�&((G����\3��N�$O�˰����r���k��#��r��p	4q˅:�9���m�Z�k��2�N7u@[�d��r]�n"�#�s�(l�K�vɽƖ�A��p7!����xh�П���E���8���[�2h�v��!�-�,LPt�*�Wr�dD@g@�}z����ɻ��7_{7;�6i�n7�y!-�ߞ��.���~�I�Y\s�B���& � �B"CN~UW`y�1NqM�la��(ʰ�7hI8��s��7���b@�m>���4�(� *@Nܗ��
{'�U�4�M*���Ȳ�m��� '�"u�B���0Pq&f|h��贿S��}����s^�'Aխ~UӉܐ��[`�7ѬS3]�E�j���@/_ �}<	�d��� ��T��!f�Ҏ!~dZ���
:XԄ^�Kh"_�L�kf�JI��EUO7)�bc�d�[\��KVӢXa�h�v���m*�e4���k
a�&�A~��w��$�7�e����;��ж#�q"'������"v
�{ey�y��V��tC/��'�[g=G��%H?��,�*+�5��	
�H�|L�`#��	f"�KP�����c5;�S[b/��)J�ږL�����'��{��}1@��=3�\�F����$5D�;y�
��<^l�pGAe=�
��?Iʃ�d�����As�O{86��i��E����g��:��MEf7�v��r?:)Q���=��ÌS(]�~���3�X�]v� r�$o����bUʍr:^�������lY]h����g�6)XjV`��S��Q����7��;�"/���O@���
K0�KG��M�1�_�=F`��L/W�\�68��]cM%_��
����K�����HU�<�������V���HS�¢��H�P���)ם��O:)m����lG���k}(PV�IJ����8Ӎ�~�vg��.��+o9�)����y5�q�0J�f��ww�G@E�|hJz�,��j�����צ�)�K�(���)�Y����A��PF�J+#�##�b�� ��~��uؓ�K��JK�����)�2���
�i��\}�����q�@�Gk�䐴���WC��S��PH*��4כ/p*���$�:�#�C��T��3�Ë�ݝ-�D��}3��1ep�ٙg�5�1#�:�B���M;�xɧ�7��2���.§�s!�tA�P��?����免m�T��!�]�]�L�!丱�U&ͪ�Ǩo� f�w�ztw�����Mh�tWX=�R�n�k� [�4�kG>��M��7�����Ÿ�Y�!sx�J �B�=�9�{U���<�ؚ����m\-l�ѫ�C�c������Q�a䝼��f��������k+�~�	̬��Ӌ���RǤV3 ���<dx�L��+S3>�/NpR����G�Jљ�R�|��������*d^\6��V��.����$�Ԙ�u�&�X�Z�,��N��×�7jo�9 ��- 9�5�qY�T�C���aѩs�j�Ѹ#F����lzd�iW��,c��[�J�Ѱ������>�b����Q"pl.:@4#qfKLN�
�Lx��L��Ȼ�JV`����qNr��?s�Awy����qB$^/���1�`Kk #;�~h+Ǯn��[���x�:��SS&2VQU�]��U2��r\b�Gl�.����6��1�Ӏ=#'��d��ps��MnĦ� ��r h�	�ާ
���Y������Z�{�U��V�W6�ѡ?�*���92�<��.��D��C�4���2z�vv�c���bq#ۻ�bv�1�ţ��b�D��^��xL�h��"8�@�<SF��8P�z*9���¹l��"�?�����%)�0$c�����e~�������</�8�[dL�@�s1~t������"ť@H�KM0�3�`�C�d=ۗ�N]��"`�(�u�Jo��/�kk;�&����s�ô7������kPɇ��P��X.��4`����`�����&�cDD�8�W����a�V����z;�� ��`��g��|�jE��*ä6\��6"���e��4V�9�������pB��R�5ua%�hn����BPS�y�_�v�";��5+��e��OP�N�%w?<:L�q;L��c1,����Mϔ��NE��k���L=�L�vC�B[�Ͼ��Q����
C�l`��-3E^�A�M��%��{bG�T�δ���q���1�c���`��vL��e:�4�����u��������2{��g�̀�����gZ�q�Sc����0SI%8��M|
��.!��&�Q�*�v� Nh���ז:yq�)��x��{"c�fx, �"��ۋwq��JgL+]͕Td�f����t*|�#8���;h�cU|��@t�p,��-�Jq������I�9Sb�߳�tf�(�]�;���/^�$`B\�'*�8lPd9�BM3V�l���Tz�)�-�1U�hGy�"e���L��U(��G1~��{��T�n�j��� ��|-���Cb�8w}T�%���wtRX����Z��>�X�p��~/x������e9�
P\u��/�{��4 N��4�u�۾5�n�j��\[˥�u��4���|b�Z=w�U�־%�^���<MW0�c�%q=�줸��Df}���Uu�!���c�]p�z�ހ�|�Wt���^����~�ʀa�%h�[P''�$��V�����	ND��A���vu-{���sK���	��e�y��g����n<�ӷ�!����Vf L7a.b�ϐ���;��]C���ݙ����m����CAC~�q�_h��O�<u������ޓ��}O�cjΣ���~mWe�Q�w6�Ha�ܧ��)j�S�P��=t��J�VdI�>6�W�ތ�c�|\�s�=rlBO�Q�t�8�������䡗,�_t��/ ���3���-�����L8��386�p	!�Ӭ�փ:�Q�e�JM�n��[���~>~��9��}У�����
=��
3P�X-��5��z����ׯ.�7��5z��Fp��,g��b���R f_j�d3�6Y������V��X�a3�|��g$E���M?V��s2�[*5,�X}<sׂ5�df?���GH]���`2pq������Bx������ˡ	fm=[���~5sd�3��PL�6�hD�;TG,��D���N����̊!z�`�"�����b|T�+	�m�E�.{�aN5��F
_�@?�(�C����{��;��+8�����0�;���V�<PC�l���HTz��6����e,�?Y���W~ZYx����# �ZG�[�,��t�_uel	���$K��{@��gX�AY8�UMB��m0F}�.͗����Q�h#~�����j:�؎ʇ�3R�p�5����)_)%q�̟����O���@Z��X'�B�H,��dN�/�m�q{��k>�ː�6]+b)c� �bz�����
-UFPa=��8 ��~�*���yT0��Q���㰂������y���Ϸ}	i�Q�A��,��N3�e��ޘ-*�ܹ>t_K�`s�u\Z�ǥ�&aJ�l>b�۶�L�R{͹9�����-��o�N�l��B��9wX�;�K�o�����A&b�c�OYA Y�\f��������8��ꕎ�!��;�n�0� {r���y