// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H5zOyy9NKxs+tpt+v7/r8wMe73SbpUIe79mJF/I5u9OwycViCWi1wUgmxCKL3iKI
KBw8nV05PcdAa4vYDTHcg4YixP0dkqJLc87a6umtOrLUG5zGYupsnrl+MSzy7WzK
/uSelvB7IOPJcpMb9y5v330x1Cg2LFupo/OncL0AcsQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 51232)
gbp+wHzyv9zPV4kt5PNgd2pX012yEtpQxFn6X4PbogpimWJhsypJgrxrRvgoGwdl
v76AHQRHkk9driftp3EfaPAnwIDjzEaNX6WVxrghFJHb7gchAhW9knw8ijy2dII1
ogk/SuivmptecsPQ8+BRzIYVysbyJA1zuzYYhDprm9ohmANMqO/EVFPqFBAe+1zK
wppiSaXJ0FqMLF7Cqbc+ODKUkDfppSGTNvNyqJkiC6P7/yboW/TswHB5GQec/uo8
CykcBIDn27InoBlDWwLIt8H8Y5XcweiK6bs7CnGKhlUUseX1KvCLOiF3pPKUUS+x
dWaaO4Nz20YsNxboixFxxboiQW5ikY2cmUMfl6FTX3r/0jMCUlpWHqszRzN9B4Cg
PVtEuCxHGC+8FN/uMwqn8QtfKgkcfMgMzKPUfwHNskpUZz3yLCivI+DxIVQMGvT/
u9uTMtBnFdsD23RRpPJO9F4xKaRAt81W7lWD7tVlstLc4stSbUaC4AJZzXC+hPym
CtGRXybKNF0wKqM1I6VR8CTt9tJkXypBhYP2kKc3dImMdTD7sg7ti0JqlCqllXTQ
7VJ9Q+TWlWZzVojGfe7aVvTlcUatdMVQ1Pm4gAAfeT0zj7OH8ehPoAdGPJo7HLRW
F3xvehJlu3o+i+qaC24ZxM2ALWEE7BSDM1lZDVQOHyvWfkd85QQMoEyKzHZeFHys
qYhLsiIwxYYjK8x3RmcFSVXpKRjVRiVtc3NdwCL5OkWNkOqBFp9OmcWzB1nq4KnH
mzRufAlup26TB9ibUhVupavfvFd4uSv8gg1j1DUSmSY7RR1719WyyrhceCdK6NK5
Z2YL0mfSx/ctvyxiaP9Z38pUee0LcptCSqOn3GhXXtoQoKzOcThj0qhRk617+eA3
kzaZM3CFsSVfM53LWAVLnUNEuYGwt5RJ8y1CZxkyiU+UzaQTjZe3tt3ctRSUVedx
+ZwbzKlDhZrgqwF1+9nQu+RNbHgpKyGceOydaDCZ3BRT+t82AtLUfPITmdX4iD96
1VLaS8rAKrkdxsuAgRokIrvmzk6F1AuFtCzAyyKVwUYF8rcr2fJ2RkbwOAxQ6ZfP
BFF+0es2jqslrJ5Px3PWqqrHk5MH9nOrdR4ovkXzNrj4QZYKdO2mt3WTlk0V1cto
SH0zcIqNPwogjzwLR6Za4k1tJgqrQL5DS6CcDxfe77gOOHCs494hKGZ8FKOy/zXe
Ll3M1bKuEC/gp0MlS94UKxvBX/mAKwfecyrUz4FH/JNMKMJia2KExIBfFFVOR6B/
0Kze9fM4bRELM93vy9Z4yKn1QG1dVv2pPie95fa3BpmbejVf3TvG3CBofsNqdVPg
OQ8XsAvUKhPyAh4SO3kfkFf7AmC1jre38zuEsT5YFo6yu8tX07hc9fJoEWZKw+7r
7lt7Ob1rvpOO0fPJW9s4/ZfOFDtdPhYVMkfAaBh5eT56d6UVUvEOmu21uEEFrmRw
awvTvGeW67z0+4G29M0xi5pmrSkoPlG8Fn2grRrF3IY0ODAcalqhEamKN3QKh7x9
qT+c2u/tni/dxRtznKkZNKtbZuJIO8MP3u+THgzeAf76rxbABy5lrFNvlwpXg4Ph
KD0m7qWVTjj4z4a1dHEJUsXqcPVZRG4TTCy2SHyTb3/dRCumCeIB5VX2VWZ9w+mv
RRye4HFV4Ykzrt+PQ9i7s3wQJrV9sAkxoJKUtHO6Oe2qE6ktjkgRnDNizvYCirqZ
iiSemHPov7sot63uD6fWFlzOvoWAxY+lYfD9b3aReYEFuVY6SqqklLedwFM5amGa
ZNFpdoM1GvXsMQE0AcfRvjZLsxdGl9oGFAk/3T8VLWbjWHceLE0x8NM2bu91gPMq
cyx37UlUSDaF4g1/0lnzZRsaRDlwh+fkds+k19fjLSJZHZtXHxHzpajAuHzZ3PY5
zWDUiqhWJZKtVRYbEnb/36EJG0OA7Rl2nOAORbNM/GAQqfxkkl3kzWV6swi06WM9
ZFxGQlh3sZiCR9dvK8KTSq/nr8ifVzfOztazlh0Jd/vAEqKSjC78oAb9xXelgc6x
oHtozBEnlgtGXDGXJHbfIZCfkKSkeqi/5SP8nQ8NFeV2uz7P7ScNxYB5Dx0TSRD2
hqkm+orqErI03vBU3Jg7oiHY/eO0yAVEEwPHCRkkwHHTl/W92Jd75QyCpHc8WK5X
tLJbBSTU8JrB907IH4LUKh88Irj0fTAvBtMZBdF14ak97fuFgsLZvNjy7u8lPDNp
ZpS+PUSShoBNQDM257PaxtTQ5AX4lWBigDdGyBtNGESL52Y5eeO1iM6h851+x1tF
lKzJtoO8MFLg0R9i4kkhdafqs7zaUURCBc79CZ1pPmuYsBpUosxcw3R5ypYPKQ51
FP0F0bPRE/9442UII4jckriE6VBCvnciUyQqgRo4dD61tcQw7BEX7zfezQZUF6Y7
4uge2vTYLvOJSaANKckvjBqG+UAxfRpgS6FbAZ4P8Du/ts9cH9D3mSMyC06bzP7K
U6KgTbbdDHFc1KGQUPhu1JwgNQZ/Q07YmT7ZxAzS7M11l7hPZ66goHuhX89CI4HS
HpNi/ZihuPMl2XVGRGQwv4d24wXMdJAInzA0lqAXUryfia9juqEj777886kUcfpS
9NvIDN8aYPjy9SZvFDKQmKS8XT1h8T4YXrivLcDI4CXIKZF+wRXGHv1TUCxioSIy
OrzZbyxouFcZoFt4iPzBwTZ/zjsaulCCz9xp1pn2JcdrV1lil0BJvgvRmc24d7fA
nIePW2RB4LW3RmBkltkiXPs67xjspXLuO/rN53zHdGsud9c/ywgap4OAYgLGWZFT
eDJXSEDE0Kzr62I2mQNnyVhe3RZ/QmDOHIMrgVcwIPNJXEPfvpw29sAm/fgRJWFq
sR4sie53RZfAMymg/AtIxtnEMqR5y8x7X9ehL7gt7NZ/g0R/Ef5WkjiUmq0252us
cNw/wvKedGXDUsbLLSmu4Q6t80L51QelxP3eM/qBl03PfxOEUysEuaHIyanwXIC1
XVnvw0BkOS7AxENFE7hct0C9Pem3vnuP3vrtKB7ctle7lwRNAibY/vFmp7XOARGK
bPNGP79dwylFRwDEVki2TXyCp5ERQyQF9QVlPHwvQvIWZLKh2NE0OC8/Q99K81dM
FtVI5SVVzob3z3Wxj/TpDJ4hb7ZQqcVXK/gpR+qqh3gsKbN7QeFk12B9q9nBLY58
1uPGvvrS1jSfAySBuX0tqLuWnLUt73xOMe76bTJEDnoJQC0ZGo+LWIAZ4fwcNf64
wvHEtSqVgusMMQpLnWgjPNetiPZJ0x05w6vPSGGBwbFKhSok7gXgGxC+vfIOcCRL
e0nGkcZkBHqbK/PWj4vAjAeCnOeI2loCGLYb+y+QRkT/X8IhrKuI2Ir4cV8ufsO4
xIHTQMq6YqLELpRrb2aVcaN8/Mr0xfkaMX/SQZ5LMbc2BwepxA1Mb5aAk9G8kksa
enYi1eg52YvG9N6sEduCQBE0rydAAmD0JPJ88v0sXp4ytDTZh1Wd/8Lb6xBIwt8m
oA57JxNYGe9r6HXfIdqA+WJJyGtwRG5jZCJg465egM+sGcBy/WXB3iHGCLg4ipqk
AXYWeL8Hz3/bQ7/xDft7EzcOtDKpS0eKpbX6A2+l+gAiENkkDWrn6aDfkcuKQa7B
3YhyvM5SH/Gh/FpIiXvSr0e6H9LVsgWC5PyqnKGNnpFhXQux+vpkct3ojba7VBd+
39no35lXDTgshO26aH5rOtV71m01IwP4PODiwtKqCd3theR1fegGM8iyd0RxHwMS
yiC876/fkHzM3/xHgzaMseJ2nHuVWDzBmgMLd2DTj+uhm7eJ7nkcbU1o0vM85d8U
Qli4+nQJUEWXjhWKYvcXPnjUT1fNYl9Bku/LVQsaH0xhXDPCdUA45PSZq/E7Dd2I
NY6PXbUzNFXBJbRkCFI0WGlyR1z9jzSEJFqc8RlpiinfLF971ERMIsI4JHn+b9t+
kTl708Lq8njttAp2HLgfXTgsyUvSAbnOVDFvQSXcKSGNCBcqfOMBs5CgKjkYVhnk
3pbRl0NTHnoUgns3ILjBvk3Bx28HxoX7zV/rl1z0adre0oJoNtdiocrpNGLqtpkg
fRoDmcLal7nmAc33JXNFHFt+VQbGLyL3kBXK9SZOTI13gw56FLBCdxR1ZsDHqYFB
MtGixzdnBKKpmCH2oz4HMRBsGv6WvznlWblme7eB7UBN4mzvz9/AHr93V4Q4phqk
YvRGgq76yTjpTXSjTImVKIAnCWfDJlb7QoaqG5/7V/+m8xHIhx9faLD+ep2cuIEI
ubCpVZ6z5SoaDQE3/DnNq1BjvoWwvVNs76DkXIAN+AFqOpChGLM3O0GT1UYinyWw
/A3TBCKE9tAKgjttn8sYfdQVaqyhRBWy9pYdXWO/jv3JoHoa+UlSyUp/cmOlEkgM
Xw/7SSCUSm/e4wkf2921ONlPUil+aIgr0nvzPpJPi/aEC5BQG9dB9B33rDkihOH/
6PLl2DQkpHLsqYOPY6JnF/WtDWxiJ5RBxyDcl+zxxZfQ70Y7jaYvhlXtUYmH5y3K
7SrRHLr0fALEF79yWe+LhP4xCINI3V5NJKxFZwUgdA4ESVNyfl9m/PeL6+H+baS3
QKAyTZp3GBTPUenf58RNy+hXKXTUh15FuoxlM6+NzVHcvAhZ0oXWilrAseto0op4
p2K9WHMGM4U3A9QjWdShwxtzBb9JdC1hGp5vNMLUMjRFUDhUkc3MWufJVxqaQtuj
IZldek0m+/S2PN46pgLTfYmye6tdpRmGgA+olV9IWpBiIIu+/l16IQkV2v0Qg2VQ
k9wYA2qCNg/P3DCcRom+iW5V3kKwdvsOAiPDn4n6Hr3jCa4/1mNTa15s9fiTL1M4
SiKQZ74cZuFObj4xcgBCov44+2J2O2czkDQlJud1VjYT3POv/OYSI55WkY0KkSKq
il8pczyRY+AWOD+aMOIOPOpuF+zCfSPzx53XFap6swXblda0xGlvHONcZEI/4Hoy
NTFWAVOj2rg7bb6Z2IjntrujtHZBSBQTp+LAFCqq+f8Kl51zEQ0jLZKai21FaW7V
V0K5ExJ6CSBVTwvJaSfsuxlqkxLxBsFAj+QjOet2QGt+86GatDr5ysMIrZ4UIq6o
BtzrXeNUPTUUH/TgG2WkiVlaRJUPP1iR+g8W8Bg5fuH2xwDLx3V+LSpmmHnr5FrO
Mnz6ro1z4L0VsRFlaX9AU+sJpj88loH/YvTVOLPppGoRSxJU1HHV7xfwkLfxIwYU
pyAMIWA5eYcatfI7rYquzV7h8bmhETh/2rWIzlRg9mjg9F6ZvhmGmI3J1ao0m5Xq
itA0xEXezY5GhbX82G0e9OVVEVgQeCnyqMMi80dfzux2FvXYtO4nENFtpzG3FRRk
tTqNcOIxiQH6iuJCpfBSHaNAgR2KGBDEQhMnu1IiE9QGnDobyDTk6uDFFWiXocwl
H36sZP9VJLTajuu3tNfR7N5W/B0W4s88KU4vzleNKcMm3EEYuGmA/a7btZsycyho
UxEfNupACnon7BmEz9V9P34X7AABj2937G+dDrqTU1WkL4ZXf4wDOL6mdxkF5Aoj
qoJ+pAWd++LSbgxWVc+v3LZzc/erIk5FNY9CA73ubD8fABFd903qyjLYcoCn7wKJ
z1h3QujNgVw0UOIjibyj1+IA0RTjYeP6QtxMIEkjD4c4IrqtuGNLIm9tpKsE8gN3
n17EqP0IfiXN1gHIUnRk2TJpKRNEoXfjtDYHDvbD21BgkIHCExzEuYlXTwyoLi9O
6NdheS/+E7PXoxm9drfavRK5edcRcONYQRrTlaSGORaQN21wLiz2KG/8yHdLxoQR
NTXF5XhCUwPeoVpj4vjlKBAHcegkhNFX8ZfQ9qvpFkZc+Os/QjIfShWMEPJ8bzFo
9fqU09emF3AG3DiTtudlzigfM10xXQEtas656wYZywca8SqolOE+mQxecEqK0B1b
nu/nkI9U4dlhK93ldOzDkwQkyhU1TTapDaXFTnwqISiXHCZdDFwJ+DOQXEnZk9yh
yDHWbWuzhroyuSr9YBTd1U0N76CoHAjUe3fUeOtn6AZhUNrfJ966dRUkIZnM/tB7
XrEICWTngLmmba47z1QVre6MNqh4j7R+1BcwN6wuJGVz7f9gmtynvmvyOMU35RYj
5GCYq9dwBN4+WGAWDYUvAsc/iDleeOo3E/Z7q4T4IBrV/1v5WxXWFwO9qrdMYNR9
HDJgI9OP3DeOv8Ljhz78uNKFMMpkB0vCXatVTMAt2mBmCUFAZg4Z1gEPjbrJBxKb
aEP9F4mB+C5vZLa3AWDLeW/jf8rBvjd0lwnSPqsa7qCaxTcw9rfqLTwMGOfmSrxE
06stqkLSkqafuKQLIYD3IlHAd4f2bfwZzzr+zUynXtRvz5PkPgrlX8ehwQXMWiLE
UXv4/MfLiNvf3qoDsd9M5lvVkvhVllwBWoGeefp1j/W5Ntw+dWGfIOgfW/pbEGCm
EkSNWPZnYcpvcBSeYD8AKuR7DHOJnJWgrRaYaK8SDmwlsQjrkoWz1TJNnKJSyEBs
8MoKM3WaSdLUOHrlbTPIKxRuvI965EQmZ4Fxfx4Lv+7K7N7YTRDUgsOU75lELKoG
bS3ZwN7V6Lj6F7quWYCeUX98rGGtY3YLUu+G3LxRiJ2RMtIwC5t4hXpgQwOirbjy
xoxbPZWvQfdH61ZMXSI5cL0pkzFn0833LMr/Jz5Ky1ePMGI9lbpPUvkQZ2cV9QiV
Uzrw+KlRgNxHsLNx3rTfgzyLI2gsI8yinIEpIXnT48N/DuKuyXPcyyViBIjRR58f
R1qX+ZGPDwdPMtOf3m7elXW7dGR46zWDMYXIe4KlKE10jPpR/Ua9K4sHLomYvRfD
aYAf0jcHC5IkyO210knUuEFdDyeFZFD+n0bm3HrQ1TQtdNVLVZLW8Q1M7hLjM2IZ
6hMObw0VKOoDKgtqKjFYXYrghU0vtwlCLh6cd+NRlTZJF5SQ69PfA9D4dpfOpkl1
MKAbkDbR1KdgskGMNqzp+OSAflRINXxFoD+CUKpxo8e6Hocmrlgruvu5Gmmva3qI
Kp0HLed+Pk+Jht0aj95SCR3/CwyRk41VSYwUgY92geghXsb6NOQvqJy5clgIuyyG
df4bfjK+2JqxoVBk5WLRlosjDfaXzWBEHwpu3iR6DYUq+b7UuPEHa0tpQy0zA0rg
XdgwCL+VQ5mNLqfDTrRp6C577td5V2uzIRxue9JnyhKVZem2sVKteusbeQXCd3OD
6DkljTBGFvNLpLzdQZaBpM6SLTMMO5fK6ruV8EGA/D5mQBQRy8SkRiHb68RHeDHD
B9ul6Eji+ue3vxPF3RhhPhrWe/XU6QPxnClrB1ptD3ge+kVJDRqXvEoerZWMXlcs
aaY5EuGDgyjEEns9GFCr27fVqf2gMLgcJyDz/OuAHEYD0B/5mf+hgvFF/4YJEJ33
hjJlvgBSx+hVlJ1/l5q205/AVbw4Fi8yOMED0DeXbKlcpV4c/KCjuT5FmIeUJii+
/5xQaNulTJZnqB2ZkHtTzS5JDXKR8fl2N6xjwaEyzTzWEV4d1rEnzZns7YyupZ10
GnkH1FLD+NMt5B2fm9PFRkotKntLDdGVaPAe7N0WI1k1PVuBwW/MEwM9vtLCs+hz
J9rzkQLsE/8dKXIj7EuwO0grRVcq9Zi0TAcRG/rYZMOGlOT0+5fQjoRe8fqvcuKL
Rfr2sNGGln/HbIqKNUqL1eYj3ekH0BWvqUDhawtxR3AhoGrzuguUXsuOlPwFzeWm
eHiDUDzw29+u42318lBjdYii0AQFp7oH8Vqpu1Tr6uhy30UX19+gvjPiPy4rOEER
0b6ca2Q4F26WFZLHmwWvU2+TGjsFjexyXdygDnEB0z9oiembbm376xEdiF6pXy8F
8UaB/rS4xXDytIXYxq1KF0kW+V8DsyYxm6VdXmA6+Zk0fJJ22dXNvmqSkJvBcYHD
LexIHQY++8yyaZAL0eiCv1xFFABDUMWUfr3nUN7U/JXontbaKnJ/JtqUv7TDUmlx
MG7h9WQpL2J331PaD/LAn4AUlGnzCiCEkeZ4ueYZ8EyM7v/BhjwIKCPi4MZL6lKQ
r6GPgqSBM6RtrQld6yaPmHa86MafuxyYY1UU+k4HVbtZNGuaohgPfA/8p2vot3F2
DCwXJKbf9UQvOxPHUTKDPxznhCQuvzdT3/NbyAVmPLruzDEs1obq6CIJ40EyNFqv
Udk1hJ9zVZnNvYNR6oqJYf21D1LsBFtQy/EKSO1jIceMFOu3jHqYsl+UBBTB9dc1
xKPhKn+tnf9OyD8VAR95pB1Ehdh0BPeoE5uOmBTFsen5l3O0VBbk5ZDUX7nefcA1
S8PggCPfJvgiu6Y8D/ojk0vzAmsJS6RaLyu+WXvhXYft2HD6WVRZwSJG17NZ5RW4
iTsLxpB7AWH6/7pLoGhDdM3AKBWN8KaPubk01y7GyGLJZL7b+I4cZL7qjHf49szZ
8sWmdFhe/XOJzWZVSJWBX9W9cvrnR11KyaNJmZvJ1epbbu5QvFL6o8NuaPtXYEoD
3WJJUk4ban4DJtA4YCII8oV9qGkf1PwjxaASITciaayeyhecKk+g0hjFq7WmaK3u
1FcE7qSBnjbBBLsyik9F841beVuOqrE3410MZ3ab9dPkodtLnF5LxESb3AIe92nF
AWBza/KkhMVCAYQkuQDihWD/wSyi+O+UExJ62NYvTOFYgBN+VF5Bra6gqi/I/h5G
Nl0/qvJnLbBEBIenBvTcNKj09F2zvNRFNL9+CGzZwTPI+M6ZU5NZHqhLLRaT8YKE
j9gxpyFTIVTrjJHTES3G4vXR0mhXYQ+1rbKBBcsoasj2dkGN4LtrEj+SqHS1YSSf
OVl4NhoJWJzYy70bMx8sIKIedNi1N03RM5e6kDgYnDnze2FwBABWhcJir2mlkGRz
RumOQs/Uj8dh1a+FuBATNEq/naT2cFfbKfszf8gxI9BqUNEAmEWVZ5CTmygLCc06
bJ+atWtLU6u4C5c5Kl7V3ahQnErXbwX4btnbDg0JKP/MiU1tc3LZFBmqlgJ7D/+K
YT1LagXkbrTQRHosJNEX1fMZCh1tBF9n5UY3zYAM2xLxTu0odbxILhiCTzeN//GF
MT6ovkHUQZaW7SBToBUWHM8/vNLy+NMgCN3hs9wKMQu9a7vp6DzVQrx9SiKY2CQR
zoI0WeDTVJiGPbvCjyOxHhjr1HV4iGPaky+9UpyCOt0/9PQawVHyCXGFX2mhVgI4
YE6hbQcyFh9E8S9NDIpTmzVgFhPntMV991CNDa8XXZ1+GzyFjciFOvyVfVXolVTV
/vcAPzgPBLytxGrf/m57/mknDrg6B+SrPM6eFkTCsjULkgCIndcB/CvATM8irGnB
2whNQFjkqJs4762HgTDNXEIRz3KBmsmPrrv15uexsruZr1lAF9HCL/cvpmtnvDRu
BPOR1Osdc0++1ijDy478QNmj1mtx1dI60fgFsqw7Q4fnkcx9ZFYMILiGhf1D3nck
CLpzu2F8FnQts3l5g2rO0jRdWvFTRf4ZTReOSud5DipWC6LUe0HuaWyvQNWTFUiN
W4dv1do7+ok82nTfK3p5IalKt4m5ZT9couOPjzXcBNoN5DV4h8bm5kLt6aVBh0Lo
OvoAAgIuOUipaEt9QfKNuyDDQ3VzTK6vVXHnkg+5N8mu/ZfpM4j6REBaIVlzoOFG
MQw/2VGjZWL4aN0eLkdr+DBSezl665t33vkDJ/OsrOKrqH72+XO0ZloYevaz6D1P
lWmndDVkqItA7ecqQvVbM/uVqygKwbcRGYl7qMI2b3/kMM4R/vD4PVs7bjh9y7IV
ONgpPj7L2s9d82A+odBmmyN26vp1frpK8LLHAehl2xHSc5mTmDxc8mG3/w6aJhWs
Q2nn2/T/wZlV/LghB0CxryGoSgYspB1c/78BwQBZxUqVoAABgZC9t8RZTmBPbsNP
RC6w4Q95ykckCKh0tqgoRAamt+UTORo9etxh7LpfENLVnT8oRX23/qVXxDzR0QLc
Tieg8iAidGqBn2gZZYKx6qSL9htFQ2PRZkYYg127rHxCNdg3ropc8qVeLlG+1KM/
VNva2byE7JSDFqPp0HJaJ9Y/w5Wjg9mGPgjV7WBhy/fZA4JUY0whMcyoTTVSQN7e
wsW6/qrymhRb8/h1an/o9cQTUmkyl2azVO5s+MGtMBgrHaWKOGQM9vJ1IdK2tlUQ
z8sVnsQdOB/y/4bQkDIxzAQDgrdFFd9AQF0AKiKFhdv3ZZ24s8iprsA/E8LtLr1U
ii64BX6Ttr/iD9PsJavedgMrjRleoYffs8JmVIrypAecLoICiDOAAF2YOV48sY1Z
Xfn9W6vFpCbcrMqx8/ihan3rbnDbCfSyWGVOfODyTjvUdpRA+pLDbf9b3XwRwY/r
ojtQ4xcLUqd2eFsP+le9FhwCPDfusI6p0KNrtWoTlAuffuQYfIcSAMvPNf7WGv/B
FnBo+CsGIAmaqi4NGWix0i6kh8GFzf2S7vQeb7eXR0bwCr59k53kWGhz+lXWSTvr
JeJs8d+hbsdUqlSoPOSo2uTyRaiqfjHYo93c9UR8rJXTpviynQc0Ir7ktCApvBrl
xThGrHk/TcNLSSG7ZDk3qk6jtcuQnsXYkkEVVUbbqDqTpjJTUeCDEaXL7r3kpFHC
iasAoVghdO3gylAsZQ0zxNc4o/lUo+EjwXNTVFBG5FaHlBHxamoeqYKn/xchLfEn
urIifbLZFijo6Ix7FAx/4arxu3HcJnnoBNbN8xHcjUoksxtHPUmRozysHtV+ZycI
FIqoETjJwFJVNhd6m48h+Uho3dMHVj7EDiPMwxhOpA4JefRXXStd9zQjRaI+oyyH
NNitq22uDrWk9OgaITaj6AbrGtQrMo1YUeMvjsTB0Lp6V6l15lKd7AanwbtrN/R5
V+L1kdv9zJikEX0b/M+FxBvgXgiEokTx/0NOcdtK1CscWopyS6BpiQPFF07+8sTf
nH2iQc97RoyXUHSHwz2v/Xlmy3eRvCwaOcNx0ATuGyBGRTCyRrmVfv4p/jiHsRvL
fE0Oo7JupwIHjyxpep2pSB2ISntHQ++MK6vSYB5p8F+Sq7i7PtEFh6s4Ehr0yN0D
9cGYfnL8FCy2oqRd3J63IlE4/83vt+ejxCvuBeO4r2feB4WgaTdmhfx0C4l5/JIE
16xM6rghxwYeZHJFRA6kXClYGvCsdVeHVcFllSXhhvoF/3Qm+Ghe9UL/j10JHeK+
21XZ06L18p7g3cspKHI827t5ICM1prdF4L3GJQBDfqGWX3cfAuZ+Pzj6CQ/EqJ9e
+UKGKop3rLFqpxkEClxNEK49KaxD9oI3nSlnl/kwh4PmKWqgsVxQf1XT3MT0roL0
nFGzSmQqfUFkDL5vJEG3+Iz2pVNtbc5ovXMhTXbxAUWxejVmuI3ckO0jfI4TMRP2
g+zgvJhcdzwR+DUyOhF3yKHoreqrXfAKhnhoJZWwhv4r5e4oWkozflFy7IvEBjEL
re8po7VmdGmKLdUJcszj5pmmiWdZOZr/vrTh84CXSW5FvpokdwrP0LdRSFvWHg2g
FV05OzGMAUpRkqBV1svRirrMyrEGtc7zD8YBlwVV+kv074rmT+PDy61w5n9zvFd5
Fus1aHEBTxEFqSwc2li0mHV49DlsKVbna4r/7uBkH3ge6EZx4qHtImYmexA3aRAz
whDrhK3QXjVY09lcRzuBTGiiLA0L99jm2JU2isuGJKKJoDqh1oYMiPtg4llMsIBo
3iw8TDbjBtvBu1+Dk9HHZMXpB9GlkbC5lyBIA0Aj8v3z0nQrDVzhcALqDbCUV7fc
DmuNjwlpfjM92tyYtVLq4vrKVELbjVwgzFgEihVLnmfGmP33vdLArWcDy8C3BurB
wzNA5EKvufS4CMVYApZwx7ItBZkju+cdt/RwnfJe7FgZbaEPWD/P1Dc9wIO2n01D
6OWCRLLrCz+3RIbPIOuTTYMcXKpRxYNq/pgpoy/7zERZPt6NmxTfXREZk+0DUrJT
3+BmfS3oxLvgo3egfQTaJWIU4HvXYXFcMnyLOPaZGuQchNTOz/rc0e0Nq2HRL69T
+5+6ZQK8qYwr5FmYEQZGjrjqEX8dUwmnfGxjj4pA3Wee+2jo7DB+lfZgL4JUzXwX
r5NwrQQ1yW1pydjC3F7eqOEqjq7mhj3GILqLht85yicwIdPw6UjL3C6FKLR8aawb
tgtAlWiAc4r9fiId/aMfbr6F4d5jIH+zzQ7VHbAWPNHXpzdyI0c0MIi3TyPHAjDa
gIm2xz3MGDurZYMpY3M4PLfZ6bI2Vg96/Gv9qk+de2iFyES+l01IUS3twOdru49s
JrsF7+excyTxCk8hDOyBtfvMeZBsHBHF8q9XU5OB7b2AIlam0h6Xv0dhrnkhLecQ
tn2pCrDnlgzEQF7l9X6i6YHhvPQ/0cFht9OHjagwiaixkwhS5MG1KJ32Tiivuwqu
qQxRPBFt+GxmdFXU6n340rceNGMuwSnvBPNXrR/00q8v3h04Eapm5G6sjYD5o5cf
dEAseF8aSotI/+Vd8nYKU5JDZjW5+U8MfzJlMrdyHVDuCyJYrJvrexmyRroFLsnR
D0g+alz00o+3Ae+E7eC06X6ZXnGnmfqjgdno7EmwOb19Yi5sOqPVPNSQdSr5hVVL
L1cKBJSKJ29el0yiKsIglLgfg2DdQ13wnVXSnKDlBvCCsfHpm6loKuoMp3VmZoId
sgaY6kMWTurCy1m+UBRTwmfiau7VhyU0j3j6Vn1DDqDYRLFEDO/8oKGObGmGRtok
eWFDBdoDEIbCxnKUUEl0q9D+AOTy4wLx9hEkCz0LwkldpBwCUW4HviFhFFx159So
tiuHBNYmDXXx97jzy3K9M0mzOEovevdgw2YDST+5qnyjx8Ujh00wjtdiYtwT+TCt
Komg4puIod5wSxojxQ/6drIS6sdppj/wPHeGmunT+/ane4x9vstCzD1jc5ujbvJP
6nQ+T5IZ6BBjKfC57QYJ/VdyZsnGqhy+ln8Cg5nFN3pVM5oIsWgQlVvZ1A5zxbIY
j3/ViVe3tnjiog1A/h75P6jkM1i9yaiqohTH3P11rSohxT+FD53TOOawhtdSumZ8
w+J4ScCN3AuEqi548XsYcNflDs5MdTuikrpaDusVrb6oqWjzu+2rRJt0qnj5xXtA
Uuw8p83DBMSN4HjzZ23wZcT1rCr+KeYfopHvogMtUk6OMsd6jng94pQcHTSXnpVu
zCi9lXak57iseAu2TCn1vuxvH2dIJffGLr1ghC2i30O8lCkTEqErKjl5aJCAM5Zm
muFi2CFZGsEBnfwQyo1I75ZQRE2fnG9XraKIyL7rwsc09ZMKFyQJvfzM/9IQJ6jO
xT9LVfb5+hgofsiYPxfqpwdygQCKJcA1s4B4FMx1ScTHCHYd5VaErIazlFCljvRH
j/ATyZwJLWOaQxQ94a3u/YdDOdx25gfzDr4UHDMq1NKpAb9FKcFOTifCkPcXF2dO
nQWxaj0pgLrc2Hdeh0lgDQ1QiRsOU3Gfqs1ZoK8lEWtfxStdrkBz3pZadj1ZcowO
zpv164dt+CNJRhs4S9ArVTDxn1bjHQkQpnUOVzLbIOS+iUiZMa2RqOlntLDHhge0
mHTrAbx5nfHKtJOcyIbtak5yw0qlK20V8i7JkGfkzDwvYaEYamEZKFXncMJE/GAF
+B8CEV0LZtfm84QrV3T27McBYDlM9wiXVsjDh0r6Dp8tdCZ9uc5Hbzd5U4sZY5fJ
7Q82jn5JkjxjlCkg5H19IMtmcTTHcO75OJbGdcM19rlcHAgKdK0MxRf9fodMQSfZ
y44jbpNNeeQA1s9fAuVDwBgIekWBcJjhsXIsSDKFwanCphPHta9zO6kFYzJBp58+
M1Q0yzF+AV5Di9385uFU/KKSDExzgkQkMGZ498/HM/64wmQm20/r1zqbG1SuuGI1
LeTbbyJub4vI4YHGRAUnWLMb+w3+axi1xaE160ykOnz3BlODGQCR6XgNFND8DBlW
HIj62Ty340xKKaPe5+HKT9xyZvDAOk+Q/2GzaJpYttbVnzC/qE2OWL/sGvsOoOYG
r9bd9xXLNoxIQofYpGAd6CPxtny4KabcaVLOXPyqk7nAIaVkpv/L3sD1IfSFLnyc
eBs2rX9a1zmbzyi201nP3tJYfrBdV/BRZ66JufZ207KV9t9dU47PZApMznYOkah7
x+6IgvbZ7gXgIUirH1vWJUP44UMZSrcWTwCHeiSbXcR2WoQsqeOpZuZCu2ABeYb4
YwNLG9f1w6X8BGpLSw66VgssClSFftEfpqSBqz9l3BeZDCrPB9mfjDK1c3RDrMRO
GJoNCLWQbzXFXu9lvbl1bkRlEzTT051OvFLxI3l9lXYkuzyxfwTpy8VQXpHveAbT
E9kVD5IOVm/4S7XMzBG31pTn9YJHijtODaZ0wZVab/Dpoh2fDIiwbw/8rMHZDKrB
I+NP8QakI/EV08hzkycluI9nxGpwvdH9HwO7jKmCgbLyEA/kUJOeWWB/FzZo6j41
ycECu9J0/iPsGTpQjh2pntqN710ii2RYzabOt6GO5hcHLuifgurRWl+QLyOFvLEp
o2Csk8Fmsj3HVI3Rit/aDUqV0tHmOKsMmImssHlabVfbNqp/lc1hVAbecze/gzkk
bHwfW90IvUaphT7Np/A281yeZtnhyEeGAM1CMmqKe5kpHpfwd79b8PifdLL2lDRU
iD1G7PqltQ6pAdk2Kw68QEvxXRl5MkMYyvYD1xukY7gERb1mVMahInqv8VZeqLW2
XAxYfLt1tEKM19S3lqE9T3R+pf10ixH3HNazewg3QS34O6PdnEoi4dhs4yXHKgj5
ljyzqxcaG1W7dPc3xlPqaNkdmrtwb6jp5cXlMZ6+HwvaP9bp4Uqe2TZVIXOCdk9T
f0y7oH4Rl4kSHbyccq1X1N1zWfmWaWDLDgQbTfdN4wsD3HubUnZbJyAsvtYdaYhq
xLvmKfgEUKo36qGe5SaQNIRnOin8KVaXTyaWKeQIxQL49QLKNodMEnQsSGLeKlc1
rhz/raRlI5BKOEb2JJOf1e2UkBGCwZfXlmAwI2iN67Jj66tzoGVukQ1y5kKn7Utm
eYf1qI4FHaJSXHWK31sXbwu3PWMz+UAQla/s+stF1/ikaFoD2vq1p0kxpn4hflj4
NkwPS7f1UT0efm1Ax88K/rE4aYpjpvtcZEyVTD7BC2fRqxDYF2XpJZeKSY+/cJ58
W1RdSTIszSskyB0FsqXNUcq2K1jmuiw4UwGxjA4jUyFmoaAWlt0H84IsWEMBfqnc
HjAj3rA4aRLwyK6BBKEdN78NhyJaK21vbOnphbCC+iEFRPjQ7ORm/l8UbxN1N33v
jce0QqpQvlxJinm4Xp8uzJasYI3UN1LM9g/JOa266twsr97ip95IXlZv8Oj4tUhB
zSYOXx75ORibsAPGhvN0SNZId/PFuecheQycWJzZLz5jVlsfRK6IRv1NC7tJCe06
HEpudv+aV4KhkM1btkSOK9s9vUXQhhFIpkgDmooTM2ra7yxT4zZ5ohCr5bgfoAut
HSaZwmk+URkuJTKFftNJZGZ2k7lysG/jTMP52OcCiSRoakJm2EbvV2inLt+is13Z
i6MEjX9lzhqWiMo3e4NSebrAKTw+IunjGeb7n+NXKPyxJyNDeJfO383VxUSzDaJw
k3oIQRSRL4B+RztaUamF1X7pDV1R+4i9rB4N4LGxYe5oJkwnrXnnU+yMBeF/R97Y
ihmUHpKXUOsOC8iLzTMoo41Elw51HLb4vAVecIXwqOUv4KPLC2OvRw/wzn4jVMJS
I5mRilgDe3cCTzpzZeVVH+DspE9VrCLZm/raZziO2e38uPKCHjMejx53K3/GrNY7
tAi3FevXWfYnp8dIYBkgy7TY/CKsruRd1qIb49qZ4Vt+irVFHNU7up6p4SO70Ng+
l0UOrQ+o6y65bMxn5U2Szhf+Lrwyr8ZXb9JljdNLJ6jioylk7QsjEidsNHGd1Acw
k6EZ84d5I7YtHLM83B1oVhm8CnA7n+b/Tp1JK6MEOEpb3zvNMAsUQbus4RqVOIrC
ej7icy3b9dwjWJbuKLl0WW2RnE2ofMeag2Ldwl4wJTl5/4pMK7UQv3zLAb9yGXHg
xOfbyS59R/C2Z8JdiZrV3/5SNIHg4yx7Uk0H9b5nLNGUV6CdNMK1JcgAAKkC52H5
pwcNOPjRKkwrzAphdeyAxaXvw/NOShMNH4T7upQi/DTs+rjOVsnFp1APq5XXmkj6
o8yRrNLeIA0FNNd9/MCmo+BDfZjWdl/Yh80Oi/BARLnyfQ3Pv6whMuG2zvMcIP/U
nvhQzhtqjU2gGMGxjAl5vvnQqanV6I7EF1PhhdpP8LoOclxq4aE7E7ao/Naxs1ei
DB6LxMtnSJ71S22l1/NvRLAy6IxEFV09mkATiMxUkiW5x5vY5AAZhBpZuQeDP+xi
0a8Ri4dLvIMS4kE1iNgcCP/n0U+WPKTfLVfjEFFWnOvyUH9ypcqW7NxiTrJm0CEU
yXcd/jrWO2eM2kxedn5joMaWSgfMRTOCkBIWPr8wyeZW6Mr6AB7JTN9aV0MGd0uv
MWnJQeEOUWYMAp0d5G4tB3OQ85zOHaCx/gxZ8Dt7iusPUAtV27PFgEleQIHOHu/3
of1HbWFMoo7TbzNeYDSGETES/qNNGO3iEbtUo6I5sYTZG60xNnpgS4JQEJeMxAwX
zd3WKeqSnaK8jWne5i6j32ptTGnjBB2ukseCtVqJ5eqaXC+91KkrwXmsZHqqEY2h
qw3Y2QIib/bW9hYy6iQNIC2Wbtcp+xBgOGWP77zfSmb0WULfhaYLP0xw92FYvKvO
BGCkg6Nc7pVRC/6sh/WHMLwy9wiAOaSMShwPgSY+I5jFwaiCAZOiRZpgPVv5ZrO/
kGGpH+bUVfyl5jS5ZwoMmtk0P8LUoBpUKxguqnoLGOo1ylpmjH9V2hCdpPnbEdHy
dNH9nDBYm4l+6BWfL5pPBpEE8dMkuRqXg28AkFgwbdjChNAacJTHZ1ipZAQZcCWs
yO001baJ4MM06X9WnteVEdhkvQNOVC9h2e6Uw3CZdWRgmCjeuCZMjOHQ6mZTVNed
WIQIpw/48p3FEZB81Cl8jhjH1K5n3NybT9HMd3psCBLLtW5FktZGOySFfxhkTRnc
KLZSzhkizRNrQDtFJ0ISmYeW10t4Jg1Iei/gVSPQRrXOpKQTJ9eK+58uZswZK+OM
X7EUDVSaMbZW88qedHTxqDnHBC3jKQdWy0XNbra2goSIkK0j1ohm2RSIyUfOCtoR
OaQ4Rc6C6owxd/HRPP4nEOW/Nt0jlzigefgPbl4QkOjxt9QrmX2RsO/kkg2Dpnzi
kjj4rr2GZnSUag2GWHdGf5/Fw/22vyJh/91YmxmPgD3zUL3Ds+YCK6aMIQYRUvUb
BVpyi7mBV2mBE5RPJRGsWpBg4OCTjSEAUq8v143XaCoZOVbzLFSt23BWBjZsnirF
45KAJEpgzLJt+cnv8p1moVB3Y0EPknYqQdrR14W84dl2GDrkTNdEi+vF4HkJvX4X
LBciAfZ0/sq4d6ouaMqk5eY9HbC9sJPaEP54b+DGGrcGbF368z2+CZdX4opMM7uk
joKABCTnydJvLh0SailX0jMnrG+qWtu+4QGfNBbg/ehQZynriWwr/6wnFKenZnuP
bF8MvFi8aa/4B+4J29tY4SRXWtSZbrQbCBJfdyo2Ax2+V4R0Uvggsi+qmY2Lypyt
XQJmgIcfyNm4pxm7CnDC7BG2IW//BFKwIVha8EISxnfd1ZGQKe5giMGgJxBn8noG
gfOPRuQp72gRXmEKZgR7aJZv4yG6Xk6kOXq4yTrHtM8sFNy3jer6UjHOUxc1X3qy
sZ8OtmF+QXopSGN8OLbG/YZqW4Rm7yz7cG4gdFVuT5SSvBpVkzAbrvzIgvGDOHLj
4CiQaSi09+uihIQ0NqHItqSd4TgIAywkqsSh8mjQ6KXBBfv7KCF9XBjskcCHBKCJ
gDMfSjFN+CZquu29UVIwqfyYYxveu4ln58Qf+lpDAOPWgOJi+8RrFJSleSpDJxHP
EPb5qZVdbfWsLekfi8IPsVwo4cO47PMqYZcn/bGesRkbdxYspU3GgwnhmWAQjzvh
nh0ZMeRIIYTah6R6VtnM3NZPeXnmMDksFepKzpyLv99Jnac0kuwWd9PfUAcvkfAm
AOk4480JNcJbHjXuaDlbrYwzGjJVlQ0bh7ddkohVLavPLqErE4VqsgXb4QtT/QIl
bzzVj648UGmtO3la14eubqHNNQLJHcIzw87sjpQGT18dcNHvpafRAcmf8wwmDBJC
vXMuvV54S15PLVzfBQtwiojBFyyS/J0d1TSH9Eak/qU0mcbHFBWuxep1QUPH9Rho
qhZ9Kw7njYmQ/3BfgyKrf7v53/0B5x7iqNkbZEcIZ2O+arkHCw9to+cWjNPqCFEn
KLAwSvdewogGO2NJZ/rzCxnqaYJgA+dvnr+8BZVrqeJIj505ggfYQcKQaoJpxodt
qUCjvDv0KwEB7VSJmBmoyUF+VjYRr6aGCkCrOApor3T0rU/iO+mxYAEqruJOSIF4
BUKzSUbFGowZOBaoVl9ucwyL+VcjNDbzz4cz1hxP1ABQoHZ9hxC1hUEuJG7bkiIu
BMR7h5xwZiRZdM4lyjvsepcMNduzsS9WdZ//drXEKsijDox377bzjEQBFewArr+t
K8nXyJMAG589451Qbt8KXQd8fhl8Z5JrF13ETNCRPpmYkqTSFZ2K4RicEmhchYwh
gBcGiydWsiTowA19XC+6p5F1nFD1dpuzknM+53f69e6ZVHazmravHyF7YVfHLi4O
FBXQmrRFdezgmE4CojxHQ5ib7R55qa7VM5p4jXRrjTrLkJFpI4641B8zhtpN5xXS
V4WirY4c/z1S3rKUZgTNg9tJYYAFQVMMWr27gSxiHlszswjMbv/6uo366kmveNoj
eZIHjnV1njO4lMmwepUuEhKq3q3zLaX7lsSYQmNgtSjh9xije/owqX7pVAJ0AxST
Sy93MP4uIVP1D0PSCW5/28RhutOuELjev9ZgwybKeujEaAZXO1N0mql/0sRzerA+
gdLAFek/ywODCckvTpkUPT0TMg7+Gkko1G9wu1TIGdpVVGuZEQfibDTweLJUS/ly
9utqt7f9fjEt4r1y52IyUwRUVcg31Y7jUbpZ1ijYJkuG57RhYKbqxQ5Fg5CAIU0V
5GlMIxTSNjgCcTncsdABiT8XRzqpHTXL4/mGkVRMM/YVsKvVbugpKVAd1m8vWYiD
rM93WDiD9pX+F7O7Fss8CWNrf/CS8Jg1Rq1G2iFW4q+4IV1P4fXphu71ie7pqBR8
jJfYuPftq2gy25VmH5c+uoBN5UocQPGwQxED5V4onNUgqvbCY1sA1w8yWpKETUcj
5YyxAm/8gLY5BgLT9gqADsnjtBR8UTp9N8Bnjq/BOX906ISy9ZzIAVUWsh9ARq1m
RM2ohbCczzl9XT0UFdNm8KXql9Ziv4jlc9xnjQ0mGWLeQ1XtqBJ4iLBrys+EwNy2
NE3Ayhld9Z4oXicDJT/Blv/0ZOEwxndciNnWhClGBVxhF7F0bO1rznv9+0A7Ij/l
PJmImRJv4N8cEEPOw0sIflfw8KenaoUZDxlQ6aEFBJ4FSjJxCVml4jo+5kbdCBsL
Q4FPaW7h1cC+VQSKeH4abWqZQ1+Gm3zlWnLkpwaEuqL1Ze4W+aP66ARyrnDvEd1Z
vgGkuh04ukeTq8FZ279Rub7DdvU5DPAKJFTnItA2ceK6pVLu/OpqSUiHcettVtS9
1Jmt+hHTxhC3FB4cdgPhy289ODa2jk+QJmYvk3qbgHS29j446isOL+oPVhQZVhZ1
jK6pN9JUbMPCHUR9+yngWmwgBf60sMsp1V1VF1eVuD7xYupmwMlLwW1+UkhOitS2
Xp9HcEbc+Bf4wbhsqPoX1AVRS8QzZ7cRxPZx/sklDO94vvLxXnt0NbDcyaC8HU8a
SH2Qn3oYKxgitOaCCsAPrSsCoMx81QqHJ/68spNive4KpBKi4plPU2BOObqHfxFl
VJRTpwYisYI51dV9YNVEfVFSo4AoEG5KNODudNCXpe8LlhDVOfIgzM9en/Ur4XdW
kxHXEtAoZnlJ9CSpJL77eP0pg8ODOfZRz5+2d7+Dm0I3yemR1ly6cdaIzEga/QJe
cuLZCBlUW2qhQUmVkvS3U/HVT3qVrQ+4O5pUWEidFQKbhVFe//p26RaWplYNtmyR
mcOQYkhPVbE1GhzqkkrcBtTbNJQJI0Vx64W9PZzD2H8QzM6BK/elf8yZmktpdDib
V9lxodE4JlDAAAzf0X3nOGvGXwBLMyrIGpT4tEDC+89tNvBewjlHNd3Gl5hc/KAy
l79c6lOthLuTWZiqdSzzLkILRFdtjhlkos8djsfyjvG0E8UC4kiUkSVz3oVFAB42
13NmujbNhbZehdlsJxIzQkp8aWFjSxH/zyAaSRqUfo+H9kBqSEwh7JZvrmRttId2
ZUBVqMGQ5Cl4a7ojRX1b0M+DZi+8BgHvt4A5b0Jf3Iqc0ZErqe7Pv9jh3Q9NQyWq
eKuaztthjbPMx23v/Irnu8MnxCbPV665whcoG0N2Ai3DJk4VETDKFazJ3kHqqPK3
XINiTCqQAbkqk8ErZvSGmPQW9ab9QwqVhYYChy09k0q2VBdbrHhEDPP6i/sTF8BM
2iWUTKoeJ/I3PPlS5pkQNz1I9ui4+5SX3j6PwfJ/bhGLjlljSOfHem/Uk2bNPN9z
FZe7gah8RCIaO3yt1P0yT1DVKUP08ZRCdWbmVLtkX/Yip3EgjAcZfKudKarzFuIT
mG5ZXmJs/FK9wHSxQVcfOjGRdnIn0+SNkY7Y3FcPzz6g5lGmJQ+++z57A0ZtzMN+
6wmaznKWGK9XOCZh7zcjPy8ng6oe+xr22ImWSy5X/gZUGMwsgrYLa42AaapHfdsw
HH6dXGgh0eOxqfuPJHrKZ3/Cr8ZoMycUQ4vfRE5sEsM1xPQ+y3P2it3u24c+NTz8
RgdB5+IvlGv99o2unqpr4LAcOwWmy/QMArun3lM1OlVYX1xmpVK3h+GPw9PGbVvZ
d/Wg4jEfIONGMmdKki63yfGzADn8clXZH7rFdqN+0rr5/0lAo2RBYDruvKRLTc8P
X/+O9PPrqvXGm9nrFdDs1Cz7/q8Lx4JoiFSwtdG9vr8DvoaajPQLJu/ddUWu8iLw
TzUcIolCY32bwQBSHa+/RYsduKpF3obULXmIEiT0tf7cpteE55szZRLELmb8WRka
Pbf4mvyjpAsnNGIoN6AjCuXkfeXEqvKSQr00NTK+h3kkKrNpbbs3rnu0ZdrPEYG1
uc6/z0RUfgh0XNsCb9kRwl2rtGFWXLbnFBJ1Kv0/LSPR2MzOkU8cM3BQNUY51Pyd
rcdPWM6aUnlco4YrveitE6Nh+juq7NpwBKQWDeVDwFO0l/yXtFmkL1Sys2rQ5VqQ
0YjkZFoRPuhkIVfYhiS2siDNyWBdMaiAGzrkoyYJXXzydTMSJs/LSfuXT0Op4U5g
fsjTg79zdPBsxnr6aABqASOvPCyqR/H/Xwiw9ultsGxjk+nbIy3+ow+mZ/PQdplo
fRf1RC0Qeo9mGHAX545r5NYPN83VwrV1rk5ERoPora2qkTCi5GCorHvOVzvxVJLq
y3dxez6DjHuQEa0IJTmDgXf6htXS06/Ns/Ipw5hg3PiakbGAn8+d26r9ySfe/huV
8JUBkqzKWfEPFmwDBHR32RrO1IZDiutX8Yy/lG3SBfzk3+8OGRhji2NEqsrt0gS1
h7cn++DqX/hD6TAgsPhupcKUY8TswMbaNUHzoeMFFs2Z8y4ILUqVVNysf/OMJ84F
RMdCEYniWd0UmE2ISfTJBsJj/7m0kiDjcWztPwU6r9vMUfmP9RC5TuOW7WaQQ2eX
YZ2HjxilzUs3Y9ixAo4qjPSo8uj4VfOQecoU3Z+JRIDS217968ajmc7OgFvM7Gvx
WNfmGaJ322YWq6b9EmeMlRLnV8dI19aud8xdijeGzRnp+kmYUowpRcZUEveVI6Z7
NF4s6agPA4vQnEfB4fxufqAmc5GgTrssoaHCzN+T3k3JS7K6f/f5Y43aD0IoPocl
LvOZ4kPnOsvikIjBRMltEIo4M8AYlnybcq+DEjr2k0v6AvuAYlHgQt9gVGoREvuz
NyZ76UHQ0r2zSLmnCpc/4uLa3Lj264UaoI/Ha59S+MzMeJLltWIHwNqUMC99edMt
BIJoC/U7PXqU2EG8LBqwKNz6gD2WFU+9lul1+/vhZyPWlwv5787cXbStaZBWtt+M
1FRJinEnQsuF3pEbZACAQnqPWa0dH3fdk+ZnJskaArJHXSm8z+kT+0f2c+Vp/es9
t7osU5HdBdNgUEs29W3bixO737UdonYF5Nf47GiDGX3HPiVtCwg54O5g0Ly6A7KJ
37ImU+/g42Otz2a8X2dOSf60IFly5ryj/iuJQFhy9B/9gtw8dZXehJUK6bIPgAdX
LZtOTagXRXvsw2NPvFJf8+qI0vZAgoyLMghlK84qZ6V6RQe+GDgdLj3+6fj0KZIc
DGfyj0IVRjx83Vyw30PGbaHBLo5xEb2arc7FJqg4gpOM/Mde4ut9WEsozMDuwFq3
yQxn0feaM0PGh6Qp9GFL1I/uA4qUOLhILaN/FeQXABzFz7+eh13d5iBWwkD0SihL
N5SjWfkL2GhTldu0FM9r78eZC84tgZJdDiGZRINFRDYEf8AoOzpjrLD0SlclRPK0
lFmLMKRC5Zb6KPGsO0W5IxCFNLHURBk9W/X6zKzrQL3Nb32cp6YfRQOEadNiJYvB
eTuVF20bYhLDNmZE+C3x5FJkOm7KZOG2lQpsKSPUnQjXEo2fnR6E2IoEIOvP+I2N
pkx7WicGTeUKkbzQ9/6TevCeudgxSWfcWWsdv+7txjz89Nc9wJ3dhcJusx2i9afx
ZUuQfPCtXax43iqBisxsXCDkvCE5TkxjipuLjl/TA58rDDN3sUIWHmL2ZDddbbYM
KUz2xnQb/PAqoB9r0l4FdtzrtylT/2Y+XAVBxgnI6ZnTmVyMcVjyiE4NpLSsjJbk
QZuj5nPcJytDZFiXD5eL5eEIkTz7t52Mby472CdaWWlojpVN73958H0d75TunxiD
Wu6tX24gRYBaQU7fy5z4yTXbU+2iqjJo30WK+jljyGobtw5ga7Slvc1igiTH5hV6
0RbRSnn4W08ms1GdLzMnOZZ3iAWWC/DHiKNKFHao/zHxQ8S5/ywiTrDrbEikNFbN
9iBBJKAmOGS86U+EDepQFQRtro0zWktMJzH9SRysZ+uOUYtndB8ONGO/G0JB0kwb
2AIhareEdMHqemjqkEc6FqQCl+TZV6e0i0RdrrMJ4oi2bX5xyVvY0hfM0MXZF4qk
l3GmnzZmjQhFjVwAtHphPIEVedHW5Udc/zN9beru0easlIOGONzvw6ZnxLecUzFt
W3/q7oqgXjtw8BobvQdoePbLqbKowFnk/2yagCSmvasJKBtdIIXx+Wnf83sWYF0D
p5xGIyezPUYE/yXn6mt2T3Z90v7FJOiIHUQv95YxItMmu4nmGa9XG63qjLA3itxj
5F5Vwb88cu6Jl2ripdcrAlHylYlK5KihVY/2OFIy0iWye5/spQEn6qgI8zfzanPo
usDgn+S1KYiKI+FRLGF3Cfj40H++Dg7U7jivVvkQzh2/dObT7DZqsEJ52YtOe3I9
K8bQu99DJZeqtVwVuLSrzeCcZfzzoZHxJDtyEZTQSgYLjBc/CSA0QaDMRL+NMuEa
vGpfzFoEHIcv2H+O0+XSWvvtxIf8G36zy+rvHXdi4ZegsW5tb9/qQUoajurmaokm
HDojoDTU7++cuxwbrchr8Bsw7lCh6HixtMMpbPc2KclNFLanCHxB64HSn7YRIXWl
h6RFCAqnk81HQSocRjCOLtPMvCmtN79kyrDYgOnWnDlVGJNId9dcSSnQB/TJuZ7/
Pi/9WwGYJNuHI6QgToObxN5Oj8luUoMUMk8Jry4pUDIDwpDcR+L4xDF4oKYLI4kr
d8U8E9WMh0iUXoDo7Kz0NYlrMvr2m8+cPQ3nXZEXn9cP0g6sL7suUVVP/ISK3MYK
b53Y1KFBklcnYvxE4/wcy4p6u9DH9xxb9Phd0aMkkKSWzzKOTwrLQnwprnMPGl3I
vgNmxSNWjHZJ3BveVr1mBGYSecSQJk838xIOg34IUzx/SGqvvcseAq6qp2gzl3kW
mrtg82ndQe501TAErLrEa6s4podJYWuKW0hgPlDz6B1LYFS5EL9cJ9BOoJg5zMgE
apDVd+IkbTr9olhp/gpkDyNwLK13miqaqRD9CL0PbUIEuMRP//13qIFOrM5OxRXw
XfEhlMmK1YM1xXNJQOKc6r50JY1Ud2U3KVaOvVxLG6Evvre/b+cjo+Z/TZ6f1JG2
eEJ0x4kVn6hJ659Eo5JDp1KUfU+QtelepRawTb3n6HGD/pEhLxWq4g20kVVbD8zF
MgOUlMogiwYGHUiYueegzFm3lOuezCS4zY8ApL8QIo8gqVunKNvmS18SKUlbUPH4
22kQ8hGMZyBtwxrrVFiQYjEjsGraD4UO/aeNo8FriExD5TzxxMA+ttWsLccShfeE
9/8vrsY5l0A6vbqRGkCKFp41j8GneRNSoeuMRFPj3jnJ9tUZ92iOkA6Q4cUuT/YR
SNaIa1vHkAvPY5kKhklFKuL1EcJRLNstAYC5UmrvkgSybXM7fG9b1EY4mXYbzrkj
09mf2iEB8DMuxiQ7tvsQivr4DVQguRL1ZLckhoFZpZbdEW19QvGYsYIX2Wa3n8X9
NUz6+DgrCcwVml14tSp2IZpeDtAwQ99e1BHbOU091ZDi0dx1nYtfFAoreLhuZfQt
cJO9qcOXw48VbVgmLcFgh0oCIbB14b7F1IIZTx6Kagpaikiq6IIfW5aOdzewkciz
+ME9HZungcR3jeUY5NCniDZrgadL2nEZSFJRISIZk2UNyFhDRD6dpLMworwdLUI0
4Z1J69c/2H1fJfW30oj40h/5OD0aYi06GJbqX6vebh+UuRBI0DUizoz5WNtOSNFl
pZwsGgr7vlVObQGAq5DHjOZcvWPTlV1MUI09QEGsatrXNEy1o0ca56r7BrgzStLC
Wf3Sy6UP77OKkj9/Dz2lzQyHcMDJBZpaz8ILSfoD2EcFbUV81JKsci1nP1aHHER+
UBSqk9gO/dCbQyXN90Oc9G1At+dJdKyWbCfFAv/JtmNAWFXgRSc699YV2xCX7WgF
vTdlUS6QGFNN5N1Dl+Y0ZJGXKquewjNb84w39ZxNigIKSyAm3t2JEnKuU4kZLgK6
Ejo6iZef7OcfWEo4UA84pzqptUAPYRysUBLHMxaIuk/Dy57pjy+mn5s9uGC6JeKZ
wcOz8yfEVXRmrHGtQ4hlRAcngXqrvfUL2yBHYGr0nmWQezpPIn0b8qXCS/PhecGk
7evKqdqtm+hO5RpKVPsfXGmDfFOK2pOFKRby+7IIUQ1hx1iLxV0EnAxwHQAaEQEE
uG7LRsBXLec8mwiXyyehQ/YKxnKGxlBg1B2oXQuFDu6QGi+G2WCuYPIShWD+TYKr
QXXkc5ax6kp9Qt+rRAKxe/B8RTFYwDF1UG81Hie2ilv8/0ywYaWp62b56UWW3MTG
j80cgpqKYrew8tD51xpnrwz3kYtOuQatF3UnPJ63VCv2P7Ygeme2R+UPnW/FftYr
NyiQpKmCA5yuvYzoY6yRlPtp3eIUwcV89wu8OitgDU5hRxcPirbLmePClWEILmkj
z48n5rOWo+OzSYSb9DvExVLc+x76LClPKitCg2q0JTMaBvqrFl0XjuFycLBn8DE8
EIYUnA3Kyxv8v8mmg+sfmvFTDSLOruT9bX4zW1Q8/3euTwUhTatN/KqkNl2SyKwL
GmfDtM0vFwPa9F+33wG5av1RQwqSCLLosc0zO058O6itRDZAtF9lBg+8VJemlraG
gcnKHdCf6+cw1LNo0VgcXAnbCtF/HLBMK6DD/GxUam9uULnMQsCQX6qFh1uehVJM
a6us6TRebijE7RhaCPG9BRktfGl7DiFLQkCQuzeMLZSlGn/Wyqg0qp5MQmm9MO8T
JrX0u4ttYfSBw0TcMH/xTOsa2tRODcZxiIAw5ZlKPqwN3GzLDaUnoC5AXNuEwcfU
K3/PX0hy0+OLabWMEA+o1Omtg2NSW66OqvBalHo3DBeAOoNjujPTEldYNReUosPb
wAEB1L1q9TWj253M6/1jcTjkVlx1OCW/1nKEC3zJcJPO55jfjuVdGxPpi3zUCkzc
++zJyaka5sUfLKSIgjhzTvkAhDYL4CMBoCH8zRSZHsGhZ/fbt5CVvlhpiVsx7a9Q
+qYCotIBbVRPdBEXpcOTTeqQXLEKBTejIHrBNEU98Rmm0B2ld6RMO3fU9deEdZzP
tUw63ek5mNY88HWJi+Qf7y0zXzRwB4SqzJWh3HdXbC8Ot7+fAth1E2DEMVvkYPqP
C63lCxzsK8FEVT3/pblV3YMirjCTWgzghBZolHb28AxMswPv9ZMgZQA50OZmHZDG
GTx4/axk9pf8rZkaIlnUbSQ4NyTcXjDQLHX9nr/GJ+nDW8AigD4tklEr5hW77DnO
aUjLfoZkgE4r3hqTgsAkn3d1uygJ1c8frbcvfUb7PqSVoLWd3/x4W2UAcalc/jSE
yHaYLAFp4q0z6rlLQFM8r7UxGEM3MqGh2zVQk8v1LnXgpCkkVdHo4dQpl4YCcLyK
tjHDMJ7p/EdpvKzB7AW8v7ObEJ1j6Vs1BPwpsfVnnBhSoNvJBYO6S6v0YCJdy0Cd
jPhMtoNuLYHmCO5QZf0UBpDlSUGUGfiuzJT6o/jR8PyEinS4l5FN5VPYR/IXk0ZZ
4t0U9sS0fwF1YxB5aWw8iOzKC5DEHGIyuGf3XQv7SPFlGTFy5c13ZhvW1v0lPbBN
7XRmEWW/mV9tsFau/vEkFuoG+BuhgFHbmEhPJje9OxVOs0DifB0DNw9QEbOiHncU
WDwGC2jeMIDdWCEqubp5qidMRVsz/mEaeBPPeb9F34US9LgUHs7dfGRHZJy+oSQw
e6cU2D0xjNQrwqNqoIuNy1I51jZd522lniWR6Sqn7XBD29gOPiNyXL1yyfM/RBpC
13uS4RN/Ayus2GO5UpxiEKtkQYKzccYC7kMNjl2Tn7pEvqLPFh2JBhC8bHop7u2l
YP0J4xoIuKP5bwsVrszQYTMS/hq4KG+BQNNEt/L9i8GxqWVig9xCjil+kU5mqqn4
E84oqLbXgZ44yL7BCsK4g9rePWvDMT079V6LkD12IdWYTnfpnzSY9jImJVLdUIWF
t/m7RywgDui4v1J5SsJuPt0BOxvKzoUTr36uLQ4Ztx0AQsL26Jyd64/qfexB8kni
vT3hp/JYXFezgUNAe+wFjouAAIZVpkVWQplw7dV5Wv0xa4nOpCM1NZBcDzEzLLRC
ro4fONzXFe7jSjp68qBkAQV/gtmtQUoMMIANFrDxO5LOuqvMoLNfZSvN1xBYj2Uh
USBWziy+YNZ7TEsQ6KZQQrgUoDoBwooFpHpVZOD0SBMTEjNI/QDuWufVNqfXSD0j
+tVatoiCP4qXmYFeq2/wJyuny2NWX9EST2ib/8jnvxd4o7UAH/3LFnq4qft68O0W
NGMrx8d4uoi5k9bFXfDwNSKyS66+xYuaysRaZOk41kbMXkEbvl6sl3R3oo5P9/IK
mblHze0iDN1PN7TQxI7K8Q/QF4U2CIr0r5Cn4S7wJdxU90eW/yXAvUaYDlvjCvV8
5euwQXd2IeImNBZQeoey/9fVF5sRQQmDgsME32PXiOlDW2KWgdSfZONrM/Oq2drC
0Q+WAiArlLk4xxfCA9CgwvgBm/DGJwm9BagdQK6kRmdXJ84YUY4Zor0Ay09a0iYo
MF5+/UbKmsYgBoj+i/X5Qx5GkUWS7gYHT4ooCgfkwQr1Y/iYAMeTK6YdUH+hg0zF
w/yLoVDps110SZIBz6J6MtlaBuQRHHaVqEJ2XmNWC++9dZpuGzpxlzonfXoQLJ3F
4m7QRbn4Bj3OBLpKKSCxDVLsOU9anLfKeqh/zNa5CH9bccpC7SVQmC2cHFiSe5G/
e7fic2ZYSlsOin4CyRldZBLiQXu1aeqkAOpY/Zsj79lCnUZliNXxzpnLp2Ajl79a
J+ss2KS1e9oD/J3lUTWb6n2j4HIV6bwn/ZepJ4d9COHQa5VRXYdS9qUSYNTbfERT
8YlRNNj3gCJRPfb6tLauQaQGaC+FVg8esViFX78TNFyg3HGOZ81maEGpBM6iR4Jg
oe71Y8h5s5fsT8FvhLz0Yj8k+X7moncpW8IH3niIR4ab8w5WcGfszxzhovkR97rU
NfeDaERGp2LseZ1s6rSuS/0eCss/2y5Ac/RRUvVUPd9RTd+LoRs0vFYHpUSnWxqD
9yvwmeDgwcqjS15QU+JW8oaqxjTest+ik7QqJULcaaFVSb/6T0J6pHGCbxeJLsI1
TO4nFxGVeDUe6MGSMuQ7mPrFis6SwwrqESw6o7g77xVjujsGzeXH5tSlLjV1tEYt
L3A/HkMK+fT4E/kvMO5R76vmfEBkD89f23co2icX7GoczHYdpRJB01tDonPqwlaU
RtcH6bMev28DWSUgtmtsNPrRzNlG6nvGEWDaeEfnNnPUMtP+l8VLh3QlsN+VxFrD
lmsPNG7Qwng374W5WxPuZFirW+/2aiahLXZHbKoHqDmcCXpf3dP+SwKKvRtvZJUS
Y6xi0PqbhdcRz7rQ3rbv/aVkgfuQ7UM5KjeNZ98YvojIecZ/b8mFkW+zX7r2t9VC
0qHkqPzSrmCeQ6UuStOeYY+pTXDxa9dhGMjrcjKX5XIcX5WRvLVVZn695DX3KDDk
N1sCCezIYy+E1SOr+GC+Id5KmApD/udqwzVBoqmEskMDTo/3akwA0dGQHhyDNe0Z
aCuZRHA1WJSTO0fdnNFKAwc0cs8h+Qy4AEldeM/lhFb8AUHnpEXi5NELcZnbm6vc
pGrZGMpLqT3CFVxx9oddVjwtNsUtMAOJkrOn/amKLkOVSDkMzPxNVydN9NZAE5A6
kdkrmLB3TC+lPs9alP9J/8EZ73H5z/2Zg9fbm1ywR2gqr9SDdjv142a3/VOSCm04
fFrCYDugS5WhF4eLlLbJ0l6gjoKeoJbjljxlfAWa9onexjGcy+dOqncikZZud6QX
zvPfhbqovI/m54YJX0UzPX/dL/wsKKFL+9zCkNLM0wyVB8/3+NoveCTdKt20tq4A
H/PLutoHZ5WmbzSdnlTJmszsgPhVFXmfz/xxF3pW96t6Uf/0rr/fI2LmWLrUkJGa
5hI9xNaUejEqQ5iRRy2fP3EvPSUSxP2X+1LdZGqVh3SnsSu3FqX6ausYJG+e5EMo
o7pqTQtAlQICQUvhxoVIQStRFaAYb4ZTx/b8YnqgNBfOO2Zugrrnplk3nhstb/lq
HA8iaYPjwbRJQ6lC+/gY0rHk+c2VvORIxpyG/LLX031r+RuWJ9Jut1G/Orun6b3K
9X4jTjPao1RFY445/KVS4Hn/j1lt2Fb6RfZ7T6ytR6pyTTQUKeZT+JavTbYkgVHD
Cdy+mW3txBznYSL5NmHOB9UqzepPqynAKR9PTm5m0Fm1L30e+dDZFF0C0Vd3JSeu
gycPS8Ls74et5VnXOKjrHfAeWyIY0iKOi08HXqwMdmv+SRzR2SlBxjokH+uQra+C
A9QMu0UqXed804xYwvMtBEQf8RM7R8ufmDBqpVUE2+DRXHmw79RBKpc4sMtlINDk
tDhnIvK29Nr6eNPSBFH0v1dlIY6TWzLV8h83hicgiW6WQlMz0RyutbDtI1nR9RVh
KzqlAdoCfyMHVQ4uaQ7ANj+WXSI6mmch3zRf6lrQU75WUZ9VQueWrRGRBcjrCXFR
3GsCd1p5OUnFRYTaO/a+7N1f5tW9bc1gH7ZweO3caNrdIYXBoiWpI+RBKsRjf5Cf
8o4iEfSpy5VLKwRZNxlB2yOz/KSwJexUbjZR/hjMN+xoftcCAFeAzloX57Zx55E4
ZRz6oZ/IcTS6+6J5U6WbGZGSORMiWEBZSwsvdtoGwP1tstH/nLC+Jl+n48d8kLDF
kt9JNI4g/nDAFqWgGrmH7MtmFrTg8DEgWuxXifuDir2bi86eBV/OlTty1ERk/9hZ
9Qp1jcgrDAu1Wyh0/fQ6k37MbY6xqsXD4Oq+gb1kraq4EO3lPnn615G7VSt8sU/8
awP6bc2GvXe8Hyti0ADWJjb5FJH4JQZhMUSwwPodxeB7NvPvwt/TcAP9exHg1/bq
cECnjTuv9G7OWqi5zyE6/ZPz33okEQSeR9dk2ucDjXxkRGfTsGXnSvetW4H3AG/k
MwgBk2ZL0RNl5kbQDdLBbCtKgXsO0bB1tfQnQ5V/9s6qHYY2Ma1H/0S2PUston7u
/gdvfPM7vIZGXBVpoYvxeRHUU8kcfTObJTrnPt/MMFtstVhmxFKeLG7/0WD6u4IP
qWC0uAc4CV1jhe4kKGfNKKI9/x2ctvj2yMZ8kBZiavZjU1AjrGQgva8dWQkq3n5A
6GkNEbxaZnXL/9RrzNXuGZXxMk4SFGJIZ1T44Mytx20LPv7odDo/D88HrPq2Y18c
70Ufs8NXETeLEnh7pLdq4u/jtke2/KjGhgTYgpXn8d61JO6KvbAL3pw8hODXHxcV
O1h9dw83X0Xncnjnb0GGwRFrIxJyJeqa7ktt/bwkt1rVhXtZDfLRmg6N+Q3oopuI
PHRhKMjS9dQFxaB+rlX79rappiclQmHzU/A6GqJbwjlKaoIrN8mWsDoUNQRGxezM
97u4mPqL4EGyNvBtxHDgOnf3oO84SXqLELmaDqdA9SrzH9V/e2XhkvATfGqQDcZa
ETdNQz2Qc3HiLOUFm4HtNMtk1ruGjzErNG5eymQN2g7N6UrJhjj9MxvOYWLAziew
XsQqRNf/EESD+4PZaTO6WFxLF6ggpPHEbHeWI5ruffGUMnDl8StuiDg0ASfHUV9N
ofJ2t+a4cSE2HguloDd/vlKS4+RHJu3xlegILH+a/n4v8/HF0JxIA9AtLV5EgJ8s
7IDn0bGnOeobWNzJnRKT6JrX/SgEXwhuQlLgDF3TNLc7Bkm5S63gZl/qIGcJgQGD
XJH/Unx6wzImZAVwpXsxJ148EeYvgb9mHriJ7LmaGhrI8IQxBU4ZguOpFXaxa3Y+
8ykRj/R3DDDZs3xFOB3fBYJsILuQ//fwKxI+Gtp4rDHsCFmdaLikdC9K+ROZxRUb
+nQd9YuXX02tc7Pw4p94gpAzaBw89snzLLDke6MA1E62t//fHa689IHqygT7rZXc
PtA5uhQtYXGBMwrxlGhgX2hCpHq4gkbL+wvpeYeo/13CTl5goVk1Tv0pDQeBx2Kl
6uQmGkVILEDVXjPmJt0NE7pBwEbpXzpgnDi/YDKEYUvFSBOjDM8j6WobwwDv+pEu
7VKmKWJb8ylEutDehbdkUnPU0d8a/jFADSYIJpvRznCOoyxzl57UlOtSaz+ARQEv
difYAPL8V9qrA8Mo2r4TkF5cnop1NTdfLO84WJfy1Jwqp6deTEbwLaDGMd8ZJ6UV
fx4hj7+37JoS1V1ne9YWum7GCr+cCHLDDojbHLrhQlY39xU+HnemTcDXp8dPqT6C
fb5P5kHCwMF1BWhupXAo+ST/LsHMLmt2mKRKv1mpRYTKzOs9GnMgZ4p6i0cc2ISK
P8P6WBFV/pkB0QvnSm23QJAkVj1QIKC3sAMNcWce1ZEiOsm69K/vmPw8LiY13ghb
zCxBQ3dZ9h19Ab8uE9Q3DUKD/eqnVVTQ1gse6ERToA/OILMcRDVXeAuR5Zwxmnni
vjA2dbqmW/EMbgh/PZLq/P9RdlFiXW14EWqAodd555bqasf5zDdQtEqizXjFRn+o
m3GVNNHNBUBxDROOpcLmtXlpMaY0GJRcpExz3kZlC2VAFpc5Flb6CcZzIliksayH
2k5LTjXSzJUbjK71/fFvu1VHgvpoPkoaEZQ91AhwMsz5hjAGeGW0I1NZmdllFaj4
xt2n4jEyIrYSIG3w6T73HnW2h5T9uffR4a3kRR7yIRE6FcgraKznAU5zZyT1Un5e
4bh8A0Jt17fGTk/wGzjgXY/jRTJlVea10EJfYWM+P334syKw67kFEnC8/abyV+jg
OwK8o1f7gCWjodWbmssDZWukmzE9QIBy9B72vsbWYv1oDGbm/Pa5dOdsdhjdmiVZ
96eQVazzruC4kCazGlStKd5nifEvtnI7FPENZiI5YtUIlKAGbwmleZFwYkeRUTHK
UPzGT4rXD9grr6T/9s5Gx+KpEL1VlrfmUwTH3RbQSmeVsbW7WUOgICypoCovHSQL
7hrroW7WwzD5agNWMJnrivNbszRdgoDXBaadbbOSG9fUkMZUBI5YgTbKXwTkNBWq
1ZXtaqOwtLcsrLM+8+f+aLa1A6la81v1DYrZ7hYB67YdONNQPmBzV8LvyPDwYJBC
g6//OaBjbQ9OaqNjA3EGGh6oZZnr11V2R16tD+8//oDb+ME0UpmHVkFnhQOHMbSt
TvZSx9+CJeQWPY1dedBujIdPVqXg5Th/+Vt9X3wHPbvYkNGX50fJOe56EH/fb/mG
QTQqf6DF1Fb8SBO2fKpO+sjn1y+RmP3L9+R7Jf8e9m++M9XGM1KcdkNnZ++Ayv+B
+wLO8y3z0W90XzmEDi6FIjybjNxq0Ay9VU2G1AzJyZPPLKOMFJJdtgw1BcN0ydSN
OK/SmJPqfR2pgwgbyboUxUq/hYjV5q8Lp75q6b/+186MhzzcZM1TxFmpXPSkXqI4
dTA2YSo70PY7vrkPy/AAOhRmMFoI6kkJx3xgY6PO2VvRzrtR75oWDdmbMQDbZ692
x005Na32vUOmx39QOPdS0YvMfOrYPbCfOoLbCRdWqjhR5lXIjEZM7tZXzkDPObM3
qscWbFAo90IrY6Uv59D7NFFiMaKjllHIYLLCGoF/gTTjhD4Fl78Yj42vzg7ZbmPM
CTHWFfUlTWeqVvpFmVpexGAxnleTSjjhdXOfZjCN3cKfEO0O/bBAf7hLFoe/FAdP
YDVbMDHJTOjPhcXHWulu7lQ8twBZzZQjKLJmXZB5JFBNPr5uaxFW2xGdPlxgc+ZY
NhDKXudmAuXT4cGej50NND9xCeXFD97ZElztSfMOpOwMMVoLZ8NT8iNx1wn2fSiI
jQUwvAxHVDZGwXSAX1Vxq0QaCTe7lPFko19BkXC8YiIq8Iem+HR3Vk2idErfUiWj
KSUpHTPKiklwpjvnNhdNIu4Hkl3tnThpzH0Bjwg/UfJ4mb+MZGH0Ibf3S4ca/q5w
FsHmKlHV/dbeSmMl9Bse1KgI58PjuVLw6Xi/M1hYazWAX+wq6t9O2B2Z93TcXHkV
/Og1UQue6V0985288oH73c1ACTAX4Lf/4pqF1P3nhF99NA1DD2zXZtQxVRNc4ZHf
vOq2LF2Y+OuoIH8iMUMR0InIt0fxt88C6WTCzIEnCqbPKAIBwCmrH2d84aQHiGE6
bbrbnLG/t1NMT4QFENpkZfLJbP68r70Ca4XGszDj/0CekgC04hpotwNNjv+1djfd
H4hbJoFdzKidary9R8m//+g3hxNm/eGXoMpBgPNEpSk22S/WJsIhmXSrNmK8phKR
kL4BPyAtVDSz4c7Q/Yw++L10aTREoopFlgVLku2ygcljsKTDFIG3vpJjOvOol3KS
T2xxwW/yRdYTizNfYMrrRKpfeUlP86XdRR+WIj8kprPjx/4ykB0L6kHTpeUxRbcq
mHeF3uan1nLwOA9c5LWEYJ9QPEVEvb7ct3GL013grTV06+U63xdLETu5fAbNN/Af
E9/4ZDb7VCpFM3Ka++vONDFY8sitzAlxjtJ8F50gqenCjH5gYXTfo3eoTJIH5MAW
qcT5MGQ/Cqcg8XM1/bycBSed8m034RYtvOqyT5z+jNFOGDaK+tGsa+ThdfOCB62Q
DCJyJ9wlw0ELOF2DtgP0uI/a1hCdzsyU0zZc5A9ub8Nv+XhM4x2c2vV962px+FQC
QQPdWFOShPZBpXj+hU7LfVgrCPO/DAv48zOJ0R0C33K0qn7e3sK8hsw/OnO0dWUF
WA1/amJBvy1Uv1yMZqSHHcCvbTZClZP5iEyvfITvfuG5mA4As+H7DxNmbZyuemA9
jhlB/baYN576dI+nS/YFq8n9pGV8PrpIPOzqknqDTC0Y7mD9ZP2uaSQbtqIGnt0p
tKJZ6Ns0XD+wKU4SPx/gi5e1fKLDjM3ebsd+Iwbuow0hs0QmNYuNNXvtGJcc/IIe
cLJn2oPj+ZZHPwEEmAFqmFZDVy/8nT/1Rk75ZEDSDpbeYSkhG5I18Nc3o4UZCvJe
zNRji21zhV/sXe9tiYxkZ30+nVbdAQUG3ry8m4dNBctzVdt8MNk8iPRDqQd8yh94
AdY8E7w+cvby0lVMzwpFbOsZeZNeoCwvXJo15f4mif9/E+qGz6Kcofz+LRy8swyK
bZ7EDz43vBvbvVGIaTs7h8oE2wGCowxD+FUdoyrF6X/+drN4dVzJupOXSaskVm8O
v2wx5M1CniaMlSXLz/85sKpsaVOrDwLfEIjSWRdkEp58I55Wr0FHSIYELrS0pjIO
CR0GVFgtAQXX0gvDd1/Zl9rxllfnWCL49x9ZATML0ZgTHhx8PnhVAz2zQrHRMPJA
IY1Rybk45pKgHp6LFTvet81HB32hjrSOC00aiJ9K+LTyxYIgTnsEsjU9EKNbvJ29
+4h/OhOHKJbBzJtAQfqzmu97vErrOSqG4uCpZcjBKYwalNQEDwUThP9lLAdnLeoo
pZ3/o1qjM9/z5KtASLInPdXKVfUe22WLJil9HmGgqq9oQz+RtFUD0iabLmP41K0A
fqQlDVsHpN6xFvIL0NQZtYVXqMxfKOKholNN4+TVaPfaCH9uKc/NkqsliBsUDSCD
UCHX28p+fPprkEtAwUXVraV+pWUmIkQWhPC9qMmgDWoeGuN59E40ALJv929icEVa
3ujS6a4HUxlvGFsH4GU5LkO2qMHhp2Xzj8DaX/T990XwZqOPpjXBYbeUZr09Y5bI
VjJkpggCewSc/S1mu0HllH244bTUmevstCdgIRZOH4ah/Myfbawe92QjIzaN2tP6
3QNpvhS5cUypK1HFM9lp62hN+groMz911IPKncyWE2fZXi4eZpAC1U52B6doCO7F
mfwQO0ZBjBS+kRsVT7Lzm8jBNbCDov90CAsjGa+o5sRD1hiktrAzydw00cwDyS9M
nH0J6/ZBCOBND4Zmp2WMMTawMA32v0NrZuT3FyxEQH7TGFr+iYv2LJNkgzq9J0nt
4Duntyc2xGGSHfvMfKwkcj/uLx2r3Q8aPpQyxIPEsNBx3hrgdDegm3Fm5lM+g9L7
RINDBLtmNzhWA70bRiw2lmJPkUIw9650wqMWxfZN95gT8hwAjOeRW8qxL+G3ijL5
1ZnNGtzUbdeSzmqN0C4t9JUFV99sOBtLBrkr8AE84rASmhNvV55+MSRDTCFc6Zoz
vLcnMecyXZ05FrVV/ifpX6bB4z1jSE4u9SMYGEDWDLLP2fHxoIawu1bio9nGak7z
NswlSlHpROs0AbuBoJFNqfVw0mkT4fXffhR3ZQQR+h69KziTkbpcNjL446v5qBcb
Tt3etJ9aRwZ1fTccjOPvUp5bXMrwND2/ePS2D3VXADqUO0qOoH+3BAHh1crdeGAN
7J74deBULRsPRwDi3PCTep6fMTWa5fzDNucs8XsKUi94N/+0fPuH1EFuq8Rc+1/w
idLHg8H4O6D9mmLeyV6G0Aha+w4mviWCX5Q2dxCU18RMV1VdUPNGI9tjr3lMcOLo
h0yg+plY/hLf8XHXbvdiB6w9wLTwjGxCMdzq994R9fI47JRXlhlj/Rkxh89HuhKD
Kd+cWXY7FxBHeH3ePD1cv6wULprg/tAmxEVuxp0hQMbEF6u3dg1h3BAJGF74lOkJ
I7lbzMJmpqUsxbrwAZjEVTt8wKl8ASR4JcSCeJvblYA6naypVsp9PBW+H/bJyp4w
SkHYxk3t+jF71p8Ea76hKz3mFNAdt/KlDlTTabgiam2YcPs/kQ8j6UK1iEWiM0ja
yXCuKn0WRFOIChMaxCcgewIQ0fdrnfzscIghhbVNi2GPEqyaJxbMpFqNt37sO6F0
732PIOOn3FXoU32KtbZgjoyxDDmQ6Y6KOowiFSHJBgdYnKeYJbwy2MGdmsLKxv5P
4l7sGiCDxl5wIkM3+FZSJnrBRploxqGG5XOsPiAXbmUBpko+xveoKuYnDBkZgidi
1sU1wRv2//R2R5QkTwJtPoI0H6kHZOqWerBuJoLlc4jrCobuYUVy0pNmD2jtfVYt
G3XYtEqsUbAZYBApXHyZ6toFI8n8LrnR7X26uQ5TkHbnWNEqMfTAzaD2BHSk1la5
WQsU/K+DCCjQ8qwZd0oG0jCGXbTU71Ou++jwyKwIx/H+NULXZL5ESsRTGobF5BJu
65REgDdsIhCBk+qHw7lZ+xIQ3IRYziBHROrLe1E1RZwdjZI7eEBbVKP48cPn9coy
YI+YLDO/ESC1Ga1IFjj+QsFTIx/lEWflsiV/ZPLk8Mp+numAHAzY8QnUDNALBmCL
uEa/aOJ1n7K8Kgxn+OXHgLr8CJDT/VZVfgW1V/AeUYPrixxIdcD7yNjLdB/1HCYY
JSPHt5NwW2raJ11ExJKuluUxL9wi1UdOAdhZtxeSKVjtIP4J93Ni4b7Phj8Lx7h7
tzTFV4eckD8mcYEOdxWMjgaebP1jEi5e5KRCKNxczyhyXTeglRyY5hsKkMmZGV7w
pBcUVho+7MJixIkdvZFMBX6TjUju0bM0/hbKFpkyFk3Ohy9vtuAQxYqVG/IIqKVM
jzzxowVM8Sk52C8o6FoFtQNPNLLUoC0lrO0l/Y6Cp2FxKv3SHJQ0FDi02zqwyG5n
fOtcCEThbn4MweqjtqiHELueDnLFdlGCMmGjFEb6GNLJFhz2uX6Ikr5BpnogGUVj
aG5x34lOsfAUzZGch3+8IC+h7KTAr4QP3BvjAt1/FWSHD82Tww1m3vT4MpvIqOpJ
S5/wOLzzeNdEU/Xj1PYzdcvP5J9d+iS+JbCNJRn6e/oMbvOiW4QElZeyNl/aAfL2
C36JGAgFiyrcPxSPqc6LKUDTQl0WiwRX6jzMdcnJ0x3+8bwEIvT/i9xEoHsqAWXG
5bSf4oUM+QxBo9GgQDz+1O+cCW9XibUhkdn9GNgAUy44r5UbQidJ6C2DVFkVsoH3
6dxxrRkLNsrKLReJEzwv28HKolajHznrtF+H1o8r+no4YNmPh62uUUjuv4NyLj+F
iK41siYWDlN/F2wG4iJKq1XqWOceGBvb4pzHSNndfhLnPO87yGQGl55zUcFSQBpP
R+fsmh78qW3Kw0wfxC4+kyNoCxvZ2HTVXIbODboZb0qMU55Iv7zN3GSUZydGwYJC
6zYNic79flxClU0DWyyZaZeVoeQ3GVSWxtHq0CXyVvFMwpD7N8IvJqEEuq4OKjne
mff8QJFD/7Gftqmg8dUJZqTjrqX8US2p8wwt0MCpBVpJqwFWqXdPvjbahB+KXIwn
uiSEQNLOlT4QPyRy0s89FtFa5KoJbrxyOpJYaZOkIwEOOspWxoF958LuHZz31TJ3
IXixpG4CMzzveVFqOQ14XA0401sx4UrBdhV/zfdCqWqagj8l4+D66XtwtFM8Kh9F
yM0p+chD3JWSac5OB6Wv/wK0UpcMjZKfGowgUhXAxoPEb5eBhdUsTW3kNmnP+zRd
2IfoUyXuMTIlJ3jcLlVa1L4Il2CNrofIlbG2nxi3enLHixQ0956YoHcUYjuLgurJ
Sy49ssQTvaw8rqBeAthvo7W+WJNdqo0yNz5XM0zTQEP1DS7kC5ooKrhorWiYHpKj
2mO1MxKGgbY4ZCKmYjPzpN7nFJ1lkO5zHdcsV0Qz9IAb4oh4jIh7/MmRyz2CJmzi
kCd6Wf8rfrnKNRGdG3pqE+BVcP+hXUnPAsIhfvme1PNyRxf7YIvKvOMRXui8oEyZ
PY3UcXxoKB8oZvCmoH4SZQeWxqwlmOJGro0rayFZrPR+mLZQJhMQ3hVv4V3ayDhE
Ru4tZP+8euNC4h73fMaYHg6gV8EKYXR1YQlmpOwgn0zT2YbIGzpf0N5HkHITOzD7
d6knkP2DZGwYY9oLJDIbngsa90z7AWfto1BLLpjlADs/iV5X/Yvw4iivg0Jk/XRf
KEbh1UWNTcd912NJunJZt8Wdj6bHCk/pzf6Mm4Q+qFB58n02kjm8bRBC3EMcnPtB
Aq6II/BNGETX2OQSdj5QKaqcuzfHkkfcRtAm1pd0jRmIQ/yNvyut7UoYCqfrC1A2
ZQRstO2IUkF6Sg3JYXc2c3zsf/y5g+jsj04U+0lZK7r4ouEbKhND7SY5x1PijlUx
bFgvtuyYj4QMvqVu1HXeM1KNwOdngh93T4wagtGVo8gi7w1RsIqizEdNIOGV7KzR
JK3LtgwCPI7XLb71UoKhN/PZ+BMjLZf8Jmn5182kMiPKEeTPsFQQNc08Muxo1s9q
w+phgJsF5SYTdO4+W+3slvKtLHuvH79lR7jTtJXVdpQUrz+wG8wmhbcqtJbER2as
8HOB4e3h9IZyoJTy/l8tJPUKDfmTCKLPZW84ZYHwNEw3YDiL41IZxMmRQ63fkeCs
236ocSJ1S+j9oTTUdF1Xoj1+uhHwdhmiiT9gpZ3eg5Q6YXANYj5BsebICztDTBSX
hESUBgfSp3qHPF6Fw9KPE0FCHQJbuNL/BOxSgc9YHYZyZ2ycbWNQoTLh8nLREonv
gEtFqsTzKyjTFNBKj0bZFvYTBxmA+6LqzDzXk6wCRjKVGGmz1QZnDXLXTW/h/lKC
3Q10wtG5UjTySfocxMofhgy0edSN94Uxz9l5nJ+Zn9iGbADW5XF4/5aTb04+4G0O
Dvqrr1E5rnytltSvPnox6+y/kqQ/6HAJKujFhTwuI/ls4tK31aOGxUhVd8NZpIqg
ng44+cxyLsfjwiFNwYVDnC3hiAPNQtI4LlQjmAVN2hoLfsEcAYzRkysTFfessnhr
6jGzhwaSwKPZVquKG72MBQMGxAoslv3CmIPqssBSNNW7Y08W1czjq2whaGIXfHcy
poB7o84xmFxQCuhzkJk2BH0p2Tgx376VvkEIRklMuCDd/c5W5AoUIwZf3rfkZxBJ
YSQZOHmxFu1W648XxEeO4QoM86HuTjBvmC0i4/6tIevXOVRMy3MI6/ymCF89G0Xv
qmTVl+wXu69IGrwK4wKe2jZALEBU4Y/NtDeex7Sb4V00UW/Az10EuE2Z2x8z+AAS
Px3idtzmK3K5Ahwr1hfbBYMHvLRCVpwEF1jEWRXsGskEz1HWdCSvpurdzQ5z/c3K
de+bF8Ada8oeKDFgRSr55n4UUg/m6AGtWTPceUVS3pe736q3NXQYG02F/Y20SAJ6
6e66ekY8jsG8sNbJh+wi/oTpJ06NHRDfjI9HRDiqWefchTPfsGfvT5gUFxcyZyiC
SuEQ4BY1hfCPsKswnLTz5Ax+wKZSLr5wO/nMCFnHtqQ8Y3BkcQ8kJxLiQ5Xvr2uW
dXMwok26ea+If+7y3k3uv5MN5P1c44oiXs4/RUmIYZpkJRE3ru4+7qvKXN1XcKS1
BMc0Khw+JhOwNPqlrZEPeiGYzauEqZkjTDqnfIuoj+Do8u1HGd8hTR6QUqT1X5VZ
55ihvJFGz767empg8eUVAU0WzMlIQr+UZi83cPSawqVzw5qRSc4CZDh6JkOd14rR
BG8GC7amGJTfD00oPgN/CPfTd+X5C7PWTsD6PB6FpARqVCtKVY+WUhXLtD52xzvv
j+K54BXHgqSk2OsxagWbDs8u6/YCPgD010bzuC7jl0kvX380EcZ6K2DwagAXeawh
f2DKb4MIxg7UJHM6i6Sgil73xCdMQXSHCWNhWMj01Pe3PW8zpqI0s7kTscptVTFO
9Gxij4Sm7h6Oi7U2t+BKtaSHb0jOOoQR00izMjYOhqyr79APCInxDg/K6JkvWQ9I
M41S57DqGGBPuSntkoHKJX8tf5BosKvw2dxL/DOS0RRnJ0UFN6wQgOqo4T0nLISV
vmFZbqlSK2jai+KqxtnPcyYPtNEBg2HLZW/tDPWXb/UiiV+gty+aGK6I+O+B4Rl+
aIWBhezZxqLixn/X5+x08jlmsCtSW05x5WLuiUzBaeNs+rKydVEwMEOC3oz3j/9/
VKYLeS6rISyQjUTFU45dbtz6qQntUlxElJS203gnVyUrs82c78tbMYWUERzLQHI6
w1IyO2GaNIy9P0Q8T8EsX6M/AszpdpLYQjBbbnlVamvvMqYvQ90wwAeeX9v2NY3z
S+ANxIX8QMTwjGGc8ITxrNRYQ6iVMiTPvMVSKtBWGY+ZjdERCE5w+8l481Vs5ixF
OJ6zpq85JQC80SNW4LRK+9sLe05/BdOh69PBFEZXPyO8GBVQtdp/NqdDseZoQvfd
vFi3TJhWqbOGQ8IjeVrnME/FYB8f9QBSsRkQo83U7FG3g8/4shK5wA/7mXWRdcGp
XaewJNiBcqHnJ2LS7Ls7uxqlHpMsdVqhQDEkW73fTVzimf2C5O9ZoC1LOHT3pY7A
bJQLvHOqEqiWTnXK5pWr53bnpQ/jD6FkaZ6svJQCutcnLoaX504Wm5pSWusc8hCQ
jw+zz4+3Lx5vaq9oJ8WU8vKPlbM310Pw9LqcCIrR7imK8ybdjQdRQ5N0plQ+va3r
hsTfwtbKdCaBOY3vK/spH4N13Tq9Ld2mxs1JTeeBhKTrJ/1L/M/vgjl3HN6822gM
S2vV4sRRqkwrtXY98Bawo56/T2VRFjExEJt2hpEFpv1EX47GecQtrc2v76Ttl6SK
3Hqv8KS+7vqtAGkJj5dtwydgFbvhJP6aEML9OV3kuqLJ5zIuBnSXVRx+yhbpjW8D
gJ23QXinwpe6AyGjkQaQ5gfqtQWp1G/hpZWyjHbVdoqNR/s4RvTGp0/oZheVQjXT
+AH21GD5+C1hfwhyQMCRi8hFfV/cnuinkpTY9p5YxtsbwWiYSI9X2+qPJaF74byE
OCXrrJWvVNxR85l2THjBLKwBoLHBQZPCXAvu7cUgyNWDzVOGck2N19Leoa8iyxrt
kmxZcZk/uuaTj78oeox9ExG022f7I4UXORGVpcKT+2z8vl8g1ySU8366O1WcEURg
Qd5q16PVod2GVpdHs41n4EmOdsueHFOnJTq5vkinFXPQxsSNrFz2t+f0WL5Ae9zA
eAP8u1jj0k3FDe5Swz5/NmUgEv3TE1kh7aKe7qaII3TO+vS00zFprJp2A1naIj4w
qb/NWSf+krfq37Jhyx10GaVPp61F5D2yxbv8rRkW+zmkeC2EdKgCJv+CancQoDrH
H0F/ActkvIduCt9NtDsMVDhEM+6AUqC6GWRAE887stYmXQ+FrbjSsOoFozvZQ69/
dddGjw+kYtfryvdapop0WOsv1qBwQ0Mj+AK0sSe+5pkXDFh4YOqreosv8Hh2GpDw
tY+96jBnHYKDr8xFhg0o8zOfxW+jtHVI9v1WOGqcl/FLa8R20U6I/r8sM87Et5KT
xgGpMFJ04x6JSBQpo6LY+nY6PBBbk55VepPRmqGbdkJWUC6h87mX977uBUF8nX7W
NtQLz0BVGaRS2qtXyB1GNrAA1KzTsOYD+9dmzI/0TEa7KNrHKdjaVhIHzaNgjTTI
NclKSWCQb1HuA1stT0/YHj7r8uo/rYy8MVHRSgjgb2QjlB+1PUjep5WbwxNiU/Dn
RMzuEm0OmjDiKLStO7Zdl/IUG0mOpJyzJXK7UiQ40xbGYcdMFjEkgIw08bkoVpKS
8yTHKRg309vT5CEMoEmB2+Q2LUYH5DRipZ7cp962kR5Zc35B674hUZpuBg9PysP9
Ah2Gm56F6XkKnGNUTh7LhX8EC1Kvs5QtAkgWHFbLXnWL/a16VVEg0izGWIC0r2dG
eDAUW+M1sDzUKIB2aPcryhfLAvJ5/O+q4hsVUW6csj+kCRjKid9pRzc9LDK9GJaN
eknYsUA4U45lKF5a8gQ+N2gmmrRFuu87zgQ8pbTiZLlYVlkYejGVuWcrl/lo4m0s
vAH2ip7ljYIqtQMNUBGDXeNO0S1y9NriY1fnDYpPGTEWkkIRM6WYaweO6ITRuR5I
/D77EDrVI89jq2C7WnD4oQ9r7dD9UoiXSDjG4wrGqoW13+iQY1kGyPtgfSjSBVOh
ZGDBpLPg1QYbD4gUTRpEC/YyApm9oDZINVP3BvuzlD81yp7yof+lhjgrshEkYIex
WruSG3JWZTyT3VA/HVB3mA6CqYGjN1GrqTrw2wrtP/s0s0IWlR0I0qiPswSUsR5L
iwjMPdkhYtsckLPvQmIe8FNetu4KUVAUSq4J8WlfZnY0Sx8FgMrq8esm2/yq/Giu
u6h+VPsFP2cBusUBphy0L7SyjszmfeyulsstH+3MlBds3Wf+Bg7pUU58bdQ0zeTq
hIYOo5oOr2/RaQ9GwmM1wIGkUg1W+F9pKNG3tw3sSwmpLSrJkyVva7zTA9p1kK6T
BgEsp0iXuLWm80mOPOWs8zqTzYTaj8GpjRdiF+/VzYPUb5STysJ1hU2PqGWrkDqw
2DON4xHgP0VTw4wXau7fTLSp1vyAvA8mzlh5MIo+TUVxSShnBFdKnuQLquqgcm3G
SWEbjanp7cV8zriAr3yZrFV22LWjx1bKMWs4IbHijo3imqMYtZghjyXgoiOtsRa/
/RPxKlKQN8IyD80IdcYBXMJtu3lLkxEawVL0J/amE+DsgeUxhokaIyjV5uugTyEs
O33nJSLZ7tK+tAEOFla5ZzC7smVylE5lIj4FAnhq3p31ouKfUKvxFculOZ4mCRYc
kdmGi/2oD0z4/gYV0zbIJPr/iJF2gssWjfJ5iAv1vpCGHdCKJICmG9IPjaPUjDx7
QugAsS407TxYPqoO+FvzBlPUdvSp72u2B4CdsnEXKGLsVcSmL+ZjZHBG+nZzmAO5
DMqlzZw4MghQI0hee+QyPLS9bcAt6U7xqOGYEiNYo46yLPOUrHcdjWT7gkMatdGa
YVMwkQDDPf8QduCY8hv6Vkdg5COK03b8PvXZBbmmQG1jGuuF3J0Nb5P9NkuO13nD
uMcTNhfCvf6y1glBf31ZXMHCTrPba31SYSywg8d6wc7vBBKAqHyM8bAn6sShQoF3
JGEzqV/srDE5jXedcYtftUYBfN//HIsRUIybM7FtRBvq+L9MNrOOL2i4IOhY4Bcs
5maTvI1ScbbzGKD5hrt2j3NJ5DYK4P4mcS9zmNRO1+pxAqGlcUl5kKHXPYaPCih1
mJyNjjOLRVOm2Z8894iw/IP6jh2ePuF7PTPpGhSGdnez6KytVG/R/VUV6/SM/nuY
/uFEjfViKMEywIyJri9zwJFQPbZAn3OJbWwpl7QLfoXNDqGabVYHiHTCBgQsKT6M
E0VzDt/1ubfqvHx6xHp2iBLBXD5balvt1bE0EUj6BJdo+IPNA/4zvUIyz3+t5yto
Wj8DMr7vIScItzw+g3cfKkz/LdpIIAoI/0MxDwAK9Tw1N0JHmwQxFkv+R1mYQ/PR
olJEkZgWVglaM0/Ve75DaY6TsIkDJ8pWZcbX3iIAukYj3H8qn3AhKbAzDZVNAZpB
esi4YvzZHfVKfQFacJf6AlzvM+sZ0ChMVctQJv2UR9Gk1YqQujKjRDGhKlb2c9UB
6pJHEOtLRCq6JLJkhBFu8hHxUQ1gdy0Y43gkQuVvzg2BlsfKbZoEXcRiQmMZB6Oz
Eu0ADGWzK8JD0DtdwNZ1yGTSjzjefXYjqTx08ZOQW3RWHBIRORLwWCgOKf7HkR/x
rDJ2pF/guOm0EE0NKQEmInFWmOk7TpaH7BrgT7XYz9+3+REW6RocCXAwC0XutGh6
D14/FwLXz92GvdeNsz+7nO8RkuCTLter9G40LuH2bQkovYcWFwPlp+ewACBrPyGL
ZS7jppmB3SN7oIBtkBhDI5oAK/KuyaBwsGu507qxeP8Wj9anlg3X7+jRwT6/geta
qYJwkLfFRxKAgIg3WXpFope4bGN6A7UVLPlX87WKEE82XzYjR7tzjagrfFB0wSHF
g31pDXx9CF/Cw8Lk0ngbS1AL47676pDimgKwoxMDFjB+LxZ0vvR+NNpZoJ6oqbhI
IhLK9J5OJITwC0vX3QY9kyXfj1gl1822lXajkVUTE+YWI6EDnM7QQ7Tyrexhh1sq
iwiuYCuTZOQAdleF+W3i5hylU/i9Iv7rK5YraCLj/UAwqS0kbdfHYIy0XFrIRynR
JSwKc8HGzA6ptieV0sDio6KrP6aMCwvH+m+cvn0x5wuWP8ze8zHSSbC30eqCZGwv
JhvFztnPSjXi7O9Z2ofQzpjfNbQVdqAWWvkT3bPCtwYnsLRKLEDoY+mbG/OSg5Mf
8m4Z7sbUV3o3UieTAPilmlw2iOOvwPubWfzYy9kZpPftmctfxmfaJrU/BP1aOONc
o5ByPe8FKl7nlUL8hmgEYBAHEg0BN65Iy08+mJ/yY7rY9fwwFFoa7Z5VMwdw+Obg
Kgx5gugjCcES6RZDP97CXZ1mCVLsFyf28p2eC6X4W0BzUyz0u4yAlglWsVcFVrDW
ptYcf98lNNKt66jVTUBjx44gA7vLkK6A1r7QCkmRzAARcoz7iO9g4GggHqO2jk0N
cONeBK6cYDG0owN8CyfpdJvH9102Yhpquc1MaXlPa5MGho0aEIgbZYg1hHfMbuDN
GtRr1m0stwV+ygoiQvuXMkR7Yn66Q61jxHHn/0KBVD/H1QtDQwuybg6tCFIjSheI
oLFwXUe9QHn8PdmlSbxBUfagoSxdz6xmEfoC6oQyfSMx776lOZGsV8VQKUNI+BN0
zfYhqcPIRYWote0ScO9NrW3cqer2qvqvaQNsrEKRhNEBZvBmUZqCwNL0BEJh3Ffj
uEruEi06M0gASShbFmdaHo9roXW1HwlhNwgDw3s0WBb2tZMLXm16z1MQaopbNNCU
K2fuSGhuKMEYNXf7xdTDb/dioqHdZvQMy3aWg2+4hnphbz1x9McqGf8dLVGbOLHK
1emGWULp2TQMTdrMudB8/h6K7r9eDVryARH07E1Y2MaptcJQw2mBLsHuM0gL5WZV
7trPrN+8+SLM5xtymdVY5UuwIj3LiCZzgWIEYhQqPTxDsliZg1dCUv20m8YjoeaR
pi5wg58Qsuvy8qYu/8vtyy/z/zBXltJdRnOKgkCKHvtvwqPALTvKg14Tf7Ervc1G
ZIR2J8+FBGNoJkrStNpei5h7oz918k5xtUpza+Fpn6KmdJgpvvUELw2CVYggf3fj
6QFrJqZu8a48Am9Dd7OLRSpgj1kaOx6USlklvwF3jf2gD0A0V9qlM/LUqsIWM86i
E8y8xnps1R0cMrcSw5rFq4HPQd00jhzCGyyvjf72h2LJi69s7tiwXRx2R3R58pmJ
V1oqRT761TRNhR139Xh1Ah/5G7qf2udMoE0uRtLlp0NXTw+CnNG7ikbXOd1Alkbc
vt3KSxAcmrTqaOolRbSH/77ywB2F2zgtFrTsuHh9219KgOVD6aL5ssEEp6kpYz6R
s/BtoxtaeLtONHwysKT8t1wtdr8r8WMutFdJje3e/8Kg6X5/NcJIfFbVj7F8a0Eq
1qYrLI/U+EX6QE/EmiFzumLVXke5Ls+iU75KApn0iIWvdRvatA17zGpG8w2TvsB2
3KX4rd5rFrriJbVal3vfDXoQhJV1+Peia0u/kzji9VRp6MKTjf5rmba/2bGfBpcn
bNsFDaZCEPec34OmiXGiY5x776YsA3KgCWkYAu8K5uOmSH1qZdWvxAu6FreqQDUH
DUV+qzmEy0ZjpvZjEIN/yJ1TAGyrK2jni66yqFrBTkWFu48nMLbsfQzM3zFYM+Wu
vO6kxl3ViYOq/rezvN91qjqo/9PALMGAqrvvOma2RJt2BBCjkdbtvk/R8xY+ytOR
WDrPnfcNkNsO4jSnms4EPV2z4FXc2k267Bea6AhzXTk7O1C5RBtEZF+MX2HFPeft
V7Zqd/9E8z4M7oVt5qhiSCz90Kr1rjp9dOTYs8GgJu4RfzTLRjRbU9VcCEqZSGjV
t2gUGCYoe10ArjdnsmV7NUBph1OLwIJAqk1BSmpVu4SRHwE6Yywgn0pcrQxAGKPg
2wrHQlGqKFcj8ezLUuQyvRoRc/kClM5PlVou+f15t67BXjq6gWsFP5z582Hu4xbn
8ke5e6dVbOSKaxRhjVwo48K2OHAQ5zHNCQHqmVFqvS1Pr+sFQM6ndo5pBcjqSt+y
U0FW8UfQ+56lFFMmTYCBJ+9b3rRPMIau5/WLvxDW+vSH8YEPEVBoKvXxcXzspqXl
U2Q65RI6FTUOw17gQnkfHggd/nL0HvvIqiRDTFmoyktng7FCY0hAwrxNTLAnHFgp
1X8AnY9RgL9FdkrCNDn4LR5oaxF61fuvTo61R5hg073YYBHu++4lmgAjO4WPH65s
oShhGQ8HGJQ+KJR3YeulVJWyqOnHfrZzyrPNFtZInbicjNIZMLggLsjBwYjGlrU9
JDH5HccR9gFmg8iLOrmpFrzfwWWIpBaHn4PKMYCpYVnAJAcJ6pm6Vi4mlLm0qA/7
dTv5qFTnh0V/vOWArXSHbtBm4xHN5fJ0KEtj3MVewIfu3ySRBuD8mu/TDJufS8LE
r2hDy1sJoTUXk/9CI2usncsdTEhUZtABSHUZHtlg36oHkikf0NBIQzHxb+i6/CTq
9+qgSmMpVDJw8NBW0R22p1HgpxkZCH3IUhUTrnKHLzXID9Q/Pf+JE8mpGMBvzJNs
+H2/ge/yVmzF9z9MtzkQSuMFHZ5PpvQVyCR9Yd1UsOlgap9+xMcTlfkqbNqOsZr9
xrVvTb96RRUjvo9myZB6ZPb3ZSdHfdDmZomFwQR8R0ANR2yJslsP3qjkqN4RlLdv
AP8zmSrwvHKVHejvp0NRIifq90KOUzvSYGt5oCXa5b6b6fFGDu1SupRIVVadcrYG
2zot/rSFfY1HRn74Zfjxnib+7U/61/M+1LKvmwx0jF209wUN7dklZsn2Wb6c2C4H
WiPEXVdOppNdlWFq2epLZIV0MXbv1c+vrEuf3tlJcTDy6y9DhiuVZ7Us7WMKCZSH
zjNYEjoJSejTUh3R4dvgSieYCrHSLYYhHWh+GdEpvnfCco5roSJ0NkFF9b5VUfim
x96n4sEuSYQk9brSDlhYCeDNnQChRW/BcUF3Tl4sAL0OSvI93PB1pqeJaqdB9Tl6
WsQLn/XfApF+Xp3ywjpAzJRvusWTCwkWskkRKWmFxAXV7tyZWrZPC0zWIUEJRmp4
T96/2K1KObM4xgC97OkJybGZlGCMK5Ms5utoVV4YYY12PinNg4SRAppUAbMMH210
nrVWVqCOwcprdtgPC6qb4h7U2Ov4JaSKso/5P2HvC5hiO5keQAjumO7Rf4qbD+Dh
TpOXOCg/N5FMDs13NwLJVFObkj4VVhfzR0t1ez43E+rNDP9oQx4gazWmqt0TbKIw
91/aS3ezOyvXRqhJqGPo5sC+Q9T10DLO7GllAOrQmqzdFFMIMy8MQTxNBWRKLLgW
TM0InlNdCxu78LvUUs1uyNXpVwz5i9NP5+iAk7DPVFProgS3wOuz3/B89XMqc3qm
L6JJG+tofSNNawx8rkxSlpzSnK8rAp5LOJhPe3iMLkPvyoSQqG1S6ihgidptcA15
e53T4Nl3xYno+07sVS2h216R2j/hbGtGDKQfi1ehjtMXv4rgpkoH6+83xRO2Xp9W
pfrsWv8JN2S0n3V5AB27pSne/d9ZvbZOxP+tppd4AJ0Fpz26knRy8MfNiYIErPPy
seCBXDawTCIaCsfzjPkCTiBu35hAEFa1Ix/aGqmqevxJUr6ZM1ezS9BkSpmE8wM+
sY7+WM7+KfHPMA52E0mSB6vsd+8bsHMY7flui0EIW1zbkPpLYlznEQ7hHR1hGECv
ogF8pJpiUkmccutL50w6ks7IxnRm5B0CRGelB3d8IyiVbz0kZW9PG6WC7DogCu7g
2ziPAbyMXHgF5LwKtITBcFQkSCwwCCnsWbhN7oSyox2ABDi4PPOBVnliBM2mS2ed
aVo0MC0tDJ5wd5A3FzgkziTS0gr1AsS7ieb5/KarLoWEETQie79n8TXGZ8ZGyB/b
jHeF+iBzNrPhrflGRpHj5qHsiv4ZGEKlN5sdYmxXvvXt4dA/hRpONnhO/Db1gLQZ
GmnBTwhzjghtqdGP1bXR8+3iR2lUyWRKf5myoAtCQ/WsKCavZWrXKFsgKhvjkEDF
qVJH9UVcIdL/qBkDyFHmXDa2brI8f1F9U9a9SmpmMeW6aDrGV1Eh9IL2ZwJ+x98J
KmFCanYLWZjOherPoasDUiUNUhZihziWt6iU9ftP4QdSELdgGp1mjDVlEWjE9ZHX
RixBv8VN7UN0vV7/lWmRZxXLI0ew6kUPDiDa3oSiEPRBW5/HjiVWlUVFe7yRxOr1
W4xk4Xfod59xR0WUnZpoEL9pjqgv/BjfHEW1gOTksQLSm/6Es7u4C7CgRzD2Lzr2
6cMNH2fxY7IsbU1Fyr8tYxx4mQelnRi5KAV0JVqOJ9AaFhu0delyTtVgxv9eJaBq
pUJpnPrQiiTTQ93ZTPM9QHdrXW9SJa56IsNXoPBa79a5UUErKvK9ltNaE8ukGGoq
cCDocFywR2gerl2D44GQ1Z92EfT1Ua3qZQkvYUv9Cr88IJAAr4iNImu5sa5+9dCo
2NAQCtcO9Z9q7nxzP3EynEG9u9o3664OD21c+NAjRHOoBvGqZKrcSjyhPlaCnrMw
tc+QOmk1QQbKw+9i5wVYav6e3m52FvPiOpSpJgLxu4PikZRkKgDqOMrXEexCysI6
OKNEdAvGzNV9fttsAUwDH3WqeJNwKp0gm1qzOaoabLH4DwiIqBCF5F3rE93+/2AG
8+7SXIA9WMF8mXstJ5Po6UQ7GjUih/GBCQvOUu/8xyabEbZ9dWsS8oonQvd8Tzf7
wUKEduszhT9XZ/Cb4zunKkQ/jEOde+/FuRX9Gt5E48WMQbWF7vZsOsNIb43HuXJK
zfOiBnRzmWZgCl+eXgv4ipKKwHagjZja/aEhTeIEfduBbu7juMUuZX5IEptyOi1U
1SWvNO4jSPwLUIvmGpn824K8GiDUhPCFB6z49r+y52aOcTS2qWeNy01iLgxyQqtp
8315pSeqObRycVZslp+6pF3iU0KegwnleFvc60kQyjZj6BCBFrTTgIHRI/fdlYDH
OerGKybbUBr+pI4w0Wh4hedx+ZwKPJwUwA6GaVarHpHNAN6/eovBYMrQaFqGqfyT
ZiHoQw11cEo8Ju4ulcL928Ix4AOXA4gsv9X2CEkgM15/tYy0OUnKyHiLqyoUMgui
dDsSeKZ6+0fDmGKhErqLCtv8mhfo4LTMPdaZ0sVADZUiZUZwNi2j5j4u1wg77Kn+
+MYpzn0OMLtpbuwpt9IionMdEyWFEdiIq4tbWM6GCZpi6GkjJv2bLRP2b/Wt4gMN
8+jaGIAKdB+iYz6NeWw5AKU4BH1lcf5xRtwhx9BrQ1CNGagKJp8TiFf0251f6+W9
scdnYwFt5raQJN9LyMxNk0HHLFWLG2z0q5xyw/bSO1eD6QjordZ+DI+sHoAtBMi2
m/UoS1oHbyA1dXghcNPH7gp9Ws5ncEY/HDZv4DE49ztNqTuOOYong/OmBbHNr2qS
qw5YxH7iHl3PYjgUHtya+Hh7esrtOBmnj7/IhmdWKLUr3GisZuUAqmeQ6hjUH5cG
L/+n+EsLk6Ilfhu9KoYHYilN2H8mkTqAxwMjric5OEyAOtfjxYQmJDL2mD15q4Mn
XZ6ICF94IxQmor7iOmGHwJEIYgw/s9bI/wyU1v7sdsDXxJugdmh4BznvMMmusNYE
d/OhChHJ+pMIt3m2jZbN7o4+eCmZwbqCMfe5KS7f78H2SlfWaH2ZcQu+ECxu6S55
zB/BwRM0oWovT9i0ZlBUMDkDL+cd8jBduGzbjSF9QDYwVCWeCRjBPaLLfIsPSVfA
pMHvjHcnWL8v0ZLOyK5/EO/MZPyYtd4aBEquEKiezxYLHh737u8aSX1d0eGQL/m9
fbpWsfljL3awHVdMmkvQGwi7V1M7v5Ze0NCDJuuslvI3zi9aSsn3pKdn7U7DcyHN
7+PB5cs4dqwGZapt0SxrXDAkLsP884+hKMZNV7pNUwMFKNNHYLuslcCu0pv7oAPJ
wG9snAlgRElZMITAJmjAMvGhvGrZ5Y7AtdJwXs7bCY0I4pqFKedWfRF3MLTf/svu
rs6xqR9VnwgLCmPQGLNqE40BODqjC9c6ibgFXoLBYzETFwPcq+MOuTe7hV3R3nTU
i8JJBE2jwFzHqFMPVAr/Fh3IuysCfYtUBZpmGLaNnaXnve15omoGLEnQKSEpp3BZ
Q0luaP323lIffpYgPREaFHXN7GRf+OFdAYpJrQP/7hjdp8UudKAeG3XbbYPlQi/Z
1Q8WCtKJQCz3v4jgeuP8JI0TYLi8T5cH42Lch054Zt4OEY8fc2O00S60hy3YdasR
ajPOxwRAdL8asolTVsMMiNmq0MUhjr+2zejaizhYRt6E4sL+62JTOASEJbxZTAcD
XECzJulqboTnh5kxY/PV1zq1lQljMyeaqJ2sJoUV+zLgguMGj8pqik1ywRRavOfN
J4gA5KHcVxrG1leJzqlN3VJ57RuYwEWy0CV6YQJ4g8cJWZQZ8KMTx3d/BE2fhDHs
ZZ2xf4uRYEJitkOlwTW3lYYLaaayXMZclwFDqu8hqybg0hEnnvnPpCQ3dKqp7D8g
gj4EqALMTbTnkUic8GAY6hSyyOqHPhb1okUs+amSonJZu6z2e3U5a+RDMP/t3dwC
NujuEH2JbtYfFo3GH+g753jVE6P9pO+dtHVyrI9dQLpZl6PM9N/Htnr+u2TlAH8a
14P/3ChEhk4CmdjpkVm0cUTOhi2eyY6bZks212TNoUREU+BkHqOyib7wqXwHMWa0
hs0VLnSLSYuxF7rFb1PhxM1lRnBMFDJyMRjoegh+U1tzgkKEZu4Llqof/V8g6ryE
lFdDLGaHlFnt31tdD7hY5fIfmIeD304OzQz3RdBDuD4hhvHgcPUbrxux1gwc/6Ic
ZtMl2+Y8wLgv0rX6zoc8Jml8fuYWIzIZoLdOXGHQgV1WvJveLBukwqDRZ499S57E
zubXpF5X0K2gE2VlkWy1Dx9Xo8DlrM7wQuTzQB1sFCD1gUBAkMsJocxqO88foNMy
55bCouwW/gorH4F5gjcRoNafDZjk54f+Q4SQESJmKbqhmBaswapLR/ODr66BIryk
8Rs/OV4wFqT4Tlb5Hml85+Ko7RFsYWMXWhA2KbZ+dASEXlp2NFDQwgQa5hd90wSu
ZRY8ah//yiMwV1jepNLIbSRe69oOsEOshvpOtKVZO4SARpKseHQY0UyqNl0Y/jFe
kJz33HhYzeLp+RUmgJApxeEQ0ypmnKyMQItQHnU2KKt07ULLUlm2PWLQRwVKZ1E6
z1u2JRSLX2OgZ1U6UxD5LtJyv+1My0HCoklrf5+gyH1KsiM2+BWaP7fqj1BljWJN
QQVaVZshMB0J9HBSHdo+7JQ4RjA/q/KUHfLjBvxe4zDqhdqBlavK5NAlOOGp8uBM
lh8COkISK8XtYeS5X74JJW63sMgaT9da0b2ma3iXC5tJZHu9gUwG8B0OToHlOIW5
L9VxtGc/SSayW7m82SyiC6d7zdDPkMKiqtEFXZmzlYHWuCzMEv3WVgOK1O4LVkMG
jcmWWWqSPstI9o66tDzjXb2srzJjcNPVRjRMtEf5OBbDN4fZzBE2xNQAGU87bTul
ngq49+LV4zgxMIw1jhVPnBG4Mst6qmg4WpHwXAcqPtdri9tOWUo4BB2ZnXDojU1k
w0Vyku//Owdgu5VpCfy9QhQVY0Ry5MZE4zhxsM7qeFKq8qAwh56C7giTqxDpf8HX
fs2VFCZGAtYKTKljS37OTeaLApzIpBWkeZLW/cT2N/0rnvdItDXQTgJkzqxQ0z57
GCM86XjWhfPZHPXFvQNxjmFcn+F0P12bGPMO1C6we+CmaKSQaJbzmlZD15sbvWXm
W4OpnrgQyISn+R6dBP6yXurLsyKMNkE5Kw0QnnvXt+OvYNb1nGFqUwCZkSO6pL4h
M7eK9lCOVdXcQ24oHpr3eoGr9prGiHlxMu4NAofCx3BLyhS+MPTe+Fx2wZcgKnYr
cpRzIOXxJFLg+KR2FafQD3dNurPdN+QFGMWzSmP2/R04rwh1MpHWGegs7F21N8Sf
RPP4tWkWw//GoPnkmRu5IdKN6+M+m11FSf8rMbrP7I2PYgMtxrNO1a5AHy330Fym
+f8rvc4OmvfcV71nvUkXHieYRqjG/3JFHTPNgh1xTr4IporQf8Na5nxdKw4hbg7g
DaTQh+mF8bTfDn5dA5wGQH0IGoboFjiEhbQn5zMPwRA8RB1a8pNgkOQK+csvLhuv
lg5Lv2IdNhKmayhG/EHo8AFmTfzbjcpEg7mw7rNKF3lPVgDxGXiv5kM/V9t36OOT
Z4HHbnHMj3mDy4Fmq16CcuBF7Ot/dHHVLIZtqckSKWDcax0sfjkad3FMnP0nzIPZ
8Q+XX2EwQquAYwUsCNTq2AQjjrDb49eVZf6p0aQQSF3Tg6QSbGKCpl+1AA/5gIR9
b/zrytKSlgrmSsPwl3/T2BFsxrFyRWt0nf8DAcyab8rn77ms1QcaZxea3nX6sRMX
Bk55T19m7ac+8W2L2VY499H2W6LpqBCtQU5rtcudKRFAuv2lljz0Ru6KXX0SZEQR
a28RVTSf77WJFlxGeksVU7YCHC/+JNQjLtpIKzCgwfq5jbM8WRX7v6AUxcLgC0z8
kG8XsNHllQdvRyJOdptOkirT1W2LurMHB8AosXrZokAjtaOdp3Vi9GtEEcFfWjwK
ccHH4/CYYfSUCZ4gU0H2wCulkNJFj1yFZCeVZM3c3T95Q8h1Nmy7ichOBm/NQ+88
QIcXquPPGb8wuSo0Xagbd7vB++dX4f6kk/vRjf0D5/pQESWUsNtitNhhml8u0mRU
0iyRJcECTfZ9fU8RJbSWHsDOgK/Y04KX4ON3UXRoGj5ChT3RntVW5rwSYxpMjohA
XkC6DKFValRZmnCGm51jxLAdkX+rZhdPnEqQNvr1R4oRNGKc6gR3vhHvBdnBcWp+
TbGcxSJMHUKDPhcWSKmKD1uHEI5gN/PpZ4RvFQ1i8X8tzL38NhisJWZVQm1YEkk3
nZV9b/RySmZxFz6OTv++/N9A/iMjhhUN67PAhrm/9Ufzwl08rjCcIrn9KaOQucMD
N0Hgmw3HqLLLoZ7jEUyjXTn47/KEvOYY1vBF1chrsU+K3SJjZNDNFvczo61Fs5RG
pT1pzvNEqnsoZNC6N0e/BgHX+JOyG3DLr5CSyx+FtB3VGAS4YT7nxnEj6EB0M1Jq
eug7gzGloXxtKIsuxCLb2JeROiEGWLqe+XXNObSxF+cG4c5yZ8OI/x8dn3Pgaej+
QmTUcmYHlPFRGizHzcz3SYvzCdKQUcaFho1ux0zblc+LBJRJn4BhPHT6Q54itc4b
k4U2/vkMx10eZjNHKhmZag3JfwxlgXy0FvAA6clXhltcaRhjXX4Yjy1QVRt+Tign
Pu1nprl7Gc7ZEncqHuMv1mq1U6hBVsjpm6S9SWPvJQiTfQ2Mlr+7Fa6B80X5t1ah
bqQshrMEBUnKwqhp7V4by+ihNnOjMT4naib1gh/rmKLOQQ54WKXJ/V/ffcJYp8o7
KhIckI2iHpyHFkWyOTFPn1chJfNovn2AU0TByrvpzWxjUBaBV/RCPby59/OU2A6f
N5QYdYdmP+j1XJiuQskTpiPOFHAZapnhrkBPY2mZvl4oAaJ3fmnBqZYDEnSTn6bB
qX4g4L8rV35he7ZI/C8nUcl4H3Awq8JfvNP55rZdeDkHVNZ8Mz52q9Fawc/51wpQ
Bk+wmjoeF9tEadpdtrE3U8vkTG9/y1tX44Y9IPj8GFxl4Fa1k7KtxjEdGcGjxbwI
c4auw7ZmFIHd/qW1tdkX0OFiohB5YhzitlJaNADPz0+QjnnroRSII5u64GRJeWSv
NCLMQ8OKK+fs76i9oZzkRX7xkE3DJL3elnYHIIfhxC/w5yGoAaY1IIxdr2PfxS02
zhmPgyPR6Zk6MwpOYUjP/IoqvGeg4KpE4nKB94+p84wGhLe6xelAjrjB5w3sKVc2
lc9p4jfq6GyBU9hzUhDpmLDJr3qw6BkvS73GqVC4QZiH1C+rQt0bGjvvDllalLA7
2hL+8WJYm81cIPYTnA1t6VaaIz34qfb6wkZt0JjrlLU4sNoX5n/8nHTjI8UmvFrz
57ngAkbWB+1XWyNnog32AlqyfBDHkNfR9svMKG3DVuW71Od0+VQzlAfY64cb6rQW
GUkxp/tS1lICfCEdHPK/X8rfJkRYmIfxPcd2BfdNkExp64Y0E/cWezN1E9mnlEeO
md82ptOhYc3g2vPFlpI0E9Inj4QoworUg2ORomXIEpwdXOiVQ66wG6ZyNSYUN3e+
XkAUMJzG4ZH3SorFB60wlD6U51T+48ZFPJtbjspwhKR4YOVukw7V7RgAfORLn4UG
mudoyf/CvCYFGgvnAKTDzp6CSGfJyhvUr++PmbgHu0PyzOApb3bwapSeYNplPniT
il/lk8P9xqUDfSDWV+qnvJysedr7IbL4XQlaqXXTFy9ZI0jYB4yJ7cCEn7QQosNp
oofUxV6jTnMxkzENBvmBqy/o+e7J3NG3WreSbqZVOb4t7XQRN46HRCXN9DXsiksE
QreJ9W3OWRMdPwSewi8ddIq0NWBUAWmJy2p8CQRDSwx+XO/3fBb5PuEDRbU+0HsZ
x3jgn/JCPAmhYZCKCZE8i1rEJSXFCCs6Oyx8DvKERbJ1x9kADvGUp9/e5J6gi4xf
jXBWVYppq5KpghfB5YIZMUMC09vSbSt4OEHbx/NZEz2yPZWMjwBl9HHW/P5tCkRp
v8KiTLpVkLrQONC9w1nFQcNY29agcxGMN7AtFHkfuUIK+enFQLb00ur+SY1KwD2i
UZlF9E5FxhOEt9Dw+K1PI/6+gRu7wtfhcNrlwaTpicSpkTJjuBPylh+Q0CqvNc03
9/AM7cKoiWTOUgLqhw1S+j6Cc8dVOT1064zDfTTOCsBhtJd4nJRZ/AmaxKUkuEks
rQIB264forra8E9tnqzbNlCdD2Ys3QvfAjDKREcgTBVCmwSnT8PDj8eOgPmesgfN
viC21kXv6+S4SibITkNTm8HKulY/FLwYaMzWOCuin9MQhYxHJk4X+xFGb+SmtATx
no1lHw6zCRCgOvnIjCwawl74Kj8c77yaH/87BOSO53yLisufsGXZoZPnt1L/Gmr1
j4ISjYRJ6mQlKQNW7PnGUmlPD2sSR1nemZoavHps0hXNN1Ow55KVRgZV7RiDfKTS
Bs/2uuw+EA3mSYuP2Gek9vCQoT5n+dz5d3ZPOTRS/F1YFBKcffwAbc5XOhq6BijH
xX7Ufa5dILXJKNXgOpaJkmG29fhfglUKwc8lhqQteWOglLazlhaM+DrHBMy1swTl
lRqvldjNwNiz9Zavjp4JNGtmV7FPNgjSfxj6GMWfToO2edmwuD/Wa8dmGYamBgMl
KRVtjP53nww/H9xJHB7rV+P9hiiymBwBt1FSglZD4/6HFHkVlrjXnDbCY9niRo8R
vdWe6WModl6HdxHWEyWitUepj8UNd9iOjZSaRJi2oOJc8qV/Vv9jTDzBY+IT4q7m
DuHCRWIOpzcCrruxew7lJNC3M/CUoInd6i7PZiGOvWGVB5eGM6OV1AkI48vL1FeD
rx5aN1id70bh0mLck3Lm+kkWZJBu4h/OAW4eI7Fu2Bf2FgrMNEiJWD7Ny1qWOHbK
sGDnM+6nLdk0rarI/lLff93b9o6G+qIiloqHyXopK7rSht4VorjmslB17lpFcm1S
yTNlJ5q2Zw5CLSAdiEOIK2Gh6mca9cOxyYnmWjtGMj91dbynsq4EmAkapGNkXdSo
Tk47nAnj1XyrG3oS72Tr+SylfA7TcwlgTJreey63Cl34KVbUiVsdCyE7sCnoDG03
KA4lD1XXKqpoAvkWGy282ybBfoyqzSfaaZ/gq7g0htJRgMSbrjuPy2w0rgd1kzk6
j9Ti5gPLnUWfg6IG8vWV70qarUft3GKUupqA9o8qqwgBsPFIb+HiEbraKV19b2D/
RifjaSibMrBloCuOVIMk0l8P+22++d15xANpArp1qypuWM0SUuCk1KKn/p+zMHmV
ulYJWRO9VuP9j7c0NOXxXvrdQrRsBuolg6jBsbejsMtZMY5uwT3B91i4lKIwK/NS
tdruksu8Lohya04qYPuX4blV+YusvTGqJf+GaomGOxlgWwbUzCia1K2uE6nNm9uA
VWE+A6CKGekOAdpkIqbObf1WLzYzdyCe4XlUuXzJYKgC10ArPUf9Px4m4YjiSoLA
EM3rkjNOvKZ4a0S9+jicRPngofDjvQkBRWz7JpuYpdGy2lQz/dZpbjO+vrMIEISr
uNUhuzJB5p3OVX/8pKDBFaYlvtB+djodLwbX6thwmu2i4sYMoalFL8BjXx2wRu6u
IGKsAomXPduZblz+uMb/9iY2NewlLaApU2OIcAZ17lVsDMUzZQiE5Tt2I/rpk9oF
VPw8RS+pkhqw02NAcuTBNMiBfG8IwD/DYVBRY+GAoeXiK7yGPV+f17CSDORdeaEx
3KRMeTHZj/uJKws42wONfglep075hzslYByuug4cZyyCxYKwql5rJnnUPLN4Cwvi
bH7A6HnwrpachJDscmZwI1Yq/R58zGh2jWcHoAEUrGmCLkAVUMpSfiUnFyzxf5Up
Y1xU70SPkvmORvs4rDfzUMzk3O2F7RbTJlG5F1iWuuMOsnYENMd5xfuMvRECZ9IS
HGTapMN+amx4O2Z7LQWCML+4FzK2Panv8vzeqlxoU+5KLMVVJ2lUqQn0pU7dHjkD
mHFhuQvUC+QG0ssHYTxU4V/RIE0Dvo1ZsGs/3QZ7SJVx1Vr1CGlNeNunyp6HVlda
pJTCopbL0y1T/y+u4o//qmak5+6TzbZc9Jo9mvCweqxEm2llMpG4PB54bA2GBJFl
AlGi+MBQD06hu+ni8pidUOaORDQLexCsjnvIkDw3g0Rios63q/jlq/ij2BpbbfRn
SJIFaUKM7zChvDQWArxeAneCpj5xS7xhsyNRxbVDtySr57t7yLPXGKLp5LPewUK7
w7JL9IaCKvZky7W+CylYumfrVv7V+5YDF3o/+Olss/2h+AU6+8VapvNodSSdsjx1
CP/jukwcnAp2TCRPPZ1gMsEJWANrn4p3fGooXrBulkRer8QNaRP/kQrd3RciL4RH
doEsPX+V7N0/2UhrNnPGFz3wgKZP2xAa9QhuJ5VyihGWMR922UezsBwQ1FM4j2ya
SXjd0RVsruxxwF2HIG6d9H/NWjezlS0K+WyunccVdYHKpDHSt9pLVqKjn/mf4JHJ
VvdGbdbkAKHhvEJb7HIZ0PgHHOElG3vm5VWjSnf37hVLGnlejdyTx/88l+3UqH7V
U5W3q3ptCd2za8xeoOjz5WQMeN25XOV90Cc41othYY/Kq5a2eDgamSgouXmA3P5C
KOppc/laNVbk7Gnz/Zqe7tYIFks+5QQ2/6pcy91hfjs3gLC56pxnF7lj/OXiV7ii
I5BdrxZqSMqDHQxCrV9mtsZ+EMOLuK1o/BYTX+dec8xnzoX3KOMUpX2b2qNAXWj9
uki6Q3RHsszFrqUkG/rKObn7LBMG+/r0M3XURNgEh9A9l4CBtoUfeui32dm8+7lb
3CcqrbNpyXCCyzerusQumJjXasXXWlvmuVmY+SsyKW/7bWJ63aUKOK7E+mCh2WD7
TuQzDXPSgZ1MpHCwi12Y2dAr2KRp2Ufw7nAu8/csvYVuB8MfVXZr43Z/OrIJJJg5
QNZb9Kg60HMHJ1yPcPmilXQl1onVHvBvVOX/XSzMw4l6DZju5/SJbPWKemX7Kk6O
OVE+4x5pKOqkFn3e6x64wj6gT/coqne3rkhABdpfqk4HoGvfybvyMFpa5zcGcmmS
V3fTUwG3PBOXqrMXEiZYCgEvoFfOugQlJ23KGznZYxBiuBGbCIhLKfXG3n/gjcoI
ZNIPZLw3U//7mOJxx1jtYXMt2fZVoG/xwo6M+0Ydv59LzcvRtgXpBbb6ieYZ4Kav
27F5Q4FThPfYH93WD6oS4Ge8LMmtChhbU+Umkwl4LdU1s/g021/aB5fFklOWxPAz
kiMYhbS7V8D12/Nr1naKsjJ+zAk3ive0ECyqsGwBj1ECzkdgh492kvYZOpUuF0J+
iIFniXaTEipuNkNSEU34gvKNfKYWYldXlltzu1oplIjBMwZ3KcDzU4/wiaDKKjCB
TtwZbbj36/nMws68Fyf8jJ7ka6lLU9cWxcIhDohu7SSHjqJpVi3BKZQVGvNmF/cv
BaMvUdddobjSCDx9+fJg9JAo4gMXyWB0B3p93rYr/butwdQ7fb+OLFv9Vmffrsqy
JvzSm64BohkmWcb3wYldU1tLAQUKQsbOcF93DNW+zrNln8daLIIe/PDIYmxbKOFc
WYE2s3K2VHLz/OcGN/bkhD9r3DTn3gdWn5hfU7aXl9nVqzgS552Q4//cUhPDANCJ
SJYBxMvED5SESBf2ZzoeQKrjMNH8GYRKCjqQVyf5Jwkc4YMKNUiej/xRPXndA3nX
m8tONjdk4069fEEMgB61c9XBtwWtDQeGRnqNZoXTGSWYTHxDFVvS1dWxiXykLjeB
vd9c6ReYeD7xd1+2llkJCvAjKwMP8u0R8TtUcHQxPve3g8MZtHyzDIx61rn0tcbc
lbgqWudgH86NCwvO0BV6slHefRkyzGqVy8cNkP4muR7B6wq9wuu2bUrx/tzP8Dgv
jW3Bqdh6am7vSdxDR75ln7gU9L9MLz/iP8qEp26sG/5/Ss8c4Hs39We9538K0wNF
7BrDIa8sgRnl/hGdlTrmribgqUhItFys+SRu3typcXg81MtRIOussq2lTD/Zux4n
ACqoXX77EgiqrpUWeWPksj/OGPYhQsWAA8mtHB/rckeCqfw5qP+f0MgTIzDURWVr
od++SXzCa3tD1LF0CzUlw+d5yJH6hzpwVMvDKko4FW6vcC+EAjr0kQCuJSNGqXpW
lPjKbpMcXR7BMeXxnqADHrYlbzv1VwUyc0oHB8aR5V+l9Ibv6Jp8J/qFJ1Xuu9/i
LZzWPApeGdIkr7n9bvjx9if/VdiBDUVzjPieKNKDyUqW0RyXfNE9qU+GQNJbmjfp
kiHK5fbS3L4ZxNMB0ZY2FORuP//n0wY8t53Ti6+8VL56uQKy1lRcGNJjgGbuUOEp
ns85kXwpVaXdzA7pBKAH9Tuj92dKPsseb8NyQSrzUGfLFqYr82aijfZ8i9Mbj1vc
TNDfvScffOb/PWOaSGX8r3NYiHtrFGMdVMM3fTA76jkkyDYbSdLD0VaG6BjvQnt4
bRPMyY1ImAh0mHfdRb5BjfHvnP9tPFmchOcQnU0g/ccOfYXXraUrBcX8QhG4b6wK
LCEvB/n0wei6TzldKZrONLlrAOi/tcMGQ8w9yHx/6e6/SxC5Vg+wMfy+AV8woRIJ
cbRMs4dhkXpHTaqp8sV9PyzZU1yenD0nPQ5JszcicM44vBH9rmAMROEZfZKPjqyT
MCIBaNyQRYjTTBuTlbKQmfTsjAiJwaFKwJTAxC18nCBmAwNoit5BLjA2pXri75tb
PfUFD0taWo7wv8GtpHdtxkfQ8huXP5oRCeQPH7pgv3g5mFOXUqdEgcOwG8JrQcFr
c6K4xOmzvvgniGtFg95A694fMU9VhYOTRzWz8MS4z0FHq4/1sPXyHZm+vfVgGoWJ
CE726fpCzhA7eBEU5QoN741H+qx6GaeMkFcvI/OZOvtawr+nIM9q00R92NIHh4mg
h1YOKva2MseDba+dd5q4rg1Jw4WFDzUt0JyXNywPpKrI6/M66nGE98WYhTG1OeMT
HmujXYyz1AyLQQszFN44LC/OOXgu+q9RwcCf5nVjmYu39PzkWdyMHq/NX6GmdN16
lBGg31ytal47MqgoeqQxJ4M3Rst5wqOoAG+b8cAYZe++5ra6poDelUAGV6aBV7R7
CERJiQJpJ20ObZafUGqYod2jcKnKlH55zYMdDFFWzFRjtL+2g8WZRsiLVHAuti4A
eo8O2SYfCY9ifHmwy2XJAdvulfPw/AtbpQ6AE6XeY7Mr56VqYYW9mq4C86TihEUS
CVhXvNQBMpOxxrtSkMHKSkIa2rXOWYTKrnRmcf7L54X9WnnT/s9VqzsYIIJJ5+X+
EpF94zile23hmspsnaDC0mqhgVFLkXlyOlh/wAdxCZFw+qNdIMA09FAsWJK2MKXL
hqFfFKBR2l4s9raHngzn5OpJlH8VZGTPJWjQl2x9gsja3rBR8OMUmz/Nt9zjG4vW
TAY0IaBujxED58lPoRDHQmAKTQEu2JtZvfaxcaw9Y5P5SCU873ptG4NNO11PG7kk
z8Ve+cL1JsFk1a3ZbTDp5vyMNTa8anZyUpSiTJNdwpUNn9XFE5h4rsD468FQ2GrG
wrXowDot1UQVgerioKq2nUINaXrNPyFkR7C/zgLM6hg/Bo+dq3hommlatqos4VHa
rXf8+I0mYd7LWm1MZ62F0pE9i+JA49Q1QLQ1DyVa20UoutFbbOgVWs43HyCvpphk
s5+Gp1HR9rx7HqQqFXRWjXLK4ZitAUrmTVcADXc9Qe6CzewigAsTjcbNuSDpk8j1
tliDokWLsabJmOUPAczHmX1UFs088N5b65hZkMdKj5T/J52nDA+HiaPD2XFrRZvD
LiSTDg3gUwWtEv6VsNmsQHBNl+0L3lgCK31J7qwJ1U+SDiOtu3Pb2nLmOl1EHTi9
wZwL39x39H28uCb5ssCrwWXo3KNuOdtmjsU9zk0cgcU0ZUdMcqqEV43wMtHjsI1+
i4d7P/PRLnxuzCtUTZh+8eSwK6YhjSlWp0FGdTLu17XKUc/UyzSKxMAVwSDntFEi
F4FRJRlVGXCVluPYKT4oDLAhvBmR0UHCi8vG4NNataBFwi8Frmo+OjkBjzLC8S8D
lPw7ipVnRtC/Hxyhp6nToYWF1F8JBk6PeG+RU10tNN5yPGVyoZZTSxEqKUQYhJWT
oKcJs+/AoO5kP1Q44qP72MwVcymiIYN+YRkYH2qa4omnRAM8uRVW39SybQKH6hsZ
Ko4UAd7EDfphIEIqKwhLZdpE5LG8u92E+0rri+vjfY/ZcjGKHCZZ0xGsM7FYfHsa
RITwGxVH3lzjMZNsb62+X8lsZ7+kcUyk8NDdkDVkdIT3Pmp11086+GQSiqU0Z0DI
8FvctKyVg5Iu4peRbE7LoBG1LrhZCS7n5CZsF8BmKnLbPnPn556WIcReJpazACbX
T38zrA/qtKZSekpgXOJr6mQKlAznwYanKH16jid9RekyN4l67jnu0KGiMuQgkhrD
9WsC/ycQVdoHuS4zbiJq+dLmspg8egb5M/RFqDtDE69iRTZkr6Ifms4XzlJiBSU0
lphQSk9bzHs8repdazQBx082ma2gLMXw4DE5RXhNOfQ7QKaWsguHukr70woJC8gT
ux0DtHZSLu6vXu1MuOZuZj041BMNAFh73wwlcO/lg03roVep7zHRCikv9STc2SCG
R4PSWXRHVdeF4bw3NdunA8fLoy/c4IaAGXEPUfmFOuJHjDM+UbA9X2dDHUsfHRKN
MxRhJlIpTgz/654Zr0AQuiIrIxQlIkRfEAGOOImCi+bhFjQQmqyomfXWdihitqaM
L76Td7uFoOiB3MsT/S1CA3HblX3XKpx1BHbzP2F7FdgYbSsand1o3JRhJNgm9yJw
eYfJXri/e4Zd3ZoM6XujN6vcWLt0dteJ58ZjwraVce/Kr4WiBZfeGsE5WiwwQt3Z
UcW99PDMsD+RtN/b8uW/XmnwMGZwsU88L2UYHix4XhvAUUHqLTnYuPaZ6eXaMhXi
o2GxRbBubf90Yc7785MNRu88cr6ypTIlSJI61cJxgRKIqs5MzTHOEGbX2cW1pOnN
1K8gT6zg2e1Vn8ikrSn1vM/gEBh5jdNHCtSJskq755qxXPnGs/X6rKUpuI7oGSPC
UyGv4OTPRTUihl3B1pzoVSq0fiTdw0JoCRAS0wKNlaCPPw19K9TKW/3ZNCFYV7QA
DaledmECJ0cEuEynUvjqvzo5nZo7eyDLDh6WArgURNl8+S2JgL+9j7ilSXxQGFrD
dtycm7RIvY+1i9q7JnyygSPbiFzaZRTZTh9mlJtnjqSqFSdvu6BnHuQJ3HJgHuxH
bTsGR3FCgX1LLGt67Ex2IIt0nwXWpjOrMY5BreILFVwLCO0EEu/CFBtGwQY3wgb5
3TX7U/561ZIOX1XueKh9cZSOu4iYLuj+kPI0jNacFlpzPLkxw1KGwiipxSL1W9UE
g1/lT7zZ64LtNNppZrCh9bo9rVT7lWAfyA5WMeGgrR8LiYFCZY7tomOx1jbFejq0
loLlKMhGhoP85sXF2UsXjFRAgbGdWf8YmvIhlp0v9J+0Sh5rLrh+gc0FsUG0z3DP
7E2ALbuWWNShd4wpDqgaffePUUrAIa7VXScIaUwmpzhglpw/bqpm/nqzIH88z23N
3jdlMmRNx1f6I5OUdG97LcZYp4MaiuyRPPJx0Xt6hgh3NRQqMjRAG2naVIDpSF1J
wLhYlswRYzxKJ82rDfWI7tH34HagXiKd3YH1gqvdWyAycoysnK8Gb1RVgp7MxY9o
SAXw1tjZHJ0nMlRFCaUcyLqKpJyqpEmIYcotPMQyRIqHeWaNKK2rniCpOD6qn4id
1+iOsfA6SJLSN+Xw+Qt8Imo460SqxbyavKzNCFe6x77Z35/DP4kbAQsHQejjSRa0
IwQQ7Ltnlsd76d9PbSE2gOO4mz/lb0fFCiF+4Cp+wMwqbfdElF+YS3Vu/wma2OZy
oSq7iU91lVUaPvLxuvN+1Nz6Cc866Zc+NW16jOjtLL9jSiBEZM9B6a09HGh5orjk
EGhGtLvGLnDeIlaj3bCcwJx3iTG6L0rFcQuaxRIkXo+hDo0lp30CJyNjwRdnrrDR
DaYi1rLew8kqYC6YIUuwYKuoOzpgQkbBfHb+wy3UirabiesZH9FGiH4P32LxFlxe
BvptcqkNcZ0jImKfvP+x2oIgwLWoOVCyimjTpE8GqlhE/QcrymGU3OfWifnLGWyw
sDFm8SYGOG+LZb+2RkbP4KvN1AkxZAbvcD3ETiFM06y2GOYQ6It9jJ8T8JdYMr8v
Gnr21TdEf9WpBebBqYT+H0etaRuoUJebUfVum7i+EAFbuUx41uaAmO2bUtXUC0fA
YFof1vMBclOAVs1pjHruq0n8pqhLPu2my7S2aFsciResu2PuyxwhuGEoPrk/PNBg
fXJhnK63sdyhUX6ovExYnxNLBeAIfySe7zthGzqQkmQCKdb0pCsPWI3PravzFIVu
0ARt1AciLGaa8eqXW62JpK2tvKcbDV7d5Qq00qMk2SQ9ZP7qHbrt2HK4wMTgDCBe
gsWBR29VjAm4E8AEjmHF+ARjU9W+qYge43DqzvLZA6o0ppwPvPSV2hMvxPFLneHv
ZQkY1lB15zabFEwTYSxJV0DilVZA7zm+wI3K+7Lxd1cklehBeg5bw53raGBQZ0Uu
5Z3k8IyMLpAd31h+6crKokO+aN+1QEE7EDe43Aa5nYxkhJXWU3pzbYi6FolcrQIs
eZjOURoCsmwYZoOydaemncLcWgzmFygLPHg6UnGttC/l1WM5TulFHI2M7kIPZJHP
mAjRLS1AGbOkGnjdPWPMKcYe9FjcZA0ZchPm4yCR6r4dOoiTblCV5BDIaqTi7QMt
wa6utyi/5ORnuu6EDkKEF6Rdv/TieeA3xBXzBKkqzzFaKW3Q5PhYHZbGcu3yVtDc
nCZFXcSpFPrjZVKZTVMmjHQi6JVVhZM5GTGkbdTAk8QTa52AV6ip0lvg7rmHlJH8
A+xQ7lBMvEU1tVTiGtlWUU0QnR/7va1O0TqSfz7iVE0pyjLK2EzRHkWivtma399N
itdlXjOZfu4E+XWaH+m/BusQIWOgGmC/qEIma3bJiCYxMaTBkl3VYpo4EM5brfVS
Ev+FY3ZfpDmcyCCnY0D1ALtMxAHGcUe4CCdrT2n6geigK4eJiCz4bUwjhkUjA8LA
3QiL3QVJAyjGrxr9pkSAeQGqmHdpTCjK0+Ut9ASi8O7F1WLxvRGypUoRKbXxUVwz
bZCAPv1NqVvyp8H44AUNjM20JlrsFx1o5RccJR3Q6cmqOj7VNLIlrcO2ejTbiiwg
+OR1adElHoYTkP7QcCtTD2o5EwDiiFHwqU0Eo9KEpmk6zrEpfZwqf0zq7GK/NPaW
AJaxqA/4xkaRGjH9uLq7rPPDjh0+ooJtfj7MY6/sDojzms0w1gNuUnw2WkixC5Mw
Waw3f+u7nwEswpKShkRNkyNtfzi2fCvPfX6dQIRaDw9jq4ebPgX6xn6nn4bBEZiE
p93eGacBbTpeBkUxkcKKzFuF2w6LYfYYuWgs9q4CHhyeJ+LB95Uhkp2BBdwwxZTZ
BIc2wdeS1S4xtd51ey0LNd3y12xDlLs8bcAlIwIuzaZYnGVZSHnTRapFQGxZMrRB
O7PbLOh3/NPr68eyOvtWTEkZkLRLOaaMPjGWHNf5ejsunOVkbyUBqYIDYcWSkmSx
0VIyt9VILXm6v4YkkvoFrL+C9zsr6baQDcBM/iSTdanMkMZQvozqDv30gmg1PE1s
PJs17G9RN/5akC3lXEcZixg7RzwY6V6OrULyjN9zQThdSzwQhBRjNKbM2yr/VygG
yTNPvUbd0pJqwPcwsJEPwWByisBp5ZLoxrVz+bcsOawy2llVzMisubDyqzjvLYt+
kfsiL3mmJxaTcGTtg89IchnsOrxZK9njkZsH79jX0DdmriD1KtCQrs0aUFyQLDzg
BsmPfMuUqnWxBoqXIhjuxck7Qy5ywPkbkhHp4fDSi7x7qPCKRO1/TqxoMhhw9o7v
VJnFOpy2elGqM0NhKliyUJuuf/3HPKCdUkcVScQPit3a+5NCNtsRKqfkKsM/yoWL
8ttWZpWZhh5VgYitHVF8at0aK+mqwp0Xd9ddXpLqt3KsF6KKEu1FmO7UP+7QR+s8
ZVRRSaQI9TTDbbgOP1BT3Pvq/F7z4DUHFXSZmBCYAm/vm4GllGeUsr76lPcfDvzQ
Qbj00n1WTc5i6TR1Uyk4mHLUB7gSwn4HwRrueyAtp8+L3DG9Pm2uIv1fpSuWk/wT
Pw0y2UQthrVEqRFTcfzezAen02d7JkcYAaaojWxrv4HO9tgOHWFqG2ww0YgudvpF
qDqq6bvWbk5gbu2177AgEjdjCGIxGUX0VGV4CJi7NwWQDhFUqYmv3kTRUH3WKyN2
Q2f4oXGT7Y758WfqRTO3bjvrnRliZCSv4Op03aFTvkmHV2oibWlV3BSRyWGCtyGo
ErS5ZITnsUx5toLA9G0/Nw3sn1tt42GmZxHHkiGo/JvH2jKQbTK4o6yZTkD2kGUu
CLc2mZzqUlLe7gfMz1dL0XLMioxmEuY0kIwwcOzvjD5+eigNaawaZ05qWJ97Pb5d
St9oHKVaxGjvWNw9BxrQCAEP3CQZPufnMmgzmwoMtsvIJF9tqVImSfYLeIlMkFk6
8J327iHgOHoOEaZHI2r8VhyPno36mDFyarmK80+e+SrTevW1WouKWikqvvIE7A6w
C7KFo8POdFT0lFNRlLD1AvXm9m40XlESEWCl9s/ttJOhAYoxmuMYUO+mPErVwSfD
X4Bf0WubxqRmqsZOfBacGsKEhy79vQDbZYTqrYmYGQwxA/GvrpJ+PDHh+hIXzUd9
StqgEAb24tG6Yvh/elv5lyTM3grZeNw/iXyRbsWTDxvWXfs+YazuSJz1MSKR2Oyx
iJ9CQ2Xb5omXOCJ5EdLEjUgWKaWz+21XDJ/QW8qMsjtS52BQuqw+1G2f8ffWKxcs
DPwCmYjvQVNVYxMSiGb7OQg6IWYfNkDWYen89OoEy2x7OYohX2zO8ASIJ5f3TGjD
5rs+uRxm1f6Szynuf3d41GbVNT9mL7RyDPD1b5SQ/7/SMRFDCcOhXRfWJDmAoh7E
Y0LbYPs+Sm8ZzQrAXBs+6GBbmEuU0b8AIT715yF8hyYq7T9+Va8yC0hYKOpDSM0S
V40my7tUi3jLZjjWC5L1LJYxezFB/0IUrTxRgEBQP7e/sZ0QRfYE3B4DgTGbAeDI
fFcqXE0EQ3isrG4BdqfKSc6VEgTXyn4FnhA+fgWTEiPmi5hsd+oqiZc1/iJsJnmE
KkIafBgqxZ08usrz2enbJg//554Lk12wwXhwYfh4mZ4bOVBr2VhNMl5GAewELeS5
QEYL2gH++t0oXgyOPhDXdTAVgPcAz0FvDTHRTGpi3+pKR6BcqUIIbKkf32X3y3Da
CxMqZb4nY/J7bnu5D7FhkByBJ0IeK3zzkuk4bCOJl3aBSC7AhaAFh4VTbrxbuCUf
1AL7EaTycWhJiVuRq0PFFu/8pW29/fE14K29PYlrMCvQtQJpZGur+6dTdX9gkh+R
OX/5P+pfimg623g/3F0n+ZFaS3lHznV6iCizTSXkaGCUqTfvOthIwVL1f1BxU9Hj
rvJ/opCTA0wvqWX4Co1PO/d346GO7MjQJMkQJG6lsH/yWR75+Fj22VsOv6igWled
H3eHRV1CLuFNcIJ3tahOB6Jx00PBsuhvS2oGxvzljgwupOyImuJU6XVKpkEiKZM1
eQbmmSxPyuX7gkhLrpNCjMr8BSkdhlrMj8xktZlwoJVn/k4pi12uqdNlMtWVnxnS
19PnfFhzbmFZFfqHM77WGAKtctHNIhRuirZjl/ZIp/1fXhR29nHUqmwtmlYaP2mO
FeCW4tunuUaeXrTJ/Opu5MFXWvi+h2lqbOHYKkh4jE/MwkzwXS/1KUPXHCB6p5Nt
UOwZXtg/M6ZuJy13IkDE3IfjeerR4Li9afs71jlcrhAf/6L2spxunI01UWuD+Jcq
dXqz5/7udCRv/LUA6QkiiuUMFIdcWGft1Vs9XT224e+ZH1ikSTVCLYxz+H/rlgn0
sS++0KBgcr9um9lOCk+o5OPasUarJycZD56pSJdJD3wXsinZBIgWSOP4Mcx+XwxV
QnUH2JwamH482X3iPQa3x+13bfDQh1GYWcV1QvlLDQLfPwc8F0y0Y3jE6caazEMA
l3IfThSncfYLWPXjGNuWY+DT8uvTYpWJLkpb6uQmYpaswsJO+tkNnbT0egAArEmv
2TRdoZAPdMaoJhrwYJg5BSMBUm3QNNpSl3M4u+rRvg+ZNsHPLb7xIvcIvXMKt8AB
Hw6ORxAY0ONH/KotFxamYtmZs0I50wFsEuKuQ1qujrfpujs6S1iMF0fOrNdH2Xno
1BWk7LHkE62jWnkREraGn7dqjidRr48SLsKMKBKuei4KoL+viWpUXJj7feQgzTeJ
YEkZN1gQlgg50e92KNxZ1rYAYPUNxjJwJDnfusE8swiKf72959aDCXBJUeYuruJm
MmWhK3nkgbejvkMkM02PJcC+Ue2PgVDId8JZt9a54ujIVHb1xmiZi2xqMiQUrdWk
KGatm72gTHNC7K69qRVKwIB0vk4Ej6f55a4jMdJw6iZNOKuSYJ08cSmC5VsqlQkn
KmVXgk0WOICslnLT/W0BpKOfSaTplgo4CTfCk2ayq5AVJ/4N0a46aos0a5azdL4G
6F4lC1X3tGkscRBwR6CFLiXK46jU9I8z6AiVqNT6NA47g0aikQ5ZJZwysM8QPuBR
zmovUjl2SzJjZn6L8c6MbVkAKh335rWpXF5o2aDfQrckmbJxL0JT8v1J3K4QYo0i
ZYVpz9z7lp0IKviNr1460/VlDxAbIWqe9g0bX4kGjqxKs5ZvjHxJw2c6ySPH9fui
ORB/3vMb8tU/+dK5rWX9FENtFRvABo/HSZKdErdcfHCy69M2yJF/xywQK4Ch3i7Z
SqhN4qi3Jo8BCdArSbxEQGh7fgDykWDntsiYG8zUL0ZeNsDx0tp8/YRTku1CtZub
TVhkHqyjjwVmXIevUCyKMAtzLOLaNjr876F0I4QuiO4K/iXJY8RGuHSAgtmqdABL
q911jhWgGuCD3dmqr5owK7maJy3C7tTG03EByoZ+YYZCfX3DqZXcUG41qtI3ffNj
7SGjhZ3zYEKMlf6OrDzEUu+Kq5QAxr/x+mm3a43N/ECg2JSiWu/CB+OC3WbZBH1G
GDZVaFGhdIPOYJelM68lw5yS3JjcUULLAlBNjikepxCItaqZEeMQnrdwX52mGrcK
+EhbMc95vslO+CnYlMgj+yv8dF+HBssEOSh6m+d+GvTlEBWEgLTeppDATnnIpYwp
YvdS6wZk1AIpJQkg8DGTp+eaMOAhc8R1yTHf8mAA3RKnMnn84EGPo5y+Ac1iiQzu
mfsJjOkv/Go2MwxLWtN2K05qwFWzl231Em7m8xYSG6hovoNXYCGrKC+IvPANFwkU
8HudqlXXAtqoAPgw+Bcryir28Do5c7STBCZx6V90RAUS1NN4dLQuoDqt6wp2SZIP
q+uV8K/f/CwW2FJMV92IqFmj2t1uIgny2GGg7oaFlmnH7JMrCJ4en+MI7qbch+kT
l4oD8QJI970oFyNLdgHnJ2/DTicCXd1x43dFcjaGMMQmBeRZ/+vqQ30SbgiQz/Es
9gNeurLjs8XScBpF0TM4dw==
`pragma protect end_protected
