��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��o?�x��@�1�7��[�.�☭Ҝ���T�2�h������ZP�I�cN�نUƃ�Ѱ�J�^�q�N�#��,�>ɪ,�<�P"g��9���*NmG�X}χ>o��B*��b��ѫA1�O�<;
�����V`�ً��Q����B��^�z`�<�Og���l��"�����ȡ0&v�S�V�疠A�׌%Żx�ud͆�ٸ2ށ��!�SL��n)�G���wHil�� `�� �ӑ��A*A{/�[[�\�a�B���A�w���m_�lr4�KΠտ�#�_s�����X�80�p"���b(�f%�/x���C�Ս$��l;X�WC�+*�1i҈��8���� J�fQ�U&�YD@��|Jd.%���#�P1��8.�T� K1�>�@I�@�{	��y����c�o�`ǽ�	�w�:�qa`/`��\Qk=�)�>��� ��o�`Ո�w#n���m�-օgq�{��I����	��f8I���E?g�<iO��C>y'Q��Lr��+|;:=9�|����[��C�|��ڴ>U� �Y��lb5���^��쪕��[�?>H�)��c�ɯj�;�3�>���3��C4ZZ+EoVϔ8\7Sw;-�Hr�'_�*rHx�H����������pfڑwa�Y)�ï0F�_�C����Ԩ��L��H��j�>\��}�{F.C�3�"^<�]�oWq\��uu����y��66�p�?��Rr���g��r�c���(�F?�Ry�T�o}s
�K I�كlq��ʜ�a�f>�ɹ�s�ոR���3ԩ�u]t&��w-n��w��3�q� �e�H�5+��tm��&�����h�p�1���˿o=�~/֬�1�l��^��4;'_�0�������ހ�Sc��&z	�sф�S!K
��
����~zU���-;m��­6�]|)&9F�x}�u
�Z/�����
X�x�h�^��+��t�ݯ,�?���k3��.s2t@V֙�VZ�Pc;E��ąp��i��� :���ٱ�=J ���-�h�Z��y��Ň�u�P���)���s�>`��1�s����������ﲚ2s���9y?�D;�2M�h�j:5F�8����nJJ����cl^��c�HS�B@�PT�N.�b��l�Q�[X�h��0
�U���皬�<�;��w7�(?��I��ܣ�Ȇ���Ų)8H�e�C�|�/�;�����[��t���-QIy	[*�$�H�M�'�1�U��%��|�2���$�6��)[xKiV�ts��c���zY�g�g7U��FTG�~����:k$h-��"A���3zʱ�u�����Ob�h=�U2�t�!/���K��jOuy��Z�����ݞ��b��_����8��]��吽?��#�ҲuX:XH$D�+"j?��e�ǳ�w�{r؁?ߣ�n��-M������em���G�IS�z��`����A�Ϲ�Ds�h%��!���9���J$�HP -�2�z�9u�y�ߒ��*v��Wv���-� ��b��/MjΪ{�Ճ�Ur�Cvƌ敽���Tk<5/-�[��yEN34��X�������`��46vGzc��YD�ޝ U�~��i�(p��~Ɇ��8�!n�>\C�[OF0�k�h��n��w6�M���
���~|g��0�� ��!��;t��'pe�avH��r[��K�3)5��!�{���q�e�m��=#��N���/ZGVM�7�b�m�,V�Z��:��(�&+^|D�M��5eXf�����_ CW���Z�U��`�&�c�����mr������4\҃��P)}t|Q����xoӋw��d�����$٦X�&�u3��0�v<c�-�C�����|4�L�_4�����L�U���w�TK�X���q`�  ��ϰ�.�%p���s�����e������=BW��s�'^b)?��Fؔ��]hÔ����~żj ��*�xa����,	�2;�M��F/��k^�����"#h�U+��vN�(���2U�5~��E�N�E��kұ��s�;E�^]��h�9���.��$t	�p��z���ʼy�eݭk�/��i�M�WYe#0�Y����<��-Kx0DK�1�Fq��5Uw�S��/gC�3���u]�`��оݹ�>�&��1b�S)�JloԎKn�;�q.;��W��+����Inݥ��gT۽�1����v�0͓Zk�R�I����t�&����DX�dCn~؎xb}�芃����Y}J�����"��JJ�m��&�E�,��{=2mp��YU����d��7�˷Yi��C��I��&�v��jsSZ�(4�~,z�S���_re*����*�>������j�5���}|K�@|���Ц����Y~R�$Ď�,E�\Zn�xt��|��K#΢7�QwK?I���N�u��g]�LgH�J��:�_u���5��}a<�bo�o��3T�4��E��R!����Jz�N�B�	��8$�r�Ew� ّ�s�=�V<�È�˙�Z��}��0wDP�.1S˿��6UB��\E�s�E	�Y,�@�������׺M�>�;F�_2$�ô�9p{RN��,��h��Ic�`���	36OV�"�l
�]�薜���'Ys~���[B���4"���^��	o+GBޠ�d�8Y�l6��1��t�gQ�S��y��v���[ADW�>�=nM��afN[��`?�������{*O��*�+s������tqC���@����2e��5�����W��4]��O�Q(2P�rHQ��d��:�b�U$��P���+3�	�XN�\�q���{�����d�O4��	�9[�wJ�Ba�>K�	E�$��4g�Z��T�t������'�.�MB��A9v͙}$�D� )�)�
	�t$�*��ĳ<	2���e\��r���Z�0Cy*�2/A�TCD��,�f�x��	����8��]�W~Ipd)6�yF��0fo6��0z6cp9�J	���i��ou������"�4J��U(}��������E��T5�e0ż��2�o���L,r�)��J+��e�N�9/��%G�K�VnI��9��h�e���y8s�� _��E�?�YA(�^50V�y��{����0X� d�t�;A��=����O��Y� D�&��2;!\�G���Zd�it��X�񭀃IC�#�MEX��}���讗ԫ��z���|�J��]Ť�m�z�h��F�
Xv	��j7Gi?V ���IN>�p������mK�� �쎨\��L{Rږ�j���@�0ҕw�:�������:ِQ���C��p�;�[�b�ۯw���󆀖��'�(���z��$��n`sF��a�* �$��Ŷ��L�7�^T3�A{:���Ky��x�l�`M	g���D{�1�YE�s��]Mߞ<��|�cȇ�9Н��/�dI\u4_������P=�Y���L�����N��y�a�MDw[N�����"-��w���B~�î�!�6��y�N�$�r�0{��U�}�P�+F=�Y�#83�`�:,�0�͋/�.pm�x�/�@N�D����@�0m�v�)�5���m�I��}R��`)Z�Qv@C���}V�ck��n�;5ꡪ�لI�6�BIે|�C�C � �@j��q$XE�B_Q�a�F��`}�d��%-�p�G|[�9��ZB��j�#��(��C�W���I〧��ы��ueu���͋W�d~
���K���w���,����7[DT��L�w�s
~�!�����N939G�'P2�Rf���-�^�����D��m�AqMq3��ڀe,I��9u��6A���j���3�Z.�e">�5�p��ym�-zɢ~��څ﹊H��vH���.B���b�������;d=C2Q�J����Ţ�B����W��L�;)��4+���Z{�����2�D���"���BLQ0��(&vE�Y_�ېI�K"��P��hi{Ȇ�[��tmP>��p�1?!&M����#Dk�,�@5r0�9M����4�Ņ<m��:�LCK�y-�c7���@�I�oc ��(�H�<��h�ᵓ!�`rd�ro��@_\ɐ=uI��ß�n�fG�	~{�kK������ľ';Ը�jGT8D������y�z$[w2g�OV�Z�[K`Bџdo����bᖺ⥹HSXE[��Ћ���;��Pwl���?��}-��h�ިy�g��$�ß��A�^n�w�Ԑ�G�����w�J/2�H$0��&ѕ6 �>q
����|���]��]��X:Q	7����h9`#�e��QA�z����Ꝉ� �4��������^F�AFޏ��W��!�b(��9����_�ɵ�J��D<�|h��u�cD��@��Tؒ�Z�����j6;�K������۰�%Q+TD�����G�	�Eפ���������>�A����?��h{�~���5��{��p,����k�}�����v�kX��3Q
+#_N^__r3�A?z�O)�S�;����5E��Y+;���snq��4�o�_`��竪=l3�Xl5x�k�g:�R�;����!������qa�t�<-�y�H?�p�8/����L�!���!�ʿFo|;WU�9U���8I��Ta�5�Z���R!���!N�h[�ٛ��PU��2��?��I�j�V�����c}��b�#܃dAS���x�S�����I�@���T����
��Ѳ	 Z[G;����U����X�)|��v�f�.���qQ��+JmJd���>>8�$�Vp�Z� ]�n����]����[����D���P��,rd������e�Zqc[k,� 	N.�@@�`���"�)��'�Ӿ�[�!OS(|K��p۹�$ VT�:�|w���ِ�K��c���uy73(F0��i|%���DE�,H���i�-f�(G���G�)W���z��oE� ��jf �pDU�t�0l���Z�W��G��șH�#y=jXkꭻK�B��sNEMew����Yu�J��g�w��5��>�M�&5-�Q��(b
�|�9�r�Bޘ7.��)*����ʎ��<»9"jw��|D5gv;}vfP*�5�+�w���UNIR� !p�2��}��%b�B=��=b�y�~`f��%<�����j�	�+��y*1m��`ާ�e����08��J��wҹ��ar�Q���H [)����řn�P��4�A:q��ꗱo�F3�����v@�T�F�P�*$N�ta=Z�����H�ZW���?*`�WnQH��-~y��0������oy�#����Uq�ό��?wU����Y�H}9c�w��:b�1�1��9�hOΑ��`׃&���3�b�\S�MKG>ia�Y��/�Z�i��b��Su�3ڙg}��Q�1�8rۅ`��}�/�Y�0��fs����F����*1�Y�ECus��'P�p����x)^"�3���tL�!���pq�BG2�TRo���o�D�ܣ��º:�C��1S}��Genf-��'4vFMr57ש 6m��qʦ��j"��2{�	o�6Ī�TwM�5�ֱ��Ĕ\oYi�4��h�;qc��-����9 �}�޾n����''��ԎkW�����7� ze:5��!��
��6(��!����?���#��j?w�_�pg]��Kc|Y�����p���}��˳6��}�]��v��dєc_�Ai��zT&Y�U��!3K�&������D�[̧�Hݛ��5��^�qU�gz��ԌV�j��*=v�fNk�����\b��J���*�N1�hV�]�V:�k�㜡@g=��rۛ���E��}Ka�t��m�����z����A:�:��-��K-^W���k�5�2���BqY�P�����Z�O�۹o$���jA}���hT?�Su��c���=�?K����8����0G-197��z3x4�4f�H��Q��dbNW�M�������M :-;,��r�ӧg鷷���zf�8�;�@}� H-zZ�m����p[R`�Y�%8:�]�?;w�5�����͔�����+�c*��V�� �m�o'�G���SncC��B�N�B`��
��D����?��Έ��l��͡��F�ei�m��p�M���)��h�X~��n�.�f��v�_`
c��]�(3��C�@�n�f��F}4��u�}?���n��r$*I�Q)�Ɛ���P:DV���
���h1�2@�ׇ�3�ߴ�t�U���O��|;�q�O�h���v�6�ˈn��-�`�
6( ��� M�o�{��{']b}j��X�7�����L���^��T�?���ԓ�gʻ�6ײL:AG�.i|y`�m	։���)g0�d����;��W�Q�V�E���!���J����������P�ZUsX!Z�o��L����QCh �[����.A0��f-k	�Xh��Z�����ⓡ�.�(Y���&<I��[��_c���p���SU<�(+Z?G�j,!r���$#�$��;���hO�ݵs��l�!��l����v�.$��v�}���<!o9b"��yC��8����J��B�"�/k�l�� K����`QǖT�)�cV�\y�;#�5���p4�2'\k;;��s��T���W� Z���=�O������yJ�3\��9R�թ9�>���mύzN;�
�����XJl�wGF��p�J���ɑ��Cz�+�����K�&_xܻ�P;\�l�˳����z��gػA�D�g�����:�U��"l�e�O���E �����V�����9`~���S�U�K�~���Q�rD]֯V�K�Q�J�2�Q>̪�,��j��R�I�̄Jn>���bp���G3"��z���G_�NW��oKq�K��.y�R�(�?P�y��/�`΋#j1w��i��|�ܘ���x�����oL!oa��S������E=l���NAc�tW�QE���7��ᏡAY8��O�}�k�R�bu��6���E���>�TS_�
:�]�M�~R�"�Ff6�C�yZv0��rd�6ܖ�⎣}&��Dϒ5�1��V"r� ��Q��,��/��a/^��*��j�=��F|��kM�;?M�*C{U���w�3�\G}�/d��I�o.��L����q���?d��S$L��)~�t҃�\q�2J�����x1�(X��:]�)�=!Y%�1�N#|�*K�<�O檴��X�sM�u��E�����2"�q�iȵH<wșx���U�M�~�`�j�$}�;��c͔w]�D��le�M��ƛ͛G�z�����^�����>xUj̑���5#T  /MC�{r�m��V�T���R��b��@�e��0Mnΐ�`Dp��]���-'6�g��S��g͛.� �ï�_o�%�>���	O��NUv�-�p�p�K��摋�	�SR�J�������_��S�͐�s�l�{�Ls���֠�(�1�?䰹F��Q�+e��t�d">>3wbv�
tN4���[�S�6oH�gz����&4���{ &��H����g	���e�uT�ڌ1"�p��+�KA�Pw�!c����l��`�y�X�F�S@ڪ4�	�bhxR�)E��tjxȘ[�H~�;,�gX���&Zc����`�,mC��c)	�l	-t��P;a�WH������v�_f������d�^��K�lz/S��{��Ɂ��kȼ>�m��&�Y9X�:"���!�t2*.-+��ɔ/EV����U�ֵe�Z❎��wN5'Bn	#�(�Cp~���%�W��Q! ��qjn��s�}�G�K��{u��`;�Td���T���C9���:Me��Yj�_�h�k�ꮔ%�;E����-(XQ�t\�u��1�\h�M#+|c���I���ɞ�Զ���ib�Qn��z�	ޮ���j����Rҧ��y�@��??ئ��6@_�*e.?�@����i�a
�ء���vB"�Z�1]1�����$
Ab�Ի��u�Zi��u��`#�,���s���?�3A��`;U����z05��Z<0ز|��M��w��2��'��j��u��"�|@���xEP���(���sbJ�q��89�ۛ{���;�6"�3P@����nT�A!���|"~��4Ե���*u�?[_� ���v��ѵC�S�݋
"�$Q�kZ�b�J��f7'\58�(X���=����YJ��C��i�⽩7�=!}���п����߯O@�X �ͧ3Ca�����6Vö@E����]H���7+�Ly��[�Ӭr�?X-ﳞ*�gx���