��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħP	�(<�%5,i v1`��Z��7#��kϟ�,����I�v�u�du�|
�����ZjGjX[�Sr��:�vH�~x`v������#�v�0r�g_5���Gn)����h�����ed���F�/^qh���G�>���= �7����wmLxĐ�jH�n[n������M���	�JF�fL��`�)Z=hZL�E���������^Q�e?
r���ʽ{�X�G�'�i���^(�C=i��� �L��uf4��*�j�����̷������:��M�z�_@�&[aMɄ; M�a�usvg�����I��o�?�$�S�*#�/�0}f
�׀&�J,uu��|�wu��0��!��m�,�
e��=ۖU�LZ_b���Yg���I+b'k���?7g�q�bD@�wР����]C'ym/#���f��Q�7����u�]�O�t`�=@��Tu�&�d��H��TM[�{̚I�;��7׍>L�Zv�zyÜn��H�k̘�v��x��q
p���⠿�-/��lH��Y�e̊�$\���LR"IT�kw��@�b!�1!�"Wt�*�I͈��'�FuBz��H(�d3m�O�����G?w1Y�"�q��Q�_����1�(~/<V�~�ɩ5��/U�c#C���X�:E����ҚK�X����~�#zz����x��Pԣ��B�6T$��%@���2����hgY��)�gP�+� ȳWq���Es��0M)5j�;���h��e�_�M�ʢ�ن��� �b\�~l�^���x�U�Jc«[�}����T4�Yx�M���F�"fp��R� .�n}Z�}�K�X���15��JyU)�T��6K���J�v��¼�i��jJ�b���k�K$�ܮ�"d*����y(O�V��3���b�1�2Z�я8��L#S��/.iDM^�����Ȥ!�rhr�(��Gz��R �(������0`f��Ns	֠�ӍX^st1ԭZ�9:����Y��G��_6��=���I������^�;����R@�Զ��)R*1�bѮ���h�j퓿=�v��P�s"}�d�׏f��%Ů�
��Y
���2\�+�����ӻ
̓"q�guЄ�9�H:����-!R�R�����4d���8[�Ѕ�)D�s�K�$Xk�XB8Z��R�I,��Z�+�i�Ҁj�$�eQ�Dt��Jw6���:E<Lo������nq�X�D1ĭق�>�q�,3E)����O�Ԭ:��~N=�\�smÎm�:qmR��O��B��j�Z��`���Tdv)M��{K��r��rc߰�0�*�QJ�n+�+_��ki�7��ە����M�Vo|h��7X� 1����F4��č{@����_%'��^�J��5�c�x%7�,UO��2����.�KʄN��ޡ�@ m���F�����=¾���?l�0��Q�mB��2T��}�A�u5�0�R�&}&T����yQ| ~h��0}����K�)��F��(x[��"�<I�-o9aI��e�-t
�/���!�+����@��^�!��Y݈?�"rz,,m�YS��W/#��\����X<��e�:���Ccc���.�Ub5���D�*ux����0�uH�ؚ��.9�'U�#��!��n©���]H��/ZL�@��|Ƿ