��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�>��,�t�Jq�%�qr��A���/4�HRN��Ί��w:p��'�˷34��>,'2��q�B�'�ri�v��B>�k����2(Ahb�I��Z
9�-��I|:$�a�^�^RB������������i3���k�����Ԓ��B1��X�}�%Z����'z�_�x64mhOm~(�� '��U�B3��H��.�6��K]v�(��`ჸ�<D������Ö \��j.o�ShL�v5��SԲ��z�өY߫�%��?�'�����"��@�_���B��
�k�7�S�b#5�	�9��K��b�3��j�BM0� ��@��b"u*C���o�˸�V��v�$���,ް6b�?Ph��lL��5�V��am�!7��!A{؂�ߢ3�"=4�Ct��B�b՜H�+O�X s�ڼ�R�O�Ū��������2�p��>�N�9�>���m �Y&LE"�i̓Z�V���6�! ���Qf���?b}R�V��p.kN��rzX�H�}��>�<7U4���� �`*g/�z�b/܄��O������i��*�������"����8�[6��XC
�	��_�HP�Ҩ�J�)o��s�4O���q�\NLY�ӵ@�,�g�hR��@���GN����� �+8�[� |
�(�GR��rJ����x�t��,4�¦���<��%�_];�E�����`���d����":���v�nñF)-*{ќ5q�/��G �Fҟ���ټϞ��
�UeY����YN����0�L�h����!�YQ��݊�����
���u�����Vl����x�҈C���gێ!�����m���y�]�!IL��n�k��B�˓��4��d�PDT�žDi�������^�E��??w�ʀ�;�4�+�e�J�Vy�Rf�T2֝���%��2j�����)�IP�zss�K��e�>�ؖԁSߔ�%��>M�Q��a�()#���Ly>s�������c�a��^���2�
������w�������,�v�ξB㗀4s��5|Q�1	�C�f3�]��zR�s�7�` �4۩nm~��*��{�kFF߉о�4��;�HT⋳;�4i�,�ݚ�P��LΛ0�g��%�{a�aJ��,aX2� �㩜+��ǡ�*4vI|;��9j�*L��|]!�g�y3��箳�C,�s�Y��o���	��[�0U� 09'���^�'�� Y�'XY
���&5�ͺ�^�*4��d�a���� .I^�
����@����_����Q���E��v.ٽp�G�WZT��b<,~�wq�>��"���I��(-K�g������z�;Mɠ�'8J"�H���������h�N'C<��ᒎ��jƫ���ԕ�I�c�K�p|�dR��!Ĵ�K��[Q�c4W��!d��A���)��k?]T��h~�ԭ-w�f�Bp��+��~'g�t�_B�;J}3O{g���L�9V����4�қQ�v�QOg�(֯�\mL ��g�~�v�)�����Y�Kp�[ͫP�.ov�yw�s��Ǥ��^�K���\ؠ�E=�r/8�,G�eKa�t�����h����j�:W�Q	G��y�E�i�����a-6��4�+�s�i��K��\6~���B�hV�3�67.�������iA�����t��R�ВӠ�q��r>6K���ם���!�/.���#W/��c7$<f+<��g��N��n�Z��qZ����Dߒp��TinL�_�䉍��0u���*L]5K b��e�f�32`Y��8D���o����ie&���b����!��swќ�0��*�����L���?~5
@.�io���U��c���O�լByK5@��cK����C�`���}�C��]�b�j�pZ�mm��f)�RoP»���=�1A�+�Q�� &1�7��v��hY��?����v��;x���"����纱�hB��1g����
�bĐ��B���3K���vޜ���P#R�.R�[�9A��
��� � Cv������+5��alB>X�B����]�ȷ�x} �P� ��6� X�q7]�-�4��4U��ˁd�.�u�DR��C�)L��y�t��W'�������$-�s���_) �2@u��ҝ �x���m�9њ�{4��b�H�p�K�v����t�������2m�.�/d��j�ҍ��9u�!-�dB��܂�y:
���YT9�#؉�s�r�4o��촌�?���h���mg���!�~������x0�:9Fs-` fs�nKp�bow����u�q�VK}�rN�F,�Ƭ�zG<m���@3�G?w� #y�K$��B��XK��Aq#�P�*5��+H[x��Q��D�r^2
�k\�C��8�����4|���#̔�{�٥�#�_�|�b_P���e�1�;����:�rr8t cZG?[:�C�k�^>�8 >��I���v�JX^�/!K����݊Lu^<�� S԰!�[�a~� ���nfe�2l�Mƾ J,k)H��M6j�_���>A�/�G	�6�zLc��R��a�Dd���2yߵ4$�K��)��.�䞂����YXfrAs���e�-M�u�`�E�n����C�ot%"|��غ�,�E���OG��>|I�~�8=d�%N�M���*�g�i����=U�����*�ޅ�fY��+5}\����Pu�s��A2Y���n �������
��Ϋz��Ħ�p�ρhnq�VE`�66�xj�P�ݸ�Y��ɍ�y�ڋ�L&�`,br���ކ��uW��m��5l����Sڶ�B2X�R_�Ɵm�n⼗c��� ���N��ZT��2@A��4�_����#���z������# 4P!�u*|�)�7D��c����fT4��w*T ͷ$�ʫF��DT�YG0���,��In._��f�y�i���^���]���[-���+g�N5�]*�1�i{�$�&���j2��k�j<���Srw
���/[��y�T�wͥ �;\|��ؓCY�!��y���?�=-��\TS��D�DO�F��ZG��Ox�.*%��w�������'6V�'s�O1��ް#,�DAW��>�V��[��F"e
��W��sy�k��Z0 e �h��$`�m����;W����{�]<�Zf�k����G��p[]c��d7c�V�����5漦h���=�*���v�1)^�5�oK����iG�\��n����'�ON� @� *��	��a������Ȣ"�=fN�X�)���I��_�8���e�ed��48�E���Lr��n��#�p��N�;g}�L�d˻��Ck�A��@���K�wBt�R���[���s'��I�X�X�x�.]Q��sg�<�K/� }X&�y��a�wW���=���-<�]�O{�ɍ�����rP&�\�)�z�7�E@/��Lb�#��Ϩe�8���(;1�f�c����q4u�j]g�5�)����[Q@9�f�ZA�sJ�7�ul���ۆ�4~\<���b�w��ܐ�¡~H��Ѹ<�M���JsTJİ}�����I�Zۘ��ێ;|	� SS�u~�������>�1Bw�,��r�'�7Q�G� ��awU.��r�~���	�m��gl�`���X� Tv��F�{��z���e��v>? �����yh
d`��h�\�R����;X;�5n��:�{��]��Ch��oV��=k��\%l�]z���V���� gI�Y-���mk���0����%#%�����X�Vj�t������HT�qd���u���H ��v'������_M�9q|�0!ޡi�h!fZ#Aop�Q�������P֞����9')�I��c�-6��<X��odZ��Fp��Qj�{*�k��Š{a�!΃.^`�b�c��5'(1�=�x �>:i�$�Ҽ>RK1�����!^�S͌���>�r�#�=Z-�P7��y��`�f� �kG����Ǒ4�� �;�-�#��i+��3��H����?���z}g���KН���懘�U2����H�jU�'s,�s�B�mD-��r��߱�X��~�j��E�欵bN����MiS7�*��8��LFaY�����z*�v5�V�@iV,�vǽr����l��v������y׏`�
ͻ� �OK��I/�>V�f'��}R��;z
K�h]hO��uM��iU�K#���h���Am?f��9���J��r�C|\����	JU��Ho�ĭ�3d��y5rZTh�T��<_�w�j~��{�=�Y���N.It�1�Y�ء�����ZK����R­\?�R�ݓ �J�T���N��ٷd����ZIW��tA	�Fu�0��/��]`�����>��홴Û&v@�Ԛ�I� � �@�� ��*�;0�p���c��3��~ȬR��5C���7��'S��NVqc�#�+��pFD�B�!���WrP��T�
��^>��7)U~m�|�A@	Tgy�C+H�y^b<,R��ˆ3���AG��F�H�M��a������|r�Hd��o��T�.�f+Ѳ�8P�5Ct'S�斤8Y�&,�­9*�x�{X�5�	G�~��}Z��5���m���=4nX����������C��k�۟=ĕ(���F�E�������A�RF��d�@�~i>�.���xS�Ub5�Oog�Kp���Һ_�ɇ��>�g���x�B�"4W&���E����m��K#Ea�'�(��8} ���<���za����@����Ӈ��+�$����-���B��r��>��u�a�u�Y��
��i���)���ԈZ8~)���l5`煣ղ��[�H�-���rq>uf�d�8�S�%��qN��I[�q��٢z��c<� ����<�)w��)4�8�@]ԓ^��� ��7�^�_QPw֎���mF�:!J���`Q�p���)o(۩���~C�����V{X鿝*e�]��/�ҖM,������[������i�<�y^�D��`��&}Թ毱�����\��&��6�MrB�1eZd�~i�Ⱥ�9�����FS�ɍ	�i��ȼ� �M=}��<V������Ju�L����w�woB���Z�2?o!��&��M_)Ô�>+Y߂5�u�� J2=D�d'uim��1����rI�4m�-�S��L��	��
�*|EW��<�~�P�O��8�I���G�>��"��
i�a{T�$�	9���\�� ��cR�%/CEux������WZ������� 'i�o\�U�ә��9�1;��E��kۅ4ac��a!@D��p�l��`�ud�u(q =<�'[w\�Ԯ���fm_=%��Zf���~�0�÷�}�#)��g�k�I�K�f����&<��T���V��_,"�ޫl�]$|2��ױ#ʹ�y�j_������a �&ٻ���m5���<@����v�[G�l_w} ��''�׸��|ס��߄	�($�u/�Kݻs+c]�T~Ie{b�B%�$�(-:T=~�Vd��ۏ���VM�3'��K�R*`^<�WY ����A`�=�����7�:�U�T�U0��q� ���J����	� j��6�=��8xI!�f�9ܯ�Ll���7~ĺZ<�Cd/��L)H��-�f���= 9�4��L��;'-�ό��B{�	{���t@PČD�.SK5]�Kgb���S��@���Q�M,3N"�Õ,�X	]����5�%l�\-�m|�{j�|�>全�u�F��<x9�o*~�!�8�l����l�����%
�|��{��5-j�r�	����ߏȌ#�C@���b䰏��I�K�
l��_��Fa9��R�	jC����� �	�؂��7�^�{�lۮ����91>l�;"M 0��NN�J���G���M&�83b_����j{f����E�S �^K�A����6LPLW1�]mN��"���B5q&�&�*Ɗ��@G?���)�o�Uc>�,��Jy����%o�M����j��1�-���/�BY���~� ��"*��&zX1BB'!������\"� YE'I~(ft�Vu�c�gA|�b�U�����:�v."��c\�bK�ү�I���i�wM�99'�&`�(�蕐�%`��-kbbS�b��kv�ua�]�
Q1����`�`o�j�9XD֬��\��~]J�
�e�0��)��UfߟT��h��1���p�C��؍��=�6Q=m����\1�X���������Z��kF������+}^�-�z|�c�2y~�����/WB	�[����=�u�����"����^�M�P��Gq/`d��oZ&X	�8��$�$���xˠq��������d[��U�ƫBn9�t�i @�����^))��Q��{�J�jgh)Tޅ�z�����mT79%���GF:�c)�ܬȑ��0^ve���~k��2�-X�C	��ߝS
U{u�� %g��pE�dz��Ғn��v��J��OO��~�����@|e�����~�վ\.=����r��);z�Z�#!OV�='D�/����>�̈������]u��H�K2�I�\��CE�'�6���z��Ն�j�\6�G�H̒F�M���'El���>��1�^���6J�?�����C0qh�-;fG���ڽ�B�bhy��i6�X�6hv�ݕ F �ԁ?;L�b�$%��f��`[;I���Ѕ!�:Y����!���И�Z���A`r��>?ʪ��.�0��ݞpw؀M\OQ��a���C��xL_\Eu�/�pgݙC���a���;uG�0.X�3z~�-���E�| �WpW�S���O
��A۽���3�С�4n��R�wm�?b�,� 
I�+W�D]�䚣���ͦ�!��[4V��	���γ�x�.b��J�	~�<�ԋ���6��~�֬�J�'ˤ�{�e�>��.'�Z����W[E;����$�Ty�M����Kvݣ�j�u4�Ҳ������k	9U�w��׺+W�����*|;<�FQ�df��B>�c��"P�j�Co&\�V^�9瞚/����*��/�R���T߳�)���$��2�PFݘq�|"nWؖ�k�t-o'���f�ƶ�Jـ����;�ͼdeU3o(P��*_��������A�s�u�sxGl���M�K��oUc��O����� ��(>?���R`f��s����]�2��X�ma���D7Ð�j�@AsO��59�����Xvi��"�ϳ9�)޵t���&{ͧ`n�B0�yQL�m��PR��ے^ �ۧt� D�������K��Dܤ��^R�XN�A.�B�#�?Du�C���Sr�qm�bѸڤ?k߶��w����{@Q`��~b�0'vb�ľ�S�\)�Ƞ��4�!Nb]�l�0j����8O�Y̉����,��l$Q�91B~ q���ά��AqZ�h萑~�si��*��}�z��+��<��i࢏u��������R�׆��Au1'���'�r`��3 �J��&�4�p����8�.���#���B?���Qu]q�bMq8cƕF��n`��@p�J<.nFR�ݶ�y�Ⱥb����i�τ6Tt�$���怢����E�ӻ��)�L%�-WVy��<��x��%njc��k��a�ؼ	�(��O^ �� Y�Z���oE���+�sL�>�u����uȧKPX�ڪ3W!���0�5d$[,���Y¬�ڝ�(0�}]Yϵ��'�x��q�v��-�""�Xs�.X��h�b�5�CK~HǑ�{(����^��꒘D]_�?�h�m9Ž��� ��͠B�ԢqO��N�J����B
�EG�Z�/��&�0��@q�	����מ�~��H�[�gR���l	��փz_�� �j9��)Q���Ґ0L����e6���BEeI �K��&�9��%�#���u�^íܞ��Ā��
�������쳉0�9J��5��(��r�՜�m<�|�Eo0c~>�i��y0��(��7��}Mp���
L˺ޓV��l���=��W�������R@?UU����ȏ�C�
�vkL{�B �J�%g�?"�����8���rca�{�ً��:F�K������0���^Z"8�����h��yPq��.qD�CIt�hm~Ůq5�fKeǰ1�����<4�Ö�b�T�=>ڶ��f��X8Ѣ�ԓ��"�m��r}����F�,���lR��lhc��0�GZ̋�Y|����.�pY�������i��U!�0=����5�7X,e�zğ�f�[��l�
BQk�Ʉ%U�,"��ߪ�駯�F�V��w��4�� 0f�'7g��%��&���~*�ck����ВΤ��ioN4��;��κD��^
wB��,h�S������!#��.^j��L�TdsT) &"z
��=e�M�^�[N�_�����Ž̍5}�����>�W��R��]��ɩ����>�0�S�FP��A�΃+M�}���М+�O��㜘�ɷ��q�d<R��Z�?�0��Ĉ��f:N�B�SÓس�~
�- ���5z�ȝ�^��ΐ����J��N���b�;#���"?pk����Wd�s4<�a�� /�z����vD�:�u�,,�kӉj����Wy��Dâ�"��g�N~�Q��~̉�4E�-I̪J�˪S*�����"�A��~:���s��MV]R������`��'��YͮP䤮�3��V�\�?�����Vp	�6�z�ḠFI]��h#�PU��2����y�I�d���o�;D55��#`z}��� . ��s�t��c�8WlW@C��$%�m��q>����+�ɴ9�}���C�ÿ>F�LN���O8�(g�-��Οم�2O�)B�?�{��T���2�����Nɭste�^����g�e�br{,
}�}�΄�'�z��&���d�#�@4/���-�ccA��=���K��^Էax���@�v���ű�j���E}u:'��0؋�2��C�\0D�"�La!�2��E��,��r�Z'�Q�&љ�g��ɿ��B|��&����p-R���m��'d�{92ܢ`��MX
а��p���o%{�'�2 ͓ݫ#��;wN&�->nǅ�'�����[x��%x�F��ZY���.�#��U&�~e����v
 x�̢�{&�N�y��H��;��p�˼��e�j���׾$2�$k����Hy6Hu�� {���
�!#fa�z���fQQ�v�6Y��;f)��:��$���F,�����X������66����.��^򔌩�nZ��,����Z��؞-�ISo^H�����[���6���2�AI��s��v�'�c��\U�͋,F��&��,�����m��k��"�|[��؛	��$A�*��%Cz�\o�Pl����RO���U�0�dda�O�{z� �r�`��K;���ǯՀI��<wS95p��&H��ˇ[���]���,<q�Ʀ�5��DYN���=�����H�3d����68